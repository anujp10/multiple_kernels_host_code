// Benchmark "kernel_10_0" written by ABC on Sun Jul 19 10:21:02 2020

module kernel_10_0 ( 
    i_10_0_31_0, i_10_0_180_0, i_10_0_185_0, i_10_0_216_0, i_10_0_277_0,
    i_10_0_278_0, i_10_0_286_0, i_10_0_324_0, i_10_0_408_0, i_10_0_424_0,
    i_10_0_427_0, i_10_0_432_0, i_10_0_433_0, i_10_0_444_0, i_10_0_465_0,
    i_10_0_514_0, i_10_0_697_0, i_10_0_954_0, i_10_0_955_0, i_10_0_956_0,
    i_10_0_957_0, i_10_0_970_0, i_10_0_994_0, i_10_0_1116_0, i_10_0_1119_0,
    i_10_0_1167_0, i_10_0_1239_0, i_10_0_1243_0, i_10_0_1244_0,
    i_10_0_1307_0, i_10_0_1540_0, i_10_0_1541_0, i_10_0_1547_0,
    i_10_0_1549_0, i_10_0_1550_0, i_10_0_1690_0, i_10_0_1758_0,
    i_10_0_1760_0, i_10_0_1818_0, i_10_0_1909_0, i_10_0_1911_0,
    i_10_0_1984_0, i_10_0_2023_0, i_10_0_2029_0, i_10_0_2434_0,
    i_10_0_2442_0, i_10_0_2443_0, i_10_0_2455_0, i_10_0_2456_0,
    i_10_0_2534_0, i_10_0_2659_0, i_10_0_2719_0, i_10_0_2821_0,
    i_10_0_2830_0, i_10_0_2880_0, i_10_0_2881_0, i_10_0_2883_0,
    i_10_0_2886_0, i_10_0_2887_0, i_10_0_2919_0, i_10_0_2920_0,
    i_10_0_3034_0, i_10_0_3075_0, i_10_0_3198_0, i_10_0_3384_0,
    i_10_0_3385_0, i_10_0_3386_0, i_10_0_3387_0, i_10_0_3388_0,
    i_10_0_3389_0, i_10_0_3437_0, i_10_0_3537_0, i_10_0_3540_0,
    i_10_0_3647_0, i_10_0_3650_0, i_10_0_3652_0, i_10_0_3685_0,
    i_10_0_3686_0, i_10_0_3720_0, i_10_0_3783_0, i_10_0_3784_0,
    i_10_0_3785_0, i_10_0_3787_0, i_10_0_3811_0, i_10_0_3812_0,
    i_10_0_3842_0, i_10_0_3847_0, i_10_0_3848_0, i_10_0_3908_0,
    i_10_0_3963_0, i_10_0_3982_0, i_10_0_3994_0, i_10_0_3995_0,
    i_10_0_4115_0, i_10_0_4172_0, i_10_0_4215_0, i_10_0_4216_0,
    i_10_0_4218_0, i_10_0_4283_0, i_10_0_4530_0,
    o_10_0_0_0  );
  input  i_10_0_31_0, i_10_0_180_0, i_10_0_185_0, i_10_0_216_0,
    i_10_0_277_0, i_10_0_278_0, i_10_0_286_0, i_10_0_324_0, i_10_0_408_0,
    i_10_0_424_0, i_10_0_427_0, i_10_0_432_0, i_10_0_433_0, i_10_0_444_0,
    i_10_0_465_0, i_10_0_514_0, i_10_0_697_0, i_10_0_954_0, i_10_0_955_0,
    i_10_0_956_0, i_10_0_957_0, i_10_0_970_0, i_10_0_994_0, i_10_0_1116_0,
    i_10_0_1119_0, i_10_0_1167_0, i_10_0_1239_0, i_10_0_1243_0,
    i_10_0_1244_0, i_10_0_1307_0, i_10_0_1540_0, i_10_0_1541_0,
    i_10_0_1547_0, i_10_0_1549_0, i_10_0_1550_0, i_10_0_1690_0,
    i_10_0_1758_0, i_10_0_1760_0, i_10_0_1818_0, i_10_0_1909_0,
    i_10_0_1911_0, i_10_0_1984_0, i_10_0_2023_0, i_10_0_2029_0,
    i_10_0_2434_0, i_10_0_2442_0, i_10_0_2443_0, i_10_0_2455_0,
    i_10_0_2456_0, i_10_0_2534_0, i_10_0_2659_0, i_10_0_2719_0,
    i_10_0_2821_0, i_10_0_2830_0, i_10_0_2880_0, i_10_0_2881_0,
    i_10_0_2883_0, i_10_0_2886_0, i_10_0_2887_0, i_10_0_2919_0,
    i_10_0_2920_0, i_10_0_3034_0, i_10_0_3075_0, i_10_0_3198_0,
    i_10_0_3384_0, i_10_0_3385_0, i_10_0_3386_0, i_10_0_3387_0,
    i_10_0_3388_0, i_10_0_3389_0, i_10_0_3437_0, i_10_0_3537_0,
    i_10_0_3540_0, i_10_0_3647_0, i_10_0_3650_0, i_10_0_3652_0,
    i_10_0_3685_0, i_10_0_3686_0, i_10_0_3720_0, i_10_0_3783_0,
    i_10_0_3784_0, i_10_0_3785_0, i_10_0_3787_0, i_10_0_3811_0,
    i_10_0_3812_0, i_10_0_3842_0, i_10_0_3847_0, i_10_0_3848_0,
    i_10_0_3908_0, i_10_0_3963_0, i_10_0_3982_0, i_10_0_3994_0,
    i_10_0_3995_0, i_10_0_4115_0, i_10_0_4172_0, i_10_0_4215_0,
    i_10_0_4216_0, i_10_0_4218_0, i_10_0_4283_0, i_10_0_4530_0;
  output o_10_0_0_0;
  assign o_10_0_0_0 = 0;
endmodule



// Benchmark "kernel_10_1" written by ABC on Sun Jul 19 10:21:03 2020

module kernel_10_1 ( 
    i_10_1_53_0, i_10_1_86_0, i_10_1_118_0, i_10_1_280_0, i_10_1_424_0,
    i_10_1_427_0, i_10_1_436_0, i_10_1_437_0, i_10_1_442_0, i_10_1_444_0,
    i_10_1_459_0, i_10_1_463_0, i_10_1_467_0, i_10_1_514_0, i_10_1_518_0,
    i_10_1_587_0, i_10_1_706_0, i_10_1_746_0, i_10_1_764_0, i_10_1_793_0,
    i_10_1_794_0, i_10_1_832_0, i_10_1_833_0, i_10_1_964_0, i_10_1_989_0,
    i_10_1_991_0, i_10_1_1054_0, i_10_1_1055_0, i_10_1_1361_0,
    i_10_1_1466_0, i_10_1_1541_0, i_10_1_1619_0, i_10_1_1684_0,
    i_10_1_1685_0, i_10_1_1768_0, i_10_1_1819_0, i_10_1_1821_0,
    i_10_1_1862_0, i_10_1_2182_0, i_10_1_2306_0, i_10_1_2330_0,
    i_10_1_2333_0, i_10_1_2336_0, i_10_1_2357_0, i_10_1_2360_0,
    i_10_1_2449_0, i_10_1_2453_0, i_10_1_2468_0, i_10_1_2478_0,
    i_10_1_2482_0, i_10_1_2515_0, i_10_1_2528_0, i_10_1_2539_0,
    i_10_1_2628_0, i_10_1_2630_0, i_10_1_2676_0, i_10_1_2681_0,
    i_10_1_2717_0, i_10_1_2728_0, i_10_1_2827_0, i_10_1_2828_0,
    i_10_1_2830_0, i_10_1_2873_0, i_10_1_2917_0, i_10_1_2918_0,
    i_10_1_2920_0, i_10_1_2921_0, i_10_1_3195_0, i_10_1_3197_0,
    i_10_1_3206_0, i_10_1_3208_0, i_10_1_3209_0, i_10_1_3353_0,
    i_10_1_3384_0, i_10_1_3403_0, i_10_1_3404_0, i_10_1_3434_0,
    i_10_1_3451_0, i_10_1_3583_0, i_10_1_3584_0, i_10_1_3587_0,
    i_10_1_3589_0, i_10_1_3610_0, i_10_1_3614_0, i_10_1_3620_0,
    i_10_1_3688_0, i_10_1_3734_0, i_10_1_3835_0, i_10_1_3836_0,
    i_10_1_3857_0, i_10_1_3920_0, i_10_1_3988_0, i_10_1_4031_0,
    i_10_1_4144_0, i_10_1_4147_0, i_10_1_4171_0, i_10_1_4192_0,
    i_10_1_4279_0, i_10_1_4577_0, i_10_1_4586_0,
    o_10_1_0_0  );
  input  i_10_1_53_0, i_10_1_86_0, i_10_1_118_0, i_10_1_280_0,
    i_10_1_424_0, i_10_1_427_0, i_10_1_436_0, i_10_1_437_0, i_10_1_442_0,
    i_10_1_444_0, i_10_1_459_0, i_10_1_463_0, i_10_1_467_0, i_10_1_514_0,
    i_10_1_518_0, i_10_1_587_0, i_10_1_706_0, i_10_1_746_0, i_10_1_764_0,
    i_10_1_793_0, i_10_1_794_0, i_10_1_832_0, i_10_1_833_0, i_10_1_964_0,
    i_10_1_989_0, i_10_1_991_0, i_10_1_1054_0, i_10_1_1055_0,
    i_10_1_1361_0, i_10_1_1466_0, i_10_1_1541_0, i_10_1_1619_0,
    i_10_1_1684_0, i_10_1_1685_0, i_10_1_1768_0, i_10_1_1819_0,
    i_10_1_1821_0, i_10_1_1862_0, i_10_1_2182_0, i_10_1_2306_0,
    i_10_1_2330_0, i_10_1_2333_0, i_10_1_2336_0, i_10_1_2357_0,
    i_10_1_2360_0, i_10_1_2449_0, i_10_1_2453_0, i_10_1_2468_0,
    i_10_1_2478_0, i_10_1_2482_0, i_10_1_2515_0, i_10_1_2528_0,
    i_10_1_2539_0, i_10_1_2628_0, i_10_1_2630_0, i_10_1_2676_0,
    i_10_1_2681_0, i_10_1_2717_0, i_10_1_2728_0, i_10_1_2827_0,
    i_10_1_2828_0, i_10_1_2830_0, i_10_1_2873_0, i_10_1_2917_0,
    i_10_1_2918_0, i_10_1_2920_0, i_10_1_2921_0, i_10_1_3195_0,
    i_10_1_3197_0, i_10_1_3206_0, i_10_1_3208_0, i_10_1_3209_0,
    i_10_1_3353_0, i_10_1_3384_0, i_10_1_3403_0, i_10_1_3404_0,
    i_10_1_3434_0, i_10_1_3451_0, i_10_1_3583_0, i_10_1_3584_0,
    i_10_1_3587_0, i_10_1_3589_0, i_10_1_3610_0, i_10_1_3614_0,
    i_10_1_3620_0, i_10_1_3688_0, i_10_1_3734_0, i_10_1_3835_0,
    i_10_1_3836_0, i_10_1_3857_0, i_10_1_3920_0, i_10_1_3988_0,
    i_10_1_4031_0, i_10_1_4144_0, i_10_1_4147_0, i_10_1_4171_0,
    i_10_1_4192_0, i_10_1_4279_0, i_10_1_4577_0, i_10_1_4586_0;
  output o_10_1_0_0;
  assign o_10_1_0_0 = 0;
endmodule



// Benchmark "kernel_10_2" written by ABC on Sun Jul 19 10:21:05 2020

module kernel_10_2 ( 
    i_10_2_171_0, i_10_2_174_0, i_10_2_175_0, i_10_2_176_0, i_10_2_216_0,
    i_10_2_217_0, i_10_2_316_0, i_10_2_317_0, i_10_2_318_0, i_10_2_321_0,
    i_10_2_322_0, i_10_2_412_0, i_10_2_429_0, i_10_2_442_0, i_10_2_467_0,
    i_10_2_797_0, i_10_2_800_0, i_10_2_892_0, i_10_2_958_0, i_10_2_959_0,
    i_10_2_1006_0, i_10_2_1026_0, i_10_2_1027_0, i_10_2_1029_0,
    i_10_2_1134_0, i_10_2_1233_0, i_10_2_1234_0, i_10_2_1235_0,
    i_10_2_1236_0, i_10_2_1237_0, i_10_2_1238_0, i_10_2_1242_0,
    i_10_2_1245_0, i_10_2_1306_0, i_10_2_1307_0, i_10_2_1579_0,
    i_10_2_1580_0, i_10_2_1651_0, i_10_2_1652_0, i_10_2_1685_0,
    i_10_2_1819_0, i_10_2_1820_0, i_10_2_1821_0, i_10_2_1951_0,
    i_10_2_1991_0, i_10_2_2184_0, i_10_2_2185_0, i_10_2_2311_0,
    i_10_2_2352_0, i_10_2_2359_0, i_10_2_2361_0, i_10_2_2364_0,
    i_10_2_2376_0, i_10_2_2410_0, i_10_2_2448_0, i_10_2_2450_0,
    i_10_2_2457_0, i_10_2_2458_0, i_10_2_2461_0, i_10_2_2462_0,
    i_10_2_2629_0, i_10_2_2631_0, i_10_2_2635_0, i_10_2_2662_0,
    i_10_2_2719_0, i_10_2_2819_0, i_10_2_2827_0, i_10_2_2829_0,
    i_10_2_2830_0, i_10_2_2918_0, i_10_2_2920_0, i_10_2_3093_0,
    i_10_2_3094_0, i_10_2_3151_0, i_10_2_3276_0, i_10_2_3388_0,
    i_10_2_3391_0, i_10_2_3402_0, i_10_2_3404_0, i_10_2_3551_0,
    i_10_2_3586_0, i_10_2_3609_0, i_10_2_3616_0, i_10_2_3647_0,
    i_10_2_3783_0, i_10_2_3784_0, i_10_2_3787_0, i_10_2_3836_0,
    i_10_2_3838_0, i_10_2_3847_0, i_10_2_3853_0, i_10_2_3855_0,
    i_10_2_3856_0, i_10_2_4127_0, i_10_2_4212_0, i_10_2_4269_0,
    i_10_2_4285_0, i_10_2_4564_0, i_10_2_4566_0, i_10_2_4567_0,
    o_10_2_0_0  );
  input  i_10_2_171_0, i_10_2_174_0, i_10_2_175_0, i_10_2_176_0,
    i_10_2_216_0, i_10_2_217_0, i_10_2_316_0, i_10_2_317_0, i_10_2_318_0,
    i_10_2_321_0, i_10_2_322_0, i_10_2_412_0, i_10_2_429_0, i_10_2_442_0,
    i_10_2_467_0, i_10_2_797_0, i_10_2_800_0, i_10_2_892_0, i_10_2_958_0,
    i_10_2_959_0, i_10_2_1006_0, i_10_2_1026_0, i_10_2_1027_0,
    i_10_2_1029_0, i_10_2_1134_0, i_10_2_1233_0, i_10_2_1234_0,
    i_10_2_1235_0, i_10_2_1236_0, i_10_2_1237_0, i_10_2_1238_0,
    i_10_2_1242_0, i_10_2_1245_0, i_10_2_1306_0, i_10_2_1307_0,
    i_10_2_1579_0, i_10_2_1580_0, i_10_2_1651_0, i_10_2_1652_0,
    i_10_2_1685_0, i_10_2_1819_0, i_10_2_1820_0, i_10_2_1821_0,
    i_10_2_1951_0, i_10_2_1991_0, i_10_2_2184_0, i_10_2_2185_0,
    i_10_2_2311_0, i_10_2_2352_0, i_10_2_2359_0, i_10_2_2361_0,
    i_10_2_2364_0, i_10_2_2376_0, i_10_2_2410_0, i_10_2_2448_0,
    i_10_2_2450_0, i_10_2_2457_0, i_10_2_2458_0, i_10_2_2461_0,
    i_10_2_2462_0, i_10_2_2629_0, i_10_2_2631_0, i_10_2_2635_0,
    i_10_2_2662_0, i_10_2_2719_0, i_10_2_2819_0, i_10_2_2827_0,
    i_10_2_2829_0, i_10_2_2830_0, i_10_2_2918_0, i_10_2_2920_0,
    i_10_2_3093_0, i_10_2_3094_0, i_10_2_3151_0, i_10_2_3276_0,
    i_10_2_3388_0, i_10_2_3391_0, i_10_2_3402_0, i_10_2_3404_0,
    i_10_2_3551_0, i_10_2_3586_0, i_10_2_3609_0, i_10_2_3616_0,
    i_10_2_3647_0, i_10_2_3783_0, i_10_2_3784_0, i_10_2_3787_0,
    i_10_2_3836_0, i_10_2_3838_0, i_10_2_3847_0, i_10_2_3853_0,
    i_10_2_3855_0, i_10_2_3856_0, i_10_2_4127_0, i_10_2_4212_0,
    i_10_2_4269_0, i_10_2_4285_0, i_10_2_4564_0, i_10_2_4566_0,
    i_10_2_4567_0;
  output o_10_2_0_0;
  assign o_10_2_0_0 = ~((~i_10_2_1029_0 & ((i_10_2_175_0 & ((~i_10_2_958_0 & ~i_10_2_2462_0 & ~i_10_2_3094_0) | (~i_10_2_2830_0 & ~i_10_2_3847_0))) | (~i_10_2_1006_0 & ~i_10_2_2185_0 & ~i_10_2_2629_0 & ~i_10_2_3093_0 & ~i_10_2_3388_0 & ~i_10_2_3391_0) | (i_10_2_797_0 & i_10_2_2364_0 & ~i_10_2_2461_0 & ~i_10_2_2631_0 & i_10_2_3838_0) | (~i_10_2_800_0 & ~i_10_2_1238_0 & ~i_10_2_2829_0 & i_10_2_3616_0 & ~i_10_2_3783_0 & ~i_10_2_4269_0))) | (i_10_2_467_0 & ((~i_10_2_2184_0 & ~i_10_2_2311_0 & ~i_10_2_2364_0 & ~i_10_2_2457_0 & ~i_10_2_2829_0 & ~i_10_2_3391_0) | (i_10_2_1652_0 & i_10_2_1819_0 & ~i_10_2_4566_0))) | (~i_10_2_797_0 & ((~i_10_2_467_0 & i_10_2_1236_0 & i_10_2_1237_0 & ~i_10_2_1579_0 & ~i_10_2_3276_0 & ~i_10_2_4566_0) | (~i_10_2_429_0 & ~i_10_2_1236_0 & ~i_10_2_2184_0 & ~i_10_2_2462_0 & ~i_10_2_2629_0 & i_10_2_2635_0 & ~i_10_2_3586_0 & ~i_10_2_4567_0))) | (~i_10_2_429_0 & ((~i_10_2_216_0 & ~i_10_2_2457_0 & ~i_10_2_2662_0 & ~i_10_2_2829_0 & ~i_10_2_3391_0 & ~i_10_2_3402_0 & i_10_2_3838_0 & ~i_10_2_4564_0) | (~i_10_2_1242_0 & i_10_2_1651_0 & ~i_10_2_3388_0 & ~i_10_2_4269_0 & ~i_10_2_4566_0))) | (~i_10_2_2311_0 & ((~i_10_2_2184_0 & ((~i_10_2_216_0 & ((~i_10_2_2185_0 & ~i_10_2_2361_0 & ~i_10_2_2461_0 & ~i_10_2_2462_0 & ~i_10_2_2629_0) | (~i_10_2_2635_0 & ~i_10_2_2827_0 & ~i_10_2_3402_0 & i_10_2_3838_0 & i_10_2_3855_0))) | (~i_10_2_1236_0 & i_10_2_1238_0 & ~i_10_2_3404_0))) | (~i_10_2_3783_0 & ((~i_10_2_467_0 & ((~i_10_2_1006_0 & ~i_10_2_1651_0 & ~i_10_2_1821_0 & ~i_10_2_2462_0 & ~i_10_2_2629_0 & ~i_10_2_2662_0 & ~i_10_2_2920_0) | (~i_10_2_800_0 & ~i_10_2_3093_0 & ~i_10_2_3388_0 & ~i_10_2_3787_0 & ~i_10_2_4212_0 & ~i_10_2_4564_0))) | (~i_10_2_800_0 & ~i_10_2_959_0 & ~i_10_2_1026_0 & ~i_10_2_1245_0 & ~i_10_2_1951_0 & ~i_10_2_1991_0 & ~i_10_2_2410_0 & ~i_10_2_3551_0 & ~i_10_2_3609_0 & ~i_10_2_3784_0))) | (~i_10_2_2359_0 & i_10_2_3647_0))) | (~i_10_2_1027_0 & ((~i_10_2_1821_0 & ~i_10_2_2184_0 & i_10_2_2827_0 & ~i_10_2_2920_0 & ~i_10_2_3609_0 & ~i_10_2_3836_0) | (~i_10_2_2364_0 & ~i_10_2_2410_0 & ~i_10_2_2829_0 & i_10_2_3616_0 & ~i_10_2_3647_0 & ~i_10_2_3856_0))) | (i_10_2_1651_0 & ((~i_10_2_174_0 & ~i_10_2_467_0 & i_10_2_1652_0 & ~i_10_2_3783_0 & ~i_10_2_3838_0) | (i_10_2_3838_0 & i_10_2_4564_0))) | (~i_10_2_2364_0 & ((~i_10_2_2376_0 & ~i_10_2_2457_0 & ~i_10_2_3551_0 & i_10_2_3836_0) | (~i_10_2_2184_0 & ~i_10_2_2185_0 & ~i_10_2_2462_0 & ~i_10_2_2829_0 & ~i_10_2_4212_0))) | (~i_10_2_3855_0 & ((~i_10_2_2461_0 & ((~i_10_2_1242_0 & ~i_10_2_2185_0 & ~i_10_2_2376_0 & ~i_10_2_2830_0 & ~i_10_2_3402_0) | (i_10_2_321_0 & ~i_10_2_3784_0))) | (i_10_2_1238_0 & ~i_10_2_2830_0))) | (~i_10_2_2185_0 & ((~i_10_2_217_0 & ~i_10_2_3551_0 & i_10_2_3609_0 & ~i_10_2_3847_0) | (i_10_2_1307_0 & ~i_10_2_3616_0 & ~i_10_2_4566_0))) | (~i_10_2_2462_0 & ((~i_10_2_892_0 & ~i_10_2_1651_0 & i_10_2_2461_0 & i_10_2_3609_0) | (i_10_2_1821_0 & ~i_10_2_2635_0 & ~i_10_2_3094_0 & ~i_10_2_3783_0 & ~i_10_2_4285_0))) | (~i_10_2_4566_0 & ((i_10_2_174_0 & ~i_10_2_958_0 & i_10_2_2829_0) | (i_10_2_2448_0 & ~i_10_2_2829_0 & ~i_10_2_3647_0))) | (i_10_2_1652_0 & ~i_10_2_2361_0 & i_10_2_3391_0) | (i_10_2_1580_0 & ~i_10_2_2635_0 & ~i_10_2_3783_0));
endmodule



// Benchmark "kernel_10_3" written by ABC on Sun Jul 19 10:21:06 2020

module kernel_10_3 ( 
    i_10_3_176_0, i_10_3_289_0, i_10_3_316_0, i_10_3_325_0, i_10_3_391_0,
    i_10_3_406_0, i_10_3_409_0, i_10_3_433_0, i_10_3_442_0, i_10_3_444_0,
    i_10_3_466_0, i_10_3_622_0, i_10_3_725_0, i_10_3_792_0, i_10_3_955_0,
    i_10_3_1000_0, i_10_3_1027_0, i_10_3_1028_0, i_10_3_1084_0,
    i_10_3_1233_0, i_10_3_1235_0, i_10_3_1244_0, i_10_3_1431_0,
    i_10_3_1432_0, i_10_3_1433_0, i_10_3_1544_0, i_10_3_1577_0,
    i_10_3_1604_0, i_10_3_1683_0, i_10_3_1684_0, i_10_3_1686_0,
    i_10_3_1687_0, i_10_3_1914_0, i_10_3_1921_0, i_10_3_1955_0,
    i_10_3_1981_0, i_10_3_2017_0, i_10_3_2179_0, i_10_3_2349_0,
    i_10_3_2350_0, i_10_3_2351_0, i_10_3_2360_0, i_10_3_2451_0,
    i_10_3_2452_0, i_10_3_2453_0, i_10_3_2530_0, i_10_3_2531_0,
    i_10_3_2567_0, i_10_3_2605_0, i_10_3_2639_0, i_10_3_2655_0,
    i_10_3_2656_0, i_10_3_2657_0, i_10_3_2728_0, i_10_3_2729_0,
    i_10_3_2736_0, i_10_3_2737_0, i_10_3_2754_0, i_10_3_2836_0,
    i_10_3_2844_0, i_10_3_2883_0, i_10_3_2920_0, i_10_3_2921_0,
    i_10_3_3069_0, i_10_3_3072_0, i_10_3_3073_0, i_10_3_3198_0,
    i_10_3_3269_0, i_10_3_3315_0, i_10_3_3330_0, i_10_3_3331_0,
    i_10_3_3332_0, i_10_3_3350_0, i_10_3_3385_0, i_10_3_3386_0,
    i_10_3_3387_0, i_10_3_3406_0, i_10_3_3458_0, i_10_3_3522_0,
    i_10_3_3555_0, i_10_3_3556_0, i_10_3_3587_0, i_10_3_3612_0,
    i_10_3_3837_0, i_10_3_3838_0, i_10_3_3839_0, i_10_3_3848_0,
    i_10_3_3853_0, i_10_3_3855_0, i_10_3_3945_0, i_10_3_4115_0,
    i_10_3_4117_0, i_10_3_4122_0, i_10_3_4150_0, i_10_3_4164_0,
    i_10_3_4172_0, i_10_3_4178_0, i_10_3_4392_0, i_10_3_4428_0,
    i_10_3_4582_0,
    o_10_3_0_0  );
  input  i_10_3_176_0, i_10_3_289_0, i_10_3_316_0, i_10_3_325_0,
    i_10_3_391_0, i_10_3_406_0, i_10_3_409_0, i_10_3_433_0, i_10_3_442_0,
    i_10_3_444_0, i_10_3_466_0, i_10_3_622_0, i_10_3_725_0, i_10_3_792_0,
    i_10_3_955_0, i_10_3_1000_0, i_10_3_1027_0, i_10_3_1028_0,
    i_10_3_1084_0, i_10_3_1233_0, i_10_3_1235_0, i_10_3_1244_0,
    i_10_3_1431_0, i_10_3_1432_0, i_10_3_1433_0, i_10_3_1544_0,
    i_10_3_1577_0, i_10_3_1604_0, i_10_3_1683_0, i_10_3_1684_0,
    i_10_3_1686_0, i_10_3_1687_0, i_10_3_1914_0, i_10_3_1921_0,
    i_10_3_1955_0, i_10_3_1981_0, i_10_3_2017_0, i_10_3_2179_0,
    i_10_3_2349_0, i_10_3_2350_0, i_10_3_2351_0, i_10_3_2360_0,
    i_10_3_2451_0, i_10_3_2452_0, i_10_3_2453_0, i_10_3_2530_0,
    i_10_3_2531_0, i_10_3_2567_0, i_10_3_2605_0, i_10_3_2639_0,
    i_10_3_2655_0, i_10_3_2656_0, i_10_3_2657_0, i_10_3_2728_0,
    i_10_3_2729_0, i_10_3_2736_0, i_10_3_2737_0, i_10_3_2754_0,
    i_10_3_2836_0, i_10_3_2844_0, i_10_3_2883_0, i_10_3_2920_0,
    i_10_3_2921_0, i_10_3_3069_0, i_10_3_3072_0, i_10_3_3073_0,
    i_10_3_3198_0, i_10_3_3269_0, i_10_3_3315_0, i_10_3_3330_0,
    i_10_3_3331_0, i_10_3_3332_0, i_10_3_3350_0, i_10_3_3385_0,
    i_10_3_3386_0, i_10_3_3387_0, i_10_3_3406_0, i_10_3_3458_0,
    i_10_3_3522_0, i_10_3_3555_0, i_10_3_3556_0, i_10_3_3587_0,
    i_10_3_3612_0, i_10_3_3837_0, i_10_3_3838_0, i_10_3_3839_0,
    i_10_3_3848_0, i_10_3_3853_0, i_10_3_3855_0, i_10_3_3945_0,
    i_10_3_4115_0, i_10_3_4117_0, i_10_3_4122_0, i_10_3_4150_0,
    i_10_3_4164_0, i_10_3_4172_0, i_10_3_4178_0, i_10_3_4392_0,
    i_10_3_4428_0, i_10_3_4582_0;
  output o_10_3_0_0;
  assign o_10_3_0_0 = 0;
endmodule



// Benchmark "kernel_10_4" written by ABC on Sun Jul 19 10:21:07 2020

module kernel_10_4 ( 
    i_10_4_63_0, i_10_4_89_0, i_10_4_144_0, i_10_4_148_0, i_10_4_263_0,
    i_10_4_283_0, i_10_4_287_0, i_10_4_329_0, i_10_4_408_0, i_10_4_424_0,
    i_10_4_427_0, i_10_4_464_0, i_10_4_532_0, i_10_4_556_0, i_10_4_796_0,
    i_10_4_933_0, i_10_4_963_0, i_10_4_1003_0, i_10_4_1058_0,
    i_10_4_1198_0, i_10_4_1267_0, i_10_4_1306_0, i_10_4_1307_0,
    i_10_4_1308_0, i_10_4_1485_0, i_10_4_1488_0, i_10_4_1489_0,
    i_10_4_1619_0, i_10_4_1653_0, i_10_4_1654_0, i_10_4_1795_0,
    i_10_4_1804_0, i_10_4_1818_0, i_10_4_1917_0, i_10_4_1929_0,
    i_10_4_1937_0, i_10_4_1948_0, i_10_4_1949_0, i_10_4_2028_0,
    i_10_4_2182_0, i_10_4_2244_0, i_10_4_2247_0, i_10_4_2336_0,
    i_10_4_2361_0, i_10_4_2364_0, i_10_4_2430_0, i_10_4_2448_0,
    i_10_4_2449_0, i_10_4_2451_0, i_10_4_2454_0, i_10_4_2469_0,
    i_10_4_2479_0, i_10_4_2513_0, i_10_4_2515_0, i_10_4_2516_0,
    i_10_4_2542_0, i_10_4_2544_0, i_10_4_2662_0, i_10_4_2663_0,
    i_10_4_2710_0, i_10_4_2713_0, i_10_4_2724_0, i_10_4_2789_0,
    i_10_4_2821_0, i_10_4_2834_0, i_10_4_3043_0, i_10_4_3070_0,
    i_10_4_3073_0, i_10_4_3235_0, i_10_4_3280_0, i_10_4_3282_0,
    i_10_4_3283_0, i_10_4_3312_0, i_10_4_3315_0, i_10_4_3384_0,
    i_10_4_3385_0, i_10_4_3401_0, i_10_4_3454_0, i_10_4_3611_0,
    i_10_4_3616_0, i_10_4_3645_0, i_10_4_3685_0, i_10_4_3725_0,
    i_10_4_3856_0, i_10_4_3888_0, i_10_4_3891_0, i_10_4_3909_0,
    i_10_4_3942_0, i_10_4_4116_0, i_10_4_4156_0, i_10_4_4237_0,
    i_10_4_4279_0, i_10_4_4287_0, i_10_4_4288_0, i_10_4_4289_0,
    i_10_4_4396_0, i_10_4_4397_0, i_10_4_4531_0, i_10_4_4582_0,
    i_10_4_4583_0,
    o_10_4_0_0  );
  input  i_10_4_63_0, i_10_4_89_0, i_10_4_144_0, i_10_4_148_0,
    i_10_4_263_0, i_10_4_283_0, i_10_4_287_0, i_10_4_329_0, i_10_4_408_0,
    i_10_4_424_0, i_10_4_427_0, i_10_4_464_0, i_10_4_532_0, i_10_4_556_0,
    i_10_4_796_0, i_10_4_933_0, i_10_4_963_0, i_10_4_1003_0, i_10_4_1058_0,
    i_10_4_1198_0, i_10_4_1267_0, i_10_4_1306_0, i_10_4_1307_0,
    i_10_4_1308_0, i_10_4_1485_0, i_10_4_1488_0, i_10_4_1489_0,
    i_10_4_1619_0, i_10_4_1653_0, i_10_4_1654_0, i_10_4_1795_0,
    i_10_4_1804_0, i_10_4_1818_0, i_10_4_1917_0, i_10_4_1929_0,
    i_10_4_1937_0, i_10_4_1948_0, i_10_4_1949_0, i_10_4_2028_0,
    i_10_4_2182_0, i_10_4_2244_0, i_10_4_2247_0, i_10_4_2336_0,
    i_10_4_2361_0, i_10_4_2364_0, i_10_4_2430_0, i_10_4_2448_0,
    i_10_4_2449_0, i_10_4_2451_0, i_10_4_2454_0, i_10_4_2469_0,
    i_10_4_2479_0, i_10_4_2513_0, i_10_4_2515_0, i_10_4_2516_0,
    i_10_4_2542_0, i_10_4_2544_0, i_10_4_2662_0, i_10_4_2663_0,
    i_10_4_2710_0, i_10_4_2713_0, i_10_4_2724_0, i_10_4_2789_0,
    i_10_4_2821_0, i_10_4_2834_0, i_10_4_3043_0, i_10_4_3070_0,
    i_10_4_3073_0, i_10_4_3235_0, i_10_4_3280_0, i_10_4_3282_0,
    i_10_4_3283_0, i_10_4_3312_0, i_10_4_3315_0, i_10_4_3384_0,
    i_10_4_3385_0, i_10_4_3401_0, i_10_4_3454_0, i_10_4_3611_0,
    i_10_4_3616_0, i_10_4_3645_0, i_10_4_3685_0, i_10_4_3725_0,
    i_10_4_3856_0, i_10_4_3888_0, i_10_4_3891_0, i_10_4_3909_0,
    i_10_4_3942_0, i_10_4_4116_0, i_10_4_4156_0, i_10_4_4237_0,
    i_10_4_4279_0, i_10_4_4287_0, i_10_4_4288_0, i_10_4_4289_0,
    i_10_4_4396_0, i_10_4_4397_0, i_10_4_4531_0, i_10_4_4582_0,
    i_10_4_4583_0;
  output o_10_4_0_0;
  assign o_10_4_0_0 = 0;
endmodule



// Benchmark "kernel_10_5" written by ABC on Sun Jul 19 10:21:08 2020

module kernel_10_5 ( 
    i_10_5_27_0, i_10_5_45_0, i_10_5_146_0, i_10_5_203_0, i_10_5_222_0,
    i_10_5_243_0, i_10_5_252_0, i_10_5_279_0, i_10_5_286_0, i_10_5_287_0,
    i_10_5_288_0, i_10_5_465_0, i_10_5_466_0, i_10_5_467_0, i_10_5_503_0,
    i_10_5_517_0, i_10_5_558_0, i_10_5_747_0, i_10_5_748_0, i_10_5_798_0,
    i_10_5_845_0, i_10_5_954_0, i_10_5_955_0, i_10_5_1026_0, i_10_5_1031_0,
    i_10_5_1197_0, i_10_5_1233_0, i_10_5_1234_0, i_10_5_1236_0,
    i_10_5_1237_0, i_10_5_1239_0, i_10_5_1240_0, i_10_5_1241_0,
    i_10_5_1242_0, i_10_5_1243_0, i_10_5_1274_0, i_10_5_1311_0,
    i_10_5_1373_0, i_10_5_1378_0, i_10_5_1616_0, i_10_5_1648_0,
    i_10_5_1649_0, i_10_5_1757_0, i_10_5_1824_0, i_10_5_1912_0,
    i_10_5_1953_0, i_10_5_1957_0, i_10_5_1961_0, i_10_5_2161_0,
    i_10_5_2178_0, i_10_5_2196_0, i_10_5_2197_0, i_10_5_2254_0,
    i_10_5_2303_0, i_10_5_2307_0, i_10_5_2354_0, i_10_5_2357_0,
    i_10_5_2449_0, i_10_5_2450_0, i_10_5_2451_0, i_10_5_2454_0,
    i_10_5_2458_0, i_10_5_2469_0, i_10_5_2470_0, i_10_5_2489_0,
    i_10_5_2605_0, i_10_5_2608_0, i_10_5_2628_0, i_10_5_2629_0,
    i_10_5_2630_0, i_10_5_2646_0, i_10_5_2680_0, i_10_5_2696_0,
    i_10_5_2701_0, i_10_5_2732_0, i_10_5_2833_0, i_10_5_2886_0,
    i_10_5_2948_0, i_10_5_2960_0, i_10_5_3267_0, i_10_5_3268_0,
    i_10_5_3279_0, i_10_5_3289_0, i_10_5_3292_0, i_10_5_3301_0,
    i_10_5_3384_0, i_10_5_3387_0, i_10_5_3473_0, i_10_5_3588_0,
    i_10_5_3589_0, i_10_5_3625_0, i_10_5_3649_0, i_10_5_3724_0,
    i_10_5_3780_0, i_10_5_3783_0, i_10_5_3853_0, i_10_5_4165_0,
    i_10_5_4319_0, i_10_5_4586_0, i_10_5_4588_0,
    o_10_5_0_0  );
  input  i_10_5_27_0, i_10_5_45_0, i_10_5_146_0, i_10_5_203_0,
    i_10_5_222_0, i_10_5_243_0, i_10_5_252_0, i_10_5_279_0, i_10_5_286_0,
    i_10_5_287_0, i_10_5_288_0, i_10_5_465_0, i_10_5_466_0, i_10_5_467_0,
    i_10_5_503_0, i_10_5_517_0, i_10_5_558_0, i_10_5_747_0, i_10_5_748_0,
    i_10_5_798_0, i_10_5_845_0, i_10_5_954_0, i_10_5_955_0, i_10_5_1026_0,
    i_10_5_1031_0, i_10_5_1197_0, i_10_5_1233_0, i_10_5_1234_0,
    i_10_5_1236_0, i_10_5_1237_0, i_10_5_1239_0, i_10_5_1240_0,
    i_10_5_1241_0, i_10_5_1242_0, i_10_5_1243_0, i_10_5_1274_0,
    i_10_5_1311_0, i_10_5_1373_0, i_10_5_1378_0, i_10_5_1616_0,
    i_10_5_1648_0, i_10_5_1649_0, i_10_5_1757_0, i_10_5_1824_0,
    i_10_5_1912_0, i_10_5_1953_0, i_10_5_1957_0, i_10_5_1961_0,
    i_10_5_2161_0, i_10_5_2178_0, i_10_5_2196_0, i_10_5_2197_0,
    i_10_5_2254_0, i_10_5_2303_0, i_10_5_2307_0, i_10_5_2354_0,
    i_10_5_2357_0, i_10_5_2449_0, i_10_5_2450_0, i_10_5_2451_0,
    i_10_5_2454_0, i_10_5_2458_0, i_10_5_2469_0, i_10_5_2470_0,
    i_10_5_2489_0, i_10_5_2605_0, i_10_5_2608_0, i_10_5_2628_0,
    i_10_5_2629_0, i_10_5_2630_0, i_10_5_2646_0, i_10_5_2680_0,
    i_10_5_2696_0, i_10_5_2701_0, i_10_5_2732_0, i_10_5_2833_0,
    i_10_5_2886_0, i_10_5_2948_0, i_10_5_2960_0, i_10_5_3267_0,
    i_10_5_3268_0, i_10_5_3279_0, i_10_5_3289_0, i_10_5_3292_0,
    i_10_5_3301_0, i_10_5_3384_0, i_10_5_3387_0, i_10_5_3473_0,
    i_10_5_3588_0, i_10_5_3589_0, i_10_5_3625_0, i_10_5_3649_0,
    i_10_5_3724_0, i_10_5_3780_0, i_10_5_3783_0, i_10_5_3853_0,
    i_10_5_4165_0, i_10_5_4319_0, i_10_5_4586_0, i_10_5_4588_0;
  output o_10_5_0_0;
  assign o_10_5_0_0 = 0;
endmodule



// Benchmark "kernel_10_6" written by ABC on Sun Jul 19 10:21:08 2020

module kernel_10_6 ( 
    i_10_6_30_0, i_10_6_51_0, i_10_6_52_0, i_10_6_53_0, i_10_6_142_0,
    i_10_6_143_0, i_10_6_151_0, i_10_6_243_0, i_10_6_252_0, i_10_6_271_0,
    i_10_6_272_0, i_10_6_350_0, i_10_6_358_0, i_10_6_430_0, i_10_6_464_0,
    i_10_6_495_0, i_10_6_514_0, i_10_6_517_0, i_10_6_518_0, i_10_6_591_0,
    i_10_6_714_0, i_10_6_754_0, i_10_6_755_0, i_10_6_799_0, i_10_6_831_0,
    i_10_6_832_0, i_10_6_970_0, i_10_6_988_0, i_10_6_997_0, i_10_6_1082_0,
    i_10_6_1166_0, i_10_6_1209_0, i_10_6_1240_0, i_10_6_1357_0,
    i_10_6_1367_0, i_10_6_1384_0, i_10_6_1446_0, i_10_6_1635_0,
    i_10_6_1636_0, i_10_6_1645_0, i_10_6_1690_0, i_10_6_1764_0,
    i_10_6_1768_0, i_10_6_1805_0, i_10_6_1808_0, i_10_6_1824_0,
    i_10_6_1825_0, i_10_6_1918_0, i_10_6_1952_0, i_10_6_1959_0,
    i_10_6_2004_0, i_10_6_2031_0, i_10_6_2182_0, i_10_6_2185_0,
    i_10_6_2247_0, i_10_6_2312_0, i_10_6_2329_0, i_10_6_2360_0,
    i_10_6_2390_0, i_10_6_2452_0, i_10_6_2510_0, i_10_6_2573_0,
    i_10_6_2602_0, i_10_6_2614_0, i_10_6_2741_0, i_10_6_2882_0,
    i_10_6_2913_0, i_10_6_2984_0, i_10_6_3122_0, i_10_6_3202_0,
    i_10_6_3315_0, i_10_6_3410_0, i_10_6_3473_0, i_10_6_3497_0,
    i_10_6_3547_0, i_10_6_3586_0, i_10_6_3587_0, i_10_6_3684_0,
    i_10_6_3688_0, i_10_6_3721_0, i_10_6_3822_0, i_10_6_3849_0,
    i_10_6_3850_0, i_10_6_3851_0, i_10_6_3854_0, i_10_6_3856_0,
    i_10_6_3878_0, i_10_6_3912_0, i_10_6_3985_0, i_10_6_4028_0,
    i_10_6_4116_0, i_10_6_4117_0, i_10_6_4119_0, i_10_6_4120_0,
    i_10_6_4121_0, i_10_6_4266_0, i_10_6_4269_0, i_10_6_4289_0,
    i_10_6_4459_0, i_10_6_4463_0,
    o_10_6_0_0  );
  input  i_10_6_30_0, i_10_6_51_0, i_10_6_52_0, i_10_6_53_0,
    i_10_6_142_0, i_10_6_143_0, i_10_6_151_0, i_10_6_243_0, i_10_6_252_0,
    i_10_6_271_0, i_10_6_272_0, i_10_6_350_0, i_10_6_358_0, i_10_6_430_0,
    i_10_6_464_0, i_10_6_495_0, i_10_6_514_0, i_10_6_517_0, i_10_6_518_0,
    i_10_6_591_0, i_10_6_714_0, i_10_6_754_0, i_10_6_755_0, i_10_6_799_0,
    i_10_6_831_0, i_10_6_832_0, i_10_6_970_0, i_10_6_988_0, i_10_6_997_0,
    i_10_6_1082_0, i_10_6_1166_0, i_10_6_1209_0, i_10_6_1240_0,
    i_10_6_1357_0, i_10_6_1367_0, i_10_6_1384_0, i_10_6_1446_0,
    i_10_6_1635_0, i_10_6_1636_0, i_10_6_1645_0, i_10_6_1690_0,
    i_10_6_1764_0, i_10_6_1768_0, i_10_6_1805_0, i_10_6_1808_0,
    i_10_6_1824_0, i_10_6_1825_0, i_10_6_1918_0, i_10_6_1952_0,
    i_10_6_1959_0, i_10_6_2004_0, i_10_6_2031_0, i_10_6_2182_0,
    i_10_6_2185_0, i_10_6_2247_0, i_10_6_2312_0, i_10_6_2329_0,
    i_10_6_2360_0, i_10_6_2390_0, i_10_6_2452_0, i_10_6_2510_0,
    i_10_6_2573_0, i_10_6_2602_0, i_10_6_2614_0, i_10_6_2741_0,
    i_10_6_2882_0, i_10_6_2913_0, i_10_6_2984_0, i_10_6_3122_0,
    i_10_6_3202_0, i_10_6_3315_0, i_10_6_3410_0, i_10_6_3473_0,
    i_10_6_3497_0, i_10_6_3547_0, i_10_6_3586_0, i_10_6_3587_0,
    i_10_6_3684_0, i_10_6_3688_0, i_10_6_3721_0, i_10_6_3822_0,
    i_10_6_3849_0, i_10_6_3850_0, i_10_6_3851_0, i_10_6_3854_0,
    i_10_6_3856_0, i_10_6_3878_0, i_10_6_3912_0, i_10_6_3985_0,
    i_10_6_4028_0, i_10_6_4116_0, i_10_6_4117_0, i_10_6_4119_0,
    i_10_6_4120_0, i_10_6_4121_0, i_10_6_4266_0, i_10_6_4269_0,
    i_10_6_4289_0, i_10_6_4459_0, i_10_6_4463_0;
  output o_10_6_0_0;
  assign o_10_6_0_0 = 0;
endmodule



// Benchmark "kernel_10_7" written by ABC on Sun Jul 19 10:21:09 2020

module kernel_10_7 ( 
    i_10_7_40_0, i_10_7_173_0, i_10_7_184_0, i_10_7_185_0, i_10_7_188_0,
    i_10_7_271_0, i_10_7_272_0, i_10_7_283_0, i_10_7_285_0, i_10_7_370_0,
    i_10_7_390_0, i_10_7_391_0, i_10_7_461_0, i_10_7_463_0, i_10_7_464_0,
    i_10_7_465_0, i_10_7_502_0, i_10_7_563_0, i_10_7_751_0, i_10_7_754_0,
    i_10_7_905_0, i_10_7_917_0, i_10_7_933_0, i_10_7_934_0, i_10_7_965_0,
    i_10_7_966_0, i_10_7_1056_0, i_10_7_1234_0, i_10_7_1235_0,
    i_10_7_1241_0, i_10_7_1312_0, i_10_7_1348_0, i_10_7_1366_0,
    i_10_7_1543_0, i_10_7_1552_0, i_10_7_1645_0, i_10_7_1652_0,
    i_10_7_1686_0, i_10_7_1714_0, i_10_7_1767_0, i_10_7_1812_0,
    i_10_7_1813_0, i_10_7_1819_0, i_10_7_1822_0, i_10_7_1907_0,
    i_10_7_1922_0, i_10_7_1950_0, i_10_7_1957_0, i_10_7_1991_0,
    i_10_7_2023_0, i_10_7_2184_0, i_10_7_2247_0, i_10_7_2309_0,
    i_10_7_2388_0, i_10_7_2451_0, i_10_7_2467_0, i_10_7_2511_0,
    i_10_7_2516_0, i_10_7_2540_0, i_10_7_2602_0, i_10_7_2617_0,
    i_10_7_2735_0, i_10_7_2743_0, i_10_7_2789_0, i_10_7_2806_0,
    i_10_7_2807_0, i_10_7_2825_0, i_10_7_2827_0, i_10_7_2980_0,
    i_10_7_3198_0, i_10_7_3200_0, i_10_7_3328_0, i_10_7_3352_0,
    i_10_7_3353_0, i_10_7_3454_0, i_10_7_3469_0, i_10_7_3470_0,
    i_10_7_3525_0, i_10_7_3582_0, i_10_7_3588_0, i_10_7_3590_0,
    i_10_7_3622_0, i_10_7_3625_0, i_10_7_3685_0, i_10_7_3723_0,
    i_10_7_3839_0, i_10_7_3855_0, i_10_7_3856_0, i_10_7_3860_0,
    i_10_7_3881_0, i_10_7_3895_0, i_10_7_3946_0, i_10_7_3950_0,
    i_10_7_4054_0, i_10_7_4113_0, i_10_7_4118_0, i_10_7_4217_0,
    i_10_7_4237_0, i_10_7_4267_0, i_10_7_4295_0,
    o_10_7_0_0  );
  input  i_10_7_40_0, i_10_7_173_0, i_10_7_184_0, i_10_7_185_0,
    i_10_7_188_0, i_10_7_271_0, i_10_7_272_0, i_10_7_283_0, i_10_7_285_0,
    i_10_7_370_0, i_10_7_390_0, i_10_7_391_0, i_10_7_461_0, i_10_7_463_0,
    i_10_7_464_0, i_10_7_465_0, i_10_7_502_0, i_10_7_563_0, i_10_7_751_0,
    i_10_7_754_0, i_10_7_905_0, i_10_7_917_0, i_10_7_933_0, i_10_7_934_0,
    i_10_7_965_0, i_10_7_966_0, i_10_7_1056_0, i_10_7_1234_0,
    i_10_7_1235_0, i_10_7_1241_0, i_10_7_1312_0, i_10_7_1348_0,
    i_10_7_1366_0, i_10_7_1543_0, i_10_7_1552_0, i_10_7_1645_0,
    i_10_7_1652_0, i_10_7_1686_0, i_10_7_1714_0, i_10_7_1767_0,
    i_10_7_1812_0, i_10_7_1813_0, i_10_7_1819_0, i_10_7_1822_0,
    i_10_7_1907_0, i_10_7_1922_0, i_10_7_1950_0, i_10_7_1957_0,
    i_10_7_1991_0, i_10_7_2023_0, i_10_7_2184_0, i_10_7_2247_0,
    i_10_7_2309_0, i_10_7_2388_0, i_10_7_2451_0, i_10_7_2467_0,
    i_10_7_2511_0, i_10_7_2516_0, i_10_7_2540_0, i_10_7_2602_0,
    i_10_7_2617_0, i_10_7_2735_0, i_10_7_2743_0, i_10_7_2789_0,
    i_10_7_2806_0, i_10_7_2807_0, i_10_7_2825_0, i_10_7_2827_0,
    i_10_7_2980_0, i_10_7_3198_0, i_10_7_3200_0, i_10_7_3328_0,
    i_10_7_3352_0, i_10_7_3353_0, i_10_7_3454_0, i_10_7_3469_0,
    i_10_7_3470_0, i_10_7_3525_0, i_10_7_3582_0, i_10_7_3588_0,
    i_10_7_3590_0, i_10_7_3622_0, i_10_7_3625_0, i_10_7_3685_0,
    i_10_7_3723_0, i_10_7_3839_0, i_10_7_3855_0, i_10_7_3856_0,
    i_10_7_3860_0, i_10_7_3881_0, i_10_7_3895_0, i_10_7_3946_0,
    i_10_7_3950_0, i_10_7_4054_0, i_10_7_4113_0, i_10_7_4118_0,
    i_10_7_4217_0, i_10_7_4237_0, i_10_7_4267_0, i_10_7_4295_0;
  output o_10_7_0_0;
  assign o_10_7_0_0 = 0;
endmodule



// Benchmark "kernel_10_8" written by ABC on Sun Jul 19 10:21:11 2020

module kernel_10_8 ( 
    i_10_8_124_0, i_10_8_174_0, i_10_8_175_0, i_10_8_176_0, i_10_8_220_0,
    i_10_8_223_0, i_10_8_283_0, i_10_8_284_0, i_10_8_328_0, i_10_8_329_0,
    i_10_8_395_0, i_10_8_433_0, i_10_8_434_0, i_10_8_442_0, i_10_8_465_0,
    i_10_8_518_0, i_10_8_565_0, i_10_8_793_0, i_10_8_907_0, i_10_8_954_0,
    i_10_8_968_0, i_10_8_991_0, i_10_8_1006_0, i_10_8_1033_0,
    i_10_8_1309_0, i_10_8_1310_0, i_10_8_1349_0, i_10_8_1367_0,
    i_10_8_1379_0, i_10_8_1439_0, i_10_8_1555_0, i_10_8_1556_0,
    i_10_8_1684_0, i_10_8_1685_0, i_10_8_1687_0, i_10_8_1768_0,
    i_10_8_1769_0, i_10_8_1810_0, i_10_8_1819_0, i_10_8_1824_0,
    i_10_8_1951_0, i_10_8_1952_0, i_10_8_2029_0, i_10_8_2185_0,
    i_10_8_2186_0, i_10_8_2201_0, i_10_8_2311_0, i_10_8_2312_0,
    i_10_8_2351_0, i_10_8_2353_0, i_10_8_2362_0, i_10_8_2410_0,
    i_10_8_2411_0, i_10_8_2449_0, i_10_8_2450_0, i_10_8_2451_0,
    i_10_8_2455_0, i_10_8_2504_0, i_10_8_2572_0, i_10_8_2603_0,
    i_10_8_2629_0, i_10_8_2632_0, i_10_8_2657_0, i_10_8_2659_0,
    i_10_8_2660_0, i_10_8_2680_0, i_10_8_2681_0, i_10_8_2705_0,
    i_10_8_2722_0, i_10_8_2723_0, i_10_8_2725_0, i_10_8_2729_0,
    i_10_8_2730_0, i_10_8_2731_0, i_10_8_2789_0, i_10_8_2829_0,
    i_10_8_2830_0, i_10_8_2923_0, i_10_8_2924_0, i_10_8_3047_0,
    i_10_8_3076_0, i_10_8_3158_0, i_10_8_3497_0, i_10_8_3609_0,
    i_10_8_3624_0, i_10_8_3650_0, i_10_8_3836_0, i_10_8_3844_0,
    i_10_8_3846_0, i_10_8_3855_0, i_10_8_3857_0, i_10_8_3912_0,
    i_10_8_3914_0, i_10_8_3986_0, i_10_8_4058_0, i_10_8_4118_0,
    i_10_8_4237_0, i_10_8_4285_0, i_10_8_4288_0, i_10_8_4289_0,
    o_10_8_0_0  );
  input  i_10_8_124_0, i_10_8_174_0, i_10_8_175_0, i_10_8_176_0,
    i_10_8_220_0, i_10_8_223_0, i_10_8_283_0, i_10_8_284_0, i_10_8_328_0,
    i_10_8_329_0, i_10_8_395_0, i_10_8_433_0, i_10_8_434_0, i_10_8_442_0,
    i_10_8_465_0, i_10_8_518_0, i_10_8_565_0, i_10_8_793_0, i_10_8_907_0,
    i_10_8_954_0, i_10_8_968_0, i_10_8_991_0, i_10_8_1006_0, i_10_8_1033_0,
    i_10_8_1309_0, i_10_8_1310_0, i_10_8_1349_0, i_10_8_1367_0,
    i_10_8_1379_0, i_10_8_1439_0, i_10_8_1555_0, i_10_8_1556_0,
    i_10_8_1684_0, i_10_8_1685_0, i_10_8_1687_0, i_10_8_1768_0,
    i_10_8_1769_0, i_10_8_1810_0, i_10_8_1819_0, i_10_8_1824_0,
    i_10_8_1951_0, i_10_8_1952_0, i_10_8_2029_0, i_10_8_2185_0,
    i_10_8_2186_0, i_10_8_2201_0, i_10_8_2311_0, i_10_8_2312_0,
    i_10_8_2351_0, i_10_8_2353_0, i_10_8_2362_0, i_10_8_2410_0,
    i_10_8_2411_0, i_10_8_2449_0, i_10_8_2450_0, i_10_8_2451_0,
    i_10_8_2455_0, i_10_8_2504_0, i_10_8_2572_0, i_10_8_2603_0,
    i_10_8_2629_0, i_10_8_2632_0, i_10_8_2657_0, i_10_8_2659_0,
    i_10_8_2660_0, i_10_8_2680_0, i_10_8_2681_0, i_10_8_2705_0,
    i_10_8_2722_0, i_10_8_2723_0, i_10_8_2725_0, i_10_8_2729_0,
    i_10_8_2730_0, i_10_8_2731_0, i_10_8_2789_0, i_10_8_2829_0,
    i_10_8_2830_0, i_10_8_2923_0, i_10_8_2924_0, i_10_8_3047_0,
    i_10_8_3076_0, i_10_8_3158_0, i_10_8_3497_0, i_10_8_3609_0,
    i_10_8_3624_0, i_10_8_3650_0, i_10_8_3836_0, i_10_8_3844_0,
    i_10_8_3846_0, i_10_8_3855_0, i_10_8_3857_0, i_10_8_3912_0,
    i_10_8_3914_0, i_10_8_3986_0, i_10_8_4058_0, i_10_8_4118_0,
    i_10_8_4237_0, i_10_8_4285_0, i_10_8_4288_0, i_10_8_4289_0;
  output o_10_8_0_0;
  assign o_10_8_0_0 = ~((~i_10_8_2680_0 & ((~i_10_8_433_0 & ((~i_10_8_434_0 & ~i_10_8_1951_0 & ~i_10_8_2186_0 & ~i_10_8_2311_0 & ~i_10_8_2411_0 & ~i_10_8_2657_0 & ~i_10_8_2723_0 & ~i_10_8_2789_0 & ~i_10_8_2829_0 & ~i_10_8_3855_0 & ~i_10_8_3857_0) | (~i_10_8_565_0 & ~i_10_8_907_0 & ~i_10_8_1349_0 & ~i_10_8_1555_0 & ~i_10_8_1810_0 & ~i_10_8_2312_0 & ~i_10_8_2504_0 & ~i_10_8_2603_0 & i_10_8_2731_0 & ~i_10_8_4058_0 & ~i_10_8_4237_0 & ~i_10_8_4288_0))) | (~i_10_8_328_0 & ~i_10_8_395_0 & ~i_10_8_991_0 & ~i_10_8_1006_0 & ~i_10_8_1952_0 & ~i_10_8_2353_0 & ~i_10_8_2504_0 & ~i_10_8_2657_0 & ~i_10_8_3076_0 & ~i_10_8_3609_0))) | (~i_10_8_907_0 & ((i_10_8_174_0 & ~i_10_8_329_0 & ~i_10_8_395_0 & ~i_10_8_1768_0 & ~i_10_8_2411_0) | (~i_10_8_124_0 & ~i_10_8_442_0 & ~i_10_8_1310_0 & ~i_10_8_1769_0 & ~i_10_8_1810_0 & ~i_10_8_1952_0 & ~i_10_8_2603_0 & ~i_10_8_2829_0 & ~i_10_8_3650_0 & ~i_10_8_3857_0 & ~i_10_8_4058_0 & ~i_10_8_4237_0))) | (~i_10_8_284_0 & ((~i_10_8_124_0 & ((~i_10_8_328_0 & ~i_10_8_434_0 & ~i_10_8_565_0 & ~i_10_8_1684_0 & ~i_10_8_2312_0 & i_10_8_2353_0 & ~i_10_8_2705_0 & ~i_10_8_2830_0) | (~i_10_8_1006_0 & i_10_8_3912_0))) | (~i_10_8_328_0 & ~i_10_8_954_0 & ~i_10_8_1768_0 & ~i_10_8_2201_0 & ~i_10_8_2603_0 & i_10_8_2629_0 & ~i_10_8_2705_0 & ~i_10_8_2731_0 & ~i_10_8_3047_0 & ~i_10_8_3836_0) | (~i_10_8_1006_0 & ~i_10_8_1951_0 & i_10_8_2680_0 & ~i_10_8_2723_0 & ~i_10_8_3076_0 & ~i_10_8_3855_0))) | (~i_10_8_2312_0 & ((~i_10_8_328_0 & ~i_10_8_2504_0 & ((~i_10_8_2410_0 & i_10_8_2450_0) | (~i_10_8_1309_0 & ~i_10_8_1555_0 & ~i_10_8_1768_0 & ~i_10_8_2186_0 & ~i_10_8_2657_0 & ~i_10_8_4058_0))) | (~i_10_8_565_0 & ((i_10_8_518_0 & ~i_10_8_1556_0 & ~i_10_8_2659_0 & ~i_10_8_2723_0 & ~i_10_8_2924_0 & ~i_10_8_4118_0) | (~i_10_8_1310_0 & i_10_8_2632_0 & ~i_10_8_2657_0 & ~i_10_8_2705_0 & ~i_10_8_2830_0 & ~i_10_8_3844_0 & ~i_10_8_4237_0))) | (~i_10_8_4237_0 & ((~i_10_8_1006_0 & ~i_10_8_1310_0 & ~i_10_8_1810_0 & ~i_10_8_2632_0 & i_10_8_2731_0 & i_10_8_3855_0) | (i_10_8_283_0 & ~i_10_8_329_0 & ~i_10_8_465_0 & ~i_10_8_991_0 & ~i_10_8_2410_0 & ~i_10_8_2455_0 & ~i_10_8_2629_0 & ~i_10_8_3650_0 & ~i_10_8_3836_0 & ~i_10_8_3986_0 & ~i_10_8_4058_0))) | (i_10_8_223_0 & i_10_8_2829_0 & i_10_8_3846_0))) | (~i_10_8_395_0 & ((i_10_8_1684_0 & ~i_10_8_2351_0 & ~i_10_8_2410_0) | (~i_10_8_991_0 & i_10_8_1687_0 & ~i_10_8_1810_0 & ~i_10_8_2353_0 & ~i_10_8_2504_0))) | (~i_10_8_434_0 & ((~i_10_8_1439_0 & ~i_10_8_1555_0 & ~i_10_8_1556_0 & ~i_10_8_2311_0 & ~i_10_8_2353_0 & ~i_10_8_2504_0 & ~i_10_8_2659_0) | (~i_10_8_1768_0 & ~i_10_8_1769_0 & ~i_10_8_2186_0 & i_10_8_4288_0))) | (~i_10_8_1310_0 & ((i_10_8_2186_0 & ~i_10_8_2729_0 & ~i_10_8_2830_0 & ~i_10_8_3855_0 & i_10_8_3857_0) | (~i_10_8_329_0 & i_10_8_793_0 & ~i_10_8_1810_0 & ~i_10_8_2353_0 & ~i_10_8_4237_0))) | (~i_10_8_1810_0 & ((~i_10_8_518_0 & ~i_10_8_954_0 & ~i_10_8_1439_0 & ~i_10_8_1768_0 & i_10_8_2632_0 & ~i_10_8_2681_0 & i_10_8_2830_0 & ~i_10_8_3047_0 & i_10_8_4118_0) | (~i_10_8_1006_0 & ~i_10_8_1555_0 & ~i_10_8_1687_0 & ~i_10_8_2185_0 & ~i_10_8_2186_0 & ~i_10_8_2351_0 & ~i_10_8_2603_0 & ~i_10_8_2657_0 & ~i_10_8_2660_0 & ~i_10_8_2722_0 & ~i_10_8_2729_0 & ~i_10_8_2829_0 & ~i_10_8_4058_0 & ~i_10_8_4289_0))) | (i_10_8_2924_0 & ((i_10_8_2186_0 & i_10_8_2504_0) | (i_10_8_2923_0 & ~i_10_8_4237_0))) | (~i_10_8_3986_0 & ((~i_10_8_2451_0 & i_10_8_2455_0 & ~i_10_8_2660_0 & i_10_8_3855_0) | (i_10_8_2632_0 & i_10_8_4288_0 & ~i_10_8_4289_0))) | (~i_10_8_283_0 & ~i_10_8_565_0 & i_10_8_1687_0 & i_10_8_2353_0 & ~i_10_8_3857_0) | (~i_10_8_991_0 & ~i_10_8_2185_0 & ~i_10_8_2632_0 & i_10_8_2722_0 & ~i_10_8_2725_0 & i_10_8_2829_0 & ~i_10_8_3855_0 & ~i_10_8_4237_0));
endmodule



// Benchmark "kernel_10_9" written by ABC on Sun Jul 19 10:21:11 2020

module kernel_10_9 ( 
    i_10_9_47_0, i_10_9_146_0, i_10_9_171_0, i_10_9_176_0, i_10_9_191_0,
    i_10_9_224_0, i_10_9_247_0, i_10_9_279_0, i_10_9_281_0, i_10_9_287_0,
    i_10_9_315_0, i_10_9_317_0, i_10_9_443_0, i_10_9_459_0, i_10_9_462_0,
    i_10_9_463_0, i_10_9_464_0, i_10_9_509_0, i_10_9_635_0, i_10_9_821_0,
    i_10_9_891_0, i_10_9_894_0, i_10_9_1029_0, i_10_9_1030_0,
    i_10_9_1031_0, i_10_9_1085_0, i_10_9_1235_0, i_10_9_1238_0,
    i_10_9_1250_0, i_10_9_1297_0, i_10_9_1298_0, i_10_9_1306_0,
    i_10_9_1631_0, i_10_9_1634_0, i_10_9_1685_0, i_10_9_1691_0,
    i_10_9_1822_0, i_10_9_1912_0, i_10_9_1981_0, i_10_9_1992_0,
    i_10_9_2027_0, i_10_9_2107_0, i_10_9_2197_0, i_10_9_2198_0,
    i_10_9_2201_0, i_10_9_2288_0, i_10_9_2334_0, i_10_9_2338_0,
    i_10_9_2352_0, i_10_9_2358_0, i_10_9_2379_0, i_10_9_2380_0,
    i_10_9_2452_0, i_10_9_2468_0, i_10_9_2470_0, i_10_9_2530_0,
    i_10_9_2567_0, i_10_9_2650_0, i_10_9_2656_0, i_10_9_2658_0,
    i_10_9_2711_0, i_10_9_2714_0, i_10_9_2728_0, i_10_9_2729_0,
    i_10_9_2740_0, i_10_9_2741_0, i_10_9_2783_0, i_10_9_2846_0,
    i_10_9_2918_0, i_10_9_2990_0, i_10_9_3046_0, i_10_9_3087_0,
    i_10_9_3313_0, i_10_9_3389_0, i_10_9_3390_0, i_10_9_3391_0,
    i_10_9_3395_0, i_10_9_3467_0, i_10_9_3502_0, i_10_9_3539_0,
    i_10_9_3557_0, i_10_9_3587_0, i_10_9_3612_0, i_10_9_3650_0,
    i_10_9_3652_0, i_10_9_3787_0, i_10_9_3838_0, i_10_9_3841_0,
    i_10_9_3847_0, i_10_9_3848_0, i_10_9_3910_0, i_10_9_3982_0,
    i_10_9_4027_0, i_10_9_4028_0, i_10_9_4113_0, i_10_9_4124_0,
    i_10_9_4172_0, i_10_9_4215_0, i_10_9_4277_0, i_10_9_4280_0,
    o_10_9_0_0  );
  input  i_10_9_47_0, i_10_9_146_0, i_10_9_171_0, i_10_9_176_0,
    i_10_9_191_0, i_10_9_224_0, i_10_9_247_0, i_10_9_279_0, i_10_9_281_0,
    i_10_9_287_0, i_10_9_315_0, i_10_9_317_0, i_10_9_443_0, i_10_9_459_0,
    i_10_9_462_0, i_10_9_463_0, i_10_9_464_0, i_10_9_509_0, i_10_9_635_0,
    i_10_9_821_0, i_10_9_891_0, i_10_9_894_0, i_10_9_1029_0, i_10_9_1030_0,
    i_10_9_1031_0, i_10_9_1085_0, i_10_9_1235_0, i_10_9_1238_0,
    i_10_9_1250_0, i_10_9_1297_0, i_10_9_1298_0, i_10_9_1306_0,
    i_10_9_1631_0, i_10_9_1634_0, i_10_9_1685_0, i_10_9_1691_0,
    i_10_9_1822_0, i_10_9_1912_0, i_10_9_1981_0, i_10_9_1992_0,
    i_10_9_2027_0, i_10_9_2107_0, i_10_9_2197_0, i_10_9_2198_0,
    i_10_9_2201_0, i_10_9_2288_0, i_10_9_2334_0, i_10_9_2338_0,
    i_10_9_2352_0, i_10_9_2358_0, i_10_9_2379_0, i_10_9_2380_0,
    i_10_9_2452_0, i_10_9_2468_0, i_10_9_2470_0, i_10_9_2530_0,
    i_10_9_2567_0, i_10_9_2650_0, i_10_9_2656_0, i_10_9_2658_0,
    i_10_9_2711_0, i_10_9_2714_0, i_10_9_2728_0, i_10_9_2729_0,
    i_10_9_2740_0, i_10_9_2741_0, i_10_9_2783_0, i_10_9_2846_0,
    i_10_9_2918_0, i_10_9_2990_0, i_10_9_3046_0, i_10_9_3087_0,
    i_10_9_3313_0, i_10_9_3389_0, i_10_9_3390_0, i_10_9_3391_0,
    i_10_9_3395_0, i_10_9_3467_0, i_10_9_3502_0, i_10_9_3539_0,
    i_10_9_3557_0, i_10_9_3587_0, i_10_9_3612_0, i_10_9_3650_0,
    i_10_9_3652_0, i_10_9_3787_0, i_10_9_3838_0, i_10_9_3841_0,
    i_10_9_3847_0, i_10_9_3848_0, i_10_9_3910_0, i_10_9_3982_0,
    i_10_9_4027_0, i_10_9_4028_0, i_10_9_4113_0, i_10_9_4124_0,
    i_10_9_4172_0, i_10_9_4215_0, i_10_9_4277_0, i_10_9_4280_0;
  output o_10_9_0_0;
  assign o_10_9_0_0 = 0;
endmodule



// Benchmark "kernel_10_10" written by ABC on Sun Jul 19 10:21:12 2020

module kernel_10_10 ( 
    i_10_10_283_0, i_10_10_285_0, i_10_10_319_0, i_10_10_426_0,
    i_10_10_435_0, i_10_10_507_0, i_10_10_622_0, i_10_10_636_0,
    i_10_10_891_0, i_10_10_897_0, i_10_10_949_0, i_10_10_950_0,
    i_10_10_1027_0, i_10_10_1029_0, i_10_10_1057_0, i_10_10_1117_0,
    i_10_10_1118_0, i_10_10_1122_0, i_10_10_1236_0, i_10_10_1243_0,
    i_10_10_1246_0, i_10_10_1247_0, i_10_10_1354_0, i_10_10_1396_0,
    i_10_10_1542_0, i_10_10_1575_0, i_10_10_1618_0, i_10_10_1648_0,
    i_10_10_1649_0, i_10_10_1691_0, i_10_10_1910_0, i_10_10_1945_0,
    i_10_10_1946_0, i_10_10_1959_0, i_10_10_1989_0, i_10_10_1992_0,
    i_10_10_2380_0, i_10_10_2454_0, i_10_10_2460_0, i_10_10_2511_0,
    i_10_10_2556_0, i_10_10_2557_0, i_10_10_2568_0, i_10_10_2608_0,
    i_10_10_2630_0, i_10_10_2631_0, i_10_10_2646_0, i_10_10_2657_0,
    i_10_10_2658_0, i_10_10_2659_0, i_10_10_2660_0, i_10_10_2710_0,
    i_10_10_2720_0, i_10_10_2727_0, i_10_10_2729_0, i_10_10_2829_0,
    i_10_10_2867_0, i_10_10_2881_0, i_10_10_2921_0, i_10_10_2923_0,
    i_10_10_3042_0, i_10_10_3045_0, i_10_10_3046_0, i_10_10_3072_0,
    i_10_10_3161_0, i_10_10_3229_0, i_10_10_3267_0, i_10_10_3269_0,
    i_10_10_3300_0, i_10_10_3336_0, i_10_10_3386_0, i_10_10_3440_0,
    i_10_10_3540_0, i_10_10_3549_0, i_10_10_3550_0, i_10_10_3551_0,
    i_10_10_3557_0, i_10_10_3620_0, i_10_10_3782_0, i_10_10_3848_0,
    i_10_10_3852_0, i_10_10_3981_0, i_10_10_4025_0, i_10_10_4026_0,
    i_10_10_4027_0, i_10_10_4118_0, i_10_10_4119_0, i_10_10_4125_0,
    i_10_10_4149_0, i_10_10_4151_0, i_10_10_4167_0, i_10_10_4191_0,
    i_10_10_4212_0, i_10_10_4213_0, i_10_10_4214_0, i_10_10_4290_0,
    i_10_10_4317_0, i_10_10_4565_0, i_10_10_4583_0, i_10_10_4584_0,
    o_10_10_0_0  );
  input  i_10_10_283_0, i_10_10_285_0, i_10_10_319_0, i_10_10_426_0,
    i_10_10_435_0, i_10_10_507_0, i_10_10_622_0, i_10_10_636_0,
    i_10_10_891_0, i_10_10_897_0, i_10_10_949_0, i_10_10_950_0,
    i_10_10_1027_0, i_10_10_1029_0, i_10_10_1057_0, i_10_10_1117_0,
    i_10_10_1118_0, i_10_10_1122_0, i_10_10_1236_0, i_10_10_1243_0,
    i_10_10_1246_0, i_10_10_1247_0, i_10_10_1354_0, i_10_10_1396_0,
    i_10_10_1542_0, i_10_10_1575_0, i_10_10_1618_0, i_10_10_1648_0,
    i_10_10_1649_0, i_10_10_1691_0, i_10_10_1910_0, i_10_10_1945_0,
    i_10_10_1946_0, i_10_10_1959_0, i_10_10_1989_0, i_10_10_1992_0,
    i_10_10_2380_0, i_10_10_2454_0, i_10_10_2460_0, i_10_10_2511_0,
    i_10_10_2556_0, i_10_10_2557_0, i_10_10_2568_0, i_10_10_2608_0,
    i_10_10_2630_0, i_10_10_2631_0, i_10_10_2646_0, i_10_10_2657_0,
    i_10_10_2658_0, i_10_10_2659_0, i_10_10_2660_0, i_10_10_2710_0,
    i_10_10_2720_0, i_10_10_2727_0, i_10_10_2729_0, i_10_10_2829_0,
    i_10_10_2867_0, i_10_10_2881_0, i_10_10_2921_0, i_10_10_2923_0,
    i_10_10_3042_0, i_10_10_3045_0, i_10_10_3046_0, i_10_10_3072_0,
    i_10_10_3161_0, i_10_10_3229_0, i_10_10_3267_0, i_10_10_3269_0,
    i_10_10_3300_0, i_10_10_3336_0, i_10_10_3386_0, i_10_10_3440_0,
    i_10_10_3540_0, i_10_10_3549_0, i_10_10_3550_0, i_10_10_3551_0,
    i_10_10_3557_0, i_10_10_3620_0, i_10_10_3782_0, i_10_10_3848_0,
    i_10_10_3852_0, i_10_10_3981_0, i_10_10_4025_0, i_10_10_4026_0,
    i_10_10_4027_0, i_10_10_4118_0, i_10_10_4119_0, i_10_10_4125_0,
    i_10_10_4149_0, i_10_10_4151_0, i_10_10_4167_0, i_10_10_4191_0,
    i_10_10_4212_0, i_10_10_4213_0, i_10_10_4214_0, i_10_10_4290_0,
    i_10_10_4317_0, i_10_10_4565_0, i_10_10_4583_0, i_10_10_4584_0;
  output o_10_10_0_0;
  assign o_10_10_0_0 = 0;
endmodule



// Benchmark "kernel_10_11" written by ABC on Sun Jul 19 10:21:13 2020

module kernel_10_11 ( 
    i_10_11_89_0, i_10_11_172_0, i_10_11_174_0, i_10_11_319_0,
    i_10_11_322_0, i_10_11_391_0, i_10_11_443_0, i_10_11_460_0,
    i_10_11_562_0, i_10_11_753_0, i_10_11_960_0, i_10_11_1048_0,
    i_10_11_1049_0, i_10_11_1088_0, i_10_11_1168_0, i_10_11_1240_0,
    i_10_11_1432_0, i_10_11_1435_0, i_10_11_1439_0, i_10_11_1545_0,
    i_10_11_1582_0, i_10_11_1583_0, i_10_11_1627_0, i_10_11_1650_0,
    i_10_11_1651_0, i_10_11_1686_0, i_10_11_1687_0, i_10_11_1689_0,
    i_10_11_1690_0, i_10_11_1691_0, i_10_11_1816_0, i_10_11_2023_0,
    i_10_11_2029_0, i_10_11_2201_0, i_10_11_2203_0, i_10_11_2353_0,
    i_10_11_2355_0, i_10_11_2356_0, i_10_11_2357_0, i_10_11_2359_0,
    i_10_11_2453_0, i_10_11_2463_0, i_10_11_2468_0, i_10_11_2471_0,
    i_10_11_2506_0, i_10_11_2542_0, i_10_11_2661_0, i_10_11_2662_0,
    i_10_11_2679_0, i_10_11_2707_0, i_10_11_2720_0, i_10_11_2733_0,
    i_10_11_2735_0, i_10_11_2784_0, i_10_11_2785_0, i_10_11_2789_0,
    i_10_11_2824_0, i_10_11_2966_0, i_10_11_3046_0, i_10_11_3070_0,
    i_10_11_3075_0, i_10_11_3238_0, i_10_11_3279_0, i_10_11_3281_0,
    i_10_11_3316_0, i_10_11_3389_0, i_10_11_3392_0, i_10_11_3431_0,
    i_10_11_3469_0, i_10_11_3525_0, i_10_11_3541_0, i_10_11_3556_0,
    i_10_11_3609_0, i_10_11_3683_0, i_10_11_3723_0, i_10_11_3724_0,
    i_10_11_3725_0, i_10_11_3727_0, i_10_11_3728_0, i_10_11_3780_0,
    i_10_11_3838_0, i_10_11_3844_0, i_10_11_3846_0, i_10_11_3847_0,
    i_10_11_3848_0, i_10_11_3946_0, i_10_11_4119_0, i_10_11_4121_0,
    i_10_11_4126_0, i_10_11_4128_0, i_10_11_4129_0, i_10_11_4207_0,
    i_10_11_4281_0, i_10_11_4282_0, i_10_11_4283_0, i_10_11_4291_0,
    i_10_11_4563_0, i_10_11_4566_0, i_10_11_4567_0, i_10_11_4583_0,
    o_10_11_0_0  );
  input  i_10_11_89_0, i_10_11_172_0, i_10_11_174_0, i_10_11_319_0,
    i_10_11_322_0, i_10_11_391_0, i_10_11_443_0, i_10_11_460_0,
    i_10_11_562_0, i_10_11_753_0, i_10_11_960_0, i_10_11_1048_0,
    i_10_11_1049_0, i_10_11_1088_0, i_10_11_1168_0, i_10_11_1240_0,
    i_10_11_1432_0, i_10_11_1435_0, i_10_11_1439_0, i_10_11_1545_0,
    i_10_11_1582_0, i_10_11_1583_0, i_10_11_1627_0, i_10_11_1650_0,
    i_10_11_1651_0, i_10_11_1686_0, i_10_11_1687_0, i_10_11_1689_0,
    i_10_11_1690_0, i_10_11_1691_0, i_10_11_1816_0, i_10_11_2023_0,
    i_10_11_2029_0, i_10_11_2201_0, i_10_11_2203_0, i_10_11_2353_0,
    i_10_11_2355_0, i_10_11_2356_0, i_10_11_2357_0, i_10_11_2359_0,
    i_10_11_2453_0, i_10_11_2463_0, i_10_11_2468_0, i_10_11_2471_0,
    i_10_11_2506_0, i_10_11_2542_0, i_10_11_2661_0, i_10_11_2662_0,
    i_10_11_2679_0, i_10_11_2707_0, i_10_11_2720_0, i_10_11_2733_0,
    i_10_11_2735_0, i_10_11_2784_0, i_10_11_2785_0, i_10_11_2789_0,
    i_10_11_2824_0, i_10_11_2966_0, i_10_11_3046_0, i_10_11_3070_0,
    i_10_11_3075_0, i_10_11_3238_0, i_10_11_3279_0, i_10_11_3281_0,
    i_10_11_3316_0, i_10_11_3389_0, i_10_11_3392_0, i_10_11_3431_0,
    i_10_11_3469_0, i_10_11_3525_0, i_10_11_3541_0, i_10_11_3556_0,
    i_10_11_3609_0, i_10_11_3683_0, i_10_11_3723_0, i_10_11_3724_0,
    i_10_11_3725_0, i_10_11_3727_0, i_10_11_3728_0, i_10_11_3780_0,
    i_10_11_3838_0, i_10_11_3844_0, i_10_11_3846_0, i_10_11_3847_0,
    i_10_11_3848_0, i_10_11_3946_0, i_10_11_4119_0, i_10_11_4121_0,
    i_10_11_4126_0, i_10_11_4128_0, i_10_11_4129_0, i_10_11_4207_0,
    i_10_11_4281_0, i_10_11_4282_0, i_10_11_4283_0, i_10_11_4291_0,
    i_10_11_4563_0, i_10_11_4566_0, i_10_11_4567_0, i_10_11_4583_0;
  output o_10_11_0_0;
  assign o_10_11_0_0 = 0;
endmodule



// Benchmark "kernel_10_12" written by ABC on Sun Jul 19 10:21:14 2020

module kernel_10_12 ( 
    i_10_12_44_0, i_10_12_147_0, i_10_12_151_0, i_10_12_177_0,
    i_10_12_430_0, i_10_12_448_0, i_10_12_518_0, i_10_12_521_0,
    i_10_12_637_0, i_10_12_714_0, i_10_12_717_0, i_10_12_735_0,
    i_10_12_798_0, i_10_12_832_0, i_10_12_903_0, i_10_12_931_0,
    i_10_12_967_0, i_10_12_970_0, i_10_12_1087_0, i_10_12_1127_0,
    i_10_12_1165_0, i_10_12_1233_0, i_10_12_1273_0, i_10_12_1306_0,
    i_10_12_1307_0, i_10_12_1310_0, i_10_12_1535_0, i_10_12_1537_0,
    i_10_12_1580_0, i_10_12_1637_0, i_10_12_1641_0, i_10_12_1709_0,
    i_10_12_1768_0, i_10_12_1795_0, i_10_12_1820_0, i_10_12_1874_0,
    i_10_12_1922_0, i_10_12_2001_0, i_10_12_2004_0, i_10_12_2028_0,
    i_10_12_2032_0, i_10_12_2186_0, i_10_12_2212_0, i_10_12_2309_0,
    i_10_12_2310_0, i_10_12_2311_0, i_10_12_2353_0, i_10_12_2354_0,
    i_10_12_2356_0, i_10_12_2389_0, i_10_12_2390_0, i_10_12_2451_0,
    i_10_12_2461_0, i_10_12_2472_0, i_10_12_2518_0, i_10_12_2631_0,
    i_10_12_2678_0, i_10_12_2680_0, i_10_12_2705_0, i_10_12_2914_0,
    i_10_12_2919_0, i_10_12_2983_0, i_10_12_2987_0, i_10_12_3014_0,
    i_10_12_3200_0, i_10_12_3234_0, i_10_12_3235_0, i_10_12_3279_0,
    i_10_12_3280_0, i_10_12_3319_0, i_10_12_3391_0, i_10_12_3470_0,
    i_10_12_3472_0, i_10_12_3473_0, i_10_12_3495_0, i_10_12_3496_0,
    i_10_12_3522_0, i_10_12_3525_0, i_10_12_3540_0, i_10_12_3541_0,
    i_10_12_3584_0, i_10_12_3588_0, i_10_12_3650_0, i_10_12_3776_0,
    i_10_12_3788_0, i_10_12_3823_0, i_10_12_3854_0, i_10_12_4013_0,
    i_10_12_4028_0, i_10_12_4051_0, i_10_12_4054_0, i_10_12_4117_0,
    i_10_12_4118_0, i_10_12_4229_0, i_10_12_4269_0, i_10_12_4282_0,
    i_10_12_4287_0, i_10_12_4291_0, i_10_12_4435_0, i_10_12_4588_0,
    o_10_12_0_0  );
  input  i_10_12_44_0, i_10_12_147_0, i_10_12_151_0, i_10_12_177_0,
    i_10_12_430_0, i_10_12_448_0, i_10_12_518_0, i_10_12_521_0,
    i_10_12_637_0, i_10_12_714_0, i_10_12_717_0, i_10_12_735_0,
    i_10_12_798_0, i_10_12_832_0, i_10_12_903_0, i_10_12_931_0,
    i_10_12_967_0, i_10_12_970_0, i_10_12_1087_0, i_10_12_1127_0,
    i_10_12_1165_0, i_10_12_1233_0, i_10_12_1273_0, i_10_12_1306_0,
    i_10_12_1307_0, i_10_12_1310_0, i_10_12_1535_0, i_10_12_1537_0,
    i_10_12_1580_0, i_10_12_1637_0, i_10_12_1641_0, i_10_12_1709_0,
    i_10_12_1768_0, i_10_12_1795_0, i_10_12_1820_0, i_10_12_1874_0,
    i_10_12_1922_0, i_10_12_2001_0, i_10_12_2004_0, i_10_12_2028_0,
    i_10_12_2032_0, i_10_12_2186_0, i_10_12_2212_0, i_10_12_2309_0,
    i_10_12_2310_0, i_10_12_2311_0, i_10_12_2353_0, i_10_12_2354_0,
    i_10_12_2356_0, i_10_12_2389_0, i_10_12_2390_0, i_10_12_2451_0,
    i_10_12_2461_0, i_10_12_2472_0, i_10_12_2518_0, i_10_12_2631_0,
    i_10_12_2678_0, i_10_12_2680_0, i_10_12_2705_0, i_10_12_2914_0,
    i_10_12_2919_0, i_10_12_2983_0, i_10_12_2987_0, i_10_12_3014_0,
    i_10_12_3200_0, i_10_12_3234_0, i_10_12_3235_0, i_10_12_3279_0,
    i_10_12_3280_0, i_10_12_3319_0, i_10_12_3391_0, i_10_12_3470_0,
    i_10_12_3472_0, i_10_12_3473_0, i_10_12_3495_0, i_10_12_3496_0,
    i_10_12_3522_0, i_10_12_3525_0, i_10_12_3540_0, i_10_12_3541_0,
    i_10_12_3584_0, i_10_12_3588_0, i_10_12_3650_0, i_10_12_3776_0,
    i_10_12_3788_0, i_10_12_3823_0, i_10_12_3854_0, i_10_12_4013_0,
    i_10_12_4028_0, i_10_12_4051_0, i_10_12_4054_0, i_10_12_4117_0,
    i_10_12_4118_0, i_10_12_4229_0, i_10_12_4269_0, i_10_12_4282_0,
    i_10_12_4287_0, i_10_12_4291_0, i_10_12_4435_0, i_10_12_4588_0;
  output o_10_12_0_0;
  assign o_10_12_0_0 = 0;
endmodule



// Benchmark "kernel_10_13" written by ABC on Sun Jul 19 10:21:15 2020

module kernel_10_13 ( 
    i_10_13_223_0, i_10_13_276_0, i_10_13_287_0, i_10_13_318_0,
    i_10_13_319_0, i_10_13_322_0, i_10_13_324_0, i_10_13_411_0,
    i_10_13_412_0, i_10_13_424_0, i_10_13_430_0, i_10_13_431_0,
    i_10_13_432_0, i_10_13_435_0, i_10_13_447_0, i_10_13_465_0,
    i_10_13_798_0, i_10_13_800_0, i_10_13_1249_0, i_10_13_1363_0,
    i_10_13_1365_0, i_10_13_1431_0, i_10_13_1437_0, i_10_13_1439_0,
    i_10_13_1546_0, i_10_13_1579_0, i_10_13_1581_0, i_10_13_1582_0,
    i_10_13_1626_0, i_10_13_1627_0, i_10_13_1653_0, i_10_13_1686_0,
    i_10_13_1687_0, i_10_13_1688_0, i_10_13_1724_0, i_10_13_1821_0,
    i_10_13_1822_0, i_10_13_1823_0, i_10_13_1911_0, i_10_13_1912_0,
    i_10_13_1995_0, i_10_13_1996_0, i_10_13_2005_0, i_10_13_2199_0,
    i_10_13_2452_0, i_10_13_2454_0, i_10_13_2466_0, i_10_13_2572_0,
    i_10_13_2604_0, i_10_13_2631_0, i_10_13_2632_0, i_10_13_2634_0,
    i_10_13_2635_0, i_10_13_2636_0, i_10_13_2705_0, i_10_13_2713_0,
    i_10_13_2722_0, i_10_13_2723_0, i_10_13_2730_0, i_10_13_2733_0,
    i_10_13_2734_0, i_10_13_2781_0, i_10_13_2826_0, i_10_13_2827_0,
    i_10_13_2828_0, i_10_13_2829_0, i_10_13_2830_0, i_10_13_2880_0,
    i_10_13_2883_0, i_10_13_2884_0, i_10_13_2885_0, i_10_13_3045_0,
    i_10_13_3070_0, i_10_13_3087_0, i_10_13_3151_0, i_10_13_3202_0,
    i_10_13_3268_0, i_10_13_3321_0, i_10_13_3387_0, i_10_13_3388_0,
    i_10_13_3543_0, i_10_13_3582_0, i_10_13_3613_0, i_10_13_3614_0,
    i_10_13_3616_0, i_10_13_3836_0, i_10_13_3837_0, i_10_13_3859_0,
    i_10_13_3912_0, i_10_13_3913_0, i_10_13_3978_0, i_10_13_3991_0,
    i_10_13_4057_0, i_10_13_4128_0, i_10_13_4129_0, i_10_13_4175_0,
    i_10_13_4281_0, i_10_13_4282_0, i_10_13_4283_0, i_10_13_4569_0,
    o_10_13_0_0  );
  input  i_10_13_223_0, i_10_13_276_0, i_10_13_287_0, i_10_13_318_0,
    i_10_13_319_0, i_10_13_322_0, i_10_13_324_0, i_10_13_411_0,
    i_10_13_412_0, i_10_13_424_0, i_10_13_430_0, i_10_13_431_0,
    i_10_13_432_0, i_10_13_435_0, i_10_13_447_0, i_10_13_465_0,
    i_10_13_798_0, i_10_13_800_0, i_10_13_1249_0, i_10_13_1363_0,
    i_10_13_1365_0, i_10_13_1431_0, i_10_13_1437_0, i_10_13_1439_0,
    i_10_13_1546_0, i_10_13_1579_0, i_10_13_1581_0, i_10_13_1582_0,
    i_10_13_1626_0, i_10_13_1627_0, i_10_13_1653_0, i_10_13_1686_0,
    i_10_13_1687_0, i_10_13_1688_0, i_10_13_1724_0, i_10_13_1821_0,
    i_10_13_1822_0, i_10_13_1823_0, i_10_13_1911_0, i_10_13_1912_0,
    i_10_13_1995_0, i_10_13_1996_0, i_10_13_2005_0, i_10_13_2199_0,
    i_10_13_2452_0, i_10_13_2454_0, i_10_13_2466_0, i_10_13_2572_0,
    i_10_13_2604_0, i_10_13_2631_0, i_10_13_2632_0, i_10_13_2634_0,
    i_10_13_2635_0, i_10_13_2636_0, i_10_13_2705_0, i_10_13_2713_0,
    i_10_13_2722_0, i_10_13_2723_0, i_10_13_2730_0, i_10_13_2733_0,
    i_10_13_2734_0, i_10_13_2781_0, i_10_13_2826_0, i_10_13_2827_0,
    i_10_13_2828_0, i_10_13_2829_0, i_10_13_2830_0, i_10_13_2880_0,
    i_10_13_2883_0, i_10_13_2884_0, i_10_13_2885_0, i_10_13_3045_0,
    i_10_13_3070_0, i_10_13_3087_0, i_10_13_3151_0, i_10_13_3202_0,
    i_10_13_3268_0, i_10_13_3321_0, i_10_13_3387_0, i_10_13_3388_0,
    i_10_13_3543_0, i_10_13_3582_0, i_10_13_3613_0, i_10_13_3614_0,
    i_10_13_3616_0, i_10_13_3836_0, i_10_13_3837_0, i_10_13_3859_0,
    i_10_13_3912_0, i_10_13_3913_0, i_10_13_3978_0, i_10_13_3991_0,
    i_10_13_4057_0, i_10_13_4128_0, i_10_13_4129_0, i_10_13_4175_0,
    i_10_13_4281_0, i_10_13_4282_0, i_10_13_4283_0, i_10_13_4569_0;
  output o_10_13_0_0;
  assign o_10_13_0_0 = ~((~i_10_13_2713_0 & ((~i_10_13_432_0 & ((~i_10_13_319_0 & i_10_13_1653_0 & ~i_10_13_2466_0 & i_10_13_3978_0) | (~i_10_13_1822_0 & ~i_10_13_2723_0 & ~i_10_13_3070_0 & ~i_10_13_3268_0 & ~i_10_13_3913_0 & ~i_10_13_3978_0 & ~i_10_13_4129_0 & ~i_10_13_4281_0))) | (~i_10_13_1431_0 & ~i_10_13_1439_0 & ~i_10_13_2828_0 & ~i_10_13_3268_0 & ~i_10_13_3837_0 & ~i_10_13_3978_0 & ~i_10_13_3991_0 & ~i_10_13_4281_0))) | (~i_10_13_319_0 & ((~i_10_13_318_0 & ~i_10_13_1821_0 & i_10_13_3837_0) | (~i_10_13_322_0 & ~i_10_13_411_0 & ~i_10_13_424_0 & ~i_10_13_800_0 & i_10_13_1653_0 & ~i_10_13_2734_0 & ~i_10_13_3045_0 & ~i_10_13_3087_0 & ~i_10_13_4282_0))) | (~i_10_13_322_0 & ((~i_10_13_424_0 & ~i_10_13_3268_0 & ~i_10_13_3582_0 & ~i_10_13_3614_0 & ~i_10_13_3837_0) | (~i_10_13_1823_0 & i_10_13_2631_0 & ~i_10_13_2734_0 & ~i_10_13_2884_0 & ~i_10_13_3070_0 & ~i_10_13_4569_0))) | (~i_10_13_1437_0 & ((~i_10_13_1626_0 & i_10_13_2829_0 & i_10_13_2830_0 & ~i_10_13_3912_0 & ~i_10_13_4128_0 & ~i_10_13_4175_0) | (~i_10_13_2452_0 & ~i_10_13_2826_0 & ~i_10_13_2828_0 & ~i_10_13_3388_0 & i_10_13_3616_0 & ~i_10_13_4281_0 & ~i_10_13_4282_0))) | (~i_10_13_4282_0 & ((~i_10_13_318_0 & ~i_10_13_1686_0 & ~i_10_13_2781_0 & ((~i_10_13_1688_0 & ~i_10_13_1912_0 & ~i_10_13_2452_0 & ~i_10_13_2454_0 & ~i_10_13_2884_0 & ~i_10_13_3268_0 & ~i_10_13_4128_0) | (~i_10_13_1431_0 & ~i_10_13_1579_0 & ~i_10_13_1626_0 & ~i_10_13_2466_0 & ~i_10_13_2885_0 & ~i_10_13_3978_0 & ~i_10_13_4283_0))) | (~i_10_13_3070_0 & (i_10_13_798_0 | (~i_10_13_424_0 & ~i_10_13_2005_0 & i_10_13_2632_0 & ~i_10_13_4129_0))))) | (~i_10_13_1822_0 & ~i_10_13_4175_0 & ((~i_10_13_1431_0 & i_10_13_2632_0 & ~i_10_13_3087_0 & ~i_10_13_3613_0) | (~i_10_13_435_0 & ~i_10_13_2604_0 & ~i_10_13_3837_0))) | (~i_10_13_2199_0 & ((~i_10_13_1582_0 & ~i_10_13_2634_0 & i_10_13_3616_0 & ~i_10_13_3978_0) | (~i_10_13_1431_0 & ~i_10_13_2883_0 & ~i_10_13_3070_0 & ~i_10_13_3582_0 & ~i_10_13_3991_0 & ~i_10_13_4283_0))) | (~i_10_13_1431_0 & ((~i_10_13_1579_0 & ~i_10_13_1823_0 & ~i_10_13_2883_0 & ~i_10_13_2884_0 & ~i_10_13_3582_0) | (i_10_13_3202_0 & ~i_10_13_3543_0 & ~i_10_13_4129_0))) | (~i_10_13_1579_0 & ((~i_10_13_318_0 & i_10_13_1687_0 & i_10_13_2466_0 & ~i_10_13_2722_0 & ~i_10_13_3388_0 & i_10_13_3582_0) | (~i_10_13_1687_0 & ~i_10_13_2883_0 & ~i_10_13_2884_0 & i_10_13_3045_0 & ~i_10_13_3087_0 & ~i_10_13_3614_0))) | (~i_10_13_1582_0 & ~i_10_13_3582_0 & ((~i_10_13_2452_0 & ~i_10_13_2466_0 & ~i_10_13_2883_0 & ~i_10_13_3070_0 & ~i_10_13_3836_0) | (i_10_13_2705_0 & ~i_10_13_3837_0))) | (i_10_13_2723_0 & ((i_10_13_1911_0 & ~i_10_13_2466_0) | (i_10_13_2713_0 & ~i_10_13_3837_0))) | (~i_10_13_4281_0 & ((i_10_13_2827_0 & ~i_10_13_2880_0 & ~i_10_13_3268_0 & ~i_10_13_3859_0) | (~i_10_13_1627_0 & ~i_10_13_3543_0 & i_10_13_3859_0 & ~i_10_13_3978_0))) | (~i_10_13_3087_0 & ~i_10_13_3614_0 & i_10_13_1912_0 & ~i_10_13_2452_0));
endmodule



// Benchmark "kernel_10_14" written by ABC on Sun Jul 19 10:21:16 2020

module kernel_10_14 ( 
    i_10_14_183_0, i_10_14_195_0, i_10_14_324_0, i_10_14_394_0,
    i_10_14_409_0, i_10_14_430_0, i_10_14_445_0, i_10_14_460_0,
    i_10_14_463_0, i_10_14_511_0, i_10_14_516_0, i_10_14_520_0,
    i_10_14_577_0, i_10_14_697_0, i_10_14_732_0, i_10_14_733_0,
    i_10_14_798_0, i_10_14_864_0, i_10_14_867_0, i_10_14_969_0,
    i_10_14_1098_0, i_10_14_1119_0, i_10_14_1120_0, i_10_14_1168_0,
    i_10_14_1239_0, i_10_14_1246_0, i_10_14_1551_0, i_10_14_1581_0,
    i_10_14_1620_0, i_10_14_1693_0, i_10_14_1696_0, i_10_14_1715_0,
    i_10_14_1756_0, i_10_14_1767_0, i_10_14_1789_0, i_10_14_1885_0,
    i_10_14_1908_0, i_10_14_1912_0, i_10_14_1948_0, i_10_14_1950_0,
    i_10_14_2085_0, i_10_14_2155_0, i_10_14_2334_0, i_10_14_2352_0,
    i_10_14_2442_0, i_10_14_2452_0, i_10_14_2453_0, i_10_14_2463_0,
    i_10_14_2481_0, i_10_14_2574_0, i_10_14_2577_0, i_10_14_2631_0,
    i_10_14_2634_0, i_10_14_2676_0, i_10_14_2680_0, i_10_14_2711_0,
    i_10_14_2830_0, i_10_14_2866_0, i_10_14_2868_0, i_10_14_2919_0,
    i_10_14_2922_0, i_10_14_2983_0, i_10_14_2984_0, i_10_14_3036_0,
    i_10_14_3047_0, i_10_14_3049_0, i_10_14_3198_0, i_10_14_3199_0,
    i_10_14_3277_0, i_10_14_3298_0, i_10_14_3312_0, i_10_14_3407_0,
    i_10_14_3540_0, i_10_14_3541_0, i_10_14_3609_0, i_10_14_3686_0,
    i_10_14_3688_0, i_10_14_3720_0, i_10_14_3724_0, i_10_14_3795_0,
    i_10_14_3921_0, i_10_14_3931_0, i_10_14_3964_0, i_10_14_3968_0,
    i_10_14_3981_0, i_10_14_3982_0, i_10_14_3984_0, i_10_14_3985_0,
    i_10_14_4155_0, i_10_14_4191_0, i_10_14_4192_0, i_10_14_4207_0,
    i_10_14_4269_0, i_10_14_4271_0, i_10_14_4273_0, i_10_14_4278_0,
    i_10_14_4279_0, i_10_14_4290_0, i_10_14_4291_0, i_10_14_4515_0,
    o_10_14_0_0  );
  input  i_10_14_183_0, i_10_14_195_0, i_10_14_324_0, i_10_14_394_0,
    i_10_14_409_0, i_10_14_430_0, i_10_14_445_0, i_10_14_460_0,
    i_10_14_463_0, i_10_14_511_0, i_10_14_516_0, i_10_14_520_0,
    i_10_14_577_0, i_10_14_697_0, i_10_14_732_0, i_10_14_733_0,
    i_10_14_798_0, i_10_14_864_0, i_10_14_867_0, i_10_14_969_0,
    i_10_14_1098_0, i_10_14_1119_0, i_10_14_1120_0, i_10_14_1168_0,
    i_10_14_1239_0, i_10_14_1246_0, i_10_14_1551_0, i_10_14_1581_0,
    i_10_14_1620_0, i_10_14_1693_0, i_10_14_1696_0, i_10_14_1715_0,
    i_10_14_1756_0, i_10_14_1767_0, i_10_14_1789_0, i_10_14_1885_0,
    i_10_14_1908_0, i_10_14_1912_0, i_10_14_1948_0, i_10_14_1950_0,
    i_10_14_2085_0, i_10_14_2155_0, i_10_14_2334_0, i_10_14_2352_0,
    i_10_14_2442_0, i_10_14_2452_0, i_10_14_2453_0, i_10_14_2463_0,
    i_10_14_2481_0, i_10_14_2574_0, i_10_14_2577_0, i_10_14_2631_0,
    i_10_14_2634_0, i_10_14_2676_0, i_10_14_2680_0, i_10_14_2711_0,
    i_10_14_2830_0, i_10_14_2866_0, i_10_14_2868_0, i_10_14_2919_0,
    i_10_14_2922_0, i_10_14_2983_0, i_10_14_2984_0, i_10_14_3036_0,
    i_10_14_3047_0, i_10_14_3049_0, i_10_14_3198_0, i_10_14_3199_0,
    i_10_14_3277_0, i_10_14_3298_0, i_10_14_3312_0, i_10_14_3407_0,
    i_10_14_3540_0, i_10_14_3541_0, i_10_14_3609_0, i_10_14_3686_0,
    i_10_14_3688_0, i_10_14_3720_0, i_10_14_3724_0, i_10_14_3795_0,
    i_10_14_3921_0, i_10_14_3931_0, i_10_14_3964_0, i_10_14_3968_0,
    i_10_14_3981_0, i_10_14_3982_0, i_10_14_3984_0, i_10_14_3985_0,
    i_10_14_4155_0, i_10_14_4191_0, i_10_14_4192_0, i_10_14_4207_0,
    i_10_14_4269_0, i_10_14_4271_0, i_10_14_4273_0, i_10_14_4278_0,
    i_10_14_4279_0, i_10_14_4290_0, i_10_14_4291_0, i_10_14_4515_0;
  output o_10_14_0_0;
  assign o_10_14_0_0 = ~((~i_10_14_520_0 & ((~i_10_14_516_0 & ~i_10_14_2922_0 & ~i_10_14_3312_0 & ~i_10_14_3609_0 & i_10_14_4273_0) | (~i_10_14_394_0 & ~i_10_14_1912_0 & ~i_10_14_4273_0))) | (~i_10_14_394_0 & ((~i_10_14_2680_0 & ~i_10_14_3609_0 & ~i_10_14_4279_0) | (~i_10_14_3049_0 & ~i_10_14_3312_0 & i_10_14_4273_0 & i_10_14_4291_0))) | (~i_10_14_1908_0 & ((i_10_14_2453_0 & ~i_10_14_4269_0) | (~i_10_14_1620_0 & i_10_14_2631_0 & ~i_10_14_3047_0 & ~i_10_14_3199_0 & i_10_14_3981_0 & ~i_10_14_4271_0))) | (~i_10_14_1620_0 & (~i_10_14_3982_0 | (~i_10_14_2452_0 & ~i_10_14_2919_0 & ~i_10_14_3049_0 & ~i_10_14_3688_0))) | (~i_10_14_3277_0 & ((~i_10_14_969_0 & i_10_14_2676_0) | (~i_10_14_3981_0 & ~i_10_14_4278_0))) | (~i_10_14_4278_0 & ((i_10_14_2453_0 & ~i_10_14_2463_0) | (~i_10_14_3984_0 & ~i_10_14_4279_0))) | i_10_14_3686_0 | (~i_10_14_2334_0 & i_10_14_2983_0 & ~i_10_14_4279_0) | (~i_10_14_460_0 & ~i_10_14_2453_0 & ~i_10_14_3049_0 & ~i_10_14_3540_0 & ~i_10_14_3688_0) | (~i_10_14_1239_0 & ~i_10_14_3312_0 & ~i_10_14_3985_0) | (~i_10_14_2634_0 & i_10_14_3036_0 & ~i_10_14_4273_0));
endmodule



// Benchmark "kernel_10_15" written by ABC on Sun Jul 19 10:21:17 2020

module kernel_10_15 ( 
    i_10_15_51_0, i_10_15_148_0, i_10_15_283_0, i_10_15_295_0,
    i_10_15_322_0, i_10_15_436_0, i_10_15_445_0, i_10_15_448_0,
    i_10_15_449_0, i_10_15_463_0, i_10_15_467_0, i_10_15_562_0,
    i_10_15_896_0, i_10_15_899_0, i_10_15_907_0, i_10_15_997_0,
    i_10_15_1033_0, i_10_15_1034_0, i_10_15_1051_0, i_10_15_1234_0,
    i_10_15_1249_0, i_10_15_1250_0, i_10_15_1446_0, i_10_15_1447_0,
    i_10_15_1619_0, i_10_15_1636_0, i_10_15_1637_0, i_10_15_1652_0,
    i_10_15_1684_0, i_10_15_1686_0, i_10_15_1687_0, i_10_15_1688_0,
    i_10_15_1690_0, i_10_15_1691_0, i_10_15_1808_0, i_10_15_1819_0,
    i_10_15_1823_0, i_10_15_1826_0, i_10_15_1910_0, i_10_15_1913_0,
    i_10_15_1960_0, i_10_15_2015_0, i_10_15_2158_0, i_10_15_2231_0,
    i_10_15_2353_0, i_10_15_2354_0, i_10_15_2355_0, i_10_15_2357_0,
    i_10_15_2365_0, i_10_15_2448_0, i_10_15_2456_0, i_10_15_2481_0,
    i_10_15_2482_0, i_10_15_2528_0, i_10_15_2535_0, i_10_15_2540_0,
    i_10_15_2546_0, i_10_15_2571_0, i_10_15_2572_0, i_10_15_2608_0,
    i_10_15_2632_0, i_10_15_2636_0, i_10_15_2654_0, i_10_15_2659_0,
    i_10_15_2662_0, i_10_15_2689_0, i_10_15_2708_0, i_10_15_2788_0,
    i_10_15_2832_0, i_10_15_2833_0, i_10_15_3038_0, i_10_15_3076_0,
    i_10_15_3196_0, i_10_15_3199_0, i_10_15_3200_0, i_10_15_3272_0,
    i_10_15_3274_0, i_10_15_3275_0, i_10_15_3278_0, i_10_15_3356_0,
    i_10_15_3384_0, i_10_15_3391_0, i_10_15_3392_0, i_10_15_3463_0,
    i_10_15_3527_0, i_10_15_3544_0, i_10_15_3721_0, i_10_15_3733_0,
    i_10_15_3859_0, i_10_15_3894_0, i_10_15_3905_0, i_10_15_3985_0,
    i_10_15_3986_0, i_10_15_3992_0, i_10_15_4030_0, i_10_15_4031_0,
    i_10_15_4118_0, i_10_15_4121_0, i_10_15_4154_0, i_10_15_4570_0,
    o_10_15_0_0  );
  input  i_10_15_51_0, i_10_15_148_0, i_10_15_283_0, i_10_15_295_0,
    i_10_15_322_0, i_10_15_436_0, i_10_15_445_0, i_10_15_448_0,
    i_10_15_449_0, i_10_15_463_0, i_10_15_467_0, i_10_15_562_0,
    i_10_15_896_0, i_10_15_899_0, i_10_15_907_0, i_10_15_997_0,
    i_10_15_1033_0, i_10_15_1034_0, i_10_15_1051_0, i_10_15_1234_0,
    i_10_15_1249_0, i_10_15_1250_0, i_10_15_1446_0, i_10_15_1447_0,
    i_10_15_1619_0, i_10_15_1636_0, i_10_15_1637_0, i_10_15_1652_0,
    i_10_15_1684_0, i_10_15_1686_0, i_10_15_1687_0, i_10_15_1688_0,
    i_10_15_1690_0, i_10_15_1691_0, i_10_15_1808_0, i_10_15_1819_0,
    i_10_15_1823_0, i_10_15_1826_0, i_10_15_1910_0, i_10_15_1913_0,
    i_10_15_1960_0, i_10_15_2015_0, i_10_15_2158_0, i_10_15_2231_0,
    i_10_15_2353_0, i_10_15_2354_0, i_10_15_2355_0, i_10_15_2357_0,
    i_10_15_2365_0, i_10_15_2448_0, i_10_15_2456_0, i_10_15_2481_0,
    i_10_15_2482_0, i_10_15_2528_0, i_10_15_2535_0, i_10_15_2540_0,
    i_10_15_2546_0, i_10_15_2571_0, i_10_15_2572_0, i_10_15_2608_0,
    i_10_15_2632_0, i_10_15_2636_0, i_10_15_2654_0, i_10_15_2659_0,
    i_10_15_2662_0, i_10_15_2689_0, i_10_15_2708_0, i_10_15_2788_0,
    i_10_15_2832_0, i_10_15_2833_0, i_10_15_3038_0, i_10_15_3076_0,
    i_10_15_3196_0, i_10_15_3199_0, i_10_15_3200_0, i_10_15_3272_0,
    i_10_15_3274_0, i_10_15_3275_0, i_10_15_3278_0, i_10_15_3356_0,
    i_10_15_3384_0, i_10_15_3391_0, i_10_15_3392_0, i_10_15_3463_0,
    i_10_15_3527_0, i_10_15_3544_0, i_10_15_3721_0, i_10_15_3733_0,
    i_10_15_3859_0, i_10_15_3894_0, i_10_15_3905_0, i_10_15_3985_0,
    i_10_15_3986_0, i_10_15_3992_0, i_10_15_4030_0, i_10_15_4031_0,
    i_10_15_4118_0, i_10_15_4121_0, i_10_15_4154_0, i_10_15_4570_0;
  output o_10_15_0_0;
  assign o_10_15_0_0 = 0;
endmodule



// Benchmark "kernel_10_16" written by ABC on Sun Jul 19 10:21:18 2020

module kernel_10_16 ( 
    i_10_16_40_0, i_10_16_149_0, i_10_16_153_0, i_10_16_175_0,
    i_10_16_183_0, i_10_16_229_0, i_10_16_265_0, i_10_16_363_0,
    i_10_16_366_0, i_10_16_406_0, i_10_16_408_0, i_10_16_437_0,
    i_10_16_448_0, i_10_16_513_0, i_10_16_670_0, i_10_16_691_0,
    i_10_16_751_0, i_10_16_906_0, i_10_16_933_0, i_10_16_1029_0,
    i_10_16_1033_0, i_10_16_1038_0, i_10_16_1135_0, i_10_16_1137_0,
    i_10_16_1138_0, i_10_16_1139_0, i_10_16_1153_0, i_10_16_1157_0,
    i_10_16_1158_0, i_10_16_1164_0, i_10_16_1165_0, i_10_16_1218_0,
    i_10_16_1219_0, i_10_16_1238_0, i_10_16_1239_0, i_10_16_1264_0,
    i_10_16_1266_0, i_10_16_1267_0, i_10_16_1305_0, i_10_16_1308_0,
    i_10_16_1310_0, i_10_16_1311_0, i_10_16_1378_0, i_10_16_1399_0,
    i_10_16_1455_0, i_10_16_1552_0, i_10_16_1554_0, i_10_16_1632_0,
    i_10_16_1647_0, i_10_16_1815_0, i_10_16_1858_0, i_10_16_1872_0,
    i_10_16_1914_0, i_10_16_1948_0, i_10_16_1956_0, i_10_16_1998_0,
    i_10_16_2019_0, i_10_16_2020_0, i_10_16_2068_0, i_10_16_2391_0,
    i_10_16_2409_0, i_10_16_2505_0, i_10_16_2508_0, i_10_16_2568_0,
    i_10_16_2589_0, i_10_16_2605_0, i_10_16_2613_0, i_10_16_2634_0,
    i_10_16_2703_0, i_10_16_2704_0, i_10_16_2705_0, i_10_16_2706_0,
    i_10_16_2707_0, i_10_16_2713_0, i_10_16_2724_0, i_10_16_2725_0,
    i_10_16_2733_0, i_10_16_2985_0, i_10_16_2986_0, i_10_16_3234_0,
    i_10_16_3293_0, i_10_16_3397_0, i_10_16_3435_0, i_10_16_3455_0,
    i_10_16_3470_0, i_10_16_3498_0, i_10_16_3541_0, i_10_16_3667_0,
    i_10_16_3717_0, i_10_16_3720_0, i_10_16_3779_0, i_10_16_3789_0,
    i_10_16_3879_0, i_10_16_4116_0, i_10_16_4117_0, i_10_16_4120_0,
    i_10_16_4140_0, i_10_16_4278_0, i_10_16_4555_0, i_10_16_4570_0,
    o_10_16_0_0  );
  input  i_10_16_40_0, i_10_16_149_0, i_10_16_153_0, i_10_16_175_0,
    i_10_16_183_0, i_10_16_229_0, i_10_16_265_0, i_10_16_363_0,
    i_10_16_366_0, i_10_16_406_0, i_10_16_408_0, i_10_16_437_0,
    i_10_16_448_0, i_10_16_513_0, i_10_16_670_0, i_10_16_691_0,
    i_10_16_751_0, i_10_16_906_0, i_10_16_933_0, i_10_16_1029_0,
    i_10_16_1033_0, i_10_16_1038_0, i_10_16_1135_0, i_10_16_1137_0,
    i_10_16_1138_0, i_10_16_1139_0, i_10_16_1153_0, i_10_16_1157_0,
    i_10_16_1158_0, i_10_16_1164_0, i_10_16_1165_0, i_10_16_1218_0,
    i_10_16_1219_0, i_10_16_1238_0, i_10_16_1239_0, i_10_16_1264_0,
    i_10_16_1266_0, i_10_16_1267_0, i_10_16_1305_0, i_10_16_1308_0,
    i_10_16_1310_0, i_10_16_1311_0, i_10_16_1378_0, i_10_16_1399_0,
    i_10_16_1455_0, i_10_16_1552_0, i_10_16_1554_0, i_10_16_1632_0,
    i_10_16_1647_0, i_10_16_1815_0, i_10_16_1858_0, i_10_16_1872_0,
    i_10_16_1914_0, i_10_16_1948_0, i_10_16_1956_0, i_10_16_1998_0,
    i_10_16_2019_0, i_10_16_2020_0, i_10_16_2068_0, i_10_16_2391_0,
    i_10_16_2409_0, i_10_16_2505_0, i_10_16_2508_0, i_10_16_2568_0,
    i_10_16_2589_0, i_10_16_2605_0, i_10_16_2613_0, i_10_16_2634_0,
    i_10_16_2703_0, i_10_16_2704_0, i_10_16_2705_0, i_10_16_2706_0,
    i_10_16_2707_0, i_10_16_2713_0, i_10_16_2724_0, i_10_16_2725_0,
    i_10_16_2733_0, i_10_16_2985_0, i_10_16_2986_0, i_10_16_3234_0,
    i_10_16_3293_0, i_10_16_3397_0, i_10_16_3435_0, i_10_16_3455_0,
    i_10_16_3470_0, i_10_16_3498_0, i_10_16_3541_0, i_10_16_3667_0,
    i_10_16_3717_0, i_10_16_3720_0, i_10_16_3779_0, i_10_16_3789_0,
    i_10_16_3879_0, i_10_16_4116_0, i_10_16_4117_0, i_10_16_4120_0,
    i_10_16_4140_0, i_10_16_4278_0, i_10_16_4555_0, i_10_16_4570_0;
  output o_10_16_0_0;
  assign o_10_16_0_0 = 0;
endmodule



// Benchmark "kernel_10_17" written by ABC on Sun Jul 19 10:21:19 2020

module kernel_10_17 ( 
    i_10_17_37_0, i_10_17_49_0, i_10_17_68_0, i_10_17_128_0, i_10_17_155_0,
    i_10_17_244_0, i_10_17_282_0, i_10_17_286_0, i_10_17_406_0,
    i_10_17_407_0, i_10_17_438_0, i_10_17_441_0, i_10_17_443_0,
    i_10_17_463_0, i_10_17_464_0, i_10_17_824_0, i_10_17_959_0,
    i_10_17_994_0, i_10_17_1001_0, i_10_17_1109_0, i_10_17_1241_0,
    i_10_17_1248_0, i_10_17_1305_0, i_10_17_1306_0, i_10_17_1310_0,
    i_10_17_1313_0, i_10_17_1432_0, i_10_17_1579_0, i_10_17_1647_0,
    i_10_17_1648_0, i_10_17_1651_0, i_10_17_1684_0, i_10_17_1688_0,
    i_10_17_1795_0, i_10_17_1800_0, i_10_17_1913_0, i_10_17_1948_0,
    i_10_17_2196_0, i_10_17_2197_0, i_10_17_2234_0, i_10_17_2246_0,
    i_10_17_2352_0, i_10_17_2354_0, i_10_17_2407_0, i_10_17_2449_0,
    i_10_17_2455_0, i_10_17_2518_0, i_10_17_2534_0, i_10_17_2606_0,
    i_10_17_2628_0, i_10_17_2677_0, i_10_17_2706_0, i_10_17_2727_0,
    i_10_17_2730_0, i_10_17_2734_0, i_10_17_2832_0, i_10_17_2880_0,
    i_10_17_3040_0, i_10_17_3199_0, i_10_17_3232_0, i_10_17_3238_0,
    i_10_17_3271_0, i_10_17_3281_0, i_10_17_3384_0, i_10_17_3386_0,
    i_10_17_3387_0, i_10_17_3388_0, i_10_17_3389_0, i_10_17_3523_0,
    i_10_17_3611_0, i_10_17_3613_0, i_10_17_3614_0, i_10_17_3649_0,
    i_10_17_3650_0, i_10_17_3652_0, i_10_17_3684_0, i_10_17_3685_0,
    i_10_17_3781_0, i_10_17_3782_0, i_10_17_3784_0, i_10_17_3787_0,
    i_10_17_3788_0, i_10_17_3800_0, i_10_17_3834_0, i_10_17_3835_0,
    i_10_17_3844_0, i_10_17_3847_0, i_10_17_3856_0, i_10_17_3860_0,
    i_10_17_4027_0, i_10_17_4120_0, i_10_17_4123_0, i_10_17_4143_0,
    i_10_17_4170_0, i_10_17_4276_0, i_10_17_4285_0, i_10_17_4286_0,
    i_10_17_4288_0, i_10_17_4289_0, i_10_17_4372_0,
    o_10_17_0_0  );
  input  i_10_17_37_0, i_10_17_49_0, i_10_17_68_0, i_10_17_128_0,
    i_10_17_155_0, i_10_17_244_0, i_10_17_282_0, i_10_17_286_0,
    i_10_17_406_0, i_10_17_407_0, i_10_17_438_0, i_10_17_441_0,
    i_10_17_443_0, i_10_17_463_0, i_10_17_464_0, i_10_17_824_0,
    i_10_17_959_0, i_10_17_994_0, i_10_17_1001_0, i_10_17_1109_0,
    i_10_17_1241_0, i_10_17_1248_0, i_10_17_1305_0, i_10_17_1306_0,
    i_10_17_1310_0, i_10_17_1313_0, i_10_17_1432_0, i_10_17_1579_0,
    i_10_17_1647_0, i_10_17_1648_0, i_10_17_1651_0, i_10_17_1684_0,
    i_10_17_1688_0, i_10_17_1795_0, i_10_17_1800_0, i_10_17_1913_0,
    i_10_17_1948_0, i_10_17_2196_0, i_10_17_2197_0, i_10_17_2234_0,
    i_10_17_2246_0, i_10_17_2352_0, i_10_17_2354_0, i_10_17_2407_0,
    i_10_17_2449_0, i_10_17_2455_0, i_10_17_2518_0, i_10_17_2534_0,
    i_10_17_2606_0, i_10_17_2628_0, i_10_17_2677_0, i_10_17_2706_0,
    i_10_17_2727_0, i_10_17_2730_0, i_10_17_2734_0, i_10_17_2832_0,
    i_10_17_2880_0, i_10_17_3040_0, i_10_17_3199_0, i_10_17_3232_0,
    i_10_17_3238_0, i_10_17_3271_0, i_10_17_3281_0, i_10_17_3384_0,
    i_10_17_3386_0, i_10_17_3387_0, i_10_17_3388_0, i_10_17_3389_0,
    i_10_17_3523_0, i_10_17_3611_0, i_10_17_3613_0, i_10_17_3614_0,
    i_10_17_3649_0, i_10_17_3650_0, i_10_17_3652_0, i_10_17_3684_0,
    i_10_17_3685_0, i_10_17_3781_0, i_10_17_3782_0, i_10_17_3784_0,
    i_10_17_3787_0, i_10_17_3788_0, i_10_17_3800_0, i_10_17_3834_0,
    i_10_17_3835_0, i_10_17_3844_0, i_10_17_3847_0, i_10_17_3856_0,
    i_10_17_3860_0, i_10_17_4027_0, i_10_17_4120_0, i_10_17_4123_0,
    i_10_17_4143_0, i_10_17_4170_0, i_10_17_4276_0, i_10_17_4285_0,
    i_10_17_4286_0, i_10_17_4288_0, i_10_17_4289_0, i_10_17_4372_0;
  output o_10_17_0_0;
  assign o_10_17_0_0 = 0;
endmodule



// Benchmark "kernel_10_18" written by ABC on Sun Jul 19 10:21:20 2020

module kernel_10_18 ( 
    i_10_18_28_0, i_10_18_171_0, i_10_18_174_0, i_10_18_175_0,
    i_10_18_176_0, i_10_18_261_0, i_10_18_267_0, i_10_18_390_0,
    i_10_18_393_0, i_10_18_409_0, i_10_18_410_0, i_10_18_411_0,
    i_10_18_412_0, i_10_18_441_0, i_10_18_442_0, i_10_18_446_0,
    i_10_18_718_0, i_10_18_793_0, i_10_18_796_0, i_10_18_960_0,
    i_10_18_1003_0, i_10_18_1005_0, i_10_18_1006_0, i_10_18_1026_0,
    i_10_18_1028_0, i_10_18_1036_0, i_10_18_1238_0, i_10_18_1242_0,
    i_10_18_1312_0, i_10_18_1431_0, i_10_18_1432_0, i_10_18_1434_0,
    i_10_18_1440_0, i_10_18_1539_0, i_10_18_1554_0, i_10_18_1575_0,
    i_10_18_1651_0, i_10_18_1652_0, i_10_18_1655_0, i_10_18_1688_0,
    i_10_18_1691_0, i_10_18_1819_0, i_10_18_1822_0, i_10_18_1824_0,
    i_10_18_1825_0, i_10_18_1947_0, i_10_18_1950_0, i_10_18_2001_0,
    i_10_18_2178_0, i_10_18_2179_0, i_10_18_2184_0, i_10_18_2185_0,
    i_10_18_2186_0, i_10_18_2355_0, i_10_18_2358_0, i_10_18_2410_0,
    i_10_18_2460_0, i_10_18_2466_0, i_10_18_2469_0, i_10_18_2565_0,
    i_10_18_2567_0, i_10_18_2605_0, i_10_18_2656_0, i_10_18_2724_0,
    i_10_18_2725_0, i_10_18_2731_0, i_10_18_2732_0, i_10_18_2735_0,
    i_10_18_2832_0, i_10_18_2883_0, i_10_18_2923_0, i_10_18_2987_0,
    i_10_18_3036_0, i_10_18_3042_0, i_10_18_3045_0, i_10_18_3069_0,
    i_10_18_3070_0, i_10_18_3095_0, i_10_18_3198_0, i_10_18_3202_0,
    i_10_18_3276_0, i_10_18_3388_0, i_10_18_3391_0, i_10_18_3467_0,
    i_10_18_3471_0, i_10_18_3522_0, i_10_18_3523_0, i_10_18_3525_0,
    i_10_18_3610_0, i_10_18_3780_0, i_10_18_3783_0, i_10_18_3788_0,
    i_10_18_3834_0, i_10_18_3838_0, i_10_18_3841_0, i_10_18_3855_0,
    i_10_18_3856_0, i_10_18_3913_0, i_10_18_4291_0, i_10_18_4292_0,
    o_10_18_0_0  );
  input  i_10_18_28_0, i_10_18_171_0, i_10_18_174_0, i_10_18_175_0,
    i_10_18_176_0, i_10_18_261_0, i_10_18_267_0, i_10_18_390_0,
    i_10_18_393_0, i_10_18_409_0, i_10_18_410_0, i_10_18_411_0,
    i_10_18_412_0, i_10_18_441_0, i_10_18_442_0, i_10_18_446_0,
    i_10_18_718_0, i_10_18_793_0, i_10_18_796_0, i_10_18_960_0,
    i_10_18_1003_0, i_10_18_1005_0, i_10_18_1006_0, i_10_18_1026_0,
    i_10_18_1028_0, i_10_18_1036_0, i_10_18_1238_0, i_10_18_1242_0,
    i_10_18_1312_0, i_10_18_1431_0, i_10_18_1432_0, i_10_18_1434_0,
    i_10_18_1440_0, i_10_18_1539_0, i_10_18_1554_0, i_10_18_1575_0,
    i_10_18_1651_0, i_10_18_1652_0, i_10_18_1655_0, i_10_18_1688_0,
    i_10_18_1691_0, i_10_18_1819_0, i_10_18_1822_0, i_10_18_1824_0,
    i_10_18_1825_0, i_10_18_1947_0, i_10_18_1950_0, i_10_18_2001_0,
    i_10_18_2178_0, i_10_18_2179_0, i_10_18_2184_0, i_10_18_2185_0,
    i_10_18_2186_0, i_10_18_2355_0, i_10_18_2358_0, i_10_18_2410_0,
    i_10_18_2460_0, i_10_18_2466_0, i_10_18_2469_0, i_10_18_2565_0,
    i_10_18_2567_0, i_10_18_2605_0, i_10_18_2656_0, i_10_18_2724_0,
    i_10_18_2725_0, i_10_18_2731_0, i_10_18_2732_0, i_10_18_2735_0,
    i_10_18_2832_0, i_10_18_2883_0, i_10_18_2923_0, i_10_18_2987_0,
    i_10_18_3036_0, i_10_18_3042_0, i_10_18_3045_0, i_10_18_3069_0,
    i_10_18_3070_0, i_10_18_3095_0, i_10_18_3198_0, i_10_18_3202_0,
    i_10_18_3276_0, i_10_18_3388_0, i_10_18_3391_0, i_10_18_3467_0,
    i_10_18_3471_0, i_10_18_3522_0, i_10_18_3523_0, i_10_18_3525_0,
    i_10_18_3610_0, i_10_18_3780_0, i_10_18_3783_0, i_10_18_3788_0,
    i_10_18_3834_0, i_10_18_3838_0, i_10_18_3841_0, i_10_18_3855_0,
    i_10_18_3856_0, i_10_18_3913_0, i_10_18_4291_0, i_10_18_4292_0;
  output o_10_18_0_0;
  assign o_10_18_0_0 = ~((~i_10_18_1026_0 & ((~i_10_18_261_0 & ((~i_10_18_390_0 & ~i_10_18_796_0 & ~i_10_18_960_0 & ~i_10_18_1238_0 & ~i_10_18_1434_0 & ~i_10_18_2179_0 & ~i_10_18_2185_0 & ~i_10_18_2186_0 & ~i_10_18_2567_0 & ~i_10_18_3095_0 & ~i_10_18_3783_0) | (~i_10_18_1554_0 & ~i_10_18_1822_0 & i_10_18_2355_0 & i_10_18_2731_0 & ~i_10_18_3202_0 & ~i_10_18_3856_0))) | (~i_10_18_1005_0 & ((~i_10_18_267_0 & ((~i_10_18_171_0 & ~i_10_18_390_0 & ~i_10_18_960_0 & ~i_10_18_1539_0 & ~i_10_18_1554_0 & ~i_10_18_2001_0 & ~i_10_18_2184_0 & ~i_10_18_2466_0 & ~i_10_18_3069_0 & i_10_18_3841_0) | (i_10_18_796_0 & ~i_10_18_1431_0 & ~i_10_18_2186_0 & ~i_10_18_2460_0 & ~i_10_18_3783_0 & ~i_10_18_3855_0))) | (~i_10_18_446_0 & ~i_10_18_1431_0 & ~i_10_18_1688_0 & i_10_18_1822_0 & ~i_10_18_2179_0 & ~i_10_18_2731_0 & ~i_10_18_3391_0) | (~i_10_18_393_0 & ~i_10_18_960_0 & ~i_10_18_1434_0 & ~i_10_18_1825_0 & ~i_10_18_2185_0 & ~i_10_18_2466_0 & ~i_10_18_2567_0 & ~i_10_18_2605_0 & ~i_10_18_2732_0 & ~i_10_18_2923_0 & ~i_10_18_3070_0 & ~i_10_18_3467_0 & ~i_10_18_3783_0 & ~i_10_18_3834_0))) | (~i_10_18_393_0 & ~i_10_18_2731_0 & ~i_10_18_3069_0 & ((~i_10_18_1431_0 & ~i_10_18_1554_0 & ~i_10_18_1947_0 & ~i_10_18_2179_0 & ~i_10_18_2987_0 & ~i_10_18_3036_0 & ~i_10_18_3095_0 & ~i_10_18_3388_0 & ~i_10_18_3391_0) | (~i_10_18_28_0 & ~i_10_18_1003_0 & ~i_10_18_1691_0 & ~i_10_18_2184_0 & ~i_10_18_2185_0 & ~i_10_18_2466_0 & ~i_10_18_2567_0 & ~i_10_18_3042_0 & ~i_10_18_3471_0 & ~i_10_18_3855_0))) | (i_10_18_175_0 & i_10_18_176_0 & ~i_10_18_1539_0 & ~i_10_18_4291_0))) | (~i_10_18_1431_0 & ((~i_10_18_267_0 & ((~i_10_18_1036_0 & ~i_10_18_1242_0 & i_10_18_1819_0 & ~i_10_18_1947_0 & ~i_10_18_2184_0 & ~i_10_18_2355_0 & ~i_10_18_2565_0 & ~i_10_18_2735_0 & ~i_10_18_3198_0) | (~i_10_18_28_0 & ~i_10_18_1028_0 & ~i_10_18_1554_0 & ~i_10_18_2178_0 & ~i_10_18_2179_0 & ~i_10_18_2185_0 & ~i_10_18_2358_0 & ~i_10_18_3045_0 & ~i_10_18_3069_0 & ~i_10_18_3388_0 & ~i_10_18_3391_0 & ~i_10_18_3471_0))) | (~i_10_18_28_0 & ((~i_10_18_393_0 & ~i_10_18_1554_0 & i_10_18_2725_0 & ~i_10_18_3042_0) | (i_10_18_442_0 & ~i_10_18_1947_0 & ~i_10_18_3045_0 & ~i_10_18_3855_0))) | (~i_10_18_2358_0 & ((~i_10_18_446_0 & i_10_18_1238_0 & ~i_10_18_1539_0 & ~i_10_18_2179_0 & ~i_10_18_2410_0 & ~i_10_18_2567_0 & ~i_10_18_2725_0 & ~i_10_18_3095_0 & ~i_10_18_3391_0) | (~i_10_18_718_0 & ~i_10_18_1006_0 & i_10_18_1691_0 & ~i_10_18_3783_0))) | (~i_10_18_1028_0 & i_10_18_1822_0 & ~i_10_18_3036_0 & ~i_10_18_3198_0 & ~i_10_18_3388_0 & ~i_10_18_3856_0))) | (~i_10_18_1432_0 & ((~i_10_18_960_0 & ((~i_10_18_1005_0 & i_10_18_1238_0 & ~i_10_18_1242_0 & ~i_10_18_2001_0 & ~i_10_18_3095_0) | (~i_10_18_1434_0 & ~i_10_18_1554_0 & ~i_10_18_1575_0 & ~i_10_18_2355_0 & ~i_10_18_2358_0 & ~i_10_18_2567_0 & ~i_10_18_3788_0 & ~i_10_18_3838_0 & ~i_10_18_3841_0 & ~i_10_18_4291_0))) | (i_10_18_1652_0 & i_10_18_1819_0 & ~i_10_18_2178_0 & ~i_10_18_2179_0 & ~i_10_18_2185_0 & ~i_10_18_3045_0))) | (~i_10_18_3042_0 & ((~i_10_18_1005_0 & ((~i_10_18_174_0 & ~i_10_18_1028_0 & ~i_10_18_1238_0 & i_10_18_1825_0 & ~i_10_18_2178_0 & ~i_10_18_2184_0 & ~i_10_18_2355_0 & ~i_10_18_3036_0 & ~i_10_18_3045_0) | (i_10_18_390_0 & ~i_10_18_1003_0 & ~i_10_18_1575_0 & ~i_10_18_2832_0 & ~i_10_18_3841_0 & ~i_10_18_3856_0))) | (~i_10_18_1539_0 & ((~i_10_18_1554_0 & ~i_10_18_2358_0 & ((~i_10_18_2355_0 & ~i_10_18_2731_0 & ~i_10_18_3036_0 & i_10_18_3202_0) | (~i_10_18_390_0 & ~i_10_18_393_0 & ~i_10_18_446_0 & ~i_10_18_718_0 & ~i_10_18_1006_0 & i_10_18_1825_0 & ~i_10_18_2178_0 & ~i_10_18_2410_0 & ~i_10_18_2460_0 & ~i_10_18_3788_0))) | (~i_10_18_28_0 & ~i_10_18_1242_0 & i_10_18_1651_0 & ~i_10_18_1947_0 & ~i_10_18_1950_0 & ~i_10_18_2001_0 & ~i_10_18_2178_0 & ~i_10_18_2460_0 & ~i_10_18_2832_0 & ~i_10_18_2987_0 & ~i_10_18_3198_0))) | (~i_10_18_3036_0 & i_10_18_3467_0 & i_10_18_3610_0))) | (~i_10_18_3855_0 & ((~i_10_18_1312_0 & ((i_10_18_442_0 & i_10_18_3467_0) | (i_10_18_1003_0 & ~i_10_18_2184_0 & ~i_10_18_2987_0 & ~i_10_18_3471_0 & ~i_10_18_3834_0))) | (~i_10_18_2656_0 & i_10_18_3388_0 & ~i_10_18_3391_0 & ~i_10_18_3783_0 & ~i_10_18_3838_0 & ~i_10_18_3841_0))) | (i_10_18_171_0 & ~i_10_18_1539_0 & ~i_10_18_2355_0 & ~i_10_18_2358_0 & i_10_18_3045_0 & ~i_10_18_3471_0));
endmodule



// Benchmark "kernel_10_19" written by ABC on Sun Jul 19 10:21:21 2020

module kernel_10_19 ( 
    i_10_19_219_0, i_10_19_220_0, i_10_19_221_0, i_10_19_269_0,
    i_10_19_282_0, i_10_19_316_0, i_10_19_320_0, i_10_19_329_0,
    i_10_19_431_0, i_10_19_436_0, i_10_19_445_0, i_10_19_446_0,
    i_10_19_464_0, i_10_19_467_0, i_10_19_518_0, i_10_19_752_0,
    i_10_19_799_0, i_10_19_853_0, i_10_19_854_0, i_10_19_899_0,
    i_10_19_956_0, i_10_19_1030_0, i_10_19_1032_0, i_10_19_1082_0,
    i_10_19_1123_0, i_10_19_1220_0, i_10_19_1249_0, i_10_19_1308_0,
    i_10_19_1309_0, i_10_19_1610_0, i_10_19_1618_0, i_10_19_1619_0,
    i_10_19_1822_0, i_10_19_1916_0, i_10_19_1997_0, i_10_19_2004_0,
    i_10_19_2021_0, i_10_19_2023_0, i_10_19_2203_0, i_10_19_2228_0,
    i_10_19_2231_0, i_10_19_2349_0, i_10_19_2350_0, i_10_19_2354_0,
    i_10_19_2365_0, i_10_19_2382_0, i_10_19_2460_0, i_10_19_2463_0,
    i_10_19_2464_0, i_10_19_2470_0, i_10_19_2472_0, i_10_19_2473_0,
    i_10_19_2634_0, i_10_19_2645_0, i_10_19_2678_0, i_10_19_2704_0,
    i_10_19_2723_0, i_10_19_2832_0, i_10_19_2833_0, i_10_19_2834_0,
    i_10_19_2886_0, i_10_19_2984_0, i_10_19_3050_0, i_10_19_3072_0,
    i_10_19_3196_0, i_10_19_3197_0, i_10_19_3278_0, i_10_19_3280_0,
    i_10_19_3283_0, i_10_19_3384_0, i_10_19_3387_0, i_10_19_3388_0,
    i_10_19_3469_0, i_10_19_3495_0, i_10_19_3496_0, i_10_19_3523_0,
    i_10_19_3544_0, i_10_19_3549_0, i_10_19_3651_0, i_10_19_3682_0,
    i_10_19_3684_0, i_10_19_3729_0, i_10_19_3732_0, i_10_19_3839_0,
    i_10_19_3842_0, i_10_19_3856_0, i_10_19_3859_0, i_10_19_3860_0,
    i_10_19_3895_0, i_10_19_3910_0, i_10_19_3913_0, i_10_19_3983_0,
    i_10_19_3988_0, i_10_19_4027_0, i_10_19_4029_0, i_10_19_4030_0,
    i_10_19_4216_0, i_10_19_4277_0, i_10_19_4283_0, i_10_19_4568_0,
    o_10_19_0_0  );
  input  i_10_19_219_0, i_10_19_220_0, i_10_19_221_0, i_10_19_269_0,
    i_10_19_282_0, i_10_19_316_0, i_10_19_320_0, i_10_19_329_0,
    i_10_19_431_0, i_10_19_436_0, i_10_19_445_0, i_10_19_446_0,
    i_10_19_464_0, i_10_19_467_0, i_10_19_518_0, i_10_19_752_0,
    i_10_19_799_0, i_10_19_853_0, i_10_19_854_0, i_10_19_899_0,
    i_10_19_956_0, i_10_19_1030_0, i_10_19_1032_0, i_10_19_1082_0,
    i_10_19_1123_0, i_10_19_1220_0, i_10_19_1249_0, i_10_19_1308_0,
    i_10_19_1309_0, i_10_19_1610_0, i_10_19_1618_0, i_10_19_1619_0,
    i_10_19_1822_0, i_10_19_1916_0, i_10_19_1997_0, i_10_19_2004_0,
    i_10_19_2021_0, i_10_19_2023_0, i_10_19_2203_0, i_10_19_2228_0,
    i_10_19_2231_0, i_10_19_2349_0, i_10_19_2350_0, i_10_19_2354_0,
    i_10_19_2365_0, i_10_19_2382_0, i_10_19_2460_0, i_10_19_2463_0,
    i_10_19_2464_0, i_10_19_2470_0, i_10_19_2472_0, i_10_19_2473_0,
    i_10_19_2634_0, i_10_19_2645_0, i_10_19_2678_0, i_10_19_2704_0,
    i_10_19_2723_0, i_10_19_2832_0, i_10_19_2833_0, i_10_19_2834_0,
    i_10_19_2886_0, i_10_19_2984_0, i_10_19_3050_0, i_10_19_3072_0,
    i_10_19_3196_0, i_10_19_3197_0, i_10_19_3278_0, i_10_19_3280_0,
    i_10_19_3283_0, i_10_19_3384_0, i_10_19_3387_0, i_10_19_3388_0,
    i_10_19_3469_0, i_10_19_3495_0, i_10_19_3496_0, i_10_19_3523_0,
    i_10_19_3544_0, i_10_19_3549_0, i_10_19_3651_0, i_10_19_3682_0,
    i_10_19_3684_0, i_10_19_3729_0, i_10_19_3732_0, i_10_19_3839_0,
    i_10_19_3842_0, i_10_19_3856_0, i_10_19_3859_0, i_10_19_3860_0,
    i_10_19_3895_0, i_10_19_3910_0, i_10_19_3913_0, i_10_19_3983_0,
    i_10_19_3988_0, i_10_19_4027_0, i_10_19_4029_0, i_10_19_4030_0,
    i_10_19_4216_0, i_10_19_4277_0, i_10_19_4283_0, i_10_19_4568_0;
  output o_10_19_0_0;
  assign o_10_19_0_0 = 0;
endmodule



// Benchmark "kernel_10_20" written by ABC on Sun Jul 19 10:21:22 2020

module kernel_10_20 ( 
    i_10_20_49_0, i_10_20_180_0, i_10_20_315_0, i_10_20_405_0,
    i_10_20_431_0, i_10_20_435_0, i_10_20_436_0, i_10_20_439_0,
    i_10_20_444_0, i_10_20_445_0, i_10_20_447_0, i_10_20_449_0,
    i_10_20_467_0, i_10_20_591_0, i_10_20_636_0, i_10_20_700_0,
    i_10_20_735_0, i_10_20_753_0, i_10_20_754_0, i_10_20_799_0,
    i_10_20_1038_0, i_10_20_1039_0, i_10_20_1040_0, i_10_20_1201_0,
    i_10_20_1236_0, i_10_20_1237_0, i_10_20_1238_0, i_10_20_1240_0,
    i_10_20_1552_0, i_10_20_1782_0, i_10_20_1821_0, i_10_20_1822_0,
    i_10_20_1824_0, i_10_20_2147_0, i_10_20_2155_0, i_10_20_2241_0,
    i_10_20_2244_0, i_10_20_2245_0, i_10_20_2307_0, i_10_20_2309_0,
    i_10_20_2310_0, i_10_20_2333_0, i_10_20_2334_0, i_10_20_2352_0,
    i_10_20_2388_0, i_10_20_2460_0, i_10_20_2470_0, i_10_20_2517_0,
    i_10_20_2542_0, i_10_20_2607_0, i_10_20_2633_0, i_10_20_2634_0,
    i_10_20_2635_0, i_10_20_2650_0, i_10_20_2651_0, i_10_20_2677_0,
    i_10_20_2703_0, i_10_20_2704_0, i_10_20_2718_0, i_10_20_2721_0,
    i_10_20_2730_0, i_10_20_2731_0, i_10_20_2732_0, i_10_20_2820_0,
    i_10_20_2830_0, i_10_20_2832_0, i_10_20_2919_0, i_10_20_3271_0,
    i_10_20_3273_0, i_10_20_3387_0, i_10_20_3388_0, i_10_20_3389_0,
    i_10_20_3500_0, i_10_20_3610_0, i_10_20_3614_0, i_10_20_3646_0,
    i_10_20_3649_0, i_10_20_3652_0, i_10_20_3684_0, i_10_20_3685_0,
    i_10_20_3783_0, i_10_20_3786_0, i_10_20_3838_0, i_10_20_3854_0,
    i_10_20_3856_0, i_10_20_3859_0, i_10_20_3881_0, i_10_20_3882_0,
    i_10_20_3982_0, i_10_20_4116_0, i_10_20_4117_0, i_10_20_4118_0,
    i_10_20_4119_0, i_10_20_4120_0, i_10_20_4188_0, i_10_20_4462_0,
    i_10_20_4485_0, i_10_20_4513_0, i_10_20_4516_0, i_10_20_4602_0,
    o_10_20_0_0  );
  input  i_10_20_49_0, i_10_20_180_0, i_10_20_315_0, i_10_20_405_0,
    i_10_20_431_0, i_10_20_435_0, i_10_20_436_0, i_10_20_439_0,
    i_10_20_444_0, i_10_20_445_0, i_10_20_447_0, i_10_20_449_0,
    i_10_20_467_0, i_10_20_591_0, i_10_20_636_0, i_10_20_700_0,
    i_10_20_735_0, i_10_20_753_0, i_10_20_754_0, i_10_20_799_0,
    i_10_20_1038_0, i_10_20_1039_0, i_10_20_1040_0, i_10_20_1201_0,
    i_10_20_1236_0, i_10_20_1237_0, i_10_20_1238_0, i_10_20_1240_0,
    i_10_20_1552_0, i_10_20_1782_0, i_10_20_1821_0, i_10_20_1822_0,
    i_10_20_1824_0, i_10_20_2147_0, i_10_20_2155_0, i_10_20_2241_0,
    i_10_20_2244_0, i_10_20_2245_0, i_10_20_2307_0, i_10_20_2309_0,
    i_10_20_2310_0, i_10_20_2333_0, i_10_20_2334_0, i_10_20_2352_0,
    i_10_20_2388_0, i_10_20_2460_0, i_10_20_2470_0, i_10_20_2517_0,
    i_10_20_2542_0, i_10_20_2607_0, i_10_20_2633_0, i_10_20_2634_0,
    i_10_20_2635_0, i_10_20_2650_0, i_10_20_2651_0, i_10_20_2677_0,
    i_10_20_2703_0, i_10_20_2704_0, i_10_20_2718_0, i_10_20_2721_0,
    i_10_20_2730_0, i_10_20_2731_0, i_10_20_2732_0, i_10_20_2820_0,
    i_10_20_2830_0, i_10_20_2832_0, i_10_20_2919_0, i_10_20_3271_0,
    i_10_20_3273_0, i_10_20_3387_0, i_10_20_3388_0, i_10_20_3389_0,
    i_10_20_3500_0, i_10_20_3610_0, i_10_20_3614_0, i_10_20_3646_0,
    i_10_20_3649_0, i_10_20_3652_0, i_10_20_3684_0, i_10_20_3685_0,
    i_10_20_3783_0, i_10_20_3786_0, i_10_20_3838_0, i_10_20_3854_0,
    i_10_20_3856_0, i_10_20_3859_0, i_10_20_3881_0, i_10_20_3882_0,
    i_10_20_3982_0, i_10_20_4116_0, i_10_20_4117_0, i_10_20_4118_0,
    i_10_20_4119_0, i_10_20_4120_0, i_10_20_4188_0, i_10_20_4462_0,
    i_10_20_4485_0, i_10_20_4513_0, i_10_20_4516_0, i_10_20_4602_0;
  output o_10_20_0_0;
  assign o_10_20_0_0 = 0;
endmodule



// Benchmark "kernel_10_21" written by ABC on Sun Jul 19 10:21:23 2020

module kernel_10_21 ( 
    i_10_21_45_0, i_10_21_185_0, i_10_21_217_0, i_10_21_281_0,
    i_10_21_282_0, i_10_21_283_0, i_10_21_284_0, i_10_21_289_0,
    i_10_21_315_0, i_10_21_405_0, i_10_21_408_0, i_10_21_435_0,
    i_10_21_436_0, i_10_21_462_0, i_10_21_463_0, i_10_21_464_0,
    i_10_21_466_0, i_10_21_892_0, i_10_21_1028_0, i_10_21_1233_0,
    i_10_21_1240_0, i_10_21_1306_0, i_10_21_1307_0, i_10_21_1311_0,
    i_10_21_1363_0, i_10_21_1432_0, i_10_21_1444_0, i_10_21_1540_0,
    i_10_21_1543_0, i_10_21_1576_0, i_10_21_1577_0, i_10_21_1648_0,
    i_10_21_1651_0, i_10_21_1655_0, i_10_21_1675_0, i_10_21_1686_0,
    i_10_21_1687_0, i_10_21_1689_0, i_10_21_1690_0, i_10_21_1819_0,
    i_10_21_1989_0, i_10_21_1990_0, i_10_21_2334_0, i_10_21_2358_0,
    i_10_21_2359_0, i_10_21_2361_0, i_10_21_2362_0, i_10_21_2380_0,
    i_10_21_2457_0, i_10_21_2467_0, i_10_21_2631_0, i_10_21_2709_0,
    i_10_21_2710_0, i_10_21_2719_0, i_10_21_2826_0, i_10_21_2829_0,
    i_10_21_2830_0, i_10_21_2831_0, i_10_21_2834_0, i_10_21_2880_0,
    i_10_21_2881_0, i_10_21_2918_0, i_10_21_2920_0, i_10_21_2921_0,
    i_10_21_3034_0, i_10_21_3037_0, i_10_21_3043_0, i_10_21_3072_0,
    i_10_21_3075_0, i_10_21_3269_0, i_10_21_3277_0, i_10_21_3280_0,
    i_10_21_3324_0, i_10_21_3327_0, i_10_21_3392_0, i_10_21_3408_0,
    i_10_21_3409_0, i_10_21_3466_0, i_10_21_3469_0, i_10_21_3611_0,
    i_10_21_3785_0, i_10_21_3835_0, i_10_21_3838_0, i_10_21_3847_0,
    i_10_21_3848_0, i_10_21_3849_0, i_10_21_3856_0, i_10_21_3857_0,
    i_10_21_3892_0, i_10_21_4116_0, i_10_21_4120_0, i_10_21_4122_0,
    i_10_21_4125_0, i_10_21_4126_0, i_10_21_4212_0, i_10_21_4213_0,
    i_10_21_4267_0, i_10_21_4276_0, i_10_21_4566_0, i_10_21_4567_0,
    o_10_21_0_0  );
  input  i_10_21_45_0, i_10_21_185_0, i_10_21_217_0, i_10_21_281_0,
    i_10_21_282_0, i_10_21_283_0, i_10_21_284_0, i_10_21_289_0,
    i_10_21_315_0, i_10_21_405_0, i_10_21_408_0, i_10_21_435_0,
    i_10_21_436_0, i_10_21_462_0, i_10_21_463_0, i_10_21_464_0,
    i_10_21_466_0, i_10_21_892_0, i_10_21_1028_0, i_10_21_1233_0,
    i_10_21_1240_0, i_10_21_1306_0, i_10_21_1307_0, i_10_21_1311_0,
    i_10_21_1363_0, i_10_21_1432_0, i_10_21_1444_0, i_10_21_1540_0,
    i_10_21_1543_0, i_10_21_1576_0, i_10_21_1577_0, i_10_21_1648_0,
    i_10_21_1651_0, i_10_21_1655_0, i_10_21_1675_0, i_10_21_1686_0,
    i_10_21_1687_0, i_10_21_1689_0, i_10_21_1690_0, i_10_21_1819_0,
    i_10_21_1989_0, i_10_21_1990_0, i_10_21_2334_0, i_10_21_2358_0,
    i_10_21_2359_0, i_10_21_2361_0, i_10_21_2362_0, i_10_21_2380_0,
    i_10_21_2457_0, i_10_21_2467_0, i_10_21_2631_0, i_10_21_2709_0,
    i_10_21_2710_0, i_10_21_2719_0, i_10_21_2826_0, i_10_21_2829_0,
    i_10_21_2830_0, i_10_21_2831_0, i_10_21_2834_0, i_10_21_2880_0,
    i_10_21_2881_0, i_10_21_2918_0, i_10_21_2920_0, i_10_21_2921_0,
    i_10_21_3034_0, i_10_21_3037_0, i_10_21_3043_0, i_10_21_3072_0,
    i_10_21_3075_0, i_10_21_3269_0, i_10_21_3277_0, i_10_21_3280_0,
    i_10_21_3324_0, i_10_21_3327_0, i_10_21_3392_0, i_10_21_3408_0,
    i_10_21_3409_0, i_10_21_3466_0, i_10_21_3469_0, i_10_21_3611_0,
    i_10_21_3785_0, i_10_21_3835_0, i_10_21_3838_0, i_10_21_3847_0,
    i_10_21_3848_0, i_10_21_3849_0, i_10_21_3856_0, i_10_21_3857_0,
    i_10_21_3892_0, i_10_21_4116_0, i_10_21_4120_0, i_10_21_4122_0,
    i_10_21_4125_0, i_10_21_4126_0, i_10_21_4212_0, i_10_21_4213_0,
    i_10_21_4267_0, i_10_21_4276_0, i_10_21_4566_0, i_10_21_4567_0;
  output o_10_21_0_0;
  assign o_10_21_0_0 = ~((~i_10_21_462_0 & ((~i_10_21_1686_0 & ~i_10_21_2710_0 & ~i_10_21_2831_0 & i_10_21_3409_0 & ~i_10_21_3849_0) | (~i_10_21_185_0 & i_10_21_2631_0 & ~i_10_21_2920_0 & ~i_10_21_4567_0))) | (~i_10_21_1240_0 & ((~i_10_21_408_0 & ~i_10_21_466_0 & ~i_10_21_1689_0 & ~i_10_21_2921_0 & ~i_10_21_3409_0 & i_10_21_3838_0 & ~i_10_21_3848_0 & i_10_21_3856_0 & ~i_10_21_4125_0) | (~i_10_21_282_0 & ~i_10_21_283_0 & ~i_10_21_3043_0 & ~i_10_21_3611_0 & ~i_10_21_3838_0 & ~i_10_21_4122_0 & ~i_10_21_4126_0))) | (~i_10_21_3785_0 & ((~i_10_21_185_0 & ((~i_10_21_892_0 & ~i_10_21_1444_0 & i_10_21_1655_0 & ~i_10_21_1990_0 & ~i_10_21_3392_0) | (i_10_21_436_0 & ~i_10_21_3269_0 & ~i_10_21_4120_0 & ~i_10_21_4566_0))) | (~i_10_21_1311_0 & ~i_10_21_4566_0 & ((i_10_21_282_0 & i_10_21_284_0 & ~i_10_21_2362_0 & ~i_10_21_2921_0 & ~i_10_21_3409_0) | (~i_10_21_289_0 & ~i_10_21_408_0 & ~i_10_21_2920_0 & ~i_10_21_3847_0 & ~i_10_21_3857_0))) | (~i_10_21_892_0 & ~i_10_21_1651_0 & ~i_10_21_1686_0 & ~i_10_21_2362_0 & ~i_10_21_3857_0) | (~i_10_21_1233_0 & i_10_21_2631_0 & i_10_21_3280_0) | (~i_10_21_284_0 & ~i_10_21_2358_0 & ~i_10_21_2829_0 & ~i_10_21_2831_0 & ~i_10_21_3072_0 & ~i_10_21_4122_0))) | (~i_10_21_1990_0 & ((~i_10_21_892_0 & ((~i_10_21_408_0 & ~i_10_21_1363_0 & ~i_10_21_2831_0 & ~i_10_21_2834_0 & ~i_10_21_3269_0 & ~i_10_21_3392_0 & ~i_10_21_4116_0 & ~i_10_21_4120_0) | (i_10_21_1240_0 & ~i_10_21_2826_0 & ~i_10_21_2830_0 & ~i_10_21_4566_0))) | (i_10_21_1651_0 & ~i_10_21_1989_0 & ~i_10_21_2709_0 & ~i_10_21_2829_0 & ~i_10_21_3043_0 & ~i_10_21_3392_0 & ~i_10_21_3409_0 & ~i_10_21_4212_0))) | (~i_10_21_408_0 & ((~i_10_21_2359_0 & ~i_10_21_2380_0 & ~i_10_21_2709_0 & ~i_10_21_2830_0 & ~i_10_21_3392_0) | (~i_10_21_217_0 & ~i_10_21_284_0 & ~i_10_21_2358_0 & ~i_10_21_3043_0 & ~i_10_21_3075_0 & ~i_10_21_3856_0))) | (~i_10_21_2359_0 & ((i_10_21_1306_0 & ~i_10_21_2361_0) | (~i_10_21_282_0 & i_10_21_1648_0 & i_10_21_4116_0))) | (~i_10_21_282_0 & ((~i_10_21_185_0 & ~i_10_21_2362_0 & ~i_10_21_2709_0 & ~i_10_21_2918_0 & ~i_10_21_3072_0 & ~i_10_21_3392_0) | (~i_10_21_284_0 & i_10_21_1686_0 & ~i_10_21_2831_0 & ~i_10_21_3269_0 & ~i_10_21_4126_0))) | (~i_10_21_1444_0 & ((~i_10_21_185_0 & ~i_10_21_2362_0 & ((~i_10_21_1989_0 & ~i_10_21_2361_0 & ~i_10_21_2831_0) | (~i_10_21_405_0 & ~i_10_21_435_0 & ~i_10_21_464_0 & ~i_10_21_2334_0 & ~i_10_21_2457_0 & ~i_10_21_2719_0 & ~i_10_21_2834_0 & ~i_10_21_3037_0 & ~i_10_21_3849_0))) | (~i_10_21_284_0 & ~i_10_21_1690_0 & ~i_10_21_2920_0 & ~i_10_21_3849_0 & i_10_21_4566_0 & i_10_21_4567_0))) | (~i_10_21_284_0 & (i_10_21_1543_0 | (~i_10_21_1651_0 & i_10_21_1690_0 & ~i_10_21_2631_0 & i_10_21_3075_0))) | (~i_10_21_4567_0 & ((i_10_21_466_0 & i_10_21_1655_0 & ~i_10_21_2829_0 & ~i_10_21_2921_0) | (i_10_21_2359_0 & ~i_10_21_2631_0 & i_10_21_2921_0 & i_10_21_3611_0 & ~i_10_21_3848_0))) | (i_10_21_281_0 & ~i_10_21_1363_0 & i_10_21_2826_0 & ~i_10_21_2920_0 & i_10_21_4116_0));
endmodule



// Benchmark "kernel_10_22" written by ABC on Sun Jul 19 10:21:24 2020

module kernel_10_22 ( 
    i_10_22_21_0, i_10_22_22_0, i_10_22_48_0, i_10_22_134_0, i_10_22_180_0,
    i_10_22_181_0, i_10_22_184_0, i_10_22_185_0, i_10_22_428_0,
    i_10_22_433_0, i_10_22_515_0, i_10_22_599_0, i_10_22_639_0,
    i_10_22_640_0, i_10_22_716_0, i_10_22_759_0, i_10_22_793_0,
    i_10_22_798_0, i_10_22_799_0, i_10_22_950_0, i_10_22_1000_0,
    i_10_22_1028_0, i_10_22_1131_0, i_10_22_1164_0, i_10_22_1171_0,
    i_10_22_1238_0, i_10_22_1246_0, i_10_22_1247_0, i_10_22_1312_0,
    i_10_22_1447_0, i_10_22_1453_0, i_10_22_1541_0, i_10_22_1607_0,
    i_10_22_1616_0, i_10_22_1632_0, i_10_22_1633_0, i_10_22_1786_0,
    i_10_22_1823_0, i_10_22_1826_0, i_10_22_1882_0, i_10_22_1909_0,
    i_10_22_1912_0, i_10_22_1992_0, i_10_22_2011_0, i_10_22_2012_0,
    i_10_22_2091_0, i_10_22_2162_0, i_10_22_2335_0, i_10_22_2349_0,
    i_10_22_2365_0, i_10_22_2383_0, i_10_22_2439_0, i_10_22_2441_0,
    i_10_22_2461_0, i_10_22_2578_0, i_10_22_2604_0, i_10_22_2608_0,
    i_10_22_2640_0, i_10_22_2649_0, i_10_22_2686_0, i_10_22_2711_0,
    i_10_22_2747_0, i_10_22_2828_0, i_10_22_2866_0, i_10_22_2885_0,
    i_10_22_2918_0, i_10_22_2922_0, i_10_22_2923_0, i_10_22_3083_0,
    i_10_22_3088_0, i_10_22_3107_0, i_10_22_3202_0, i_10_22_3226_0,
    i_10_22_3234_0, i_10_22_3439_0, i_10_22_3537_0, i_10_22_3538_0,
    i_10_22_3623_0, i_10_22_3650_0, i_10_22_3721_0, i_10_22_3786_0,
    i_10_22_3787_0, i_10_22_3788_0, i_10_22_3835_0, i_10_22_3836_0,
    i_10_22_3889_0, i_10_22_3892_0, i_10_22_3963_0, i_10_22_3964_0,
    i_10_22_4152_0, i_10_22_4157_0, i_10_22_4185_0, i_10_22_4186_0,
    i_10_22_4188_0, i_10_22_4190_0, i_10_22_4217_0, i_10_22_4287_0,
    i_10_22_4435_0, i_10_22_4457_0, i_10_22_4462_0,
    o_10_22_0_0  );
  input  i_10_22_21_0, i_10_22_22_0, i_10_22_48_0, i_10_22_134_0,
    i_10_22_180_0, i_10_22_181_0, i_10_22_184_0, i_10_22_185_0,
    i_10_22_428_0, i_10_22_433_0, i_10_22_515_0, i_10_22_599_0,
    i_10_22_639_0, i_10_22_640_0, i_10_22_716_0, i_10_22_759_0,
    i_10_22_793_0, i_10_22_798_0, i_10_22_799_0, i_10_22_950_0,
    i_10_22_1000_0, i_10_22_1028_0, i_10_22_1131_0, i_10_22_1164_0,
    i_10_22_1171_0, i_10_22_1238_0, i_10_22_1246_0, i_10_22_1247_0,
    i_10_22_1312_0, i_10_22_1447_0, i_10_22_1453_0, i_10_22_1541_0,
    i_10_22_1607_0, i_10_22_1616_0, i_10_22_1632_0, i_10_22_1633_0,
    i_10_22_1786_0, i_10_22_1823_0, i_10_22_1826_0, i_10_22_1882_0,
    i_10_22_1909_0, i_10_22_1912_0, i_10_22_1992_0, i_10_22_2011_0,
    i_10_22_2012_0, i_10_22_2091_0, i_10_22_2162_0, i_10_22_2335_0,
    i_10_22_2349_0, i_10_22_2365_0, i_10_22_2383_0, i_10_22_2439_0,
    i_10_22_2441_0, i_10_22_2461_0, i_10_22_2578_0, i_10_22_2604_0,
    i_10_22_2608_0, i_10_22_2640_0, i_10_22_2649_0, i_10_22_2686_0,
    i_10_22_2711_0, i_10_22_2747_0, i_10_22_2828_0, i_10_22_2866_0,
    i_10_22_2885_0, i_10_22_2918_0, i_10_22_2922_0, i_10_22_2923_0,
    i_10_22_3083_0, i_10_22_3088_0, i_10_22_3107_0, i_10_22_3202_0,
    i_10_22_3226_0, i_10_22_3234_0, i_10_22_3439_0, i_10_22_3537_0,
    i_10_22_3538_0, i_10_22_3623_0, i_10_22_3650_0, i_10_22_3721_0,
    i_10_22_3786_0, i_10_22_3787_0, i_10_22_3788_0, i_10_22_3835_0,
    i_10_22_3836_0, i_10_22_3889_0, i_10_22_3892_0, i_10_22_3963_0,
    i_10_22_3964_0, i_10_22_4152_0, i_10_22_4157_0, i_10_22_4185_0,
    i_10_22_4186_0, i_10_22_4188_0, i_10_22_4190_0, i_10_22_4217_0,
    i_10_22_4287_0, i_10_22_4435_0, i_10_22_4457_0, i_10_22_4462_0;
  output o_10_22_0_0;
  assign o_10_22_0_0 = 0;
endmodule



// Benchmark "kernel_10_23" written by ABC on Sun Jul 19 10:21:25 2020

module kernel_10_23 ( 
    i_10_23_224_0, i_10_23_293_0, i_10_23_409_0, i_10_23_410_0,
    i_10_23_444_0, i_10_23_445_0, i_10_23_447_0, i_10_23_643_0,
    i_10_23_646_0, i_10_23_797_0, i_10_23_1000_0, i_10_23_1123_0,
    i_10_23_1172_0, i_10_23_1216_0, i_10_23_1264_0, i_10_23_1313_0,
    i_10_23_1348_0, i_10_23_1543_0, i_10_23_1578_0, i_10_23_1579_0,
    i_10_23_1580_0, i_10_23_1582_0, i_10_23_1583_0, i_10_23_1648_0,
    i_10_23_1724_0, i_10_23_1810_0, i_10_23_1821_0, i_10_23_1826_0,
    i_10_23_1991_0, i_10_23_1994_0, i_10_23_2023_0, i_10_23_2352_0,
    i_10_23_2354_0, i_10_23_2360_0, i_10_23_2363_0, i_10_23_2365_0,
    i_10_23_2366_0, i_10_23_2380_0, i_10_23_2381_0, i_10_23_2384_0,
    i_10_23_2453_0, i_10_23_2466_0, i_10_23_2656_0, i_10_23_2657_0,
    i_10_23_2700_0, i_10_23_2708_0, i_10_23_2711_0, i_10_23_2714_0,
    i_10_23_2717_0, i_10_23_2718_0, i_10_23_2719_0, i_10_23_2720_0,
    i_10_23_2723_0, i_10_23_2729_0, i_10_23_2730_0, i_10_23_2732_0,
    i_10_23_2734_0, i_10_23_2735_0, i_10_23_2828_0, i_10_23_2831_0,
    i_10_23_3038_0, i_10_23_3230_0, i_10_23_3287_0, i_10_23_3290_0,
    i_10_23_3301_0, i_10_23_3302_0, i_10_23_3384_0, i_10_23_3388_0,
    i_10_23_3389_0, i_10_23_3403_0, i_10_23_3406_0, i_10_23_3430_0,
    i_10_23_3461_0, i_10_23_3467_0, i_10_23_3520_0, i_10_23_3523_0,
    i_10_23_3524_0, i_10_23_3587_0, i_10_23_3611_0, i_10_23_3614_0,
    i_10_23_3650_0, i_10_23_3689_0, i_10_23_3728_0, i_10_23_3785_0,
    i_10_23_3852_0, i_10_23_3855_0, i_10_23_3857_0, i_10_23_3893_0,
    i_10_23_3923_0, i_10_23_3994_0, i_10_23_4118_0, i_10_23_4120_0,
    i_10_23_4121_0, i_10_23_4169_0, i_10_23_4271_0, i_10_23_4273_0,
    i_10_23_4275_0, i_10_23_4289_0, i_10_23_4461_0, i_10_23_4571_0,
    o_10_23_0_0  );
  input  i_10_23_224_0, i_10_23_293_0, i_10_23_409_0, i_10_23_410_0,
    i_10_23_444_0, i_10_23_445_0, i_10_23_447_0, i_10_23_643_0,
    i_10_23_646_0, i_10_23_797_0, i_10_23_1000_0, i_10_23_1123_0,
    i_10_23_1172_0, i_10_23_1216_0, i_10_23_1264_0, i_10_23_1313_0,
    i_10_23_1348_0, i_10_23_1543_0, i_10_23_1578_0, i_10_23_1579_0,
    i_10_23_1580_0, i_10_23_1582_0, i_10_23_1583_0, i_10_23_1648_0,
    i_10_23_1724_0, i_10_23_1810_0, i_10_23_1821_0, i_10_23_1826_0,
    i_10_23_1991_0, i_10_23_1994_0, i_10_23_2023_0, i_10_23_2352_0,
    i_10_23_2354_0, i_10_23_2360_0, i_10_23_2363_0, i_10_23_2365_0,
    i_10_23_2366_0, i_10_23_2380_0, i_10_23_2381_0, i_10_23_2384_0,
    i_10_23_2453_0, i_10_23_2466_0, i_10_23_2656_0, i_10_23_2657_0,
    i_10_23_2700_0, i_10_23_2708_0, i_10_23_2711_0, i_10_23_2714_0,
    i_10_23_2717_0, i_10_23_2718_0, i_10_23_2719_0, i_10_23_2720_0,
    i_10_23_2723_0, i_10_23_2729_0, i_10_23_2730_0, i_10_23_2732_0,
    i_10_23_2734_0, i_10_23_2735_0, i_10_23_2828_0, i_10_23_2831_0,
    i_10_23_3038_0, i_10_23_3230_0, i_10_23_3287_0, i_10_23_3290_0,
    i_10_23_3301_0, i_10_23_3302_0, i_10_23_3384_0, i_10_23_3388_0,
    i_10_23_3389_0, i_10_23_3403_0, i_10_23_3406_0, i_10_23_3430_0,
    i_10_23_3461_0, i_10_23_3467_0, i_10_23_3520_0, i_10_23_3523_0,
    i_10_23_3524_0, i_10_23_3587_0, i_10_23_3611_0, i_10_23_3614_0,
    i_10_23_3650_0, i_10_23_3689_0, i_10_23_3728_0, i_10_23_3785_0,
    i_10_23_3852_0, i_10_23_3855_0, i_10_23_3857_0, i_10_23_3893_0,
    i_10_23_3923_0, i_10_23_3994_0, i_10_23_4118_0, i_10_23_4120_0,
    i_10_23_4121_0, i_10_23_4169_0, i_10_23_4271_0, i_10_23_4273_0,
    i_10_23_4275_0, i_10_23_4289_0, i_10_23_4461_0, i_10_23_4571_0;
  output o_10_23_0_0;
  assign o_10_23_0_0 = 0;
endmodule



// Benchmark "kernel_10_24" written by ABC on Sun Jul 19 10:21:26 2020

module kernel_10_24 ( 
    i_10_24_82_0, i_10_24_181_0, i_10_24_210_0, i_10_24_216_0,
    i_10_24_217_0, i_10_24_221_0, i_10_24_271_0, i_10_24_274_0,
    i_10_24_275_0, i_10_24_281_0, i_10_24_406_0, i_10_24_409_0,
    i_10_24_437_0, i_10_24_449_0, i_10_24_482_0, i_10_24_508_0,
    i_10_24_826_0, i_10_24_892_0, i_10_24_944_0, i_10_24_963_0,
    i_10_24_1060_0, i_10_24_1080_0, i_10_24_1117_0, i_10_24_1242_0,
    i_10_24_1243_0, i_10_24_1248_0, i_10_24_1249_0, i_10_24_1310_0,
    i_10_24_1354_0, i_10_24_1355_0, i_10_24_1359_0, i_10_24_1360_0,
    i_10_24_1575_0, i_10_24_1576_0, i_10_24_1603_0, i_10_24_1617_0,
    i_10_24_1688_0, i_10_24_1765_0, i_10_24_1786_0, i_10_24_1881_0,
    i_10_24_1903_0, i_10_24_1922_0, i_10_24_2020_0, i_10_24_2197_0,
    i_10_24_2331_0, i_10_24_2332_0, i_10_24_2367_0, i_10_24_2450_0,
    i_10_24_2502_0, i_10_24_2540_0, i_10_24_2631_0, i_10_24_2638_0,
    i_10_24_2646_0, i_10_24_2647_0, i_10_24_2704_0, i_10_24_2728_0,
    i_10_24_2862_0, i_10_24_2869_0, i_10_24_2872_0, i_10_24_2916_0,
    i_10_24_2919_0, i_10_24_2920_0, i_10_24_2953_0, i_10_24_3054_0,
    i_10_24_3195_0, i_10_24_3262_0, i_10_24_3384_0, i_10_24_3550_0,
    i_10_24_3610_0, i_10_24_3611_0, i_10_24_3720_0, i_10_24_3721_0,
    i_10_24_3846_0, i_10_24_3847_0, i_10_24_3848_0, i_10_24_3851_0,
    i_10_24_3856_0, i_10_24_3884_0, i_10_24_3888_0, i_10_24_3889_0,
    i_10_24_3915_0, i_10_24_3960_0, i_10_24_3961_0, i_10_24_3963_0,
    i_10_24_3964_0, i_10_24_4023_0, i_10_24_4024_0, i_10_24_4025_0,
    i_10_24_4118_0, i_10_24_4177_0, i_10_24_4185_0, i_10_24_4186_0,
    i_10_24_4188_0, i_10_24_4287_0, i_10_24_4325_0, i_10_24_4420_0,
    i_10_24_4428_0, i_10_24_4510_0, i_10_24_4527_0, i_10_24_4600_0,
    o_10_24_0_0  );
  input  i_10_24_82_0, i_10_24_181_0, i_10_24_210_0, i_10_24_216_0,
    i_10_24_217_0, i_10_24_221_0, i_10_24_271_0, i_10_24_274_0,
    i_10_24_275_0, i_10_24_281_0, i_10_24_406_0, i_10_24_409_0,
    i_10_24_437_0, i_10_24_449_0, i_10_24_482_0, i_10_24_508_0,
    i_10_24_826_0, i_10_24_892_0, i_10_24_944_0, i_10_24_963_0,
    i_10_24_1060_0, i_10_24_1080_0, i_10_24_1117_0, i_10_24_1242_0,
    i_10_24_1243_0, i_10_24_1248_0, i_10_24_1249_0, i_10_24_1310_0,
    i_10_24_1354_0, i_10_24_1355_0, i_10_24_1359_0, i_10_24_1360_0,
    i_10_24_1575_0, i_10_24_1576_0, i_10_24_1603_0, i_10_24_1617_0,
    i_10_24_1688_0, i_10_24_1765_0, i_10_24_1786_0, i_10_24_1881_0,
    i_10_24_1903_0, i_10_24_1922_0, i_10_24_2020_0, i_10_24_2197_0,
    i_10_24_2331_0, i_10_24_2332_0, i_10_24_2367_0, i_10_24_2450_0,
    i_10_24_2502_0, i_10_24_2540_0, i_10_24_2631_0, i_10_24_2638_0,
    i_10_24_2646_0, i_10_24_2647_0, i_10_24_2704_0, i_10_24_2728_0,
    i_10_24_2862_0, i_10_24_2869_0, i_10_24_2872_0, i_10_24_2916_0,
    i_10_24_2919_0, i_10_24_2920_0, i_10_24_2953_0, i_10_24_3054_0,
    i_10_24_3195_0, i_10_24_3262_0, i_10_24_3384_0, i_10_24_3550_0,
    i_10_24_3610_0, i_10_24_3611_0, i_10_24_3720_0, i_10_24_3721_0,
    i_10_24_3846_0, i_10_24_3847_0, i_10_24_3848_0, i_10_24_3851_0,
    i_10_24_3856_0, i_10_24_3884_0, i_10_24_3888_0, i_10_24_3889_0,
    i_10_24_3915_0, i_10_24_3960_0, i_10_24_3961_0, i_10_24_3963_0,
    i_10_24_3964_0, i_10_24_4023_0, i_10_24_4024_0, i_10_24_4025_0,
    i_10_24_4118_0, i_10_24_4177_0, i_10_24_4185_0, i_10_24_4186_0,
    i_10_24_4188_0, i_10_24_4287_0, i_10_24_4325_0, i_10_24_4420_0,
    i_10_24_4428_0, i_10_24_4510_0, i_10_24_4527_0, i_10_24_4600_0;
  output o_10_24_0_0;
  assign o_10_24_0_0 = 0;
endmodule



// Benchmark "kernel_10_25" written by ABC on Sun Jul 19 10:21:27 2020

module kernel_10_25 ( 
    i_10_25_35_0, i_10_25_172_0, i_10_25_174_0, i_10_25_175_0,
    i_10_25_176_0, i_10_25_178_0, i_10_25_183_0, i_10_25_220_0,
    i_10_25_221_0, i_10_25_272_0, i_10_25_285_0, i_10_25_286_0,
    i_10_25_328_0, i_10_25_410_0, i_10_25_429_0, i_10_25_460_0,
    i_10_25_711_0, i_10_25_795_0, i_10_25_796_0, i_10_25_907_0,
    i_10_25_961_0, i_10_25_999_0, i_10_25_1006_0, i_10_25_1168_0,
    i_10_25_1169_0, i_10_25_1236_0, i_10_25_1244_0, i_10_25_1263_0,
    i_10_25_1580_0, i_10_25_1583_0, i_10_25_1654_0, i_10_25_1686_0,
    i_10_25_1689_0, i_10_25_1691_0, i_10_25_1821_0, i_10_25_1822_0,
    i_10_25_1823_0, i_10_25_1910_0, i_10_25_1913_0, i_10_25_2022_0,
    i_10_25_2349_0, i_10_25_2350_0, i_10_25_2351_0, i_10_25_2352_0,
    i_10_25_2353_0, i_10_25_2354_0, i_10_25_2379_0, i_10_25_2407_0,
    i_10_25_2409_0, i_10_25_2410_0, i_10_25_2451_0, i_10_25_2452_0,
    i_10_25_2453_0, i_10_25_2681_0, i_10_25_2703_0, i_10_25_2708_0,
    i_10_25_2711_0, i_10_25_2714_0, i_10_25_2722_0, i_10_25_2725_0,
    i_10_25_2733_0, i_10_25_2734_0, i_10_25_2735_0, i_10_25_2828_0,
    i_10_25_3036_0, i_10_25_3153_0, i_10_25_3165_0, i_10_25_3195_0,
    i_10_25_3196_0, i_10_25_3202_0, i_10_25_3231_0, i_10_25_3237_0,
    i_10_25_3279_0, i_10_25_3281_0, i_10_25_3325_0, i_10_25_3388_0,
    i_10_25_3613_0, i_10_25_3614_0, i_10_25_3616_0, i_10_25_3646_0,
    i_10_25_3649_0, i_10_25_3723_0, i_10_25_3724_0, i_10_25_3781_0,
    i_10_25_3838_0, i_10_25_3839_0, i_10_25_3846_0, i_10_25_3856_0,
    i_10_25_3857_0, i_10_25_3859_0, i_10_25_3883_0, i_10_25_3895_0,
    i_10_25_3913_0, i_10_25_3991_0, i_10_25_4120_0, i_10_25_4121_0,
    i_10_25_4129_0, i_10_25_4174_0, i_10_25_4269_0, i_10_25_4283_0,
    o_10_25_0_0  );
  input  i_10_25_35_0, i_10_25_172_0, i_10_25_174_0, i_10_25_175_0,
    i_10_25_176_0, i_10_25_178_0, i_10_25_183_0, i_10_25_220_0,
    i_10_25_221_0, i_10_25_272_0, i_10_25_285_0, i_10_25_286_0,
    i_10_25_328_0, i_10_25_410_0, i_10_25_429_0, i_10_25_460_0,
    i_10_25_711_0, i_10_25_795_0, i_10_25_796_0, i_10_25_907_0,
    i_10_25_961_0, i_10_25_999_0, i_10_25_1006_0, i_10_25_1168_0,
    i_10_25_1169_0, i_10_25_1236_0, i_10_25_1244_0, i_10_25_1263_0,
    i_10_25_1580_0, i_10_25_1583_0, i_10_25_1654_0, i_10_25_1686_0,
    i_10_25_1689_0, i_10_25_1691_0, i_10_25_1821_0, i_10_25_1822_0,
    i_10_25_1823_0, i_10_25_1910_0, i_10_25_1913_0, i_10_25_2022_0,
    i_10_25_2349_0, i_10_25_2350_0, i_10_25_2351_0, i_10_25_2352_0,
    i_10_25_2353_0, i_10_25_2354_0, i_10_25_2379_0, i_10_25_2407_0,
    i_10_25_2409_0, i_10_25_2410_0, i_10_25_2451_0, i_10_25_2452_0,
    i_10_25_2453_0, i_10_25_2681_0, i_10_25_2703_0, i_10_25_2708_0,
    i_10_25_2711_0, i_10_25_2714_0, i_10_25_2722_0, i_10_25_2725_0,
    i_10_25_2733_0, i_10_25_2734_0, i_10_25_2735_0, i_10_25_2828_0,
    i_10_25_3036_0, i_10_25_3153_0, i_10_25_3165_0, i_10_25_3195_0,
    i_10_25_3196_0, i_10_25_3202_0, i_10_25_3231_0, i_10_25_3237_0,
    i_10_25_3279_0, i_10_25_3281_0, i_10_25_3325_0, i_10_25_3388_0,
    i_10_25_3613_0, i_10_25_3614_0, i_10_25_3616_0, i_10_25_3646_0,
    i_10_25_3649_0, i_10_25_3723_0, i_10_25_3724_0, i_10_25_3781_0,
    i_10_25_3838_0, i_10_25_3839_0, i_10_25_3846_0, i_10_25_3856_0,
    i_10_25_3857_0, i_10_25_3859_0, i_10_25_3883_0, i_10_25_3895_0,
    i_10_25_3913_0, i_10_25_3991_0, i_10_25_4120_0, i_10_25_4121_0,
    i_10_25_4129_0, i_10_25_4174_0, i_10_25_4269_0, i_10_25_4283_0;
  output o_10_25_0_0;
  assign o_10_25_0_0 = ~((~i_10_25_286_0 & ((~i_10_25_172_0 & ~i_10_25_1821_0 & ~i_10_25_3895_0 & ~i_10_25_3913_0 & ~i_10_25_3991_0) | (~i_10_25_410_0 & ~i_10_25_1168_0 & ~i_10_25_1822_0 & ~i_10_25_2733_0 & ~i_10_25_3279_0 & ~i_10_25_4120_0))) | (~i_10_25_172_0 & ((~i_10_25_1654_0 & ~i_10_25_2349_0 & ~i_10_25_2452_0 & ~i_10_25_2681_0 & ~i_10_25_3231_0 & ~i_10_25_3237_0) | (~i_10_25_220_0 & ~i_10_25_1168_0 & ~i_10_25_1583_0 & ~i_10_25_2703_0 & ~i_10_25_3165_0 & ~i_10_25_3846_0 & ~i_10_25_3991_0))) | (~i_10_25_220_0 & ((~i_10_25_410_0 & ~i_10_25_1821_0 & ~i_10_25_2708_0 & ~i_10_25_3165_0 & ~i_10_25_3237_0 & ~i_10_25_3781_0) | (~i_10_25_176_0 & ~i_10_25_1913_0 & i_10_25_2349_0 & ~i_10_25_2703_0 & ~i_10_25_2725_0 & ~i_10_25_2828_0 & ~i_10_25_3649_0 & i_10_25_3838_0 & ~i_10_25_4120_0))) | (~i_10_25_3165_0 & ((~i_10_25_711_0 & ((~i_10_25_174_0 & ((~i_10_25_796_0 & ~i_10_25_907_0 & ~i_10_25_1168_0 & ~i_10_25_2451_0 & ~i_10_25_2725_0) | (~i_10_25_1236_0 & ~i_10_25_2351_0 & ~i_10_25_3196_0 & ~i_10_25_3895_0 & ~i_10_25_3991_0))) | (~i_10_25_410_0 & ((~i_10_25_2350_0 & ~i_10_25_2703_0 & i_10_25_2722_0 & ~i_10_25_3781_0 & ~i_10_25_3839_0) | (~i_10_25_175_0 & ~i_10_25_2734_0 & ~i_10_25_3195_0 & ~i_10_25_3237_0 & ~i_10_25_3991_0 & ~i_10_25_4174_0))) | (~i_10_25_3281_0 & ~i_10_25_3991_0 & ((~i_10_25_795_0 & ~i_10_25_999_0 & ~i_10_25_1691_0 & i_10_25_2452_0 & ~i_10_25_2708_0) | (~i_10_25_460_0 & ~i_10_25_1168_0 & ~i_10_25_1654_0 & ~i_10_25_2022_0 & ~i_10_25_2714_0))))) | (~i_10_25_3237_0 & ((~i_10_25_174_0 & ~i_10_25_1169_0 & ~i_10_25_1583_0 & ~i_10_25_2451_0 & ~i_10_25_2711_0) | (~i_10_25_460_0 & ~i_10_25_907_0 & ~i_10_25_1823_0 & ~i_10_25_2022_0 & ~i_10_25_3036_0 & ~i_10_25_3195_0 & ~i_10_25_3231_0))) | (~i_10_25_221_0 & ~i_10_25_795_0 & ~i_10_25_2708_0 & ~i_10_25_3196_0 & ~i_10_25_3616_0 & ~i_10_25_3839_0 & ~i_10_25_3846_0 & ~i_10_25_4269_0))) | (~i_10_25_174_0 & ~i_10_25_2711_0 & ((~i_10_25_907_0 & ~i_10_25_1691_0 & ~i_10_25_2352_0 & ~i_10_25_3195_0 & i_10_25_3646_0) | (~i_10_25_796_0 & ~i_10_25_2022_0 & ~i_10_25_3838_0 & ~i_10_25_3839_0))) | (~i_10_25_175_0 & ((~i_10_25_1236_0 & ~i_10_25_2735_0 & i_10_25_3281_0) | (~i_10_25_907_0 & ~i_10_25_1244_0 & ~i_10_25_1910_0 & ~i_10_25_2451_0 & ~i_10_25_3281_0 & ~i_10_25_4174_0))) | (~i_10_25_1821_0 & ((~i_10_25_1168_0 & ~i_10_25_1236_0 & ~i_10_25_1580_0 & ~i_10_25_2453_0 & ~i_10_25_3196_0 & ~i_10_25_3279_0) | (~i_10_25_328_0 & ~i_10_25_3388_0 & i_10_25_3859_0))) | (~i_10_25_1168_0 & ((~i_10_25_183_0 & ~i_10_25_460_0 & ~i_10_25_2349_0 & i_10_25_2452_0 & ~i_10_25_2733_0 & ~i_10_25_3231_0 & ~i_10_25_3614_0 & ~i_10_25_3616_0) | (~i_10_25_999_0 & ~i_10_25_1823_0 & ~i_10_25_2451_0 & ~i_10_25_3913_0 & ~i_10_25_3991_0 & ~i_10_25_4283_0))) | (~i_10_25_1236_0 & ((~i_10_25_1910_0 & ~i_10_25_2451_0 & ~i_10_25_2452_0 & ~i_10_25_2733_0 & ~i_10_25_3279_0 & i_10_25_4121_0) | (~i_10_25_711_0 & ~i_10_25_1823_0 & ~i_10_25_2022_0 & i_10_25_3616_0 & ~i_10_25_3913_0 & ~i_10_25_4269_0))) | (~i_10_25_2451_0 & ((~i_10_25_796_0 & ~i_10_25_2452_0 & ~i_10_25_3196_0 & ~i_10_25_3913_0) | (~i_10_25_2453_0 & ~i_10_25_3036_0 & ~i_10_25_3613_0 & ~i_10_25_3846_0 & ~i_10_25_4174_0))) | (~i_10_25_3838_0 & ~i_10_25_3895_0 & ((~i_10_25_429_0 & ~i_10_25_2353_0 & ~i_10_25_2722_0 & i_10_25_3388_0) | (i_10_25_2708_0 & ~i_10_25_4129_0))) | (~i_10_25_2733_0 & i_10_25_3202_0 & ~i_10_25_3781_0 & i_10_25_3839_0 & ~i_10_25_3859_0));
endmodule



// Benchmark "kernel_10_26" written by ABC on Sun Jul 19 10:21:29 2020

module kernel_10_26 ( 
    i_10_26_174_0, i_10_26_176_0, i_10_26_286_0, i_10_26_293_0,
    i_10_26_296_0, i_10_26_326_0, i_10_26_328_0, i_10_26_394_0,
    i_10_26_429_0, i_10_26_444_0, i_10_26_445_0, i_10_26_447_0,
    i_10_26_448_0, i_10_26_465_0, i_10_26_792_0, i_10_26_798_0,
    i_10_26_799_0, i_10_26_955_0, i_10_26_1002_0, i_10_26_1032_0,
    i_10_26_1034_0, i_10_26_1240_0, i_10_26_1241_0, i_10_26_1265_0,
    i_10_26_1305_0, i_10_26_1306_0, i_10_26_1309_0, i_10_26_1651_0,
    i_10_26_1819_0, i_10_26_1821_0, i_10_26_1826_0, i_10_26_1911_0,
    i_10_26_1989_0, i_10_26_1995_0, i_10_26_1996_0, i_10_26_2311_0,
    i_10_26_2349_0, i_10_26_2351_0, i_10_26_2357_0, i_10_26_2364_0,
    i_10_26_2452_0, i_10_26_2571_0, i_10_26_2655_0, i_10_26_2656_0,
    i_10_26_2657_0, i_10_26_2658_0, i_10_26_2659_0, i_10_26_2703_0,
    i_10_26_2704_0, i_10_26_2714_0, i_10_26_2727_0, i_10_26_2728_0,
    i_10_26_2730_0, i_10_26_2731_0, i_10_26_2732_0, i_10_26_2787_0,
    i_10_26_2788_0, i_10_26_2819_0, i_10_26_2884_0, i_10_26_2985_0,
    i_10_26_2987_0, i_10_26_3039_0, i_10_26_3045_0, i_10_26_3046_0,
    i_10_26_3048_0, i_10_26_3049_0, i_10_26_3075_0, i_10_26_3076_0,
    i_10_26_3091_0, i_10_26_3094_0, i_10_26_3195_0, i_10_26_3198_0,
    i_10_26_3271_0, i_10_26_3272_0, i_10_26_3298_0, i_10_26_3326_0,
    i_10_26_3405_0, i_10_26_3407_0, i_10_26_3408_0, i_10_26_3409_0,
    i_10_26_3472_0, i_10_26_3613_0, i_10_26_3646_0, i_10_26_3855_0,
    i_10_26_3857_0, i_10_26_3860_0, i_10_26_3983_0, i_10_26_3985_0,
    i_10_26_3986_0, i_10_26_4115_0, i_10_26_4116_0, i_10_26_4117_0,
    i_10_26_4128_0, i_10_26_4216_0, i_10_26_4269_0, i_10_26_4270_0,
    i_10_26_4271_0, i_10_26_4278_0, i_10_26_4288_0, i_10_26_4568_0,
    o_10_26_0_0  );
  input  i_10_26_174_0, i_10_26_176_0, i_10_26_286_0, i_10_26_293_0,
    i_10_26_296_0, i_10_26_326_0, i_10_26_328_0, i_10_26_394_0,
    i_10_26_429_0, i_10_26_444_0, i_10_26_445_0, i_10_26_447_0,
    i_10_26_448_0, i_10_26_465_0, i_10_26_792_0, i_10_26_798_0,
    i_10_26_799_0, i_10_26_955_0, i_10_26_1002_0, i_10_26_1032_0,
    i_10_26_1034_0, i_10_26_1240_0, i_10_26_1241_0, i_10_26_1265_0,
    i_10_26_1305_0, i_10_26_1306_0, i_10_26_1309_0, i_10_26_1651_0,
    i_10_26_1819_0, i_10_26_1821_0, i_10_26_1826_0, i_10_26_1911_0,
    i_10_26_1989_0, i_10_26_1995_0, i_10_26_1996_0, i_10_26_2311_0,
    i_10_26_2349_0, i_10_26_2351_0, i_10_26_2357_0, i_10_26_2364_0,
    i_10_26_2452_0, i_10_26_2571_0, i_10_26_2655_0, i_10_26_2656_0,
    i_10_26_2657_0, i_10_26_2658_0, i_10_26_2659_0, i_10_26_2703_0,
    i_10_26_2704_0, i_10_26_2714_0, i_10_26_2727_0, i_10_26_2728_0,
    i_10_26_2730_0, i_10_26_2731_0, i_10_26_2732_0, i_10_26_2787_0,
    i_10_26_2788_0, i_10_26_2819_0, i_10_26_2884_0, i_10_26_2985_0,
    i_10_26_2987_0, i_10_26_3039_0, i_10_26_3045_0, i_10_26_3046_0,
    i_10_26_3048_0, i_10_26_3049_0, i_10_26_3075_0, i_10_26_3076_0,
    i_10_26_3091_0, i_10_26_3094_0, i_10_26_3195_0, i_10_26_3198_0,
    i_10_26_3271_0, i_10_26_3272_0, i_10_26_3298_0, i_10_26_3326_0,
    i_10_26_3405_0, i_10_26_3407_0, i_10_26_3408_0, i_10_26_3409_0,
    i_10_26_3472_0, i_10_26_3613_0, i_10_26_3646_0, i_10_26_3855_0,
    i_10_26_3857_0, i_10_26_3860_0, i_10_26_3983_0, i_10_26_3985_0,
    i_10_26_3986_0, i_10_26_4115_0, i_10_26_4116_0, i_10_26_4117_0,
    i_10_26_4128_0, i_10_26_4216_0, i_10_26_4269_0, i_10_26_4270_0,
    i_10_26_4271_0, i_10_26_4278_0, i_10_26_4288_0, i_10_26_4568_0;
  output o_10_26_0_0;
  assign o_10_26_0_0 = ~((~i_10_26_2311_0 & ((~i_10_26_286_0 & ~i_10_26_326_0 & ((i_10_26_1651_0 & ~i_10_26_2658_0 & ~i_10_26_3048_0 & ~i_10_26_3195_0 & ~i_10_26_3407_0 & ~i_10_26_3855_0) | (~i_10_26_445_0 & ~i_10_26_1826_0 & ~i_10_26_2364_0 & i_10_26_2452_0 & i_10_26_3409_0 & ~i_10_26_4288_0))) | (~i_10_26_955_0 & ~i_10_26_3049_0 & ~i_10_26_4128_0 & ((~i_10_26_1240_0 & ~i_10_26_2659_0 & ~i_10_26_2819_0 & ~i_10_26_3094_0 & ~i_10_26_3198_0 & ~i_10_26_3405_0 & ~i_10_26_3986_0 & ~i_10_26_4216_0 & ~i_10_26_4271_0) | (~i_10_26_429_0 & ~i_10_26_792_0 & ~i_10_26_1265_0 & ~i_10_26_1651_0 & ~i_10_26_1821_0 & ~i_10_26_3046_0 & ~i_10_26_3091_0 & ~i_10_26_4288_0))) | (i_10_26_4117_0 & ((~i_10_26_1995_0 & ~i_10_26_1996_0 & ~i_10_26_2819_0 & ~i_10_26_3046_0 & ~i_10_26_3076_0 & ~i_10_26_3271_0 & ~i_10_26_3405_0 & ~i_10_26_3472_0) | (i_10_26_465_0 & ~i_10_26_1034_0 & i_10_26_2728_0 & ~i_10_26_3983_0 & ~i_10_26_4568_0))))) | (~i_10_26_1032_0 & ((~i_10_26_326_0 & ~i_10_26_3855_0 & ((~i_10_26_444_0 & i_10_26_1306_0 & ~i_10_26_1911_0 & ~i_10_26_2819_0 & ~i_10_26_3094_0 & ~i_10_26_2349_0 & ~i_10_26_2452_0) | (~i_10_26_394_0 & ~i_10_26_1240_0 & ~i_10_26_1241_0 & ~i_10_26_1989_0 & ~i_10_26_1996_0 & ~i_10_26_3405_0 & ~i_10_26_3646_0))) | (~i_10_26_394_0 & ~i_10_26_3048_0 & ~i_10_26_3983_0 & ((~i_10_26_1821_0 & i_10_26_1826_0 & ~i_10_26_1911_0 & ~i_10_26_1996_0 & ~i_10_26_2730_0 & ~i_10_26_3076_0 & ~i_10_26_4128_0) | (i_10_26_465_0 & ~i_10_26_2349_0 & ~i_10_26_2656_0 & ~i_10_26_3049_0 & ~i_10_26_3091_0 & ~i_10_26_4216_0))) | (~i_10_26_1002_0 & ~i_10_26_1821_0 & ~i_10_26_1996_0 & ~i_10_26_2656_0 & ~i_10_26_2703_0 & ~i_10_26_3075_0 & ~i_10_26_3091_0 & ~i_10_26_3272_0 & ~i_10_26_3405_0 & ~i_10_26_3985_0 & ~i_10_26_3986_0))) | (~i_10_26_3049_0 & ((~i_10_26_394_0 & ((~i_10_26_1309_0 & ~i_10_26_2351_0 & ~i_10_26_2364_0 & ~i_10_26_2658_0 & ~i_10_26_2728_0 & ~i_10_26_2819_0 & ~i_10_26_3091_0 & ~i_10_26_3646_0 & ~i_10_26_3857_0) | (i_10_26_2730_0 & i_10_26_2732_0 & ~i_10_26_3048_0 & ~i_10_26_3271_0 & ~i_10_26_3409_0 & ~i_10_26_3613_0 & ~i_10_26_3985_0))) | (~i_10_26_1911_0 & ((i_10_26_1309_0 & i_10_26_2357_0 & ~i_10_26_2788_0) | (~i_10_26_293_0 & ~i_10_26_444_0 & ~i_10_26_1821_0 & ~i_10_26_1989_0 & ~i_10_26_2349_0 & i_10_26_2732_0 & ~i_10_26_3048_0 & ~i_10_26_3075_0 & ~i_10_26_3094_0 & ~i_10_26_3195_0))) | (i_10_26_444_0 & i_10_26_1819_0 & ~i_10_26_2452_0 & ~i_10_26_2658_0) | (i_10_26_448_0 & ~i_10_26_2659_0 & ~i_10_26_3048_0 & ~i_10_26_4116_0) | (~i_10_26_2657_0 & ~i_10_26_2714_0 & i_10_26_3613_0 & ~i_10_26_3855_0 & ~i_10_26_3985_0 & ~i_10_26_4216_0 & ~i_10_26_4288_0))) | (~i_10_26_3409_0 & ((i_10_26_445_0 & ((~i_10_26_792_0 & i_10_26_2452_0 & i_10_26_3195_0 & ~i_10_26_3857_0) | (~i_10_26_955_0 & i_10_26_4117_0 & ~i_10_26_4288_0))) | (~i_10_26_3045_0 & ((~i_10_26_1241_0 & ~i_10_26_1306_0 & ~i_10_26_3075_0 & ~i_10_26_3076_0 & ~i_10_26_3407_0 & i_10_26_4116_0) | (i_10_26_465_0 & ~i_10_26_2357_0 & ~i_10_26_2788_0 & ~i_10_26_3405_0 & ~i_10_26_3985_0 & ~i_10_26_4117_0))))) | (~i_10_26_792_0 & ((i_10_26_1651_0 & ~i_10_26_3198_0 & i_10_26_3855_0 & ~i_10_26_4115_0 & i_10_26_4116_0) | (~i_10_26_328_0 & ~i_10_26_444_0 & ~i_10_26_2657_0 & ~i_10_26_2884_0 & ~i_10_26_3045_0 & ~i_10_26_3046_0 & ~i_10_26_3195_0 & ~i_10_26_3408_0 & ~i_10_26_3857_0 & ~i_10_26_4116_0 & ~i_10_26_4288_0))) | (~i_10_26_328_0 & ((~i_10_26_429_0 & ~i_10_26_1306_0 & ~i_10_26_1309_0 & i_10_26_1911_0 & ~i_10_26_3857_0) | (~i_10_26_1240_0 & ~i_10_26_1265_0 & i_10_26_1306_0 & ~i_10_26_1819_0 & ~i_10_26_1911_0 & ~i_10_26_3075_0 & ~i_10_26_3855_0 & ~i_10_26_3983_0 & ~i_10_26_4216_0))) | (~i_10_26_3076_0 & ((~i_10_26_429_0 & ~i_10_26_1996_0 & ~i_10_26_3195_0 & ((i_10_26_286_0 & ~i_10_26_1989_0 & ~i_10_26_2659_0 & ~i_10_26_3048_0 & ~i_10_26_3075_0 & ~i_10_26_3857_0 & ~i_10_26_4115_0) | (~i_10_26_1034_0 & ~i_10_26_2655_0 & ~i_10_26_2819_0 & ~i_10_26_3045_0 & ~i_10_26_3046_0 & ~i_10_26_3094_0 & ~i_10_26_4216_0))) | (i_10_26_2730_0 & ~i_10_26_3045_0 & ~i_10_26_3046_0 & ~i_10_26_3048_0 & ~i_10_26_3407_0 & ~i_10_26_3983_0) | (~i_10_26_3094_0 & ~i_10_26_3857_0 & i_10_26_4270_0))) | (i_10_26_2351_0 & ((~i_10_26_955_0 & i_10_26_1651_0 & ~i_10_26_2819_0 & ~i_10_26_3045_0) | (i_10_26_1265_0 & ~i_10_26_2349_0 & i_10_26_4117_0))) | (~i_10_26_2452_0 & ~i_10_26_2819_0 & ((i_10_26_1306_0 & ~i_10_26_1911_0 & i_10_26_3613_0 & i_10_26_3857_0 & ~i_10_26_3860_0) | (~i_10_26_296_0 & ~i_10_26_2658_0 & ~i_10_26_3046_0 & ~i_10_26_3048_0 & ~i_10_26_3094_0 & ~i_10_26_3195_0 & ~i_10_26_3646_0 & ~i_10_26_3986_0 & ~i_10_26_4117_0))) | (~i_10_26_3075_0 & ((~i_10_26_1265_0 & ~i_10_26_1309_0 & ~i_10_26_1996_0 & ~i_10_26_2571_0 & ~i_10_26_2655_0 & ~i_10_26_2788_0 & ~i_10_26_2884_0 & ~i_10_26_3091_0 & ~i_10_26_3405_0 & ~i_10_26_3408_0) | (~i_10_26_3048_0 & ~i_10_26_3271_0 & i_10_26_4278_0))) | (i_10_26_4288_0 & ((i_10_26_2657_0 & ~i_10_26_3271_0 & ~i_10_26_3405_0 & i_10_26_3613_0 & ~i_10_26_3986_0) | (i_10_26_3198_0 & ~i_10_26_3857_0 & i_10_26_4117_0))) | (i_10_26_1819_0 & i_10_26_2730_0 & i_10_26_2731_0 & ~i_10_26_3091_0 & ~i_10_26_3195_0 & ~i_10_26_3407_0));
endmodule



// Benchmark "kernel_10_27" written by ABC on Sun Jul 19 10:21:29 2020

module kernel_10_27 ( 
    i_10_27_40_0, i_10_27_229_0, i_10_27_230_0, i_10_27_271_0,
    i_10_27_272_0, i_10_27_319_0, i_10_27_423_0, i_10_27_427_0,
    i_10_27_430_0, i_10_27_433_0, i_10_27_449_0, i_10_27_464_0,
    i_10_27_543_0, i_10_27_741_0, i_10_27_751_0, i_10_27_877_0,
    i_10_27_1027_0, i_10_27_1054_0, i_10_27_1111_0, i_10_27_1252_0,
    i_10_27_1265_0, i_10_27_1311_0, i_10_27_1348_0, i_10_27_1354_0,
    i_10_27_1361_0, i_10_27_1364_0, i_10_27_1416_0, i_10_27_1492_0,
    i_10_27_1545_0, i_10_27_1552_0, i_10_27_1554_0, i_10_27_1579_0,
    i_10_27_1642_0, i_10_27_1650_0, i_10_27_1651_0, i_10_27_1652_0,
    i_10_27_1888_0, i_10_27_1909_0, i_10_27_1948_0, i_10_27_2161_0,
    i_10_27_2167_0, i_10_27_2168_0, i_10_27_2185_0, i_10_27_2186_0,
    i_10_27_2453_0, i_10_27_2458_0, i_10_27_2516_0, i_10_27_2641_0,
    i_10_27_2658_0, i_10_27_2663_0, i_10_27_2731_0, i_10_27_2732_0,
    i_10_27_2821_0, i_10_27_2865_0, i_10_27_2869_0, i_10_27_2885_0,
    i_10_27_2912_0, i_10_27_2917_0, i_10_27_2919_0, i_10_27_2924_0,
    i_10_27_2957_0, i_10_27_2983_0, i_10_27_3040_0, i_10_27_3201_0,
    i_10_27_3203_0, i_10_27_3270_0, i_10_27_3307_0, i_10_27_3325_0,
    i_10_27_3469_0, i_10_27_3472_0, i_10_27_3521_0, i_10_27_3523_0,
    i_10_27_3526_0, i_10_27_3540_0, i_10_27_3541_0, i_10_27_3544_0,
    i_10_27_3614_0, i_10_27_3718_0, i_10_27_3781_0, i_10_27_3786_0,
    i_10_27_3828_0, i_10_27_3852_0, i_10_27_3890_0, i_10_27_3910_0,
    i_10_27_3947_0, i_10_27_3988_0, i_10_27_3990_0, i_10_27_4008_0,
    i_10_27_4013_0, i_10_27_4054_0, i_10_27_4116_0, i_10_27_4117_0,
    i_10_27_4149_0, i_10_27_4152_0, i_10_27_4154_0, i_10_27_4190_0,
    i_10_27_4272_0, i_10_27_4285_0, i_10_27_4570_0, i_10_27_4595_0,
    o_10_27_0_0  );
  input  i_10_27_40_0, i_10_27_229_0, i_10_27_230_0, i_10_27_271_0,
    i_10_27_272_0, i_10_27_319_0, i_10_27_423_0, i_10_27_427_0,
    i_10_27_430_0, i_10_27_433_0, i_10_27_449_0, i_10_27_464_0,
    i_10_27_543_0, i_10_27_741_0, i_10_27_751_0, i_10_27_877_0,
    i_10_27_1027_0, i_10_27_1054_0, i_10_27_1111_0, i_10_27_1252_0,
    i_10_27_1265_0, i_10_27_1311_0, i_10_27_1348_0, i_10_27_1354_0,
    i_10_27_1361_0, i_10_27_1364_0, i_10_27_1416_0, i_10_27_1492_0,
    i_10_27_1545_0, i_10_27_1552_0, i_10_27_1554_0, i_10_27_1579_0,
    i_10_27_1642_0, i_10_27_1650_0, i_10_27_1651_0, i_10_27_1652_0,
    i_10_27_1888_0, i_10_27_1909_0, i_10_27_1948_0, i_10_27_2161_0,
    i_10_27_2167_0, i_10_27_2168_0, i_10_27_2185_0, i_10_27_2186_0,
    i_10_27_2453_0, i_10_27_2458_0, i_10_27_2516_0, i_10_27_2641_0,
    i_10_27_2658_0, i_10_27_2663_0, i_10_27_2731_0, i_10_27_2732_0,
    i_10_27_2821_0, i_10_27_2865_0, i_10_27_2869_0, i_10_27_2885_0,
    i_10_27_2912_0, i_10_27_2917_0, i_10_27_2919_0, i_10_27_2924_0,
    i_10_27_2957_0, i_10_27_2983_0, i_10_27_3040_0, i_10_27_3201_0,
    i_10_27_3203_0, i_10_27_3270_0, i_10_27_3307_0, i_10_27_3325_0,
    i_10_27_3469_0, i_10_27_3472_0, i_10_27_3521_0, i_10_27_3523_0,
    i_10_27_3526_0, i_10_27_3540_0, i_10_27_3541_0, i_10_27_3544_0,
    i_10_27_3614_0, i_10_27_3718_0, i_10_27_3781_0, i_10_27_3786_0,
    i_10_27_3828_0, i_10_27_3852_0, i_10_27_3890_0, i_10_27_3910_0,
    i_10_27_3947_0, i_10_27_3988_0, i_10_27_3990_0, i_10_27_4008_0,
    i_10_27_4013_0, i_10_27_4054_0, i_10_27_4116_0, i_10_27_4117_0,
    i_10_27_4149_0, i_10_27_4152_0, i_10_27_4154_0, i_10_27_4190_0,
    i_10_27_4272_0, i_10_27_4285_0, i_10_27_4570_0, i_10_27_4595_0;
  output o_10_27_0_0;
  assign o_10_27_0_0 = 0;
endmodule



// Benchmark "kernel_10_28" written by ABC on Sun Jul 19 10:21:31 2020

module kernel_10_28 ( 
    i_10_28_89_0, i_10_28_171_0, i_10_28_221_0, i_10_28_222_0,
    i_10_28_223_0, i_10_28_224_0, i_10_28_285_0, i_10_28_287_0,
    i_10_28_318_0, i_10_28_319_0, i_10_28_323_0, i_10_28_432_0,
    i_10_28_433_0, i_10_28_444_0, i_10_28_445_0, i_10_28_446_0,
    i_10_28_449_0, i_10_28_506_0, i_10_28_719_0, i_10_28_752_0,
    i_10_28_795_0, i_10_28_1037_0, i_10_28_1236_0, i_10_28_1238_0,
    i_10_28_1242_0, i_10_28_1243_0, i_10_28_1244_0, i_10_28_1246_0,
    i_10_28_1647_0, i_10_28_1650_0, i_10_28_1651_0, i_10_28_1652_0,
    i_10_28_1653_0, i_10_28_1819_0, i_10_28_1821_0, i_10_28_1824_0,
    i_10_28_1825_0, i_10_28_1989_0, i_10_28_2338_0, i_10_28_2359_0,
    i_10_28_2362_0, i_10_28_2467_0, i_10_28_2468_0, i_10_28_2629_0,
    i_10_28_2631_0, i_10_28_2633_0, i_10_28_2635_0, i_10_28_2645_0,
    i_10_28_2657_0, i_10_28_2658_0, i_10_28_2659_0, i_10_28_2660_0,
    i_10_28_2678_0, i_10_28_2720_0, i_10_28_2785_0, i_10_28_2788_0,
    i_10_28_2821_0, i_10_28_2888_0, i_10_28_2919_0, i_10_28_2920_0,
    i_10_28_2922_0, i_10_28_2924_0, i_10_28_2981_0, i_10_28_3033_0,
    i_10_28_3034_0, i_10_28_3150_0, i_10_28_3151_0, i_10_28_3152_0,
    i_10_28_3154_0, i_10_28_3155_0, i_10_28_3156_0, i_10_28_3157_0,
    i_10_28_3195_0, i_10_28_3274_0, i_10_28_3278_0, i_10_28_3385_0,
    i_10_28_3408_0, i_10_28_3587_0, i_10_28_3685_0, i_10_28_3780_0,
    i_10_28_3782_0, i_10_28_3788_0, i_10_28_3834_0, i_10_28_3835_0,
    i_10_28_3836_0, i_10_28_3839_0, i_10_28_3847_0, i_10_28_3848_0,
    i_10_28_3853_0, i_10_28_3854_0, i_10_28_3856_0, i_10_28_3857_0,
    i_10_28_3860_0, i_10_28_4116_0, i_10_28_4129_0, i_10_28_4565_0,
    i_10_28_4567_0, i_10_28_4568_0, i_10_28_4570_0, i_10_28_4571_0,
    o_10_28_0_0  );
  input  i_10_28_89_0, i_10_28_171_0, i_10_28_221_0, i_10_28_222_0,
    i_10_28_223_0, i_10_28_224_0, i_10_28_285_0, i_10_28_287_0,
    i_10_28_318_0, i_10_28_319_0, i_10_28_323_0, i_10_28_432_0,
    i_10_28_433_0, i_10_28_444_0, i_10_28_445_0, i_10_28_446_0,
    i_10_28_449_0, i_10_28_506_0, i_10_28_719_0, i_10_28_752_0,
    i_10_28_795_0, i_10_28_1037_0, i_10_28_1236_0, i_10_28_1238_0,
    i_10_28_1242_0, i_10_28_1243_0, i_10_28_1244_0, i_10_28_1246_0,
    i_10_28_1647_0, i_10_28_1650_0, i_10_28_1651_0, i_10_28_1652_0,
    i_10_28_1653_0, i_10_28_1819_0, i_10_28_1821_0, i_10_28_1824_0,
    i_10_28_1825_0, i_10_28_1989_0, i_10_28_2338_0, i_10_28_2359_0,
    i_10_28_2362_0, i_10_28_2467_0, i_10_28_2468_0, i_10_28_2629_0,
    i_10_28_2631_0, i_10_28_2633_0, i_10_28_2635_0, i_10_28_2645_0,
    i_10_28_2657_0, i_10_28_2658_0, i_10_28_2659_0, i_10_28_2660_0,
    i_10_28_2678_0, i_10_28_2720_0, i_10_28_2785_0, i_10_28_2788_0,
    i_10_28_2821_0, i_10_28_2888_0, i_10_28_2919_0, i_10_28_2920_0,
    i_10_28_2922_0, i_10_28_2924_0, i_10_28_2981_0, i_10_28_3033_0,
    i_10_28_3034_0, i_10_28_3150_0, i_10_28_3151_0, i_10_28_3152_0,
    i_10_28_3154_0, i_10_28_3155_0, i_10_28_3156_0, i_10_28_3157_0,
    i_10_28_3195_0, i_10_28_3274_0, i_10_28_3278_0, i_10_28_3385_0,
    i_10_28_3408_0, i_10_28_3587_0, i_10_28_3685_0, i_10_28_3780_0,
    i_10_28_3782_0, i_10_28_3788_0, i_10_28_3834_0, i_10_28_3835_0,
    i_10_28_3836_0, i_10_28_3839_0, i_10_28_3847_0, i_10_28_3848_0,
    i_10_28_3853_0, i_10_28_3854_0, i_10_28_3856_0, i_10_28_3857_0,
    i_10_28_3860_0, i_10_28_4116_0, i_10_28_4129_0, i_10_28_4565_0,
    i_10_28_4567_0, i_10_28_4568_0, i_10_28_4570_0, i_10_28_4571_0;
  output o_10_28_0_0;
  assign o_10_28_0_0 = ~((~i_10_28_222_0 & ((~i_10_28_2919_0 & ~i_10_28_3034_0 & ~i_10_28_3788_0 & ~i_10_28_3856_0 & ~i_10_28_3860_0 & i_10_28_4116_0) | (~i_10_28_433_0 & ~i_10_28_752_0 & i_10_28_2660_0 & ~i_10_28_2678_0 & ~i_10_28_2924_0 & ~i_10_28_3834_0 & ~i_10_28_3839_0 & ~i_10_28_4567_0))) | (i_10_28_445_0 & ((~i_10_28_2629_0 & ~i_10_28_2631_0 & ~i_10_28_2633_0 & ~i_10_28_2922_0 & ~i_10_28_2924_0 & ~i_10_28_3033_0 & ~i_10_28_3782_0) | (~i_10_28_795_0 & ~i_10_28_1244_0 & ~i_10_28_1653_0 & ~i_10_28_3034_0 & ~i_10_28_3385_0 & ~i_10_28_3836_0 & ~i_10_28_3839_0 & ~i_10_28_3848_0))) | (~i_10_28_719_0 & ((~i_10_28_1246_0 & ~i_10_28_2359_0 & ~i_10_28_2633_0 & ~i_10_28_2919_0 & ~i_10_28_2920_0 & ~i_10_28_3685_0 & ~i_10_28_3839_0 & ~i_10_28_3857_0) | (~i_10_28_1037_0 & ~i_10_28_1243_0 & ~i_10_28_1647_0 & ~i_10_28_2635_0 & ~i_10_28_2924_0 & ~i_10_28_3780_0 & ~i_10_28_3860_0))) | (~i_10_28_1037_0 & ((~i_10_28_287_0 & ~i_10_28_1238_0 & ~i_10_28_1242_0 & ~i_10_28_2922_0 & ~i_10_28_3274_0 & i_10_28_3835_0) | (~i_10_28_89_0 & ~i_10_28_1647_0 & ~i_10_28_1653_0 & ~i_10_28_2359_0 & ~i_10_28_2645_0 & ~i_10_28_3195_0 & ~i_10_28_4567_0 & ~i_10_28_4570_0 & ~i_10_28_4571_0))) | (~i_10_28_3857_0 & ((~i_10_28_3848_0 & ((~i_10_28_221_0 & ~i_10_28_2919_0 & ((~i_10_28_1238_0 & ~i_10_28_1650_0 & ~i_10_28_2629_0 & ~i_10_28_3839_0 & ~i_10_28_4565_0) | (~i_10_28_1236_0 & ~i_10_28_1243_0 & ~i_10_28_2645_0 & ~i_10_28_2920_0 & ~i_10_28_3195_0 & ~i_10_28_3685_0 & ~i_10_28_3854_0 & ~i_10_28_4567_0))) | (~i_10_28_1653_0 & ~i_10_28_1824_0 & ~i_10_28_1825_0 & ~i_10_28_2362_0 & ~i_10_28_2660_0 & ~i_10_28_3034_0 & ~i_10_28_3780_0 & ~i_10_28_3839_0))) | (~i_10_28_446_0 & ~i_10_28_752_0 & ~i_10_28_1236_0 & ~i_10_28_1244_0 & ~i_10_28_3033_0 & ~i_10_28_3274_0 & ~i_10_28_3685_0 & ~i_10_28_3780_0))) | (~i_10_28_1244_0 & ((~i_10_28_221_0 & ((~i_10_28_752_0 & ~i_10_28_1651_0 & ~i_10_28_2660_0 & ~i_10_28_2922_0 & ~i_10_28_3834_0 & ~i_10_28_3839_0 & ~i_10_28_4116_0) | (~i_10_28_224_0 & ~i_10_28_1243_0 & ~i_10_28_1647_0 & ~i_10_28_1653_0 & ~i_10_28_3274_0 & ~i_10_28_4565_0))) | (~i_10_28_224_0 & ((~i_10_28_752_0 & ~i_10_28_1647_0 & ~i_10_28_1821_0 & ~i_10_28_1989_0 & ~i_10_28_2338_0 & ~i_10_28_2924_0 & ~i_10_28_3780_0) | (i_10_28_1819_0 & ~i_10_28_2362_0 & ~i_10_28_2629_0 & ~i_10_28_3854_0 & ~i_10_28_4570_0))) | (~i_10_28_2645_0 & ((~i_10_28_1242_0 & ~i_10_28_1246_0 & ~i_10_28_2338_0 & ~i_10_28_2631_0 & ~i_10_28_2981_0 & ~i_10_28_3788_0 & i_10_28_4567_0) | (~i_10_28_223_0 & ~i_10_28_1243_0 & ~i_10_28_2924_0 & ~i_10_28_4565_0 & ~i_10_28_4568_0))) | (i_10_28_2468_0 & ~i_10_28_3033_0 & ~i_10_28_3853_0))) | (~i_10_28_2629_0 & ((i_10_28_3587_0 & ~i_10_28_3860_0) | (i_10_28_2678_0 & ~i_10_28_4129_0))) | (~i_10_28_3034_0 & ((i_10_28_1825_0 & ~i_10_28_2338_0 & i_10_28_3835_0 & ~i_10_28_3854_0) | (i_10_28_171_0 & ~i_10_28_1238_0 & ~i_10_28_2359_0 & ~i_10_28_2924_0 & i_10_28_3856_0 & ~i_10_28_4116_0))) | (~i_10_28_2924_0 & ((i_10_28_2659_0 & ~i_10_28_2920_0 & ~i_10_28_2981_0 & ~i_10_28_3788_0 & ~i_10_28_3848_0) | (i_10_28_795_0 & ~i_10_28_1652_0 & ~i_10_28_2720_0 & ~i_10_28_3033_0 & ~i_10_28_3839_0 & i_10_28_4565_0))) | (~i_10_28_3274_0 & ((~i_10_28_1652_0 & ((~i_10_28_1651_0 & i_10_28_1653_0 & ~i_10_28_2362_0 & ~i_10_28_3848_0) | (~i_10_28_2633_0 & i_10_28_3848_0 & ~i_10_28_3860_0 & ~i_10_28_4565_0))) | (~i_10_28_224_0 & ~i_10_28_445_0 & ~i_10_28_1246_0 & ~i_10_28_2645_0 & ~i_10_28_3385_0 & ~i_10_28_3780_0 & ~i_10_28_3782_0 & ~i_10_28_3848_0 & ~i_10_28_4565_0))) | (~i_10_28_1650_0 & i_10_28_2981_0 & i_10_28_3839_0) | (i_10_28_2678_0 & ~i_10_28_3782_0 & ~i_10_28_3856_0 & ~i_10_28_4567_0));
endmodule



// Benchmark "kernel_10_29" written by ABC on Sun Jul 19 10:21:32 2020

module kernel_10_29 ( 
    i_10_29_174_0, i_10_29_179_0, i_10_29_223_0, i_10_29_243_0,
    i_10_29_256_0, i_10_29_257_0, i_10_29_286_0, i_10_29_318_0,
    i_10_29_319_0, i_10_29_321_0, i_10_29_323_0, i_10_29_387_0,
    i_10_29_435_0, i_10_29_436_0, i_10_29_443_0, i_10_29_447_0,
    i_10_29_561_0, i_10_29_907_0, i_10_29_997_0, i_10_29_1003_0,
    i_10_29_1004_0, i_10_29_1040_0, i_10_29_1042_0, i_10_29_1043_0,
    i_10_29_1263_0, i_10_29_1308_0, i_10_29_1344_0, i_10_29_1347_0,
    i_10_29_1435_0, i_10_29_1444_0, i_10_29_1542_0, i_10_29_1543_0,
    i_10_29_1544_0, i_10_29_1576_0, i_10_29_1578_0, i_10_29_1579_0,
    i_10_29_1580_0, i_10_29_1582_0, i_10_29_1611_0, i_10_29_1636_0,
    i_10_29_1654_0, i_10_29_1689_0, i_10_29_1691_0, i_10_29_1768_0,
    i_10_29_1816_0, i_10_29_1821_0, i_10_29_1822_0, i_10_29_1913_0,
    i_10_29_1956_0, i_10_29_1984_0, i_10_29_2003_0, i_10_29_2019_0,
    i_10_29_2083_0, i_10_29_2291_0, i_10_29_2436_0, i_10_29_2451_0,
    i_10_29_2453_0, i_10_29_2514_0, i_10_29_2515_0, i_10_29_2631_0,
    i_10_29_2656_0, i_10_29_2703_0, i_10_29_2704_0, i_10_29_2716_0,
    i_10_29_2826_0, i_10_29_2882_0, i_10_29_2920_0, i_10_29_2960_0,
    i_10_29_3036_0, i_10_29_3277_0, i_10_29_3289_0, i_10_29_3298_0,
    i_10_29_3431_0, i_10_29_3473_0, i_10_29_3541_0, i_10_29_3544_0,
    i_10_29_3614_0, i_10_29_3649_0, i_10_29_3729_0, i_10_29_3784_0,
    i_10_29_3786_0, i_10_29_3787_0, i_10_29_3837_0, i_10_29_3848_0,
    i_10_29_3856_0, i_10_29_3912_0, i_10_29_3946_0, i_10_29_3982_0,
    i_10_29_4114_0, i_10_29_4115_0, i_10_29_4171_0, i_10_29_4172_0,
    i_10_29_4175_0, i_10_29_4233_0, i_10_29_4234_0, i_10_29_4279_0,
    i_10_29_4459_0, i_10_29_4462_0, i_10_29_4568_0, i_10_29_4571_0,
    o_10_29_0_0  );
  input  i_10_29_174_0, i_10_29_179_0, i_10_29_223_0, i_10_29_243_0,
    i_10_29_256_0, i_10_29_257_0, i_10_29_286_0, i_10_29_318_0,
    i_10_29_319_0, i_10_29_321_0, i_10_29_323_0, i_10_29_387_0,
    i_10_29_435_0, i_10_29_436_0, i_10_29_443_0, i_10_29_447_0,
    i_10_29_561_0, i_10_29_907_0, i_10_29_997_0, i_10_29_1003_0,
    i_10_29_1004_0, i_10_29_1040_0, i_10_29_1042_0, i_10_29_1043_0,
    i_10_29_1263_0, i_10_29_1308_0, i_10_29_1344_0, i_10_29_1347_0,
    i_10_29_1435_0, i_10_29_1444_0, i_10_29_1542_0, i_10_29_1543_0,
    i_10_29_1544_0, i_10_29_1576_0, i_10_29_1578_0, i_10_29_1579_0,
    i_10_29_1580_0, i_10_29_1582_0, i_10_29_1611_0, i_10_29_1636_0,
    i_10_29_1654_0, i_10_29_1689_0, i_10_29_1691_0, i_10_29_1768_0,
    i_10_29_1816_0, i_10_29_1821_0, i_10_29_1822_0, i_10_29_1913_0,
    i_10_29_1956_0, i_10_29_1984_0, i_10_29_2003_0, i_10_29_2019_0,
    i_10_29_2083_0, i_10_29_2291_0, i_10_29_2436_0, i_10_29_2451_0,
    i_10_29_2453_0, i_10_29_2514_0, i_10_29_2515_0, i_10_29_2631_0,
    i_10_29_2656_0, i_10_29_2703_0, i_10_29_2704_0, i_10_29_2716_0,
    i_10_29_2826_0, i_10_29_2882_0, i_10_29_2920_0, i_10_29_2960_0,
    i_10_29_3036_0, i_10_29_3277_0, i_10_29_3289_0, i_10_29_3298_0,
    i_10_29_3431_0, i_10_29_3473_0, i_10_29_3541_0, i_10_29_3544_0,
    i_10_29_3614_0, i_10_29_3649_0, i_10_29_3729_0, i_10_29_3784_0,
    i_10_29_3786_0, i_10_29_3787_0, i_10_29_3837_0, i_10_29_3848_0,
    i_10_29_3856_0, i_10_29_3912_0, i_10_29_3946_0, i_10_29_3982_0,
    i_10_29_4114_0, i_10_29_4115_0, i_10_29_4171_0, i_10_29_4172_0,
    i_10_29_4175_0, i_10_29_4233_0, i_10_29_4234_0, i_10_29_4279_0,
    i_10_29_4459_0, i_10_29_4462_0, i_10_29_4568_0, i_10_29_4571_0;
  output o_10_29_0_0;
  assign o_10_29_0_0 = 0;
endmodule



// Benchmark "kernel_10_30" written by ABC on Sun Jul 19 10:21:33 2020

module kernel_10_30 ( 
    i_10_30_86_0, i_10_30_88_0, i_10_30_89_0, i_10_30_280_0, i_10_30_284_0,
    i_10_30_330_0, i_10_30_393_0, i_10_30_394_0, i_10_30_395_0,
    i_10_30_413_0, i_10_30_431_0, i_10_30_437_0, i_10_30_459_0,
    i_10_30_462_0, i_10_30_463_0, i_10_30_464_0, i_10_30_700_0,
    i_10_30_996_0, i_10_30_1033_0, i_10_30_1039_0, i_10_30_1041_0,
    i_10_30_1168_0, i_10_30_1237_0, i_10_30_1245_0, i_10_30_1246_0,
    i_10_30_1247_0, i_10_30_1248_0, i_10_30_1249_0, i_10_30_1250_0,
    i_10_30_1313_0, i_10_30_1367_0, i_10_30_1384_0, i_10_30_1385_0,
    i_10_30_1582_0, i_10_30_1649_0, i_10_30_1716_0, i_10_30_1717_0,
    i_10_30_1735_0, i_10_30_1768_0, i_10_30_1769_0, i_10_30_1823_0,
    i_10_30_1912_0, i_10_30_1913_0, i_10_30_2005_0, i_10_30_2006_0,
    i_10_30_2201_0, i_10_30_2350_0, i_10_30_2354_0, i_10_30_2355_0,
    i_10_30_2356_0, i_10_30_2357_0, i_10_30_2361_0, i_10_30_2383_0,
    i_10_30_2438_0, i_10_30_2449_0, i_10_30_2451_0, i_10_30_2452_0,
    i_10_30_2455_0, i_10_30_2456_0, i_10_30_2516_0, i_10_30_2653_0,
    i_10_30_2681_0, i_10_30_2728_0, i_10_30_2918_0, i_10_30_2920_0,
    i_10_30_3041_0, i_10_30_3043_0, i_10_30_3076_0, i_10_30_3094_0,
    i_10_30_3200_0, i_10_30_3270_0, i_10_30_3280_0, i_10_30_3386_0,
    i_10_30_3387_0, i_10_30_3544_0, i_10_30_3611_0, i_10_30_3612_0,
    i_10_30_3613_0, i_10_30_3614_0, i_10_30_3615_0, i_10_30_3617_0,
    i_10_30_3781_0, i_10_30_3783_0, i_10_30_3787_0, i_10_30_3788_0,
    i_10_30_3836_0, i_10_30_3837_0, i_10_30_3838_0, i_10_30_3839_0,
    i_10_30_3846_0, i_10_30_3855_0, i_10_30_3856_0, i_10_30_3857_0,
    i_10_30_3886_0, i_10_30_3887_0, i_10_30_4120_0, i_10_30_4130_0,
    i_10_30_4219_0, i_10_30_4291_0, i_10_30_4292_0,
    o_10_30_0_0  );
  input  i_10_30_86_0, i_10_30_88_0, i_10_30_89_0, i_10_30_280_0,
    i_10_30_284_0, i_10_30_330_0, i_10_30_393_0, i_10_30_394_0,
    i_10_30_395_0, i_10_30_413_0, i_10_30_431_0, i_10_30_437_0,
    i_10_30_459_0, i_10_30_462_0, i_10_30_463_0, i_10_30_464_0,
    i_10_30_700_0, i_10_30_996_0, i_10_30_1033_0, i_10_30_1039_0,
    i_10_30_1041_0, i_10_30_1168_0, i_10_30_1237_0, i_10_30_1245_0,
    i_10_30_1246_0, i_10_30_1247_0, i_10_30_1248_0, i_10_30_1249_0,
    i_10_30_1250_0, i_10_30_1313_0, i_10_30_1367_0, i_10_30_1384_0,
    i_10_30_1385_0, i_10_30_1582_0, i_10_30_1649_0, i_10_30_1716_0,
    i_10_30_1717_0, i_10_30_1735_0, i_10_30_1768_0, i_10_30_1769_0,
    i_10_30_1823_0, i_10_30_1912_0, i_10_30_1913_0, i_10_30_2005_0,
    i_10_30_2006_0, i_10_30_2201_0, i_10_30_2350_0, i_10_30_2354_0,
    i_10_30_2355_0, i_10_30_2356_0, i_10_30_2357_0, i_10_30_2361_0,
    i_10_30_2383_0, i_10_30_2438_0, i_10_30_2449_0, i_10_30_2451_0,
    i_10_30_2452_0, i_10_30_2455_0, i_10_30_2456_0, i_10_30_2516_0,
    i_10_30_2653_0, i_10_30_2681_0, i_10_30_2728_0, i_10_30_2918_0,
    i_10_30_2920_0, i_10_30_3041_0, i_10_30_3043_0, i_10_30_3076_0,
    i_10_30_3094_0, i_10_30_3200_0, i_10_30_3270_0, i_10_30_3280_0,
    i_10_30_3386_0, i_10_30_3387_0, i_10_30_3544_0, i_10_30_3611_0,
    i_10_30_3612_0, i_10_30_3613_0, i_10_30_3614_0, i_10_30_3615_0,
    i_10_30_3617_0, i_10_30_3781_0, i_10_30_3783_0, i_10_30_3787_0,
    i_10_30_3788_0, i_10_30_3836_0, i_10_30_3837_0, i_10_30_3838_0,
    i_10_30_3839_0, i_10_30_3846_0, i_10_30_3855_0, i_10_30_3856_0,
    i_10_30_3857_0, i_10_30_3886_0, i_10_30_3887_0, i_10_30_4120_0,
    i_10_30_4130_0, i_10_30_4219_0, i_10_30_4291_0, i_10_30_4292_0;
  output o_10_30_0_0;
  assign o_10_30_0_0 = ~((~i_10_30_3200_0 & ((~i_10_30_393_0 & ~i_10_30_2006_0 & ~i_10_30_2456_0 & ((~i_10_30_996_0 & ~i_10_30_1041_0 & ~i_10_30_1250_0 & ~i_10_30_3611_0 & ~i_10_30_3836_0) | (~i_10_30_1039_0 & ~i_10_30_3837_0 & ~i_10_30_4292_0))) | (~i_10_30_394_0 & ((~i_10_30_86_0 & i_10_30_463_0 & ~i_10_30_1248_0 & ~i_10_30_1250_0 & ~i_10_30_1313_0 & ~i_10_30_3839_0) | (~i_10_30_89_0 & ~i_10_30_1041_0 & ~i_10_30_1249_0 & ~i_10_30_1913_0 & ~i_10_30_2681_0 & ~i_10_30_3857_0))) | (~i_10_30_462_0 & ~i_10_30_463_0 & ~i_10_30_700_0 & ~i_10_30_3617_0 & ~i_10_30_3783_0) | (~i_10_30_88_0 & i_10_30_464_0 & i_10_30_3280_0 & ~i_10_30_3386_0 & ~i_10_30_3615_0 & i_10_30_4120_0))) | (~i_10_30_1367_0 & ((~i_10_30_393_0 & ~i_10_30_395_0 & ((~i_10_30_89_0 & ~i_10_30_1768_0 & ~i_10_30_1769_0 & ~i_10_30_2005_0 & ~i_10_30_2452_0 & i_10_30_2456_0 & ~i_10_30_3611_0) | (~i_10_30_1245_0 & ~i_10_30_2920_0 & ~i_10_30_3781_0 & ~i_10_30_3839_0 & ~i_10_30_4292_0))) | (i_10_30_1249_0 & ((~i_10_30_996_0 & ~i_10_30_2006_0 & ~i_10_30_2201_0 & ~i_10_30_3836_0 & ~i_10_30_3837_0 & ~i_10_30_4130_0) | (~i_10_30_1168_0 & ~i_10_30_2449_0 & i_10_30_2452_0 & ~i_10_30_3617_0 & ~i_10_30_4219_0))) | (~i_10_30_1168_0 & ~i_10_30_3270_0 & ~i_10_30_3613_0 & ((~i_10_30_431_0 & ~i_10_30_3837_0) | (~i_10_30_437_0 & ~i_10_30_1735_0 & ~i_10_30_2361_0 & ~i_10_30_2449_0 & ~i_10_30_3544_0 & ~i_10_30_3612_0 & ~i_10_30_3783_0 & ~i_10_30_3846_0))) | (~i_10_30_462_0 & i_10_30_463_0 & ~i_10_30_3386_0 & i_10_30_3781_0 & ~i_10_30_3837_0))) | (~i_10_30_89_0 & ((~i_10_30_462_0 & ~i_10_30_463_0 & ~i_10_30_700_0 & ~i_10_30_1913_0 & ~i_10_30_2005_0 & ~i_10_30_2006_0 & ~i_10_30_3781_0) | (~i_10_30_395_0 & ~i_10_30_1168_0 & ~i_10_30_1649_0 & ~i_10_30_2383_0 & ~i_10_30_2456_0 & ~i_10_30_3041_0 & ~i_10_30_3611_0 & ~i_10_30_3615_0 & ~i_10_30_3617_0 & ~i_10_30_3855_0 & ~i_10_30_3856_0))) | (~i_10_30_1039_0 & ((~i_10_30_413_0 & ~i_10_30_437_0 & ~i_10_30_996_0 & ~i_10_30_1168_0 & ~i_10_30_1735_0 & ~i_10_30_2918_0 & ~i_10_30_3837_0 & ~i_10_30_3838_0) | (~i_10_30_462_0 & ~i_10_30_1250_0 & ~i_10_30_2456_0 & ~i_10_30_3094_0 & ~i_10_30_3783_0 & ~i_10_30_3839_0))) | (~i_10_30_437_0 & ((~i_10_30_462_0 & ~i_10_30_464_0 & ~i_10_30_700_0 & i_10_30_1313_0) | (~i_10_30_1246_0 & ~i_10_30_1735_0 & ~i_10_30_1768_0 & ~i_10_30_2681_0 & ~i_10_30_3094_0 & ~i_10_30_3614_0 & ~i_10_30_3617_0 & ~i_10_30_4130_0))) | (~i_10_30_464_0 & ~i_10_30_3837_0 & ((~i_10_30_88_0 & ~i_10_30_1823_0 & ~i_10_30_3614_0) | (i_10_30_2456_0 & i_10_30_4120_0))) | (~i_10_30_3094_0 & ((~i_10_30_88_0 & ((i_10_30_2452_0 & i_10_30_2455_0 & ~i_10_30_2728_0 & ~i_10_30_3386_0 & ~i_10_30_3617_0 & ~i_10_30_3846_0 & ~i_10_30_4130_0) | (i_10_30_462_0 & ~i_10_30_996_0 & ~i_10_30_2005_0 & ~i_10_30_2006_0 & ~i_10_30_2201_0 & ~i_10_30_2449_0 & ~i_10_30_3783_0 & ~i_10_30_4292_0))) | (~i_10_30_996_0 & ~i_10_30_1735_0 & ~i_10_30_2449_0 & ~i_10_30_3617_0 & ~i_10_30_3783_0 & i_10_30_2728_0 & ~i_10_30_3041_0) | (~i_10_30_1250_0 & ~i_10_30_2455_0 & i_10_30_3787_0 & ~i_10_30_4292_0) | (~i_10_30_284_0 & i_10_30_1033_0 & ~i_10_30_2681_0 & ~i_10_30_2920_0 & ~i_10_30_3836_0))) | (~i_10_30_1246_0 & i_10_30_1649_0 & i_10_30_2350_0) | (~i_10_30_462_0 & i_10_30_1246_0 & ~i_10_30_1823_0 & i_10_30_3836_0 & ~i_10_30_4130_0));
endmodule



// Benchmark "kernel_10_31" written by ABC on Sun Jul 19 10:21:34 2020

module kernel_10_31 ( 
    i_10_31_32_0, i_10_31_88_0, i_10_31_133_0, i_10_31_151_0,
    i_10_31_266_0, i_10_31_349_0, i_10_31_364_0, i_10_31_393_0,
    i_10_31_394_0, i_10_31_431_0, i_10_31_464_0, i_10_31_465_0,
    i_10_31_466_0, i_10_31_566_0, i_10_31_591_0, i_10_31_592_0,
    i_10_31_673_0, i_10_31_674_0, i_10_31_750_0, i_10_31_754_0,
    i_10_31_770_0, i_10_31_798_0, i_10_31_952_0, i_10_31_953_0,
    i_10_31_976_0, i_10_31_996_0, i_10_31_1033_0, i_10_31_1052_0,
    i_10_31_1059_0, i_10_31_1235_0, i_10_31_1236_0, i_10_31_1238_0,
    i_10_31_1241_0, i_10_31_1312_0, i_10_31_1358_0, i_10_31_1382_0,
    i_10_31_1457_0, i_10_31_1491_0, i_10_31_1619_0, i_10_31_1822_0,
    i_10_31_1867_0, i_10_31_1906_0, i_10_31_1912_0, i_10_31_1913_0,
    i_10_31_1914_0, i_10_31_1952_0, i_10_31_1957_0, i_10_31_1958_0,
    i_10_31_1960_0, i_10_31_1987_0, i_10_31_2095_0, i_10_31_2275_0,
    i_10_31_2276_0, i_10_31_2362_0, i_10_31_2465_0, i_10_31_2481_0,
    i_10_31_2508_0, i_10_31_2516_0, i_10_31_2572_0, i_10_31_2644_0,
    i_10_31_2661_0, i_10_31_2662_0, i_10_31_2678_0, i_10_31_2712_0,
    i_10_31_2744_0, i_10_31_2782_0, i_10_31_2786_0, i_10_31_2914_0,
    i_10_31_2916_0, i_10_31_2948_0, i_10_31_2956_0, i_10_31_2960_0,
    i_10_31_3093_0, i_10_31_3175_0, i_10_31_3176_0, i_10_31_3198_0,
    i_10_31_3199_0, i_10_31_3362_0, i_10_31_3446_0, i_10_31_3451_0,
    i_10_31_3470_0, i_10_31_3472_0, i_10_31_3473_0, i_10_31_3495_0,
    i_10_31_3508_0, i_10_31_3614_0, i_10_31_3622_0, i_10_31_3642_0,
    i_10_31_3643_0, i_10_31_3649_0, i_10_31_3652_0, i_10_31_3858_0,
    i_10_31_3860_0, i_10_31_3885_0, i_10_31_4056_0, i_10_31_4057_0,
    i_10_31_4058_0, i_10_31_4129_0, i_10_31_4287_0, i_10_31_4526_0,
    o_10_31_0_0  );
  input  i_10_31_32_0, i_10_31_88_0, i_10_31_133_0, i_10_31_151_0,
    i_10_31_266_0, i_10_31_349_0, i_10_31_364_0, i_10_31_393_0,
    i_10_31_394_0, i_10_31_431_0, i_10_31_464_0, i_10_31_465_0,
    i_10_31_466_0, i_10_31_566_0, i_10_31_591_0, i_10_31_592_0,
    i_10_31_673_0, i_10_31_674_0, i_10_31_750_0, i_10_31_754_0,
    i_10_31_770_0, i_10_31_798_0, i_10_31_952_0, i_10_31_953_0,
    i_10_31_976_0, i_10_31_996_0, i_10_31_1033_0, i_10_31_1052_0,
    i_10_31_1059_0, i_10_31_1235_0, i_10_31_1236_0, i_10_31_1238_0,
    i_10_31_1241_0, i_10_31_1312_0, i_10_31_1358_0, i_10_31_1382_0,
    i_10_31_1457_0, i_10_31_1491_0, i_10_31_1619_0, i_10_31_1822_0,
    i_10_31_1867_0, i_10_31_1906_0, i_10_31_1912_0, i_10_31_1913_0,
    i_10_31_1914_0, i_10_31_1952_0, i_10_31_1957_0, i_10_31_1958_0,
    i_10_31_1960_0, i_10_31_1987_0, i_10_31_2095_0, i_10_31_2275_0,
    i_10_31_2276_0, i_10_31_2362_0, i_10_31_2465_0, i_10_31_2481_0,
    i_10_31_2508_0, i_10_31_2516_0, i_10_31_2572_0, i_10_31_2644_0,
    i_10_31_2661_0, i_10_31_2662_0, i_10_31_2678_0, i_10_31_2712_0,
    i_10_31_2744_0, i_10_31_2782_0, i_10_31_2786_0, i_10_31_2914_0,
    i_10_31_2916_0, i_10_31_2948_0, i_10_31_2956_0, i_10_31_2960_0,
    i_10_31_3093_0, i_10_31_3175_0, i_10_31_3176_0, i_10_31_3198_0,
    i_10_31_3199_0, i_10_31_3362_0, i_10_31_3446_0, i_10_31_3451_0,
    i_10_31_3470_0, i_10_31_3472_0, i_10_31_3473_0, i_10_31_3495_0,
    i_10_31_3508_0, i_10_31_3614_0, i_10_31_3622_0, i_10_31_3642_0,
    i_10_31_3643_0, i_10_31_3649_0, i_10_31_3652_0, i_10_31_3858_0,
    i_10_31_3860_0, i_10_31_3885_0, i_10_31_4056_0, i_10_31_4057_0,
    i_10_31_4058_0, i_10_31_4129_0, i_10_31_4287_0, i_10_31_4526_0;
  output o_10_31_0_0;
  assign o_10_31_0_0 = ~((~i_10_31_1235_0 & ((~i_10_31_1241_0 & ((~i_10_31_466_0 & ((~i_10_31_2678_0 & ((~i_10_31_3614_0 & ((~i_10_31_32_0 & ~i_10_31_2644_0 & ((~i_10_31_266_0 & ~i_10_31_1491_0 & i_10_31_1822_0 & ~i_10_31_3198_0 & ~i_10_31_3649_0 & ~i_10_31_3860_0) | (~i_10_31_464_0 & ~i_10_31_1312_0 & ~i_10_31_1822_0 & ~i_10_31_1952_0 & ~i_10_31_2508_0 & ~i_10_31_2572_0 & ~i_10_31_2712_0 & ~i_10_31_3199_0 & ~i_10_31_3470_0 & ~i_10_31_3858_0 & ~i_10_31_4129_0))) | (~i_10_31_798_0 & ~i_10_31_3199_0 & i_10_31_3649_0 & ~i_10_31_3652_0))) | (~i_10_31_464_0 & ~i_10_31_4287_0 & ((~i_10_31_88_0 & ~i_10_31_151_0 & ~i_10_31_1312_0 & ~i_10_31_1952_0 & ~i_10_31_2465_0 & ~i_10_31_2508_0 & ~i_10_31_2786_0 & ~i_10_31_3198_0 & ~i_10_31_3199_0) | (~i_10_31_1033_0 & i_10_31_1822_0 & ~i_10_31_2362_0 & ~i_10_31_2782_0 & ~i_10_31_3508_0 & ~i_10_31_3858_0))))) | (~i_10_31_3470_0 & ((~i_10_31_151_0 & i_10_31_1033_0 & ~i_10_31_1238_0 & ~i_10_31_2644_0 & ~i_10_31_2786_0 & ~i_10_31_2916_0 & ~i_10_31_3858_0 & ~i_10_31_3860_0) | (~i_10_31_465_0 & i_10_31_1236_0 & ~i_10_31_3198_0 & ~i_10_31_4056_0))) | (~i_10_31_464_0 & ~i_10_31_1033_0 & ~i_10_31_1491_0 & i_10_31_1822_0 & ~i_10_31_3614_0 & ~i_10_31_3649_0 & ~i_10_31_4129_0))) | (~i_10_31_465_0 & i_10_31_1236_0 & ~i_10_31_3614_0 & ((~i_10_31_151_0 & ~i_10_31_393_0 & ~i_10_31_1491_0 & ~i_10_31_2782_0) | (~i_10_31_4056_0 & ~i_10_31_4287_0))) | (~i_10_31_3652_0 & ((i_10_31_1912_0 & ~i_10_31_2782_0) | (~i_10_31_88_0 & ~i_10_31_464_0 & ~i_10_31_2508_0 & ~i_10_31_2572_0 & ~i_10_31_3198_0 & i_10_31_4129_0 & ~i_10_31_4287_0))))) | (~i_10_31_465_0 & ((~i_10_31_464_0 & ~i_10_31_1033_0 & ~i_10_31_1236_0 & ~i_10_31_1822_0 & ~i_10_31_2362_0 & ~i_10_31_2661_0 & ~i_10_31_2782_0 & ~i_10_31_2786_0 & i_10_31_3652_0 & ~i_10_31_3858_0 & ~i_10_31_3860_0) | (i_10_31_464_0 & i_10_31_2916_0 & ~i_10_31_3199_0 & ~i_10_31_4287_0))) | (i_10_31_754_0 & ~i_10_31_2572_0 & ((~i_10_31_466_0 & ~i_10_31_2508_0 & ~i_10_31_3649_0) | (~i_10_31_151_0 & ~i_10_31_798_0 & ~i_10_31_1238_0 & ~i_10_31_1914_0 & ~i_10_31_3858_0 & ~i_10_31_3860_0 & ~i_10_31_2678_0 & ~i_10_31_3198_0))) | (~i_10_31_798_0 & ((~i_10_31_464_0 & ~i_10_31_1033_0 & ~i_10_31_1312_0 & ~i_10_31_1822_0 & ~i_10_31_1952_0 & ~i_10_31_2362_0 & ~i_10_31_2662_0 & ~i_10_31_2678_0 & ~i_10_31_2712_0 & ~i_10_31_3470_0 & ~i_10_31_3614_0 & ~i_10_31_3649_0 & ~i_10_31_3652_0 & ~i_10_31_3860_0) | (~i_10_31_466_0 & i_10_31_1913_0 & ~i_10_31_3198_0 & ~i_10_31_3199_0 & ~i_10_31_4129_0))) | (~i_10_31_464_0 & ((~i_10_31_393_0 & ~i_10_31_431_0 & ~i_10_31_466_0 & ~i_10_31_1312_0 & ~i_10_31_1491_0 & ~i_10_31_2362_0 & ~i_10_31_2508_0 & ~i_10_31_2644_0 & ~i_10_31_2661_0 & ~i_10_31_2678_0 & ~i_10_31_3198_0 & ~i_10_31_3199_0 & ~i_10_31_3470_0 & ~i_10_31_4129_0) | (i_10_31_2916_0 & i_10_31_3199_0 & ~i_10_31_3652_0 & ~i_10_31_3858_0 & ~i_10_31_4287_0))) | (~i_10_31_466_0 & ~i_10_31_2362_0 & ((~i_10_31_266_0 & i_10_31_1822_0 & i_10_31_2916_0 & i_10_31_3649_0 & ~i_10_31_3652_0 & i_10_31_4287_0) | (~i_10_31_1822_0 & ~i_10_31_2786_0 & ~i_10_31_3198_0 & i_10_31_3199_0 & ~i_10_31_3649_0 & ~i_10_31_4287_0))) | (i_10_31_1912_0 & ((i_10_31_798_0 & i_10_31_1236_0 & i_10_31_3198_0 & ~i_10_31_3473_0) | (~i_10_31_32_0 & ~i_10_31_566_0 & ~i_10_31_1312_0 & ~i_10_31_1914_0 & ~i_10_31_2712_0 & ~i_10_31_2782_0 & ~i_10_31_3198_0 & ~i_10_31_4129_0))))) | (~i_10_31_3858_0 & ((i_10_31_1033_0 & ~i_10_31_1822_0 & ((~i_10_31_151_0 & ~i_10_31_465_0 & ~i_10_31_466_0 & ~i_10_31_1238_0 & ~i_10_31_2572_0 & ~i_10_31_2661_0 & ~i_10_31_3470_0) | (~i_10_31_32_0 & i_10_31_151_0 & i_10_31_1312_0 & ~i_10_31_3860_0))) | (~i_10_31_1241_0 & ((~i_10_31_465_0 & ~i_10_31_2782_0 & ((~i_10_31_464_0 & ~i_10_31_2916_0 & ~i_10_31_3093_0 & i_10_31_3198_0 & ~i_10_31_3470_0 & ~i_10_31_3649_0) | (i_10_31_754_0 & ~i_10_31_1491_0 & i_10_31_1822_0 & i_10_31_3652_0))) | (~i_10_31_151_0 & ~i_10_31_2362_0 & ~i_10_31_2481_0 & i_10_31_3495_0 & ~i_10_31_3652_0 & ~i_10_31_4056_0))) | (~i_10_31_151_0 & i_10_31_1913_0 & ((~i_10_31_466_0 & i_10_31_1912_0 & ~i_10_31_2678_0) | (~i_10_31_2362_0 & i_10_31_3198_0 & ~i_10_31_4057_0 & ~i_10_31_4287_0))) | (~i_10_31_1238_0 & ((~i_10_31_431_0 & i_10_31_798_0 & i_10_31_1236_0 & ~i_10_31_1914_0 & ~i_10_31_2916_0 & ~i_10_31_3199_0 & ~i_10_31_3508_0 & ~i_10_31_4056_0) | (~i_10_31_754_0 & i_10_31_996_0 & ~i_10_31_1491_0 & ~i_10_31_2362_0 & ~i_10_31_4287_0))) | (~i_10_31_466_0 & i_10_31_1312_0 & i_10_31_2362_0 & ~i_10_31_2662_0 & ~i_10_31_2786_0 & ~i_10_31_3199_0) | (~i_10_31_750_0 & i_10_31_2662_0 & ~i_10_31_3508_0 & ~i_10_31_3614_0 & ~i_10_31_3649_0 & ~i_10_31_3860_0 & ~i_10_31_4129_0 & i_10_31_4287_0))) | (~i_10_31_3860_0 & ((~i_10_31_151_0 & i_10_31_754_0 & ~i_10_31_4129_0 & ((~i_10_31_464_0 & ~i_10_31_466_0 & i_10_31_1312_0 & ~i_10_31_2678_0) | (~i_10_31_1241_0 & ~i_10_31_1491_0 & ~i_10_31_2362_0 & ~i_10_31_3198_0 & ~i_10_31_4056_0))) | (~i_10_31_1241_0 & ((~i_10_31_1033_0 & i_10_31_2362_0 & ~i_10_31_2662_0 & i_10_31_3614_0 & i_10_31_3649_0 & i_10_31_3652_0) | (i_10_31_466_0 & i_10_31_1913_0 & ~i_10_31_1914_0 & ~i_10_31_3093_0 & ~i_10_31_3198_0 & ~i_10_31_3652_0))) | (i_10_31_996_0 & ((~i_10_31_2508_0 & ~i_10_31_2782_0 & ~i_10_31_3614_0 & ((~i_10_31_798_0 & ~i_10_31_1822_0 & ~i_10_31_1914_0 & i_10_31_2661_0 & ~i_10_31_3093_0) | (~i_10_31_466_0 & ~i_10_31_2916_0 & ~i_10_31_3199_0))) | (~i_10_31_464_0 & ~i_10_31_1238_0 & i_10_31_1822_0 & ~i_10_31_2678_0 & ~i_10_31_2786_0 & ~i_10_31_3093_0))) | (i_10_31_798_0 & i_10_31_1312_0 & ~i_10_31_2661_0 & ~i_10_31_3649_0 & i_10_31_3858_0))) | (~i_10_31_431_0 & ((~i_10_31_464_0 & ~i_10_31_1238_0 & i_10_31_1913_0 & ~i_10_31_2662_0) | (~i_10_31_466_0 & ~i_10_31_1952_0 & i_10_31_2481_0 & ~i_10_31_3649_0 & ~i_10_31_4129_0))) | (i_10_31_1822_0 & ((i_10_31_2465_0 & ~i_10_31_2644_0 & ~i_10_31_2786_0 & ~i_10_31_3614_0) | (~i_10_31_464_0 & i_10_31_465_0 & ~i_10_31_1491_0 & ~i_10_31_2661_0 & ~i_10_31_3199_0 & ~i_10_31_3649_0 & ~i_10_31_4056_0))) | (~i_10_31_1491_0 & ~i_10_31_4129_0 & ((~i_10_31_466_0 & i_10_31_3495_0) | (i_10_31_2481_0 & ~i_10_31_2508_0 & ~i_10_31_2644_0 & ~i_10_31_2678_0 & ~i_10_31_3649_0))) | (~i_10_31_1238_0 & ((~i_10_31_465_0 & ((~i_10_31_466_0 & i_10_31_798_0 & ~i_10_31_1952_0 & ~i_10_31_2362_0 & ~i_10_31_2508_0 & ~i_10_31_2678_0 & ~i_10_31_2712_0 & ~i_10_31_3649_0) | (i_10_31_1913_0 & ~i_10_31_2662_0 & i_10_31_3199_0 & ~i_10_31_3652_0))) | (i_10_31_1913_0 & (i_10_31_2916_0 | (~i_10_31_2662_0 & ~i_10_31_3614_0) | (~i_10_31_466_0 & i_10_31_3649_0))))) | (i_10_31_1912_0 & ((~i_10_31_88_0 & ~i_10_31_465_0 & ~i_10_31_566_0 & ~i_10_31_1312_0 & ~i_10_31_2661_0 & ~i_10_31_2782_0 & ~i_10_31_3199_0 & ~i_10_31_3470_0) | (~i_10_31_1241_0 & ~i_10_31_2678_0 & ~i_10_31_3198_0 & i_10_31_3652_0))) | (~i_10_31_1241_0 & ((~i_10_31_2662_0 & i_10_31_2678_0 & i_10_31_3472_0) | (~i_10_31_3649_0 & ~i_10_31_4056_0 & i_10_31_1236_0 & i_10_31_3495_0))) | (i_10_31_3495_0 & ((i_10_31_1952_0 & ~i_10_31_2508_0 & ~i_10_31_2678_0) | (i_10_31_2362_0 & ~i_10_31_2786_0 & i_10_31_4129_0))));
endmodule



// Benchmark "kernel_10_32" written by ABC on Sun Jul 19 10:21:35 2020

module kernel_10_32 ( 
    i_10_32_82_0, i_10_32_217_0, i_10_32_263_0, i_10_32_283_0,
    i_10_32_285_0, i_10_32_288_0, i_10_32_289_0, i_10_32_318_0,
    i_10_32_319_0, i_10_32_320_0, i_10_32_322_0, i_10_32_323_0,
    i_10_32_390_0, i_10_32_464_0, i_10_32_497_0, i_10_32_558_0,
    i_10_32_559_0, i_10_32_640_0, i_10_32_755_0, i_10_32_798_0,
    i_10_32_896_0, i_10_32_1000_0, i_10_32_1007_0, i_10_32_1027_0,
    i_10_32_1030_0, i_10_32_1234_0, i_10_32_1236_0, i_10_32_1308_0,
    i_10_32_1454_0, i_10_32_1575_0, i_10_32_1578_0, i_10_32_1579_0,
    i_10_32_1655_0, i_10_32_1691_0, i_10_32_1767_0, i_10_32_1819_0,
    i_10_32_1823_0, i_10_32_1909_0, i_10_32_1989_0, i_10_32_1993_0,
    i_10_32_2153_0, i_10_32_2196_0, i_10_32_2200_0, i_10_32_2297_0,
    i_10_32_2361_0, i_10_32_2364_0, i_10_32_2448_0, i_10_32_2514_0,
    i_10_32_2558_0, i_10_32_2566_0, i_10_32_2603_0, i_10_32_2631_0,
    i_10_32_2632_0, i_10_32_2647_0, i_10_32_2702_0, i_10_32_2711_0,
    i_10_32_2719_0, i_10_32_2723_0, i_10_32_2728_0, i_10_32_2730_0,
    i_10_32_2827_0, i_10_32_2831_0, i_10_32_2888_0, i_10_32_2917_0,
    i_10_32_2921_0, i_10_32_3073_0, i_10_32_3160_0, i_10_32_3234_0,
    i_10_32_3276_0, i_10_32_3385_0, i_10_32_3388_0, i_10_32_3523_0,
    i_10_32_3541_0, i_10_32_3543_0, i_10_32_3558_0, i_10_32_3565_0,
    i_10_32_3613_0, i_10_32_3720_0, i_10_32_3721_0, i_10_32_3785_0,
    i_10_32_3852_0, i_10_32_3889_0, i_10_32_3986_0, i_10_32_4023_0,
    i_10_32_4024_0, i_10_32_4096_0, i_10_32_4117_0, i_10_32_4119_0,
    i_10_32_4122_0, i_10_32_4123_0, i_10_32_4126_0, i_10_32_4153_0,
    i_10_32_4167_0, i_10_32_4168_0, i_10_32_4170_0, i_10_32_4171_0,
    i_10_32_4174_0, i_10_32_4275_0, i_10_32_4285_0, i_10_32_4571_0,
    o_10_32_0_0  );
  input  i_10_32_82_0, i_10_32_217_0, i_10_32_263_0, i_10_32_283_0,
    i_10_32_285_0, i_10_32_288_0, i_10_32_289_0, i_10_32_318_0,
    i_10_32_319_0, i_10_32_320_0, i_10_32_322_0, i_10_32_323_0,
    i_10_32_390_0, i_10_32_464_0, i_10_32_497_0, i_10_32_558_0,
    i_10_32_559_0, i_10_32_640_0, i_10_32_755_0, i_10_32_798_0,
    i_10_32_896_0, i_10_32_1000_0, i_10_32_1007_0, i_10_32_1027_0,
    i_10_32_1030_0, i_10_32_1234_0, i_10_32_1236_0, i_10_32_1308_0,
    i_10_32_1454_0, i_10_32_1575_0, i_10_32_1578_0, i_10_32_1579_0,
    i_10_32_1655_0, i_10_32_1691_0, i_10_32_1767_0, i_10_32_1819_0,
    i_10_32_1823_0, i_10_32_1909_0, i_10_32_1989_0, i_10_32_1993_0,
    i_10_32_2153_0, i_10_32_2196_0, i_10_32_2200_0, i_10_32_2297_0,
    i_10_32_2361_0, i_10_32_2364_0, i_10_32_2448_0, i_10_32_2514_0,
    i_10_32_2558_0, i_10_32_2566_0, i_10_32_2603_0, i_10_32_2631_0,
    i_10_32_2632_0, i_10_32_2647_0, i_10_32_2702_0, i_10_32_2711_0,
    i_10_32_2719_0, i_10_32_2723_0, i_10_32_2728_0, i_10_32_2730_0,
    i_10_32_2827_0, i_10_32_2831_0, i_10_32_2888_0, i_10_32_2917_0,
    i_10_32_2921_0, i_10_32_3073_0, i_10_32_3160_0, i_10_32_3234_0,
    i_10_32_3276_0, i_10_32_3385_0, i_10_32_3388_0, i_10_32_3523_0,
    i_10_32_3541_0, i_10_32_3543_0, i_10_32_3558_0, i_10_32_3565_0,
    i_10_32_3613_0, i_10_32_3720_0, i_10_32_3721_0, i_10_32_3785_0,
    i_10_32_3852_0, i_10_32_3889_0, i_10_32_3986_0, i_10_32_4023_0,
    i_10_32_4024_0, i_10_32_4096_0, i_10_32_4117_0, i_10_32_4119_0,
    i_10_32_4122_0, i_10_32_4123_0, i_10_32_4126_0, i_10_32_4153_0,
    i_10_32_4167_0, i_10_32_4168_0, i_10_32_4170_0, i_10_32_4171_0,
    i_10_32_4174_0, i_10_32_4275_0, i_10_32_4285_0, i_10_32_4571_0;
  output o_10_32_0_0;
  assign o_10_32_0_0 = 0;
endmodule



// Benchmark "kernel_10_33" written by ABC on Sun Jul 19 10:21:36 2020

module kernel_10_33 ( 
    i_10_33_279_0, i_10_33_441_0, i_10_33_442_0, i_10_33_445_0,
    i_10_33_446_0, i_10_33_469_0, i_10_33_590_0, i_10_33_733_0,
    i_10_33_736_0, i_10_33_737_0, i_10_33_784_0, i_10_33_901_0,
    i_10_33_932_0, i_10_33_1031_0, i_10_33_1043_0, i_10_33_1120_0,
    i_10_33_1240_0, i_10_33_1249_0, i_10_33_1343_0, i_10_33_1391_0,
    i_10_33_1552_0, i_10_33_1683_0, i_10_33_1685_0, i_10_33_1690_0,
    i_10_33_1765_0, i_10_33_1766_0, i_10_33_1822_0, i_10_33_1888_0,
    i_10_33_1909_0, i_10_33_1912_0, i_10_33_1913_0, i_10_33_2243_0,
    i_10_33_2380_0, i_10_33_2462_0, i_10_33_2464_0, i_10_33_2476_0,
    i_10_33_2514_0, i_10_33_2542_0, i_10_33_2543_0, i_10_33_2571_0,
    i_10_33_2635_0, i_10_33_2644_0, i_10_33_2645_0, i_10_33_2653_0,
    i_10_33_2654_0, i_10_33_2663_0, i_10_33_2701_0, i_10_33_2710_0,
    i_10_33_2719_0, i_10_33_2727_0, i_10_33_2728_0, i_10_33_2729_0,
    i_10_33_2731_0, i_10_33_2732_0, i_10_33_2734_0, i_10_33_2737_0,
    i_10_33_2820_0, i_10_33_2831_0, i_10_33_2920_0, i_10_33_2923_0,
    i_10_33_2983_0, i_10_33_3033_0, i_10_33_3048_0, i_10_33_3076_0,
    i_10_33_3114_0, i_10_33_3201_0, i_10_33_3202_0, i_10_33_3279_0,
    i_10_33_3352_0, i_10_33_3353_0, i_10_33_3356_0, i_10_33_3390_0,
    i_10_33_3391_0, i_10_33_3392_0, i_10_33_3522_0, i_10_33_3538_0,
    i_10_33_3551_0, i_10_33_3612_0, i_10_33_3614_0, i_10_33_3616_0,
    i_10_33_3800_0, i_10_33_3839_0, i_10_33_3841_0, i_10_33_3859_0,
    i_10_33_3860_0, i_10_33_3887_0, i_10_33_3923_0, i_10_33_3981_0,
    i_10_33_4124_0, i_10_33_4154_0, i_10_33_4156_0, i_10_33_4183_0,
    i_10_33_4238_0, i_10_33_4270_0, i_10_33_4273_0, i_10_33_4288_0,
    i_10_33_4459_0, i_10_33_4568_0, i_10_33_4570_0, i_10_33_4594_0,
    o_10_33_0_0  );
  input  i_10_33_279_0, i_10_33_441_0, i_10_33_442_0, i_10_33_445_0,
    i_10_33_446_0, i_10_33_469_0, i_10_33_590_0, i_10_33_733_0,
    i_10_33_736_0, i_10_33_737_0, i_10_33_784_0, i_10_33_901_0,
    i_10_33_932_0, i_10_33_1031_0, i_10_33_1043_0, i_10_33_1120_0,
    i_10_33_1240_0, i_10_33_1249_0, i_10_33_1343_0, i_10_33_1391_0,
    i_10_33_1552_0, i_10_33_1683_0, i_10_33_1685_0, i_10_33_1690_0,
    i_10_33_1765_0, i_10_33_1766_0, i_10_33_1822_0, i_10_33_1888_0,
    i_10_33_1909_0, i_10_33_1912_0, i_10_33_1913_0, i_10_33_2243_0,
    i_10_33_2380_0, i_10_33_2462_0, i_10_33_2464_0, i_10_33_2476_0,
    i_10_33_2514_0, i_10_33_2542_0, i_10_33_2543_0, i_10_33_2571_0,
    i_10_33_2635_0, i_10_33_2644_0, i_10_33_2645_0, i_10_33_2653_0,
    i_10_33_2654_0, i_10_33_2663_0, i_10_33_2701_0, i_10_33_2710_0,
    i_10_33_2719_0, i_10_33_2727_0, i_10_33_2728_0, i_10_33_2729_0,
    i_10_33_2731_0, i_10_33_2732_0, i_10_33_2734_0, i_10_33_2737_0,
    i_10_33_2820_0, i_10_33_2831_0, i_10_33_2920_0, i_10_33_2923_0,
    i_10_33_2983_0, i_10_33_3033_0, i_10_33_3048_0, i_10_33_3076_0,
    i_10_33_3114_0, i_10_33_3201_0, i_10_33_3202_0, i_10_33_3279_0,
    i_10_33_3352_0, i_10_33_3353_0, i_10_33_3356_0, i_10_33_3390_0,
    i_10_33_3391_0, i_10_33_3392_0, i_10_33_3522_0, i_10_33_3538_0,
    i_10_33_3551_0, i_10_33_3612_0, i_10_33_3614_0, i_10_33_3616_0,
    i_10_33_3800_0, i_10_33_3839_0, i_10_33_3841_0, i_10_33_3859_0,
    i_10_33_3860_0, i_10_33_3887_0, i_10_33_3923_0, i_10_33_3981_0,
    i_10_33_4124_0, i_10_33_4154_0, i_10_33_4156_0, i_10_33_4183_0,
    i_10_33_4238_0, i_10_33_4270_0, i_10_33_4273_0, i_10_33_4288_0,
    i_10_33_4459_0, i_10_33_4568_0, i_10_33_4570_0, i_10_33_4594_0;
  output o_10_33_0_0;
  assign o_10_33_0_0 = 0;
endmodule



// Benchmark "kernel_10_34" written by ABC on Sun Jul 19 10:21:36 2020

module kernel_10_34 ( 
    i_10_34_14_0, i_10_34_41_0, i_10_34_175_0, i_10_34_176_0,
    i_10_34_260_0, i_10_34_266_0, i_10_34_320_0, i_10_34_388_0,
    i_10_34_429_0, i_10_34_500_0, i_10_34_508_0, i_10_34_509_0,
    i_10_34_559_0, i_10_34_714_0, i_10_34_718_0, i_10_34_866_0,
    i_10_34_956_0, i_10_34_993_0, i_10_34_1055_0, i_10_34_1112_0,
    i_10_34_1115_0, i_10_34_1207_0, i_10_34_1211_0, i_10_34_1220_0,
    i_10_34_1236_0, i_10_34_1301_0, i_10_34_1360_0, i_10_34_1366_0,
    i_10_34_1379_0, i_10_34_1380_0, i_10_34_1541_0, i_10_34_1544_0,
    i_10_34_1621_0, i_10_34_1634_0, i_10_34_1650_0, i_10_34_1685_0,
    i_10_34_1687_0, i_10_34_1691_0, i_10_34_1733_0, i_10_34_1802_0,
    i_10_34_1877_0, i_10_34_1920_0, i_10_34_1921_0, i_10_34_1981_0,
    i_10_34_1985_0, i_10_34_2003_0, i_10_34_2027_0, i_10_34_2030_0,
    i_10_34_2036_0, i_10_34_2089_0, i_10_34_2204_0, i_10_34_2341_0,
    i_10_34_2359_0, i_10_34_2372_0, i_10_34_2383_0, i_10_34_2467_0,
    i_10_34_2471_0, i_10_34_2558_0, i_10_34_2576_0, i_10_34_2596_0,
    i_10_34_2734_0, i_10_34_2836_0, i_10_34_2839_0, i_10_34_2849_0,
    i_10_34_2851_0, i_10_34_2864_0, i_10_34_2867_0, i_10_34_2963_0,
    i_10_34_2966_0, i_10_34_2972_0, i_10_34_2975_0, i_10_34_3223_0,
    i_10_34_3313_0, i_10_34_3352_0, i_10_34_3353_0, i_10_34_3388_0,
    i_10_34_3466_0, i_10_34_3485_0, i_10_34_3506_0, i_10_34_3519_0,
    i_10_34_3541_0, i_10_34_3542_0, i_10_34_3545_0, i_10_34_3611_0,
    i_10_34_3794_0, i_10_34_3841_0, i_10_34_3842_0, i_10_34_3856_0,
    i_10_34_3908_0, i_10_34_3943_0, i_10_34_4027_0, i_10_34_4028_0,
    i_10_34_4118_0, i_10_34_4127_0, i_10_34_4148_0, i_10_34_4153_0,
    i_10_34_4169_0, i_10_34_4205_0, i_10_34_4287_0, i_10_34_4395_0,
    o_10_34_0_0  );
  input  i_10_34_14_0, i_10_34_41_0, i_10_34_175_0, i_10_34_176_0,
    i_10_34_260_0, i_10_34_266_0, i_10_34_320_0, i_10_34_388_0,
    i_10_34_429_0, i_10_34_500_0, i_10_34_508_0, i_10_34_509_0,
    i_10_34_559_0, i_10_34_714_0, i_10_34_718_0, i_10_34_866_0,
    i_10_34_956_0, i_10_34_993_0, i_10_34_1055_0, i_10_34_1112_0,
    i_10_34_1115_0, i_10_34_1207_0, i_10_34_1211_0, i_10_34_1220_0,
    i_10_34_1236_0, i_10_34_1301_0, i_10_34_1360_0, i_10_34_1366_0,
    i_10_34_1379_0, i_10_34_1380_0, i_10_34_1541_0, i_10_34_1544_0,
    i_10_34_1621_0, i_10_34_1634_0, i_10_34_1650_0, i_10_34_1685_0,
    i_10_34_1687_0, i_10_34_1691_0, i_10_34_1733_0, i_10_34_1802_0,
    i_10_34_1877_0, i_10_34_1920_0, i_10_34_1921_0, i_10_34_1981_0,
    i_10_34_1985_0, i_10_34_2003_0, i_10_34_2027_0, i_10_34_2030_0,
    i_10_34_2036_0, i_10_34_2089_0, i_10_34_2204_0, i_10_34_2341_0,
    i_10_34_2359_0, i_10_34_2372_0, i_10_34_2383_0, i_10_34_2467_0,
    i_10_34_2471_0, i_10_34_2558_0, i_10_34_2576_0, i_10_34_2596_0,
    i_10_34_2734_0, i_10_34_2836_0, i_10_34_2839_0, i_10_34_2849_0,
    i_10_34_2851_0, i_10_34_2864_0, i_10_34_2867_0, i_10_34_2963_0,
    i_10_34_2966_0, i_10_34_2972_0, i_10_34_2975_0, i_10_34_3223_0,
    i_10_34_3313_0, i_10_34_3352_0, i_10_34_3353_0, i_10_34_3388_0,
    i_10_34_3466_0, i_10_34_3485_0, i_10_34_3506_0, i_10_34_3519_0,
    i_10_34_3541_0, i_10_34_3542_0, i_10_34_3545_0, i_10_34_3611_0,
    i_10_34_3794_0, i_10_34_3841_0, i_10_34_3842_0, i_10_34_3856_0,
    i_10_34_3908_0, i_10_34_3943_0, i_10_34_4027_0, i_10_34_4028_0,
    i_10_34_4118_0, i_10_34_4127_0, i_10_34_4148_0, i_10_34_4153_0,
    i_10_34_4169_0, i_10_34_4205_0, i_10_34_4287_0, i_10_34_4395_0;
  output o_10_34_0_0;
  assign o_10_34_0_0 = 0;
endmodule



// Benchmark "kernel_10_35" written by ABC on Sun Jul 19 10:21:37 2020

module kernel_10_35 ( 
    i_10_35_174_0, i_10_35_176_0, i_10_35_407_0, i_10_35_409_0,
    i_10_35_443_0, i_10_35_520_0, i_10_35_697_0, i_10_35_798_0,
    i_10_35_799_0, i_10_35_956_0, i_10_35_958_0, i_10_35_998_0,
    i_10_35_1032_0, i_10_35_1246_0, i_10_35_1248_0, i_10_35_1249_0,
    i_10_35_1250_0, i_10_35_1308_0, i_10_35_1309_0, i_10_35_1310_0,
    i_10_35_1311_0, i_10_35_1432_0, i_10_35_1439_0, i_10_35_1552_0,
    i_10_35_1619_0, i_10_35_1650_0, i_10_35_1651_0, i_10_35_1687_0,
    i_10_35_1690_0, i_10_35_1691_0, i_10_35_1821_0, i_10_35_1822_0,
    i_10_35_1825_0, i_10_35_1996_0, i_10_35_2021_0, i_10_35_2023_0,
    i_10_35_2201_0, i_10_35_2365_0, i_10_35_2366_0, i_10_35_2451_0,
    i_10_35_2452_0, i_10_35_2463_0, i_10_35_2464_0, i_10_35_2470_0,
    i_10_35_2473_0, i_10_35_2514_0, i_10_35_2571_0, i_10_35_2702_0,
    i_10_35_2705_0, i_10_35_2711_0, i_10_35_2722_0, i_10_35_2725_0,
    i_10_35_2829_0, i_10_35_2832_0, i_10_35_2833_0, i_10_35_2920_0,
    i_10_35_2923_0, i_10_35_2924_0, i_10_35_3072_0, i_10_35_3074_0,
    i_10_35_3075_0, i_10_35_3112_0, i_10_35_3199_0, i_10_35_3270_0,
    i_10_35_3273_0, i_10_35_3277_0, i_10_35_3284_0, i_10_35_3386_0,
    i_10_35_3407_0, i_10_35_3408_0, i_10_35_3586_0, i_10_35_3609_0,
    i_10_35_3612_0, i_10_35_3613_0, i_10_35_3614_0, i_10_35_3615_0,
    i_10_35_3732_0, i_10_35_3733_0, i_10_35_3734_0, i_10_35_3780_0,
    i_10_35_3781_0, i_10_35_3782_0, i_10_35_3786_0, i_10_35_3787_0,
    i_10_35_3788_0, i_10_35_3841_0, i_10_35_3856_0, i_10_35_4029_0,
    i_10_35_4114_0, i_10_35_4116_0, i_10_35_4125_0, i_10_35_4130_0,
    i_10_35_4216_0, i_10_35_4217_0, i_10_35_4218_0, i_10_35_4269_0,
    i_10_35_4275_0, i_10_35_4290_0, i_10_35_4564_0, i_10_35_4565_0,
    o_10_35_0_0  );
  input  i_10_35_174_0, i_10_35_176_0, i_10_35_407_0, i_10_35_409_0,
    i_10_35_443_0, i_10_35_520_0, i_10_35_697_0, i_10_35_798_0,
    i_10_35_799_0, i_10_35_956_0, i_10_35_958_0, i_10_35_998_0,
    i_10_35_1032_0, i_10_35_1246_0, i_10_35_1248_0, i_10_35_1249_0,
    i_10_35_1250_0, i_10_35_1308_0, i_10_35_1309_0, i_10_35_1310_0,
    i_10_35_1311_0, i_10_35_1432_0, i_10_35_1439_0, i_10_35_1552_0,
    i_10_35_1619_0, i_10_35_1650_0, i_10_35_1651_0, i_10_35_1687_0,
    i_10_35_1690_0, i_10_35_1691_0, i_10_35_1821_0, i_10_35_1822_0,
    i_10_35_1825_0, i_10_35_1996_0, i_10_35_2021_0, i_10_35_2023_0,
    i_10_35_2201_0, i_10_35_2365_0, i_10_35_2366_0, i_10_35_2451_0,
    i_10_35_2452_0, i_10_35_2463_0, i_10_35_2464_0, i_10_35_2470_0,
    i_10_35_2473_0, i_10_35_2514_0, i_10_35_2571_0, i_10_35_2702_0,
    i_10_35_2705_0, i_10_35_2711_0, i_10_35_2722_0, i_10_35_2725_0,
    i_10_35_2829_0, i_10_35_2832_0, i_10_35_2833_0, i_10_35_2920_0,
    i_10_35_2923_0, i_10_35_2924_0, i_10_35_3072_0, i_10_35_3074_0,
    i_10_35_3075_0, i_10_35_3112_0, i_10_35_3199_0, i_10_35_3270_0,
    i_10_35_3273_0, i_10_35_3277_0, i_10_35_3284_0, i_10_35_3386_0,
    i_10_35_3407_0, i_10_35_3408_0, i_10_35_3586_0, i_10_35_3609_0,
    i_10_35_3612_0, i_10_35_3613_0, i_10_35_3614_0, i_10_35_3615_0,
    i_10_35_3732_0, i_10_35_3733_0, i_10_35_3734_0, i_10_35_3780_0,
    i_10_35_3781_0, i_10_35_3782_0, i_10_35_3786_0, i_10_35_3787_0,
    i_10_35_3788_0, i_10_35_3841_0, i_10_35_3856_0, i_10_35_4029_0,
    i_10_35_4114_0, i_10_35_4116_0, i_10_35_4125_0, i_10_35_4130_0,
    i_10_35_4216_0, i_10_35_4217_0, i_10_35_4218_0, i_10_35_4269_0,
    i_10_35_4275_0, i_10_35_4290_0, i_10_35_4564_0, i_10_35_4565_0;
  output o_10_35_0_0;
  assign o_10_35_0_0 = ~(~i_10_35_4130_0 | ~i_10_35_3733_0 | ~i_10_35_3734_0 | ~i_10_35_2832_0 | ~i_10_35_3732_0 | ~i_10_35_176_0 | ~i_10_35_1249_0);
endmodule



// Benchmark "kernel_10_36" written by ABC on Sun Jul 19 10:21:38 2020

module kernel_10_36 ( 
    i_10_36_32_0, i_10_36_34_0, i_10_36_173_0, i_10_36_224_0,
    i_10_36_245_0, i_10_36_247_0, i_10_36_248_0, i_10_36_253_0,
    i_10_36_254_0, i_10_36_260_0, i_10_36_266_0, i_10_36_434_0,
    i_10_36_496_0, i_10_36_542_0, i_10_36_716_0, i_10_36_717_0,
    i_10_36_793_0, i_10_36_795_0, i_10_36_799_0, i_10_36_901_0,
    i_10_36_956_0, i_10_36_1030_0, i_10_36_1234_0, i_10_36_1236_0,
    i_10_36_1237_0, i_10_36_1238_0, i_10_36_1246_0, i_10_36_1247_0,
    i_10_36_1310_0, i_10_36_1325_0, i_10_36_1349_0, i_10_36_1435_0,
    i_10_36_1436_0, i_10_36_1437_0, i_10_36_1439_0, i_10_36_1543_0,
    i_10_36_1579_0, i_10_36_1580_0, i_10_36_1583_0, i_10_36_1653_0,
    i_10_36_1654_0, i_10_36_1655_0, i_10_36_1685_0, i_10_36_1686_0,
    i_10_36_1688_0, i_10_36_1689_0, i_10_36_1690_0, i_10_36_1909_0,
    i_10_36_1937_0, i_10_36_1948_0, i_10_36_1949_0, i_10_36_1954_0,
    i_10_36_2365_0, i_10_36_2387_0, i_10_36_2449_0, i_10_36_2454_0,
    i_10_36_2474_0, i_10_36_2477_0, i_10_36_2511_0, i_10_36_2531_0,
    i_10_36_2532_0, i_10_36_2540_0, i_10_36_2601_0, i_10_36_2660_0,
    i_10_36_2661_0, i_10_36_2730_0, i_10_36_2735_0, i_10_36_2881_0,
    i_10_36_2885_0, i_10_36_2918_0, i_10_36_3072_0, i_10_36_3197_0,
    i_10_36_3199_0, i_10_36_3201_0, i_10_36_3233_0, i_10_36_3281_0,
    i_10_36_3295_0, i_10_36_3332_0, i_10_36_3341_0, i_10_36_3493_0,
    i_10_36_3522_0, i_10_36_3523_0, i_10_36_3545_0, i_10_36_3586_0,
    i_10_36_3611_0, i_10_36_3646_0, i_10_36_3733_0, i_10_36_3784_0,
    i_10_36_3809_0, i_10_36_3841_0, i_10_36_3842_0, i_10_36_3883_0,
    i_10_36_3983_0, i_10_36_3997_0, i_10_36_4007_0, i_10_36_4116_0,
    i_10_36_4126_0, i_10_36_4367_0, i_10_36_4385_0, i_10_36_4585_0,
    o_10_36_0_0  );
  input  i_10_36_32_0, i_10_36_34_0, i_10_36_173_0, i_10_36_224_0,
    i_10_36_245_0, i_10_36_247_0, i_10_36_248_0, i_10_36_253_0,
    i_10_36_254_0, i_10_36_260_0, i_10_36_266_0, i_10_36_434_0,
    i_10_36_496_0, i_10_36_542_0, i_10_36_716_0, i_10_36_717_0,
    i_10_36_793_0, i_10_36_795_0, i_10_36_799_0, i_10_36_901_0,
    i_10_36_956_0, i_10_36_1030_0, i_10_36_1234_0, i_10_36_1236_0,
    i_10_36_1237_0, i_10_36_1238_0, i_10_36_1246_0, i_10_36_1247_0,
    i_10_36_1310_0, i_10_36_1325_0, i_10_36_1349_0, i_10_36_1435_0,
    i_10_36_1436_0, i_10_36_1437_0, i_10_36_1439_0, i_10_36_1543_0,
    i_10_36_1579_0, i_10_36_1580_0, i_10_36_1583_0, i_10_36_1653_0,
    i_10_36_1654_0, i_10_36_1655_0, i_10_36_1685_0, i_10_36_1686_0,
    i_10_36_1688_0, i_10_36_1689_0, i_10_36_1690_0, i_10_36_1909_0,
    i_10_36_1937_0, i_10_36_1948_0, i_10_36_1949_0, i_10_36_1954_0,
    i_10_36_2365_0, i_10_36_2387_0, i_10_36_2449_0, i_10_36_2454_0,
    i_10_36_2474_0, i_10_36_2477_0, i_10_36_2511_0, i_10_36_2531_0,
    i_10_36_2532_0, i_10_36_2540_0, i_10_36_2601_0, i_10_36_2660_0,
    i_10_36_2661_0, i_10_36_2730_0, i_10_36_2735_0, i_10_36_2881_0,
    i_10_36_2885_0, i_10_36_2918_0, i_10_36_3072_0, i_10_36_3197_0,
    i_10_36_3199_0, i_10_36_3201_0, i_10_36_3233_0, i_10_36_3281_0,
    i_10_36_3295_0, i_10_36_3332_0, i_10_36_3341_0, i_10_36_3493_0,
    i_10_36_3522_0, i_10_36_3523_0, i_10_36_3545_0, i_10_36_3586_0,
    i_10_36_3611_0, i_10_36_3646_0, i_10_36_3733_0, i_10_36_3784_0,
    i_10_36_3809_0, i_10_36_3841_0, i_10_36_3842_0, i_10_36_3883_0,
    i_10_36_3983_0, i_10_36_3997_0, i_10_36_4007_0, i_10_36_4116_0,
    i_10_36_4126_0, i_10_36_4367_0, i_10_36_4385_0, i_10_36_4585_0;
  output o_10_36_0_0;
  assign o_10_36_0_0 = 0;
endmodule



// Benchmark "kernel_10_37" written by ABC on Sun Jul 19 10:21:40 2020

module kernel_10_37 ( 
    i_10_37_176_0, i_10_37_251_0, i_10_37_282_0, i_10_37_283_0,
    i_10_37_284_0, i_10_37_289_0, i_10_37_320_0, i_10_37_329_0,
    i_10_37_425_0, i_10_37_434_0, i_10_37_442_0, i_10_37_458_0,
    i_10_37_460_0, i_10_37_461_0, i_10_37_464_0, i_10_37_749_0,
    i_10_37_755_0, i_10_37_792_0, i_10_37_796_0, i_10_37_965_0,
    i_10_37_1238_0, i_10_37_1239_0, i_10_37_1242_0, i_10_37_1243_0,
    i_10_37_1250_0, i_10_37_1310_0, i_10_37_1575_0, i_10_37_1576_0,
    i_10_37_1655_0, i_10_37_1681_0, i_10_37_1686_0, i_10_37_1687_0,
    i_10_37_1688_0, i_10_37_1768_0, i_10_37_1819_0, i_10_37_1823_0,
    i_10_37_1824_0, i_10_37_1990_0, i_10_37_1991_0, i_10_37_2197_0,
    i_10_37_2351_0, i_10_37_2353_0, i_10_37_2354_0, i_10_37_2359_0,
    i_10_37_2361_0, i_10_37_2362_0, i_10_37_2363_0, i_10_37_2449_0,
    i_10_37_2452_0, i_10_37_2453_0, i_10_37_2467_0, i_10_37_2468_0,
    i_10_37_2474_0, i_10_37_2632_0, i_10_37_2633_0, i_10_37_2657_0,
    i_10_37_2674_0, i_10_37_2710_0, i_10_37_2782_0, i_10_37_2783_0,
    i_10_37_2830_0, i_10_37_2919_0, i_10_37_3043_0, i_10_37_3044_0,
    i_10_37_3088_0, i_10_37_3151_0, i_10_37_3199_0, i_10_37_3271_0,
    i_10_37_3273_0, i_10_37_3277_0, i_10_37_3388_0, i_10_37_3406_0,
    i_10_37_3409_0, i_10_37_3467_0, i_10_37_3496_0, i_10_37_3550_0,
    i_10_37_3587_0, i_10_37_3610_0, i_10_37_3617_0, i_10_37_3648_0,
    i_10_37_3785_0, i_10_37_3786_0, i_10_37_3838_0, i_10_37_3850_0,
    i_10_37_3853_0, i_10_37_3856_0, i_10_37_3857_0, i_10_37_3858_0,
    i_10_37_3888_0, i_10_37_3889_0, i_10_37_3949_0, i_10_37_3991_0,
    i_10_37_4050_0, i_10_37_4115_0, i_10_37_4117_0, i_10_37_4121_0,
    i_10_37_4267_0, i_10_37_4288_0, i_10_37_4289_0, i_10_37_4568_0,
    o_10_37_0_0  );
  input  i_10_37_176_0, i_10_37_251_0, i_10_37_282_0, i_10_37_283_0,
    i_10_37_284_0, i_10_37_289_0, i_10_37_320_0, i_10_37_329_0,
    i_10_37_425_0, i_10_37_434_0, i_10_37_442_0, i_10_37_458_0,
    i_10_37_460_0, i_10_37_461_0, i_10_37_464_0, i_10_37_749_0,
    i_10_37_755_0, i_10_37_792_0, i_10_37_796_0, i_10_37_965_0,
    i_10_37_1238_0, i_10_37_1239_0, i_10_37_1242_0, i_10_37_1243_0,
    i_10_37_1250_0, i_10_37_1310_0, i_10_37_1575_0, i_10_37_1576_0,
    i_10_37_1655_0, i_10_37_1681_0, i_10_37_1686_0, i_10_37_1687_0,
    i_10_37_1688_0, i_10_37_1768_0, i_10_37_1819_0, i_10_37_1823_0,
    i_10_37_1824_0, i_10_37_1990_0, i_10_37_1991_0, i_10_37_2197_0,
    i_10_37_2351_0, i_10_37_2353_0, i_10_37_2354_0, i_10_37_2359_0,
    i_10_37_2361_0, i_10_37_2362_0, i_10_37_2363_0, i_10_37_2449_0,
    i_10_37_2452_0, i_10_37_2453_0, i_10_37_2467_0, i_10_37_2468_0,
    i_10_37_2474_0, i_10_37_2632_0, i_10_37_2633_0, i_10_37_2657_0,
    i_10_37_2674_0, i_10_37_2710_0, i_10_37_2782_0, i_10_37_2783_0,
    i_10_37_2830_0, i_10_37_2919_0, i_10_37_3043_0, i_10_37_3044_0,
    i_10_37_3088_0, i_10_37_3151_0, i_10_37_3199_0, i_10_37_3271_0,
    i_10_37_3273_0, i_10_37_3277_0, i_10_37_3388_0, i_10_37_3406_0,
    i_10_37_3409_0, i_10_37_3467_0, i_10_37_3496_0, i_10_37_3550_0,
    i_10_37_3587_0, i_10_37_3610_0, i_10_37_3617_0, i_10_37_3648_0,
    i_10_37_3785_0, i_10_37_3786_0, i_10_37_3838_0, i_10_37_3850_0,
    i_10_37_3853_0, i_10_37_3856_0, i_10_37_3857_0, i_10_37_3858_0,
    i_10_37_3888_0, i_10_37_3889_0, i_10_37_3949_0, i_10_37_3991_0,
    i_10_37_4050_0, i_10_37_4115_0, i_10_37_4117_0, i_10_37_4121_0,
    i_10_37_4267_0, i_10_37_4288_0, i_10_37_4289_0, i_10_37_4568_0;
  output o_10_37_0_0;
  assign o_10_37_0_0 = ~((~i_10_37_282_0 & ((~i_10_37_460_0 & i_10_37_1687_0 & ~i_10_37_2474_0 & ~i_10_37_4050_0 & i_10_37_4115_0) | (~i_10_37_458_0 & ~i_10_37_1239_0 & ~i_10_37_1655_0 & ~i_10_37_2453_0 & i_10_37_3199_0 & ~i_10_37_4121_0 & ~i_10_37_4568_0))) | (i_10_37_460_0 & ((~i_10_37_284_0 & ~i_10_37_1824_0 & i_10_37_2632_0 & i_10_37_2783_0 & ~i_10_37_3838_0) | (~i_10_37_320_0 & ~i_10_37_2351_0 & ~i_10_37_2830_0 & ~i_10_37_3043_0 & ~i_10_37_4050_0))) | (~i_10_37_3786_0 & ((~i_10_37_251_0 & ~i_10_37_3550_0 & ((~i_10_37_284_0 & ~i_10_37_1310_0 & ~i_10_37_1991_0 & ~i_10_37_2354_0 & ~i_10_37_3044_0 & ~i_10_37_4050_0) | (~i_10_37_176_0 & ~i_10_37_2474_0 & ~i_10_37_2674_0 & ~i_10_37_2783_0 & ~i_10_37_3088_0 & ~i_10_37_3648_0 & ~i_10_37_3785_0 & ~i_10_37_4288_0))) | (~i_10_37_425_0 & ~i_10_37_442_0 & ~i_10_37_755_0 & ~i_10_37_1310_0 & ~i_10_37_3273_0 & ~i_10_37_3617_0 & ~i_10_37_3850_0 & ~i_10_37_3853_0 & ~i_10_37_3991_0))) | (~i_10_37_284_0 & ((~i_10_37_2452_0 & ~i_10_37_3043_0 & ~i_10_37_3838_0 & ~i_10_37_4117_0) | (~i_10_37_251_0 & ~i_10_37_755_0 & ~i_10_37_1990_0 & i_10_37_2632_0 & ~i_10_37_3088_0 & ~i_10_37_4568_0))) | (i_10_37_1819_0 & ((~i_10_37_251_0 & ~i_10_37_1990_0 & ~i_10_37_1991_0 & ~i_10_37_2674_0 & ~i_10_37_3467_0) | (~i_10_37_2197_0 & ~i_10_37_2452_0 & ~i_10_37_2453_0 & ~i_10_37_2468_0 & ~i_10_37_3785_0 & ~i_10_37_3838_0 & ~i_10_37_4568_0))) | (~i_10_37_1990_0 & ((~i_10_37_251_0 & ~i_10_37_2361_0 & ~i_10_37_2453_0 & ~i_10_37_2782_0 & ~i_10_37_3857_0) | (~i_10_37_2363_0 & i_10_37_3406_0 & ~i_10_37_3785_0 & ~i_10_37_3991_0 & i_10_37_4288_0))) | (~i_10_37_2361_0 & ((~i_10_37_2363_0 & ((~i_10_37_289_0 & ~i_10_37_458_0 & ~i_10_37_2362_0 & ~i_10_37_2453_0 & ~i_10_37_2919_0 & ~i_10_37_3199_0 & ~i_10_37_3467_0 & ~i_10_37_3853_0 & ~i_10_37_4050_0) | (~i_10_37_460_0 & ~i_10_37_755_0 & ~i_10_37_1239_0 & ~i_10_37_1250_0 & ~i_10_37_2657_0 & ~i_10_37_3388_0 & ~i_10_37_4568_0))) | (~i_10_37_1991_0 & ~i_10_37_2783_0 & ~i_10_37_2919_0 & ~i_10_37_3785_0 & ~i_10_37_3857_0 & ~i_10_37_3991_0 & ~i_10_37_4050_0))) | (~i_10_37_1823_0 & ((~i_10_37_251_0 & ((~i_10_37_1250_0 & ~i_10_37_1768_0 & ~i_10_37_2362_0 & ~i_10_37_2467_0 & ~i_10_37_2710_0) | (i_10_37_2353_0 & ~i_10_37_3850_0))) | (~i_10_37_4117_0 & ((~i_10_37_2362_0 & ~i_10_37_2453_0 & i_10_37_2830_0 & ~i_10_37_3043_0) | (i_10_37_796_0 & ~i_10_37_1250_0 & ~i_10_37_1655_0 & ~i_10_37_1824_0 & ~i_10_37_3550_0 & ~i_10_37_3587_0 & ~i_10_37_4289_0))))) | (i_10_37_329_0 & i_10_37_2632_0) | (i_10_37_1239_0 & i_10_37_1310_0 & i_10_37_2474_0 & ~i_10_37_3043_0) | (~i_10_37_1243_0 & i_10_37_2633_0 & ~i_10_37_2782_0 & ~i_10_37_3273_0 & i_10_37_3409_0 & ~i_10_37_3550_0) | (i_10_37_792_0 & ~i_10_37_796_0 & i_10_37_3648_0) | (~i_10_37_2452_0 & ~i_10_37_2453_0 & i_10_37_3277_0 & ~i_10_37_3838_0) | (i_10_37_3273_0 & ~i_10_37_3785_0 & i_10_37_3858_0) | (~i_10_37_1819_0 & i_10_37_2197_0 & ~i_10_37_2632_0 & ~i_10_37_2633_0 & ~i_10_37_3277_0 & ~i_10_37_3467_0 & ~i_10_37_3850_0 & ~i_10_37_3858_0 & ~i_10_37_3889_0) | (~i_10_37_251_0 & i_10_37_1687_0 & ~i_10_37_2363_0 & ~i_10_37_3991_0 & ~i_10_37_4115_0));
endmodule



// Benchmark "kernel_10_38" written by ABC on Sun Jul 19 10:21:41 2020

module kernel_10_38 ( 
    i_10_38_125_0, i_10_38_172_0, i_10_38_173_0, i_10_38_174_0,
    i_10_38_175_0, i_10_38_222_0, i_10_38_224_0, i_10_38_269_0,
    i_10_38_393_0, i_10_38_394_0, i_10_38_405_0, i_10_38_409_0,
    i_10_38_410_0, i_10_38_413_0, i_10_38_429_0, i_10_38_430_0,
    i_10_38_431_0, i_10_38_433_0, i_10_38_439_0, i_10_38_440_0,
    i_10_38_445_0, i_10_38_447_0, i_10_38_460_0, i_10_38_462_0,
    i_10_38_566_0, i_10_38_957_0, i_10_38_1006_0, i_10_38_1241_0,
    i_10_38_1309_0, i_10_38_1448_0, i_10_38_1550_0, i_10_38_1556_0,
    i_10_38_1637_0, i_10_38_1649_0, i_10_38_1651_0, i_10_38_1652_0,
    i_10_38_1653_0, i_10_38_1654_0, i_10_38_1655_0, i_10_38_1823_0,
    i_10_38_1825_0, i_10_38_1826_0, i_10_38_2006_0, i_10_38_2351_0,
    i_10_38_2354_0, i_10_38_2355_0, i_10_38_2356_0, i_10_38_2357_0,
    i_10_38_2358_0, i_10_38_2366_0, i_10_38_2448_0, i_10_38_2458_0,
    i_10_38_2572_0, i_10_38_2629_0, i_10_38_2632_0, i_10_38_2681_0,
    i_10_38_2700_0, i_10_38_2705_0, i_10_38_2706_0, i_10_38_2707_0,
    i_10_38_2708_0, i_10_38_2716_0, i_10_38_2718_0, i_10_38_2721_0,
    i_10_38_2723_0, i_10_38_2725_0, i_10_38_2728_0, i_10_38_2730_0,
    i_10_38_2731_0, i_10_38_2732_0, i_10_38_2735_0, i_10_38_2832_0,
    i_10_38_2833_0, i_10_38_2834_0, i_10_38_2881_0, i_10_38_2884_0,
    i_10_38_2985_0, i_10_38_3076_0, i_10_38_3087_0, i_10_38_3091_0,
    i_10_38_3093_0, i_10_38_3094_0, i_10_38_3095_0, i_10_38_3155_0,
    i_10_38_3198_0, i_10_38_3281_0, i_10_38_3391_0, i_10_38_3408_0,
    i_10_38_3611_0, i_10_38_3612_0, i_10_38_3615_0, i_10_38_3811_0,
    i_10_38_3835_0, i_10_38_3838_0, i_10_38_3839_0, i_10_38_3853_0,
    i_10_38_4120_0, i_10_38_4126_0, i_10_38_4127_0, i_10_38_4128_0,
    o_10_38_0_0  );
  input  i_10_38_125_0, i_10_38_172_0, i_10_38_173_0, i_10_38_174_0,
    i_10_38_175_0, i_10_38_222_0, i_10_38_224_0, i_10_38_269_0,
    i_10_38_393_0, i_10_38_394_0, i_10_38_405_0, i_10_38_409_0,
    i_10_38_410_0, i_10_38_413_0, i_10_38_429_0, i_10_38_430_0,
    i_10_38_431_0, i_10_38_433_0, i_10_38_439_0, i_10_38_440_0,
    i_10_38_445_0, i_10_38_447_0, i_10_38_460_0, i_10_38_462_0,
    i_10_38_566_0, i_10_38_957_0, i_10_38_1006_0, i_10_38_1241_0,
    i_10_38_1309_0, i_10_38_1448_0, i_10_38_1550_0, i_10_38_1556_0,
    i_10_38_1637_0, i_10_38_1649_0, i_10_38_1651_0, i_10_38_1652_0,
    i_10_38_1653_0, i_10_38_1654_0, i_10_38_1655_0, i_10_38_1823_0,
    i_10_38_1825_0, i_10_38_1826_0, i_10_38_2006_0, i_10_38_2351_0,
    i_10_38_2354_0, i_10_38_2355_0, i_10_38_2356_0, i_10_38_2357_0,
    i_10_38_2358_0, i_10_38_2366_0, i_10_38_2448_0, i_10_38_2458_0,
    i_10_38_2572_0, i_10_38_2629_0, i_10_38_2632_0, i_10_38_2681_0,
    i_10_38_2700_0, i_10_38_2705_0, i_10_38_2706_0, i_10_38_2707_0,
    i_10_38_2708_0, i_10_38_2716_0, i_10_38_2718_0, i_10_38_2721_0,
    i_10_38_2723_0, i_10_38_2725_0, i_10_38_2728_0, i_10_38_2730_0,
    i_10_38_2731_0, i_10_38_2732_0, i_10_38_2735_0, i_10_38_2832_0,
    i_10_38_2833_0, i_10_38_2834_0, i_10_38_2881_0, i_10_38_2884_0,
    i_10_38_2985_0, i_10_38_3076_0, i_10_38_3087_0, i_10_38_3091_0,
    i_10_38_3093_0, i_10_38_3094_0, i_10_38_3095_0, i_10_38_3155_0,
    i_10_38_3198_0, i_10_38_3281_0, i_10_38_3391_0, i_10_38_3408_0,
    i_10_38_3611_0, i_10_38_3612_0, i_10_38_3615_0, i_10_38_3811_0,
    i_10_38_3835_0, i_10_38_3838_0, i_10_38_3839_0, i_10_38_3853_0,
    i_10_38_4120_0, i_10_38_4126_0, i_10_38_4127_0, i_10_38_4128_0;
  output o_10_38_0_0;
  assign o_10_38_0_0 = ~((~i_10_38_957_0 & ((~i_10_38_125_0 & ((~i_10_38_409_0 & ~i_10_38_433_0 & ~i_10_38_445_0 & ~i_10_38_1556_0 & ~i_10_38_1649_0 & ~i_10_38_2358_0 & ~i_10_38_2632_0 & ~i_10_38_3093_0 & ~i_10_38_3095_0 & ~i_10_38_3408_0 & ~i_10_38_3612_0) | (~i_10_38_462_0 & ~i_10_38_1550_0 & ~i_10_38_1825_0 & ~i_10_38_2728_0 & ~i_10_38_2884_0 & ~i_10_38_3198_0 & ~i_10_38_3391_0 & ~i_10_38_4120_0 & ~i_10_38_4128_0))) | (~i_10_38_462_0 & ((~i_10_38_430_0 & ~i_10_38_431_0 & ~i_10_38_1550_0 & ~i_10_38_1823_0 & ~i_10_38_2718_0 & ~i_10_38_2723_0 & ~i_10_38_2881_0 & ~i_10_38_3093_0 & ~i_10_38_3281_0) | (~i_10_38_440_0 & ~i_10_38_1649_0 & ~i_10_38_2716_0 & ~i_10_38_2884_0 & ~i_10_38_3198_0 & i_10_38_3838_0 & ~i_10_38_4128_0))) | (~i_10_38_3093_0 & ((i_10_38_1653_0 & ~i_10_38_3087_0 & ~i_10_38_3094_0) | (~i_10_38_2632_0 & ~i_10_38_2716_0 & i_10_38_2731_0 & ~i_10_38_2735_0 & ~i_10_38_3198_0 & ~i_10_38_3611_0 & ~i_10_38_3615_0))) | (~i_10_38_433_0 & i_10_38_462_0 & ~i_10_38_1550_0 & i_10_38_1651_0 & ~i_10_38_3198_0) | (i_10_38_1652_0 & i_10_38_2700_0 & ~i_10_38_3839_0) | (~i_10_38_429_0 & i_10_38_460_0 & ~i_10_38_1823_0 & ~i_10_38_2458_0 & ~i_10_38_2881_0 & ~i_10_38_3091_0 & ~i_10_38_3612_0 & ~i_10_38_4128_0))) | (~i_10_38_3095_0 & ((~i_10_38_175_0 & ~i_10_38_3093_0 & ((~i_10_38_393_0 & ~i_10_38_1241_0 & i_10_38_1825_0 & ~i_10_38_2458_0 & ~i_10_38_2718_0 & ~i_10_38_2985_0 & ~i_10_38_3087_0) | (i_10_38_1654_0 & ~i_10_38_2356_0 & ~i_10_38_3198_0 & ~i_10_38_3611_0))) | (~i_10_38_429_0 & (i_10_38_4127_0 | (i_10_38_1241_0 & ~i_10_38_2006_0 & ~i_10_38_2881_0 & ~i_10_38_3087_0 & ~i_10_38_3091_0 & ~i_10_38_3094_0))) | (~i_10_38_433_0 & ((~i_10_38_447_0 & ~i_10_38_460_0 & ~i_10_38_462_0 & ~i_10_38_1550_0 & i_10_38_1651_0 & ~i_10_38_2700_0) | (~i_10_38_439_0 & ~i_10_38_1823_0 & i_10_38_1825_0 & ~i_10_38_2006_0 & ~i_10_38_2723_0 & ~i_10_38_2728_0 & ~i_10_38_3838_0))) | (~i_10_38_445_0 & i_10_38_2357_0 & ~i_10_38_3087_0) | (~i_10_38_394_0 & ~i_10_38_566_0 & ~i_10_38_1309_0 & ~i_10_38_2458_0 & ~i_10_38_2629_0 & ~i_10_38_3391_0 & ~i_10_38_3408_0 & ~i_10_38_3611_0 & i_10_38_3838_0))) | (~i_10_38_393_0 & ((~i_10_38_433_0 & ~i_10_38_1550_0 & ~i_10_38_1826_0 & ~i_10_38_2006_0 & i_10_38_2354_0 & ~i_10_38_2681_0) | (~i_10_38_409_0 & ~i_10_38_1309_0 & ~i_10_38_2358_0 & ~i_10_38_2458_0 & ~i_10_38_2632_0 & ~i_10_38_2725_0 & ~i_10_38_2735_0 & ~i_10_38_2884_0 & ~i_10_38_3198_0 & ~i_10_38_3612_0))) | (~i_10_38_440_0 & ((i_10_38_224_0 & i_10_38_1825_0) | (~i_10_38_173_0 & ~i_10_38_429_0 & ~i_10_38_433_0 & ~i_10_38_445_0 & ~i_10_38_1823_0 & ~i_10_38_2884_0 & ~i_10_38_3198_0 & ~i_10_38_3838_0 & ~i_10_38_4120_0))) | (~i_10_38_429_0 & ((i_10_38_1655_0 & i_10_38_2354_0 & ~i_10_38_2881_0) | (i_10_38_2718_0 & i_10_38_2731_0 & ~i_10_38_2884_0 & ~i_10_38_3391_0 & ~i_10_38_3612_0))) | (~i_10_38_431_0 & ((~i_10_38_433_0 & ((~i_10_38_430_0 & i_10_38_1823_0 & ~i_10_38_1826_0 & ~i_10_38_2358_0 & ~i_10_38_3087_0 & ~i_10_38_3094_0 & ~i_10_38_2448_0 & ~i_10_38_2632_0) | (i_10_38_2448_0 & ~i_10_38_2884_0 & ~i_10_38_3198_0 & i_10_38_3611_0))) | (~i_10_38_1309_0 & ~i_10_38_1823_0 & ~i_10_38_2728_0 & ~i_10_38_3087_0 & ~i_10_38_3198_0 & i_10_38_3853_0))) | (~i_10_38_445_0 & ((~i_10_38_2730_0 & i_10_38_2731_0 & ~i_10_38_3091_0 & ~i_10_38_3391_0 & ~i_10_38_3835_0) | (~i_10_38_172_0 & ~i_10_38_462_0 & ~i_10_38_1309_0 & i_10_38_1649_0 & ~i_10_38_3839_0))) | (~i_10_38_1550_0 & ((i_10_38_1652_0 & i_10_38_2705_0) | (i_10_38_460_0 & ~i_10_38_462_0 & i_10_38_1651_0 & i_10_38_2700_0 & ~i_10_38_2728_0))) | (~i_10_38_462_0 & ((i_10_38_173_0 & ~i_10_38_2354_0 & ~i_10_38_2458_0 & ~i_10_38_3094_0) | (i_10_38_1651_0 & ~i_10_38_1823_0 & ~i_10_38_2723_0 & ~i_10_38_2884_0 & ~i_10_38_3612_0 & ~i_10_38_3838_0 & ~i_10_38_3853_0))) | (i_10_38_1652_0 & ((~i_10_38_1823_0 & i_10_38_2700_0) | (~i_10_38_2458_0 & i_10_38_2718_0 & i_10_38_2721_0 & ~i_10_38_4128_0))) | (~i_10_38_3087_0 & ((~i_10_38_2358_0 & i_10_38_2728_0 & i_10_38_2732_0 & ~i_10_38_3091_0 & ~i_10_38_3094_0) | (~i_10_38_394_0 & i_10_38_2832_0 & i_10_38_2833_0 & ~i_10_38_3198_0))) | (~i_10_38_3198_0 & ((i_10_38_409_0 & i_10_38_462_0 & ~i_10_38_2728_0) | (i_10_38_172_0 & i_10_38_3611_0 & ~i_10_38_4126_0))) | (i_10_38_172_0 & ((i_10_38_1309_0 & ~i_10_38_1652_0) | (i_10_38_175_0 & ~i_10_38_409_0 & ~i_10_38_4128_0))) | (i_10_38_410_0 & i_10_38_1655_0 & ~i_10_38_2355_0) | (~i_10_38_1309_0 & ~i_10_38_2735_0 & i_10_38_2834_0) | (i_10_38_2706_0 & ~i_10_38_3093_0) | (i_10_38_1653_0 & i_10_38_1654_0 & ~i_10_38_2632_0 & ~i_10_38_2832_0 & ~i_10_38_3611_0) | (i_10_38_1649_0 & i_10_38_2700_0 & i_10_38_3838_0) | (i_10_38_2351_0 & ~i_10_38_2721_0 & ~i_10_38_3281_0 & ~i_10_38_3838_0));
endmodule



// Benchmark "kernel_10_39" written by ABC on Sun Jul 19 10:21:43 2020

module kernel_10_39 ( 
    i_10_39_172_0, i_10_39_174_0, i_10_39_176_0, i_10_39_260_0,
    i_10_39_268_0, i_10_39_269_0, i_10_39_284_0, i_10_39_328_0,
    i_10_39_329_0, i_10_39_394_0, i_10_39_408_0, i_10_39_409_0,
    i_10_39_410_0, i_10_39_425_0, i_10_39_436_0, i_10_39_510_0,
    i_10_39_514_0, i_10_39_794_0, i_10_39_796_0, i_10_39_797_0,
    i_10_39_798_0, i_10_39_799_0, i_10_39_800_0, i_10_39_1006_0,
    i_10_39_1029_0, i_10_39_1261_0, i_10_39_1264_0, i_10_39_1308_0,
    i_10_39_1309_0, i_10_39_1438_0, i_10_39_1439_0, i_10_39_1546_0,
    i_10_39_1628_0, i_10_39_1651_0, i_10_39_1655_0, i_10_39_1691_0,
    i_10_39_1727_0, i_10_39_1821_0, i_10_39_1822_0, i_10_39_1823_0,
    i_10_39_1825_0, i_10_39_1912_0, i_10_39_1996_0, i_10_39_2254_0,
    i_10_39_2364_0, i_10_39_2451_0, i_10_39_2461_0, i_10_39_2463_0,
    i_10_39_2470_0, i_10_39_2473_0, i_10_39_2573_0, i_10_39_2634_0,
    i_10_39_2635_0, i_10_39_2636_0, i_10_39_2659_0, i_10_39_2704_0,
    i_10_39_2717_0, i_10_39_2720_0, i_10_39_2722_0, i_10_39_2723_0,
    i_10_39_2725_0, i_10_39_2730_0, i_10_39_2731_0, i_10_39_2826_0,
    i_10_39_2830_0, i_10_39_2832_0, i_10_39_2884_0, i_10_39_2885_0,
    i_10_39_3077_0, i_10_39_3087_0, i_10_39_3088_0, i_10_39_3153_0,
    i_10_39_3195_0, i_10_39_3196_0, i_10_39_3197_0, i_10_39_3200_0,
    i_10_39_3280_0, i_10_39_3329_0, i_10_39_3388_0, i_10_39_3389_0,
    i_10_39_3409_0, i_10_39_3473_0, i_10_39_3586_0, i_10_39_3610_0,
    i_10_39_3611_0, i_10_39_3614_0, i_10_39_3616_0, i_10_39_3648_0,
    i_10_39_3651_0, i_10_39_3652_0, i_10_39_3860_0, i_10_39_4126_0,
    i_10_39_4271_0, i_10_39_4289_0, i_10_39_4564_0, i_10_39_4565_0,
    i_10_39_4567_0, i_10_39_4568_0, i_10_39_4570_0, i_10_39_4571_0,
    o_10_39_0_0  );
  input  i_10_39_172_0, i_10_39_174_0, i_10_39_176_0, i_10_39_260_0,
    i_10_39_268_0, i_10_39_269_0, i_10_39_284_0, i_10_39_328_0,
    i_10_39_329_0, i_10_39_394_0, i_10_39_408_0, i_10_39_409_0,
    i_10_39_410_0, i_10_39_425_0, i_10_39_436_0, i_10_39_510_0,
    i_10_39_514_0, i_10_39_794_0, i_10_39_796_0, i_10_39_797_0,
    i_10_39_798_0, i_10_39_799_0, i_10_39_800_0, i_10_39_1006_0,
    i_10_39_1029_0, i_10_39_1261_0, i_10_39_1264_0, i_10_39_1308_0,
    i_10_39_1309_0, i_10_39_1438_0, i_10_39_1439_0, i_10_39_1546_0,
    i_10_39_1628_0, i_10_39_1651_0, i_10_39_1655_0, i_10_39_1691_0,
    i_10_39_1727_0, i_10_39_1821_0, i_10_39_1822_0, i_10_39_1823_0,
    i_10_39_1825_0, i_10_39_1912_0, i_10_39_1996_0, i_10_39_2254_0,
    i_10_39_2364_0, i_10_39_2451_0, i_10_39_2461_0, i_10_39_2463_0,
    i_10_39_2470_0, i_10_39_2473_0, i_10_39_2573_0, i_10_39_2634_0,
    i_10_39_2635_0, i_10_39_2636_0, i_10_39_2659_0, i_10_39_2704_0,
    i_10_39_2717_0, i_10_39_2720_0, i_10_39_2722_0, i_10_39_2723_0,
    i_10_39_2725_0, i_10_39_2730_0, i_10_39_2731_0, i_10_39_2826_0,
    i_10_39_2830_0, i_10_39_2832_0, i_10_39_2884_0, i_10_39_2885_0,
    i_10_39_3077_0, i_10_39_3087_0, i_10_39_3088_0, i_10_39_3153_0,
    i_10_39_3195_0, i_10_39_3196_0, i_10_39_3197_0, i_10_39_3200_0,
    i_10_39_3280_0, i_10_39_3329_0, i_10_39_3388_0, i_10_39_3389_0,
    i_10_39_3409_0, i_10_39_3473_0, i_10_39_3586_0, i_10_39_3610_0,
    i_10_39_3611_0, i_10_39_3614_0, i_10_39_3616_0, i_10_39_3648_0,
    i_10_39_3651_0, i_10_39_3652_0, i_10_39_3860_0, i_10_39_4126_0,
    i_10_39_4271_0, i_10_39_4289_0, i_10_39_4564_0, i_10_39_4565_0,
    i_10_39_4567_0, i_10_39_4568_0, i_10_39_4570_0, i_10_39_4571_0;
  output o_10_39_0_0;
  assign o_10_39_0_0 = ~((i_10_39_172_0 & ((~i_10_39_1821_0 & ~i_10_39_4126_0) | (i_10_39_1822_0 & ~i_10_39_3586_0 & ~i_10_39_3611_0 & ~i_10_39_3651_0 & ~i_10_39_4568_0))) | (~i_10_39_260_0 & ((~i_10_39_1006_0 & ~i_10_39_1821_0 & ~i_10_39_2470_0 & ~i_10_39_2473_0 & ~i_10_39_2659_0 & ~i_10_39_2722_0 & ~i_10_39_2885_0 & ~i_10_39_3088_0 & ~i_10_39_3195_0 & ~i_10_39_3197_0) | (~i_10_39_268_0 & ~i_10_39_1029_0 & ~i_10_39_1823_0 & ~i_10_39_2451_0 & ~i_10_39_2573_0 & ~i_10_39_2884_0 & ~i_10_39_3087_0 & ~i_10_39_3610_0 & ~i_10_39_3648_0 & ~i_10_39_4564_0))) | (~i_10_39_269_0 & ((~i_10_39_1438_0 & i_10_39_2722_0 & ~i_10_39_3196_0 & ~i_10_39_3648_0) | (~i_10_39_268_0 & ~i_10_39_408_0 & ~i_10_39_799_0 & i_10_39_1825_0 & ~i_10_39_3087_0 & i_10_39_3388_0 & ~i_10_39_3651_0))) | (~i_10_39_284_0 & ((~i_10_39_799_0 & ~i_10_39_1439_0 & i_10_39_2730_0 & ~i_10_39_3195_0 & ~i_10_39_3388_0 & ~i_10_39_3610_0) | (i_10_39_1821_0 & i_10_39_1822_0 & i_10_39_1912_0 & ~i_10_39_2470_0 & i_10_39_2659_0 & ~i_10_39_3087_0 & ~i_10_39_4289_0))) | (~i_10_39_436_0 & ((~i_10_39_799_0 & ~i_10_39_1823_0 & ~i_10_39_2573_0 & ~i_10_39_2722_0 & ~i_10_39_2884_0 & i_10_39_3389_0 & ~i_10_39_3611_0) | (~i_10_39_268_0 & ~i_10_39_1029_0 & ~i_10_39_1628_0 & ~i_10_39_2364_0 & i_10_39_2636_0 & ~i_10_39_2659_0 & ~i_10_39_2832_0 & ~i_10_39_3586_0 & ~i_10_39_3860_0))) | (i_10_39_799_0 & (i_10_39_1912_0 | (~i_10_39_3280_0 & i_10_39_3616_0 & ~i_10_39_3860_0 & ~i_10_39_4567_0))) | (~i_10_39_1308_0 & ((~i_10_39_1438_0 & ~i_10_39_1822_0 & ~i_10_39_1823_0 & ~i_10_39_3087_0) | (i_10_39_1825_0 & ~i_10_39_3196_0 & i_10_39_3610_0))) | (~i_10_39_1546_0 & ((~i_10_39_1823_0 & ~i_10_39_1825_0 & i_10_39_3388_0) | (i_10_39_796_0 & ~i_10_39_1438_0 & ~i_10_39_1439_0 & ~i_10_39_2885_0 & ~i_10_39_3195_0 & ~i_10_39_3648_0))) | (~i_10_39_1439_0 & ~i_10_39_3195_0 & ((~i_10_39_1821_0 & ~i_10_39_1822_0 & ~i_10_39_3196_0 & ~i_10_39_3280_0 & ~i_10_39_3610_0) | (i_10_39_3389_0 & ~i_10_39_3860_0))) | (~i_10_39_3088_0 & ((~i_10_39_2451_0 & ((~i_10_39_268_0 & ((~i_10_39_794_0 & ~i_10_39_797_0 & ~i_10_39_1006_0 & ~i_10_39_1309_0 & ~i_10_39_1821_0 & ~i_10_39_2573_0) | (~i_10_39_172_0 & ~i_10_39_176_0 & ~i_10_39_1628_0 & ~i_10_39_1651_0 & ~i_10_39_2473_0 & ~i_10_39_2720_0 & ~i_10_39_2730_0 & i_10_39_3200_0 & ~i_10_39_3610_0))) | (~i_10_39_1006_0 & ~i_10_39_3087_0 & ((~i_10_39_1628_0 & i_10_39_1825_0 & i_10_39_3616_0) | (~i_10_39_1309_0 & ~i_10_39_1651_0 & ~i_10_39_2884_0 & ~i_10_39_3197_0 & ~i_10_39_3648_0))))) | (i_10_39_514_0 & ~i_10_39_1029_0 & ~i_10_39_1438_0 & ~i_10_39_3196_0) | (i_10_39_798_0 & ~i_10_39_2473_0 & ~i_10_39_3611_0) | (~i_10_39_394_0 & i_10_39_436_0 & ~i_10_39_798_0 & ~i_10_39_1823_0 & i_10_39_2473_0 & i_10_39_2731_0 & i_10_39_3610_0 & ~i_10_39_3614_0 & ~i_10_39_4271_0))) | (~i_10_39_1438_0 & ((~i_10_39_1912_0 & ~i_10_39_2451_0 & i_10_39_2830_0 & ~i_10_39_3473_0) | (~i_10_39_1821_0 & ~i_10_39_1822_0 & ~i_10_39_3586_0 & ~i_10_39_3614_0 & ~i_10_39_4567_0))) | (i_10_39_1822_0 & ((i_10_39_2722_0 & ~i_10_39_2731_0 & i_10_39_3610_0) | (~i_10_39_1309_0 & ~i_10_39_1823_0 & ~i_10_39_2884_0 & ~i_10_39_2885_0 & i_10_39_3196_0 & ~i_10_39_4567_0))) | (~i_10_39_2473_0 & ((i_10_39_2730_0 & i_10_39_2731_0 & ~i_10_39_3200_0 & ~i_10_39_4126_0) | (i_10_39_1308_0 & i_10_39_1309_0 & i_10_39_2832_0 & ~i_10_39_4567_0 & ~i_10_39_4568_0))) | (i_10_39_4564_0 & ((~i_10_39_3196_0 & i_10_39_3648_0 & i_10_39_4289_0) | (i_10_39_1651_0 & ~i_10_39_3610_0 & ~i_10_39_3648_0 & ~i_10_39_4565_0))) | (~i_10_39_268_0 & ~i_10_39_1628_0 & i_10_39_2725_0) | (i_10_39_797_0 & ~i_10_39_2885_0 & i_10_39_3611_0 & ~i_10_39_3614_0) | (~i_10_39_1655_0 & i_10_39_2364_0 & ~i_10_39_2470_0 & i_10_39_3652_0));
endmodule



// Benchmark "kernel_10_40" written by ABC on Sun Jul 19 10:21:44 2020

module kernel_10_40 ( 
    i_10_40_118_0, i_10_40_171_0, i_10_40_172_0, i_10_40_175_0,
    i_10_40_216_0, i_10_40_217_0, i_10_40_218_0, i_10_40_220_0,
    i_10_40_221_0, i_10_40_224_0, i_10_40_243_0, i_10_40_244_0,
    i_10_40_245_0, i_10_40_280_0, i_10_40_329_0, i_10_40_390_0,
    i_10_40_405_0, i_10_40_406_0, i_10_40_409_0, i_10_40_447_0,
    i_10_40_711_0, i_10_40_712_0, i_10_40_799_0, i_10_40_898_0,
    i_10_40_967_0, i_10_40_991_0, i_10_40_1029_0, i_10_40_1030_0,
    i_10_40_1233_0, i_10_40_1241_0, i_10_40_1306_0, i_10_40_1434_0,
    i_10_40_1441_0, i_10_40_1648_0, i_10_40_1649_0, i_10_40_1651_0,
    i_10_40_1683_0, i_10_40_1821_0, i_10_40_1824_0, i_10_40_1990_0,
    i_10_40_2351_0, i_10_40_2353_0, i_10_40_2354_0, i_10_40_2363_0,
    i_10_40_2451_0, i_10_40_2473_0, i_10_40_2628_0, i_10_40_2632_0,
    i_10_40_2635_0, i_10_40_2654_0, i_10_40_2656_0, i_10_40_2709_0,
    i_10_40_2717_0, i_10_40_2718_0, i_10_40_2735_0, i_10_40_2826_0,
    i_10_40_2827_0, i_10_40_2831_0, i_10_40_2832_0, i_10_40_2833_0,
    i_10_40_2834_0, i_10_40_2920_0, i_10_40_2921_0, i_10_40_2924_0,
    i_10_40_2986_0, i_10_40_3034_0, i_10_40_3151_0, i_10_40_3152_0,
    i_10_40_3153_0, i_10_40_3162_0, i_10_40_3163_0, i_10_40_3198_0,
    i_10_40_3322_0, i_10_40_3329_0, i_10_40_3389_0, i_10_40_3406_0,
    i_10_40_3466_0, i_10_40_3472_0, i_10_40_3547_0, i_10_40_3610_0,
    i_10_40_3611_0, i_10_40_3613_0, i_10_40_3647_0, i_10_40_3733_0,
    i_10_40_3782_0, i_10_40_3837_0, i_10_40_3839_0, i_10_40_3856_0,
    i_10_40_3912_0, i_10_40_3983_0, i_10_40_4113_0, i_10_40_4114_0,
    i_10_40_4115_0, i_10_40_4116_0, i_10_40_4117_0, i_10_40_4129_0,
    i_10_40_4271_0, i_10_40_4287_0, i_10_40_4288_0, i_10_40_4289_0,
    o_10_40_0_0  );
  input  i_10_40_118_0, i_10_40_171_0, i_10_40_172_0, i_10_40_175_0,
    i_10_40_216_0, i_10_40_217_0, i_10_40_218_0, i_10_40_220_0,
    i_10_40_221_0, i_10_40_224_0, i_10_40_243_0, i_10_40_244_0,
    i_10_40_245_0, i_10_40_280_0, i_10_40_329_0, i_10_40_390_0,
    i_10_40_405_0, i_10_40_406_0, i_10_40_409_0, i_10_40_447_0,
    i_10_40_711_0, i_10_40_712_0, i_10_40_799_0, i_10_40_898_0,
    i_10_40_967_0, i_10_40_991_0, i_10_40_1029_0, i_10_40_1030_0,
    i_10_40_1233_0, i_10_40_1241_0, i_10_40_1306_0, i_10_40_1434_0,
    i_10_40_1441_0, i_10_40_1648_0, i_10_40_1649_0, i_10_40_1651_0,
    i_10_40_1683_0, i_10_40_1821_0, i_10_40_1824_0, i_10_40_1990_0,
    i_10_40_2351_0, i_10_40_2353_0, i_10_40_2354_0, i_10_40_2363_0,
    i_10_40_2451_0, i_10_40_2473_0, i_10_40_2628_0, i_10_40_2632_0,
    i_10_40_2635_0, i_10_40_2654_0, i_10_40_2656_0, i_10_40_2709_0,
    i_10_40_2717_0, i_10_40_2718_0, i_10_40_2735_0, i_10_40_2826_0,
    i_10_40_2827_0, i_10_40_2831_0, i_10_40_2832_0, i_10_40_2833_0,
    i_10_40_2834_0, i_10_40_2920_0, i_10_40_2921_0, i_10_40_2924_0,
    i_10_40_2986_0, i_10_40_3034_0, i_10_40_3151_0, i_10_40_3152_0,
    i_10_40_3153_0, i_10_40_3162_0, i_10_40_3163_0, i_10_40_3198_0,
    i_10_40_3322_0, i_10_40_3329_0, i_10_40_3389_0, i_10_40_3406_0,
    i_10_40_3466_0, i_10_40_3472_0, i_10_40_3547_0, i_10_40_3610_0,
    i_10_40_3611_0, i_10_40_3613_0, i_10_40_3647_0, i_10_40_3733_0,
    i_10_40_3782_0, i_10_40_3837_0, i_10_40_3839_0, i_10_40_3856_0,
    i_10_40_3912_0, i_10_40_3983_0, i_10_40_4113_0, i_10_40_4114_0,
    i_10_40_4115_0, i_10_40_4116_0, i_10_40_4117_0, i_10_40_4129_0,
    i_10_40_4271_0, i_10_40_4287_0, i_10_40_4288_0, i_10_40_4289_0;
  output o_10_40_0_0;
  assign o_10_40_0_0 = ~((~i_10_40_216_0 & ((~i_10_40_244_0 & ~i_10_40_409_0 & ~i_10_40_898_0 & ~i_10_40_2920_0 & ~i_10_40_3162_0 & ~i_10_40_3163_0 & ~i_10_40_3611_0 & ~i_10_40_3856_0) | (~i_10_40_171_0 & ~i_10_40_217_0 & ~i_10_40_218_0 & ~i_10_40_406_0 & ~i_10_40_712_0 & ~i_10_40_2834_0 & ~i_10_40_2921_0 & ~i_10_40_3613_0 & ~i_10_40_3837_0 & ~i_10_40_3912_0))) | (~i_10_40_2833_0 & ((~i_10_40_409_0 & ((~i_10_40_217_0 & ((~i_10_40_1651_0 & ~i_10_40_2656_0) | (~i_10_40_244_0 & ~i_10_40_1030_0 & i_10_40_2628_0 & ~i_10_40_2920_0 & i_10_40_4114_0))) | (~i_10_40_175_0 & ~i_10_40_218_0 & ~i_10_40_406_0 & ~i_10_40_1649_0 & ~i_10_40_1683_0 & i_10_40_2628_0 & ~i_10_40_2826_0))) | (~i_10_40_2656_0 & ((~i_10_40_243_0 & ~i_10_40_245_0 & ~i_10_40_712_0 & ~i_10_40_2635_0 & ~i_10_40_3406_0 & ~i_10_40_3610_0) | (~i_10_40_898_0 & ~i_10_40_1648_0 & i_10_40_1651_0 & ~i_10_40_2921_0 & i_10_40_3613_0 & ~i_10_40_4113_0))) | (~i_10_40_220_0 & ~i_10_40_1441_0 & i_10_40_2831_0 & ~i_10_40_3611_0))) | (~i_10_40_224_0 & ~i_10_40_3198_0 & ((~i_10_40_243_0 & ~i_10_40_245_0 & ~i_10_40_280_0 & ~i_10_40_898_0 & ~i_10_40_3162_0 & ~i_10_40_3163_0 & ~i_10_40_1683_0 & i_10_40_2635_0) | (~i_10_40_175_0 & ~i_10_40_220_0 & ~i_10_40_244_0 & ~i_10_40_991_0 & ~i_10_40_1306_0 & ~i_10_40_1441_0 & ~i_10_40_1649_0 & ~i_10_40_2826_0 & ~i_10_40_3837_0 & ~i_10_40_4288_0))) | (~i_10_40_175_0 & ((~i_10_40_172_0 & ~i_10_40_1648_0 & ~i_10_40_1649_0 & ~i_10_40_1651_0 & i_10_40_3389_0) | (~i_10_40_218_0 & ~i_10_40_220_0 & ~i_10_40_712_0 & ~i_10_40_2363_0 & ~i_10_40_3163_0 & ~i_10_40_3406_0 & ~i_10_40_3912_0 & ~i_10_40_4117_0))) | (~i_10_40_218_0 & ~i_10_40_3912_0 & ((~i_10_40_221_0 & ~i_10_40_243_0 & ~i_10_40_405_0 & ~i_10_40_898_0 & ~i_10_40_1306_0 & ~i_10_40_1648_0 & ~i_10_40_1990_0 & ~i_10_40_2921_0 & ~i_10_40_3613_0) | (~i_10_40_711_0 & ~i_10_40_1030_0 & ~i_10_40_2831_0 & ~i_10_40_3782_0 & ~i_10_40_4114_0 & ~i_10_40_4115_0 & i_10_40_4288_0))) | (~i_10_40_220_0 & ((~i_10_40_1651_0 & ~i_10_40_1821_0 & ~i_10_40_2717_0 & i_10_40_2831_0 & ~i_10_40_3163_0 & ~i_10_40_3782_0) | (~i_10_40_221_0 & ~i_10_40_1649_0 & i_10_40_2632_0 & ~i_10_40_4113_0 & ~i_10_40_4115_0 & ~i_10_40_4129_0))) | (~i_10_40_712_0 & ((~i_10_40_711_0 & i_10_40_1306_0 & ~i_10_40_1441_0 & i_10_40_2656_0 & ~i_10_40_2832_0 & ~i_10_40_3983_0) | (~i_10_40_405_0 & ~i_10_40_2451_0 & ~i_10_40_2635_0 & ~i_10_40_2924_0 & ~i_10_40_3162_0 & ~i_10_40_3163_0 & i_10_40_4116_0 & i_10_40_4117_0 & ~i_10_40_4289_0))) | (~i_10_40_991_0 & ~i_10_40_1651_0 & ((~i_10_40_221_0 & ~i_10_40_967_0 & ~i_10_40_1648_0 & ~i_10_40_1821_0 & i_10_40_2656_0 & ~i_10_40_2921_0) | (~i_10_40_898_0 & ~i_10_40_2363_0 & ~i_10_40_3162_0 & ~i_10_40_3611_0 & ~i_10_40_3839_0 & ~i_10_40_4114_0 & ~i_10_40_4116_0))) | (i_10_40_2834_0 & ((~i_10_40_2831_0 & ~i_10_40_2986_0 & ~i_10_40_3406_0 & i_10_40_3613_0) | (~i_10_40_2832_0 & i_10_40_3198_0 & ~i_10_40_4129_0))));
endmodule



// Benchmark "kernel_10_41" written by ABC on Sun Jul 19 10:21:45 2020

module kernel_10_41 ( 
    i_10_41_27_0, i_10_41_68_0, i_10_41_86_0, i_10_41_103_0, i_10_41_176_0,
    i_10_41_178_0, i_10_41_215_0, i_10_41_224_0, i_10_41_248_0,
    i_10_41_425_0, i_10_41_562_0, i_10_41_565_0, i_10_41_566_0,
    i_10_41_586_0, i_10_41_824_0, i_10_41_960_0, i_10_41_989_0,
    i_10_41_1000_0, i_10_41_1001_0, i_10_41_1004_0, i_10_41_1101_0,
    i_10_41_1223_0, i_10_41_1238_0, i_10_41_1240_0, i_10_41_1349_0,
    i_10_41_1367_0, i_10_41_1439_0, i_10_41_1544_0, i_10_41_1547_0,
    i_10_41_1583_0, i_10_41_1651_0, i_10_41_1652_0, i_10_41_1687_0,
    i_10_41_1715_0, i_10_41_1766_0, i_10_41_1772_0, i_10_41_1778_0,
    i_10_41_1988_0, i_10_41_1991_0, i_10_41_1997_0, i_10_41_2000_0,
    i_10_41_2006_0, i_10_41_2023_0, i_10_41_2033_0, i_10_41_2348_0,
    i_10_41_2449_0, i_10_41_2453_0, i_10_41_2509_0, i_10_41_2510_0,
    i_10_41_2539_0, i_10_41_2567_0, i_10_41_2570_0, i_10_41_2571_0,
    i_10_41_2609_0, i_10_41_2636_0, i_10_41_2641_0, i_10_41_2644_0,
    i_10_41_2645_0, i_10_41_2720_0, i_10_41_2744_0, i_10_41_2834_0,
    i_10_41_2848_0, i_10_41_2849_0, i_10_41_2851_0, i_10_41_2966_0,
    i_10_41_2968_0, i_10_41_2999_0, i_10_41_3002_0, i_10_41_3041_0,
    i_10_41_3071_0, i_10_41_3074_0, i_10_41_3230_0, i_10_41_3238_0,
    i_10_41_3299_0, i_10_41_3307_0, i_10_41_3308_0, i_10_41_3409_0,
    i_10_41_3470_0, i_10_41_3506_0, i_10_41_3544_0, i_10_41_3545_0,
    i_10_41_3611_0, i_10_41_3797_0, i_10_41_3852_0, i_10_41_3853_0,
    i_10_41_3856_0, i_10_41_3923_0, i_10_41_3944_0, i_10_41_3989_0,
    i_10_41_4027_0, i_10_41_4129_0, i_10_41_4130_0, i_10_41_4148_0,
    i_10_41_4175_0, i_10_41_4217_0, i_10_41_4237_0, i_10_41_4238_0,
    i_10_41_4436_0, i_10_41_4461_0, i_10_41_4463_0,
    o_10_41_0_0  );
  input  i_10_41_27_0, i_10_41_68_0, i_10_41_86_0, i_10_41_103_0,
    i_10_41_176_0, i_10_41_178_0, i_10_41_215_0, i_10_41_224_0,
    i_10_41_248_0, i_10_41_425_0, i_10_41_562_0, i_10_41_565_0,
    i_10_41_566_0, i_10_41_586_0, i_10_41_824_0, i_10_41_960_0,
    i_10_41_989_0, i_10_41_1000_0, i_10_41_1001_0, i_10_41_1004_0,
    i_10_41_1101_0, i_10_41_1223_0, i_10_41_1238_0, i_10_41_1240_0,
    i_10_41_1349_0, i_10_41_1367_0, i_10_41_1439_0, i_10_41_1544_0,
    i_10_41_1547_0, i_10_41_1583_0, i_10_41_1651_0, i_10_41_1652_0,
    i_10_41_1687_0, i_10_41_1715_0, i_10_41_1766_0, i_10_41_1772_0,
    i_10_41_1778_0, i_10_41_1988_0, i_10_41_1991_0, i_10_41_1997_0,
    i_10_41_2000_0, i_10_41_2006_0, i_10_41_2023_0, i_10_41_2033_0,
    i_10_41_2348_0, i_10_41_2449_0, i_10_41_2453_0, i_10_41_2509_0,
    i_10_41_2510_0, i_10_41_2539_0, i_10_41_2567_0, i_10_41_2570_0,
    i_10_41_2571_0, i_10_41_2609_0, i_10_41_2636_0, i_10_41_2641_0,
    i_10_41_2644_0, i_10_41_2645_0, i_10_41_2720_0, i_10_41_2744_0,
    i_10_41_2834_0, i_10_41_2848_0, i_10_41_2849_0, i_10_41_2851_0,
    i_10_41_2966_0, i_10_41_2968_0, i_10_41_2999_0, i_10_41_3002_0,
    i_10_41_3041_0, i_10_41_3071_0, i_10_41_3074_0, i_10_41_3230_0,
    i_10_41_3238_0, i_10_41_3299_0, i_10_41_3307_0, i_10_41_3308_0,
    i_10_41_3409_0, i_10_41_3470_0, i_10_41_3506_0, i_10_41_3544_0,
    i_10_41_3545_0, i_10_41_3611_0, i_10_41_3797_0, i_10_41_3852_0,
    i_10_41_3853_0, i_10_41_3856_0, i_10_41_3923_0, i_10_41_3944_0,
    i_10_41_3989_0, i_10_41_4027_0, i_10_41_4129_0, i_10_41_4130_0,
    i_10_41_4148_0, i_10_41_4175_0, i_10_41_4217_0, i_10_41_4237_0,
    i_10_41_4238_0, i_10_41_4436_0, i_10_41_4461_0, i_10_41_4463_0;
  output o_10_41_0_0;
  assign o_10_41_0_0 = 0;
endmodule



// Benchmark "kernel_10_42" written by ABC on Sun Jul 19 10:21:46 2020

module kernel_10_42 ( 
    i_10_42_30_0, i_10_42_34_0, i_10_42_117_0, i_10_42_256_0,
    i_10_42_260_0, i_10_42_390_0, i_10_42_391_0, i_10_42_395_0,
    i_10_42_565_0, i_10_42_714_0, i_10_42_717_0, i_10_42_800_0,
    i_10_42_954_0, i_10_42_955_0, i_10_42_956_0, i_10_42_957_0,
    i_10_42_958_0, i_10_42_959_0, i_10_42_1030_0, i_10_42_1235_0,
    i_10_42_1245_0, i_10_42_1366_0, i_10_42_1439_0, i_10_42_1445_0,
    i_10_42_1450_0, i_10_42_1576_0, i_10_42_1579_0, i_10_42_1582_0,
    i_10_42_1619_0, i_10_42_1653_0, i_10_42_1691_0, i_10_42_1823_0,
    i_10_42_1826_0, i_10_42_2029_0, i_10_42_2030_0, i_10_42_2086_0,
    i_10_42_2197_0, i_10_42_2200_0, i_10_42_2201_0, i_10_42_2352_0,
    i_10_42_2353_0, i_10_42_2357_0, i_10_42_2383_0, i_10_42_2470_0,
    i_10_42_2536_0, i_10_42_2608_0, i_10_42_2614_0, i_10_42_2615_0,
    i_10_42_2632_0, i_10_42_2705_0, i_10_42_2707_0, i_10_42_2725_0,
    i_10_42_2869_0, i_10_42_3037_0, i_10_42_3039_0, i_10_42_3072_0,
    i_10_42_3196_0, i_10_42_3201_0, i_10_42_3202_0, i_10_42_3270_0,
    i_10_42_3391_0, i_10_42_3408_0, i_10_42_3469_0, i_10_42_3590_0,
    i_10_42_3612_0, i_10_42_3616_0, i_10_42_3617_0, i_10_42_3645_0,
    i_10_42_3646_0, i_10_42_3647_0, i_10_42_3649_0, i_10_42_3650_0,
    i_10_42_3651_0, i_10_42_3652_0, i_10_42_3653_0, i_10_42_3726_0,
    i_10_42_3729_0, i_10_42_3783_0, i_10_42_3784_0, i_10_42_3785_0,
    i_10_42_3786_0, i_10_42_3787_0, i_10_42_3788_0, i_10_42_3811_0,
    i_10_42_3837_0, i_10_42_3843_0, i_10_42_3844_0, i_10_42_3847_0,
    i_10_42_3856_0, i_10_42_3857_0, i_10_42_3914_0, i_10_42_4012_0,
    i_10_42_4116_0, i_10_42_4117_0, i_10_42_4118_0, i_10_42_4119_0,
    i_10_42_4120_0, i_10_42_4267_0, i_10_42_4564_0, i_10_42_4565_0,
    o_10_42_0_0  );
  input  i_10_42_30_0, i_10_42_34_0, i_10_42_117_0, i_10_42_256_0,
    i_10_42_260_0, i_10_42_390_0, i_10_42_391_0, i_10_42_395_0,
    i_10_42_565_0, i_10_42_714_0, i_10_42_717_0, i_10_42_800_0,
    i_10_42_954_0, i_10_42_955_0, i_10_42_956_0, i_10_42_957_0,
    i_10_42_958_0, i_10_42_959_0, i_10_42_1030_0, i_10_42_1235_0,
    i_10_42_1245_0, i_10_42_1366_0, i_10_42_1439_0, i_10_42_1445_0,
    i_10_42_1450_0, i_10_42_1576_0, i_10_42_1579_0, i_10_42_1582_0,
    i_10_42_1619_0, i_10_42_1653_0, i_10_42_1691_0, i_10_42_1823_0,
    i_10_42_1826_0, i_10_42_2029_0, i_10_42_2030_0, i_10_42_2086_0,
    i_10_42_2197_0, i_10_42_2200_0, i_10_42_2201_0, i_10_42_2352_0,
    i_10_42_2353_0, i_10_42_2357_0, i_10_42_2383_0, i_10_42_2470_0,
    i_10_42_2536_0, i_10_42_2608_0, i_10_42_2614_0, i_10_42_2615_0,
    i_10_42_2632_0, i_10_42_2705_0, i_10_42_2707_0, i_10_42_2725_0,
    i_10_42_2869_0, i_10_42_3037_0, i_10_42_3039_0, i_10_42_3072_0,
    i_10_42_3196_0, i_10_42_3201_0, i_10_42_3202_0, i_10_42_3270_0,
    i_10_42_3391_0, i_10_42_3408_0, i_10_42_3469_0, i_10_42_3590_0,
    i_10_42_3612_0, i_10_42_3616_0, i_10_42_3617_0, i_10_42_3645_0,
    i_10_42_3646_0, i_10_42_3647_0, i_10_42_3649_0, i_10_42_3650_0,
    i_10_42_3651_0, i_10_42_3652_0, i_10_42_3653_0, i_10_42_3726_0,
    i_10_42_3729_0, i_10_42_3783_0, i_10_42_3784_0, i_10_42_3785_0,
    i_10_42_3786_0, i_10_42_3787_0, i_10_42_3788_0, i_10_42_3811_0,
    i_10_42_3837_0, i_10_42_3843_0, i_10_42_3844_0, i_10_42_3847_0,
    i_10_42_3856_0, i_10_42_3857_0, i_10_42_3914_0, i_10_42_4012_0,
    i_10_42_4116_0, i_10_42_4117_0, i_10_42_4118_0, i_10_42_4119_0,
    i_10_42_4120_0, i_10_42_4267_0, i_10_42_4564_0, i_10_42_4565_0;
  output o_10_42_0_0;
  assign o_10_42_0_0 = 0;
endmodule



// Benchmark "kernel_10_43" written by ABC on Sun Jul 19 10:21:47 2020

module kernel_10_43 ( 
    i_10_43_27_0, i_10_43_28_0, i_10_43_48_0, i_10_43_117_0, i_10_43_118_0,
    i_10_43_121_0, i_10_43_218_0, i_10_43_315_0, i_10_43_317_0,
    i_10_43_388_0, i_10_43_390_0, i_10_43_391_0, i_10_43_445_0,
    i_10_43_463_0, i_10_43_748_0, i_10_43_892_0, i_10_43_946_0,
    i_10_43_956_0, i_10_43_958_0, i_10_43_1162_0, i_10_43_1234_0,
    i_10_43_1237_0, i_10_43_1261_0, i_10_43_1305_0, i_10_43_1309_0,
    i_10_43_1354_0, i_10_43_1362_0, i_10_43_1377_0, i_10_43_1445_0,
    i_10_43_1451_0, i_10_43_1576_0, i_10_43_1611_0, i_10_43_1613_0,
    i_10_43_1640_0, i_10_43_1732_0, i_10_43_1804_0, i_10_43_1820_0,
    i_10_43_1821_0, i_10_43_1873_0, i_10_43_1882_0, i_10_43_1899_0,
    i_10_43_1915_0, i_10_43_1917_0, i_10_43_1918_0, i_10_43_1944_0,
    i_10_43_1946_0, i_10_43_1991_0, i_10_43_2081_0, i_10_43_2155_0,
    i_10_43_2179_0, i_10_43_2180_0, i_10_43_2241_0, i_10_43_2358_0,
    i_10_43_2380_0, i_10_43_2468_0, i_10_43_2504_0, i_10_43_2629_0,
    i_10_43_2630_0, i_10_43_2631_0, i_10_43_2781_0, i_10_43_2782_0,
    i_10_43_2818_0, i_10_43_2819_0, i_10_43_2881_0, i_10_43_2882_0,
    i_10_43_3036_0, i_10_43_3038_0, i_10_43_3073_0, i_10_43_3281_0,
    i_10_43_3430_0, i_10_43_3465_0, i_10_43_3537_0, i_10_43_3582_0,
    i_10_43_3614_0, i_10_43_3645_0, i_10_43_3646_0, i_10_43_3647_0,
    i_10_43_3649_0, i_10_43_3650_0, i_10_43_3782_0, i_10_43_3784_0,
    i_10_43_3785_0, i_10_43_3842_0, i_10_43_3979_0, i_10_43_4050_0,
    i_10_43_4115_0, i_10_43_4123_0, i_10_43_4126_0, i_10_43_4217_0,
    i_10_43_4220_0, i_10_43_4261_0, i_10_43_4268_0, i_10_43_4277_0,
    i_10_43_4279_0, i_10_43_4292_0, i_10_43_4302_0, i_10_43_4527_0,
    i_10_43_4528_0, i_10_43_4529_0, i_10_43_4583_0,
    o_10_43_0_0  );
  input  i_10_43_27_0, i_10_43_28_0, i_10_43_48_0, i_10_43_117_0,
    i_10_43_118_0, i_10_43_121_0, i_10_43_218_0, i_10_43_315_0,
    i_10_43_317_0, i_10_43_388_0, i_10_43_390_0, i_10_43_391_0,
    i_10_43_445_0, i_10_43_463_0, i_10_43_748_0, i_10_43_892_0,
    i_10_43_946_0, i_10_43_956_0, i_10_43_958_0, i_10_43_1162_0,
    i_10_43_1234_0, i_10_43_1237_0, i_10_43_1261_0, i_10_43_1305_0,
    i_10_43_1309_0, i_10_43_1354_0, i_10_43_1362_0, i_10_43_1377_0,
    i_10_43_1445_0, i_10_43_1451_0, i_10_43_1576_0, i_10_43_1611_0,
    i_10_43_1613_0, i_10_43_1640_0, i_10_43_1732_0, i_10_43_1804_0,
    i_10_43_1820_0, i_10_43_1821_0, i_10_43_1873_0, i_10_43_1882_0,
    i_10_43_1899_0, i_10_43_1915_0, i_10_43_1917_0, i_10_43_1918_0,
    i_10_43_1944_0, i_10_43_1946_0, i_10_43_1991_0, i_10_43_2081_0,
    i_10_43_2155_0, i_10_43_2179_0, i_10_43_2180_0, i_10_43_2241_0,
    i_10_43_2358_0, i_10_43_2380_0, i_10_43_2468_0, i_10_43_2504_0,
    i_10_43_2629_0, i_10_43_2630_0, i_10_43_2631_0, i_10_43_2781_0,
    i_10_43_2782_0, i_10_43_2818_0, i_10_43_2819_0, i_10_43_2881_0,
    i_10_43_2882_0, i_10_43_3036_0, i_10_43_3038_0, i_10_43_3073_0,
    i_10_43_3281_0, i_10_43_3430_0, i_10_43_3465_0, i_10_43_3537_0,
    i_10_43_3582_0, i_10_43_3614_0, i_10_43_3645_0, i_10_43_3646_0,
    i_10_43_3647_0, i_10_43_3649_0, i_10_43_3650_0, i_10_43_3782_0,
    i_10_43_3784_0, i_10_43_3785_0, i_10_43_3842_0, i_10_43_3979_0,
    i_10_43_4050_0, i_10_43_4115_0, i_10_43_4123_0, i_10_43_4126_0,
    i_10_43_4217_0, i_10_43_4220_0, i_10_43_4261_0, i_10_43_4268_0,
    i_10_43_4277_0, i_10_43_4279_0, i_10_43_4292_0, i_10_43_4302_0,
    i_10_43_4527_0, i_10_43_4528_0, i_10_43_4529_0, i_10_43_4583_0;
  output o_10_43_0_0;
  assign o_10_43_0_0 = 0;
endmodule



// Benchmark "kernel_10_44" written by ABC on Sun Jul 19 10:21:47 2020

module kernel_10_44 ( 
    i_10_44_41_0, i_10_44_45_0, i_10_44_73_0, i_10_44_148_0, i_10_44_149_0,
    i_10_44_188_0, i_10_44_286_0, i_10_44_296_0, i_10_44_316_0,
    i_10_44_319_0, i_10_44_372_0, i_10_44_438_0, i_10_44_448_0,
    i_10_44_463_0, i_10_44_501_0, i_10_44_502_0, i_10_44_724_0,
    i_10_44_752_0, i_10_44_826_0, i_10_44_844_0, i_10_44_934_0,
    i_10_44_1036_0, i_10_44_1083_0, i_10_44_1085_0, i_10_44_1088_0,
    i_10_44_1166_0, i_10_44_1268_0, i_10_44_1307_0, i_10_44_1327_0,
    i_10_44_1338_0, i_10_44_1354_0, i_10_44_1534_0, i_10_44_1545_0,
    i_10_44_1555_0, i_10_44_1616_0, i_10_44_1655_0, i_10_44_1686_0,
    i_10_44_1689_0, i_10_44_1821_0, i_10_44_1872_0, i_10_44_1909_0,
    i_10_44_1910_0, i_10_44_1911_0, i_10_44_1914_0, i_10_44_1918_0,
    i_10_44_1958_0, i_10_44_1986_0, i_10_44_2093_0, i_10_44_2157_0,
    i_10_44_2166_0, i_10_44_2245_0, i_10_44_2246_0, i_10_44_2284_0,
    i_10_44_2352_0, i_10_44_2357_0, i_10_44_2380_0, i_10_44_2491_0,
    i_10_44_2560_0, i_10_44_2563_0, i_10_44_2569_0, i_10_44_2613_0,
    i_10_44_2629_0, i_10_44_2678_0, i_10_44_2697_0, i_10_44_2731_0,
    i_10_44_2734_0, i_10_44_2782_0, i_10_44_2865_0, i_10_44_2960_0,
    i_10_44_2993_0, i_10_44_3011_0, i_10_44_3012_0, i_10_44_3034_0,
    i_10_44_3036_0, i_10_44_3040_0, i_10_44_3070_0, i_10_44_3084_0,
    i_10_44_3091_0, i_10_44_3235_0, i_10_44_3264_0, i_10_44_3308_0,
    i_10_44_3317_0, i_10_44_3433_0, i_10_44_3436_0, i_10_44_3471_0,
    i_10_44_3540_0, i_10_44_3541_0, i_10_44_3617_0, i_10_44_3624_0,
    i_10_44_3641_0, i_10_44_3668_0, i_10_44_3853_0, i_10_44_3882_0,
    i_10_44_3892_0, i_10_44_4073_0, i_10_44_4157_0, i_10_44_4267_0,
    i_10_44_4534_0, i_10_44_4535_0, i_10_44_4565_0,
    o_10_44_0_0  );
  input  i_10_44_41_0, i_10_44_45_0, i_10_44_73_0, i_10_44_148_0,
    i_10_44_149_0, i_10_44_188_0, i_10_44_286_0, i_10_44_296_0,
    i_10_44_316_0, i_10_44_319_0, i_10_44_372_0, i_10_44_438_0,
    i_10_44_448_0, i_10_44_463_0, i_10_44_501_0, i_10_44_502_0,
    i_10_44_724_0, i_10_44_752_0, i_10_44_826_0, i_10_44_844_0,
    i_10_44_934_0, i_10_44_1036_0, i_10_44_1083_0, i_10_44_1085_0,
    i_10_44_1088_0, i_10_44_1166_0, i_10_44_1268_0, i_10_44_1307_0,
    i_10_44_1327_0, i_10_44_1338_0, i_10_44_1354_0, i_10_44_1534_0,
    i_10_44_1545_0, i_10_44_1555_0, i_10_44_1616_0, i_10_44_1655_0,
    i_10_44_1686_0, i_10_44_1689_0, i_10_44_1821_0, i_10_44_1872_0,
    i_10_44_1909_0, i_10_44_1910_0, i_10_44_1911_0, i_10_44_1914_0,
    i_10_44_1918_0, i_10_44_1958_0, i_10_44_1986_0, i_10_44_2093_0,
    i_10_44_2157_0, i_10_44_2166_0, i_10_44_2245_0, i_10_44_2246_0,
    i_10_44_2284_0, i_10_44_2352_0, i_10_44_2357_0, i_10_44_2380_0,
    i_10_44_2491_0, i_10_44_2560_0, i_10_44_2563_0, i_10_44_2569_0,
    i_10_44_2613_0, i_10_44_2629_0, i_10_44_2678_0, i_10_44_2697_0,
    i_10_44_2731_0, i_10_44_2734_0, i_10_44_2782_0, i_10_44_2865_0,
    i_10_44_2960_0, i_10_44_2993_0, i_10_44_3011_0, i_10_44_3012_0,
    i_10_44_3034_0, i_10_44_3036_0, i_10_44_3040_0, i_10_44_3070_0,
    i_10_44_3084_0, i_10_44_3091_0, i_10_44_3235_0, i_10_44_3264_0,
    i_10_44_3308_0, i_10_44_3317_0, i_10_44_3433_0, i_10_44_3436_0,
    i_10_44_3471_0, i_10_44_3540_0, i_10_44_3541_0, i_10_44_3617_0,
    i_10_44_3624_0, i_10_44_3641_0, i_10_44_3668_0, i_10_44_3853_0,
    i_10_44_3882_0, i_10_44_3892_0, i_10_44_4073_0, i_10_44_4157_0,
    i_10_44_4267_0, i_10_44_4534_0, i_10_44_4535_0, i_10_44_4565_0;
  output o_10_44_0_0;
  assign o_10_44_0_0 = 0;
endmodule



// Benchmark "kernel_10_45" written by ABC on Sun Jul 19 10:21:48 2020

module kernel_10_45 ( 
    i_10_45_30_0, i_10_45_33_0, i_10_45_34_0, i_10_45_121_0, i_10_45_123_0,
    i_10_45_124_0, i_10_45_132_0, i_10_45_146_0, i_10_45_157_0,
    i_10_45_183_0, i_10_45_184_0, i_10_45_185_0, i_10_45_248_0,
    i_10_45_269_0, i_10_45_317_0, i_10_45_320_0, i_10_45_431_0,
    i_10_45_444_0, i_10_45_449_0, i_10_45_462_0, i_10_45_466_0,
    i_10_45_758_0, i_10_45_921_0, i_10_45_958_0, i_10_45_1003_0,
    i_10_45_1005_0, i_10_45_1013_0, i_10_45_1015_0, i_10_45_1029_0,
    i_10_45_1048_0, i_10_45_1050_0, i_10_45_1308_0, i_10_45_1365_0,
    i_10_45_1370_0, i_10_45_1383_0, i_10_45_1500_0, i_10_45_1546_0,
    i_10_45_1579_0, i_10_45_1612_0, i_10_45_1613_0, i_10_45_1617_0,
    i_10_45_1651_0, i_10_45_1733_0, i_10_45_1767_0, i_10_45_1768_0,
    i_10_45_1906_0, i_10_45_1911_0, i_10_45_1912_0, i_10_45_1913_0,
    i_10_45_1942_0, i_10_45_1950_0, i_10_45_1951_0, i_10_45_1956_0,
    i_10_45_1957_0, i_10_45_1959_0, i_10_45_1981_0, i_10_45_2000_0,
    i_10_45_2038_0, i_10_45_2041_0, i_10_45_2094_0, i_10_45_2201_0,
    i_10_45_2562_0, i_10_45_2570_0, i_10_45_2659_0, i_10_45_2660_0,
    i_10_45_2721_0, i_10_45_2725_0, i_10_45_2787_0, i_10_45_2833_0,
    i_10_45_2834_0, i_10_45_2883_0, i_10_45_2921_0, i_10_45_2990_0,
    i_10_45_3012_0, i_10_45_3013_0, i_10_45_3202_0, i_10_45_3298_0,
    i_10_45_3299_0, i_10_45_3326_0, i_10_45_3392_0, i_10_45_3473_0,
    i_10_45_3558_0, i_10_45_3589_0, i_10_45_3617_0, i_10_45_3624_0,
    i_10_45_3840_0, i_10_45_3841_0, i_10_45_3855_0, i_10_45_3858_0,
    i_10_45_3945_0, i_10_45_3980_0, i_10_45_3995_0, i_10_45_4053_0,
    i_10_45_4116_0, i_10_45_4183_0, i_10_45_4288_0, i_10_45_4299_0,
    i_10_45_4547_0, i_10_45_4569_0, i_10_45_4593_0,
    o_10_45_0_0  );
  input  i_10_45_30_0, i_10_45_33_0, i_10_45_34_0, i_10_45_121_0,
    i_10_45_123_0, i_10_45_124_0, i_10_45_132_0, i_10_45_146_0,
    i_10_45_157_0, i_10_45_183_0, i_10_45_184_0, i_10_45_185_0,
    i_10_45_248_0, i_10_45_269_0, i_10_45_317_0, i_10_45_320_0,
    i_10_45_431_0, i_10_45_444_0, i_10_45_449_0, i_10_45_462_0,
    i_10_45_466_0, i_10_45_758_0, i_10_45_921_0, i_10_45_958_0,
    i_10_45_1003_0, i_10_45_1005_0, i_10_45_1013_0, i_10_45_1015_0,
    i_10_45_1029_0, i_10_45_1048_0, i_10_45_1050_0, i_10_45_1308_0,
    i_10_45_1365_0, i_10_45_1370_0, i_10_45_1383_0, i_10_45_1500_0,
    i_10_45_1546_0, i_10_45_1579_0, i_10_45_1612_0, i_10_45_1613_0,
    i_10_45_1617_0, i_10_45_1651_0, i_10_45_1733_0, i_10_45_1767_0,
    i_10_45_1768_0, i_10_45_1906_0, i_10_45_1911_0, i_10_45_1912_0,
    i_10_45_1913_0, i_10_45_1942_0, i_10_45_1950_0, i_10_45_1951_0,
    i_10_45_1956_0, i_10_45_1957_0, i_10_45_1959_0, i_10_45_1981_0,
    i_10_45_2000_0, i_10_45_2038_0, i_10_45_2041_0, i_10_45_2094_0,
    i_10_45_2201_0, i_10_45_2562_0, i_10_45_2570_0, i_10_45_2659_0,
    i_10_45_2660_0, i_10_45_2721_0, i_10_45_2725_0, i_10_45_2787_0,
    i_10_45_2833_0, i_10_45_2834_0, i_10_45_2883_0, i_10_45_2921_0,
    i_10_45_2990_0, i_10_45_3012_0, i_10_45_3013_0, i_10_45_3202_0,
    i_10_45_3298_0, i_10_45_3299_0, i_10_45_3326_0, i_10_45_3392_0,
    i_10_45_3473_0, i_10_45_3558_0, i_10_45_3589_0, i_10_45_3617_0,
    i_10_45_3624_0, i_10_45_3840_0, i_10_45_3841_0, i_10_45_3855_0,
    i_10_45_3858_0, i_10_45_3945_0, i_10_45_3980_0, i_10_45_3995_0,
    i_10_45_4053_0, i_10_45_4116_0, i_10_45_4183_0, i_10_45_4288_0,
    i_10_45_4299_0, i_10_45_4547_0, i_10_45_4569_0, i_10_45_4593_0;
  output o_10_45_0_0;
  assign o_10_45_0_0 = 0;
endmodule



// Benchmark "kernel_10_46" written by ABC on Sun Jul 19 10:21:49 2020

module kernel_10_46 ( 
    i_10_46_38_0, i_10_46_149_0, i_10_46_155_0, i_10_46_171_0,
    i_10_46_172_0, i_10_46_178_0, i_10_46_218_0, i_10_46_244_0,
    i_10_46_245_0, i_10_46_248_0, i_10_46_280_0, i_10_46_286_0,
    i_10_46_287_0, i_10_46_317_0, i_10_46_328_0, i_10_46_329_0,
    i_10_46_332_0, i_10_46_440_0, i_10_46_443_0, i_10_46_465_0,
    i_10_46_749_0, i_10_46_796_0, i_10_46_797_0, i_10_46_901_0,
    i_10_46_991_0, i_10_46_1028_0, i_10_46_1234_0, i_10_46_1244_0,
    i_10_46_1247_0, i_10_46_1265_0, i_10_46_1307_0, i_10_46_1309_0,
    i_10_46_1577_0, i_10_46_1579_0, i_10_46_1580_0, i_10_46_1595_0,
    i_10_46_1648_0, i_10_46_1649_0, i_10_46_1652_0, i_10_46_1690_0,
    i_10_46_1691_0, i_10_46_1811_0, i_10_46_1819_0, i_10_46_1824_0,
    i_10_46_1946_0, i_10_46_2018_0, i_10_46_2024_0, i_10_46_2197_0,
    i_10_46_2201_0, i_10_46_2312_0, i_10_46_2350_0, i_10_46_2351_0,
    i_10_46_2353_0, i_10_46_2354_0, i_10_46_2406_0, i_10_46_2467_0,
    i_10_46_2470_0, i_10_46_2503_0, i_10_46_2602_0, i_10_46_2603_0,
    i_10_46_2606_0, i_10_46_2634_0, i_10_46_2660_0, i_10_46_2710_0,
    i_10_46_2711_0, i_10_46_2729_0, i_10_46_2731_0, i_10_46_2827_0,
    i_10_46_2830_0, i_10_46_2831_0, i_10_46_2834_0, i_10_46_3161_0,
    i_10_46_3196_0, i_10_46_3197_0, i_10_46_3278_0, i_10_46_3583_0,
    i_10_46_3585_0, i_10_46_3586_0, i_10_46_3613_0, i_10_46_3650_0,
    i_10_46_3686_0, i_10_46_3781_0, i_10_46_3786_0, i_10_46_3809_0,
    i_10_46_3835_0, i_10_46_3841_0, i_10_46_3848_0, i_10_46_3889_0,
    i_10_46_3908_0, i_10_46_4114_0, i_10_46_4115_0, i_10_46_4172_0,
    i_10_46_4277_0, i_10_46_4285_0, i_10_46_4286_0, i_10_46_4288_0,
    i_10_46_4289_0, i_10_46_4291_0, i_10_46_4565_0, i_10_46_4570_0,
    o_10_46_0_0  );
  input  i_10_46_38_0, i_10_46_149_0, i_10_46_155_0, i_10_46_171_0,
    i_10_46_172_0, i_10_46_178_0, i_10_46_218_0, i_10_46_244_0,
    i_10_46_245_0, i_10_46_248_0, i_10_46_280_0, i_10_46_286_0,
    i_10_46_287_0, i_10_46_317_0, i_10_46_328_0, i_10_46_329_0,
    i_10_46_332_0, i_10_46_440_0, i_10_46_443_0, i_10_46_465_0,
    i_10_46_749_0, i_10_46_796_0, i_10_46_797_0, i_10_46_901_0,
    i_10_46_991_0, i_10_46_1028_0, i_10_46_1234_0, i_10_46_1244_0,
    i_10_46_1247_0, i_10_46_1265_0, i_10_46_1307_0, i_10_46_1309_0,
    i_10_46_1577_0, i_10_46_1579_0, i_10_46_1580_0, i_10_46_1595_0,
    i_10_46_1648_0, i_10_46_1649_0, i_10_46_1652_0, i_10_46_1690_0,
    i_10_46_1691_0, i_10_46_1811_0, i_10_46_1819_0, i_10_46_1824_0,
    i_10_46_1946_0, i_10_46_2018_0, i_10_46_2024_0, i_10_46_2197_0,
    i_10_46_2201_0, i_10_46_2312_0, i_10_46_2350_0, i_10_46_2351_0,
    i_10_46_2353_0, i_10_46_2354_0, i_10_46_2406_0, i_10_46_2467_0,
    i_10_46_2470_0, i_10_46_2503_0, i_10_46_2602_0, i_10_46_2603_0,
    i_10_46_2606_0, i_10_46_2634_0, i_10_46_2660_0, i_10_46_2710_0,
    i_10_46_2711_0, i_10_46_2729_0, i_10_46_2731_0, i_10_46_2827_0,
    i_10_46_2830_0, i_10_46_2831_0, i_10_46_2834_0, i_10_46_3161_0,
    i_10_46_3196_0, i_10_46_3197_0, i_10_46_3278_0, i_10_46_3583_0,
    i_10_46_3585_0, i_10_46_3586_0, i_10_46_3613_0, i_10_46_3650_0,
    i_10_46_3686_0, i_10_46_3781_0, i_10_46_3786_0, i_10_46_3809_0,
    i_10_46_3835_0, i_10_46_3841_0, i_10_46_3848_0, i_10_46_3889_0,
    i_10_46_3908_0, i_10_46_4114_0, i_10_46_4115_0, i_10_46_4172_0,
    i_10_46_4277_0, i_10_46_4285_0, i_10_46_4286_0, i_10_46_4288_0,
    i_10_46_4289_0, i_10_46_4291_0, i_10_46_4565_0, i_10_46_4570_0;
  output o_10_46_0_0;
  assign o_10_46_0_0 = ~((~i_10_46_2603_0 & ((~i_10_46_245_0 & ((~i_10_46_1265_0 & ~i_10_46_1580_0 & ~i_10_46_1691_0 & ~i_10_46_1811_0) | (~i_10_46_287_0 & ~i_10_46_901_0 & ~i_10_46_1649_0 & ~i_10_46_1824_0 & ~i_10_46_2312_0 & i_10_46_2351_0))) | (~i_10_46_248_0 & ((~i_10_46_749_0 & i_10_46_2634_0) | (~i_10_46_901_0 & ~i_10_46_1307_0 & ~i_10_46_1652_0 & ~i_10_46_4286_0))) | (~i_10_46_2606_0 & ((~i_10_46_329_0 & ((~i_10_46_244_0 & ~i_10_46_1824_0 & ~i_10_46_4114_0) | (~i_10_46_1648_0 & ~i_10_46_2024_0 & ~i_10_46_2503_0 & ~i_10_46_2602_0 & ~i_10_46_3781_0 & ~i_10_46_4277_0))) | (~i_10_46_1028_0 & ~i_10_46_1811_0 & ~i_10_46_3686_0 & ~i_10_46_4115_0))) | (~i_10_46_2602_0 & ((~i_10_46_2351_0 & ((i_10_46_280_0 & ~i_10_46_443_0 & ~i_10_46_3586_0 & ~i_10_46_3650_0) | (~i_10_46_749_0 & ~i_10_46_797_0 & ~i_10_46_1247_0 & ~i_10_46_3278_0 & ~i_10_46_3781_0 & ~i_10_46_3786_0 & ~i_10_46_4277_0))) | (~i_10_46_328_0 & ~i_10_46_1244_0 & ~i_10_46_1690_0 & ~i_10_46_2201_0 & ~i_10_46_2660_0 & ~i_10_46_2710_0 & ~i_10_46_4277_0))) | (i_10_46_244_0 & ~i_10_46_1577_0 & ~i_10_46_2197_0 & ~i_10_46_2350_0 & ~i_10_46_2354_0 & ~i_10_46_3686_0 & ~i_10_46_3841_0))) | (~i_10_46_1579_0 & ((~i_10_46_245_0 & ~i_10_46_328_0 & ~i_10_46_1811_0 & ~i_10_46_2312_0 & ~i_10_46_2602_0 & ~i_10_46_3161_0 & ~i_10_46_3841_0) | (~i_10_46_178_0 & ~i_10_46_280_0 & ~i_10_46_2350_0 & ~i_10_46_3650_0 & ~i_10_46_4565_0))) | (~i_10_46_245_0 & ((~i_10_46_443_0 & i_10_46_1579_0 & ~i_10_46_2312_0 & ~i_10_46_2827_0 & i_10_46_2831_0) | (~i_10_46_440_0 & ~i_10_46_796_0 & ~i_10_46_1247_0 & i_10_46_1580_0 & ~i_10_46_2503_0 & ~i_10_46_3613_0 & i_10_46_3650_0 & ~i_10_46_3908_0))) | (~i_10_46_2602_0 & ((~i_10_46_1649_0 & ~i_10_46_2312_0 & ~i_10_46_2831_0 & i_10_46_3583_0 & ~i_10_46_3686_0) | (~i_10_46_149_0 & ~i_10_46_1244_0 & i_10_46_1819_0 & ~i_10_46_2731_0 & i_10_46_3781_0 & i_10_46_4114_0))) | (i_10_46_286_0 & ~i_10_46_2606_0 & i_10_46_3686_0) | (~i_10_46_1309_0 & ~i_10_46_1652_0 & i_10_46_1824_0 & ~i_10_46_2729_0 & ~i_10_46_3841_0) | (i_10_46_149_0 & i_10_46_2731_0 & ~i_10_46_4115_0));
endmodule



// Benchmark "kernel_10_47" written by ABC on Sun Jul 19 10:21:51 2020

module kernel_10_47 ( 
    i_10_47_174_0, i_10_47_175_0, i_10_47_177_0, i_10_47_244_0,
    i_10_47_245_0, i_10_47_247_0, i_10_47_276_0, i_10_47_289_0,
    i_10_47_290_0, i_10_47_292_0, i_10_47_293_0, i_10_47_361_0,
    i_10_47_364_0, i_10_47_405_0, i_10_47_406_0, i_10_47_409_0,
    i_10_47_410_0, i_10_47_411_0, i_10_47_412_0, i_10_47_435_0,
    i_10_47_445_0, i_10_47_456_0, i_10_47_460_0, i_10_47_461_0,
    i_10_47_463_0, i_10_47_467_0, i_10_47_510_0, i_10_47_749_0,
    i_10_47_792_0, i_10_47_796_0, i_10_47_797_0, i_10_47_799_0,
    i_10_47_800_0, i_10_47_1269_0, i_10_47_1306_0, i_10_47_1359_0,
    i_10_47_1441_0, i_10_47_1442_0, i_10_47_1649_0, i_10_47_1655_0,
    i_10_47_1819_0, i_10_47_1822_0, i_10_47_1910_0, i_10_47_1992_0,
    i_10_47_2178_0, i_10_47_2359_0, i_10_47_2360_0, i_10_47_2361_0,
    i_10_47_2448_0, i_10_47_2467_0, i_10_47_2468_0, i_10_47_2628_0,
    i_10_47_2630_0, i_10_47_2631_0, i_10_47_2632_0, i_10_47_2658_0,
    i_10_47_2659_0, i_10_47_2661_0, i_10_47_2673_0, i_10_47_2680_0,
    i_10_47_2702_0, i_10_47_2731_0, i_10_47_2781_0, i_10_47_2783_0,
    i_10_47_2784_0, i_10_47_2882_0, i_10_47_2980_0, i_10_47_3044_0,
    i_10_47_3069_0, i_10_47_3070_0, i_10_47_3071_0, i_10_47_3073_0,
    i_10_47_3074_0, i_10_47_3277_0, i_10_47_3278_0, i_10_47_3321_0,
    i_10_47_3323_0, i_10_47_3328_0, i_10_47_3384_0, i_10_47_3392_0,
    i_10_47_3523_0, i_10_47_3610_0, i_10_47_3613_0, i_10_47_3787_0,
    i_10_47_3788_0, i_10_47_3807_0, i_10_47_3808_0, i_10_47_3849_0,
    i_10_47_3855_0, i_10_47_3858_0, i_10_47_3983_0, i_10_47_3994_0,
    i_10_47_4119_0, i_10_47_4270_0, i_10_47_4285_0, i_10_47_4288_0,
    i_10_47_4289_0, i_10_47_4291_0, i_10_47_4292_0, i_10_47_4564_0,
    o_10_47_0_0  );
  input  i_10_47_174_0, i_10_47_175_0, i_10_47_177_0, i_10_47_244_0,
    i_10_47_245_0, i_10_47_247_0, i_10_47_276_0, i_10_47_289_0,
    i_10_47_290_0, i_10_47_292_0, i_10_47_293_0, i_10_47_361_0,
    i_10_47_364_0, i_10_47_405_0, i_10_47_406_0, i_10_47_409_0,
    i_10_47_410_0, i_10_47_411_0, i_10_47_412_0, i_10_47_435_0,
    i_10_47_445_0, i_10_47_456_0, i_10_47_460_0, i_10_47_461_0,
    i_10_47_463_0, i_10_47_467_0, i_10_47_510_0, i_10_47_749_0,
    i_10_47_792_0, i_10_47_796_0, i_10_47_797_0, i_10_47_799_0,
    i_10_47_800_0, i_10_47_1269_0, i_10_47_1306_0, i_10_47_1359_0,
    i_10_47_1441_0, i_10_47_1442_0, i_10_47_1649_0, i_10_47_1655_0,
    i_10_47_1819_0, i_10_47_1822_0, i_10_47_1910_0, i_10_47_1992_0,
    i_10_47_2178_0, i_10_47_2359_0, i_10_47_2360_0, i_10_47_2361_0,
    i_10_47_2448_0, i_10_47_2467_0, i_10_47_2468_0, i_10_47_2628_0,
    i_10_47_2630_0, i_10_47_2631_0, i_10_47_2632_0, i_10_47_2658_0,
    i_10_47_2659_0, i_10_47_2661_0, i_10_47_2673_0, i_10_47_2680_0,
    i_10_47_2702_0, i_10_47_2731_0, i_10_47_2781_0, i_10_47_2783_0,
    i_10_47_2784_0, i_10_47_2882_0, i_10_47_2980_0, i_10_47_3044_0,
    i_10_47_3069_0, i_10_47_3070_0, i_10_47_3071_0, i_10_47_3073_0,
    i_10_47_3074_0, i_10_47_3277_0, i_10_47_3278_0, i_10_47_3321_0,
    i_10_47_3323_0, i_10_47_3328_0, i_10_47_3384_0, i_10_47_3392_0,
    i_10_47_3523_0, i_10_47_3610_0, i_10_47_3613_0, i_10_47_3787_0,
    i_10_47_3788_0, i_10_47_3807_0, i_10_47_3808_0, i_10_47_3849_0,
    i_10_47_3855_0, i_10_47_3858_0, i_10_47_3983_0, i_10_47_3994_0,
    i_10_47_4119_0, i_10_47_4270_0, i_10_47_4285_0, i_10_47_4288_0,
    i_10_47_4289_0, i_10_47_4291_0, i_10_47_4292_0, i_10_47_4564_0;
  output o_10_47_0_0;
  assign o_10_47_0_0 = ~((~i_10_47_177_0 & ~i_10_47_3073_0 & ((~i_10_47_799_0 & ~i_10_47_1359_0 & ~i_10_47_1655_0 & ~i_10_47_2361_0 & ~i_10_47_2448_0 & ~i_10_47_2702_0 & ~i_10_47_3384_0) | (~i_10_47_174_0 & ~i_10_47_175_0 & ~i_10_47_244_0 & ~i_10_47_293_0 & ~i_10_47_3855_0))) | (~i_10_47_175_0 & ((~i_10_47_405_0 & ~i_10_47_412_0 & i_10_47_1819_0 & ~i_10_47_2468_0 & ~i_10_47_3613_0) | (~i_10_47_411_0 & ~i_10_47_796_0 & ~i_10_47_2783_0 & ~i_10_47_3071_0 & ~i_10_47_3074_0 & i_10_47_4119_0))) | (i_10_47_244_0 & ((~i_10_47_289_0 & ~i_10_47_290_0 & ~i_10_47_799_0 & i_10_47_1306_0 & ~i_10_47_2361_0 & ~i_10_47_3787_0) | (~i_10_47_463_0 & ~i_10_47_1306_0 & ~i_10_47_1819_0 & ~i_10_47_3070_0 & ~i_10_47_3613_0 & ~i_10_47_4564_0))) | (~i_10_47_247_0 & ((~i_10_47_245_0 & ~i_10_47_289_0 & ~i_10_47_410_0 & ~i_10_47_800_0 & ~i_10_47_2784_0 & ~i_10_47_3994_0) | (~i_10_47_409_0 & ~i_10_47_1306_0 & ~i_10_47_1992_0 & i_10_47_3788_0 & ~i_10_47_4119_0))) | (~i_10_47_3074_0 & ((~i_10_47_292_0 & ~i_10_47_409_0 & ((~i_10_47_411_0 & ~i_10_47_2361_0 & ~i_10_47_3071_0) | (~i_10_47_406_0 & ~i_10_47_456_0 & ~i_10_47_3787_0))) | (~i_10_47_3044_0 & ((~i_10_47_289_0 & ~i_10_47_412_0 & ~i_10_47_463_0 & ~i_10_47_2784_0 & ~i_10_47_3994_0 & ~i_10_47_2361_0 & ~i_10_47_2783_0) | (~i_10_47_290_0 & ~i_10_47_411_0 & ~i_10_47_2680_0 & ~i_10_47_3070_0 & ~i_10_47_3071_0 & ~i_10_47_3392_0 & ~i_10_47_4119_0 & ~i_10_47_4564_0))) | (~i_10_47_456_0 & i_10_47_463_0 & i_10_47_3858_0))) | (~i_10_47_293_0 & ~i_10_47_1442_0 & ((~i_10_47_244_0 & ~i_10_47_406_0 & ~i_10_47_409_0 & ~i_10_47_799_0 & ~i_10_47_2781_0 & ~i_10_47_3613_0) | (~i_10_47_1441_0 & i_10_47_1819_0 & ~i_10_47_2361_0 & ~i_10_47_3788_0))) | (~i_10_47_797_0 & ((~i_10_47_2361_0 & i_10_47_4270_0) | (~i_10_47_2630_0 & ~i_10_47_2702_0 & ~i_10_47_2784_0 & ~i_10_47_3071_0 & i_10_47_3613_0 & ~i_10_47_3787_0 & ~i_10_47_4564_0))) | (~i_10_47_800_0 & ((~i_10_47_2784_0 & ~i_10_47_3070_0 & ~i_10_47_3384_0 & ~i_10_47_3523_0 & ~i_10_47_3787_0) | (~i_10_47_409_0 & i_10_47_2659_0 & ~i_10_47_4119_0))) | (i_10_47_445_0 & ((i_10_47_2731_0 & (i_10_47_456_0 | i_10_47_2661_0)) | (i_10_47_463_0 & ~i_10_47_796_0 & ~i_10_47_4119_0))) | (~i_10_47_463_0 & i_10_47_1649_0 & i_10_47_2632_0 & i_10_47_3855_0 & i_10_47_3858_0));
endmodule



// Benchmark "kernel_10_48" written by ABC on Sun Jul 19 10:21:52 2020

module kernel_10_48 ( 
    i_10_48_174_0, i_10_48_180_0, i_10_48_248_0, i_10_48_287_0,
    i_10_48_327_0, i_10_48_369_0, i_10_48_448_0, i_10_48_586_0,
    i_10_48_588_0, i_10_48_633_0, i_10_48_781_0, i_10_48_782_0,
    i_10_48_795_0, i_10_48_798_0, i_10_48_799_0, i_10_48_904_0,
    i_10_48_1087_0, i_10_48_1235_0, i_10_48_1241_0, i_10_48_1249_0,
    i_10_48_1362_0, i_10_48_1363_0, i_10_48_1450_0, i_10_48_1453_0,
    i_10_48_1454_0, i_10_48_1490_0, i_10_48_1551_0, i_10_48_1555_0,
    i_10_48_1577_0, i_10_48_1646_0, i_10_48_1789_0, i_10_48_1882_0,
    i_10_48_1911_0, i_10_48_1914_0, i_10_48_1979_0, i_10_48_2028_0,
    i_10_48_2082_0, i_10_48_2085_0, i_10_48_2155_0, i_10_48_2158_0,
    i_10_48_2159_0, i_10_48_2241_0, i_10_48_2261_0, i_10_48_2264_0,
    i_10_48_2310_0, i_10_48_2322_0, i_10_48_2337_0, i_10_48_2353_0,
    i_10_48_2383_0, i_10_48_2385_0, i_10_48_2407_0, i_10_48_2411_0,
    i_10_48_2442_0, i_10_48_2443_0, i_10_48_2449_0, i_10_48_2451_0,
    i_10_48_2452_0, i_10_48_2517_0, i_10_48_2518_0, i_10_48_2539_0,
    i_10_48_2572_0, i_10_48_2573_0, i_10_48_2648_0, i_10_48_2703_0,
    i_10_48_2707_0, i_10_48_2921_0, i_10_48_2924_0, i_10_48_2954_0,
    i_10_48_2957_0, i_10_48_3101_0, i_10_48_3228_0, i_10_48_3360_0,
    i_10_48_3390_0, i_10_48_3492_0, i_10_48_3499_0, i_10_48_3525_0,
    i_10_48_3577_0, i_10_48_3613_0, i_10_48_3618_0, i_10_48_3649_0,
    i_10_48_3784_0, i_10_48_3837_0, i_10_48_3838_0, i_10_48_3850_0,
    i_10_48_3856_0, i_10_48_3895_0, i_10_48_3963_0, i_10_48_3964_0,
    i_10_48_3983_0, i_10_48_4120_0, i_10_48_4188_0, i_10_48_4273_0,
    i_10_48_4289_0, i_10_48_4423_0, i_10_48_4458_0, i_10_48_4461_0,
    i_10_48_4513_0, i_10_48_4525_0, i_10_48_4566_0, i_10_48_4569_0,
    o_10_48_0_0  );
  input  i_10_48_174_0, i_10_48_180_0, i_10_48_248_0, i_10_48_287_0,
    i_10_48_327_0, i_10_48_369_0, i_10_48_448_0, i_10_48_586_0,
    i_10_48_588_0, i_10_48_633_0, i_10_48_781_0, i_10_48_782_0,
    i_10_48_795_0, i_10_48_798_0, i_10_48_799_0, i_10_48_904_0,
    i_10_48_1087_0, i_10_48_1235_0, i_10_48_1241_0, i_10_48_1249_0,
    i_10_48_1362_0, i_10_48_1363_0, i_10_48_1450_0, i_10_48_1453_0,
    i_10_48_1454_0, i_10_48_1490_0, i_10_48_1551_0, i_10_48_1555_0,
    i_10_48_1577_0, i_10_48_1646_0, i_10_48_1789_0, i_10_48_1882_0,
    i_10_48_1911_0, i_10_48_1914_0, i_10_48_1979_0, i_10_48_2028_0,
    i_10_48_2082_0, i_10_48_2085_0, i_10_48_2155_0, i_10_48_2158_0,
    i_10_48_2159_0, i_10_48_2241_0, i_10_48_2261_0, i_10_48_2264_0,
    i_10_48_2310_0, i_10_48_2322_0, i_10_48_2337_0, i_10_48_2353_0,
    i_10_48_2383_0, i_10_48_2385_0, i_10_48_2407_0, i_10_48_2411_0,
    i_10_48_2442_0, i_10_48_2443_0, i_10_48_2449_0, i_10_48_2451_0,
    i_10_48_2452_0, i_10_48_2517_0, i_10_48_2518_0, i_10_48_2539_0,
    i_10_48_2572_0, i_10_48_2573_0, i_10_48_2648_0, i_10_48_2703_0,
    i_10_48_2707_0, i_10_48_2921_0, i_10_48_2924_0, i_10_48_2954_0,
    i_10_48_2957_0, i_10_48_3101_0, i_10_48_3228_0, i_10_48_3360_0,
    i_10_48_3390_0, i_10_48_3492_0, i_10_48_3499_0, i_10_48_3525_0,
    i_10_48_3577_0, i_10_48_3613_0, i_10_48_3618_0, i_10_48_3649_0,
    i_10_48_3784_0, i_10_48_3837_0, i_10_48_3838_0, i_10_48_3850_0,
    i_10_48_3856_0, i_10_48_3895_0, i_10_48_3963_0, i_10_48_3964_0,
    i_10_48_3983_0, i_10_48_4120_0, i_10_48_4188_0, i_10_48_4273_0,
    i_10_48_4289_0, i_10_48_4423_0, i_10_48_4458_0, i_10_48_4461_0,
    i_10_48_4513_0, i_10_48_4525_0, i_10_48_4566_0, i_10_48_4569_0;
  output o_10_48_0_0;
  assign o_10_48_0_0 = 0;
endmodule



// Benchmark "kernel_10_49" written by ABC on Sun Jul 19 10:21:53 2020

module kernel_10_49 ( 
    i_10_49_30_0, i_10_49_117_0, i_10_49_171_0, i_10_49_172_0,
    i_10_49_173_0, i_10_49_174_0, i_10_49_175_0, i_10_49_285_0,
    i_10_49_315_0, i_10_49_318_0, i_10_49_325_0, i_10_49_424_0,
    i_10_49_427_0, i_10_49_432_0, i_10_49_448_0, i_10_49_796_0,
    i_10_49_797_0, i_10_49_800_0, i_10_49_955_0, i_10_49_957_0,
    i_10_49_958_0, i_10_49_959_0, i_10_49_968_0, i_10_49_1002_0,
    i_10_49_1028_0, i_10_49_1029_0, i_10_49_1308_0, i_10_49_1311_0,
    i_10_49_1361_0, i_10_49_1614_0, i_10_49_1617_0, i_10_49_1652_0,
    i_10_49_1821_0, i_10_49_1944_0, i_10_49_1945_0, i_10_49_1956_0,
    i_10_49_2016_0, i_10_49_2178_0, i_10_49_2179_0, i_10_49_2181_0,
    i_10_49_2184_0, i_10_49_2308_0, i_10_49_2354_0, i_10_49_2358_0,
    i_10_49_2359_0, i_10_49_2361_0, i_10_49_2362_0, i_10_49_2448_0,
    i_10_49_2457_0, i_10_49_2613_0, i_10_49_2628_0, i_10_49_2629_0,
    i_10_49_2631_0, i_10_49_2635_0, i_10_49_2700_0, i_10_49_2701_0,
    i_10_49_2702_0, i_10_49_2718_0, i_10_49_2782_0, i_10_49_2823_0,
    i_10_49_2826_0, i_10_49_2885_0, i_10_49_3033_0, i_10_49_3034_0,
    i_10_49_3036_0, i_10_49_3037_0, i_10_49_3041_0, i_10_49_3045_0,
    i_10_49_3046_0, i_10_49_3087_0, i_10_49_3151_0, i_10_49_3195_0,
    i_10_49_3196_0, i_10_49_3197_0, i_10_49_3271_0, i_10_49_3278_0,
    i_10_49_3403_0, i_10_49_3616_0, i_10_49_3645_0, i_10_49_3648_0,
    i_10_49_3649_0, i_10_49_3650_0, i_10_49_3651_0, i_10_49_3652_0,
    i_10_49_3780_0, i_10_49_3786_0, i_10_49_3838_0, i_10_49_3852_0,
    i_10_49_3853_0, i_10_49_3855_0, i_10_49_3856_0, i_10_49_3858_0,
    i_10_49_4050_0, i_10_49_4122_0, i_10_49_4123_0, i_10_49_4266_0,
    i_10_49_4288_0, i_10_49_4458_0, i_10_49_4459_0, i_10_49_4571_0,
    o_10_49_0_0  );
  input  i_10_49_30_0, i_10_49_117_0, i_10_49_171_0, i_10_49_172_0,
    i_10_49_173_0, i_10_49_174_0, i_10_49_175_0, i_10_49_285_0,
    i_10_49_315_0, i_10_49_318_0, i_10_49_325_0, i_10_49_424_0,
    i_10_49_427_0, i_10_49_432_0, i_10_49_448_0, i_10_49_796_0,
    i_10_49_797_0, i_10_49_800_0, i_10_49_955_0, i_10_49_957_0,
    i_10_49_958_0, i_10_49_959_0, i_10_49_968_0, i_10_49_1002_0,
    i_10_49_1028_0, i_10_49_1029_0, i_10_49_1308_0, i_10_49_1311_0,
    i_10_49_1361_0, i_10_49_1614_0, i_10_49_1617_0, i_10_49_1652_0,
    i_10_49_1821_0, i_10_49_1944_0, i_10_49_1945_0, i_10_49_1956_0,
    i_10_49_2016_0, i_10_49_2178_0, i_10_49_2179_0, i_10_49_2181_0,
    i_10_49_2184_0, i_10_49_2308_0, i_10_49_2354_0, i_10_49_2358_0,
    i_10_49_2359_0, i_10_49_2361_0, i_10_49_2362_0, i_10_49_2448_0,
    i_10_49_2457_0, i_10_49_2613_0, i_10_49_2628_0, i_10_49_2629_0,
    i_10_49_2631_0, i_10_49_2635_0, i_10_49_2700_0, i_10_49_2701_0,
    i_10_49_2702_0, i_10_49_2718_0, i_10_49_2782_0, i_10_49_2823_0,
    i_10_49_2826_0, i_10_49_2885_0, i_10_49_3033_0, i_10_49_3034_0,
    i_10_49_3036_0, i_10_49_3037_0, i_10_49_3041_0, i_10_49_3045_0,
    i_10_49_3046_0, i_10_49_3087_0, i_10_49_3151_0, i_10_49_3195_0,
    i_10_49_3196_0, i_10_49_3197_0, i_10_49_3271_0, i_10_49_3278_0,
    i_10_49_3403_0, i_10_49_3616_0, i_10_49_3645_0, i_10_49_3648_0,
    i_10_49_3649_0, i_10_49_3650_0, i_10_49_3651_0, i_10_49_3652_0,
    i_10_49_3780_0, i_10_49_3786_0, i_10_49_3838_0, i_10_49_3852_0,
    i_10_49_3853_0, i_10_49_3855_0, i_10_49_3856_0, i_10_49_3858_0,
    i_10_49_4050_0, i_10_49_4122_0, i_10_49_4123_0, i_10_49_4266_0,
    i_10_49_4288_0, i_10_49_4458_0, i_10_49_4459_0, i_10_49_4571_0;
  output o_10_49_0_0;
  assign o_10_49_0_0 = ~((~i_10_49_117_0 & ~i_10_49_3271_0 & ((~i_10_49_1614_0 & ~i_10_49_2178_0 & ~i_10_49_2181_0 & ~i_10_49_2361_0 & ~i_10_49_3045_0 & ~i_10_49_3046_0 & ~i_10_49_3858_0) | (~i_10_49_955_0 & ~i_10_49_958_0 & ~i_10_49_1002_0 & ~i_10_49_1311_0 & ~i_10_49_2457_0 & ~i_10_49_4288_0))) | (~i_10_49_424_0 & ((~i_10_49_957_0 & ~i_10_49_1311_0 & ~i_10_49_2178_0 & ~i_10_49_2179_0 & ~i_10_49_3403_0 & ~i_10_49_3652_0) | (~i_10_49_2826_0 & ~i_10_49_3036_0 & ~i_10_49_3780_0 & ~i_10_49_3853_0))) | (~i_10_49_957_0 & ((~i_10_49_174_0 & i_10_49_1821_0 & ~i_10_49_2362_0 & ~i_10_49_2826_0 & ~i_10_49_3033_0 & i_10_49_3853_0) | (~i_10_49_30_0 & ~i_10_49_1617_0 & ~i_10_49_1945_0 & ~i_10_49_2179_0 & ~i_10_49_2358_0 & ~i_10_49_3852_0 & ~i_10_49_4050_0))) | (~i_10_49_959_0 & ((i_10_49_172_0 & ~i_10_49_2629_0) | (~i_10_49_1029_0 & ~i_10_49_2178_0 & ~i_10_49_3195_0 & ~i_10_49_3780_0 & ~i_10_49_3855_0 & ~i_10_49_4050_0 & ~i_10_49_4122_0))) | (~i_10_49_1029_0 & ((~i_10_49_30_0 & i_10_49_1821_0 & ~i_10_49_2629_0 & i_10_49_2631_0 & ~i_10_49_2823_0) | (~i_10_49_2362_0 & ~i_10_49_2613_0 & ~i_10_49_2718_0 & ~i_10_49_3650_0 & ~i_10_49_3780_0 & ~i_10_49_4050_0 & ~i_10_49_4288_0))) | (~i_10_49_30_0 & ~i_10_49_1944_0 & ((~i_10_49_1028_0 & ~i_10_49_1945_0 & ~i_10_49_2181_0 & ~i_10_49_2184_0 & ~i_10_49_2359_0 & ~i_10_49_2362_0 & ~i_10_49_2718_0 & ~i_10_49_2826_0 & ~i_10_49_3197_0) | (~i_10_49_427_0 & ~i_10_49_3036_0 & ~i_10_49_3195_0 & ~i_10_49_3196_0 & ~i_10_49_3403_0 & ~i_10_49_3780_0 & ~i_10_49_4288_0))) | (~i_10_49_1028_0 & ~i_10_49_1614_0 & ((~i_10_49_432_0 & ~i_10_49_2613_0 & ~i_10_49_3046_0 & ~i_10_49_3648_0 & ~i_10_49_3650_0 & ~i_10_49_3652_0) | (~i_10_49_1821_0 & ~i_10_49_2628_0 & ~i_10_49_3034_0 & ~i_10_49_3786_0))) | (~i_10_49_3034_0 & ((i_10_49_3041_0 & ~i_10_49_3855_0) | (~i_10_49_2613_0 & ~i_10_49_3045_0 & ~i_10_49_3786_0 & i_10_49_3858_0))) | (~i_10_49_1311_0 & i_10_49_1652_0 & ~i_10_49_2179_0 & ~i_10_49_3786_0) | (i_10_49_173_0 & ~i_10_49_2457_0) | (i_10_49_1308_0 & i_10_49_3041_0 & ~i_10_49_3648_0 & i_10_49_3651_0) | (~i_10_49_3037_0 & i_10_49_3197_0 & i_10_49_3652_0 & i_10_49_3838_0 & i_10_49_3855_0) | (~i_10_49_2631_0 & ~i_10_49_3033_0 & ~i_10_49_3856_0 & i_10_49_3858_0) | (~i_10_49_4050_0 & ~i_10_49_4122_0 & i_10_49_797_0 & ~i_10_49_955_0));
endmodule



// Benchmark "kernel_10_50" written by ABC on Sun Jul 19 10:21:54 2020

module kernel_10_50 ( 
    i_10_50_171_0, i_10_50_172_0, i_10_50_178_0, i_10_50_223_0,
    i_10_50_254_0, i_10_50_270_0, i_10_50_279_0, i_10_50_282_0,
    i_10_50_289_0, i_10_50_317_0, i_10_50_391_0, i_10_50_392_0,
    i_10_50_395_0, i_10_50_409_0, i_10_50_410_0, i_10_50_447_0,
    i_10_50_461_0, i_10_50_464_0, i_10_50_715_0, i_10_50_793_0,
    i_10_50_799_0, i_10_50_956_0, i_10_50_992_0, i_10_50_1027_0,
    i_10_50_1028_0, i_10_50_1030_0, i_10_50_1243_0, i_10_50_1244_0,
    i_10_50_1305_0, i_10_50_1360_0, i_10_50_1433_0, i_10_50_1435_0,
    i_10_50_1436_0, i_10_50_1489_0, i_10_50_1540_0, i_10_50_1541_0,
    i_10_50_1543_0, i_10_50_1544_0, i_10_50_1576_0, i_10_50_1577_0,
    i_10_50_1580_0, i_10_50_1647_0, i_10_50_1655_0, i_10_50_1684_0,
    i_10_50_1685_0, i_10_50_1688_0, i_10_50_1690_0, i_10_50_1820_0,
    i_10_50_1822_0, i_10_50_1823_0, i_10_50_2027_0, i_10_50_2030_0,
    i_10_50_2352_0, i_10_50_2381_0, i_10_50_2470_0, i_10_50_2530_0,
    i_10_50_2628_0, i_10_50_2630_0, i_10_50_2631_0, i_10_50_2632_0,
    i_10_50_2633_0, i_10_50_2634_0, i_10_50_2658_0, i_10_50_2659_0,
    i_10_50_2732_0, i_10_50_2782_0, i_10_50_2834_0, i_10_50_2846_0,
    i_10_50_2963_0, i_10_50_3035_0, i_10_50_3044_0, i_10_50_3071_0,
    i_10_50_3073_0, i_10_50_3155_0, i_10_50_3160_0, i_10_50_3199_0,
    i_10_50_3203_0, i_10_50_3269_0, i_10_50_3332_0, i_10_50_3386_0,
    i_10_50_3391_0, i_10_50_3473_0, i_10_50_3494_0, i_10_50_3522_0,
    i_10_50_3583_0, i_10_50_3586_0, i_10_50_3780_0, i_10_50_3781_0,
    i_10_50_3787_0, i_10_50_3788_0, i_10_50_3838_0, i_10_50_3839_0,
    i_10_50_3841_0, i_10_50_3848_0, i_10_50_3853_0, i_10_50_3982_0,
    i_10_50_4172_0, i_10_50_4277_0, i_10_50_4280_0, i_10_50_4287_0,
    o_10_50_0_0  );
  input  i_10_50_171_0, i_10_50_172_0, i_10_50_178_0, i_10_50_223_0,
    i_10_50_254_0, i_10_50_270_0, i_10_50_279_0, i_10_50_282_0,
    i_10_50_289_0, i_10_50_317_0, i_10_50_391_0, i_10_50_392_0,
    i_10_50_395_0, i_10_50_409_0, i_10_50_410_0, i_10_50_447_0,
    i_10_50_461_0, i_10_50_464_0, i_10_50_715_0, i_10_50_793_0,
    i_10_50_799_0, i_10_50_956_0, i_10_50_992_0, i_10_50_1027_0,
    i_10_50_1028_0, i_10_50_1030_0, i_10_50_1243_0, i_10_50_1244_0,
    i_10_50_1305_0, i_10_50_1360_0, i_10_50_1433_0, i_10_50_1435_0,
    i_10_50_1436_0, i_10_50_1489_0, i_10_50_1540_0, i_10_50_1541_0,
    i_10_50_1543_0, i_10_50_1544_0, i_10_50_1576_0, i_10_50_1577_0,
    i_10_50_1580_0, i_10_50_1647_0, i_10_50_1655_0, i_10_50_1684_0,
    i_10_50_1685_0, i_10_50_1688_0, i_10_50_1690_0, i_10_50_1820_0,
    i_10_50_1822_0, i_10_50_1823_0, i_10_50_2027_0, i_10_50_2030_0,
    i_10_50_2352_0, i_10_50_2381_0, i_10_50_2470_0, i_10_50_2530_0,
    i_10_50_2628_0, i_10_50_2630_0, i_10_50_2631_0, i_10_50_2632_0,
    i_10_50_2633_0, i_10_50_2634_0, i_10_50_2658_0, i_10_50_2659_0,
    i_10_50_2732_0, i_10_50_2782_0, i_10_50_2834_0, i_10_50_2846_0,
    i_10_50_2963_0, i_10_50_3035_0, i_10_50_3044_0, i_10_50_3071_0,
    i_10_50_3073_0, i_10_50_3155_0, i_10_50_3160_0, i_10_50_3199_0,
    i_10_50_3203_0, i_10_50_3269_0, i_10_50_3332_0, i_10_50_3386_0,
    i_10_50_3391_0, i_10_50_3473_0, i_10_50_3494_0, i_10_50_3522_0,
    i_10_50_3583_0, i_10_50_3586_0, i_10_50_3780_0, i_10_50_3781_0,
    i_10_50_3787_0, i_10_50_3788_0, i_10_50_3838_0, i_10_50_3839_0,
    i_10_50_3841_0, i_10_50_3848_0, i_10_50_3853_0, i_10_50_3982_0,
    i_10_50_4172_0, i_10_50_4277_0, i_10_50_4280_0, i_10_50_4287_0;
  output o_10_50_0_0;
  assign o_10_50_0_0 = ~((~i_10_50_254_0 & ((~i_10_50_392_0 & ((~i_10_50_317_0 & ~i_10_50_1244_0 & ~i_10_50_1544_0 & ~i_10_50_3071_0 & ~i_10_50_4277_0) | (~i_10_50_178_0 & i_10_50_279_0 & ~i_10_50_461_0 & ~i_10_50_2027_0 & ~i_10_50_2634_0 & i_10_50_3386_0 & ~i_10_50_4280_0 & ~i_10_50_4287_0))) | (~i_10_50_4277_0 & ((~i_10_50_1028_0 & ~i_10_50_1822_0 & ~i_10_50_2633_0 & ~i_10_50_2834_0 & ~i_10_50_3848_0 & ~i_10_50_4172_0) | (~i_10_50_1647_0 & i_10_50_3044_0 & i_10_50_3848_0 & ~i_10_50_4280_0))))) | (~i_10_50_956_0 & ((~i_10_50_1028_0 & i_10_50_1030_0 & ~i_10_50_2732_0 & ~i_10_50_3044_0 & ~i_10_50_3386_0) | (~i_10_50_395_0 & ~i_10_50_1433_0 & ~i_10_50_1543_0 & i_10_50_2632_0 & ~i_10_50_3787_0))) | (~i_10_50_395_0 & ((~i_10_50_1028_0 & i_10_50_1435_0 & ~i_10_50_2782_0 & ~i_10_50_4277_0) | (~i_10_50_1027_0 & i_10_50_1688_0 & ~i_10_50_3044_0 & ~i_10_50_3071_0 & ~i_10_50_4280_0))) | (~i_10_50_1684_0 & ((~i_10_50_1541_0 & ~i_10_50_2630_0 & ~i_10_50_3199_0 & ~i_10_50_3391_0) | (~i_10_50_172_0 & ~i_10_50_1543_0 & ~i_10_50_1823_0 & ~i_10_50_3071_0 & ~i_10_50_3838_0 & ~i_10_50_4280_0))) | (~i_10_50_1541_0 & ((~i_10_50_1540_0 & ~i_10_50_1647_0 & ~i_10_50_2030_0 & i_10_50_2352_0) | (i_10_50_1305_0 & ~i_10_50_1823_0 & i_10_50_2381_0) | (~i_10_50_1244_0 & i_10_50_2634_0) | (~i_10_50_1028_0 & ~i_10_50_1544_0 & ~i_10_50_1685_0 & ~i_10_50_3203_0) | (~i_10_50_410_0 & i_10_50_1244_0 & ~i_10_50_1433_0 & i_10_50_2628_0 & ~i_10_50_3841_0))) | (~i_10_50_1577_0 & i_10_50_3848_0 & i_10_50_4277_0));
endmodule



// Benchmark "kernel_10_51" written by ABC on Sun Jul 19 10:21:55 2020

module kernel_10_51 ( 
    i_10_51_174_0, i_10_51_279_0, i_10_51_280_0, i_10_51_316_0,
    i_10_51_318_0, i_10_51_319_0, i_10_51_330_0, i_10_51_331_0,
    i_10_51_393_0, i_10_51_409_0, i_10_51_425_0, i_10_51_432_0,
    i_10_51_625_0, i_10_51_712_0, i_10_51_749_0, i_10_51_864_0,
    i_10_51_901_0, i_10_51_902_0, i_10_51_958_0, i_10_51_1030_0,
    i_10_51_1036_0, i_10_51_1037_0, i_10_51_1045_0, i_10_51_1046_0,
    i_10_51_1080_0, i_10_51_1081_0, i_10_51_1084_0, i_10_51_1152_0,
    i_10_51_1153_0, i_10_51_1299_0, i_10_51_1306_0, i_10_51_1347_0,
    i_10_51_1378_0, i_10_51_1433_0, i_10_51_1434_0, i_10_51_1435_0,
    i_10_51_1450_0, i_10_51_1451_0, i_10_51_1541_0, i_10_51_1542_0,
    i_10_51_1543_0, i_10_51_1545_0, i_10_51_1611_0, i_10_51_1623_0,
    i_10_51_1626_0, i_10_51_1629_0, i_10_51_1630_0, i_10_51_1631_0,
    i_10_51_1683_0, i_10_51_1686_0, i_10_51_1714_0, i_10_51_1818_0,
    i_10_51_1914_0, i_10_51_1915_0, i_10_51_1956_0, i_10_51_2199_0,
    i_10_51_2200_0, i_10_51_2201_0, i_10_51_2349_0, i_10_51_2350_0,
    i_10_51_2355_0, i_10_51_2356_0, i_10_51_2471_0, i_10_51_2565_0,
    i_10_51_2635_0, i_10_51_2677_0, i_10_51_2706_0, i_10_51_2716_0,
    i_10_51_2719_0, i_10_51_2721_0, i_10_51_2833_0, i_10_51_2866_0,
    i_10_51_2881_0, i_10_51_3073_0, i_10_51_3223_0, i_10_51_3276_0,
    i_10_51_3333_0, i_10_51_3384_0, i_10_51_3388_0, i_10_51_3504_0,
    i_10_51_3609_0, i_10_51_3615_0, i_10_51_3649_0, i_10_51_3807_0,
    i_10_51_3841_0, i_10_51_3854_0, i_10_51_3859_0, i_10_51_3860_0,
    i_10_51_3908_0, i_10_51_3925_0, i_10_51_3946_0, i_10_51_3979_0,
    i_10_51_3980_0, i_10_51_4025_0, i_10_51_4173_0, i_10_51_4275_0,
    i_10_51_4276_0, i_10_51_4277_0, i_10_51_4278_0, i_10_51_4281_0,
    o_10_51_0_0  );
  input  i_10_51_174_0, i_10_51_279_0, i_10_51_280_0, i_10_51_316_0,
    i_10_51_318_0, i_10_51_319_0, i_10_51_330_0, i_10_51_331_0,
    i_10_51_393_0, i_10_51_409_0, i_10_51_425_0, i_10_51_432_0,
    i_10_51_625_0, i_10_51_712_0, i_10_51_749_0, i_10_51_864_0,
    i_10_51_901_0, i_10_51_902_0, i_10_51_958_0, i_10_51_1030_0,
    i_10_51_1036_0, i_10_51_1037_0, i_10_51_1045_0, i_10_51_1046_0,
    i_10_51_1080_0, i_10_51_1081_0, i_10_51_1084_0, i_10_51_1152_0,
    i_10_51_1153_0, i_10_51_1299_0, i_10_51_1306_0, i_10_51_1347_0,
    i_10_51_1378_0, i_10_51_1433_0, i_10_51_1434_0, i_10_51_1435_0,
    i_10_51_1450_0, i_10_51_1451_0, i_10_51_1541_0, i_10_51_1542_0,
    i_10_51_1543_0, i_10_51_1545_0, i_10_51_1611_0, i_10_51_1623_0,
    i_10_51_1626_0, i_10_51_1629_0, i_10_51_1630_0, i_10_51_1631_0,
    i_10_51_1683_0, i_10_51_1686_0, i_10_51_1714_0, i_10_51_1818_0,
    i_10_51_1914_0, i_10_51_1915_0, i_10_51_1956_0, i_10_51_2199_0,
    i_10_51_2200_0, i_10_51_2201_0, i_10_51_2349_0, i_10_51_2350_0,
    i_10_51_2355_0, i_10_51_2356_0, i_10_51_2471_0, i_10_51_2565_0,
    i_10_51_2635_0, i_10_51_2677_0, i_10_51_2706_0, i_10_51_2716_0,
    i_10_51_2719_0, i_10_51_2721_0, i_10_51_2833_0, i_10_51_2866_0,
    i_10_51_2881_0, i_10_51_3073_0, i_10_51_3223_0, i_10_51_3276_0,
    i_10_51_3333_0, i_10_51_3384_0, i_10_51_3388_0, i_10_51_3504_0,
    i_10_51_3609_0, i_10_51_3615_0, i_10_51_3649_0, i_10_51_3807_0,
    i_10_51_3841_0, i_10_51_3854_0, i_10_51_3859_0, i_10_51_3860_0,
    i_10_51_3908_0, i_10_51_3925_0, i_10_51_3946_0, i_10_51_3979_0,
    i_10_51_3980_0, i_10_51_4025_0, i_10_51_4173_0, i_10_51_4275_0,
    i_10_51_4276_0, i_10_51_4277_0, i_10_51_4278_0, i_10_51_4281_0;
  output o_10_51_0_0;
  assign o_10_51_0_0 = 0;
endmodule



// Benchmark "kernel_10_52" written by ABC on Sun Jul 19 10:21:56 2020

module kernel_10_52 ( 
    i_10_52_70_0, i_10_52_175_0, i_10_52_178_0, i_10_52_179_0,
    i_10_52_250_0, i_10_52_267_0, i_10_52_269_0, i_10_52_279_0,
    i_10_52_280_0, i_10_52_319_0, i_10_52_323_0, i_10_52_500_0,
    i_10_52_503_0, i_10_52_513_0, i_10_52_514_0, i_10_52_591_0,
    i_10_52_629_0, i_10_52_799_0, i_10_52_907_0, i_10_52_931_0,
    i_10_52_932_0, i_10_52_969_0, i_10_52_1011_0, i_10_52_1029_0,
    i_10_52_1116_0, i_10_52_1223_0, i_10_52_1238_0, i_10_52_1240_0,
    i_10_52_1241_0, i_10_52_1304_0, i_10_52_1309_0, i_10_52_1311_0,
    i_10_52_1313_0, i_10_52_1348_0, i_10_52_1349_0, i_10_52_1436_0,
    i_10_52_1437_0, i_10_52_1438_0, i_10_52_1547_0, i_10_52_1563_0,
    i_10_52_1628_0, i_10_52_1687_0, i_10_52_1689_0, i_10_52_1705_0,
    i_10_52_1808_0, i_10_52_1822_0, i_10_52_1885_0, i_10_52_1908_0,
    i_10_52_1909_0, i_10_52_1960_0, i_10_52_2006_0, i_10_52_2023_0,
    i_10_52_2030_0, i_10_52_2113_0, i_10_52_2322_0, i_10_52_2345_0,
    i_10_52_2348_0, i_10_52_2370_0, i_10_52_2436_0, i_10_52_2451_0,
    i_10_52_2455_0, i_10_52_2456_0, i_10_52_2471_0, i_10_52_2633_0,
    i_10_52_2641_0, i_10_52_2649_0, i_10_52_2663_0, i_10_52_2714_0,
    i_10_52_2725_0, i_10_52_2834_0, i_10_52_2851_0, i_10_52_2883_0,
    i_10_52_2884_0, i_10_52_2887_0, i_10_52_2896_0, i_10_52_2919_0,
    i_10_52_2923_0, i_10_52_3058_0, i_10_52_3077_0, i_10_52_3266_0,
    i_10_52_3270_0, i_10_52_3326_0, i_10_52_3338_0, i_10_52_3469_0,
    i_10_52_3473_0, i_10_52_3590_0, i_10_52_3611_0, i_10_52_3615_0,
    i_10_52_3787_0, i_10_52_3963_0, i_10_52_3991_0, i_10_52_4000_0,
    i_10_52_4011_0, i_10_52_4129_0, i_10_52_4156_0, i_10_52_4175_0,
    i_10_52_4219_0, i_10_52_4273_0, i_10_52_4422_0, i_10_52_4597_0,
    o_10_52_0_0  );
  input  i_10_52_70_0, i_10_52_175_0, i_10_52_178_0, i_10_52_179_0,
    i_10_52_250_0, i_10_52_267_0, i_10_52_269_0, i_10_52_279_0,
    i_10_52_280_0, i_10_52_319_0, i_10_52_323_0, i_10_52_500_0,
    i_10_52_503_0, i_10_52_513_0, i_10_52_514_0, i_10_52_591_0,
    i_10_52_629_0, i_10_52_799_0, i_10_52_907_0, i_10_52_931_0,
    i_10_52_932_0, i_10_52_969_0, i_10_52_1011_0, i_10_52_1029_0,
    i_10_52_1116_0, i_10_52_1223_0, i_10_52_1238_0, i_10_52_1240_0,
    i_10_52_1241_0, i_10_52_1304_0, i_10_52_1309_0, i_10_52_1311_0,
    i_10_52_1313_0, i_10_52_1348_0, i_10_52_1349_0, i_10_52_1436_0,
    i_10_52_1437_0, i_10_52_1438_0, i_10_52_1547_0, i_10_52_1563_0,
    i_10_52_1628_0, i_10_52_1687_0, i_10_52_1689_0, i_10_52_1705_0,
    i_10_52_1808_0, i_10_52_1822_0, i_10_52_1885_0, i_10_52_1908_0,
    i_10_52_1909_0, i_10_52_1960_0, i_10_52_2006_0, i_10_52_2023_0,
    i_10_52_2030_0, i_10_52_2113_0, i_10_52_2322_0, i_10_52_2345_0,
    i_10_52_2348_0, i_10_52_2370_0, i_10_52_2436_0, i_10_52_2451_0,
    i_10_52_2455_0, i_10_52_2456_0, i_10_52_2471_0, i_10_52_2633_0,
    i_10_52_2641_0, i_10_52_2649_0, i_10_52_2663_0, i_10_52_2714_0,
    i_10_52_2725_0, i_10_52_2834_0, i_10_52_2851_0, i_10_52_2883_0,
    i_10_52_2884_0, i_10_52_2887_0, i_10_52_2896_0, i_10_52_2919_0,
    i_10_52_2923_0, i_10_52_3058_0, i_10_52_3077_0, i_10_52_3266_0,
    i_10_52_3270_0, i_10_52_3326_0, i_10_52_3338_0, i_10_52_3469_0,
    i_10_52_3473_0, i_10_52_3590_0, i_10_52_3611_0, i_10_52_3615_0,
    i_10_52_3787_0, i_10_52_3963_0, i_10_52_3991_0, i_10_52_4000_0,
    i_10_52_4011_0, i_10_52_4129_0, i_10_52_4156_0, i_10_52_4175_0,
    i_10_52_4219_0, i_10_52_4273_0, i_10_52_4422_0, i_10_52_4597_0;
  output o_10_52_0_0;
  assign o_10_52_0_0 = 0;
endmodule



// Benchmark "kernel_10_53" written by ABC on Sun Jul 19 10:21:57 2020

module kernel_10_53 ( 
    i_10_53_48_0, i_10_53_135_0, i_10_53_146_0, i_10_53_175_0,
    i_10_53_187_0, i_10_53_216_0, i_10_53_218_0, i_10_53_444_0,
    i_10_53_544_0, i_10_53_792_0, i_10_53_793_0, i_10_53_796_0,
    i_10_53_820_0, i_10_53_981_0, i_10_53_1138_0, i_10_53_1153_0,
    i_10_53_1233_0, i_10_53_1242_0, i_10_53_1245_0, i_10_53_1306_0,
    i_10_53_1307_0, i_10_53_1434_0, i_10_53_1443_0, i_10_53_1444_0,
    i_10_53_1445_0, i_10_53_1485_0, i_10_53_1539_0, i_10_53_1540_0,
    i_10_53_1542_0, i_10_53_1557_0, i_10_53_1575_0, i_10_53_1582_0,
    i_10_53_1632_0, i_10_53_1649_0, i_10_53_1651_0, i_10_53_1791_0,
    i_10_53_1911_0, i_10_53_1912_0, i_10_53_1913_0, i_10_53_1921_0,
    i_10_53_2088_0, i_10_53_2200_0, i_10_53_2214_0, i_10_53_2349_0,
    i_10_53_2352_0, i_10_53_2448_0, i_10_53_2449_0, i_10_53_2469_0,
    i_10_53_2538_0, i_10_53_2604_0, i_10_53_2608_0, i_10_53_2629_0,
    i_10_53_2630_0, i_10_53_2631_0, i_10_53_2632_0, i_10_53_2635_0,
    i_10_53_2658_0, i_10_53_2677_0, i_10_53_2700_0, i_10_53_2703_0,
    i_10_53_2718_0, i_10_53_2721_0, i_10_53_2727_0, i_10_53_2729_0,
    i_10_53_2737_0, i_10_53_2817_0, i_10_53_2828_0, i_10_53_2829_0,
    i_10_53_2910_0, i_10_53_3045_0, i_10_53_3199_0, i_10_53_3231_0,
    i_10_53_3276_0, i_10_53_3280_0, i_10_53_3297_0, i_10_53_3298_0,
    i_10_53_3388_0, i_10_53_3431_0, i_10_53_3505_0, i_10_53_3609_0,
    i_10_53_3612_0, i_10_53_3645_0, i_10_53_3702_0, i_10_53_3729_0,
    i_10_53_3781_0, i_10_53_3783_0, i_10_53_3838_0, i_10_53_3840_0,
    i_10_53_3847_0, i_10_53_3848_0, i_10_53_3852_0, i_10_53_3854_0,
    i_10_53_3874_0, i_10_53_4128_0, i_10_53_4219_0, i_10_53_4266_0,
    i_10_53_4269_0, i_10_53_4276_0, i_10_53_4277_0, i_10_53_4288_0,
    o_10_53_0_0  );
  input  i_10_53_48_0, i_10_53_135_0, i_10_53_146_0, i_10_53_175_0,
    i_10_53_187_0, i_10_53_216_0, i_10_53_218_0, i_10_53_444_0,
    i_10_53_544_0, i_10_53_792_0, i_10_53_793_0, i_10_53_796_0,
    i_10_53_820_0, i_10_53_981_0, i_10_53_1138_0, i_10_53_1153_0,
    i_10_53_1233_0, i_10_53_1242_0, i_10_53_1245_0, i_10_53_1306_0,
    i_10_53_1307_0, i_10_53_1434_0, i_10_53_1443_0, i_10_53_1444_0,
    i_10_53_1445_0, i_10_53_1485_0, i_10_53_1539_0, i_10_53_1540_0,
    i_10_53_1542_0, i_10_53_1557_0, i_10_53_1575_0, i_10_53_1582_0,
    i_10_53_1632_0, i_10_53_1649_0, i_10_53_1651_0, i_10_53_1791_0,
    i_10_53_1911_0, i_10_53_1912_0, i_10_53_1913_0, i_10_53_1921_0,
    i_10_53_2088_0, i_10_53_2200_0, i_10_53_2214_0, i_10_53_2349_0,
    i_10_53_2352_0, i_10_53_2448_0, i_10_53_2449_0, i_10_53_2469_0,
    i_10_53_2538_0, i_10_53_2604_0, i_10_53_2608_0, i_10_53_2629_0,
    i_10_53_2630_0, i_10_53_2631_0, i_10_53_2632_0, i_10_53_2635_0,
    i_10_53_2658_0, i_10_53_2677_0, i_10_53_2700_0, i_10_53_2703_0,
    i_10_53_2718_0, i_10_53_2721_0, i_10_53_2727_0, i_10_53_2729_0,
    i_10_53_2737_0, i_10_53_2817_0, i_10_53_2828_0, i_10_53_2829_0,
    i_10_53_2910_0, i_10_53_3045_0, i_10_53_3199_0, i_10_53_3231_0,
    i_10_53_3276_0, i_10_53_3280_0, i_10_53_3297_0, i_10_53_3298_0,
    i_10_53_3388_0, i_10_53_3431_0, i_10_53_3505_0, i_10_53_3609_0,
    i_10_53_3612_0, i_10_53_3645_0, i_10_53_3702_0, i_10_53_3729_0,
    i_10_53_3781_0, i_10_53_3783_0, i_10_53_3838_0, i_10_53_3840_0,
    i_10_53_3847_0, i_10_53_3848_0, i_10_53_3852_0, i_10_53_3854_0,
    i_10_53_3874_0, i_10_53_4128_0, i_10_53_4219_0, i_10_53_4266_0,
    i_10_53_4269_0, i_10_53_4276_0, i_10_53_4277_0, i_10_53_4288_0;
  output o_10_53_0_0;
  assign o_10_53_0_0 = 0;
endmodule



// Benchmark "kernel_10_54" written by ABC on Sun Jul 19 10:21:58 2020

module kernel_10_54 ( 
    i_10_54_184_0, i_10_54_185_0, i_10_54_188_0, i_10_54_210_0,
    i_10_54_211_0, i_10_54_213_0, i_10_54_220_0, i_10_54_251_0,
    i_10_54_405_0, i_10_54_432_0, i_10_54_441_0, i_10_54_466_0,
    i_10_54_498_0, i_10_54_516_0, i_10_54_577_0, i_10_54_578_0,
    i_10_54_586_0, i_10_54_594_0, i_10_54_694_0, i_10_54_699_0,
    i_10_54_800_0, i_10_54_928_0, i_10_54_960_0, i_10_54_969_0,
    i_10_54_987_0, i_10_54_1065_0, i_10_54_1138_0, i_10_54_1167_0,
    i_10_54_1204_0, i_10_54_1255_0, i_10_54_1256_0, i_10_54_1435_0,
    i_10_54_1545_0, i_10_54_1605_0, i_10_54_1650_0, i_10_54_1758_0,
    i_10_54_1759_0, i_10_54_1826_0, i_10_54_1884_0, i_10_54_1911_0,
    i_10_54_1978_0, i_10_54_1986_0, i_10_54_2158_0, i_10_54_2254_0,
    i_10_54_2323_0, i_10_54_2349_0, i_10_54_2352_0, i_10_54_2360_0,
    i_10_54_2403_0, i_10_54_2455_0, i_10_54_2502_0, i_10_54_2506_0,
    i_10_54_2507_0, i_10_54_2589_0, i_10_54_2598_0, i_10_54_2604_0,
    i_10_54_2632_0, i_10_54_2640_0, i_10_54_2649_0, i_10_54_2663_0,
    i_10_54_2676_0, i_10_54_2701_0, i_10_54_2708_0, i_10_54_2716_0,
    i_10_54_2875_0, i_10_54_2924_0, i_10_54_2983_0, i_10_54_3033_0,
    i_10_54_3051_0, i_10_54_3052_0, i_10_54_3054_0, i_10_54_3268_0,
    i_10_54_3270_0, i_10_54_3271_0, i_10_54_3273_0, i_10_54_3299_0,
    i_10_54_3300_0, i_10_54_3492_0, i_10_54_3493_0, i_10_54_3540_0,
    i_10_54_3541_0, i_10_54_3683_0, i_10_54_3850_0, i_10_54_3888_0,
    i_10_54_3963_0, i_10_54_4090_0, i_10_54_4130_0, i_10_54_4188_0,
    i_10_54_4219_0, i_10_54_4220_0, i_10_54_4230_0, i_10_54_4233_0,
    i_10_54_4234_0, i_10_54_4279_0, i_10_54_4459_0, i_10_54_4461_0,
    i_10_54_4513_0, i_10_54_4564_0, i_10_54_4565_0, i_10_54_4571_0,
    o_10_54_0_0  );
  input  i_10_54_184_0, i_10_54_185_0, i_10_54_188_0, i_10_54_210_0,
    i_10_54_211_0, i_10_54_213_0, i_10_54_220_0, i_10_54_251_0,
    i_10_54_405_0, i_10_54_432_0, i_10_54_441_0, i_10_54_466_0,
    i_10_54_498_0, i_10_54_516_0, i_10_54_577_0, i_10_54_578_0,
    i_10_54_586_0, i_10_54_594_0, i_10_54_694_0, i_10_54_699_0,
    i_10_54_800_0, i_10_54_928_0, i_10_54_960_0, i_10_54_969_0,
    i_10_54_987_0, i_10_54_1065_0, i_10_54_1138_0, i_10_54_1167_0,
    i_10_54_1204_0, i_10_54_1255_0, i_10_54_1256_0, i_10_54_1435_0,
    i_10_54_1545_0, i_10_54_1605_0, i_10_54_1650_0, i_10_54_1758_0,
    i_10_54_1759_0, i_10_54_1826_0, i_10_54_1884_0, i_10_54_1911_0,
    i_10_54_1978_0, i_10_54_1986_0, i_10_54_2158_0, i_10_54_2254_0,
    i_10_54_2323_0, i_10_54_2349_0, i_10_54_2352_0, i_10_54_2360_0,
    i_10_54_2403_0, i_10_54_2455_0, i_10_54_2502_0, i_10_54_2506_0,
    i_10_54_2507_0, i_10_54_2589_0, i_10_54_2598_0, i_10_54_2604_0,
    i_10_54_2632_0, i_10_54_2640_0, i_10_54_2649_0, i_10_54_2663_0,
    i_10_54_2676_0, i_10_54_2701_0, i_10_54_2708_0, i_10_54_2716_0,
    i_10_54_2875_0, i_10_54_2924_0, i_10_54_2983_0, i_10_54_3033_0,
    i_10_54_3051_0, i_10_54_3052_0, i_10_54_3054_0, i_10_54_3268_0,
    i_10_54_3270_0, i_10_54_3271_0, i_10_54_3273_0, i_10_54_3299_0,
    i_10_54_3300_0, i_10_54_3492_0, i_10_54_3493_0, i_10_54_3540_0,
    i_10_54_3541_0, i_10_54_3683_0, i_10_54_3850_0, i_10_54_3888_0,
    i_10_54_3963_0, i_10_54_4090_0, i_10_54_4130_0, i_10_54_4188_0,
    i_10_54_4219_0, i_10_54_4220_0, i_10_54_4230_0, i_10_54_4233_0,
    i_10_54_4234_0, i_10_54_4279_0, i_10_54_4459_0, i_10_54_4461_0,
    i_10_54_4513_0, i_10_54_4564_0, i_10_54_4565_0, i_10_54_4571_0;
  output o_10_54_0_0;
  assign o_10_54_0_0 = 0;
endmodule



// Benchmark "kernel_10_55" written by ABC on Sun Jul 19 10:21:58 2020

module kernel_10_55 ( 
    i_10_55_29_0, i_10_55_89_0, i_10_55_120_0, i_10_55_387_0,
    i_10_55_388_0, i_10_55_390_0, i_10_55_391_0, i_10_55_426_0,
    i_10_55_459_0, i_10_55_460_0, i_10_55_461_0, i_10_55_558_0,
    i_10_55_559_0, i_10_55_689_0, i_10_55_747_0, i_10_55_748_0,
    i_10_55_750_0, i_10_55_752_0, i_10_55_919_0, i_10_55_985_0,
    i_10_55_999_0, i_10_55_1048_0, i_10_55_1053_0, i_10_55_1054_0,
    i_10_55_1236_0, i_10_55_1237_0, i_10_55_1305_0, i_10_55_1309_0,
    i_10_55_1362_0, i_10_55_1381_0, i_10_55_1455_0, i_10_55_1578_0,
    i_10_55_1611_0, i_10_55_1612_0, i_10_55_1613_0, i_10_55_1643_0,
    i_10_55_1764_0, i_10_55_1765_0, i_10_55_1822_0, i_10_55_1826_0,
    i_10_55_1945_0, i_10_55_1947_0, i_10_55_1953_0, i_10_55_1954_0,
    i_10_55_1996_0, i_10_55_2062_0, i_10_55_2108_0, i_10_55_2179_0,
    i_10_55_2406_0, i_10_55_2413_0, i_10_55_2455_0, i_10_55_2456_0,
    i_10_55_2478_0, i_10_55_2613_0, i_10_55_2655_0, i_10_55_2659_0,
    i_10_55_2661_0, i_10_55_2688_0, i_10_55_2689_0, i_10_55_2710_0,
    i_10_55_2730_0, i_10_55_2817_0, i_10_55_2911_0, i_10_55_3036_0,
    i_10_55_3037_0, i_10_55_3043_0, i_10_55_3076_0, i_10_55_3090_0,
    i_10_55_3195_0, i_10_55_3196_0, i_10_55_3348_0, i_10_55_3349_0,
    i_10_55_3352_0, i_10_55_3469_0, i_10_55_3470_0, i_10_55_3585_0,
    i_10_55_3618_0, i_10_55_3619_0, i_10_55_3620_0, i_10_55_3637_0,
    i_10_55_3645_0, i_10_55_3646_0, i_10_55_3647_0, i_10_55_3732_0,
    i_10_55_3853_0, i_10_55_3854_0, i_10_55_3879_0, i_10_55_3880_0,
    i_10_55_3942_0, i_10_55_3988_0, i_10_55_4025_0, i_10_55_4028_0,
    i_10_55_4029_0, i_10_55_4030_0, i_10_55_4051_0, i_10_55_4053_0,
    i_10_55_4275_0, i_10_55_4341_0, i_10_55_4530_0, i_10_55_4586_0,
    o_10_55_0_0  );
  input  i_10_55_29_0, i_10_55_89_0, i_10_55_120_0, i_10_55_387_0,
    i_10_55_388_0, i_10_55_390_0, i_10_55_391_0, i_10_55_426_0,
    i_10_55_459_0, i_10_55_460_0, i_10_55_461_0, i_10_55_558_0,
    i_10_55_559_0, i_10_55_689_0, i_10_55_747_0, i_10_55_748_0,
    i_10_55_750_0, i_10_55_752_0, i_10_55_919_0, i_10_55_985_0,
    i_10_55_999_0, i_10_55_1048_0, i_10_55_1053_0, i_10_55_1054_0,
    i_10_55_1236_0, i_10_55_1237_0, i_10_55_1305_0, i_10_55_1309_0,
    i_10_55_1362_0, i_10_55_1381_0, i_10_55_1455_0, i_10_55_1578_0,
    i_10_55_1611_0, i_10_55_1612_0, i_10_55_1613_0, i_10_55_1643_0,
    i_10_55_1764_0, i_10_55_1765_0, i_10_55_1822_0, i_10_55_1826_0,
    i_10_55_1945_0, i_10_55_1947_0, i_10_55_1953_0, i_10_55_1954_0,
    i_10_55_1996_0, i_10_55_2062_0, i_10_55_2108_0, i_10_55_2179_0,
    i_10_55_2406_0, i_10_55_2413_0, i_10_55_2455_0, i_10_55_2456_0,
    i_10_55_2478_0, i_10_55_2613_0, i_10_55_2655_0, i_10_55_2659_0,
    i_10_55_2661_0, i_10_55_2688_0, i_10_55_2689_0, i_10_55_2710_0,
    i_10_55_2730_0, i_10_55_2817_0, i_10_55_2911_0, i_10_55_3036_0,
    i_10_55_3037_0, i_10_55_3043_0, i_10_55_3076_0, i_10_55_3090_0,
    i_10_55_3195_0, i_10_55_3196_0, i_10_55_3348_0, i_10_55_3349_0,
    i_10_55_3352_0, i_10_55_3469_0, i_10_55_3470_0, i_10_55_3585_0,
    i_10_55_3618_0, i_10_55_3619_0, i_10_55_3620_0, i_10_55_3637_0,
    i_10_55_3645_0, i_10_55_3646_0, i_10_55_3647_0, i_10_55_3732_0,
    i_10_55_3853_0, i_10_55_3854_0, i_10_55_3879_0, i_10_55_3880_0,
    i_10_55_3942_0, i_10_55_3988_0, i_10_55_4025_0, i_10_55_4028_0,
    i_10_55_4029_0, i_10_55_4030_0, i_10_55_4051_0, i_10_55_4053_0,
    i_10_55_4275_0, i_10_55_4341_0, i_10_55_4530_0, i_10_55_4586_0;
  output o_10_55_0_0;
  assign o_10_55_0_0 = 0;
endmodule



// Benchmark "kernel_10_56" written by ABC on Sun Jul 19 10:21:59 2020

module kernel_10_56 ( 
    i_10_56_27_0, i_10_56_33_0, i_10_56_34_0, i_10_56_52_0, i_10_56_172_0,
    i_10_56_178_0, i_10_56_224_0, i_10_56_258_0, i_10_56_282_0,
    i_10_56_366_0, i_10_56_390_0, i_10_56_408_0, i_10_56_409_0,
    i_10_56_442_0, i_10_56_445_0, i_10_56_498_0, i_10_56_502_0,
    i_10_56_541_0, i_10_56_602_0, i_10_56_798_0, i_10_56_954_0,
    i_10_56_958_0, i_10_56_960_0, i_10_56_990_0, i_10_56_991_0,
    i_10_56_992_0, i_10_56_1033_0, i_10_56_1083_0, i_10_56_1088_0,
    i_10_56_1164_0, i_10_56_1250_0, i_10_56_1305_0, i_10_56_1306_0,
    i_10_56_1308_0, i_10_56_1309_0, i_10_56_1381_0, i_10_56_1443_0,
    i_10_56_1545_0, i_10_56_1686_0, i_10_56_1715_0, i_10_56_1770_0,
    i_10_56_1813_0, i_10_56_1854_0, i_10_56_1908_0, i_10_56_2005_0,
    i_10_56_2006_0, i_10_56_2254_0, i_10_56_2353_0, i_10_56_2380_0,
    i_10_56_2460_0, i_10_56_2536_0, i_10_56_2606_0, i_10_56_2632_0,
    i_10_56_2634_0, i_10_56_2704_0, i_10_56_2714_0, i_10_56_2722_0,
    i_10_56_2731_0, i_10_56_2742_0, i_10_56_2826_0, i_10_56_2829_0,
    i_10_56_2884_0, i_10_56_2920_0, i_10_56_2923_0, i_10_56_2986_0,
    i_10_56_3033_0, i_10_56_3072_0, i_10_56_3076_0, i_10_56_3165_0,
    i_10_56_3200_0, i_10_56_3201_0, i_10_56_3282_0, i_10_56_3298_0,
    i_10_56_3330_0, i_10_56_3333_0, i_10_56_3336_0, i_10_56_3405_0,
    i_10_56_3406_0, i_10_56_3408_0, i_10_56_3441_0, i_10_56_3466_0,
    i_10_56_3609_0, i_10_56_3612_0, i_10_56_3616_0, i_10_56_3618_0,
    i_10_56_3624_0, i_10_56_3625_0, i_10_56_3649_0, i_10_56_3652_0,
    i_10_56_3653_0, i_10_56_3780_0, i_10_56_3783_0, i_10_56_3784_0,
    i_10_56_3844_0, i_10_56_3847_0, i_10_56_3853_0, i_10_56_3947_0,
    i_10_56_4126_0, i_10_56_4288_0, i_10_56_4567_0,
    o_10_56_0_0  );
  input  i_10_56_27_0, i_10_56_33_0, i_10_56_34_0, i_10_56_52_0,
    i_10_56_172_0, i_10_56_178_0, i_10_56_224_0, i_10_56_258_0,
    i_10_56_282_0, i_10_56_366_0, i_10_56_390_0, i_10_56_408_0,
    i_10_56_409_0, i_10_56_442_0, i_10_56_445_0, i_10_56_498_0,
    i_10_56_502_0, i_10_56_541_0, i_10_56_602_0, i_10_56_798_0,
    i_10_56_954_0, i_10_56_958_0, i_10_56_960_0, i_10_56_990_0,
    i_10_56_991_0, i_10_56_992_0, i_10_56_1033_0, i_10_56_1083_0,
    i_10_56_1088_0, i_10_56_1164_0, i_10_56_1250_0, i_10_56_1305_0,
    i_10_56_1306_0, i_10_56_1308_0, i_10_56_1309_0, i_10_56_1381_0,
    i_10_56_1443_0, i_10_56_1545_0, i_10_56_1686_0, i_10_56_1715_0,
    i_10_56_1770_0, i_10_56_1813_0, i_10_56_1854_0, i_10_56_1908_0,
    i_10_56_2005_0, i_10_56_2006_0, i_10_56_2254_0, i_10_56_2353_0,
    i_10_56_2380_0, i_10_56_2460_0, i_10_56_2536_0, i_10_56_2606_0,
    i_10_56_2632_0, i_10_56_2634_0, i_10_56_2704_0, i_10_56_2714_0,
    i_10_56_2722_0, i_10_56_2731_0, i_10_56_2742_0, i_10_56_2826_0,
    i_10_56_2829_0, i_10_56_2884_0, i_10_56_2920_0, i_10_56_2923_0,
    i_10_56_2986_0, i_10_56_3033_0, i_10_56_3072_0, i_10_56_3076_0,
    i_10_56_3165_0, i_10_56_3200_0, i_10_56_3201_0, i_10_56_3282_0,
    i_10_56_3298_0, i_10_56_3330_0, i_10_56_3333_0, i_10_56_3336_0,
    i_10_56_3405_0, i_10_56_3406_0, i_10_56_3408_0, i_10_56_3441_0,
    i_10_56_3466_0, i_10_56_3609_0, i_10_56_3612_0, i_10_56_3616_0,
    i_10_56_3618_0, i_10_56_3624_0, i_10_56_3625_0, i_10_56_3649_0,
    i_10_56_3652_0, i_10_56_3653_0, i_10_56_3780_0, i_10_56_3783_0,
    i_10_56_3784_0, i_10_56_3844_0, i_10_56_3847_0, i_10_56_3853_0,
    i_10_56_3947_0, i_10_56_4126_0, i_10_56_4288_0, i_10_56_4567_0;
  output o_10_56_0_0;
  assign o_10_56_0_0 = 0;
endmodule



// Benchmark "kernel_10_57" written by ABC on Sun Jul 19 10:22:00 2020

module kernel_10_57 ( 
    i_10_57_52_0, i_10_57_178_0, i_10_57_224_0, i_10_57_275_0,
    i_10_57_277_0, i_10_57_281_0, i_10_57_283_0, i_10_57_287_0,
    i_10_57_408_0, i_10_57_446_0, i_10_57_730_0, i_10_57_797_0,
    i_10_57_898_0, i_10_57_958_0, i_10_57_996_0, i_10_57_997_0,
    i_10_57_1033_0, i_10_57_1034_0, i_10_57_1247_0, i_10_57_1306_0,
    i_10_57_1311_0, i_10_57_1363_0, i_10_57_1543_0, i_10_57_1553_0,
    i_10_57_1579_0, i_10_57_1626_0, i_10_57_1654_0, i_10_57_1689_0,
    i_10_57_1690_0, i_10_57_1736_0, i_10_57_1819_0, i_10_57_1820_0,
    i_10_57_1821_0, i_10_57_1822_0, i_10_57_1826_0, i_10_57_1909_0,
    i_10_57_1912_0, i_10_57_1996_0, i_10_57_1997_0, i_10_57_2019_0,
    i_10_57_2028_0, i_10_57_2031_0, i_10_57_2352_0, i_10_57_2353_0,
    i_10_57_2355_0, i_10_57_2449_0, i_10_57_2452_0, i_10_57_2454_0,
    i_10_57_2455_0, i_10_57_2474_0, i_10_57_2565_0, i_10_57_2568_0,
    i_10_57_2572_0, i_10_57_2662_0, i_10_57_2705_0, i_10_57_2716_0,
    i_10_57_2717_0, i_10_57_2721_0, i_10_57_2725_0, i_10_57_2732_0,
    i_10_57_2734_0, i_10_57_2880_0, i_10_57_2884_0, i_10_57_2917_0,
    i_10_57_2918_0, i_10_57_2920_0, i_10_57_2964_0, i_10_57_3038_0,
    i_10_57_3049_0, i_10_57_3054_0, i_10_57_3197_0, i_10_57_3277_0,
    i_10_57_3384_0, i_10_57_3385_0, i_10_57_3388_0, i_10_57_3391_0,
    i_10_57_3405_0, i_10_57_3406_0, i_10_57_3501_0, i_10_57_3525_0,
    i_10_57_3589_0, i_10_57_3610_0, i_10_57_3613_0, i_10_57_3614_0,
    i_10_57_3617_0, i_10_57_3653_0, i_10_57_3720_0, i_10_57_3780_0,
    i_10_57_3781_0, i_10_57_3784_0, i_10_57_3834_0, i_10_57_3837_0,
    i_10_57_3839_0, i_10_57_3857_0, i_10_57_3896_0, i_10_57_3982_0,
    i_10_57_4030_0, i_10_57_4266_0, i_10_57_4291_0, i_10_57_4567_0,
    o_10_57_0_0  );
  input  i_10_57_52_0, i_10_57_178_0, i_10_57_224_0, i_10_57_275_0,
    i_10_57_277_0, i_10_57_281_0, i_10_57_283_0, i_10_57_287_0,
    i_10_57_408_0, i_10_57_446_0, i_10_57_730_0, i_10_57_797_0,
    i_10_57_898_0, i_10_57_958_0, i_10_57_996_0, i_10_57_997_0,
    i_10_57_1033_0, i_10_57_1034_0, i_10_57_1247_0, i_10_57_1306_0,
    i_10_57_1311_0, i_10_57_1363_0, i_10_57_1543_0, i_10_57_1553_0,
    i_10_57_1579_0, i_10_57_1626_0, i_10_57_1654_0, i_10_57_1689_0,
    i_10_57_1690_0, i_10_57_1736_0, i_10_57_1819_0, i_10_57_1820_0,
    i_10_57_1821_0, i_10_57_1822_0, i_10_57_1826_0, i_10_57_1909_0,
    i_10_57_1912_0, i_10_57_1996_0, i_10_57_1997_0, i_10_57_2019_0,
    i_10_57_2028_0, i_10_57_2031_0, i_10_57_2352_0, i_10_57_2353_0,
    i_10_57_2355_0, i_10_57_2449_0, i_10_57_2452_0, i_10_57_2454_0,
    i_10_57_2455_0, i_10_57_2474_0, i_10_57_2565_0, i_10_57_2568_0,
    i_10_57_2572_0, i_10_57_2662_0, i_10_57_2705_0, i_10_57_2716_0,
    i_10_57_2717_0, i_10_57_2721_0, i_10_57_2725_0, i_10_57_2732_0,
    i_10_57_2734_0, i_10_57_2880_0, i_10_57_2884_0, i_10_57_2917_0,
    i_10_57_2918_0, i_10_57_2920_0, i_10_57_2964_0, i_10_57_3038_0,
    i_10_57_3049_0, i_10_57_3054_0, i_10_57_3197_0, i_10_57_3277_0,
    i_10_57_3384_0, i_10_57_3385_0, i_10_57_3388_0, i_10_57_3391_0,
    i_10_57_3405_0, i_10_57_3406_0, i_10_57_3501_0, i_10_57_3525_0,
    i_10_57_3589_0, i_10_57_3610_0, i_10_57_3613_0, i_10_57_3614_0,
    i_10_57_3617_0, i_10_57_3653_0, i_10_57_3720_0, i_10_57_3780_0,
    i_10_57_3781_0, i_10_57_3784_0, i_10_57_3834_0, i_10_57_3837_0,
    i_10_57_3839_0, i_10_57_3857_0, i_10_57_3896_0, i_10_57_3982_0,
    i_10_57_4030_0, i_10_57_4266_0, i_10_57_4291_0, i_10_57_4567_0;
  output o_10_57_0_0;
  assign o_10_57_0_0 = 0;
endmodule



// Benchmark "kernel_10_58" written by ABC on Sun Jul 19 10:22:02 2020

module kernel_10_58 ( 
    i_10_58_174_0, i_10_58_179_0, i_10_58_279_0, i_10_58_280_0,
    i_10_58_290_0, i_10_58_317_0, i_10_58_328_0, i_10_58_406_0,
    i_10_58_407_0, i_10_58_443_0, i_10_58_712_0, i_10_58_713_0,
    i_10_58_748_0, i_10_58_749_0, i_10_58_797_0, i_10_58_893_0,
    i_10_58_955_0, i_10_58_1000_0, i_10_58_1001_0, i_10_58_1033_0,
    i_10_58_1308_0, i_10_58_1309_0, i_10_58_1310_0, i_10_58_1360_0,
    i_10_58_1540_0, i_10_58_1541_0, i_10_58_1647_0, i_10_58_1649_0,
    i_10_58_1651_0, i_10_58_1652_0, i_10_58_1683_0, i_10_58_1684_0,
    i_10_58_1685_0, i_10_58_1687_0, i_10_58_1688_0, i_10_58_1721_0,
    i_10_58_1729_0, i_10_58_1819_0, i_10_58_1820_0, i_10_58_1826_0,
    i_10_58_1946_0, i_10_58_1949_0, i_10_58_1989_0, i_10_58_1999_0,
    i_10_58_2180_0, i_10_58_2198_0, i_10_58_2351_0, i_10_58_2354_0,
    i_10_58_2358_0, i_10_58_2377_0, i_10_58_2449_0, i_10_58_2450_0,
    i_10_58_2452_0, i_10_58_2632_0, i_10_58_2674_0, i_10_58_2716_0,
    i_10_58_2720_0, i_10_58_2723_0, i_10_58_2738_0, i_10_58_2782_0,
    i_10_58_2785_0, i_10_58_2828_0, i_10_58_2829_0, i_10_58_2917_0,
    i_10_58_2918_0, i_10_58_3034_0, i_10_58_3035_0, i_10_58_3036_0,
    i_10_58_3037_0, i_10_58_3038_0, i_10_58_3042_0, i_10_58_3043_0,
    i_10_58_3087_0, i_10_58_3153_0, i_10_58_3406_0, i_10_58_3407_0,
    i_10_58_3550_0, i_10_58_3613_0, i_10_58_3614_0, i_10_58_3648_0,
    i_10_58_3650_0, i_10_58_3834_0, i_10_58_3838_0, i_10_58_3847_0,
    i_10_58_3848_0, i_10_58_3852_0, i_10_58_3854_0, i_10_58_3856_0,
    i_10_58_3857_0, i_10_58_3907_0, i_10_58_3910_0, i_10_58_3992_0,
    i_10_58_4113_0, i_10_58_4122_0, i_10_58_4125_0, i_10_58_4564_0,
    i_10_58_4565_0, i_10_58_4566_0, i_10_58_4567_0, i_10_58_4568_0,
    o_10_58_0_0  );
  input  i_10_58_174_0, i_10_58_179_0, i_10_58_279_0, i_10_58_280_0,
    i_10_58_290_0, i_10_58_317_0, i_10_58_328_0, i_10_58_406_0,
    i_10_58_407_0, i_10_58_443_0, i_10_58_712_0, i_10_58_713_0,
    i_10_58_748_0, i_10_58_749_0, i_10_58_797_0, i_10_58_893_0,
    i_10_58_955_0, i_10_58_1000_0, i_10_58_1001_0, i_10_58_1033_0,
    i_10_58_1308_0, i_10_58_1309_0, i_10_58_1310_0, i_10_58_1360_0,
    i_10_58_1540_0, i_10_58_1541_0, i_10_58_1647_0, i_10_58_1649_0,
    i_10_58_1651_0, i_10_58_1652_0, i_10_58_1683_0, i_10_58_1684_0,
    i_10_58_1685_0, i_10_58_1687_0, i_10_58_1688_0, i_10_58_1721_0,
    i_10_58_1729_0, i_10_58_1819_0, i_10_58_1820_0, i_10_58_1826_0,
    i_10_58_1946_0, i_10_58_1949_0, i_10_58_1989_0, i_10_58_1999_0,
    i_10_58_2180_0, i_10_58_2198_0, i_10_58_2351_0, i_10_58_2354_0,
    i_10_58_2358_0, i_10_58_2377_0, i_10_58_2449_0, i_10_58_2450_0,
    i_10_58_2452_0, i_10_58_2632_0, i_10_58_2674_0, i_10_58_2716_0,
    i_10_58_2720_0, i_10_58_2723_0, i_10_58_2738_0, i_10_58_2782_0,
    i_10_58_2785_0, i_10_58_2828_0, i_10_58_2829_0, i_10_58_2917_0,
    i_10_58_2918_0, i_10_58_3034_0, i_10_58_3035_0, i_10_58_3036_0,
    i_10_58_3037_0, i_10_58_3038_0, i_10_58_3042_0, i_10_58_3043_0,
    i_10_58_3087_0, i_10_58_3153_0, i_10_58_3406_0, i_10_58_3407_0,
    i_10_58_3550_0, i_10_58_3613_0, i_10_58_3614_0, i_10_58_3648_0,
    i_10_58_3650_0, i_10_58_3834_0, i_10_58_3838_0, i_10_58_3847_0,
    i_10_58_3848_0, i_10_58_3852_0, i_10_58_3854_0, i_10_58_3856_0,
    i_10_58_3857_0, i_10_58_3907_0, i_10_58_3910_0, i_10_58_3992_0,
    i_10_58_4113_0, i_10_58_4122_0, i_10_58_4125_0, i_10_58_4564_0,
    i_10_58_4565_0, i_10_58_4566_0, i_10_58_4567_0, i_10_58_4568_0;
  output o_10_58_0_0;
  assign o_10_58_0_0 = ~((i_10_58_174_0 & ((~i_10_58_1688_0 & ~i_10_58_2452_0 & i_10_58_3406_0) | (~i_10_58_407_0 & ~i_10_58_748_0 & ~i_10_58_1651_0 & ~i_10_58_1685_0 & ~i_10_58_1729_0 & ~i_10_58_2785_0 & ~i_10_58_2828_0 & ~i_10_58_3038_0 & ~i_10_58_3407_0 & ~i_10_58_3907_0))) | (~i_10_58_280_0 & ((~i_10_58_1540_0 & i_10_58_1683_0 & ~i_10_58_1688_0 & i_10_58_1819_0 & i_10_58_3406_0 & ~i_10_58_3650_0) | (~i_10_58_713_0 & ~i_10_58_1687_0 & ~i_10_58_2180_0 & ~i_10_58_3838_0 & ~i_10_58_3907_0 & ~i_10_58_3992_0 & ~i_10_58_4113_0))) | (~i_10_58_1684_0 & ((~i_10_58_179_0 & ((~i_10_58_317_0 & ~i_10_58_1033_0 & ~i_10_58_1540_0 & ~i_10_58_1649_0 & ~i_10_58_1999_0 & ~i_10_58_3407_0 & ~i_10_58_3614_0) | (~i_10_58_1652_0 & ~i_10_58_2723_0 & ~i_10_58_3038_0 & ~i_10_58_3406_0 & i_10_58_3838_0 & ~i_10_58_3910_0))) | (~i_10_58_2716_0 & ((~i_10_58_328_0 & ((~i_10_58_1647_0 & ~i_10_58_1688_0 & ~i_10_58_1999_0 & ~i_10_58_2829_0 & ~i_10_58_3034_0 & ~i_10_58_3857_0 & ~i_10_58_3907_0) | (~i_10_58_713_0 & ~i_10_58_1826_0 & ~i_10_58_2198_0 & ~i_10_58_2354_0 & ~i_10_58_2452_0 & ~i_10_58_4113_0))) | (~i_10_58_749_0 & i_10_58_1308_0 & ~i_10_58_1540_0 & ~i_10_58_1826_0 & ~i_10_58_2351_0))) | (~i_10_58_1652_0 & (i_10_58_4125_0 | (~i_10_58_797_0 & ~i_10_58_1308_0 & ~i_10_58_3037_0 & i_10_58_3614_0))) | (~i_10_58_1683_0 & ((~i_10_58_713_0 & ~i_10_58_749_0 & ~i_10_58_1649_0 & i_10_58_3854_0) | (~i_10_58_712_0 & i_10_58_3852_0 & ~i_10_58_3907_0))))) | (~i_10_58_3406_0 & ((~i_10_58_174_0 & ((~i_10_58_179_0 & ~i_10_58_797_0 & ~i_10_58_1826_0 & ~i_10_58_2351_0 & ~i_10_58_2450_0 & i_10_58_3037_0 & ~i_10_58_3847_0) | (~i_10_58_748_0 & ~i_10_58_749_0 & ~i_10_58_955_0 & ~i_10_58_1001_0 & ~i_10_58_1310_0 & ~i_10_58_1652_0 & ~i_10_58_2449_0 & ~i_10_58_2674_0 & ~i_10_58_2782_0 & ~i_10_58_2785_0 & ~i_10_58_3034_0 & ~i_10_58_3035_0 & ~i_10_58_3907_0 & ~i_10_58_4568_0))) | (~i_10_58_749_0 & ((~i_10_58_1649_0 & ~i_10_58_1687_0 & ~i_10_58_2716_0 & i_10_58_3037_0) | (~i_10_58_179_0 & ~i_10_58_712_0 & ~i_10_58_797_0 & ~i_10_58_1541_0 & ~i_10_58_2723_0 & ~i_10_58_3613_0 & ~i_10_58_3857_0 & ~i_10_58_4122_0))) | (i_10_58_1826_0 & i_10_58_2785_0 & ~i_10_58_3910_0))) | (~i_10_58_955_0 & ((~i_10_58_317_0 & ~i_10_58_713_0 & ~i_10_58_748_0 & ~i_10_58_1033_0 & ~i_10_58_1310_0 & ~i_10_58_1647_0 & i_10_58_1819_0 & ~i_10_58_2828_0 & ~i_10_58_3037_0) | (~i_10_58_712_0 & ~i_10_58_1541_0 & i_10_58_2358_0 & ~i_10_58_3648_0 & ~i_10_58_3848_0))) | (~i_10_58_317_0 & ((~i_10_58_1651_0 & ~i_10_58_1685_0 & i_10_58_2354_0 & ~i_10_58_2716_0 & ~i_10_58_2723_0) | (~i_10_58_712_0 & ~i_10_58_1309_0 & ~i_10_58_1541_0 & i_10_58_1651_0 & i_10_58_1652_0 & ~i_10_58_1683_0 & ~i_10_58_1729_0 & ~i_10_58_2452_0 & ~i_10_58_3613_0 & ~i_10_58_4565_0 & ~i_10_58_4567_0))) | (~i_10_58_712_0 & ((~i_10_58_748_0 & ~i_10_58_797_0 & i_10_58_1308_0 & ~i_10_58_1688_0 & ~i_10_58_2723_0 & ~i_10_58_3407_0) | (~i_10_58_1540_0 & ~i_10_58_2180_0 & i_10_58_2632_0 & ~i_10_58_2716_0 & ~i_10_58_2720_0 & ~i_10_58_3856_0 & ~i_10_58_3907_0))) | (~i_10_58_713_0 & ((i_10_58_1826_0 & i_10_58_2782_0 & ~i_10_58_3614_0 & ~i_10_58_3907_0) | (~i_10_58_748_0 & ~i_10_58_1308_0 & i_10_58_1819_0 & ~i_10_58_2198_0 & ~i_10_58_2716_0 & ~i_10_58_3038_0 & ~i_10_58_3407_0 & ~i_10_58_3648_0 & ~i_10_58_4122_0))) | (~i_10_58_749_0 & ((~i_10_58_3613_0 & ((~i_10_58_1647_0 & ~i_10_58_1729_0 & ~i_10_58_2716_0 & i_10_58_3034_0) | (~i_10_58_1688_0 & ~i_10_58_2198_0 & ~i_10_58_2452_0 & ~i_10_58_3407_0 & ~i_10_58_3992_0))) | (~i_10_58_3838_0 & i_10_58_4568_0))) | (~i_10_58_1652_0 & ((i_10_58_2829_0 & i_10_58_3648_0) | (i_10_58_1033_0 & i_10_58_3650_0) | (~i_10_58_174_0 & ~i_10_58_1310_0 & ~i_10_58_1683_0 & i_10_58_2716_0 & i_10_58_3406_0 & ~i_10_58_3857_0))) | (i_10_58_179_0 & i_10_58_2785_0 & i_10_58_3037_0 & ~i_10_58_3613_0));
endmodule



// Benchmark "kernel_10_59" written by ABC on Sun Jul 19 10:22:02 2020

module kernel_10_59 ( 
    i_10_59_150_0, i_10_59_180_0, i_10_59_286_0, i_10_59_319_0,
    i_10_59_461_0, i_10_59_588_0, i_10_59_592_0, i_10_59_633_0,
    i_10_59_692_0, i_10_59_735_0, i_10_59_798_0, i_10_59_799_0,
    i_10_59_828_0, i_10_59_831_0, i_10_59_929_0, i_10_59_961_0,
    i_10_59_962_0, i_10_59_1040_0, i_10_59_1041_0, i_10_59_1120_0,
    i_10_59_1167_0, i_10_59_1180_0, i_10_59_1306_0, i_10_59_1344_0,
    i_10_59_1346_0, i_10_59_1365_0, i_10_59_1366_0, i_10_59_1554_0,
    i_10_59_1570_0, i_10_59_1648_0, i_10_59_1744_0, i_10_59_1769_0,
    i_10_59_1771_0, i_10_59_1785_0, i_10_59_1788_0, i_10_59_1791_0,
    i_10_59_2011_0, i_10_59_2012_0, i_10_59_2025_0, i_10_59_2142_0,
    i_10_59_2380_0, i_10_59_2389_0, i_10_59_2437_0, i_10_59_2438_0,
    i_10_59_2452_0, i_10_59_2478_0, i_10_59_2479_0, i_10_59_2480_0,
    i_10_59_2542_0, i_10_59_2636_0, i_10_59_2652_0, i_10_59_2713_0,
    i_10_59_2818_0, i_10_59_2828_0, i_10_59_2831_0, i_10_59_2844_0,
    i_10_59_2848_0, i_10_59_2883_0, i_10_59_2910_0, i_10_59_2911_0,
    i_10_59_2922_0, i_10_59_2923_0, i_10_59_2938_0, i_10_59_2958_0,
    i_10_59_2959_0, i_10_59_2978_0, i_10_59_2986_0, i_10_59_3046_0,
    i_10_59_3118_0, i_10_59_3211_0, i_10_59_3228_0, i_10_59_3387_0,
    i_10_59_3390_0, i_10_59_3404_0, i_10_59_3408_0, i_10_59_3468_0,
    i_10_59_3525_0, i_10_59_3539_0, i_10_59_3585_0, i_10_59_3598_0,
    i_10_59_3605_0, i_10_59_3772_0, i_10_59_3808_0, i_10_59_3809_0,
    i_10_59_3894_0, i_10_59_3905_0, i_10_59_3918_0, i_10_59_3964_0,
    i_10_59_3967_0, i_10_59_3969_0, i_10_59_3991_0, i_10_59_3994_0,
    i_10_59_4012_0, i_10_59_4013_0, i_10_59_4294_0, i_10_59_4387_0,
    i_10_59_4440_0, i_10_59_4455_0, i_10_59_4535_0, i_10_59_4598_0,
    o_10_59_0_0  );
  input  i_10_59_150_0, i_10_59_180_0, i_10_59_286_0, i_10_59_319_0,
    i_10_59_461_0, i_10_59_588_0, i_10_59_592_0, i_10_59_633_0,
    i_10_59_692_0, i_10_59_735_0, i_10_59_798_0, i_10_59_799_0,
    i_10_59_828_0, i_10_59_831_0, i_10_59_929_0, i_10_59_961_0,
    i_10_59_962_0, i_10_59_1040_0, i_10_59_1041_0, i_10_59_1120_0,
    i_10_59_1167_0, i_10_59_1180_0, i_10_59_1306_0, i_10_59_1344_0,
    i_10_59_1346_0, i_10_59_1365_0, i_10_59_1366_0, i_10_59_1554_0,
    i_10_59_1570_0, i_10_59_1648_0, i_10_59_1744_0, i_10_59_1769_0,
    i_10_59_1771_0, i_10_59_1785_0, i_10_59_1788_0, i_10_59_1791_0,
    i_10_59_2011_0, i_10_59_2012_0, i_10_59_2025_0, i_10_59_2142_0,
    i_10_59_2380_0, i_10_59_2389_0, i_10_59_2437_0, i_10_59_2438_0,
    i_10_59_2452_0, i_10_59_2478_0, i_10_59_2479_0, i_10_59_2480_0,
    i_10_59_2542_0, i_10_59_2636_0, i_10_59_2652_0, i_10_59_2713_0,
    i_10_59_2818_0, i_10_59_2828_0, i_10_59_2831_0, i_10_59_2844_0,
    i_10_59_2848_0, i_10_59_2883_0, i_10_59_2910_0, i_10_59_2911_0,
    i_10_59_2922_0, i_10_59_2923_0, i_10_59_2938_0, i_10_59_2958_0,
    i_10_59_2959_0, i_10_59_2978_0, i_10_59_2986_0, i_10_59_3046_0,
    i_10_59_3118_0, i_10_59_3211_0, i_10_59_3228_0, i_10_59_3387_0,
    i_10_59_3390_0, i_10_59_3404_0, i_10_59_3408_0, i_10_59_3468_0,
    i_10_59_3525_0, i_10_59_3539_0, i_10_59_3585_0, i_10_59_3598_0,
    i_10_59_3605_0, i_10_59_3772_0, i_10_59_3808_0, i_10_59_3809_0,
    i_10_59_3894_0, i_10_59_3905_0, i_10_59_3918_0, i_10_59_3964_0,
    i_10_59_3967_0, i_10_59_3969_0, i_10_59_3991_0, i_10_59_3994_0,
    i_10_59_4012_0, i_10_59_4013_0, i_10_59_4294_0, i_10_59_4387_0,
    i_10_59_4440_0, i_10_59_4455_0, i_10_59_4535_0, i_10_59_4598_0;
  output o_10_59_0_0;
  assign o_10_59_0_0 = 0;
endmodule



// Benchmark "kernel_10_60" written by ABC on Sun Jul 19 10:22:03 2020

module kernel_10_60 ( 
    i_10_60_51_0, i_10_60_246_0, i_10_60_247_0, i_10_60_254_0,
    i_10_60_287_0, i_10_60_290_0, i_10_60_315_0, i_10_60_316_0,
    i_10_60_319_0, i_10_60_320_0, i_10_60_327_0, i_10_60_392_0,
    i_10_60_393_0, i_10_60_467_0, i_10_60_908_0, i_10_60_1055_0,
    i_10_60_1083_0, i_10_60_1160_0, i_10_60_1234_0, i_10_60_1235_0,
    i_10_60_1238_0, i_10_60_1242_0, i_10_60_1245_0, i_10_60_1308_0,
    i_10_60_1362_0, i_10_60_1432_0, i_10_60_1441_0, i_10_60_1444_0,
    i_10_60_1540_0, i_10_60_1551_0, i_10_60_1575_0, i_10_60_1576_0,
    i_10_60_1577_0, i_10_60_1622_0, i_10_60_1655_0, i_10_60_1730_0,
    i_10_60_1800_0, i_10_60_1911_0, i_10_60_1981_0, i_10_60_1982_0,
    i_10_60_2196_0, i_10_60_2197_0, i_10_60_2338_0, i_10_60_2349_0,
    i_10_60_2352_0, i_10_60_2353_0, i_10_60_2354_0, i_10_60_2448_0,
    i_10_60_2457_0, i_10_60_2515_0, i_10_60_2516_0, i_10_60_2563_0,
    i_10_60_2567_0, i_10_60_2608_0, i_10_60_2629_0, i_10_60_2701_0,
    i_10_60_2712_0, i_10_60_2713_0, i_10_60_2731_0, i_10_60_2820_0,
    i_10_60_2827_0, i_10_60_2845_0, i_10_60_2955_0, i_10_60_2961_0,
    i_10_60_2962_0, i_10_60_3042_0, i_10_60_3070_0, i_10_60_3071_0,
    i_10_60_3277_0, i_10_60_3278_0, i_10_60_3353_0, i_10_60_3384_0,
    i_10_60_3470_0, i_10_60_3538_0, i_10_60_3557_0, i_10_60_3584_0,
    i_10_60_3610_0, i_10_60_3611_0, i_10_60_3723_0, i_10_60_3835_0,
    i_10_60_3836_0, i_10_60_3838_0, i_10_60_3857_0, i_10_60_3906_0,
    i_10_60_4030_0, i_10_60_4062_0, i_10_60_4113_0, i_10_60_4114_0,
    i_10_60_4122_0, i_10_60_4123_0, i_10_60_4127_0, i_10_60_4151_0,
    i_10_60_4168_0, i_10_60_4169_0, i_10_60_4191_0, i_10_60_4275_0,
    i_10_60_4278_0, i_10_60_4289_0, i_10_60_4581_0, i_10_60_4582_0,
    o_10_60_0_0  );
  input  i_10_60_51_0, i_10_60_246_0, i_10_60_247_0, i_10_60_254_0,
    i_10_60_287_0, i_10_60_290_0, i_10_60_315_0, i_10_60_316_0,
    i_10_60_319_0, i_10_60_320_0, i_10_60_327_0, i_10_60_392_0,
    i_10_60_393_0, i_10_60_467_0, i_10_60_908_0, i_10_60_1055_0,
    i_10_60_1083_0, i_10_60_1160_0, i_10_60_1234_0, i_10_60_1235_0,
    i_10_60_1238_0, i_10_60_1242_0, i_10_60_1245_0, i_10_60_1308_0,
    i_10_60_1362_0, i_10_60_1432_0, i_10_60_1441_0, i_10_60_1444_0,
    i_10_60_1540_0, i_10_60_1551_0, i_10_60_1575_0, i_10_60_1576_0,
    i_10_60_1577_0, i_10_60_1622_0, i_10_60_1655_0, i_10_60_1730_0,
    i_10_60_1800_0, i_10_60_1911_0, i_10_60_1981_0, i_10_60_1982_0,
    i_10_60_2196_0, i_10_60_2197_0, i_10_60_2338_0, i_10_60_2349_0,
    i_10_60_2352_0, i_10_60_2353_0, i_10_60_2354_0, i_10_60_2448_0,
    i_10_60_2457_0, i_10_60_2515_0, i_10_60_2516_0, i_10_60_2563_0,
    i_10_60_2567_0, i_10_60_2608_0, i_10_60_2629_0, i_10_60_2701_0,
    i_10_60_2712_0, i_10_60_2713_0, i_10_60_2731_0, i_10_60_2820_0,
    i_10_60_2827_0, i_10_60_2845_0, i_10_60_2955_0, i_10_60_2961_0,
    i_10_60_2962_0, i_10_60_3042_0, i_10_60_3070_0, i_10_60_3071_0,
    i_10_60_3277_0, i_10_60_3278_0, i_10_60_3353_0, i_10_60_3384_0,
    i_10_60_3470_0, i_10_60_3538_0, i_10_60_3557_0, i_10_60_3584_0,
    i_10_60_3610_0, i_10_60_3611_0, i_10_60_3723_0, i_10_60_3835_0,
    i_10_60_3836_0, i_10_60_3838_0, i_10_60_3857_0, i_10_60_3906_0,
    i_10_60_4030_0, i_10_60_4062_0, i_10_60_4113_0, i_10_60_4114_0,
    i_10_60_4122_0, i_10_60_4123_0, i_10_60_4127_0, i_10_60_4151_0,
    i_10_60_4168_0, i_10_60_4169_0, i_10_60_4191_0, i_10_60_4275_0,
    i_10_60_4278_0, i_10_60_4289_0, i_10_60_4581_0, i_10_60_4582_0;
  output o_10_60_0_0;
  assign o_10_60_0_0 = 0;
endmodule



// Benchmark "kernel_10_61" written by ABC on Sun Jul 19 10:22:04 2020

module kernel_10_61 ( 
    i_10_61_122_0, i_10_61_148_0, i_10_61_277_0, i_10_61_289_0,
    i_10_61_326_0, i_10_61_370_0, i_10_61_412_0, i_10_61_413_0,
    i_10_61_463_0, i_10_61_505_0, i_10_61_640_0, i_10_61_733_0,
    i_10_61_959_0, i_10_61_1009_0, i_10_61_1019_0, i_10_61_1054_0,
    i_10_61_1055_0, i_10_61_1156_0, i_10_61_1202_0, i_10_61_1243_0,
    i_10_61_1265_0, i_10_61_1287_0, i_10_61_1382_0, i_10_61_1456_0,
    i_10_61_1499_0, i_10_61_1540_0, i_10_61_1547_0, i_10_61_1611_0,
    i_10_61_1615_0, i_10_61_1622_0, i_10_61_1625_0, i_10_61_1648_0,
    i_10_61_1730_0, i_10_61_1747_0, i_10_61_1783_0, i_10_61_1819_0,
    i_10_61_1936_0, i_10_61_2018_0, i_10_61_2027_0, i_10_61_2156_0,
    i_10_61_2197_0, i_10_61_2200_0, i_10_61_2332_0, i_10_61_2336_0,
    i_10_61_2351_0, i_10_61_2359_0, i_10_61_2360_0, i_10_61_2372_0,
    i_10_61_2432_0, i_10_61_2435_0, i_10_61_2455_0, i_10_61_2513_0,
    i_10_61_2525_0, i_10_61_2605_0, i_10_61_2606_0, i_10_61_2630_0,
    i_10_61_2632_0, i_10_61_2824_0, i_10_61_2827_0, i_10_61_2837_0,
    i_10_61_2847_0, i_10_61_2864_0, i_10_61_2920_0, i_10_61_2975_0,
    i_10_61_2993_0, i_10_61_3280_0, i_10_61_3281_0, i_10_61_3298_0,
    i_10_61_3314_0, i_10_61_3317_0, i_10_61_3402_0, i_10_61_3403_0,
    i_10_61_3440_0, i_10_61_3469_0, i_10_61_3540_0, i_10_61_3565_0,
    i_10_61_3613_0, i_10_61_3616_0, i_10_61_3721_0, i_10_61_3800_0,
    i_10_61_3835_0, i_10_61_3836_0, i_10_61_3839_0, i_10_61_3842_0,
    i_10_61_3858_0, i_10_61_3898_0, i_10_61_3944_0, i_10_61_3982_0,
    i_10_61_3998_0, i_10_61_4087_0, i_10_61_4088_0, i_10_61_4130_0,
    i_10_61_4151_0, i_10_61_4156_0, i_10_61_4243_0, i_10_61_4267_0,
    i_10_61_4276_0, i_10_61_4277_0, i_10_61_4367_0, i_10_61_4595_0,
    o_10_61_0_0  );
  input  i_10_61_122_0, i_10_61_148_0, i_10_61_277_0, i_10_61_289_0,
    i_10_61_326_0, i_10_61_370_0, i_10_61_412_0, i_10_61_413_0,
    i_10_61_463_0, i_10_61_505_0, i_10_61_640_0, i_10_61_733_0,
    i_10_61_959_0, i_10_61_1009_0, i_10_61_1019_0, i_10_61_1054_0,
    i_10_61_1055_0, i_10_61_1156_0, i_10_61_1202_0, i_10_61_1243_0,
    i_10_61_1265_0, i_10_61_1287_0, i_10_61_1382_0, i_10_61_1456_0,
    i_10_61_1499_0, i_10_61_1540_0, i_10_61_1547_0, i_10_61_1611_0,
    i_10_61_1615_0, i_10_61_1622_0, i_10_61_1625_0, i_10_61_1648_0,
    i_10_61_1730_0, i_10_61_1747_0, i_10_61_1783_0, i_10_61_1819_0,
    i_10_61_1936_0, i_10_61_2018_0, i_10_61_2027_0, i_10_61_2156_0,
    i_10_61_2197_0, i_10_61_2200_0, i_10_61_2332_0, i_10_61_2336_0,
    i_10_61_2351_0, i_10_61_2359_0, i_10_61_2360_0, i_10_61_2372_0,
    i_10_61_2432_0, i_10_61_2435_0, i_10_61_2455_0, i_10_61_2513_0,
    i_10_61_2525_0, i_10_61_2605_0, i_10_61_2606_0, i_10_61_2630_0,
    i_10_61_2632_0, i_10_61_2824_0, i_10_61_2827_0, i_10_61_2837_0,
    i_10_61_2847_0, i_10_61_2864_0, i_10_61_2920_0, i_10_61_2975_0,
    i_10_61_2993_0, i_10_61_3280_0, i_10_61_3281_0, i_10_61_3298_0,
    i_10_61_3314_0, i_10_61_3317_0, i_10_61_3402_0, i_10_61_3403_0,
    i_10_61_3440_0, i_10_61_3469_0, i_10_61_3540_0, i_10_61_3565_0,
    i_10_61_3613_0, i_10_61_3616_0, i_10_61_3721_0, i_10_61_3800_0,
    i_10_61_3835_0, i_10_61_3836_0, i_10_61_3839_0, i_10_61_3842_0,
    i_10_61_3858_0, i_10_61_3898_0, i_10_61_3944_0, i_10_61_3982_0,
    i_10_61_3998_0, i_10_61_4087_0, i_10_61_4088_0, i_10_61_4130_0,
    i_10_61_4151_0, i_10_61_4156_0, i_10_61_4243_0, i_10_61_4267_0,
    i_10_61_4276_0, i_10_61_4277_0, i_10_61_4367_0, i_10_61_4595_0;
  output o_10_61_0_0;
  assign o_10_61_0_0 = 0;
endmodule



// Benchmark "kernel_10_62" written by ABC on Sun Jul 19 10:22:05 2020

module kernel_10_62 ( 
    i_10_62_221_0, i_10_62_243_0, i_10_62_244_0, i_10_62_250_0,
    i_10_62_281_0, i_10_62_283_0, i_10_62_286_0, i_10_62_322_0,
    i_10_62_323_0, i_10_62_439_0, i_10_62_467_0, i_10_62_755_0,
    i_10_62_796_0, i_10_62_799_0, i_10_62_800_0, i_10_62_904_0,
    i_10_62_991_0, i_10_62_992_0, i_10_62_1033_0, i_10_62_1034_0,
    i_10_62_1233_0, i_10_62_1237_0, i_10_62_1238_0, i_10_62_1240_0,
    i_10_62_1241_0, i_10_62_1300_0, i_10_62_1309_0, i_10_62_1432_0,
    i_10_62_1437_0, i_10_62_1438_0, i_10_62_1578_0, i_10_62_1579_0,
    i_10_62_1583_0, i_10_62_1651_0, i_10_62_1653_0, i_10_62_1655_0,
    i_10_62_1686_0, i_10_62_1816_0, i_10_62_1817_0, i_10_62_1823_0,
    i_10_62_1912_0, i_10_62_1913_0, i_10_62_2185_0, i_10_62_2306_0,
    i_10_62_2351_0, i_10_62_2362_0, i_10_62_2363_0, i_10_62_2448_0,
    i_10_62_2473_0, i_10_62_2608_0, i_10_62_2631_0, i_10_62_2662_0,
    i_10_62_2705_0, i_10_62_2719_0, i_10_62_2728_0, i_10_62_2734_0,
    i_10_62_2735_0, i_10_62_2785_0, i_10_62_2786_0, i_10_62_2828_0,
    i_10_62_2833_0, i_10_62_2834_0, i_10_62_2888_0, i_10_62_2924_0,
    i_10_62_2986_0, i_10_62_3154_0, i_10_62_3163_0, i_10_62_3196_0,
    i_10_62_3197_0, i_10_62_3322_0, i_10_62_3388_0, i_10_62_3406_0,
    i_10_62_3407_0, i_10_62_3588_0, i_10_62_3589_0, i_10_62_3590_0,
    i_10_62_3613_0, i_10_62_3616_0, i_10_62_3617_0, i_10_62_3646_0,
    i_10_62_3652_0, i_10_62_3682_0, i_10_62_3838_0, i_10_62_3839_0,
    i_10_62_3840_0, i_10_62_3841_0, i_10_62_3856_0, i_10_62_3983_0,
    i_10_62_3984_0, i_10_62_3991_0, i_10_62_3992_0, i_10_62_4028_0,
    i_10_62_4117_0, i_10_62_4118_0, i_10_62_4120_0, i_10_62_4130_0,
    i_10_62_4270_0, i_10_62_4271_0, i_10_62_4290_0, i_10_62_4567_0,
    o_10_62_0_0  );
  input  i_10_62_221_0, i_10_62_243_0, i_10_62_244_0, i_10_62_250_0,
    i_10_62_281_0, i_10_62_283_0, i_10_62_286_0, i_10_62_322_0,
    i_10_62_323_0, i_10_62_439_0, i_10_62_467_0, i_10_62_755_0,
    i_10_62_796_0, i_10_62_799_0, i_10_62_800_0, i_10_62_904_0,
    i_10_62_991_0, i_10_62_992_0, i_10_62_1033_0, i_10_62_1034_0,
    i_10_62_1233_0, i_10_62_1237_0, i_10_62_1238_0, i_10_62_1240_0,
    i_10_62_1241_0, i_10_62_1300_0, i_10_62_1309_0, i_10_62_1432_0,
    i_10_62_1437_0, i_10_62_1438_0, i_10_62_1578_0, i_10_62_1579_0,
    i_10_62_1583_0, i_10_62_1651_0, i_10_62_1653_0, i_10_62_1655_0,
    i_10_62_1686_0, i_10_62_1816_0, i_10_62_1817_0, i_10_62_1823_0,
    i_10_62_1912_0, i_10_62_1913_0, i_10_62_2185_0, i_10_62_2306_0,
    i_10_62_2351_0, i_10_62_2362_0, i_10_62_2363_0, i_10_62_2448_0,
    i_10_62_2473_0, i_10_62_2608_0, i_10_62_2631_0, i_10_62_2662_0,
    i_10_62_2705_0, i_10_62_2719_0, i_10_62_2728_0, i_10_62_2734_0,
    i_10_62_2735_0, i_10_62_2785_0, i_10_62_2786_0, i_10_62_2828_0,
    i_10_62_2833_0, i_10_62_2834_0, i_10_62_2888_0, i_10_62_2924_0,
    i_10_62_2986_0, i_10_62_3154_0, i_10_62_3163_0, i_10_62_3196_0,
    i_10_62_3197_0, i_10_62_3322_0, i_10_62_3388_0, i_10_62_3406_0,
    i_10_62_3407_0, i_10_62_3588_0, i_10_62_3589_0, i_10_62_3590_0,
    i_10_62_3613_0, i_10_62_3616_0, i_10_62_3617_0, i_10_62_3646_0,
    i_10_62_3652_0, i_10_62_3682_0, i_10_62_3838_0, i_10_62_3839_0,
    i_10_62_3840_0, i_10_62_3841_0, i_10_62_3856_0, i_10_62_3983_0,
    i_10_62_3984_0, i_10_62_3991_0, i_10_62_3992_0, i_10_62_4028_0,
    i_10_62_4117_0, i_10_62_4118_0, i_10_62_4120_0, i_10_62_4130_0,
    i_10_62_4270_0, i_10_62_4271_0, i_10_62_4290_0, i_10_62_4567_0;
  output o_10_62_0_0;
  assign o_10_62_0_0 = ~((~i_10_62_992_0 & ((~i_10_62_244_0 & ((~i_10_62_323_0 & ~i_10_62_1033_0 & ~i_10_62_3197_0) | (~i_10_62_439_0 & ~i_10_62_2306_0 & ~i_10_62_2734_0 & ~i_10_62_2785_0 & ~i_10_62_3682_0 & ~i_10_62_3991_0))) | (~i_10_62_439_0 & ~i_10_62_2363_0 & ~i_10_62_3163_0 & ~i_10_62_3646_0 & ~i_10_62_3991_0))) | (i_10_62_800_0 & (i_10_62_4290_0 | (~i_10_62_221_0 & ~i_10_62_1583_0 & ~i_10_62_2828_0 & i_10_62_2924_0 & ~i_10_62_3838_0))) | (~i_10_62_991_0 & ((~i_10_62_1309_0 & i_10_62_1655_0 & ~i_10_62_2833_0 & ~i_10_62_2986_0 & ~i_10_62_3163_0) | (~i_10_62_322_0 & ~i_10_62_2185_0 & ~i_10_62_3407_0 & ~i_10_62_3839_0 & ~i_10_62_3992_0 & ~i_10_62_4567_0))) | (~i_10_62_1034_0 & ((~i_10_62_755_0 & ~i_10_62_904_0 & ~i_10_62_1817_0 & i_10_62_2631_0 & i_10_62_2834_0) | (~i_10_62_1309_0 & ~i_10_62_1579_0 & ~i_10_62_2306_0 & ~i_10_62_2735_0 & ~i_10_62_3992_0))) | (~i_10_62_1816_0 & ((~i_10_62_250_0 & ~i_10_62_2363_0 & ~i_10_62_2735_0 & ~i_10_62_2924_0 & ~i_10_62_3197_0 & ~i_10_62_3682_0) | (~i_10_62_243_0 & ~i_10_62_2306_0 & ~i_10_62_3406_0 & ~i_10_62_3992_0))) | (~i_10_62_1823_0 & ((i_10_62_1655_0 & ~i_10_62_1817_0 & ~i_10_62_2631_0 & ~i_10_62_3196_0) | (~i_10_62_1583_0 & ~i_10_62_2608_0 & ~i_10_62_2662_0 & ~i_10_62_3682_0))) | (~i_10_62_2735_0 & ~i_10_62_4120_0 & ((i_10_62_796_0 & ~i_10_62_1578_0 & i_10_62_2924_0) | (~i_10_62_796_0 & ~i_10_62_3407_0 & i_10_62_3646_0 & ~i_10_62_3682_0 & ~i_10_62_3984_0))) | (i_10_62_2924_0 & ((~i_10_62_439_0 & ~i_10_62_1432_0 & i_10_62_2631_0 & ~i_10_62_3163_0) | (i_10_62_3840_0 & ~i_10_62_4117_0))) | (~i_10_62_3196_0 & ((i_10_62_2828_0 & ~i_10_62_3613_0 & ~i_10_62_3992_0) | (i_10_62_1686_0 & ~i_10_62_2363_0 & ~i_10_62_3991_0 & i_10_62_4028_0))) | (~i_10_62_3991_0 & ((~i_10_62_2362_0 & i_10_62_3617_0 & ~i_10_62_3839_0) | (~i_10_62_3388_0 & ~i_10_62_3406_0 & i_10_62_3652_0 & ~i_10_62_4130_0))) | (i_10_62_1913_0 & i_10_62_2728_0) | (~i_10_62_3838_0 & i_10_62_4270_0));
endmodule



// Benchmark "kernel_10_63" written by ABC on Sun Jul 19 10:22:06 2020

module kernel_10_63 ( 
    i_10_63_174_0, i_10_63_216_0, i_10_63_220_0, i_10_63_246_0,
    i_10_63_292_0, i_10_63_293_0, i_10_63_328_0, i_10_63_329_0,
    i_10_63_410_0, i_10_63_443_0, i_10_63_445_0, i_10_63_465_0,
    i_10_63_645_0, i_10_63_897_0, i_10_63_898_0, i_10_63_899_0,
    i_10_63_1168_0, i_10_63_1239_0, i_10_63_1240_0, i_10_63_1308_0,
    i_10_63_1362_0, i_10_63_1366_0, i_10_63_1444_0, i_10_63_1579_0,
    i_10_63_1648_0, i_10_63_1650_0, i_10_63_1654_0, i_10_63_1675_0,
    i_10_63_1684_0, i_10_63_1685_0, i_10_63_1825_0, i_10_63_1915_0,
    i_10_63_1952_0, i_10_63_1995_0, i_10_63_1996_0, i_10_63_2337_0,
    i_10_63_2350_0, i_10_63_2352_0, i_10_63_2364_0, i_10_63_2365_0,
    i_10_63_2382_0, i_10_63_2383_0, i_10_63_2408_0, i_10_63_2411_0,
    i_10_63_2451_0, i_10_63_2470_0, i_10_63_2481_0, i_10_63_2572_0,
    i_10_63_2631_0, i_10_63_2632_0, i_10_63_2656_0, i_10_63_2658_0,
    i_10_63_2661_0, i_10_63_2706_0, i_10_63_2707_0, i_10_63_2716_0,
    i_10_63_2721_0, i_10_63_2731_0, i_10_63_2734_0, i_10_63_2821_0,
    i_10_63_2824_0, i_10_63_2831_0, i_10_63_2884_0, i_10_63_2919_0,
    i_10_63_2920_0, i_10_63_2923_0, i_10_63_3034_0, i_10_63_3035_0,
    i_10_63_3036_0, i_10_63_3153_0, i_10_63_3196_0, i_10_63_3199_0,
    i_10_63_3202_0, i_10_63_3270_0, i_10_63_3273_0, i_10_63_3279_0,
    i_10_63_3282_0, i_10_63_3283_0, i_10_63_3388_0, i_10_63_3404_0,
    i_10_63_3433_0, i_10_63_3469_0, i_10_63_3472_0, i_10_63_3519_0,
    i_10_63_3522_0, i_10_63_3647_0, i_10_63_3648_0, i_10_63_3651_0,
    i_10_63_3653_0, i_10_63_3783_0, i_10_63_3785_0, i_10_63_3835_0,
    i_10_63_3847_0, i_10_63_3848_0, i_10_63_3985_0, i_10_63_4116_0,
    i_10_63_4119_0, i_10_63_4120_0, i_10_63_4283_0, i_10_63_4291_0,
    o_10_63_0_0  );
  input  i_10_63_174_0, i_10_63_216_0, i_10_63_220_0, i_10_63_246_0,
    i_10_63_292_0, i_10_63_293_0, i_10_63_328_0, i_10_63_329_0,
    i_10_63_410_0, i_10_63_443_0, i_10_63_445_0, i_10_63_465_0,
    i_10_63_645_0, i_10_63_897_0, i_10_63_898_0, i_10_63_899_0,
    i_10_63_1168_0, i_10_63_1239_0, i_10_63_1240_0, i_10_63_1308_0,
    i_10_63_1362_0, i_10_63_1366_0, i_10_63_1444_0, i_10_63_1579_0,
    i_10_63_1648_0, i_10_63_1650_0, i_10_63_1654_0, i_10_63_1675_0,
    i_10_63_1684_0, i_10_63_1685_0, i_10_63_1825_0, i_10_63_1915_0,
    i_10_63_1952_0, i_10_63_1995_0, i_10_63_1996_0, i_10_63_2337_0,
    i_10_63_2350_0, i_10_63_2352_0, i_10_63_2364_0, i_10_63_2365_0,
    i_10_63_2382_0, i_10_63_2383_0, i_10_63_2408_0, i_10_63_2411_0,
    i_10_63_2451_0, i_10_63_2470_0, i_10_63_2481_0, i_10_63_2572_0,
    i_10_63_2631_0, i_10_63_2632_0, i_10_63_2656_0, i_10_63_2658_0,
    i_10_63_2661_0, i_10_63_2706_0, i_10_63_2707_0, i_10_63_2716_0,
    i_10_63_2721_0, i_10_63_2731_0, i_10_63_2734_0, i_10_63_2821_0,
    i_10_63_2824_0, i_10_63_2831_0, i_10_63_2884_0, i_10_63_2919_0,
    i_10_63_2920_0, i_10_63_2923_0, i_10_63_3034_0, i_10_63_3035_0,
    i_10_63_3036_0, i_10_63_3153_0, i_10_63_3196_0, i_10_63_3199_0,
    i_10_63_3202_0, i_10_63_3270_0, i_10_63_3273_0, i_10_63_3279_0,
    i_10_63_3282_0, i_10_63_3283_0, i_10_63_3388_0, i_10_63_3404_0,
    i_10_63_3433_0, i_10_63_3469_0, i_10_63_3472_0, i_10_63_3519_0,
    i_10_63_3522_0, i_10_63_3647_0, i_10_63_3648_0, i_10_63_3651_0,
    i_10_63_3653_0, i_10_63_3783_0, i_10_63_3785_0, i_10_63_3835_0,
    i_10_63_3847_0, i_10_63_3848_0, i_10_63_3985_0, i_10_63_4116_0,
    i_10_63_4119_0, i_10_63_4120_0, i_10_63_4283_0, i_10_63_4291_0;
  output o_10_63_0_0;
  assign o_10_63_0_0 = ~((~i_10_63_3835_0 & ((~i_10_63_246_0 & ((~i_10_63_292_0 & ~i_10_63_293_0 & ~i_10_63_898_0 & ~i_10_63_2408_0 & ~i_10_63_2656_0 & i_10_63_3847_0) | (~i_10_63_443_0 & i_10_63_2631_0 & ~i_10_63_3036_0 & ~i_10_63_3270_0 & ~i_10_63_3522_0 & ~i_10_63_3785_0 & ~i_10_63_3848_0))) | (~i_10_63_899_0 & ~i_10_63_1650_0 & ~i_10_63_2658_0 & ~i_10_63_2707_0 & ~i_10_63_2923_0 & ~i_10_63_3647_0) | (~i_10_63_1444_0 & ~i_10_63_2408_0 & ~i_10_63_2631_0 & ~i_10_63_2632_0 & ~i_10_63_2721_0 & i_10_63_2919_0 & ~i_10_63_3270_0 & i_10_63_3785_0))) | (~i_10_63_216_0 & ((~i_10_63_220_0 & ((~i_10_63_1444_0 & ~i_10_63_2631_0 & i_10_63_3847_0) | (~i_10_63_2451_0 & ~i_10_63_2721_0 & i_10_63_3848_0))) | (~i_10_63_293_0 & ((~i_10_63_328_0 & ~i_10_63_1650_0 & ~i_10_63_1996_0 & ~i_10_63_2383_0 & ~i_10_63_3519_0) | (~i_10_63_329_0 & ~i_10_63_2352_0 & ~i_10_63_2364_0 & ~i_10_63_2411_0 & ~i_10_63_2572_0 & ~i_10_63_2631_0 & ~i_10_63_2658_0 & ~i_10_63_3270_0 & ~i_10_63_3785_0 & ~i_10_63_3847_0))) | (~i_10_63_445_0 & ((~i_10_63_292_0 & ~i_10_63_328_0 & ~i_10_63_1996_0 & ~i_10_63_2631_0 & ~i_10_63_2632_0 & ~i_10_63_3522_0) | (~i_10_63_1995_0 & ~i_10_63_2364_0 & ~i_10_63_2365_0 & ~i_10_63_3647_0 & ~i_10_63_3648_0 & ~i_10_63_4116_0))) | (i_10_63_2632_0 & ((~i_10_63_329_0 & ~i_10_63_898_0 & ~i_10_63_1684_0 & ~i_10_63_2337_0 & ~i_10_63_2350_0) | (i_10_63_1579_0 & ~i_10_63_2408_0 & ~i_10_63_3035_0 & ~i_10_63_3847_0))))) | (~i_10_63_329_0 & ((i_10_63_1952_0 & ~i_10_63_2707_0 & ~i_10_63_2923_0) | (~i_10_63_898_0 & ~i_10_63_1444_0 & ~i_10_63_1648_0 & ~i_10_63_1996_0 & ~i_10_63_2337_0 & ~i_10_63_2451_0 & ~i_10_63_3196_0 & ~i_10_63_3270_0 & ~i_10_63_3433_0 & ~i_10_63_3985_0))) | (~i_10_63_1579_0 & ((~i_10_63_443_0 & i_10_63_2632_0 & i_10_63_2920_0 & ~i_10_63_2923_0 & ~i_10_63_3270_0 & ~i_10_63_3519_0) | (~i_10_63_174_0 & i_10_63_1648_0 & i_10_63_1650_0 & ~i_10_63_1684_0 & ~i_10_63_2350_0 & ~i_10_63_3279_0 & ~i_10_63_3647_0))) | (~i_10_63_174_0 & ((~i_10_63_2352_0 & ~i_10_63_2451_0 & ~i_10_63_2656_0 & i_10_63_4116_0) | (~i_10_63_443_0 & ~i_10_63_2365_0 & ~i_10_63_3522_0 & i_10_63_4120_0))) | (i_10_63_1654_0 & i_10_63_4116_0 & ((~i_10_63_1444_0 & ~i_10_63_2656_0) | (~i_10_63_292_0 & ~i_10_63_293_0 & ~i_10_63_2408_0 & ~i_10_63_2919_0 & ~i_10_63_3199_0))) | (~i_10_63_292_0 & ((~i_10_63_443_0 & ~i_10_63_1444_0 & ~i_10_63_1996_0 & i_10_63_2658_0 & i_10_63_2661_0 & ~i_10_63_3270_0) | (~i_10_63_410_0 & ~i_10_63_1684_0 & i_10_63_1825_0 & ~i_10_63_2408_0 & ~i_10_63_2481_0 & ~i_10_63_2734_0 & ~i_10_63_3273_0))) | (~i_10_63_2364_0 & ((~i_10_63_293_0 & ~i_10_63_3273_0 & ((~i_10_63_1366_0 & ~i_10_63_2350_0 & ~i_10_63_2383_0 & ~i_10_63_2656_0 & ~i_10_63_2919_0 & ~i_10_63_3199_0) | (~i_10_63_220_0 & ~i_10_63_899_0 & ~i_10_63_1685_0 & ~i_10_63_3270_0 & ~i_10_63_3519_0 & ~i_10_63_1952_0 & ~i_10_63_2408_0))) | (~i_10_63_645_0 & ~i_10_63_1444_0 & i_10_63_1825_0 & ~i_10_63_2352_0 & ~i_10_63_2716_0 & i_10_63_2923_0))) | (~i_10_63_2706_0 & ((~i_10_63_1685_0 & ~i_10_63_2656_0 & i_10_63_3647_0) | (~i_10_63_3388_0 & ~i_10_63_3519_0 & i_10_63_4119_0 & i_10_63_4120_0))) | (~i_10_63_3270_0 & ((i_10_63_1825_0 & i_10_63_3196_0) | (i_10_63_3036_0 & ~i_10_63_3647_0))) | (~i_10_63_4120_0 & ((~i_10_63_2631_0 & i_10_63_3648_0 & i_10_63_3835_0 & ~i_10_63_3847_0) | (~i_10_63_2383_0 & ~i_10_63_2661_0 & i_10_63_4291_0))) | (~i_10_63_2352_0 & i_10_63_2408_0 & ~i_10_63_2481_0 & i_10_63_2631_0 & ~i_10_63_2923_0) | (i_10_63_1579_0 & i_10_63_2821_0 & ~i_10_63_3519_0) | (i_10_63_2884_0 & i_10_63_3647_0) | (~i_10_63_2337_0 & i_10_63_3034_0 & ~i_10_63_3785_0));
endmodule



// Benchmark "kernel_10_64" written by ABC on Sun Jul 19 10:22:07 2020

module kernel_10_64 ( 
    i_10_64_34_0, i_10_64_65_0, i_10_64_172_0, i_10_64_224_0,
    i_10_64_281_0, i_10_64_284_0, i_10_64_330_0, i_10_64_331_0,
    i_10_64_442_0, i_10_64_448_0, i_10_64_541_0, i_10_64_542_0,
    i_10_64_544_0, i_10_64_545_0, i_10_64_596_0, i_10_64_712_0,
    i_10_64_713_0, i_10_64_715_0, i_10_64_736_0, i_10_64_794_0,
    i_10_64_797_0, i_10_64_955_0, i_10_64_956_0, i_10_64_990_0,
    i_10_64_1084_0, i_10_64_1241_0, i_10_64_1247_0, i_10_64_1249_0,
    i_10_64_1309_0, i_10_64_1514_0, i_10_64_1561_0, i_10_64_1562_0,
    i_10_64_1578_0, i_10_64_1579_0, i_10_64_1580_0, i_10_64_1615_0,
    i_10_64_1616_0, i_10_64_1650_0, i_10_64_1687_0, i_10_64_1691_0,
    i_10_64_1765_0, i_10_64_1819_0, i_10_64_1821_0, i_10_64_1824_0,
    i_10_64_1825_0, i_10_64_1954_0, i_10_64_2156_0, i_10_64_2164_0,
    i_10_64_2355_0, i_10_64_2361_0, i_10_64_2362_0, i_10_64_2364_0,
    i_10_64_2365_0, i_10_64_2432_0, i_10_64_2435_0, i_10_64_2470_0,
    i_10_64_2603_0, i_10_64_2634_0, i_10_64_2662_0, i_10_64_2728_0,
    i_10_64_2729_0, i_10_64_2817_0, i_10_64_2820_0, i_10_64_2867_0,
    i_10_64_2979_0, i_10_64_2982_0, i_10_64_3076_0, i_10_64_3077_0,
    i_10_64_3116_0, i_10_64_3232_0, i_10_64_3233_0, i_10_64_3235_0,
    i_10_64_3239_0, i_10_64_3316_0, i_10_64_3385_0, i_10_64_3386_0,
    i_10_64_3407_0, i_10_64_3410_0, i_10_64_3431_0, i_10_64_3590_0,
    i_10_64_3611_0, i_10_64_3683_0, i_10_64_3728_0, i_10_64_3808_0,
    i_10_64_3844_0, i_10_64_3845_0, i_10_64_3906_0, i_10_64_3907_0,
    i_10_64_3994_0, i_10_64_4008_0, i_10_64_4064_0, i_10_64_4100_0,
    i_10_64_4117_0, i_10_64_4217_0, i_10_64_4220_0, i_10_64_4267_0,
    i_10_64_4289_0, i_10_64_4292_0, i_10_64_4475_0, i_10_64_4564_0,
    o_10_64_0_0  );
  input  i_10_64_34_0, i_10_64_65_0, i_10_64_172_0, i_10_64_224_0,
    i_10_64_281_0, i_10_64_284_0, i_10_64_330_0, i_10_64_331_0,
    i_10_64_442_0, i_10_64_448_0, i_10_64_541_0, i_10_64_542_0,
    i_10_64_544_0, i_10_64_545_0, i_10_64_596_0, i_10_64_712_0,
    i_10_64_713_0, i_10_64_715_0, i_10_64_736_0, i_10_64_794_0,
    i_10_64_797_0, i_10_64_955_0, i_10_64_956_0, i_10_64_990_0,
    i_10_64_1084_0, i_10_64_1241_0, i_10_64_1247_0, i_10_64_1249_0,
    i_10_64_1309_0, i_10_64_1514_0, i_10_64_1561_0, i_10_64_1562_0,
    i_10_64_1578_0, i_10_64_1579_0, i_10_64_1580_0, i_10_64_1615_0,
    i_10_64_1616_0, i_10_64_1650_0, i_10_64_1687_0, i_10_64_1691_0,
    i_10_64_1765_0, i_10_64_1819_0, i_10_64_1821_0, i_10_64_1824_0,
    i_10_64_1825_0, i_10_64_1954_0, i_10_64_2156_0, i_10_64_2164_0,
    i_10_64_2355_0, i_10_64_2361_0, i_10_64_2362_0, i_10_64_2364_0,
    i_10_64_2365_0, i_10_64_2432_0, i_10_64_2435_0, i_10_64_2470_0,
    i_10_64_2603_0, i_10_64_2634_0, i_10_64_2662_0, i_10_64_2728_0,
    i_10_64_2729_0, i_10_64_2817_0, i_10_64_2820_0, i_10_64_2867_0,
    i_10_64_2979_0, i_10_64_2982_0, i_10_64_3076_0, i_10_64_3077_0,
    i_10_64_3116_0, i_10_64_3232_0, i_10_64_3233_0, i_10_64_3235_0,
    i_10_64_3239_0, i_10_64_3316_0, i_10_64_3385_0, i_10_64_3386_0,
    i_10_64_3407_0, i_10_64_3410_0, i_10_64_3431_0, i_10_64_3590_0,
    i_10_64_3611_0, i_10_64_3683_0, i_10_64_3728_0, i_10_64_3808_0,
    i_10_64_3844_0, i_10_64_3845_0, i_10_64_3906_0, i_10_64_3907_0,
    i_10_64_3994_0, i_10_64_4008_0, i_10_64_4064_0, i_10_64_4100_0,
    i_10_64_4117_0, i_10_64_4217_0, i_10_64_4220_0, i_10_64_4267_0,
    i_10_64_4289_0, i_10_64_4292_0, i_10_64_4475_0, i_10_64_4564_0;
  output o_10_64_0_0;
  assign o_10_64_0_0 = 0;
endmodule



// Benchmark "kernel_10_65" written by ABC on Sun Jul 19 10:22:09 2020

module kernel_10_65 ( 
    i_10_65_29_0, i_10_65_49_0, i_10_65_50_0, i_10_65_171_0, i_10_65_224_0,
    i_10_65_263_0, i_10_65_277_0, i_10_65_316_0, i_10_65_317_0,
    i_10_65_319_0, i_10_65_320_0, i_10_65_322_0, i_10_65_326_0,
    i_10_65_346_0, i_10_65_362_0, i_10_65_388_0, i_10_65_433_0,
    i_10_65_434_0, i_10_65_437_0, i_10_65_440_0, i_10_65_441_0,
    i_10_65_442_0, i_10_65_448_0, i_10_65_715_0, i_10_65_716_0,
    i_10_65_800_0, i_10_65_947_0, i_10_65_991_0, i_10_65_992_0,
    i_10_65_1001_0, i_10_65_1004_0, i_10_65_1046_0, i_10_65_1084_0,
    i_10_65_1085_0, i_10_65_1135_0, i_10_65_1136_0, i_10_65_1163_0,
    i_10_65_1217_0, i_10_65_1220_0, i_10_65_1238_0, i_10_65_1239_0,
    i_10_65_1306_0, i_10_65_1307_0, i_10_65_1342_0, i_10_65_1346_0,
    i_10_65_1379_0, i_10_65_1432_0, i_10_65_1544_0, i_10_65_1547_0,
    i_10_65_1613_0, i_10_65_1652_0, i_10_65_1653_0, i_10_65_1823_0,
    i_10_65_2000_0, i_10_65_2201_0, i_10_65_2203_0, i_10_65_2204_0,
    i_10_65_2351_0, i_10_65_2354_0, i_10_65_2357_0, i_10_65_2360_0,
    i_10_65_2362_0, i_10_65_2380_0, i_10_65_2450_0, i_10_65_2630_0,
    i_10_65_2675_0, i_10_65_2711_0, i_10_65_2713_0, i_10_65_2720_0,
    i_10_65_2723_0, i_10_65_2724_0, i_10_65_2783_0, i_10_65_2818_0,
    i_10_65_2819_0, i_10_65_2822_0, i_10_65_2832_0, i_10_65_2882_0,
    i_10_65_2884_0, i_10_65_2918_0, i_10_65_2921_0, i_10_65_2980_0,
    i_10_65_2983_0, i_10_65_3092_0, i_10_65_3152_0, i_10_65_3156_0,
    i_10_65_3202_0, i_10_65_3203_0, i_10_65_3278_0, i_10_65_3281_0,
    i_10_65_3584_0, i_10_65_3586_0, i_10_65_3615_0, i_10_65_3835_0,
    i_10_65_3838_0, i_10_65_3841_0, i_10_65_3893_0, i_10_65_3980_0,
    i_10_65_3983_0, i_10_65_4280_0, i_10_65_4283_0,
    o_10_65_0_0  );
  input  i_10_65_29_0, i_10_65_49_0, i_10_65_50_0, i_10_65_171_0,
    i_10_65_224_0, i_10_65_263_0, i_10_65_277_0, i_10_65_316_0,
    i_10_65_317_0, i_10_65_319_0, i_10_65_320_0, i_10_65_322_0,
    i_10_65_326_0, i_10_65_346_0, i_10_65_362_0, i_10_65_388_0,
    i_10_65_433_0, i_10_65_434_0, i_10_65_437_0, i_10_65_440_0,
    i_10_65_441_0, i_10_65_442_0, i_10_65_448_0, i_10_65_715_0,
    i_10_65_716_0, i_10_65_800_0, i_10_65_947_0, i_10_65_991_0,
    i_10_65_992_0, i_10_65_1001_0, i_10_65_1004_0, i_10_65_1046_0,
    i_10_65_1084_0, i_10_65_1085_0, i_10_65_1135_0, i_10_65_1136_0,
    i_10_65_1163_0, i_10_65_1217_0, i_10_65_1220_0, i_10_65_1238_0,
    i_10_65_1239_0, i_10_65_1306_0, i_10_65_1307_0, i_10_65_1342_0,
    i_10_65_1346_0, i_10_65_1379_0, i_10_65_1432_0, i_10_65_1544_0,
    i_10_65_1547_0, i_10_65_1613_0, i_10_65_1652_0, i_10_65_1653_0,
    i_10_65_1823_0, i_10_65_2000_0, i_10_65_2201_0, i_10_65_2203_0,
    i_10_65_2204_0, i_10_65_2351_0, i_10_65_2354_0, i_10_65_2357_0,
    i_10_65_2360_0, i_10_65_2362_0, i_10_65_2380_0, i_10_65_2450_0,
    i_10_65_2630_0, i_10_65_2675_0, i_10_65_2711_0, i_10_65_2713_0,
    i_10_65_2720_0, i_10_65_2723_0, i_10_65_2724_0, i_10_65_2783_0,
    i_10_65_2818_0, i_10_65_2819_0, i_10_65_2822_0, i_10_65_2832_0,
    i_10_65_2882_0, i_10_65_2884_0, i_10_65_2918_0, i_10_65_2921_0,
    i_10_65_2980_0, i_10_65_2983_0, i_10_65_3092_0, i_10_65_3152_0,
    i_10_65_3156_0, i_10_65_3202_0, i_10_65_3203_0, i_10_65_3278_0,
    i_10_65_3281_0, i_10_65_3584_0, i_10_65_3586_0, i_10_65_3615_0,
    i_10_65_3835_0, i_10_65_3838_0, i_10_65_3841_0, i_10_65_3893_0,
    i_10_65_3980_0, i_10_65_3983_0, i_10_65_4280_0, i_10_65_4283_0;
  output o_10_65_0_0;
  assign o_10_65_0_0 = ~((~i_10_65_316_0 & ((~i_10_65_29_0 & ~i_10_65_317_0 & ~i_10_65_434_0 & ~i_10_65_800_0 & ~i_10_65_2819_0 & i_10_65_2921_0) | (~i_10_65_1004_0 & ~i_10_65_1544_0 & ~i_10_65_2675_0 & i_10_65_3586_0 & ~i_10_65_3835_0 & ~i_10_65_3980_0 & ~i_10_65_3983_0))) | (~i_10_65_322_0 & ((~i_10_65_263_0 & ~i_10_65_317_0 & ~i_10_65_388_0 & ~i_10_65_716_0 & ~i_10_65_1084_0 & ~i_10_65_1544_0 & ~i_10_65_3278_0 & ~i_10_65_3980_0) | (i_10_65_992_0 & ~i_10_65_2351_0 & i_10_65_3584_0 & i_10_65_3983_0))) | (~i_10_65_263_0 & ((i_10_65_224_0 & ~i_10_65_320_0 & ~i_10_65_1307_0 & ~i_10_65_3983_0) | (~i_10_65_1085_0 & ~i_10_65_2204_0 & ~i_10_65_2354_0 & ~i_10_65_2724_0 & ~i_10_65_2783_0 & ~i_10_65_2818_0 & ~i_10_65_2819_0 & ~i_10_65_3203_0 & ~i_10_65_4280_0))) | (~i_10_65_2819_0 & ((~i_10_65_29_0 & ((~i_10_65_991_0 & ~i_10_65_1001_0 & ~i_10_65_1547_0 & ~i_10_65_2203_0 & ~i_10_65_2380_0 & ~i_10_65_2713_0 & ~i_10_65_2882_0 & ~i_10_65_3980_0) | (~i_10_65_224_0 & ~i_10_65_320_0 & ~i_10_65_433_0 & ~i_10_65_440_0 & i_10_65_1306_0 & ~i_10_65_2822_0 & ~i_10_65_4283_0))) | (~i_10_65_991_0 & ((~i_10_65_320_0 & ~i_10_65_388_0 & ~i_10_65_2000_0 & ~i_10_65_2450_0 & ~i_10_65_2783_0 & ~i_10_65_3584_0 & ~i_10_65_3893_0) | (~i_10_65_319_0 & ~i_10_65_434_0 & ~i_10_65_1001_0 & ~i_10_65_2675_0 & ~i_10_65_2980_0 & ~i_10_65_3841_0 & ~i_10_65_3980_0 & ~i_10_65_4283_0))))) | (~i_10_65_433_0 & ~i_10_65_2882_0 & ((~i_10_65_992_0 & ~i_10_65_1004_0 & ~i_10_65_1544_0 & ~i_10_65_1613_0 & ~i_10_65_2201_0 & ~i_10_65_2362_0 & ~i_10_65_2818_0 & ~i_10_65_3092_0 & ~i_10_65_4280_0) | (~i_10_65_1085_0 & ~i_10_65_1823_0 & ~i_10_65_2723_0 & ~i_10_65_3203_0 & ~i_10_65_3586_0 & ~i_10_65_3838_0 & ~i_10_65_4283_0))) | (~i_10_65_434_0 & ~i_10_65_3838_0 & ((~i_10_65_317_0 & ~i_10_65_326_0 & ~i_10_65_1004_0 & ~i_10_65_1547_0 & ~i_10_65_2783_0 & ~i_10_65_2822_0) | (~i_10_65_2354_0 & ~i_10_65_2357_0 & ~i_10_65_3584_0 & ~i_10_65_3983_0))) | (~i_10_65_317_0 & ((~i_10_65_1306_0 & ~i_10_65_1823_0 & ~i_10_65_2000_0 & ~i_10_65_2201_0 & ~i_10_65_2822_0 & ~i_10_65_3980_0) | (~i_10_65_1307_0 & ~i_10_65_1346_0 & ~i_10_65_2357_0 & ~i_10_65_2980_0 & ~i_10_65_3278_0 & i_10_65_3983_0 & ~i_10_65_4280_0))) | (i_10_65_1652_0 & ((~i_10_65_29_0 & ~i_10_65_437_0 & ~i_10_65_991_0 & ~i_10_65_1547_0 & i_10_65_1823_0 & ~i_10_65_2380_0 & ~i_10_65_3835_0) | (i_10_65_2362_0 & ~i_10_65_3980_0))) | (i_10_65_2724_0 & ~i_10_65_2822_0 & i_10_65_2832_0 & ~i_10_65_2983_0 & ~i_10_65_3835_0));
endmodule



// Benchmark "kernel_10_66" written by ABC on Sun Jul 19 10:22:09 2020

module kernel_10_66 ( 
    i_10_66_28_0, i_10_66_29_0, i_10_66_117_0, i_10_66_118_0,
    i_10_66_121_0, i_10_66_180_0, i_10_66_181_0, i_10_66_262_0,
    i_10_66_266_0, i_10_66_348_0, i_10_66_390_0, i_10_66_435_0,
    i_10_66_441_0, i_10_66_442_0, i_10_66_444_0, i_10_66_460_0,
    i_10_66_461_0, i_10_66_559_0, i_10_66_560_0, i_10_66_562_0,
    i_10_66_599_0, i_10_66_795_0, i_10_66_999_0, i_10_66_1027_0,
    i_10_66_1119_0, i_10_66_1165_0, i_10_66_1305_0, i_10_66_1357_0,
    i_10_66_1359_0, i_10_66_1360_0, i_10_66_1363_0, i_10_66_1366_0,
    i_10_66_1401_0, i_10_66_1477_0, i_10_66_1612_0, i_10_66_1652_0,
    i_10_66_1683_0, i_10_66_1691_0, i_10_66_1821_0, i_10_66_1908_0,
    i_10_66_1920_0, i_10_66_1947_0, i_10_66_1956_0, i_10_66_2309_0,
    i_10_66_2408_0, i_10_66_2452_0, i_10_66_2455_0, i_10_66_2482_0,
    i_10_66_2654_0, i_10_66_2656_0, i_10_66_2657_0, i_10_66_2658_0,
    i_10_66_2659_0, i_10_66_2703_0, i_10_66_2725_0, i_10_66_2744_0,
    i_10_66_2754_0, i_10_66_2755_0, i_10_66_2826_0, i_10_66_2828_0,
    i_10_66_3036_0, i_10_66_3203_0, i_10_66_3235_0, i_10_66_3268_0,
    i_10_66_3271_0, i_10_66_3284_0, i_10_66_3305_0, i_10_66_3349_0,
    i_10_66_3392_0, i_10_66_3473_0, i_10_66_3480_0, i_10_66_3494_0,
    i_10_66_3497_0, i_10_66_3561_0, i_10_66_3585_0, i_10_66_3586_0,
    i_10_66_3587_0, i_10_66_3589_0, i_10_66_3609_0, i_10_66_3610_0,
    i_10_66_3614_0, i_10_66_3620_0, i_10_66_3625_0, i_10_66_3646_0,
    i_10_66_3648_0, i_10_66_3649_0, i_10_66_3702_0, i_10_66_3788_0,
    i_10_66_3838_0, i_10_66_3853_0, i_10_66_3882_0, i_10_66_3883_0,
    i_10_66_3983_0, i_10_66_3985_0, i_10_66_4054_0, i_10_66_4055_0,
    i_10_66_4057_0, i_10_66_4118_0, i_10_66_4144_0, i_10_66_4145_0,
    o_10_66_0_0  );
  input  i_10_66_28_0, i_10_66_29_0, i_10_66_117_0, i_10_66_118_0,
    i_10_66_121_0, i_10_66_180_0, i_10_66_181_0, i_10_66_262_0,
    i_10_66_266_0, i_10_66_348_0, i_10_66_390_0, i_10_66_435_0,
    i_10_66_441_0, i_10_66_442_0, i_10_66_444_0, i_10_66_460_0,
    i_10_66_461_0, i_10_66_559_0, i_10_66_560_0, i_10_66_562_0,
    i_10_66_599_0, i_10_66_795_0, i_10_66_999_0, i_10_66_1027_0,
    i_10_66_1119_0, i_10_66_1165_0, i_10_66_1305_0, i_10_66_1357_0,
    i_10_66_1359_0, i_10_66_1360_0, i_10_66_1363_0, i_10_66_1366_0,
    i_10_66_1401_0, i_10_66_1477_0, i_10_66_1612_0, i_10_66_1652_0,
    i_10_66_1683_0, i_10_66_1691_0, i_10_66_1821_0, i_10_66_1908_0,
    i_10_66_1920_0, i_10_66_1947_0, i_10_66_1956_0, i_10_66_2309_0,
    i_10_66_2408_0, i_10_66_2452_0, i_10_66_2455_0, i_10_66_2482_0,
    i_10_66_2654_0, i_10_66_2656_0, i_10_66_2657_0, i_10_66_2658_0,
    i_10_66_2659_0, i_10_66_2703_0, i_10_66_2725_0, i_10_66_2744_0,
    i_10_66_2754_0, i_10_66_2755_0, i_10_66_2826_0, i_10_66_2828_0,
    i_10_66_3036_0, i_10_66_3203_0, i_10_66_3235_0, i_10_66_3268_0,
    i_10_66_3271_0, i_10_66_3284_0, i_10_66_3305_0, i_10_66_3349_0,
    i_10_66_3392_0, i_10_66_3473_0, i_10_66_3480_0, i_10_66_3494_0,
    i_10_66_3497_0, i_10_66_3561_0, i_10_66_3585_0, i_10_66_3586_0,
    i_10_66_3587_0, i_10_66_3589_0, i_10_66_3609_0, i_10_66_3610_0,
    i_10_66_3614_0, i_10_66_3620_0, i_10_66_3625_0, i_10_66_3646_0,
    i_10_66_3648_0, i_10_66_3649_0, i_10_66_3702_0, i_10_66_3788_0,
    i_10_66_3838_0, i_10_66_3853_0, i_10_66_3882_0, i_10_66_3883_0,
    i_10_66_3983_0, i_10_66_3985_0, i_10_66_4054_0, i_10_66_4055_0,
    i_10_66_4057_0, i_10_66_4118_0, i_10_66_4144_0, i_10_66_4145_0;
  output o_10_66_0_0;
  assign o_10_66_0_0 = 0;
endmodule



// Benchmark "kernel_10_67" written by ABC on Sun Jul 19 10:22:10 2020

module kernel_10_67 ( 
    i_10_67_144_0, i_10_67_146_0, i_10_67_219_0, i_10_67_223_0,
    i_10_67_387_0, i_10_67_388_0, i_10_67_423_0, i_10_67_424_0,
    i_10_67_425_0, i_10_67_426_0, i_10_67_427_0, i_10_67_445_0,
    i_10_67_460_0, i_10_67_462_0, i_10_67_463_0, i_10_67_507_0,
    i_10_67_508_0, i_10_67_693_0, i_10_67_711_0, i_10_67_747_0,
    i_10_67_795_0, i_10_67_796_0, i_10_67_900_0, i_10_67_995_0,
    i_10_67_1234_0, i_10_67_1243_0, i_10_67_1246_0, i_10_67_1248_0,
    i_10_67_1260_0, i_10_67_1305_0, i_10_67_1341_0, i_10_67_1485_0,
    i_10_67_1683_0, i_10_67_1819_0, i_10_67_1823_0, i_10_67_1825_0,
    i_10_67_1911_0, i_10_67_1999_0, i_10_67_2019_0, i_10_67_2241_0,
    i_10_67_2350_0, i_10_67_2351_0, i_10_67_2352_0, i_10_67_2353_0,
    i_10_67_2354_0, i_10_67_2356_0, i_10_67_2450_0, i_10_67_2451_0,
    i_10_67_2452_0, i_10_67_2538_0, i_10_67_2543_0, i_10_67_2678_0,
    i_10_67_2700_0, i_10_67_2701_0, i_10_67_2702_0, i_10_67_2710_0,
    i_10_67_2716_0, i_10_67_2820_0, i_10_67_2916_0, i_10_67_3037_0,
    i_10_67_3087_0, i_10_67_3088_0, i_10_67_3091_0, i_10_67_3114_0,
    i_10_67_3198_0, i_10_67_3237_0, i_10_67_3276_0, i_10_67_3277_0,
    i_10_67_3280_0, i_10_67_3312_0, i_10_67_3408_0, i_10_67_3409_0,
    i_10_67_3465_0, i_10_67_3538_0, i_10_67_3582_0, i_10_67_3583_0,
    i_10_67_3585_0, i_10_67_3586_0, i_10_67_3612_0, i_10_67_3613_0,
    i_10_67_3648_0, i_10_67_3682_0, i_10_67_3717_0, i_10_67_3780_0,
    i_10_67_3781_0, i_10_67_3786_0, i_10_67_3807_0, i_10_67_3808_0,
    i_10_67_3834_0, i_10_67_3835_0, i_10_67_3838_0, i_10_67_3841_0,
    i_10_67_3850_0, i_10_67_3857_0, i_10_67_3860_0, i_10_67_3985_0,
    i_10_67_4117_0, i_10_67_4169_0, i_10_67_4284_0, i_10_67_4290_0,
    o_10_67_0_0  );
  input  i_10_67_144_0, i_10_67_146_0, i_10_67_219_0, i_10_67_223_0,
    i_10_67_387_0, i_10_67_388_0, i_10_67_423_0, i_10_67_424_0,
    i_10_67_425_0, i_10_67_426_0, i_10_67_427_0, i_10_67_445_0,
    i_10_67_460_0, i_10_67_462_0, i_10_67_463_0, i_10_67_507_0,
    i_10_67_508_0, i_10_67_693_0, i_10_67_711_0, i_10_67_747_0,
    i_10_67_795_0, i_10_67_796_0, i_10_67_900_0, i_10_67_995_0,
    i_10_67_1234_0, i_10_67_1243_0, i_10_67_1246_0, i_10_67_1248_0,
    i_10_67_1260_0, i_10_67_1305_0, i_10_67_1341_0, i_10_67_1485_0,
    i_10_67_1683_0, i_10_67_1819_0, i_10_67_1823_0, i_10_67_1825_0,
    i_10_67_1911_0, i_10_67_1999_0, i_10_67_2019_0, i_10_67_2241_0,
    i_10_67_2350_0, i_10_67_2351_0, i_10_67_2352_0, i_10_67_2353_0,
    i_10_67_2354_0, i_10_67_2356_0, i_10_67_2450_0, i_10_67_2451_0,
    i_10_67_2452_0, i_10_67_2538_0, i_10_67_2543_0, i_10_67_2678_0,
    i_10_67_2700_0, i_10_67_2701_0, i_10_67_2702_0, i_10_67_2710_0,
    i_10_67_2716_0, i_10_67_2820_0, i_10_67_2916_0, i_10_67_3037_0,
    i_10_67_3087_0, i_10_67_3088_0, i_10_67_3091_0, i_10_67_3114_0,
    i_10_67_3198_0, i_10_67_3237_0, i_10_67_3276_0, i_10_67_3277_0,
    i_10_67_3280_0, i_10_67_3312_0, i_10_67_3408_0, i_10_67_3409_0,
    i_10_67_3465_0, i_10_67_3538_0, i_10_67_3582_0, i_10_67_3583_0,
    i_10_67_3585_0, i_10_67_3586_0, i_10_67_3612_0, i_10_67_3613_0,
    i_10_67_3648_0, i_10_67_3682_0, i_10_67_3717_0, i_10_67_3780_0,
    i_10_67_3781_0, i_10_67_3786_0, i_10_67_3807_0, i_10_67_3808_0,
    i_10_67_3834_0, i_10_67_3835_0, i_10_67_3838_0, i_10_67_3841_0,
    i_10_67_3850_0, i_10_67_3857_0, i_10_67_3860_0, i_10_67_3985_0,
    i_10_67_4117_0, i_10_67_4169_0, i_10_67_4284_0, i_10_67_4290_0;
  output o_10_67_0_0;
  assign o_10_67_0_0 = ~((~i_10_67_223_0 & ((~i_10_67_219_0 & (~i_10_67_424_0 | (i_10_67_460_0 & ~i_10_67_1341_0 & ~i_10_67_2356_0 & ~i_10_67_3276_0 & ~i_10_67_3465_0))) | (~i_10_67_423_0 & ~i_10_67_747_0 & ~i_10_67_795_0))) | (~i_10_67_387_0 & ((~i_10_67_1485_0 & ~i_10_67_1999_0 & ~i_10_67_2820_0) | (~i_10_67_711_0 & ~i_10_67_3312_0 & ~i_10_67_3613_0))) | (~i_10_67_900_0 & ~i_10_67_3091_0 & ((~i_10_67_795_0 & ~i_10_67_1999_0) | (~i_10_67_460_0 & ~i_10_67_1248_0 & ~i_10_67_1911_0 & ~i_10_67_3841_0 & ~i_10_67_3860_0 & ~i_10_67_3985_0))) | (~i_10_67_1683_0 & ((~i_10_67_463_0 & ~i_10_67_1825_0 & i_10_67_3835_0) | (~i_10_67_1234_0 & ~i_10_67_1485_0 & i_10_67_3857_0))) | (~i_10_67_1825_0 & ((~i_10_67_711_0 & i_10_67_1819_0 & ~i_10_67_3237_0 & ~i_10_67_3277_0) | (~i_10_67_2350_0 & ~i_10_67_2710_0 & ~i_10_67_3648_0 & ~i_10_67_3834_0 & ~i_10_67_3860_0))) | (i_10_67_1260_0 & ~i_10_67_2450_0 & ~i_10_67_3087_0) | (~i_10_67_445_0 & ~i_10_67_3280_0 & ~i_10_67_3613_0 & ~i_10_67_3860_0) | (~i_10_67_144_0 & ~i_10_67_388_0 & ~i_10_67_3237_0 & ~i_10_67_3857_0) | (~i_10_67_423_0 & i_10_67_3985_0) | (~i_10_67_146_0 & ~i_10_67_426_0 & ~i_10_67_995_0 & ~i_10_67_1819_0 & ~i_10_67_3312_0 & ~i_10_67_3838_0 & ~i_10_67_4117_0 & ~i_10_67_4290_0));
endmodule



// Benchmark "kernel_10_68" written by ABC on Sun Jul 19 10:22:11 2020

module kernel_10_68 ( 
    i_10_68_42_0, i_10_68_67_0, i_10_68_68_0, i_10_68_150_0, i_10_68_174_0,
    i_10_68_183_0, i_10_68_324_0, i_10_68_364_0, i_10_68_405_0,
    i_10_68_426_0, i_10_68_441_0, i_10_68_443_0, i_10_68_445_0,
    i_10_68_733_0, i_10_68_734_0, i_10_68_793_0, i_10_68_880_0,
    i_10_68_1119_0, i_10_68_1237_0, i_10_68_1243_0, i_10_68_1308_0,
    i_10_68_1309_0, i_10_68_1380_0, i_10_68_1609_0, i_10_68_1617_0,
    i_10_68_1618_0, i_10_68_1648_0, i_10_68_1649_0, i_10_68_1650_0,
    i_10_68_1689_0, i_10_68_1910_0, i_10_68_1960_0, i_10_68_1995_0,
    i_10_68_1996_0, i_10_68_2082_0, i_10_68_2355_0, i_10_68_2380_0,
    i_10_68_2448_0, i_10_68_2449_0, i_10_68_2450_0, i_10_68_2451_0,
    i_10_68_2452_0, i_10_68_2460_0, i_10_68_2511_0, i_10_68_2589_0,
    i_10_68_2590_0, i_10_68_2659_0, i_10_68_2701_0, i_10_68_2705_0,
    i_10_68_2708_0, i_10_68_2715_0, i_10_68_2716_0, i_10_68_2718_0,
    i_10_68_2730_0, i_10_68_2734_0, i_10_68_2787_0, i_10_68_2788_0,
    i_10_68_2828_0, i_10_68_2982_0, i_10_68_3048_0, i_10_68_3049_0,
    i_10_68_3171_0, i_10_68_3199_0, i_10_68_3271_0, i_10_68_3279_0,
    i_10_68_3289_0, i_10_68_3292_0, i_10_68_3391_0, i_10_68_3392_0,
    i_10_68_3471_0, i_10_68_3589_0, i_10_68_3609_0, i_10_68_3610_0,
    i_10_68_3611_0, i_10_68_3648_0, i_10_68_3649_0, i_10_68_3684_0,
    i_10_68_3720_0, i_10_68_3814_0, i_10_68_3815_0, i_10_68_3834_0,
    i_10_68_3837_0, i_10_68_3838_0, i_10_68_3855_0, i_10_68_3882_0,
    i_10_68_3893_0, i_10_68_3945_0, i_10_68_3987_0, i_10_68_4118_0,
    i_10_68_4182_0, i_10_68_4216_0, i_10_68_4218_0, i_10_68_4233_0,
    i_10_68_4234_0, i_10_68_4236_0, i_10_68_4237_0, i_10_68_4425_0,
    i_10_68_4426_0, i_10_68_4506_0, i_10_68_4507_0,
    o_10_68_0_0  );
  input  i_10_68_42_0, i_10_68_67_0, i_10_68_68_0, i_10_68_150_0,
    i_10_68_174_0, i_10_68_183_0, i_10_68_324_0, i_10_68_364_0,
    i_10_68_405_0, i_10_68_426_0, i_10_68_441_0, i_10_68_443_0,
    i_10_68_445_0, i_10_68_733_0, i_10_68_734_0, i_10_68_793_0,
    i_10_68_880_0, i_10_68_1119_0, i_10_68_1237_0, i_10_68_1243_0,
    i_10_68_1308_0, i_10_68_1309_0, i_10_68_1380_0, i_10_68_1609_0,
    i_10_68_1617_0, i_10_68_1618_0, i_10_68_1648_0, i_10_68_1649_0,
    i_10_68_1650_0, i_10_68_1689_0, i_10_68_1910_0, i_10_68_1960_0,
    i_10_68_1995_0, i_10_68_1996_0, i_10_68_2082_0, i_10_68_2355_0,
    i_10_68_2380_0, i_10_68_2448_0, i_10_68_2449_0, i_10_68_2450_0,
    i_10_68_2451_0, i_10_68_2452_0, i_10_68_2460_0, i_10_68_2511_0,
    i_10_68_2589_0, i_10_68_2590_0, i_10_68_2659_0, i_10_68_2701_0,
    i_10_68_2705_0, i_10_68_2708_0, i_10_68_2715_0, i_10_68_2716_0,
    i_10_68_2718_0, i_10_68_2730_0, i_10_68_2734_0, i_10_68_2787_0,
    i_10_68_2788_0, i_10_68_2828_0, i_10_68_2982_0, i_10_68_3048_0,
    i_10_68_3049_0, i_10_68_3171_0, i_10_68_3199_0, i_10_68_3271_0,
    i_10_68_3279_0, i_10_68_3289_0, i_10_68_3292_0, i_10_68_3391_0,
    i_10_68_3392_0, i_10_68_3471_0, i_10_68_3589_0, i_10_68_3609_0,
    i_10_68_3610_0, i_10_68_3611_0, i_10_68_3648_0, i_10_68_3649_0,
    i_10_68_3684_0, i_10_68_3720_0, i_10_68_3814_0, i_10_68_3815_0,
    i_10_68_3834_0, i_10_68_3837_0, i_10_68_3838_0, i_10_68_3855_0,
    i_10_68_3882_0, i_10_68_3893_0, i_10_68_3945_0, i_10_68_3987_0,
    i_10_68_4118_0, i_10_68_4182_0, i_10_68_4216_0, i_10_68_4218_0,
    i_10_68_4233_0, i_10_68_4234_0, i_10_68_4236_0, i_10_68_4237_0,
    i_10_68_4425_0, i_10_68_4426_0, i_10_68_4506_0, i_10_68_4507_0;
  output o_10_68_0_0;
  assign o_10_68_0_0 = 0;
endmodule



// Benchmark "kernel_10_69" written by ABC on Sun Jul 19 10:22:12 2020

module kernel_10_69 ( 
    i_10_69_27_0, i_10_69_28_0, i_10_69_122_0, i_10_69_171_0,
    i_10_69_190_0, i_10_69_239_0, i_10_69_292_0, i_10_69_369_0,
    i_10_69_387_0, i_10_69_430_0, i_10_69_465_0, i_10_69_512_0,
    i_10_69_546_0, i_10_69_547_0, i_10_69_711_0, i_10_69_717_0,
    i_10_69_759_0, i_10_69_907_0, i_10_69_1040_0, i_10_69_1120_0,
    i_10_69_1121_0, i_10_69_1179_0, i_10_69_1251_0, i_10_69_1273_0,
    i_10_69_1310_0, i_10_69_1345_0, i_10_69_1352_0, i_10_69_1380_0,
    i_10_69_1441_0, i_10_69_1545_0, i_10_69_1548_0, i_10_69_1578_0,
    i_10_69_1614_0, i_10_69_1616_0, i_10_69_1620_0, i_10_69_1632_0,
    i_10_69_1654_0, i_10_69_1803_0, i_10_69_2047_0, i_10_69_2160_0,
    i_10_69_2178_0, i_10_69_2180_0, i_10_69_2209_0, i_10_69_2290_0,
    i_10_69_2349_0, i_10_69_2352_0, i_10_69_2372_0, i_10_69_2448_0,
    i_10_69_2449_0, i_10_69_2452_0, i_10_69_2632_0, i_10_69_2686_0,
    i_10_69_2725_0, i_10_69_2829_0, i_10_69_2830_0, i_10_69_2834_0,
    i_10_69_2885_0, i_10_69_2922_0, i_10_69_2935_0, i_10_69_2936_0,
    i_10_69_3034_0, i_10_69_3035_0, i_10_69_3038_0, i_10_69_3046_0,
    i_10_69_3067_0, i_10_69_3231_0, i_10_69_3274_0, i_10_69_3291_0,
    i_10_69_3292_0, i_10_69_3293_0, i_10_69_3523_0, i_10_69_3554_0,
    i_10_69_3611_0, i_10_69_3612_0, i_10_69_3615_0, i_10_69_3621_0,
    i_10_69_3637_0, i_10_69_3685_0, i_10_69_3699_0, i_10_69_3703_0,
    i_10_69_3784_0, i_10_69_3786_0, i_10_69_3787_0, i_10_69_3859_0,
    i_10_69_3961_0, i_10_69_3965_0, i_10_69_4052_0, i_10_69_4091_0,
    i_10_69_4126_0, i_10_69_4153_0, i_10_69_4231_0, i_10_69_4233_0,
    i_10_69_4286_0, i_10_69_4304_0, i_10_69_4309_0, i_10_69_4310_0,
    i_10_69_4503_0, i_10_69_4529_0, i_10_69_4591_0, i_10_69_4592_0,
    o_10_69_0_0  );
  input  i_10_69_27_0, i_10_69_28_0, i_10_69_122_0, i_10_69_171_0,
    i_10_69_190_0, i_10_69_239_0, i_10_69_292_0, i_10_69_369_0,
    i_10_69_387_0, i_10_69_430_0, i_10_69_465_0, i_10_69_512_0,
    i_10_69_546_0, i_10_69_547_0, i_10_69_711_0, i_10_69_717_0,
    i_10_69_759_0, i_10_69_907_0, i_10_69_1040_0, i_10_69_1120_0,
    i_10_69_1121_0, i_10_69_1179_0, i_10_69_1251_0, i_10_69_1273_0,
    i_10_69_1310_0, i_10_69_1345_0, i_10_69_1352_0, i_10_69_1380_0,
    i_10_69_1441_0, i_10_69_1545_0, i_10_69_1548_0, i_10_69_1578_0,
    i_10_69_1614_0, i_10_69_1616_0, i_10_69_1620_0, i_10_69_1632_0,
    i_10_69_1654_0, i_10_69_1803_0, i_10_69_2047_0, i_10_69_2160_0,
    i_10_69_2178_0, i_10_69_2180_0, i_10_69_2209_0, i_10_69_2290_0,
    i_10_69_2349_0, i_10_69_2352_0, i_10_69_2372_0, i_10_69_2448_0,
    i_10_69_2449_0, i_10_69_2452_0, i_10_69_2632_0, i_10_69_2686_0,
    i_10_69_2725_0, i_10_69_2829_0, i_10_69_2830_0, i_10_69_2834_0,
    i_10_69_2885_0, i_10_69_2922_0, i_10_69_2935_0, i_10_69_2936_0,
    i_10_69_3034_0, i_10_69_3035_0, i_10_69_3038_0, i_10_69_3046_0,
    i_10_69_3067_0, i_10_69_3231_0, i_10_69_3274_0, i_10_69_3291_0,
    i_10_69_3292_0, i_10_69_3293_0, i_10_69_3523_0, i_10_69_3554_0,
    i_10_69_3611_0, i_10_69_3612_0, i_10_69_3615_0, i_10_69_3621_0,
    i_10_69_3637_0, i_10_69_3685_0, i_10_69_3699_0, i_10_69_3703_0,
    i_10_69_3784_0, i_10_69_3786_0, i_10_69_3787_0, i_10_69_3859_0,
    i_10_69_3961_0, i_10_69_3965_0, i_10_69_4052_0, i_10_69_4091_0,
    i_10_69_4126_0, i_10_69_4153_0, i_10_69_4231_0, i_10_69_4233_0,
    i_10_69_4286_0, i_10_69_4304_0, i_10_69_4309_0, i_10_69_4310_0,
    i_10_69_4503_0, i_10_69_4529_0, i_10_69_4591_0, i_10_69_4592_0;
  output o_10_69_0_0;
  assign o_10_69_0_0 = 0;
endmodule



// Benchmark "kernel_10_70" written by ABC on Sun Jul 19 10:22:13 2020

module kernel_10_70 ( 
    i_10_70_37_0, i_10_70_40_0, i_10_70_52_0, i_10_70_247_0, i_10_70_286_0,
    i_10_70_315_0, i_10_70_316_0, i_10_70_320_0, i_10_70_321_0,
    i_10_70_322_0, i_10_70_323_0, i_10_70_408_0, i_10_70_409_0,
    i_10_70_410_0, i_10_70_430_0, i_10_70_439_0, i_10_70_691_0,
    i_10_70_832_0, i_10_70_833_0, i_10_70_994_0, i_10_70_1027_0,
    i_10_70_1030_0, i_10_70_1031_0, i_10_70_1040_0, i_10_70_1048_0,
    i_10_70_1082_0, i_10_70_1164_0, i_10_70_1165_0, i_10_70_1166_0,
    i_10_70_1223_0, i_10_70_1233_0, i_10_70_1243_0, i_10_70_1265_0,
    i_10_70_1267_0, i_10_70_1268_0, i_10_70_1344_0, i_10_70_1345_0,
    i_10_70_1543_0, i_10_70_1544_0, i_10_70_1575_0, i_10_70_1578_0,
    i_10_70_1580_0, i_10_70_1650_0, i_10_70_1651_0, i_10_70_1654_0,
    i_10_70_1713_0, i_10_70_1825_0, i_10_70_1914_0, i_10_70_2017_0,
    i_10_70_2024_0, i_10_70_2204_0, i_10_70_2242_0, i_10_70_2251_0,
    i_10_70_2364_0, i_10_70_2459_0, i_10_70_2607_0, i_10_70_2657_0,
    i_10_70_2661_0, i_10_70_2662_0, i_10_70_2703_0, i_10_70_2704_0,
    i_10_70_2705_0, i_10_70_2707_0, i_10_70_2724_0, i_10_70_2833_0,
    i_10_70_2880_0, i_10_70_2982_0, i_10_70_2983_0, i_10_70_3069_0,
    i_10_70_3237_0, i_10_70_3279_0, i_10_70_3280_0, i_10_70_3288_0,
    i_10_70_3496_0, i_10_70_3497_0, i_10_70_3523_0, i_10_70_3525_0,
    i_10_70_3526_0, i_10_70_3615_0, i_10_70_3787_0, i_10_70_3788_0,
    i_10_70_3852_0, i_10_70_3856_0, i_10_70_3910_0, i_10_70_3913_0,
    i_10_70_3987_0, i_10_70_4116_0, i_10_70_4117_0, i_10_70_4118_0,
    i_10_70_4119_0, i_10_70_4125_0, i_10_70_4129_0, i_10_70_4170_0,
    i_10_70_4173_0, i_10_70_4215_0, i_10_70_4226_0, i_10_70_4272_0,
    i_10_70_4275_0, i_10_70_4565_0, i_10_70_4568_0,
    o_10_70_0_0  );
  input  i_10_70_37_0, i_10_70_40_0, i_10_70_52_0, i_10_70_247_0,
    i_10_70_286_0, i_10_70_315_0, i_10_70_316_0, i_10_70_320_0,
    i_10_70_321_0, i_10_70_322_0, i_10_70_323_0, i_10_70_408_0,
    i_10_70_409_0, i_10_70_410_0, i_10_70_430_0, i_10_70_439_0,
    i_10_70_691_0, i_10_70_832_0, i_10_70_833_0, i_10_70_994_0,
    i_10_70_1027_0, i_10_70_1030_0, i_10_70_1031_0, i_10_70_1040_0,
    i_10_70_1048_0, i_10_70_1082_0, i_10_70_1164_0, i_10_70_1165_0,
    i_10_70_1166_0, i_10_70_1223_0, i_10_70_1233_0, i_10_70_1243_0,
    i_10_70_1265_0, i_10_70_1267_0, i_10_70_1268_0, i_10_70_1344_0,
    i_10_70_1345_0, i_10_70_1543_0, i_10_70_1544_0, i_10_70_1575_0,
    i_10_70_1578_0, i_10_70_1580_0, i_10_70_1650_0, i_10_70_1651_0,
    i_10_70_1654_0, i_10_70_1713_0, i_10_70_1825_0, i_10_70_1914_0,
    i_10_70_2017_0, i_10_70_2024_0, i_10_70_2204_0, i_10_70_2242_0,
    i_10_70_2251_0, i_10_70_2364_0, i_10_70_2459_0, i_10_70_2607_0,
    i_10_70_2657_0, i_10_70_2661_0, i_10_70_2662_0, i_10_70_2703_0,
    i_10_70_2704_0, i_10_70_2705_0, i_10_70_2707_0, i_10_70_2724_0,
    i_10_70_2833_0, i_10_70_2880_0, i_10_70_2982_0, i_10_70_2983_0,
    i_10_70_3069_0, i_10_70_3237_0, i_10_70_3279_0, i_10_70_3280_0,
    i_10_70_3288_0, i_10_70_3496_0, i_10_70_3497_0, i_10_70_3523_0,
    i_10_70_3525_0, i_10_70_3526_0, i_10_70_3615_0, i_10_70_3787_0,
    i_10_70_3788_0, i_10_70_3852_0, i_10_70_3856_0, i_10_70_3910_0,
    i_10_70_3913_0, i_10_70_3987_0, i_10_70_4116_0, i_10_70_4117_0,
    i_10_70_4118_0, i_10_70_4119_0, i_10_70_4125_0, i_10_70_4129_0,
    i_10_70_4170_0, i_10_70_4173_0, i_10_70_4215_0, i_10_70_4226_0,
    i_10_70_4272_0, i_10_70_4275_0, i_10_70_4565_0, i_10_70_4568_0;
  output o_10_70_0_0;
  assign o_10_70_0_0 = 0;
endmodule



// Benchmark "kernel_10_71" written by ABC on Sun Jul 19 10:22:14 2020

module kernel_10_71 ( 
    i_10_71_29_0, i_10_71_118_0, i_10_71_259_0, i_10_71_260_0,
    i_10_71_280_0, i_10_71_317_0, i_10_71_331_0, i_10_71_332_0,
    i_10_71_373_0, i_10_71_387_0, i_10_71_388_0, i_10_71_391_0,
    i_10_71_439_0, i_10_71_462_0, i_10_71_517_0, i_10_71_518_0,
    i_10_71_959_0, i_10_71_967_0, i_10_71_1031_0, i_10_71_1043_0,
    i_10_71_1057_0, i_10_71_1058_0, i_10_71_1083_0, i_10_71_1084_0,
    i_10_71_1139_0, i_10_71_1233_0, i_10_71_1234_0, i_10_71_1235_0,
    i_10_71_1237_0, i_10_71_1238_0, i_10_71_1240_0, i_10_71_1291_0,
    i_10_71_1312_0, i_10_71_1431_0, i_10_71_1433_0, i_10_71_1539_0,
    i_10_71_1540_0, i_10_71_1576_0, i_10_71_1577_0, i_10_71_1621_0,
    i_10_71_1654_0, i_10_71_1717_0, i_10_71_1764_0, i_10_71_1768_0,
    i_10_71_1769_0, i_10_71_1822_0, i_10_71_1824_0, i_10_71_1825_0,
    i_10_71_1826_0, i_10_71_1958_0, i_10_71_1980_0, i_10_71_1981_0,
    i_10_71_1984_0, i_10_71_2017_0, i_10_71_2020_0, i_10_71_2351_0,
    i_10_71_2356_0, i_10_71_2452_0, i_10_71_2471_0, i_10_71_2546_0,
    i_10_71_2565_0, i_10_71_2566_0, i_10_71_2581_0, i_10_71_2628_0,
    i_10_71_2631_0, i_10_71_2632_0, i_10_71_2635_0, i_10_71_2659_0,
    i_10_71_2704_0, i_10_71_2705_0, i_10_71_2713_0, i_10_71_2734_0,
    i_10_71_2824_0, i_10_71_2830_0, i_10_71_2921_0, i_10_71_3035_0,
    i_10_71_3039_0, i_10_71_3050_0, i_10_71_3073_0, i_10_71_3196_0,
    i_10_71_3323_0, i_10_71_3586_0, i_10_71_3612_0, i_10_71_3619_0,
    i_10_71_3620_0, i_10_71_3720_0, i_10_71_3786_0, i_10_71_3910_0,
    i_10_71_3947_0, i_10_71_3983_0, i_10_71_4004_0, i_10_71_4051_0,
    i_10_71_4054_0, i_10_71_4123_0, i_10_71_4168_0, i_10_71_4169_0,
    i_10_71_4171_0, i_10_71_4192_0, i_10_71_4282_0, i_10_71_4530_0,
    o_10_71_0_0  );
  input  i_10_71_29_0, i_10_71_118_0, i_10_71_259_0, i_10_71_260_0,
    i_10_71_280_0, i_10_71_317_0, i_10_71_331_0, i_10_71_332_0,
    i_10_71_373_0, i_10_71_387_0, i_10_71_388_0, i_10_71_391_0,
    i_10_71_439_0, i_10_71_462_0, i_10_71_517_0, i_10_71_518_0,
    i_10_71_959_0, i_10_71_967_0, i_10_71_1031_0, i_10_71_1043_0,
    i_10_71_1057_0, i_10_71_1058_0, i_10_71_1083_0, i_10_71_1084_0,
    i_10_71_1139_0, i_10_71_1233_0, i_10_71_1234_0, i_10_71_1235_0,
    i_10_71_1237_0, i_10_71_1238_0, i_10_71_1240_0, i_10_71_1291_0,
    i_10_71_1312_0, i_10_71_1431_0, i_10_71_1433_0, i_10_71_1539_0,
    i_10_71_1540_0, i_10_71_1576_0, i_10_71_1577_0, i_10_71_1621_0,
    i_10_71_1654_0, i_10_71_1717_0, i_10_71_1764_0, i_10_71_1768_0,
    i_10_71_1769_0, i_10_71_1822_0, i_10_71_1824_0, i_10_71_1825_0,
    i_10_71_1826_0, i_10_71_1958_0, i_10_71_1980_0, i_10_71_1981_0,
    i_10_71_1984_0, i_10_71_2017_0, i_10_71_2020_0, i_10_71_2351_0,
    i_10_71_2356_0, i_10_71_2452_0, i_10_71_2471_0, i_10_71_2546_0,
    i_10_71_2565_0, i_10_71_2566_0, i_10_71_2581_0, i_10_71_2628_0,
    i_10_71_2631_0, i_10_71_2632_0, i_10_71_2635_0, i_10_71_2659_0,
    i_10_71_2704_0, i_10_71_2705_0, i_10_71_2713_0, i_10_71_2734_0,
    i_10_71_2824_0, i_10_71_2830_0, i_10_71_2921_0, i_10_71_3035_0,
    i_10_71_3039_0, i_10_71_3050_0, i_10_71_3073_0, i_10_71_3196_0,
    i_10_71_3323_0, i_10_71_3586_0, i_10_71_3612_0, i_10_71_3619_0,
    i_10_71_3620_0, i_10_71_3720_0, i_10_71_3786_0, i_10_71_3910_0,
    i_10_71_3947_0, i_10_71_3983_0, i_10_71_4004_0, i_10_71_4051_0,
    i_10_71_4054_0, i_10_71_4123_0, i_10_71_4168_0, i_10_71_4169_0,
    i_10_71_4171_0, i_10_71_4192_0, i_10_71_4282_0, i_10_71_4530_0;
  output o_10_71_0_0;
  assign o_10_71_0_0 = 0;
endmodule



// Benchmark "kernel_10_72" written by ABC on Sun Jul 19 10:22:15 2020

module kernel_10_72 ( 
    i_10_72_174_0, i_10_72_183_0, i_10_72_408_0, i_10_72_424_0,
    i_10_72_447_0, i_10_72_515_0, i_10_72_517_0, i_10_72_637_0,
    i_10_72_798_0, i_10_72_903_0, i_10_72_962_0, i_10_72_967_0,
    i_10_72_968_0, i_10_72_996_0, i_10_72_1032_0, i_10_72_1087_0,
    i_10_72_1236_0, i_10_72_1237_0, i_10_72_1238_0, i_10_72_1246_0,
    i_10_72_1247_0, i_10_72_1249_0, i_10_72_1250_0, i_10_72_1491_0,
    i_10_72_1544_0, i_10_72_1619_0, i_10_72_1647_0, i_10_72_1689_0,
    i_10_72_1821_0, i_10_72_1823_0, i_10_72_1825_0, i_10_72_1912_0,
    i_10_72_1945_0, i_10_72_2008_0, i_10_72_2311_0, i_10_72_2382_0,
    i_10_72_2383_0, i_10_72_2450_0, i_10_72_2452_0, i_10_72_2453_0,
    i_10_72_2470_0, i_10_72_2471_0, i_10_72_2643_0, i_10_72_2644_0,
    i_10_72_2681_0, i_10_72_2715_0, i_10_72_2716_0, i_10_72_2721_0,
    i_10_72_2722_0, i_10_72_2730_0, i_10_72_2732_0, i_10_72_2733_0,
    i_10_72_2785_0, i_10_72_2827_0, i_10_72_2833_0, i_10_72_2834_0,
    i_10_72_2880_0, i_10_72_2917_0, i_10_72_2920_0, i_10_72_2921_0,
    i_10_72_3035_0, i_10_72_3043_0, i_10_72_3044_0, i_10_72_3069_0,
    i_10_72_3072_0, i_10_72_3164_0, i_10_72_3199_0, i_10_72_3282_0,
    i_10_72_3387_0, i_10_72_3390_0, i_10_72_3391_0, i_10_72_3406_0,
    i_10_72_3468_0, i_10_72_3495_0, i_10_72_3496_0, i_10_72_3506_0,
    i_10_72_3526_0, i_10_72_3583_0, i_10_72_3586_0, i_10_72_3587_0,
    i_10_72_3589_0, i_10_72_3613_0, i_10_72_3616_0, i_10_72_3617_0,
    i_10_72_3648_0, i_10_72_3652_0, i_10_72_3653_0, i_10_72_3783_0,
    i_10_72_3784_0, i_10_72_3785_0, i_10_72_3786_0, i_10_72_3854_0,
    i_10_72_3878_0, i_10_72_4115_0, i_10_72_4126_0, i_10_72_4213_0,
    i_10_72_4218_0, i_10_72_4272_0, i_10_72_4273_0, i_10_72_4568_0,
    o_10_72_0_0  );
  input  i_10_72_174_0, i_10_72_183_0, i_10_72_408_0, i_10_72_424_0,
    i_10_72_447_0, i_10_72_515_0, i_10_72_517_0, i_10_72_637_0,
    i_10_72_798_0, i_10_72_903_0, i_10_72_962_0, i_10_72_967_0,
    i_10_72_968_0, i_10_72_996_0, i_10_72_1032_0, i_10_72_1087_0,
    i_10_72_1236_0, i_10_72_1237_0, i_10_72_1238_0, i_10_72_1246_0,
    i_10_72_1247_0, i_10_72_1249_0, i_10_72_1250_0, i_10_72_1491_0,
    i_10_72_1544_0, i_10_72_1619_0, i_10_72_1647_0, i_10_72_1689_0,
    i_10_72_1821_0, i_10_72_1823_0, i_10_72_1825_0, i_10_72_1912_0,
    i_10_72_1945_0, i_10_72_2008_0, i_10_72_2311_0, i_10_72_2382_0,
    i_10_72_2383_0, i_10_72_2450_0, i_10_72_2452_0, i_10_72_2453_0,
    i_10_72_2470_0, i_10_72_2471_0, i_10_72_2643_0, i_10_72_2644_0,
    i_10_72_2681_0, i_10_72_2715_0, i_10_72_2716_0, i_10_72_2721_0,
    i_10_72_2722_0, i_10_72_2730_0, i_10_72_2732_0, i_10_72_2733_0,
    i_10_72_2785_0, i_10_72_2827_0, i_10_72_2833_0, i_10_72_2834_0,
    i_10_72_2880_0, i_10_72_2917_0, i_10_72_2920_0, i_10_72_2921_0,
    i_10_72_3035_0, i_10_72_3043_0, i_10_72_3044_0, i_10_72_3069_0,
    i_10_72_3072_0, i_10_72_3164_0, i_10_72_3199_0, i_10_72_3282_0,
    i_10_72_3387_0, i_10_72_3390_0, i_10_72_3391_0, i_10_72_3406_0,
    i_10_72_3468_0, i_10_72_3495_0, i_10_72_3496_0, i_10_72_3506_0,
    i_10_72_3526_0, i_10_72_3583_0, i_10_72_3586_0, i_10_72_3587_0,
    i_10_72_3589_0, i_10_72_3613_0, i_10_72_3616_0, i_10_72_3617_0,
    i_10_72_3648_0, i_10_72_3652_0, i_10_72_3653_0, i_10_72_3783_0,
    i_10_72_3784_0, i_10_72_3785_0, i_10_72_3786_0, i_10_72_3854_0,
    i_10_72_3878_0, i_10_72_4115_0, i_10_72_4126_0, i_10_72_4213_0,
    i_10_72_4218_0, i_10_72_4272_0, i_10_72_4273_0, i_10_72_4568_0;
  output o_10_72_0_0;
  assign o_10_72_0_0 = 0;
endmodule



// Benchmark "kernel_10_73" written by ABC on Sun Jul 19 10:22:16 2020

module kernel_10_73 ( 
    i_10_73_270_0, i_10_73_273_0, i_10_73_282_0, i_10_73_283_0,
    i_10_73_284_0, i_10_73_289_0, i_10_73_290_0, i_10_73_293_0,
    i_10_73_315_0, i_10_73_391_0, i_10_73_408_0, i_10_73_411_0,
    i_10_73_424_0, i_10_73_425_0, i_10_73_441_0, i_10_73_442_0,
    i_10_73_794_0, i_10_73_1163_0, i_10_73_1310_0, i_10_73_1360_0,
    i_10_73_1361_0, i_10_73_1444_0, i_10_73_1445_0, i_10_73_1540_0,
    i_10_73_1543_0, i_10_73_1575_0, i_10_73_1577_0, i_10_73_1579_0,
    i_10_73_1649_0, i_10_73_1650_0, i_10_73_1651_0, i_10_73_1688_0,
    i_10_73_1721_0, i_10_73_1818_0, i_10_73_1819_0, i_10_73_1821_0,
    i_10_73_1946_0, i_10_73_1991_0, i_10_73_1993_0, i_10_73_2183_0,
    i_10_73_2197_0, i_10_73_2350_0, i_10_73_2353_0, i_10_73_2358_0,
    i_10_73_2359_0, i_10_73_2458_0, i_10_73_2471_0, i_10_73_2629_0,
    i_10_73_2630_0, i_10_73_2632_0, i_10_73_2634_0, i_10_73_2656_0,
    i_10_73_2657_0, i_10_73_2659_0, i_10_73_2660_0, i_10_73_2674_0,
    i_10_73_2675_0, i_10_73_2700_0, i_10_73_2703_0, i_10_73_2710_0,
    i_10_73_2711_0, i_10_73_2719_0, i_10_73_2721_0, i_10_73_2722_0,
    i_10_73_2724_0, i_10_73_2828_0, i_10_73_2829_0, i_10_73_2830_0,
    i_10_73_2885_0, i_10_73_2983_0, i_10_73_3043_0, i_10_73_3088_0,
    i_10_73_3089_0, i_10_73_3201_0, i_10_73_3232_0, i_10_73_3233_0,
    i_10_73_3328_0, i_10_73_3349_0, i_10_73_3350_0, i_10_73_3390_0,
    i_10_73_3431_0, i_10_73_3523_0, i_10_73_3527_0, i_10_73_3549_0,
    i_10_73_3586_0, i_10_73_3587_0, i_10_73_3609_0, i_10_73_3610_0,
    i_10_73_3835_0, i_10_73_3845_0, i_10_73_3859_0, i_10_73_3944_0,
    i_10_73_3983_0, i_10_73_4052_0, i_10_73_4168_0, i_10_73_4169_0,
    i_10_73_4275_0, i_10_73_4284_0, i_10_73_4567_0, i_10_73_4568_0,
    o_10_73_0_0  );
  input  i_10_73_270_0, i_10_73_273_0, i_10_73_282_0, i_10_73_283_0,
    i_10_73_284_0, i_10_73_289_0, i_10_73_290_0, i_10_73_293_0,
    i_10_73_315_0, i_10_73_391_0, i_10_73_408_0, i_10_73_411_0,
    i_10_73_424_0, i_10_73_425_0, i_10_73_441_0, i_10_73_442_0,
    i_10_73_794_0, i_10_73_1163_0, i_10_73_1310_0, i_10_73_1360_0,
    i_10_73_1361_0, i_10_73_1444_0, i_10_73_1445_0, i_10_73_1540_0,
    i_10_73_1543_0, i_10_73_1575_0, i_10_73_1577_0, i_10_73_1579_0,
    i_10_73_1649_0, i_10_73_1650_0, i_10_73_1651_0, i_10_73_1688_0,
    i_10_73_1721_0, i_10_73_1818_0, i_10_73_1819_0, i_10_73_1821_0,
    i_10_73_1946_0, i_10_73_1991_0, i_10_73_1993_0, i_10_73_2183_0,
    i_10_73_2197_0, i_10_73_2350_0, i_10_73_2353_0, i_10_73_2358_0,
    i_10_73_2359_0, i_10_73_2458_0, i_10_73_2471_0, i_10_73_2629_0,
    i_10_73_2630_0, i_10_73_2632_0, i_10_73_2634_0, i_10_73_2656_0,
    i_10_73_2657_0, i_10_73_2659_0, i_10_73_2660_0, i_10_73_2674_0,
    i_10_73_2675_0, i_10_73_2700_0, i_10_73_2703_0, i_10_73_2710_0,
    i_10_73_2711_0, i_10_73_2719_0, i_10_73_2721_0, i_10_73_2722_0,
    i_10_73_2724_0, i_10_73_2828_0, i_10_73_2829_0, i_10_73_2830_0,
    i_10_73_2885_0, i_10_73_2983_0, i_10_73_3043_0, i_10_73_3088_0,
    i_10_73_3089_0, i_10_73_3201_0, i_10_73_3232_0, i_10_73_3233_0,
    i_10_73_3328_0, i_10_73_3349_0, i_10_73_3350_0, i_10_73_3390_0,
    i_10_73_3431_0, i_10_73_3523_0, i_10_73_3527_0, i_10_73_3549_0,
    i_10_73_3586_0, i_10_73_3587_0, i_10_73_3609_0, i_10_73_3610_0,
    i_10_73_3835_0, i_10_73_3845_0, i_10_73_3859_0, i_10_73_3944_0,
    i_10_73_3983_0, i_10_73_4052_0, i_10_73_4168_0, i_10_73_4169_0,
    i_10_73_4275_0, i_10_73_4284_0, i_10_73_4567_0, i_10_73_4568_0;
  output o_10_73_0_0;
  assign o_10_73_0_0 = ~((~i_10_73_282_0 & ((~i_10_73_284_0 & ~i_10_73_293_0 & i_10_73_1819_0 & ~i_10_73_2656_0 & ~i_10_73_2674_0) | (~i_10_73_289_0 & ~i_10_73_1163_0 & ~i_10_73_1444_0 & ~i_10_73_2660_0 & ~i_10_73_3201_0 & ~i_10_73_3845_0 & ~i_10_73_4052_0))) | (~i_10_73_3088_0 & ((~i_10_73_290_0 & ((~i_10_73_425_0 & ~i_10_73_1991_0 & ~i_10_73_2722_0 & ~i_10_73_2829_0) | (~i_10_73_284_0 & ~i_10_73_441_0 & ~i_10_73_1445_0 & ~i_10_73_2358_0 & ~i_10_73_3089_0 & ~i_10_73_3233_0 & ~i_10_73_3944_0))) | (~i_10_73_3233_0 & ((i_10_73_442_0 & ~i_10_73_1649_0 & ~i_10_73_2710_0 & ~i_10_73_2828_0) | (~i_10_73_3089_0 & ~i_10_73_3586_0 & ~i_10_73_3587_0 & ~i_10_73_4567_0))))) | (~i_10_73_293_0 & ((~i_10_73_391_0 & ~i_10_73_1444_0 & ~i_10_73_1445_0 & ~i_10_73_1993_0 & ~i_10_73_2471_0 & ~i_10_73_2657_0 & ~i_10_73_2719_0 & ~i_10_73_3549_0) | (~i_10_73_1361_0 & ~i_10_73_2660_0 & ~i_10_73_2674_0 & ~i_10_73_3089_0 & ~i_10_73_4567_0))) | (~i_10_73_3549_0 & ((~i_10_73_284_0 & ((~i_10_73_425_0 & i_10_73_1818_0) | (~i_10_73_2675_0 & ~i_10_73_2724_0 & ~i_10_73_2830_0 & ~i_10_73_3523_0 & ~i_10_73_4052_0))) | (~i_10_73_289_0 & ~i_10_73_411_0 & ~i_10_73_425_0 & ~i_10_73_442_0 & ~i_10_73_1444_0 & ~i_10_73_1445_0))) | (~i_10_73_1821_0 & ((~i_10_73_1360_0 & ~i_10_73_1361_0 & ~i_10_73_1445_0 & i_10_73_1649_0 & ~i_10_73_2471_0 & ~i_10_73_2710_0) | (~i_10_73_1310_0 & i_10_73_1651_0 & ~i_10_73_3586_0 & ~i_10_73_4052_0))) | (~i_10_73_2711_0 & ((~i_10_73_284_0 & i_10_73_441_0 & ~i_10_73_3232_0 & i_10_73_3610_0) | (~i_10_73_2656_0 & ~i_10_73_2659_0 & ~i_10_73_2660_0 & ~i_10_73_2719_0 & ~i_10_73_3201_0 & ~i_10_73_4052_0))) | (~i_10_73_424_0 & ~i_10_73_1991_0 & ~i_10_73_3527_0 & i_10_73_3835_0) | (~i_10_73_2634_0 & ~i_10_73_2657_0 & ~i_10_73_2719_0 & ~i_10_73_2830_0 & ~i_10_73_3232_0 & i_10_73_3859_0) | (~i_10_73_1444_0 & i_10_73_2656_0 & i_10_73_2660_0 & ~i_10_73_3089_0 & i_10_73_3983_0) | (i_10_73_2358_0 & i_10_73_2630_0 & ~i_10_73_3043_0 & i_10_73_4568_0));
endmodule



// Benchmark "kernel_10_74" written by ABC on Sun Jul 19 10:22:17 2020

module kernel_10_74 ( 
    i_10_74_26_0, i_10_74_208_0, i_10_74_248_0, i_10_74_257_0,
    i_10_74_272_0, i_10_74_275_0, i_10_74_391_0, i_10_74_394_0,
    i_10_74_408_0, i_10_74_443_0, i_10_74_445_0, i_10_74_520_0,
    i_10_74_716_0, i_10_74_729_0, i_10_74_797_0, i_10_74_799_0,
    i_10_74_955_0, i_10_74_970_0, i_10_74_971_0, i_10_74_1037_0,
    i_10_74_1235_0, i_10_74_1243_0, i_10_74_1244_0, i_10_74_1246_0,
    i_10_74_1247_0, i_10_74_1310_0, i_10_74_1541_0, i_10_74_1544_0,
    i_10_74_1550_0, i_10_74_1552_0, i_10_74_1655_0, i_10_74_1688_0,
    i_10_74_1759_0, i_10_74_1909_0, i_10_74_1910_0, i_10_74_1911_0,
    i_10_74_1957_0, i_10_74_2008_0, i_10_74_2027_0, i_10_74_2155_0,
    i_10_74_2180_0, i_10_74_2242_0, i_10_74_2334_0, i_10_74_2336_0,
    i_10_74_2339_0, i_10_74_2379_0, i_10_74_2405_0, i_10_74_2411_0,
    i_10_74_2441_0, i_10_74_2442_0, i_10_74_2456_0, i_10_74_2506_0,
    i_10_74_2531_0, i_10_74_2534_0, i_10_74_2629_0, i_10_74_2637_0,
    i_10_74_2638_0, i_10_74_2640_0, i_10_74_2647_0, i_10_74_2702_0,
    i_10_74_2723_0, i_10_74_2729_0, i_10_74_2866_0, i_10_74_2920_0,
    i_10_74_2954_0, i_10_74_3033_0, i_10_74_3034_0, i_10_74_3036_0,
    i_10_74_3074_0, i_10_74_3197_0, i_10_74_3205_0, i_10_74_3224_0,
    i_10_74_3226_0, i_10_74_3286_0, i_10_74_3331_0, i_10_74_3332_0,
    i_10_74_3585_0, i_10_74_3650_0, i_10_74_3787_0, i_10_74_3817_0,
    i_10_74_3851_0, i_10_74_3860_0, i_10_74_3944_0, i_10_74_3965_0,
    i_10_74_4113_0, i_10_74_4117_0, i_10_74_4118_0, i_10_74_4185_0,
    i_10_74_4186_0, i_10_74_4188_0, i_10_74_4267_0, i_10_74_4268_0,
    i_10_74_4270_0, i_10_74_4271_0, i_10_74_4286_0, i_10_74_4289_0,
    i_10_74_4514_0, i_10_74_4528_0, i_10_74_4564_0, i_10_74_4566_0,
    o_10_74_0_0  );
  input  i_10_74_26_0, i_10_74_208_0, i_10_74_248_0, i_10_74_257_0,
    i_10_74_272_0, i_10_74_275_0, i_10_74_391_0, i_10_74_394_0,
    i_10_74_408_0, i_10_74_443_0, i_10_74_445_0, i_10_74_520_0,
    i_10_74_716_0, i_10_74_729_0, i_10_74_797_0, i_10_74_799_0,
    i_10_74_955_0, i_10_74_970_0, i_10_74_971_0, i_10_74_1037_0,
    i_10_74_1235_0, i_10_74_1243_0, i_10_74_1244_0, i_10_74_1246_0,
    i_10_74_1247_0, i_10_74_1310_0, i_10_74_1541_0, i_10_74_1544_0,
    i_10_74_1550_0, i_10_74_1552_0, i_10_74_1655_0, i_10_74_1688_0,
    i_10_74_1759_0, i_10_74_1909_0, i_10_74_1910_0, i_10_74_1911_0,
    i_10_74_1957_0, i_10_74_2008_0, i_10_74_2027_0, i_10_74_2155_0,
    i_10_74_2180_0, i_10_74_2242_0, i_10_74_2334_0, i_10_74_2336_0,
    i_10_74_2339_0, i_10_74_2379_0, i_10_74_2405_0, i_10_74_2411_0,
    i_10_74_2441_0, i_10_74_2442_0, i_10_74_2456_0, i_10_74_2506_0,
    i_10_74_2531_0, i_10_74_2534_0, i_10_74_2629_0, i_10_74_2637_0,
    i_10_74_2638_0, i_10_74_2640_0, i_10_74_2647_0, i_10_74_2702_0,
    i_10_74_2723_0, i_10_74_2729_0, i_10_74_2866_0, i_10_74_2920_0,
    i_10_74_2954_0, i_10_74_3033_0, i_10_74_3034_0, i_10_74_3036_0,
    i_10_74_3074_0, i_10_74_3197_0, i_10_74_3205_0, i_10_74_3224_0,
    i_10_74_3226_0, i_10_74_3286_0, i_10_74_3331_0, i_10_74_3332_0,
    i_10_74_3585_0, i_10_74_3650_0, i_10_74_3787_0, i_10_74_3817_0,
    i_10_74_3851_0, i_10_74_3860_0, i_10_74_3944_0, i_10_74_3965_0,
    i_10_74_4113_0, i_10_74_4117_0, i_10_74_4118_0, i_10_74_4185_0,
    i_10_74_4186_0, i_10_74_4188_0, i_10_74_4267_0, i_10_74_4268_0,
    i_10_74_4270_0, i_10_74_4271_0, i_10_74_4286_0, i_10_74_4289_0,
    i_10_74_4514_0, i_10_74_4528_0, i_10_74_4564_0, i_10_74_4566_0;
  output o_10_74_0_0;
  assign o_10_74_0_0 = 0;
endmodule



// Benchmark "kernel_10_75" written by ABC on Sun Jul 19 10:22:18 2020

module kernel_10_75 ( 
    i_10_75_38_0, i_10_75_49_0, i_10_75_66_0, i_10_75_69_0, i_10_75_155_0,
    i_10_75_191_0, i_10_75_194_0, i_10_75_218_0, i_10_75_237_0,
    i_10_75_246_0, i_10_75_425_0, i_10_75_442_0, i_10_75_460_0,
    i_10_75_595_0, i_10_75_621_0, i_10_75_794_0, i_10_75_958_0,
    i_10_75_995_0, i_10_75_1026_0, i_10_75_1245_0, i_10_75_1246_0,
    i_10_75_1299_0, i_10_75_1310_0, i_10_75_1314_0, i_10_75_1445_0,
    i_10_75_1485_0, i_10_75_1549_0, i_10_75_1550_0, i_10_75_1559_0,
    i_10_75_1798_0, i_10_75_1823_0, i_10_75_1854_0, i_10_75_1876_0,
    i_10_75_2036_0, i_10_75_2198_0, i_10_75_2324_0, i_10_75_2350_0,
    i_10_75_2351_0, i_10_75_2353_0, i_10_75_2448_0, i_10_75_2449_0,
    i_10_75_2450_0, i_10_75_2453_0, i_10_75_2474_0, i_10_75_2475_0,
    i_10_75_2530_0, i_10_75_2531_0, i_10_75_2532_0, i_10_75_2569_0,
    i_10_75_2603_0, i_10_75_2674_0, i_10_75_2707_0, i_10_75_2710_0,
    i_10_75_2713_0, i_10_75_2727_0, i_10_75_2804_0, i_10_75_2818_0,
    i_10_75_2888_0, i_10_75_2909_0, i_10_75_2980_0, i_10_75_2983_0,
    i_10_75_2984_0, i_10_75_2989_0, i_10_75_2992_0, i_10_75_3076_0,
    i_10_75_3077_0, i_10_75_3198_0, i_10_75_3206_0, i_10_75_3277_0,
    i_10_75_3278_0, i_10_75_3303_0, i_10_75_3333_0, i_10_75_3462_0,
    i_10_75_3468_0, i_10_75_3469_0, i_10_75_3470_0, i_10_75_3501_0,
    i_10_75_3503_0, i_10_75_3522_0, i_10_75_3523_0, i_10_75_3524_0,
    i_10_75_3541_0, i_10_75_3613_0, i_10_75_3649_0, i_10_75_3774_0,
    i_10_75_3783_0, i_10_75_3853_0, i_10_75_3854_0, i_10_75_3857_0,
    i_10_75_3859_0, i_10_75_3860_0, i_10_75_3911_0, i_10_75_3926_0,
    i_10_75_4005_0, i_10_75_4214_0, i_10_75_4249_0, i_10_75_4277_0,
    i_10_75_4291_0, i_10_75_4457_0, i_10_75_4559_0,
    o_10_75_0_0  );
  input  i_10_75_38_0, i_10_75_49_0, i_10_75_66_0, i_10_75_69_0,
    i_10_75_155_0, i_10_75_191_0, i_10_75_194_0, i_10_75_218_0,
    i_10_75_237_0, i_10_75_246_0, i_10_75_425_0, i_10_75_442_0,
    i_10_75_460_0, i_10_75_595_0, i_10_75_621_0, i_10_75_794_0,
    i_10_75_958_0, i_10_75_995_0, i_10_75_1026_0, i_10_75_1245_0,
    i_10_75_1246_0, i_10_75_1299_0, i_10_75_1310_0, i_10_75_1314_0,
    i_10_75_1445_0, i_10_75_1485_0, i_10_75_1549_0, i_10_75_1550_0,
    i_10_75_1559_0, i_10_75_1798_0, i_10_75_1823_0, i_10_75_1854_0,
    i_10_75_1876_0, i_10_75_2036_0, i_10_75_2198_0, i_10_75_2324_0,
    i_10_75_2350_0, i_10_75_2351_0, i_10_75_2353_0, i_10_75_2448_0,
    i_10_75_2449_0, i_10_75_2450_0, i_10_75_2453_0, i_10_75_2474_0,
    i_10_75_2475_0, i_10_75_2530_0, i_10_75_2531_0, i_10_75_2532_0,
    i_10_75_2569_0, i_10_75_2603_0, i_10_75_2674_0, i_10_75_2707_0,
    i_10_75_2710_0, i_10_75_2713_0, i_10_75_2727_0, i_10_75_2804_0,
    i_10_75_2818_0, i_10_75_2888_0, i_10_75_2909_0, i_10_75_2980_0,
    i_10_75_2983_0, i_10_75_2984_0, i_10_75_2989_0, i_10_75_2992_0,
    i_10_75_3076_0, i_10_75_3077_0, i_10_75_3198_0, i_10_75_3206_0,
    i_10_75_3277_0, i_10_75_3278_0, i_10_75_3303_0, i_10_75_3333_0,
    i_10_75_3462_0, i_10_75_3468_0, i_10_75_3469_0, i_10_75_3470_0,
    i_10_75_3501_0, i_10_75_3503_0, i_10_75_3522_0, i_10_75_3523_0,
    i_10_75_3524_0, i_10_75_3541_0, i_10_75_3613_0, i_10_75_3649_0,
    i_10_75_3774_0, i_10_75_3783_0, i_10_75_3853_0, i_10_75_3854_0,
    i_10_75_3857_0, i_10_75_3859_0, i_10_75_3860_0, i_10_75_3911_0,
    i_10_75_3926_0, i_10_75_4005_0, i_10_75_4214_0, i_10_75_4249_0,
    i_10_75_4277_0, i_10_75_4291_0, i_10_75_4457_0, i_10_75_4559_0;
  output o_10_75_0_0;
  assign o_10_75_0_0 = 0;
endmodule



// Benchmark "kernel_10_76" written by ABC on Sun Jul 19 10:22:19 2020

module kernel_10_76 ( 
    i_10_76_40_0, i_10_76_174_0, i_10_76_175_0, i_10_76_178_0,
    i_10_76_244_0, i_10_76_284_0, i_10_76_285_0, i_10_76_316_0,
    i_10_76_317_0, i_10_76_395_0, i_10_76_405_0, i_10_76_406_0,
    i_10_76_410_0, i_10_76_438_0, i_10_76_447_0, i_10_76_448_0,
    i_10_76_449_0, i_10_76_463_0, i_10_76_464_0, i_10_76_533_0,
    i_10_76_626_0, i_10_76_718_0, i_10_76_719_0, i_10_76_752_0,
    i_10_76_755_0, i_10_76_958_0, i_10_76_959_0, i_10_76_969_0,
    i_10_76_990_0, i_10_76_991_0, i_10_76_994_0, i_10_76_1051_0,
    i_10_76_1123_0, i_10_76_1233_0, i_10_76_1238_0, i_10_76_1344_0,
    i_10_76_1433_0, i_10_76_1445_0, i_10_76_1539_0, i_10_76_1546_0,
    i_10_76_1621_0, i_10_76_1622_0, i_10_76_1626_0, i_10_76_1635_0,
    i_10_76_1652_0, i_10_76_1685_0, i_10_76_1766_0, i_10_76_1825_0,
    i_10_76_2003_0, i_10_76_2019_0, i_10_76_2164_0, i_10_76_2355_0,
    i_10_76_2356_0, i_10_76_2359_0, i_10_76_2362_0, i_10_76_2514_0,
    i_10_76_2539_0, i_10_76_2562_0, i_10_76_2563_0, i_10_76_2570_0,
    i_10_76_2604_0, i_10_76_2632_0, i_10_76_2676_0, i_10_76_2706_0,
    i_10_76_2733_0, i_10_76_2734_0, i_10_76_2781_0, i_10_76_2866_0,
    i_10_76_2884_0, i_10_76_3046_0, i_10_76_3069_0, i_10_76_3070_0,
    i_10_76_3072_0, i_10_76_3073_0, i_10_76_3074_0, i_10_76_3279_0,
    i_10_76_3283_0, i_10_76_3284_0, i_10_76_3387_0, i_10_76_3540_0,
    i_10_76_3583_0, i_10_76_3648_0, i_10_76_3651_0, i_10_76_3811_0,
    i_10_76_3812_0, i_10_76_3840_0, i_10_76_3987_0, i_10_76_3988_0,
    i_10_76_4114_0, i_10_76_4115_0, i_10_76_4121_0, i_10_76_4129_0,
    i_10_76_4150_0, i_10_76_4151_0, i_10_76_4172_0, i_10_76_4174_0,
    i_10_76_4216_0, i_10_76_4276_0, i_10_76_4279_0, i_10_76_4571_0,
    o_10_76_0_0  );
  input  i_10_76_40_0, i_10_76_174_0, i_10_76_175_0, i_10_76_178_0,
    i_10_76_244_0, i_10_76_284_0, i_10_76_285_0, i_10_76_316_0,
    i_10_76_317_0, i_10_76_395_0, i_10_76_405_0, i_10_76_406_0,
    i_10_76_410_0, i_10_76_438_0, i_10_76_447_0, i_10_76_448_0,
    i_10_76_449_0, i_10_76_463_0, i_10_76_464_0, i_10_76_533_0,
    i_10_76_626_0, i_10_76_718_0, i_10_76_719_0, i_10_76_752_0,
    i_10_76_755_0, i_10_76_958_0, i_10_76_959_0, i_10_76_969_0,
    i_10_76_990_0, i_10_76_991_0, i_10_76_994_0, i_10_76_1051_0,
    i_10_76_1123_0, i_10_76_1233_0, i_10_76_1238_0, i_10_76_1344_0,
    i_10_76_1433_0, i_10_76_1445_0, i_10_76_1539_0, i_10_76_1546_0,
    i_10_76_1621_0, i_10_76_1622_0, i_10_76_1626_0, i_10_76_1635_0,
    i_10_76_1652_0, i_10_76_1685_0, i_10_76_1766_0, i_10_76_1825_0,
    i_10_76_2003_0, i_10_76_2019_0, i_10_76_2164_0, i_10_76_2355_0,
    i_10_76_2356_0, i_10_76_2359_0, i_10_76_2362_0, i_10_76_2514_0,
    i_10_76_2539_0, i_10_76_2562_0, i_10_76_2563_0, i_10_76_2570_0,
    i_10_76_2604_0, i_10_76_2632_0, i_10_76_2676_0, i_10_76_2706_0,
    i_10_76_2733_0, i_10_76_2734_0, i_10_76_2781_0, i_10_76_2866_0,
    i_10_76_2884_0, i_10_76_3046_0, i_10_76_3069_0, i_10_76_3070_0,
    i_10_76_3072_0, i_10_76_3073_0, i_10_76_3074_0, i_10_76_3279_0,
    i_10_76_3283_0, i_10_76_3284_0, i_10_76_3387_0, i_10_76_3540_0,
    i_10_76_3583_0, i_10_76_3648_0, i_10_76_3651_0, i_10_76_3811_0,
    i_10_76_3812_0, i_10_76_3840_0, i_10_76_3987_0, i_10_76_3988_0,
    i_10_76_4114_0, i_10_76_4115_0, i_10_76_4121_0, i_10_76_4129_0,
    i_10_76_4150_0, i_10_76_4151_0, i_10_76_4172_0, i_10_76_4174_0,
    i_10_76_4216_0, i_10_76_4276_0, i_10_76_4279_0, i_10_76_4571_0;
  output o_10_76_0_0;
  assign o_10_76_0_0 = 0;
endmodule



// Benchmark "kernel_10_77" written by ABC on Sun Jul 19 10:22:19 2020

module kernel_10_77 ( 
    i_10_77_71_0, i_10_77_83_0, i_10_77_217_0, i_10_77_254_0,
    i_10_77_277_0, i_10_77_320_0, i_10_77_322_0, i_10_77_388_0,
    i_10_77_409_0, i_10_77_423_0, i_10_77_424_0, i_10_77_425_0,
    i_10_77_427_0, i_10_77_428_0, i_10_77_434_0, i_10_77_532_0,
    i_10_77_693_0, i_10_77_904_0, i_10_77_991_0, i_10_77_1028_0,
    i_10_77_1033_0, i_10_77_1040_0, i_10_77_1043_0, i_10_77_1117_0,
    i_10_77_1171_0, i_10_77_1197_0, i_10_77_1308_0, i_10_77_1399_0,
    i_10_77_1400_0, i_10_77_1577_0, i_10_77_1733_0, i_10_77_1741_0,
    i_10_77_1766_0, i_10_77_1768_0, i_10_77_1822_0, i_10_77_1910_0,
    i_10_77_1944_0, i_10_77_1948_0, i_10_77_1985_0, i_10_77_1991_0,
    i_10_77_1993_0, i_10_77_2023_0, i_10_77_2377_0, i_10_77_2383_0,
    i_10_77_2454_0, i_10_77_2455_0, i_10_77_2458_0, i_10_77_2476_0,
    i_10_77_2557_0, i_10_77_2558_0, i_10_77_2560_0, i_10_77_2569_0,
    i_10_77_2635_0, i_10_77_2647_0, i_10_77_2648_0, i_10_77_2650_0,
    i_10_77_2658_0, i_10_77_2659_0, i_10_77_2711_0, i_10_77_2714_0,
    i_10_77_2720_0, i_10_77_2721_0, i_10_77_2722_0, i_10_77_2881_0,
    i_10_77_2885_0, i_10_77_2923_0, i_10_77_3071_0, i_10_77_3088_0,
    i_10_77_3092_0, i_10_77_3195_0, i_10_77_3203_0, i_10_77_3278_0,
    i_10_77_3353_0, i_10_77_3385_0, i_10_77_3386_0, i_10_77_3387_0,
    i_10_77_3389_0, i_10_77_3405_0, i_10_77_3440_0, i_10_77_3547_0,
    i_10_77_3548_0, i_10_77_3550_0, i_10_77_3610_0, i_10_77_3611_0,
    i_10_77_3834_0, i_10_77_3841_0, i_10_77_3855_0, i_10_77_3856_0,
    i_10_77_3979_0, i_10_77_3989_0, i_10_77_4024_0, i_10_77_4025_0,
    i_10_77_4027_0, i_10_77_4029_0, i_10_77_4030_0, i_10_77_4128_0,
    i_10_77_4171_0, i_10_77_4456_0, i_10_77_4578_0, i_10_77_4590_0,
    o_10_77_0_0  );
  input  i_10_77_71_0, i_10_77_83_0, i_10_77_217_0, i_10_77_254_0,
    i_10_77_277_0, i_10_77_320_0, i_10_77_322_0, i_10_77_388_0,
    i_10_77_409_0, i_10_77_423_0, i_10_77_424_0, i_10_77_425_0,
    i_10_77_427_0, i_10_77_428_0, i_10_77_434_0, i_10_77_532_0,
    i_10_77_693_0, i_10_77_904_0, i_10_77_991_0, i_10_77_1028_0,
    i_10_77_1033_0, i_10_77_1040_0, i_10_77_1043_0, i_10_77_1117_0,
    i_10_77_1171_0, i_10_77_1197_0, i_10_77_1308_0, i_10_77_1399_0,
    i_10_77_1400_0, i_10_77_1577_0, i_10_77_1733_0, i_10_77_1741_0,
    i_10_77_1766_0, i_10_77_1768_0, i_10_77_1822_0, i_10_77_1910_0,
    i_10_77_1944_0, i_10_77_1948_0, i_10_77_1985_0, i_10_77_1991_0,
    i_10_77_1993_0, i_10_77_2023_0, i_10_77_2377_0, i_10_77_2383_0,
    i_10_77_2454_0, i_10_77_2455_0, i_10_77_2458_0, i_10_77_2476_0,
    i_10_77_2557_0, i_10_77_2558_0, i_10_77_2560_0, i_10_77_2569_0,
    i_10_77_2635_0, i_10_77_2647_0, i_10_77_2648_0, i_10_77_2650_0,
    i_10_77_2658_0, i_10_77_2659_0, i_10_77_2711_0, i_10_77_2714_0,
    i_10_77_2720_0, i_10_77_2721_0, i_10_77_2722_0, i_10_77_2881_0,
    i_10_77_2885_0, i_10_77_2923_0, i_10_77_3071_0, i_10_77_3088_0,
    i_10_77_3092_0, i_10_77_3195_0, i_10_77_3203_0, i_10_77_3278_0,
    i_10_77_3353_0, i_10_77_3385_0, i_10_77_3386_0, i_10_77_3387_0,
    i_10_77_3389_0, i_10_77_3405_0, i_10_77_3440_0, i_10_77_3547_0,
    i_10_77_3548_0, i_10_77_3550_0, i_10_77_3610_0, i_10_77_3611_0,
    i_10_77_3834_0, i_10_77_3841_0, i_10_77_3855_0, i_10_77_3856_0,
    i_10_77_3979_0, i_10_77_3989_0, i_10_77_4024_0, i_10_77_4025_0,
    i_10_77_4027_0, i_10_77_4029_0, i_10_77_4030_0, i_10_77_4128_0,
    i_10_77_4171_0, i_10_77_4456_0, i_10_77_4578_0, i_10_77_4590_0;
  output o_10_77_0_0;
  assign o_10_77_0_0 = 0;
endmodule



// Benchmark "kernel_10_78" written by ABC on Sun Jul 19 10:22:20 2020

module kernel_10_78 ( 
    i_10_78_15_0, i_10_78_117_0, i_10_78_118_0, i_10_78_121_0,
    i_10_78_140_0, i_10_78_265_0, i_10_78_282_0, i_10_78_328_0,
    i_10_78_449_0, i_10_78_513_0, i_10_78_562_0, i_10_78_634_0,
    i_10_78_718_0, i_10_78_930_0, i_10_78_958_0, i_10_78_959_0,
    i_10_78_963_0, i_10_78_1033_0, i_10_78_1162_0, i_10_78_1163_0,
    i_10_78_1206_0, i_10_78_1239_0, i_10_78_1362_0, i_10_78_1380_0,
    i_10_78_1451_0, i_10_78_1533_0, i_10_78_1634_0, i_10_78_1642_0,
    i_10_78_1654_0, i_10_78_1686_0, i_10_78_1687_0, i_10_78_1688_0,
    i_10_78_1722_0, i_10_78_1723_0, i_10_78_1724_0, i_10_78_1729_0,
    i_10_78_1730_0, i_10_78_1795_0, i_10_78_1821_0, i_10_78_1914_0,
    i_10_78_1948_0, i_10_78_2057_0, i_10_78_2065_0, i_10_78_2066_0,
    i_10_78_2241_0, i_10_78_2244_0, i_10_78_2349_0, i_10_78_2350_0,
    i_10_78_2365_0, i_10_78_2390_0, i_10_78_2468_0, i_10_78_2469_0,
    i_10_78_2517_0, i_10_78_2541_0, i_10_78_2542_0, i_10_78_2544_0,
    i_10_78_2607_0, i_10_78_2608_0, i_10_78_2614_0, i_10_78_2615_0,
    i_10_78_2666_0, i_10_78_2715_0, i_10_78_2721_0, i_10_78_2722_0,
    i_10_78_2741_0, i_10_78_2995_0, i_10_78_3035_0, i_10_78_3036_0,
    i_10_78_3070_0, i_10_78_3390_0, i_10_78_3391_0, i_10_78_3392_0,
    i_10_78_3449_0, i_10_78_3451_0, i_10_78_3492_0, i_10_78_3493_0,
    i_10_78_3496_0, i_10_78_3525_0, i_10_78_3541_0, i_10_78_3544_0,
    i_10_78_3613_0, i_10_78_3648_0, i_10_78_3652_0, i_10_78_3719_0,
    i_10_78_3777_0, i_10_78_3853_0, i_10_78_3854_0, i_10_78_3878_0,
    i_10_78_3913_0, i_10_78_3983_0, i_10_78_4114_0, i_10_78_4115_0,
    i_10_78_4116_0, i_10_78_4129_0, i_10_78_4131_0, i_10_78_4290_0,
    i_10_78_4450_0, i_10_78_4458_0, i_10_78_4459_0, i_10_78_4531_0,
    o_10_78_0_0  );
  input  i_10_78_15_0, i_10_78_117_0, i_10_78_118_0, i_10_78_121_0,
    i_10_78_140_0, i_10_78_265_0, i_10_78_282_0, i_10_78_328_0,
    i_10_78_449_0, i_10_78_513_0, i_10_78_562_0, i_10_78_634_0,
    i_10_78_718_0, i_10_78_930_0, i_10_78_958_0, i_10_78_959_0,
    i_10_78_963_0, i_10_78_1033_0, i_10_78_1162_0, i_10_78_1163_0,
    i_10_78_1206_0, i_10_78_1239_0, i_10_78_1362_0, i_10_78_1380_0,
    i_10_78_1451_0, i_10_78_1533_0, i_10_78_1634_0, i_10_78_1642_0,
    i_10_78_1654_0, i_10_78_1686_0, i_10_78_1687_0, i_10_78_1688_0,
    i_10_78_1722_0, i_10_78_1723_0, i_10_78_1724_0, i_10_78_1729_0,
    i_10_78_1730_0, i_10_78_1795_0, i_10_78_1821_0, i_10_78_1914_0,
    i_10_78_1948_0, i_10_78_2057_0, i_10_78_2065_0, i_10_78_2066_0,
    i_10_78_2241_0, i_10_78_2244_0, i_10_78_2349_0, i_10_78_2350_0,
    i_10_78_2365_0, i_10_78_2390_0, i_10_78_2468_0, i_10_78_2469_0,
    i_10_78_2517_0, i_10_78_2541_0, i_10_78_2542_0, i_10_78_2544_0,
    i_10_78_2607_0, i_10_78_2608_0, i_10_78_2614_0, i_10_78_2615_0,
    i_10_78_2666_0, i_10_78_2715_0, i_10_78_2721_0, i_10_78_2722_0,
    i_10_78_2741_0, i_10_78_2995_0, i_10_78_3035_0, i_10_78_3036_0,
    i_10_78_3070_0, i_10_78_3390_0, i_10_78_3391_0, i_10_78_3392_0,
    i_10_78_3449_0, i_10_78_3451_0, i_10_78_3492_0, i_10_78_3493_0,
    i_10_78_3496_0, i_10_78_3525_0, i_10_78_3541_0, i_10_78_3544_0,
    i_10_78_3613_0, i_10_78_3648_0, i_10_78_3652_0, i_10_78_3719_0,
    i_10_78_3777_0, i_10_78_3853_0, i_10_78_3854_0, i_10_78_3878_0,
    i_10_78_3913_0, i_10_78_3983_0, i_10_78_4114_0, i_10_78_4115_0,
    i_10_78_4116_0, i_10_78_4129_0, i_10_78_4131_0, i_10_78_4290_0,
    i_10_78_4450_0, i_10_78_4458_0, i_10_78_4459_0, i_10_78_4531_0;
  output o_10_78_0_0;
  assign o_10_78_0_0 = 0;
endmodule



// Benchmark "kernel_10_79" written by ABC on Sun Jul 19 10:22:21 2020

module kernel_10_79 ( 
    i_10_79_175_0, i_10_79_187_0, i_10_79_246_0, i_10_79_249_0,
    i_10_79_265_0, i_10_79_283_0, i_10_79_411_0, i_10_79_412_0,
    i_10_79_430_0, i_10_79_431_0, i_10_79_440_0, i_10_79_444_0,
    i_10_79_446_0, i_10_79_457_0, i_10_79_509_0, i_10_79_518_0,
    i_10_79_521_0, i_10_79_797_0, i_10_79_956_0, i_10_79_957_0,
    i_10_79_958_0, i_10_79_959_0, i_10_79_967_0, i_10_79_997_0,
    i_10_79_1006_0, i_10_79_1007_0, i_10_79_1052_0, i_10_79_1138_0,
    i_10_79_1140_0, i_10_79_1247_0, i_10_79_1248_0, i_10_79_1493_0,
    i_10_79_1555_0, i_10_79_1556_0, i_10_79_1653_0, i_10_79_1691_0,
    i_10_79_1823_0, i_10_79_1913_0, i_10_79_1987_0, i_10_79_2005_0,
    i_10_79_2006_0, i_10_79_2350_0, i_10_79_2353_0, i_10_79_2364_0,
    i_10_79_2452_0, i_10_79_2474_0, i_10_79_2509_0, i_10_79_2607_0,
    i_10_79_2656_0, i_10_79_2662_0, i_10_79_2681_0, i_10_79_2706_0,
    i_10_79_2716_0, i_10_79_2717_0, i_10_79_2721_0, i_10_79_2732_0,
    i_10_79_2734_0, i_10_79_2735_0, i_10_79_2852_0, i_10_79_2880_0,
    i_10_79_2884_0, i_10_79_2885_0, i_10_79_2887_0, i_10_79_2922_0,
    i_10_79_3039_0, i_10_79_3093_0, i_10_79_3094_0, i_10_79_3095_0,
    i_10_79_3281_0, i_10_79_3355_0, i_10_79_3387_0, i_10_79_3388_0,
    i_10_79_3389_0, i_10_79_3406_0, i_10_79_3409_0, i_10_79_3472_0,
    i_10_79_3473_0, i_10_79_3497_0, i_10_79_3585_0, i_10_79_3587_0,
    i_10_79_3613_0, i_10_79_3646_0, i_10_79_3648_0, i_10_79_3649_0,
    i_10_79_3651_0, i_10_79_3784_0, i_10_79_3785_0, i_10_79_3786_0,
    i_10_79_3787_0, i_10_79_3788_0, i_10_79_3836_0, i_10_79_3847_0,
    i_10_79_3850_0, i_10_79_3851_0, i_10_79_3913_0, i_10_79_3914_0,
    i_10_79_3983_0, i_10_79_3986_0, i_10_79_4116_0, i_10_79_4117_0,
    o_10_79_0_0  );
  input  i_10_79_175_0, i_10_79_187_0, i_10_79_246_0, i_10_79_249_0,
    i_10_79_265_0, i_10_79_283_0, i_10_79_411_0, i_10_79_412_0,
    i_10_79_430_0, i_10_79_431_0, i_10_79_440_0, i_10_79_444_0,
    i_10_79_446_0, i_10_79_457_0, i_10_79_509_0, i_10_79_518_0,
    i_10_79_521_0, i_10_79_797_0, i_10_79_956_0, i_10_79_957_0,
    i_10_79_958_0, i_10_79_959_0, i_10_79_967_0, i_10_79_997_0,
    i_10_79_1006_0, i_10_79_1007_0, i_10_79_1052_0, i_10_79_1138_0,
    i_10_79_1140_0, i_10_79_1247_0, i_10_79_1248_0, i_10_79_1493_0,
    i_10_79_1555_0, i_10_79_1556_0, i_10_79_1653_0, i_10_79_1691_0,
    i_10_79_1823_0, i_10_79_1913_0, i_10_79_1987_0, i_10_79_2005_0,
    i_10_79_2006_0, i_10_79_2350_0, i_10_79_2353_0, i_10_79_2364_0,
    i_10_79_2452_0, i_10_79_2474_0, i_10_79_2509_0, i_10_79_2607_0,
    i_10_79_2656_0, i_10_79_2662_0, i_10_79_2681_0, i_10_79_2706_0,
    i_10_79_2716_0, i_10_79_2717_0, i_10_79_2721_0, i_10_79_2732_0,
    i_10_79_2734_0, i_10_79_2735_0, i_10_79_2852_0, i_10_79_2880_0,
    i_10_79_2884_0, i_10_79_2885_0, i_10_79_2887_0, i_10_79_2922_0,
    i_10_79_3039_0, i_10_79_3093_0, i_10_79_3094_0, i_10_79_3095_0,
    i_10_79_3281_0, i_10_79_3355_0, i_10_79_3387_0, i_10_79_3388_0,
    i_10_79_3389_0, i_10_79_3406_0, i_10_79_3409_0, i_10_79_3472_0,
    i_10_79_3473_0, i_10_79_3497_0, i_10_79_3585_0, i_10_79_3587_0,
    i_10_79_3613_0, i_10_79_3646_0, i_10_79_3648_0, i_10_79_3649_0,
    i_10_79_3651_0, i_10_79_3784_0, i_10_79_3785_0, i_10_79_3786_0,
    i_10_79_3787_0, i_10_79_3788_0, i_10_79_3836_0, i_10_79_3847_0,
    i_10_79_3850_0, i_10_79_3851_0, i_10_79_3913_0, i_10_79_3914_0,
    i_10_79_3983_0, i_10_79_3986_0, i_10_79_4116_0, i_10_79_4117_0;
  output o_10_79_0_0;
  assign o_10_79_0_0 = ~((~i_10_79_3281_0 & ((~i_10_79_175_0 & ((~i_10_79_2452_0 & ~i_10_79_2656_0 & ~i_10_79_2735_0 & ~i_10_79_3094_0 & i_10_79_3387_0 & i_10_79_3388_0 & ~i_10_79_3473_0) | (~i_10_79_457_0 & ~i_10_79_518_0 & ~i_10_79_1007_0 & ~i_10_79_2662_0 & ~i_10_79_3093_0 & ~i_10_79_3406_0 & ~i_10_79_3913_0))) | (i_10_79_249_0 & ~i_10_79_446_0 & ~i_10_79_1493_0 & ~i_10_79_2656_0) | (~i_10_79_431_0 & ~i_10_79_440_0 & ~i_10_79_2452_0 & ~i_10_79_3409_0 & ~i_10_79_3472_0 & ~i_10_79_3473_0 & ~i_10_79_3497_0))) | (i_10_79_430_0 & ((~i_10_79_521_0 & ~i_10_79_958_0 & ~i_10_79_1007_0 & ~i_10_79_2681_0 & ~i_10_79_2734_0 & ~i_10_79_3388_0 & ~i_10_79_3409_0) | (i_10_79_1248_0 & ~i_10_79_1555_0 & ~i_10_79_2474_0 & ~i_10_79_3094_0 & ~i_10_79_3613_0 & ~i_10_79_3913_0))) | (~i_10_79_2717_0 & ((~i_10_79_430_0 & ((~i_10_79_1006_0 & ~i_10_79_2735_0 & i_10_79_2884_0 & ~i_10_79_3389_0 & ~i_10_79_3983_0) | (~i_10_79_1556_0 & ~i_10_79_2681_0 & ~i_10_79_2884_0 & ~i_10_79_3986_0))) | (~i_10_79_2681_0 & ((~i_10_79_1493_0 & ~i_10_79_1653_0 & ~i_10_79_2474_0 & ~i_10_79_2716_0 & ~i_10_79_2735_0 & ~i_10_79_3497_0 & ~i_10_79_3613_0) | (~i_10_79_431_0 & ~i_10_79_797_0 & ~i_10_79_1555_0 & ~i_10_79_2005_0 & ~i_10_79_2006_0 & ~i_10_79_2922_0 & ~i_10_79_3406_0 & ~i_10_79_3914_0))) | (~i_10_79_440_0 & ~i_10_79_2735_0 & ~i_10_79_2884_0 & i_10_79_2922_0 & ~i_10_79_3983_0))) | (~i_10_79_2880_0 & ((~i_10_79_440_0 & ((~i_10_79_265_0 & ~i_10_79_2006_0 & ~i_10_79_3473_0 & i_10_79_3649_0) | (~i_10_79_444_0 & ~i_10_79_1555_0 & ~i_10_79_1823_0 & ~i_10_79_2474_0 & ~i_10_79_3094_0 & ~i_10_79_3472_0 & ~i_10_79_3986_0))) | (~i_10_79_457_0 & ~i_10_79_959_0 & ~i_10_79_967_0 & ~i_10_79_1006_0 & ~i_10_79_1493_0 & ~i_10_79_1556_0 & ~i_10_79_2006_0 & ~i_10_79_2350_0 & ~i_10_79_3094_0 & ~i_10_79_3095_0 & ~i_10_79_3406_0 & ~i_10_79_3497_0 & ~i_10_79_3646_0 & ~i_10_79_3851_0 & ~i_10_79_3913_0 & ~i_10_79_3914_0))) | (~i_10_79_2716_0 & ((~i_10_79_1555_0 & i_10_79_3093_0 & ~i_10_79_3094_0 & ~i_10_79_3986_0) | (~i_10_79_1006_0 & ~i_10_79_1493_0 & ~i_10_79_1556_0 & ~i_10_79_2885_0 & ~i_10_79_2887_0 & ~i_10_79_3649_0 & ~i_10_79_3651_0 & ~i_10_79_3913_0 & ~i_10_79_4117_0))) | (~i_10_79_446_0 & ~i_10_79_457_0 & i_10_79_2364_0 & i_10_79_2656_0) | (~i_10_79_431_0 & ~i_10_79_956_0 & ~i_10_79_958_0 & ~i_10_79_1007_0 & ~i_10_79_1913_0 & ~i_10_79_2734_0 & ~i_10_79_2885_0 & ~i_10_79_2887_0 & ~i_10_79_3786_0 & ~i_10_79_3913_0));
endmodule



// Benchmark "kernel_10_80" written by ABC on Sun Jul 19 10:22:22 2020

module kernel_10_80 ( 
    i_10_80_52_0, i_10_80_224_0, i_10_80_293_0, i_10_80_319_0,
    i_10_80_425_0, i_10_80_427_0, i_10_80_464_0, i_10_80_694_0,
    i_10_80_793_0, i_10_80_845_0, i_10_80_849_0, i_10_80_927_0,
    i_10_80_1000_0, i_10_80_1037_0, i_10_80_1045_0, i_10_80_1118_0,
    i_10_80_1299_0, i_10_80_1341_0, i_10_80_1342_0, i_10_80_1343_0,
    i_10_80_1352_0, i_10_80_1438_0, i_10_80_1450_0, i_10_80_1549_0,
    i_10_80_1550_0, i_10_80_1553_0, i_10_80_1616_0, i_10_80_1652_0,
    i_10_80_1715_0, i_10_80_1728_0, i_10_80_1742_0, i_10_80_1766_0,
    i_10_80_1822_0, i_10_80_1873_0, i_10_80_1909_0, i_10_80_1910_0,
    i_10_80_1913_0, i_10_80_1946_0, i_10_80_2091_0, i_10_80_2183_0,
    i_10_80_2185_0, i_10_80_2186_0, i_10_80_2209_0, i_10_80_2305_0,
    i_10_80_2309_0, i_10_80_2312_0, i_10_80_2448_0, i_10_80_2450_0,
    i_10_80_2453_0, i_10_80_2464_0, i_10_80_2479_0, i_10_80_2480_0,
    i_10_80_2566_0, i_10_80_2640_0, i_10_80_2648_0, i_10_80_2663_0,
    i_10_80_2674_0, i_10_80_2677_0, i_10_80_2725_0, i_10_80_2740_0,
    i_10_80_2741_0, i_10_80_2831_0, i_10_80_2880_0, i_10_80_2881_0,
    i_10_80_2882_0, i_10_80_2918_0, i_10_80_2920_0, i_10_80_3052_0,
    i_10_80_3091_0, i_10_80_3201_0, i_10_80_3203_0, i_10_80_3268_0,
    i_10_80_3276_0, i_10_80_3277_0, i_10_80_3278_0, i_10_80_3350_0,
    i_10_80_3406_0, i_10_80_3410_0, i_10_80_3431_0, i_10_80_3602_0,
    i_10_80_3604_0, i_10_80_3704_0, i_10_80_3796_0, i_10_80_3828_0,
    i_10_80_3889_0, i_10_80_3901_0, i_10_80_3902_0, i_10_80_3979_0,
    i_10_80_3980_0, i_10_80_3983_0, i_10_80_4029_0, i_10_80_4099_0,
    i_10_80_4115_0, i_10_80_4124_0, i_10_80_4127_0, i_10_80_4175_0,
    i_10_80_4270_0, i_10_80_4564_0, i_10_80_4591_0, i_10_80_4594_0,
    o_10_80_0_0  );
  input  i_10_80_52_0, i_10_80_224_0, i_10_80_293_0, i_10_80_319_0,
    i_10_80_425_0, i_10_80_427_0, i_10_80_464_0, i_10_80_694_0,
    i_10_80_793_0, i_10_80_845_0, i_10_80_849_0, i_10_80_927_0,
    i_10_80_1000_0, i_10_80_1037_0, i_10_80_1045_0, i_10_80_1118_0,
    i_10_80_1299_0, i_10_80_1341_0, i_10_80_1342_0, i_10_80_1343_0,
    i_10_80_1352_0, i_10_80_1438_0, i_10_80_1450_0, i_10_80_1549_0,
    i_10_80_1550_0, i_10_80_1553_0, i_10_80_1616_0, i_10_80_1652_0,
    i_10_80_1715_0, i_10_80_1728_0, i_10_80_1742_0, i_10_80_1766_0,
    i_10_80_1822_0, i_10_80_1873_0, i_10_80_1909_0, i_10_80_1910_0,
    i_10_80_1913_0, i_10_80_1946_0, i_10_80_2091_0, i_10_80_2183_0,
    i_10_80_2185_0, i_10_80_2186_0, i_10_80_2209_0, i_10_80_2305_0,
    i_10_80_2309_0, i_10_80_2312_0, i_10_80_2448_0, i_10_80_2450_0,
    i_10_80_2453_0, i_10_80_2464_0, i_10_80_2479_0, i_10_80_2480_0,
    i_10_80_2566_0, i_10_80_2640_0, i_10_80_2648_0, i_10_80_2663_0,
    i_10_80_2674_0, i_10_80_2677_0, i_10_80_2725_0, i_10_80_2740_0,
    i_10_80_2741_0, i_10_80_2831_0, i_10_80_2880_0, i_10_80_2881_0,
    i_10_80_2882_0, i_10_80_2918_0, i_10_80_2920_0, i_10_80_3052_0,
    i_10_80_3091_0, i_10_80_3201_0, i_10_80_3203_0, i_10_80_3268_0,
    i_10_80_3276_0, i_10_80_3277_0, i_10_80_3278_0, i_10_80_3350_0,
    i_10_80_3406_0, i_10_80_3410_0, i_10_80_3431_0, i_10_80_3602_0,
    i_10_80_3604_0, i_10_80_3704_0, i_10_80_3796_0, i_10_80_3828_0,
    i_10_80_3889_0, i_10_80_3901_0, i_10_80_3902_0, i_10_80_3979_0,
    i_10_80_3980_0, i_10_80_3983_0, i_10_80_4029_0, i_10_80_4099_0,
    i_10_80_4115_0, i_10_80_4124_0, i_10_80_4127_0, i_10_80_4175_0,
    i_10_80_4270_0, i_10_80_4564_0, i_10_80_4591_0, i_10_80_4594_0;
  output o_10_80_0_0;
  assign o_10_80_0_0 = 0;
endmodule



// Benchmark "kernel_10_81" written by ABC on Sun Jul 19 10:22:23 2020

module kernel_10_81 ( 
    i_10_81_76_0, i_10_81_124_0, i_10_81_179_0, i_10_81_183_0,
    i_10_81_184_0, i_10_81_247_0, i_10_81_260_0, i_10_81_281_0,
    i_10_81_317_0, i_10_81_318_0, i_10_81_319_0, i_10_81_320_0,
    i_10_81_322_0, i_10_81_323_0, i_10_81_376_0, i_10_81_394_0,
    i_10_81_410_0, i_10_81_430_0, i_10_81_435_0, i_10_81_436_0,
    i_10_81_467_0, i_10_81_629_0, i_10_81_692_0, i_10_81_1032_0,
    i_10_81_1045_0, i_10_81_1083_0, i_10_81_1138_0, i_10_81_1158_0,
    i_10_81_1160_0, i_10_81_1166_0, i_10_81_1169_0, i_10_81_1240_0,
    i_10_81_1241_0, i_10_81_1268_0, i_10_81_1305_0, i_10_81_1312_0,
    i_10_81_1341_0, i_10_81_1366_0, i_10_81_1385_0, i_10_81_1542_0,
    i_10_81_1547_0, i_10_81_1713_0, i_10_81_1821_0, i_10_81_1851_0,
    i_10_81_1852_0, i_10_81_1879_0, i_10_81_1880_0, i_10_81_1912_0,
    i_10_81_1913_0, i_10_81_2059_0, i_10_81_2202_0, i_10_81_2203_0,
    i_10_81_2204_0, i_10_81_2355_0, i_10_81_2356_0, i_10_81_2380_0,
    i_10_81_2456_0, i_10_81_2542_0, i_10_81_2543_0, i_10_81_2580_0,
    i_10_81_2581_0, i_10_81_2582_0, i_10_81_2605_0, i_10_81_2608_0,
    i_10_81_2609_0, i_10_81_2636_0, i_10_81_2681_0, i_10_81_2705_0,
    i_10_81_2717_0, i_10_81_2725_0, i_10_81_2786_0, i_10_81_2834_0,
    i_10_81_2842_0, i_10_81_2884_0, i_10_81_2919_0, i_10_81_2986_0,
    i_10_81_2987_0, i_10_81_3072_0, i_10_81_3073_0, i_10_81_3198_0,
    i_10_81_3237_0, i_10_81_3283_0, i_10_81_3302_0, i_10_81_3391_0,
    i_10_81_3472_0, i_10_81_3589_0, i_10_81_3610_0, i_10_81_3911_0,
    i_10_81_3944_0, i_10_81_3948_0, i_10_81_3979_0, i_10_81_4028_0,
    i_10_81_4116_0, i_10_81_4117_0, i_10_81_4121_0, i_10_81_4126_0,
    i_10_81_4174_0, i_10_81_4281_0, i_10_81_4282_0, i_10_81_4288_0,
    o_10_81_0_0  );
  input  i_10_81_76_0, i_10_81_124_0, i_10_81_179_0, i_10_81_183_0,
    i_10_81_184_0, i_10_81_247_0, i_10_81_260_0, i_10_81_281_0,
    i_10_81_317_0, i_10_81_318_0, i_10_81_319_0, i_10_81_320_0,
    i_10_81_322_0, i_10_81_323_0, i_10_81_376_0, i_10_81_394_0,
    i_10_81_410_0, i_10_81_430_0, i_10_81_435_0, i_10_81_436_0,
    i_10_81_467_0, i_10_81_629_0, i_10_81_692_0, i_10_81_1032_0,
    i_10_81_1045_0, i_10_81_1083_0, i_10_81_1138_0, i_10_81_1158_0,
    i_10_81_1160_0, i_10_81_1166_0, i_10_81_1169_0, i_10_81_1240_0,
    i_10_81_1241_0, i_10_81_1268_0, i_10_81_1305_0, i_10_81_1312_0,
    i_10_81_1341_0, i_10_81_1366_0, i_10_81_1385_0, i_10_81_1542_0,
    i_10_81_1547_0, i_10_81_1713_0, i_10_81_1821_0, i_10_81_1851_0,
    i_10_81_1852_0, i_10_81_1879_0, i_10_81_1880_0, i_10_81_1912_0,
    i_10_81_1913_0, i_10_81_2059_0, i_10_81_2202_0, i_10_81_2203_0,
    i_10_81_2204_0, i_10_81_2355_0, i_10_81_2356_0, i_10_81_2380_0,
    i_10_81_2456_0, i_10_81_2542_0, i_10_81_2543_0, i_10_81_2580_0,
    i_10_81_2581_0, i_10_81_2582_0, i_10_81_2605_0, i_10_81_2608_0,
    i_10_81_2609_0, i_10_81_2636_0, i_10_81_2681_0, i_10_81_2705_0,
    i_10_81_2717_0, i_10_81_2725_0, i_10_81_2786_0, i_10_81_2834_0,
    i_10_81_2842_0, i_10_81_2884_0, i_10_81_2919_0, i_10_81_2986_0,
    i_10_81_2987_0, i_10_81_3072_0, i_10_81_3073_0, i_10_81_3198_0,
    i_10_81_3237_0, i_10_81_3283_0, i_10_81_3302_0, i_10_81_3391_0,
    i_10_81_3472_0, i_10_81_3589_0, i_10_81_3610_0, i_10_81_3911_0,
    i_10_81_3944_0, i_10_81_3948_0, i_10_81_3979_0, i_10_81_4028_0,
    i_10_81_4116_0, i_10_81_4117_0, i_10_81_4121_0, i_10_81_4126_0,
    i_10_81_4174_0, i_10_81_4281_0, i_10_81_4282_0, i_10_81_4288_0;
  output o_10_81_0_0;
  assign o_10_81_0_0 = 0;
endmodule



// Benchmark "kernel_10_82" written by ABC on Sun Jul 19 10:22:24 2020

module kernel_10_82 ( 
    i_10_82_244_0, i_10_82_247_0, i_10_82_265_0, i_10_82_279_0,
    i_10_82_316_0, i_10_82_320_0, i_10_82_406_0, i_10_82_460_0,
    i_10_82_467_0, i_10_82_755_0, i_10_82_820_0, i_10_82_960_0,
    i_10_82_997_0, i_10_82_1084_0, i_10_82_1236_0, i_10_82_1313_0,
    i_10_82_1345_0, i_10_82_1346_0, i_10_82_1348_0, i_10_82_1360_0,
    i_10_82_1543_0, i_10_82_1552_0, i_10_82_1580_0, i_10_82_1583_0,
    i_10_82_1630_0, i_10_82_1648_0, i_10_82_1649_0, i_10_82_1654_0,
    i_10_82_1655_0, i_10_82_1683_0, i_10_82_1713_0, i_10_82_1768_0,
    i_10_82_1800_0, i_10_82_1824_0, i_10_82_1825_0, i_10_82_1912_0,
    i_10_82_1988_0, i_10_82_2025_0, i_10_82_2182_0, i_10_82_2197_0,
    i_10_82_2198_0, i_10_82_2312_0, i_10_82_2361_0, i_10_82_2384_0,
    i_10_82_2457_0, i_10_82_2458_0, i_10_82_2468_0, i_10_82_2470_0,
    i_10_82_2565_0, i_10_82_2659_0, i_10_82_2660_0, i_10_82_2673_0,
    i_10_82_2701_0, i_10_82_2709_0, i_10_82_2710_0, i_10_82_2719_0,
    i_10_82_2720_0, i_10_82_2723_0, i_10_82_2729_0, i_10_82_2730_0,
    i_10_82_2735_0, i_10_82_2757_0, i_10_82_2882_0, i_10_82_2884_0,
    i_10_82_2887_0, i_10_82_2920_0, i_10_82_3046_0, i_10_82_3049_0,
    i_10_82_3268_0, i_10_82_3279_0, i_10_82_3280_0, i_10_82_3312_0,
    i_10_82_3325_0, i_10_82_3406_0, i_10_82_3407_0, i_10_82_3410_0,
    i_10_82_3541_0, i_10_82_3545_0, i_10_82_3585_0, i_10_82_3586_0,
    i_10_82_3610_0, i_10_82_3614_0, i_10_82_3650_0, i_10_82_3784_0,
    i_10_82_3808_0, i_10_82_3838_0, i_10_82_3847_0, i_10_82_3848_0,
    i_10_82_3854_0, i_10_82_3857_0, i_10_82_3994_0, i_10_82_4113_0,
    i_10_82_4116_0, i_10_82_4117_0, i_10_82_4118_0, i_10_82_4273_0,
    i_10_82_4285_0, i_10_82_4291_0, i_10_82_4568_0, i_10_82_4590_0,
    o_10_82_0_0  );
  input  i_10_82_244_0, i_10_82_247_0, i_10_82_265_0, i_10_82_279_0,
    i_10_82_316_0, i_10_82_320_0, i_10_82_406_0, i_10_82_460_0,
    i_10_82_467_0, i_10_82_755_0, i_10_82_820_0, i_10_82_960_0,
    i_10_82_997_0, i_10_82_1084_0, i_10_82_1236_0, i_10_82_1313_0,
    i_10_82_1345_0, i_10_82_1346_0, i_10_82_1348_0, i_10_82_1360_0,
    i_10_82_1543_0, i_10_82_1552_0, i_10_82_1580_0, i_10_82_1583_0,
    i_10_82_1630_0, i_10_82_1648_0, i_10_82_1649_0, i_10_82_1654_0,
    i_10_82_1655_0, i_10_82_1683_0, i_10_82_1713_0, i_10_82_1768_0,
    i_10_82_1800_0, i_10_82_1824_0, i_10_82_1825_0, i_10_82_1912_0,
    i_10_82_1988_0, i_10_82_2025_0, i_10_82_2182_0, i_10_82_2197_0,
    i_10_82_2198_0, i_10_82_2312_0, i_10_82_2361_0, i_10_82_2384_0,
    i_10_82_2457_0, i_10_82_2458_0, i_10_82_2468_0, i_10_82_2470_0,
    i_10_82_2565_0, i_10_82_2659_0, i_10_82_2660_0, i_10_82_2673_0,
    i_10_82_2701_0, i_10_82_2709_0, i_10_82_2710_0, i_10_82_2719_0,
    i_10_82_2720_0, i_10_82_2723_0, i_10_82_2729_0, i_10_82_2730_0,
    i_10_82_2735_0, i_10_82_2757_0, i_10_82_2882_0, i_10_82_2884_0,
    i_10_82_2887_0, i_10_82_2920_0, i_10_82_3046_0, i_10_82_3049_0,
    i_10_82_3268_0, i_10_82_3279_0, i_10_82_3280_0, i_10_82_3312_0,
    i_10_82_3325_0, i_10_82_3406_0, i_10_82_3407_0, i_10_82_3410_0,
    i_10_82_3541_0, i_10_82_3545_0, i_10_82_3585_0, i_10_82_3586_0,
    i_10_82_3610_0, i_10_82_3614_0, i_10_82_3650_0, i_10_82_3784_0,
    i_10_82_3808_0, i_10_82_3838_0, i_10_82_3847_0, i_10_82_3848_0,
    i_10_82_3854_0, i_10_82_3857_0, i_10_82_3994_0, i_10_82_4113_0,
    i_10_82_4116_0, i_10_82_4117_0, i_10_82_4118_0, i_10_82_4273_0,
    i_10_82_4285_0, i_10_82_4291_0, i_10_82_4568_0, i_10_82_4590_0;
  output o_10_82_0_0;
  assign o_10_82_0_0 = 0;
endmodule



// Benchmark "kernel_10_83" written by ABC on Sun Jul 19 10:22:24 2020

module kernel_10_83 ( 
    i_10_83_82_0, i_10_83_117_0, i_10_83_118_0, i_10_83_120_0,
    i_10_83_172_0, i_10_83_173_0, i_10_83_174_0, i_10_83_175_0,
    i_10_83_247_0, i_10_83_280_0, i_10_83_281_0, i_10_83_315_0,
    i_10_83_322_0, i_10_83_444_0, i_10_83_447_0, i_10_83_499_0,
    i_10_83_515_0, i_10_83_564_0, i_10_83_740_0, i_10_83_758_0,
    i_10_83_932_0, i_10_83_1238_0, i_10_83_1245_0, i_10_83_1306_0,
    i_10_83_1308_0, i_10_83_1311_0, i_10_83_1312_0, i_10_83_1361_0,
    i_10_83_1542_0, i_10_83_1611_0, i_10_83_1620_0, i_10_83_1648_0,
    i_10_83_1683_0, i_10_83_1821_0, i_10_83_1822_0, i_10_83_1918_0,
    i_10_83_1944_0, i_10_83_1945_0, i_10_83_1946_0, i_10_83_1947_0,
    i_10_83_1948_0, i_10_83_1951_0, i_10_83_1956_0, i_10_83_2023_0,
    i_10_83_2179_0, i_10_83_2243_0, i_10_83_2356_0, i_10_83_2380_0,
    i_10_83_2432_0, i_10_83_2460_0, i_10_83_2466_0, i_10_83_2511_0,
    i_10_83_2631_0, i_10_83_2635_0, i_10_83_2655_0, i_10_83_2656_0,
    i_10_83_2673_0, i_10_83_2674_0, i_10_83_2703_0, i_10_83_2711_0,
    i_10_83_2713_0, i_10_83_2716_0, i_10_83_2722_0, i_10_83_2727_0,
    i_10_83_2729_0, i_10_83_2819_0, i_10_83_2831_0, i_10_83_2885_0,
    i_10_83_2987_0, i_10_83_3036_0, i_10_83_3046_0, i_10_83_3089_0,
    i_10_83_3268_0, i_10_83_3278_0, i_10_83_3281_0, i_10_83_3284_0,
    i_10_83_3286_0, i_10_83_3296_0, i_10_83_3523_0, i_10_83_3524_0,
    i_10_83_3561_0, i_10_83_3614_0, i_10_83_3618_0, i_10_83_3649_0,
    i_10_83_3838_0, i_10_83_3854_0, i_10_83_3860_0, i_10_83_4023_0,
    i_10_83_4050_0, i_10_83_4117_0, i_10_83_4129_0, i_10_83_4174_0,
    i_10_83_4283_0, i_10_83_4286_0, i_10_83_4352_0, i_10_83_4460_0,
    i_10_83_4558_0, i_10_83_4559_0, i_10_83_4568_0, i_10_83_4569_0,
    o_10_83_0_0  );
  input  i_10_83_82_0, i_10_83_117_0, i_10_83_118_0, i_10_83_120_0,
    i_10_83_172_0, i_10_83_173_0, i_10_83_174_0, i_10_83_175_0,
    i_10_83_247_0, i_10_83_280_0, i_10_83_281_0, i_10_83_315_0,
    i_10_83_322_0, i_10_83_444_0, i_10_83_447_0, i_10_83_499_0,
    i_10_83_515_0, i_10_83_564_0, i_10_83_740_0, i_10_83_758_0,
    i_10_83_932_0, i_10_83_1238_0, i_10_83_1245_0, i_10_83_1306_0,
    i_10_83_1308_0, i_10_83_1311_0, i_10_83_1312_0, i_10_83_1361_0,
    i_10_83_1542_0, i_10_83_1611_0, i_10_83_1620_0, i_10_83_1648_0,
    i_10_83_1683_0, i_10_83_1821_0, i_10_83_1822_0, i_10_83_1918_0,
    i_10_83_1944_0, i_10_83_1945_0, i_10_83_1946_0, i_10_83_1947_0,
    i_10_83_1948_0, i_10_83_1951_0, i_10_83_1956_0, i_10_83_2023_0,
    i_10_83_2179_0, i_10_83_2243_0, i_10_83_2356_0, i_10_83_2380_0,
    i_10_83_2432_0, i_10_83_2460_0, i_10_83_2466_0, i_10_83_2511_0,
    i_10_83_2631_0, i_10_83_2635_0, i_10_83_2655_0, i_10_83_2656_0,
    i_10_83_2673_0, i_10_83_2674_0, i_10_83_2703_0, i_10_83_2711_0,
    i_10_83_2713_0, i_10_83_2716_0, i_10_83_2722_0, i_10_83_2727_0,
    i_10_83_2729_0, i_10_83_2819_0, i_10_83_2831_0, i_10_83_2885_0,
    i_10_83_2987_0, i_10_83_3036_0, i_10_83_3046_0, i_10_83_3089_0,
    i_10_83_3268_0, i_10_83_3278_0, i_10_83_3281_0, i_10_83_3284_0,
    i_10_83_3286_0, i_10_83_3296_0, i_10_83_3523_0, i_10_83_3524_0,
    i_10_83_3561_0, i_10_83_3614_0, i_10_83_3618_0, i_10_83_3649_0,
    i_10_83_3838_0, i_10_83_3854_0, i_10_83_3860_0, i_10_83_4023_0,
    i_10_83_4050_0, i_10_83_4117_0, i_10_83_4129_0, i_10_83_4174_0,
    i_10_83_4283_0, i_10_83_4286_0, i_10_83_4352_0, i_10_83_4460_0,
    i_10_83_4558_0, i_10_83_4559_0, i_10_83_4568_0, i_10_83_4569_0;
  output o_10_83_0_0;
  assign o_10_83_0_0 = 0;
endmodule



// Benchmark "kernel_10_84" written by ABC on Sun Jul 19 10:22:25 2020

module kernel_10_84 ( 
    i_10_84_221_0, i_10_84_240_0, i_10_84_283_0, i_10_84_296_0,
    i_10_84_413_0, i_10_84_438_0, i_10_84_445_0, i_10_84_446_0,
    i_10_84_465_0, i_10_84_466_0, i_10_84_799_0, i_10_84_827_0,
    i_10_84_897_0, i_10_84_993_0, i_10_84_996_0, i_10_84_1033_0,
    i_10_84_1034_0, i_10_84_1085_0, i_10_84_1153_0, i_10_84_1174_0,
    i_10_84_1175_0, i_10_84_1205_0, i_10_84_1233_0, i_10_84_1234_0,
    i_10_84_1238_0, i_10_84_1246_0, i_10_84_1247_0, i_10_84_1248_0,
    i_10_84_1308_0, i_10_84_1349_0, i_10_84_1363_0, i_10_84_1555_0,
    i_10_84_1556_0, i_10_84_1610_0, i_10_84_1627_0, i_10_84_1648_0,
    i_10_84_1687_0, i_10_84_1818_0, i_10_84_1819_0, i_10_84_1825_0,
    i_10_84_1950_0, i_10_84_2002_0, i_10_84_2003_0, i_10_84_2350_0,
    i_10_84_2351_0, i_10_84_2357_0, i_10_84_2364_0, i_10_84_2384_0,
    i_10_84_2411_0, i_10_84_2449_0, i_10_84_2465_0, i_10_84_2519_0,
    i_10_84_2540_0, i_10_84_2542_0, i_10_84_2543_0, i_10_84_2545_0,
    i_10_84_2572_0, i_10_84_2573_0, i_10_84_2634_0, i_10_84_2635_0,
    i_10_84_2708_0, i_10_84_2712_0, i_10_84_2730_0, i_10_84_2818_0,
    i_10_84_2830_0, i_10_84_2880_0, i_10_84_2887_0, i_10_84_2917_0,
    i_10_84_2918_0, i_10_84_2921_0, i_10_84_2922_0, i_10_84_2956_0,
    i_10_84_3039_0, i_10_84_3049_0, i_10_84_3090_0, i_10_84_3091_0,
    i_10_84_3162_0, i_10_84_3163_0, i_10_84_3277_0, i_10_84_3356_0,
    i_10_84_3390_0, i_10_84_3392_0, i_10_84_3446_0, i_10_84_3586_0,
    i_10_84_3613_0, i_10_84_3688_0, i_10_84_3689_0, i_10_84_3717_0,
    i_10_84_3734_0, i_10_84_3786_0, i_10_84_3850_0, i_10_84_3859_0,
    i_10_84_3892_0, i_10_84_4168_0, i_10_84_4267_0, i_10_84_4276_0,
    i_10_84_4277_0, i_10_84_4279_0, i_10_84_4568_0, i_10_84_4571_0,
    o_10_84_0_0  );
  input  i_10_84_221_0, i_10_84_240_0, i_10_84_283_0, i_10_84_296_0,
    i_10_84_413_0, i_10_84_438_0, i_10_84_445_0, i_10_84_446_0,
    i_10_84_465_0, i_10_84_466_0, i_10_84_799_0, i_10_84_827_0,
    i_10_84_897_0, i_10_84_993_0, i_10_84_996_0, i_10_84_1033_0,
    i_10_84_1034_0, i_10_84_1085_0, i_10_84_1153_0, i_10_84_1174_0,
    i_10_84_1175_0, i_10_84_1205_0, i_10_84_1233_0, i_10_84_1234_0,
    i_10_84_1238_0, i_10_84_1246_0, i_10_84_1247_0, i_10_84_1248_0,
    i_10_84_1308_0, i_10_84_1349_0, i_10_84_1363_0, i_10_84_1555_0,
    i_10_84_1556_0, i_10_84_1610_0, i_10_84_1627_0, i_10_84_1648_0,
    i_10_84_1687_0, i_10_84_1818_0, i_10_84_1819_0, i_10_84_1825_0,
    i_10_84_1950_0, i_10_84_2002_0, i_10_84_2003_0, i_10_84_2350_0,
    i_10_84_2351_0, i_10_84_2357_0, i_10_84_2364_0, i_10_84_2384_0,
    i_10_84_2411_0, i_10_84_2449_0, i_10_84_2465_0, i_10_84_2519_0,
    i_10_84_2540_0, i_10_84_2542_0, i_10_84_2543_0, i_10_84_2545_0,
    i_10_84_2572_0, i_10_84_2573_0, i_10_84_2634_0, i_10_84_2635_0,
    i_10_84_2708_0, i_10_84_2712_0, i_10_84_2730_0, i_10_84_2818_0,
    i_10_84_2830_0, i_10_84_2880_0, i_10_84_2887_0, i_10_84_2917_0,
    i_10_84_2918_0, i_10_84_2921_0, i_10_84_2922_0, i_10_84_2956_0,
    i_10_84_3039_0, i_10_84_3049_0, i_10_84_3090_0, i_10_84_3091_0,
    i_10_84_3162_0, i_10_84_3163_0, i_10_84_3277_0, i_10_84_3356_0,
    i_10_84_3390_0, i_10_84_3392_0, i_10_84_3446_0, i_10_84_3586_0,
    i_10_84_3613_0, i_10_84_3688_0, i_10_84_3689_0, i_10_84_3717_0,
    i_10_84_3734_0, i_10_84_3786_0, i_10_84_3850_0, i_10_84_3859_0,
    i_10_84_3892_0, i_10_84_4168_0, i_10_84_4267_0, i_10_84_4276_0,
    i_10_84_4277_0, i_10_84_4279_0, i_10_84_4568_0, i_10_84_4571_0;
  output o_10_84_0_0;
  assign o_10_84_0_0 = 0;
endmodule



// Benchmark "kernel_10_85" written by ABC on Sun Jul 19 10:22:27 2020

module kernel_10_85 ( 
    i_10_85_64_0, i_10_85_253_0, i_10_85_254_0, i_10_85_316_0,
    i_10_85_328_0, i_10_85_388_0, i_10_85_390_0, i_10_85_391_0,
    i_10_85_435_0, i_10_85_442_0, i_10_85_443_0, i_10_85_444_0,
    i_10_85_466_0, i_10_85_467_0, i_10_85_504_0, i_10_85_512_0,
    i_10_85_793_0, i_10_85_796_0, i_10_85_800_0, i_10_85_1002_0,
    i_10_85_1027_0, i_10_85_1028_0, i_10_85_1033_0, i_10_85_1034_0,
    i_10_85_1343_0, i_10_85_1433_0, i_10_85_1436_0, i_10_85_1442_0,
    i_10_85_1445_0, i_10_85_1539_0, i_10_85_1540_0, i_10_85_1541_0,
    i_10_85_1576_0, i_10_85_1579_0, i_10_85_1580_0, i_10_85_1620_0,
    i_10_85_1650_0, i_10_85_1688_0, i_10_85_1689_0, i_10_85_1690_0,
    i_10_85_1818_0, i_10_85_1819_0, i_10_85_1823_0, i_10_85_1910_0,
    i_10_85_1984_0, i_10_85_1988_0, i_10_85_1995_0, i_10_85_2198_0,
    i_10_85_2305_0, i_10_85_2306_0, i_10_85_2349_0, i_10_85_2363_0,
    i_10_85_2380_0, i_10_85_2530_0, i_10_85_2531_0, i_10_85_2603_0,
    i_10_85_2655_0, i_10_85_2677_0, i_10_85_2712_0, i_10_85_2721_0,
    i_10_85_2723_0, i_10_85_2735_0, i_10_85_2829_0, i_10_85_2830_0,
    i_10_85_2862_0, i_10_85_2863_0, i_10_85_2885_0, i_10_85_2924_0,
    i_10_85_3036_0, i_10_85_3088_0, i_10_85_3199_0, i_10_85_3201_0,
    i_10_85_3202_0, i_10_85_3270_0, i_10_85_3277_0, i_10_85_3278_0,
    i_10_85_3298_0, i_10_85_3321_0, i_10_85_3325_0, i_10_85_3386_0,
    i_10_85_3392_0, i_10_85_3406_0, i_10_85_3407_0, i_10_85_3614_0,
    i_10_85_3781_0, i_10_85_3782_0, i_10_85_3783_0, i_10_85_3784_0,
    i_10_85_3837_0, i_10_85_3853_0, i_10_85_3943_0, i_10_85_3979_0,
    i_10_85_3980_0, i_10_85_4006_0, i_10_85_4116_0, i_10_85_4286_0,
    i_10_85_4287_0, i_10_85_4565_0, i_10_85_4591_0, i_10_85_4592_0,
    o_10_85_0_0  );
  input  i_10_85_64_0, i_10_85_253_0, i_10_85_254_0, i_10_85_316_0,
    i_10_85_328_0, i_10_85_388_0, i_10_85_390_0, i_10_85_391_0,
    i_10_85_435_0, i_10_85_442_0, i_10_85_443_0, i_10_85_444_0,
    i_10_85_466_0, i_10_85_467_0, i_10_85_504_0, i_10_85_512_0,
    i_10_85_793_0, i_10_85_796_0, i_10_85_800_0, i_10_85_1002_0,
    i_10_85_1027_0, i_10_85_1028_0, i_10_85_1033_0, i_10_85_1034_0,
    i_10_85_1343_0, i_10_85_1433_0, i_10_85_1436_0, i_10_85_1442_0,
    i_10_85_1445_0, i_10_85_1539_0, i_10_85_1540_0, i_10_85_1541_0,
    i_10_85_1576_0, i_10_85_1579_0, i_10_85_1580_0, i_10_85_1620_0,
    i_10_85_1650_0, i_10_85_1688_0, i_10_85_1689_0, i_10_85_1690_0,
    i_10_85_1818_0, i_10_85_1819_0, i_10_85_1823_0, i_10_85_1910_0,
    i_10_85_1984_0, i_10_85_1988_0, i_10_85_1995_0, i_10_85_2198_0,
    i_10_85_2305_0, i_10_85_2306_0, i_10_85_2349_0, i_10_85_2363_0,
    i_10_85_2380_0, i_10_85_2530_0, i_10_85_2531_0, i_10_85_2603_0,
    i_10_85_2655_0, i_10_85_2677_0, i_10_85_2712_0, i_10_85_2721_0,
    i_10_85_2723_0, i_10_85_2735_0, i_10_85_2829_0, i_10_85_2830_0,
    i_10_85_2862_0, i_10_85_2863_0, i_10_85_2885_0, i_10_85_2924_0,
    i_10_85_3036_0, i_10_85_3088_0, i_10_85_3199_0, i_10_85_3201_0,
    i_10_85_3202_0, i_10_85_3270_0, i_10_85_3277_0, i_10_85_3278_0,
    i_10_85_3298_0, i_10_85_3321_0, i_10_85_3325_0, i_10_85_3386_0,
    i_10_85_3392_0, i_10_85_3406_0, i_10_85_3407_0, i_10_85_3614_0,
    i_10_85_3781_0, i_10_85_3782_0, i_10_85_3783_0, i_10_85_3784_0,
    i_10_85_3837_0, i_10_85_3853_0, i_10_85_3943_0, i_10_85_3979_0,
    i_10_85_3980_0, i_10_85_4006_0, i_10_85_4116_0, i_10_85_4286_0,
    i_10_85_4287_0, i_10_85_4565_0, i_10_85_4591_0, i_10_85_4592_0;
  output o_10_85_0_0;
  assign o_10_85_0_0 = ~((~i_10_85_3614_0 & ((~i_10_85_1002_0 & ~i_10_85_3979_0 & ((~i_10_85_467_0 & ~i_10_85_1541_0 & i_10_85_1819_0 & ~i_10_85_3270_0 & ~i_10_85_3406_0 & i_10_85_3853_0) | (~i_10_85_3837_0 & i_10_85_4287_0))) | (~i_10_85_1540_0 & ~i_10_85_2198_0 & ((~i_10_85_2306_0 & ~i_10_85_3088_0 & ~i_10_85_3277_0 & ~i_10_85_3783_0) | (~i_10_85_466_0 & ~i_10_85_1620_0 & ~i_10_85_2305_0 & ~i_10_85_2924_0 & ~i_10_85_3386_0 & ~i_10_85_3784_0 & ~i_10_85_3980_0))) | (~i_10_85_1688_0 & ~i_10_85_2305_0 & ~i_10_85_2603_0 & ~i_10_85_2655_0 & ~i_10_85_2677_0 & ~i_10_85_2721_0 & ~i_10_85_2885_0 & ~i_10_85_3270_0 & i_10_85_3853_0))) | (~i_10_85_1539_0 & ((~i_10_85_388_0 & ~i_10_85_1027_0 & ~i_10_85_1028_0 & ~i_10_85_1433_0 & ~i_10_85_1995_0 & ~i_10_85_2885_0 & ~i_10_85_3088_0) | (~i_10_85_390_0 & i_10_85_467_0 & ~i_10_85_1541_0 & ~i_10_85_1910_0 & ~i_10_85_2712_0 & ~i_10_85_2735_0 & ~i_10_85_3407_0))) | (~i_10_85_2885_0 & ((~i_10_85_388_0 & ((~i_10_85_316_0 & ~i_10_85_1027_0 & ~i_10_85_1028_0 & ~i_10_85_1995_0 & ~i_10_85_3278_0) | (~i_10_85_1541_0 & i_10_85_1689_0 & i_10_85_1819_0 & ~i_10_85_2924_0 & ~i_10_85_3853_0))) | (~i_10_85_316_0 & ~i_10_85_1540_0 & ~i_10_85_1910_0 & ((~i_10_85_796_0 & ~i_10_85_1541_0 & ~i_10_85_1580_0 & ~i_10_85_2306_0 & ~i_10_85_2603_0) | (~i_10_85_1576_0 & ~i_10_85_3036_0 & ~i_10_85_3201_0 & ~i_10_85_3784_0))))) | (~i_10_85_1433_0 & ((~i_10_85_467_0 & ~i_10_85_1343_0 & ~i_10_85_1620_0 & ~i_10_85_1688_0 & i_10_85_1819_0 & ~i_10_85_2603_0) | (~i_10_85_1028_0 & i_10_85_1576_0 & ~i_10_85_2305_0 & ~i_10_85_2723_0 & ~i_10_85_2735_0 & ~i_10_85_3277_0))) | (~i_10_85_3386_0 & ((~i_10_85_467_0 & ((~i_10_85_390_0 & i_10_85_2723_0 & i_10_85_3614_0 & ~i_10_85_3784_0) | (~i_10_85_1033_0 & i_10_85_1579_0 & ~i_10_85_1620_0 & ~i_10_85_2198_0 & ~i_10_85_2924_0 & ~i_10_85_3202_0 & ~i_10_85_3270_0 & ~i_10_85_3407_0 & ~i_10_85_4286_0))) | (~i_10_85_254_0 & ~i_10_85_435_0 & i_10_85_796_0 & ~i_10_85_1995_0))) | (~i_10_85_254_0 & ((~i_10_85_390_0 & ~i_10_85_1541_0 & ~i_10_85_2349_0 & ~i_10_85_3201_0 & ~i_10_85_3392_0 & ~i_10_85_3406_0 & ~i_10_85_3781_0) | (~i_10_85_391_0 & ~i_10_85_1689_0 & i_10_85_1818_0 & i_10_85_2349_0 & ~i_10_85_4286_0))) | (~i_10_85_4286_0 & ((~i_10_85_1580_0 & ((~i_10_85_1027_0 & ~i_10_85_1540_0 & ~i_10_85_3199_0 & ~i_10_85_3392_0) | (~i_10_85_316_0 & ~i_10_85_3202_0 & ~i_10_85_3783_0 & i_10_85_3837_0))) | (~i_10_85_390_0 & ~i_10_85_1688_0 & ~i_10_85_2305_0 & ~i_10_85_2603_0 & ~i_10_85_3277_0 & ~i_10_85_3278_0 & ~i_10_85_3782_0))) | (i_10_85_3270_0 & ~i_10_85_3782_0 & (i_10_85_4116_0 | (i_10_85_1579_0 & ~i_10_85_3202_0 & i_10_85_3853_0))) | (i_10_85_1688_0 & i_10_85_2830_0));
endmodule



// Benchmark "kernel_10_86" written by ABC on Sun Jul 19 10:22:28 2020

module kernel_10_86 ( 
    i_10_86_174_0, i_10_86_220_0, i_10_86_221_0, i_10_86_245_0,
    i_10_86_287_0, i_10_86_328_0, i_10_86_408_0, i_10_86_409_0,
    i_10_86_410_0, i_10_86_441_0, i_10_86_442_0, i_10_86_508_0,
    i_10_86_509_0, i_10_86_797_0, i_10_86_892_0, i_10_86_958_0,
    i_10_86_994_0, i_10_86_1026_0, i_10_86_1027_0, i_10_86_1028_0,
    i_10_86_1242_0, i_10_86_1262_0, i_10_86_1305_0, i_10_86_1432_0,
    i_10_86_1541_0, i_10_86_1620_0, i_10_86_1621_0, i_10_86_1685_0,
    i_10_86_1691_0, i_10_86_1819_0, i_10_86_1820_0, i_10_86_1821_0,
    i_10_86_1909_0, i_10_86_1990_0, i_10_86_2161_0, i_10_86_2353_0,
    i_10_86_2356_0, i_10_86_2359_0, i_10_86_2362_0, i_10_86_2448_0,
    i_10_86_2450_0, i_10_86_2566_0, i_10_86_2628_0, i_10_86_2629_0,
    i_10_86_2630_0, i_10_86_2631_0, i_10_86_2632_0, i_10_86_2633_0,
    i_10_86_2635_0, i_10_86_2719_0, i_10_86_2722_0, i_10_86_2729_0,
    i_10_86_2781_0, i_10_86_2785_0, i_10_86_2817_0, i_10_86_2818_0,
    i_10_86_2826_0, i_10_86_2827_0, i_10_86_2828_0, i_10_86_2834_0,
    i_10_86_2880_0, i_10_86_2881_0, i_10_86_2882_0, i_10_86_2884_0,
    i_10_86_2921_0, i_10_86_2923_0, i_10_86_2924_0, i_10_86_3069_0,
    i_10_86_3070_0, i_10_86_3088_0, i_10_86_3199_0, i_10_86_3272_0,
    i_10_86_3384_0, i_10_86_3407_0, i_10_86_3523_0, i_10_86_3555_0,
    i_10_86_3583_0, i_10_86_3584_0, i_10_86_3585_0, i_10_86_3610_0,
    i_10_86_3612_0, i_10_86_3780_0, i_10_86_3783_0, i_10_86_3785_0,
    i_10_86_3838_0, i_10_86_3839_0, i_10_86_3844_0, i_10_86_3846_0,
    i_10_86_3852_0, i_10_86_3889_0, i_10_86_4114_0, i_10_86_4116_0,
    i_10_86_4122_0, i_10_86_4123_0, i_10_86_4126_0, i_10_86_4168_0,
    i_10_86_4214_0, i_10_86_4566_0, i_10_86_4590_0, i_10_86_4591_0,
    o_10_86_0_0  );
  input  i_10_86_174_0, i_10_86_220_0, i_10_86_221_0, i_10_86_245_0,
    i_10_86_287_0, i_10_86_328_0, i_10_86_408_0, i_10_86_409_0,
    i_10_86_410_0, i_10_86_441_0, i_10_86_442_0, i_10_86_508_0,
    i_10_86_509_0, i_10_86_797_0, i_10_86_892_0, i_10_86_958_0,
    i_10_86_994_0, i_10_86_1026_0, i_10_86_1027_0, i_10_86_1028_0,
    i_10_86_1242_0, i_10_86_1262_0, i_10_86_1305_0, i_10_86_1432_0,
    i_10_86_1541_0, i_10_86_1620_0, i_10_86_1621_0, i_10_86_1685_0,
    i_10_86_1691_0, i_10_86_1819_0, i_10_86_1820_0, i_10_86_1821_0,
    i_10_86_1909_0, i_10_86_1990_0, i_10_86_2161_0, i_10_86_2353_0,
    i_10_86_2356_0, i_10_86_2359_0, i_10_86_2362_0, i_10_86_2448_0,
    i_10_86_2450_0, i_10_86_2566_0, i_10_86_2628_0, i_10_86_2629_0,
    i_10_86_2630_0, i_10_86_2631_0, i_10_86_2632_0, i_10_86_2633_0,
    i_10_86_2635_0, i_10_86_2719_0, i_10_86_2722_0, i_10_86_2729_0,
    i_10_86_2781_0, i_10_86_2785_0, i_10_86_2817_0, i_10_86_2818_0,
    i_10_86_2826_0, i_10_86_2827_0, i_10_86_2828_0, i_10_86_2834_0,
    i_10_86_2880_0, i_10_86_2881_0, i_10_86_2882_0, i_10_86_2884_0,
    i_10_86_2921_0, i_10_86_2923_0, i_10_86_2924_0, i_10_86_3069_0,
    i_10_86_3070_0, i_10_86_3088_0, i_10_86_3199_0, i_10_86_3272_0,
    i_10_86_3384_0, i_10_86_3407_0, i_10_86_3523_0, i_10_86_3555_0,
    i_10_86_3583_0, i_10_86_3584_0, i_10_86_3585_0, i_10_86_3610_0,
    i_10_86_3612_0, i_10_86_3780_0, i_10_86_3783_0, i_10_86_3785_0,
    i_10_86_3838_0, i_10_86_3839_0, i_10_86_3844_0, i_10_86_3846_0,
    i_10_86_3852_0, i_10_86_3889_0, i_10_86_4114_0, i_10_86_4116_0,
    i_10_86_4122_0, i_10_86_4123_0, i_10_86_4126_0, i_10_86_4168_0,
    i_10_86_4214_0, i_10_86_4566_0, i_10_86_4590_0, i_10_86_4591_0;
  output o_10_86_0_0;
  assign o_10_86_0_0 = ~((~i_10_86_2566_0 & ((~i_10_86_174_0 & ((~i_10_86_220_0 & ~i_10_86_410_0 & ~i_10_86_1027_0 & ~i_10_86_1541_0 & ~i_10_86_1620_0 & ~i_10_86_3070_0) | (~i_10_86_408_0 & ~i_10_86_2630_0 & ~i_10_86_2632_0 & ~i_10_86_2781_0 & ~i_10_86_2921_0 & ~i_10_86_3523_0 & ~i_10_86_3780_0 & ~i_10_86_3846_0 & ~i_10_86_4168_0))) | (~i_10_86_1026_0 & i_10_86_2828_0 & ~i_10_86_2884_0) | (~i_10_86_1541_0 & i_10_86_2632_0 & ~i_10_86_2729_0 & ~i_10_86_2828_0 & i_10_86_2923_0 & ~i_10_86_3070_0))) | (~i_10_86_4114_0 & ((~i_10_86_220_0 & ((i_10_86_1819_0 & ~i_10_86_2722_0 & ~i_10_86_2781_0 & ~i_10_86_2785_0 & ~i_10_86_3199_0 & ~i_10_86_4123_0) | (~i_10_86_410_0 & ~i_10_86_1432_0 & ~i_10_86_2834_0 & i_10_86_3852_0 & ~i_10_86_4116_0 & ~i_10_86_4126_0))) | (~i_10_86_245_0 & i_10_86_1691_0 & i_10_86_2921_0 & ~i_10_86_4123_0))) | (~i_10_86_245_0 & ((i_10_86_442_0 & ~i_10_86_1685_0 & ~i_10_86_3523_0 & ~i_10_86_3838_0) | (~i_10_86_408_0 & ~i_10_86_1621_0 & ~i_10_86_2353_0 & ~i_10_86_2356_0 & ~i_10_86_2448_0 & ~i_10_86_2722_0 & ~i_10_86_2781_0 & ~i_10_86_3069_0 & ~i_10_86_3070_0 & ~i_10_86_3407_0 & ~i_10_86_4126_0 & ~i_10_86_4214_0))) | (~i_10_86_1242_0 & ((~i_10_86_994_0 & ~i_10_86_1821_0 & ~i_10_86_3272_0 & i_10_86_3407_0 & ~i_10_86_3838_0 & ~i_10_86_3839_0) | (~i_10_86_797_0 & ~i_10_86_1685_0 & ~i_10_86_1990_0 & ~i_10_86_2834_0 & ~i_10_86_3069_0 & ~i_10_86_3612_0 & ~i_10_86_4126_0 & ~i_10_86_4168_0 & ~i_10_86_4214_0 & ~i_10_86_4566_0))) | (i_10_86_2827_0 & ((~i_10_86_1541_0 & ~i_10_86_1990_0 & i_10_86_2362_0 & ~i_10_86_2448_0) | (~i_10_86_2359_0 & ~i_10_86_4122_0))) | (~i_10_86_2359_0 & ((~i_10_86_1541_0 & ~i_10_86_1620_0 & ~i_10_86_2923_0 & ~i_10_86_3780_0 & i_10_86_4116_0 & ~i_10_86_4123_0) | (i_10_86_408_0 & ~i_10_86_1432_0 & ~i_10_86_2635_0 & ~i_10_86_2834_0 & ~i_10_86_3846_0 & ~i_10_86_4566_0))) | (~i_10_86_409_0 & ((~i_10_86_1541_0 & ~i_10_86_4214_0 & ((~i_10_86_1026_0 & i_10_86_1821_0 & ~i_10_86_1990_0 & ~i_10_86_3272_0 & ~i_10_86_4122_0) | (~i_10_86_2353_0 & ~i_10_86_3069_0 & ~i_10_86_3785_0 & ~i_10_86_3846_0 & ~i_10_86_4123_0))) | (~i_10_86_1685_0 & ~i_10_86_1819_0 & ~i_10_86_2834_0 & i_10_86_2924_0 & ~i_10_86_3384_0 & ~i_10_86_3783_0))) | (~i_10_86_1990_0 & ((~i_10_86_3612_0 & ~i_10_86_4126_0 & ~i_10_86_1028_0 & i_10_86_2450_0) | (~i_10_86_2630_0 & ~i_10_86_2632_0 & ~i_10_86_2729_0 & ~i_10_86_2834_0 & ~i_10_86_3069_0 & ~i_10_86_3780_0 & ~i_10_86_3783_0 & ~i_10_86_3785_0 & ~i_10_86_4123_0 & ~i_10_86_4168_0))) | (~i_10_86_3384_0 & ((i_10_86_2630_0 & ~i_10_86_2722_0 & i_10_86_2729_0 & ~i_10_86_3783_0) | (~i_10_86_2923_0 & ~i_10_86_3070_0 & ~i_10_86_3583_0 & i_10_86_3612_0 & ~i_10_86_3785_0))) | (~i_10_86_3070_0 & ((i_10_86_328_0 & ~i_10_86_2362_0) | (i_10_86_2353_0 & i_10_86_3844_0 & ~i_10_86_3846_0) | (~i_10_86_892_0 & ~i_10_86_1027_0 & ~i_10_86_1621_0 & ~i_10_86_3199_0 & ~i_10_86_4122_0))));
endmodule



// Benchmark "kernel_10_87" written by ABC on Sun Jul 19 10:22:29 2020

module kernel_10_87 ( 
    i_10_87_182_0, i_10_87_220_0, i_10_87_247_0, i_10_87_285_0,
    i_10_87_290_0, i_10_87_328_0, i_10_87_329_0, i_10_87_371_0,
    i_10_87_407_0, i_10_87_623_0, i_10_87_729_0, i_10_87_730_0,
    i_10_87_731_0, i_10_87_733_0, i_10_87_754_0, i_10_87_796_0,
    i_10_87_797_0, i_10_87_899_0, i_10_87_1030_0, i_10_87_1031_0,
    i_10_87_1219_0, i_10_87_1264_0, i_10_87_1267_0, i_10_87_1306_0,
    i_10_87_1307_0, i_10_87_1308_0, i_10_87_1312_0, i_10_87_1345_0,
    i_10_87_1349_0, i_10_87_1441_0, i_10_87_1442_0, i_10_87_1913_0,
    i_10_87_1987_0, i_10_87_2017_0, i_10_87_2019_0, i_10_87_2020_0,
    i_10_87_2197_0, i_10_87_2201_0, i_10_87_2324_0, i_10_87_2358_0,
    i_10_87_2386_0, i_10_87_2461_0, i_10_87_2463_0, i_10_87_2464_0,
    i_10_87_2467_0, i_10_87_2471_0, i_10_87_2628_0, i_10_87_2631_0,
    i_10_87_2632_0, i_10_87_2656_0, i_10_87_2704_0, i_10_87_2722_0,
    i_10_87_2785_0, i_10_87_2804_0, i_10_87_2827_0, i_10_87_2870_0,
    i_10_87_2916_0, i_10_87_2917_0, i_10_87_2918_0, i_10_87_2919_0,
    i_10_87_2920_0, i_10_87_2922_0, i_10_87_2984_0, i_10_87_3035_0,
    i_10_87_3070_0, i_10_87_3196_0, i_10_87_3203_0, i_10_87_3390_0,
    i_10_87_3402_0, i_10_87_3430_0, i_10_87_3519_0, i_10_87_3522_0,
    i_10_87_3588_0, i_10_87_3609_0, i_10_87_3611_0, i_10_87_3614_0,
    i_10_87_3645_0, i_10_87_3647_0, i_10_87_3648_0, i_10_87_3649_0,
    i_10_87_3734_0, i_10_87_3783_0, i_10_87_3787_0, i_10_87_3788_0,
    i_10_87_3842_0, i_10_87_3853_0, i_10_87_3855_0, i_10_87_4028_0,
    i_10_87_4113_0, i_10_87_4167_0, i_10_87_4170_0, i_10_87_4171_0,
    i_10_87_4172_0, i_10_87_4212_0, i_10_87_4215_0, i_10_87_4216_0,
    i_10_87_4217_0, i_10_87_4288_0, i_10_87_4289_0, i_10_87_4462_0,
    o_10_87_0_0  );
  input  i_10_87_182_0, i_10_87_220_0, i_10_87_247_0, i_10_87_285_0,
    i_10_87_290_0, i_10_87_328_0, i_10_87_329_0, i_10_87_371_0,
    i_10_87_407_0, i_10_87_623_0, i_10_87_729_0, i_10_87_730_0,
    i_10_87_731_0, i_10_87_733_0, i_10_87_754_0, i_10_87_796_0,
    i_10_87_797_0, i_10_87_899_0, i_10_87_1030_0, i_10_87_1031_0,
    i_10_87_1219_0, i_10_87_1264_0, i_10_87_1267_0, i_10_87_1306_0,
    i_10_87_1307_0, i_10_87_1308_0, i_10_87_1312_0, i_10_87_1345_0,
    i_10_87_1349_0, i_10_87_1441_0, i_10_87_1442_0, i_10_87_1913_0,
    i_10_87_1987_0, i_10_87_2017_0, i_10_87_2019_0, i_10_87_2020_0,
    i_10_87_2197_0, i_10_87_2201_0, i_10_87_2324_0, i_10_87_2358_0,
    i_10_87_2386_0, i_10_87_2461_0, i_10_87_2463_0, i_10_87_2464_0,
    i_10_87_2467_0, i_10_87_2471_0, i_10_87_2628_0, i_10_87_2631_0,
    i_10_87_2632_0, i_10_87_2656_0, i_10_87_2704_0, i_10_87_2722_0,
    i_10_87_2785_0, i_10_87_2804_0, i_10_87_2827_0, i_10_87_2870_0,
    i_10_87_2916_0, i_10_87_2917_0, i_10_87_2918_0, i_10_87_2919_0,
    i_10_87_2920_0, i_10_87_2922_0, i_10_87_2984_0, i_10_87_3035_0,
    i_10_87_3070_0, i_10_87_3196_0, i_10_87_3203_0, i_10_87_3390_0,
    i_10_87_3402_0, i_10_87_3430_0, i_10_87_3519_0, i_10_87_3522_0,
    i_10_87_3588_0, i_10_87_3609_0, i_10_87_3611_0, i_10_87_3614_0,
    i_10_87_3645_0, i_10_87_3647_0, i_10_87_3648_0, i_10_87_3649_0,
    i_10_87_3734_0, i_10_87_3783_0, i_10_87_3787_0, i_10_87_3788_0,
    i_10_87_3842_0, i_10_87_3853_0, i_10_87_3855_0, i_10_87_4028_0,
    i_10_87_4113_0, i_10_87_4167_0, i_10_87_4170_0, i_10_87_4171_0,
    i_10_87_4172_0, i_10_87_4212_0, i_10_87_4215_0, i_10_87_4216_0,
    i_10_87_4217_0, i_10_87_4288_0, i_10_87_4289_0, i_10_87_4462_0;
  output o_10_87_0_0;
  assign o_10_87_0_0 = 0;
endmodule



// Benchmark "kernel_10_88" written by ABC on Sun Jul 19 10:22:30 2020

module kernel_10_88 ( 
    i_10_88_86_0, i_10_88_174_0, i_10_88_177_0, i_10_88_179_0,
    i_10_88_264_0, i_10_88_284_0, i_10_88_409_0, i_10_88_413_0,
    i_10_88_536_0, i_10_88_635_0, i_10_88_754_0, i_10_88_797_0,
    i_10_88_961_0, i_10_88_964_0, i_10_88_994_0, i_10_88_996_0,
    i_10_88_1028_0, i_10_88_1160_0, i_10_88_1238_0, i_10_88_1241_0,
    i_10_88_1274_0, i_10_88_1310_0, i_10_88_1345_0, i_10_88_1346_0,
    i_10_88_1360_0, i_10_88_1361_0, i_10_88_1364_0, i_10_88_1436_0,
    i_10_88_1438_0, i_10_88_1439_0, i_10_88_1542_0, i_10_88_1547_0,
    i_10_88_1549_0, i_10_88_1555_0, i_10_88_1582_0, i_10_88_1625_0,
    i_10_88_1627_0, i_10_88_1628_0, i_10_88_1650_0, i_10_88_1736_0,
    i_10_88_1821_0, i_10_88_1823_0, i_10_88_1994_0, i_10_88_2023_0,
    i_10_88_2024_0, i_10_88_2032_0, i_10_88_2033_0, i_10_88_2201_0,
    i_10_88_2324_0, i_10_88_2350_0, i_10_88_2364_0, i_10_88_2453_0,
    i_10_88_2456_0, i_10_88_2507_0, i_10_88_2516_0, i_10_88_2609_0,
    i_10_88_2628_0, i_10_88_2632_0, i_10_88_2656_0, i_10_88_2674_0,
    i_10_88_2678_0, i_10_88_2711_0, i_10_88_2717_0, i_10_88_2732_0,
    i_10_88_2734_0, i_10_88_2783_0, i_10_88_2789_0, i_10_88_2829_0,
    i_10_88_2831_0, i_10_88_2850_0, i_10_88_2884_0, i_10_88_2885_0,
    i_10_88_2967_0, i_10_88_2968_0, i_10_88_2969_0, i_10_88_3047_0,
    i_10_88_3074_0, i_10_88_3077_0, i_10_88_3091_0, i_10_88_3199_0,
    i_10_88_3277_0, i_10_88_3290_0, i_10_88_3337_0, i_10_88_3431_0,
    i_10_88_3434_0, i_10_88_3470_0, i_10_88_3494_0, i_10_88_3507_0,
    i_10_88_3584_0, i_10_88_3652_0, i_10_88_3841_0, i_10_88_3850_0,
    i_10_88_3860_0, i_10_88_4051_0, i_10_88_4130_0, i_10_88_4175_0,
    i_10_88_4262_0, i_10_88_4292_0, i_10_88_4460_0, i_10_88_4586_0,
    o_10_88_0_0  );
  input  i_10_88_86_0, i_10_88_174_0, i_10_88_177_0, i_10_88_179_0,
    i_10_88_264_0, i_10_88_284_0, i_10_88_409_0, i_10_88_413_0,
    i_10_88_536_0, i_10_88_635_0, i_10_88_754_0, i_10_88_797_0,
    i_10_88_961_0, i_10_88_964_0, i_10_88_994_0, i_10_88_996_0,
    i_10_88_1028_0, i_10_88_1160_0, i_10_88_1238_0, i_10_88_1241_0,
    i_10_88_1274_0, i_10_88_1310_0, i_10_88_1345_0, i_10_88_1346_0,
    i_10_88_1360_0, i_10_88_1361_0, i_10_88_1364_0, i_10_88_1436_0,
    i_10_88_1438_0, i_10_88_1439_0, i_10_88_1542_0, i_10_88_1547_0,
    i_10_88_1549_0, i_10_88_1555_0, i_10_88_1582_0, i_10_88_1625_0,
    i_10_88_1627_0, i_10_88_1628_0, i_10_88_1650_0, i_10_88_1736_0,
    i_10_88_1821_0, i_10_88_1823_0, i_10_88_1994_0, i_10_88_2023_0,
    i_10_88_2024_0, i_10_88_2032_0, i_10_88_2033_0, i_10_88_2201_0,
    i_10_88_2324_0, i_10_88_2350_0, i_10_88_2364_0, i_10_88_2453_0,
    i_10_88_2456_0, i_10_88_2507_0, i_10_88_2516_0, i_10_88_2609_0,
    i_10_88_2628_0, i_10_88_2632_0, i_10_88_2656_0, i_10_88_2674_0,
    i_10_88_2678_0, i_10_88_2711_0, i_10_88_2717_0, i_10_88_2732_0,
    i_10_88_2734_0, i_10_88_2783_0, i_10_88_2789_0, i_10_88_2829_0,
    i_10_88_2831_0, i_10_88_2850_0, i_10_88_2884_0, i_10_88_2885_0,
    i_10_88_2967_0, i_10_88_2968_0, i_10_88_2969_0, i_10_88_3047_0,
    i_10_88_3074_0, i_10_88_3077_0, i_10_88_3091_0, i_10_88_3199_0,
    i_10_88_3277_0, i_10_88_3290_0, i_10_88_3337_0, i_10_88_3431_0,
    i_10_88_3434_0, i_10_88_3470_0, i_10_88_3494_0, i_10_88_3507_0,
    i_10_88_3584_0, i_10_88_3652_0, i_10_88_3841_0, i_10_88_3850_0,
    i_10_88_3860_0, i_10_88_4051_0, i_10_88_4130_0, i_10_88_4175_0,
    i_10_88_4262_0, i_10_88_4292_0, i_10_88_4460_0, i_10_88_4586_0;
  output o_10_88_0_0;
  assign o_10_88_0_0 = 0;
endmodule



// Benchmark "kernel_10_89" written by ABC on Sun Jul 19 10:22:31 2020

module kernel_10_89 ( 
    i_10_89_68_0, i_10_89_263_0, i_10_89_270_0, i_10_89_273_0,
    i_10_89_274_0, i_10_89_282_0, i_10_89_283_0, i_10_89_284_0,
    i_10_89_287_0, i_10_89_315_0, i_10_89_317_0, i_10_89_318_0,
    i_10_89_319_0, i_10_89_320_0, i_10_89_322_0, i_10_89_323_0,
    i_10_89_391_0, i_10_89_392_0, i_10_89_410_0, i_10_89_442_0,
    i_10_89_443_0, i_10_89_559_0, i_10_89_560_0, i_10_89_991_0,
    i_10_89_1001_0, i_10_89_1004_0, i_10_89_1085_0, i_10_89_1111_0,
    i_10_89_1138_0, i_10_89_1235_0, i_10_89_1238_0, i_10_89_1307_0,
    i_10_89_1309_0, i_10_89_1310_0, i_10_89_1311_0, i_10_89_1360_0,
    i_10_89_1379_0, i_10_89_1433_0, i_10_89_1436_0, i_10_89_1442_0,
    i_10_89_1544_0, i_10_89_1546_0, i_10_89_1547_0, i_10_89_1580_0,
    i_10_89_1651_0, i_10_89_1652_0, i_10_89_1730_0, i_10_89_1825_0,
    i_10_89_1826_0, i_10_89_2000_0, i_10_89_2024_0, i_10_89_2312_0,
    i_10_89_2352_0, i_10_89_2354_0, i_10_89_2356_0, i_10_89_2449_0,
    i_10_89_2468_0, i_10_89_2538_0, i_10_89_2558_0, i_10_89_2567_0,
    i_10_89_2605_0, i_10_89_2615_0, i_10_89_2632_0, i_10_89_2703_0,
    i_10_89_2704_0, i_10_89_2707_0, i_10_89_2713_0, i_10_89_2719_0,
    i_10_89_2723_0, i_10_89_2727_0, i_10_89_2728_0, i_10_89_2731_0,
    i_10_89_2833_0, i_10_89_2834_0, i_10_89_3044_0, i_10_89_3072_0,
    i_10_89_3268_0, i_10_89_3467_0, i_10_89_3542_0, i_10_89_3545_0,
    i_10_89_3584_0, i_10_89_3647_0, i_10_89_3650_0, i_10_89_3653_0,
    i_10_89_3775_0, i_10_89_3785_0, i_10_89_3839_0, i_10_89_3840_0,
    i_10_89_3859_0, i_10_89_3980_0, i_10_89_3983_0, i_10_89_3986_0,
    i_10_89_4114_0, i_10_89_4115_0, i_10_89_4116_0, i_10_89_4117_0,
    i_10_89_4121_0, i_10_89_4283_0, i_10_89_4285_0, i_10_89_4288_0,
    o_10_89_0_0  );
  input  i_10_89_68_0, i_10_89_263_0, i_10_89_270_0, i_10_89_273_0,
    i_10_89_274_0, i_10_89_282_0, i_10_89_283_0, i_10_89_284_0,
    i_10_89_287_0, i_10_89_315_0, i_10_89_317_0, i_10_89_318_0,
    i_10_89_319_0, i_10_89_320_0, i_10_89_322_0, i_10_89_323_0,
    i_10_89_391_0, i_10_89_392_0, i_10_89_410_0, i_10_89_442_0,
    i_10_89_443_0, i_10_89_559_0, i_10_89_560_0, i_10_89_991_0,
    i_10_89_1001_0, i_10_89_1004_0, i_10_89_1085_0, i_10_89_1111_0,
    i_10_89_1138_0, i_10_89_1235_0, i_10_89_1238_0, i_10_89_1307_0,
    i_10_89_1309_0, i_10_89_1310_0, i_10_89_1311_0, i_10_89_1360_0,
    i_10_89_1379_0, i_10_89_1433_0, i_10_89_1436_0, i_10_89_1442_0,
    i_10_89_1544_0, i_10_89_1546_0, i_10_89_1547_0, i_10_89_1580_0,
    i_10_89_1651_0, i_10_89_1652_0, i_10_89_1730_0, i_10_89_1825_0,
    i_10_89_1826_0, i_10_89_2000_0, i_10_89_2024_0, i_10_89_2312_0,
    i_10_89_2352_0, i_10_89_2354_0, i_10_89_2356_0, i_10_89_2449_0,
    i_10_89_2468_0, i_10_89_2538_0, i_10_89_2558_0, i_10_89_2567_0,
    i_10_89_2605_0, i_10_89_2615_0, i_10_89_2632_0, i_10_89_2703_0,
    i_10_89_2704_0, i_10_89_2707_0, i_10_89_2713_0, i_10_89_2719_0,
    i_10_89_2723_0, i_10_89_2727_0, i_10_89_2728_0, i_10_89_2731_0,
    i_10_89_2833_0, i_10_89_2834_0, i_10_89_3044_0, i_10_89_3072_0,
    i_10_89_3268_0, i_10_89_3467_0, i_10_89_3542_0, i_10_89_3545_0,
    i_10_89_3584_0, i_10_89_3647_0, i_10_89_3650_0, i_10_89_3653_0,
    i_10_89_3775_0, i_10_89_3785_0, i_10_89_3839_0, i_10_89_3840_0,
    i_10_89_3859_0, i_10_89_3980_0, i_10_89_3983_0, i_10_89_3986_0,
    i_10_89_4114_0, i_10_89_4115_0, i_10_89_4116_0, i_10_89_4117_0,
    i_10_89_4121_0, i_10_89_4283_0, i_10_89_4285_0, i_10_89_4288_0;
  output o_10_89_0_0;
  assign o_10_89_0_0 = ~((~i_10_89_284_0 & ((~i_10_89_323_0 & ~i_10_89_1085_0 & i_10_89_1651_0 & ~i_10_89_2312_0) | (~i_10_89_1307_0 & ~i_10_89_1547_0 & ~i_10_89_2468_0 & ~i_10_89_3983_0))) | (~i_10_89_392_0 & ((~i_10_89_1001_0 & ((~i_10_89_391_0 & ~i_10_89_1580_0 & i_10_89_2731_0) | (~i_10_89_1085_0 & ~i_10_89_1309_0 & ~i_10_89_1547_0 & ~i_10_89_2352_0 & ~i_10_89_2468_0 & ~i_10_89_2615_0 & ~i_10_89_3980_0))) | (~i_10_89_1360_0 & ((~i_10_89_560_0 & ~i_10_89_1004_0 & ~i_10_89_2024_0 & ~i_10_89_2312_0 & ~i_10_89_2356_0 & ~i_10_89_2615_0 & ~i_10_89_2707_0 & ~i_10_89_3044_0) | (~i_10_89_263_0 & ~i_10_89_1546_0 & ~i_10_89_2000_0 & ~i_10_89_2468_0 & ~i_10_89_3839_0 & ~i_10_89_3983_0 & ~i_10_89_3986_0 & ~i_10_89_4283_0))))) | (~i_10_89_3545_0 & ((~i_10_89_263_0 & ((~i_10_89_317_0 & ~i_10_89_443_0 & ~i_10_89_2312_0 & ~i_10_89_2728_0 & ~i_10_89_3467_0 & i_10_89_3840_0) | (~i_10_89_320_0 & ~i_10_89_1004_0 & ~i_10_89_1307_0 & ~i_10_89_2356_0 & ~i_10_89_3647_0 & ~i_10_89_3983_0))) | (~i_10_89_560_0 & ((i_10_89_991_0 & ~i_10_89_1310_0) | (~i_10_89_320_0 & ~i_10_89_410_0 & ~i_10_89_1004_0 & ~i_10_89_1433_0 & ~i_10_89_1580_0 & ~i_10_89_3542_0 & ~i_10_89_4121_0))) | (~i_10_89_2024_0 & ((~i_10_89_287_0 & ~i_10_89_323_0 & ~i_10_89_1360_0 & ~i_10_89_1544_0 & ~i_10_89_1651_0 & ~i_10_89_2731_0 & ~i_10_89_3467_0 & ~i_10_89_3647_0 & ~i_10_89_3983_0) | (~i_10_89_559_0 & ~i_10_89_1085_0 & ~i_10_89_1310_0 & ~i_10_89_2000_0 & i_10_89_2352_0 & ~i_10_89_3542_0 & ~i_10_89_3650_0 & ~i_10_89_4283_0))))) | (~i_10_89_317_0 & ((~i_10_89_442_0 & ~i_10_89_1360_0 & ~i_10_89_1580_0 & ~i_10_89_2354_0 & ~i_10_89_3467_0 & ~i_10_89_3986_0) | (~i_10_89_283_0 & ~i_10_89_1436_0 & ~i_10_89_2713_0 & ~i_10_89_3650_0 & ~i_10_89_4115_0))) | (~i_10_89_283_0 & ((i_10_89_318_0 & ~i_10_89_322_0 & i_10_89_3980_0) | (~i_10_89_1436_0 & i_10_89_1826_0 & ~i_10_89_2356_0 & ~i_10_89_2723_0 & ~i_10_89_3840_0 & ~i_10_89_3980_0))) | (~i_10_89_323_0 & (i_10_89_2833_0 | (i_10_89_2312_0 & i_10_89_3840_0))) | (~i_10_89_3467_0 & ((~i_10_89_1085_0 & ((~i_10_89_991_0 & ~i_10_89_1547_0 & i_10_89_1826_0 & ~i_10_89_3542_0 & ~i_10_89_3653_0) | (i_10_89_4116_0 & i_10_89_4117_0))) | (~i_10_89_2312_0 & ((~i_10_89_320_0 & ~i_10_89_1004_0 & i_10_89_2354_0 & ~i_10_89_2834_0 & ~i_10_89_3980_0) | (i_10_89_1652_0 & i_10_89_2356_0 & ~i_10_89_3647_0 & ~i_10_89_3650_0 & ~i_10_89_4288_0))))) | (i_10_89_4115_0 & ((i_10_89_1310_0 & ~i_10_89_2000_0 & ~i_10_89_2024_0 & i_10_89_4121_0) | (i_10_89_3859_0 & ~i_10_89_3986_0 & i_10_89_4117_0 & ~i_10_89_4288_0))) | (~i_10_89_4288_0 & ((i_10_89_2703_0 & i_10_89_2834_0 & ~i_10_89_3044_0) | (~i_10_89_1307_0 & ~i_10_89_1310_0 & i_10_89_2632_0 & ~i_10_89_2703_0 & ~i_10_89_3983_0))) | (~i_10_89_3983_0 & ((i_10_89_282_0 & i_10_89_287_0 & ~i_10_89_319_0 & ~i_10_89_3542_0) | (i_10_89_410_0 & i_10_89_2356_0 & ~i_10_89_3839_0))) | (i_10_89_443_0 & ~i_10_89_1238_0 & ~i_10_89_1433_0 & ~i_10_89_2719_0 & ~i_10_89_3980_0 & ~i_10_89_4121_0));
endmodule



// Benchmark "kernel_10_90" written by ABC on Sun Jul 19 10:22:32 2020

module kernel_10_90 ( 
    i_10_90_31_0, i_10_90_32_0, i_10_90_175_0, i_10_90_190_0,
    i_10_90_221_0, i_10_90_330_0, i_10_90_331_0, i_10_90_387_0,
    i_10_90_390_0, i_10_90_391_0, i_10_90_432_0, i_10_90_463_0,
    i_10_90_946_0, i_10_90_990_0, i_10_90_1037_0, i_10_90_1056_0,
    i_10_90_1081_0, i_10_90_1116_0, i_10_90_1233_0, i_10_90_1242_0,
    i_10_90_1243_0, i_10_90_1366_0, i_10_90_1432_0, i_10_90_1652_0,
    i_10_90_1654_0, i_10_90_1655_0, i_10_90_1730_0, i_10_90_1913_0,
    i_10_90_1921_0, i_10_90_1945_0, i_10_90_1949_0, i_10_90_1954_0,
    i_10_90_1992_0, i_10_90_2182_0, i_10_90_2304_0, i_10_90_2349_0,
    i_10_90_2350_0, i_10_90_2381_0, i_10_90_2449_0, i_10_90_2450_0,
    i_10_90_2466_0, i_10_90_2467_0, i_10_90_2469_0, i_10_90_2529_0,
    i_10_90_2602_0, i_10_90_2606_0, i_10_90_2629_0, i_10_90_2636_0,
    i_10_90_2701_0, i_10_90_2705_0, i_10_90_2721_0, i_10_90_2722_0,
    i_10_90_2725_0, i_10_90_2953_0, i_10_90_2979_0, i_10_90_3034_0,
    i_10_90_3035_0, i_10_90_3044_0, i_10_90_3074_0, i_10_90_3095_0,
    i_10_90_3231_0, i_10_90_3233_0, i_10_90_3277_0, i_10_90_3281_0,
    i_10_90_3312_0, i_10_90_3385_0, i_10_90_3402_0, i_10_90_3434_0,
    i_10_90_3466_0, i_10_90_3586_0, i_10_90_3587_0, i_10_90_3590_0,
    i_10_90_3610_0, i_10_90_3614_0, i_10_90_3646_0, i_10_90_3648_0,
    i_10_90_3649_0, i_10_90_3721_0, i_10_90_3839_0, i_10_90_3841_0,
    i_10_90_3852_0, i_10_90_3856_0, i_10_90_3857_0, i_10_90_3978_0,
    i_10_90_3979_0, i_10_90_3980_0, i_10_90_3982_0, i_10_90_3987_0,
    i_10_90_3991_0, i_10_90_4026_0, i_10_90_4027_0, i_10_90_4028_0,
    i_10_90_4051_0, i_10_90_4053_0, i_10_90_4266_0, i_10_90_4275_0,
    i_10_90_4276_0, i_10_90_4277_0, i_10_90_4287_0, i_10_90_4554_0,
    o_10_90_0_0  );
  input  i_10_90_31_0, i_10_90_32_0, i_10_90_175_0, i_10_90_190_0,
    i_10_90_221_0, i_10_90_330_0, i_10_90_331_0, i_10_90_387_0,
    i_10_90_390_0, i_10_90_391_0, i_10_90_432_0, i_10_90_463_0,
    i_10_90_946_0, i_10_90_990_0, i_10_90_1037_0, i_10_90_1056_0,
    i_10_90_1081_0, i_10_90_1116_0, i_10_90_1233_0, i_10_90_1242_0,
    i_10_90_1243_0, i_10_90_1366_0, i_10_90_1432_0, i_10_90_1652_0,
    i_10_90_1654_0, i_10_90_1655_0, i_10_90_1730_0, i_10_90_1913_0,
    i_10_90_1921_0, i_10_90_1945_0, i_10_90_1949_0, i_10_90_1954_0,
    i_10_90_1992_0, i_10_90_2182_0, i_10_90_2304_0, i_10_90_2349_0,
    i_10_90_2350_0, i_10_90_2381_0, i_10_90_2449_0, i_10_90_2450_0,
    i_10_90_2466_0, i_10_90_2467_0, i_10_90_2469_0, i_10_90_2529_0,
    i_10_90_2602_0, i_10_90_2606_0, i_10_90_2629_0, i_10_90_2636_0,
    i_10_90_2701_0, i_10_90_2705_0, i_10_90_2721_0, i_10_90_2722_0,
    i_10_90_2725_0, i_10_90_2953_0, i_10_90_2979_0, i_10_90_3034_0,
    i_10_90_3035_0, i_10_90_3044_0, i_10_90_3074_0, i_10_90_3095_0,
    i_10_90_3231_0, i_10_90_3233_0, i_10_90_3277_0, i_10_90_3281_0,
    i_10_90_3312_0, i_10_90_3385_0, i_10_90_3402_0, i_10_90_3434_0,
    i_10_90_3466_0, i_10_90_3586_0, i_10_90_3587_0, i_10_90_3590_0,
    i_10_90_3610_0, i_10_90_3614_0, i_10_90_3646_0, i_10_90_3648_0,
    i_10_90_3649_0, i_10_90_3721_0, i_10_90_3839_0, i_10_90_3841_0,
    i_10_90_3852_0, i_10_90_3856_0, i_10_90_3857_0, i_10_90_3978_0,
    i_10_90_3979_0, i_10_90_3980_0, i_10_90_3982_0, i_10_90_3987_0,
    i_10_90_3991_0, i_10_90_4026_0, i_10_90_4027_0, i_10_90_4028_0,
    i_10_90_4051_0, i_10_90_4053_0, i_10_90_4266_0, i_10_90_4275_0,
    i_10_90_4276_0, i_10_90_4277_0, i_10_90_4287_0, i_10_90_4554_0;
  output o_10_90_0_0;
  assign o_10_90_0_0 = 0;
endmodule



// Benchmark "kernel_10_91" written by ABC on Sun Jul 19 10:22:32 2020

module kernel_10_91 ( 
    i_10_91_173_0, i_10_91_266_0, i_10_91_283_0, i_10_91_316_0,
    i_10_91_387_0, i_10_91_438_0, i_10_91_447_0, i_10_91_578_0,
    i_10_91_697_0, i_10_91_698_0, i_10_91_733_0, i_10_91_734_0,
    i_10_91_754_0, i_10_91_928_0, i_10_91_997_0, i_10_91_1040_0,
    i_10_91_1043_0, i_10_91_1138_0, i_10_91_1167_0, i_10_91_1205_0,
    i_10_91_1234_0, i_10_91_1237_0, i_10_91_1309_0, i_10_91_1344_0,
    i_10_91_1346_0, i_10_91_1384_0, i_10_91_1403_0, i_10_91_1550_0,
    i_10_91_1552_0, i_10_91_1553_0, i_10_91_1745_0, i_10_91_1766_0,
    i_10_91_1825_0, i_10_91_1910_0, i_10_91_1958_0, i_10_91_2092_0,
    i_10_91_2159_0, i_10_91_2209_0, i_10_91_2330_0, i_10_91_2361_0,
    i_10_91_2377_0, i_10_91_2450_0, i_10_91_2452_0, i_10_91_2527_0,
    i_10_91_2539_0, i_10_91_2540_0, i_10_91_2543_0, i_10_91_2616_0,
    i_10_91_2630_0, i_10_91_2632_0, i_10_91_2660_0, i_10_91_2677_0,
    i_10_91_2714_0, i_10_91_2731_0, i_10_91_2755_0, i_10_91_2817_0,
    i_10_91_2818_0, i_10_91_2882_0, i_10_91_2920_0, i_10_91_3041_0,
    i_10_91_3047_0, i_10_91_3074_0, i_10_91_3087_0, i_10_91_3088_0,
    i_10_91_3089_0, i_10_91_3092_0, i_10_91_3198_0, i_10_91_3199_0,
    i_10_91_3280_0, i_10_91_3330_0, i_10_91_3331_0, i_10_91_3350_0,
    i_10_91_3353_0, i_10_91_3359_0, i_10_91_3404_0, i_10_91_3405_0,
    i_10_91_3503_0, i_10_91_3524_0, i_10_91_3539_0, i_10_91_3551_0,
    i_10_91_3555_0, i_10_91_3614_0, i_10_91_3859_0, i_10_91_3860_0,
    i_10_91_3899_0, i_10_91_3983_0, i_10_91_3992_0, i_10_91_4057_0,
    i_10_91_4167_0, i_10_91_4271_0, i_10_91_4282_0, i_10_91_4292_0,
    i_10_91_4376_0, i_10_91_4379_0, i_10_91_4382_0, i_10_91_4554_0,
    i_10_91_4568_0, i_10_91_4574_0, i_10_91_4576_0, i_10_91_4577_0,
    o_10_91_0_0  );
  input  i_10_91_173_0, i_10_91_266_0, i_10_91_283_0, i_10_91_316_0,
    i_10_91_387_0, i_10_91_438_0, i_10_91_447_0, i_10_91_578_0,
    i_10_91_697_0, i_10_91_698_0, i_10_91_733_0, i_10_91_734_0,
    i_10_91_754_0, i_10_91_928_0, i_10_91_997_0, i_10_91_1040_0,
    i_10_91_1043_0, i_10_91_1138_0, i_10_91_1167_0, i_10_91_1205_0,
    i_10_91_1234_0, i_10_91_1237_0, i_10_91_1309_0, i_10_91_1344_0,
    i_10_91_1346_0, i_10_91_1384_0, i_10_91_1403_0, i_10_91_1550_0,
    i_10_91_1552_0, i_10_91_1553_0, i_10_91_1745_0, i_10_91_1766_0,
    i_10_91_1825_0, i_10_91_1910_0, i_10_91_1958_0, i_10_91_2092_0,
    i_10_91_2159_0, i_10_91_2209_0, i_10_91_2330_0, i_10_91_2361_0,
    i_10_91_2377_0, i_10_91_2450_0, i_10_91_2452_0, i_10_91_2527_0,
    i_10_91_2539_0, i_10_91_2540_0, i_10_91_2543_0, i_10_91_2616_0,
    i_10_91_2630_0, i_10_91_2632_0, i_10_91_2660_0, i_10_91_2677_0,
    i_10_91_2714_0, i_10_91_2731_0, i_10_91_2755_0, i_10_91_2817_0,
    i_10_91_2818_0, i_10_91_2882_0, i_10_91_2920_0, i_10_91_3041_0,
    i_10_91_3047_0, i_10_91_3074_0, i_10_91_3087_0, i_10_91_3088_0,
    i_10_91_3089_0, i_10_91_3092_0, i_10_91_3198_0, i_10_91_3199_0,
    i_10_91_3280_0, i_10_91_3330_0, i_10_91_3331_0, i_10_91_3350_0,
    i_10_91_3353_0, i_10_91_3359_0, i_10_91_3404_0, i_10_91_3405_0,
    i_10_91_3503_0, i_10_91_3524_0, i_10_91_3539_0, i_10_91_3551_0,
    i_10_91_3555_0, i_10_91_3614_0, i_10_91_3859_0, i_10_91_3860_0,
    i_10_91_3899_0, i_10_91_3983_0, i_10_91_3992_0, i_10_91_4057_0,
    i_10_91_4167_0, i_10_91_4271_0, i_10_91_4282_0, i_10_91_4292_0,
    i_10_91_4376_0, i_10_91_4379_0, i_10_91_4382_0, i_10_91_4554_0,
    i_10_91_4568_0, i_10_91_4574_0, i_10_91_4576_0, i_10_91_4577_0;
  output o_10_91_0_0;
  assign o_10_91_0_0 = 0;
endmodule



// Benchmark "kernel_10_92" written by ABC on Sun Jul 19 10:22:33 2020

module kernel_10_92 ( 
    i_10_92_27_0, i_10_92_156_0, i_10_92_180_0, i_10_92_258_0,
    i_10_92_267_0, i_10_92_268_0, i_10_92_280_0, i_10_92_292_0,
    i_10_92_331_0, i_10_92_348_0, i_10_92_363_0, i_10_92_425_0,
    i_10_92_444_0, i_10_92_446_0, i_10_92_449_0, i_10_92_562_0,
    i_10_92_564_0, i_10_92_565_0, i_10_92_669_0, i_10_92_910_0,
    i_10_92_918_0, i_10_92_933_0, i_10_92_958_0, i_10_92_988_0,
    i_10_92_999_0, i_10_92_1000_0, i_10_92_1047_0, i_10_92_1052_0,
    i_10_92_1105_0, i_10_92_1305_0, i_10_92_1306_0, i_10_92_1311_0,
    i_10_92_1326_0, i_10_92_1457_0, i_10_92_1614_0, i_10_92_1615_0,
    i_10_92_1684_0, i_10_92_1685_0, i_10_92_1818_0, i_10_92_1899_0,
    i_10_92_1942_0, i_10_92_1948_0, i_10_92_1992_0, i_10_92_2001_0,
    i_10_92_2020_0, i_10_92_2079_0, i_10_92_2142_0, i_10_92_2182_0,
    i_10_92_2186_0, i_10_92_2239_0, i_10_92_2326_0, i_10_92_2350_0,
    i_10_92_2351_0, i_10_92_2352_0, i_10_92_2409_0, i_10_92_2452_0,
    i_10_92_2469_0, i_10_92_2582_0, i_10_92_2605_0, i_10_92_2611_0,
    i_10_92_2614_0, i_10_92_2615_0, i_10_92_2703_0, i_10_92_2754_0,
    i_10_92_2787_0, i_10_92_3009_0, i_10_92_3039_0, i_10_92_3069_0,
    i_10_92_3090_0, i_10_92_3195_0, i_10_92_3283_0, i_10_92_3297_0,
    i_10_92_3301_0, i_10_92_3325_0, i_10_92_3448_0, i_10_92_3495_0,
    i_10_92_3499_0, i_10_92_3558_0, i_10_92_3561_0, i_10_92_3588_0,
    i_10_92_3589_0, i_10_92_3609_0, i_10_92_3610_0, i_10_92_3637_0,
    i_10_92_3695_0, i_10_92_3699_0, i_10_92_3852_0, i_10_92_3882_0,
    i_10_92_3945_0, i_10_92_3982_0, i_10_92_4027_0, i_10_92_4050_0,
    i_10_92_4067_0, i_10_92_4186_0, i_10_92_4293_0, i_10_92_4372_0,
    i_10_92_4373_0, i_10_92_4449_0, i_10_92_4457_0, i_10_92_4530_0,
    o_10_92_0_0  );
  input  i_10_92_27_0, i_10_92_156_0, i_10_92_180_0, i_10_92_258_0,
    i_10_92_267_0, i_10_92_268_0, i_10_92_280_0, i_10_92_292_0,
    i_10_92_331_0, i_10_92_348_0, i_10_92_363_0, i_10_92_425_0,
    i_10_92_444_0, i_10_92_446_0, i_10_92_449_0, i_10_92_562_0,
    i_10_92_564_0, i_10_92_565_0, i_10_92_669_0, i_10_92_910_0,
    i_10_92_918_0, i_10_92_933_0, i_10_92_958_0, i_10_92_988_0,
    i_10_92_999_0, i_10_92_1000_0, i_10_92_1047_0, i_10_92_1052_0,
    i_10_92_1105_0, i_10_92_1305_0, i_10_92_1306_0, i_10_92_1311_0,
    i_10_92_1326_0, i_10_92_1457_0, i_10_92_1614_0, i_10_92_1615_0,
    i_10_92_1684_0, i_10_92_1685_0, i_10_92_1818_0, i_10_92_1899_0,
    i_10_92_1942_0, i_10_92_1948_0, i_10_92_1992_0, i_10_92_2001_0,
    i_10_92_2020_0, i_10_92_2079_0, i_10_92_2142_0, i_10_92_2182_0,
    i_10_92_2186_0, i_10_92_2239_0, i_10_92_2326_0, i_10_92_2350_0,
    i_10_92_2351_0, i_10_92_2352_0, i_10_92_2409_0, i_10_92_2452_0,
    i_10_92_2469_0, i_10_92_2582_0, i_10_92_2605_0, i_10_92_2611_0,
    i_10_92_2614_0, i_10_92_2615_0, i_10_92_2703_0, i_10_92_2754_0,
    i_10_92_2787_0, i_10_92_3009_0, i_10_92_3039_0, i_10_92_3069_0,
    i_10_92_3090_0, i_10_92_3195_0, i_10_92_3283_0, i_10_92_3297_0,
    i_10_92_3301_0, i_10_92_3325_0, i_10_92_3448_0, i_10_92_3495_0,
    i_10_92_3499_0, i_10_92_3558_0, i_10_92_3561_0, i_10_92_3588_0,
    i_10_92_3589_0, i_10_92_3609_0, i_10_92_3610_0, i_10_92_3637_0,
    i_10_92_3695_0, i_10_92_3699_0, i_10_92_3852_0, i_10_92_3882_0,
    i_10_92_3945_0, i_10_92_3982_0, i_10_92_4027_0, i_10_92_4050_0,
    i_10_92_4067_0, i_10_92_4186_0, i_10_92_4293_0, i_10_92_4372_0,
    i_10_92_4373_0, i_10_92_4449_0, i_10_92_4457_0, i_10_92_4530_0;
  output o_10_92_0_0;
  assign o_10_92_0_0 = 0;
endmodule



// Benchmark "kernel_10_93" written by ABC on Sun Jul 19 10:22:35 2020

module kernel_10_93 ( 
    i_10_93_82_0, i_10_93_221_0, i_10_93_281_0, i_10_93_283_0,
    i_10_93_409_0, i_10_93_423_0, i_10_93_424_0, i_10_93_446_0,
    i_10_93_448_0, i_10_93_495_0, i_10_93_505_0, i_10_93_513_0,
    i_10_93_794_0, i_10_93_964_0, i_10_93_1236_0, i_10_93_1240_0,
    i_10_93_1260_0, i_10_93_1309_0, i_10_93_1342_0, i_10_93_1359_0,
    i_10_93_1377_0, i_10_93_1444_0, i_10_93_1446_0, i_10_93_1450_0,
    i_10_93_1540_0, i_10_93_1582_0, i_10_93_1655_0, i_10_93_1683_0,
    i_10_93_1819_0, i_10_93_1820_0, i_10_93_1821_0, i_10_93_1913_0,
    i_10_93_1944_0, i_10_93_1945_0, i_10_93_1989_0, i_10_93_2026_0,
    i_10_93_2331_0, i_10_93_2353_0, i_10_93_2364_0, i_10_93_2377_0,
    i_10_93_2380_0, i_10_93_2403_0, i_10_93_2404_0, i_10_93_2502_0,
    i_10_93_2503_0, i_10_93_2504_0, i_10_93_2628_0, i_10_93_2632_0,
    i_10_93_2637_0, i_10_93_2638_0, i_10_93_2655_0, i_10_93_2658_0,
    i_10_93_2673_0, i_10_93_2674_0, i_10_93_2675_0, i_10_93_2711_0,
    i_10_93_2718_0, i_10_93_2722_0, i_10_93_2724_0, i_10_93_2727_0,
    i_10_93_2728_0, i_10_93_2781_0, i_10_93_2827_0, i_10_93_2830_0,
    i_10_93_2831_0, i_10_93_2881_0, i_10_93_2920_0, i_10_93_2979_0,
    i_10_93_2980_0, i_10_93_3042_0, i_10_93_3070_0, i_10_93_3073_0,
    i_10_93_3076_0, i_10_93_3151_0, i_10_93_3195_0, i_10_93_3198_0,
    i_10_93_3385_0, i_10_93_3586_0, i_10_93_3609_0, i_10_93_3780_0,
    i_10_93_3781_0, i_10_93_3835_0, i_10_93_3837_0, i_10_93_3838_0,
    i_10_93_3841_0, i_10_93_3843_0, i_10_93_3852_0, i_10_93_3889_0,
    i_10_93_3979_0, i_10_93_3980_0, i_10_93_4054_0, i_10_93_4118_0,
    i_10_93_4122_0, i_10_93_4123_0, i_10_93_4126_0, i_10_93_4289_0,
    i_10_93_4564_0, i_10_93_4567_0, i_10_93_4568_0, i_10_93_4570_0,
    o_10_93_0_0  );
  input  i_10_93_82_0, i_10_93_221_0, i_10_93_281_0, i_10_93_283_0,
    i_10_93_409_0, i_10_93_423_0, i_10_93_424_0, i_10_93_446_0,
    i_10_93_448_0, i_10_93_495_0, i_10_93_505_0, i_10_93_513_0,
    i_10_93_794_0, i_10_93_964_0, i_10_93_1236_0, i_10_93_1240_0,
    i_10_93_1260_0, i_10_93_1309_0, i_10_93_1342_0, i_10_93_1359_0,
    i_10_93_1377_0, i_10_93_1444_0, i_10_93_1446_0, i_10_93_1450_0,
    i_10_93_1540_0, i_10_93_1582_0, i_10_93_1655_0, i_10_93_1683_0,
    i_10_93_1819_0, i_10_93_1820_0, i_10_93_1821_0, i_10_93_1913_0,
    i_10_93_1944_0, i_10_93_1945_0, i_10_93_1989_0, i_10_93_2026_0,
    i_10_93_2331_0, i_10_93_2353_0, i_10_93_2364_0, i_10_93_2377_0,
    i_10_93_2380_0, i_10_93_2403_0, i_10_93_2404_0, i_10_93_2502_0,
    i_10_93_2503_0, i_10_93_2504_0, i_10_93_2628_0, i_10_93_2632_0,
    i_10_93_2637_0, i_10_93_2638_0, i_10_93_2655_0, i_10_93_2658_0,
    i_10_93_2673_0, i_10_93_2674_0, i_10_93_2675_0, i_10_93_2711_0,
    i_10_93_2718_0, i_10_93_2722_0, i_10_93_2724_0, i_10_93_2727_0,
    i_10_93_2728_0, i_10_93_2781_0, i_10_93_2827_0, i_10_93_2830_0,
    i_10_93_2831_0, i_10_93_2881_0, i_10_93_2920_0, i_10_93_2979_0,
    i_10_93_2980_0, i_10_93_3042_0, i_10_93_3070_0, i_10_93_3073_0,
    i_10_93_3076_0, i_10_93_3151_0, i_10_93_3195_0, i_10_93_3198_0,
    i_10_93_3385_0, i_10_93_3586_0, i_10_93_3609_0, i_10_93_3780_0,
    i_10_93_3781_0, i_10_93_3835_0, i_10_93_3837_0, i_10_93_3838_0,
    i_10_93_3841_0, i_10_93_3843_0, i_10_93_3852_0, i_10_93_3889_0,
    i_10_93_3979_0, i_10_93_3980_0, i_10_93_4054_0, i_10_93_4118_0,
    i_10_93_4122_0, i_10_93_4123_0, i_10_93_4126_0, i_10_93_4289_0,
    i_10_93_4564_0, i_10_93_4567_0, i_10_93_4568_0, i_10_93_4570_0;
  output o_10_93_0_0;
  assign o_10_93_0_0 = ~((~i_10_93_409_0 & ~i_10_93_3843_0 & ((~i_10_93_513_0 & ~i_10_93_1540_0 & ~i_10_93_2364_0 & ~i_10_93_2403_0 & ~i_10_93_2504_0 & ~i_10_93_2637_0 & ~i_10_93_2638_0 & ~i_10_93_3195_0) | (~i_10_93_424_0 & ~i_10_93_1260_0 & ~i_10_93_1446_0 & ~i_10_93_1913_0 & ~i_10_93_1944_0 & ~i_10_93_1945_0 & ~i_10_93_2377_0 & ~i_10_93_2502_0 & ~i_10_93_3889_0 & ~i_10_93_4054_0))) | (~i_10_93_1444_0 & ((~i_10_93_2718_0 & ((~i_10_93_424_0 & ((~i_10_93_423_0 & ~i_10_93_1913_0 & ~i_10_93_1945_0 & ~i_10_93_2380_0 & ~i_10_93_2728_0 & ~i_10_93_3042_0 & ~i_10_93_4122_0) | (~i_10_93_1446_0 & ~i_10_93_1944_0 & ~i_10_93_2502_0 & ~i_10_93_2503_0 & ~i_10_93_2628_0 & ~i_10_93_3837_0 & ~i_10_93_4567_0))) | (i_10_93_794_0 & ~i_10_93_1683_0 & ~i_10_93_1945_0 & ~i_10_93_2377_0 & ~i_10_93_2504_0 & ~i_10_93_2658_0 & ~i_10_93_2673_0))) | (~i_10_93_513_0 & ~i_10_93_1236_0 & ~i_10_93_1683_0 & ~i_10_93_1989_0 & ~i_10_93_2404_0 & ~i_10_93_2502_0 & ~i_10_93_2637_0 & ~i_10_93_2827_0) | (~i_10_93_82_0 & ~i_10_93_964_0 & ~i_10_93_1260_0 & ~i_10_93_1582_0 & ~i_10_93_2380_0 & ~i_10_93_2504_0 & ~i_10_93_2673_0 & ~i_10_93_2980_0 & ~i_10_93_3042_0 & ~i_10_93_4568_0))) | (~i_10_93_513_0 & ((~i_10_93_446_0 & i_10_93_2632_0 & ~i_10_93_2637_0 & ~i_10_93_2673_0 & ~i_10_93_2674_0 & ~i_10_93_2724_0 & ~i_10_93_2727_0) | (~i_10_93_1240_0 & ~i_10_93_2404_0 & ~i_10_93_2502_0 & ~i_10_93_2658_0 & ~i_10_93_2831_0))) | (~i_10_93_1944_0 & ((~i_10_93_1359_0 & ((~i_10_93_2658_0 & ((~i_10_93_446_0 & ((~i_10_93_964_0 & ~i_10_93_1236_0 & ~i_10_93_1309_0 & ~i_10_93_2504_0 & ~i_10_93_2637_0 & ~i_10_93_2331_0 & ~i_10_93_2403_0) | (~i_10_93_1819_0 & ~i_10_93_1945_0 & i_10_93_2632_0 & ~i_10_93_2830_0 & ~i_10_93_3586_0))) | (~i_10_93_283_0 & ~i_10_93_2380_0 & ~i_10_93_2404_0 & ~i_10_93_2655_0 & i_10_93_3889_0))) | (~i_10_93_964_0 & ~i_10_93_1236_0 & ~i_10_93_1260_0 & ~i_10_93_2353_0 & ~i_10_93_2377_0 & ~i_10_93_2502_0 & ~i_10_93_2674_0 & ~i_10_93_2711_0))) | (~i_10_93_2403_0 & ~i_10_93_2637_0 & ~i_10_93_2722_0 & ~i_10_93_2979_0 & i_10_93_3838_0))) | (~i_10_93_964_0 & ((~i_10_93_2404_0 & ~i_10_93_2658_0 & ~i_10_93_2673_0 & ~i_10_93_2781_0 & ~i_10_93_2920_0 & ~i_10_93_3586_0 & ~i_10_93_4123_0) | (~i_10_93_1945_0 & ~i_10_93_2502_0 & ~i_10_93_2638_0 & ~i_10_93_2674_0 & ~i_10_93_2979_0 & i_10_93_4289_0))) | (~i_10_93_1446_0 & ((~i_10_93_2403_0 & ~i_10_93_2673_0 & ~i_10_93_2728_0 & i_10_93_3609_0) | (~i_10_93_2637_0 & ~i_10_93_2674_0 & ~i_10_93_2675_0 & ~i_10_93_2727_0 & i_10_93_3385_0 & ~i_10_93_4568_0))) | (i_10_93_2632_0 & ~i_10_93_2658_0 & i_10_93_3609_0) | (~i_10_93_1240_0 & ~i_10_93_2728_0 & ~i_10_93_2980_0 & i_10_93_3835_0) | (~i_10_93_1913_0 & i_10_93_1945_0 & ~i_10_93_2503_0 & i_10_93_2504_0 & ~i_10_93_2920_0 & ~i_10_93_3979_0) | (~i_10_93_2674_0 & i_10_93_2675_0 & i_10_93_3979_0 & ~i_10_93_4567_0));
endmodule



// Benchmark "kernel_10_94" written by ABC on Sun Jul 19 10:22:36 2020

module kernel_10_94 ( 
    i_10_94_12_0, i_10_94_63_0, i_10_94_64_0, i_10_94_77_0, i_10_94_172_0,
    i_10_94_174_0, i_10_94_175_0, i_10_94_208_0, i_10_94_223_0,
    i_10_94_244_0, i_10_94_286_0, i_10_94_315_0, i_10_94_318_0,
    i_10_94_406_0, i_10_94_594_0, i_10_94_639_0, i_10_94_733_0,
    i_10_94_891_0, i_10_94_946_0, i_10_94_999_0, i_10_94_1000_0,
    i_10_94_1041_0, i_10_94_1060_0, i_10_94_1174_0, i_10_94_1239_0,
    i_10_94_1241_0, i_10_94_1242_0, i_10_94_1244_0, i_10_94_1264_0,
    i_10_94_1267_0, i_10_94_1268_0, i_10_94_1367_0, i_10_94_1382_0,
    i_10_94_1545_0, i_10_94_1579_0, i_10_94_1593_0, i_10_94_1611_0,
    i_10_94_1633_0, i_10_94_1653_0, i_10_94_1654_0, i_10_94_1696_0,
    i_10_94_1883_0, i_10_94_1912_0, i_10_94_1919_0, i_10_94_1953_0,
    i_10_94_1989_0, i_10_94_1998_0, i_10_94_2106_0, i_10_94_2203_0,
    i_10_94_2236_0, i_10_94_2245_0, i_10_94_2246_0, i_10_94_2254_0,
    i_10_94_2448_0, i_10_94_2459_0, i_10_94_2475_0, i_10_94_2502_0,
    i_10_94_2514_0, i_10_94_2541_0, i_10_94_2565_0, i_10_94_2611_0,
    i_10_94_2633_0, i_10_94_2659_0, i_10_94_2662_0, i_10_94_2663_0,
    i_10_94_2676_0, i_10_94_2730_0, i_10_94_2782_0, i_10_94_2807_0,
    i_10_94_2882_0, i_10_94_3198_0, i_10_94_3202_0, i_10_94_3454_0,
    i_10_94_3537_0, i_10_94_3540_0, i_10_94_3618_0, i_10_94_3700_0,
    i_10_94_3771_0, i_10_94_3847_0, i_10_94_3852_0, i_10_94_3854_0,
    i_10_94_3857_0, i_10_94_3881_0, i_10_94_3897_0, i_10_94_3901_0,
    i_10_94_3978_0, i_10_94_4118_0, i_10_94_4150_0, i_10_94_4152_0,
    i_10_94_4153_0, i_10_94_4155_0, i_10_94_4158_0, i_10_94_4173_0,
    i_10_94_4174_0, i_10_94_4213_0, i_10_94_4266_0, i_10_94_4410_0,
    i_10_94_4431_0, i_10_94_4438_0, i_10_94_4528_0,
    o_10_94_0_0  );
  input  i_10_94_12_0, i_10_94_63_0, i_10_94_64_0, i_10_94_77_0,
    i_10_94_172_0, i_10_94_174_0, i_10_94_175_0, i_10_94_208_0,
    i_10_94_223_0, i_10_94_244_0, i_10_94_286_0, i_10_94_315_0,
    i_10_94_318_0, i_10_94_406_0, i_10_94_594_0, i_10_94_639_0,
    i_10_94_733_0, i_10_94_891_0, i_10_94_946_0, i_10_94_999_0,
    i_10_94_1000_0, i_10_94_1041_0, i_10_94_1060_0, i_10_94_1174_0,
    i_10_94_1239_0, i_10_94_1241_0, i_10_94_1242_0, i_10_94_1244_0,
    i_10_94_1264_0, i_10_94_1267_0, i_10_94_1268_0, i_10_94_1367_0,
    i_10_94_1382_0, i_10_94_1545_0, i_10_94_1579_0, i_10_94_1593_0,
    i_10_94_1611_0, i_10_94_1633_0, i_10_94_1653_0, i_10_94_1654_0,
    i_10_94_1696_0, i_10_94_1883_0, i_10_94_1912_0, i_10_94_1919_0,
    i_10_94_1953_0, i_10_94_1989_0, i_10_94_1998_0, i_10_94_2106_0,
    i_10_94_2203_0, i_10_94_2236_0, i_10_94_2245_0, i_10_94_2246_0,
    i_10_94_2254_0, i_10_94_2448_0, i_10_94_2459_0, i_10_94_2475_0,
    i_10_94_2502_0, i_10_94_2514_0, i_10_94_2541_0, i_10_94_2565_0,
    i_10_94_2611_0, i_10_94_2633_0, i_10_94_2659_0, i_10_94_2662_0,
    i_10_94_2663_0, i_10_94_2676_0, i_10_94_2730_0, i_10_94_2782_0,
    i_10_94_2807_0, i_10_94_2882_0, i_10_94_3198_0, i_10_94_3202_0,
    i_10_94_3454_0, i_10_94_3537_0, i_10_94_3540_0, i_10_94_3618_0,
    i_10_94_3700_0, i_10_94_3771_0, i_10_94_3847_0, i_10_94_3852_0,
    i_10_94_3854_0, i_10_94_3857_0, i_10_94_3881_0, i_10_94_3897_0,
    i_10_94_3901_0, i_10_94_3978_0, i_10_94_4118_0, i_10_94_4150_0,
    i_10_94_4152_0, i_10_94_4153_0, i_10_94_4155_0, i_10_94_4158_0,
    i_10_94_4173_0, i_10_94_4174_0, i_10_94_4213_0, i_10_94_4266_0,
    i_10_94_4410_0, i_10_94_4431_0, i_10_94_4438_0, i_10_94_4528_0;
  output o_10_94_0_0;
  assign o_10_94_0_0 = 0;
endmodule



// Benchmark "kernel_10_95" written by ABC on Sun Jul 19 10:22:36 2020

module kernel_10_95 ( 
    i_10_95_146_0, i_10_95_280_0, i_10_95_315_0, i_10_95_316_0,
    i_10_95_318_0, i_10_95_319_0, i_10_95_406_0, i_10_95_411_0,
    i_10_95_412_0, i_10_95_427_0, i_10_95_441_0, i_10_95_442_0,
    i_10_95_444_0, i_10_95_445_0, i_10_95_448_0, i_10_95_460_0,
    i_10_95_461_0, i_10_95_462_0, i_10_95_588_0, i_10_95_712_0,
    i_10_95_715_0, i_10_95_716_0, i_10_95_747_0, i_10_95_793_0,
    i_10_95_795_0, i_10_95_796_0, i_10_95_798_0, i_10_95_828_0,
    i_10_95_927_0, i_10_95_963_0, i_10_95_966_0, i_10_95_967_0,
    i_10_95_993_0, i_10_95_1002_0, i_10_95_1003_0, i_10_95_1116_0,
    i_10_95_1234_0, i_10_95_1235_0, i_10_95_1341_0, i_10_95_1344_0,
    i_10_95_1444_0, i_10_95_1649_0, i_10_95_1650_0, i_10_95_1651_0,
    i_10_95_1652_0, i_10_95_1685_0, i_10_95_1686_0, i_10_95_1687_0,
    i_10_95_1818_0, i_10_95_1821_0, i_10_95_1945_0, i_10_95_1949_0,
    i_10_95_2154_0, i_10_95_2181_0, i_10_95_2334_0, i_10_95_2335_0,
    i_10_95_2337_0, i_10_95_2338_0, i_10_95_2350_0, i_10_95_2379_0,
    i_10_95_2383_0, i_10_95_2407_0, i_10_95_2449_0, i_10_95_2451_0,
    i_10_95_2452_0, i_10_95_2473_0, i_10_95_2474_0, i_10_95_2629_0,
    i_10_95_2631_0, i_10_95_2632_0, i_10_95_2634_0, i_10_95_2658_0,
    i_10_95_2661_0, i_10_95_2662_0, i_10_95_2712_0, i_10_95_2733_0,
    i_10_95_2734_0, i_10_95_2784_0, i_10_95_2826_0, i_10_95_2880_0,
    i_10_95_2917_0, i_10_95_2984_0, i_10_95_3039_0, i_10_95_3270_0,
    i_10_95_3387_0, i_10_95_3402_0, i_10_95_3405_0, i_10_95_3582_0,
    i_10_95_3583_0, i_10_95_3585_0, i_10_95_3586_0, i_10_95_3589_0,
    i_10_95_3590_0, i_10_95_3613_0, i_10_95_3727_0, i_10_95_3787_0,
    i_10_95_4266_0, i_10_95_4284_0, i_10_95_4285_0, i_10_95_4459_0,
    o_10_95_0_0  );
  input  i_10_95_146_0, i_10_95_280_0, i_10_95_315_0, i_10_95_316_0,
    i_10_95_318_0, i_10_95_319_0, i_10_95_406_0, i_10_95_411_0,
    i_10_95_412_0, i_10_95_427_0, i_10_95_441_0, i_10_95_442_0,
    i_10_95_444_0, i_10_95_445_0, i_10_95_448_0, i_10_95_460_0,
    i_10_95_461_0, i_10_95_462_0, i_10_95_588_0, i_10_95_712_0,
    i_10_95_715_0, i_10_95_716_0, i_10_95_747_0, i_10_95_793_0,
    i_10_95_795_0, i_10_95_796_0, i_10_95_798_0, i_10_95_828_0,
    i_10_95_927_0, i_10_95_963_0, i_10_95_966_0, i_10_95_967_0,
    i_10_95_993_0, i_10_95_1002_0, i_10_95_1003_0, i_10_95_1116_0,
    i_10_95_1234_0, i_10_95_1235_0, i_10_95_1341_0, i_10_95_1344_0,
    i_10_95_1444_0, i_10_95_1649_0, i_10_95_1650_0, i_10_95_1651_0,
    i_10_95_1652_0, i_10_95_1685_0, i_10_95_1686_0, i_10_95_1687_0,
    i_10_95_1818_0, i_10_95_1821_0, i_10_95_1945_0, i_10_95_1949_0,
    i_10_95_2154_0, i_10_95_2181_0, i_10_95_2334_0, i_10_95_2335_0,
    i_10_95_2337_0, i_10_95_2338_0, i_10_95_2350_0, i_10_95_2379_0,
    i_10_95_2383_0, i_10_95_2407_0, i_10_95_2449_0, i_10_95_2451_0,
    i_10_95_2452_0, i_10_95_2473_0, i_10_95_2474_0, i_10_95_2629_0,
    i_10_95_2631_0, i_10_95_2632_0, i_10_95_2634_0, i_10_95_2658_0,
    i_10_95_2661_0, i_10_95_2662_0, i_10_95_2712_0, i_10_95_2733_0,
    i_10_95_2734_0, i_10_95_2784_0, i_10_95_2826_0, i_10_95_2880_0,
    i_10_95_2917_0, i_10_95_2984_0, i_10_95_3039_0, i_10_95_3270_0,
    i_10_95_3387_0, i_10_95_3402_0, i_10_95_3405_0, i_10_95_3582_0,
    i_10_95_3583_0, i_10_95_3585_0, i_10_95_3586_0, i_10_95_3589_0,
    i_10_95_3590_0, i_10_95_3613_0, i_10_95_3727_0, i_10_95_3787_0,
    i_10_95_4266_0, i_10_95_4284_0, i_10_95_4285_0, i_10_95_4459_0;
  output o_10_95_0_0;
  assign o_10_95_0_0 = 0;
endmodule



// Benchmark "kernel_10_96" written by ABC on Sun Jul 19 10:22:38 2020

module kernel_10_96 ( 
    i_10_96_174_0, i_10_96_175_0, i_10_96_176_0, i_10_96_177_0,
    i_10_96_221_0, i_10_96_224_0, i_10_96_283_0, i_10_96_328_0,
    i_10_96_329_0, i_10_96_331_0, i_10_96_391_0, i_10_96_408_0,
    i_10_96_410_0, i_10_96_428_0, i_10_96_797_0, i_10_96_898_0,
    i_10_96_1236_0, i_10_96_1238_0, i_10_96_1544_0, i_10_96_1552_0,
    i_10_96_1555_0, i_10_96_1579_0, i_10_96_1650_0, i_10_96_1655_0,
    i_10_96_1690_0, i_10_96_1769_0, i_10_96_1821_0, i_10_96_1822_0,
    i_10_96_1823_0, i_10_96_1945_0, i_10_96_1997_0, i_10_96_2024_0,
    i_10_96_2026_0, i_10_96_2311_0, i_10_96_2352_0, i_10_96_2353_0,
    i_10_96_2354_0, i_10_96_2356_0, i_10_96_2410_0, i_10_96_2453_0,
    i_10_96_2467_0, i_10_96_2468_0, i_10_96_2473_0, i_10_96_2603_0,
    i_10_96_2631_0, i_10_96_2632_0, i_10_96_2633_0, i_10_96_2656_0,
    i_10_96_2680_0, i_10_96_2706_0, i_10_96_2707_0, i_10_96_2783_0,
    i_10_96_2785_0, i_10_96_2786_0, i_10_96_2827_0, i_10_96_2828_0,
    i_10_96_2830_0, i_10_96_2920_0, i_10_96_2923_0, i_10_96_2924_0,
    i_10_96_3038_0, i_10_96_3044_0, i_10_96_3152_0, i_10_96_3153_0,
    i_10_96_3156_0, i_10_96_3157_0, i_10_96_3201_0, i_10_96_3387_0,
    i_10_96_3389_0, i_10_96_3583_0, i_10_96_3584_0, i_10_96_3612_0,
    i_10_96_3613_0, i_10_96_3614_0, i_10_96_3844_0, i_10_96_3846_0,
    i_10_96_3847_0, i_10_96_3848_0, i_10_96_3851_0, i_10_96_3852_0,
    i_10_96_3856_0, i_10_96_3991_0, i_10_96_3992_0, i_10_96_4119_0,
    i_10_96_4122_0, i_10_96_4125_0, i_10_96_4129_0, i_10_96_4130_0,
    i_10_96_4269_0, i_10_96_4270_0, i_10_96_4271_0, i_10_96_4276_0,
    i_10_96_4277_0, i_10_96_4286_0, i_10_96_4288_0, i_10_96_4289_0,
    i_10_96_4563_0, i_10_96_4564_0, i_10_96_4567_0, i_10_96_4568_0,
    o_10_96_0_0  );
  input  i_10_96_174_0, i_10_96_175_0, i_10_96_176_0, i_10_96_177_0,
    i_10_96_221_0, i_10_96_224_0, i_10_96_283_0, i_10_96_328_0,
    i_10_96_329_0, i_10_96_331_0, i_10_96_391_0, i_10_96_408_0,
    i_10_96_410_0, i_10_96_428_0, i_10_96_797_0, i_10_96_898_0,
    i_10_96_1236_0, i_10_96_1238_0, i_10_96_1544_0, i_10_96_1552_0,
    i_10_96_1555_0, i_10_96_1579_0, i_10_96_1650_0, i_10_96_1655_0,
    i_10_96_1690_0, i_10_96_1769_0, i_10_96_1821_0, i_10_96_1822_0,
    i_10_96_1823_0, i_10_96_1945_0, i_10_96_1997_0, i_10_96_2024_0,
    i_10_96_2026_0, i_10_96_2311_0, i_10_96_2352_0, i_10_96_2353_0,
    i_10_96_2354_0, i_10_96_2356_0, i_10_96_2410_0, i_10_96_2453_0,
    i_10_96_2467_0, i_10_96_2468_0, i_10_96_2473_0, i_10_96_2603_0,
    i_10_96_2631_0, i_10_96_2632_0, i_10_96_2633_0, i_10_96_2656_0,
    i_10_96_2680_0, i_10_96_2706_0, i_10_96_2707_0, i_10_96_2783_0,
    i_10_96_2785_0, i_10_96_2786_0, i_10_96_2827_0, i_10_96_2828_0,
    i_10_96_2830_0, i_10_96_2920_0, i_10_96_2923_0, i_10_96_2924_0,
    i_10_96_3038_0, i_10_96_3044_0, i_10_96_3152_0, i_10_96_3153_0,
    i_10_96_3156_0, i_10_96_3157_0, i_10_96_3201_0, i_10_96_3387_0,
    i_10_96_3389_0, i_10_96_3583_0, i_10_96_3584_0, i_10_96_3612_0,
    i_10_96_3613_0, i_10_96_3614_0, i_10_96_3844_0, i_10_96_3846_0,
    i_10_96_3847_0, i_10_96_3848_0, i_10_96_3851_0, i_10_96_3852_0,
    i_10_96_3856_0, i_10_96_3991_0, i_10_96_3992_0, i_10_96_4119_0,
    i_10_96_4122_0, i_10_96_4125_0, i_10_96_4129_0, i_10_96_4130_0,
    i_10_96_4269_0, i_10_96_4270_0, i_10_96_4271_0, i_10_96_4276_0,
    i_10_96_4277_0, i_10_96_4286_0, i_10_96_4288_0, i_10_96_4289_0,
    i_10_96_4563_0, i_10_96_4564_0, i_10_96_4567_0, i_10_96_4568_0;
  output o_10_96_0_0;
  assign o_10_96_0_0 = ~((~i_10_96_797_0 & ((~i_10_96_1650_0 & ~i_10_96_1655_0 & i_10_96_1822_0 & ~i_10_96_2468_0 & ~i_10_96_2473_0 & ~i_10_96_2786_0 & ~i_10_96_2923_0 & ~i_10_96_3038_0 & ~i_10_96_3852_0) | (i_10_96_1555_0 & ~i_10_96_3612_0 & ~i_10_96_4288_0))) | (~i_10_96_176_0 & ((~i_10_96_175_0 & ((~i_10_96_1823_0 & ~i_10_96_1997_0 & ~i_10_96_2656_0 & ~i_10_96_2920_0) | (~i_10_96_1236_0 & ~i_10_96_1945_0 & i_10_96_2785_0 & ~i_10_96_2828_0 & ~i_10_96_4130_0))) | (~i_10_96_428_0 & ~i_10_96_1236_0 & ~i_10_96_1238_0 & ~i_10_96_2631_0 & i_10_96_2920_0 & i_10_96_2923_0 & ~i_10_96_3851_0) | (~i_10_96_1650_0 & ~i_10_96_1821_0 & ~i_10_96_1945_0 & ~i_10_96_1997_0 & ~i_10_96_2024_0 & ~i_10_96_2453_0 & ~i_10_96_2786_0 & ~i_10_96_3584_0 & ~i_10_96_4122_0))) | (i_10_96_1579_0 & ((~i_10_96_175_0 & i_10_96_1544_0 & i_10_96_1650_0) | (~i_10_96_1655_0 & i_10_96_2632_0))) | (~i_10_96_1579_0 & ((i_10_96_1650_0 & i_10_96_1821_0 & ~i_10_96_3583_0 & i_10_96_3852_0) | (~i_10_96_175_0 & ~i_10_96_1822_0 & ~i_10_96_1823_0 & ~i_10_96_2707_0 & ~i_10_96_3613_0 & ~i_10_96_3852_0 & ~i_10_96_4130_0))) | (~i_10_96_410_0 & ((~i_10_96_4130_0 & ((~i_10_96_175_0 & ~i_10_96_2024_0 & ((~i_10_96_2467_0 & ~i_10_96_2783_0 & ~i_10_96_3856_0) | (~i_10_96_221_0 & ~i_10_96_898_0 & ~i_10_96_2468_0 & ~i_10_96_3583_0 & ~i_10_96_4567_0))) | (~i_10_96_2783_0 & ~i_10_96_3612_0 & i_10_96_3852_0 & i_10_96_3856_0))) | (~i_10_96_2783_0 & ((~i_10_96_283_0 & ~i_10_96_1544_0 & i_10_96_1823_0 & ~i_10_96_2467_0 & ~i_10_96_2707_0 & ~i_10_96_2786_0 & ~i_10_96_2920_0 & ~i_10_96_2923_0) | (i_10_96_2633_0 & i_10_96_2656_0 & ~i_10_96_3844_0 & ~i_10_96_4289_0))) | (~i_10_96_1945_0 & ~i_10_96_2311_0 & i_10_96_2631_0 & ~i_10_96_2920_0 & i_10_96_3856_0) | (~i_10_96_221_0 & ~i_10_96_408_0 & ~i_10_96_1238_0 & ~i_10_96_3583_0 & ~i_10_96_3614_0 & ~i_10_96_4129_0))) | (~i_10_96_1238_0 & ((~i_10_96_174_0 & ~i_10_96_224_0 & ~i_10_96_1823_0 & ~i_10_96_1945_0 & ~i_10_96_2468_0 & ~i_10_96_2786_0 & i_10_96_3613_0) | (~i_10_96_3583_0 & i_10_96_4269_0))) | (~i_10_96_1655_0 & ((i_10_96_2631_0 & ~i_10_96_2783_0 & ~i_10_96_2920_0) | (~i_10_96_224_0 & i_10_96_391_0 & ~i_10_96_1821_0 & ~i_10_96_3614_0 & ~i_10_96_4130_0))) | (~i_10_96_224_0 & ((~i_10_96_2024_0 & i_10_96_2354_0 & ~i_10_96_2467_0 & ~i_10_96_2828_0 & ~i_10_96_3613_0) | (~i_10_96_1823_0 & ~i_10_96_2453_0 & ~i_10_96_2786_0 & ~i_10_96_3044_0 & ~i_10_96_3584_0 & i_10_96_4125_0))) | (i_10_96_391_0 & (~i_10_96_3584_0 | (i_10_96_4270_0 & i_10_96_4288_0))) | (~i_10_96_1769_0 & ~i_10_96_2467_0 & ((~i_10_96_2603_0 & ~i_10_96_2785_0 & ~i_10_96_2830_0 & ~i_10_96_3584_0 & ~i_10_96_3612_0 & ~i_10_96_3992_0 & ~i_10_96_4129_0 & ~i_10_96_4130_0) | (~i_10_96_408_0 & ~i_10_96_3044_0 & i_10_96_3844_0 & ~i_10_96_4286_0 & ~i_10_96_4288_0))) | (~i_10_96_408_0 & ((~i_10_96_177_0 & ~i_10_96_1822_0 & ~i_10_96_1823_0 & ~i_10_96_2473_0 & ~i_10_96_2783_0 & ~i_10_96_2785_0 & ~i_10_96_3614_0 & ~i_10_96_4125_0) | (i_10_96_2830_0 & i_10_96_4567_0))) | (i_10_96_1821_0 & ((~i_10_96_2352_0 & ~i_10_96_3201_0 & ~i_10_96_3583_0 & ~i_10_96_3992_0 & i_10_96_4119_0 & ~i_10_96_4129_0) | (i_10_96_174_0 & i_10_96_175_0 & ~i_10_96_2468_0 & ~i_10_96_2707_0 & ~i_10_96_2783_0 & ~i_10_96_2924_0 & ~i_10_96_3044_0 & ~i_10_96_3584_0 & ~i_10_96_3852_0 & ~i_10_96_4269_0))) | (~i_10_96_2786_0 & ((~i_10_96_1823_0 & i_10_96_2356_0 & ~i_10_96_2631_0 & ~i_10_96_2785_0 & ~i_10_96_3584_0) | (~i_10_96_221_0 & ~i_10_96_391_0 & ~i_10_96_4130_0 & i_10_96_4288_0))) | (i_10_96_328_0 & i_10_96_3201_0) | (i_10_96_2603_0 & i_10_96_2633_0 & i_10_96_3612_0) | (~i_10_96_2024_0 & i_10_96_3389_0 & ~i_10_96_3613_0 & i_10_96_4288_0) | (~i_10_96_4130_0 & i_10_96_4276_0) | (~i_10_96_1822_0 & ~i_10_96_1997_0 & i_10_96_2923_0 & ~i_10_96_3992_0 & i_10_96_4289_0));
endmodule



// Benchmark "kernel_10_97" written by ABC on Sun Jul 19 10:22:39 2020

module kernel_10_97 ( 
    i_10_97_49_0, i_10_97_123_0, i_10_97_124_0, i_10_97_171_0,
    i_10_97_217_0, i_10_97_218_0, i_10_97_244_0, i_10_97_293_0,
    i_10_97_317_0, i_10_97_320_0, i_10_97_325_0, i_10_97_431_0,
    i_10_97_432_0, i_10_97_462_0, i_10_97_512_0, i_10_97_990_0,
    i_10_97_1084_0, i_10_97_1306_0, i_10_97_1450_0, i_10_97_1576_0,
    i_10_97_1577_0, i_10_97_1619_0, i_10_97_1621_0, i_10_97_1649_0,
    i_10_97_1685_0, i_10_97_1687_0, i_10_97_1767_0, i_10_97_1820_0,
    i_10_97_1823_0, i_10_97_1990_0, i_10_97_1991_0, i_10_97_2003_0,
    i_10_97_2312_0, i_10_97_2351_0, i_10_97_2359_0, i_10_97_2360_0,
    i_10_97_2362_0, i_10_97_2363_0, i_10_97_2377_0, i_10_97_2449_0,
    i_10_97_2462_0, i_10_97_2468_0, i_10_97_2510_0, i_10_97_2628_0,
    i_10_97_2636_0, i_10_97_2639_0, i_10_97_2681_0, i_10_97_2711_0,
    i_10_97_2712_0, i_10_97_2713_0, i_10_97_2723_0, i_10_97_2731_0,
    i_10_97_2828_0, i_10_97_2831_0, i_10_97_2881_0, i_10_97_2882_0,
    i_10_97_2916_0, i_10_97_2917_0, i_10_97_2918_0, i_10_97_2919_0,
    i_10_97_2921_0, i_10_97_2924_0, i_10_97_3069_0, i_10_97_3198_0,
    i_10_97_3200_0, i_10_97_3269_0, i_10_97_3273_0, i_10_97_3289_0,
    i_10_97_3290_0, i_10_97_3402_0, i_10_97_3404_0, i_10_97_3406_0,
    i_10_97_3407_0, i_10_97_3538_0, i_10_97_3610_0, i_10_97_3611_0,
    i_10_97_3648_0, i_10_97_3649_0, i_10_97_3731_0, i_10_97_3734_0,
    i_10_97_3787_0, i_10_97_3788_0, i_10_97_3815_0, i_10_97_3835_0,
    i_10_97_3846_0, i_10_97_3910_0, i_10_97_3981_0, i_10_97_3982_0,
    i_10_97_3983_0, i_10_97_3986_0, i_10_97_3991_0, i_10_97_4027_0,
    i_10_97_4028_0, i_10_97_4030_0, i_10_97_4031_0, i_10_97_4121_0,
    i_10_97_4127_0, i_10_97_4214_0, i_10_97_4274_0, i_10_97_4290_0,
    o_10_97_0_0  );
  input  i_10_97_49_0, i_10_97_123_0, i_10_97_124_0, i_10_97_171_0,
    i_10_97_217_0, i_10_97_218_0, i_10_97_244_0, i_10_97_293_0,
    i_10_97_317_0, i_10_97_320_0, i_10_97_325_0, i_10_97_431_0,
    i_10_97_432_0, i_10_97_462_0, i_10_97_512_0, i_10_97_990_0,
    i_10_97_1084_0, i_10_97_1306_0, i_10_97_1450_0, i_10_97_1576_0,
    i_10_97_1577_0, i_10_97_1619_0, i_10_97_1621_0, i_10_97_1649_0,
    i_10_97_1685_0, i_10_97_1687_0, i_10_97_1767_0, i_10_97_1820_0,
    i_10_97_1823_0, i_10_97_1990_0, i_10_97_1991_0, i_10_97_2003_0,
    i_10_97_2312_0, i_10_97_2351_0, i_10_97_2359_0, i_10_97_2360_0,
    i_10_97_2362_0, i_10_97_2363_0, i_10_97_2377_0, i_10_97_2449_0,
    i_10_97_2462_0, i_10_97_2468_0, i_10_97_2510_0, i_10_97_2628_0,
    i_10_97_2636_0, i_10_97_2639_0, i_10_97_2681_0, i_10_97_2711_0,
    i_10_97_2712_0, i_10_97_2713_0, i_10_97_2723_0, i_10_97_2731_0,
    i_10_97_2828_0, i_10_97_2831_0, i_10_97_2881_0, i_10_97_2882_0,
    i_10_97_2916_0, i_10_97_2917_0, i_10_97_2918_0, i_10_97_2919_0,
    i_10_97_2921_0, i_10_97_2924_0, i_10_97_3069_0, i_10_97_3198_0,
    i_10_97_3200_0, i_10_97_3269_0, i_10_97_3273_0, i_10_97_3289_0,
    i_10_97_3290_0, i_10_97_3402_0, i_10_97_3404_0, i_10_97_3406_0,
    i_10_97_3407_0, i_10_97_3538_0, i_10_97_3610_0, i_10_97_3611_0,
    i_10_97_3648_0, i_10_97_3649_0, i_10_97_3731_0, i_10_97_3734_0,
    i_10_97_3787_0, i_10_97_3788_0, i_10_97_3815_0, i_10_97_3835_0,
    i_10_97_3846_0, i_10_97_3910_0, i_10_97_3981_0, i_10_97_3982_0,
    i_10_97_3983_0, i_10_97_3986_0, i_10_97_3991_0, i_10_97_4027_0,
    i_10_97_4028_0, i_10_97_4030_0, i_10_97_4031_0, i_10_97_4121_0,
    i_10_97_4127_0, i_10_97_4214_0, i_10_97_4274_0, i_10_97_4290_0;
  output o_10_97_0_0;
  assign o_10_97_0_0 = 0;
endmodule



// Benchmark "kernel_10_98" written by ABC on Sun Jul 19 10:22:40 2020

module kernel_10_98 ( 
    i_10_98_48_0, i_10_98_173_0, i_10_98_181_0, i_10_98_223_0,
    i_10_98_287_0, i_10_98_319_0, i_10_98_320_0, i_10_98_347_0,
    i_10_98_393_0, i_10_98_442_0, i_10_98_445_0, i_10_98_448_0,
    i_10_98_463_0, i_10_98_716_0, i_10_98_719_0, i_10_98_793_0,
    i_10_98_799_0, i_10_98_827_0, i_10_98_832_0, i_10_98_963_0,
    i_10_98_964_0, i_10_98_967_0, i_10_98_1081_0, i_10_98_1085_0,
    i_10_98_1238_0, i_10_98_1248_0, i_10_98_1249_0, i_10_98_1309_0,
    i_10_98_1313_0, i_10_98_1364_0, i_10_98_1367_0, i_10_98_1438_0,
    i_10_98_1575_0, i_10_98_1579_0, i_10_98_1616_0, i_10_98_1641_0,
    i_10_98_1642_0, i_10_98_1648_0, i_10_98_1685_0, i_10_98_1687_0,
    i_10_98_1689_0, i_10_98_1821_0, i_10_98_1908_0, i_10_98_1916_0,
    i_10_98_1948_0, i_10_98_2020_0, i_10_98_2455_0, i_10_98_2470_0,
    i_10_98_2508_0, i_10_98_2520_0, i_10_98_2604_0, i_10_98_2634_0,
    i_10_98_2704_0, i_10_98_2714_0, i_10_98_2726_0, i_10_98_2729_0,
    i_10_98_2828_0, i_10_98_2884_0, i_10_98_2885_0, i_10_98_2888_0,
    i_10_98_2916_0, i_10_98_2923_0, i_10_98_2924_0, i_10_98_2958_0,
    i_10_98_3037_0, i_10_98_3196_0, i_10_98_3270_0, i_10_98_3284_0,
    i_10_98_3384_0, i_10_98_3388_0, i_10_98_3429_0, i_10_98_3446_0,
    i_10_98_3505_0, i_10_98_3522_0, i_10_98_3523_0, i_10_98_3559_0,
    i_10_98_3561_0, i_10_98_3563_0, i_10_98_3589_0, i_10_98_3614_0,
    i_10_98_3650_0, i_10_98_3651_0, i_10_98_3652_0, i_10_98_3810_0,
    i_10_98_3811_0, i_10_98_3859_0, i_10_98_3860_0, i_10_98_3948_0,
    i_10_98_3949_0, i_10_98_3978_0, i_10_98_3981_0, i_10_98_4050_0,
    i_10_98_4114_0, i_10_98_4117_0, i_10_98_4204_0, i_10_98_4217_0,
    i_10_98_4284_0, i_10_98_4288_0, i_10_98_4291_0, i_10_98_4292_0,
    o_10_98_0_0  );
  input  i_10_98_48_0, i_10_98_173_0, i_10_98_181_0, i_10_98_223_0,
    i_10_98_287_0, i_10_98_319_0, i_10_98_320_0, i_10_98_347_0,
    i_10_98_393_0, i_10_98_442_0, i_10_98_445_0, i_10_98_448_0,
    i_10_98_463_0, i_10_98_716_0, i_10_98_719_0, i_10_98_793_0,
    i_10_98_799_0, i_10_98_827_0, i_10_98_832_0, i_10_98_963_0,
    i_10_98_964_0, i_10_98_967_0, i_10_98_1081_0, i_10_98_1085_0,
    i_10_98_1238_0, i_10_98_1248_0, i_10_98_1249_0, i_10_98_1309_0,
    i_10_98_1313_0, i_10_98_1364_0, i_10_98_1367_0, i_10_98_1438_0,
    i_10_98_1575_0, i_10_98_1579_0, i_10_98_1616_0, i_10_98_1641_0,
    i_10_98_1642_0, i_10_98_1648_0, i_10_98_1685_0, i_10_98_1687_0,
    i_10_98_1689_0, i_10_98_1821_0, i_10_98_1908_0, i_10_98_1916_0,
    i_10_98_1948_0, i_10_98_2020_0, i_10_98_2455_0, i_10_98_2470_0,
    i_10_98_2508_0, i_10_98_2520_0, i_10_98_2604_0, i_10_98_2634_0,
    i_10_98_2704_0, i_10_98_2714_0, i_10_98_2726_0, i_10_98_2729_0,
    i_10_98_2828_0, i_10_98_2884_0, i_10_98_2885_0, i_10_98_2888_0,
    i_10_98_2916_0, i_10_98_2923_0, i_10_98_2924_0, i_10_98_2958_0,
    i_10_98_3037_0, i_10_98_3196_0, i_10_98_3270_0, i_10_98_3284_0,
    i_10_98_3384_0, i_10_98_3388_0, i_10_98_3429_0, i_10_98_3446_0,
    i_10_98_3505_0, i_10_98_3522_0, i_10_98_3523_0, i_10_98_3559_0,
    i_10_98_3561_0, i_10_98_3563_0, i_10_98_3589_0, i_10_98_3614_0,
    i_10_98_3650_0, i_10_98_3651_0, i_10_98_3652_0, i_10_98_3810_0,
    i_10_98_3811_0, i_10_98_3859_0, i_10_98_3860_0, i_10_98_3948_0,
    i_10_98_3949_0, i_10_98_3978_0, i_10_98_3981_0, i_10_98_4050_0,
    i_10_98_4114_0, i_10_98_4117_0, i_10_98_4204_0, i_10_98_4217_0,
    i_10_98_4284_0, i_10_98_4288_0, i_10_98_4291_0, i_10_98_4292_0;
  output o_10_98_0_0;
  assign o_10_98_0_0 = 0;
endmodule



// Benchmark "kernel_10_99" written by ABC on Sun Jul 19 10:22:41 2020

module kernel_10_99 ( 
    i_10_99_39_0, i_10_99_121_0, i_10_99_148_0, i_10_99_149_0,
    i_10_99_157_0, i_10_99_188_0, i_10_99_244_0, i_10_99_256_0,
    i_10_99_257_0, i_10_99_271_0, i_10_99_394_0, i_10_99_395_0,
    i_10_99_445_0, i_10_99_544_0, i_10_99_585_0, i_10_99_598_0,
    i_10_99_601_0, i_10_99_602_0, i_10_99_688_0, i_10_99_734_0,
    i_10_99_800_0, i_10_99_880_0, i_10_99_1003_0, i_10_99_1013_0,
    i_10_99_1154_0, i_10_99_1241_0, i_10_99_1242_0, i_10_99_1249_0,
    i_10_99_1281_0, i_10_99_1438_0, i_10_99_1441_0, i_10_99_1516_0,
    i_10_99_1542_0, i_10_99_1544_0, i_10_99_1560_0, i_10_99_1565_0,
    i_10_99_1580_0, i_10_99_1612_0, i_10_99_1615_0, i_10_99_1616_0,
    i_10_99_1686_0, i_10_99_1819_0, i_10_99_1822_0, i_10_99_1823_0,
    i_10_99_1885_0, i_10_99_1920_0, i_10_99_1959_0, i_10_99_1961_0,
    i_10_99_2020_0, i_10_99_2023_0, i_10_99_2349_0, i_10_99_2350_0,
    i_10_99_2353_0, i_10_99_2354_0, i_10_99_2408_0, i_10_99_2518_0,
    i_10_99_2532_0, i_10_99_2535_0, i_10_99_2536_0, i_10_99_2537_0,
    i_10_99_2629_0, i_10_99_2632_0, i_10_99_2634_0, i_10_99_2696_0,
    i_10_99_2713_0, i_10_99_2734_0, i_10_99_2735_0, i_10_99_2821_0,
    i_10_99_2833_0, i_10_99_2870_0, i_10_99_2884_0, i_10_99_2984_0,
    i_10_99_3199_0, i_10_99_3269_0, i_10_99_3392_0, i_10_99_3431_0,
    i_10_99_3433_0, i_10_99_3496_0, i_10_99_3524_0, i_10_99_3582_0,
    i_10_99_3609_0, i_10_99_3784_0, i_10_99_3881_0, i_10_99_3944_0,
    i_10_99_3982_0, i_10_99_4013_0, i_10_99_4113_0, i_10_99_4114_0,
    i_10_99_4117_0, i_10_99_4175_0, i_10_99_4178_0, i_10_99_4186_0,
    i_10_99_4214_0, i_10_99_4267_0, i_10_99_4270_0, i_10_99_4273_0,
    i_10_99_4522_0, i_10_99_4564_0, i_10_99_4565_0, i_10_99_4566_0,
    o_10_99_0_0  );
  input  i_10_99_39_0, i_10_99_121_0, i_10_99_148_0, i_10_99_149_0,
    i_10_99_157_0, i_10_99_188_0, i_10_99_244_0, i_10_99_256_0,
    i_10_99_257_0, i_10_99_271_0, i_10_99_394_0, i_10_99_395_0,
    i_10_99_445_0, i_10_99_544_0, i_10_99_585_0, i_10_99_598_0,
    i_10_99_601_0, i_10_99_602_0, i_10_99_688_0, i_10_99_734_0,
    i_10_99_800_0, i_10_99_880_0, i_10_99_1003_0, i_10_99_1013_0,
    i_10_99_1154_0, i_10_99_1241_0, i_10_99_1242_0, i_10_99_1249_0,
    i_10_99_1281_0, i_10_99_1438_0, i_10_99_1441_0, i_10_99_1516_0,
    i_10_99_1542_0, i_10_99_1544_0, i_10_99_1560_0, i_10_99_1565_0,
    i_10_99_1580_0, i_10_99_1612_0, i_10_99_1615_0, i_10_99_1616_0,
    i_10_99_1686_0, i_10_99_1819_0, i_10_99_1822_0, i_10_99_1823_0,
    i_10_99_1885_0, i_10_99_1920_0, i_10_99_1959_0, i_10_99_1961_0,
    i_10_99_2020_0, i_10_99_2023_0, i_10_99_2349_0, i_10_99_2350_0,
    i_10_99_2353_0, i_10_99_2354_0, i_10_99_2408_0, i_10_99_2518_0,
    i_10_99_2532_0, i_10_99_2535_0, i_10_99_2536_0, i_10_99_2537_0,
    i_10_99_2629_0, i_10_99_2632_0, i_10_99_2634_0, i_10_99_2696_0,
    i_10_99_2713_0, i_10_99_2734_0, i_10_99_2735_0, i_10_99_2821_0,
    i_10_99_2833_0, i_10_99_2870_0, i_10_99_2884_0, i_10_99_2984_0,
    i_10_99_3199_0, i_10_99_3269_0, i_10_99_3392_0, i_10_99_3431_0,
    i_10_99_3433_0, i_10_99_3496_0, i_10_99_3524_0, i_10_99_3582_0,
    i_10_99_3609_0, i_10_99_3784_0, i_10_99_3881_0, i_10_99_3944_0,
    i_10_99_3982_0, i_10_99_4013_0, i_10_99_4113_0, i_10_99_4114_0,
    i_10_99_4117_0, i_10_99_4175_0, i_10_99_4178_0, i_10_99_4186_0,
    i_10_99_4214_0, i_10_99_4267_0, i_10_99_4270_0, i_10_99_4273_0,
    i_10_99_4522_0, i_10_99_4564_0, i_10_99_4565_0, i_10_99_4566_0;
  output o_10_99_0_0;
  assign o_10_99_0_0 = ~((~i_10_99_1438_0 & ((~i_10_99_244_0 & ~i_10_99_1612_0 & ((~i_10_99_1580_0 & ~i_10_99_1615_0 & ~i_10_99_1819_0 & ~i_10_99_2353_0 & ~i_10_99_2833_0 & ~i_10_99_3431_0) | (~i_10_99_2354_0 & ~i_10_99_3199_0 & ~i_10_99_3269_0 & ~i_10_99_3392_0 & i_10_99_4565_0))) | (~i_10_99_4270_0 & ((~i_10_99_256_0 & ((~i_10_99_2629_0 & ~i_10_99_2833_0 & ~i_10_99_3431_0 & ~i_10_99_3582_0 & i_10_99_4114_0 & ~i_10_99_4267_0) | (~i_10_99_148_0 & ~i_10_99_257_0 & ~i_10_99_395_0 & i_10_99_1819_0 & ~i_10_99_2023_0 & ~i_10_99_4273_0))) | (i_10_99_1823_0 & ~i_10_99_2629_0 & ~i_10_99_3433_0 & ~i_10_99_4214_0 & ~i_10_99_4565_0 & ~i_10_99_4566_0))) | (~i_10_99_257_0 & ~i_10_99_1003_0 & ~i_10_99_1686_0 & ~i_10_99_2632_0 & ~i_10_99_3199_0 & ~i_10_99_3269_0 & ~i_10_99_3433_0 & ~i_10_99_3582_0 & ~i_10_99_4267_0) | (~i_10_99_121_0 & ~i_10_99_1542_0 & ~i_10_99_1544_0 & ~i_10_99_2353_0 & ~i_10_99_3982_0 & ~i_10_99_4117_0) | (~i_10_99_2629_0 & i_10_99_2632_0 & ~i_10_99_2735_0 & ~i_10_99_2833_0 & ~i_10_99_2984_0 & ~i_10_99_4114_0 & ~i_10_99_4565_0))) | (~i_10_99_2629_0 & ((~i_10_99_148_0 & ((~i_10_99_395_0 & ~i_10_99_1242_0 & ~i_10_99_1249_0 & i_10_99_1686_0 & ~i_10_99_2354_0 & ~i_10_99_4175_0) | (~i_10_99_257_0 & ~i_10_99_394_0 & ~i_10_99_1544_0 & i_10_99_2354_0 & ~i_10_99_2634_0 & ~i_10_99_2735_0 & ~i_10_99_3609_0 & ~i_10_99_4113_0 & ~i_10_99_4267_0 & ~i_10_99_4564_0))) | (~i_10_99_121_0 & ~i_10_99_244_0 & ~i_10_99_1542_0 & ~i_10_99_1580_0 & ~i_10_99_2408_0 & ~i_10_99_3784_0 & ~i_10_99_3982_0 & ~i_10_99_4175_0))) | (~i_10_99_121_0 & ((~i_10_99_1544_0 & ~i_10_99_2353_0 & ~i_10_99_2833_0 & ~i_10_99_3199_0 & i_10_99_4113_0) | (~i_10_99_244_0 & ~i_10_99_1542_0 & ~i_10_99_1580_0 & ~i_10_99_3269_0 & ~i_10_99_3392_0 & ~i_10_99_3431_0 & ~i_10_99_4175_0 & ~i_10_99_4564_0))) | (~i_10_99_2349_0 & ((~i_10_99_3433_0 & ((~i_10_99_244_0 & ((~i_10_99_257_0 & i_10_99_2735_0 & ~i_10_99_3392_0 & ~i_10_99_4270_0) | (~i_10_99_800_0 & ~i_10_99_2353_0 & ~i_10_99_4267_0 & ~i_10_99_4273_0))) | (~i_10_99_1542_0 & ~i_10_99_1544_0 & ~i_10_99_1612_0 & ~i_10_99_1819_0 & ~i_10_99_2833_0 & ~i_10_99_3496_0 & ~i_10_99_3609_0 & ~i_10_99_3982_0 & ~i_10_99_4565_0 & ~i_10_99_4566_0))) | (~i_10_99_1542_0 & ~i_10_99_1615_0 & ~i_10_99_2354_0 & ~i_10_99_3199_0 & ~i_10_99_3431_0) | (~i_10_99_1242_0 & ~i_10_99_1580_0 & ~i_10_99_3609_0 & ~i_10_99_4270_0 & ~i_10_99_4566_0))) | (~i_10_99_1544_0 & ((~i_10_99_1242_0 & ((~i_10_99_2020_0 & ~i_10_99_2350_0 & ~i_10_99_2354_0 & ~i_10_99_4117_0) | (i_10_99_1686_0 & i_10_99_1819_0 & ~i_10_99_1822_0 & ~i_10_99_3582_0 & ~i_10_99_4565_0))) | (~i_10_99_1003_0 & ~i_10_99_1249_0 & ~i_10_99_1542_0 & ~i_10_99_2353_0 & ~i_10_99_2408_0 & ~i_10_99_3496_0 & ~i_10_99_4113_0))) | (~i_10_99_4566_0 & ((~i_10_99_257_0 & ~i_10_99_4175_0 & ((~i_10_99_1542_0 & ~i_10_99_1615_0 & ~i_10_99_2353_0 & ~i_10_99_4267_0 & ~i_10_99_4270_0) | (~i_10_99_2350_0 & ~i_10_99_2408_0 & i_10_99_2634_0 & ~i_10_99_4565_0))) | (~i_10_99_1615_0 & ~i_10_99_2350_0 & ~i_10_99_2884_0 & i_10_99_3524_0))) | (~i_10_99_3609_0 & ((~i_10_99_1542_0 & ((~i_10_99_1686_0 & ((~i_10_99_395_0 & ~i_10_99_2020_0 & ~i_10_99_2408_0 & ~i_10_99_2884_0 & ~i_10_99_2984_0 & ~i_10_99_3784_0 & ~i_10_99_4267_0) | (~i_10_99_257_0 & ~i_10_99_1249_0 & ~i_10_99_2350_0 & ~i_10_99_3524_0 & ~i_10_99_4175_0 & ~i_10_99_4565_0))) | (i_10_99_1819_0 & ~i_10_99_2354_0 & ~i_10_99_3392_0 & ~i_10_99_3524_0 & ~i_10_99_4113_0))) | (i_10_99_2821_0 & i_10_99_3524_0 & ~i_10_99_3982_0))) | (~i_10_99_257_0 & ((i_10_99_1249_0 & ~i_10_99_1823_0 & ~i_10_99_2350_0 & ~i_10_99_3392_0 & ~i_10_99_3433_0) | (i_10_99_148_0 & ~i_10_99_1580_0 & i_10_99_4114_0))) | (~i_10_99_2354_0 & ((i_10_99_1822_0 & ((~i_10_99_1249_0 & ~i_10_99_1580_0 & ~i_10_99_2350_0) | (~i_10_99_1823_0 & i_10_99_3433_0))) | (~i_10_99_1819_0 & i_10_99_2353_0 & ~i_10_99_2884_0 & ~i_10_99_3431_0 & ~i_10_99_3784_0 & ~i_10_99_4273_0 & ~i_10_99_4565_0))) | (~i_10_99_1249_0 & ~i_10_99_1580_0 & (i_10_99_2821_0 | (~i_10_99_2023_0 & ~i_10_99_2884_0 & i_10_99_3582_0 & ~i_10_99_4565_0))) | (~i_10_99_2984_0 & ~i_10_99_3433_0 & i_10_99_3496_0) | (i_10_99_2634_0 & i_10_99_2734_0 & i_10_99_3524_0) | (i_10_99_2023_0 & i_10_99_2408_0 & i_10_99_4566_0));
endmodule



// Benchmark "kernel_10_100" written by ABC on Sun Jul 19 10:22:43 2020

module kernel_10_100 ( 
    i_10_100_27_0, i_10_100_251_0, i_10_100_406_0, i_10_100_408_0,
    i_10_100_432_0, i_10_100_441_0, i_10_100_444_0, i_10_100_445_0,
    i_10_100_730_0, i_10_100_755_0, i_10_100_954_0, i_10_100_1000_0,
    i_10_100_1001_0, i_10_100_1005_0, i_10_100_1083_0, i_10_100_1234_0,
    i_10_100_1235_0, i_10_100_1241_0, i_10_100_1274_0, i_10_100_1307_0,
    i_10_100_1310_0, i_10_100_1313_0, i_10_100_1546_0, i_10_100_1547_0,
    i_10_100_1549_0, i_10_100_1550_0, i_10_100_1552_0, i_10_100_1612_0,
    i_10_100_1613_0, i_10_100_1649_0, i_10_100_1655_0, i_10_100_1677_0,
    i_10_100_1684_0, i_10_100_1690_0, i_10_100_1720_0, i_10_100_1823_0,
    i_10_100_1944_0, i_10_100_1945_0, i_10_100_1946_0, i_10_100_2083_0,
    i_10_100_2152_0, i_10_100_2179_0, i_10_100_2180_0, i_10_100_2200_0,
    i_10_100_2201_0, i_10_100_2306_0, i_10_100_2380_0, i_10_100_2405_0,
    i_10_100_2407_0, i_10_100_2449_0, i_10_100_2453_0, i_10_100_2459_0,
    i_10_100_2472_0, i_10_100_2474_0, i_10_100_2632_0, i_10_100_2654_0,
    i_10_100_2722_0, i_10_100_2723_0, i_10_100_2731_0, i_10_100_2741_0,
    i_10_100_2826_0, i_10_100_2827_0, i_10_100_2830_0, i_10_100_2831_0,
    i_10_100_2885_0, i_10_100_2917_0, i_10_100_2952_0, i_10_100_2953_0,
    i_10_100_3051_0, i_10_100_3054_0, i_10_100_3055_0, i_10_100_3167_0,
    i_10_100_3277_0, i_10_100_3281_0, i_10_100_3298_0, i_10_100_3387_0,
    i_10_100_3391_0, i_10_100_3392_0, i_10_100_3467_0, i_10_100_3470_0,
    i_10_100_3472_0, i_10_100_3584_0, i_10_100_3587_0, i_10_100_3611_0,
    i_10_100_3612_0, i_10_100_3650_0, i_10_100_3838_0, i_10_100_3854_0,
    i_10_100_3855_0, i_10_100_3859_0, i_10_100_3990_0, i_10_100_3991_0,
    i_10_100_3992_0, i_10_100_4052_0, i_10_100_4054_0, i_10_100_4113_0,
    i_10_100_4117_0, i_10_100_4214_0, i_10_100_4230_0, i_10_100_4266_0,
    o_10_100_0_0  );
  input  i_10_100_27_0, i_10_100_251_0, i_10_100_406_0, i_10_100_408_0,
    i_10_100_432_0, i_10_100_441_0, i_10_100_444_0, i_10_100_445_0,
    i_10_100_730_0, i_10_100_755_0, i_10_100_954_0, i_10_100_1000_0,
    i_10_100_1001_0, i_10_100_1005_0, i_10_100_1083_0, i_10_100_1234_0,
    i_10_100_1235_0, i_10_100_1241_0, i_10_100_1274_0, i_10_100_1307_0,
    i_10_100_1310_0, i_10_100_1313_0, i_10_100_1546_0, i_10_100_1547_0,
    i_10_100_1549_0, i_10_100_1550_0, i_10_100_1552_0, i_10_100_1612_0,
    i_10_100_1613_0, i_10_100_1649_0, i_10_100_1655_0, i_10_100_1677_0,
    i_10_100_1684_0, i_10_100_1690_0, i_10_100_1720_0, i_10_100_1823_0,
    i_10_100_1944_0, i_10_100_1945_0, i_10_100_1946_0, i_10_100_2083_0,
    i_10_100_2152_0, i_10_100_2179_0, i_10_100_2180_0, i_10_100_2200_0,
    i_10_100_2201_0, i_10_100_2306_0, i_10_100_2380_0, i_10_100_2405_0,
    i_10_100_2407_0, i_10_100_2449_0, i_10_100_2453_0, i_10_100_2459_0,
    i_10_100_2472_0, i_10_100_2474_0, i_10_100_2632_0, i_10_100_2654_0,
    i_10_100_2722_0, i_10_100_2723_0, i_10_100_2731_0, i_10_100_2741_0,
    i_10_100_2826_0, i_10_100_2827_0, i_10_100_2830_0, i_10_100_2831_0,
    i_10_100_2885_0, i_10_100_2917_0, i_10_100_2952_0, i_10_100_2953_0,
    i_10_100_3051_0, i_10_100_3054_0, i_10_100_3055_0, i_10_100_3167_0,
    i_10_100_3277_0, i_10_100_3281_0, i_10_100_3298_0, i_10_100_3387_0,
    i_10_100_3391_0, i_10_100_3392_0, i_10_100_3467_0, i_10_100_3470_0,
    i_10_100_3472_0, i_10_100_3584_0, i_10_100_3587_0, i_10_100_3611_0,
    i_10_100_3612_0, i_10_100_3650_0, i_10_100_3838_0, i_10_100_3854_0,
    i_10_100_3855_0, i_10_100_3859_0, i_10_100_3990_0, i_10_100_3991_0,
    i_10_100_3992_0, i_10_100_4052_0, i_10_100_4054_0, i_10_100_4113_0,
    i_10_100_4117_0, i_10_100_4214_0, i_10_100_4230_0, i_10_100_4266_0;
  output o_10_100_0_0;
  assign o_10_100_0_0 = ~((~i_10_100_27_0 & ((~i_10_100_1234_0 & ~i_10_100_1946_0 & ~i_10_100_2405_0 & ~i_10_100_3167_0 & ~i_10_100_3611_0) | (~i_10_100_1001_0 & ~i_10_100_1612_0 & ~i_10_100_1945_0 & ~i_10_100_2453_0 & i_10_100_3854_0))) | (~i_10_100_406_0 & ((~i_10_100_1307_0 & ~i_10_100_1823_0 & ~i_10_100_1945_0) | (~i_10_100_1005_0 & ~i_10_100_1234_0 & ~i_10_100_1552_0 & ~i_10_100_1613_0 & ~i_10_100_1690_0 & ~i_10_100_3167_0 & ~i_10_100_4230_0))) | (~i_10_100_444_0 & ((~i_10_100_445_0 & ~i_10_100_755_0 & ~i_10_100_1945_0 & ~i_10_100_3472_0) | (~i_10_100_1613_0 & ~i_10_100_2180_0 & ~i_10_100_2453_0 & ~i_10_100_2827_0 & ~i_10_100_3277_0 & ~i_10_100_3612_0))) | (~i_10_100_2200_0 & ~i_10_100_4230_0 & ((~i_10_100_445_0 & ~i_10_100_2405_0) | (~i_10_100_1005_0 & ~i_10_100_2306_0 & ~i_10_100_2472_0 & ~i_10_100_3467_0 & ~i_10_100_3990_0 & ~i_10_100_4052_0))) | (~i_10_100_2201_0 & (i_10_100_2831_0 | (~i_10_100_441_0 & ~i_10_100_1005_0 & ~i_10_100_1313_0 & ~i_10_100_1613_0 & ~i_10_100_3467_0 & ~i_10_100_3611_0 & ~i_10_100_4054_0))) | (~i_10_100_2306_0 & ~i_10_100_3472_0 & ((~i_10_100_1000_0 & ~i_10_100_2453_0 & ~i_10_100_3584_0) | (~i_10_100_1083_0 & ~i_10_100_2180_0 & ~i_10_100_3838_0))) | (~i_10_100_1005_0 & ~i_10_100_1944_0 & ((~i_10_100_3990_0 & ((~i_10_100_1001_0 & ~i_10_100_3838_0) | (~i_10_100_954_0 & i_10_100_2449_0 & ~i_10_100_4266_0))) | (i_10_100_1549_0 & ~i_10_100_1823_0 & ~i_10_100_3584_0))) | (i_10_100_1649_0 & i_10_100_2917_0) | (~i_10_100_1612_0 & ~i_10_100_1655_0 & i_10_100_1945_0 & ~i_10_100_3587_0 & ~i_10_100_4266_0) | (~i_10_100_1310_0 & ~i_10_100_1547_0 & ~i_10_100_1649_0 & ~i_10_100_2179_0 & ~i_10_100_3612_0 & ~i_10_100_3855_0 & ~i_10_100_4113_0));
endmodule



// Benchmark "kernel_10_101" written by ABC on Sun Jul 19 10:22:44 2020

module kernel_10_101 ( 
    i_10_101_36_0, i_10_101_37_0, i_10_101_155_0, i_10_101_172_0,
    i_10_101_175_0, i_10_101_176_0, i_10_101_221_0, i_10_101_281_0,
    i_10_101_282_0, i_10_101_296_0, i_10_101_315_0, i_10_101_316_0,
    i_10_101_390_0, i_10_101_434_0, i_10_101_438_0, i_10_101_442_0,
    i_10_101_793_0, i_10_101_796_0, i_10_101_797_0, i_10_101_800_0,
    i_10_101_899_0, i_10_101_990_0, i_10_101_996_0, i_10_101_1085_0,
    i_10_101_1153_0, i_10_101_1237_0, i_10_101_1238_0, i_10_101_1239_0,
    i_10_101_1306_0, i_10_101_1341_0, i_10_101_1345_0, i_10_101_1349_0,
    i_10_101_1441_0, i_10_101_1551_0, i_10_101_1654_0, i_10_101_1655_0,
    i_10_101_1676_0, i_10_101_1686_0, i_10_101_1825_0, i_10_101_1910_0,
    i_10_101_1944_0, i_10_101_2005_0, i_10_101_2019_0, i_10_101_2352_0,
    i_10_101_2356_0, i_10_101_2365_0, i_10_101_2514_0, i_10_101_2628_0,
    i_10_101_2629_0, i_10_101_2630_0, i_10_101_2631_0, i_10_101_2632_0,
    i_10_101_2633_0, i_10_101_2636_0, i_10_101_2657_0, i_10_101_2661_0,
    i_10_101_2673_0, i_10_101_2703_0, i_10_101_2704_0, i_10_101_2705_0,
    i_10_101_2711_0, i_10_101_2729_0, i_10_101_2783_0, i_10_101_2829_0,
    i_10_101_2831_0, i_10_101_2885_0, i_10_101_2916_0, i_10_101_2923_0,
    i_10_101_2984_0, i_10_101_3034_0, i_10_101_3035_0, i_10_101_3069_0,
    i_10_101_3070_0, i_10_101_3198_0, i_10_101_3234_0, i_10_101_3270_0,
    i_10_101_3280_0, i_10_101_3384_0, i_10_101_3522_0, i_10_101_3540_0,
    i_10_101_3583_0, i_10_101_3609_0, i_10_101_3612_0, i_10_101_3613_0,
    i_10_101_3647_0, i_10_101_3837_0, i_10_101_3839_0, i_10_101_3853_0,
    i_10_101_3855_0, i_10_101_3856_0, i_10_101_3860_0, i_10_101_3872_0,
    i_10_101_4122_0, i_10_101_4123_0, i_10_101_4125_0, i_10_101_4126_0,
    i_10_101_4167_0, i_10_101_4168_0, i_10_101_4287_0, i_10_101_4566_0,
    o_10_101_0_0  );
  input  i_10_101_36_0, i_10_101_37_0, i_10_101_155_0, i_10_101_172_0,
    i_10_101_175_0, i_10_101_176_0, i_10_101_221_0, i_10_101_281_0,
    i_10_101_282_0, i_10_101_296_0, i_10_101_315_0, i_10_101_316_0,
    i_10_101_390_0, i_10_101_434_0, i_10_101_438_0, i_10_101_442_0,
    i_10_101_793_0, i_10_101_796_0, i_10_101_797_0, i_10_101_800_0,
    i_10_101_899_0, i_10_101_990_0, i_10_101_996_0, i_10_101_1085_0,
    i_10_101_1153_0, i_10_101_1237_0, i_10_101_1238_0, i_10_101_1239_0,
    i_10_101_1306_0, i_10_101_1341_0, i_10_101_1345_0, i_10_101_1349_0,
    i_10_101_1441_0, i_10_101_1551_0, i_10_101_1654_0, i_10_101_1655_0,
    i_10_101_1676_0, i_10_101_1686_0, i_10_101_1825_0, i_10_101_1910_0,
    i_10_101_1944_0, i_10_101_2005_0, i_10_101_2019_0, i_10_101_2352_0,
    i_10_101_2356_0, i_10_101_2365_0, i_10_101_2514_0, i_10_101_2628_0,
    i_10_101_2629_0, i_10_101_2630_0, i_10_101_2631_0, i_10_101_2632_0,
    i_10_101_2633_0, i_10_101_2636_0, i_10_101_2657_0, i_10_101_2661_0,
    i_10_101_2673_0, i_10_101_2703_0, i_10_101_2704_0, i_10_101_2705_0,
    i_10_101_2711_0, i_10_101_2729_0, i_10_101_2783_0, i_10_101_2829_0,
    i_10_101_2831_0, i_10_101_2885_0, i_10_101_2916_0, i_10_101_2923_0,
    i_10_101_2984_0, i_10_101_3034_0, i_10_101_3035_0, i_10_101_3069_0,
    i_10_101_3070_0, i_10_101_3198_0, i_10_101_3234_0, i_10_101_3270_0,
    i_10_101_3280_0, i_10_101_3384_0, i_10_101_3522_0, i_10_101_3540_0,
    i_10_101_3583_0, i_10_101_3609_0, i_10_101_3612_0, i_10_101_3613_0,
    i_10_101_3647_0, i_10_101_3837_0, i_10_101_3839_0, i_10_101_3853_0,
    i_10_101_3855_0, i_10_101_3856_0, i_10_101_3860_0, i_10_101_3872_0,
    i_10_101_4122_0, i_10_101_4123_0, i_10_101_4125_0, i_10_101_4126_0,
    i_10_101_4167_0, i_10_101_4168_0, i_10_101_4287_0, i_10_101_4566_0;
  output o_10_101_0_0;
  assign o_10_101_0_0 = ~((~i_10_101_4126_0 & ((~i_10_101_175_0 & ((~i_10_101_390_0 & ~i_10_101_1237_0 & ~i_10_101_1441_0 & ~i_10_101_2356_0 & ~i_10_101_2673_0 & ~i_10_101_2704_0 & ~i_10_101_3035_0 & ~i_10_101_3540_0) | (~i_10_101_442_0 & ~i_10_101_793_0 & ~i_10_101_2636_0 & i_10_101_3613_0 & ~i_10_101_3853_0 & ~i_10_101_3855_0 & ~i_10_101_4168_0))) | (~i_10_101_282_0 & ~i_10_101_2661_0 & ~i_10_101_2829_0 & ~i_10_101_2831_0 & ~i_10_101_2916_0 & ~i_10_101_3069_0 & ~i_10_101_4122_0) | (~i_10_101_1237_0 & i_10_101_1306_0 & ~i_10_101_1441_0 & ~i_10_101_3612_0 & ~i_10_101_3839_0 & ~i_10_101_4125_0) | (~i_10_101_172_0 & ~i_10_101_1345_0 & ~i_10_101_1349_0 & i_10_101_2703_0 & ~i_10_101_3070_0 & ~i_10_101_3613_0 & ~i_10_101_4123_0 & ~i_10_101_4287_0))) | (~i_10_101_2019_0 & ((~i_10_101_315_0 & ((~i_10_101_996_0 & ~i_10_101_1349_0 & ~i_10_101_2705_0 & ~i_10_101_3070_0 & ~i_10_101_4122_0) | (~i_10_101_296_0 & ~i_10_101_438_0 & ~i_10_101_4123_0 & ~i_10_101_4125_0))) | (~i_10_101_3069_0 & ~i_10_101_3855_0 & ((~i_10_101_797_0 & ~i_10_101_1341_0 & ~i_10_101_2704_0 & ~i_10_101_2729_0 & ~i_10_101_2831_0 & ~i_10_101_2885_0 & ~i_10_101_2916_0 & ~i_10_101_4122_0) | (~i_10_101_2631_0 & ~i_10_101_2829_0 & ~i_10_101_3839_0 & ~i_10_101_3856_0 & ~i_10_101_4125_0 & ~i_10_101_4167_0))) | (~i_10_101_172_0 & (i_10_101_2630_0 | (~i_10_101_2831_0 & ((~i_10_101_282_0 & ~i_10_101_1825_0 & i_10_101_2628_0) | (~i_10_101_996_0 & i_10_101_2632_0))))) | (i_10_101_2633_0 & ~i_10_101_3540_0 & i_10_101_3856_0))) | (~i_10_101_1306_0 & ((~i_10_101_990_0 & ~i_10_101_1551_0 & ~i_10_101_2783_0 & ~i_10_101_2831_0 & ~i_10_101_3070_0 & ~i_10_101_3612_0 & ~i_10_101_3860_0 & ~i_10_101_4122_0) | (~i_10_101_1345_0 & ~i_10_101_1441_0 & ~i_10_101_2661_0 & ~i_10_101_2711_0 & ~i_10_101_3034_0 & ~i_10_101_3198_0 & ~i_10_101_3384_0 & ~i_10_101_4125_0 & ~i_10_101_4287_0))) | (~i_10_101_390_0 & ((~i_10_101_1345_0 & ((~i_10_101_2705_0 & ~i_10_101_3070_0 & ~i_10_101_4122_0 & ~i_10_101_4125_0) | (~i_10_101_176_0 & ~i_10_101_796_0 & ~i_10_101_1825_0 & ~i_10_101_4123_0 & ~i_10_101_4287_0 & ~i_10_101_2703_0 & ~i_10_101_3540_0))) | (~i_10_101_1825_0 & ~i_10_101_2005_0 & ~i_10_101_2831_0 & ~i_10_101_3384_0 & i_10_101_3612_0 & ~i_10_101_3856_0 & ~i_10_101_4125_0))) | (~i_10_101_4122_0 & ((i_10_101_1825_0 & i_10_101_2628_0 & i_10_101_2629_0 & ~i_10_101_2729_0) | (~i_10_101_1085_0 & ~i_10_101_1349_0 & ~i_10_101_2783_0 & ~i_10_101_3280_0 & ~i_10_101_3522_0 & ~i_10_101_3647_0 & ~i_10_101_4125_0 & ~i_10_101_4168_0))) | (i_10_101_434_0 & ~i_10_101_1341_0 & ~i_10_101_2630_0 & ~i_10_101_2661_0 & ~i_10_101_3069_0) | (i_10_101_2923_0 & i_10_101_3198_0 & ~i_10_101_3270_0) | (~i_10_101_2365_0 & i_10_101_2631_0 & i_10_101_3384_0 & ~i_10_101_3839_0 & i_10_101_3853_0 & i_10_101_3856_0));
endmodule



// Benchmark "kernel_10_102" written by ABC on Sun Jul 19 10:22:45 2020

module kernel_10_102 ( 
    i_10_102_27_0, i_10_102_31_0, i_10_102_81_0, i_10_102_121_0,
    i_10_102_126_0, i_10_102_172_0, i_10_102_174_0, i_10_102_181_0,
    i_10_102_182_0, i_10_102_281_0, i_10_102_282_0, i_10_102_324_0,
    i_10_102_370_0, i_10_102_373_0, i_10_102_387_0, i_10_102_432_0,
    i_10_102_433_0, i_10_102_445_0, i_10_102_495_0, i_10_102_516_0,
    i_10_102_684_0, i_10_102_931_0, i_10_102_957_0, i_10_102_960_0,
    i_10_102_961_0, i_10_102_1086_0, i_10_102_1233_0, i_10_102_1236_0,
    i_10_102_1237_0, i_10_102_1324_0, i_10_102_1362_0, i_10_102_1364_0,
    i_10_102_1432_0, i_10_102_1530_0, i_10_102_1543_0, i_10_102_1548_0,
    i_10_102_1683_0, i_10_102_1687_0, i_10_102_1822_0, i_10_102_1824_0,
    i_10_102_1825_0, i_10_102_1917_0, i_10_102_1936_0, i_10_102_1939_0,
    i_10_102_1944_0, i_10_102_1945_0, i_10_102_1948_0, i_10_102_1949_0,
    i_10_102_1954_0, i_10_102_2025_0, i_10_102_2179_0, i_10_102_2304_0,
    i_10_102_2305_0, i_10_102_2329_0, i_10_102_2361_0, i_10_102_2377_0,
    i_10_102_2403_0, i_10_102_2453_0, i_10_102_2539_0, i_10_102_2556_0,
    i_10_102_2612_0, i_10_102_2820_0, i_10_102_2827_0, i_10_102_2828_0,
    i_10_102_2910_0, i_10_102_2911_0, i_10_102_3007_0, i_10_102_3042_0,
    i_10_102_3087_0, i_10_102_3088_0, i_10_102_3234_0, i_10_102_3313_0,
    i_10_102_3351_0, i_10_102_3438_0, i_10_102_3439_0, i_10_102_3447_0,
    i_10_102_3465_0, i_10_102_3466_0, i_10_102_3519_0, i_10_102_3582_0,
    i_10_102_3585_0, i_10_102_3615_0, i_10_102_3649_0, i_10_102_3786_0,
    i_10_102_3856_0, i_10_102_3942_0, i_10_102_3943_0, i_10_102_3945_0,
    i_10_102_3982_0, i_10_102_4023_0, i_10_102_4027_0, i_10_102_4230_0,
    i_10_102_4232_0, i_10_102_4369_0, i_10_102_4437_0, i_10_102_4446_0,
    i_10_102_4528_0, i_10_102_4529_0, i_10_102_4566_0, i_10_102_4581_0,
    o_10_102_0_0  );
  input  i_10_102_27_0, i_10_102_31_0, i_10_102_81_0, i_10_102_121_0,
    i_10_102_126_0, i_10_102_172_0, i_10_102_174_0, i_10_102_181_0,
    i_10_102_182_0, i_10_102_281_0, i_10_102_282_0, i_10_102_324_0,
    i_10_102_370_0, i_10_102_373_0, i_10_102_387_0, i_10_102_432_0,
    i_10_102_433_0, i_10_102_445_0, i_10_102_495_0, i_10_102_516_0,
    i_10_102_684_0, i_10_102_931_0, i_10_102_957_0, i_10_102_960_0,
    i_10_102_961_0, i_10_102_1086_0, i_10_102_1233_0, i_10_102_1236_0,
    i_10_102_1237_0, i_10_102_1324_0, i_10_102_1362_0, i_10_102_1364_0,
    i_10_102_1432_0, i_10_102_1530_0, i_10_102_1543_0, i_10_102_1548_0,
    i_10_102_1683_0, i_10_102_1687_0, i_10_102_1822_0, i_10_102_1824_0,
    i_10_102_1825_0, i_10_102_1917_0, i_10_102_1936_0, i_10_102_1939_0,
    i_10_102_1944_0, i_10_102_1945_0, i_10_102_1948_0, i_10_102_1949_0,
    i_10_102_1954_0, i_10_102_2025_0, i_10_102_2179_0, i_10_102_2304_0,
    i_10_102_2305_0, i_10_102_2329_0, i_10_102_2361_0, i_10_102_2377_0,
    i_10_102_2403_0, i_10_102_2453_0, i_10_102_2539_0, i_10_102_2556_0,
    i_10_102_2612_0, i_10_102_2820_0, i_10_102_2827_0, i_10_102_2828_0,
    i_10_102_2910_0, i_10_102_2911_0, i_10_102_3007_0, i_10_102_3042_0,
    i_10_102_3087_0, i_10_102_3088_0, i_10_102_3234_0, i_10_102_3313_0,
    i_10_102_3351_0, i_10_102_3438_0, i_10_102_3439_0, i_10_102_3447_0,
    i_10_102_3465_0, i_10_102_3466_0, i_10_102_3519_0, i_10_102_3582_0,
    i_10_102_3585_0, i_10_102_3615_0, i_10_102_3649_0, i_10_102_3786_0,
    i_10_102_3856_0, i_10_102_3942_0, i_10_102_3943_0, i_10_102_3945_0,
    i_10_102_3982_0, i_10_102_4023_0, i_10_102_4027_0, i_10_102_4230_0,
    i_10_102_4232_0, i_10_102_4369_0, i_10_102_4437_0, i_10_102_4446_0,
    i_10_102_4528_0, i_10_102_4529_0, i_10_102_4566_0, i_10_102_4581_0;
  output o_10_102_0_0;
  assign o_10_102_0_0 = ~(i_10_102_174_0 | (~i_10_102_3087_0 & ~i_10_102_3088_0) | (~i_10_102_27_0 & ~i_10_102_1233_0) | (~i_10_102_387_0 & i_10_102_1822_0 & ~i_10_102_2612_0) | (~i_10_102_957_0 & ~i_10_102_960_0 & ~i_10_102_961_0 & ~i_10_102_2453_0));
endmodule



// Benchmark "kernel_10_103" written by ABC on Sun Jul 19 10:22:46 2020

module kernel_10_103 ( 
    i_10_103_216_0, i_10_103_218_0, i_10_103_247_0, i_10_103_279_0,
    i_10_103_284_0, i_10_103_319_0, i_10_103_429_0, i_10_103_430_0,
    i_10_103_435_0, i_10_103_438_0, i_10_103_439_0, i_10_103_449_0,
    i_10_103_463_0, i_10_103_466_0, i_10_103_748_0, i_10_103_961_0,
    i_10_103_993_0, i_10_103_996_0, i_10_103_1059_0, i_10_103_1238_0,
    i_10_103_1250_0, i_10_103_1354_0, i_10_103_1357_0, i_10_103_1556_0,
    i_10_103_1684_0, i_10_103_1685_0, i_10_103_1756_0, i_10_103_1818_0,
    i_10_103_1821_0, i_10_103_1824_0, i_10_103_1825_0, i_10_103_1912_0,
    i_10_103_1916_0, i_10_103_1947_0, i_10_103_1990_0, i_10_103_2312_0,
    i_10_103_2353_0, i_10_103_2355_0, i_10_103_2373_0, i_10_103_2451_0,
    i_10_103_2452_0, i_10_103_2454_0, i_10_103_2469_0, i_10_103_2514_0,
    i_10_103_2516_0, i_10_103_2546_0, i_10_103_2659_0, i_10_103_2660_0,
    i_10_103_2701_0, i_10_103_2704_0, i_10_103_2711_0, i_10_103_2720_0,
    i_10_103_2728_0, i_10_103_2729_0, i_10_103_2820_0, i_10_103_2821_0,
    i_10_103_2884_0, i_10_103_3039_0, i_10_103_3049_0, i_10_103_3093_0,
    i_10_103_3094_0, i_10_103_3174_0, i_10_103_3195_0, i_10_103_3235_0,
    i_10_103_3271_0, i_10_103_3279_0, i_10_103_3280_0, i_10_103_3281_0,
    i_10_103_3282_0, i_10_103_3283_0, i_10_103_3292_0, i_10_103_3318_0,
    i_10_103_3384_0, i_10_103_3385_0, i_10_103_3388_0, i_10_103_3389_0,
    i_10_103_3390_0, i_10_103_3525_0, i_10_103_3526_0, i_10_103_3616_0,
    i_10_103_3617_0, i_10_103_3685_0, i_10_103_3702_0, i_10_103_3705_0,
    i_10_103_3850_0, i_10_103_3857_0, i_10_103_3859_0, i_10_103_3885_0,
    i_10_103_3902_0, i_10_103_3946_0, i_10_103_4027_0, i_10_103_4031_0,
    i_10_103_4056_0, i_10_103_4116_0, i_10_103_4117_0, i_10_103_4213_0,
    i_10_103_4271_0, i_10_103_4567_0, i_10_103_4568_0, i_10_103_4589_0,
    o_10_103_0_0  );
  input  i_10_103_216_0, i_10_103_218_0, i_10_103_247_0, i_10_103_279_0,
    i_10_103_284_0, i_10_103_319_0, i_10_103_429_0, i_10_103_430_0,
    i_10_103_435_0, i_10_103_438_0, i_10_103_439_0, i_10_103_449_0,
    i_10_103_463_0, i_10_103_466_0, i_10_103_748_0, i_10_103_961_0,
    i_10_103_993_0, i_10_103_996_0, i_10_103_1059_0, i_10_103_1238_0,
    i_10_103_1250_0, i_10_103_1354_0, i_10_103_1357_0, i_10_103_1556_0,
    i_10_103_1684_0, i_10_103_1685_0, i_10_103_1756_0, i_10_103_1818_0,
    i_10_103_1821_0, i_10_103_1824_0, i_10_103_1825_0, i_10_103_1912_0,
    i_10_103_1916_0, i_10_103_1947_0, i_10_103_1990_0, i_10_103_2312_0,
    i_10_103_2353_0, i_10_103_2355_0, i_10_103_2373_0, i_10_103_2451_0,
    i_10_103_2452_0, i_10_103_2454_0, i_10_103_2469_0, i_10_103_2514_0,
    i_10_103_2516_0, i_10_103_2546_0, i_10_103_2659_0, i_10_103_2660_0,
    i_10_103_2701_0, i_10_103_2704_0, i_10_103_2711_0, i_10_103_2720_0,
    i_10_103_2728_0, i_10_103_2729_0, i_10_103_2820_0, i_10_103_2821_0,
    i_10_103_2884_0, i_10_103_3039_0, i_10_103_3049_0, i_10_103_3093_0,
    i_10_103_3094_0, i_10_103_3174_0, i_10_103_3195_0, i_10_103_3235_0,
    i_10_103_3271_0, i_10_103_3279_0, i_10_103_3280_0, i_10_103_3281_0,
    i_10_103_3282_0, i_10_103_3283_0, i_10_103_3292_0, i_10_103_3318_0,
    i_10_103_3384_0, i_10_103_3385_0, i_10_103_3388_0, i_10_103_3389_0,
    i_10_103_3390_0, i_10_103_3525_0, i_10_103_3526_0, i_10_103_3616_0,
    i_10_103_3617_0, i_10_103_3685_0, i_10_103_3702_0, i_10_103_3705_0,
    i_10_103_3850_0, i_10_103_3857_0, i_10_103_3859_0, i_10_103_3885_0,
    i_10_103_3902_0, i_10_103_3946_0, i_10_103_4027_0, i_10_103_4031_0,
    i_10_103_4056_0, i_10_103_4116_0, i_10_103_4117_0, i_10_103_4213_0,
    i_10_103_4271_0, i_10_103_4567_0, i_10_103_4568_0, i_10_103_4589_0;
  output o_10_103_0_0;
  assign o_10_103_0_0 = 0;
endmodule



// Benchmark "kernel_10_104" written by ABC on Sun Jul 19 10:22:46 2020

module kernel_10_104 ( 
    i_10_104_117_0, i_10_104_118_0, i_10_104_220_0, i_10_104_315_0,
    i_10_104_316_0, i_10_104_387_0, i_10_104_388_0, i_10_104_389_0,
    i_10_104_391_0, i_10_104_394_0, i_10_104_408_0, i_10_104_427_0,
    i_10_104_436_0, i_10_104_462_0, i_10_104_532_0, i_10_104_795_0,
    i_10_104_819_0, i_10_104_824_0, i_10_104_958_0, i_10_104_999_0,
    i_10_104_1000_0, i_10_104_1026_0, i_10_104_1080_0, i_10_104_1236_0,
    i_10_104_1296_0, i_10_104_1305_0, i_10_104_1306_0, i_10_104_1308_0,
    i_10_104_1378_0, i_10_104_1431_0, i_10_104_1448_0, i_10_104_1543_0,
    i_10_104_1575_0, i_10_104_1576_0, i_10_104_1578_0, i_10_104_1621_0,
    i_10_104_1651_0, i_10_104_1683_0, i_10_104_1684_0, i_10_104_1685_0,
    i_10_104_1729_0, i_10_104_1732_0, i_10_104_1733_0, i_10_104_1764_0,
    i_10_104_1819_0, i_10_104_2022_0, i_10_104_2028_0, i_10_104_2200_0,
    i_10_104_2203_0, i_10_104_2204_0, i_10_104_2250_0, i_10_104_2352_0,
    i_10_104_2377_0, i_10_104_2405_0, i_10_104_2410_0, i_10_104_2452_0,
    i_10_104_2454_0, i_10_104_2455_0, i_10_104_2467_0, i_10_104_2540_0,
    i_10_104_2556_0, i_10_104_2565_0, i_10_104_2628_0, i_10_104_2629_0,
    i_10_104_2719_0, i_10_104_2727_0, i_10_104_2729_0, i_10_104_2781_0,
    i_10_104_2782_0, i_10_104_2785_0, i_10_104_2863_0, i_10_104_2880_0,
    i_10_104_2980_0, i_10_104_3042_0, i_10_104_3195_0, i_10_104_3313_0,
    i_10_104_3389_0, i_10_104_3392_0, i_10_104_3466_0, i_10_104_3469_0,
    i_10_104_3501_0, i_10_104_3522_0, i_10_104_3550_0, i_10_104_3559_0,
    i_10_104_3582_0, i_10_104_3583_0, i_10_104_3840_0, i_10_104_3841_0,
    i_10_104_3857_0, i_10_104_4006_0, i_10_104_4023_0, i_10_104_4024_0,
    i_10_104_4113_0, i_10_104_4115_0, i_10_104_4117_0, i_10_104_4118_0,
    i_10_104_4204_0, i_10_104_4275_0, i_10_104_4289_0, i_10_104_4581_0,
    o_10_104_0_0  );
  input  i_10_104_117_0, i_10_104_118_0, i_10_104_220_0, i_10_104_315_0,
    i_10_104_316_0, i_10_104_387_0, i_10_104_388_0, i_10_104_389_0,
    i_10_104_391_0, i_10_104_394_0, i_10_104_408_0, i_10_104_427_0,
    i_10_104_436_0, i_10_104_462_0, i_10_104_532_0, i_10_104_795_0,
    i_10_104_819_0, i_10_104_824_0, i_10_104_958_0, i_10_104_999_0,
    i_10_104_1000_0, i_10_104_1026_0, i_10_104_1080_0, i_10_104_1236_0,
    i_10_104_1296_0, i_10_104_1305_0, i_10_104_1306_0, i_10_104_1308_0,
    i_10_104_1378_0, i_10_104_1431_0, i_10_104_1448_0, i_10_104_1543_0,
    i_10_104_1575_0, i_10_104_1576_0, i_10_104_1578_0, i_10_104_1621_0,
    i_10_104_1651_0, i_10_104_1683_0, i_10_104_1684_0, i_10_104_1685_0,
    i_10_104_1729_0, i_10_104_1732_0, i_10_104_1733_0, i_10_104_1764_0,
    i_10_104_1819_0, i_10_104_2022_0, i_10_104_2028_0, i_10_104_2200_0,
    i_10_104_2203_0, i_10_104_2204_0, i_10_104_2250_0, i_10_104_2352_0,
    i_10_104_2377_0, i_10_104_2405_0, i_10_104_2410_0, i_10_104_2452_0,
    i_10_104_2454_0, i_10_104_2455_0, i_10_104_2467_0, i_10_104_2540_0,
    i_10_104_2556_0, i_10_104_2565_0, i_10_104_2628_0, i_10_104_2629_0,
    i_10_104_2719_0, i_10_104_2727_0, i_10_104_2729_0, i_10_104_2781_0,
    i_10_104_2782_0, i_10_104_2785_0, i_10_104_2863_0, i_10_104_2880_0,
    i_10_104_2980_0, i_10_104_3042_0, i_10_104_3195_0, i_10_104_3313_0,
    i_10_104_3389_0, i_10_104_3392_0, i_10_104_3466_0, i_10_104_3469_0,
    i_10_104_3501_0, i_10_104_3522_0, i_10_104_3550_0, i_10_104_3559_0,
    i_10_104_3582_0, i_10_104_3583_0, i_10_104_3840_0, i_10_104_3841_0,
    i_10_104_3857_0, i_10_104_4006_0, i_10_104_4023_0, i_10_104_4024_0,
    i_10_104_4113_0, i_10_104_4115_0, i_10_104_4117_0, i_10_104_4118_0,
    i_10_104_4204_0, i_10_104_4275_0, i_10_104_4289_0, i_10_104_4581_0;
  output o_10_104_0_0;
  assign o_10_104_0_0 = 0;
endmodule



// Benchmark "kernel_10_105" written by ABC on Sun Jul 19 10:22:47 2020

module kernel_10_105 ( 
    i_10_105_37_0, i_10_105_256_0, i_10_105_283_0, i_10_105_318_0,
    i_10_105_322_0, i_10_105_324_0, i_10_105_325_0, i_10_105_328_0,
    i_10_105_405_0, i_10_105_441_0, i_10_105_444_0, i_10_105_460_0,
    i_10_105_464_0, i_10_105_588_0, i_10_105_894_0, i_10_105_954_0,
    i_10_105_993_0, i_10_105_1003_0, i_10_105_1031_0, i_10_105_1086_0,
    i_10_105_1241_0, i_10_105_1377_0, i_10_105_1378_0, i_10_105_1435_0,
    i_10_105_1542_0, i_10_105_1543_0, i_10_105_1546_0, i_10_105_1579_0,
    i_10_105_1580_0, i_10_105_1581_0, i_10_105_1582_0, i_10_105_1596_0,
    i_10_105_1612_0, i_10_105_1647_0, i_10_105_1648_0, i_10_105_1649_0,
    i_10_105_1654_0, i_10_105_1689_0, i_10_105_1768_0, i_10_105_1822_0,
    i_10_105_1824_0, i_10_105_1825_0, i_10_105_1947_0, i_10_105_1948_0,
    i_10_105_1992_0, i_10_105_1995_0, i_10_105_2200_0, i_10_105_2203_0,
    i_10_105_2242_0, i_10_105_2309_0, i_10_105_2330_0, i_10_105_2352_0,
    i_10_105_2353_0, i_10_105_2356_0, i_10_105_2364_0, i_10_105_2452_0,
    i_10_105_2453_0, i_10_105_2454_0, i_10_105_2455_0, i_10_105_2458_0,
    i_10_105_2471_0, i_10_105_2473_0, i_10_105_2541_0, i_10_105_2604_0,
    i_10_105_2607_0, i_10_105_2658_0, i_10_105_2714_0, i_10_105_2787_0,
    i_10_105_2829_0, i_10_105_2831_0, i_10_105_2917_0, i_10_105_2982_0,
    i_10_105_3270_0, i_10_105_3274_0, i_10_105_3281_0, i_10_105_3282_0,
    i_10_105_3525_0, i_10_105_3526_0, i_10_105_3614_0, i_10_105_3616_0,
    i_10_105_3683_0, i_10_105_3780_0, i_10_105_3787_0, i_10_105_3840_0,
    i_10_105_3841_0, i_10_105_3848_0, i_10_105_3854_0, i_10_105_3857_0,
    i_10_105_3859_0, i_10_105_3891_0, i_10_105_3893_0, i_10_105_3979_0,
    i_10_105_3982_0, i_10_105_4233_0, i_10_105_4287_0, i_10_105_4292_0,
    i_10_105_4456_0, i_10_105_4459_0, i_10_105_4566_0, i_10_105_4570_0,
    o_10_105_0_0  );
  input  i_10_105_37_0, i_10_105_256_0, i_10_105_283_0, i_10_105_318_0,
    i_10_105_322_0, i_10_105_324_0, i_10_105_325_0, i_10_105_328_0,
    i_10_105_405_0, i_10_105_441_0, i_10_105_444_0, i_10_105_460_0,
    i_10_105_464_0, i_10_105_588_0, i_10_105_894_0, i_10_105_954_0,
    i_10_105_993_0, i_10_105_1003_0, i_10_105_1031_0, i_10_105_1086_0,
    i_10_105_1241_0, i_10_105_1377_0, i_10_105_1378_0, i_10_105_1435_0,
    i_10_105_1542_0, i_10_105_1543_0, i_10_105_1546_0, i_10_105_1579_0,
    i_10_105_1580_0, i_10_105_1581_0, i_10_105_1582_0, i_10_105_1596_0,
    i_10_105_1612_0, i_10_105_1647_0, i_10_105_1648_0, i_10_105_1649_0,
    i_10_105_1654_0, i_10_105_1689_0, i_10_105_1768_0, i_10_105_1822_0,
    i_10_105_1824_0, i_10_105_1825_0, i_10_105_1947_0, i_10_105_1948_0,
    i_10_105_1992_0, i_10_105_1995_0, i_10_105_2200_0, i_10_105_2203_0,
    i_10_105_2242_0, i_10_105_2309_0, i_10_105_2330_0, i_10_105_2352_0,
    i_10_105_2353_0, i_10_105_2356_0, i_10_105_2364_0, i_10_105_2452_0,
    i_10_105_2453_0, i_10_105_2454_0, i_10_105_2455_0, i_10_105_2458_0,
    i_10_105_2471_0, i_10_105_2473_0, i_10_105_2541_0, i_10_105_2604_0,
    i_10_105_2607_0, i_10_105_2658_0, i_10_105_2714_0, i_10_105_2787_0,
    i_10_105_2829_0, i_10_105_2831_0, i_10_105_2917_0, i_10_105_2982_0,
    i_10_105_3270_0, i_10_105_3274_0, i_10_105_3281_0, i_10_105_3282_0,
    i_10_105_3525_0, i_10_105_3526_0, i_10_105_3614_0, i_10_105_3616_0,
    i_10_105_3683_0, i_10_105_3780_0, i_10_105_3787_0, i_10_105_3840_0,
    i_10_105_3841_0, i_10_105_3848_0, i_10_105_3854_0, i_10_105_3857_0,
    i_10_105_3859_0, i_10_105_3891_0, i_10_105_3893_0, i_10_105_3979_0,
    i_10_105_3982_0, i_10_105_4233_0, i_10_105_4287_0, i_10_105_4292_0,
    i_10_105_4456_0, i_10_105_4459_0, i_10_105_4566_0, i_10_105_4570_0;
  output o_10_105_0_0;
  assign o_10_105_0_0 = 0;
endmodule



// Benchmark "kernel_10_106" written by ABC on Sun Jul 19 10:22:49 2020

module kernel_10_106 ( 
    i_10_106_175_0, i_10_106_268_0, i_10_106_280_0, i_10_106_285_0,
    i_10_106_296_0, i_10_106_316_0, i_10_106_317_0, i_10_106_327_0,
    i_10_106_328_0, i_10_106_329_0, i_10_106_409_0, i_10_106_439_0,
    i_10_106_443_0, i_10_106_453_0, i_10_106_516_0, i_10_106_520_0,
    i_10_106_749_0, i_10_106_800_0, i_10_106_999_0, i_10_106_1080_0,
    i_10_106_1081_0, i_10_106_1217_0, i_10_106_1233_0, i_10_106_1234_0,
    i_10_106_1238_0, i_10_106_1263_0, i_10_106_1264_0, i_10_106_1265_0,
    i_10_106_1366_0, i_10_106_1438_0, i_10_106_1439_0, i_10_106_1448_0,
    i_10_106_1546_0, i_10_106_1615_0, i_10_106_1684_0, i_10_106_1687_0,
    i_10_106_1688_0, i_10_106_1818_0, i_10_106_1819_0, i_10_106_1821_0,
    i_10_106_1822_0, i_10_106_1826_0, i_10_106_2337_0, i_10_106_2351_0,
    i_10_106_2352_0, i_10_106_2353_0, i_10_106_2354_0, i_10_106_2408_0,
    i_10_106_2461_0, i_10_106_2470_0, i_10_106_2606_0, i_10_106_2655_0,
    i_10_106_2658_0, i_10_106_2659_0, i_10_106_2660_0, i_10_106_2680_0,
    i_10_106_2707_0, i_10_106_2722_0, i_10_106_2723_0, i_10_106_2729_0,
    i_10_106_2827_0, i_10_106_2828_0, i_10_106_2831_0, i_10_106_2885_0,
    i_10_106_2979_0, i_10_106_2980_0, i_10_106_2981_0, i_10_106_2985_0,
    i_10_106_2986_0, i_10_106_2987_0, i_10_106_3070_0, i_10_106_3074_0,
    i_10_106_3157_0, i_10_106_3158_0, i_10_106_3198_0, i_10_106_3199_0,
    i_10_106_3200_0, i_10_106_3201_0, i_10_106_3274_0, i_10_106_3280_0,
    i_10_106_3281_0, i_10_106_3384_0, i_10_106_3385_0, i_10_106_3388_0,
    i_10_106_3493_0, i_10_106_3496_0, i_10_106_3497_0, i_10_106_3522_0,
    i_10_106_3583_0, i_10_106_3837_0, i_10_106_3851_0, i_10_106_3858_0,
    i_10_106_3872_0, i_10_106_3896_0, i_10_106_3906_0, i_10_106_3979_0,
    i_10_106_4266_0, i_10_106_4270_0, i_10_106_4277_0, i_10_106_4279_0,
    o_10_106_0_0  );
  input  i_10_106_175_0, i_10_106_268_0, i_10_106_280_0, i_10_106_285_0,
    i_10_106_296_0, i_10_106_316_0, i_10_106_317_0, i_10_106_327_0,
    i_10_106_328_0, i_10_106_329_0, i_10_106_409_0, i_10_106_439_0,
    i_10_106_443_0, i_10_106_453_0, i_10_106_516_0, i_10_106_520_0,
    i_10_106_749_0, i_10_106_800_0, i_10_106_999_0, i_10_106_1080_0,
    i_10_106_1081_0, i_10_106_1217_0, i_10_106_1233_0, i_10_106_1234_0,
    i_10_106_1238_0, i_10_106_1263_0, i_10_106_1264_0, i_10_106_1265_0,
    i_10_106_1366_0, i_10_106_1438_0, i_10_106_1439_0, i_10_106_1448_0,
    i_10_106_1546_0, i_10_106_1615_0, i_10_106_1684_0, i_10_106_1687_0,
    i_10_106_1688_0, i_10_106_1818_0, i_10_106_1819_0, i_10_106_1821_0,
    i_10_106_1822_0, i_10_106_1826_0, i_10_106_2337_0, i_10_106_2351_0,
    i_10_106_2352_0, i_10_106_2353_0, i_10_106_2354_0, i_10_106_2408_0,
    i_10_106_2461_0, i_10_106_2470_0, i_10_106_2606_0, i_10_106_2655_0,
    i_10_106_2658_0, i_10_106_2659_0, i_10_106_2660_0, i_10_106_2680_0,
    i_10_106_2707_0, i_10_106_2722_0, i_10_106_2723_0, i_10_106_2729_0,
    i_10_106_2827_0, i_10_106_2828_0, i_10_106_2831_0, i_10_106_2885_0,
    i_10_106_2979_0, i_10_106_2980_0, i_10_106_2981_0, i_10_106_2985_0,
    i_10_106_2986_0, i_10_106_2987_0, i_10_106_3070_0, i_10_106_3074_0,
    i_10_106_3157_0, i_10_106_3158_0, i_10_106_3198_0, i_10_106_3199_0,
    i_10_106_3200_0, i_10_106_3201_0, i_10_106_3274_0, i_10_106_3280_0,
    i_10_106_3281_0, i_10_106_3384_0, i_10_106_3385_0, i_10_106_3388_0,
    i_10_106_3493_0, i_10_106_3496_0, i_10_106_3497_0, i_10_106_3522_0,
    i_10_106_3583_0, i_10_106_3837_0, i_10_106_3851_0, i_10_106_3858_0,
    i_10_106_3872_0, i_10_106_3896_0, i_10_106_3906_0, i_10_106_3979_0,
    i_10_106_4266_0, i_10_106_4270_0, i_10_106_4277_0, i_10_106_4279_0;
  output o_10_106_0_0;
  assign o_10_106_0_0 = ~((i_10_106_175_0 & ~i_10_106_3896_0 & ((i_10_106_516_0 & i_10_106_1818_0 & ~i_10_106_2828_0) | (~i_10_106_1366_0 & ~i_10_106_1821_0 & ~i_10_106_2606_0 & ~i_10_106_2723_0 & ~i_10_106_2729_0 & ~i_10_106_2981_0 & ~i_10_106_4270_0))) | (~i_10_106_329_0 & ((~i_10_106_327_0 & ~i_10_106_2827_0 & ~i_10_106_2980_0 & ~i_10_106_2986_0 & ~i_10_106_3201_0 & ~i_10_106_3497_0) | (~i_10_106_328_0 & ~i_10_106_1081_0 & ~i_10_106_2337_0 & ~i_10_106_2658_0 & i_10_106_3979_0))) | (~i_10_106_327_0 & ((~i_10_106_317_0 & ~i_10_106_409_0 & ~i_10_106_800_0 & ~i_10_106_1615_0 & ~i_10_106_2606_0 & ~i_10_106_2986_0 & ~i_10_106_3384_0) | (~i_10_106_749_0 & ~i_10_106_1264_0 & ~i_10_106_2337_0 & ~i_10_106_2354_0 & ~i_10_106_3388_0 & ~i_10_106_3496_0 & ~i_10_106_3906_0))) | (~i_10_106_3497_0 & ((~i_10_106_1263_0 & ((~i_10_106_1080_0 & ~i_10_106_2707_0 & ~i_10_106_4277_0 & ((~i_10_106_296_0 & ~i_10_106_2352_0 & ~i_10_106_2408_0 & ~i_10_106_2680_0 & ~i_10_106_3274_0) | (~i_10_106_1265_0 & ~i_10_106_2985_0 & ~i_10_106_3851_0))) | (~i_10_106_316_0 & ~i_10_106_1265_0 & ~i_10_106_1822_0 & ~i_10_106_2337_0 & ~i_10_106_2408_0 & ~i_10_106_2461_0 & ~i_10_106_2986_0))) | (~i_10_106_3496_0 & ((~i_10_106_409_0 & ~i_10_106_2353_0 & ~i_10_106_2828_0 & ~i_10_106_3198_0 & ~i_10_106_3385_0 & ~i_10_106_3906_0) | (~i_10_106_1081_0 & ~i_10_106_1265_0 & ~i_10_106_1821_0 & ~i_10_106_2680_0 & ~i_10_106_2707_0 & ~i_10_106_2985_0 & ~i_10_106_3979_0))))) | (~i_10_106_3496_0 & ((~i_10_106_1081_0 & ((~i_10_106_1264_0 & ~i_10_106_1265_0 & ~i_10_106_2680_0 & ~i_10_106_2979_0 & ~i_10_106_2981_0 & ~i_10_106_2986_0) | (i_10_106_516_0 & ~i_10_106_1263_0 & ~i_10_106_2351_0 & ~i_10_106_2722_0 & ~i_10_106_2723_0 & ~i_10_106_2729_0 & ~i_10_106_3274_0))) | (~i_10_106_285_0 & ~i_10_106_520_0 & ~i_10_106_2660_0 & ~i_10_106_2831_0 & ~i_10_106_2979_0 & ~i_10_106_3906_0))) | (i_10_106_3280_0 & ((i_10_106_439_0 & ~i_10_106_2986_0 & ~i_10_106_3281_0) | (~i_10_106_2828_0 & i_10_106_3522_0 & ~i_10_106_3906_0))));
endmodule



// Benchmark "kernel_10_107" written by ABC on Sun Jul 19 10:22:50 2020

module kernel_10_107 ( 
    i_10_107_176_0, i_10_107_187_0, i_10_107_283_0, i_10_107_319_0,
    i_10_107_390_0, i_10_107_391_0, i_10_107_392_0, i_10_107_405_0,
    i_10_107_409_0, i_10_107_424_0, i_10_107_426_0, i_10_107_427_0,
    i_10_107_433_0, i_10_107_434_0, i_10_107_459_0, i_10_107_462_0,
    i_10_107_794_0, i_10_107_991_0, i_10_107_1026_0, i_10_107_1027_0,
    i_10_107_1031_0, i_10_107_1043_0, i_10_107_1081_0, i_10_107_1135_0,
    i_10_107_1306_0, i_10_107_1442_0, i_10_107_1540_0, i_10_107_1541_0,
    i_10_107_1548_0, i_10_107_1575_0, i_10_107_1577_0, i_10_107_1651_0,
    i_10_107_1683_0, i_10_107_1684_0, i_10_107_1685_0, i_10_107_1769_0,
    i_10_107_1825_0, i_10_107_1990_0, i_10_107_2349_0, i_10_107_2353_0,
    i_10_107_2356_0, i_10_107_2360_0, i_10_107_2404_0, i_10_107_2448_0,
    i_10_107_2631_0, i_10_107_2632_0, i_10_107_2633_0, i_10_107_2673_0,
    i_10_107_2674_0, i_10_107_2675_0, i_10_107_2681_0, i_10_107_2701_0,
    i_10_107_2703_0, i_10_107_2723_0, i_10_107_2727_0, i_10_107_2783_0,
    i_10_107_2887_0, i_10_107_2918_0, i_10_107_2921_0, i_10_107_3069_0,
    i_10_107_3071_0, i_10_107_3073_0, i_10_107_3152_0, i_10_107_3153_0,
    i_10_107_3156_0, i_10_107_3158_0, i_10_107_3268_0, i_10_107_3269_0,
    i_10_107_3322_0, i_10_107_3328_0, i_10_107_3330_0, i_10_107_3406_0,
    i_10_107_3585_0, i_10_107_3586_0, i_10_107_3612_0, i_10_107_3614_0,
    i_10_107_3616_0, i_10_107_3649_0, i_10_107_3780_0, i_10_107_3782_0,
    i_10_107_3783_0, i_10_107_3784_0, i_10_107_3785_0, i_10_107_3835_0,
    i_10_107_3837_0, i_10_107_3838_0, i_10_107_3839_0, i_10_107_3855_0,
    i_10_107_3856_0, i_10_107_3857_0, i_10_107_3980_0, i_10_107_4117_0,
    i_10_107_4118_0, i_10_107_4119_0, i_10_107_4120_0, i_10_107_4121_0,
    i_10_107_4266_0, i_10_107_4276_0, i_10_107_4288_0, i_10_107_4567_0,
    o_10_107_0_0  );
  input  i_10_107_176_0, i_10_107_187_0, i_10_107_283_0, i_10_107_319_0,
    i_10_107_390_0, i_10_107_391_0, i_10_107_392_0, i_10_107_405_0,
    i_10_107_409_0, i_10_107_424_0, i_10_107_426_0, i_10_107_427_0,
    i_10_107_433_0, i_10_107_434_0, i_10_107_459_0, i_10_107_462_0,
    i_10_107_794_0, i_10_107_991_0, i_10_107_1026_0, i_10_107_1027_0,
    i_10_107_1031_0, i_10_107_1043_0, i_10_107_1081_0, i_10_107_1135_0,
    i_10_107_1306_0, i_10_107_1442_0, i_10_107_1540_0, i_10_107_1541_0,
    i_10_107_1548_0, i_10_107_1575_0, i_10_107_1577_0, i_10_107_1651_0,
    i_10_107_1683_0, i_10_107_1684_0, i_10_107_1685_0, i_10_107_1769_0,
    i_10_107_1825_0, i_10_107_1990_0, i_10_107_2349_0, i_10_107_2353_0,
    i_10_107_2356_0, i_10_107_2360_0, i_10_107_2404_0, i_10_107_2448_0,
    i_10_107_2631_0, i_10_107_2632_0, i_10_107_2633_0, i_10_107_2673_0,
    i_10_107_2674_0, i_10_107_2675_0, i_10_107_2681_0, i_10_107_2701_0,
    i_10_107_2703_0, i_10_107_2723_0, i_10_107_2727_0, i_10_107_2783_0,
    i_10_107_2887_0, i_10_107_2918_0, i_10_107_2921_0, i_10_107_3069_0,
    i_10_107_3071_0, i_10_107_3073_0, i_10_107_3152_0, i_10_107_3153_0,
    i_10_107_3156_0, i_10_107_3158_0, i_10_107_3268_0, i_10_107_3269_0,
    i_10_107_3322_0, i_10_107_3328_0, i_10_107_3330_0, i_10_107_3406_0,
    i_10_107_3585_0, i_10_107_3586_0, i_10_107_3612_0, i_10_107_3614_0,
    i_10_107_3616_0, i_10_107_3649_0, i_10_107_3780_0, i_10_107_3782_0,
    i_10_107_3783_0, i_10_107_3784_0, i_10_107_3785_0, i_10_107_3835_0,
    i_10_107_3837_0, i_10_107_3838_0, i_10_107_3839_0, i_10_107_3855_0,
    i_10_107_3856_0, i_10_107_3857_0, i_10_107_3980_0, i_10_107_4117_0,
    i_10_107_4118_0, i_10_107_4119_0, i_10_107_4120_0, i_10_107_4121_0,
    i_10_107_4266_0, i_10_107_4276_0, i_10_107_4288_0, i_10_107_4567_0;
  output o_10_107_0_0;
  assign o_10_107_0_0 = ~((~i_10_107_3783_0 & ((i_10_107_283_0 & ~i_10_107_1541_0 & ((~i_10_107_187_0 & ~i_10_107_391_0 & ~i_10_107_1575_0 & ~i_10_107_1769_0 & ~i_10_107_2349_0 & ~i_10_107_3069_0) | (~i_10_107_1026_0 & ~i_10_107_1027_0 & ~i_10_107_3614_0 & ~i_10_107_3616_0 & ~i_10_107_3857_0 & ~i_10_107_4266_0))) | (~i_10_107_409_0 & ~i_10_107_2727_0 & ~i_10_107_4276_0 & ((~i_10_107_1027_0 & ~i_10_107_1540_0 & ~i_10_107_1769_0 & ~i_10_107_2681_0 & ~i_10_107_3069_0 & ~i_10_107_3269_0 & i_10_107_3835_0) | (~i_10_107_392_0 & ~i_10_107_462_0 & ~i_10_107_1306_0 & ~i_10_107_1548_0 & ~i_10_107_3612_0 & ~i_10_107_3614_0 & ~i_10_107_4118_0 & ~i_10_107_4121_0))) | (i_10_107_3586_0 & i_10_107_3784_0) | (~i_10_107_426_0 & ~i_10_107_1540_0 & ~i_10_107_1684_0 & ~i_10_107_1769_0 & i_10_107_2632_0 & ~i_10_107_2723_0 & ~i_10_107_3585_0 & ~i_10_107_4266_0))) | (~i_10_107_187_0 & ((~i_10_107_391_0 & ~i_10_107_1027_0 & i_10_107_4120_0) | (~i_10_107_1043_0 & ~i_10_107_1540_0 & ~i_10_107_1685_0 & ~i_10_107_3069_0 & ~i_10_107_3614_0 & ~i_10_107_3649_0 & ~i_10_107_4266_0))) | (~i_10_107_283_0 & ((~i_10_107_1026_0 & ~i_10_107_1685_0 & ~i_10_107_3073_0 & ~i_10_107_3782_0 & ~i_10_107_3855_0) | (~i_10_107_390_0 & ~i_10_107_1577_0 & ~i_10_107_1684_0 & ~i_10_107_2448_0 & ~i_10_107_3614_0 & ~i_10_107_3780_0 & ~i_10_107_4276_0))) | (~i_10_107_1043_0 & ((~i_10_107_794_0 & ~i_10_107_1540_0 & i_10_107_2631_0 & i_10_107_2727_0 & ~i_10_107_3073_0 & ~i_10_107_3585_0) | (~i_10_107_1026_0 & ~i_10_107_1541_0 & ~i_10_107_1683_0 & ~i_10_107_1769_0 & ~i_10_107_3784_0 & ~i_10_107_3855_0))) | (~i_10_107_3785_0 & ((i_10_107_1306_0 & ~i_10_107_1575_0 & ((~i_10_107_1540_0 & ~i_10_107_3268_0 & ~i_10_107_3857_0) | (~i_10_107_1683_0 & i_10_107_4288_0))) | (~i_10_107_3069_0 & ((~i_10_107_1541_0 & ~i_10_107_1684_0 & ~i_10_107_3073_0 & i_10_107_3585_0) | (i_10_107_2356_0 & ~i_10_107_2360_0 & ~i_10_107_3782_0 & ~i_10_107_4288_0))))) | (~i_10_107_3071_0 & ((~i_10_107_3069_0 & ~i_10_107_3406_0 & ~i_10_107_3855_0 & i_10_107_4120_0) | (~i_10_107_1027_0 & ~i_10_107_1651_0 & i_10_107_1825_0 & ~i_10_107_3614_0 & ~i_10_107_3856_0 & ~i_10_107_4276_0))) | (~i_10_107_3069_0 & ((~i_10_107_1027_0 & ((~i_10_107_427_0 & ~i_10_107_1081_0 & ~i_10_107_2703_0 & ~i_10_107_2921_0 & ~i_10_107_3649_0 & i_10_107_3835_0) | (~i_10_107_1540_0 & ~i_10_107_3612_0 & ~i_10_107_3838_0 & ~i_10_107_3839_0))) | (~i_10_107_3612_0 & ((~i_10_107_459_0 & ~i_10_107_1306_0 & ~i_10_107_1540_0 & ~i_10_107_2353_0 & ~i_10_107_2448_0 & i_10_107_4117_0) | (~i_10_107_1031_0 & i_10_107_2356_0 & ~i_10_107_3268_0 & ~i_10_107_3856_0 & i_10_107_4288_0))) | (~i_10_107_462_0 & ~i_10_107_1683_0 & ~i_10_107_1684_0 & ~i_10_107_2349_0 & ~i_10_107_3269_0 & ~i_10_107_3614_0 & i_10_107_3649_0 & ~i_10_107_3839_0))) | (i_10_107_459_0 & ~i_10_107_1540_0 & ~i_10_107_1769_0 & i_10_107_3586_0) | (i_10_107_427_0 & ~i_10_107_2632_0 & ~i_10_107_3614_0) | (i_10_107_2681_0 & ~i_10_107_3835_0 & ~i_10_107_3857_0) | (~i_10_107_1541_0 & i_10_107_2918_0 & ~i_10_107_3586_0 & ~i_10_107_3780_0 & ~i_10_107_4276_0) | (~i_10_107_390_0 & ~i_10_107_409_0 & ~i_10_107_426_0 & ~i_10_107_1685_0 & i_10_107_2632_0 & ~i_10_107_3855_0 & ~i_10_107_4118_0 & ~i_10_107_4288_0));
endmodule



// Benchmark "kernel_10_108" written by ABC on Sun Jul 19 10:22:51 2020

module kernel_10_108 ( 
    i_10_108_123_0, i_10_108_153_0, i_10_108_171_0, i_10_108_175_0,
    i_10_108_244_0, i_10_108_248_0, i_10_108_434_0, i_10_108_436_0,
    i_10_108_519_0, i_10_108_799_0, i_10_108_963_0, i_10_108_1036_0,
    i_10_108_1120_0, i_10_108_1234_0, i_10_108_1306_0, i_10_108_1308_0,
    i_10_108_1363_0, i_10_108_1365_0, i_10_108_1431_0, i_10_108_1447_0,
    i_10_108_1554_0, i_10_108_1612_0, i_10_108_1653_0, i_10_108_1654_0,
    i_10_108_1655_0, i_10_108_1687_0, i_10_108_1690_0, i_10_108_1820_0,
    i_10_108_1821_0, i_10_108_1944_0, i_10_108_1945_0, i_10_108_1950_0,
    i_10_108_1953_0, i_10_108_2199_0, i_10_108_2200_0, i_10_108_2204_0,
    i_10_108_2307_0, i_10_108_2361_0, i_10_108_2407_0, i_10_108_2470_0,
    i_10_108_2514_0, i_10_108_2607_0, i_10_108_2630_0, i_10_108_2636_0,
    i_10_108_2660_0, i_10_108_2679_0, i_10_108_2701_0, i_10_108_2722_0,
    i_10_108_2724_0, i_10_108_2725_0, i_10_108_2726_0, i_10_108_2727_0,
    i_10_108_2821_0, i_10_108_2874_0, i_10_108_2885_0, i_10_108_2923_0,
    i_10_108_2994_0, i_10_108_3036_0, i_10_108_3072_0, i_10_108_3073_0,
    i_10_108_3090_0, i_10_108_3195_0, i_10_108_3198_0, i_10_108_3203_0,
    i_10_108_3278_0, i_10_108_3282_0, i_10_108_3298_0, i_10_108_3388_0,
    i_10_108_3429_0, i_10_108_3430_0, i_10_108_3436_0, i_10_108_3467_0,
    i_10_108_3468_0, i_10_108_3471_0, i_10_108_3472_0, i_10_108_3498_0,
    i_10_108_3522_0, i_10_108_3612_0, i_10_108_3621_0, i_10_108_3646_0,
    i_10_108_3648_0, i_10_108_3649_0, i_10_108_3651_0, i_10_108_3723_0,
    i_10_108_3726_0, i_10_108_3783_0, i_10_108_3834_0, i_10_108_3853_0,
    i_10_108_3855_0, i_10_108_3859_0, i_10_108_3860_0, i_10_108_3909_0,
    i_10_108_3983_0, i_10_108_4171_0, i_10_108_4174_0, i_10_108_4213_0,
    i_10_108_4216_0, i_10_108_4273_0, i_10_108_4277_0, i_10_108_4291_0,
    o_10_108_0_0  );
  input  i_10_108_123_0, i_10_108_153_0, i_10_108_171_0, i_10_108_175_0,
    i_10_108_244_0, i_10_108_248_0, i_10_108_434_0, i_10_108_436_0,
    i_10_108_519_0, i_10_108_799_0, i_10_108_963_0, i_10_108_1036_0,
    i_10_108_1120_0, i_10_108_1234_0, i_10_108_1306_0, i_10_108_1308_0,
    i_10_108_1363_0, i_10_108_1365_0, i_10_108_1431_0, i_10_108_1447_0,
    i_10_108_1554_0, i_10_108_1612_0, i_10_108_1653_0, i_10_108_1654_0,
    i_10_108_1655_0, i_10_108_1687_0, i_10_108_1690_0, i_10_108_1820_0,
    i_10_108_1821_0, i_10_108_1944_0, i_10_108_1945_0, i_10_108_1950_0,
    i_10_108_1953_0, i_10_108_2199_0, i_10_108_2200_0, i_10_108_2204_0,
    i_10_108_2307_0, i_10_108_2361_0, i_10_108_2407_0, i_10_108_2470_0,
    i_10_108_2514_0, i_10_108_2607_0, i_10_108_2630_0, i_10_108_2636_0,
    i_10_108_2660_0, i_10_108_2679_0, i_10_108_2701_0, i_10_108_2722_0,
    i_10_108_2724_0, i_10_108_2725_0, i_10_108_2726_0, i_10_108_2727_0,
    i_10_108_2821_0, i_10_108_2874_0, i_10_108_2885_0, i_10_108_2923_0,
    i_10_108_2994_0, i_10_108_3036_0, i_10_108_3072_0, i_10_108_3073_0,
    i_10_108_3090_0, i_10_108_3195_0, i_10_108_3198_0, i_10_108_3203_0,
    i_10_108_3278_0, i_10_108_3282_0, i_10_108_3298_0, i_10_108_3388_0,
    i_10_108_3429_0, i_10_108_3430_0, i_10_108_3436_0, i_10_108_3467_0,
    i_10_108_3468_0, i_10_108_3471_0, i_10_108_3472_0, i_10_108_3498_0,
    i_10_108_3522_0, i_10_108_3612_0, i_10_108_3621_0, i_10_108_3646_0,
    i_10_108_3648_0, i_10_108_3649_0, i_10_108_3651_0, i_10_108_3723_0,
    i_10_108_3726_0, i_10_108_3783_0, i_10_108_3834_0, i_10_108_3853_0,
    i_10_108_3855_0, i_10_108_3859_0, i_10_108_3860_0, i_10_108_3909_0,
    i_10_108_3983_0, i_10_108_4171_0, i_10_108_4174_0, i_10_108_4213_0,
    i_10_108_4216_0, i_10_108_4273_0, i_10_108_4277_0, i_10_108_4291_0;
  output o_10_108_0_0;
  assign o_10_108_0_0 = 0;
endmodule



// Benchmark "kernel_10_109" written by ABC on Sun Jul 19 10:22:52 2020

module kernel_10_109 ( 
    i_10_109_39_0, i_10_109_63_0, i_10_109_64_0, i_10_109_172_0,
    i_10_109_316_0, i_10_109_405_0, i_10_109_408_0, i_10_109_409_0,
    i_10_109_432_0, i_10_109_433_0, i_10_109_436_0, i_10_109_659_0,
    i_10_109_712_0, i_10_109_796_0, i_10_109_797_0, i_10_109_990_0,
    i_10_109_991_0, i_10_109_993_0, i_10_109_1026_0, i_10_109_1154_0,
    i_10_109_1234_0, i_10_109_1238_0, i_10_109_1306_0, i_10_109_1359_0,
    i_10_109_1360_0, i_10_109_1362_0, i_10_109_1433_0, i_10_109_1442_0,
    i_10_109_1539_0, i_10_109_1541_0, i_10_109_1542_0, i_10_109_1544_0,
    i_10_109_1621_0, i_10_109_1622_0, i_10_109_1683_0, i_10_109_1685_0,
    i_10_109_1687_0, i_10_109_1688_0, i_10_109_1711_0, i_10_109_1992_0,
    i_10_109_2016_0, i_10_109_2017_0, i_10_109_2179_0, i_10_109_2197_0,
    i_10_109_2352_0, i_10_109_2359_0, i_10_109_2362_0, i_10_109_2363_0,
    i_10_109_2512_0, i_10_109_2566_0, i_10_109_2628_0, i_10_109_2659_0,
    i_10_109_2718_0, i_10_109_2730_0, i_10_109_2781_0, i_10_109_2829_0,
    i_10_109_2837_0, i_10_109_2872_0, i_10_109_3042_0, i_10_109_3044_0,
    i_10_109_3069_0, i_10_109_3070_0, i_10_109_3071_0, i_10_109_3073_0,
    i_10_109_3074_0, i_10_109_3195_0, i_10_109_3268_0, i_10_109_3331_0,
    i_10_109_3332_0, i_10_109_3384_0, i_10_109_3538_0, i_10_109_3541_0,
    i_10_109_3612_0, i_10_109_3785_0, i_10_109_3807_0, i_10_109_3808_0,
    i_10_109_3838_0, i_10_109_3839_0, i_10_109_3850_0, i_10_109_3853_0,
    i_10_109_3855_0, i_10_109_3857_0, i_10_109_3880_0, i_10_109_3980_0,
    i_10_109_3991_0, i_10_109_4113_0, i_10_109_4114_0, i_10_109_4115_0,
    i_10_109_4116_0, i_10_109_4122_0, i_10_109_4172_0, i_10_109_4175_0,
    i_10_109_4230_0, i_10_109_4275_0, i_10_109_4285_0, i_10_109_4292_0,
    i_10_109_4437_0, i_10_109_4567_0, i_10_109_4568_0, i_10_109_4569_0,
    o_10_109_0_0  );
  input  i_10_109_39_0, i_10_109_63_0, i_10_109_64_0, i_10_109_172_0,
    i_10_109_316_0, i_10_109_405_0, i_10_109_408_0, i_10_109_409_0,
    i_10_109_432_0, i_10_109_433_0, i_10_109_436_0, i_10_109_659_0,
    i_10_109_712_0, i_10_109_796_0, i_10_109_797_0, i_10_109_990_0,
    i_10_109_991_0, i_10_109_993_0, i_10_109_1026_0, i_10_109_1154_0,
    i_10_109_1234_0, i_10_109_1238_0, i_10_109_1306_0, i_10_109_1359_0,
    i_10_109_1360_0, i_10_109_1362_0, i_10_109_1433_0, i_10_109_1442_0,
    i_10_109_1539_0, i_10_109_1541_0, i_10_109_1542_0, i_10_109_1544_0,
    i_10_109_1621_0, i_10_109_1622_0, i_10_109_1683_0, i_10_109_1685_0,
    i_10_109_1687_0, i_10_109_1688_0, i_10_109_1711_0, i_10_109_1992_0,
    i_10_109_2016_0, i_10_109_2017_0, i_10_109_2179_0, i_10_109_2197_0,
    i_10_109_2352_0, i_10_109_2359_0, i_10_109_2362_0, i_10_109_2363_0,
    i_10_109_2512_0, i_10_109_2566_0, i_10_109_2628_0, i_10_109_2659_0,
    i_10_109_2718_0, i_10_109_2730_0, i_10_109_2781_0, i_10_109_2829_0,
    i_10_109_2837_0, i_10_109_2872_0, i_10_109_3042_0, i_10_109_3044_0,
    i_10_109_3069_0, i_10_109_3070_0, i_10_109_3071_0, i_10_109_3073_0,
    i_10_109_3074_0, i_10_109_3195_0, i_10_109_3268_0, i_10_109_3331_0,
    i_10_109_3332_0, i_10_109_3384_0, i_10_109_3538_0, i_10_109_3541_0,
    i_10_109_3612_0, i_10_109_3785_0, i_10_109_3807_0, i_10_109_3808_0,
    i_10_109_3838_0, i_10_109_3839_0, i_10_109_3850_0, i_10_109_3853_0,
    i_10_109_3855_0, i_10_109_3857_0, i_10_109_3880_0, i_10_109_3980_0,
    i_10_109_3991_0, i_10_109_4113_0, i_10_109_4114_0, i_10_109_4115_0,
    i_10_109_4116_0, i_10_109_4122_0, i_10_109_4172_0, i_10_109_4175_0,
    i_10_109_4230_0, i_10_109_4275_0, i_10_109_4285_0, i_10_109_4292_0,
    i_10_109_4437_0, i_10_109_4567_0, i_10_109_4568_0, i_10_109_4569_0;
  output o_10_109_0_0;
  assign o_10_109_0_0 = 0;
endmodule



// Benchmark "kernel_10_110" written by ABC on Sun Jul 19 10:22:53 2020

module kernel_10_110 ( 
    i_10_110_31_0, i_10_110_37_0, i_10_110_178_0, i_10_110_218_0,
    i_10_110_220_0, i_10_110_224_0, i_10_110_319_0, i_10_110_406_0,
    i_10_110_407_0, i_10_110_448_0, i_10_110_514_0, i_10_110_602_0,
    i_10_110_711_0, i_10_110_713_0, i_10_110_714_0, i_10_110_732_0,
    i_10_110_794_0, i_10_110_797_0, i_10_110_800_0, i_10_110_828_0,
    i_10_110_830_0, i_10_110_963_0, i_10_110_1239_0, i_10_110_1363_0,
    i_10_110_1454_0, i_10_110_1579_0, i_10_110_1647_0, i_10_110_1649_0,
    i_10_110_1683_0, i_10_110_1684_0, i_10_110_1685_0, i_10_110_1687_0,
    i_10_110_1688_0, i_10_110_1691_0, i_10_110_1719_0, i_10_110_1765_0,
    i_10_110_1766_0, i_10_110_1801_0, i_10_110_1802_0, i_10_110_1805_0,
    i_10_110_1821_0, i_10_110_1915_0, i_10_110_1939_0, i_10_110_2096_0,
    i_10_110_2307_0, i_10_110_2308_0, i_10_110_2448_0, i_10_110_2449_0,
    i_10_110_2450_0, i_10_110_2468_0, i_10_110_2539_0, i_10_110_2542_0,
    i_10_110_2659_0, i_10_110_2723_0, i_10_110_2725_0, i_10_110_2726_0,
    i_10_110_2728_0, i_10_110_2734_0, i_10_110_2781_0, i_10_110_2782_0,
    i_10_110_2784_0, i_10_110_2788_0, i_10_110_2820_0, i_10_110_2832_0,
    i_10_110_2985_0, i_10_110_3199_0, i_10_110_3270_0, i_10_110_3279_0,
    i_10_110_3280_0, i_10_110_3281_0, i_10_110_3283_0, i_10_110_3291_0,
    i_10_110_3325_0, i_10_110_3384_0, i_10_110_3390_0, i_10_110_3406_0,
    i_10_110_3409_0, i_10_110_3430_0, i_10_110_3494_0, i_10_110_3523_0,
    i_10_110_3539_0, i_10_110_3616_0, i_10_110_3649_0, i_10_110_3725_0,
    i_10_110_3727_0, i_10_110_3781_0, i_10_110_3852_0, i_10_110_3854_0,
    i_10_110_3857_0, i_10_110_3858_0, i_10_110_3906_0, i_10_110_3982_0,
    i_10_110_4054_0, i_10_110_4121_0, i_10_110_4238_0, i_10_110_4268_0,
    i_10_110_4285_0, i_10_110_4286_0, i_10_110_4289_0, i_10_110_4477_0,
    o_10_110_0_0  );
  input  i_10_110_31_0, i_10_110_37_0, i_10_110_178_0, i_10_110_218_0,
    i_10_110_220_0, i_10_110_224_0, i_10_110_319_0, i_10_110_406_0,
    i_10_110_407_0, i_10_110_448_0, i_10_110_514_0, i_10_110_602_0,
    i_10_110_711_0, i_10_110_713_0, i_10_110_714_0, i_10_110_732_0,
    i_10_110_794_0, i_10_110_797_0, i_10_110_800_0, i_10_110_828_0,
    i_10_110_830_0, i_10_110_963_0, i_10_110_1239_0, i_10_110_1363_0,
    i_10_110_1454_0, i_10_110_1579_0, i_10_110_1647_0, i_10_110_1649_0,
    i_10_110_1683_0, i_10_110_1684_0, i_10_110_1685_0, i_10_110_1687_0,
    i_10_110_1688_0, i_10_110_1691_0, i_10_110_1719_0, i_10_110_1765_0,
    i_10_110_1766_0, i_10_110_1801_0, i_10_110_1802_0, i_10_110_1805_0,
    i_10_110_1821_0, i_10_110_1915_0, i_10_110_1939_0, i_10_110_2096_0,
    i_10_110_2307_0, i_10_110_2308_0, i_10_110_2448_0, i_10_110_2449_0,
    i_10_110_2450_0, i_10_110_2468_0, i_10_110_2539_0, i_10_110_2542_0,
    i_10_110_2659_0, i_10_110_2723_0, i_10_110_2725_0, i_10_110_2726_0,
    i_10_110_2728_0, i_10_110_2734_0, i_10_110_2781_0, i_10_110_2782_0,
    i_10_110_2784_0, i_10_110_2788_0, i_10_110_2820_0, i_10_110_2832_0,
    i_10_110_2985_0, i_10_110_3199_0, i_10_110_3270_0, i_10_110_3279_0,
    i_10_110_3280_0, i_10_110_3281_0, i_10_110_3283_0, i_10_110_3291_0,
    i_10_110_3325_0, i_10_110_3384_0, i_10_110_3390_0, i_10_110_3406_0,
    i_10_110_3409_0, i_10_110_3430_0, i_10_110_3494_0, i_10_110_3523_0,
    i_10_110_3539_0, i_10_110_3616_0, i_10_110_3649_0, i_10_110_3725_0,
    i_10_110_3727_0, i_10_110_3781_0, i_10_110_3852_0, i_10_110_3854_0,
    i_10_110_3857_0, i_10_110_3858_0, i_10_110_3906_0, i_10_110_3982_0,
    i_10_110_4054_0, i_10_110_4121_0, i_10_110_4238_0, i_10_110_4268_0,
    i_10_110_4285_0, i_10_110_4286_0, i_10_110_4289_0, i_10_110_4477_0;
  output o_10_110_0_0;
  assign o_10_110_0_0 = 0;
endmodule



// Benchmark "kernel_10_111" written by ABC on Sun Jul 19 10:22:53 2020

module kernel_10_111 ( 
    i_10_111_171_0, i_10_111_174_0, i_10_111_175_0, i_10_111_177_0,
    i_10_111_178_0, i_10_111_179_0, i_10_111_248_0, i_10_111_281_0,
    i_10_111_284_0, i_10_111_293_0, i_10_111_315_0, i_10_111_316_0,
    i_10_111_318_0, i_10_111_319_0, i_10_111_409_0, i_10_111_411_0,
    i_10_111_412_0, i_10_111_459_0, i_10_111_466_0, i_10_111_797_0,
    i_10_111_799_0, i_10_111_957_0, i_10_111_994_0, i_10_111_1087_0,
    i_10_111_1156_0, i_10_111_1237_0, i_10_111_1238_0, i_10_111_1240_0,
    i_10_111_1250_0, i_10_111_1268_0, i_10_111_1313_0, i_10_111_1344_0,
    i_10_111_1347_0, i_10_111_1348_0, i_10_111_1442_0, i_10_111_1445_0,
    i_10_111_1577_0, i_10_111_1580_0, i_10_111_1685_0, i_10_111_1686_0,
    i_10_111_1714_0, i_10_111_1821_0, i_10_111_1825_0, i_10_111_1872_0,
    i_10_111_1874_0, i_10_111_1995_0, i_10_111_2198_0, i_10_111_2334_0,
    i_10_111_2358_0, i_10_111_2365_0, i_10_111_2472_0, i_10_111_2517_0,
    i_10_111_2518_0, i_10_111_2519_0, i_10_111_2605_0, i_10_111_2629_0,
    i_10_111_2631_0, i_10_111_2632_0, i_10_111_2634_0, i_10_111_2635_0,
    i_10_111_2636_0, i_10_111_2674_0, i_10_111_2700_0, i_10_111_2704_0,
    i_10_111_2710_0, i_10_111_2711_0, i_10_111_2723_0, i_10_111_2724_0,
    i_10_111_2781_0, i_10_111_2782_0, i_10_111_2785_0, i_10_111_2832_0,
    i_10_111_3072_0, i_10_111_3073_0, i_10_111_3201_0, i_10_111_3279_0,
    i_10_111_3319_0, i_10_111_3385_0, i_10_111_3431_0, i_10_111_3497_0,
    i_10_111_3543_0, i_10_111_3562_0, i_10_111_3586_0, i_10_111_3611_0,
    i_10_111_3617_0, i_10_111_3841_0, i_10_111_3893_0, i_10_111_3942_0,
    i_10_111_3943_0, i_10_111_4116_0, i_10_111_4117_0, i_10_111_4118_0,
    i_10_111_4120_0, i_10_111_4121_0, i_10_111_4128_0, i_10_111_4129_0,
    i_10_111_4130_0, i_10_111_4173_0, i_10_111_4281_0, i_10_111_4291_0,
    o_10_111_0_0  );
  input  i_10_111_171_0, i_10_111_174_0, i_10_111_175_0, i_10_111_177_0,
    i_10_111_178_0, i_10_111_179_0, i_10_111_248_0, i_10_111_281_0,
    i_10_111_284_0, i_10_111_293_0, i_10_111_315_0, i_10_111_316_0,
    i_10_111_318_0, i_10_111_319_0, i_10_111_409_0, i_10_111_411_0,
    i_10_111_412_0, i_10_111_459_0, i_10_111_466_0, i_10_111_797_0,
    i_10_111_799_0, i_10_111_957_0, i_10_111_994_0, i_10_111_1087_0,
    i_10_111_1156_0, i_10_111_1237_0, i_10_111_1238_0, i_10_111_1240_0,
    i_10_111_1250_0, i_10_111_1268_0, i_10_111_1313_0, i_10_111_1344_0,
    i_10_111_1347_0, i_10_111_1348_0, i_10_111_1442_0, i_10_111_1445_0,
    i_10_111_1577_0, i_10_111_1580_0, i_10_111_1685_0, i_10_111_1686_0,
    i_10_111_1714_0, i_10_111_1821_0, i_10_111_1825_0, i_10_111_1872_0,
    i_10_111_1874_0, i_10_111_1995_0, i_10_111_2198_0, i_10_111_2334_0,
    i_10_111_2358_0, i_10_111_2365_0, i_10_111_2472_0, i_10_111_2517_0,
    i_10_111_2518_0, i_10_111_2519_0, i_10_111_2605_0, i_10_111_2629_0,
    i_10_111_2631_0, i_10_111_2632_0, i_10_111_2634_0, i_10_111_2635_0,
    i_10_111_2636_0, i_10_111_2674_0, i_10_111_2700_0, i_10_111_2704_0,
    i_10_111_2710_0, i_10_111_2711_0, i_10_111_2723_0, i_10_111_2724_0,
    i_10_111_2781_0, i_10_111_2782_0, i_10_111_2785_0, i_10_111_2832_0,
    i_10_111_3072_0, i_10_111_3073_0, i_10_111_3201_0, i_10_111_3279_0,
    i_10_111_3319_0, i_10_111_3385_0, i_10_111_3431_0, i_10_111_3497_0,
    i_10_111_3543_0, i_10_111_3562_0, i_10_111_3586_0, i_10_111_3611_0,
    i_10_111_3617_0, i_10_111_3841_0, i_10_111_3893_0, i_10_111_3942_0,
    i_10_111_3943_0, i_10_111_4116_0, i_10_111_4117_0, i_10_111_4118_0,
    i_10_111_4120_0, i_10_111_4121_0, i_10_111_4128_0, i_10_111_4129_0,
    i_10_111_4130_0, i_10_111_4173_0, i_10_111_4281_0, i_10_111_4291_0;
  output o_10_111_0_0;
  assign o_10_111_0_0 = 0;
endmodule



// Benchmark "kernel_10_112" written by ABC on Sun Jul 19 10:22:54 2020

module kernel_10_112 ( 
    i_10_112_41_0, i_10_112_64_0, i_10_112_216_0, i_10_112_317_0,
    i_10_112_431_0, i_10_112_433_0, i_10_112_437_0, i_10_112_442_0,
    i_10_112_443_0, i_10_112_538_0, i_10_112_895_0, i_10_112_992_0,
    i_10_112_1034_0, i_10_112_1119_0, i_10_112_1239_0, i_10_112_1308_0,
    i_10_112_1309_0, i_10_112_1311_0, i_10_112_1378_0, i_10_112_1456_0,
    i_10_112_1653_0, i_10_112_1655_0, i_10_112_1676_0, i_10_112_1683_0,
    i_10_112_1684_0, i_10_112_1690_0, i_10_112_1809_0, i_10_112_1822_0,
    i_10_112_1824_0, i_10_112_1950_0, i_10_112_2110_0, i_10_112_2202_0,
    i_10_112_2261_0, i_10_112_2359_0, i_10_112_2361_0, i_10_112_2461_0,
    i_10_112_2467_0, i_10_112_2572_0, i_10_112_2641_0, i_10_112_2658_0,
    i_10_112_2659_0, i_10_112_2710_0, i_10_112_2726_0, i_10_112_2727_0,
    i_10_112_2733_0, i_10_112_2826_0, i_10_112_2827_0, i_10_112_2829_0,
    i_10_112_2830_0, i_10_112_2831_0, i_10_112_2835_0, i_10_112_2852_0,
    i_10_112_2920_0, i_10_112_2982_0, i_10_112_2993_0, i_10_112_3042_0,
    i_10_112_3048_0, i_10_112_3073_0, i_10_112_3093_0, i_10_112_3197_0,
    i_10_112_3198_0, i_10_112_3199_0, i_10_112_3200_0, i_10_112_3271_0,
    i_10_112_3454_0, i_10_112_3541_0, i_10_112_3561_0, i_10_112_3609_0,
    i_10_112_3612_0, i_10_112_3703_0, i_10_112_3775_0, i_10_112_3838_0,
    i_10_112_3839_0, i_10_112_3854_0, i_10_112_3855_0, i_10_112_3856_0,
    i_10_112_3859_0, i_10_112_3860_0, i_10_112_3990_0, i_10_112_3991_0,
    i_10_112_4029_0, i_10_112_4030_0, i_10_112_4031_0, i_10_112_4116_0,
    i_10_112_4117_0, i_10_112_4119_0, i_10_112_4120_0, i_10_112_4129_0,
    i_10_112_4159_0, i_10_112_4171_0, i_10_112_4172_0, i_10_112_4173_0,
    i_10_112_4174_0, i_10_112_4232_0, i_10_112_4279_0, i_10_112_4290_0,
    i_10_112_4439_0, i_10_112_4529_0, i_10_112_4564_0, i_10_112_4597_0,
    o_10_112_0_0  );
  input  i_10_112_41_0, i_10_112_64_0, i_10_112_216_0, i_10_112_317_0,
    i_10_112_431_0, i_10_112_433_0, i_10_112_437_0, i_10_112_442_0,
    i_10_112_443_0, i_10_112_538_0, i_10_112_895_0, i_10_112_992_0,
    i_10_112_1034_0, i_10_112_1119_0, i_10_112_1239_0, i_10_112_1308_0,
    i_10_112_1309_0, i_10_112_1311_0, i_10_112_1378_0, i_10_112_1456_0,
    i_10_112_1653_0, i_10_112_1655_0, i_10_112_1676_0, i_10_112_1683_0,
    i_10_112_1684_0, i_10_112_1690_0, i_10_112_1809_0, i_10_112_1822_0,
    i_10_112_1824_0, i_10_112_1950_0, i_10_112_2110_0, i_10_112_2202_0,
    i_10_112_2261_0, i_10_112_2359_0, i_10_112_2361_0, i_10_112_2461_0,
    i_10_112_2467_0, i_10_112_2572_0, i_10_112_2641_0, i_10_112_2658_0,
    i_10_112_2659_0, i_10_112_2710_0, i_10_112_2726_0, i_10_112_2727_0,
    i_10_112_2733_0, i_10_112_2826_0, i_10_112_2827_0, i_10_112_2829_0,
    i_10_112_2830_0, i_10_112_2831_0, i_10_112_2835_0, i_10_112_2852_0,
    i_10_112_2920_0, i_10_112_2982_0, i_10_112_2993_0, i_10_112_3042_0,
    i_10_112_3048_0, i_10_112_3073_0, i_10_112_3093_0, i_10_112_3197_0,
    i_10_112_3198_0, i_10_112_3199_0, i_10_112_3200_0, i_10_112_3271_0,
    i_10_112_3454_0, i_10_112_3541_0, i_10_112_3561_0, i_10_112_3609_0,
    i_10_112_3612_0, i_10_112_3703_0, i_10_112_3775_0, i_10_112_3838_0,
    i_10_112_3839_0, i_10_112_3854_0, i_10_112_3855_0, i_10_112_3856_0,
    i_10_112_3859_0, i_10_112_3860_0, i_10_112_3990_0, i_10_112_3991_0,
    i_10_112_4029_0, i_10_112_4030_0, i_10_112_4031_0, i_10_112_4116_0,
    i_10_112_4117_0, i_10_112_4119_0, i_10_112_4120_0, i_10_112_4129_0,
    i_10_112_4159_0, i_10_112_4171_0, i_10_112_4172_0, i_10_112_4173_0,
    i_10_112_4174_0, i_10_112_4232_0, i_10_112_4279_0, i_10_112_4290_0,
    i_10_112_4439_0, i_10_112_4529_0, i_10_112_4564_0, i_10_112_4597_0;
  output o_10_112_0_0;
  assign o_10_112_0_0 = 0;
endmodule



// Benchmark "kernel_10_113" written by ABC on Sun Jul 19 10:22:56 2020

module kernel_10_113 ( 
    i_10_113_35_0, i_10_113_124_0, i_10_113_178_0, i_10_113_249_0,
    i_10_113_282_0, i_10_113_283_0, i_10_113_284_0, i_10_113_286_0,
    i_10_113_319_0, i_10_113_322_0, i_10_113_324_0, i_10_113_408_0,
    i_10_113_409_0, i_10_113_430_0, i_10_113_437_0, i_10_113_444_0,
    i_10_113_445_0, i_10_113_446_0, i_10_113_460_0, i_10_113_967_0,
    i_10_113_993_0, i_10_113_1000_0, i_10_113_1002_0, i_10_113_1005_0,
    i_10_113_1006_0, i_10_113_1233_0, i_10_113_1237_0, i_10_113_1247_0,
    i_10_113_1249_0, i_10_113_1310_0, i_10_113_1576_0, i_10_113_1582_0,
    i_10_113_1617_0, i_10_113_1650_0, i_10_113_1818_0, i_10_113_1819_0,
    i_10_113_1821_0, i_10_113_1822_0, i_10_113_1823_0, i_10_113_1912_0,
    i_10_113_1913_0, i_10_113_1950_0, i_10_113_1951_0, i_10_113_2179_0,
    i_10_113_2180_0, i_10_113_2184_0, i_10_113_2334_0, i_10_113_2338_0,
    i_10_113_2349_0, i_10_113_2381_0, i_10_113_2382_0, i_10_113_2383_0,
    i_10_113_2407_0, i_10_113_2409_0, i_10_113_2410_0, i_10_113_2449_0,
    i_10_113_2454_0, i_10_113_2629_0, i_10_113_2635_0, i_10_113_2636_0,
    i_10_113_2655_0, i_10_113_2679_0, i_10_113_2706_0, i_10_113_2710_0,
    i_10_113_2716_0, i_10_113_2728_0, i_10_113_2730_0, i_10_113_2829_0,
    i_10_113_2917_0, i_10_113_3039_0, i_10_113_3049_0, i_10_113_3094_0,
    i_10_113_3095_0, i_10_113_3153_0, i_10_113_3154_0, i_10_113_3155_0,
    i_10_113_3198_0, i_10_113_3200_0, i_10_113_3237_0, i_10_113_3269_0,
    i_10_113_3270_0, i_10_113_3280_0, i_10_113_3388_0, i_10_113_3389_0,
    i_10_113_3390_0, i_10_113_3404_0, i_10_113_3405_0, i_10_113_3526_0,
    i_10_113_3582_0, i_10_113_3613_0, i_10_113_3616_0, i_10_113_3783_0,
    i_10_113_3837_0, i_10_113_3838_0, i_10_113_3839_0, i_10_113_3847_0,
    i_10_113_3853_0, i_10_113_3856_0, i_10_113_4120_0, i_10_113_4268_0,
    o_10_113_0_0  );
  input  i_10_113_35_0, i_10_113_124_0, i_10_113_178_0, i_10_113_249_0,
    i_10_113_282_0, i_10_113_283_0, i_10_113_284_0, i_10_113_286_0,
    i_10_113_319_0, i_10_113_322_0, i_10_113_324_0, i_10_113_408_0,
    i_10_113_409_0, i_10_113_430_0, i_10_113_437_0, i_10_113_444_0,
    i_10_113_445_0, i_10_113_446_0, i_10_113_460_0, i_10_113_967_0,
    i_10_113_993_0, i_10_113_1000_0, i_10_113_1002_0, i_10_113_1005_0,
    i_10_113_1006_0, i_10_113_1233_0, i_10_113_1237_0, i_10_113_1247_0,
    i_10_113_1249_0, i_10_113_1310_0, i_10_113_1576_0, i_10_113_1582_0,
    i_10_113_1617_0, i_10_113_1650_0, i_10_113_1818_0, i_10_113_1819_0,
    i_10_113_1821_0, i_10_113_1822_0, i_10_113_1823_0, i_10_113_1912_0,
    i_10_113_1913_0, i_10_113_1950_0, i_10_113_1951_0, i_10_113_2179_0,
    i_10_113_2180_0, i_10_113_2184_0, i_10_113_2334_0, i_10_113_2338_0,
    i_10_113_2349_0, i_10_113_2381_0, i_10_113_2382_0, i_10_113_2383_0,
    i_10_113_2407_0, i_10_113_2409_0, i_10_113_2410_0, i_10_113_2449_0,
    i_10_113_2454_0, i_10_113_2629_0, i_10_113_2635_0, i_10_113_2636_0,
    i_10_113_2655_0, i_10_113_2679_0, i_10_113_2706_0, i_10_113_2710_0,
    i_10_113_2716_0, i_10_113_2728_0, i_10_113_2730_0, i_10_113_2829_0,
    i_10_113_2917_0, i_10_113_3039_0, i_10_113_3049_0, i_10_113_3094_0,
    i_10_113_3095_0, i_10_113_3153_0, i_10_113_3154_0, i_10_113_3155_0,
    i_10_113_3198_0, i_10_113_3200_0, i_10_113_3237_0, i_10_113_3269_0,
    i_10_113_3270_0, i_10_113_3280_0, i_10_113_3388_0, i_10_113_3389_0,
    i_10_113_3390_0, i_10_113_3404_0, i_10_113_3405_0, i_10_113_3526_0,
    i_10_113_3582_0, i_10_113_3613_0, i_10_113_3616_0, i_10_113_3783_0,
    i_10_113_3837_0, i_10_113_3838_0, i_10_113_3839_0, i_10_113_3847_0,
    i_10_113_3853_0, i_10_113_3856_0, i_10_113_4120_0, i_10_113_4268_0;
  output o_10_113_0_0;
  assign o_10_113_0_0 = ~((~i_10_113_35_0 & ((~i_10_113_1002_0 & i_10_113_1819_0 & ~i_10_113_2179_0 & ~i_10_113_2338_0 & ~i_10_113_2349_0) | (~i_10_113_1006_0 & ~i_10_113_1617_0 & ~i_10_113_2180_0 & ~i_10_113_2381_0 & ~i_10_113_2383_0 & ~i_10_113_3198_0 & ~i_10_113_3270_0))) | (~i_10_113_3405_0 & ((~i_10_113_124_0 & ~i_10_113_1576_0 & ~i_10_113_2407_0 & ((~i_10_113_2184_0 & ~i_10_113_2381_0 & ~i_10_113_2383_0 & ~i_10_113_2409_0 & ~i_10_113_2706_0 & ~i_10_113_3200_0) | (~i_10_113_1582_0 & ~i_10_113_1950_0 & ~i_10_113_2179_0 & ~i_10_113_2382_0 & ~i_10_113_2829_0 & ~i_10_113_2917_0 & ~i_10_113_3095_0 & ~i_10_113_3616_0))) | (~i_10_113_2184_0 & ((~i_10_113_324_0 & i_10_113_460_0 & ~i_10_113_2381_0 & ~i_10_113_2706_0 & ~i_10_113_2917_0 & ~i_10_113_3095_0 & ~i_10_113_3200_0) | (i_10_113_1237_0 & ~i_10_113_2635_0 & ~i_10_113_2636_0 & ~i_10_113_2679_0 & ~i_10_113_3269_0))))) | (~i_10_113_445_0 & ((~i_10_113_1576_0 & ~i_10_113_1950_0 & ~i_10_113_2179_0 & ~i_10_113_2410_0 & ~i_10_113_3200_0) | (~i_10_113_1247_0 & ~i_10_113_1617_0 & ~i_10_113_1823_0 & ~i_10_113_2636_0 & ~i_10_113_2829_0 & ~i_10_113_3390_0 & i_10_113_3616_0))) | (~i_10_113_446_0 & ((~i_10_113_444_0 & ~i_10_113_1822_0 & ~i_10_113_1823_0 & ~i_10_113_1950_0 & ~i_10_113_1951_0 & ~i_10_113_2179_0) | (i_10_113_460_0 & ~i_10_113_1006_0 & ~i_10_113_1821_0 & ~i_10_113_2349_0))) | (~i_10_113_444_0 & ~i_10_113_3856_0 & ((~i_10_113_1822_0 & i_10_113_2180_0 & ~i_10_113_2410_0) | (~i_10_113_1006_0 & i_10_113_2636_0 & ~i_10_113_3095_0 & ~i_10_113_4268_0))) | (~i_10_113_3783_0 & ((~i_10_113_1006_0 & ((i_10_113_445_0 & ~i_10_113_460_0 & ~i_10_113_1000_0 & ~i_10_113_1650_0 & ~i_10_113_2409_0 & ~i_10_113_2679_0 & ~i_10_113_3095_0) | (i_10_113_460_0 & ~i_10_113_967_0 & ~i_10_113_2184_0 & ~i_10_113_2338_0 & ~i_10_113_2716_0 & ~i_10_113_3269_0))) | (i_10_113_409_0 & ~i_10_113_2409_0) | (~i_10_113_1951_0 & ~i_10_113_2179_0 & ~i_10_113_1582_0 & ~i_10_113_1650_0 & ~i_10_113_2180_0 & ~i_10_113_2410_0 & ~i_10_113_3094_0 & ~i_10_113_3237_0))) | (i_10_113_460_0 & ((~i_10_113_2635_0 & i_10_113_2728_0 & ~i_10_113_3838_0) | (~i_10_113_1000_0 & ~i_10_113_2180_0 & ~i_10_113_3039_0 & i_10_113_3613_0 & i_10_113_3853_0))) | (~i_10_113_3839_0 & ((~i_10_113_1310_0 & ~i_10_113_2179_0 & ~i_10_113_2410_0 & i_10_113_2635_0 & ~i_10_113_3389_0 & ~i_10_113_3613_0 & ~i_10_113_3838_0) | (~i_10_113_324_0 & ~i_10_113_1000_0 & ~i_10_113_2635_0 & ~i_10_113_3270_0 & ~i_10_113_3847_0 & i_10_113_3853_0))) | (i_10_113_286_0 & i_10_113_1249_0 & ~i_10_113_1951_0) | (i_10_113_283_0 & ~i_10_113_1950_0 & ~i_10_113_2180_0 & ~i_10_113_2338_0 & ~i_10_113_3095_0) | (i_10_113_3389_0 & ~i_10_113_3837_0));
endmodule



// Benchmark "kernel_10_114" written by ABC on Sun Jul 19 10:22:56 2020

module kernel_10_114 ( 
    i_10_114_27_0, i_10_114_28_0, i_10_114_30_0, i_10_114_291_0,
    i_10_114_319_0, i_10_114_435_0, i_10_114_495_0, i_10_114_712_0,
    i_10_114_720_0, i_10_114_821_0, i_10_114_895_0, i_10_114_1026_0,
    i_10_114_1234_0, i_10_114_1236_0, i_10_114_1237_0, i_10_114_1278_0,
    i_10_114_1308_0, i_10_114_1362_0, i_10_114_1432_0, i_10_114_1434_0,
    i_10_114_1435_0, i_10_114_1539_0, i_10_114_1540_0, i_10_114_1547_0,
    i_10_114_1647_0, i_10_114_1653_0, i_10_114_1683_0, i_10_114_1684_0,
    i_10_114_1765_0, i_10_114_1805_0, i_10_114_1912_0, i_10_114_1920_0,
    i_10_114_1985_0, i_10_114_2178_0, i_10_114_2179_0, i_10_114_2224_0,
    i_10_114_2308_0, i_10_114_2349_0, i_10_114_2352_0, i_10_114_2361_0,
    i_10_114_2431_0, i_10_114_2451_0, i_10_114_2529_0, i_10_114_2566_0,
    i_10_114_2610_0, i_10_114_2628_0, i_10_114_2650_0, i_10_114_2659_0,
    i_10_114_2691_0, i_10_114_2713_0, i_10_114_2718_0, i_10_114_2722_0,
    i_10_114_2736_0, i_10_114_2743_0, i_10_114_2923_0, i_10_114_2924_0,
    i_10_114_2926_0, i_10_114_2927_0, i_10_114_2934_0, i_10_114_2943_0,
    i_10_114_2944_0, i_10_114_3037_0, i_10_114_3078_0, i_10_114_3199_0,
    i_10_114_3200_0, i_10_114_3279_0, i_10_114_3391_0, i_10_114_3392_0,
    i_10_114_3406_0, i_10_114_3408_0, i_10_114_3465_0, i_10_114_3466_0,
    i_10_114_3523_0, i_10_114_3610_0, i_10_114_3612_0, i_10_114_3613_0,
    i_10_114_3614_0, i_10_114_3645_0, i_10_114_3650_0, i_10_114_3681_0,
    i_10_114_3682_0, i_10_114_3744_0, i_10_114_3781_0, i_10_114_3782_0,
    i_10_114_3783_0, i_10_114_3807_0, i_10_114_3817_0, i_10_114_3855_0,
    i_10_114_3856_0, i_10_114_3857_0, i_10_114_3888_0, i_10_114_4005_0,
    i_10_114_4006_0, i_10_114_4027_0, i_10_114_4114_0, i_10_114_4117_0,
    i_10_114_4219_0, i_10_114_4275_0, i_10_114_4276_0, i_10_114_4284_0,
    o_10_114_0_0  );
  input  i_10_114_27_0, i_10_114_28_0, i_10_114_30_0, i_10_114_291_0,
    i_10_114_319_0, i_10_114_435_0, i_10_114_495_0, i_10_114_712_0,
    i_10_114_720_0, i_10_114_821_0, i_10_114_895_0, i_10_114_1026_0,
    i_10_114_1234_0, i_10_114_1236_0, i_10_114_1237_0, i_10_114_1278_0,
    i_10_114_1308_0, i_10_114_1362_0, i_10_114_1432_0, i_10_114_1434_0,
    i_10_114_1435_0, i_10_114_1539_0, i_10_114_1540_0, i_10_114_1547_0,
    i_10_114_1647_0, i_10_114_1653_0, i_10_114_1683_0, i_10_114_1684_0,
    i_10_114_1765_0, i_10_114_1805_0, i_10_114_1912_0, i_10_114_1920_0,
    i_10_114_1985_0, i_10_114_2178_0, i_10_114_2179_0, i_10_114_2224_0,
    i_10_114_2308_0, i_10_114_2349_0, i_10_114_2352_0, i_10_114_2361_0,
    i_10_114_2431_0, i_10_114_2451_0, i_10_114_2529_0, i_10_114_2566_0,
    i_10_114_2610_0, i_10_114_2628_0, i_10_114_2650_0, i_10_114_2659_0,
    i_10_114_2691_0, i_10_114_2713_0, i_10_114_2718_0, i_10_114_2722_0,
    i_10_114_2736_0, i_10_114_2743_0, i_10_114_2923_0, i_10_114_2924_0,
    i_10_114_2926_0, i_10_114_2927_0, i_10_114_2934_0, i_10_114_2943_0,
    i_10_114_2944_0, i_10_114_3037_0, i_10_114_3078_0, i_10_114_3199_0,
    i_10_114_3200_0, i_10_114_3279_0, i_10_114_3391_0, i_10_114_3392_0,
    i_10_114_3406_0, i_10_114_3408_0, i_10_114_3465_0, i_10_114_3466_0,
    i_10_114_3523_0, i_10_114_3610_0, i_10_114_3612_0, i_10_114_3613_0,
    i_10_114_3614_0, i_10_114_3645_0, i_10_114_3650_0, i_10_114_3681_0,
    i_10_114_3682_0, i_10_114_3744_0, i_10_114_3781_0, i_10_114_3782_0,
    i_10_114_3783_0, i_10_114_3807_0, i_10_114_3817_0, i_10_114_3855_0,
    i_10_114_3856_0, i_10_114_3857_0, i_10_114_3888_0, i_10_114_4005_0,
    i_10_114_4006_0, i_10_114_4027_0, i_10_114_4114_0, i_10_114_4117_0,
    i_10_114_4219_0, i_10_114_4275_0, i_10_114_4276_0, i_10_114_4284_0;
  output o_10_114_0_0;
  assign o_10_114_0_0 = 0;
endmodule



// Benchmark "kernel_10_115" written by ABC on Sun Jul 19 10:22:57 2020

module kernel_10_115 ( 
    i_10_115_45_0, i_10_115_46_0, i_10_115_48_0, i_10_115_49_0,
    i_10_115_175_0, i_10_115_217_0, i_10_115_247_0, i_10_115_285_0,
    i_10_115_289_0, i_10_115_291_0, i_10_115_405_0, i_10_115_406_0,
    i_10_115_407_0, i_10_115_412_0, i_10_115_442_0, i_10_115_443_0,
    i_10_115_463_0, i_10_115_465_0, i_10_115_797_0, i_10_115_799_0,
    i_10_115_999_0, i_10_115_1002_0, i_10_115_1030_0, i_10_115_1035_0,
    i_10_115_1234_0, i_10_115_1238_0, i_10_115_1363_0, i_10_115_1436_0,
    i_10_115_1655_0, i_10_115_1688_0, i_10_115_1821_0, i_10_115_1909_0,
    i_10_115_1914_0, i_10_115_1915_0, i_10_115_1993_0, i_10_115_1994_0,
    i_10_115_2186_0, i_10_115_2362_0, i_10_115_2365_0, i_10_115_2449_0,
    i_10_115_2458_0, i_10_115_2460_0, i_10_115_2468_0, i_10_115_2471_0,
    i_10_115_2473_0, i_10_115_2474_0, i_10_115_2481_0, i_10_115_2546_0,
    i_10_115_2572_0, i_10_115_2608_0, i_10_115_2650_0, i_10_115_2661_0,
    i_10_115_2662_0, i_10_115_2674_0, i_10_115_2710_0, i_10_115_2711_0,
    i_10_115_2718_0, i_10_115_2720_0, i_10_115_2723_0, i_10_115_2781_0,
    i_10_115_2820_0, i_10_115_2920_0, i_10_115_2921_0, i_10_115_2924_0,
    i_10_115_3070_0, i_10_115_3195_0, i_10_115_3267_0, i_10_115_3268_0,
    i_10_115_3276_0, i_10_115_3388_0, i_10_115_3389_0, i_10_115_3390_0,
    i_10_115_3402_0, i_10_115_3406_0, i_10_115_3407_0, i_10_115_3467_0,
    i_10_115_3587_0, i_10_115_3611_0, i_10_115_3619_0, i_10_115_3688_0,
    i_10_115_3734_0, i_10_115_3842_0, i_10_115_3851_0, i_10_115_3852_0,
    i_10_115_3858_0, i_10_115_3859_0, i_10_115_3910_0, i_10_115_3929_0,
    i_10_115_3981_0, i_10_115_3982_0, i_10_115_4117_0, i_10_115_4119_0,
    i_10_115_4120_0, i_10_115_4121_0, i_10_115_4126_0, i_10_115_4129_0,
    i_10_115_4290_0, i_10_115_4291_0, i_10_115_4292_0, i_10_115_4459_0,
    o_10_115_0_0  );
  input  i_10_115_45_0, i_10_115_46_0, i_10_115_48_0, i_10_115_49_0,
    i_10_115_175_0, i_10_115_217_0, i_10_115_247_0, i_10_115_285_0,
    i_10_115_289_0, i_10_115_291_0, i_10_115_405_0, i_10_115_406_0,
    i_10_115_407_0, i_10_115_412_0, i_10_115_442_0, i_10_115_443_0,
    i_10_115_463_0, i_10_115_465_0, i_10_115_797_0, i_10_115_799_0,
    i_10_115_999_0, i_10_115_1002_0, i_10_115_1030_0, i_10_115_1035_0,
    i_10_115_1234_0, i_10_115_1238_0, i_10_115_1363_0, i_10_115_1436_0,
    i_10_115_1655_0, i_10_115_1688_0, i_10_115_1821_0, i_10_115_1909_0,
    i_10_115_1914_0, i_10_115_1915_0, i_10_115_1993_0, i_10_115_1994_0,
    i_10_115_2186_0, i_10_115_2362_0, i_10_115_2365_0, i_10_115_2449_0,
    i_10_115_2458_0, i_10_115_2460_0, i_10_115_2468_0, i_10_115_2471_0,
    i_10_115_2473_0, i_10_115_2474_0, i_10_115_2481_0, i_10_115_2546_0,
    i_10_115_2572_0, i_10_115_2608_0, i_10_115_2650_0, i_10_115_2661_0,
    i_10_115_2662_0, i_10_115_2674_0, i_10_115_2710_0, i_10_115_2711_0,
    i_10_115_2718_0, i_10_115_2720_0, i_10_115_2723_0, i_10_115_2781_0,
    i_10_115_2820_0, i_10_115_2920_0, i_10_115_2921_0, i_10_115_2924_0,
    i_10_115_3070_0, i_10_115_3195_0, i_10_115_3267_0, i_10_115_3268_0,
    i_10_115_3276_0, i_10_115_3388_0, i_10_115_3389_0, i_10_115_3390_0,
    i_10_115_3402_0, i_10_115_3406_0, i_10_115_3407_0, i_10_115_3467_0,
    i_10_115_3587_0, i_10_115_3611_0, i_10_115_3619_0, i_10_115_3688_0,
    i_10_115_3734_0, i_10_115_3842_0, i_10_115_3851_0, i_10_115_3852_0,
    i_10_115_3858_0, i_10_115_3859_0, i_10_115_3910_0, i_10_115_3929_0,
    i_10_115_3981_0, i_10_115_3982_0, i_10_115_4117_0, i_10_115_4119_0,
    i_10_115_4120_0, i_10_115_4121_0, i_10_115_4126_0, i_10_115_4129_0,
    i_10_115_4290_0, i_10_115_4291_0, i_10_115_4292_0, i_10_115_4459_0;
  output o_10_115_0_0;
  assign o_10_115_0_0 = 0;
endmodule



// Benchmark "kernel_10_116" written by ABC on Sun Jul 19 10:22:58 2020

module kernel_10_116 ( 
    i_10_116_174_0, i_10_116_175_0, i_10_116_177_0, i_10_116_260_0,
    i_10_116_268_0, i_10_116_283_0, i_10_116_294_0, i_10_116_321_0,
    i_10_116_363_0, i_10_116_438_0, i_10_116_439_0, i_10_116_459_0,
    i_10_116_465_0, i_10_116_466_0, i_10_116_510_0, i_10_116_597_0,
    i_10_116_749_0, i_10_116_897_0, i_10_116_993_0, i_10_116_1005_0,
    i_10_116_1033_0, i_10_116_1034_0, i_10_116_1138_0, i_10_116_1236_0,
    i_10_116_1239_0, i_10_116_1299_0, i_10_116_1306_0, i_10_116_1311_0,
    i_10_116_1312_0, i_10_116_1347_0, i_10_116_1365_0, i_10_116_1445_0,
    i_10_116_1446_0, i_10_116_1455_0, i_10_116_1822_0, i_10_116_2022_0,
    i_10_116_2112_0, i_10_116_2253_0, i_10_116_2265_0, i_10_116_2293_0,
    i_10_116_2352_0, i_10_116_2353_0, i_10_116_2364_0, i_10_116_2365_0,
    i_10_116_2452_0, i_10_116_2454_0, i_10_116_2455_0, i_10_116_2474_0,
    i_10_116_2479_0, i_10_116_2568_0, i_10_116_2571_0, i_10_116_2604_0,
    i_10_116_2643_0, i_10_116_2663_0, i_10_116_2680_0, i_10_116_2712_0,
    i_10_116_2715_0, i_10_116_2734_0, i_10_116_2784_0, i_10_116_2882_0,
    i_10_116_2884_0, i_10_116_2959_0, i_10_116_3045_0, i_10_116_3048_0,
    i_10_116_3072_0, i_10_116_3075_0, i_10_116_3198_0, i_10_116_3237_0,
    i_10_116_3273_0, i_10_116_3275_0, i_10_116_3282_0, i_10_116_3318_0,
    i_10_116_3336_0, i_10_116_3354_0, i_10_116_3388_0, i_10_116_3390_0,
    i_10_116_3392_0, i_10_116_3407_0, i_10_116_3470_0, i_10_116_3538_0,
    i_10_116_3543_0, i_10_116_3559_0, i_10_116_3561_0, i_10_116_3585_0,
    i_10_116_3813_0, i_10_116_3837_0, i_10_116_3845_0, i_10_116_3859_0,
    i_10_116_3903_0, i_10_116_3984_0, i_10_116_3985_0, i_10_116_3988_0,
    i_10_116_4056_0, i_10_116_4117_0, i_10_116_4120_0, i_10_116_4128_0,
    i_10_116_4173_0, i_10_116_4236_0, i_10_116_4292_0, i_10_116_4434_0,
    o_10_116_0_0  );
  input  i_10_116_174_0, i_10_116_175_0, i_10_116_177_0, i_10_116_260_0,
    i_10_116_268_0, i_10_116_283_0, i_10_116_294_0, i_10_116_321_0,
    i_10_116_363_0, i_10_116_438_0, i_10_116_439_0, i_10_116_459_0,
    i_10_116_465_0, i_10_116_466_0, i_10_116_510_0, i_10_116_597_0,
    i_10_116_749_0, i_10_116_897_0, i_10_116_993_0, i_10_116_1005_0,
    i_10_116_1033_0, i_10_116_1034_0, i_10_116_1138_0, i_10_116_1236_0,
    i_10_116_1239_0, i_10_116_1299_0, i_10_116_1306_0, i_10_116_1311_0,
    i_10_116_1312_0, i_10_116_1347_0, i_10_116_1365_0, i_10_116_1445_0,
    i_10_116_1446_0, i_10_116_1455_0, i_10_116_1822_0, i_10_116_2022_0,
    i_10_116_2112_0, i_10_116_2253_0, i_10_116_2265_0, i_10_116_2293_0,
    i_10_116_2352_0, i_10_116_2353_0, i_10_116_2364_0, i_10_116_2365_0,
    i_10_116_2452_0, i_10_116_2454_0, i_10_116_2455_0, i_10_116_2474_0,
    i_10_116_2479_0, i_10_116_2568_0, i_10_116_2571_0, i_10_116_2604_0,
    i_10_116_2643_0, i_10_116_2663_0, i_10_116_2680_0, i_10_116_2712_0,
    i_10_116_2715_0, i_10_116_2734_0, i_10_116_2784_0, i_10_116_2882_0,
    i_10_116_2884_0, i_10_116_2959_0, i_10_116_3045_0, i_10_116_3048_0,
    i_10_116_3072_0, i_10_116_3075_0, i_10_116_3198_0, i_10_116_3237_0,
    i_10_116_3273_0, i_10_116_3275_0, i_10_116_3282_0, i_10_116_3318_0,
    i_10_116_3336_0, i_10_116_3354_0, i_10_116_3388_0, i_10_116_3390_0,
    i_10_116_3392_0, i_10_116_3407_0, i_10_116_3470_0, i_10_116_3538_0,
    i_10_116_3543_0, i_10_116_3559_0, i_10_116_3561_0, i_10_116_3585_0,
    i_10_116_3813_0, i_10_116_3837_0, i_10_116_3845_0, i_10_116_3859_0,
    i_10_116_3903_0, i_10_116_3984_0, i_10_116_3985_0, i_10_116_3988_0,
    i_10_116_4056_0, i_10_116_4117_0, i_10_116_4120_0, i_10_116_4128_0,
    i_10_116_4173_0, i_10_116_4236_0, i_10_116_4292_0, i_10_116_4434_0;
  output o_10_116_0_0;
  assign o_10_116_0_0 = ~((~i_10_116_294_0 & ((~i_10_116_897_0 & ~i_10_116_1822_0 & ~i_10_116_2022_0 & ~i_10_116_2604_0 & ~i_10_116_3543_0 & ~i_10_116_3985_0) | (~i_10_116_2571_0 & ~i_10_116_2643_0 & ~i_10_116_3075_0 & i_10_116_3388_0 & ~i_10_116_4056_0))) | (~i_10_116_1005_0 & ((i_10_116_1311_0 & ~i_10_116_3237_0 & ~i_10_116_3273_0) | (~i_10_116_3072_0 & ~i_10_116_3392_0 & ~i_10_116_3585_0 & ~i_10_116_4128_0))) | (~i_10_116_2365_0 & ((~i_10_116_1306_0 & i_10_116_2364_0 & i_10_116_2454_0) | (i_10_116_1822_0 & ~i_10_116_2022_0 & ~i_10_116_2712_0 & ~i_10_116_3072_0 & ~i_10_116_4236_0 & ~i_10_116_4292_0))) | (~i_10_116_1446_0 & ((~i_10_116_2571_0 & ((~i_10_116_1347_0 & ~i_10_116_3282_0 & ~i_10_116_3390_0 & ~i_10_116_3392_0 & ~i_10_116_3984_0) | (~i_10_116_260_0 & ~i_10_116_3072_0 & ~i_10_116_4128_0 & ~i_10_116_4236_0))) | (~i_10_116_2364_0 & ~i_10_116_2455_0 & ~i_10_116_3538_0 & i_10_116_3837_0 & ~i_10_116_3985_0 & ~i_10_116_4173_0))) | (~i_10_116_2364_0 & ((~i_10_116_897_0 & ~i_10_116_1239_0 & ~i_10_116_3198_0 & i_10_116_3837_0) | (~i_10_116_3075_0 & ~i_10_116_3273_0 & ~i_10_116_3543_0 & ~i_10_116_4173_0))) | (~i_10_116_897_0 & ((~i_10_116_2715_0 & ~i_10_116_3075_0 & ~i_10_116_3275_0 & ~i_10_116_3390_0) | (i_10_116_2680_0 & ~i_10_116_4056_0))) | (~i_10_116_2643_0 & ((~i_10_116_2479_0 & i_10_116_2680_0 & ~i_10_116_3585_0) | (~i_10_116_459_0 & ~i_10_116_2784_0 & i_10_116_3392_0 & ~i_10_116_3985_0 & i_10_116_4128_0 & ~i_10_116_4173_0))) | (~i_10_116_3407_0 & ((i_10_116_3859_0 & ((~i_10_116_1365_0 & i_10_116_2734_0 & ~i_10_116_3045_0 & i_10_116_3390_0) | (~i_10_116_175_0 & ~i_10_116_438_0 & ~i_10_116_993_0 & ~i_10_116_2353_0 & ~i_10_116_3984_0))) | (~i_10_116_2352_0 & ~i_10_116_2712_0 & ~i_10_116_4173_0))) | (i_10_116_465_0 & i_10_116_1365_0) | (i_10_116_260_0 & i_10_116_1311_0 & ~i_10_116_3275_0) | (i_10_116_1312_0 & ~i_10_116_3845_0 & i_10_116_4120_0));
endmodule



// Benchmark "kernel_10_117" written by ABC on Sun Jul 19 10:22:59 2020

module kernel_10_117 ( 
    i_10_117_161_0, i_10_117_222_0, i_10_117_224_0, i_10_117_251_0,
    i_10_117_293_0, i_10_117_295_0, i_10_117_296_0, i_10_117_409_0,
    i_10_117_410_0, i_10_117_412_0, i_10_117_436_0, i_10_117_448_0,
    i_10_117_449_0, i_10_117_462_0, i_10_117_467_0, i_10_117_629_0,
    i_10_117_800_0, i_10_117_898_0, i_10_117_899_0, i_10_117_997_0,
    i_10_117_1033_0, i_10_117_1034_0, i_10_117_1051_0, i_10_117_1239_0,
    i_10_117_1263_0, i_10_117_1309_0, i_10_117_1365_0, i_10_117_1435_0,
    i_10_117_1650_0, i_10_117_1652_0, i_10_117_1654_0, i_10_117_1655_0,
    i_10_117_1687_0, i_10_117_1816_0, i_10_117_1817_0, i_10_117_1818_0,
    i_10_117_1912_0, i_10_117_1950_0, i_10_117_1997_0, i_10_117_2360_0,
    i_10_117_2362_0, i_10_117_2383_0, i_10_117_2455_0, i_10_117_2470_0,
    i_10_117_2471_0, i_10_117_2472_0, i_10_117_2516_0, i_10_117_2654_0,
    i_10_117_2658_0, i_10_117_2661_0, i_10_117_2662_0, i_10_117_2680_0,
    i_10_117_2720_0, i_10_117_2724_0, i_10_117_2725_0, i_10_117_2734_0,
    i_10_117_2735_0, i_10_117_2833_0, i_10_117_2924_0, i_10_117_2986_0,
    i_10_117_3153_0, i_10_117_3154_0, i_10_117_3155_0, i_10_117_3157_0,
    i_10_117_3166_0, i_10_117_3281_0, i_10_117_3544_0, i_10_117_3561_0,
    i_10_117_3586_0, i_10_117_3589_0, i_10_117_3616_0, i_10_117_3617_0,
    i_10_117_3720_0, i_10_117_3733_0, i_10_117_3734_0, i_10_117_3784_0,
    i_10_117_3813_0, i_10_117_3814_0, i_10_117_3815_0, i_10_117_3834_0,
    i_10_117_3835_0, i_10_117_3836_0, i_10_117_3840_0, i_10_117_3841_0,
    i_10_117_3842_0, i_10_117_4117_0, i_10_117_4121_0, i_10_117_4129_0,
    i_10_117_4130_0, i_10_117_4173_0, i_10_117_4174_0, i_10_117_4219_0,
    i_10_117_4220_0, i_10_117_4266_0, i_10_117_4267_0, i_10_117_4270_0,
    i_10_117_4289_0, i_10_117_4290_0, i_10_117_4292_0, i_10_117_4566_0,
    o_10_117_0_0  );
  input  i_10_117_161_0, i_10_117_222_0, i_10_117_224_0, i_10_117_251_0,
    i_10_117_293_0, i_10_117_295_0, i_10_117_296_0, i_10_117_409_0,
    i_10_117_410_0, i_10_117_412_0, i_10_117_436_0, i_10_117_448_0,
    i_10_117_449_0, i_10_117_462_0, i_10_117_467_0, i_10_117_629_0,
    i_10_117_800_0, i_10_117_898_0, i_10_117_899_0, i_10_117_997_0,
    i_10_117_1033_0, i_10_117_1034_0, i_10_117_1051_0, i_10_117_1239_0,
    i_10_117_1263_0, i_10_117_1309_0, i_10_117_1365_0, i_10_117_1435_0,
    i_10_117_1650_0, i_10_117_1652_0, i_10_117_1654_0, i_10_117_1655_0,
    i_10_117_1687_0, i_10_117_1816_0, i_10_117_1817_0, i_10_117_1818_0,
    i_10_117_1912_0, i_10_117_1950_0, i_10_117_1997_0, i_10_117_2360_0,
    i_10_117_2362_0, i_10_117_2383_0, i_10_117_2455_0, i_10_117_2470_0,
    i_10_117_2471_0, i_10_117_2472_0, i_10_117_2516_0, i_10_117_2654_0,
    i_10_117_2658_0, i_10_117_2661_0, i_10_117_2662_0, i_10_117_2680_0,
    i_10_117_2720_0, i_10_117_2724_0, i_10_117_2725_0, i_10_117_2734_0,
    i_10_117_2735_0, i_10_117_2833_0, i_10_117_2924_0, i_10_117_2986_0,
    i_10_117_3153_0, i_10_117_3154_0, i_10_117_3155_0, i_10_117_3157_0,
    i_10_117_3166_0, i_10_117_3281_0, i_10_117_3544_0, i_10_117_3561_0,
    i_10_117_3586_0, i_10_117_3589_0, i_10_117_3616_0, i_10_117_3617_0,
    i_10_117_3720_0, i_10_117_3733_0, i_10_117_3734_0, i_10_117_3784_0,
    i_10_117_3813_0, i_10_117_3814_0, i_10_117_3815_0, i_10_117_3834_0,
    i_10_117_3835_0, i_10_117_3836_0, i_10_117_3840_0, i_10_117_3841_0,
    i_10_117_3842_0, i_10_117_4117_0, i_10_117_4121_0, i_10_117_4129_0,
    i_10_117_4130_0, i_10_117_4173_0, i_10_117_4174_0, i_10_117_4219_0,
    i_10_117_4220_0, i_10_117_4266_0, i_10_117_4267_0, i_10_117_4270_0,
    i_10_117_4289_0, i_10_117_4290_0, i_10_117_4292_0, i_10_117_4566_0;
  output o_10_117_0_0;
  assign o_10_117_0_0 = ~((~i_10_117_293_0 & ((~i_10_117_295_0 & ~i_10_117_3166_0 & ((~i_10_117_251_0 & ~i_10_117_296_0 & ~i_10_117_1816_0 & ~i_10_117_2362_0 & ~i_10_117_3734_0) | (~i_10_117_410_0 & ~i_10_117_1034_0 & ~i_10_117_1365_0 & ~i_10_117_3617_0 & ~i_10_117_4130_0))) | (~i_10_117_410_0 & ((~i_10_117_1034_0 & ~i_10_117_2735_0 & ~i_10_117_4129_0) | (~i_10_117_409_0 & ~i_10_117_899_0 & ~i_10_117_1817_0 & ~i_10_117_2383_0 & ~i_10_117_2734_0 & ~i_10_117_2986_0 & ~i_10_117_4219_0))) | (~i_10_117_4130_0 & ~i_10_117_4220_0 & ((~i_10_117_997_0 & ~i_10_117_1950_0 & i_10_117_2734_0 & ~i_10_117_3733_0) | (~i_10_117_2735_0 & ~i_10_117_4129_0 & ~i_10_117_222_0 & ~i_10_117_2383_0))) | (~i_10_117_1365_0 & ~i_10_117_2734_0 & ~i_10_117_3734_0 & ~i_10_117_3784_0 & i_10_117_4566_0))) | (~i_10_117_222_0 & ((i_10_117_1435_0 & i_10_117_1687_0) | (~i_10_117_1654_0 & i_10_117_3784_0 & i_10_117_4566_0))) | (~i_10_117_251_0 & ((i_10_117_2658_0 & i_10_117_2725_0 & ~i_10_117_3166_0 & i_10_117_4121_0 & ~i_10_117_4130_0) | (~i_10_117_1239_0 & ~i_10_117_2360_0 & ~i_10_117_2680_0 & ~i_10_117_3589_0 & ~i_10_117_4219_0 & ~i_10_117_4289_0 & ~i_10_117_4292_0))) | (~i_10_117_899_0 & ((~i_10_117_410_0 & ~i_10_117_1034_0 & ~i_10_117_1263_0 & ~i_10_117_1654_0 & ~i_10_117_2986_0 & ~i_10_117_3834_0) | (~i_10_117_412_0 & ~i_10_117_436_0 & ~i_10_117_467_0 & ~i_10_117_2720_0 & i_10_117_3841_0 & i_10_117_3842_0))) | (i_10_117_1435_0 & (i_10_117_4566_0 | (i_10_117_1687_0 & ~i_10_117_2455_0))) | (~i_10_117_1655_0 & ((~i_10_117_2661_0 & i_10_117_2833_0 & ~i_10_117_4292_0) | (~i_10_117_224_0 & i_10_117_3784_0 & i_10_117_4566_0))) | (~i_10_117_4130_0 & ((i_10_117_1650_0 & ~i_10_117_2661_0 & i_10_117_3617_0 & ~i_10_117_3836_0) | (~i_10_117_1033_0 & ~i_10_117_1239_0 & ~i_10_117_2360_0 & ~i_10_117_2724_0 & ~i_10_117_2725_0 & ~i_10_117_3586_0 & ~i_10_117_3841_0))) | (~i_10_117_409_0 & ~i_10_117_2455_0 & i_10_117_3586_0 & i_10_117_4117_0));
endmodule



// Benchmark "kernel_10_118" written by ABC on Sun Jul 19 10:23:00 2020

module kernel_10_118 ( 
    i_10_118_155_0, i_10_118_157_0, i_10_118_174_0, i_10_118_180_0,
    i_10_118_248_0, i_10_118_281_0, i_10_118_317_0, i_10_118_413_0,
    i_10_118_428_0, i_10_118_442_0, i_10_118_443_0, i_10_118_444_0,
    i_10_118_445_0, i_10_118_463_0, i_10_118_464_0, i_10_118_497_0,
    i_10_118_689_0, i_10_118_799_0, i_10_118_800_0, i_10_118_820_0,
    i_10_118_997_0, i_10_118_1235_0, i_10_118_1237_0, i_10_118_1248_0,
    i_10_118_1306_0, i_10_118_1354_0, i_10_118_1359_0, i_10_118_1489_0,
    i_10_118_1543_0, i_10_118_1577_0, i_10_118_1580_0, i_10_118_1683_0,
    i_10_118_1684_0, i_10_118_1685_0, i_10_118_1686_0, i_10_118_1688_0,
    i_10_118_1689_0, i_10_118_1914_0, i_10_118_1916_0, i_10_118_1946_0,
    i_10_118_2019_0, i_10_118_2020_0, i_10_118_2026_0, i_10_118_2351_0,
    i_10_118_2358_0, i_10_118_2365_0, i_10_118_2378_0, i_10_118_2467_0,
    i_10_118_2470_0, i_10_118_2515_0, i_10_118_2632_0, i_10_118_2662_0,
    i_10_118_2704_0, i_10_118_2705_0, i_10_118_2710_0, i_10_118_2723_0,
    i_10_118_2727_0, i_10_118_2728_0, i_10_118_2735_0, i_10_118_2979_0,
    i_10_118_2986_0, i_10_118_2987_0, i_10_118_3033_0, i_10_118_3036_0,
    i_10_118_3202_0, i_10_118_3269_0, i_10_118_3274_0, i_10_118_3277_0,
    i_10_118_3280_0, i_10_118_3281_0, i_10_118_3314_0, i_10_118_3384_0,
    i_10_118_3387_0, i_10_118_3522_0, i_10_118_3611_0, i_10_118_3614_0,
    i_10_118_3728_0, i_10_118_3787_0, i_10_118_3800_0, i_10_118_3836_0,
    i_10_118_3896_0, i_10_118_3946_0, i_10_118_4114_0, i_10_118_4116_0,
    i_10_118_4118_0, i_10_118_4123_0, i_10_118_4124_0, i_10_118_4126_0,
    i_10_118_4127_0, i_10_118_4168_0, i_10_118_4169_0, i_10_118_4171_0,
    i_10_118_4172_0, i_10_118_4173_0, i_10_118_4270_0, i_10_118_4280_0,
    i_10_118_4283_0, i_10_118_4284_0, i_10_118_4291_0, i_10_118_4415_0,
    o_10_118_0_0  );
  input  i_10_118_155_0, i_10_118_157_0, i_10_118_174_0, i_10_118_180_0,
    i_10_118_248_0, i_10_118_281_0, i_10_118_317_0, i_10_118_413_0,
    i_10_118_428_0, i_10_118_442_0, i_10_118_443_0, i_10_118_444_0,
    i_10_118_445_0, i_10_118_463_0, i_10_118_464_0, i_10_118_497_0,
    i_10_118_689_0, i_10_118_799_0, i_10_118_800_0, i_10_118_820_0,
    i_10_118_997_0, i_10_118_1235_0, i_10_118_1237_0, i_10_118_1248_0,
    i_10_118_1306_0, i_10_118_1354_0, i_10_118_1359_0, i_10_118_1489_0,
    i_10_118_1543_0, i_10_118_1577_0, i_10_118_1580_0, i_10_118_1683_0,
    i_10_118_1684_0, i_10_118_1685_0, i_10_118_1686_0, i_10_118_1688_0,
    i_10_118_1689_0, i_10_118_1914_0, i_10_118_1916_0, i_10_118_1946_0,
    i_10_118_2019_0, i_10_118_2020_0, i_10_118_2026_0, i_10_118_2351_0,
    i_10_118_2358_0, i_10_118_2365_0, i_10_118_2378_0, i_10_118_2467_0,
    i_10_118_2470_0, i_10_118_2515_0, i_10_118_2632_0, i_10_118_2662_0,
    i_10_118_2704_0, i_10_118_2705_0, i_10_118_2710_0, i_10_118_2723_0,
    i_10_118_2727_0, i_10_118_2728_0, i_10_118_2735_0, i_10_118_2979_0,
    i_10_118_2986_0, i_10_118_2987_0, i_10_118_3033_0, i_10_118_3036_0,
    i_10_118_3202_0, i_10_118_3269_0, i_10_118_3274_0, i_10_118_3277_0,
    i_10_118_3280_0, i_10_118_3281_0, i_10_118_3314_0, i_10_118_3384_0,
    i_10_118_3387_0, i_10_118_3522_0, i_10_118_3611_0, i_10_118_3614_0,
    i_10_118_3728_0, i_10_118_3787_0, i_10_118_3800_0, i_10_118_3836_0,
    i_10_118_3896_0, i_10_118_3946_0, i_10_118_4114_0, i_10_118_4116_0,
    i_10_118_4118_0, i_10_118_4123_0, i_10_118_4124_0, i_10_118_4126_0,
    i_10_118_4127_0, i_10_118_4168_0, i_10_118_4169_0, i_10_118_4171_0,
    i_10_118_4172_0, i_10_118_4173_0, i_10_118_4270_0, i_10_118_4280_0,
    i_10_118_4283_0, i_10_118_4284_0, i_10_118_4291_0, i_10_118_4415_0;
  output o_10_118_0_0;
  assign o_10_118_0_0 = 0;
endmodule



// Benchmark "kernel_10_119" written by ABC on Sun Jul 19 10:23:01 2020

module kernel_10_119 ( 
    i_10_119_250_0, i_10_119_286_0, i_10_119_446_0, i_10_119_448_0,
    i_10_119_462_0, i_10_119_754_0, i_10_119_755_0, i_10_119_795_0,
    i_10_119_796_0, i_10_119_904_0, i_10_119_955_0, i_10_119_956_0,
    i_10_119_957_0, i_10_119_958_0, i_10_119_997_0, i_10_119_1235_0,
    i_10_119_1240_0, i_10_119_1552_0, i_10_119_1654_0, i_10_119_1684_0,
    i_10_119_1686_0, i_10_119_1687_0, i_10_119_1911_0, i_10_119_1912_0,
    i_10_119_1994_0, i_10_119_2312_0, i_10_119_2357_0, i_10_119_2358_0,
    i_10_119_2359_0, i_10_119_2360_0, i_10_119_2383_0, i_10_119_2407_0,
    i_10_119_2437_0, i_10_119_2460_0, i_10_119_2464_0, i_10_119_2467_0,
    i_10_119_2468_0, i_10_119_2470_0, i_10_119_2536_0, i_10_119_2542_0,
    i_10_119_2604_0, i_10_119_2630_0, i_10_119_2631_0, i_10_119_2635_0,
    i_10_119_2660_0, i_10_119_2680_0, i_10_119_2701_0, i_10_119_2722_0,
    i_10_119_2723_0, i_10_119_2728_0, i_10_119_2729_0, i_10_119_2731_0,
    i_10_119_2781_0, i_10_119_2917_0, i_10_119_2918_0, i_10_119_2921_0,
    i_10_119_2923_0, i_10_119_2924_0, i_10_119_3041_0, i_10_119_3197_0,
    i_10_119_3201_0, i_10_119_3277_0, i_10_119_3387_0, i_10_119_3405_0,
    i_10_119_3406_0, i_10_119_3467_0, i_10_119_3494_0, i_10_119_3523_0,
    i_10_119_3583_0, i_10_119_3612_0, i_10_119_3614_0, i_10_119_3705_0,
    i_10_119_3732_0, i_10_119_3783_0, i_10_119_3784_0, i_10_119_3785_0,
    i_10_119_3786_0, i_10_119_3807_0, i_10_119_3838_0, i_10_119_3847_0,
    i_10_119_3851_0, i_10_119_3895_0, i_10_119_3980_0, i_10_119_4113_0,
    i_10_119_4114_0, i_10_119_4116_0, i_10_119_4117_0, i_10_119_4169_0,
    i_10_119_4267_0, i_10_119_4270_0, i_10_119_4274_0, i_10_119_4282_0,
    i_10_119_4283_0, i_10_119_4289_0, i_10_119_4292_0, i_10_119_4569_0,
    i_10_119_4570_0, i_10_119_4571_0, i_10_119_4580_0, i_10_119_4585_0,
    o_10_119_0_0  );
  input  i_10_119_250_0, i_10_119_286_0, i_10_119_446_0, i_10_119_448_0,
    i_10_119_462_0, i_10_119_754_0, i_10_119_755_0, i_10_119_795_0,
    i_10_119_796_0, i_10_119_904_0, i_10_119_955_0, i_10_119_956_0,
    i_10_119_957_0, i_10_119_958_0, i_10_119_997_0, i_10_119_1235_0,
    i_10_119_1240_0, i_10_119_1552_0, i_10_119_1654_0, i_10_119_1684_0,
    i_10_119_1686_0, i_10_119_1687_0, i_10_119_1911_0, i_10_119_1912_0,
    i_10_119_1994_0, i_10_119_2312_0, i_10_119_2357_0, i_10_119_2358_0,
    i_10_119_2359_0, i_10_119_2360_0, i_10_119_2383_0, i_10_119_2407_0,
    i_10_119_2437_0, i_10_119_2460_0, i_10_119_2464_0, i_10_119_2467_0,
    i_10_119_2468_0, i_10_119_2470_0, i_10_119_2536_0, i_10_119_2542_0,
    i_10_119_2604_0, i_10_119_2630_0, i_10_119_2631_0, i_10_119_2635_0,
    i_10_119_2660_0, i_10_119_2680_0, i_10_119_2701_0, i_10_119_2722_0,
    i_10_119_2723_0, i_10_119_2728_0, i_10_119_2729_0, i_10_119_2731_0,
    i_10_119_2781_0, i_10_119_2917_0, i_10_119_2918_0, i_10_119_2921_0,
    i_10_119_2923_0, i_10_119_2924_0, i_10_119_3041_0, i_10_119_3197_0,
    i_10_119_3201_0, i_10_119_3277_0, i_10_119_3387_0, i_10_119_3405_0,
    i_10_119_3406_0, i_10_119_3467_0, i_10_119_3494_0, i_10_119_3523_0,
    i_10_119_3583_0, i_10_119_3612_0, i_10_119_3614_0, i_10_119_3705_0,
    i_10_119_3732_0, i_10_119_3783_0, i_10_119_3784_0, i_10_119_3785_0,
    i_10_119_3786_0, i_10_119_3807_0, i_10_119_3838_0, i_10_119_3847_0,
    i_10_119_3851_0, i_10_119_3895_0, i_10_119_3980_0, i_10_119_4113_0,
    i_10_119_4114_0, i_10_119_4116_0, i_10_119_4117_0, i_10_119_4169_0,
    i_10_119_4267_0, i_10_119_4270_0, i_10_119_4274_0, i_10_119_4282_0,
    i_10_119_4283_0, i_10_119_4289_0, i_10_119_4292_0, i_10_119_4569_0,
    i_10_119_4570_0, i_10_119_4571_0, i_10_119_4580_0, i_10_119_4585_0;
  output o_10_119_0_0;
  assign o_10_119_0_0 = 0;
endmodule



// Benchmark "kernel_10_120" written by ABC on Sun Jul 19 10:23:03 2020

module kernel_10_120 ( 
    i_10_120_28_0, i_10_120_119_0, i_10_120_122_0, i_10_120_172_0,
    i_10_120_174_0, i_10_120_175_0, i_10_120_280_0, i_10_120_281_0,
    i_10_120_424_0, i_10_120_425_0, i_10_120_432_0, i_10_120_433_0,
    i_10_120_434_0, i_10_120_436_0, i_10_120_437_0, i_10_120_449_0,
    i_10_120_459_0, i_10_120_992_0, i_10_120_1044_0, i_10_120_1045_0,
    i_10_120_1197_0, i_10_120_1233_0, i_10_120_1236_0, i_10_120_1239_0,
    i_10_120_1305_0, i_10_120_1308_0, i_10_120_1309_0, i_10_120_1310_0,
    i_10_120_1312_0, i_10_120_1540_0, i_10_120_1580_0, i_10_120_1612_0,
    i_10_120_1651_0, i_10_120_1652_0, i_10_120_1686_0, i_10_120_1687_0,
    i_10_120_1688_0, i_10_120_1689_0, i_10_120_1824_0, i_10_120_1946_0,
    i_10_120_1991_0, i_10_120_2030_0, i_10_120_2179_0, i_10_120_2204_0,
    i_10_120_2349_0, i_10_120_2350_0, i_10_120_2359_0, i_10_120_2360_0,
    i_10_120_2362_0, i_10_120_2377_0, i_10_120_2448_0, i_10_120_2457_0,
    i_10_120_2512_0, i_10_120_2513_0, i_10_120_2628_0, i_10_120_2629_0,
    i_10_120_2630_0, i_10_120_2633_0, i_10_120_2636_0, i_10_120_2659_0,
    i_10_120_2660_0, i_10_120_2663_0, i_10_120_2675_0, i_10_120_2723_0,
    i_10_120_2830_0, i_10_120_2831_0, i_10_120_2832_0, i_10_120_2917_0,
    i_10_120_2919_0, i_10_120_2983_0, i_10_120_3046_0, i_10_120_3050_0,
    i_10_120_3087_0, i_10_120_3323_0, i_10_120_3326_0, i_10_120_3350_0,
    i_10_120_3392_0, i_10_120_3402_0, i_10_120_3403_0, i_10_120_3404_0,
    i_10_120_3406_0, i_10_120_3551_0, i_10_120_3614_0, i_10_120_3650_0,
    i_10_120_3782_0, i_10_120_3785_0, i_10_120_3834_0, i_10_120_3836_0,
    i_10_120_3838_0, i_10_120_3848_0, i_10_120_3853_0, i_10_120_3854_0,
    i_10_120_3855_0, i_10_120_3856_0, i_10_120_3858_0, i_10_120_3980_0,
    i_10_120_3988_0, i_10_120_4028_0, i_10_120_4216_0, i_10_120_4266_0,
    o_10_120_0_0  );
  input  i_10_120_28_0, i_10_120_119_0, i_10_120_122_0, i_10_120_172_0,
    i_10_120_174_0, i_10_120_175_0, i_10_120_280_0, i_10_120_281_0,
    i_10_120_424_0, i_10_120_425_0, i_10_120_432_0, i_10_120_433_0,
    i_10_120_434_0, i_10_120_436_0, i_10_120_437_0, i_10_120_449_0,
    i_10_120_459_0, i_10_120_992_0, i_10_120_1044_0, i_10_120_1045_0,
    i_10_120_1197_0, i_10_120_1233_0, i_10_120_1236_0, i_10_120_1239_0,
    i_10_120_1305_0, i_10_120_1308_0, i_10_120_1309_0, i_10_120_1310_0,
    i_10_120_1312_0, i_10_120_1540_0, i_10_120_1580_0, i_10_120_1612_0,
    i_10_120_1651_0, i_10_120_1652_0, i_10_120_1686_0, i_10_120_1687_0,
    i_10_120_1688_0, i_10_120_1689_0, i_10_120_1824_0, i_10_120_1946_0,
    i_10_120_1991_0, i_10_120_2030_0, i_10_120_2179_0, i_10_120_2204_0,
    i_10_120_2349_0, i_10_120_2350_0, i_10_120_2359_0, i_10_120_2360_0,
    i_10_120_2362_0, i_10_120_2377_0, i_10_120_2448_0, i_10_120_2457_0,
    i_10_120_2512_0, i_10_120_2513_0, i_10_120_2628_0, i_10_120_2629_0,
    i_10_120_2630_0, i_10_120_2633_0, i_10_120_2636_0, i_10_120_2659_0,
    i_10_120_2660_0, i_10_120_2663_0, i_10_120_2675_0, i_10_120_2723_0,
    i_10_120_2830_0, i_10_120_2831_0, i_10_120_2832_0, i_10_120_2917_0,
    i_10_120_2919_0, i_10_120_2983_0, i_10_120_3046_0, i_10_120_3050_0,
    i_10_120_3087_0, i_10_120_3323_0, i_10_120_3326_0, i_10_120_3350_0,
    i_10_120_3392_0, i_10_120_3402_0, i_10_120_3403_0, i_10_120_3404_0,
    i_10_120_3406_0, i_10_120_3551_0, i_10_120_3614_0, i_10_120_3650_0,
    i_10_120_3782_0, i_10_120_3785_0, i_10_120_3834_0, i_10_120_3836_0,
    i_10_120_3838_0, i_10_120_3848_0, i_10_120_3853_0, i_10_120_3854_0,
    i_10_120_3855_0, i_10_120_3856_0, i_10_120_3858_0, i_10_120_3980_0,
    i_10_120_3988_0, i_10_120_4028_0, i_10_120_4216_0, i_10_120_4266_0;
  output o_10_120_0_0;
  assign o_10_120_0_0 = ~((~i_10_120_28_0 & ((i_10_120_174_0 & ~i_10_120_425_0 & ~i_10_120_2675_0) | (~i_10_120_122_0 & ~i_10_120_436_0 & ~i_10_120_437_0 & i_10_120_1309_0 & i_10_120_1310_0 & ~i_10_120_1946_0 & ~i_10_120_2359_0 & ~i_10_120_2633_0 & ~i_10_120_3046_0 & ~i_10_120_3404_0))) | (~i_10_120_2179_0 & ((~i_10_120_432_0 & ((i_10_120_174_0 & ~i_10_120_2919_0 & ~i_10_120_3404_0) | (~i_10_120_424_0 & i_10_120_1824_0 & ~i_10_120_2675_0 & ~i_10_120_3406_0))) | (i_10_120_2636_0 & ((i_10_120_1946_0 & i_10_120_2350_0) | (~i_10_120_434_0 & ~i_10_120_2663_0 & i_10_120_2983_0 & ~i_10_120_3551_0))) | (~i_10_120_437_0 & i_10_120_1236_0 & ~i_10_120_1689_0) | (~i_10_120_2377_0 & ~i_10_120_2630_0 & ~i_10_120_2663_0 & ~i_10_120_2831_0 & ~i_10_120_3785_0))) | (~i_10_120_424_0 & ((~i_10_120_1308_0 & ~i_10_120_1309_0 & ~i_10_120_2360_0 & ~i_10_120_2675_0 & ~i_10_120_3404_0) | (~i_10_120_3650_0 & i_10_120_4266_0))) | (~i_10_120_122_0 & ((~i_10_120_434_0 & ((i_10_120_459_0 & ~i_10_120_1612_0 & ~i_10_120_2359_0 & ~i_10_120_2675_0 & ~i_10_120_2832_0) | (~i_10_120_992_0 & ~i_10_120_2630_0 & i_10_120_3614_0 & i_10_120_3836_0 & ~i_10_120_4216_0))) | (~i_10_120_436_0 & ~i_10_120_449_0 & ~i_10_120_1612_0 & ~i_10_120_2349_0 & ~i_10_120_2360_0 & ~i_10_120_2630_0 & ~i_10_120_3046_0 & ~i_10_120_3402_0 & ~i_10_120_4216_0) | (~i_10_120_2362_0 & ~i_10_120_2629_0 & i_10_120_2831_0 & ~i_10_120_3855_0 & i_10_120_4028_0))) | (~i_10_120_1612_0 & ((~i_10_120_175_0 & ~i_10_120_992_0 & i_10_120_2636_0 & ~i_10_120_2659_0 & ~i_10_120_2660_0 & ~i_10_120_2675_0 & ~i_10_120_3087_0 & ~i_10_120_3650_0) | (~i_10_120_1310_0 & ~i_10_120_2359_0 & ~i_10_120_2362_0 & ~i_10_120_2831_0 & ~i_10_120_3050_0 & i_10_120_3853_0 & ~i_10_120_3988_0))) | (~i_10_120_992_0 & ((i_10_120_1652_0 & ~i_10_120_2629_0 & ~i_10_120_2630_0 & ~i_10_120_2675_0 & ~i_10_120_3087_0) | (~i_10_120_1652_0 & ~i_10_120_1824_0 & ~i_10_120_1946_0 & ~i_10_120_2377_0 & ~i_10_120_2628_0 & ~i_10_120_3614_0 & ~i_10_120_3856_0))) | (~i_10_120_2359_0 & ((~i_10_120_1651_0 & ((~i_10_120_437_0 & ~i_10_120_3406_0 & ~i_10_120_3614_0 & i_10_120_3855_0) | (~i_10_120_1824_0 & ~i_10_120_2630_0 & ~i_10_120_2675_0 & ~i_10_120_2830_0 & ~i_10_120_3785_0 & ~i_10_120_3980_0))) | (~i_10_120_2659_0 & i_10_120_2660_0 & ~i_10_120_2675_0 & ~i_10_120_2917_0 & ~i_10_120_3551_0 & ~i_10_120_3858_0))) | (~i_10_120_2629_0 & ((~i_10_120_2830_0 & ~i_10_120_3392_0 & i_10_120_3403_0) | (~i_10_120_2663_0 & i_10_120_2723_0 & i_10_120_3855_0))) | (~i_10_120_2630_0 & ((~i_10_120_1310_0 & ~i_10_120_2457_0 & ~i_10_120_2660_0 & ~i_10_120_3087_0 & ~i_10_120_3614_0) | (~i_10_120_1580_0 & ~i_10_120_2633_0 & ~i_10_120_2919_0 & ~i_10_120_3046_0 & ~i_10_120_3050_0 & ~i_10_120_3853_0 & ~i_10_120_3988_0))) | (~i_10_120_1309_0 & ((~i_10_120_1310_0 & ~i_10_120_4216_0 & ((~i_10_120_1686_0 & ~i_10_120_2636_0 & ~i_10_120_2663_0 & ~i_10_120_2917_0 & ~i_10_120_3980_0) | (~i_10_120_174_0 & ~i_10_120_425_0 & ~i_10_120_3855_0 & ~i_10_120_3858_0 & ~i_10_120_4028_0))) | (i_10_120_449_0 & ~i_10_120_3551_0 & ~i_10_120_3838_0 & ~i_10_120_3980_0))) | (~i_10_120_3406_0 & ((i_10_120_280_0 & i_10_120_281_0 & ~i_10_120_2377_0 & ~i_10_120_2675_0) | (~i_10_120_1540_0 & i_10_120_1687_0 & ~i_10_120_3854_0 & ~i_10_120_3856_0))) | (i_10_120_2349_0 & i_10_120_2917_0) | (i_10_120_2983_0 & i_10_120_3050_0 & i_10_120_3392_0) | (i_10_120_175_0 & ~i_10_120_1312_0 & ~i_10_120_2360_0 & ~i_10_120_3614_0) | (~i_10_120_2349_0 & ~i_10_120_2659_0 & ~i_10_120_2660_0 & i_10_120_3403_0 & ~i_10_120_3404_0 & ~i_10_120_3980_0));
endmodule



// Benchmark "kernel_10_121" written by ABC on Sun Jul 19 10:23:04 2020

module kernel_10_121 ( 
    i_10_121_176_0, i_10_121_219_0, i_10_121_220_0, i_10_121_283_0,
    i_10_121_284_0, i_10_121_285_0, i_10_121_316_0, i_10_121_317_0,
    i_10_121_443_0, i_10_121_446_0, i_10_121_447_0, i_10_121_459_0,
    i_10_121_460_0, i_10_121_462_0, i_10_121_465_0, i_10_121_623_0,
    i_10_121_793_0, i_10_121_794_0, i_10_121_796_0, i_10_121_797_0,
    i_10_121_799_0, i_10_121_962_0, i_10_121_1026_0, i_10_121_1032_0,
    i_10_121_1033_0, i_10_121_1081_0, i_10_121_1084_0, i_10_121_1235_0,
    i_10_121_1313_0, i_10_121_1546_0, i_10_121_1575_0, i_10_121_1577_0,
    i_10_121_1620_0, i_10_121_1765_0, i_10_121_1819_0, i_10_121_1820_0,
    i_10_121_1822_0, i_10_121_1825_0, i_10_121_1826_0, i_10_121_1913_0,
    i_10_121_2025_0, i_10_121_2026_0, i_10_121_2197_0, i_10_121_2199_0,
    i_10_121_2200_0, i_10_121_2350_0, i_10_121_2351_0, i_10_121_2352_0,
    i_10_121_2353_0, i_10_121_2354_0, i_10_121_2362_0, i_10_121_2380_0,
    i_10_121_2448_0, i_10_121_2450_0, i_10_121_2456_0, i_10_121_2631_0,
    i_10_121_2633_0, i_10_121_2660_0, i_10_121_2712_0, i_10_121_2722_0,
    i_10_121_2723_0, i_10_121_2727_0, i_10_121_2728_0, i_10_121_2730_0,
    i_10_121_2732_0, i_10_121_2827_0, i_10_121_2917_0, i_10_121_2920_0,
    i_10_121_2921_0, i_10_121_2924_0, i_10_121_2980_0, i_10_121_3075_0,
    i_10_121_3152_0, i_10_121_3203_0, i_10_121_3281_0, i_10_121_3384_0,
    i_10_121_3389_0, i_10_121_3391_0, i_10_121_3407_0, i_10_121_3616_0,
    i_10_121_3617_0, i_10_121_3648_0, i_10_121_3787_0, i_10_121_3839_0,
    i_10_121_3847_0, i_10_121_3857_0, i_10_121_3858_0, i_10_121_3860_0,
    i_10_121_3906_0, i_10_121_3907_0, i_10_121_4051_0, i_10_121_4118_0,
    i_10_121_4275_0, i_10_121_4276_0, i_10_121_4277_0, i_10_121_4284_0,
    i_10_121_4288_0, i_10_121_4564_0, i_10_121_4569_0, i_10_121_4570_0,
    o_10_121_0_0  );
  input  i_10_121_176_0, i_10_121_219_0, i_10_121_220_0, i_10_121_283_0,
    i_10_121_284_0, i_10_121_285_0, i_10_121_316_0, i_10_121_317_0,
    i_10_121_443_0, i_10_121_446_0, i_10_121_447_0, i_10_121_459_0,
    i_10_121_460_0, i_10_121_462_0, i_10_121_465_0, i_10_121_623_0,
    i_10_121_793_0, i_10_121_794_0, i_10_121_796_0, i_10_121_797_0,
    i_10_121_799_0, i_10_121_962_0, i_10_121_1026_0, i_10_121_1032_0,
    i_10_121_1033_0, i_10_121_1081_0, i_10_121_1084_0, i_10_121_1235_0,
    i_10_121_1313_0, i_10_121_1546_0, i_10_121_1575_0, i_10_121_1577_0,
    i_10_121_1620_0, i_10_121_1765_0, i_10_121_1819_0, i_10_121_1820_0,
    i_10_121_1822_0, i_10_121_1825_0, i_10_121_1826_0, i_10_121_1913_0,
    i_10_121_2025_0, i_10_121_2026_0, i_10_121_2197_0, i_10_121_2199_0,
    i_10_121_2200_0, i_10_121_2350_0, i_10_121_2351_0, i_10_121_2352_0,
    i_10_121_2353_0, i_10_121_2354_0, i_10_121_2362_0, i_10_121_2380_0,
    i_10_121_2448_0, i_10_121_2450_0, i_10_121_2456_0, i_10_121_2631_0,
    i_10_121_2633_0, i_10_121_2660_0, i_10_121_2712_0, i_10_121_2722_0,
    i_10_121_2723_0, i_10_121_2727_0, i_10_121_2728_0, i_10_121_2730_0,
    i_10_121_2732_0, i_10_121_2827_0, i_10_121_2917_0, i_10_121_2920_0,
    i_10_121_2921_0, i_10_121_2924_0, i_10_121_2980_0, i_10_121_3075_0,
    i_10_121_3152_0, i_10_121_3203_0, i_10_121_3281_0, i_10_121_3384_0,
    i_10_121_3389_0, i_10_121_3391_0, i_10_121_3407_0, i_10_121_3616_0,
    i_10_121_3617_0, i_10_121_3648_0, i_10_121_3787_0, i_10_121_3839_0,
    i_10_121_3847_0, i_10_121_3857_0, i_10_121_3858_0, i_10_121_3860_0,
    i_10_121_3906_0, i_10_121_3907_0, i_10_121_4051_0, i_10_121_4118_0,
    i_10_121_4275_0, i_10_121_4276_0, i_10_121_4277_0, i_10_121_4284_0,
    i_10_121_4288_0, i_10_121_4564_0, i_10_121_4569_0, i_10_121_4570_0;
  output o_10_121_0_0;
  assign o_10_121_0_0 = ~((~i_10_121_1081_0 & ((~i_10_121_285_0 & ((~i_10_121_316_0 & ~i_10_121_1032_0 & ~i_10_121_1620_0 & ~i_10_121_2362_0 & ~i_10_121_2722_0 & i_10_121_3839_0 & ~i_10_121_3907_0) | (~i_10_121_2199_0 & ~i_10_121_2352_0 & ~i_10_121_3075_0 & ~i_10_121_3391_0 & ~i_10_121_4275_0 & ~i_10_121_4277_0))) | (~i_10_121_3906_0 & ((~i_10_121_462_0 & ~i_10_121_1032_0 & ~i_10_121_1235_0 & ~i_10_121_2350_0 & ~i_10_121_2354_0) | (~i_10_121_443_0 & i_10_121_794_0 & ~i_10_121_4277_0))) | (~i_10_121_1026_0 & ~i_10_121_1033_0 & ~i_10_121_1822_0 & i_10_121_1826_0 & ~i_10_121_3203_0))) | (~i_10_121_317_0 & ((~i_10_121_2199_0 & i_10_121_2350_0 & ~i_10_121_2723_0 & ~i_10_121_2728_0 & ~i_10_121_3281_0) | (~i_10_121_1026_0 & ~i_10_121_1033_0 & ~i_10_121_316_0 & ~i_10_121_465_0 & ~i_10_121_1577_0 & ~i_10_121_1620_0 & ~i_10_121_2362_0 & ~i_10_121_2722_0 & ~i_10_121_3906_0))) | (~i_10_121_1575_0 & ((i_10_121_1819_0 & ~i_10_121_1913_0 & ~i_10_121_2352_0 & ~i_10_121_2712_0 & ~i_10_121_2732_0 & ~i_10_121_3384_0 & ~i_10_121_3787_0) | (~i_10_121_316_0 & ~i_10_121_1546_0 & ~i_10_121_2353_0 & ~i_10_121_2354_0 & ~i_10_121_3075_0 & ~i_10_121_3648_0 & ~i_10_121_3907_0))) | (~i_10_121_316_0 & ((i_10_121_1826_0 & i_10_121_2353_0 & ~i_10_121_2362_0 & ~i_10_121_3203_0) | (~i_10_121_1026_0 & ~i_10_121_1620_0 & ~i_10_121_1913_0 & ~i_10_121_3075_0 & ~i_10_121_3787_0 & ~i_10_121_3857_0 & ~i_10_121_3906_0 & ~i_10_121_4276_0 & ~i_10_121_4277_0))) | (~i_10_121_1546_0 & i_10_121_2353_0 & ((~i_10_121_962_0 & ~i_10_121_2197_0 & i_10_121_2354_0 & ~i_10_121_2660_0 & ~i_10_121_3281_0 & ~i_10_121_4276_0) | (~i_10_121_1033_0 & ~i_10_121_1913_0 & ~i_10_121_2351_0 & ~i_10_121_3075_0 & ~i_10_121_4275_0 & ~i_10_121_4277_0 & ~i_10_121_4284_0))) | (~i_10_121_1033_0 & ((i_10_121_1819_0 & i_10_121_2450_0 & ~i_10_121_2712_0 & ~i_10_121_3847_0 & ~i_10_121_3906_0) | (~i_10_121_2197_0 & ~i_10_121_2350_0 & ~i_10_121_2353_0 & ~i_10_121_3075_0 & ~i_10_121_4275_0 & ~i_10_121_4277_0))) | (~i_10_121_1822_0 & ((i_10_121_796_0 & ~i_10_121_2199_0 & ~i_10_121_2351_0) | (i_10_121_2450_0 & ~i_10_121_4276_0 & ~i_10_121_4277_0 & i_10_121_4288_0))) | (~i_10_121_2362_0 & ((i_10_121_2730_0 & i_10_121_3391_0 & i_10_121_3860_0) | (~i_10_121_1577_0 & ~i_10_121_2354_0 & ~i_10_121_2450_0 & ~i_10_121_2727_0 & ~i_10_121_2920_0 & ~i_10_121_3075_0 & ~i_10_121_3847_0 & ~i_10_121_3906_0 & ~i_10_121_4275_0))) | (~i_10_121_2732_0 & ((~i_10_121_1032_0 & ~i_10_121_1913_0 & ~i_10_121_2633_0 & ~i_10_121_2727_0 & i_10_121_2827_0 & ~i_10_121_2920_0 & ~i_10_121_3391_0 & ~i_10_121_3857_0) | (i_10_121_465_0 & ~i_10_121_2350_0 & ~i_10_121_2921_0 & ~i_10_121_3407_0 & i_10_121_3858_0 & ~i_10_121_4275_0))) | (~i_10_121_3847_0 & ((~i_10_121_4275_0 & ((~i_10_121_219_0 & ~i_10_121_797_0 & i_10_121_1313_0 & i_10_121_1826_0 & ~i_10_121_2380_0 & ~i_10_121_2712_0) | (i_10_121_1575_0 & ~i_10_121_2200_0 & ~i_10_121_2660_0 & ~i_10_121_2827_0 & ~i_10_121_3391_0))) | (i_10_121_220_0 & ~i_10_121_283_0 & i_10_121_1032_0 & ~i_10_121_3858_0))) | (~i_10_121_283_0 & ((i_10_121_1825_0 & ~i_10_121_2200_0 & ~i_10_121_3648_0) | (~i_10_121_1620_0 & i_10_121_2730_0 & i_10_121_3858_0 & ~i_10_121_3906_0 & ~i_10_121_3907_0))) | (i_10_121_797_0 & ~i_10_121_2200_0 & ~i_10_121_2351_0 & ~i_10_121_3075_0) | (~i_10_121_1826_0 & ~i_10_121_2352_0 & i_10_121_3281_0 & ~i_10_121_3389_0 & i_10_121_3391_0 & i_10_121_3857_0));
endmodule



// Benchmark "kernel_10_122" written by ABC on Sun Jul 19 10:23:05 2020

module kernel_10_122 ( 
    i_10_122_31_0, i_10_122_153_0, i_10_122_171_0, i_10_122_223_0,
    i_10_122_279_0, i_10_122_282_0, i_10_122_285_0, i_10_122_327_0,
    i_10_122_329_0, i_10_122_413_0, i_10_122_444_0, i_10_122_445_0,
    i_10_122_463_0, i_10_122_513_0, i_10_122_594_0, i_10_122_633_0,
    i_10_122_750_0, i_10_122_795_0, i_10_122_797_0, i_10_122_799_0,
    i_10_122_800_0, i_10_122_900_0, i_10_122_955_0, i_10_122_1236_0,
    i_10_122_1241_0, i_10_122_1245_0, i_10_122_1306_0, i_10_122_1309_0,
    i_10_122_1313_0, i_10_122_1435_0, i_10_122_1491_0, i_10_122_1580_0,
    i_10_122_1654_0, i_10_122_1683_0, i_10_122_1686_0, i_10_122_1791_0,
    i_10_122_1911_0, i_10_122_1936_0, i_10_122_1951_0, i_10_122_1998_0,
    i_10_122_2028_0, i_10_122_2183_0, i_10_122_2325_0, i_10_122_2349_0,
    i_10_122_2376_0, i_10_122_2451_0, i_10_122_2452_0, i_10_122_2455_0,
    i_10_122_2469_0, i_10_122_2506_0, i_10_122_2632_0, i_10_122_2634_0,
    i_10_122_2635_0, i_10_122_2636_0, i_10_122_2659_0, i_10_122_2661_0,
    i_10_122_2673_0, i_10_122_2679_0, i_10_122_2709_0, i_10_122_2712_0,
    i_10_122_2721_0, i_10_122_2722_0, i_10_122_2725_0, i_10_122_2727_0,
    i_10_122_2733_0, i_10_122_2781_0, i_10_122_2820_0, i_10_122_2910_0,
    i_10_122_3070_0, i_10_122_3071_0, i_10_122_3088_0, i_10_122_3279_0,
    i_10_122_3283_0, i_10_122_3297_0, i_10_122_3451_0, i_10_122_3492_0,
    i_10_122_3495_0, i_10_122_3585_0, i_10_122_3587_0, i_10_122_3612_0,
    i_10_122_3619_0, i_10_122_3645_0, i_10_122_3649_0, i_10_122_3724_0,
    i_10_122_3780_0, i_10_122_3781_0, i_10_122_3783_0, i_10_122_3786_0,
    i_10_122_3853_0, i_10_122_3870_0, i_10_122_3873_0, i_10_122_3912_0,
    i_10_122_3945_0, i_10_122_4114_0, i_10_122_4150_0, i_10_122_4188_0,
    i_10_122_4267_0, i_10_122_4269_0, i_10_122_4270_0, i_10_122_4461_0,
    o_10_122_0_0  );
  input  i_10_122_31_0, i_10_122_153_0, i_10_122_171_0, i_10_122_223_0,
    i_10_122_279_0, i_10_122_282_0, i_10_122_285_0, i_10_122_327_0,
    i_10_122_329_0, i_10_122_413_0, i_10_122_444_0, i_10_122_445_0,
    i_10_122_463_0, i_10_122_513_0, i_10_122_594_0, i_10_122_633_0,
    i_10_122_750_0, i_10_122_795_0, i_10_122_797_0, i_10_122_799_0,
    i_10_122_800_0, i_10_122_900_0, i_10_122_955_0, i_10_122_1236_0,
    i_10_122_1241_0, i_10_122_1245_0, i_10_122_1306_0, i_10_122_1309_0,
    i_10_122_1313_0, i_10_122_1435_0, i_10_122_1491_0, i_10_122_1580_0,
    i_10_122_1654_0, i_10_122_1683_0, i_10_122_1686_0, i_10_122_1791_0,
    i_10_122_1911_0, i_10_122_1936_0, i_10_122_1951_0, i_10_122_1998_0,
    i_10_122_2028_0, i_10_122_2183_0, i_10_122_2325_0, i_10_122_2349_0,
    i_10_122_2376_0, i_10_122_2451_0, i_10_122_2452_0, i_10_122_2455_0,
    i_10_122_2469_0, i_10_122_2506_0, i_10_122_2632_0, i_10_122_2634_0,
    i_10_122_2635_0, i_10_122_2636_0, i_10_122_2659_0, i_10_122_2661_0,
    i_10_122_2673_0, i_10_122_2679_0, i_10_122_2709_0, i_10_122_2712_0,
    i_10_122_2721_0, i_10_122_2722_0, i_10_122_2725_0, i_10_122_2727_0,
    i_10_122_2733_0, i_10_122_2781_0, i_10_122_2820_0, i_10_122_2910_0,
    i_10_122_3070_0, i_10_122_3071_0, i_10_122_3088_0, i_10_122_3279_0,
    i_10_122_3283_0, i_10_122_3297_0, i_10_122_3451_0, i_10_122_3492_0,
    i_10_122_3495_0, i_10_122_3585_0, i_10_122_3587_0, i_10_122_3612_0,
    i_10_122_3619_0, i_10_122_3645_0, i_10_122_3649_0, i_10_122_3724_0,
    i_10_122_3780_0, i_10_122_3781_0, i_10_122_3783_0, i_10_122_3786_0,
    i_10_122_3853_0, i_10_122_3870_0, i_10_122_3873_0, i_10_122_3912_0,
    i_10_122_3945_0, i_10_122_4114_0, i_10_122_4150_0, i_10_122_4188_0,
    i_10_122_4267_0, i_10_122_4269_0, i_10_122_4270_0, i_10_122_4461_0;
  output o_10_122_0_0;
  assign o_10_122_0_0 = 0;
endmodule



// Benchmark "kernel_10_123" written by ABC on Sun Jul 19 10:23:06 2020

module kernel_10_123 ( 
    i_10_123_395_0, i_10_123_405_0, i_10_123_725_0, i_10_123_728_0,
    i_10_123_799_0, i_10_123_820_0, i_10_123_928_0, i_10_123_929_0,
    i_10_123_957_0, i_10_123_958_0, i_10_123_959_0, i_10_123_961_0,
    i_10_123_989_0, i_10_123_1027_0, i_10_123_1028_0, i_10_123_1116_0,
    i_10_123_1119_0, i_10_123_1165_0, i_10_123_1239_0, i_10_123_1305_0,
    i_10_123_1311_0, i_10_123_1352_0, i_10_123_1359_0, i_10_123_1360_0,
    i_10_123_1363_0, i_10_123_1364_0, i_10_123_1394_0, i_10_123_1605_0,
    i_10_123_1606_0, i_10_123_1618_0, i_10_123_1621_0, i_10_123_1698_0,
    i_10_123_1699_0, i_10_123_1768_0, i_10_123_1786_0, i_10_123_1822_0,
    i_10_123_1823_0, i_10_123_1954_0, i_10_123_2008_0, i_10_123_2196_0,
    i_10_123_2243_0, i_10_123_2350_0, i_10_123_2353_0, i_10_123_2446_0,
    i_10_123_2452_0, i_10_123_2641_0, i_10_123_2700_0, i_10_123_2703_0,
    i_10_123_2828_0, i_10_123_2831_0, i_10_123_2856_0, i_10_123_2857_0,
    i_10_123_2868_0, i_10_123_2872_0, i_10_123_2916_0, i_10_123_2917_0,
    i_10_123_2919_0, i_10_123_2920_0, i_10_123_2921_0, i_10_123_2924_0,
    i_10_123_2935_0, i_10_123_3037_0, i_10_123_3038_0, i_10_123_3070_0,
    i_10_123_3225_0, i_10_123_3226_0, i_10_123_3234_0, i_10_123_3271_0,
    i_10_123_3306_0, i_10_123_3316_0, i_10_123_3317_0, i_10_123_3385_0,
    i_10_123_3404_0, i_10_123_3451_0, i_10_123_3455_0, i_10_123_3542_0,
    i_10_123_3543_0, i_10_123_3556_0, i_10_123_3596_0, i_10_123_3720_0,
    i_10_123_3721_0, i_10_123_3726_0, i_10_123_3727_0, i_10_123_3836_0,
    i_10_123_3848_0, i_10_123_3860_0, i_10_123_3920_0, i_10_123_3960_0,
    i_10_123_3961_0, i_10_123_3962_0, i_10_123_3964_0, i_10_123_3965_0,
    i_10_123_4136_0, i_10_123_4143_0, i_10_123_4217_0, i_10_123_4323_0,
    i_10_123_4529_0, i_10_123_4568_0, i_10_123_4574_0, i_10_123_4591_0,
    o_10_123_0_0  );
  input  i_10_123_395_0, i_10_123_405_0, i_10_123_725_0, i_10_123_728_0,
    i_10_123_799_0, i_10_123_820_0, i_10_123_928_0, i_10_123_929_0,
    i_10_123_957_0, i_10_123_958_0, i_10_123_959_0, i_10_123_961_0,
    i_10_123_989_0, i_10_123_1027_0, i_10_123_1028_0, i_10_123_1116_0,
    i_10_123_1119_0, i_10_123_1165_0, i_10_123_1239_0, i_10_123_1305_0,
    i_10_123_1311_0, i_10_123_1352_0, i_10_123_1359_0, i_10_123_1360_0,
    i_10_123_1363_0, i_10_123_1364_0, i_10_123_1394_0, i_10_123_1605_0,
    i_10_123_1606_0, i_10_123_1618_0, i_10_123_1621_0, i_10_123_1698_0,
    i_10_123_1699_0, i_10_123_1768_0, i_10_123_1786_0, i_10_123_1822_0,
    i_10_123_1823_0, i_10_123_1954_0, i_10_123_2008_0, i_10_123_2196_0,
    i_10_123_2243_0, i_10_123_2350_0, i_10_123_2353_0, i_10_123_2446_0,
    i_10_123_2452_0, i_10_123_2641_0, i_10_123_2700_0, i_10_123_2703_0,
    i_10_123_2828_0, i_10_123_2831_0, i_10_123_2856_0, i_10_123_2857_0,
    i_10_123_2868_0, i_10_123_2872_0, i_10_123_2916_0, i_10_123_2917_0,
    i_10_123_2919_0, i_10_123_2920_0, i_10_123_2921_0, i_10_123_2924_0,
    i_10_123_2935_0, i_10_123_3037_0, i_10_123_3038_0, i_10_123_3070_0,
    i_10_123_3225_0, i_10_123_3226_0, i_10_123_3234_0, i_10_123_3271_0,
    i_10_123_3306_0, i_10_123_3316_0, i_10_123_3317_0, i_10_123_3385_0,
    i_10_123_3404_0, i_10_123_3451_0, i_10_123_3455_0, i_10_123_3542_0,
    i_10_123_3543_0, i_10_123_3556_0, i_10_123_3596_0, i_10_123_3720_0,
    i_10_123_3721_0, i_10_123_3726_0, i_10_123_3727_0, i_10_123_3836_0,
    i_10_123_3848_0, i_10_123_3860_0, i_10_123_3920_0, i_10_123_3960_0,
    i_10_123_3961_0, i_10_123_3962_0, i_10_123_3964_0, i_10_123_3965_0,
    i_10_123_4136_0, i_10_123_4143_0, i_10_123_4217_0, i_10_123_4323_0,
    i_10_123_4529_0, i_10_123_4568_0, i_10_123_4574_0, i_10_123_4591_0;
  output o_10_123_0_0;
  assign o_10_123_0_0 = 0;
endmodule



// Benchmark "kernel_10_124" written by ABC on Sun Jul 19 10:23:07 2020

module kernel_10_124 ( 
    i_10_124_146_0, i_10_124_176_0, i_10_124_275_0, i_10_124_282_0,
    i_10_124_316_0, i_10_124_388_0, i_10_124_389_0, i_10_124_406_0,
    i_10_124_424_0, i_10_124_425_0, i_10_124_433_0, i_10_124_434_0,
    i_10_124_441_0, i_10_124_443_0, i_10_124_463_0, i_10_124_464_0,
    i_10_124_505_0, i_10_124_506_0, i_10_124_751_0, i_10_124_797_0,
    i_10_124_992_0, i_10_124_1028_0, i_10_124_1030_0, i_10_124_1037_0,
    i_10_124_1235_0, i_10_124_1238_0, i_10_124_1305_0, i_10_124_1313_0,
    i_10_124_1342_0, i_10_124_1343_0, i_10_124_1360_0, i_10_124_1361_0,
    i_10_124_1445_0, i_10_124_1578_0, i_10_124_1579_0, i_10_124_1580_0,
    i_10_124_1648_0, i_10_124_1650_0, i_10_124_1651_0, i_10_124_1652_0,
    i_10_124_1653_0, i_10_124_1688_0, i_10_124_1818_0, i_10_124_1821_0,
    i_10_124_2183_0, i_10_124_2197_0, i_10_124_2324_0, i_10_124_2353_0,
    i_10_124_2356_0, i_10_124_2379_0, i_10_124_2456_0, i_10_124_2471_0,
    i_10_124_2629_0, i_10_124_2630_0, i_10_124_2655_0, i_10_124_2656_0,
    i_10_124_2659_0, i_10_124_2660_0, i_10_124_2675_0, i_10_124_2711_0,
    i_10_124_2732_0, i_10_124_2919_0, i_10_124_3043_0, i_10_124_3070_0,
    i_10_124_3071_0, i_10_124_3072_0, i_10_124_3087_0, i_10_124_3088_0,
    i_10_124_3089_0, i_10_124_3353_0, i_10_124_3385_0, i_10_124_3388_0,
    i_10_124_3389_0, i_10_124_3403_0, i_10_124_3404_0, i_10_124_3406_0,
    i_10_124_3467_0, i_10_124_3523_0, i_10_124_3526_0, i_10_124_3584_0,
    i_10_124_3586_0, i_10_124_3614_0, i_10_124_3782_0, i_10_124_3784_0,
    i_10_124_3837_0, i_10_124_3838_0, i_10_124_3850_0, i_10_124_3855_0,
    i_10_124_3859_0, i_10_124_3875_0, i_10_124_3890_0, i_10_124_3944_0,
    i_10_124_3991_0, i_10_124_3992_0, i_10_124_3994_0, i_10_124_4052_0,
    i_10_124_4114_0, i_10_124_4115_0, i_10_124_4288_0, i_10_124_4291_0,
    o_10_124_0_0  );
  input  i_10_124_146_0, i_10_124_176_0, i_10_124_275_0, i_10_124_282_0,
    i_10_124_316_0, i_10_124_388_0, i_10_124_389_0, i_10_124_406_0,
    i_10_124_424_0, i_10_124_425_0, i_10_124_433_0, i_10_124_434_0,
    i_10_124_441_0, i_10_124_443_0, i_10_124_463_0, i_10_124_464_0,
    i_10_124_505_0, i_10_124_506_0, i_10_124_751_0, i_10_124_797_0,
    i_10_124_992_0, i_10_124_1028_0, i_10_124_1030_0, i_10_124_1037_0,
    i_10_124_1235_0, i_10_124_1238_0, i_10_124_1305_0, i_10_124_1313_0,
    i_10_124_1342_0, i_10_124_1343_0, i_10_124_1360_0, i_10_124_1361_0,
    i_10_124_1445_0, i_10_124_1578_0, i_10_124_1579_0, i_10_124_1580_0,
    i_10_124_1648_0, i_10_124_1650_0, i_10_124_1651_0, i_10_124_1652_0,
    i_10_124_1653_0, i_10_124_1688_0, i_10_124_1818_0, i_10_124_1821_0,
    i_10_124_2183_0, i_10_124_2197_0, i_10_124_2324_0, i_10_124_2353_0,
    i_10_124_2356_0, i_10_124_2379_0, i_10_124_2456_0, i_10_124_2471_0,
    i_10_124_2629_0, i_10_124_2630_0, i_10_124_2655_0, i_10_124_2656_0,
    i_10_124_2659_0, i_10_124_2660_0, i_10_124_2675_0, i_10_124_2711_0,
    i_10_124_2732_0, i_10_124_2919_0, i_10_124_3043_0, i_10_124_3070_0,
    i_10_124_3071_0, i_10_124_3072_0, i_10_124_3087_0, i_10_124_3088_0,
    i_10_124_3089_0, i_10_124_3353_0, i_10_124_3385_0, i_10_124_3388_0,
    i_10_124_3389_0, i_10_124_3403_0, i_10_124_3404_0, i_10_124_3406_0,
    i_10_124_3467_0, i_10_124_3523_0, i_10_124_3526_0, i_10_124_3584_0,
    i_10_124_3586_0, i_10_124_3614_0, i_10_124_3782_0, i_10_124_3784_0,
    i_10_124_3837_0, i_10_124_3838_0, i_10_124_3850_0, i_10_124_3855_0,
    i_10_124_3859_0, i_10_124_3875_0, i_10_124_3890_0, i_10_124_3944_0,
    i_10_124_3991_0, i_10_124_3992_0, i_10_124_3994_0, i_10_124_4052_0,
    i_10_124_4114_0, i_10_124_4115_0, i_10_124_4288_0, i_10_124_4291_0;
  output o_10_124_0_0;
  assign o_10_124_0_0 = ~((~i_10_124_282_0 & ((~i_10_124_434_0 & i_10_124_443_0 & ~i_10_124_3586_0 & ~i_10_124_3944_0) | (~i_10_124_389_0 & ~i_10_124_797_0 & ~i_10_124_2324_0 & ~i_10_124_3088_0 & ~i_10_124_3089_0 & ~i_10_124_3850_0 & ~i_10_124_3991_0 & ~i_10_124_3992_0))) | (~i_10_124_388_0 & ((~i_10_124_434_0 & ~i_10_124_1238_0 & ~i_10_124_2379_0 & ~i_10_124_2659_0 & ~i_10_124_3526_0 & ~i_10_124_3784_0) | (~i_10_124_1028_0 & ~i_10_124_2324_0 & ~i_10_124_2471_0 & i_10_124_3855_0 & ~i_10_124_4052_0))) | (~i_10_124_425_0 & ((~i_10_124_1235_0 & i_10_124_3523_0) | (~i_10_124_389_0 & ~i_10_124_2324_0 & ~i_10_124_3088_0 & ~i_10_124_3584_0))) | (~i_10_124_1342_0 & ((~i_10_124_2656_0 & ~i_10_124_2675_0 & ~i_10_124_3404_0) | (~i_10_124_146_0 & ~i_10_124_1361_0 & i_10_124_2656_0 & ~i_10_124_2711_0 & ~i_10_124_4052_0))) | (~i_10_124_4291_0 & ((~i_10_124_1360_0 & ((i_10_124_1652_0 & ~i_10_124_2711_0 & ~i_10_124_3850_0) | (~i_10_124_424_0 & ~i_10_124_992_0 & ~i_10_124_1361_0 & ~i_10_124_2324_0 & ~i_10_124_3784_0 & ~i_10_124_3859_0 & ~i_10_124_3944_0))) | (i_10_124_316_0 & ~i_10_124_2711_0))) | (~i_10_124_146_0 & ((~i_10_124_3087_0 & ~i_10_124_3088_0 & ~i_10_124_3992_0 & ((~i_10_124_176_0 & ~i_10_124_1028_0 & ~i_10_124_2324_0 & ~i_10_124_2379_0 & ~i_10_124_2456_0) | (~i_10_124_406_0 & ~i_10_124_3089_0 & ~i_10_124_3406_0 & ~i_10_124_4115_0))) | (~i_10_124_316_0 & ~i_10_124_434_0 & ~i_10_124_1361_0 & ~i_10_124_3385_0 & ~i_10_124_3994_0))) | (~i_10_124_1238_0 & i_10_124_1818_0 & ~i_10_124_2711_0) | (~i_10_124_3070_0 & ~i_10_124_3089_0 & ~i_10_124_3389_0 & ~i_10_124_3584_0 & ~i_10_124_4288_0));
endmodule



// Benchmark "kernel_10_125" written by ABC on Sun Jul 19 10:23:08 2020

module kernel_10_125 ( 
    i_10_125_31_0, i_10_125_32_0, i_10_125_53_0, i_10_125_86_0,
    i_10_125_178_0, i_10_125_179_0, i_10_125_329_0, i_10_125_409_0,
    i_10_125_463_0, i_10_125_465_0, i_10_125_466_0, i_10_125_467_0,
    i_10_125_507_0, i_10_125_518_0, i_10_125_628_0, i_10_125_729_0,
    i_10_125_799_0, i_10_125_955_0, i_10_125_956_0, i_10_125_1005_0,
    i_10_125_1034_0, i_10_125_1235_0, i_10_125_1238_0, i_10_125_1241_0,
    i_10_125_1247_0, i_10_125_1305_0, i_10_125_1310_0, i_10_125_1348_0,
    i_10_125_1444_0, i_10_125_1445_0, i_10_125_1653_0, i_10_125_1717_0,
    i_10_125_1718_0, i_10_125_1765_0, i_10_125_1818_0, i_10_125_1821_0,
    i_10_125_1929_0, i_10_125_1948_0, i_10_125_2022_0, i_10_125_2023_0,
    i_10_125_2181_0, i_10_125_2252_0, i_10_125_2254_0, i_10_125_2326_0,
    i_10_125_2356_0, i_10_125_2357_0, i_10_125_2410_0, i_10_125_2456_0,
    i_10_125_2467_0, i_10_125_2469_0, i_10_125_2472_0, i_10_125_2514_0,
    i_10_125_2515_0, i_10_125_2516_0, i_10_125_2519_0, i_10_125_2570_0,
    i_10_125_2631_0, i_10_125_2632_0, i_10_125_2678_0, i_10_125_2681_0,
    i_10_125_2704_0, i_10_125_2705_0, i_10_125_2713_0, i_10_125_2714_0,
    i_10_125_2717_0, i_10_125_2722_0, i_10_125_2760_0, i_10_125_2784_0,
    i_10_125_2788_0, i_10_125_2830_0, i_10_125_2831_0, i_10_125_2832_0,
    i_10_125_2884_0, i_10_125_3072_0, i_10_125_3073_0, i_10_125_3201_0,
    i_10_125_3281_0, i_10_125_3283_0, i_10_125_3386_0, i_10_125_3390_0,
    i_10_125_3391_0, i_10_125_3392_0, i_10_125_3444_0, i_10_125_3500_0,
    i_10_125_3507_0, i_10_125_3586_0, i_10_125_3587_0, i_10_125_3589_0,
    i_10_125_3590_0, i_10_125_3616_0, i_10_125_3617_0, i_10_125_3648_0,
    i_10_125_3781_0, i_10_125_3782_0, i_10_125_3844_0, i_10_125_3845_0,
    i_10_125_3858_0, i_10_125_4115_0, i_10_125_4129_0, i_10_125_4568_0,
    o_10_125_0_0  );
  input  i_10_125_31_0, i_10_125_32_0, i_10_125_53_0, i_10_125_86_0,
    i_10_125_178_0, i_10_125_179_0, i_10_125_329_0, i_10_125_409_0,
    i_10_125_463_0, i_10_125_465_0, i_10_125_466_0, i_10_125_467_0,
    i_10_125_507_0, i_10_125_518_0, i_10_125_628_0, i_10_125_729_0,
    i_10_125_799_0, i_10_125_955_0, i_10_125_956_0, i_10_125_1005_0,
    i_10_125_1034_0, i_10_125_1235_0, i_10_125_1238_0, i_10_125_1241_0,
    i_10_125_1247_0, i_10_125_1305_0, i_10_125_1310_0, i_10_125_1348_0,
    i_10_125_1444_0, i_10_125_1445_0, i_10_125_1653_0, i_10_125_1717_0,
    i_10_125_1718_0, i_10_125_1765_0, i_10_125_1818_0, i_10_125_1821_0,
    i_10_125_1929_0, i_10_125_1948_0, i_10_125_2022_0, i_10_125_2023_0,
    i_10_125_2181_0, i_10_125_2252_0, i_10_125_2254_0, i_10_125_2326_0,
    i_10_125_2356_0, i_10_125_2357_0, i_10_125_2410_0, i_10_125_2456_0,
    i_10_125_2467_0, i_10_125_2469_0, i_10_125_2472_0, i_10_125_2514_0,
    i_10_125_2515_0, i_10_125_2516_0, i_10_125_2519_0, i_10_125_2570_0,
    i_10_125_2631_0, i_10_125_2632_0, i_10_125_2678_0, i_10_125_2681_0,
    i_10_125_2704_0, i_10_125_2705_0, i_10_125_2713_0, i_10_125_2714_0,
    i_10_125_2717_0, i_10_125_2722_0, i_10_125_2760_0, i_10_125_2784_0,
    i_10_125_2788_0, i_10_125_2830_0, i_10_125_2831_0, i_10_125_2832_0,
    i_10_125_2884_0, i_10_125_3072_0, i_10_125_3073_0, i_10_125_3201_0,
    i_10_125_3281_0, i_10_125_3283_0, i_10_125_3386_0, i_10_125_3390_0,
    i_10_125_3391_0, i_10_125_3392_0, i_10_125_3444_0, i_10_125_3500_0,
    i_10_125_3507_0, i_10_125_3586_0, i_10_125_3587_0, i_10_125_3589_0,
    i_10_125_3590_0, i_10_125_3616_0, i_10_125_3617_0, i_10_125_3648_0,
    i_10_125_3781_0, i_10_125_3782_0, i_10_125_3844_0, i_10_125_3845_0,
    i_10_125_3858_0, i_10_125_4115_0, i_10_125_4129_0, i_10_125_4568_0;
  output o_10_125_0_0;
  assign o_10_125_0_0 = 0;
endmodule



// Benchmark "kernel_10_126" written by ABC on Sun Jul 19 10:23:08 2020

module kernel_10_126 ( 
    i_10_126_57_0, i_10_126_171_0, i_10_126_184_0, i_10_126_223_0,
    i_10_126_247_0, i_10_126_271_0, i_10_126_327_0, i_10_126_390_0,
    i_10_126_424_0, i_10_126_436_0, i_10_126_442_0, i_10_126_443_0,
    i_10_126_445_0, i_10_126_463_0, i_10_126_464_0, i_10_126_589_0,
    i_10_126_717_0, i_10_126_993_0, i_10_126_1035_0, i_10_126_1041_0,
    i_10_126_1057_0, i_10_126_1111_0, i_10_126_1207_0, i_10_126_1210_0,
    i_10_126_1246_0, i_10_126_1264_0, i_10_126_1381_0, i_10_126_1399_0,
    i_10_126_1400_0, i_10_126_1453_0, i_10_126_1541_0, i_10_126_1614_0,
    i_10_126_1632_0, i_10_126_1633_0, i_10_126_1650_0, i_10_126_1655_0,
    i_10_126_1688_0, i_10_126_1692_0, i_10_126_1764_0, i_10_126_1765_0,
    i_10_126_1766_0, i_10_126_1794_0, i_10_126_1820_0, i_10_126_1893_0,
    i_10_126_1938_0, i_10_126_1988_0, i_10_126_2031_0, i_10_126_2032_0,
    i_10_126_2068_0, i_10_126_2208_0, i_10_126_2244_0, i_10_126_2259_0,
    i_10_126_2308_0, i_10_126_2309_0, i_10_126_2311_0, i_10_126_2353_0,
    i_10_126_2387_0, i_10_126_2388_0, i_10_126_2452_0, i_10_126_2523_0,
    i_10_126_2559_0, i_10_126_2658_0, i_10_126_2662_0, i_10_126_2676_0,
    i_10_126_2704_0, i_10_126_2820_0, i_10_126_3010_0, i_10_126_3046_0,
    i_10_126_3073_0, i_10_126_3117_0, i_10_126_3209_0, i_10_126_3277_0,
    i_10_126_3327_0, i_10_126_3451_0, i_10_126_3466_0, i_10_126_3494_0,
    i_10_126_3497_0, i_10_126_3526_0, i_10_126_3540_0, i_10_126_3570_0,
    i_10_126_3577_0, i_10_126_3578_0, i_10_126_3616_0, i_10_126_3639_0,
    i_10_126_3688_0, i_10_126_3725_0, i_10_126_3780_0, i_10_126_3787_0,
    i_10_126_3838_0, i_10_126_3855_0, i_10_126_3942_0, i_10_126_3946_0,
    i_10_126_3981_0, i_10_126_4174_0, i_10_126_4192_0, i_10_126_4193_0,
    i_10_126_4263_0, i_10_126_4282_0, i_10_126_4567_0, i_10_126_4574_0,
    o_10_126_0_0  );
  input  i_10_126_57_0, i_10_126_171_0, i_10_126_184_0, i_10_126_223_0,
    i_10_126_247_0, i_10_126_271_0, i_10_126_327_0, i_10_126_390_0,
    i_10_126_424_0, i_10_126_436_0, i_10_126_442_0, i_10_126_443_0,
    i_10_126_445_0, i_10_126_463_0, i_10_126_464_0, i_10_126_589_0,
    i_10_126_717_0, i_10_126_993_0, i_10_126_1035_0, i_10_126_1041_0,
    i_10_126_1057_0, i_10_126_1111_0, i_10_126_1207_0, i_10_126_1210_0,
    i_10_126_1246_0, i_10_126_1264_0, i_10_126_1381_0, i_10_126_1399_0,
    i_10_126_1400_0, i_10_126_1453_0, i_10_126_1541_0, i_10_126_1614_0,
    i_10_126_1632_0, i_10_126_1633_0, i_10_126_1650_0, i_10_126_1655_0,
    i_10_126_1688_0, i_10_126_1692_0, i_10_126_1764_0, i_10_126_1765_0,
    i_10_126_1766_0, i_10_126_1794_0, i_10_126_1820_0, i_10_126_1893_0,
    i_10_126_1938_0, i_10_126_1988_0, i_10_126_2031_0, i_10_126_2032_0,
    i_10_126_2068_0, i_10_126_2208_0, i_10_126_2244_0, i_10_126_2259_0,
    i_10_126_2308_0, i_10_126_2309_0, i_10_126_2311_0, i_10_126_2353_0,
    i_10_126_2387_0, i_10_126_2388_0, i_10_126_2452_0, i_10_126_2523_0,
    i_10_126_2559_0, i_10_126_2658_0, i_10_126_2662_0, i_10_126_2676_0,
    i_10_126_2704_0, i_10_126_2820_0, i_10_126_3010_0, i_10_126_3046_0,
    i_10_126_3073_0, i_10_126_3117_0, i_10_126_3209_0, i_10_126_3277_0,
    i_10_126_3327_0, i_10_126_3451_0, i_10_126_3466_0, i_10_126_3494_0,
    i_10_126_3497_0, i_10_126_3526_0, i_10_126_3540_0, i_10_126_3570_0,
    i_10_126_3577_0, i_10_126_3578_0, i_10_126_3616_0, i_10_126_3639_0,
    i_10_126_3688_0, i_10_126_3725_0, i_10_126_3780_0, i_10_126_3787_0,
    i_10_126_3838_0, i_10_126_3855_0, i_10_126_3942_0, i_10_126_3946_0,
    i_10_126_3981_0, i_10_126_4174_0, i_10_126_4192_0, i_10_126_4193_0,
    i_10_126_4263_0, i_10_126_4282_0, i_10_126_4567_0, i_10_126_4574_0;
  output o_10_126_0_0;
  assign o_10_126_0_0 = 0;
endmodule



// Benchmark "kernel_10_127" written by ABC on Sun Jul 19 10:23:10 2020

module kernel_10_127 ( 
    i_10_127_145_0, i_10_127_146_0, i_10_127_172_0, i_10_127_173_0,
    i_10_127_176_0, i_10_127_217_0, i_10_127_222_0, i_10_127_224_0,
    i_10_127_262_0, i_10_127_284_0, i_10_127_432_0, i_10_127_442_0,
    i_10_127_443_0, i_10_127_444_0, i_10_127_445_0, i_10_127_446_0,
    i_10_127_455_0, i_10_127_461_0, i_10_127_514_0, i_10_127_515_0,
    i_10_127_793_0, i_10_127_794_0, i_10_127_796_0, i_10_127_797_0,
    i_10_127_965_0, i_10_127_967_0, i_10_127_968_0, i_10_127_1085_0,
    i_10_127_1242_0, i_10_127_1305_0, i_10_127_1360_0, i_10_127_1361_0,
    i_10_127_1364_0, i_10_127_1575_0, i_10_127_1576_0, i_10_127_1577_0,
    i_10_127_1631_0, i_10_127_1649_0, i_10_127_1651_0, i_10_127_1652_0,
    i_10_127_1688_0, i_10_127_1819_0, i_10_127_1820_0, i_10_127_1821_0,
    i_10_127_1822_0, i_10_127_1823_0, i_10_127_1824_0, i_10_127_1945_0,
    i_10_127_1999_0, i_10_127_2243_0, i_10_127_2350_0, i_10_127_2355_0,
    i_10_127_2379_0, i_10_127_2380_0, i_10_127_2448_0, i_10_127_2453_0,
    i_10_127_2458_0, i_10_127_2462_0, i_10_127_2503_0, i_10_127_2504_0,
    i_10_127_2629_0, i_10_127_2674_0, i_10_127_2675_0, i_10_127_2681_0,
    i_10_127_2701_0, i_10_127_2718_0, i_10_127_2719_0, i_10_127_2726_0,
    i_10_127_2734_0, i_10_127_2827_0, i_10_127_2828_0, i_10_127_2830_0,
    i_10_127_2908_0, i_10_127_3046_0, i_10_127_3232_0, i_10_127_3233_0,
    i_10_127_3387_0, i_10_127_3389_0, i_10_127_3494_0, i_10_127_3520_0,
    i_10_127_3524_0, i_10_127_3584_0, i_10_127_3587_0, i_10_127_3610_0,
    i_10_127_3613_0, i_10_127_3784_0, i_10_127_3809_0, i_10_127_3839_0,
    i_10_127_3846_0, i_10_127_3853_0, i_10_127_3858_0, i_10_127_3890_0,
    i_10_127_3913_0, i_10_127_3943_0, i_10_127_4130_0, i_10_127_4268_0,
    i_10_127_4287_0, i_10_127_4288_0, i_10_127_4291_0, i_10_127_4565_0,
    o_10_127_0_0  );
  input  i_10_127_145_0, i_10_127_146_0, i_10_127_172_0, i_10_127_173_0,
    i_10_127_176_0, i_10_127_217_0, i_10_127_222_0, i_10_127_224_0,
    i_10_127_262_0, i_10_127_284_0, i_10_127_432_0, i_10_127_442_0,
    i_10_127_443_0, i_10_127_444_0, i_10_127_445_0, i_10_127_446_0,
    i_10_127_455_0, i_10_127_461_0, i_10_127_514_0, i_10_127_515_0,
    i_10_127_793_0, i_10_127_794_0, i_10_127_796_0, i_10_127_797_0,
    i_10_127_965_0, i_10_127_967_0, i_10_127_968_0, i_10_127_1085_0,
    i_10_127_1242_0, i_10_127_1305_0, i_10_127_1360_0, i_10_127_1361_0,
    i_10_127_1364_0, i_10_127_1575_0, i_10_127_1576_0, i_10_127_1577_0,
    i_10_127_1631_0, i_10_127_1649_0, i_10_127_1651_0, i_10_127_1652_0,
    i_10_127_1688_0, i_10_127_1819_0, i_10_127_1820_0, i_10_127_1821_0,
    i_10_127_1822_0, i_10_127_1823_0, i_10_127_1824_0, i_10_127_1945_0,
    i_10_127_1999_0, i_10_127_2243_0, i_10_127_2350_0, i_10_127_2355_0,
    i_10_127_2379_0, i_10_127_2380_0, i_10_127_2448_0, i_10_127_2453_0,
    i_10_127_2458_0, i_10_127_2462_0, i_10_127_2503_0, i_10_127_2504_0,
    i_10_127_2629_0, i_10_127_2674_0, i_10_127_2675_0, i_10_127_2681_0,
    i_10_127_2701_0, i_10_127_2718_0, i_10_127_2719_0, i_10_127_2726_0,
    i_10_127_2734_0, i_10_127_2827_0, i_10_127_2828_0, i_10_127_2830_0,
    i_10_127_2908_0, i_10_127_3046_0, i_10_127_3232_0, i_10_127_3233_0,
    i_10_127_3387_0, i_10_127_3389_0, i_10_127_3494_0, i_10_127_3520_0,
    i_10_127_3524_0, i_10_127_3584_0, i_10_127_3587_0, i_10_127_3610_0,
    i_10_127_3613_0, i_10_127_3784_0, i_10_127_3809_0, i_10_127_3839_0,
    i_10_127_3846_0, i_10_127_3853_0, i_10_127_3858_0, i_10_127_3890_0,
    i_10_127_3913_0, i_10_127_3943_0, i_10_127_4130_0, i_10_127_4268_0,
    i_10_127_4287_0, i_10_127_4288_0, i_10_127_4291_0, i_10_127_4565_0;
  output o_10_127_0_0;
  assign o_10_127_0_0 = ~((~i_10_127_4130_0 & ((~i_10_127_172_0 & ((~i_10_127_514_0 & ~i_10_127_796_0 & ~i_10_127_1823_0 & ~i_10_127_2674_0 & ~i_10_127_3232_0 & ~i_10_127_3524_0) | (~i_10_127_443_0 & ~i_10_127_444_0 & ~i_10_127_1360_0 & ~i_10_127_1824_0 & ~i_10_127_2350_0 & ~i_10_127_3046_0 & ~i_10_127_3913_0))) | (i_10_127_172_0 & ~i_10_127_444_0 & ~i_10_127_515_0 & ~i_10_127_2718_0 & ~i_10_127_3232_0 & ~i_10_127_3610_0) | (~i_10_127_446_0 & i_10_127_2734_0 & i_10_127_3839_0))) | (~i_10_127_173_0 & ((~i_10_127_146_0 & ~i_10_127_445_0 & ~i_10_127_1361_0 & ~i_10_127_2380_0 & ~i_10_127_2681_0 & ~i_10_127_3232_0) | (~i_10_127_145_0 & ~i_10_127_1649_0 & ~i_10_127_1823_0 & ~i_10_127_2504_0 & ~i_10_127_2718_0 & ~i_10_127_3494_0 & ~i_10_127_3839_0 & ~i_10_127_3890_0 & ~i_10_127_3913_0 & ~i_10_127_3943_0))) | (~i_10_127_145_0 & ((i_10_127_444_0 & ~i_10_127_1577_0 & ~i_10_127_2504_0 & ~i_10_127_3233_0 & i_10_127_3853_0) | (~i_10_127_224_0 & ~i_10_127_455_0 & ~i_10_127_965_0 & ~i_10_127_1085_0 & ~i_10_127_1360_0 & ~i_10_127_1649_0 & ~i_10_127_2448_0 & ~i_10_127_2734_0 & ~i_10_127_3494_0 & ~i_10_127_3524_0 & ~i_10_127_3784_0 & ~i_10_127_3890_0 & ~i_10_127_3913_0))) | (~i_10_127_968_0 & ((~i_10_127_146_0 & ((~i_10_127_796_0 & ~i_10_127_1652_0 & ~i_10_127_1820_0 & ~i_10_127_3524_0 & ~i_10_127_3784_0 & ~i_10_127_2675_0 & ~i_10_127_3387_0) | (~i_10_127_1242_0 & ~i_10_127_1361_0 & ~i_10_127_2380_0 & ~i_10_127_2453_0 & ~i_10_127_2462_0 & ~i_10_127_3232_0 & ~i_10_127_3233_0 & ~i_10_127_3613_0 & ~i_10_127_3858_0))) | (~i_10_127_1651_0 & ~i_10_127_1652_0 & ~i_10_127_2503_0 & ~i_10_127_2681_0 & ~i_10_127_3233_0 & ~i_10_127_3587_0) | (~i_10_127_797_0 & ~i_10_127_1361_0 & i_10_127_1819_0 & ~i_10_127_2675_0 & ~i_10_127_3839_0))) | (~i_10_127_176_0 & ~i_10_127_1364_0 & ((~i_10_127_514_0 & ~i_10_127_515_0 & ~i_10_127_2462_0 & ~i_10_127_2503_0 & ~i_10_127_3233_0 & i_10_127_3610_0 & ~i_10_127_3890_0 & ~i_10_127_4268_0) | (~i_10_127_461_0 & ~i_10_127_967_0 & ~i_10_127_1688_0 & ~i_10_127_3494_0 & ~i_10_127_4565_0))) | (~i_10_127_3233_0 & ((~i_10_127_446_0 & ((i_10_127_284_0 & ~i_10_127_793_0 & i_10_127_1305_0 & i_10_127_1823_0) | (~i_10_127_796_0 & ~i_10_127_1360_0 & i_10_127_1820_0 & ~i_10_127_3913_0))) | (~i_10_127_965_0 & ~i_10_127_1819_0 & ~i_10_127_1823_0 & ~i_10_127_2503_0 & ~i_10_127_2504_0 & ~i_10_127_3839_0 & ~i_10_127_3943_0 & ~i_10_127_4268_0 & ~i_10_127_4291_0))) | (~i_10_127_794_0 & ((i_10_127_432_0 & i_10_127_1820_0) | (~i_10_127_3046_0 & ~i_10_127_3913_0 & ~i_10_127_2453_0 & i_10_127_2681_0))) | (~i_10_127_1688_0 & ((~i_10_127_443_0 & ~i_10_127_1822_0 & ~i_10_127_3520_0) | (~i_10_127_793_0 & i_10_127_2830_0 & ~i_10_127_3839_0))) | (~i_10_127_3232_0 & ((~i_10_127_444_0 & ~i_10_127_797_0 & ~i_10_127_965_0 & ~i_10_127_2453_0 & ~i_10_127_2629_0) | (~i_10_127_514_0 & ~i_10_127_2674_0 & ~i_10_127_2726_0 & i_10_127_2828_0))) | (~i_10_127_797_0 & ((~i_10_127_2719_0 & ~i_10_127_2734_0 & i_10_127_3784_0) | (i_10_127_1824_0 & ~i_10_127_3858_0) | (~i_10_127_445_0 & ~i_10_127_796_0 & i_10_127_3613_0 & i_10_127_4130_0))) | (~i_10_127_461_0 & i_10_127_514_0 & i_10_127_1576_0) | (i_10_127_262_0 & ~i_10_127_1999_0 & i_10_127_3610_0 & i_10_127_3858_0));
endmodule



// Benchmark "kernel_10_128" written by ABC on Sun Jul 19 10:23:11 2020

module kernel_10_128 ( 
    i_10_128_244_0, i_10_128_281_0, i_10_128_282_0, i_10_128_284_0,
    i_10_128_288_0, i_10_128_289_0, i_10_128_315_0, i_10_128_319_0,
    i_10_128_412_0, i_10_128_435_0, i_10_128_449_0, i_10_128_461_0,
    i_10_128_462_0, i_10_128_464_0, i_10_128_467_0, i_10_128_500_0,
    i_10_128_735_0, i_10_128_792_0, i_10_128_797_0, i_10_128_1118_0,
    i_10_128_1234_0, i_10_128_1235_0, i_10_128_1238_0, i_10_128_1243_0,
    i_10_128_1244_0, i_10_128_1245_0, i_10_128_1273_0, i_10_128_1307_0,
    i_10_128_1361_0, i_10_128_1451_0, i_10_128_1583_0, i_10_128_1651_0,
    i_10_128_1652_0, i_10_128_1687_0, i_10_128_1688_0, i_10_128_1818_0,
    i_10_128_1819_0, i_10_128_1820_0, i_10_128_1822_0, i_10_128_1910_0,
    i_10_128_1945_0, i_10_128_1946_0, i_10_128_1949_0, i_10_128_1951_0,
    i_10_128_1989_0, i_10_128_1990_0, i_10_128_2178_0, i_10_128_2333_0,
    i_10_128_2352_0, i_10_128_2353_0, i_10_128_2356_0, i_10_128_2364_0,
    i_10_128_2376_0, i_10_128_2407_0, i_10_128_2408_0, i_10_128_2441_0,
    i_10_128_2454_0, i_10_128_2455_0, i_10_128_2459_0, i_10_128_2470_0,
    i_10_128_2673_0, i_10_128_2679_0, i_10_128_2700_0, i_10_128_2704_0,
    i_10_128_2709_0, i_10_128_2882_0, i_10_128_2918_0, i_10_128_2921_0,
    i_10_128_2924_0, i_10_128_3267_0, i_10_128_3268_0, i_10_128_3269_0,
    i_10_128_3276_0, i_10_128_3277_0, i_10_128_3278_0, i_10_128_3280_0,
    i_10_128_3281_0, i_10_128_3384_0, i_10_128_3386_0, i_10_128_3406_0,
    i_10_128_3497_0, i_10_128_3586_0, i_10_128_3615_0, i_10_128_3645_0,
    i_10_128_3682_0, i_10_128_3728_0, i_10_128_3784_0, i_10_128_3839_0,
    i_10_128_3846_0, i_10_128_3858_0, i_10_128_3859_0, i_10_128_3894_0,
    i_10_128_3895_0, i_10_128_3984_0, i_10_128_4054_0, i_10_128_4116_0,
    i_10_128_4117_0, i_10_128_4119_0, i_10_128_4457_0, i_10_128_4568_0,
    o_10_128_0_0  );
  input  i_10_128_244_0, i_10_128_281_0, i_10_128_282_0, i_10_128_284_0,
    i_10_128_288_0, i_10_128_289_0, i_10_128_315_0, i_10_128_319_0,
    i_10_128_412_0, i_10_128_435_0, i_10_128_449_0, i_10_128_461_0,
    i_10_128_462_0, i_10_128_464_0, i_10_128_467_0, i_10_128_500_0,
    i_10_128_735_0, i_10_128_792_0, i_10_128_797_0, i_10_128_1118_0,
    i_10_128_1234_0, i_10_128_1235_0, i_10_128_1238_0, i_10_128_1243_0,
    i_10_128_1244_0, i_10_128_1245_0, i_10_128_1273_0, i_10_128_1307_0,
    i_10_128_1361_0, i_10_128_1451_0, i_10_128_1583_0, i_10_128_1651_0,
    i_10_128_1652_0, i_10_128_1687_0, i_10_128_1688_0, i_10_128_1818_0,
    i_10_128_1819_0, i_10_128_1820_0, i_10_128_1822_0, i_10_128_1910_0,
    i_10_128_1945_0, i_10_128_1946_0, i_10_128_1949_0, i_10_128_1951_0,
    i_10_128_1989_0, i_10_128_1990_0, i_10_128_2178_0, i_10_128_2333_0,
    i_10_128_2352_0, i_10_128_2353_0, i_10_128_2356_0, i_10_128_2364_0,
    i_10_128_2376_0, i_10_128_2407_0, i_10_128_2408_0, i_10_128_2441_0,
    i_10_128_2454_0, i_10_128_2455_0, i_10_128_2459_0, i_10_128_2470_0,
    i_10_128_2673_0, i_10_128_2679_0, i_10_128_2700_0, i_10_128_2704_0,
    i_10_128_2709_0, i_10_128_2882_0, i_10_128_2918_0, i_10_128_2921_0,
    i_10_128_2924_0, i_10_128_3267_0, i_10_128_3268_0, i_10_128_3269_0,
    i_10_128_3276_0, i_10_128_3277_0, i_10_128_3278_0, i_10_128_3280_0,
    i_10_128_3281_0, i_10_128_3384_0, i_10_128_3386_0, i_10_128_3406_0,
    i_10_128_3497_0, i_10_128_3586_0, i_10_128_3615_0, i_10_128_3645_0,
    i_10_128_3682_0, i_10_128_3728_0, i_10_128_3784_0, i_10_128_3839_0,
    i_10_128_3846_0, i_10_128_3858_0, i_10_128_3859_0, i_10_128_3894_0,
    i_10_128_3895_0, i_10_128_3984_0, i_10_128_4054_0, i_10_128_4116_0,
    i_10_128_4117_0, i_10_128_4119_0, i_10_128_4457_0, i_10_128_4568_0;
  output o_10_128_0_0;
  assign o_10_128_0_0 = 0;
endmodule



// Benchmark "kernel_10_129" written by ABC on Sun Jul 19 10:23:11 2020

module kernel_10_129 ( 
    i_10_129_51_0, i_10_129_52_0, i_10_129_153_0, i_10_129_156_0,
    i_10_129_181_0, i_10_129_237_0, i_10_129_251_0, i_10_129_283_0,
    i_10_129_293_0, i_10_129_327_0, i_10_129_354_0, i_10_129_355_0,
    i_10_129_357_0, i_10_129_589_0, i_10_129_633_0, i_10_129_636_0,
    i_10_129_687_0, i_10_129_688_0, i_10_129_732_0, i_10_129_828_0,
    i_10_129_930_0, i_10_129_993_0, i_10_129_1135_0, i_10_129_1161_0,
    i_10_129_1209_0, i_10_129_1234_0, i_10_129_1290_0, i_10_129_1306_0,
    i_10_129_1380_0, i_10_129_1530_0, i_10_129_1531_0, i_10_129_1533_0,
    i_10_129_1534_0, i_10_129_1543_0, i_10_129_1560_0, i_10_129_1561_0,
    i_10_129_1632_0, i_10_129_1651_0, i_10_129_1686_0, i_10_129_1791_0,
    i_10_129_1800_0, i_10_129_1801_0, i_10_129_1848_0, i_10_129_1912_0,
    i_10_129_1918_0, i_10_129_2163_0, i_10_129_2200_0, i_10_129_2253_0,
    i_10_129_2256_0, i_10_129_2442_0, i_10_129_2450_0, i_10_129_2529_0,
    i_10_129_2604_0, i_10_129_2632_0, i_10_129_2674_0, i_10_129_2713_0,
    i_10_129_2715_0, i_10_129_2716_0, i_10_129_2724_0, i_10_129_2775_0,
    i_10_129_2832_0, i_10_129_2979_0, i_10_129_2982_0, i_10_129_3096_0,
    i_10_129_3099_0, i_10_129_3196_0, i_10_129_3198_0, i_10_129_3199_0,
    i_10_129_3280_0, i_10_129_3282_0, i_10_129_3289_0, i_10_129_3291_0,
    i_10_129_3315_0, i_10_129_3325_0, i_10_129_3387_0, i_10_129_3388_0,
    i_10_129_3390_0, i_10_129_3391_0, i_10_129_3465_0, i_10_129_3564_0,
    i_10_129_3577_0, i_10_129_3609_0, i_10_129_3610_0, i_10_129_3645_0,
    i_10_129_3646_0, i_10_129_3648_0, i_10_129_3702_0, i_10_129_3703_0,
    i_10_129_3774_0, i_10_129_3780_0, i_10_129_3783_0, i_10_129_3786_0,
    i_10_129_3857_0, i_10_129_3870_0, i_10_129_3873_0, i_10_129_3996_0,
    i_10_129_4131_0, i_10_129_4226_0, i_10_129_4461_0, i_10_129_4582_0,
    o_10_129_0_0  );
  input  i_10_129_51_0, i_10_129_52_0, i_10_129_153_0, i_10_129_156_0,
    i_10_129_181_0, i_10_129_237_0, i_10_129_251_0, i_10_129_283_0,
    i_10_129_293_0, i_10_129_327_0, i_10_129_354_0, i_10_129_355_0,
    i_10_129_357_0, i_10_129_589_0, i_10_129_633_0, i_10_129_636_0,
    i_10_129_687_0, i_10_129_688_0, i_10_129_732_0, i_10_129_828_0,
    i_10_129_930_0, i_10_129_993_0, i_10_129_1135_0, i_10_129_1161_0,
    i_10_129_1209_0, i_10_129_1234_0, i_10_129_1290_0, i_10_129_1306_0,
    i_10_129_1380_0, i_10_129_1530_0, i_10_129_1531_0, i_10_129_1533_0,
    i_10_129_1534_0, i_10_129_1543_0, i_10_129_1560_0, i_10_129_1561_0,
    i_10_129_1632_0, i_10_129_1651_0, i_10_129_1686_0, i_10_129_1791_0,
    i_10_129_1800_0, i_10_129_1801_0, i_10_129_1848_0, i_10_129_1912_0,
    i_10_129_1918_0, i_10_129_2163_0, i_10_129_2200_0, i_10_129_2253_0,
    i_10_129_2256_0, i_10_129_2442_0, i_10_129_2450_0, i_10_129_2529_0,
    i_10_129_2604_0, i_10_129_2632_0, i_10_129_2674_0, i_10_129_2713_0,
    i_10_129_2715_0, i_10_129_2716_0, i_10_129_2724_0, i_10_129_2775_0,
    i_10_129_2832_0, i_10_129_2979_0, i_10_129_2982_0, i_10_129_3096_0,
    i_10_129_3099_0, i_10_129_3196_0, i_10_129_3198_0, i_10_129_3199_0,
    i_10_129_3280_0, i_10_129_3282_0, i_10_129_3289_0, i_10_129_3291_0,
    i_10_129_3315_0, i_10_129_3325_0, i_10_129_3387_0, i_10_129_3388_0,
    i_10_129_3390_0, i_10_129_3391_0, i_10_129_3465_0, i_10_129_3564_0,
    i_10_129_3577_0, i_10_129_3609_0, i_10_129_3610_0, i_10_129_3645_0,
    i_10_129_3646_0, i_10_129_3648_0, i_10_129_3702_0, i_10_129_3703_0,
    i_10_129_3774_0, i_10_129_3780_0, i_10_129_3783_0, i_10_129_3786_0,
    i_10_129_3857_0, i_10_129_3870_0, i_10_129_3873_0, i_10_129_3996_0,
    i_10_129_4131_0, i_10_129_4226_0, i_10_129_4461_0, i_10_129_4582_0;
  output o_10_129_0_0;
  assign o_10_129_0_0 = 0;
endmodule



// Benchmark "kernel_10_130" written by ABC on Sun Jul 19 10:23:12 2020

module kernel_10_130 ( 
    i_10_130_51_0, i_10_130_293_0, i_10_130_391_0, i_10_130_427_0,
    i_10_130_428_0, i_10_130_433_0, i_10_130_447_0, i_10_130_449_0,
    i_10_130_465_0, i_10_130_613_0, i_10_130_714_0, i_10_130_750_0,
    i_10_130_893_0, i_10_130_984_0, i_10_130_993_0, i_10_130_1012_0,
    i_10_130_1029_0, i_10_130_1034_0, i_10_130_1170_0, i_10_130_1171_0,
    i_10_130_1239_0, i_10_130_1242_0, i_10_130_1244_0, i_10_130_1245_0,
    i_10_130_1246_0, i_10_130_1247_0, i_10_130_1248_0, i_10_130_1249_0,
    i_10_130_1445_0, i_10_130_1447_0, i_10_130_1542_0, i_10_130_1632_0,
    i_10_130_1650_0, i_10_130_1653_0, i_10_130_1654_0, i_10_130_1756_0,
    i_10_130_1758_0, i_10_130_1759_0, i_10_130_1819_0, i_10_130_1823_0,
    i_10_130_2012_0, i_10_130_2181_0, i_10_130_2203_0, i_10_130_2207_0,
    i_10_130_2225_0, i_10_130_2307_0, i_10_130_2362_0, i_10_130_2454_0,
    i_10_130_2470_0, i_10_130_2471_0, i_10_130_2473_0, i_10_130_2532_0,
    i_10_130_2628_0, i_10_130_2655_0, i_10_130_2660_0, i_10_130_2686_0,
    i_10_130_2916_0, i_10_130_3033_0, i_10_130_3034_0, i_10_130_3037_0,
    i_10_130_3041_0, i_10_130_3166_0, i_10_130_3169_0, i_10_130_3172_0,
    i_10_130_3307_0, i_10_130_3334_0, i_10_130_3386_0, i_10_130_3429_0,
    i_10_130_3469_0, i_10_130_3586_0, i_10_130_3590_0, i_10_130_3617_0,
    i_10_130_3684_0, i_10_130_3685_0, i_10_130_3687_0, i_10_130_3688_0,
    i_10_130_3717_0, i_10_130_3729_0, i_10_130_3780_0, i_10_130_3784_0,
    i_10_130_3786_0, i_10_130_3829_0, i_10_130_3844_0, i_10_130_4008_0,
    i_10_130_4011_0, i_10_130_4066_0, i_10_130_4117_0, i_10_130_4118_0,
    i_10_130_4174_0, i_10_130_4175_0, i_10_130_4188_0, i_10_130_4219_0,
    i_10_130_4260_0, i_10_130_4261_0, i_10_130_4269_0, i_10_130_4276_0,
    i_10_130_4287_0, i_10_130_4477_0, i_10_130_4569_0, i_10_130_4597_0,
    o_10_130_0_0  );
  input  i_10_130_51_0, i_10_130_293_0, i_10_130_391_0, i_10_130_427_0,
    i_10_130_428_0, i_10_130_433_0, i_10_130_447_0, i_10_130_449_0,
    i_10_130_465_0, i_10_130_613_0, i_10_130_714_0, i_10_130_750_0,
    i_10_130_893_0, i_10_130_984_0, i_10_130_993_0, i_10_130_1012_0,
    i_10_130_1029_0, i_10_130_1034_0, i_10_130_1170_0, i_10_130_1171_0,
    i_10_130_1239_0, i_10_130_1242_0, i_10_130_1244_0, i_10_130_1245_0,
    i_10_130_1246_0, i_10_130_1247_0, i_10_130_1248_0, i_10_130_1249_0,
    i_10_130_1445_0, i_10_130_1447_0, i_10_130_1542_0, i_10_130_1632_0,
    i_10_130_1650_0, i_10_130_1653_0, i_10_130_1654_0, i_10_130_1756_0,
    i_10_130_1758_0, i_10_130_1759_0, i_10_130_1819_0, i_10_130_1823_0,
    i_10_130_2012_0, i_10_130_2181_0, i_10_130_2203_0, i_10_130_2207_0,
    i_10_130_2225_0, i_10_130_2307_0, i_10_130_2362_0, i_10_130_2454_0,
    i_10_130_2470_0, i_10_130_2471_0, i_10_130_2473_0, i_10_130_2532_0,
    i_10_130_2628_0, i_10_130_2655_0, i_10_130_2660_0, i_10_130_2686_0,
    i_10_130_2916_0, i_10_130_3033_0, i_10_130_3034_0, i_10_130_3037_0,
    i_10_130_3041_0, i_10_130_3166_0, i_10_130_3169_0, i_10_130_3172_0,
    i_10_130_3307_0, i_10_130_3334_0, i_10_130_3386_0, i_10_130_3429_0,
    i_10_130_3469_0, i_10_130_3586_0, i_10_130_3590_0, i_10_130_3617_0,
    i_10_130_3684_0, i_10_130_3685_0, i_10_130_3687_0, i_10_130_3688_0,
    i_10_130_3717_0, i_10_130_3729_0, i_10_130_3780_0, i_10_130_3784_0,
    i_10_130_3786_0, i_10_130_3829_0, i_10_130_3844_0, i_10_130_4008_0,
    i_10_130_4011_0, i_10_130_4066_0, i_10_130_4117_0, i_10_130_4118_0,
    i_10_130_4174_0, i_10_130_4175_0, i_10_130_4188_0, i_10_130_4219_0,
    i_10_130_4260_0, i_10_130_4261_0, i_10_130_4269_0, i_10_130_4276_0,
    i_10_130_4287_0, i_10_130_4477_0, i_10_130_4569_0, i_10_130_4597_0;
  output o_10_130_0_0;
  assign o_10_130_0_0 = 0;
endmodule



// Benchmark "kernel_10_131" written by ABC on Sun Jul 19 10:23:13 2020

module kernel_10_131 ( 
    i_10_131_48_0, i_10_131_118_0, i_10_131_136_0, i_10_131_171_0,
    i_10_131_182_0, i_10_131_246_0, i_10_131_282_0, i_10_131_283_0,
    i_10_131_285_0, i_10_131_286_0, i_10_131_291_0, i_10_131_292_0,
    i_10_131_293_0, i_10_131_315_0, i_10_131_330_0, i_10_131_390_0,
    i_10_131_391_0, i_10_131_407_0, i_10_131_409_0, i_10_131_410_0,
    i_10_131_448_0, i_10_131_625_0, i_10_131_634_0, i_10_131_689_0,
    i_10_131_792_0, i_10_131_826_0, i_10_131_957_0, i_10_131_963_0,
    i_10_131_967_0, i_10_131_993_0, i_10_131_1051_0, i_10_131_1052_0,
    i_10_131_1163_0, i_10_131_1266_0, i_10_131_1267_0, i_10_131_1302_0,
    i_10_131_1306_0, i_10_131_1435_0, i_10_131_1444_0, i_10_131_1488_0,
    i_10_131_1579_0, i_10_131_1581_0, i_10_131_1618_0, i_10_131_1649_0,
    i_10_131_1653_0, i_10_131_1683_0, i_10_131_1684_0, i_10_131_1800_0,
    i_10_131_2004_0, i_10_131_2025_0, i_10_131_2082_0, i_10_131_2202_0,
    i_10_131_2203_0, i_10_131_2353_0, i_10_131_2355_0, i_10_131_2361_0,
    i_10_131_2377_0, i_10_131_2455_0, i_10_131_2475_0, i_10_131_2541_0,
    i_10_131_2566_0, i_10_131_2572_0, i_10_131_2605_0, i_10_131_2607_0,
    i_10_131_2608_0, i_10_131_2611_0, i_10_131_2634_0, i_10_131_2677_0,
    i_10_131_2679_0, i_10_131_2709_0, i_10_131_2712_0, i_10_131_2718_0,
    i_10_131_2719_0, i_10_131_2725_0, i_10_131_2734_0, i_10_131_2782_0,
    i_10_131_2985_0, i_10_131_3198_0, i_10_131_3199_0, i_10_131_3235_0,
    i_10_131_3282_0, i_10_131_3288_0, i_10_131_3387_0, i_10_131_3388_0,
    i_10_131_3433_0, i_10_131_3471_0, i_10_131_3585_0, i_10_131_3609_0,
    i_10_131_3647_0, i_10_131_3721_0, i_10_131_3859_0, i_10_131_3860_0,
    i_10_131_4030_0, i_10_131_4113_0, i_10_131_4116_0, i_10_131_4275_0,
    i_10_131_4276_0, i_10_131_4280_0, i_10_131_4459_0, i_10_131_4566_0,
    o_10_131_0_0  );
  input  i_10_131_48_0, i_10_131_118_0, i_10_131_136_0, i_10_131_171_0,
    i_10_131_182_0, i_10_131_246_0, i_10_131_282_0, i_10_131_283_0,
    i_10_131_285_0, i_10_131_286_0, i_10_131_291_0, i_10_131_292_0,
    i_10_131_293_0, i_10_131_315_0, i_10_131_330_0, i_10_131_390_0,
    i_10_131_391_0, i_10_131_407_0, i_10_131_409_0, i_10_131_410_0,
    i_10_131_448_0, i_10_131_625_0, i_10_131_634_0, i_10_131_689_0,
    i_10_131_792_0, i_10_131_826_0, i_10_131_957_0, i_10_131_963_0,
    i_10_131_967_0, i_10_131_993_0, i_10_131_1051_0, i_10_131_1052_0,
    i_10_131_1163_0, i_10_131_1266_0, i_10_131_1267_0, i_10_131_1302_0,
    i_10_131_1306_0, i_10_131_1435_0, i_10_131_1444_0, i_10_131_1488_0,
    i_10_131_1579_0, i_10_131_1581_0, i_10_131_1618_0, i_10_131_1649_0,
    i_10_131_1653_0, i_10_131_1683_0, i_10_131_1684_0, i_10_131_1800_0,
    i_10_131_2004_0, i_10_131_2025_0, i_10_131_2082_0, i_10_131_2202_0,
    i_10_131_2203_0, i_10_131_2353_0, i_10_131_2355_0, i_10_131_2361_0,
    i_10_131_2377_0, i_10_131_2455_0, i_10_131_2475_0, i_10_131_2541_0,
    i_10_131_2566_0, i_10_131_2572_0, i_10_131_2605_0, i_10_131_2607_0,
    i_10_131_2608_0, i_10_131_2611_0, i_10_131_2634_0, i_10_131_2677_0,
    i_10_131_2679_0, i_10_131_2709_0, i_10_131_2712_0, i_10_131_2718_0,
    i_10_131_2719_0, i_10_131_2725_0, i_10_131_2734_0, i_10_131_2782_0,
    i_10_131_2985_0, i_10_131_3198_0, i_10_131_3199_0, i_10_131_3235_0,
    i_10_131_3282_0, i_10_131_3288_0, i_10_131_3387_0, i_10_131_3388_0,
    i_10_131_3433_0, i_10_131_3471_0, i_10_131_3585_0, i_10_131_3609_0,
    i_10_131_3647_0, i_10_131_3721_0, i_10_131_3859_0, i_10_131_3860_0,
    i_10_131_4030_0, i_10_131_4113_0, i_10_131_4116_0, i_10_131_4275_0,
    i_10_131_4276_0, i_10_131_4280_0, i_10_131_4459_0, i_10_131_4566_0;
  output o_10_131_0_0;
  assign o_10_131_0_0 = 0;
endmodule



// Benchmark "kernel_10_132" written by ABC on Sun Jul 19 10:23:14 2020

module kernel_10_132 ( 
    i_10_132_222_0, i_10_132_223_0, i_10_132_224_0, i_10_132_271_0,
    i_10_132_327_0, i_10_132_328_0, i_10_132_332_0, i_10_132_407_0,
    i_10_132_430_0, i_10_132_433_0, i_10_132_435_0, i_10_132_438_0,
    i_10_132_439_0, i_10_132_507_0, i_10_132_699_0, i_10_132_955_0,
    i_10_132_996_0, i_10_132_997_0, i_10_132_1001_0, i_10_132_1005_0,
    i_10_132_1138_0, i_10_132_1237_0, i_10_132_1238_0, i_10_132_1246_0,
    i_10_132_1247_0, i_10_132_1249_0, i_10_132_1264_0, i_10_132_1307_0,
    i_10_132_1309_0, i_10_132_1310_0, i_10_132_1312_0, i_10_132_1438_0,
    i_10_132_1554_0, i_10_132_1654_0, i_10_132_1688_0, i_10_132_1818_0,
    i_10_132_2020_0, i_10_132_2158_0, i_10_132_2407_0, i_10_132_2508_0,
    i_10_132_2509_0, i_10_132_2629_0, i_10_132_2630_0, i_10_132_2634_0,
    i_10_132_2635_0, i_10_132_2657_0, i_10_132_2661_0, i_10_132_2679_0,
    i_10_132_2680_0, i_10_132_2681_0, i_10_132_2720_0, i_10_132_2724_0,
    i_10_132_2783_0, i_10_132_2820_0, i_10_132_2823_0, i_10_132_2826_0,
    i_10_132_2827_0, i_10_132_2828_0, i_10_132_2831_0, i_10_132_2881_0,
    i_10_132_2882_0, i_10_132_2980_0, i_10_132_2982_0, i_10_132_2985_0,
    i_10_132_3041_0, i_10_132_3072_0, i_10_132_3199_0, i_10_132_3271_0,
    i_10_132_3328_0, i_10_132_3387_0, i_10_132_3388_0, i_10_132_3390_0,
    i_10_132_3391_0, i_10_132_3408_0, i_10_132_3496_0, i_10_132_3614_0,
    i_10_132_3646_0, i_10_132_3648_0, i_10_132_3652_0, i_10_132_3682_0,
    i_10_132_3729_0, i_10_132_3780_0, i_10_132_3781_0, i_10_132_3846_0,
    i_10_132_3848_0, i_10_132_3850_0, i_10_132_3852_0, i_10_132_3853_0,
    i_10_132_3855_0, i_10_132_3859_0, i_10_132_3981_0, i_10_132_3982_0,
    i_10_132_3984_0, i_10_132_3985_0, i_10_132_3986_0, i_10_132_4056_0,
    i_10_132_4129_0, i_10_132_4238_0, i_10_132_4288_0, i_10_132_4289_0,
    o_10_132_0_0  );
  input  i_10_132_222_0, i_10_132_223_0, i_10_132_224_0, i_10_132_271_0,
    i_10_132_327_0, i_10_132_328_0, i_10_132_332_0, i_10_132_407_0,
    i_10_132_430_0, i_10_132_433_0, i_10_132_435_0, i_10_132_438_0,
    i_10_132_439_0, i_10_132_507_0, i_10_132_699_0, i_10_132_955_0,
    i_10_132_996_0, i_10_132_997_0, i_10_132_1001_0, i_10_132_1005_0,
    i_10_132_1138_0, i_10_132_1237_0, i_10_132_1238_0, i_10_132_1246_0,
    i_10_132_1247_0, i_10_132_1249_0, i_10_132_1264_0, i_10_132_1307_0,
    i_10_132_1309_0, i_10_132_1310_0, i_10_132_1312_0, i_10_132_1438_0,
    i_10_132_1554_0, i_10_132_1654_0, i_10_132_1688_0, i_10_132_1818_0,
    i_10_132_2020_0, i_10_132_2158_0, i_10_132_2407_0, i_10_132_2508_0,
    i_10_132_2509_0, i_10_132_2629_0, i_10_132_2630_0, i_10_132_2634_0,
    i_10_132_2635_0, i_10_132_2657_0, i_10_132_2661_0, i_10_132_2679_0,
    i_10_132_2680_0, i_10_132_2681_0, i_10_132_2720_0, i_10_132_2724_0,
    i_10_132_2783_0, i_10_132_2820_0, i_10_132_2823_0, i_10_132_2826_0,
    i_10_132_2827_0, i_10_132_2828_0, i_10_132_2831_0, i_10_132_2881_0,
    i_10_132_2882_0, i_10_132_2980_0, i_10_132_2982_0, i_10_132_2985_0,
    i_10_132_3041_0, i_10_132_3072_0, i_10_132_3199_0, i_10_132_3271_0,
    i_10_132_3328_0, i_10_132_3387_0, i_10_132_3388_0, i_10_132_3390_0,
    i_10_132_3391_0, i_10_132_3408_0, i_10_132_3496_0, i_10_132_3614_0,
    i_10_132_3646_0, i_10_132_3648_0, i_10_132_3652_0, i_10_132_3682_0,
    i_10_132_3729_0, i_10_132_3780_0, i_10_132_3781_0, i_10_132_3846_0,
    i_10_132_3848_0, i_10_132_3850_0, i_10_132_3852_0, i_10_132_3853_0,
    i_10_132_3855_0, i_10_132_3859_0, i_10_132_3981_0, i_10_132_3982_0,
    i_10_132_3984_0, i_10_132_3985_0, i_10_132_3986_0, i_10_132_4056_0,
    i_10_132_4129_0, i_10_132_4238_0, i_10_132_4288_0, i_10_132_4289_0;
  output o_10_132_0_0;
  assign o_10_132_0_0 = ~((~i_10_132_332_0 & ((~i_10_132_328_0 & ((~i_10_132_438_0 & ~i_10_132_2679_0 & ~i_10_132_3496_0 & ~i_10_132_3781_0) | (~i_10_132_1264_0 & ~i_10_132_2407_0 & ~i_10_132_2982_0 & ~i_10_132_2985_0 & ~i_10_132_3984_0))) | (~i_10_132_996_0 & ~i_10_132_2657_0 & ~i_10_132_2679_0 & ~i_10_132_2820_0 & ~i_10_132_3982_0 & ~i_10_132_4238_0))) | (~i_10_132_2508_0 & ((~i_10_132_433_0 & ((~i_10_132_407_0 & ~i_10_132_1001_0 & ~i_10_132_2679_0 & ~i_10_132_2823_0 & ~i_10_132_2982_0 & ~i_10_132_3496_0) | (~i_10_132_435_0 & ~i_10_132_997_0 & ~i_10_132_1438_0 & ~i_10_132_3614_0 & ~i_10_132_3981_0 & ~i_10_132_4129_0 & ~i_10_132_4238_0))) | (~i_10_132_327_0 & ~i_10_132_996_0 & ~i_10_132_2657_0 & ~i_10_132_2680_0 & ~i_10_132_2724_0 & ~i_10_132_2827_0 & ~i_10_132_4129_0) | (~i_10_132_1264_0 & ~i_10_132_1654_0 & ~i_10_132_2985_0 & ~i_10_132_3984_0 & ~i_10_132_3985_0))) | (~i_10_132_2982_0 & ((~i_10_132_327_0 & ((~i_10_132_224_0 & ~i_10_132_1654_0 & ~i_10_132_2629_0 & ~i_10_132_2634_0 & ~i_10_132_2831_0) | (~i_10_132_1264_0 & ~i_10_132_2509_0 & ~i_10_132_2661_0 & ~i_10_132_3985_0))) | (~i_10_132_996_0 & i_10_132_2657_0 & ~i_10_132_2820_0 & ~i_10_132_3982_0))) | (~i_10_132_2820_0 & ((~i_10_132_223_0 & ~i_10_132_430_0 & ~i_10_132_1554_0 & ~i_10_132_2720_0 & ~i_10_132_2783_0 & ~i_10_132_3496_0 & ~i_10_132_3614_0 & ~i_10_132_3984_0) | (~i_10_132_2657_0 & i_10_132_2828_0 & ~i_10_132_3041_0 & ~i_10_132_3646_0 & ~i_10_132_4129_0 & ~i_10_132_4238_0))) | (~i_10_132_4129_0 & ((~i_10_132_2831_0 & i_10_132_3390_0 & i_10_132_3496_0) | (~i_10_132_997_0 & ~i_10_132_2681_0 & ~i_10_132_2827_0 & ~i_10_132_2985_0 & ~i_10_132_3652_0))) | (~i_10_132_439_0 & ~i_10_132_2635_0 & ~i_10_132_2680_0 & i_10_132_3853_0));
endmodule



// Benchmark "kernel_10_133" written by ABC on Sun Jul 19 10:23:16 2020

module kernel_10_133 ( 
    i_10_133_176_0, i_10_133_178_0, i_10_133_247_0, i_10_133_283_0,
    i_10_133_284_0, i_10_133_286_0, i_10_133_322_0, i_10_133_323_0,
    i_10_133_327_0, i_10_133_407_0, i_10_133_441_0, i_10_133_447_0,
    i_10_133_461_0, i_10_133_504_0, i_10_133_509_0, i_10_133_511_0,
    i_10_133_796_0, i_10_133_957_0, i_10_133_1039_0, i_10_133_1043_0,
    i_10_133_1235_0, i_10_133_1237_0, i_10_133_1246_0, i_10_133_1345_0,
    i_10_133_1346_0, i_10_133_1442_0, i_10_133_1578_0, i_10_133_1649_0,
    i_10_133_1655_0, i_10_133_1683_0, i_10_133_1727_0, i_10_133_1768_0,
    i_10_133_1823_0, i_10_133_1910_0, i_10_133_1912_0, i_10_133_1913_0,
    i_10_133_1951_0, i_10_133_2000_0, i_10_133_2005_0, i_10_133_2028_0,
    i_10_133_2186_0, i_10_133_2361_0, i_10_133_2364_0, i_10_133_2365_0,
    i_10_133_2450_0, i_10_133_2452_0, i_10_133_2453_0, i_10_133_2569_0,
    i_10_133_2632_0, i_10_133_2710_0, i_10_133_2723_0, i_10_133_2735_0,
    i_10_133_2884_0, i_10_133_2916_0, i_10_133_3151_0, i_10_133_3195_0,
    i_10_133_3268_0, i_10_133_3271_0, i_10_133_3274_0, i_10_133_3277_0,
    i_10_133_3278_0, i_10_133_3279_0, i_10_133_3280_0, i_10_133_3281_0,
    i_10_133_3283_0, i_10_133_3322_0, i_10_133_3384_0, i_10_133_3392_0,
    i_10_133_3402_0, i_10_133_3407_0, i_10_133_3520_0, i_10_133_3521_0,
    i_10_133_3537_0, i_10_133_3542_0, i_10_133_3613_0, i_10_133_3614_0,
    i_10_133_3647_0, i_10_133_3648_0, i_10_133_3649_0, i_10_133_3784_0,
    i_10_133_3785_0, i_10_133_3786_0, i_10_133_3787_0, i_10_133_3837_0,
    i_10_133_3846_0, i_10_133_3858_0, i_10_133_3859_0, i_10_133_3894_0,
    i_10_133_3895_0, i_10_133_3896_0, i_10_133_3912_0, i_10_133_3913_0,
    i_10_133_3914_0, i_10_133_4126_0, i_10_133_4281_0, i_10_133_4283_0,
    i_10_133_4288_0, i_10_133_4290_0, i_10_133_4292_0, i_10_133_4565_0,
    o_10_133_0_0  );
  input  i_10_133_176_0, i_10_133_178_0, i_10_133_247_0, i_10_133_283_0,
    i_10_133_284_0, i_10_133_286_0, i_10_133_322_0, i_10_133_323_0,
    i_10_133_327_0, i_10_133_407_0, i_10_133_441_0, i_10_133_447_0,
    i_10_133_461_0, i_10_133_504_0, i_10_133_509_0, i_10_133_511_0,
    i_10_133_796_0, i_10_133_957_0, i_10_133_1039_0, i_10_133_1043_0,
    i_10_133_1235_0, i_10_133_1237_0, i_10_133_1246_0, i_10_133_1345_0,
    i_10_133_1346_0, i_10_133_1442_0, i_10_133_1578_0, i_10_133_1649_0,
    i_10_133_1655_0, i_10_133_1683_0, i_10_133_1727_0, i_10_133_1768_0,
    i_10_133_1823_0, i_10_133_1910_0, i_10_133_1912_0, i_10_133_1913_0,
    i_10_133_1951_0, i_10_133_2000_0, i_10_133_2005_0, i_10_133_2028_0,
    i_10_133_2186_0, i_10_133_2361_0, i_10_133_2364_0, i_10_133_2365_0,
    i_10_133_2450_0, i_10_133_2452_0, i_10_133_2453_0, i_10_133_2569_0,
    i_10_133_2632_0, i_10_133_2710_0, i_10_133_2723_0, i_10_133_2735_0,
    i_10_133_2884_0, i_10_133_2916_0, i_10_133_3151_0, i_10_133_3195_0,
    i_10_133_3268_0, i_10_133_3271_0, i_10_133_3274_0, i_10_133_3277_0,
    i_10_133_3278_0, i_10_133_3279_0, i_10_133_3280_0, i_10_133_3281_0,
    i_10_133_3283_0, i_10_133_3322_0, i_10_133_3384_0, i_10_133_3392_0,
    i_10_133_3402_0, i_10_133_3407_0, i_10_133_3520_0, i_10_133_3521_0,
    i_10_133_3537_0, i_10_133_3542_0, i_10_133_3613_0, i_10_133_3614_0,
    i_10_133_3647_0, i_10_133_3648_0, i_10_133_3649_0, i_10_133_3784_0,
    i_10_133_3785_0, i_10_133_3786_0, i_10_133_3787_0, i_10_133_3837_0,
    i_10_133_3846_0, i_10_133_3858_0, i_10_133_3859_0, i_10_133_3894_0,
    i_10_133_3895_0, i_10_133_3896_0, i_10_133_3912_0, i_10_133_3913_0,
    i_10_133_3914_0, i_10_133_4126_0, i_10_133_4281_0, i_10_133_4283_0,
    i_10_133_4288_0, i_10_133_4290_0, i_10_133_4292_0, i_10_133_4565_0;
  output o_10_133_0_0;
  assign o_10_133_0_0 = ~((~i_10_133_176_0 & ((~i_10_133_178_0 & ~i_10_133_1346_0 & ~i_10_133_2710_0 & ~i_10_133_2723_0 & ~i_10_133_3613_0 & ~i_10_133_3895_0 & ~i_10_133_4290_0) | (~i_10_133_407_0 & ~i_10_133_3195_0 & ~i_10_133_3384_0 & ~i_10_133_3407_0 & ~i_10_133_3542_0 & i_10_133_3649_0 & ~i_10_133_3894_0 & ~i_10_133_4292_0))) | (~i_10_133_178_0 & ((~i_10_133_322_0 & ~i_10_133_447_0 & ~i_10_133_461_0 & ~i_10_133_1910_0 & ~i_10_133_1913_0 & ~i_10_133_3278_0 & ~i_10_133_3402_0 & ~i_10_133_3520_0 & ~i_10_133_3914_0 & ~i_10_133_4126_0 & ~i_10_133_4283_0) | (i_10_133_1578_0 & ~i_10_133_3277_0 & i_10_133_3613_0 & ~i_10_133_3913_0 & ~i_10_133_4290_0))) | (~i_10_133_2005_0 & ((~i_10_133_283_0 & ~i_10_133_3912_0 & ((~i_10_133_407_0 & ~i_10_133_1951_0 & ~i_10_133_2453_0 & i_10_133_2632_0 & ~i_10_133_2884_0 & ~i_10_133_3278_0) | (~i_10_133_1246_0 & ~i_10_133_2450_0 & ~i_10_133_2723_0 & ~i_10_133_2735_0 & ~i_10_133_3402_0 & ~i_10_133_3407_0 & ~i_10_133_3520_0 & ~i_10_133_3537_0 & ~i_10_133_3914_0))) | (~i_10_133_1235_0 & ~i_10_133_4281_0 & ((~i_10_133_1043_0 & ~i_10_133_1345_0 & ~i_10_133_1346_0 & ~i_10_133_1823_0 & ~i_10_133_2452_0 & ~i_10_133_3392_0 & ~i_10_133_3407_0 & ~i_10_133_3537_0 & ~i_10_133_3614_0 & ~i_10_133_4283_0) | (~i_10_133_461_0 & ~i_10_133_2884_0 & ~i_10_133_3384_0 & ~i_10_133_3896_0 & ~i_10_133_4292_0))))) | (~i_10_133_4288_0 & ((~i_10_133_284_0 & ~i_10_133_3895_0 & ((~i_10_133_2710_0 & i_10_133_3384_0) | (~i_10_133_1246_0 & i_10_133_2710_0 & ~i_10_133_3614_0 & ~i_10_133_3837_0))) | (~i_10_133_796_0 & ~i_10_133_957_0 & ~i_10_133_2735_0 & i_10_133_2884_0 & ~i_10_133_3277_0 & ~i_10_133_3281_0 & ~i_10_133_3894_0) | (~i_10_133_323_0 & ~i_10_133_1039_0 & ~i_10_133_1043_0 & ~i_10_133_1912_0 & ~i_10_133_2884_0 & ~i_10_133_3283_0 & ~i_10_133_3521_0 & ~i_10_133_3914_0 & ~i_10_133_4290_0))) | (~i_10_133_3914_0 & ((~i_10_133_1043_0 & ((~i_10_133_322_0 & ~i_10_133_1346_0 & ~i_10_133_2365_0 & ~i_10_133_2710_0 & ~i_10_133_2723_0 & ~i_10_133_3277_0 & ~i_10_133_3281_0 & ~i_10_133_3859_0 & ~i_10_133_3894_0 & ~i_10_133_3895_0 & ~i_10_133_3913_0) | (~i_10_133_247_0 & ~i_10_133_407_0 & ~i_10_133_2450_0 & i_10_133_3281_0 & ~i_10_133_3520_0 & i_10_133_3859_0 & ~i_10_133_4126_0 & ~i_10_133_4281_0))) | (~i_10_133_1039_0 & ~i_10_133_1246_0 & ~i_10_133_1345_0 & ~i_10_133_1910_0 & ~i_10_133_2000_0 & ~i_10_133_2028_0 & ~i_10_133_2365_0 & ~i_10_133_2450_0 & ~i_10_133_2453_0 & ~i_10_133_3268_0 & ~i_10_133_3407_0 & ~i_10_133_3520_0 & ~i_10_133_3537_0 & ~i_10_133_3912_0 & ~i_10_133_4283_0))) | (~i_10_133_4283_0 & ((~i_10_133_247_0 & ((~i_10_133_1235_0 & ~i_10_133_1768_0 & ~i_10_133_1823_0 & ~i_10_133_2710_0 & ~i_10_133_2735_0 & ~i_10_133_3279_0 & ~i_10_133_3542_0 & ~i_10_133_3913_0) | (~i_10_133_322_0 & ~i_10_133_1237_0 & ~i_10_133_1912_0 & ~i_10_133_2000_0 & ~i_10_133_2028_0 & ~i_10_133_2453_0 & ~i_10_133_3281_0 & ~i_10_133_3613_0 & ~i_10_133_3785_0 & ~i_10_133_4292_0))) | (~i_10_133_322_0 & ~i_10_133_1235_0 & ~i_10_133_1237_0 & ~i_10_133_3521_0 & ~i_10_133_3537_0 & ~i_10_133_3542_0 & ~i_10_133_3896_0 & ~i_10_133_3912_0 & ~i_10_133_3913_0 & i_10_133_4292_0))) | (~i_10_133_407_0 & ~i_10_133_2884_0 & ((~i_10_133_286_0 & ~i_10_133_1951_0 & ~i_10_133_2028_0 & ~i_10_133_2453_0 & ~i_10_133_2735_0 & ~i_10_133_3392_0 & ~i_10_133_3859_0 & i_10_133_4290_0) | (~i_10_133_323_0 & ~i_10_133_1246_0 & ~i_10_133_1683_0 & ~i_10_133_1823_0 & ~i_10_133_2000_0 & ~i_10_133_2916_0 & ~i_10_133_3195_0 & ~i_10_133_3271_0 & ~i_10_133_3647_0 & ~i_10_133_4126_0 & ~i_10_133_4290_0))) | (~i_10_133_2453_0 & ((i_10_133_2361_0 & ~i_10_133_3542_0) | (~i_10_133_3277_0 & ~i_10_133_3614_0 & i_10_133_3859_0 & ~i_10_133_4281_0 & ~i_10_133_4290_0))) | (~i_10_133_3278_0 & ((i_10_133_3268_0 & i_10_133_3407_0) | (~i_10_133_1910_0 & ~i_10_133_2028_0 & ~i_10_133_3195_0 & ~i_10_133_3280_0 & ~i_10_133_3520_0 & ~i_10_133_3894_0 & ~i_10_133_3896_0 & ~i_10_133_3913_0 & ~i_10_133_4292_0))) | (~i_10_133_3614_0 & ((i_10_133_2710_0 & i_10_133_3402_0 & i_10_133_3407_0) | (~i_10_133_3279_0 & ~i_10_133_3894_0 & ~i_10_133_3913_0 & i_10_133_4565_0))) | (~i_10_133_4292_0 & ((i_10_133_286_0 & ~i_10_133_3280_0 & i_10_133_3846_0) | (i_10_133_247_0 & ~i_10_133_2450_0 & ~i_10_133_3837_0 & ~i_10_133_3913_0))) | (~i_10_133_322_0 & ~i_10_133_1235_0 & ~i_10_133_2632_0 & i_10_133_3280_0 & ~i_10_133_4281_0 & i_10_133_4288_0 & ~i_10_133_4290_0));
endmodule



// Benchmark "kernel_10_134" written by ABC on Sun Jul 19 10:23:16 2020

module kernel_10_134 ( 
    i_10_134_31_0, i_10_134_37_0, i_10_134_67_0, i_10_134_117_0,
    i_10_134_125_0, i_10_134_259_0, i_10_134_264_0, i_10_134_266_0,
    i_10_134_284_0, i_10_134_317_0, i_10_134_394_0, i_10_134_405_0,
    i_10_134_406_0, i_10_134_688_0, i_10_134_715_0, i_10_134_756_0,
    i_10_134_865_0, i_10_134_866_0, i_10_134_952_0, i_10_134_991_0,
    i_10_134_993_0, i_10_134_1054_0, i_10_134_1084_0, i_10_134_1135_0,
    i_10_134_1136_0, i_10_134_1267_0, i_10_134_1269_0, i_10_134_1281_0,
    i_10_134_1378_0, i_10_134_1438_0, i_10_134_1439_0, i_10_134_1554_0,
    i_10_134_1577_0, i_10_134_1579_0, i_10_134_1582_0, i_10_134_1583_0,
    i_10_134_1687_0, i_10_134_1803_0, i_10_134_1810_0, i_10_134_1811_0,
    i_10_134_1818_0, i_10_134_1846_0, i_10_134_1909_0, i_10_134_1910_0,
    i_10_134_1912_0, i_10_134_1986_0, i_10_134_2017_0, i_10_134_2018_0,
    i_10_134_2185_0, i_10_134_2263_0, i_10_134_2351_0, i_10_134_2353_0,
    i_10_134_2383_0, i_10_134_2404_0, i_10_134_2473_0, i_10_134_2474_0,
    i_10_134_2487_0, i_10_134_2519_0, i_10_134_2536_0, i_10_134_2563_0,
    i_10_134_2578_0, i_10_134_2586_0, i_10_134_2596_0, i_10_134_2607_0,
    i_10_134_2608_0, i_10_134_2702_0, i_10_134_2722_0, i_10_134_2725_0,
    i_10_134_2726_0, i_10_134_2734_0, i_10_134_2735_0, i_10_134_2787_0,
    i_10_134_2809_0, i_10_134_2881_0, i_10_134_2884_0, i_10_134_2885_0,
    i_10_134_2955_0, i_10_134_2983_0, i_10_134_2993_0, i_10_134_3043_0,
    i_10_134_3048_0, i_10_134_3282_0, i_10_134_3283_0, i_10_134_3284_0,
    i_10_134_3356_0, i_10_134_3394_0, i_10_134_3395_0, i_10_134_3562_0,
    i_10_134_3609_0, i_10_134_3841_0, i_10_134_3985_0, i_10_134_4031_0,
    i_10_134_4063_0, i_10_134_4292_0, i_10_134_4377_0, i_10_134_4378_0,
    i_10_134_4397_0, i_10_134_4434_0, i_10_134_4588_0, i_10_134_4589_0,
    o_10_134_0_0  );
  input  i_10_134_31_0, i_10_134_37_0, i_10_134_67_0, i_10_134_117_0,
    i_10_134_125_0, i_10_134_259_0, i_10_134_264_0, i_10_134_266_0,
    i_10_134_284_0, i_10_134_317_0, i_10_134_394_0, i_10_134_405_0,
    i_10_134_406_0, i_10_134_688_0, i_10_134_715_0, i_10_134_756_0,
    i_10_134_865_0, i_10_134_866_0, i_10_134_952_0, i_10_134_991_0,
    i_10_134_993_0, i_10_134_1054_0, i_10_134_1084_0, i_10_134_1135_0,
    i_10_134_1136_0, i_10_134_1267_0, i_10_134_1269_0, i_10_134_1281_0,
    i_10_134_1378_0, i_10_134_1438_0, i_10_134_1439_0, i_10_134_1554_0,
    i_10_134_1577_0, i_10_134_1579_0, i_10_134_1582_0, i_10_134_1583_0,
    i_10_134_1687_0, i_10_134_1803_0, i_10_134_1810_0, i_10_134_1811_0,
    i_10_134_1818_0, i_10_134_1846_0, i_10_134_1909_0, i_10_134_1910_0,
    i_10_134_1912_0, i_10_134_1986_0, i_10_134_2017_0, i_10_134_2018_0,
    i_10_134_2185_0, i_10_134_2263_0, i_10_134_2351_0, i_10_134_2353_0,
    i_10_134_2383_0, i_10_134_2404_0, i_10_134_2473_0, i_10_134_2474_0,
    i_10_134_2487_0, i_10_134_2519_0, i_10_134_2536_0, i_10_134_2563_0,
    i_10_134_2578_0, i_10_134_2586_0, i_10_134_2596_0, i_10_134_2607_0,
    i_10_134_2608_0, i_10_134_2702_0, i_10_134_2722_0, i_10_134_2725_0,
    i_10_134_2726_0, i_10_134_2734_0, i_10_134_2735_0, i_10_134_2787_0,
    i_10_134_2809_0, i_10_134_2881_0, i_10_134_2884_0, i_10_134_2885_0,
    i_10_134_2955_0, i_10_134_2983_0, i_10_134_2993_0, i_10_134_3043_0,
    i_10_134_3048_0, i_10_134_3282_0, i_10_134_3283_0, i_10_134_3284_0,
    i_10_134_3356_0, i_10_134_3394_0, i_10_134_3395_0, i_10_134_3562_0,
    i_10_134_3609_0, i_10_134_3841_0, i_10_134_3985_0, i_10_134_4031_0,
    i_10_134_4063_0, i_10_134_4292_0, i_10_134_4377_0, i_10_134_4378_0,
    i_10_134_4397_0, i_10_134_4434_0, i_10_134_4588_0, i_10_134_4589_0;
  output o_10_134_0_0;
  assign o_10_134_0_0 = 0;
endmodule



// Benchmark "kernel_10_135" written by ABC on Sun Jul 19 10:23:17 2020

module kernel_10_135 ( 
    i_10_135_52_0, i_10_135_171_0, i_10_135_173_0, i_10_135_176_0,
    i_10_135_178_0, i_10_135_179_0, i_10_135_221_0, i_10_135_222_0,
    i_10_135_224_0, i_10_135_279_0, i_10_135_296_0, i_10_135_328_0,
    i_10_135_329_0, i_10_135_390_0, i_10_135_391_0, i_10_135_394_0,
    i_10_135_439_0, i_10_135_446_0, i_10_135_449_0, i_10_135_515_0,
    i_10_135_516_0, i_10_135_517_0, i_10_135_518_0, i_10_135_521_0,
    i_10_135_596_0, i_10_135_957_0, i_10_135_959_0, i_10_135_998_0,
    i_10_135_1138_0, i_10_135_1160_0, i_10_135_1265_0, i_10_135_1268_0,
    i_10_135_1445_0, i_10_135_1636_0, i_10_135_1651_0, i_10_135_1652_0,
    i_10_135_1686_0, i_10_135_1687_0, i_10_135_1817_0, i_10_135_1819_0,
    i_10_135_1821_0, i_10_135_1877_0, i_10_135_2026_0, i_10_135_2179_0,
    i_10_135_2201_0, i_10_135_2255_0, i_10_135_2330_0, i_10_135_2353_0,
    i_10_135_2354_0, i_10_135_2364_0, i_10_135_2515_0, i_10_135_2631_0,
    i_10_135_2636_0, i_10_135_2675_0, i_10_135_2678_0, i_10_135_2681_0,
    i_10_135_2705_0, i_10_135_2706_0, i_10_135_2725_0, i_10_135_2821_0,
    i_10_135_2825_0, i_10_135_2829_0, i_10_135_2920_0, i_10_135_2980_0,
    i_10_135_2984_0, i_10_135_3035_0, i_10_135_3036_0, i_10_135_3038_0,
    i_10_135_3199_0, i_10_135_3275_0, i_10_135_3281_0, i_10_135_3290_0,
    i_10_135_3293_0, i_10_135_3494_0, i_10_135_3497_0, i_10_135_3523_0,
    i_10_135_3524_0, i_10_135_3527_0, i_10_135_3583_0, i_10_135_3616_0,
    i_10_135_3781_0, i_10_135_3782_0, i_10_135_3784_0, i_10_135_3785_0,
    i_10_135_3787_0, i_10_135_3788_0, i_10_135_3800_0, i_10_135_3910_0,
    i_10_135_3911_0, i_10_135_3913_0, i_10_135_3914_0, i_10_135_3950_0,
    i_10_135_4120_0, i_10_135_4121_0, i_10_135_4127_0, i_10_135_4130_0,
    i_10_135_4238_0, i_10_135_4268_0, i_10_135_4280_0, i_10_135_4463_0,
    o_10_135_0_0  );
  input  i_10_135_52_0, i_10_135_171_0, i_10_135_173_0, i_10_135_176_0,
    i_10_135_178_0, i_10_135_179_0, i_10_135_221_0, i_10_135_222_0,
    i_10_135_224_0, i_10_135_279_0, i_10_135_296_0, i_10_135_328_0,
    i_10_135_329_0, i_10_135_390_0, i_10_135_391_0, i_10_135_394_0,
    i_10_135_439_0, i_10_135_446_0, i_10_135_449_0, i_10_135_515_0,
    i_10_135_516_0, i_10_135_517_0, i_10_135_518_0, i_10_135_521_0,
    i_10_135_596_0, i_10_135_957_0, i_10_135_959_0, i_10_135_998_0,
    i_10_135_1138_0, i_10_135_1160_0, i_10_135_1265_0, i_10_135_1268_0,
    i_10_135_1445_0, i_10_135_1636_0, i_10_135_1651_0, i_10_135_1652_0,
    i_10_135_1686_0, i_10_135_1687_0, i_10_135_1817_0, i_10_135_1819_0,
    i_10_135_1821_0, i_10_135_1877_0, i_10_135_2026_0, i_10_135_2179_0,
    i_10_135_2201_0, i_10_135_2255_0, i_10_135_2330_0, i_10_135_2353_0,
    i_10_135_2354_0, i_10_135_2364_0, i_10_135_2515_0, i_10_135_2631_0,
    i_10_135_2636_0, i_10_135_2675_0, i_10_135_2678_0, i_10_135_2681_0,
    i_10_135_2705_0, i_10_135_2706_0, i_10_135_2725_0, i_10_135_2821_0,
    i_10_135_2825_0, i_10_135_2829_0, i_10_135_2920_0, i_10_135_2980_0,
    i_10_135_2984_0, i_10_135_3035_0, i_10_135_3036_0, i_10_135_3038_0,
    i_10_135_3199_0, i_10_135_3275_0, i_10_135_3281_0, i_10_135_3290_0,
    i_10_135_3293_0, i_10_135_3494_0, i_10_135_3497_0, i_10_135_3523_0,
    i_10_135_3524_0, i_10_135_3527_0, i_10_135_3583_0, i_10_135_3616_0,
    i_10_135_3781_0, i_10_135_3782_0, i_10_135_3784_0, i_10_135_3785_0,
    i_10_135_3787_0, i_10_135_3788_0, i_10_135_3800_0, i_10_135_3910_0,
    i_10_135_3911_0, i_10_135_3913_0, i_10_135_3914_0, i_10_135_3950_0,
    i_10_135_4120_0, i_10_135_4121_0, i_10_135_4127_0, i_10_135_4130_0,
    i_10_135_4238_0, i_10_135_4268_0, i_10_135_4280_0, i_10_135_4463_0;
  output o_10_135_0_0;
  assign o_10_135_0_0 = ~((~i_10_135_1877_0 & ((~i_10_135_222_0 & ~i_10_135_4280_0 & ((~i_10_135_329_0 & ~i_10_135_515_0 & ~i_10_135_1817_0 & ~i_10_135_2201_0 & ~i_10_135_2330_0 & ~i_10_135_2678_0 & ~i_10_135_2821_0 & ~i_10_135_2829_0 & ~i_10_135_3524_0 & ~i_10_135_3527_0 & ~i_10_135_3910_0 & ~i_10_135_3950_0) | (~i_10_135_279_0 & i_10_135_516_0 & ~i_10_135_2675_0 & ~i_10_135_3494_0 & ~i_10_135_4121_0))) | (~i_10_135_2984_0 & ((i_10_135_2353_0 & ~i_10_135_2678_0 & ~i_10_135_3911_0 & ~i_10_135_4120_0 & i_10_135_4127_0) | (~i_10_135_296_0 & ~i_10_135_998_0 & ~i_10_135_1687_0 & ~i_10_135_2179_0 & i_10_135_2706_0 & ~i_10_135_3527_0 & ~i_10_135_4238_0))) | (~i_10_135_173_0 & ~i_10_135_957_0 & ~i_10_135_1265_0 & ~i_10_135_2330_0 & ~i_10_135_2364_0 & ~i_10_135_2705_0 & ~i_10_135_3494_0 & ~i_10_135_3497_0 & ~i_10_135_3523_0 & ~i_10_135_3911_0 & ~i_10_135_3950_0))) | (~i_10_135_4268_0 & ((~i_10_135_224_0 & ((~i_10_135_221_0 & ~i_10_135_279_0 & ~i_10_135_394_0 & ~i_10_135_1265_0 & ~i_10_135_1821_0 & ~i_10_135_2821_0 & ~i_10_135_2920_0 & ~i_10_135_3275_0 & ~i_10_135_3527_0 & ~i_10_135_3616_0 & ~i_10_135_3914_0 & ~i_10_135_3950_0) | (~i_10_135_515_0 & ~i_10_135_521_0 & ~i_10_135_957_0 & ~i_10_135_2706_0 & ~i_10_135_3523_0 & ~i_10_135_3524_0 & ~i_10_135_4120_0))) | (~i_10_135_176_0 & ~i_10_135_1268_0 & i_10_135_2636_0 & ~i_10_135_2706_0 & ~i_10_135_2825_0 & ~i_10_135_3035_0 & ~i_10_135_3497_0 & ~i_10_135_3524_0 & ~i_10_135_4127_0 & ~i_10_135_4280_0))) | (~i_10_135_521_0 & ((~i_10_135_176_0 & ((~i_10_135_329_0 & ~i_10_135_2636_0 & ~i_10_135_2706_0 & ~i_10_135_2920_0 & ~i_10_135_2980_0 & ~i_10_135_2984_0) | (~i_10_135_998_0 & ~i_10_135_2675_0 & ~i_10_135_2678_0 & ~i_10_135_2705_0 & ~i_10_135_3524_0 & ~i_10_135_3527_0))) | (~i_10_135_279_0 & ~i_10_135_998_0 & ~i_10_135_2354_0 & ~i_10_135_2675_0 & ~i_10_135_3281_0 & ~i_10_135_3524_0 & ~i_10_135_4280_0))) | (~i_10_135_1265_0 & ((~i_10_135_173_0 & ~i_10_135_178_0 & ~i_10_135_518_0 & ~i_10_135_1445_0 & ~i_10_135_2825_0 & ~i_10_135_3038_0) | (~i_10_135_1821_0 & i_10_135_2631_0 & i_10_135_2675_0 & ~i_10_135_2920_0 & ~i_10_135_2984_0 & ~i_10_135_3524_0 & ~i_10_135_3910_0))) | (~i_10_135_173_0 & ((~i_10_135_2636_0 & i_10_135_3035_0 & ~i_10_135_3281_0) | (~i_10_135_515_0 & ~i_10_135_2330_0 & ~i_10_135_2725_0 & ~i_10_135_2825_0 & ~i_10_135_2984_0 & ~i_10_135_3523_0 & ~i_10_135_3914_0))) | (~i_10_135_518_0 & ((~i_10_135_515_0 & ~i_10_135_2330_0 & ~i_10_135_2354_0 & ~i_10_135_3281_0 & ~i_10_135_3524_0 & ~i_10_135_3527_0) | (~i_10_135_1445_0 & ~i_10_135_2725_0 & ~i_10_135_3523_0 & ~i_10_135_4127_0))) | (~i_10_135_515_0 & ((~i_10_135_998_0 & ~i_10_135_2353_0 & ~i_10_135_2984_0 & i_10_135_3199_0 & ~i_10_135_3275_0 & ~i_10_135_3583_0 & ~i_10_135_3914_0) | (i_10_135_3785_0 & i_10_135_4127_0))) | (~i_10_135_1819_0 & ~i_10_135_3583_0 & ((~i_10_135_516_0 & ~i_10_135_2364_0 & ~i_10_135_2705_0 & ~i_10_135_2725_0 & ~i_10_135_2821_0 & ~i_10_135_2920_0 & ~i_10_135_3497_0 & ~i_10_135_3524_0) | (~i_10_135_1821_0 & ~i_10_135_2636_0 & i_10_135_2920_0 & i_10_135_4127_0))) | (i_10_135_4268_0 & (i_10_135_959_0 | (i_10_135_3616_0 & i_10_135_4280_0))) | (i_10_135_279_0 & ~i_10_135_296_0 & ~i_10_135_957_0 & ~i_10_135_2675_0 & ~i_10_135_2681_0 & ~i_10_135_2920_0 & ~i_10_135_2980_0 & ~i_10_135_3524_0 & ~i_10_135_3527_0 & ~i_10_135_3910_0));
endmodule



// Benchmark "kernel_10_136" written by ABC on Sun Jul 19 10:23:19 2020

module kernel_10_136 ( 
    i_10_136_174_0, i_10_136_219_0, i_10_136_286_0, i_10_136_318_0,
    i_10_136_328_0, i_10_136_424_0, i_10_136_444_0, i_10_136_446_0,
    i_10_136_793_0, i_10_136_799_0, i_10_136_896_0, i_10_136_955_0,
    i_10_136_1032_0, i_10_136_1033_0, i_10_136_1308_0, i_10_136_1437_0,
    i_10_136_1542_0, i_10_136_1583_0, i_10_136_1650_0, i_10_136_1688_0,
    i_10_136_1765_0, i_10_136_1821_0, i_10_136_1822_0, i_10_136_1912_0,
    i_10_136_1913_0, i_10_136_1995_0, i_10_136_2178_0, i_10_136_2179_0,
    i_10_136_2180_0, i_10_136_2305_0, i_10_136_2306_0, i_10_136_2326_0,
    i_10_136_2350_0, i_10_136_2351_0, i_10_136_2352_0, i_10_136_2353_0,
    i_10_136_2361_0, i_10_136_2382_0, i_10_136_2404_0, i_10_136_2452_0,
    i_10_136_2502_0, i_10_136_2571_0, i_10_136_2633_0, i_10_136_2636_0,
    i_10_136_2673_0, i_10_136_2705_0, i_10_136_2714_0, i_10_136_2727_0,
    i_10_136_2728_0, i_10_136_2729_0, i_10_136_2733_0, i_10_136_2734_0,
    i_10_136_2735_0, i_10_136_2826_0, i_10_136_2827_0, i_10_136_2830_0,
    i_10_136_2832_0, i_10_136_2922_0, i_10_136_3070_0, i_10_136_3153_0,
    i_10_136_3155_0, i_10_136_3162_0, i_10_136_3196_0, i_10_136_3199_0,
    i_10_136_3202_0, i_10_136_3268_0, i_10_136_3270_0, i_10_136_3277_0,
    i_10_136_3326_0, i_10_136_3385_0, i_10_136_3388_0, i_10_136_3389_0,
    i_10_136_3390_0, i_10_136_3470_0, i_10_136_3612_0, i_10_136_3613_0,
    i_10_136_3649_0, i_10_136_3652_0, i_10_136_3683_0, i_10_136_3732_0,
    i_10_136_3780_0, i_10_136_3782_0, i_10_136_3834_0, i_10_136_3857_0,
    i_10_136_3907_0, i_10_136_3982_0, i_10_136_4050_0, i_10_136_4051_0,
    i_10_136_4119_0, i_10_136_4128_0, i_10_136_4129_0, i_10_136_4130_0,
    i_10_136_4168_0, i_10_136_4169_0, i_10_136_4219_0, i_10_136_4270_0,
    i_10_136_4281_0, i_10_136_4288_0, i_10_136_4566_0, i_10_136_4569_0,
    o_10_136_0_0  );
  input  i_10_136_174_0, i_10_136_219_0, i_10_136_286_0, i_10_136_318_0,
    i_10_136_328_0, i_10_136_424_0, i_10_136_444_0, i_10_136_446_0,
    i_10_136_793_0, i_10_136_799_0, i_10_136_896_0, i_10_136_955_0,
    i_10_136_1032_0, i_10_136_1033_0, i_10_136_1308_0, i_10_136_1437_0,
    i_10_136_1542_0, i_10_136_1583_0, i_10_136_1650_0, i_10_136_1688_0,
    i_10_136_1765_0, i_10_136_1821_0, i_10_136_1822_0, i_10_136_1912_0,
    i_10_136_1913_0, i_10_136_1995_0, i_10_136_2178_0, i_10_136_2179_0,
    i_10_136_2180_0, i_10_136_2305_0, i_10_136_2306_0, i_10_136_2326_0,
    i_10_136_2350_0, i_10_136_2351_0, i_10_136_2352_0, i_10_136_2353_0,
    i_10_136_2361_0, i_10_136_2382_0, i_10_136_2404_0, i_10_136_2452_0,
    i_10_136_2502_0, i_10_136_2571_0, i_10_136_2633_0, i_10_136_2636_0,
    i_10_136_2673_0, i_10_136_2705_0, i_10_136_2714_0, i_10_136_2727_0,
    i_10_136_2728_0, i_10_136_2729_0, i_10_136_2733_0, i_10_136_2734_0,
    i_10_136_2735_0, i_10_136_2826_0, i_10_136_2827_0, i_10_136_2830_0,
    i_10_136_2832_0, i_10_136_2922_0, i_10_136_3070_0, i_10_136_3153_0,
    i_10_136_3155_0, i_10_136_3162_0, i_10_136_3196_0, i_10_136_3199_0,
    i_10_136_3202_0, i_10_136_3268_0, i_10_136_3270_0, i_10_136_3277_0,
    i_10_136_3326_0, i_10_136_3385_0, i_10_136_3388_0, i_10_136_3389_0,
    i_10_136_3390_0, i_10_136_3470_0, i_10_136_3612_0, i_10_136_3613_0,
    i_10_136_3649_0, i_10_136_3652_0, i_10_136_3683_0, i_10_136_3732_0,
    i_10_136_3780_0, i_10_136_3782_0, i_10_136_3834_0, i_10_136_3857_0,
    i_10_136_3907_0, i_10_136_3982_0, i_10_136_4050_0, i_10_136_4051_0,
    i_10_136_4119_0, i_10_136_4128_0, i_10_136_4129_0, i_10_136_4130_0,
    i_10_136_4168_0, i_10_136_4169_0, i_10_136_4219_0, i_10_136_4270_0,
    i_10_136_4281_0, i_10_136_4288_0, i_10_136_4566_0, i_10_136_4569_0;
  output o_10_136_0_0;
  assign o_10_136_0_0 = ~((~i_10_136_318_0 & ((i_10_136_286_0 & ~i_10_136_1032_0 & i_10_136_2452_0 & ~i_10_136_4050_0) | (~i_10_136_219_0 & ~i_10_136_424_0 & ~i_10_136_444_0 & ~i_10_136_793_0 & ~i_10_136_955_0 & ~i_10_136_1437_0 & ~i_10_136_1583_0 & ~i_10_136_2179_0 & ~i_10_136_2727_0 & ~i_10_136_2922_0 & ~i_10_136_3070_0 & ~i_10_136_3683_0 & ~i_10_136_4130_0))) | (~i_10_136_424_0 & ((~i_10_136_446_0 & ~i_10_136_2305_0 & ~i_10_136_2452_0 & i_10_136_2729_0 & ~i_10_136_2922_0 & ~i_10_136_3782_0 & ~i_10_136_4050_0) | (~i_10_136_1822_0 & i_10_136_2353_0 & ~i_10_136_2714_0 & ~i_10_136_3070_0 & ~i_10_136_3683_0 & ~i_10_136_4281_0))) | (~i_10_136_1032_0 & ((~i_10_136_446_0 & ~i_10_136_3199_0 & i_10_136_3907_0) | (i_10_136_174_0 & ~i_10_136_1308_0 & ~i_10_136_1688_0 & i_10_136_2452_0 & i_10_136_3612_0 & ~i_10_136_4050_0))) | (~i_10_136_4128_0 & ((~i_10_136_2180_0 & ((~i_10_136_1033_0 & ~i_10_136_2305_0 & ~i_10_136_2728_0 & ~i_10_136_3199_0 & ((~i_10_136_1688_0 & ~i_10_136_2352_0 & ~i_10_136_2361_0 & ~i_10_136_2452_0 & ~i_10_136_2502_0 & ~i_10_136_3470_0 & ~i_10_136_3612_0 & ~i_10_136_3857_0) | (~i_10_136_174_0 & ~i_10_136_2178_0 & ~i_10_136_2727_0 & ~i_10_136_2827_0 & ~i_10_136_2830_0 & ~i_10_136_3070_0 & ~i_10_136_3782_0 & ~i_10_136_4050_0 & ~i_10_136_4129_0))) | (~i_10_136_2178_0 & ((~i_10_136_2361_0 & ~i_10_136_2733_0 & i_10_136_2922_0 & ~i_10_136_3202_0 & ~i_10_136_3277_0) | (~i_10_136_1308_0 & ~i_10_136_1821_0 & ~i_10_136_2306_0 & ~i_10_136_2705_0 & ~i_10_136_2734_0 & ~i_10_136_3613_0))) | (~i_10_136_1821_0 & ((~i_10_136_2179_0 & ~i_10_136_2306_0 & ~i_10_136_2727_0 & ~i_10_136_3202_0 & ~i_10_136_3683_0 & ~i_10_136_4130_0 & ~i_10_136_3389_0 & ~i_10_136_3612_0) | (~i_10_136_1650_0 & ~i_10_136_3070_0 & i_10_136_3389_0 & ~i_10_136_4281_0))))) | (~i_10_136_1437_0 & ~i_10_136_2673_0 & ((~i_10_136_955_0 & ~i_10_136_2179_0 & ~i_10_136_2306_0 & i_10_136_4270_0) | (~i_10_136_219_0 & ~i_10_136_1821_0 & ~i_10_136_2452_0 & ~i_10_136_2827_0 & ~i_10_136_3070_0 & ~i_10_136_3389_0 & ~i_10_136_3470_0 & ~i_10_136_3683_0 & ~i_10_136_4051_0 & ~i_10_136_4288_0))) | (~i_10_136_444_0 & ~i_10_136_1650_0 & ~i_10_136_1995_0 & ~i_10_136_2178_0 & ~i_10_136_2305_0 & ~i_10_136_2306_0 & ~i_10_136_2832_0 & ~i_10_136_3199_0 & ~i_10_136_3270_0 & ~i_10_136_3683_0 & ~i_10_136_3780_0 & ~i_10_136_3982_0 & ~i_10_136_4050_0 & ~i_10_136_4281_0))) | (~i_10_136_174_0 & ((~i_10_136_1688_0 & ~i_10_136_2179_0 & i_10_136_2826_0 & i_10_136_2827_0 & ~i_10_136_4051_0 & ~i_10_136_4119_0) | (~i_10_136_1033_0 & ~i_10_136_1308_0 & ~i_10_136_2326_0 & ~i_10_136_2705_0 & ~i_10_136_2727_0 & ~i_10_136_3196_0 & ~i_10_136_3270_0 & ~i_10_136_3649_0 & ~i_10_136_4270_0))) | (~i_10_136_3196_0 & ((~i_10_136_219_0 & ~i_10_136_3612_0 & ~i_10_136_3613_0 & ((~i_10_136_1437_0 & ~i_10_136_1821_0 & ~i_10_136_2180_0 & ~i_10_136_2714_0 & ~i_10_136_3834_0 & ~i_10_136_4129_0) | (~i_10_136_955_0 & ~i_10_136_1308_0 & ~i_10_136_2179_0 & ~i_10_136_2502_0 & ~i_10_136_2571_0 & ~i_10_136_3683_0 & ~i_10_136_3780_0 & ~i_10_136_4219_0))) | (~i_10_136_799_0 & ~i_10_136_1308_0 & ~i_10_136_1437_0 & ~i_10_136_2180_0 & ~i_10_136_2305_0 & ~i_10_136_2306_0 & ~i_10_136_2361_0 & ~i_10_136_2633_0 & ~i_10_136_2922_0 & ~i_10_136_3162_0 & ~i_10_136_4050_0 & ~i_10_136_4051_0))) | (~i_10_136_2178_0 & ((~i_10_136_3683_0 & ((~i_10_136_1308_0 & ((~i_10_136_1821_0 & ~i_10_136_2306_0 & ~i_10_136_2571_0 & ~i_10_136_3199_0) | (~i_10_136_1437_0 & ~i_10_136_1995_0 & ~i_10_136_2179_0 & ~i_10_136_2180_0 & ~i_10_136_2350_0 & ~i_10_136_2452_0 & ~i_10_136_3070_0 & ~i_10_136_3613_0))) | (~i_10_136_444_0 & ~i_10_136_1437_0 & ~i_10_136_1822_0 & ~i_10_136_3649_0 & ~i_10_136_3732_0 & ~i_10_136_4130_0 & ~i_10_136_4281_0))) | (i_10_136_446_0 & ~i_10_136_2305_0 & ~i_10_136_2571_0 & ~i_10_136_2832_0 & ~i_10_136_3268_0 & ~i_10_136_3390_0 & ~i_10_136_3652_0 & ~i_10_136_3782_0 & ~i_10_136_3982_0 & ~i_10_136_4051_0 & ~i_10_136_4219_0))) | (i_10_136_2636_0 & ((~i_10_136_444_0 & ((~i_10_136_2306_0 & ~i_10_136_3732_0 & ~i_10_136_3780_0 & ~i_10_136_4050_0 & i_10_136_4119_0 & ~i_10_136_4281_0) | (~i_10_136_4288_0 & i_10_136_4569_0))) | (i_10_136_2353_0 & i_10_136_4270_0 & ~i_10_136_4566_0))) | (~i_10_136_2306_0 & (i_10_136_328_0 | (~i_10_136_2305_0 & ~i_10_136_2350_0 & i_10_136_2826_0 & ~i_10_136_4051_0 & ~i_10_136_4219_0 & ~i_10_136_3070_0 & ~i_10_136_3982_0))) | (~i_10_136_2305_0 & ((~i_10_136_1033_0 & ~i_10_136_2180_0 & i_10_136_2827_0 & ~i_10_136_3780_0) | (~i_10_136_955_0 & ~i_10_136_1542_0 & ~i_10_136_1995_0 & i_10_136_3388_0 & ~i_10_136_3389_0 & ~i_10_136_3857_0))) | (~i_10_136_1821_0 & ~i_10_136_2452_0 & ~i_10_136_3070_0 & i_10_136_3385_0 & i_10_136_3613_0 & ~i_10_136_3652_0) | (~i_10_136_793_0 & i_10_136_3683_0 & i_10_136_4270_0) | (~i_10_136_1437_0 & ~i_10_136_1688_0 & i_10_136_2353_0 & ~i_10_136_2705_0 & ~i_10_136_3390_0 & ~i_10_136_4051_0 & ~i_10_136_4270_0));
endmodule



// Benchmark "kernel_10_137" written by ABC on Sun Jul 19 10:23:20 2020

module kernel_10_137 ( 
    i_10_137_37_0, i_10_137_148_0, i_10_137_222_0, i_10_137_223_0,
    i_10_137_325_0, i_10_137_352_0, i_10_137_445_0, i_10_137_459_0,
    i_10_137_462_0, i_10_137_520_0, i_10_137_586_0, i_10_137_587_0,
    i_10_137_594_0, i_10_137_729_0, i_10_137_730_0, i_10_137_749_0,
    i_10_137_795_0, i_10_137_834_0, i_10_137_846_0, i_10_137_892_0,
    i_10_137_955_0, i_10_137_956_0, i_10_137_1026_0, i_10_137_1027_0,
    i_10_137_1039_0, i_10_137_1042_0, i_10_137_1117_0, i_10_137_1118_0,
    i_10_137_1161_0, i_10_137_1185_0, i_10_137_1333_0, i_10_137_1342_0,
    i_10_137_1344_0, i_10_137_1353_0, i_10_137_1362_0, i_10_137_1371_0,
    i_10_137_1574_0, i_10_137_1579_0, i_10_137_1650_0, i_10_137_1767_0,
    i_10_137_1801_0, i_10_137_1802_0, i_10_137_1810_0, i_10_137_1818_0,
    i_10_137_1819_0, i_10_137_1821_0, i_10_137_1875_0, i_10_137_1956_0,
    i_10_137_2200_0, i_10_137_2338_0, i_10_137_2351_0, i_10_137_2405_0,
    i_10_137_2451_0, i_10_137_2462_0, i_10_137_2512_0, i_10_137_2538_0,
    i_10_137_2543_0, i_10_137_2556_0, i_10_137_2568_0, i_10_137_2679_0,
    i_10_137_2704_0, i_10_137_2730_0, i_10_137_2754_0, i_10_137_2829_0,
    i_10_137_2830_0, i_10_137_2882_0, i_10_137_2922_0, i_10_137_2955_0,
    i_10_137_2992_0, i_10_137_3047_0, i_10_137_3049_0, i_10_137_3228_0,
    i_10_137_3267_0, i_10_137_3272_0, i_10_137_3384_0, i_10_137_3432_0,
    i_10_137_3433_0, i_10_137_3481_0, i_10_137_3519_0, i_10_137_3520_0,
    i_10_137_3522_0, i_10_137_3583_0, i_10_137_3584_0, i_10_137_3609_0,
    i_10_137_3614_0, i_10_137_3684_0, i_10_137_3723_0, i_10_137_3725_0,
    i_10_137_3857_0, i_10_137_4005_0, i_10_137_4006_0, i_10_137_4007_0,
    i_10_137_4118_0, i_10_137_4236_0, i_10_137_4285_0, i_10_137_4287_0,
    i_10_137_4324_0, i_10_137_4425_0, i_10_137_4488_0, i_10_137_4566_0,
    o_10_137_0_0  );
  input  i_10_137_37_0, i_10_137_148_0, i_10_137_222_0, i_10_137_223_0,
    i_10_137_325_0, i_10_137_352_0, i_10_137_445_0, i_10_137_459_0,
    i_10_137_462_0, i_10_137_520_0, i_10_137_586_0, i_10_137_587_0,
    i_10_137_594_0, i_10_137_729_0, i_10_137_730_0, i_10_137_749_0,
    i_10_137_795_0, i_10_137_834_0, i_10_137_846_0, i_10_137_892_0,
    i_10_137_955_0, i_10_137_956_0, i_10_137_1026_0, i_10_137_1027_0,
    i_10_137_1039_0, i_10_137_1042_0, i_10_137_1117_0, i_10_137_1118_0,
    i_10_137_1161_0, i_10_137_1185_0, i_10_137_1333_0, i_10_137_1342_0,
    i_10_137_1344_0, i_10_137_1353_0, i_10_137_1362_0, i_10_137_1371_0,
    i_10_137_1574_0, i_10_137_1579_0, i_10_137_1650_0, i_10_137_1767_0,
    i_10_137_1801_0, i_10_137_1802_0, i_10_137_1810_0, i_10_137_1818_0,
    i_10_137_1819_0, i_10_137_1821_0, i_10_137_1875_0, i_10_137_1956_0,
    i_10_137_2200_0, i_10_137_2338_0, i_10_137_2351_0, i_10_137_2405_0,
    i_10_137_2451_0, i_10_137_2462_0, i_10_137_2512_0, i_10_137_2538_0,
    i_10_137_2543_0, i_10_137_2556_0, i_10_137_2568_0, i_10_137_2679_0,
    i_10_137_2704_0, i_10_137_2730_0, i_10_137_2754_0, i_10_137_2829_0,
    i_10_137_2830_0, i_10_137_2882_0, i_10_137_2922_0, i_10_137_2955_0,
    i_10_137_2992_0, i_10_137_3047_0, i_10_137_3049_0, i_10_137_3228_0,
    i_10_137_3267_0, i_10_137_3272_0, i_10_137_3384_0, i_10_137_3432_0,
    i_10_137_3433_0, i_10_137_3481_0, i_10_137_3519_0, i_10_137_3520_0,
    i_10_137_3522_0, i_10_137_3583_0, i_10_137_3584_0, i_10_137_3609_0,
    i_10_137_3614_0, i_10_137_3684_0, i_10_137_3723_0, i_10_137_3725_0,
    i_10_137_3857_0, i_10_137_4005_0, i_10_137_4006_0, i_10_137_4007_0,
    i_10_137_4118_0, i_10_137_4236_0, i_10_137_4285_0, i_10_137_4287_0,
    i_10_137_4324_0, i_10_137_4425_0, i_10_137_4488_0, i_10_137_4566_0;
  output o_10_137_0_0;
  assign o_10_137_0_0 = 0;
endmodule



// Benchmark "kernel_10_138" written by ABC on Sun Jul 19 10:23:20 2020

module kernel_10_138 ( 
    i_10_138_34_0, i_10_138_171_0, i_10_138_178_0, i_10_138_250_0,
    i_10_138_283_0, i_10_138_318_0, i_10_138_392_0, i_10_138_409_0,
    i_10_138_410_0, i_10_138_441_0, i_10_138_448_0, i_10_138_449_0,
    i_10_138_514_0, i_10_138_751_0, i_10_138_963_0, i_10_138_1034_0,
    i_10_138_1080_0, i_10_138_1242_0, i_10_138_1246_0, i_10_138_1248_0,
    i_10_138_1249_0, i_10_138_1308_0, i_10_138_1547_0, i_10_138_1575_0,
    i_10_138_1578_0, i_10_138_1651_0, i_10_138_1760_0, i_10_138_1823_0,
    i_10_138_1915_0, i_10_138_2006_0, i_10_138_2022_0, i_10_138_2359_0,
    i_10_138_2411_0, i_10_138_2470_0, i_10_138_2473_0, i_10_138_2474_0,
    i_10_138_2537_0, i_10_138_2654_0, i_10_138_2659_0, i_10_138_2681_0,
    i_10_138_2710_0, i_10_138_2728_0, i_10_138_2729_0, i_10_138_2730_0,
    i_10_138_2833_0, i_10_138_2869_0, i_10_138_2920_0, i_10_138_2921_0,
    i_10_138_3034_0, i_10_138_3036_0, i_10_138_3037_0, i_10_138_3038_0,
    i_10_138_3039_0, i_10_138_3162_0, i_10_138_3199_0, i_10_138_3200_0,
    i_10_138_3202_0, i_10_138_3279_0, i_10_138_3281_0, i_10_138_3284_0,
    i_10_138_3338_0, i_10_138_3384_0, i_10_138_3386_0, i_10_138_3389_0,
    i_10_138_3403_0, i_10_138_3408_0, i_10_138_3433_0, i_10_138_3434_0,
    i_10_138_3466_0, i_10_138_3496_0, i_10_138_3522_0, i_10_138_3526_0,
    i_10_138_3612_0, i_10_138_3614_0, i_10_138_3648_0, i_10_138_3727_0,
    i_10_138_3733_0, i_10_138_3782_0, i_10_138_3783_0, i_10_138_3784_0,
    i_10_138_3785_0, i_10_138_3787_0, i_10_138_3835_0, i_10_138_3836_0,
    i_10_138_3844_0, i_10_138_3846_0, i_10_138_3848_0, i_10_138_3855_0,
    i_10_138_3856_0, i_10_138_3857_0, i_10_138_3860_0, i_10_138_3983_0,
    i_10_138_4120_0, i_10_138_4121_0, i_10_138_4220_0, i_10_138_4286_0,
    i_10_138_4289_0, i_10_138_4567_0, i_10_138_4568_0, i_10_138_4569_0,
    o_10_138_0_0  );
  input  i_10_138_34_0, i_10_138_171_0, i_10_138_178_0, i_10_138_250_0,
    i_10_138_283_0, i_10_138_318_0, i_10_138_392_0, i_10_138_409_0,
    i_10_138_410_0, i_10_138_441_0, i_10_138_448_0, i_10_138_449_0,
    i_10_138_514_0, i_10_138_751_0, i_10_138_963_0, i_10_138_1034_0,
    i_10_138_1080_0, i_10_138_1242_0, i_10_138_1246_0, i_10_138_1248_0,
    i_10_138_1249_0, i_10_138_1308_0, i_10_138_1547_0, i_10_138_1575_0,
    i_10_138_1578_0, i_10_138_1651_0, i_10_138_1760_0, i_10_138_1823_0,
    i_10_138_1915_0, i_10_138_2006_0, i_10_138_2022_0, i_10_138_2359_0,
    i_10_138_2411_0, i_10_138_2470_0, i_10_138_2473_0, i_10_138_2474_0,
    i_10_138_2537_0, i_10_138_2654_0, i_10_138_2659_0, i_10_138_2681_0,
    i_10_138_2710_0, i_10_138_2728_0, i_10_138_2729_0, i_10_138_2730_0,
    i_10_138_2833_0, i_10_138_2869_0, i_10_138_2920_0, i_10_138_2921_0,
    i_10_138_3034_0, i_10_138_3036_0, i_10_138_3037_0, i_10_138_3038_0,
    i_10_138_3039_0, i_10_138_3162_0, i_10_138_3199_0, i_10_138_3200_0,
    i_10_138_3202_0, i_10_138_3279_0, i_10_138_3281_0, i_10_138_3284_0,
    i_10_138_3338_0, i_10_138_3384_0, i_10_138_3386_0, i_10_138_3389_0,
    i_10_138_3403_0, i_10_138_3408_0, i_10_138_3433_0, i_10_138_3434_0,
    i_10_138_3466_0, i_10_138_3496_0, i_10_138_3522_0, i_10_138_3526_0,
    i_10_138_3612_0, i_10_138_3614_0, i_10_138_3648_0, i_10_138_3727_0,
    i_10_138_3733_0, i_10_138_3782_0, i_10_138_3783_0, i_10_138_3784_0,
    i_10_138_3785_0, i_10_138_3787_0, i_10_138_3835_0, i_10_138_3836_0,
    i_10_138_3844_0, i_10_138_3846_0, i_10_138_3848_0, i_10_138_3855_0,
    i_10_138_3856_0, i_10_138_3857_0, i_10_138_3860_0, i_10_138_3983_0,
    i_10_138_4120_0, i_10_138_4121_0, i_10_138_4220_0, i_10_138_4286_0,
    i_10_138_4289_0, i_10_138_4567_0, i_10_138_4568_0, i_10_138_4569_0;
  output o_10_138_0_0;
  assign o_10_138_0_0 = 0;
endmodule



// Benchmark "kernel_10_139" written by ABC on Sun Jul 19 10:23:22 2020

module kernel_10_139 ( 
    i_10_139_174_0, i_10_139_223_0, i_10_139_249_0, i_10_139_264_0,
    i_10_139_268_0, i_10_139_282_0, i_10_139_285_0, i_10_139_390_0,
    i_10_139_391_0, i_10_139_406_0, i_10_139_408_0, i_10_139_433_0,
    i_10_139_436_0, i_10_139_437_0, i_10_139_439_0, i_10_139_440_0,
    i_10_139_443_0, i_10_139_447_0, i_10_139_449_0, i_10_139_509_0,
    i_10_139_931_0, i_10_139_957_0, i_10_139_991_0, i_10_139_994_0,
    i_10_139_997_0, i_10_139_998_0, i_10_139_1002_0, i_10_139_1307_0,
    i_10_139_1308_0, i_10_139_1309_0, i_10_139_1349_0, i_10_139_1383_0,
    i_10_139_1435_0, i_10_139_1650_0, i_10_139_1654_0, i_10_139_1713_0,
    i_10_139_1823_0, i_10_139_1909_0, i_10_139_1910_0, i_10_139_1911_0,
    i_10_139_1912_0, i_10_139_1913_0, i_10_139_1915_0, i_10_139_2094_0,
    i_10_139_2184_0, i_10_139_2185_0, i_10_139_2201_0, i_10_139_2350_0,
    i_10_139_2361_0, i_10_139_2364_0, i_10_139_2451_0, i_10_139_2452_0,
    i_10_139_2464_0, i_10_139_2469_0, i_10_139_2508_0, i_10_139_2509_0,
    i_10_139_2604_0, i_10_139_2616_0, i_10_139_2617_0, i_10_139_2635_0,
    i_10_139_2680_0, i_10_139_2701_0, i_10_139_2705_0, i_10_139_2717_0,
    i_10_139_2731_0, i_10_139_2734_0, i_10_139_2817_0, i_10_139_2820_0,
    i_10_139_2821_0, i_10_139_2832_0, i_10_139_2885_0, i_10_139_2886_0,
    i_10_139_2887_0, i_10_139_2917_0, i_10_139_2919_0, i_10_139_3014_0,
    i_10_139_3195_0, i_10_139_3275_0, i_10_139_3281_0, i_10_139_3471_0,
    i_10_139_3472_0, i_10_139_3497_0, i_10_139_3706_0, i_10_139_3787_0,
    i_10_139_3837_0, i_10_139_3838_0, i_10_139_3850_0, i_10_139_3854_0,
    i_10_139_3859_0, i_10_139_3982_0, i_10_139_3984_0, i_10_139_3985_0,
    i_10_139_3986_0, i_10_139_4117_0, i_10_139_4118_0, i_10_139_4119_0,
    i_10_139_4236_0, i_10_139_4238_0, i_10_139_4533_0, i_10_139_4568_0,
    o_10_139_0_0  );
  input  i_10_139_174_0, i_10_139_223_0, i_10_139_249_0, i_10_139_264_0,
    i_10_139_268_0, i_10_139_282_0, i_10_139_285_0, i_10_139_390_0,
    i_10_139_391_0, i_10_139_406_0, i_10_139_408_0, i_10_139_433_0,
    i_10_139_436_0, i_10_139_437_0, i_10_139_439_0, i_10_139_440_0,
    i_10_139_443_0, i_10_139_447_0, i_10_139_449_0, i_10_139_509_0,
    i_10_139_931_0, i_10_139_957_0, i_10_139_991_0, i_10_139_994_0,
    i_10_139_997_0, i_10_139_998_0, i_10_139_1002_0, i_10_139_1307_0,
    i_10_139_1308_0, i_10_139_1309_0, i_10_139_1349_0, i_10_139_1383_0,
    i_10_139_1435_0, i_10_139_1650_0, i_10_139_1654_0, i_10_139_1713_0,
    i_10_139_1823_0, i_10_139_1909_0, i_10_139_1910_0, i_10_139_1911_0,
    i_10_139_1912_0, i_10_139_1913_0, i_10_139_1915_0, i_10_139_2094_0,
    i_10_139_2184_0, i_10_139_2185_0, i_10_139_2201_0, i_10_139_2350_0,
    i_10_139_2361_0, i_10_139_2364_0, i_10_139_2451_0, i_10_139_2452_0,
    i_10_139_2464_0, i_10_139_2469_0, i_10_139_2508_0, i_10_139_2509_0,
    i_10_139_2604_0, i_10_139_2616_0, i_10_139_2617_0, i_10_139_2635_0,
    i_10_139_2680_0, i_10_139_2701_0, i_10_139_2705_0, i_10_139_2717_0,
    i_10_139_2731_0, i_10_139_2734_0, i_10_139_2817_0, i_10_139_2820_0,
    i_10_139_2821_0, i_10_139_2832_0, i_10_139_2885_0, i_10_139_2886_0,
    i_10_139_2887_0, i_10_139_2917_0, i_10_139_2919_0, i_10_139_3014_0,
    i_10_139_3195_0, i_10_139_3275_0, i_10_139_3281_0, i_10_139_3471_0,
    i_10_139_3472_0, i_10_139_3497_0, i_10_139_3706_0, i_10_139_3787_0,
    i_10_139_3837_0, i_10_139_3838_0, i_10_139_3850_0, i_10_139_3854_0,
    i_10_139_3859_0, i_10_139_3982_0, i_10_139_3984_0, i_10_139_3985_0,
    i_10_139_3986_0, i_10_139_4117_0, i_10_139_4118_0, i_10_139_4119_0,
    i_10_139_4236_0, i_10_139_4238_0, i_10_139_4533_0, i_10_139_4568_0;
  output o_10_139_0_0;
  assign o_10_139_0_0 = ~((~i_10_139_264_0 & ((~i_10_139_268_0 & ((~i_10_139_439_0 & ~i_10_139_1002_0 & ~i_10_139_1349_0 & ~i_10_139_1915_0 & ~i_10_139_2184_0 & ~i_10_139_3195_0 & ~i_10_139_3859_0) | (~i_10_139_998_0 & ~i_10_139_1912_0 & ~i_10_139_2469_0 & ~i_10_139_2820_0 & i_10_139_3838_0 & ~i_10_139_3850_0 & i_10_139_3982_0 & ~i_10_139_4568_0))) | (~i_10_139_1909_0 & ~i_10_139_3854_0 & ((~i_10_139_390_0 & ~i_10_139_1913_0 & ~i_10_139_2469_0 & ~i_10_139_2508_0 & ~i_10_139_2734_0) | (~i_10_139_406_0 & ~i_10_139_1912_0 & ~i_10_139_1915_0 & ~i_10_139_2509_0 & ~i_10_139_2604_0 & ~i_10_139_2705_0 & ~i_10_139_3471_0 & ~i_10_139_4236_0))) | (~i_10_139_390_0 & ~i_10_139_2508_0 & ((~i_10_139_285_0 & ~i_10_139_1910_0 & ~i_10_139_2464_0 & ~i_10_139_2617_0 & ~i_10_139_2885_0 & ~i_10_139_3985_0) | (~i_10_139_2821_0 & ~i_10_139_3471_0 & ~i_10_139_3986_0))) | (~i_10_139_440_0 & ~i_10_139_998_0 & i_10_139_1309_0 & ~i_10_139_2616_0 & ~i_10_139_2821_0 & ~i_10_139_2885_0 & ~i_10_139_2887_0) | (~i_10_139_1912_0 & ~i_10_139_2201_0 & ~i_10_139_2361_0 & i_10_139_2451_0 & ~i_10_139_3982_0))) | (~i_10_139_3472_0 & ((~i_10_139_391_0 & ((~i_10_139_1307_0 & ~i_10_139_2201_0 & ~i_10_139_2508_0 & ~i_10_139_2616_0 & ~i_10_139_3195_0 & i_10_139_3982_0 & ~i_10_139_3984_0) | (~i_10_139_390_0 & ~i_10_139_408_0 & ~i_10_139_2734_0 & ~i_10_139_2886_0 & ~i_10_139_3281_0 & ~i_10_139_3837_0 & ~i_10_139_3854_0 & ~i_10_139_4118_0))) | (~i_10_139_2887_0 & ((~i_10_139_437_0 & ~i_10_139_2469_0 & ~i_10_139_3471_0 & ~i_10_139_3982_0) | (~i_10_139_449_0 & ~i_10_139_1915_0 & ~i_10_139_2201_0 & ~i_10_139_2451_0 & ~i_10_139_2617_0 & ~i_10_139_2820_0 & ~i_10_139_2821_0 & ~i_10_139_3850_0 & ~i_10_139_3984_0 & ~i_10_139_4119_0))))) | (~i_10_139_390_0 & ~i_10_139_3195_0 & ((~i_10_139_1307_0 & ~i_10_139_1912_0 & ~i_10_139_2185_0 & ~i_10_139_2604_0 & ~i_10_139_2717_0 & ~i_10_139_3984_0 & ~i_10_139_3985_0) | (i_10_139_439_0 & ~i_10_139_2452_0 & ~i_10_139_2509_0 & ~i_10_139_3838_0 & ~i_10_139_3986_0))) | (~i_10_139_2616_0 & ((~i_10_139_997_0 & ~i_10_139_1307_0 & ~i_10_139_1823_0 & i_10_139_2701_0 & i_10_139_2705_0 & ~i_10_139_3471_0) | (~i_10_139_1002_0 & ~i_10_139_2509_0 & ~i_10_139_2617_0 & ~i_10_139_2886_0 & ~i_10_139_2887_0 & ~i_10_139_3982_0 & ~i_10_139_3985_0))) | (i_10_139_4117_0 & ((~i_10_139_1308_0 & i_10_139_1654_0 & ~i_10_139_2452_0 & ~i_10_139_2919_0) | (~i_10_139_436_0 & ~i_10_139_3837_0))) | (~i_10_139_439_0 & ~i_10_139_3471_0 & ~i_10_139_3497_0 & ~i_10_139_3982_0));
endmodule



// Benchmark "kernel_10_140" written by ABC on Sun Jul 19 10:23:23 2020

module kernel_10_140 ( 
    i_10_140_29_0, i_10_140_117_0, i_10_140_124_0, i_10_140_154_0,
    i_10_140_181_0, i_10_140_182_0, i_10_140_183_0, i_10_140_219_0,
    i_10_140_253_0, i_10_140_257_0, i_10_140_261_0, i_10_140_264_0,
    i_10_140_318_0, i_10_140_410_0, i_10_140_427_0, i_10_140_460_0,
    i_10_140_461_0, i_10_140_463_0, i_10_140_464_0, i_10_140_904_0,
    i_10_140_946_0, i_10_140_949_0, i_10_140_958_0, i_10_140_959_0,
    i_10_140_1219_0, i_10_140_1246_0, i_10_140_1267_0, i_10_140_1297_0,
    i_10_140_1305_0, i_10_140_1306_0, i_10_140_1311_0, i_10_140_1313_0,
    i_10_140_1359_0, i_10_140_1361_0, i_10_140_1363_0, i_10_140_1364_0,
    i_10_140_1539_0, i_10_140_1540_0, i_10_140_1553_0, i_10_140_1683_0,
    i_10_140_1687_0, i_10_140_1940_0, i_10_140_1942_0, i_10_140_1980_0,
    i_10_140_2001_0, i_10_140_2202_0, i_10_140_2235_0, i_10_140_2304_0,
    i_10_140_2349_0, i_10_140_2350_0, i_10_140_2362_0, i_10_140_2376_0,
    i_10_140_2382_0, i_10_140_2383_0, i_10_140_2411_0, i_10_140_2448_0,
    i_10_140_2452_0, i_10_140_2453_0, i_10_140_2468_0, i_10_140_2514_0,
    i_10_140_2529_0, i_10_140_2530_0, i_10_140_2614_0, i_10_140_2615_0,
    i_10_140_2631_0, i_10_140_2636_0, i_10_140_2657_0, i_10_140_2738_0,
    i_10_140_2785_0, i_10_140_2832_0, i_10_140_2881_0, i_10_140_2920_0,
    i_10_140_2921_0, i_10_140_3073_0, i_10_140_3197_0, i_10_140_3278_0,
    i_10_140_3315_0, i_10_140_3408_0, i_10_140_3469_0, i_10_140_3609_0,
    i_10_140_3610_0, i_10_140_3611_0, i_10_140_3617_0, i_10_140_3647_0,
    i_10_140_3834_0, i_10_140_3838_0, i_10_140_3853_0, i_10_140_4050_0,
    i_10_140_4114_0, i_10_140_4117_0, i_10_140_4125_0, i_10_140_4129_0,
    i_10_140_4186_0, i_10_140_4217_0, i_10_140_4288_0, i_10_140_4289_0,
    i_10_140_4291_0, i_10_140_4563_0, i_10_140_4564_0, i_10_140_4567_0,
    o_10_140_0_0  );
  input  i_10_140_29_0, i_10_140_117_0, i_10_140_124_0, i_10_140_154_0,
    i_10_140_181_0, i_10_140_182_0, i_10_140_183_0, i_10_140_219_0,
    i_10_140_253_0, i_10_140_257_0, i_10_140_261_0, i_10_140_264_0,
    i_10_140_318_0, i_10_140_410_0, i_10_140_427_0, i_10_140_460_0,
    i_10_140_461_0, i_10_140_463_0, i_10_140_464_0, i_10_140_904_0,
    i_10_140_946_0, i_10_140_949_0, i_10_140_958_0, i_10_140_959_0,
    i_10_140_1219_0, i_10_140_1246_0, i_10_140_1267_0, i_10_140_1297_0,
    i_10_140_1305_0, i_10_140_1306_0, i_10_140_1311_0, i_10_140_1313_0,
    i_10_140_1359_0, i_10_140_1361_0, i_10_140_1363_0, i_10_140_1364_0,
    i_10_140_1539_0, i_10_140_1540_0, i_10_140_1553_0, i_10_140_1683_0,
    i_10_140_1687_0, i_10_140_1940_0, i_10_140_1942_0, i_10_140_1980_0,
    i_10_140_2001_0, i_10_140_2202_0, i_10_140_2235_0, i_10_140_2304_0,
    i_10_140_2349_0, i_10_140_2350_0, i_10_140_2362_0, i_10_140_2376_0,
    i_10_140_2382_0, i_10_140_2383_0, i_10_140_2411_0, i_10_140_2448_0,
    i_10_140_2452_0, i_10_140_2453_0, i_10_140_2468_0, i_10_140_2514_0,
    i_10_140_2529_0, i_10_140_2530_0, i_10_140_2614_0, i_10_140_2615_0,
    i_10_140_2631_0, i_10_140_2636_0, i_10_140_2657_0, i_10_140_2738_0,
    i_10_140_2785_0, i_10_140_2832_0, i_10_140_2881_0, i_10_140_2920_0,
    i_10_140_2921_0, i_10_140_3073_0, i_10_140_3197_0, i_10_140_3278_0,
    i_10_140_3315_0, i_10_140_3408_0, i_10_140_3469_0, i_10_140_3609_0,
    i_10_140_3610_0, i_10_140_3611_0, i_10_140_3617_0, i_10_140_3647_0,
    i_10_140_3834_0, i_10_140_3838_0, i_10_140_3853_0, i_10_140_4050_0,
    i_10_140_4114_0, i_10_140_4117_0, i_10_140_4125_0, i_10_140_4129_0,
    i_10_140_4186_0, i_10_140_4217_0, i_10_140_4288_0, i_10_140_4289_0,
    i_10_140_4291_0, i_10_140_4563_0, i_10_140_4564_0, i_10_140_4567_0;
  output o_10_140_0_0;
  assign o_10_140_0_0 = 0;
endmodule



// Benchmark "kernel_10_141" written by ABC on Sun Jul 19 10:23:23 2020

module kernel_10_141 ( 
    i_10_141_136_0, i_10_141_172_0, i_10_141_183_0, i_10_141_253_0,
    i_10_141_318_0, i_10_141_321_0, i_10_141_328_0, i_10_141_409_0,
    i_10_141_430_0, i_10_141_436_0, i_10_141_459_0, i_10_141_460_0,
    i_10_141_585_0, i_10_141_586_0, i_10_141_795_0, i_10_141_919_0,
    i_10_141_996_0, i_10_141_997_0, i_10_141_1039_0, i_10_141_1041_0,
    i_10_141_1042_0, i_10_141_1086_0, i_10_141_1087_0, i_10_141_1163_0,
    i_10_141_1238_0, i_10_141_1240_0, i_10_141_1241_0, i_10_141_1307_0,
    i_10_141_1308_0, i_10_141_1345_0, i_10_141_1361_0, i_10_141_1439_0,
    i_10_141_1551_0, i_10_141_1615_0, i_10_141_1630_0, i_10_141_1633_0,
    i_10_141_1651_0, i_10_141_1690_0, i_10_141_1691_0, i_10_141_1719_0,
    i_10_141_1729_0, i_10_141_1818_0, i_10_141_1873_0, i_10_141_1881_0,
    i_10_141_1911_0, i_10_141_2000_0, i_10_141_2233_0, i_10_141_2354_0,
    i_10_141_2407_0, i_10_141_2468_0, i_10_141_2473_0, i_10_141_2509_0,
    i_10_141_2566_0, i_10_141_2606_0, i_10_141_2718_0, i_10_141_2720_0,
    i_10_141_2787_0, i_10_141_2826_0, i_10_141_2827_0, i_10_141_2830_0,
    i_10_141_2833_0, i_10_141_2834_0, i_10_141_2908_0, i_10_141_2911_0,
    i_10_141_2920_0, i_10_141_3038_0, i_10_141_3070_0, i_10_141_3071_0,
    i_10_141_3116_0, i_10_141_3279_0, i_10_141_3406_0, i_10_141_3447_0,
    i_10_141_3587_0, i_10_141_3588_0, i_10_141_3589_0, i_10_141_3613_0,
    i_10_141_3615_0, i_10_141_3616_0, i_10_141_3622_0, i_10_141_3650_0,
    i_10_141_3774_0, i_10_141_3780_0, i_10_141_3782_0, i_10_141_3798_0,
    i_10_141_3840_0, i_10_141_3860_0, i_10_141_3891_0, i_10_141_3894_0,
    i_10_141_3895_0, i_10_141_4096_0, i_10_141_4115_0, i_10_141_4131_0,
    i_10_141_4230_0, i_10_141_4261_0, i_10_141_4312_0, i_10_141_4460_0,
    i_10_141_4519_0, i_10_141_4529_0, i_10_141_4567_0, i_10_141_4585_0,
    o_10_141_0_0  );
  input  i_10_141_136_0, i_10_141_172_0, i_10_141_183_0, i_10_141_253_0,
    i_10_141_318_0, i_10_141_321_0, i_10_141_328_0, i_10_141_409_0,
    i_10_141_430_0, i_10_141_436_0, i_10_141_459_0, i_10_141_460_0,
    i_10_141_585_0, i_10_141_586_0, i_10_141_795_0, i_10_141_919_0,
    i_10_141_996_0, i_10_141_997_0, i_10_141_1039_0, i_10_141_1041_0,
    i_10_141_1042_0, i_10_141_1086_0, i_10_141_1087_0, i_10_141_1163_0,
    i_10_141_1238_0, i_10_141_1240_0, i_10_141_1241_0, i_10_141_1307_0,
    i_10_141_1308_0, i_10_141_1345_0, i_10_141_1361_0, i_10_141_1439_0,
    i_10_141_1551_0, i_10_141_1615_0, i_10_141_1630_0, i_10_141_1633_0,
    i_10_141_1651_0, i_10_141_1690_0, i_10_141_1691_0, i_10_141_1719_0,
    i_10_141_1729_0, i_10_141_1818_0, i_10_141_1873_0, i_10_141_1881_0,
    i_10_141_1911_0, i_10_141_2000_0, i_10_141_2233_0, i_10_141_2354_0,
    i_10_141_2407_0, i_10_141_2468_0, i_10_141_2473_0, i_10_141_2509_0,
    i_10_141_2566_0, i_10_141_2606_0, i_10_141_2718_0, i_10_141_2720_0,
    i_10_141_2787_0, i_10_141_2826_0, i_10_141_2827_0, i_10_141_2830_0,
    i_10_141_2833_0, i_10_141_2834_0, i_10_141_2908_0, i_10_141_2911_0,
    i_10_141_2920_0, i_10_141_3038_0, i_10_141_3070_0, i_10_141_3071_0,
    i_10_141_3116_0, i_10_141_3279_0, i_10_141_3406_0, i_10_141_3447_0,
    i_10_141_3587_0, i_10_141_3588_0, i_10_141_3589_0, i_10_141_3613_0,
    i_10_141_3615_0, i_10_141_3616_0, i_10_141_3622_0, i_10_141_3650_0,
    i_10_141_3774_0, i_10_141_3780_0, i_10_141_3782_0, i_10_141_3798_0,
    i_10_141_3840_0, i_10_141_3860_0, i_10_141_3891_0, i_10_141_3894_0,
    i_10_141_3895_0, i_10_141_4096_0, i_10_141_4115_0, i_10_141_4131_0,
    i_10_141_4230_0, i_10_141_4261_0, i_10_141_4312_0, i_10_141_4460_0,
    i_10_141_4519_0, i_10_141_4529_0, i_10_141_4567_0, i_10_141_4585_0;
  output o_10_141_0_0;
  assign o_10_141_0_0 = 0;
endmodule



// Benchmark "kernel_10_142" written by ABC on Sun Jul 19 10:23:25 2020

module kernel_10_142 ( 
    i_10_142_171_0, i_10_142_175_0, i_10_142_279_0, i_10_142_280_0,
    i_10_142_281_0, i_10_142_282_0, i_10_142_283_0, i_10_142_284_0,
    i_10_142_286_0, i_10_142_429_0, i_10_142_445_0, i_10_142_460_0,
    i_10_142_506_0, i_10_142_517_0, i_10_142_518_0, i_10_142_519_0,
    i_10_142_794_0, i_10_142_799_0, i_10_142_967_0, i_10_142_968_0,
    i_10_142_1032_0, i_10_142_1037_0, i_10_142_1238_0, i_10_142_1349_0,
    i_10_142_1491_0, i_10_142_1550_0, i_10_142_1580_0, i_10_142_1650_0,
    i_10_142_1681_0, i_10_142_1686_0, i_10_142_1687_0, i_10_142_1688_0,
    i_10_142_1821_0, i_10_142_1822_0, i_10_142_1823_0, i_10_142_2001_0,
    i_10_142_2004_0, i_10_142_2152_0, i_10_142_2304_0, i_10_142_2305_0,
    i_10_142_2306_0, i_10_142_2351_0, i_10_142_2354_0, i_10_142_2364_0,
    i_10_142_2452_0, i_10_142_2467_0, i_10_142_2571_0, i_10_142_2630_0,
    i_10_142_2632_0, i_10_142_2655_0, i_10_142_2658_0, i_10_142_2659_0,
    i_10_142_2701_0, i_10_142_2715_0, i_10_142_2717_0, i_10_142_2721_0,
    i_10_142_2831_0, i_10_142_2883_0, i_10_142_2884_0, i_10_142_2920_0,
    i_10_142_2922_0, i_10_142_3043_0, i_10_142_3070_0, i_10_142_3071_0,
    i_10_142_3151_0, i_10_142_3165_0, i_10_142_3267_0, i_10_142_3270_0,
    i_10_142_3271_0, i_10_142_3280_0, i_10_142_3388_0, i_10_142_3389_0,
    i_10_142_3390_0, i_10_142_3404_0, i_10_142_3406_0, i_10_142_3408_0,
    i_10_142_3582_0, i_10_142_3612_0, i_10_142_3614_0, i_10_142_3784_0,
    i_10_142_3786_0, i_10_142_3787_0, i_10_142_3839_0, i_10_142_3841_0,
    i_10_142_3852_0, i_10_142_3853_0, i_10_142_3857_0, i_10_142_3889_0,
    i_10_142_3890_0, i_10_142_3912_0, i_10_142_3913_0, i_10_142_3914_0,
    i_10_142_4117_0, i_10_142_4130_0, i_10_142_4287_0, i_10_142_4288_0,
    i_10_142_4289_0, i_10_142_4290_0, i_10_142_4563_0, i_10_142_4570_0,
    o_10_142_0_0  );
  input  i_10_142_171_0, i_10_142_175_0, i_10_142_279_0, i_10_142_280_0,
    i_10_142_281_0, i_10_142_282_0, i_10_142_283_0, i_10_142_284_0,
    i_10_142_286_0, i_10_142_429_0, i_10_142_445_0, i_10_142_460_0,
    i_10_142_506_0, i_10_142_517_0, i_10_142_518_0, i_10_142_519_0,
    i_10_142_794_0, i_10_142_799_0, i_10_142_967_0, i_10_142_968_0,
    i_10_142_1032_0, i_10_142_1037_0, i_10_142_1238_0, i_10_142_1349_0,
    i_10_142_1491_0, i_10_142_1550_0, i_10_142_1580_0, i_10_142_1650_0,
    i_10_142_1681_0, i_10_142_1686_0, i_10_142_1687_0, i_10_142_1688_0,
    i_10_142_1821_0, i_10_142_1822_0, i_10_142_1823_0, i_10_142_2001_0,
    i_10_142_2004_0, i_10_142_2152_0, i_10_142_2304_0, i_10_142_2305_0,
    i_10_142_2306_0, i_10_142_2351_0, i_10_142_2354_0, i_10_142_2364_0,
    i_10_142_2452_0, i_10_142_2467_0, i_10_142_2571_0, i_10_142_2630_0,
    i_10_142_2632_0, i_10_142_2655_0, i_10_142_2658_0, i_10_142_2659_0,
    i_10_142_2701_0, i_10_142_2715_0, i_10_142_2717_0, i_10_142_2721_0,
    i_10_142_2831_0, i_10_142_2883_0, i_10_142_2884_0, i_10_142_2920_0,
    i_10_142_2922_0, i_10_142_3043_0, i_10_142_3070_0, i_10_142_3071_0,
    i_10_142_3151_0, i_10_142_3165_0, i_10_142_3267_0, i_10_142_3270_0,
    i_10_142_3271_0, i_10_142_3280_0, i_10_142_3388_0, i_10_142_3389_0,
    i_10_142_3390_0, i_10_142_3404_0, i_10_142_3406_0, i_10_142_3408_0,
    i_10_142_3582_0, i_10_142_3612_0, i_10_142_3614_0, i_10_142_3784_0,
    i_10_142_3786_0, i_10_142_3787_0, i_10_142_3839_0, i_10_142_3841_0,
    i_10_142_3852_0, i_10_142_3853_0, i_10_142_3857_0, i_10_142_3889_0,
    i_10_142_3890_0, i_10_142_3912_0, i_10_142_3913_0, i_10_142_3914_0,
    i_10_142_4117_0, i_10_142_4130_0, i_10_142_4287_0, i_10_142_4288_0,
    i_10_142_4289_0, i_10_142_4290_0, i_10_142_4563_0, i_10_142_4570_0;
  output o_10_142_0_0;
  assign o_10_142_0_0 = ~((i_10_142_171_0 & ((~i_10_142_460_0 & ~i_10_142_968_0 & ~i_10_142_1687_0 & ~i_10_142_2883_0 & ~i_10_142_3852_0 & ~i_10_142_3914_0) | (~i_10_142_1491_0 & ~i_10_142_2004_0 & ~i_10_142_3165_0 & ~i_10_142_3270_0 & ~i_10_142_3786_0 & ~i_10_142_3889_0 & ~i_10_142_3913_0 & ~i_10_142_4130_0))) | (~i_10_142_2305_0 & ((~i_10_142_171_0 & ((~i_10_142_519_0 & ~i_10_142_1688_0 & ~i_10_142_1822_0 & ~i_10_142_3784_0 & ~i_10_142_3890_0) | (~i_10_142_1032_0 & ~i_10_142_2632_0 & ~i_10_142_2658_0 & ~i_10_142_3165_0 & ~i_10_142_3280_0 & ~i_10_142_3388_0 & ~i_10_142_3612_0 & ~i_10_142_4130_0 & ~i_10_142_4287_0))) | (~i_10_142_967_0 & ~i_10_142_3913_0 & ((i_10_142_280_0 & i_10_142_794_0) | (~i_10_142_2004_0 & ~i_10_142_2883_0 & ~i_10_142_2884_0 & ~i_10_142_3165_0 & ~i_10_142_3267_0 & ~i_10_142_3271_0 & ~i_10_142_3389_0 & ~i_10_142_3890_0))) | (i_10_142_3852_0 & ~i_10_142_3912_0))) | (~i_10_142_175_0 & ((~i_10_142_2715_0 & ~i_10_142_2884_0 & i_10_142_2922_0 & ~i_10_142_3070_0 & ~i_10_142_3271_0 & ~i_10_142_3280_0 & ~i_10_142_3857_0 & ~i_10_142_3890_0) | (~i_10_142_1686_0 & i_10_142_2721_0 & ~i_10_142_3165_0 & ~i_10_142_3404_0 & ~i_10_142_3912_0))) | (i_10_142_284_0 & ((i_10_142_283_0 & ~i_10_142_967_0 & ~i_10_142_2571_0 & ~i_10_142_3404_0 & ~i_10_142_3912_0) | (~i_10_142_2452_0 & ~i_10_142_4290_0))) | (~i_10_142_3913_0 & ((~i_10_142_429_0 & ((i_10_142_518_0 & ~i_10_142_1037_0 & ~i_10_142_1550_0 & ~i_10_142_1650_0 & ~i_10_142_2452_0 & ~i_10_142_3839_0) | (i_10_142_2831_0 & ~i_10_142_2922_0 & ~i_10_142_3841_0 & ~i_10_142_3890_0))) | (~i_10_142_460_0 & ~i_10_142_517_0 & ~i_10_142_1686_0 & i_10_142_1823_0 & ~i_10_142_2004_0 & ~i_10_142_2831_0 & ~i_10_142_2920_0 & ~i_10_142_3271_0 & ~i_10_142_3890_0))) | (~i_10_142_3841_0 & ((~i_10_142_519_0 & ((~i_10_142_517_0 & ~i_10_142_1491_0 & ~i_10_142_1550_0 & ~i_10_142_1650_0 & ~i_10_142_1688_0 & ~i_10_142_2351_0 & ~i_10_142_2883_0 & ~i_10_142_3614_0 & ~i_10_142_3857_0 & ~i_10_142_3889_0) | (~i_10_142_968_0 & ~i_10_142_2452_0 & ~i_10_142_2884_0 & ~i_10_142_3280_0 & ~i_10_142_3406_0 & ~i_10_142_3582_0 & ~i_10_142_3787_0 & ~i_10_142_4563_0))) | (i_10_142_799_0 & ~i_10_142_1688_0 & ~i_10_142_1821_0 & ~i_10_142_1822_0 & ~i_10_142_3912_0 & ~i_10_142_4563_0))) | (~i_10_142_517_0 & ((~i_10_142_1650_0 & ~i_10_142_2004_0 & ~i_10_142_2571_0 & ~i_10_142_2701_0 & ~i_10_142_2715_0 & ~i_10_142_3388_0 & ~i_10_142_3857_0 & ~i_10_142_3889_0 & ~i_10_142_3914_0 & ~i_10_142_4130_0) | (~i_10_142_2884_0 & ~i_10_142_3271_0 & ~i_10_142_3390_0 & ~i_10_142_3912_0 & i_10_142_4287_0 & ~i_10_142_4289_0))) | (~i_10_142_794_0 & ((i_10_142_280_0 & ~i_10_142_2304_0) | (i_10_142_282_0 & ~i_10_142_1491_0 & ~i_10_142_2884_0 & ~i_10_142_4130_0))) | (~i_10_142_968_0 & ((~i_10_142_1491_0 & ~i_10_142_2304_0 & ~i_10_142_2883_0 & ~i_10_142_2920_0 & ~i_10_142_3280_0 & ~i_10_142_3839_0 & ~i_10_142_3889_0) | (~i_10_142_2884_0 & ~i_10_142_3614_0 & ~i_10_142_4130_0 & i_10_142_4287_0 & i_10_142_4289_0))) | (~i_10_142_1686_0 & ((~i_10_142_799_0 & ~i_10_142_1823_0 & ~i_10_142_2717_0 & ~i_10_142_3270_0 & i_10_142_3389_0) | (~i_10_142_2701_0 & ~i_10_142_2715_0 & ~i_10_142_2884_0 & i_10_142_3280_0 & ~i_10_142_3612_0))) | (~i_10_142_2883_0 & ((~i_10_142_2004_0 & ((i_10_142_3043_0 & ~i_10_142_3165_0) | (i_10_142_1686_0 & ~i_10_142_1821_0 & ~i_10_142_2701_0 & ~i_10_142_3071_0 & ~i_10_142_4570_0))) | (~i_10_142_1037_0 & i_10_142_1238_0 & ~i_10_142_1491_0 & ~i_10_142_2717_0 & ~i_10_142_3267_0))) | (~i_10_142_1491_0 & ((~i_10_142_1580_0 & ~i_10_142_3165_0 & ~i_10_142_3271_0 & i_10_142_3853_0 & ~i_10_142_3889_0 & ~i_10_142_3912_0) | (i_10_142_460_0 & ~i_10_142_967_0 & ~i_10_142_1687_0 & ~i_10_142_1688_0 & ~i_10_142_2884_0 & ~i_10_142_4289_0 & ~i_10_142_4290_0))) | (~i_10_142_279_0 & i_10_142_799_0 & ~i_10_142_1238_0 & i_10_142_3389_0 & ~i_10_142_3390_0 & i_10_142_4288_0 & ~i_10_142_4290_0));
endmodule



// Benchmark "kernel_10_143" written by ABC on Sun Jul 19 10:23:26 2020

module kernel_10_143 ( 
    i_10_143_173_0, i_10_143_176_0, i_10_143_245_0, i_10_143_272_0,
    i_10_143_275_0, i_10_143_283_0, i_10_143_316_0, i_10_143_317_0,
    i_10_143_319_0, i_10_143_320_0, i_10_143_391_0, i_10_143_413_0,
    i_10_143_434_0, i_10_143_445_0, i_10_143_461_0, i_10_143_464_0,
    i_10_143_716_0, i_10_143_749_0, i_10_143_752_0, i_10_143_794_0,
    i_10_143_797_0, i_10_143_892_0, i_10_143_893_0, i_10_143_992_0,
    i_10_143_995_0, i_10_143_1084_0, i_10_143_1154_0, i_10_143_1305_0,
    i_10_143_1310_0, i_10_143_1313_0, i_10_143_1342_0, i_10_143_1343_0,
    i_10_143_1346_0, i_10_143_1360_0, i_10_143_1361_0, i_10_143_1442_0,
    i_10_143_1622_0, i_10_143_1648_0, i_10_143_1652_0, i_10_143_1684_0,
    i_10_143_1685_0, i_10_143_1712_0, i_10_143_1823_0, i_10_143_1874_0,
    i_10_143_1916_0, i_10_143_1990_0, i_10_143_2017_0, i_10_143_2018_0,
    i_10_143_2198_0, i_10_143_2359_0, i_10_143_2381_0, i_10_143_2432_0,
    i_10_143_2468_0, i_10_143_2469_0, i_10_143_2470_0, i_10_143_2628_0,
    i_10_143_2630_0, i_10_143_2631_0, i_10_143_2632_0, i_10_143_2633_0,
    i_10_143_2636_0, i_10_143_2659_0, i_10_143_2674_0, i_10_143_2702_0,
    i_10_143_2711_0, i_10_143_2722_0, i_10_143_2782_0, i_10_143_2783_0,
    i_10_143_2827_0, i_10_143_2828_0, i_10_143_3044_0, i_10_143_3070_0,
    i_10_143_3071_0, i_10_143_3272_0, i_10_143_3278_0, i_10_143_3326_0,
    i_10_143_3328_0, i_10_143_3329_0, i_10_143_3392_0, i_10_143_3467_0,
    i_10_143_3523_0, i_10_143_3647_0, i_10_143_3837_0, i_10_143_3847_0,
    i_10_143_3848_0, i_10_143_3853_0, i_10_143_3854_0, i_10_143_3991_0,
    i_10_143_4114_0, i_10_143_4116_0, i_10_143_4117_0, i_10_143_4121_0,
    i_10_143_4127_0, i_10_143_4169_0, i_10_143_4276_0, i_10_143_4277_0,
    i_10_143_4286_0, i_10_143_4292_0, i_10_143_4568_0, i_10_143_4571_0,
    o_10_143_0_0  );
  input  i_10_143_173_0, i_10_143_176_0, i_10_143_245_0, i_10_143_272_0,
    i_10_143_275_0, i_10_143_283_0, i_10_143_316_0, i_10_143_317_0,
    i_10_143_319_0, i_10_143_320_0, i_10_143_391_0, i_10_143_413_0,
    i_10_143_434_0, i_10_143_445_0, i_10_143_461_0, i_10_143_464_0,
    i_10_143_716_0, i_10_143_749_0, i_10_143_752_0, i_10_143_794_0,
    i_10_143_797_0, i_10_143_892_0, i_10_143_893_0, i_10_143_992_0,
    i_10_143_995_0, i_10_143_1084_0, i_10_143_1154_0, i_10_143_1305_0,
    i_10_143_1310_0, i_10_143_1313_0, i_10_143_1342_0, i_10_143_1343_0,
    i_10_143_1346_0, i_10_143_1360_0, i_10_143_1361_0, i_10_143_1442_0,
    i_10_143_1622_0, i_10_143_1648_0, i_10_143_1652_0, i_10_143_1684_0,
    i_10_143_1685_0, i_10_143_1712_0, i_10_143_1823_0, i_10_143_1874_0,
    i_10_143_1916_0, i_10_143_1990_0, i_10_143_2017_0, i_10_143_2018_0,
    i_10_143_2198_0, i_10_143_2359_0, i_10_143_2381_0, i_10_143_2432_0,
    i_10_143_2468_0, i_10_143_2469_0, i_10_143_2470_0, i_10_143_2628_0,
    i_10_143_2630_0, i_10_143_2631_0, i_10_143_2632_0, i_10_143_2633_0,
    i_10_143_2636_0, i_10_143_2659_0, i_10_143_2674_0, i_10_143_2702_0,
    i_10_143_2711_0, i_10_143_2722_0, i_10_143_2782_0, i_10_143_2783_0,
    i_10_143_2827_0, i_10_143_2828_0, i_10_143_3044_0, i_10_143_3070_0,
    i_10_143_3071_0, i_10_143_3272_0, i_10_143_3278_0, i_10_143_3326_0,
    i_10_143_3328_0, i_10_143_3329_0, i_10_143_3392_0, i_10_143_3467_0,
    i_10_143_3523_0, i_10_143_3647_0, i_10_143_3837_0, i_10_143_3847_0,
    i_10_143_3848_0, i_10_143_3853_0, i_10_143_3854_0, i_10_143_3991_0,
    i_10_143_4114_0, i_10_143_4116_0, i_10_143_4117_0, i_10_143_4121_0,
    i_10_143_4127_0, i_10_143_4169_0, i_10_143_4276_0, i_10_143_4277_0,
    i_10_143_4286_0, i_10_143_4292_0, i_10_143_4568_0, i_10_143_4571_0;
  output o_10_143_0_0;
  assign o_10_143_0_0 = ~((~i_10_143_317_0 & ((~i_10_143_892_0 & ~i_10_143_1342_0 & ~i_10_143_1622_0 & ~i_10_143_1874_0 & ~i_10_143_1990_0 & ~i_10_143_3837_0 & ~i_10_143_3848_0 & ~i_10_143_4169_0) | (~i_10_143_1442_0 & i_10_143_4571_0))) | (~i_10_143_319_0 & ((~i_10_143_283_0 & ~i_10_143_995_0 & ~i_10_143_1990_0 & ~i_10_143_3071_0 & ~i_10_143_3837_0 & i_10_143_3991_0) | (~i_10_143_2782_0 & i_10_143_4114_0 & i_10_143_4116_0))) | (~i_10_143_391_0 & ((i_10_143_1342_0 & i_10_143_2631_0) | (~i_10_143_245_0 & ~i_10_143_1622_0 & i_10_143_1652_0 & ~i_10_143_2018_0 & ~i_10_143_2782_0))) | (~i_10_143_4169_0 & ((~i_10_143_2018_0 & ((~i_10_143_413_0 & ((i_10_143_1305_0 & ~i_10_143_1442_0 & ~i_10_143_2468_0) | (~i_10_143_1361_0 & ~i_10_143_2783_0 & ~i_10_143_3071_0 & i_10_143_3392_0))) | (~i_10_143_992_0 & ~i_10_143_2017_0 & ~i_10_143_2198_0 & ~i_10_143_2711_0 & ~i_10_143_3070_0 & ~i_10_143_3854_0))) | (~i_10_143_1084_0 & ((~i_10_143_1342_0 & i_10_143_1684_0 & ~i_10_143_2017_0 & ~i_10_143_2702_0 & ~i_10_143_2722_0 & ~i_10_143_2828_0 & ~i_10_143_3467_0 & ~i_10_143_4276_0) | (~i_10_143_1343_0 & ~i_10_143_1874_0 & ~i_10_143_1990_0 & ~i_10_143_3523_0 & ~i_10_143_3847_0 & ~i_10_143_3848_0 & ~i_10_143_4277_0))) | (~i_10_143_1346_0 & ~i_10_143_2017_0 & ~i_10_143_2702_0 & ~i_10_143_2711_0 & ~i_10_143_4117_0 & ~i_10_143_4277_0))) | (~i_10_143_1874_0 & ((i_10_143_2628_0 & ~i_10_143_3991_0 & ~i_10_143_4116_0 & ~i_10_143_4127_0 & ~i_10_143_4277_0) | (i_10_143_1823_0 & i_10_143_2631_0 & i_10_143_4292_0))) | (~i_10_143_1990_0 & ((i_10_143_319_0 & i_10_143_892_0 & i_10_143_3991_0) | (~i_10_143_316_0 & ~i_10_143_464_0 & ~i_10_143_1310_0 & ~i_10_143_2018_0 & ~i_10_143_2468_0 & ~i_10_143_3071_0 & ~i_10_143_3647_0 & ~i_10_143_3837_0 & ~i_10_143_4116_0 & ~i_10_143_4127_0))) | (i_10_143_2632_0 & ~i_10_143_3991_0 & ((~i_10_143_316_0 & i_10_143_2722_0 & ~i_10_143_4116_0) | (~i_10_143_320_0 & i_10_143_2631_0 & i_10_143_4286_0))) | (~i_10_143_316_0 & ((~i_10_143_1346_0 & ~i_10_143_2017_0 & ~i_10_143_2711_0 & ~i_10_143_3071_0 & ~i_10_143_4277_0) | (i_10_143_3991_0 & i_10_143_4292_0))) | (i_10_143_391_0 & i_10_143_2470_0 & ~i_10_143_2702_0 & ~i_10_143_4276_0 & ~i_10_143_4277_0));
endmodule



// Benchmark "kernel_10_144" written by ABC on Sun Jul 19 10:23:27 2020

module kernel_10_144 ( 
    i_10_144_145_0, i_10_144_177_0, i_10_144_246_0, i_10_144_252_0,
    i_10_144_282_0, i_10_144_315_0, i_10_144_316_0, i_10_144_322_0,
    i_10_144_327_0, i_10_144_443_0, i_10_144_444_0, i_10_144_498_0,
    i_10_144_501_0, i_10_144_504_0, i_10_144_505_0, i_10_144_508_0,
    i_10_144_712_0, i_10_144_1059_0, i_10_144_1084_0, i_10_144_1236_0,
    i_10_144_1239_0, i_10_144_1241_0, i_10_144_1299_0, i_10_144_1302_0,
    i_10_144_1312_0, i_10_144_1363_0, i_10_144_1434_0, i_10_144_1444_0,
    i_10_144_1542_0, i_10_144_1576_0, i_10_144_1578_0, i_10_144_1618_0,
    i_10_144_1623_0, i_10_144_1686_0, i_10_144_1688_0, i_10_144_1689_0,
    i_10_144_1731_0, i_10_144_1734_0, i_10_144_1803_0, i_10_144_1820_0,
    i_10_144_1822_0, i_10_144_1823_0, i_10_144_1978_0, i_10_144_2028_0,
    i_10_144_2031_0, i_10_144_2202_0, i_10_144_2376_0, i_10_144_2451_0,
    i_10_144_2455_0, i_10_144_2466_0, i_10_144_2469_0, i_10_144_2470_0,
    i_10_144_2472_0, i_10_144_2568_0, i_10_144_2700_0, i_10_144_2715_0,
    i_10_144_2721_0, i_10_144_2725_0, i_10_144_2733_0, i_10_144_2826_0,
    i_10_144_2832_0, i_10_144_2964_0, i_10_144_2967_0, i_10_144_3196_0,
    i_10_144_3268_0, i_10_144_3277_0, i_10_144_3279_0, i_10_144_3281_0,
    i_10_144_3282_0, i_10_144_3283_0, i_10_144_3315_0, i_10_144_3318_0,
    i_10_144_3325_0, i_10_144_3327_0, i_10_144_3385_0, i_10_144_3501_0,
    i_10_144_3504_0, i_10_144_3543_0, i_10_144_3544_0, i_10_144_3582_0,
    i_10_144_3585_0, i_10_144_3588_0, i_10_144_3646_0, i_10_144_3651_0,
    i_10_144_3781_0, i_10_144_3795_0, i_10_144_3840_0, i_10_144_3909_0,
    i_10_144_4030_0, i_10_144_4114_0, i_10_144_4119_0, i_10_144_4266_0,
    i_10_144_4269_0, i_10_144_4272_0, i_10_144_4281_0, i_10_144_4290_0,
    i_10_144_4548_0, i_10_144_4567_0, i_10_144_4570_0, i_10_144_4585_0,
    o_10_144_0_0  );
  input  i_10_144_145_0, i_10_144_177_0, i_10_144_246_0, i_10_144_252_0,
    i_10_144_282_0, i_10_144_315_0, i_10_144_316_0, i_10_144_322_0,
    i_10_144_327_0, i_10_144_443_0, i_10_144_444_0, i_10_144_498_0,
    i_10_144_501_0, i_10_144_504_0, i_10_144_505_0, i_10_144_508_0,
    i_10_144_712_0, i_10_144_1059_0, i_10_144_1084_0, i_10_144_1236_0,
    i_10_144_1239_0, i_10_144_1241_0, i_10_144_1299_0, i_10_144_1302_0,
    i_10_144_1312_0, i_10_144_1363_0, i_10_144_1434_0, i_10_144_1444_0,
    i_10_144_1542_0, i_10_144_1576_0, i_10_144_1578_0, i_10_144_1618_0,
    i_10_144_1623_0, i_10_144_1686_0, i_10_144_1688_0, i_10_144_1689_0,
    i_10_144_1731_0, i_10_144_1734_0, i_10_144_1803_0, i_10_144_1820_0,
    i_10_144_1822_0, i_10_144_1823_0, i_10_144_1978_0, i_10_144_2028_0,
    i_10_144_2031_0, i_10_144_2202_0, i_10_144_2376_0, i_10_144_2451_0,
    i_10_144_2455_0, i_10_144_2466_0, i_10_144_2469_0, i_10_144_2470_0,
    i_10_144_2472_0, i_10_144_2568_0, i_10_144_2700_0, i_10_144_2715_0,
    i_10_144_2721_0, i_10_144_2725_0, i_10_144_2733_0, i_10_144_2826_0,
    i_10_144_2832_0, i_10_144_2964_0, i_10_144_2967_0, i_10_144_3196_0,
    i_10_144_3268_0, i_10_144_3277_0, i_10_144_3279_0, i_10_144_3281_0,
    i_10_144_3282_0, i_10_144_3283_0, i_10_144_3315_0, i_10_144_3318_0,
    i_10_144_3325_0, i_10_144_3327_0, i_10_144_3385_0, i_10_144_3501_0,
    i_10_144_3504_0, i_10_144_3543_0, i_10_144_3544_0, i_10_144_3582_0,
    i_10_144_3585_0, i_10_144_3588_0, i_10_144_3646_0, i_10_144_3651_0,
    i_10_144_3781_0, i_10_144_3795_0, i_10_144_3840_0, i_10_144_3909_0,
    i_10_144_4030_0, i_10_144_4114_0, i_10_144_4119_0, i_10_144_4266_0,
    i_10_144_4269_0, i_10_144_4272_0, i_10_144_4281_0, i_10_144_4290_0,
    i_10_144_4548_0, i_10_144_4567_0, i_10_144_4570_0, i_10_144_4585_0;
  output o_10_144_0_0;
  assign o_10_144_0_0 = ~((~i_10_144_145_0 & ((~i_10_144_1434_0 & ((~i_10_144_2715_0 & ~i_10_144_3282_0 & ~i_10_144_3283_0 & ~i_10_144_3501_0) | (~i_10_144_443_0 & ~i_10_144_1734_0 & ~i_10_144_2721_0 & ~i_10_144_2733_0 & ~i_10_144_3504_0 & ~i_10_144_4266_0))) | (~i_10_144_177_0 & ~i_10_144_282_0 & ~i_10_144_1731_0 & ~i_10_144_3646_0 & ~i_10_144_4114_0 & ~i_10_144_4272_0))) | (~i_10_144_1444_0 & ((i_10_144_1236_0 & ~i_10_144_1689_0 & ~i_10_144_1822_0 & ~i_10_144_2725_0 & ~i_10_144_3385_0 & ~i_10_144_3504_0 & ~i_10_144_4030_0) | (~i_10_144_2715_0 & ~i_10_144_3268_0 & ~i_10_144_3585_0 & ~i_10_144_4272_0))) | (~i_10_144_1618_0 & ((~i_10_144_1689_0 & ~i_10_144_2451_0 & ~i_10_144_2466_0 & ~i_10_144_3543_0 & ~i_10_144_4119_0) | (i_10_144_2472_0 & i_10_144_2733_0 & ~i_10_144_3281_0 & ~i_10_144_3282_0 & ~i_10_144_4266_0 & ~i_10_144_4281_0))) | (~i_10_144_1822_0 & ((i_10_144_282_0 & i_10_144_1578_0 & ~i_10_144_3283_0 & ~i_10_144_3501_0 & ~i_10_144_3504_0) | (~i_10_144_443_0 & ~i_10_144_712_0 & ~i_10_144_2028_0 & ~i_10_144_2202_0 & ~i_10_144_3196_0 & ~i_10_144_3315_0 & ~i_10_144_3318_0 & ~i_10_144_3543_0))) | (~i_10_144_1241_0 & ((~i_10_144_443_0 & ~i_10_144_3501_0 & ((~i_10_144_1084_0 & ~i_10_144_1542_0 & ~i_10_144_1689_0 & ~i_10_144_3196_0 & ~i_10_144_3543_0) | (~i_10_144_1734_0 & ~i_10_144_2568_0 & ~i_10_144_2721_0 & ~i_10_144_3315_0 & ~i_10_144_3504_0 & ~i_10_144_4269_0))) | (~i_10_144_3277_0 & ~i_10_144_3283_0 & i_10_144_4030_0 & ~i_10_144_4290_0))) | (~i_10_144_1734_0 & ~i_10_144_3909_0 & ((~i_10_144_2469_0 & ~i_10_144_3582_0 & ~i_10_144_4272_0) | (~i_10_144_444_0 & i_10_144_1241_0 & ~i_10_144_3279_0 & ~i_10_144_3282_0 & ~i_10_144_3501_0 & ~i_10_144_4266_0 & ~i_10_144_4290_0))) | (i_10_144_1820_0 & ((~i_10_144_3279_0 & ((~i_10_144_1686_0 & ~i_10_144_1688_0 & ~i_10_144_2466_0) | (i_10_144_3781_0 & ~i_10_144_4281_0))) | (i_10_144_1084_0 & ~i_10_144_1236_0))) | (~i_10_144_2028_0 & ~i_10_144_2469_0 & ~i_10_144_2721_0 & ~i_10_144_2725_0 & ~i_10_144_3585_0) | (~i_10_144_2715_0 & ~i_10_144_3282_0 & ~i_10_144_3385_0 & ~i_10_144_3582_0 & ~i_10_144_3588_0));
endmodule



// Benchmark "kernel_10_145" written by ABC on Sun Jul 19 10:23:28 2020

module kernel_10_145 ( 
    i_10_145_21_0, i_10_145_22_0, i_10_145_58_0, i_10_145_89_0,
    i_10_145_181_0, i_10_145_213_0, i_10_145_277_0, i_10_145_280_0,
    i_10_145_388_0, i_10_145_445_0, i_10_145_500_0, i_10_145_507_0,
    i_10_145_584_0, i_10_145_595_0, i_10_145_597_0, i_10_145_598_0,
    i_10_145_659_0, i_10_145_679_0, i_10_145_729_0, i_10_145_967_0,
    i_10_145_1011_0, i_10_145_1187_0, i_10_145_1201_0, i_10_145_1326_0,
    i_10_145_1327_0, i_10_145_1345_0, i_10_145_1366_0, i_10_145_1444_0,
    i_10_145_1480_0, i_10_145_1488_0, i_10_145_1526_0, i_10_145_1536_0,
    i_10_145_1543_0, i_10_145_1548_0, i_10_145_1614_0, i_10_145_1624_0,
    i_10_145_1651_0, i_10_145_1652_0, i_10_145_1713_0, i_10_145_1750_0,
    i_10_145_1761_0, i_10_145_1789_0, i_10_145_1826_0, i_10_145_1875_0,
    i_10_145_1919_0, i_10_145_1930_0, i_10_145_2001_0, i_10_145_2152_0,
    i_10_145_2226_0, i_10_145_2227_0, i_10_145_2272_0, i_10_145_2507_0,
    i_10_145_2601_0, i_10_145_2604_0, i_10_145_2653_0, i_10_145_2667_0,
    i_10_145_2668_0, i_10_145_2732_0, i_10_145_2767_0, i_10_145_2803_0,
    i_10_145_2877_0, i_10_145_2879_0, i_10_145_2953_0, i_10_145_2963_0,
    i_10_145_3028_0, i_10_145_3029_0, i_10_145_3040_0, i_10_145_3043_0,
    i_10_145_3057_0, i_10_145_3135_0, i_10_145_3189_0, i_10_145_3190_0,
    i_10_145_3191_0, i_10_145_3201_0, i_10_145_3224_0, i_10_145_3297_0,
    i_10_145_3402_0, i_10_145_3403_0, i_10_145_3544_0, i_10_145_3604_0,
    i_10_145_3610_0, i_10_145_3616_0, i_10_145_3723_0, i_10_145_3724_0,
    i_10_145_3729_0, i_10_145_3838_0, i_10_145_3863_0, i_10_145_3922_0,
    i_10_145_3975_0, i_10_145_4068_0, i_10_145_4069_0, i_10_145_4182_0,
    i_10_145_4218_0, i_10_145_4407_0, i_10_145_4446_0, i_10_145_4447_0,
    i_10_145_4455_0, i_10_145_4459_0, i_10_145_4516_0, i_10_145_4517_0,
    o_10_145_0_0  );
  input  i_10_145_21_0, i_10_145_22_0, i_10_145_58_0, i_10_145_89_0,
    i_10_145_181_0, i_10_145_213_0, i_10_145_277_0, i_10_145_280_0,
    i_10_145_388_0, i_10_145_445_0, i_10_145_500_0, i_10_145_507_0,
    i_10_145_584_0, i_10_145_595_0, i_10_145_597_0, i_10_145_598_0,
    i_10_145_659_0, i_10_145_679_0, i_10_145_729_0, i_10_145_967_0,
    i_10_145_1011_0, i_10_145_1187_0, i_10_145_1201_0, i_10_145_1326_0,
    i_10_145_1327_0, i_10_145_1345_0, i_10_145_1366_0, i_10_145_1444_0,
    i_10_145_1480_0, i_10_145_1488_0, i_10_145_1526_0, i_10_145_1536_0,
    i_10_145_1543_0, i_10_145_1548_0, i_10_145_1614_0, i_10_145_1624_0,
    i_10_145_1651_0, i_10_145_1652_0, i_10_145_1713_0, i_10_145_1750_0,
    i_10_145_1761_0, i_10_145_1789_0, i_10_145_1826_0, i_10_145_1875_0,
    i_10_145_1919_0, i_10_145_1930_0, i_10_145_2001_0, i_10_145_2152_0,
    i_10_145_2226_0, i_10_145_2227_0, i_10_145_2272_0, i_10_145_2507_0,
    i_10_145_2601_0, i_10_145_2604_0, i_10_145_2653_0, i_10_145_2667_0,
    i_10_145_2668_0, i_10_145_2732_0, i_10_145_2767_0, i_10_145_2803_0,
    i_10_145_2877_0, i_10_145_2879_0, i_10_145_2953_0, i_10_145_2963_0,
    i_10_145_3028_0, i_10_145_3029_0, i_10_145_3040_0, i_10_145_3043_0,
    i_10_145_3057_0, i_10_145_3135_0, i_10_145_3189_0, i_10_145_3190_0,
    i_10_145_3191_0, i_10_145_3201_0, i_10_145_3224_0, i_10_145_3297_0,
    i_10_145_3402_0, i_10_145_3403_0, i_10_145_3544_0, i_10_145_3604_0,
    i_10_145_3610_0, i_10_145_3616_0, i_10_145_3723_0, i_10_145_3724_0,
    i_10_145_3729_0, i_10_145_3838_0, i_10_145_3863_0, i_10_145_3922_0,
    i_10_145_3975_0, i_10_145_4068_0, i_10_145_4069_0, i_10_145_4182_0,
    i_10_145_4218_0, i_10_145_4407_0, i_10_145_4446_0, i_10_145_4447_0,
    i_10_145_4455_0, i_10_145_4459_0, i_10_145_4516_0, i_10_145_4517_0;
  output o_10_145_0_0;
  assign o_10_145_0_0 = 0;
endmodule



// Benchmark "kernel_10_146" written by ABC on Sun Jul 19 10:23:29 2020

module kernel_10_146 ( 
    i_10_146_43_0, i_10_146_176_0, i_10_146_178_0, i_10_146_283_0,
    i_10_146_284_0, i_10_146_287_0, i_10_146_293_0, i_10_146_315_0,
    i_10_146_316_0, i_10_146_317_0, i_10_146_390_0, i_10_146_426_0,
    i_10_146_429_0, i_10_146_435_0, i_10_146_436_0, i_10_146_445_0,
    i_10_146_499_0, i_10_146_588_0, i_10_146_589_0, i_10_146_693_0,
    i_10_146_694_0, i_10_146_928_0, i_10_146_990_0, i_10_146_991_0,
    i_10_146_1033_0, i_10_146_1233_0, i_10_146_1234_0, i_10_146_1235_0,
    i_10_146_1238_0, i_10_146_1309_0, i_10_146_1310_0, i_10_146_1445_0,
    i_10_146_1541_0, i_10_146_1581_0, i_10_146_1685_0, i_10_146_1688_0,
    i_10_146_1764_0, i_10_146_1821_0, i_10_146_1823_0, i_10_146_1909_0,
    i_10_146_1910_0, i_10_146_2353_0, i_10_146_2449_0, i_10_146_2451_0,
    i_10_146_2452_0, i_10_146_2460_0, i_10_146_2463_0, i_10_146_2467_0,
    i_10_146_2468_0, i_10_146_2514_0, i_10_146_2634_0, i_10_146_2733_0,
    i_10_146_2817_0, i_10_146_2831_0, i_10_146_2880_0, i_10_146_2881_0,
    i_10_146_2883_0, i_10_146_2884_0, i_10_146_2919_0, i_10_146_2920_0,
    i_10_146_2921_0, i_10_146_2979_0, i_10_146_2980_0, i_10_146_3090_0,
    i_10_146_3091_0, i_10_146_3159_0, i_10_146_3169_0, i_10_146_3199_0,
    i_10_146_3200_0, i_10_146_3356_0, i_10_146_3388_0, i_10_146_3445_0,
    i_10_146_3446_0, i_10_146_3519_0, i_10_146_3520_0, i_10_146_3522_0,
    i_10_146_3613_0, i_10_146_3614_0, i_10_146_3699_0, i_10_146_3703_0,
    i_10_146_3826_0, i_10_146_3850_0, i_10_146_3853_0, i_10_146_3889_0,
    i_10_146_3890_0, i_10_146_3898_0, i_10_146_3899_0, i_10_146_3905_0,
    i_10_146_3906_0, i_10_146_3984_0, i_10_146_4026_0, i_10_146_4028_0,
    i_10_146_4031_0, i_10_146_4052_0, i_10_146_4097_0, i_10_146_4216_0,
    i_10_146_4531_0, i_10_146_4591_0, i_10_146_4592_0, i_10_146_4594_0,
    o_10_146_0_0  );
  input  i_10_146_43_0, i_10_146_176_0, i_10_146_178_0, i_10_146_283_0,
    i_10_146_284_0, i_10_146_287_0, i_10_146_293_0, i_10_146_315_0,
    i_10_146_316_0, i_10_146_317_0, i_10_146_390_0, i_10_146_426_0,
    i_10_146_429_0, i_10_146_435_0, i_10_146_436_0, i_10_146_445_0,
    i_10_146_499_0, i_10_146_588_0, i_10_146_589_0, i_10_146_693_0,
    i_10_146_694_0, i_10_146_928_0, i_10_146_990_0, i_10_146_991_0,
    i_10_146_1033_0, i_10_146_1233_0, i_10_146_1234_0, i_10_146_1235_0,
    i_10_146_1238_0, i_10_146_1309_0, i_10_146_1310_0, i_10_146_1445_0,
    i_10_146_1541_0, i_10_146_1581_0, i_10_146_1685_0, i_10_146_1688_0,
    i_10_146_1764_0, i_10_146_1821_0, i_10_146_1823_0, i_10_146_1909_0,
    i_10_146_1910_0, i_10_146_2353_0, i_10_146_2449_0, i_10_146_2451_0,
    i_10_146_2452_0, i_10_146_2460_0, i_10_146_2463_0, i_10_146_2467_0,
    i_10_146_2468_0, i_10_146_2514_0, i_10_146_2634_0, i_10_146_2733_0,
    i_10_146_2817_0, i_10_146_2831_0, i_10_146_2880_0, i_10_146_2881_0,
    i_10_146_2883_0, i_10_146_2884_0, i_10_146_2919_0, i_10_146_2920_0,
    i_10_146_2921_0, i_10_146_2979_0, i_10_146_2980_0, i_10_146_3090_0,
    i_10_146_3091_0, i_10_146_3159_0, i_10_146_3169_0, i_10_146_3199_0,
    i_10_146_3200_0, i_10_146_3356_0, i_10_146_3388_0, i_10_146_3445_0,
    i_10_146_3446_0, i_10_146_3519_0, i_10_146_3520_0, i_10_146_3522_0,
    i_10_146_3613_0, i_10_146_3614_0, i_10_146_3699_0, i_10_146_3703_0,
    i_10_146_3826_0, i_10_146_3850_0, i_10_146_3853_0, i_10_146_3889_0,
    i_10_146_3890_0, i_10_146_3898_0, i_10_146_3899_0, i_10_146_3905_0,
    i_10_146_3906_0, i_10_146_3984_0, i_10_146_4026_0, i_10_146_4028_0,
    i_10_146_4031_0, i_10_146_4052_0, i_10_146_4097_0, i_10_146_4216_0,
    i_10_146_4531_0, i_10_146_4591_0, i_10_146_4592_0, i_10_146_4594_0;
  output o_10_146_0_0;
  assign o_10_146_0_0 = 0;
endmodule



// Benchmark "kernel_10_147" written by ABC on Sun Jul 19 10:23:30 2020

module kernel_10_147 ( 
    i_10_147_176_0, i_10_147_218_0, i_10_147_221_0, i_10_147_270_0,
    i_10_147_275_0, i_10_147_285_0, i_10_147_319_0, i_10_147_435_0,
    i_10_147_442_0, i_10_147_464_0, i_10_147_506_0, i_10_147_507_0,
    i_10_147_955_0, i_10_147_956_0, i_10_147_959_0, i_10_147_961_0,
    i_10_147_1027_0, i_10_147_1028_0, i_10_147_1030_0, i_10_147_1031_0,
    i_10_147_1034_0, i_10_147_1086_0, i_10_147_1087_0, i_10_147_1134_0,
    i_10_147_1141_0, i_10_147_1237_0, i_10_147_1246_0, i_10_147_1307_0,
    i_10_147_1308_0, i_10_147_1540_0, i_10_147_1541_0, i_10_147_1543_0,
    i_10_147_1552_0, i_10_147_1553_0, i_10_147_1580_0, i_10_147_1649_0,
    i_10_147_1691_0, i_10_147_1820_0, i_10_147_1826_0, i_10_147_1994_0,
    i_10_147_2201_0, i_10_147_2204_0, i_10_147_2358_0, i_10_147_2363_0,
    i_10_147_2365_0, i_10_147_2461_0, i_10_147_2464_0, i_10_147_2466_0,
    i_10_147_2470_0, i_10_147_2628_0, i_10_147_2663_0, i_10_147_2674_0,
    i_10_147_2678_0, i_10_147_2700_0, i_10_147_2701_0, i_10_147_2722_0,
    i_10_147_2723_0, i_10_147_2833_0, i_10_147_2834_0, i_10_147_2885_0,
    i_10_147_2924_0, i_10_147_3196_0, i_10_147_3197_0, i_10_147_3199_0,
    i_10_147_3202_0, i_10_147_3203_0, i_10_147_3268_0, i_10_147_3280_0,
    i_10_147_3323_0, i_10_147_3392_0, i_10_147_3403_0, i_10_147_3466_0,
    i_10_147_3469_0, i_10_147_3470_0, i_10_147_3522_0, i_10_147_3583_0,
    i_10_147_3586_0, i_10_147_3587_0, i_10_147_3589_0, i_10_147_3731_0,
    i_10_147_3781_0, i_10_147_3782_0, i_10_147_3784_0, i_10_147_3785_0,
    i_10_147_3786_0, i_10_147_3787_0, i_10_147_3788_0, i_10_147_3844_0,
    i_10_147_3849_0, i_10_147_3854_0, i_10_147_3856_0, i_10_147_3857_0,
    i_10_147_3859_0, i_10_147_3860_0, i_10_147_3979_0, i_10_147_3980_0,
    i_10_147_3982_0, i_10_147_4121_0, i_10_147_4291_0, i_10_147_4567_0,
    o_10_147_0_0  );
  input  i_10_147_176_0, i_10_147_218_0, i_10_147_221_0, i_10_147_270_0,
    i_10_147_275_0, i_10_147_285_0, i_10_147_319_0, i_10_147_435_0,
    i_10_147_442_0, i_10_147_464_0, i_10_147_506_0, i_10_147_507_0,
    i_10_147_955_0, i_10_147_956_0, i_10_147_959_0, i_10_147_961_0,
    i_10_147_1027_0, i_10_147_1028_0, i_10_147_1030_0, i_10_147_1031_0,
    i_10_147_1034_0, i_10_147_1086_0, i_10_147_1087_0, i_10_147_1134_0,
    i_10_147_1141_0, i_10_147_1237_0, i_10_147_1246_0, i_10_147_1307_0,
    i_10_147_1308_0, i_10_147_1540_0, i_10_147_1541_0, i_10_147_1543_0,
    i_10_147_1552_0, i_10_147_1553_0, i_10_147_1580_0, i_10_147_1649_0,
    i_10_147_1691_0, i_10_147_1820_0, i_10_147_1826_0, i_10_147_1994_0,
    i_10_147_2201_0, i_10_147_2204_0, i_10_147_2358_0, i_10_147_2363_0,
    i_10_147_2365_0, i_10_147_2461_0, i_10_147_2464_0, i_10_147_2466_0,
    i_10_147_2470_0, i_10_147_2628_0, i_10_147_2663_0, i_10_147_2674_0,
    i_10_147_2678_0, i_10_147_2700_0, i_10_147_2701_0, i_10_147_2722_0,
    i_10_147_2723_0, i_10_147_2833_0, i_10_147_2834_0, i_10_147_2885_0,
    i_10_147_2924_0, i_10_147_3196_0, i_10_147_3197_0, i_10_147_3199_0,
    i_10_147_3202_0, i_10_147_3203_0, i_10_147_3268_0, i_10_147_3280_0,
    i_10_147_3323_0, i_10_147_3392_0, i_10_147_3403_0, i_10_147_3466_0,
    i_10_147_3469_0, i_10_147_3470_0, i_10_147_3522_0, i_10_147_3583_0,
    i_10_147_3586_0, i_10_147_3587_0, i_10_147_3589_0, i_10_147_3731_0,
    i_10_147_3781_0, i_10_147_3782_0, i_10_147_3784_0, i_10_147_3785_0,
    i_10_147_3786_0, i_10_147_3787_0, i_10_147_3788_0, i_10_147_3844_0,
    i_10_147_3849_0, i_10_147_3854_0, i_10_147_3856_0, i_10_147_3857_0,
    i_10_147_3859_0, i_10_147_3860_0, i_10_147_3979_0, i_10_147_3980_0,
    i_10_147_3982_0, i_10_147_4121_0, i_10_147_4291_0, i_10_147_4567_0;
  output o_10_147_0_0;
  assign o_10_147_0_0 = ~((~i_10_147_221_0 & ~i_10_147_2365_0 & ((~i_10_147_176_0 & ~i_10_147_319_0 & ~i_10_147_955_0 & ~i_10_147_1031_0 & ~i_10_147_3522_0 & ~i_10_147_3583_0 & ~i_10_147_3849_0) | (~i_10_147_1028_0 & ~i_10_147_1541_0 & ~i_10_147_3788_0 & ~i_10_147_3854_0))) | (~i_10_147_176_0 & ((~i_10_147_956_0 & ~i_10_147_1691_0 & ~i_10_147_2924_0 & ~i_10_147_3782_0 & ~i_10_147_3857_0) | (~i_10_147_1246_0 & i_10_147_2201_0 & ~i_10_147_3787_0 & i_10_147_3857_0 & ~i_10_147_3860_0))) | (~i_10_147_955_0 & ((~i_10_147_956_0 & ~i_10_147_1034_0 & ~i_10_147_2201_0 & ~i_10_147_2461_0 & ~i_10_147_3392_0 & ~i_10_147_3844_0) | (~i_10_147_2464_0 & i_10_147_3586_0 & i_10_147_3982_0))) | (~i_10_147_1027_0 & ~i_10_147_3196_0 & ((~i_10_147_1543_0 & ~i_10_147_1580_0 & ~i_10_147_2464_0 & ~i_10_147_2663_0 & ~i_10_147_3202_0 & ~i_10_147_3403_0) | (~i_10_147_3392_0 & ~i_10_147_3857_0 & i_10_147_4291_0))) | (~i_10_147_1031_0 & ((~i_10_147_1030_0 & ((~i_10_147_956_0 & ~i_10_147_3787_0 & ~i_10_147_3788_0) | (~i_10_147_1541_0 & ~i_10_147_1691_0 & i_10_147_3202_0 & ~i_10_147_4291_0))) | (i_10_147_1030_0 & ~i_10_147_1580_0 & i_10_147_2363_0 & ~i_10_147_2461_0))) | (~i_10_147_3403_0 & ((~i_10_147_1246_0 & ((~i_10_147_464_0 & ~i_10_147_1691_0 & ~i_10_147_3199_0 & ~i_10_147_3203_0 & ~i_10_147_3587_0 & ~i_10_147_3844_0) | (~i_10_147_285_0 & ~i_10_147_1553_0 & ~i_10_147_3786_0 & ~i_10_147_3787_0 & ~i_10_147_3788_0 & i_10_147_3854_0 & ~i_10_147_3980_0))) | (~i_10_147_442_0 & ~i_10_147_1543_0 & ~i_10_147_2201_0 & ~i_10_147_2204_0 & ~i_10_147_2663_0 & i_10_147_3202_0))) | (~i_10_147_1553_0 & ~i_10_147_3784_0 & ((~i_10_147_1541_0 & i_10_147_1691_0 & ~i_10_147_2363_0 & ~i_10_147_2461_0 & ~i_10_147_2722_0 & ~i_10_147_3466_0 & ~i_10_147_3844_0) | (~i_10_147_218_0 & ~i_10_147_2358_0 & i_10_147_2924_0 & ~i_10_147_3280_0 & ~i_10_147_3860_0 & i_10_147_4291_0))) | (~i_10_147_3787_0 & ((~i_10_147_1580_0 & i_10_147_2628_0 & ~i_10_147_2663_0 & ~i_10_147_3392_0) | (~i_10_147_2924_0 & ~i_10_147_3587_0 & i_10_147_3980_0))));
endmodule



// Benchmark "kernel_10_148" written by ABC on Sun Jul 19 10:23:31 2020

module kernel_10_148 ( 
    i_10_148_178_0, i_10_148_283_0, i_10_148_327_0, i_10_148_406_0,
    i_10_148_429_0, i_10_148_446_0, i_10_148_461_0, i_10_148_463_0,
    i_10_148_464_0, i_10_148_465_0, i_10_148_466_0, i_10_148_467_0,
    i_10_148_498_0, i_10_148_795_0, i_10_148_796_0, i_10_148_994_0,
    i_10_148_1123_0, i_10_148_1236_0, i_10_148_1237_0, i_10_148_1238_0,
    i_10_148_1240_0, i_10_148_1241_0, i_10_148_1491_0, i_10_148_1575_0,
    i_10_148_1650_0, i_10_148_1651_0, i_10_148_1683_0, i_10_148_1685_0,
    i_10_148_1689_0, i_10_148_1690_0, i_10_148_1914_0, i_10_148_1915_0,
    i_10_148_1948_0, i_10_148_2001_0, i_10_148_2005_0, i_10_148_2028_0,
    i_10_148_2244_0, i_10_148_2351_0, i_10_148_2353_0, i_10_148_2355_0,
    i_10_148_2356_0, i_10_148_2357_0, i_10_148_2359_0, i_10_148_2362_0,
    i_10_148_2363_0, i_10_148_2364_0, i_10_148_2451_0, i_10_148_2452_0,
    i_10_148_2453_0, i_10_148_2466_0, i_10_148_2478_0, i_10_148_2515_0,
    i_10_148_2565_0, i_10_148_2571_0, i_10_148_2677_0, i_10_148_2728_0,
    i_10_148_2781_0, i_10_148_2784_0, i_10_148_2823_0, i_10_148_2826_0,
    i_10_148_2827_0, i_10_148_2828_0, i_10_148_2869_0, i_10_148_3271_0,
    i_10_148_3273_0, i_10_148_3278_0, i_10_148_3279_0, i_10_148_3280_0,
    i_10_148_3281_0, i_10_148_3282_0, i_10_148_3283_0, i_10_148_3328_0,
    i_10_148_3430_0, i_10_148_3466_0, i_10_148_3471_0, i_10_148_3544_0,
    i_10_148_3582_0, i_10_148_3585_0, i_10_148_3586_0, i_10_148_3587_0,
    i_10_148_3590_0, i_10_148_3610_0, i_10_148_3684_0, i_10_148_3685_0,
    i_10_148_3721_0, i_10_148_3781_0, i_10_148_3788_0, i_10_148_3845_0,
    i_10_148_3983_0, i_10_148_4114_0, i_10_148_4119_0, i_10_148_4120_0,
    i_10_148_4128_0, i_10_148_4174_0, i_10_148_4269_0, i_10_148_4272_0,
    i_10_148_4287_0, i_10_148_4290_0, i_10_148_4291_0, i_10_148_4584_0,
    o_10_148_0_0  );
  input  i_10_148_178_0, i_10_148_283_0, i_10_148_327_0, i_10_148_406_0,
    i_10_148_429_0, i_10_148_446_0, i_10_148_461_0, i_10_148_463_0,
    i_10_148_464_0, i_10_148_465_0, i_10_148_466_0, i_10_148_467_0,
    i_10_148_498_0, i_10_148_795_0, i_10_148_796_0, i_10_148_994_0,
    i_10_148_1123_0, i_10_148_1236_0, i_10_148_1237_0, i_10_148_1238_0,
    i_10_148_1240_0, i_10_148_1241_0, i_10_148_1491_0, i_10_148_1575_0,
    i_10_148_1650_0, i_10_148_1651_0, i_10_148_1683_0, i_10_148_1685_0,
    i_10_148_1689_0, i_10_148_1690_0, i_10_148_1914_0, i_10_148_1915_0,
    i_10_148_1948_0, i_10_148_2001_0, i_10_148_2005_0, i_10_148_2028_0,
    i_10_148_2244_0, i_10_148_2351_0, i_10_148_2353_0, i_10_148_2355_0,
    i_10_148_2356_0, i_10_148_2357_0, i_10_148_2359_0, i_10_148_2362_0,
    i_10_148_2363_0, i_10_148_2364_0, i_10_148_2451_0, i_10_148_2452_0,
    i_10_148_2453_0, i_10_148_2466_0, i_10_148_2478_0, i_10_148_2515_0,
    i_10_148_2565_0, i_10_148_2571_0, i_10_148_2677_0, i_10_148_2728_0,
    i_10_148_2781_0, i_10_148_2784_0, i_10_148_2823_0, i_10_148_2826_0,
    i_10_148_2827_0, i_10_148_2828_0, i_10_148_2869_0, i_10_148_3271_0,
    i_10_148_3273_0, i_10_148_3278_0, i_10_148_3279_0, i_10_148_3280_0,
    i_10_148_3281_0, i_10_148_3282_0, i_10_148_3283_0, i_10_148_3328_0,
    i_10_148_3430_0, i_10_148_3466_0, i_10_148_3471_0, i_10_148_3544_0,
    i_10_148_3582_0, i_10_148_3585_0, i_10_148_3586_0, i_10_148_3587_0,
    i_10_148_3590_0, i_10_148_3610_0, i_10_148_3684_0, i_10_148_3685_0,
    i_10_148_3721_0, i_10_148_3781_0, i_10_148_3788_0, i_10_148_3845_0,
    i_10_148_3983_0, i_10_148_4114_0, i_10_148_4119_0, i_10_148_4120_0,
    i_10_148_4128_0, i_10_148_4174_0, i_10_148_4269_0, i_10_148_4272_0,
    i_10_148_4287_0, i_10_148_4290_0, i_10_148_4291_0, i_10_148_4584_0;
  output o_10_148_0_0;
  assign o_10_148_0_0 = 0;
endmodule



// Benchmark "kernel_10_149" written by ABC on Sun Jul 19 10:23:32 2020

module kernel_10_149 ( 
    i_10_149_29_0, i_10_149_86_0, i_10_149_122_0, i_10_149_280_0,
    i_10_149_435_0, i_10_149_438_0, i_10_149_503_0, i_10_149_585_0,
    i_10_149_739_0, i_10_149_751_0, i_10_149_800_0, i_10_149_853_0,
    i_10_149_854_0, i_10_149_930_0, i_10_149_995_0, i_10_149_1006_0,
    i_10_149_1054_0, i_10_149_1223_0, i_10_149_1234_0, i_10_149_1239_0,
    i_10_149_1354_0, i_10_149_1579_0, i_10_149_1733_0, i_10_149_1736_0,
    i_10_149_1807_0, i_10_149_1819_0, i_10_149_1914_0, i_10_149_1916_0,
    i_10_149_1919_0, i_10_149_1925_0, i_10_149_1981_0, i_10_149_1995_0,
    i_10_149_1996_0, i_10_149_2002_0, i_10_149_2093_0, i_10_149_2096_0,
    i_10_149_2306_0, i_10_149_2354_0, i_10_149_2362_0, i_10_149_2452_0,
    i_10_149_2470_0, i_10_149_2475_0, i_10_149_2542_0, i_10_149_2543_0,
    i_10_149_2567_0, i_10_149_2573_0, i_10_149_2629_0, i_10_149_2641_0,
    i_10_149_2704_0, i_10_149_2724_0, i_10_149_2725_0, i_10_149_2801_0,
    i_10_149_2828_0, i_10_149_2831_0, i_10_149_2882_0, i_10_149_2883_0,
    i_10_149_2884_0, i_10_149_2917_0, i_10_149_2919_0, i_10_149_3082_0,
    i_10_149_3088_0, i_10_149_3090_0, i_10_149_3091_0, i_10_149_3124_0,
    i_10_149_3173_0, i_10_149_3278_0, i_10_149_3281_0, i_10_149_3353_0,
    i_10_149_3385_0, i_10_149_3406_0, i_10_149_3407_0, i_10_149_3409_0,
    i_10_149_3465_0, i_10_149_3473_0, i_10_149_3508_0, i_10_149_3586_0,
    i_10_149_3612_0, i_10_149_3650_0, i_10_149_3685_0, i_10_149_3686_0,
    i_10_149_3702_0, i_10_149_3748_0, i_10_149_3786_0, i_10_149_3832_0,
    i_10_149_3834_0, i_10_149_3849_0, i_10_149_3853_0, i_10_149_3901_0,
    i_10_149_3984_0, i_10_149_3988_0, i_10_149_4029_0, i_10_149_4030_0,
    i_10_149_4128_0, i_10_149_4130_0, i_10_149_4211_0, i_10_149_4216_0,
    i_10_149_4236_0, i_10_149_4272_0, i_10_149_4289_0, i_10_149_4566_0,
    o_10_149_0_0  );
  input  i_10_149_29_0, i_10_149_86_0, i_10_149_122_0, i_10_149_280_0,
    i_10_149_435_0, i_10_149_438_0, i_10_149_503_0, i_10_149_585_0,
    i_10_149_739_0, i_10_149_751_0, i_10_149_800_0, i_10_149_853_0,
    i_10_149_854_0, i_10_149_930_0, i_10_149_995_0, i_10_149_1006_0,
    i_10_149_1054_0, i_10_149_1223_0, i_10_149_1234_0, i_10_149_1239_0,
    i_10_149_1354_0, i_10_149_1579_0, i_10_149_1733_0, i_10_149_1736_0,
    i_10_149_1807_0, i_10_149_1819_0, i_10_149_1914_0, i_10_149_1916_0,
    i_10_149_1919_0, i_10_149_1925_0, i_10_149_1981_0, i_10_149_1995_0,
    i_10_149_1996_0, i_10_149_2002_0, i_10_149_2093_0, i_10_149_2096_0,
    i_10_149_2306_0, i_10_149_2354_0, i_10_149_2362_0, i_10_149_2452_0,
    i_10_149_2470_0, i_10_149_2475_0, i_10_149_2542_0, i_10_149_2543_0,
    i_10_149_2567_0, i_10_149_2573_0, i_10_149_2629_0, i_10_149_2641_0,
    i_10_149_2704_0, i_10_149_2724_0, i_10_149_2725_0, i_10_149_2801_0,
    i_10_149_2828_0, i_10_149_2831_0, i_10_149_2882_0, i_10_149_2883_0,
    i_10_149_2884_0, i_10_149_2917_0, i_10_149_2919_0, i_10_149_3082_0,
    i_10_149_3088_0, i_10_149_3090_0, i_10_149_3091_0, i_10_149_3124_0,
    i_10_149_3173_0, i_10_149_3278_0, i_10_149_3281_0, i_10_149_3353_0,
    i_10_149_3385_0, i_10_149_3406_0, i_10_149_3407_0, i_10_149_3409_0,
    i_10_149_3465_0, i_10_149_3473_0, i_10_149_3508_0, i_10_149_3586_0,
    i_10_149_3612_0, i_10_149_3650_0, i_10_149_3685_0, i_10_149_3686_0,
    i_10_149_3702_0, i_10_149_3748_0, i_10_149_3786_0, i_10_149_3832_0,
    i_10_149_3834_0, i_10_149_3849_0, i_10_149_3853_0, i_10_149_3901_0,
    i_10_149_3984_0, i_10_149_3988_0, i_10_149_4029_0, i_10_149_4030_0,
    i_10_149_4128_0, i_10_149_4130_0, i_10_149_4211_0, i_10_149_4216_0,
    i_10_149_4236_0, i_10_149_4272_0, i_10_149_4289_0, i_10_149_4566_0;
  output o_10_149_0_0;
  assign o_10_149_0_0 = 0;
endmodule



// Benchmark "kernel_10_150" written by ABC on Sun Jul 19 10:23:33 2020

module kernel_10_150 ( 
    i_10_150_263_0, i_10_150_280_0, i_10_150_282_0, i_10_150_327_0,
    i_10_150_393_0, i_10_150_411_0, i_10_150_438_0, i_10_150_509_0,
    i_10_150_511_0, i_10_150_512_0, i_10_150_718_0, i_10_150_961_0,
    i_10_150_1026_0, i_10_150_1035_0, i_10_150_1135_0, i_10_150_1239_0,
    i_10_150_1431_0, i_10_150_1576_0, i_10_150_1683_0, i_10_150_1684_0,
    i_10_150_1686_0, i_10_150_1689_0, i_10_150_1690_0, i_10_150_1821_0,
    i_10_150_1822_0, i_10_150_1825_0, i_10_150_1980_0, i_10_150_1998_0,
    i_10_150_2001_0, i_10_150_2006_0, i_10_150_2025_0, i_10_150_2028_0,
    i_10_150_2032_0, i_10_150_2199_0, i_10_150_2361_0, i_10_150_2362_0,
    i_10_150_2364_0, i_10_150_2365_0, i_10_150_2407_0, i_10_150_2452_0,
    i_10_150_2461_0, i_10_150_2466_0, i_10_150_2469_0, i_10_150_2506_0,
    i_10_150_2630_0, i_10_150_2658_0, i_10_150_2659_0, i_10_150_2680_0,
    i_10_150_2700_0, i_10_150_2701_0, i_10_150_2703_0, i_10_150_2704_0,
    i_10_150_2716_0, i_10_150_2718_0, i_10_150_2719_0, i_10_150_2727_0,
    i_10_150_2730_0, i_10_150_2733_0, i_10_150_2734_0, i_10_150_2785_0,
    i_10_150_2788_0, i_10_150_2827_0, i_10_150_2831_0, i_10_150_2885_0,
    i_10_150_3037_0, i_10_150_3153_0, i_10_150_3154_0, i_10_150_3195_0,
    i_10_150_3196_0, i_10_150_3198_0, i_10_150_3277_0, i_10_150_3279_0,
    i_10_150_3280_0, i_10_150_3283_0, i_10_150_3312_0, i_10_150_3386_0,
    i_10_150_3388_0, i_10_150_3391_0, i_10_150_3465_0, i_10_150_3468_0,
    i_10_150_3507_0, i_10_150_3588_0, i_10_150_3646_0, i_10_150_3647_0,
    i_10_150_3650_0, i_10_150_3684_0, i_10_150_3783_0, i_10_150_3786_0,
    i_10_150_3840_0, i_10_150_3846_0, i_10_150_3982_0, i_10_150_3983_0,
    i_10_150_4116_0, i_10_150_4117_0, i_10_150_4120_0, i_10_150_4126_0,
    i_10_150_4266_0, i_10_150_4281_0, i_10_150_4290_0, i_10_150_4570_0,
    o_10_150_0_0  );
  input  i_10_150_263_0, i_10_150_280_0, i_10_150_282_0, i_10_150_327_0,
    i_10_150_393_0, i_10_150_411_0, i_10_150_438_0, i_10_150_509_0,
    i_10_150_511_0, i_10_150_512_0, i_10_150_718_0, i_10_150_961_0,
    i_10_150_1026_0, i_10_150_1035_0, i_10_150_1135_0, i_10_150_1239_0,
    i_10_150_1431_0, i_10_150_1576_0, i_10_150_1683_0, i_10_150_1684_0,
    i_10_150_1686_0, i_10_150_1689_0, i_10_150_1690_0, i_10_150_1821_0,
    i_10_150_1822_0, i_10_150_1825_0, i_10_150_1980_0, i_10_150_1998_0,
    i_10_150_2001_0, i_10_150_2006_0, i_10_150_2025_0, i_10_150_2028_0,
    i_10_150_2032_0, i_10_150_2199_0, i_10_150_2361_0, i_10_150_2362_0,
    i_10_150_2364_0, i_10_150_2365_0, i_10_150_2407_0, i_10_150_2452_0,
    i_10_150_2461_0, i_10_150_2466_0, i_10_150_2469_0, i_10_150_2506_0,
    i_10_150_2630_0, i_10_150_2658_0, i_10_150_2659_0, i_10_150_2680_0,
    i_10_150_2700_0, i_10_150_2701_0, i_10_150_2703_0, i_10_150_2704_0,
    i_10_150_2716_0, i_10_150_2718_0, i_10_150_2719_0, i_10_150_2727_0,
    i_10_150_2730_0, i_10_150_2733_0, i_10_150_2734_0, i_10_150_2785_0,
    i_10_150_2788_0, i_10_150_2827_0, i_10_150_2831_0, i_10_150_2885_0,
    i_10_150_3037_0, i_10_150_3153_0, i_10_150_3154_0, i_10_150_3195_0,
    i_10_150_3196_0, i_10_150_3198_0, i_10_150_3277_0, i_10_150_3279_0,
    i_10_150_3280_0, i_10_150_3283_0, i_10_150_3312_0, i_10_150_3386_0,
    i_10_150_3388_0, i_10_150_3391_0, i_10_150_3465_0, i_10_150_3468_0,
    i_10_150_3507_0, i_10_150_3588_0, i_10_150_3646_0, i_10_150_3647_0,
    i_10_150_3650_0, i_10_150_3684_0, i_10_150_3783_0, i_10_150_3786_0,
    i_10_150_3840_0, i_10_150_3846_0, i_10_150_3982_0, i_10_150_3983_0,
    i_10_150_4116_0, i_10_150_4117_0, i_10_150_4120_0, i_10_150_4126_0,
    i_10_150_4266_0, i_10_150_4281_0, i_10_150_4290_0, i_10_150_4570_0;
  output o_10_150_0_0;
  assign o_10_150_0_0 = ~((i_10_150_263_0 & ((~i_10_150_2785_0 & i_10_150_3650_0) | (i_10_150_2407_0 & ~i_10_150_4266_0))) | (~i_10_150_1026_0 & ((~i_10_150_393_0 & ~i_10_150_1576_0 & ~i_10_150_1683_0 & ~i_10_150_2199_0 & ~i_10_150_2785_0 & ~i_10_150_3283_0 & ~i_10_150_3388_0 & ~i_10_150_3465_0) | (~i_10_150_1684_0 & ~i_10_150_2452_0 & ~i_10_150_2469_0 & ~i_10_150_3391_0 & ~i_10_150_3840_0))) | (~i_10_150_2469_0 & ((~i_10_150_393_0 & ((i_10_150_1825_0 & ~i_10_150_2001_0 & ~i_10_150_2006_0 & ~i_10_150_3312_0 & ~i_10_150_3465_0 & ~i_10_150_3588_0) | (~i_10_150_1686_0 & ~i_10_150_1690_0 & ~i_10_150_3507_0 & ~i_10_150_3983_0 & ~i_10_150_4116_0 & ~i_10_150_4266_0 & ~i_10_150_4281_0))) | (~i_10_150_1998_0 & ~i_10_150_2831_0 & ((~i_10_150_718_0 & i_10_150_1821_0 & i_10_150_1822_0 & ~i_10_150_2199_0 & ~i_10_150_3283_0 & ~i_10_150_3386_0 & ~i_10_150_3646_0 & ~i_10_150_3840_0 & ~i_10_150_4266_0) | (~i_10_150_2006_0 & ~i_10_150_2466_0 & ~i_10_150_2734_0 & ~i_10_150_3037_0 & ~i_10_150_3507_0 & ~i_10_150_4281_0))) | (~i_10_150_438_0 & ~i_10_150_2025_0 & ~i_10_150_2032_0 & ~i_10_150_2716_0 & i_10_150_3037_0))) | (~i_10_150_4281_0 & ((~i_10_150_1431_0 & ((~i_10_150_1689_0 & ~i_10_150_2032_0 & ~i_10_150_2466_0 & ~i_10_150_3283_0) | (i_10_150_280_0 & ~i_10_150_1576_0 & ~i_10_150_1822_0 & ~i_10_150_2727_0 & ~i_10_150_3465_0))) | (~i_10_150_1689_0 & ~i_10_150_2452_0 & ~i_10_150_2703_0 & ~i_10_150_2719_0 & ~i_10_150_2727_0 & ~i_10_150_2733_0 & ~i_10_150_3846_0) | (~i_10_150_1998_0 & ~i_10_150_2716_0 & ~i_10_150_3312_0 & ~i_10_150_3391_0 & ~i_10_150_3507_0 & i_10_150_3588_0 & ~i_10_150_3840_0 & ~i_10_150_4126_0))) | (~i_10_150_1689_0 & ((i_10_150_1821_0 & i_10_150_2630_0) | (~i_10_150_1239_0 & ~i_10_150_1686_0 & ~i_10_150_2032_0 & ~i_10_150_2659_0 & ~i_10_150_3280_0 & ~i_10_150_3312_0 & ~i_10_150_3468_0))) | (~i_10_150_2730_0 & ((~i_10_150_1684_0 & i_10_150_3386_0 & ~i_10_150_3588_0) | (i_10_150_3037_0 & ~i_10_150_3507_0 & i_10_150_3982_0 & ~i_10_150_3983_0 & i_10_150_4117_0))) | (~i_10_150_3279_0 & ((~i_10_150_2733_0 & ((i_10_150_438_0 & ~i_10_150_2659_0) | (~i_10_150_1998_0 & ~i_10_150_2831_0 & ~i_10_150_3277_0 & ~i_10_150_3312_0 & ~i_10_150_3588_0))) | (i_10_150_2658_0 & ~i_10_150_4120_0 & i_10_150_4290_0) | (~i_10_150_1822_0 & ~i_10_150_2630_0 & ~i_10_150_2701_0 & ~i_10_150_3386_0 & ~i_10_150_3983_0 & ~i_10_150_4266_0 & ~i_10_150_4290_0))) | (~i_10_150_3283_0 & ((i_10_150_2452_0 & ~i_10_150_2727_0 & ~i_10_150_3650_0 & i_10_150_3982_0) | (~i_10_150_2006_0 & i_10_150_3037_0 & ~i_10_150_3507_0 & ~i_10_150_3840_0 & i_10_150_4281_0))) | (~i_10_150_2006_0 & ((~i_10_150_961_0 & ~i_10_150_2025_0 & ~i_10_150_2028_0 & i_10_150_2701_0 & ~i_10_150_3391_0 & ~i_10_150_3684_0 & ~i_10_150_4120_0) | (i_10_150_2885_0 & i_10_150_3198_0 & ~i_10_150_3840_0 & ~i_10_150_4290_0))) | (i_10_150_2407_0 & ~i_10_150_2452_0 & ~i_10_150_3280_0 & ~i_10_150_4290_0) | (~i_10_150_2199_0 & i_10_150_3388_0 & ~i_10_150_4117_0 & i_10_150_4120_0));
endmodule



// Benchmark "kernel_10_151" written by ABC on Sun Jul 19 10:23:35 2020

module kernel_10_151 ( 
    i_10_151_48_0, i_10_151_82_0, i_10_151_216_0, i_10_151_219_0,
    i_10_151_245_0, i_10_151_270_0, i_10_151_280_0, i_10_151_281_0,
    i_10_151_282_0, i_10_151_283_0, i_10_151_322_0, i_10_151_405_0,
    i_10_151_424_0, i_10_151_435_0, i_10_151_436_0, i_10_151_459_0,
    i_10_151_460_0, i_10_151_467_0, i_10_151_891_0, i_10_151_902_0,
    i_10_151_1026_0, i_10_151_1163_0, i_10_151_1236_0, i_10_151_1263_0,
    i_10_151_1307_0, i_10_151_1432_0, i_10_151_1433_0, i_10_151_1441_0,
    i_10_151_1444_0, i_10_151_1485_0, i_10_151_1539_0, i_10_151_1540_0,
    i_10_151_1579_0, i_10_151_1652_0, i_10_151_1687_0, i_10_151_1688_0,
    i_10_151_1767_0, i_10_151_1768_0, i_10_151_1824_0, i_10_151_1825_0,
    i_10_151_1826_0, i_10_151_1911_0, i_10_151_1912_0, i_10_151_2200_0,
    i_10_151_2325_0, i_10_151_2351_0, i_10_151_2449_0, i_10_151_2628_0,
    i_10_151_2631_0, i_10_151_2637_0, i_10_151_2655_0, i_10_151_2656_0,
    i_10_151_2658_0, i_10_151_2659_0, i_10_151_2660_0, i_10_151_2673_0,
    i_10_151_2674_0, i_10_151_2700_0, i_10_151_2702_0, i_10_151_2718_0,
    i_10_151_2719_0, i_10_151_2720_0, i_10_151_2721_0, i_10_151_2722_0,
    i_10_151_2723_0, i_10_151_2729_0, i_10_151_2781_0, i_10_151_2826_0,
    i_10_151_2884_0, i_10_151_2885_0, i_10_151_2921_0, i_10_151_2985_0,
    i_10_151_3033_0, i_10_151_3045_0, i_10_151_3070_0, i_10_151_3071_0,
    i_10_151_3154_0, i_10_151_3159_0, i_10_151_3196_0, i_10_151_3326_0,
    i_10_151_3388_0, i_10_151_3391_0, i_10_151_3405_0, i_10_151_3470_0,
    i_10_151_3522_0, i_10_151_3523_0, i_10_151_3645_0, i_10_151_3682_0,
    i_10_151_3782_0, i_10_151_3847_0, i_10_151_3855_0, i_10_151_3856_0,
    i_10_151_3857_0, i_10_151_3906_0, i_10_151_3907_0, i_10_151_3979_0,
    i_10_151_4117_0, i_10_151_4118_0, i_10_151_4123_0, i_10_151_4287_0,
    o_10_151_0_0  );
  input  i_10_151_48_0, i_10_151_82_0, i_10_151_216_0, i_10_151_219_0,
    i_10_151_245_0, i_10_151_270_0, i_10_151_280_0, i_10_151_281_0,
    i_10_151_282_0, i_10_151_283_0, i_10_151_322_0, i_10_151_405_0,
    i_10_151_424_0, i_10_151_435_0, i_10_151_436_0, i_10_151_459_0,
    i_10_151_460_0, i_10_151_467_0, i_10_151_891_0, i_10_151_902_0,
    i_10_151_1026_0, i_10_151_1163_0, i_10_151_1236_0, i_10_151_1263_0,
    i_10_151_1307_0, i_10_151_1432_0, i_10_151_1433_0, i_10_151_1441_0,
    i_10_151_1444_0, i_10_151_1485_0, i_10_151_1539_0, i_10_151_1540_0,
    i_10_151_1579_0, i_10_151_1652_0, i_10_151_1687_0, i_10_151_1688_0,
    i_10_151_1767_0, i_10_151_1768_0, i_10_151_1824_0, i_10_151_1825_0,
    i_10_151_1826_0, i_10_151_1911_0, i_10_151_1912_0, i_10_151_2200_0,
    i_10_151_2325_0, i_10_151_2351_0, i_10_151_2449_0, i_10_151_2628_0,
    i_10_151_2631_0, i_10_151_2637_0, i_10_151_2655_0, i_10_151_2656_0,
    i_10_151_2658_0, i_10_151_2659_0, i_10_151_2660_0, i_10_151_2673_0,
    i_10_151_2674_0, i_10_151_2700_0, i_10_151_2702_0, i_10_151_2718_0,
    i_10_151_2719_0, i_10_151_2720_0, i_10_151_2721_0, i_10_151_2722_0,
    i_10_151_2723_0, i_10_151_2729_0, i_10_151_2781_0, i_10_151_2826_0,
    i_10_151_2884_0, i_10_151_2885_0, i_10_151_2921_0, i_10_151_2985_0,
    i_10_151_3033_0, i_10_151_3045_0, i_10_151_3070_0, i_10_151_3071_0,
    i_10_151_3154_0, i_10_151_3159_0, i_10_151_3196_0, i_10_151_3326_0,
    i_10_151_3388_0, i_10_151_3391_0, i_10_151_3405_0, i_10_151_3470_0,
    i_10_151_3522_0, i_10_151_3523_0, i_10_151_3645_0, i_10_151_3682_0,
    i_10_151_3782_0, i_10_151_3847_0, i_10_151_3855_0, i_10_151_3856_0,
    i_10_151_3857_0, i_10_151_3906_0, i_10_151_3907_0, i_10_151_3979_0,
    i_10_151_4117_0, i_10_151_4118_0, i_10_151_4123_0, i_10_151_4287_0;
  output o_10_151_0_0;
  assign o_10_151_0_0 = ~((~i_10_151_82_0 & ((~i_10_151_216_0 & ~i_10_151_283_0 & ~i_10_151_902_0 & i_10_151_2656_0 & ~i_10_151_3856_0) | (~i_10_151_1912_0 & ~i_10_151_3855_0 & ~i_10_151_3907_0))) | (~i_10_151_216_0 & ((~i_10_151_1444_0 & ~i_10_151_1767_0 & ~i_10_151_2655_0 & ~i_10_151_2674_0 & ~i_10_151_2720_0 & ~i_10_151_2985_0) | (~i_10_151_219_0 & ~i_10_151_1263_0 & ~i_10_151_1485_0 & ~i_10_151_1768_0 & ~i_10_151_3045_0 & ~i_10_151_3907_0 & ~i_10_151_4287_0))) | (~i_10_151_424_0 & ((~i_10_151_1026_0 & ~i_10_151_1263_0 & ~i_10_151_2325_0 & ~i_10_151_2637_0 & ~i_10_151_3391_0 & i_10_151_3855_0 & ~i_10_151_3906_0 & ~i_10_151_3907_0) | (i_10_151_1767_0 & ~i_10_151_1768_0 & i_10_151_4287_0))) | (~i_10_151_1263_0 & ((i_10_151_467_0 & ~i_10_151_2718_0 & ~i_10_151_2719_0 & ~i_10_151_3847_0) | (~i_10_151_2659_0 & ~i_10_151_3045_0 & ~i_10_151_3856_0))) | (~i_10_151_1485_0 & ((~i_10_151_1912_0 & ~i_10_151_2637_0 & ~i_10_151_2722_0 & ~i_10_151_2884_0) | (~i_10_151_435_0 & ~i_10_151_1444_0 & ~i_10_151_2723_0 & ~i_10_151_3196_0 & ~i_10_151_3522_0 & ~i_10_151_4123_0 & ~i_10_151_4287_0))) | (~i_10_151_1444_0 & ((~i_10_151_282_0 & i_10_151_283_0 & ~i_10_151_1826_0 & ~i_10_151_2655_0) | (~i_10_151_283_0 & ~i_10_151_2885_0 & ~i_10_151_3405_0 & ~i_10_151_3855_0 & i_10_151_4118_0))) | (~i_10_151_1911_0 & ((~i_10_151_436_0 & ~i_10_151_2637_0 & ~i_10_151_2826_0 & ~i_10_151_3159_0 & ~i_10_151_3522_0 & ~i_10_151_3523_0) | (i_10_151_1236_0 & ~i_10_151_1652_0 & ~i_10_151_3391_0 & i_10_151_3857_0))) | (~i_10_151_3855_0 & ((~i_10_151_1432_0 & ~i_10_151_1688_0 & ~i_10_151_1767_0 & ~i_10_151_2449_0 & ~i_10_151_2921_0 & ~i_10_151_3159_0) | (~i_10_151_460_0 & ~i_10_151_1825_0 & i_10_151_2722_0 & ~i_10_151_3857_0 & ~i_10_151_3907_0))) | (~i_10_151_2658_0 & ~i_10_151_2721_0) | (i_10_151_1825_0 & i_10_151_3033_0 & ~i_10_151_3388_0) | (~i_10_151_2719_0 & i_10_151_3045_0 & ~i_10_151_3856_0));
endmodule



// Benchmark "kernel_10_152" written by ABC on Sun Jul 19 10:23:35 2020

module kernel_10_152 ( 
    i_10_152_153_0, i_10_152_175_0, i_10_152_220_0, i_10_152_257_0,
    i_10_152_315_0, i_10_152_316_0, i_10_152_392_0, i_10_152_432_0,
    i_10_152_437_0, i_10_152_464_0, i_10_152_561_0, i_10_152_588_0,
    i_10_152_799_0, i_10_152_1034_0, i_10_152_1039_0, i_10_152_1087_0,
    i_10_152_1234_0, i_10_152_1236_0, i_10_152_1239_0, i_10_152_1310_0,
    i_10_152_1355_0, i_10_152_1385_0, i_10_152_1432_0, i_10_152_1436_0,
    i_10_152_1448_0, i_10_152_1542_0, i_10_152_1543_0, i_10_152_1549_0,
    i_10_152_1551_0, i_10_152_1576_0, i_10_152_1655_0, i_10_152_1686_0,
    i_10_152_1687_0, i_10_152_1729_0, i_10_152_1732_0, i_10_152_1824_0,
    i_10_152_1826_0, i_10_152_1880_0, i_10_152_1951_0, i_10_152_1982_0,
    i_10_152_1984_0, i_10_152_1987_0, i_10_152_2107_0, i_10_152_2108_0,
    i_10_152_2158_0, i_10_152_2204_0, i_10_152_2331_0, i_10_152_2338_0,
    i_10_152_2352_0, i_10_152_2364_0, i_10_152_2383_0, i_10_152_2468_0,
    i_10_152_2538_0, i_10_152_2541_0, i_10_152_2632_0, i_10_152_2640_0,
    i_10_152_2731_0, i_10_152_2734_0, i_10_152_2820_0, i_10_152_2826_0,
    i_10_152_2827_0, i_10_152_2831_0, i_10_152_2881_0, i_10_152_2884_0,
    i_10_152_3043_0, i_10_152_3070_0, i_10_152_3071_0, i_10_152_3074_0,
    i_10_152_3075_0, i_10_152_3271_0, i_10_152_3277_0, i_10_152_3278_0,
    i_10_152_3282_0, i_10_152_3318_0, i_10_152_3354_0, i_10_152_3384_0,
    i_10_152_3433_0, i_10_152_3471_0, i_10_152_3540_0, i_10_152_3541_0,
    i_10_152_3542_0, i_10_152_3645_0, i_10_152_3652_0, i_10_152_3811_0,
    i_10_152_3851_0, i_10_152_3944_0, i_10_152_4086_0, i_10_152_4127_0,
    i_10_152_4172_0, i_10_152_4173_0, i_10_152_4174_0, i_10_152_4175_0,
    i_10_152_4219_0, i_10_152_4279_0, i_10_152_4280_0, i_10_152_4281_0,
    i_10_152_4282_0, i_10_152_4459_0, i_10_152_4533_0, i_10_152_4568_0,
    o_10_152_0_0  );
  input  i_10_152_153_0, i_10_152_175_0, i_10_152_220_0, i_10_152_257_0,
    i_10_152_315_0, i_10_152_316_0, i_10_152_392_0, i_10_152_432_0,
    i_10_152_437_0, i_10_152_464_0, i_10_152_561_0, i_10_152_588_0,
    i_10_152_799_0, i_10_152_1034_0, i_10_152_1039_0, i_10_152_1087_0,
    i_10_152_1234_0, i_10_152_1236_0, i_10_152_1239_0, i_10_152_1310_0,
    i_10_152_1355_0, i_10_152_1385_0, i_10_152_1432_0, i_10_152_1436_0,
    i_10_152_1448_0, i_10_152_1542_0, i_10_152_1543_0, i_10_152_1549_0,
    i_10_152_1551_0, i_10_152_1576_0, i_10_152_1655_0, i_10_152_1686_0,
    i_10_152_1687_0, i_10_152_1729_0, i_10_152_1732_0, i_10_152_1824_0,
    i_10_152_1826_0, i_10_152_1880_0, i_10_152_1951_0, i_10_152_1982_0,
    i_10_152_1984_0, i_10_152_1987_0, i_10_152_2107_0, i_10_152_2108_0,
    i_10_152_2158_0, i_10_152_2204_0, i_10_152_2331_0, i_10_152_2338_0,
    i_10_152_2352_0, i_10_152_2364_0, i_10_152_2383_0, i_10_152_2468_0,
    i_10_152_2538_0, i_10_152_2541_0, i_10_152_2632_0, i_10_152_2640_0,
    i_10_152_2731_0, i_10_152_2734_0, i_10_152_2820_0, i_10_152_2826_0,
    i_10_152_2827_0, i_10_152_2831_0, i_10_152_2881_0, i_10_152_2884_0,
    i_10_152_3043_0, i_10_152_3070_0, i_10_152_3071_0, i_10_152_3074_0,
    i_10_152_3075_0, i_10_152_3271_0, i_10_152_3277_0, i_10_152_3278_0,
    i_10_152_3282_0, i_10_152_3318_0, i_10_152_3354_0, i_10_152_3384_0,
    i_10_152_3433_0, i_10_152_3471_0, i_10_152_3540_0, i_10_152_3541_0,
    i_10_152_3542_0, i_10_152_3645_0, i_10_152_3652_0, i_10_152_3811_0,
    i_10_152_3851_0, i_10_152_3944_0, i_10_152_4086_0, i_10_152_4127_0,
    i_10_152_4172_0, i_10_152_4173_0, i_10_152_4174_0, i_10_152_4175_0,
    i_10_152_4219_0, i_10_152_4279_0, i_10_152_4280_0, i_10_152_4281_0,
    i_10_152_4282_0, i_10_152_4459_0, i_10_152_4533_0, i_10_152_4568_0;
  output o_10_152_0_0;
  assign o_10_152_0_0 = 0;
endmodule



// Benchmark "kernel_10_153" written by ABC on Sun Jul 19 10:23:36 2020

module kernel_10_153 ( 
    i_10_153_171_0, i_10_153_244_0, i_10_153_245_0, i_10_153_253_0,
    i_10_153_254_0, i_10_153_279_0, i_10_153_283_0, i_10_153_284_0,
    i_10_153_329_0, i_10_153_392_0, i_10_153_434_0, i_10_153_441_0,
    i_10_153_442_0, i_10_153_443_0, i_10_153_514_0, i_10_153_515_0,
    i_10_153_542_0, i_10_153_712_0, i_10_153_713_0, i_10_153_748_0,
    i_10_153_793_0, i_10_153_794_0, i_10_153_797_0, i_10_153_956_0,
    i_10_153_1000_0, i_10_153_1027_0, i_10_153_1028_0, i_10_153_1162_0,
    i_10_153_1234_0, i_10_153_1235_0, i_10_153_1237_0, i_10_153_1243_0,
    i_10_153_1244_0, i_10_153_1306_0, i_10_153_1310_0, i_10_153_1347_0,
    i_10_153_1540_0, i_10_153_1541_0, i_10_153_1549_0, i_10_153_1580_0,
    i_10_153_1650_0, i_10_153_1655_0, i_10_153_1684_0, i_10_153_1687_0,
    i_10_153_1688_0, i_10_153_1821_0, i_10_153_1823_0, i_10_153_2305_0,
    i_10_153_2306_0, i_10_153_2333_0, i_10_153_2349_0, i_10_153_2359_0,
    i_10_153_2361_0, i_10_153_2377_0, i_10_153_2452_0, i_10_153_2467_0,
    i_10_153_2512_0, i_10_153_2531_0, i_10_153_2603_0, i_10_153_2629_0,
    i_10_153_2632_0, i_10_153_2657_0, i_10_153_2660_0, i_10_153_2701_0,
    i_10_153_2711_0, i_10_153_2730_0, i_10_153_2732_0, i_10_153_2783_0,
    i_10_153_2827_0, i_10_153_3072_0, i_10_153_3073_0, i_10_153_3074_0,
    i_10_153_3196_0, i_10_153_3199_0, i_10_153_3200_0, i_10_153_3332_0,
    i_10_153_3384_0, i_10_153_3385_0, i_10_153_3388_0, i_10_153_3391_0,
    i_10_153_3409_0, i_10_153_3586_0, i_10_153_3587_0, i_10_153_3613_0,
    i_10_153_3614_0, i_10_153_3650_0, i_10_153_3781_0, i_10_153_3782_0,
    i_10_153_3784_0, i_10_153_3785_0, i_10_153_3788_0, i_10_153_3835_0,
    i_10_153_3838_0, i_10_153_3841_0, i_10_153_3842_0, i_10_153_4115_0,
    i_10_153_4123_0, i_10_153_4125_0, i_10_153_4126_0, i_10_153_4565_0,
    o_10_153_0_0  );
  input  i_10_153_171_0, i_10_153_244_0, i_10_153_245_0, i_10_153_253_0,
    i_10_153_254_0, i_10_153_279_0, i_10_153_283_0, i_10_153_284_0,
    i_10_153_329_0, i_10_153_392_0, i_10_153_434_0, i_10_153_441_0,
    i_10_153_442_0, i_10_153_443_0, i_10_153_514_0, i_10_153_515_0,
    i_10_153_542_0, i_10_153_712_0, i_10_153_713_0, i_10_153_748_0,
    i_10_153_793_0, i_10_153_794_0, i_10_153_797_0, i_10_153_956_0,
    i_10_153_1000_0, i_10_153_1027_0, i_10_153_1028_0, i_10_153_1162_0,
    i_10_153_1234_0, i_10_153_1235_0, i_10_153_1237_0, i_10_153_1243_0,
    i_10_153_1244_0, i_10_153_1306_0, i_10_153_1310_0, i_10_153_1347_0,
    i_10_153_1540_0, i_10_153_1541_0, i_10_153_1549_0, i_10_153_1580_0,
    i_10_153_1650_0, i_10_153_1655_0, i_10_153_1684_0, i_10_153_1687_0,
    i_10_153_1688_0, i_10_153_1821_0, i_10_153_1823_0, i_10_153_2305_0,
    i_10_153_2306_0, i_10_153_2333_0, i_10_153_2349_0, i_10_153_2359_0,
    i_10_153_2361_0, i_10_153_2377_0, i_10_153_2452_0, i_10_153_2467_0,
    i_10_153_2512_0, i_10_153_2531_0, i_10_153_2603_0, i_10_153_2629_0,
    i_10_153_2632_0, i_10_153_2657_0, i_10_153_2660_0, i_10_153_2701_0,
    i_10_153_2711_0, i_10_153_2730_0, i_10_153_2732_0, i_10_153_2783_0,
    i_10_153_2827_0, i_10_153_3072_0, i_10_153_3073_0, i_10_153_3074_0,
    i_10_153_3196_0, i_10_153_3199_0, i_10_153_3200_0, i_10_153_3332_0,
    i_10_153_3384_0, i_10_153_3385_0, i_10_153_3388_0, i_10_153_3391_0,
    i_10_153_3409_0, i_10_153_3586_0, i_10_153_3587_0, i_10_153_3613_0,
    i_10_153_3614_0, i_10_153_3650_0, i_10_153_3781_0, i_10_153_3782_0,
    i_10_153_3784_0, i_10_153_3785_0, i_10_153_3788_0, i_10_153_3835_0,
    i_10_153_3838_0, i_10_153_3841_0, i_10_153_3842_0, i_10_153_4115_0,
    i_10_153_4123_0, i_10_153_4125_0, i_10_153_4126_0, i_10_153_4565_0;
  output o_10_153_0_0;
  assign o_10_153_0_0 = 0;
endmodule



// Benchmark "kernel_10_154" written by ABC on Sun Jul 19 10:23:38 2020

module kernel_10_154 ( 
    i_10_154_27_0, i_10_154_187_0, i_10_154_188_0, i_10_154_223_0,
    i_10_154_284_0, i_10_154_315_0, i_10_154_316_0, i_10_154_317_0,
    i_10_154_323_0, i_10_154_329_0, i_10_154_409_0, i_10_154_445_0,
    i_10_154_446_0, i_10_154_458_0, i_10_154_515_0, i_10_154_793_0,
    i_10_154_797_0, i_10_154_798_0, i_10_154_800_0, i_10_154_954_0,
    i_10_154_966_0, i_10_154_1001_0, i_10_154_1028_0, i_10_154_1234_0,
    i_10_154_1309_0, i_10_154_1310_0, i_10_154_1345_0, i_10_154_1432_0,
    i_10_154_1444_0, i_10_154_1547_0, i_10_154_1555_0, i_10_154_1582_0,
    i_10_154_1583_0, i_10_154_1648_0, i_10_154_1822_0, i_10_154_1823_0,
    i_10_154_1952_0, i_10_154_2179_0, i_10_154_2353_0, i_10_154_2354_0,
    i_10_154_2356_0, i_10_154_2357_0, i_10_154_2363_0, i_10_154_2381_0,
    i_10_154_2450_0, i_10_154_2453_0, i_10_154_2632_0, i_10_154_2659_0,
    i_10_154_2702_0, i_10_154_2707_0, i_10_154_2718_0, i_10_154_2719_0,
    i_10_154_2720_0, i_10_154_2722_0, i_10_154_2828_0, i_10_154_2833_0,
    i_10_154_2884_0, i_10_154_2920_0, i_10_154_2923_0, i_10_154_2924_0,
    i_10_154_3037_0, i_10_154_3070_0, i_10_154_3071_0, i_10_154_3152_0,
    i_10_154_3277_0, i_10_154_3278_0, i_10_154_3281_0, i_10_154_3324_0,
    i_10_154_3390_0, i_10_154_3391_0, i_10_154_3466_0, i_10_154_3467_0,
    i_10_154_3519_0, i_10_154_3586_0, i_10_154_3612_0, i_10_154_3613_0,
    i_10_154_3614_0, i_10_154_3617_0, i_10_154_3653_0, i_10_154_3780_0,
    i_10_154_3781_0, i_10_154_3784_0, i_10_154_3786_0, i_10_154_3788_0,
    i_10_154_3835_0, i_10_154_3837_0, i_10_154_3838_0, i_10_154_3848_0,
    i_10_154_3856_0, i_10_154_3857_0, i_10_154_3890_0, i_10_154_3907_0,
    i_10_154_4114_0, i_10_154_4115_0, i_10_154_4282_0, i_10_154_4283_0,
    i_10_154_4287_0, i_10_154_4288_0, i_10_154_4289_0, i_10_154_4564_0,
    o_10_154_0_0  );
  input  i_10_154_27_0, i_10_154_187_0, i_10_154_188_0, i_10_154_223_0,
    i_10_154_284_0, i_10_154_315_0, i_10_154_316_0, i_10_154_317_0,
    i_10_154_323_0, i_10_154_329_0, i_10_154_409_0, i_10_154_445_0,
    i_10_154_446_0, i_10_154_458_0, i_10_154_515_0, i_10_154_793_0,
    i_10_154_797_0, i_10_154_798_0, i_10_154_800_0, i_10_154_954_0,
    i_10_154_966_0, i_10_154_1001_0, i_10_154_1028_0, i_10_154_1234_0,
    i_10_154_1309_0, i_10_154_1310_0, i_10_154_1345_0, i_10_154_1432_0,
    i_10_154_1444_0, i_10_154_1547_0, i_10_154_1555_0, i_10_154_1582_0,
    i_10_154_1583_0, i_10_154_1648_0, i_10_154_1822_0, i_10_154_1823_0,
    i_10_154_1952_0, i_10_154_2179_0, i_10_154_2353_0, i_10_154_2354_0,
    i_10_154_2356_0, i_10_154_2357_0, i_10_154_2363_0, i_10_154_2381_0,
    i_10_154_2450_0, i_10_154_2453_0, i_10_154_2632_0, i_10_154_2659_0,
    i_10_154_2702_0, i_10_154_2707_0, i_10_154_2718_0, i_10_154_2719_0,
    i_10_154_2720_0, i_10_154_2722_0, i_10_154_2828_0, i_10_154_2833_0,
    i_10_154_2884_0, i_10_154_2920_0, i_10_154_2923_0, i_10_154_2924_0,
    i_10_154_3037_0, i_10_154_3070_0, i_10_154_3071_0, i_10_154_3152_0,
    i_10_154_3277_0, i_10_154_3278_0, i_10_154_3281_0, i_10_154_3324_0,
    i_10_154_3390_0, i_10_154_3391_0, i_10_154_3466_0, i_10_154_3467_0,
    i_10_154_3519_0, i_10_154_3586_0, i_10_154_3612_0, i_10_154_3613_0,
    i_10_154_3614_0, i_10_154_3617_0, i_10_154_3653_0, i_10_154_3780_0,
    i_10_154_3781_0, i_10_154_3784_0, i_10_154_3786_0, i_10_154_3788_0,
    i_10_154_3835_0, i_10_154_3837_0, i_10_154_3838_0, i_10_154_3848_0,
    i_10_154_3856_0, i_10_154_3857_0, i_10_154_3890_0, i_10_154_3907_0,
    i_10_154_4114_0, i_10_154_4115_0, i_10_154_4282_0, i_10_154_4283_0,
    i_10_154_4287_0, i_10_154_4288_0, i_10_154_4289_0, i_10_154_4564_0;
  output o_10_154_0_0;
  assign o_10_154_0_0 = ~((~i_10_154_2179_0 & ((~i_10_154_458_0 & ((~i_10_154_3784_0 & ((~i_10_154_284_0 & ~i_10_154_3835_0 & i_10_154_3856_0 & ((~i_10_154_954_0 & ~i_10_154_1582_0 & ~i_10_154_2356_0 & ~i_10_154_2722_0) | (~i_10_154_1234_0 & ~i_10_154_1583_0 & ~i_10_154_2884_0))) | (~i_10_154_2707_0 & i_10_154_2828_0 & ~i_10_154_3780_0))) | (~i_10_154_446_0 & ~i_10_154_954_0 & ~i_10_154_1001_0 & ~i_10_154_1583_0 & ~i_10_154_1648_0 & ~i_10_154_2833_0 & ~i_10_154_2920_0 & ~i_10_154_2924_0 & ~i_10_154_3466_0 & ~i_10_154_3614_0 & ~i_10_154_3788_0 & ~i_10_154_4564_0))) | (~i_10_154_1028_0 & ~i_10_154_2453_0 & ((~i_10_154_1001_0 & ~i_10_154_3390_0 & ~i_10_154_3612_0 & ~i_10_154_3613_0 & ~i_10_154_3653_0 & ~i_10_154_3857_0) | (~i_10_154_1310_0 & ~i_10_154_1547_0 & ~i_10_154_1648_0 & i_10_154_3788_0 & i_10_154_4114_0))) | (~i_10_154_3281_0 & ~i_10_154_3786_0 & ((~i_10_154_800_0 & ~i_10_154_1309_0 & ~i_10_154_1310_0 & ~i_10_154_2722_0 & ~i_10_154_2828_0 & ~i_10_154_3070_0 & ~i_10_154_3391_0 & ~i_10_154_3835_0) | (~i_10_154_1582_0 & ~i_10_154_1823_0 & ~i_10_154_2363_0 & ~i_10_154_3466_0 & ~i_10_154_3614_0 & ~i_10_154_3617_0 & ~i_10_154_3780_0 & ~i_10_154_4282_0))) | (~i_10_154_1309_0 & ~i_10_154_3467_0 & ((~i_10_154_793_0 & i_10_154_2632_0 & i_10_154_2923_0 & ~i_10_154_3037_0 & ~i_10_154_3071_0) | (~i_10_154_3612_0 & ~i_10_154_3614_0 & ~i_10_154_3857_0 & ~i_10_154_4114_0))) | (~i_10_154_2354_0 & i_10_154_4288_0))) | (~i_10_154_458_0 & ((i_10_154_1345_0 & ~i_10_154_3612_0) | (~i_10_154_800_0 & ~i_10_154_2453_0 & ~i_10_154_2884_0 & ~i_10_154_3391_0 & ~i_10_154_3467_0 & ~i_10_154_3586_0 & ~i_10_154_3613_0 & ~i_10_154_3781_0 & ~i_10_154_3788_0))) | (i_10_154_793_0 & ((i_10_154_3281_0 & i_10_154_3519_0) | (~i_10_154_3281_0 & ~i_10_154_3614_0 & ~i_10_154_3788_0 & ~i_10_154_3837_0))) | (~i_10_154_1310_0 & ((~i_10_154_954_0 & ((~i_10_154_793_0 & ~i_10_154_2450_0 & ~i_10_154_2920_0 & ~i_10_154_2924_0 & ~i_10_154_3391_0 & ~i_10_154_3612_0) | (~i_10_154_187_0 & ~i_10_154_188_0 & ~i_10_154_2707_0 & i_10_154_3391_0 & ~i_10_154_3653_0))) | (~i_10_154_1309_0 & ~i_10_154_1823_0 & ~i_10_154_2356_0 & ~i_10_154_3070_0 & ~i_10_154_3617_0 & i_10_154_3781_0) | (~i_10_154_27_0 & ~i_10_154_1648_0 & ~i_10_154_3781_0 & i_10_154_3835_0 & ~i_10_154_3856_0))) | (~i_10_154_27_0 & ((i_10_154_1952_0 & ~i_10_154_2884_0 & ~i_10_154_3467_0 & ~i_10_154_3613_0 & ~i_10_154_3614_0 & ~i_10_154_3784_0) | (~i_10_154_187_0 & ~i_10_154_1028_0 & ~i_10_154_1555_0 & ~i_10_154_1583_0 & ~i_10_154_2363_0 & i_10_154_2722_0 & ~i_10_154_3037_0 & ~i_10_154_3466_0 & i_10_154_3856_0))) | (~i_10_154_187_0 & ((~i_10_154_317_0 & i_10_154_800_0 & ~i_10_154_1582_0 & ~i_10_154_1583_0 & ~i_10_154_1648_0 & ~i_10_154_2357_0 & ~i_10_154_2833_0 & ~i_10_154_3037_0 & ~i_10_154_3467_0) | (i_10_154_798_0 & ~i_10_154_2707_0 & ~i_10_154_3653_0 & ~i_10_154_3786_0))) | (~i_10_154_1547_0 & ((~i_10_154_1823_0 & ~i_10_154_2356_0 & ~i_10_154_2357_0 & ~i_10_154_2833_0 & ~i_10_154_3617_0 & i_10_154_3653_0 & ~i_10_154_3835_0 & ~i_10_154_3837_0 & ~i_10_154_4115_0) | (~i_10_154_1432_0 & i_10_154_2353_0 & ~i_10_154_3781_0 & ~i_10_154_3838_0 & ~i_10_154_3848_0 & ~i_10_154_4283_0))) | (~i_10_154_4282_0 & ((~i_10_154_1432_0 & ~i_10_154_1583_0 & ((~i_10_154_1582_0 & i_10_154_1822_0 & i_10_154_3037_0 & ~i_10_154_3586_0 & ~i_10_154_3614_0) | (~i_10_154_323_0 & ~i_10_154_1952_0 & ~i_10_154_2353_0 & ~i_10_154_2453_0 & ~i_10_154_3037_0 & ~i_10_154_3781_0 & ~i_10_154_3856_0))) | (~i_10_154_1234_0 & ~i_10_154_3613_0 & ~i_10_154_3614_0 & ~i_10_154_3781_0 & i_10_154_3835_0) | (~i_10_154_223_0 & i_10_154_2632_0 & ~i_10_154_3037_0 & ~i_10_154_3070_0 & i_10_154_3612_0 & ~i_10_154_3835_0))) | (~i_10_154_1822_0 & ((~i_10_154_3653_0 & ~i_10_154_3786_0 & i_10_154_27_0 & ~i_10_154_3613_0) | (~i_10_154_798_0 & ~i_10_154_1345_0 & ~i_10_154_1583_0 & ~i_10_154_1823_0 & ~i_10_154_2356_0 & ~i_10_154_2659_0 & ~i_10_154_2707_0 & ~i_10_154_2923_0 & ~i_10_154_3586_0 & ~i_10_154_4115_0))) | (~i_10_154_3612_0 & ((i_10_154_458_0 & ~i_10_154_1648_0 & ~i_10_154_2923_0 & ~i_10_154_3281_0 & ~i_10_154_3613_0 & ~i_10_154_3780_0) | (i_10_154_1234_0 & ~i_10_154_3467_0 & i_10_154_3848_0 & ~i_10_154_4114_0))) | (~i_10_154_3784_0 & ~i_10_154_3857_0 & ((i_10_154_2354_0 & ~i_10_154_3391_0 & ~i_10_154_3613_0 & ~i_10_154_3786_0 & i_10_154_3835_0) | (i_10_154_446_0 & i_10_154_797_0 & ~i_10_154_4283_0))) | (~i_10_154_1028_0 & ~i_10_154_1823_0 & i_10_154_2720_0) | (~i_10_154_2450_0 & ~i_10_154_3653_0 & ~i_10_154_3788_0 & i_10_154_4289_0));
endmodule



// Benchmark "kernel_10_155" written by ABC on Sun Jul 19 10:23:39 2020

module kernel_10_155 ( 
    i_10_155_177_0, i_10_155_246_0, i_10_155_249_0, i_10_155_252_0,
    i_10_155_264_0, i_10_155_318_0, i_10_155_320_0, i_10_155_321_0,
    i_10_155_322_0, i_10_155_327_0, i_10_155_413_0, i_10_155_462_0,
    i_10_155_933_0, i_10_155_1002_0, i_10_155_1007_0, i_10_155_1030_0,
    i_10_155_1032_0, i_10_155_1107_0, i_10_155_1110_0, i_10_155_1299_0,
    i_10_155_1302_0, i_10_155_1307_0, i_10_155_1431_0, i_10_155_1434_0,
    i_10_155_1437_0, i_10_155_1545_0, i_10_155_1581_0, i_10_155_1626_0,
    i_10_155_1654_0, i_10_155_1686_0, i_10_155_1731_0, i_10_155_1734_0,
    i_10_155_1735_0, i_10_155_1764_0, i_10_155_1806_0, i_10_155_1818_0,
    i_10_155_1821_0, i_10_155_1823_0, i_10_155_1983_0, i_10_155_1986_0,
    i_10_155_2031_0, i_10_155_2202_0, i_10_155_2349_0, i_10_155_2350_0,
    i_10_155_2351_0, i_10_155_2353_0, i_10_155_2358_0, i_10_155_2450_0,
    i_10_155_2472_0, i_10_155_2565_0, i_10_155_2568_0, i_10_155_2571_0,
    i_10_155_2604_0, i_10_155_2617_0, i_10_155_2663_0, i_10_155_2676_0,
    i_10_155_2680_0, i_10_155_2708_0, i_10_155_2712_0, i_10_155_2722_0,
    i_10_155_2734_0, i_10_155_2760_0, i_10_155_2826_0, i_10_155_2828_0,
    i_10_155_2847_0, i_10_155_2850_0, i_10_155_2920_0, i_10_155_2924_0,
    i_10_155_3045_0, i_10_155_3072_0, i_10_155_3073_0, i_10_155_3075_0,
    i_10_155_3202_0, i_10_155_3280_0, i_10_155_3390_0, i_10_155_3391_0,
    i_10_155_3434_0, i_10_155_3525_0, i_10_155_3540_0, i_10_155_3543_0,
    i_10_155_3544_0, i_10_155_3585_0, i_10_155_3617_0, i_10_155_3622_0,
    i_10_155_3645_0, i_10_155_3650_0, i_10_155_3787_0, i_10_155_3837_0,
    i_10_155_3854_0, i_10_155_3990_0, i_10_155_4029_0, i_10_155_4113_0,
    i_10_155_4115_0, i_10_155_4116_0, i_10_155_4117_0, i_10_155_4128_0,
    i_10_155_4168_0, i_10_155_4273_0, i_10_155_4584_0, i_10_155_4588_0,
    o_10_155_0_0  );
  input  i_10_155_177_0, i_10_155_246_0, i_10_155_249_0, i_10_155_252_0,
    i_10_155_264_0, i_10_155_318_0, i_10_155_320_0, i_10_155_321_0,
    i_10_155_322_0, i_10_155_327_0, i_10_155_413_0, i_10_155_462_0,
    i_10_155_933_0, i_10_155_1002_0, i_10_155_1007_0, i_10_155_1030_0,
    i_10_155_1032_0, i_10_155_1107_0, i_10_155_1110_0, i_10_155_1299_0,
    i_10_155_1302_0, i_10_155_1307_0, i_10_155_1431_0, i_10_155_1434_0,
    i_10_155_1437_0, i_10_155_1545_0, i_10_155_1581_0, i_10_155_1626_0,
    i_10_155_1654_0, i_10_155_1686_0, i_10_155_1731_0, i_10_155_1734_0,
    i_10_155_1735_0, i_10_155_1764_0, i_10_155_1806_0, i_10_155_1818_0,
    i_10_155_1821_0, i_10_155_1823_0, i_10_155_1983_0, i_10_155_1986_0,
    i_10_155_2031_0, i_10_155_2202_0, i_10_155_2349_0, i_10_155_2350_0,
    i_10_155_2351_0, i_10_155_2353_0, i_10_155_2358_0, i_10_155_2450_0,
    i_10_155_2472_0, i_10_155_2565_0, i_10_155_2568_0, i_10_155_2571_0,
    i_10_155_2604_0, i_10_155_2617_0, i_10_155_2663_0, i_10_155_2676_0,
    i_10_155_2680_0, i_10_155_2708_0, i_10_155_2712_0, i_10_155_2722_0,
    i_10_155_2734_0, i_10_155_2760_0, i_10_155_2826_0, i_10_155_2828_0,
    i_10_155_2847_0, i_10_155_2850_0, i_10_155_2920_0, i_10_155_2924_0,
    i_10_155_3045_0, i_10_155_3072_0, i_10_155_3073_0, i_10_155_3075_0,
    i_10_155_3202_0, i_10_155_3280_0, i_10_155_3390_0, i_10_155_3391_0,
    i_10_155_3434_0, i_10_155_3525_0, i_10_155_3540_0, i_10_155_3543_0,
    i_10_155_3544_0, i_10_155_3585_0, i_10_155_3617_0, i_10_155_3622_0,
    i_10_155_3645_0, i_10_155_3650_0, i_10_155_3787_0, i_10_155_3837_0,
    i_10_155_3854_0, i_10_155_3990_0, i_10_155_4029_0, i_10_155_4113_0,
    i_10_155_4115_0, i_10_155_4116_0, i_10_155_4117_0, i_10_155_4128_0,
    i_10_155_4168_0, i_10_155_4273_0, i_10_155_4584_0, i_10_155_4588_0;
  output o_10_155_0_0;
  assign o_10_155_0_0 = ~((~i_10_155_1626_0 & ((~i_10_155_264_0 & ~i_10_155_2571_0) | (~i_10_155_2031_0 & ~i_10_155_2708_0 & ~i_10_155_3075_0))) | (~i_10_155_2031_0 & ((~i_10_155_2350_0 & ~i_10_155_2571_0 & ~i_10_155_2680_0 & ~i_10_155_3990_0) | (~i_10_155_1735_0 & ~i_10_155_2734_0 & ~i_10_155_3787_0 & ~i_10_155_4273_0))) | (~i_10_155_4029_0 & i_10_155_4273_0 & ((~i_10_155_3073_0 & i_10_155_3544_0) | (~i_10_155_1734_0 & ~i_10_155_2450_0 & i_10_155_3391_0 & ~i_10_155_4168_0))) | ~i_10_155_3280_0 | (i_10_155_4117_0 & ~i_10_155_4128_0));
endmodule



// Benchmark "kernel_10_156" written by ABC on Sun Jul 19 10:23:40 2020

module kernel_10_156 ( 
    i_10_156_182_0, i_10_156_248_0, i_10_156_249_0, i_10_156_271_0,
    i_10_156_280_0, i_10_156_286_0, i_10_156_317_0, i_10_156_327_0,
    i_10_156_328_0, i_10_156_408_0, i_10_156_428_0, i_10_156_434_0,
    i_10_156_443_0, i_10_156_448_0, i_10_156_796_0, i_10_156_825_0,
    i_10_156_1029_0, i_10_156_1031_0, i_10_156_1033_0, i_10_156_1034_0,
    i_10_156_1118_0, i_10_156_1245_0, i_10_156_1441_0, i_10_156_1443_0,
    i_10_156_1492_0, i_10_156_1554_0, i_10_156_1582_0, i_10_156_1650_0,
    i_10_156_1675_0, i_10_156_1680_0, i_10_156_1682_0, i_10_156_1686_0,
    i_10_156_1818_0, i_10_156_1820_0, i_10_156_1822_0, i_10_156_1826_0,
    i_10_156_1909_0, i_10_156_1911_0, i_10_156_1947_0, i_10_156_2311_0,
    i_10_156_2354_0, i_10_156_2358_0, i_10_156_2407_0, i_10_156_2449_0,
    i_10_156_2450_0, i_10_156_2470_0, i_10_156_2471_0, i_10_156_2473_0,
    i_10_156_2633_0, i_10_156_2657_0, i_10_156_2658_0, i_10_156_2662_0,
    i_10_156_2704_0, i_10_156_2709_0, i_10_156_2710_0, i_10_156_2711_0,
    i_10_156_2714_0, i_10_156_2717_0, i_10_156_2722_0, i_10_156_2723_0,
    i_10_156_2731_0, i_10_156_2732_0, i_10_156_2826_0, i_10_156_2828_0,
    i_10_156_2872_0, i_10_156_2917_0, i_10_156_2918_0, i_10_156_2919_0,
    i_10_156_2921_0, i_10_156_3034_0, i_10_156_3035_0, i_10_156_3036_0,
    i_10_156_3163_0, i_10_156_3196_0, i_10_156_3199_0, i_10_156_3283_0,
    i_10_156_3326_0, i_10_156_3389_0, i_10_156_3392_0, i_10_156_3436_0,
    i_10_156_3470_0, i_10_156_3471_0, i_10_156_3585_0, i_10_156_3586_0,
    i_10_156_3588_0, i_10_156_3589_0, i_10_156_3647_0, i_10_156_3783_0,
    i_10_156_3854_0, i_10_156_3894_0, i_10_156_3947_0, i_10_156_3984_0,
    i_10_156_3985_0, i_10_156_3991_0, i_10_156_4121_0, i_10_156_4126_0,
    i_10_156_4216_0, i_10_156_4279_0, i_10_156_4284_0, i_10_156_4566_0,
    o_10_156_0_0  );
  input  i_10_156_182_0, i_10_156_248_0, i_10_156_249_0, i_10_156_271_0,
    i_10_156_280_0, i_10_156_286_0, i_10_156_317_0, i_10_156_327_0,
    i_10_156_328_0, i_10_156_408_0, i_10_156_428_0, i_10_156_434_0,
    i_10_156_443_0, i_10_156_448_0, i_10_156_796_0, i_10_156_825_0,
    i_10_156_1029_0, i_10_156_1031_0, i_10_156_1033_0, i_10_156_1034_0,
    i_10_156_1118_0, i_10_156_1245_0, i_10_156_1441_0, i_10_156_1443_0,
    i_10_156_1492_0, i_10_156_1554_0, i_10_156_1582_0, i_10_156_1650_0,
    i_10_156_1675_0, i_10_156_1680_0, i_10_156_1682_0, i_10_156_1686_0,
    i_10_156_1818_0, i_10_156_1820_0, i_10_156_1822_0, i_10_156_1826_0,
    i_10_156_1909_0, i_10_156_1911_0, i_10_156_1947_0, i_10_156_2311_0,
    i_10_156_2354_0, i_10_156_2358_0, i_10_156_2407_0, i_10_156_2449_0,
    i_10_156_2450_0, i_10_156_2470_0, i_10_156_2471_0, i_10_156_2473_0,
    i_10_156_2633_0, i_10_156_2657_0, i_10_156_2658_0, i_10_156_2662_0,
    i_10_156_2704_0, i_10_156_2709_0, i_10_156_2710_0, i_10_156_2711_0,
    i_10_156_2714_0, i_10_156_2717_0, i_10_156_2722_0, i_10_156_2723_0,
    i_10_156_2731_0, i_10_156_2732_0, i_10_156_2826_0, i_10_156_2828_0,
    i_10_156_2872_0, i_10_156_2917_0, i_10_156_2918_0, i_10_156_2919_0,
    i_10_156_2921_0, i_10_156_3034_0, i_10_156_3035_0, i_10_156_3036_0,
    i_10_156_3163_0, i_10_156_3196_0, i_10_156_3199_0, i_10_156_3283_0,
    i_10_156_3326_0, i_10_156_3389_0, i_10_156_3392_0, i_10_156_3436_0,
    i_10_156_3470_0, i_10_156_3471_0, i_10_156_3585_0, i_10_156_3586_0,
    i_10_156_3588_0, i_10_156_3589_0, i_10_156_3647_0, i_10_156_3783_0,
    i_10_156_3854_0, i_10_156_3894_0, i_10_156_3947_0, i_10_156_3984_0,
    i_10_156_3985_0, i_10_156_3991_0, i_10_156_4121_0, i_10_156_4126_0,
    i_10_156_4216_0, i_10_156_4279_0, i_10_156_4284_0, i_10_156_4566_0;
  output o_10_156_0_0;
  assign o_10_156_0_0 = 0;
endmodule



// Benchmark "kernel_10_157" written by ABC on Sun Jul 19 10:23:41 2020

module kernel_10_157 ( 
    i_10_157_40_0, i_10_157_64_0, i_10_157_67_0, i_10_157_151_0,
    i_10_157_181_0, i_10_157_221_0, i_10_157_223_0, i_10_157_271_0,
    i_10_157_283_0, i_10_157_290_0, i_10_157_319_0, i_10_157_320_0,
    i_10_157_362_0, i_10_157_412_0, i_10_157_424_0, i_10_157_432_0,
    i_10_157_437_0, i_10_157_444_0, i_10_157_448_0, i_10_157_496_0,
    i_10_157_559_0, i_10_157_635_0, i_10_157_718_0, i_10_157_900_0,
    i_10_157_907_0, i_10_157_927_0, i_10_157_928_0, i_10_157_958_0,
    i_10_157_990_0, i_10_157_1009_0, i_10_157_1200_0, i_10_157_1236_0,
    i_10_157_1238_0, i_10_157_1241_0, i_10_157_1272_0, i_10_157_1275_0,
    i_10_157_1278_0, i_10_157_1310_0, i_10_157_1363_0, i_10_157_1364_0,
    i_10_157_1491_0, i_10_157_1579_0, i_10_157_1705_0, i_10_157_1783_0,
    i_10_157_1824_0, i_10_157_1849_0, i_10_157_1940_0, i_10_157_1943_0,
    i_10_157_2003_0, i_10_157_2052_0, i_10_157_2089_0, i_10_157_2264_0,
    i_10_157_2338_0, i_10_157_2350_0, i_10_157_2385_0, i_10_157_2452_0,
    i_10_157_2455_0, i_10_157_2476_0, i_10_157_2512_0, i_10_157_2596_0,
    i_10_157_2711_0, i_10_157_2714_0, i_10_157_2783_0, i_10_157_2830_0,
    i_10_157_2831_0, i_10_157_2910_0, i_10_157_2953_0, i_10_157_3011_0,
    i_10_157_3045_0, i_10_157_3050_0, i_10_157_3163_0, i_10_157_3198_0,
    i_10_157_3273_0, i_10_157_3275_0, i_10_157_3276_0, i_10_157_3281_0,
    i_10_157_3284_0, i_10_157_3286_0, i_10_157_3317_0, i_10_157_3386_0,
    i_10_157_3391_0, i_10_157_3469_0, i_10_157_3584_0, i_10_157_3585_0,
    i_10_157_3612_0, i_10_157_3648_0, i_10_157_3649_0, i_10_157_3682_0,
    i_10_157_3856_0, i_10_157_3860_0, i_10_157_3947_0, i_10_157_4050_0,
    i_10_157_4126_0, i_10_157_4157_0, i_10_157_4162_0, i_10_157_4192_0,
    i_10_157_4217_0, i_10_157_4282_0, i_10_157_4307_0, i_10_157_4519_0,
    o_10_157_0_0  );
  input  i_10_157_40_0, i_10_157_64_0, i_10_157_67_0, i_10_157_151_0,
    i_10_157_181_0, i_10_157_221_0, i_10_157_223_0, i_10_157_271_0,
    i_10_157_283_0, i_10_157_290_0, i_10_157_319_0, i_10_157_320_0,
    i_10_157_362_0, i_10_157_412_0, i_10_157_424_0, i_10_157_432_0,
    i_10_157_437_0, i_10_157_444_0, i_10_157_448_0, i_10_157_496_0,
    i_10_157_559_0, i_10_157_635_0, i_10_157_718_0, i_10_157_900_0,
    i_10_157_907_0, i_10_157_927_0, i_10_157_928_0, i_10_157_958_0,
    i_10_157_990_0, i_10_157_1009_0, i_10_157_1200_0, i_10_157_1236_0,
    i_10_157_1238_0, i_10_157_1241_0, i_10_157_1272_0, i_10_157_1275_0,
    i_10_157_1278_0, i_10_157_1310_0, i_10_157_1363_0, i_10_157_1364_0,
    i_10_157_1491_0, i_10_157_1579_0, i_10_157_1705_0, i_10_157_1783_0,
    i_10_157_1824_0, i_10_157_1849_0, i_10_157_1940_0, i_10_157_1943_0,
    i_10_157_2003_0, i_10_157_2052_0, i_10_157_2089_0, i_10_157_2264_0,
    i_10_157_2338_0, i_10_157_2350_0, i_10_157_2385_0, i_10_157_2452_0,
    i_10_157_2455_0, i_10_157_2476_0, i_10_157_2512_0, i_10_157_2596_0,
    i_10_157_2711_0, i_10_157_2714_0, i_10_157_2783_0, i_10_157_2830_0,
    i_10_157_2831_0, i_10_157_2910_0, i_10_157_2953_0, i_10_157_3011_0,
    i_10_157_3045_0, i_10_157_3050_0, i_10_157_3163_0, i_10_157_3198_0,
    i_10_157_3273_0, i_10_157_3275_0, i_10_157_3276_0, i_10_157_3281_0,
    i_10_157_3284_0, i_10_157_3286_0, i_10_157_3317_0, i_10_157_3386_0,
    i_10_157_3391_0, i_10_157_3469_0, i_10_157_3584_0, i_10_157_3585_0,
    i_10_157_3612_0, i_10_157_3648_0, i_10_157_3649_0, i_10_157_3682_0,
    i_10_157_3856_0, i_10_157_3860_0, i_10_157_3947_0, i_10_157_4050_0,
    i_10_157_4126_0, i_10_157_4157_0, i_10_157_4162_0, i_10_157_4192_0,
    i_10_157_4217_0, i_10_157_4282_0, i_10_157_4307_0, i_10_157_4519_0;
  output o_10_157_0_0;
  assign o_10_157_0_0 = 0;
endmodule



// Benchmark "kernel_10_158" written by ABC on Sun Jul 19 10:23:42 2020

module kernel_10_158 ( 
    i_10_158_172_0, i_10_158_223_0, i_10_158_245_0, i_10_158_251_0,
    i_10_158_254_0, i_10_158_282_0, i_10_158_284_0, i_10_158_390_0,
    i_10_158_406_0, i_10_158_426_0, i_10_158_441_0, i_10_158_443_0,
    i_10_158_459_0, i_10_158_460_0, i_10_158_463_0, i_10_158_747_0,
    i_10_158_748_0, i_10_158_749_0, i_10_158_793_0, i_10_158_794_0,
    i_10_158_796_0, i_10_158_797_0, i_10_158_1004_0, i_10_158_1026_0,
    i_10_158_1027_0, i_10_158_1033_0, i_10_158_1240_0, i_10_158_1306_0,
    i_10_158_1310_0, i_10_158_1365_0, i_10_158_1432_0, i_10_158_1433_0,
    i_10_158_1539_0, i_10_158_1540_0, i_10_158_1541_0, i_10_158_1543_0,
    i_10_158_1544_0, i_10_158_1576_0, i_10_158_1649_0, i_10_158_1683_0,
    i_10_158_1687_0, i_10_158_1821_0, i_10_158_1822_0, i_10_158_1954_0,
    i_10_158_2180_0, i_10_158_2351_0, i_10_158_2361_0, i_10_158_2450_0,
    i_10_158_2453_0, i_10_158_2461_0, i_10_158_2572_0, i_10_158_2628_0,
    i_10_158_2657_0, i_10_158_2674_0, i_10_158_2675_0, i_10_158_2701_0,
    i_10_158_2720_0, i_10_158_2733_0, i_10_158_2734_0, i_10_158_2817_0,
    i_10_158_2818_0, i_10_158_2821_0, i_10_158_2884_0, i_10_158_2923_0,
    i_10_158_2924_0, i_10_158_3035_0, i_10_158_3048_0, i_10_158_3049_0,
    i_10_158_3069_0, i_10_158_3070_0, i_10_158_3198_0, i_10_158_3199_0,
    i_10_158_3200_0, i_10_158_3270_0, i_10_158_3331_0, i_10_158_3405_0,
    i_10_158_3522_0, i_10_158_3525_0, i_10_158_3611_0, i_10_158_3612_0,
    i_10_158_3685_0, i_10_158_3686_0, i_10_158_3780_0, i_10_158_3782_0,
    i_10_158_3783_0, i_10_158_3784_0, i_10_158_3785_0, i_10_158_3837_0,
    i_10_158_3838_0, i_10_158_3842_0, i_10_158_3857_0, i_10_158_3858_0,
    i_10_158_3859_0, i_10_158_4117_0, i_10_158_4120_0, i_10_158_4121_0,
    i_10_158_4266_0, i_10_158_4269_0, i_10_158_4276_0, i_10_158_4568_0,
    o_10_158_0_0  );
  input  i_10_158_172_0, i_10_158_223_0, i_10_158_245_0, i_10_158_251_0,
    i_10_158_254_0, i_10_158_282_0, i_10_158_284_0, i_10_158_390_0,
    i_10_158_406_0, i_10_158_426_0, i_10_158_441_0, i_10_158_443_0,
    i_10_158_459_0, i_10_158_460_0, i_10_158_463_0, i_10_158_747_0,
    i_10_158_748_0, i_10_158_749_0, i_10_158_793_0, i_10_158_794_0,
    i_10_158_796_0, i_10_158_797_0, i_10_158_1004_0, i_10_158_1026_0,
    i_10_158_1027_0, i_10_158_1033_0, i_10_158_1240_0, i_10_158_1306_0,
    i_10_158_1310_0, i_10_158_1365_0, i_10_158_1432_0, i_10_158_1433_0,
    i_10_158_1539_0, i_10_158_1540_0, i_10_158_1541_0, i_10_158_1543_0,
    i_10_158_1544_0, i_10_158_1576_0, i_10_158_1649_0, i_10_158_1683_0,
    i_10_158_1687_0, i_10_158_1821_0, i_10_158_1822_0, i_10_158_1954_0,
    i_10_158_2180_0, i_10_158_2351_0, i_10_158_2361_0, i_10_158_2450_0,
    i_10_158_2453_0, i_10_158_2461_0, i_10_158_2572_0, i_10_158_2628_0,
    i_10_158_2657_0, i_10_158_2674_0, i_10_158_2675_0, i_10_158_2701_0,
    i_10_158_2720_0, i_10_158_2733_0, i_10_158_2734_0, i_10_158_2817_0,
    i_10_158_2818_0, i_10_158_2821_0, i_10_158_2884_0, i_10_158_2923_0,
    i_10_158_2924_0, i_10_158_3035_0, i_10_158_3048_0, i_10_158_3049_0,
    i_10_158_3069_0, i_10_158_3070_0, i_10_158_3198_0, i_10_158_3199_0,
    i_10_158_3200_0, i_10_158_3270_0, i_10_158_3331_0, i_10_158_3405_0,
    i_10_158_3522_0, i_10_158_3525_0, i_10_158_3611_0, i_10_158_3612_0,
    i_10_158_3685_0, i_10_158_3686_0, i_10_158_3780_0, i_10_158_3782_0,
    i_10_158_3783_0, i_10_158_3784_0, i_10_158_3785_0, i_10_158_3837_0,
    i_10_158_3838_0, i_10_158_3842_0, i_10_158_3857_0, i_10_158_3858_0,
    i_10_158_3859_0, i_10_158_4117_0, i_10_158_4120_0, i_10_158_4121_0,
    i_10_158_4266_0, i_10_158_4269_0, i_10_158_4276_0, i_10_158_4568_0;
  output o_10_158_0_0;
  assign o_10_158_0_0 = ~((~i_10_158_2180_0 & ((~i_10_158_390_0 & ~i_10_158_4266_0 & ((~i_10_158_463_0 & ~i_10_158_1687_0 & ~i_10_158_2817_0) | (~i_10_158_748_0 & ~i_10_158_749_0 & ~i_10_158_797_0 & i_10_158_1687_0 & ~i_10_158_2453_0 & ~i_10_158_2733_0 & ~i_10_158_2734_0 & ~i_10_158_3780_0))) | (~i_10_158_1365_0 & ~i_10_158_1683_0 & ~i_10_158_3782_0 & i_10_158_3842_0 & ~i_10_158_3859_0 & ~i_10_158_4269_0))) | (~i_10_158_460_0 & ((~i_10_158_3782_0 & ~i_10_158_3837_0 & i_10_158_3857_0) | (~i_10_158_748_0 & ~i_10_158_1027_0 & ~i_10_158_1240_0 & ~i_10_158_1310_0 & ~i_10_158_3049_0 & ~i_10_158_3405_0 & ~i_10_158_3857_0))) | (~i_10_158_748_0 & ~i_10_158_1821_0 & ((~i_10_158_1365_0 & ~i_10_158_1543_0 & ~i_10_158_1576_0 & ~i_10_158_3070_0 & ~i_10_158_3785_0) | (~i_10_158_796_0 & ~i_10_158_1026_0 & ~i_10_158_1541_0 & ~i_10_158_3842_0))) | (~i_10_158_1033_0 & ~i_10_158_3858_0 & ((~i_10_158_749_0 & ~i_10_158_1649_0 & ~i_10_158_1683_0 & i_10_158_3842_0 & ~i_10_158_3857_0) | (~i_10_158_443_0 & ~i_10_158_1541_0 & ~i_10_158_2351_0 & ~i_10_158_2733_0 & ~i_10_158_3611_0 & ~i_10_158_3780_0 & ~i_10_158_4269_0))) | (~i_10_158_1365_0 & ((~i_10_158_282_0 & ~i_10_158_1027_0 & ~i_10_158_3198_0) | (~i_10_158_1310_0 & ~i_10_158_1543_0 & ~i_10_158_1544_0 & ~i_10_158_3069_0 & ~i_10_158_3612_0 & ~i_10_158_3780_0))) | (~i_10_158_1027_0 & ((~i_10_158_1026_0 & i_10_158_1306_0 & ~i_10_158_1540_0 & i_10_158_3035_0 & ~i_10_158_3069_0 & ~i_10_158_3405_0) | (i_10_158_172_0 & i_10_158_4120_0))) | (~i_10_158_1649_0 & ((~i_10_158_1540_0 & ~i_10_158_1576_0 & ~i_10_158_3198_0 & ~i_10_158_3405_0 & ~i_10_158_3782_0 & ~i_10_158_3785_0) | (~i_10_158_254_0 & ~i_10_158_1539_0 & ~i_10_158_2924_0 & ~i_10_158_3048_0 & ~i_10_158_3049_0 & ~i_10_158_3069_0 & ~i_10_158_3686_0 & ~i_10_158_3842_0))) | (~i_10_158_3070_0 & ((~i_10_158_1539_0 & ((~i_10_158_2453_0 & ~i_10_158_3035_0 & ~i_10_158_3199_0 & ~i_10_158_3782_0 & ~i_10_158_3785_0) | (~i_10_158_3612_0 & ~i_10_158_3783_0 & ~i_10_158_3784_0 & i_10_158_3858_0))) | (~i_10_158_223_0 & ~i_10_158_1240_0 & ~i_10_158_3049_0 & ~i_10_158_3069_0 & ~i_10_158_3783_0 & ~i_10_158_3785_0))) | (~i_10_158_1540_0 & ((i_10_158_459_0 & i_10_158_460_0 & i_10_158_793_0 & ~i_10_158_3270_0) | (i_10_158_282_0 & ~i_10_158_1543_0 & ~i_10_158_2733_0 & ~i_10_158_3783_0))));
endmodule



// Benchmark "kernel_10_159" written by ABC on Sun Jul 19 10:23:44 2020

module kernel_10_159 ( 
    i_10_159_29_0, i_10_159_172_0, i_10_159_273_0, i_10_159_284_0,
    i_10_159_388_0, i_10_159_409_0, i_10_159_410_0, i_10_159_442_0,
    i_10_159_459_0, i_10_159_508_0, i_10_159_511_0, i_10_159_512_0,
    i_10_159_796_0, i_10_159_800_0, i_10_159_958_0, i_10_159_1001_0,
    i_10_159_1004_0, i_10_159_1034_0, i_10_159_1081_0, i_10_159_1267_0,
    i_10_159_1433_0, i_10_159_1439_0, i_10_159_1576_0, i_10_159_1654_0,
    i_10_159_1655_0, i_10_159_1683_0, i_10_159_1690_0, i_10_159_1691_0,
    i_10_159_1736_0, i_10_159_1821_0, i_10_159_1822_0, i_10_159_1823_0,
    i_10_159_1824_0, i_10_159_1825_0, i_10_159_1913_0, i_10_159_1916_0,
    i_10_159_1946_0, i_10_159_2006_0, i_10_159_2030_0, i_10_159_2033_0,
    i_10_159_2381_0, i_10_159_2408_0, i_10_159_2449_0, i_10_159_2455_0,
    i_10_159_2472_0, i_10_159_2474_0, i_10_159_2608_0, i_10_159_2634_0,
    i_10_159_2635_0, i_10_159_2675_0, i_10_159_2722_0, i_10_159_2723_0,
    i_10_159_2730_0, i_10_159_2734_0, i_10_159_2735_0, i_10_159_2830_0,
    i_10_159_2831_0, i_10_159_2833_0, i_10_159_2885_0, i_10_159_2887_0,
    i_10_159_2922_0, i_10_159_2923_0, i_10_159_2986_0, i_10_159_3035_0,
    i_10_159_3049_0, i_10_159_3088_0, i_10_159_3320_0, i_10_159_3323_0,
    i_10_159_3384_0, i_10_159_3385_0, i_10_159_3386_0, i_10_159_3388_0,
    i_10_159_3389_0, i_10_159_3437_0, i_10_159_3470_0, i_10_159_3473_0,
    i_10_159_3509_0, i_10_159_3539_0, i_10_159_3584_0, i_10_159_3587_0,
    i_10_159_3590_0, i_10_159_3617_0, i_10_159_3784_0, i_10_159_3837_0,
    i_10_159_3839_0, i_10_159_3841_0, i_10_159_3842_0, i_10_159_3843_0,
    i_10_159_3853_0, i_10_159_3860_0, i_10_159_3890_0, i_10_159_3980_0,
    i_10_159_4114_0, i_10_159_4115_0, i_10_159_4174_0, i_10_159_4268_0,
    i_10_159_4271_0, i_10_159_4274_0, i_10_159_4287_0, i_10_159_4568_0,
    o_10_159_0_0  );
  input  i_10_159_29_0, i_10_159_172_0, i_10_159_273_0, i_10_159_284_0,
    i_10_159_388_0, i_10_159_409_0, i_10_159_410_0, i_10_159_442_0,
    i_10_159_459_0, i_10_159_508_0, i_10_159_511_0, i_10_159_512_0,
    i_10_159_796_0, i_10_159_800_0, i_10_159_958_0, i_10_159_1001_0,
    i_10_159_1004_0, i_10_159_1034_0, i_10_159_1081_0, i_10_159_1267_0,
    i_10_159_1433_0, i_10_159_1439_0, i_10_159_1576_0, i_10_159_1654_0,
    i_10_159_1655_0, i_10_159_1683_0, i_10_159_1690_0, i_10_159_1691_0,
    i_10_159_1736_0, i_10_159_1821_0, i_10_159_1822_0, i_10_159_1823_0,
    i_10_159_1824_0, i_10_159_1825_0, i_10_159_1913_0, i_10_159_1916_0,
    i_10_159_1946_0, i_10_159_2006_0, i_10_159_2030_0, i_10_159_2033_0,
    i_10_159_2381_0, i_10_159_2408_0, i_10_159_2449_0, i_10_159_2455_0,
    i_10_159_2472_0, i_10_159_2474_0, i_10_159_2608_0, i_10_159_2634_0,
    i_10_159_2635_0, i_10_159_2675_0, i_10_159_2722_0, i_10_159_2723_0,
    i_10_159_2730_0, i_10_159_2734_0, i_10_159_2735_0, i_10_159_2830_0,
    i_10_159_2831_0, i_10_159_2833_0, i_10_159_2885_0, i_10_159_2887_0,
    i_10_159_2922_0, i_10_159_2923_0, i_10_159_2986_0, i_10_159_3035_0,
    i_10_159_3049_0, i_10_159_3088_0, i_10_159_3320_0, i_10_159_3323_0,
    i_10_159_3384_0, i_10_159_3385_0, i_10_159_3386_0, i_10_159_3388_0,
    i_10_159_3389_0, i_10_159_3437_0, i_10_159_3470_0, i_10_159_3473_0,
    i_10_159_3509_0, i_10_159_3539_0, i_10_159_3584_0, i_10_159_3587_0,
    i_10_159_3590_0, i_10_159_3617_0, i_10_159_3784_0, i_10_159_3837_0,
    i_10_159_3839_0, i_10_159_3841_0, i_10_159_3842_0, i_10_159_3843_0,
    i_10_159_3853_0, i_10_159_3860_0, i_10_159_3890_0, i_10_159_3980_0,
    i_10_159_4114_0, i_10_159_4115_0, i_10_159_4174_0, i_10_159_4268_0,
    i_10_159_4271_0, i_10_159_4274_0, i_10_159_4287_0, i_10_159_4568_0;
  output o_10_159_0_0;
  assign o_10_159_0_0 = ~((~i_10_159_3509_0 & ((~i_10_159_388_0 & ((~i_10_159_442_0 & i_10_159_1654_0 & ~i_10_159_1690_0 & ~i_10_159_1736_0 & ~i_10_159_2006_0 & ~i_10_159_2887_0 & ~i_10_159_4114_0) | (~i_10_159_796_0 & ~i_10_159_1001_0 & i_10_159_1823_0 & ~i_10_159_2408_0 & ~i_10_159_2472_0 & ~i_10_159_2885_0 & ~i_10_159_3843_0 & ~i_10_159_4268_0 & ~i_10_159_4271_0 & ~i_10_159_4274_0))) | (~i_10_159_1433_0 & ((~i_10_159_409_0 & ~i_10_159_1001_0 & i_10_159_2830_0 & ~i_10_159_3320_0 & ~i_10_159_3473_0 & ~i_10_159_3590_0) | (~i_10_159_1690_0 & ~i_10_159_2735_0 & ~i_10_159_3035_0 & ~i_10_159_3584_0 & ~i_10_159_3839_0 & ~i_10_159_3890_0 & ~i_10_159_4174_0 & ~i_10_159_4268_0))) | (~i_10_159_1001_0 & ~i_10_159_2735_0 & ~i_10_159_2885_0 & ((~i_10_159_1821_0 & ~i_10_159_1823_0 & ~i_10_159_2381_0 & ~i_10_159_2408_0) | (~i_10_159_29_0 & ~i_10_159_1004_0 & ~i_10_159_1946_0 & ~i_10_159_2006_0 & ~i_10_159_2734_0 & ~i_10_159_3320_0 & ~i_10_159_4268_0 & ~i_10_159_4271_0 & ~i_10_159_4568_0))) | (~i_10_159_3980_0 & ((~i_10_159_1690_0 & i_10_159_1824_0 & ~i_10_159_1946_0 & ~i_10_159_3035_0 & ~i_10_159_3473_0 & ~i_10_159_3587_0 & ~i_10_159_3784_0) | (~i_10_159_1439_0 & ~i_10_159_1825_0 & ~i_10_159_2006_0 & i_10_159_2635_0 & ~i_10_159_3470_0 & ~i_10_159_3841_0 & ~i_10_159_4268_0 & ~i_10_159_4274_0))))) | (~i_10_159_2885_0 & ((~i_10_159_459_0 & ((~i_10_159_1001_0 & ~i_10_159_1034_0 & i_10_159_1576_0 & ~i_10_159_3539_0 & ~i_10_159_3587_0 & ~i_10_159_3590_0) | (~i_10_159_1690_0 & ~i_10_159_2474_0 & ~i_10_159_3470_0 & i_10_159_3837_0 & ~i_10_159_3980_0 & ~i_10_159_4174_0))) | (~i_10_159_284_0 & ~i_10_159_796_0 & ~i_10_159_1655_0 & ~i_10_159_2381_0 & ~i_10_159_3473_0 & ~i_10_159_3584_0 & ~i_10_159_3841_0 & ~i_10_159_3842_0 & ~i_10_159_3853_0 & ~i_10_159_3980_0 & ~i_10_159_4568_0))) | (~i_10_159_1001_0 & ((i_10_159_800_0 & ((i_10_159_459_0 & ~i_10_159_1690_0 & ~i_10_159_2986_0) | (~i_10_159_1736_0 & ~i_10_159_2006_0 & i_10_159_3388_0 & ~i_10_159_4271_0))) | (~i_10_159_1034_0 & ~i_10_159_2474_0 & ((~i_10_159_1823_0 & ~i_10_159_2734_0 & ~i_10_159_3584_0 & ~i_10_159_3784_0) | (~i_10_159_2472_0 & ~i_10_159_2735_0 & ~i_10_159_3320_0 & ~i_10_159_3539_0 & i_10_159_3837_0 & ~i_10_159_4568_0))) | (~i_10_159_2033_0 & ((i_10_159_1654_0 & i_10_159_4114_0) | (i_10_159_442_0 & ~i_10_159_1823_0 & ~i_10_159_2006_0 & ~i_10_159_3088_0 & ~i_10_159_3473_0 & ~i_10_159_3890_0 & ~i_10_159_4174_0))) | (~i_10_159_796_0 & ~i_10_159_958_0 & ~i_10_159_1822_0 & ~i_10_159_1825_0 & ~i_10_159_3035_0 & ~i_10_159_3842_0))) | (~i_10_159_2474_0 & ~i_10_159_4268_0 & ((i_10_159_800_0 & ~i_10_159_3088_0 & ~i_10_159_3470_0) | (~i_10_159_1433_0 & ~i_10_159_2449_0 & ~i_10_159_2986_0 & ~i_10_159_3035_0 & ~i_10_159_3839_0 & i_10_159_4568_0))) | (~i_10_159_3839_0 & ((i_10_159_3784_0 & i_10_159_4174_0) | (i_10_159_2923_0 & ~i_10_159_3980_0 & ~i_10_159_4271_0))) | (~i_10_159_3980_0 & ((~i_10_159_2033_0 & i_10_159_2723_0 & ~i_10_159_2735_0 & ~i_10_159_3473_0) | (i_10_159_1825_0 & ~i_10_159_2730_0 & i_10_159_2922_0 & ~i_10_159_3890_0 & i_10_159_4568_0))) | (~i_10_159_1691_0 & ~i_10_159_1824_0 & ~i_10_159_2408_0 & i_10_159_3437_0) | (~i_10_159_1576_0 & ~i_10_159_1683_0 & ~i_10_159_1823_0 & i_10_159_3388_0 & ~i_10_159_3470_0) | (i_10_159_2634_0 & i_10_159_2722_0 & ~i_10_159_3590_0) | (i_10_159_2830_0 & i_10_159_2887_0 & i_10_159_3837_0) | (~i_10_159_1821_0 & i_10_159_4114_0 & i_10_159_4568_0));
endmodule



// Benchmark "kernel_10_160" written by ABC on Sun Jul 19 10:23:44 2020

module kernel_10_160 ( 
    i_10_160_34_0, i_10_160_153_0, i_10_160_220_0, i_10_160_248_0,
    i_10_160_256_0, i_10_160_272_0, i_10_160_286_0, i_10_160_327_0,
    i_10_160_330_0, i_10_160_358_0, i_10_160_466_0, i_10_160_495_0,
    i_10_160_504_0, i_10_160_513_0, i_10_160_637_0, i_10_160_711_0,
    i_10_160_954_0, i_10_160_963_0, i_10_160_1026_0, i_10_160_1031_0,
    i_10_160_1032_0, i_10_160_1162_0, i_10_160_1165_0, i_10_160_1241_0,
    i_10_160_1242_0, i_10_160_1309_0, i_10_160_1545_0, i_10_160_1546_0,
    i_10_160_1561_0, i_10_160_1635_0, i_10_160_1651_0, i_10_160_1690_0,
    i_10_160_1691_0, i_10_160_1794_0, i_10_160_1821_0, i_10_160_1823_0,
    i_10_160_1909_0, i_10_160_1947_0, i_10_160_1984_0, i_10_160_2182_0,
    i_10_160_2256_0, i_10_160_2257_0, i_10_160_2323_0, i_10_160_2353_0,
    i_10_160_2385_0, i_10_160_2386_0, i_10_160_2455_0, i_10_160_2629_0,
    i_10_160_2633_0, i_10_160_2824_0, i_10_160_2833_0, i_10_160_2871_0,
    i_10_160_2893_0, i_10_160_2923_0, i_10_160_2924_0, i_10_160_2953_0,
    i_10_160_2986_0, i_10_160_3036_0, i_10_160_3037_0, i_10_160_3069_0,
    i_10_160_3073_0, i_10_160_3202_0, i_10_160_3203_0, i_10_160_3234_0,
    i_10_160_3291_0, i_10_160_3385_0, i_10_160_3387_0, i_10_160_3390_0,
    i_10_160_3409_0, i_10_160_3465_0, i_10_160_3492_0, i_10_160_3537_0,
    i_10_160_3580_0, i_10_160_3612_0, i_10_160_3682_0, i_10_160_3683_0,
    i_10_160_3730_0, i_10_160_3732_0, i_10_160_3774_0, i_10_160_3786_0,
    i_10_160_3787_0, i_10_160_3801_0, i_10_160_3807_0, i_10_160_3826_0,
    i_10_160_3844_0, i_10_160_3858_0, i_10_160_3860_0, i_10_160_3992_0,
    i_10_160_4009_0, i_10_160_4117_0, i_10_160_4134_0, i_10_160_4216_0,
    i_10_160_4219_0, i_10_160_4263_0, i_10_160_4264_0, i_10_160_4305_0,
    i_10_160_4436_0, i_10_160_4486_0, i_10_160_4567_0, i_10_160_4584_0,
    o_10_160_0_0  );
  input  i_10_160_34_0, i_10_160_153_0, i_10_160_220_0, i_10_160_248_0,
    i_10_160_256_0, i_10_160_272_0, i_10_160_286_0, i_10_160_327_0,
    i_10_160_330_0, i_10_160_358_0, i_10_160_466_0, i_10_160_495_0,
    i_10_160_504_0, i_10_160_513_0, i_10_160_637_0, i_10_160_711_0,
    i_10_160_954_0, i_10_160_963_0, i_10_160_1026_0, i_10_160_1031_0,
    i_10_160_1032_0, i_10_160_1162_0, i_10_160_1165_0, i_10_160_1241_0,
    i_10_160_1242_0, i_10_160_1309_0, i_10_160_1545_0, i_10_160_1546_0,
    i_10_160_1561_0, i_10_160_1635_0, i_10_160_1651_0, i_10_160_1690_0,
    i_10_160_1691_0, i_10_160_1794_0, i_10_160_1821_0, i_10_160_1823_0,
    i_10_160_1909_0, i_10_160_1947_0, i_10_160_1984_0, i_10_160_2182_0,
    i_10_160_2256_0, i_10_160_2257_0, i_10_160_2323_0, i_10_160_2353_0,
    i_10_160_2385_0, i_10_160_2386_0, i_10_160_2455_0, i_10_160_2629_0,
    i_10_160_2633_0, i_10_160_2824_0, i_10_160_2833_0, i_10_160_2871_0,
    i_10_160_2893_0, i_10_160_2923_0, i_10_160_2924_0, i_10_160_2953_0,
    i_10_160_2986_0, i_10_160_3036_0, i_10_160_3037_0, i_10_160_3069_0,
    i_10_160_3073_0, i_10_160_3202_0, i_10_160_3203_0, i_10_160_3234_0,
    i_10_160_3291_0, i_10_160_3385_0, i_10_160_3387_0, i_10_160_3390_0,
    i_10_160_3409_0, i_10_160_3465_0, i_10_160_3492_0, i_10_160_3537_0,
    i_10_160_3580_0, i_10_160_3612_0, i_10_160_3682_0, i_10_160_3683_0,
    i_10_160_3730_0, i_10_160_3732_0, i_10_160_3774_0, i_10_160_3786_0,
    i_10_160_3787_0, i_10_160_3801_0, i_10_160_3807_0, i_10_160_3826_0,
    i_10_160_3844_0, i_10_160_3858_0, i_10_160_3860_0, i_10_160_3992_0,
    i_10_160_4009_0, i_10_160_4117_0, i_10_160_4134_0, i_10_160_4216_0,
    i_10_160_4219_0, i_10_160_4263_0, i_10_160_4264_0, i_10_160_4305_0,
    i_10_160_4436_0, i_10_160_4486_0, i_10_160_4567_0, i_10_160_4584_0;
  output o_10_160_0_0;
  assign o_10_160_0_0 = 0;
endmodule



// Benchmark "kernel_10_161" written by ABC on Sun Jul 19 10:23:46 2020

module kernel_10_161 ( 
    i_10_161_185_0, i_10_161_221_0, i_10_161_254_0, i_10_161_269_0,
    i_10_161_279_0, i_10_161_280_0, i_10_161_281_0, i_10_161_282_0,
    i_10_161_285_0, i_10_161_319_0, i_10_161_320_0, i_10_161_321_0,
    i_10_161_327_0, i_10_161_328_0, i_10_161_438_0, i_10_161_439_0,
    i_10_161_443_0, i_10_161_445_0, i_10_161_446_0, i_10_161_462_0,
    i_10_161_463_0, i_10_161_464_0, i_10_161_466_0, i_10_161_467_0,
    i_10_161_511_0, i_10_161_1030_0, i_10_161_1037_0, i_10_161_1240_0,
    i_10_161_1244_0, i_10_161_1245_0, i_10_161_1247_0, i_10_161_1248_0,
    i_10_161_1250_0, i_10_161_1363_0, i_10_161_1365_0, i_10_161_1546_0,
    i_10_161_1552_0, i_10_161_1554_0, i_10_161_1690_0, i_10_161_1819_0,
    i_10_161_1821_0, i_10_161_1822_0, i_10_161_1823_0, i_10_161_1945_0,
    i_10_161_1952_0, i_10_161_2185_0, i_10_161_2306_0, i_10_161_2323_0,
    i_10_161_2351_0, i_10_161_2353_0, i_10_161_2354_0, i_10_161_2355_0,
    i_10_161_2356_0, i_10_161_2467_0, i_10_161_2470_0, i_10_161_2515_0,
    i_10_161_2617_0, i_10_161_2630_0, i_10_161_2632_0, i_10_161_2634_0,
    i_10_161_2654_0, i_10_161_2662_0, i_10_161_2720_0, i_10_161_2724_0,
    i_10_161_2734_0, i_10_161_2735_0, i_10_161_2833_0, i_10_161_2887_0,
    i_10_161_2916_0, i_10_161_2919_0, i_10_161_2920_0, i_10_161_2921_0,
    i_10_161_2924_0, i_10_161_2986_0, i_10_161_3037_0, i_10_161_3038_0,
    i_10_161_3093_0, i_10_161_3154_0, i_10_161_3155_0, i_10_161_3163_0,
    i_10_161_3196_0, i_10_161_3197_0, i_10_161_3198_0, i_10_161_3199_0,
    i_10_161_3200_0, i_10_161_3281_0, i_10_161_3283_0, i_10_161_3328_0,
    i_10_161_3390_0, i_10_161_3407_0, i_10_161_3611_0, i_10_161_3650_0,
    i_10_161_3785_0, i_10_161_3838_0, i_10_161_3839_0, i_10_161_3842_0,
    i_10_161_4183_0, i_10_161_4569_0, i_10_161_4570_0, i_10_161_4571_0,
    o_10_161_0_0  );
  input  i_10_161_185_0, i_10_161_221_0, i_10_161_254_0, i_10_161_269_0,
    i_10_161_279_0, i_10_161_280_0, i_10_161_281_0, i_10_161_282_0,
    i_10_161_285_0, i_10_161_319_0, i_10_161_320_0, i_10_161_321_0,
    i_10_161_327_0, i_10_161_328_0, i_10_161_438_0, i_10_161_439_0,
    i_10_161_443_0, i_10_161_445_0, i_10_161_446_0, i_10_161_462_0,
    i_10_161_463_0, i_10_161_464_0, i_10_161_466_0, i_10_161_467_0,
    i_10_161_511_0, i_10_161_1030_0, i_10_161_1037_0, i_10_161_1240_0,
    i_10_161_1244_0, i_10_161_1245_0, i_10_161_1247_0, i_10_161_1248_0,
    i_10_161_1250_0, i_10_161_1363_0, i_10_161_1365_0, i_10_161_1546_0,
    i_10_161_1552_0, i_10_161_1554_0, i_10_161_1690_0, i_10_161_1819_0,
    i_10_161_1821_0, i_10_161_1822_0, i_10_161_1823_0, i_10_161_1945_0,
    i_10_161_1952_0, i_10_161_2185_0, i_10_161_2306_0, i_10_161_2323_0,
    i_10_161_2351_0, i_10_161_2353_0, i_10_161_2354_0, i_10_161_2355_0,
    i_10_161_2356_0, i_10_161_2467_0, i_10_161_2470_0, i_10_161_2515_0,
    i_10_161_2617_0, i_10_161_2630_0, i_10_161_2632_0, i_10_161_2634_0,
    i_10_161_2654_0, i_10_161_2662_0, i_10_161_2720_0, i_10_161_2724_0,
    i_10_161_2734_0, i_10_161_2735_0, i_10_161_2833_0, i_10_161_2887_0,
    i_10_161_2916_0, i_10_161_2919_0, i_10_161_2920_0, i_10_161_2921_0,
    i_10_161_2924_0, i_10_161_2986_0, i_10_161_3037_0, i_10_161_3038_0,
    i_10_161_3093_0, i_10_161_3154_0, i_10_161_3155_0, i_10_161_3163_0,
    i_10_161_3196_0, i_10_161_3197_0, i_10_161_3198_0, i_10_161_3199_0,
    i_10_161_3200_0, i_10_161_3281_0, i_10_161_3283_0, i_10_161_3328_0,
    i_10_161_3390_0, i_10_161_3407_0, i_10_161_3611_0, i_10_161_3650_0,
    i_10_161_3785_0, i_10_161_3838_0, i_10_161_3839_0, i_10_161_3842_0,
    i_10_161_4183_0, i_10_161_4569_0, i_10_161_4570_0, i_10_161_4571_0;
  output o_10_161_0_0;
  assign o_10_161_0_0 = ~((~i_10_161_439_0 & ((~i_10_161_1247_0 & ~i_10_161_1819_0 & i_10_161_1821_0 & ~i_10_161_2916_0 & ~i_10_161_3199_0 & ~i_10_161_3200_0) | (~i_10_161_254_0 & ~i_10_161_446_0 & ~i_10_161_467_0 & ~i_10_161_1037_0 & ~i_10_161_1244_0 & ~i_10_161_1245_0 & ~i_10_161_1363_0 & ~i_10_161_1365_0 & ~i_10_161_3093_0 & ~i_10_161_3650_0))) | (~i_10_161_1823_0 & ((i_10_161_463_0 & ((~i_10_161_269_0 & ~i_10_161_1244_0 & ~i_10_161_1363_0 & ~i_10_161_1365_0 & ~i_10_161_3198_0 & ~i_10_161_3199_0) | (~i_10_161_279_0 & ~i_10_161_281_0 & ~i_10_161_1690_0 & ~i_10_161_1821_0 & ~i_10_161_2617_0 & ~i_10_161_2724_0 & ~i_10_161_3283_0 & ~i_10_161_4571_0))) | (~i_10_161_2306_0 & i_10_161_2353_0) | (~i_10_161_254_0 & ~i_10_161_462_0 & ~i_10_161_463_0 & i_10_161_2916_0 & ~i_10_161_3038_0 & ~i_10_161_3093_0) | (i_10_161_280_0 & ~i_10_161_464_0 & ~i_10_161_1250_0 & ~i_10_161_2920_0 & ~i_10_161_4569_0))) | (~i_10_161_1037_0 & ((~i_10_161_254_0 & ~i_10_161_3093_0 & ((~i_10_161_445_0 & i_10_161_2920_0 & ~i_10_161_3038_0 & i_10_161_3197_0 & ~i_10_161_3198_0 & ~i_10_161_3281_0) | (~i_10_161_221_0 & ~i_10_161_446_0 & ~i_10_161_1245_0 & ~i_10_161_1365_0 & ~i_10_161_2355_0 & ~i_10_161_2735_0 & ~i_10_161_3839_0))) | (~i_10_161_3200_0 & ((~i_10_161_2634_0 & ~i_10_161_3197_0 & ~i_10_161_3198_0 & ~i_10_161_3650_0) | (~i_10_161_445_0 & ~i_10_161_2470_0 & ~i_10_161_3611_0 & ~i_10_161_4569_0))) | (~i_10_161_1365_0 & ~i_10_161_1821_0 & ~i_10_161_1822_0 & ~i_10_161_2323_0 & ~i_10_161_2354_0 & ~i_10_161_2724_0 & ~i_10_161_2735_0 & ~i_10_161_3196_0))) | (~i_10_161_1365_0 & ((~i_10_161_221_0 & ~i_10_161_1822_0 & ((~i_10_161_1247_0 & ~i_10_161_2617_0 & ~i_10_161_2735_0 & ~i_10_161_3197_0) | (~i_10_161_269_0 & ~i_10_161_280_0 & i_10_161_439_0 & ~i_10_161_1821_0 & ~i_10_161_3281_0))) | (~i_10_161_2306_0 & ((~i_10_161_2734_0 & ~i_10_161_2920_0 & ~i_10_161_2921_0 & ~i_10_161_3650_0) | (~i_10_161_185_0 & ~i_10_161_445_0 & ~i_10_161_1244_0 & ~i_10_161_1245_0 & ~i_10_161_1247_0 & ~i_10_161_1248_0 & ~i_10_161_2632_0 & ~i_10_161_2986_0 & i_10_161_3838_0 & i_10_161_3839_0))) | (~i_10_161_269_0 & ~i_10_161_1250_0 & ~i_10_161_2920_0 & ~i_10_161_2921_0 & ~i_10_161_3163_0 & ~i_10_161_3197_0 & ~i_10_161_3198_0))) | (i_10_161_1240_0 & ((i_10_161_2833_0 & ~i_10_161_2924_0) | (~i_10_161_3196_0 & ~i_10_161_3199_0 & ~i_10_161_3839_0))) | (~i_10_161_1244_0 & ((~i_10_161_221_0 & i_10_161_464_0 & ~i_10_161_466_0 & ~i_10_161_3197_0 & ~i_10_161_3198_0 & ~i_10_161_2916_0 & i_10_161_2921_0) | (~i_10_161_2734_0 & i_10_161_2919_0 & ~i_10_161_3200_0 & ~i_10_161_3650_0 & ~i_10_161_3838_0))) | (~i_10_161_3407_0 & ((~i_10_161_2185_0 & ((~i_10_161_1247_0 & ~i_10_161_1248_0 & ~i_10_161_1250_0 & ~i_10_161_2617_0 & ~i_10_161_2920_0 & ~i_10_161_3038_0) | (~i_10_161_3200_0 & i_10_161_3281_0 & ~i_10_161_3785_0))) | (~i_10_161_464_0 & ~i_10_161_3093_0 & ~i_10_161_3199_0) | (~i_10_161_285_0 & ~i_10_161_467_0 & ~i_10_161_1030_0 & ~i_10_161_1245_0 & ~i_10_161_1363_0 & ~i_10_161_2921_0 & ~i_10_161_3838_0))) | (~i_10_161_3650_0 & (i_10_161_1945_0 | (~i_10_161_1822_0 & i_10_161_2470_0))) | (i_10_161_328_0 & ~i_10_161_3196_0) | (~i_10_161_2634_0 & ~i_10_161_2921_0 & i_10_161_4570_0) | (i_10_161_1030_0 & ~i_10_161_2734_0 & ~i_10_161_3200_0 & ~i_10_161_4570_0));
endmodule



// Benchmark "kernel_10_162" written by ABC on Sun Jul 19 10:23:47 2020

module kernel_10_162 ( 
    i_10_162_30_0, i_10_162_123_0, i_10_162_174_0, i_10_162_178_0,
    i_10_162_183_0, i_10_162_221_0, i_10_162_429_0, i_10_162_430_0,
    i_10_162_464_0, i_10_162_500_0, i_10_162_535_0, i_10_162_564_0,
    i_10_162_898_0, i_10_162_951_0, i_10_162_996_0, i_10_162_1033_0,
    i_10_162_1114_0, i_10_162_1119_0, i_10_162_1237_0, i_10_162_1241_0,
    i_10_162_1309_0, i_10_162_1312_0, i_10_162_1345_0, i_10_162_1349_0,
    i_10_162_1489_0, i_10_162_1541_0, i_10_162_1542_0, i_10_162_1576_0,
    i_10_162_1618_0, i_10_162_1623_0, i_10_162_1624_0, i_10_162_1683_0,
    i_10_162_1684_0, i_10_162_1686_0, i_10_162_1768_0, i_10_162_1770_0,
    i_10_162_1824_0, i_10_162_1908_0, i_10_162_1912_0, i_10_162_1957_0,
    i_10_162_2004_0, i_10_162_2348_0, i_10_162_2364_0, i_10_162_2471_0,
    i_10_162_2515_0, i_10_162_2517_0, i_10_162_2519_0, i_10_162_2562_0,
    i_10_162_2567_0, i_10_162_2651_0, i_10_162_2652_0, i_10_162_2653_0,
    i_10_162_2658_0, i_10_162_2662_0, i_10_162_2715_0, i_10_162_2716_0,
    i_10_162_2722_0, i_10_162_2723_0, i_10_162_2725_0, i_10_162_2829_0,
    i_10_162_2830_0, i_10_162_2919_0, i_10_162_2966_0, i_10_162_2980_0,
    i_10_162_3071_0, i_10_162_3090_0, i_10_162_3093_0, i_10_162_3094_0,
    i_10_162_3166_0, i_10_162_3198_0, i_10_162_3199_0, i_10_162_3407_0,
    i_10_162_3410_0, i_10_162_3434_0, i_10_162_3472_0, i_10_162_3611_0,
    i_10_162_3612_0, i_10_162_3615_0, i_10_162_3624_0, i_10_162_3702_0,
    i_10_162_3705_0, i_10_162_3723_0, i_10_162_3797_0, i_10_162_3837_0,
    i_10_162_3855_0, i_10_162_3857_0, i_10_162_3883_0, i_10_162_3922_0,
    i_10_162_3982_0, i_10_162_3985_0, i_10_162_4026_0, i_10_162_4114_0,
    i_10_162_4117_0, i_10_162_4156_0, i_10_162_4175_0, i_10_162_4219_0,
    i_10_162_4236_0, i_10_162_4270_0, i_10_162_4425_0, i_10_162_4582_0,
    o_10_162_0_0  );
  input  i_10_162_30_0, i_10_162_123_0, i_10_162_174_0, i_10_162_178_0,
    i_10_162_183_0, i_10_162_221_0, i_10_162_429_0, i_10_162_430_0,
    i_10_162_464_0, i_10_162_500_0, i_10_162_535_0, i_10_162_564_0,
    i_10_162_898_0, i_10_162_951_0, i_10_162_996_0, i_10_162_1033_0,
    i_10_162_1114_0, i_10_162_1119_0, i_10_162_1237_0, i_10_162_1241_0,
    i_10_162_1309_0, i_10_162_1312_0, i_10_162_1345_0, i_10_162_1349_0,
    i_10_162_1489_0, i_10_162_1541_0, i_10_162_1542_0, i_10_162_1576_0,
    i_10_162_1618_0, i_10_162_1623_0, i_10_162_1624_0, i_10_162_1683_0,
    i_10_162_1684_0, i_10_162_1686_0, i_10_162_1768_0, i_10_162_1770_0,
    i_10_162_1824_0, i_10_162_1908_0, i_10_162_1912_0, i_10_162_1957_0,
    i_10_162_2004_0, i_10_162_2348_0, i_10_162_2364_0, i_10_162_2471_0,
    i_10_162_2515_0, i_10_162_2517_0, i_10_162_2519_0, i_10_162_2562_0,
    i_10_162_2567_0, i_10_162_2651_0, i_10_162_2652_0, i_10_162_2653_0,
    i_10_162_2658_0, i_10_162_2662_0, i_10_162_2715_0, i_10_162_2716_0,
    i_10_162_2722_0, i_10_162_2723_0, i_10_162_2725_0, i_10_162_2829_0,
    i_10_162_2830_0, i_10_162_2919_0, i_10_162_2966_0, i_10_162_2980_0,
    i_10_162_3071_0, i_10_162_3090_0, i_10_162_3093_0, i_10_162_3094_0,
    i_10_162_3166_0, i_10_162_3198_0, i_10_162_3199_0, i_10_162_3407_0,
    i_10_162_3410_0, i_10_162_3434_0, i_10_162_3472_0, i_10_162_3611_0,
    i_10_162_3612_0, i_10_162_3615_0, i_10_162_3624_0, i_10_162_3702_0,
    i_10_162_3705_0, i_10_162_3723_0, i_10_162_3797_0, i_10_162_3837_0,
    i_10_162_3855_0, i_10_162_3857_0, i_10_162_3883_0, i_10_162_3922_0,
    i_10_162_3982_0, i_10_162_3985_0, i_10_162_4026_0, i_10_162_4114_0,
    i_10_162_4117_0, i_10_162_4156_0, i_10_162_4175_0, i_10_162_4219_0,
    i_10_162_4236_0, i_10_162_4270_0, i_10_162_4425_0, i_10_162_4582_0;
  output o_10_162_0_0;
  assign o_10_162_0_0 = 0;
endmodule



// Benchmark "kernel_10_163" written by ABC on Sun Jul 19 10:23:48 2020

module kernel_10_163 ( 
    i_10_163_322_0, i_10_163_393_0, i_10_163_409_0, i_10_163_429_0,
    i_10_163_437_0, i_10_163_438_0, i_10_163_442_0, i_10_163_445_0,
    i_10_163_447_0, i_10_163_460_0, i_10_163_589_0, i_10_163_699_0,
    i_10_163_700_0, i_10_163_732_0, i_10_163_733_0, i_10_163_736_0,
    i_10_163_750_0, i_10_163_795_0, i_10_163_827_0, i_10_163_956_0,
    i_10_163_960_0, i_10_163_994_0, i_10_163_995_0, i_10_163_997_0,
    i_10_163_1060_0, i_10_163_1237_0, i_10_163_1238_0, i_10_163_1240_0,
    i_10_163_1241_0, i_10_163_1308_0, i_10_163_1343_0, i_10_163_1346_0,
    i_10_163_1576_0, i_10_163_1651_0, i_10_163_1684_0, i_10_163_1685_0,
    i_10_163_1688_0, i_10_163_1957_0, i_10_163_2184_0, i_10_163_2185_0,
    i_10_163_2364_0, i_10_163_2461_0, i_10_163_2463_0, i_10_163_2469_0,
    i_10_163_2470_0, i_10_163_2473_0, i_10_163_2632_0, i_10_163_2635_0,
    i_10_163_2659_0, i_10_163_2660_0, i_10_163_2698_0, i_10_163_2701_0,
    i_10_163_2702_0, i_10_163_2727_0, i_10_163_2728_0, i_10_163_2735_0,
    i_10_163_2821_0, i_10_163_2883_0, i_10_163_2884_0, i_10_163_2885_0,
    i_10_163_2886_0, i_10_163_2887_0, i_10_163_2888_0, i_10_163_2920_0,
    i_10_163_2922_0, i_10_163_2958_0, i_10_163_2959_0, i_10_163_3036_0,
    i_10_163_3037_0, i_10_163_3038_0, i_10_163_3198_0, i_10_163_3201_0,
    i_10_163_3202_0, i_10_163_3271_0, i_10_163_3279_0, i_10_163_3282_0,
    i_10_163_3283_0, i_10_163_3354_0, i_10_163_3406_0, i_10_163_3522_0,
    i_10_163_3543_0, i_10_163_3544_0, i_10_163_3588_0, i_10_163_3612_0,
    i_10_163_3702_0, i_10_163_3784_0, i_10_163_3787_0, i_10_163_3814_0,
    i_10_163_3837_0, i_10_163_3853_0, i_10_163_3854_0, i_10_163_3981_0,
    i_10_163_3984_0, i_10_163_3985_0, i_10_163_3989_0, i_10_163_4028_0,
    i_10_163_4119_0, i_10_163_4273_0, i_10_163_4285_0, i_10_163_4519_0,
    o_10_163_0_0  );
  input  i_10_163_322_0, i_10_163_393_0, i_10_163_409_0, i_10_163_429_0,
    i_10_163_437_0, i_10_163_438_0, i_10_163_442_0, i_10_163_445_0,
    i_10_163_447_0, i_10_163_460_0, i_10_163_589_0, i_10_163_699_0,
    i_10_163_700_0, i_10_163_732_0, i_10_163_733_0, i_10_163_736_0,
    i_10_163_750_0, i_10_163_795_0, i_10_163_827_0, i_10_163_956_0,
    i_10_163_960_0, i_10_163_994_0, i_10_163_995_0, i_10_163_997_0,
    i_10_163_1060_0, i_10_163_1237_0, i_10_163_1238_0, i_10_163_1240_0,
    i_10_163_1241_0, i_10_163_1308_0, i_10_163_1343_0, i_10_163_1346_0,
    i_10_163_1576_0, i_10_163_1651_0, i_10_163_1684_0, i_10_163_1685_0,
    i_10_163_1688_0, i_10_163_1957_0, i_10_163_2184_0, i_10_163_2185_0,
    i_10_163_2364_0, i_10_163_2461_0, i_10_163_2463_0, i_10_163_2469_0,
    i_10_163_2470_0, i_10_163_2473_0, i_10_163_2632_0, i_10_163_2635_0,
    i_10_163_2659_0, i_10_163_2660_0, i_10_163_2698_0, i_10_163_2701_0,
    i_10_163_2702_0, i_10_163_2727_0, i_10_163_2728_0, i_10_163_2735_0,
    i_10_163_2821_0, i_10_163_2883_0, i_10_163_2884_0, i_10_163_2885_0,
    i_10_163_2886_0, i_10_163_2887_0, i_10_163_2888_0, i_10_163_2920_0,
    i_10_163_2922_0, i_10_163_2958_0, i_10_163_2959_0, i_10_163_3036_0,
    i_10_163_3037_0, i_10_163_3038_0, i_10_163_3198_0, i_10_163_3201_0,
    i_10_163_3202_0, i_10_163_3271_0, i_10_163_3279_0, i_10_163_3282_0,
    i_10_163_3283_0, i_10_163_3354_0, i_10_163_3406_0, i_10_163_3522_0,
    i_10_163_3543_0, i_10_163_3544_0, i_10_163_3588_0, i_10_163_3612_0,
    i_10_163_3702_0, i_10_163_3784_0, i_10_163_3787_0, i_10_163_3814_0,
    i_10_163_3837_0, i_10_163_3853_0, i_10_163_3854_0, i_10_163_3981_0,
    i_10_163_3984_0, i_10_163_3985_0, i_10_163_3989_0, i_10_163_4028_0,
    i_10_163_4119_0, i_10_163_4273_0, i_10_163_4285_0, i_10_163_4519_0;
  output o_10_163_0_0;
  assign o_10_163_0_0 = 0;
endmodule



// Benchmark "kernel_10_164" written by ABC on Sun Jul 19 10:23:49 2020

module kernel_10_164 ( 
    i_10_164_46_0, i_10_164_223_0, i_10_164_243_0, i_10_164_244_0,
    i_10_164_245_0, i_10_164_285_0, i_10_164_315_0, i_10_164_316_0,
    i_10_164_360_0, i_10_164_445_0, i_10_164_712_0, i_10_164_956_0,
    i_10_164_1026_0, i_10_164_1028_0, i_10_164_1044_0, i_10_164_1235_0,
    i_10_164_1243_0, i_10_164_1308_0, i_10_164_1309_0, i_10_164_1539_0,
    i_10_164_1540_0, i_10_164_1541_0, i_10_164_1576_0, i_10_164_1579_0,
    i_10_164_1649_0, i_10_164_1650_0, i_10_164_1651_0, i_10_164_1683_0,
    i_10_164_1685_0, i_10_164_1686_0, i_10_164_1955_0, i_10_164_2016_0,
    i_10_164_2178_0, i_10_164_2179_0, i_10_164_2180_0, i_10_164_2199_0,
    i_10_164_2304_0, i_10_164_2305_0, i_10_164_2307_0, i_10_164_2351_0,
    i_10_164_2353_0, i_10_164_2354_0, i_10_164_2451_0, i_10_164_2452_0,
    i_10_164_2455_0, i_10_164_2470_0, i_10_164_2471_0, i_10_164_2545_0,
    i_10_164_2569_0, i_10_164_2601_0, i_10_164_2602_0, i_10_164_2605_0,
    i_10_164_2662_0, i_10_164_2678_0, i_10_164_2703_0, i_10_164_2704_0,
    i_10_164_2719_0, i_10_164_2726_0, i_10_164_2728_0, i_10_164_2730_0,
    i_10_164_2738_0, i_10_164_2826_0, i_10_164_2827_0, i_10_164_3071_0,
    i_10_164_3196_0, i_10_164_3199_0, i_10_164_3200_0, i_10_164_3270_0,
    i_10_164_3331_0, i_10_164_3403_0, i_10_164_3405_0, i_10_164_3406_0,
    i_10_164_3493_0, i_10_164_3583_0, i_10_164_3585_0, i_10_164_3586_0,
    i_10_164_3588_0, i_10_164_3612_0, i_10_164_3613_0, i_10_164_3614_0,
    i_10_164_3615_0, i_10_164_3616_0, i_10_164_3646_0, i_10_164_3647_0,
    i_10_164_3720_0, i_10_164_3780_0, i_10_164_3781_0, i_10_164_3782_0,
    i_10_164_3783_0, i_10_164_3784_0, i_10_164_3785_0, i_10_164_3834_0,
    i_10_164_3844_0, i_10_164_3857_0, i_10_164_3909_0, i_10_164_4114_0,
    i_10_164_4115_0, i_10_164_4169_0, i_10_164_4171_0, i_10_164_4212_0,
    o_10_164_0_0  );
  input  i_10_164_46_0, i_10_164_223_0, i_10_164_243_0, i_10_164_244_0,
    i_10_164_245_0, i_10_164_285_0, i_10_164_315_0, i_10_164_316_0,
    i_10_164_360_0, i_10_164_445_0, i_10_164_712_0, i_10_164_956_0,
    i_10_164_1026_0, i_10_164_1028_0, i_10_164_1044_0, i_10_164_1235_0,
    i_10_164_1243_0, i_10_164_1308_0, i_10_164_1309_0, i_10_164_1539_0,
    i_10_164_1540_0, i_10_164_1541_0, i_10_164_1576_0, i_10_164_1579_0,
    i_10_164_1649_0, i_10_164_1650_0, i_10_164_1651_0, i_10_164_1683_0,
    i_10_164_1685_0, i_10_164_1686_0, i_10_164_1955_0, i_10_164_2016_0,
    i_10_164_2178_0, i_10_164_2179_0, i_10_164_2180_0, i_10_164_2199_0,
    i_10_164_2304_0, i_10_164_2305_0, i_10_164_2307_0, i_10_164_2351_0,
    i_10_164_2353_0, i_10_164_2354_0, i_10_164_2451_0, i_10_164_2452_0,
    i_10_164_2455_0, i_10_164_2470_0, i_10_164_2471_0, i_10_164_2545_0,
    i_10_164_2569_0, i_10_164_2601_0, i_10_164_2602_0, i_10_164_2605_0,
    i_10_164_2662_0, i_10_164_2678_0, i_10_164_2703_0, i_10_164_2704_0,
    i_10_164_2719_0, i_10_164_2726_0, i_10_164_2728_0, i_10_164_2730_0,
    i_10_164_2738_0, i_10_164_2826_0, i_10_164_2827_0, i_10_164_3071_0,
    i_10_164_3196_0, i_10_164_3199_0, i_10_164_3200_0, i_10_164_3270_0,
    i_10_164_3331_0, i_10_164_3403_0, i_10_164_3405_0, i_10_164_3406_0,
    i_10_164_3493_0, i_10_164_3583_0, i_10_164_3585_0, i_10_164_3586_0,
    i_10_164_3588_0, i_10_164_3612_0, i_10_164_3613_0, i_10_164_3614_0,
    i_10_164_3615_0, i_10_164_3616_0, i_10_164_3646_0, i_10_164_3647_0,
    i_10_164_3720_0, i_10_164_3780_0, i_10_164_3781_0, i_10_164_3782_0,
    i_10_164_3783_0, i_10_164_3784_0, i_10_164_3785_0, i_10_164_3834_0,
    i_10_164_3844_0, i_10_164_3857_0, i_10_164_3909_0, i_10_164_4114_0,
    i_10_164_4115_0, i_10_164_4169_0, i_10_164_4171_0, i_10_164_4212_0;
  output o_10_164_0_0;
  assign o_10_164_0_0 = 0;
endmodule



// Benchmark "kernel_10_165" written by ABC on Sun Jul 19 10:23:50 2020

module kernel_10_165 ( 
    i_10_165_31_0, i_10_165_42_0, i_10_165_223_0, i_10_165_255_0,
    i_10_165_263_0, i_10_165_284_0, i_10_165_390_0, i_10_165_409_0,
    i_10_165_428_0, i_10_165_446_0, i_10_165_448_0, i_10_165_459_0,
    i_10_165_460_0, i_10_165_501_0, i_10_165_504_0, i_10_165_733_0,
    i_10_165_993_0, i_10_165_999_0, i_10_165_1001_0, i_10_165_1002_0,
    i_10_165_1180_0, i_10_165_1235_0, i_10_165_1238_0, i_10_165_1246_0,
    i_10_165_1542_0, i_10_165_1551_0, i_10_165_1552_0, i_10_165_1578_0,
    i_10_165_1582_0, i_10_165_1583_0, i_10_165_1623_0, i_10_165_1649_0,
    i_10_165_1651_0, i_10_165_1684_0, i_10_165_1731_0, i_10_165_1732_0,
    i_10_165_1734_0, i_10_165_1764_0, i_10_165_1806_0, i_10_165_1813_0,
    i_10_165_1823_0, i_10_165_1981_0, i_10_165_1983_0, i_10_165_1991_0,
    i_10_165_2154_0, i_10_165_2304_0, i_10_165_2352_0, i_10_165_2353_0,
    i_10_165_2377_0, i_10_165_2378_0, i_10_165_2379_0, i_10_165_2455_0,
    i_10_165_2456_0, i_10_165_2565_0, i_10_165_2567_0, i_10_165_2568_0,
    i_10_165_2658_0, i_10_165_2661_0, i_10_165_2701_0, i_10_165_2727_0,
    i_10_165_2829_0, i_10_165_2881_0, i_10_165_2884_0, i_10_165_2952_0,
    i_10_165_2953_0, i_10_165_2982_0, i_10_165_3033_0, i_10_165_3054_0,
    i_10_165_3232_0, i_10_165_3277_0, i_10_165_3316_0, i_10_165_3318_0,
    i_10_165_3384_0, i_10_165_3472_0, i_10_165_3538_0, i_10_165_3610_0,
    i_10_165_3614_0, i_10_165_3616_0, i_10_165_3782_0, i_10_165_3835_0,
    i_10_165_3851_0, i_10_165_3906_0, i_10_165_3978_0, i_10_165_3979_0,
    i_10_165_3988_0, i_10_165_4114_0, i_10_165_4116_0, i_10_165_4117_0,
    i_10_165_4124_0, i_10_165_4266_0, i_10_165_4267_0, i_10_165_4269_0,
    i_10_165_4272_0, i_10_165_4275_0, i_10_165_4278_0, i_10_165_4281_0,
    i_10_165_4287_0, i_10_165_4288_0, i_10_165_4290_0, i_10_165_4566_0,
    o_10_165_0_0  );
  input  i_10_165_31_0, i_10_165_42_0, i_10_165_223_0, i_10_165_255_0,
    i_10_165_263_0, i_10_165_284_0, i_10_165_390_0, i_10_165_409_0,
    i_10_165_428_0, i_10_165_446_0, i_10_165_448_0, i_10_165_459_0,
    i_10_165_460_0, i_10_165_501_0, i_10_165_504_0, i_10_165_733_0,
    i_10_165_993_0, i_10_165_999_0, i_10_165_1001_0, i_10_165_1002_0,
    i_10_165_1180_0, i_10_165_1235_0, i_10_165_1238_0, i_10_165_1246_0,
    i_10_165_1542_0, i_10_165_1551_0, i_10_165_1552_0, i_10_165_1578_0,
    i_10_165_1582_0, i_10_165_1583_0, i_10_165_1623_0, i_10_165_1649_0,
    i_10_165_1651_0, i_10_165_1684_0, i_10_165_1731_0, i_10_165_1732_0,
    i_10_165_1734_0, i_10_165_1764_0, i_10_165_1806_0, i_10_165_1813_0,
    i_10_165_1823_0, i_10_165_1981_0, i_10_165_1983_0, i_10_165_1991_0,
    i_10_165_2154_0, i_10_165_2304_0, i_10_165_2352_0, i_10_165_2353_0,
    i_10_165_2377_0, i_10_165_2378_0, i_10_165_2379_0, i_10_165_2455_0,
    i_10_165_2456_0, i_10_165_2565_0, i_10_165_2567_0, i_10_165_2568_0,
    i_10_165_2658_0, i_10_165_2661_0, i_10_165_2701_0, i_10_165_2727_0,
    i_10_165_2829_0, i_10_165_2881_0, i_10_165_2884_0, i_10_165_2952_0,
    i_10_165_2953_0, i_10_165_2982_0, i_10_165_3033_0, i_10_165_3054_0,
    i_10_165_3232_0, i_10_165_3277_0, i_10_165_3316_0, i_10_165_3318_0,
    i_10_165_3384_0, i_10_165_3472_0, i_10_165_3538_0, i_10_165_3610_0,
    i_10_165_3614_0, i_10_165_3616_0, i_10_165_3782_0, i_10_165_3835_0,
    i_10_165_3851_0, i_10_165_3906_0, i_10_165_3978_0, i_10_165_3979_0,
    i_10_165_3988_0, i_10_165_4114_0, i_10_165_4116_0, i_10_165_4117_0,
    i_10_165_4124_0, i_10_165_4266_0, i_10_165_4267_0, i_10_165_4269_0,
    i_10_165_4272_0, i_10_165_4275_0, i_10_165_4278_0, i_10_165_4281_0,
    i_10_165_4287_0, i_10_165_4288_0, i_10_165_4290_0, i_10_165_4566_0;
  output o_10_165_0_0;
  assign o_10_165_0_0 = ~((~i_10_165_999_0 & ((~i_10_165_1002_0 & ~i_10_165_1238_0 & i_10_165_1582_0 & ~i_10_165_1731_0 & ~i_10_165_2378_0) | (~i_10_165_263_0 & ~i_10_165_1578_0 & ~i_10_165_4278_0))) | (~i_10_165_1552_0 & ((~i_10_165_255_0 & ~i_10_165_459_0 & ~i_10_165_460_0 & ~i_10_165_1649_0 & i_10_165_1684_0 & ~i_10_165_2378_0 & ~i_10_165_2568_0 & ~i_10_165_3978_0 & ~i_10_165_3979_0) | (~i_10_165_1623_0 & ~i_10_165_1684_0 & ~i_10_165_3782_0 & ~i_10_165_3906_0 & i_10_165_3978_0 & ~i_10_165_4281_0))) | (~i_10_165_2353_0 & ((i_10_165_1551_0 & ~i_10_165_1651_0 & ~i_10_165_1731_0) | (i_10_165_1651_0 & ~i_10_165_1732_0 & ~i_10_165_2352_0 & ~i_10_165_2884_0))) | (i_10_165_3835_0 & ((~i_10_165_1582_0 & ~i_10_165_1731_0 & ~i_10_165_1732_0 & ~i_10_165_2377_0 & ~i_10_165_2379_0 & ~i_10_165_2565_0) | (i_10_165_1552_0 & ~i_10_165_2378_0 & ~i_10_165_3316_0 & ~i_10_165_4290_0))) | (~i_10_165_1731_0 & ~i_10_165_4278_0 & ((~i_10_165_1542_0 & ~i_10_165_2565_0 & ~i_10_165_2568_0 & ~i_10_165_3906_0 & ~i_10_165_3978_0) | (~i_10_165_1551_0 & ~i_10_165_4124_0 & ~i_10_165_4287_0 & ~i_10_165_4288_0))) | (~i_10_165_1732_0 & ((~i_10_165_2304_0 & ~i_10_165_2568_0 & ~i_10_165_3316_0 & ~i_10_165_3384_0 & ~i_10_165_3472_0 & ~i_10_165_3538_0 & ~i_10_165_3851_0 & ~i_10_165_3979_0) | (~i_10_165_2565_0 & ~i_10_165_3978_0 & ~i_10_165_4272_0 & ~i_10_165_4288_0))) | (~i_10_165_2377_0 & ((~i_10_165_1583_0 & ~i_10_165_3316_0 & i_10_165_3614_0) | (~i_10_165_2568_0 & ~i_10_165_2881_0 & ~i_10_165_3277_0 & ~i_10_165_4269_0))));
endmodule



// Benchmark "kernel_10_166" written by ABC on Sun Jul 19 10:23:51 2020

module kernel_10_166 ( 
    i_10_166_174_0, i_10_166_175_0, i_10_166_179_0, i_10_166_220_0,
    i_10_166_262_0, i_10_166_282_0, i_10_166_283_0, i_10_166_321_0,
    i_10_166_322_0, i_10_166_450_0, i_10_166_711_0, i_10_166_797_0,
    i_10_166_799_0, i_10_166_957_0, i_10_166_958_0, i_10_166_960_0,
    i_10_166_967_0, i_10_166_999_0, i_10_166_1000_0, i_10_166_1083_0,
    i_10_166_1135_0, i_10_166_1169_0, i_10_166_1237_0, i_10_166_1240_0,
    i_10_166_1308_0, i_10_166_1310_0, i_10_166_1438_0, i_10_166_1679_0,
    i_10_166_1684_0, i_10_166_1687_0, i_10_166_1688_0, i_10_166_1819_0,
    i_10_166_1821_0, i_10_166_1822_0, i_10_166_1909_0, i_10_166_1911_0,
    i_10_166_1944_0, i_10_166_1945_0, i_10_166_1946_0, i_10_166_2184_0,
    i_10_166_2185_0, i_10_166_2203_0, i_10_166_2331_0, i_10_166_2350_0,
    i_10_166_2352_0, i_10_166_2353_0, i_10_166_2356_0, i_10_166_2376_0,
    i_10_166_2377_0, i_10_166_2404_0, i_10_166_2449_0, i_10_166_2452_0,
    i_10_166_2470_0, i_10_166_2502_0, i_10_166_2504_0, i_10_166_2711_0,
    i_10_166_2713_0, i_10_166_2716_0, i_10_166_2729_0, i_10_166_2734_0,
    i_10_166_2788_0, i_10_166_2880_0, i_10_166_2881_0, i_10_166_2885_0,
    i_10_166_2923_0, i_10_166_3034_0, i_10_166_3036_0, i_10_166_3042_0,
    i_10_166_3044_0, i_10_166_3150_0, i_10_166_3279_0, i_10_166_3280_0,
    i_10_166_3493_0, i_10_166_3610_0, i_10_166_3614_0, i_10_166_3687_0,
    i_10_166_3783_0, i_10_166_3786_0, i_10_166_3838_0, i_10_166_3840_0,
    i_10_166_3841_0, i_10_166_3843_0, i_10_166_3847_0, i_10_166_3851_0,
    i_10_166_3860_0, i_10_166_3877_0, i_10_166_3889_0, i_10_166_3978_0,
    i_10_166_3979_0, i_10_166_4050_0, i_10_166_4117_0, i_10_166_4122_0,
    i_10_166_4123_0, i_10_166_4129_0, i_10_166_4290_0, i_10_166_4291_0,
    i_10_166_4292_0, i_10_166_4564_0, i_10_166_4566_0, i_10_166_4567_0,
    o_10_166_0_0  );
  input  i_10_166_174_0, i_10_166_175_0, i_10_166_179_0, i_10_166_220_0,
    i_10_166_262_0, i_10_166_282_0, i_10_166_283_0, i_10_166_321_0,
    i_10_166_322_0, i_10_166_450_0, i_10_166_711_0, i_10_166_797_0,
    i_10_166_799_0, i_10_166_957_0, i_10_166_958_0, i_10_166_960_0,
    i_10_166_967_0, i_10_166_999_0, i_10_166_1000_0, i_10_166_1083_0,
    i_10_166_1135_0, i_10_166_1169_0, i_10_166_1237_0, i_10_166_1240_0,
    i_10_166_1308_0, i_10_166_1310_0, i_10_166_1438_0, i_10_166_1679_0,
    i_10_166_1684_0, i_10_166_1687_0, i_10_166_1688_0, i_10_166_1819_0,
    i_10_166_1821_0, i_10_166_1822_0, i_10_166_1909_0, i_10_166_1911_0,
    i_10_166_1944_0, i_10_166_1945_0, i_10_166_1946_0, i_10_166_2184_0,
    i_10_166_2185_0, i_10_166_2203_0, i_10_166_2331_0, i_10_166_2350_0,
    i_10_166_2352_0, i_10_166_2353_0, i_10_166_2356_0, i_10_166_2376_0,
    i_10_166_2377_0, i_10_166_2404_0, i_10_166_2449_0, i_10_166_2452_0,
    i_10_166_2470_0, i_10_166_2502_0, i_10_166_2504_0, i_10_166_2711_0,
    i_10_166_2713_0, i_10_166_2716_0, i_10_166_2729_0, i_10_166_2734_0,
    i_10_166_2788_0, i_10_166_2880_0, i_10_166_2881_0, i_10_166_2885_0,
    i_10_166_2923_0, i_10_166_3034_0, i_10_166_3036_0, i_10_166_3042_0,
    i_10_166_3044_0, i_10_166_3150_0, i_10_166_3279_0, i_10_166_3280_0,
    i_10_166_3493_0, i_10_166_3610_0, i_10_166_3614_0, i_10_166_3687_0,
    i_10_166_3783_0, i_10_166_3786_0, i_10_166_3838_0, i_10_166_3840_0,
    i_10_166_3841_0, i_10_166_3843_0, i_10_166_3847_0, i_10_166_3851_0,
    i_10_166_3860_0, i_10_166_3877_0, i_10_166_3889_0, i_10_166_3978_0,
    i_10_166_3979_0, i_10_166_4050_0, i_10_166_4117_0, i_10_166_4122_0,
    i_10_166_4123_0, i_10_166_4129_0, i_10_166_4290_0, i_10_166_4291_0,
    i_10_166_4292_0, i_10_166_4564_0, i_10_166_4566_0, i_10_166_4567_0;
  output o_10_166_0_0;
  assign o_10_166_0_0 = ~((~i_10_166_282_0 & ((~i_10_166_322_0 & ~i_10_166_958_0 & ~i_10_166_1821_0 & ~i_10_166_1944_0 & ~i_10_166_1945_0 & ~i_10_166_1946_0 & ~i_10_166_2711_0 & ~i_10_166_3042_0 & ~i_10_166_3493_0 & ~i_10_166_3843_0 & ~i_10_166_3978_0 & ~i_10_166_4122_0) | (~i_10_166_2185_0 & ~i_10_166_2352_0 & ~i_10_166_2377_0 & ~i_10_166_3786_0 & i_10_166_3847_0 & ~i_10_166_4567_0))) | (~i_10_166_450_0 & ((i_10_166_174_0 & i_10_166_1821_0 & ~i_10_166_2502_0 & ~i_10_166_3838_0 & ~i_10_166_3978_0 & ~i_10_166_4290_0) | (~i_10_166_958_0 & ~i_10_166_960_0 & ~i_10_166_999_0 & ~i_10_166_1240_0 & ~i_10_166_2376_0 & ~i_10_166_2504_0 & ~i_10_166_3687_0 & ~i_10_166_3843_0 & ~i_10_166_3979_0 & ~i_10_166_4291_0 & ~i_10_166_4564_0))) | (~i_10_166_2377_0 & ((i_10_166_799_0 & ((~i_10_166_999_0 & ~i_10_166_1438_0 & ~i_10_166_2185_0 & ~i_10_166_2502_0 & ~i_10_166_3860_0) | (~i_10_166_958_0 & ~i_10_166_1944_0 & ~i_10_166_2184_0 & ~i_10_166_4564_0))) | (~i_10_166_4123_0 & ((~i_10_166_957_0 & ~i_10_166_2376_0 & ((~i_10_166_262_0 & ~i_10_166_3687_0 & ~i_10_166_3786_0 & i_10_166_3838_0) | (~i_10_166_960_0 & ~i_10_166_1438_0 & ~i_10_166_1945_0 & ~i_10_166_2184_0 & ~i_10_166_2504_0 & ~i_10_166_3036_0 & ~i_10_166_4122_0))) | (~i_10_166_960_0 & ~i_10_166_1944_0 & ~i_10_166_2404_0 & i_10_166_3280_0))) | (~i_10_166_1000_0 & ~i_10_166_3614_0 & ~i_10_166_3786_0 & ~i_10_166_3889_0 & i_10_166_4129_0))) | (~i_10_166_2729_0 & ((~i_10_166_999_0 & ((~i_10_166_960_0 & ~i_10_166_1944_0 & i_10_166_2881_0 & i_10_166_3610_0 & ~i_10_166_3847_0) | (~i_10_166_1169_0 & ~i_10_166_1438_0 & ~i_10_166_1822_0 & ~i_10_166_2184_0 & ~i_10_166_2356_0 & ~i_10_166_2376_0 & ~i_10_166_2470_0 & ~i_10_166_3889_0 & ~i_10_166_4567_0))) | (~i_10_166_3036_0 & i_10_166_3687_0 & i_10_166_3838_0))) | (~i_10_166_1240_0 & ((~i_10_166_2350_0 & i_10_166_2352_0 & i_10_166_2880_0 & ~i_10_166_3851_0) | (~i_10_166_175_0 & ~i_10_166_179_0 & ~i_10_166_2184_0 & ~i_10_166_2185_0 & i_10_166_2203_0 & ~i_10_166_2404_0 & ~i_10_166_2504_0 & ~i_10_166_3042_0 & ~i_10_166_3044_0 & ~i_10_166_4567_0))) | (~i_10_166_3847_0 & ((i_10_166_1819_0 & ((i_10_166_1684_0 & ~i_10_166_1945_0) | (~i_10_166_1000_0 & ~i_10_166_1944_0 & ~i_10_166_2184_0 & ~i_10_166_2331_0 & ~i_10_166_3843_0))) | (~i_10_166_1909_0 & ~i_10_166_1911_0 & i_10_166_2350_0 & i_10_166_3610_0 & ~i_10_166_4050_0 & ~i_10_166_4566_0))) | (~i_10_166_1000_0 & ((~i_10_166_967_0 & ~i_10_166_1083_0 & i_10_166_1822_0 & ~i_10_166_2185_0 & ~i_10_166_2352_0 & ~i_10_166_2356_0 & ~i_10_166_2502_0 & ~i_10_166_3044_0 & ~i_10_166_4122_0) | (i_10_166_2356_0 & ~i_10_166_2404_0 & ~i_10_166_4117_0 & ~i_10_166_4123_0 & i_10_166_4566_0))) | (~i_10_166_2376_0 & ((~i_10_166_960_0 & ~i_10_166_4123_0 & ((~i_10_166_2350_0 & ~i_10_166_2502_0 & ~i_10_166_3687_0 & ~i_10_166_3786_0 & ~i_10_166_3889_0 & i_10_166_4566_0) | (~i_10_166_321_0 & ~i_10_166_967_0 & ~i_10_166_1438_0 & ~i_10_166_1822_0 & ~i_10_166_1945_0 & ~i_10_166_2788_0 & ~i_10_166_3036_0 & ~i_10_166_4290_0 & ~i_10_166_4566_0))) | (~i_10_166_1946_0 & ((~i_10_166_1821_0 & i_10_166_2711_0 & ~i_10_166_3042_0 & ~i_10_166_3786_0 & ~i_10_166_4564_0) | (~i_10_166_797_0 & i_10_166_1822_0 & ~i_10_166_2203_0 & ~i_10_166_2352_0 & ~i_10_166_3860_0 & ~i_10_166_3978_0 & ~i_10_166_3979_0 & ~i_10_166_4566_0))) | (~i_10_166_3978_0 & ((~i_10_166_957_0 & ~i_10_166_967_0 & i_10_166_2353_0 & ~i_10_166_3034_0 & ~i_10_166_3851_0 & ~i_10_166_3979_0 & ~i_10_166_4292_0 & ~i_10_166_4566_0) | (~i_10_166_1688_0 & ~i_10_166_2404_0 & ~i_10_166_2502_0 & ~i_10_166_3036_0 & ~i_10_166_4050_0 & i_10_166_4117_0 & ~i_10_166_4564_0 & ~i_10_166_4567_0))))) | (~i_10_166_283_0 & ~i_10_166_960_0 & ~i_10_166_1169_0 & i_10_166_1308_0 & i_10_166_3841_0) | (i_10_166_1240_0 & ~i_10_166_1944_0 & ~i_10_166_2185_0 & ~i_10_166_3979_0 & ~i_10_166_4566_0 & ~i_10_166_2504_0 & ~i_10_166_2881_0) | (i_10_166_3840_0 & ~i_10_166_3843_0 & ~i_10_166_3978_0 & ~i_10_166_4050_0 & ~i_10_166_4567_0));
endmodule



// Benchmark "kernel_10_167" written by ABC on Sun Jul 19 10:23:53 2020

module kernel_10_167 ( 
    i_10_167_33_0, i_10_167_174_0, i_10_167_175_0, i_10_167_178_0,
    i_10_167_285_0, i_10_167_286_0, i_10_167_332_0, i_10_167_390_0,
    i_10_167_442_0, i_10_167_447_0, i_10_167_448_0, i_10_167_459_0,
    i_10_167_460_0, i_10_167_467_0, i_10_167_800_0, i_10_167_1029_0,
    i_10_167_1034_0, i_10_167_1237_0, i_10_167_1238_0, i_10_167_1239_0,
    i_10_167_1308_0, i_10_167_1309_0, i_10_167_1545_0, i_10_167_1619_0,
    i_10_167_1648_0, i_10_167_1651_0, i_10_167_1687_0, i_10_167_1767_0,
    i_10_167_1769_0, i_10_167_1824_0, i_10_167_1825_0, i_10_167_1912_0,
    i_10_167_1950_0, i_10_167_1951_0, i_10_167_1952_0, i_10_167_1961_0,
    i_10_167_2004_0, i_10_167_2019_0, i_10_167_2185_0, i_10_167_2186_0,
    i_10_167_2436_0, i_10_167_2455_0, i_10_167_2515_0, i_10_167_2516_0,
    i_10_167_2631_0, i_10_167_2634_0, i_10_167_2635_0, i_10_167_2656_0,
    i_10_167_2707_0, i_10_167_2708_0, i_10_167_2710_0, i_10_167_2718_0,
    i_10_167_2723_0, i_10_167_2731_0, i_10_167_2757_0, i_10_167_2782_0,
    i_10_167_2788_0, i_10_167_2827_0, i_10_167_3036_0, i_10_167_3037_0,
    i_10_167_3040_0, i_10_167_3093_0, i_10_167_3094_0, i_10_167_3095_0,
    i_10_167_3198_0, i_10_167_3199_0, i_10_167_3202_0, i_10_167_3277_0,
    i_10_167_3278_0, i_10_167_3279_0, i_10_167_3280_0, i_10_167_3328_0,
    i_10_167_3407_0, i_10_167_3433_0, i_10_167_3466_0, i_10_167_3468_0,
    i_10_167_3469_0, i_10_167_3494_0, i_10_167_3496_0, i_10_167_3610_0,
    i_10_167_3613_0, i_10_167_3614_0, i_10_167_3650_0, i_10_167_3652_0,
    i_10_167_3702_0, i_10_167_3783_0, i_10_167_3784_0, i_10_167_3786_0,
    i_10_167_3838_0, i_10_167_3842_0, i_10_167_3855_0, i_10_167_3856_0,
    i_10_167_3857_0, i_10_167_3985_0, i_10_167_3991_0, i_10_167_4126_0,
    i_10_167_4129_0, i_10_167_4130_0, i_10_167_4273_0, i_10_167_4565_0,
    o_10_167_0_0  );
  input  i_10_167_33_0, i_10_167_174_0, i_10_167_175_0, i_10_167_178_0,
    i_10_167_285_0, i_10_167_286_0, i_10_167_332_0, i_10_167_390_0,
    i_10_167_442_0, i_10_167_447_0, i_10_167_448_0, i_10_167_459_0,
    i_10_167_460_0, i_10_167_467_0, i_10_167_800_0, i_10_167_1029_0,
    i_10_167_1034_0, i_10_167_1237_0, i_10_167_1238_0, i_10_167_1239_0,
    i_10_167_1308_0, i_10_167_1309_0, i_10_167_1545_0, i_10_167_1619_0,
    i_10_167_1648_0, i_10_167_1651_0, i_10_167_1687_0, i_10_167_1767_0,
    i_10_167_1769_0, i_10_167_1824_0, i_10_167_1825_0, i_10_167_1912_0,
    i_10_167_1950_0, i_10_167_1951_0, i_10_167_1952_0, i_10_167_1961_0,
    i_10_167_2004_0, i_10_167_2019_0, i_10_167_2185_0, i_10_167_2186_0,
    i_10_167_2436_0, i_10_167_2455_0, i_10_167_2515_0, i_10_167_2516_0,
    i_10_167_2631_0, i_10_167_2634_0, i_10_167_2635_0, i_10_167_2656_0,
    i_10_167_2707_0, i_10_167_2708_0, i_10_167_2710_0, i_10_167_2718_0,
    i_10_167_2723_0, i_10_167_2731_0, i_10_167_2757_0, i_10_167_2782_0,
    i_10_167_2788_0, i_10_167_2827_0, i_10_167_3036_0, i_10_167_3037_0,
    i_10_167_3040_0, i_10_167_3093_0, i_10_167_3094_0, i_10_167_3095_0,
    i_10_167_3198_0, i_10_167_3199_0, i_10_167_3202_0, i_10_167_3277_0,
    i_10_167_3278_0, i_10_167_3279_0, i_10_167_3280_0, i_10_167_3328_0,
    i_10_167_3407_0, i_10_167_3433_0, i_10_167_3466_0, i_10_167_3468_0,
    i_10_167_3469_0, i_10_167_3494_0, i_10_167_3496_0, i_10_167_3610_0,
    i_10_167_3613_0, i_10_167_3614_0, i_10_167_3650_0, i_10_167_3652_0,
    i_10_167_3702_0, i_10_167_3783_0, i_10_167_3784_0, i_10_167_3786_0,
    i_10_167_3838_0, i_10_167_3842_0, i_10_167_3855_0, i_10_167_3856_0,
    i_10_167_3857_0, i_10_167_3985_0, i_10_167_3991_0, i_10_167_4126_0,
    i_10_167_4129_0, i_10_167_4130_0, i_10_167_4273_0, i_10_167_4565_0;
  output o_10_167_0_0;
  assign o_10_167_0_0 = ~((~i_10_167_467_0 & (i_10_167_1824_0 | (~i_10_167_332_0 & i_10_167_390_0 & ~i_10_167_3652_0 & ~i_10_167_3838_0 & ~i_10_167_3842_0))) | (~i_10_167_1619_0 & (~i_10_167_2634_0 | ~i_10_167_3093_0)) | (~i_10_167_2827_0 & ((~i_10_167_390_0 & ~i_10_167_2631_0 & ~i_10_167_3407_0) | (~i_10_167_447_0 & ~i_10_167_3094_0 & ~i_10_167_3783_0 & i_10_167_3855_0))) | (~i_10_167_3279_0 & ((~i_10_167_1308_0 & ~i_10_167_2185_0) | (~i_10_167_3094_0 & ~i_10_167_3856_0))) | (i_10_167_1825_0 & ~i_10_167_3650_0 & ~i_10_167_3784_0) | (i_10_167_285_0 & ~i_10_167_3855_0) | (i_10_167_4126_0 & ~i_10_167_4273_0) | (~i_10_167_3985_0 & ~i_10_167_4565_0));
endmodule



// Benchmark "kernel_10_168" written by ABC on Sun Jul 19 10:23:53 2020

module kernel_10_168 ( 
    i_10_168_30_0, i_10_168_69_0, i_10_168_193_0, i_10_168_279_0,
    i_10_168_285_0, i_10_168_387_0, i_10_168_390_0, i_10_168_393_0,
    i_10_168_426_0, i_10_168_445_0, i_10_168_462_0, i_10_168_463_0,
    i_10_168_465_0, i_10_168_480_0, i_10_168_759_0, i_10_168_826_0,
    i_10_168_950_0, i_10_168_1029_0, i_10_168_1030_0, i_10_168_1031_0,
    i_10_168_1034_0, i_10_168_1260_0, i_10_168_1261_0, i_10_168_1262_0,
    i_10_168_1308_0, i_10_168_1353_0, i_10_168_1435_0, i_10_168_1498_0,
    i_10_168_1548_0, i_10_168_1579_0, i_10_168_1581_0, i_10_168_1617_0,
    i_10_168_1623_0, i_10_168_1650_0, i_10_168_1687_0, i_10_168_1691_0,
    i_10_168_1743_0, i_10_168_1756_0, i_10_168_1759_0, i_10_168_1803_0,
    i_10_168_1918_0, i_10_168_2164_0, i_10_168_2196_0, i_10_168_2198_0,
    i_10_168_2307_0, i_10_168_2311_0, i_10_168_2312_0, i_10_168_2338_0,
    i_10_168_2351_0, i_10_168_2352_0, i_10_168_2362_0, i_10_168_2433_0,
    i_10_168_2457_0, i_10_168_2460_0, i_10_168_2472_0, i_10_168_2559_0,
    i_10_168_2565_0, i_10_168_2568_0, i_10_168_2631_0, i_10_168_2634_0,
    i_10_168_2661_0, i_10_168_2830_0, i_10_168_2845_0, i_10_168_2865_0,
    i_10_168_3072_0, i_10_168_3201_0, i_10_168_3202_0, i_10_168_3267_0,
    i_10_168_3268_0, i_10_168_3333_0, i_10_168_3334_0, i_10_168_3392_0,
    i_10_168_3406_0, i_10_168_3465_0, i_10_168_3468_0, i_10_168_3609_0,
    i_10_168_3612_0, i_10_168_3615_0, i_10_168_3681_0, i_10_168_3685_0,
    i_10_168_3686_0, i_10_168_3688_0, i_10_168_3706_0, i_10_168_3727_0,
    i_10_168_3777_0, i_10_168_3781_0, i_10_168_3843_0, i_10_168_3844_0,
    i_10_168_3993_0, i_10_168_4098_0, i_10_168_4113_0, i_10_168_4121_0,
    i_10_168_4175_0, i_10_168_4218_0, i_10_168_4236_0, i_10_168_4290_0,
    i_10_168_4458_0, i_10_168_4477_0, i_10_168_4478_0, i_10_168_4561_0,
    o_10_168_0_0  );
  input  i_10_168_30_0, i_10_168_69_0, i_10_168_193_0, i_10_168_279_0,
    i_10_168_285_0, i_10_168_387_0, i_10_168_390_0, i_10_168_393_0,
    i_10_168_426_0, i_10_168_445_0, i_10_168_462_0, i_10_168_463_0,
    i_10_168_465_0, i_10_168_480_0, i_10_168_759_0, i_10_168_826_0,
    i_10_168_950_0, i_10_168_1029_0, i_10_168_1030_0, i_10_168_1031_0,
    i_10_168_1034_0, i_10_168_1260_0, i_10_168_1261_0, i_10_168_1262_0,
    i_10_168_1308_0, i_10_168_1353_0, i_10_168_1435_0, i_10_168_1498_0,
    i_10_168_1548_0, i_10_168_1579_0, i_10_168_1581_0, i_10_168_1617_0,
    i_10_168_1623_0, i_10_168_1650_0, i_10_168_1687_0, i_10_168_1691_0,
    i_10_168_1743_0, i_10_168_1756_0, i_10_168_1759_0, i_10_168_1803_0,
    i_10_168_1918_0, i_10_168_2164_0, i_10_168_2196_0, i_10_168_2198_0,
    i_10_168_2307_0, i_10_168_2311_0, i_10_168_2312_0, i_10_168_2338_0,
    i_10_168_2351_0, i_10_168_2352_0, i_10_168_2362_0, i_10_168_2433_0,
    i_10_168_2457_0, i_10_168_2460_0, i_10_168_2472_0, i_10_168_2559_0,
    i_10_168_2565_0, i_10_168_2568_0, i_10_168_2631_0, i_10_168_2634_0,
    i_10_168_2661_0, i_10_168_2830_0, i_10_168_2845_0, i_10_168_2865_0,
    i_10_168_3072_0, i_10_168_3201_0, i_10_168_3202_0, i_10_168_3267_0,
    i_10_168_3268_0, i_10_168_3333_0, i_10_168_3334_0, i_10_168_3392_0,
    i_10_168_3406_0, i_10_168_3465_0, i_10_168_3468_0, i_10_168_3609_0,
    i_10_168_3612_0, i_10_168_3615_0, i_10_168_3681_0, i_10_168_3685_0,
    i_10_168_3686_0, i_10_168_3688_0, i_10_168_3706_0, i_10_168_3727_0,
    i_10_168_3777_0, i_10_168_3781_0, i_10_168_3843_0, i_10_168_3844_0,
    i_10_168_3993_0, i_10_168_4098_0, i_10_168_4113_0, i_10_168_4121_0,
    i_10_168_4175_0, i_10_168_4218_0, i_10_168_4236_0, i_10_168_4290_0,
    i_10_168_4458_0, i_10_168_4477_0, i_10_168_4478_0, i_10_168_4561_0;
  output o_10_168_0_0;
  assign o_10_168_0_0 = 0;
endmodule



// Benchmark "kernel_10_169" written by ABC on Sun Jul 19 10:23:55 2020

module kernel_10_169 ( 
    i_10_169_172_0, i_10_169_178_0, i_10_169_279_0, i_10_169_280_0,
    i_10_169_282_0, i_10_169_423_0, i_10_169_428_0, i_10_169_429_0,
    i_10_169_430_0, i_10_169_433_0, i_10_169_435_0, i_10_169_436_0,
    i_10_169_438_0, i_10_169_439_0, i_10_169_440_0, i_10_169_441_0,
    i_10_169_447_0, i_10_169_465_0, i_10_169_507_0, i_10_169_717_0,
    i_10_169_748_0, i_10_169_751_0, i_10_169_793_0, i_10_169_800_0,
    i_10_169_1137_0, i_10_169_1138_0, i_10_169_1237_0, i_10_169_1238_0,
    i_10_169_1249_0, i_10_169_1305_0, i_10_169_1306_0, i_10_169_1308_0,
    i_10_169_1309_0, i_10_169_1579_0, i_10_169_1647_0, i_10_169_1683_0,
    i_10_169_1687_0, i_10_169_1819_0, i_10_169_1820_0, i_10_169_1823_0,
    i_10_169_2350_0, i_10_169_2351_0, i_10_169_2352_0, i_10_169_2353_0,
    i_10_169_2354_0, i_10_169_2453_0, i_10_169_2514_0, i_10_169_2516_0,
    i_10_169_2629_0, i_10_169_2634_0, i_10_169_2636_0, i_10_169_2703_0,
    i_10_169_2704_0, i_10_169_2706_0, i_10_169_2715_0, i_10_169_2718_0,
    i_10_169_2884_0, i_10_169_2885_0, i_10_169_2980_0, i_10_169_2986_0,
    i_10_169_3034_0, i_10_169_3036_0, i_10_169_3087_0, i_10_169_3093_0,
    i_10_169_3094_0, i_10_169_3154_0, i_10_169_3155_0, i_10_169_3165_0,
    i_10_169_3196_0, i_10_169_3198_0, i_10_169_3199_0, i_10_169_3200_0,
    i_10_169_3321_0, i_10_169_3322_0, i_10_169_3384_0, i_10_169_3405_0,
    i_10_169_3406_0, i_10_169_3407_0, i_10_169_3408_0, i_10_169_3409_0,
    i_10_169_3610_0, i_10_169_3613_0, i_10_169_3614_0, i_10_169_3615_0,
    i_10_169_3650_0, i_10_169_3702_0, i_10_169_3780_0, i_10_169_3782_0,
    i_10_169_3788_0, i_10_169_3837_0, i_10_169_3846_0, i_10_169_3856_0,
    i_10_169_3859_0, i_10_169_3982_0, i_10_169_4115_0, i_10_169_4273_0,
    i_10_169_4288_0, i_10_169_4564_0, i_10_169_4565_0, i_10_169_4568_0,
    o_10_169_0_0  );
  input  i_10_169_172_0, i_10_169_178_0, i_10_169_279_0, i_10_169_280_0,
    i_10_169_282_0, i_10_169_423_0, i_10_169_428_0, i_10_169_429_0,
    i_10_169_430_0, i_10_169_433_0, i_10_169_435_0, i_10_169_436_0,
    i_10_169_438_0, i_10_169_439_0, i_10_169_440_0, i_10_169_441_0,
    i_10_169_447_0, i_10_169_465_0, i_10_169_507_0, i_10_169_717_0,
    i_10_169_748_0, i_10_169_751_0, i_10_169_793_0, i_10_169_800_0,
    i_10_169_1137_0, i_10_169_1138_0, i_10_169_1237_0, i_10_169_1238_0,
    i_10_169_1249_0, i_10_169_1305_0, i_10_169_1306_0, i_10_169_1308_0,
    i_10_169_1309_0, i_10_169_1579_0, i_10_169_1647_0, i_10_169_1683_0,
    i_10_169_1687_0, i_10_169_1819_0, i_10_169_1820_0, i_10_169_1823_0,
    i_10_169_2350_0, i_10_169_2351_0, i_10_169_2352_0, i_10_169_2353_0,
    i_10_169_2354_0, i_10_169_2453_0, i_10_169_2514_0, i_10_169_2516_0,
    i_10_169_2629_0, i_10_169_2634_0, i_10_169_2636_0, i_10_169_2703_0,
    i_10_169_2704_0, i_10_169_2706_0, i_10_169_2715_0, i_10_169_2718_0,
    i_10_169_2884_0, i_10_169_2885_0, i_10_169_2980_0, i_10_169_2986_0,
    i_10_169_3034_0, i_10_169_3036_0, i_10_169_3087_0, i_10_169_3093_0,
    i_10_169_3094_0, i_10_169_3154_0, i_10_169_3155_0, i_10_169_3165_0,
    i_10_169_3196_0, i_10_169_3198_0, i_10_169_3199_0, i_10_169_3200_0,
    i_10_169_3321_0, i_10_169_3322_0, i_10_169_3384_0, i_10_169_3405_0,
    i_10_169_3406_0, i_10_169_3407_0, i_10_169_3408_0, i_10_169_3409_0,
    i_10_169_3610_0, i_10_169_3613_0, i_10_169_3614_0, i_10_169_3615_0,
    i_10_169_3650_0, i_10_169_3702_0, i_10_169_3780_0, i_10_169_3782_0,
    i_10_169_3788_0, i_10_169_3837_0, i_10_169_3846_0, i_10_169_3856_0,
    i_10_169_3859_0, i_10_169_3982_0, i_10_169_4115_0, i_10_169_4273_0,
    i_10_169_4288_0, i_10_169_4564_0, i_10_169_4565_0, i_10_169_4568_0;
  output o_10_169_0_0;
  assign o_10_169_0_0 = ~((~i_10_169_438_0 & ((~i_10_169_433_0 & ((~i_10_169_440_0 & ~i_10_169_1647_0 & i_10_169_1823_0 & ~i_10_169_2884_0 & ~i_10_169_3384_0 & ~i_10_169_3408_0 & ~i_10_169_3982_0 & ~i_10_169_4115_0) | (~i_10_169_439_0 & ~i_10_169_1579_0 & ~i_10_169_2715_0 & ~i_10_169_3034_0 & ~i_10_169_3198_0 & ~i_10_169_3200_0 & ~i_10_169_3780_0 & ~i_10_169_4568_0))) | (~i_10_169_439_0 & ((~i_10_169_435_0 & ((~i_10_169_429_0 & ~i_10_169_1579_0 & ~i_10_169_1819_0 & ~i_10_169_1823_0 & ~i_10_169_2885_0 & ~i_10_169_3034_0 & ~i_10_169_3165_0 & ~i_10_169_3199_0) | (~i_10_169_423_0 & ~i_10_169_436_0 & ~i_10_169_748_0 & ~i_10_169_2629_0 & ~i_10_169_2715_0 & ~i_10_169_2884_0 & ~i_10_169_3087_0 & ~i_10_169_3196_0 & ~i_10_169_3405_0 & ~i_10_169_3407_0))) | (~i_10_169_440_0 & ~i_10_169_1305_0 & ~i_10_169_1308_0 & ~i_10_169_2453_0 & ~i_10_169_3199_0 & ~i_10_169_3408_0 & ~i_10_169_3614_0) | (i_10_169_282_0 & ~i_10_169_1309_0 & ~i_10_169_3409_0 & ~i_10_169_3780_0 & ~i_10_169_4115_0))) | (~i_10_169_436_0 & i_10_169_2351_0 & ~i_10_169_3780_0 & ~i_10_169_3982_0))) | (~i_10_169_439_0 & ((~i_10_169_423_0 & ((~i_10_169_441_0 & ~i_10_169_748_0 & i_10_169_2353_0 & ~i_10_169_2453_0 & ~i_10_169_2980_0 & ~i_10_169_3200_0) | (i_10_169_428_0 & ~i_10_169_1823_0 & ~i_10_169_3196_0 & i_10_169_3614_0))) | (~i_10_169_751_0 & ((~i_10_169_440_0 & i_10_169_1579_0 & i_10_169_2354_0 & ~i_10_169_3093_0) | (~i_10_169_2986_0 & ~i_10_169_3087_0 & ~i_10_169_3196_0 & ~i_10_169_3198_0 & ~i_10_169_3859_0 & ~i_10_169_3982_0 & i_10_169_4115_0))) | (~i_10_169_1305_0 & ((i_10_169_1249_0 & ~i_10_169_2715_0 & ~i_10_169_3034_0 & ~i_10_169_3615_0) | (~i_10_169_1647_0 & ~i_10_169_2634_0 & ~i_10_169_2986_0 & ~i_10_169_3165_0 & ~i_10_169_3196_0 & ~i_10_169_3198_0 & ~i_10_169_3406_0 & ~i_10_169_3856_0))) | (~i_10_169_3405_0 & ((~i_10_169_430_0 & ~i_10_169_435_0 & ~i_10_169_2885_0 & ~i_10_169_3087_0 & ~i_10_169_3610_0 & ~i_10_169_3780_0 & ~i_10_169_3782_0 & ~i_10_169_3837_0) | (~i_10_169_2884_0 & i_10_169_4568_0))) | (~i_10_169_429_0 & ~i_10_169_436_0 & ~i_10_169_1647_0 & ~i_10_169_1683_0 & ~i_10_169_3613_0 & ~i_10_169_3614_0 & i_10_169_3788_0))) | (~i_10_169_430_0 & ~i_10_169_465_0 & ((~i_10_169_178_0 & ~i_10_169_441_0 & ~i_10_169_1687_0 & ~i_10_169_2634_0 & ~i_10_169_2884_0 & ~i_10_169_2986_0 & ~i_10_169_3087_0 & ~i_10_169_3610_0 & ~i_10_169_3650_0 & ~i_10_169_3837_0) | (~i_10_169_440_0 & ~i_10_169_751_0 & ~i_10_169_793_0 & ~i_10_169_1237_0 & ~i_10_169_1306_0 & ~i_10_169_2885_0 & ~i_10_169_3165_0 & ~i_10_169_3196_0 & ~i_10_169_3615_0 & ~i_10_169_3982_0))) | (~i_10_169_435_0 & ((~i_10_169_440_0 & ~i_10_169_1308_0 & ~i_10_169_1647_0 & i_10_169_2350_0 & ~i_10_169_2980_0 & ~i_10_169_3409_0) | (~i_10_169_436_0 & ~i_10_169_748_0 & ~i_10_169_1305_0 & i_10_169_1819_0 & ~i_10_169_2884_0 & ~i_10_169_3614_0 & ~i_10_169_3782_0))) | (~i_10_169_440_0 & ~i_10_169_3087_0 & ((i_10_169_793_0 & ~i_10_169_3196_0 & ~i_10_169_3610_0 & ~i_10_169_3782_0) | (i_10_169_279_0 & ~i_10_169_429_0 & ~i_10_169_1309_0 & ~i_10_169_2885_0 & i_10_169_4288_0))) | (~i_10_169_2634_0 & ((~i_10_169_279_0 & ~i_10_169_447_0 & ~i_10_169_1308_0 & ~i_10_169_1820_0 & ~i_10_169_3982_0 & i_10_169_4115_0 & ~i_10_169_3610_0 & ~i_10_169_3613_0) | (i_10_169_1309_0 & i_10_169_4564_0))) | (i_10_169_4115_0 & ((i_10_169_2453_0 & ~i_10_169_2629_0 & ~i_10_169_3610_0 & ~i_10_169_3846_0) | (i_10_169_4288_0 & i_10_169_4565_0))) | (~i_10_169_428_0 & ~i_10_169_748_0 & i_10_169_1820_0 & ~i_10_169_2353_0 & ~i_10_169_2703_0 & ~i_10_169_2885_0 & ~i_10_169_3036_0 & ~i_10_169_3094_0 & ~i_10_169_3782_0) | (i_10_169_172_0 & ~i_10_169_3200_0 & ~i_10_169_3405_0 & i_10_169_4568_0));
endmodule



// Benchmark "kernel_10_170" written by ABC on Sun Jul 19 10:23:56 2020

module kernel_10_170 ( 
    i_10_170_51_0, i_10_170_83_0, i_10_170_223_0, i_10_170_280_0,
    i_10_170_281_0, i_10_170_282_0, i_10_170_286_0, i_10_170_289_0,
    i_10_170_394_0, i_10_170_430_0, i_10_170_512_0, i_10_170_516_0,
    i_10_170_743_0, i_10_170_751_0, i_10_170_823_0, i_10_170_824_0,
    i_10_170_852_0, i_10_170_896_0, i_10_170_1003_0, i_10_170_1030_0,
    i_10_170_1031_0, i_10_170_1112_0, i_10_170_1219_0, i_10_170_1300_0,
    i_10_170_1306_0, i_10_170_1309_0, i_10_170_1345_0, i_10_170_1346_0,
    i_10_170_1349_0, i_10_170_1357_0, i_10_170_1435_0, i_10_170_1439_0,
    i_10_170_1445_0, i_10_170_1493_0, i_10_170_1544_0, i_10_170_1556_0,
    i_10_170_1607_0, i_10_170_1652_0, i_10_170_1654_0, i_10_170_1803_0,
    i_10_170_1804_0, i_10_170_1820_0, i_10_170_1915_0, i_10_170_1996_0,
    i_10_170_1997_0, i_10_170_2184_0, i_10_170_2185_0, i_10_170_2291_0,
    i_10_170_2380_0, i_10_170_2444_0, i_10_170_2566_0, i_10_170_2567_0,
    i_10_170_2570_0, i_10_170_2604_0, i_10_170_2644_0, i_10_170_2674_0,
    i_10_170_2712_0, i_10_170_2713_0, i_10_170_2714_0, i_10_170_2730_0,
    i_10_170_2734_0, i_10_170_2742_0, i_10_170_2827_0, i_10_170_2867_0,
    i_10_170_2882_0, i_10_170_2965_0, i_10_170_2990_0, i_10_170_3046_0,
    i_10_170_3091_0, i_10_170_3162_0, i_10_170_3197_0, i_10_170_3391_0,
    i_10_170_3505_0, i_10_170_3558_0, i_10_170_3609_0, i_10_170_3653_0,
    i_10_170_3797_0, i_10_170_3841_0, i_10_170_3842_0, i_10_170_3859_0,
    i_10_170_3892_0, i_10_170_3893_0, i_10_170_3979_0, i_10_170_4026_0,
    i_10_170_4027_0, i_10_170_4028_0, i_10_170_4030_0, i_10_170_4129_0,
    i_10_170_4153_0, i_10_170_4154_0, i_10_170_4175_0, i_10_170_4193_0,
    i_10_170_4208_0, i_10_170_4237_0, i_10_170_4271_0, i_10_170_4278_0,
    i_10_170_4400_0, i_10_170_4455_0, i_10_170_4535_0, i_10_170_4553_0,
    o_10_170_0_0  );
  input  i_10_170_51_0, i_10_170_83_0, i_10_170_223_0, i_10_170_280_0,
    i_10_170_281_0, i_10_170_282_0, i_10_170_286_0, i_10_170_289_0,
    i_10_170_394_0, i_10_170_430_0, i_10_170_512_0, i_10_170_516_0,
    i_10_170_743_0, i_10_170_751_0, i_10_170_823_0, i_10_170_824_0,
    i_10_170_852_0, i_10_170_896_0, i_10_170_1003_0, i_10_170_1030_0,
    i_10_170_1031_0, i_10_170_1112_0, i_10_170_1219_0, i_10_170_1300_0,
    i_10_170_1306_0, i_10_170_1309_0, i_10_170_1345_0, i_10_170_1346_0,
    i_10_170_1349_0, i_10_170_1357_0, i_10_170_1435_0, i_10_170_1439_0,
    i_10_170_1445_0, i_10_170_1493_0, i_10_170_1544_0, i_10_170_1556_0,
    i_10_170_1607_0, i_10_170_1652_0, i_10_170_1654_0, i_10_170_1803_0,
    i_10_170_1804_0, i_10_170_1820_0, i_10_170_1915_0, i_10_170_1996_0,
    i_10_170_1997_0, i_10_170_2184_0, i_10_170_2185_0, i_10_170_2291_0,
    i_10_170_2380_0, i_10_170_2444_0, i_10_170_2566_0, i_10_170_2567_0,
    i_10_170_2570_0, i_10_170_2604_0, i_10_170_2644_0, i_10_170_2674_0,
    i_10_170_2712_0, i_10_170_2713_0, i_10_170_2714_0, i_10_170_2730_0,
    i_10_170_2734_0, i_10_170_2742_0, i_10_170_2827_0, i_10_170_2867_0,
    i_10_170_2882_0, i_10_170_2965_0, i_10_170_2990_0, i_10_170_3046_0,
    i_10_170_3091_0, i_10_170_3162_0, i_10_170_3197_0, i_10_170_3391_0,
    i_10_170_3505_0, i_10_170_3558_0, i_10_170_3609_0, i_10_170_3653_0,
    i_10_170_3797_0, i_10_170_3841_0, i_10_170_3842_0, i_10_170_3859_0,
    i_10_170_3892_0, i_10_170_3893_0, i_10_170_3979_0, i_10_170_4026_0,
    i_10_170_4027_0, i_10_170_4028_0, i_10_170_4030_0, i_10_170_4129_0,
    i_10_170_4153_0, i_10_170_4154_0, i_10_170_4175_0, i_10_170_4193_0,
    i_10_170_4208_0, i_10_170_4237_0, i_10_170_4271_0, i_10_170_4278_0,
    i_10_170_4400_0, i_10_170_4455_0, i_10_170_4535_0, i_10_170_4553_0;
  output o_10_170_0_0;
  assign o_10_170_0_0 = 0;
endmodule



// Benchmark "kernel_10_171" written by ABC on Sun Jul 19 10:23:57 2020

module kernel_10_171 ( 
    i_10_171_177_0, i_10_171_184_0, i_10_171_220_0, i_10_171_223_0,
    i_10_171_291_0, i_10_171_321_0, i_10_171_329_0, i_10_171_394_0,
    i_10_171_411_0, i_10_171_426_0, i_10_171_427_0, i_10_171_430_0,
    i_10_171_444_0, i_10_171_448_0, i_10_171_467_0, i_10_171_511_0,
    i_10_171_693_0, i_10_171_694_0, i_10_171_730_0, i_10_171_733_0,
    i_10_171_796_0, i_10_171_797_0, i_10_171_800_0, i_10_171_961_0,
    i_10_171_970_0, i_10_171_999_0, i_10_171_1233_0, i_10_171_1234_0,
    i_10_171_1235_0, i_10_171_1238_0, i_10_171_1243_0, i_10_171_1363_0,
    i_10_171_1548_0, i_10_171_1549_0, i_10_171_1552_0, i_10_171_1578_0,
    i_10_171_1617_0, i_10_171_1734_0, i_10_171_1821_0, i_10_171_1823_0,
    i_10_171_1909_0, i_10_171_1912_0, i_10_171_1990_0, i_10_171_2358_0,
    i_10_171_2361_0, i_10_171_2362_0, i_10_171_2364_0, i_10_171_2365_0,
    i_10_171_2376_0, i_10_171_2383_0, i_10_171_2448_0, i_10_171_2716_0,
    i_10_171_2719_0, i_10_171_2823_0, i_10_171_2827_0, i_10_171_2829_0,
    i_10_171_2883_0, i_10_171_2884_0, i_10_171_2917_0, i_10_171_2953_0,
    i_10_171_2980_0, i_10_171_2982_0, i_10_171_2985_0, i_10_171_3034_0,
    i_10_171_3036_0, i_10_171_3038_0, i_10_171_3153_0, i_10_171_3154_0,
    i_10_171_3200_0, i_10_171_3273_0, i_10_171_3276_0, i_10_171_3279_0,
    i_10_171_3281_0, i_10_171_3282_0, i_10_171_3283_0, i_10_171_3324_0,
    i_10_171_3326_0, i_10_171_3784_0, i_10_171_3850_0, i_10_171_3852_0,
    i_10_171_3853_0, i_10_171_3855_0, i_10_171_3858_0, i_10_171_3859_0,
    i_10_171_3860_0, i_10_171_3888_0, i_10_171_3895_0, i_10_171_3912_0,
    i_10_171_3978_0, i_10_171_3979_0, i_10_171_3981_0, i_10_171_3982_0,
    i_10_171_3984_0, i_10_171_3985_0, i_10_171_3990_0, i_10_171_4113_0,
    i_10_171_4121_0, i_10_171_4281_0, i_10_171_4292_0, i_10_171_4570_0,
    o_10_171_0_0  );
  input  i_10_171_177_0, i_10_171_184_0, i_10_171_220_0, i_10_171_223_0,
    i_10_171_291_0, i_10_171_321_0, i_10_171_329_0, i_10_171_394_0,
    i_10_171_411_0, i_10_171_426_0, i_10_171_427_0, i_10_171_430_0,
    i_10_171_444_0, i_10_171_448_0, i_10_171_467_0, i_10_171_511_0,
    i_10_171_693_0, i_10_171_694_0, i_10_171_730_0, i_10_171_733_0,
    i_10_171_796_0, i_10_171_797_0, i_10_171_800_0, i_10_171_961_0,
    i_10_171_970_0, i_10_171_999_0, i_10_171_1233_0, i_10_171_1234_0,
    i_10_171_1235_0, i_10_171_1238_0, i_10_171_1243_0, i_10_171_1363_0,
    i_10_171_1548_0, i_10_171_1549_0, i_10_171_1552_0, i_10_171_1578_0,
    i_10_171_1617_0, i_10_171_1734_0, i_10_171_1821_0, i_10_171_1823_0,
    i_10_171_1909_0, i_10_171_1912_0, i_10_171_1990_0, i_10_171_2358_0,
    i_10_171_2361_0, i_10_171_2362_0, i_10_171_2364_0, i_10_171_2365_0,
    i_10_171_2376_0, i_10_171_2383_0, i_10_171_2448_0, i_10_171_2716_0,
    i_10_171_2719_0, i_10_171_2823_0, i_10_171_2827_0, i_10_171_2829_0,
    i_10_171_2883_0, i_10_171_2884_0, i_10_171_2917_0, i_10_171_2953_0,
    i_10_171_2980_0, i_10_171_2982_0, i_10_171_2985_0, i_10_171_3034_0,
    i_10_171_3036_0, i_10_171_3038_0, i_10_171_3153_0, i_10_171_3154_0,
    i_10_171_3200_0, i_10_171_3273_0, i_10_171_3276_0, i_10_171_3279_0,
    i_10_171_3281_0, i_10_171_3282_0, i_10_171_3283_0, i_10_171_3324_0,
    i_10_171_3326_0, i_10_171_3784_0, i_10_171_3850_0, i_10_171_3852_0,
    i_10_171_3853_0, i_10_171_3855_0, i_10_171_3858_0, i_10_171_3859_0,
    i_10_171_3860_0, i_10_171_3888_0, i_10_171_3895_0, i_10_171_3912_0,
    i_10_171_3978_0, i_10_171_3979_0, i_10_171_3981_0, i_10_171_3982_0,
    i_10_171_3984_0, i_10_171_3985_0, i_10_171_3990_0, i_10_171_4113_0,
    i_10_171_4121_0, i_10_171_4281_0, i_10_171_4292_0, i_10_171_4570_0;
  output o_10_171_0_0;
  assign o_10_171_0_0 = ~((~i_10_171_321_0 & ((~i_10_171_329_0 & ~i_10_171_394_0 & ~i_10_171_694_0 & ~i_10_171_1548_0 & ~i_10_171_1617_0 & ~i_10_171_1734_0 & ~i_10_171_2376_0 & ~i_10_171_2980_0 & ~i_10_171_2982_0 & ~i_10_171_2985_0) | (~i_10_171_796_0 & ~i_10_171_999_0 & ~i_10_171_1552_0 & i_10_171_3855_0))) | (~i_10_171_970_0 & ((~i_10_171_427_0 & ((~i_10_171_329_0 & ((~i_10_171_444_0 & ~i_10_171_467_0 & ~i_10_171_693_0 & ~i_10_171_1990_0 & ~i_10_171_2823_0 & ~i_10_171_2883_0 & ~i_10_171_3276_0 & ~i_10_171_4281_0) | (~i_10_171_426_0 & ~i_10_171_1578_0 & ~i_10_171_1912_0 & ~i_10_171_2376_0 & ~i_10_171_2827_0 & ~i_10_171_3888_0 & ~i_10_171_3912_0 & ~i_10_171_3981_0 & ~i_10_171_3990_0 & ~i_10_171_4570_0))) | (~i_10_171_426_0 & ~i_10_171_430_0 & ~i_10_171_999_0 & ~i_10_171_2719_0 & ~i_10_171_2823_0 & ~i_10_171_3276_0 & ~i_10_171_3850_0 & ~i_10_171_3888_0 & ~i_10_171_3981_0 & ~i_10_171_3982_0 & ~i_10_171_3985_0))) | (~i_10_171_2985_0 & ((~i_10_171_1548_0 & ~i_10_171_1552_0 & ~i_10_171_1734_0 & ~i_10_171_2883_0 & ~i_10_171_2982_0 & ~i_10_171_3912_0 & ~i_10_171_3981_0) | (~i_10_171_693_0 & ~i_10_171_2980_0 & ~i_10_171_3283_0 & ~i_10_171_3895_0 & ~i_10_171_3978_0 & ~i_10_171_3982_0))))) | (~i_10_171_3985_0 & ((~i_10_171_430_0 & ((~i_10_171_467_0 & ~i_10_171_961_0 & ~i_10_171_1549_0 & ~i_10_171_2884_0 & ~i_10_171_2985_0 & ~i_10_171_3282_0 & ~i_10_171_3982_0) | (~i_10_171_797_0 & ~i_10_171_999_0 & ~i_10_171_3912_0 & ~i_10_171_3978_0 & ~i_10_171_3990_0))) | (~i_10_171_1549_0 & ~i_10_171_2823_0 & i_10_171_2982_0 & ~i_10_171_3034_0 & ~i_10_171_3850_0 & ~i_10_171_3981_0))) | (~i_10_171_3912_0 & ((~i_10_171_1552_0 & ~i_10_171_3034_0 & ((~i_10_171_223_0 & ~i_10_171_693_0 & ~i_10_171_1734_0 & ~i_10_171_2716_0 & ~i_10_171_3888_0 & ~i_10_171_3895_0 & ~i_10_171_3979_0 & ~i_10_171_3984_0) | (~i_10_171_426_0 & ~i_10_171_427_0 & ~i_10_171_2448_0 & ~i_10_171_2827_0 & ~i_10_171_2884_0 & ~i_10_171_2980_0 & ~i_10_171_3982_0 & ~i_10_171_3990_0 & ~i_10_171_4292_0))) | (~i_10_171_2448_0 & ~i_10_171_2716_0 & ~i_10_171_2827_0 & ~i_10_171_2980_0 & ~i_10_171_3273_0 & ~i_10_171_3281_0 & ~i_10_171_3282_0 & ~i_10_171_3858_0 & ~i_10_171_3888_0 & ~i_10_171_3979_0 & ~i_10_171_4292_0))) | (~i_10_171_2883_0 & ((~i_10_171_2448_0 & ((i_10_171_467_0 & ~i_10_171_1821_0 & ~i_10_171_2383_0 & ~i_10_171_2716_0 & ~i_10_171_3282_0 & ~i_10_171_3888_0 & ~i_10_171_4281_0) | (~i_10_171_448_0 & ~i_10_171_1734_0 & ~i_10_171_3038_0 & ~i_10_171_3279_0 & i_10_171_4292_0 & ~i_10_171_4570_0))) | (~i_10_171_2823_0 & i_10_171_3859_0 & ~i_10_171_4281_0) | (i_10_171_2719_0 & i_10_171_3858_0 & ~i_10_171_3990_0))) | (~i_10_171_1734_0 & ((~i_10_171_394_0 & ~i_10_171_694_0 & i_10_171_1235_0 & ~i_10_171_2985_0) | (~i_10_171_444_0 & ~i_10_171_796_0 & ~i_10_171_2719_0 & ~i_10_171_3850_0 & ~i_10_171_3981_0 & ~i_10_171_3990_0 & ~i_10_171_4281_0))) | (~i_10_171_3984_0 & ((i_10_171_1233_0 & i_10_171_1238_0 & ~i_10_171_1548_0 & ~i_10_171_2376_0 & i_10_171_3852_0) | (~i_10_171_3850_0 & i_10_171_3859_0 & i_10_171_3888_0 & ~i_10_171_3990_0))));
endmodule



// Benchmark "kernel_10_172" written by ABC on Sun Jul 19 10:23:58 2020

module kernel_10_172 ( 
    i_10_172_70_0, i_10_172_71_0, i_10_172_157_0, i_10_172_185_0,
    i_10_172_283_0, i_10_172_285_0, i_10_172_286_0, i_10_172_316_0,
    i_10_172_434_0, i_10_172_445_0, i_10_172_447_0, i_10_172_562_0,
    i_10_172_563_0, i_10_172_953_0, i_10_172_1045_0, i_10_172_1080_0,
    i_10_172_1081_0, i_10_172_1160_0, i_10_172_1236_0, i_10_172_1237_0,
    i_10_172_1238_0, i_10_172_1267_0, i_10_172_1363_0, i_10_172_1544_0,
    i_10_172_1555_0, i_10_172_1577_0, i_10_172_1614_0, i_10_172_1627_0,
    i_10_172_1642_0, i_10_172_1654_0, i_10_172_1772_0, i_10_172_1922_0,
    i_10_172_2017_0, i_10_172_2159_0, i_10_172_2203_0, i_10_172_2240_0,
    i_10_172_2354_0, i_10_172_2356_0, i_10_172_2357_0, i_10_172_2361_0,
    i_10_172_2364_0, i_10_172_2365_0, i_10_172_2407_0, i_10_172_2436_0,
    i_10_172_2451_0, i_10_172_2452_0, i_10_172_2458_0, i_10_172_2461_0,
    i_10_172_2463_0, i_10_172_2464_0, i_10_172_2516_0, i_10_172_2518_0,
    i_10_172_2564_0, i_10_172_2570_0, i_10_172_2573_0, i_10_172_2602_0,
    i_10_172_2607_0, i_10_172_2633_0, i_10_172_2656_0, i_10_172_2658_0,
    i_10_172_2717_0, i_10_172_2826_0, i_10_172_2829_0, i_10_172_2830_0,
    i_10_172_2831_0, i_10_172_2834_0, i_10_172_2885_0, i_10_172_3036_0,
    i_10_172_3046_0, i_10_172_3074_0, i_10_172_3160_0, i_10_172_3199_0,
    i_10_172_3392_0, i_10_172_3519_0, i_10_172_3545_0, i_10_172_3563_0,
    i_10_172_3585_0, i_10_172_3586_0, i_10_172_3613_0, i_10_172_3721_0,
    i_10_172_3722_0, i_10_172_3788_0, i_10_172_3842_0, i_10_172_3850_0,
    i_10_172_3856_0, i_10_172_3857_0, i_10_172_3907_0, i_10_172_3923_0,
    i_10_172_3988_0, i_10_172_4120_0, i_10_172_4122_0, i_10_172_4123_0,
    i_10_172_4168_0, i_10_172_4169_0, i_10_172_4282_0, i_10_172_4283_0,
    i_10_172_4310_0, i_10_172_4435_0, i_10_172_4521_0, i_10_172_4565_0,
    o_10_172_0_0  );
  input  i_10_172_70_0, i_10_172_71_0, i_10_172_157_0, i_10_172_185_0,
    i_10_172_283_0, i_10_172_285_0, i_10_172_286_0, i_10_172_316_0,
    i_10_172_434_0, i_10_172_445_0, i_10_172_447_0, i_10_172_562_0,
    i_10_172_563_0, i_10_172_953_0, i_10_172_1045_0, i_10_172_1080_0,
    i_10_172_1081_0, i_10_172_1160_0, i_10_172_1236_0, i_10_172_1237_0,
    i_10_172_1238_0, i_10_172_1267_0, i_10_172_1363_0, i_10_172_1544_0,
    i_10_172_1555_0, i_10_172_1577_0, i_10_172_1614_0, i_10_172_1627_0,
    i_10_172_1642_0, i_10_172_1654_0, i_10_172_1772_0, i_10_172_1922_0,
    i_10_172_2017_0, i_10_172_2159_0, i_10_172_2203_0, i_10_172_2240_0,
    i_10_172_2354_0, i_10_172_2356_0, i_10_172_2357_0, i_10_172_2361_0,
    i_10_172_2364_0, i_10_172_2365_0, i_10_172_2407_0, i_10_172_2436_0,
    i_10_172_2451_0, i_10_172_2452_0, i_10_172_2458_0, i_10_172_2461_0,
    i_10_172_2463_0, i_10_172_2464_0, i_10_172_2516_0, i_10_172_2518_0,
    i_10_172_2564_0, i_10_172_2570_0, i_10_172_2573_0, i_10_172_2602_0,
    i_10_172_2607_0, i_10_172_2633_0, i_10_172_2656_0, i_10_172_2658_0,
    i_10_172_2717_0, i_10_172_2826_0, i_10_172_2829_0, i_10_172_2830_0,
    i_10_172_2831_0, i_10_172_2834_0, i_10_172_2885_0, i_10_172_3036_0,
    i_10_172_3046_0, i_10_172_3074_0, i_10_172_3160_0, i_10_172_3199_0,
    i_10_172_3392_0, i_10_172_3519_0, i_10_172_3545_0, i_10_172_3563_0,
    i_10_172_3585_0, i_10_172_3586_0, i_10_172_3613_0, i_10_172_3721_0,
    i_10_172_3722_0, i_10_172_3788_0, i_10_172_3842_0, i_10_172_3850_0,
    i_10_172_3856_0, i_10_172_3857_0, i_10_172_3907_0, i_10_172_3923_0,
    i_10_172_3988_0, i_10_172_4120_0, i_10_172_4122_0, i_10_172_4123_0,
    i_10_172_4168_0, i_10_172_4169_0, i_10_172_4282_0, i_10_172_4283_0,
    i_10_172_4310_0, i_10_172_4435_0, i_10_172_4521_0, i_10_172_4565_0;
  output o_10_172_0_0;
  assign o_10_172_0_0 = 0;
endmodule



// Benchmark "kernel_10_173" written by ABC on Sun Jul 19 10:23:58 2020

module kernel_10_173 ( 
    i_10_173_133_0, i_10_173_221_0, i_10_173_257_0, i_10_173_263_0,
    i_10_173_269_0, i_10_173_282_0, i_10_173_405_0, i_10_173_409_0,
    i_10_173_442_0, i_10_173_566_0, i_10_173_626_0, i_10_173_793_0,
    i_10_173_1003_0, i_10_173_1004_0, i_10_173_1007_0, i_10_173_1016_0,
    i_10_173_1052_0, i_10_173_1106_0, i_10_173_1213_0, i_10_173_1234_0,
    i_10_173_1235_0, i_10_173_1237_0, i_10_173_1238_0, i_10_173_1267_0,
    i_10_173_1300_0, i_10_173_1303_0, i_10_173_1304_0, i_10_173_1305_0,
    i_10_173_1345_0, i_10_173_1540_0, i_10_173_1628_0, i_10_173_1683_0,
    i_10_173_1685_0, i_10_173_1686_0, i_10_173_1728_0, i_10_173_1729_0,
    i_10_173_1769_0, i_10_173_1771_0, i_10_173_1804_0, i_10_173_1823_0,
    i_10_173_1922_0, i_10_173_2006_0, i_10_173_2200_0, i_10_173_2362_0,
    i_10_173_2365_0, i_10_173_2436_0, i_10_173_2449_0, i_10_173_2453_0,
    i_10_173_2461_0, i_10_173_2563_0, i_10_173_2564_0, i_10_173_2607_0,
    i_10_173_2608_0, i_10_173_2631_0, i_10_173_2636_0, i_10_173_2658_0,
    i_10_173_2660_0, i_10_173_2711_0, i_10_173_2716_0, i_10_173_2734_0,
    i_10_173_2759_0, i_10_173_2762_0, i_10_173_2824_0, i_10_173_2831_0,
    i_10_173_2845_0, i_10_173_2870_0, i_10_173_2962_0, i_10_173_2963_0,
    i_10_173_3033_0, i_10_173_3036_0, i_10_173_3185_0, i_10_173_3200_0,
    i_10_173_3317_0, i_10_173_3389_0, i_10_173_3473_0, i_10_173_3526_0,
    i_10_173_3538_0, i_10_173_3540_0, i_10_173_3541_0, i_10_173_3542_0,
    i_10_173_3614_0, i_10_173_3702_0, i_10_173_3838_0, i_10_173_3839_0,
    i_10_173_3840_0, i_10_173_3843_0, i_10_173_3844_0, i_10_173_3858_0,
    i_10_173_3913_0, i_10_173_3986_0, i_10_173_4118_0, i_10_173_4151_0,
    i_10_173_4168_0, i_10_173_4169_0, i_10_173_4266_0, i_10_173_4274_0,
    i_10_173_4287_0, i_10_173_4428_0, i_10_173_4553_0, i_10_173_4565_0,
    o_10_173_0_0  );
  input  i_10_173_133_0, i_10_173_221_0, i_10_173_257_0, i_10_173_263_0,
    i_10_173_269_0, i_10_173_282_0, i_10_173_405_0, i_10_173_409_0,
    i_10_173_442_0, i_10_173_566_0, i_10_173_626_0, i_10_173_793_0,
    i_10_173_1003_0, i_10_173_1004_0, i_10_173_1007_0, i_10_173_1016_0,
    i_10_173_1052_0, i_10_173_1106_0, i_10_173_1213_0, i_10_173_1234_0,
    i_10_173_1235_0, i_10_173_1237_0, i_10_173_1238_0, i_10_173_1267_0,
    i_10_173_1300_0, i_10_173_1303_0, i_10_173_1304_0, i_10_173_1305_0,
    i_10_173_1345_0, i_10_173_1540_0, i_10_173_1628_0, i_10_173_1683_0,
    i_10_173_1685_0, i_10_173_1686_0, i_10_173_1728_0, i_10_173_1729_0,
    i_10_173_1769_0, i_10_173_1771_0, i_10_173_1804_0, i_10_173_1823_0,
    i_10_173_1922_0, i_10_173_2006_0, i_10_173_2200_0, i_10_173_2362_0,
    i_10_173_2365_0, i_10_173_2436_0, i_10_173_2449_0, i_10_173_2453_0,
    i_10_173_2461_0, i_10_173_2563_0, i_10_173_2564_0, i_10_173_2607_0,
    i_10_173_2608_0, i_10_173_2631_0, i_10_173_2636_0, i_10_173_2658_0,
    i_10_173_2660_0, i_10_173_2711_0, i_10_173_2716_0, i_10_173_2734_0,
    i_10_173_2759_0, i_10_173_2762_0, i_10_173_2824_0, i_10_173_2831_0,
    i_10_173_2845_0, i_10_173_2870_0, i_10_173_2962_0, i_10_173_2963_0,
    i_10_173_3033_0, i_10_173_3036_0, i_10_173_3185_0, i_10_173_3200_0,
    i_10_173_3317_0, i_10_173_3389_0, i_10_173_3473_0, i_10_173_3526_0,
    i_10_173_3538_0, i_10_173_3540_0, i_10_173_3541_0, i_10_173_3542_0,
    i_10_173_3614_0, i_10_173_3702_0, i_10_173_3838_0, i_10_173_3839_0,
    i_10_173_3840_0, i_10_173_3843_0, i_10_173_3844_0, i_10_173_3858_0,
    i_10_173_3913_0, i_10_173_3986_0, i_10_173_4118_0, i_10_173_4151_0,
    i_10_173_4168_0, i_10_173_4169_0, i_10_173_4266_0, i_10_173_4274_0,
    i_10_173_4287_0, i_10_173_4428_0, i_10_173_4553_0, i_10_173_4565_0;
  output o_10_173_0_0;
  assign o_10_173_0_0 = 0;
endmodule



// Benchmark "kernel_10_174" written by ABC on Sun Jul 19 10:23:59 2020

module kernel_10_174 ( 
    i_10_174_89_0, i_10_174_177_0, i_10_174_179_0, i_10_174_267_0,
    i_10_174_283_0, i_10_174_317_0, i_10_174_389_0, i_10_174_390_0,
    i_10_174_407_0, i_10_174_441_0, i_10_174_460_0, i_10_174_713_0,
    i_10_174_795_0, i_10_174_993_0, i_10_174_1003_0, i_10_174_1121_0,
    i_10_174_1260_0, i_10_174_1360_0, i_10_174_1431_0, i_10_174_1540_0,
    i_10_174_1552_0, i_10_174_1683_0, i_10_174_1684_0, i_10_174_1685_0,
    i_10_174_1687_0, i_10_174_1688_0, i_10_174_1740_0, i_10_174_1771_0,
    i_10_174_1800_0, i_10_174_1801_0, i_10_174_1803_0, i_10_174_1804_0,
    i_10_174_1819_0, i_10_174_1821_0, i_10_174_1981_0, i_10_174_2000_0,
    i_10_174_2365_0, i_10_174_2449_0, i_10_174_2452_0, i_10_174_2539_0,
    i_10_174_2543_0, i_10_174_2565_0, i_10_174_2566_0, i_10_174_2608_0,
    i_10_174_2629_0, i_10_174_2631_0, i_10_174_2657_0, i_10_174_2673_0,
    i_10_174_2700_0, i_10_174_2702_0, i_10_174_2703_0, i_10_174_2704_0,
    i_10_174_2705_0, i_10_174_2709_0, i_10_174_2710_0, i_10_174_2713_0,
    i_10_174_2728_0, i_10_174_2729_0, i_10_174_2737_0, i_10_174_2782_0,
    i_10_174_2785_0, i_10_174_2786_0, i_10_174_2821_0, i_10_174_2828_0,
    i_10_174_2829_0, i_10_174_3040_0, i_10_174_3043_0, i_10_174_3073_0,
    i_10_174_3091_0, i_10_174_3114_0, i_10_174_3166_0, i_10_174_3233_0,
    i_10_174_3281_0, i_10_174_3385_0, i_10_174_3386_0, i_10_174_3388_0,
    i_10_174_3406_0, i_10_174_3407_0, i_10_174_3410_0, i_10_174_3542_0,
    i_10_174_3584_0, i_10_174_3645_0, i_10_174_3647_0, i_10_174_3648_0,
    i_10_174_3649_0, i_10_174_3650_0, i_10_174_3652_0, i_10_174_3811_0,
    i_10_174_3834_0, i_10_174_3837_0, i_10_174_3855_0, i_10_174_3902_0,
    i_10_174_3904_0, i_10_174_3906_0, i_10_174_4025_0, i_10_174_4115_0,
    i_10_174_4214_0, i_10_174_4290_0, i_10_174_4291_0, i_10_174_4568_0,
    o_10_174_0_0  );
  input  i_10_174_89_0, i_10_174_177_0, i_10_174_179_0, i_10_174_267_0,
    i_10_174_283_0, i_10_174_317_0, i_10_174_389_0, i_10_174_390_0,
    i_10_174_407_0, i_10_174_441_0, i_10_174_460_0, i_10_174_713_0,
    i_10_174_795_0, i_10_174_993_0, i_10_174_1003_0, i_10_174_1121_0,
    i_10_174_1260_0, i_10_174_1360_0, i_10_174_1431_0, i_10_174_1540_0,
    i_10_174_1552_0, i_10_174_1683_0, i_10_174_1684_0, i_10_174_1685_0,
    i_10_174_1687_0, i_10_174_1688_0, i_10_174_1740_0, i_10_174_1771_0,
    i_10_174_1800_0, i_10_174_1801_0, i_10_174_1803_0, i_10_174_1804_0,
    i_10_174_1819_0, i_10_174_1821_0, i_10_174_1981_0, i_10_174_2000_0,
    i_10_174_2365_0, i_10_174_2449_0, i_10_174_2452_0, i_10_174_2539_0,
    i_10_174_2543_0, i_10_174_2565_0, i_10_174_2566_0, i_10_174_2608_0,
    i_10_174_2629_0, i_10_174_2631_0, i_10_174_2657_0, i_10_174_2673_0,
    i_10_174_2700_0, i_10_174_2702_0, i_10_174_2703_0, i_10_174_2704_0,
    i_10_174_2705_0, i_10_174_2709_0, i_10_174_2710_0, i_10_174_2713_0,
    i_10_174_2728_0, i_10_174_2729_0, i_10_174_2737_0, i_10_174_2782_0,
    i_10_174_2785_0, i_10_174_2786_0, i_10_174_2821_0, i_10_174_2828_0,
    i_10_174_2829_0, i_10_174_3040_0, i_10_174_3043_0, i_10_174_3073_0,
    i_10_174_3091_0, i_10_174_3114_0, i_10_174_3166_0, i_10_174_3233_0,
    i_10_174_3281_0, i_10_174_3385_0, i_10_174_3386_0, i_10_174_3388_0,
    i_10_174_3406_0, i_10_174_3407_0, i_10_174_3410_0, i_10_174_3542_0,
    i_10_174_3584_0, i_10_174_3645_0, i_10_174_3647_0, i_10_174_3648_0,
    i_10_174_3649_0, i_10_174_3650_0, i_10_174_3652_0, i_10_174_3811_0,
    i_10_174_3834_0, i_10_174_3837_0, i_10_174_3855_0, i_10_174_3902_0,
    i_10_174_3904_0, i_10_174_3906_0, i_10_174_4025_0, i_10_174_4115_0,
    i_10_174_4214_0, i_10_174_4290_0, i_10_174_4291_0, i_10_174_4568_0;
  output o_10_174_0_0;
  assign o_10_174_0_0 = 0;
endmodule



// Benchmark "kernel_10_175" written by ABC on Sun Jul 19 10:24:00 2020

module kernel_10_175 ( 
    i_10_175_221_0, i_10_175_248_0, i_10_175_280_0, i_10_175_281_0,
    i_10_175_284_0, i_10_175_328_0, i_10_175_388_0, i_10_175_391_0,
    i_10_175_536_0, i_10_175_621_0, i_10_175_635_0, i_10_175_639_0,
    i_10_175_659_0, i_10_175_716_0, i_10_175_722_0, i_10_175_946_0,
    i_10_175_967_0, i_10_175_998_0, i_10_175_1237_0, i_10_175_1296_0,
    i_10_175_1305_0, i_10_175_1378_0, i_10_175_1453_0, i_10_175_1540_0,
    i_10_175_1544_0, i_10_175_1546_0, i_10_175_1562_0, i_10_175_1565_0,
    i_10_175_1617_0, i_10_175_1705_0, i_10_175_1809_0, i_10_175_1877_0,
    i_10_175_1917_0, i_10_175_1999_0, i_10_175_2000_0, i_10_175_2008_0,
    i_10_175_2020_0, i_10_175_2021_0, i_10_175_2039_0, i_10_175_2054_0,
    i_10_175_2057_0, i_10_175_2109_0, i_10_175_2183_0, i_10_175_2305_0,
    i_10_175_2306_0, i_10_175_2326_0, i_10_175_2452_0, i_10_175_2454_0,
    i_10_175_2455_0, i_10_175_2456_0, i_10_175_2507_0, i_10_175_2515_0,
    i_10_175_2557_0, i_10_175_2602_0, i_10_175_2605_0, i_10_175_2663_0,
    i_10_175_2674_0, i_10_175_2675_0, i_10_175_2848_0, i_10_175_2909_0,
    i_10_175_2911_0, i_10_175_2953_0, i_10_175_2961_0, i_10_175_3073_0,
    i_10_175_3106_0, i_10_175_3203_0, i_10_175_3278_0, i_10_175_3284_0,
    i_10_175_3285_0, i_10_175_3376_0, i_10_175_3386_0, i_10_175_3410_0,
    i_10_175_3431_0, i_10_175_3604_0, i_10_175_3609_0, i_10_175_3699_0,
    i_10_175_3777_0, i_10_175_3785_0, i_10_175_3788_0, i_10_175_3857_0,
    i_10_175_3902_0, i_10_175_3919_0, i_10_175_3947_0, i_10_175_3979_0,
    i_10_175_4023_0, i_10_175_4024_0, i_10_175_4025_0, i_10_175_4114_0,
    i_10_175_4117_0, i_10_175_4122_0, i_10_175_4123_0, i_10_175_4149_0,
    i_10_175_4150_0, i_10_175_4216_0, i_10_175_4220_0, i_10_175_4267_0,
    i_10_175_4275_0, i_10_175_4411_0, i_10_175_4522_0, i_10_175_4523_0,
    o_10_175_0_0  );
  input  i_10_175_221_0, i_10_175_248_0, i_10_175_280_0, i_10_175_281_0,
    i_10_175_284_0, i_10_175_328_0, i_10_175_388_0, i_10_175_391_0,
    i_10_175_536_0, i_10_175_621_0, i_10_175_635_0, i_10_175_639_0,
    i_10_175_659_0, i_10_175_716_0, i_10_175_722_0, i_10_175_946_0,
    i_10_175_967_0, i_10_175_998_0, i_10_175_1237_0, i_10_175_1296_0,
    i_10_175_1305_0, i_10_175_1378_0, i_10_175_1453_0, i_10_175_1540_0,
    i_10_175_1544_0, i_10_175_1546_0, i_10_175_1562_0, i_10_175_1565_0,
    i_10_175_1617_0, i_10_175_1705_0, i_10_175_1809_0, i_10_175_1877_0,
    i_10_175_1917_0, i_10_175_1999_0, i_10_175_2000_0, i_10_175_2008_0,
    i_10_175_2020_0, i_10_175_2021_0, i_10_175_2039_0, i_10_175_2054_0,
    i_10_175_2057_0, i_10_175_2109_0, i_10_175_2183_0, i_10_175_2305_0,
    i_10_175_2306_0, i_10_175_2326_0, i_10_175_2452_0, i_10_175_2454_0,
    i_10_175_2455_0, i_10_175_2456_0, i_10_175_2507_0, i_10_175_2515_0,
    i_10_175_2557_0, i_10_175_2602_0, i_10_175_2605_0, i_10_175_2663_0,
    i_10_175_2674_0, i_10_175_2675_0, i_10_175_2848_0, i_10_175_2909_0,
    i_10_175_2911_0, i_10_175_2953_0, i_10_175_2961_0, i_10_175_3073_0,
    i_10_175_3106_0, i_10_175_3203_0, i_10_175_3278_0, i_10_175_3284_0,
    i_10_175_3285_0, i_10_175_3376_0, i_10_175_3386_0, i_10_175_3410_0,
    i_10_175_3431_0, i_10_175_3604_0, i_10_175_3609_0, i_10_175_3699_0,
    i_10_175_3777_0, i_10_175_3785_0, i_10_175_3788_0, i_10_175_3857_0,
    i_10_175_3902_0, i_10_175_3919_0, i_10_175_3947_0, i_10_175_3979_0,
    i_10_175_4023_0, i_10_175_4024_0, i_10_175_4025_0, i_10_175_4114_0,
    i_10_175_4117_0, i_10_175_4122_0, i_10_175_4123_0, i_10_175_4149_0,
    i_10_175_4150_0, i_10_175_4216_0, i_10_175_4220_0, i_10_175_4267_0,
    i_10_175_4275_0, i_10_175_4411_0, i_10_175_4522_0, i_10_175_4523_0;
  output o_10_175_0_0;
  assign o_10_175_0_0 = 0;
endmodule



// Benchmark "kernel_10_176" written by ABC on Sun Jul 19 10:24:01 2020

module kernel_10_176 ( 
    i_10_176_34_0, i_10_176_121_0, i_10_176_122_0, i_10_176_124_0,
    i_10_176_132_0, i_10_176_133_0, i_10_176_177_0, i_10_176_178_0,
    i_10_176_183_0, i_10_176_331_0, i_10_176_367_0, i_10_176_374_0,
    i_10_176_386_0, i_10_176_429_0, i_10_176_437_0, i_10_176_439_0,
    i_10_176_440_0, i_10_176_462_0, i_10_176_599_0, i_10_176_600_0,
    i_10_176_602_0, i_10_176_634_0, i_10_176_754_0, i_10_176_755_0,
    i_10_176_906_0, i_10_176_967_0, i_10_176_971_0, i_10_176_1160_0,
    i_10_176_1240_0, i_10_176_1483_0, i_10_176_1499_0, i_10_176_1543_0,
    i_10_176_1627_0, i_10_176_1644_0, i_10_176_1645_0, i_10_176_1700_0,
    i_10_176_1727_0, i_10_176_1765_0, i_10_176_1781_0, i_10_176_1795_0,
    i_10_176_1796_0, i_10_176_1826_0, i_10_176_1913_0, i_10_176_2004_0,
    i_10_176_2060_0, i_10_176_2095_0, i_10_176_2245_0, i_10_176_2246_0,
    i_10_176_2248_0, i_10_176_2470_0, i_10_176_2473_0, i_10_176_2474_0,
    i_10_176_2512_0, i_10_176_2516_0, i_10_176_2534_0, i_10_176_2571_0,
    i_10_176_2572_0, i_10_176_2633_0, i_10_176_2708_0, i_10_176_2715_0,
    i_10_176_2789_0, i_10_176_2913_0, i_10_176_2914_0, i_10_176_2915_0,
    i_10_176_2958_0, i_10_176_2983_0, i_10_176_2984_0, i_10_176_3069_0,
    i_10_176_3095_0, i_10_176_3229_0, i_10_176_3356_0, i_10_176_3431_0,
    i_10_176_3451_0, i_10_176_3452_0, i_10_176_3471_0, i_10_176_3472_0,
    i_10_176_3473_0, i_10_176_3496_0, i_10_176_3545_0, i_10_176_3586_0,
    i_10_176_3589_0, i_10_176_3590_0, i_10_176_3603_0, i_10_176_3624_0,
    i_10_176_3625_0, i_10_176_3856_0, i_10_176_3857_0, i_10_176_3885_0,
    i_10_176_3949_0, i_10_176_3950_0, i_10_176_3979_0, i_10_176_4004_0,
    i_10_176_4058_0, i_10_176_4117_0, i_10_176_4120_0, i_10_176_4171_0,
    i_10_176_4265_0, i_10_176_4291_0, i_10_176_4426_0, i_10_176_4481_0,
    o_10_176_0_0  );
  input  i_10_176_34_0, i_10_176_121_0, i_10_176_122_0, i_10_176_124_0,
    i_10_176_132_0, i_10_176_133_0, i_10_176_177_0, i_10_176_178_0,
    i_10_176_183_0, i_10_176_331_0, i_10_176_367_0, i_10_176_374_0,
    i_10_176_386_0, i_10_176_429_0, i_10_176_437_0, i_10_176_439_0,
    i_10_176_440_0, i_10_176_462_0, i_10_176_599_0, i_10_176_600_0,
    i_10_176_602_0, i_10_176_634_0, i_10_176_754_0, i_10_176_755_0,
    i_10_176_906_0, i_10_176_967_0, i_10_176_971_0, i_10_176_1160_0,
    i_10_176_1240_0, i_10_176_1483_0, i_10_176_1499_0, i_10_176_1543_0,
    i_10_176_1627_0, i_10_176_1644_0, i_10_176_1645_0, i_10_176_1700_0,
    i_10_176_1727_0, i_10_176_1765_0, i_10_176_1781_0, i_10_176_1795_0,
    i_10_176_1796_0, i_10_176_1826_0, i_10_176_1913_0, i_10_176_2004_0,
    i_10_176_2060_0, i_10_176_2095_0, i_10_176_2245_0, i_10_176_2246_0,
    i_10_176_2248_0, i_10_176_2470_0, i_10_176_2473_0, i_10_176_2474_0,
    i_10_176_2512_0, i_10_176_2516_0, i_10_176_2534_0, i_10_176_2571_0,
    i_10_176_2572_0, i_10_176_2633_0, i_10_176_2708_0, i_10_176_2715_0,
    i_10_176_2789_0, i_10_176_2913_0, i_10_176_2914_0, i_10_176_2915_0,
    i_10_176_2958_0, i_10_176_2983_0, i_10_176_2984_0, i_10_176_3069_0,
    i_10_176_3095_0, i_10_176_3229_0, i_10_176_3356_0, i_10_176_3431_0,
    i_10_176_3451_0, i_10_176_3452_0, i_10_176_3471_0, i_10_176_3472_0,
    i_10_176_3473_0, i_10_176_3496_0, i_10_176_3545_0, i_10_176_3586_0,
    i_10_176_3589_0, i_10_176_3590_0, i_10_176_3603_0, i_10_176_3624_0,
    i_10_176_3625_0, i_10_176_3856_0, i_10_176_3857_0, i_10_176_3885_0,
    i_10_176_3949_0, i_10_176_3950_0, i_10_176_3979_0, i_10_176_4004_0,
    i_10_176_4058_0, i_10_176_4117_0, i_10_176_4120_0, i_10_176_4171_0,
    i_10_176_4265_0, i_10_176_4291_0, i_10_176_4426_0, i_10_176_4481_0;
  output o_10_176_0_0;
  assign o_10_176_0_0 = 0;
endmodule



// Benchmark "kernel_10_177" written by ABC on Sun Jul 19 10:24:02 2020

module kernel_10_177 ( 
    i_10_177_317_0, i_10_177_325_0, i_10_177_372_0, i_10_177_373_0,
    i_10_177_376_0, i_10_177_388_0, i_10_177_405_0, i_10_177_434_0,
    i_10_177_444_0, i_10_177_446_0, i_10_177_447_0, i_10_177_448_0,
    i_10_177_459_0, i_10_177_462_0, i_10_177_466_0, i_10_177_467_0,
    i_10_177_578_0, i_10_177_736_0, i_10_177_737_0, i_10_177_792_0,
    i_10_177_793_0, i_10_177_794_0, i_10_177_799_0, i_10_177_800_0,
    i_10_177_970_0, i_10_177_1002_0, i_10_177_1003_0, i_10_177_1006_0,
    i_10_177_1116_0, i_10_177_1163_0, i_10_177_1183_0, i_10_177_1242_0,
    i_10_177_1305_0, i_10_177_1306_0, i_10_177_1315_0, i_10_177_1344_0,
    i_10_177_1363_0, i_10_177_1441_0, i_10_177_1442_0, i_10_177_1543_0,
    i_10_177_1549_0, i_10_177_1642_0, i_10_177_1729_0, i_10_177_1730_0,
    i_10_177_1823_0, i_10_177_1826_0, i_10_177_1910_0, i_10_177_1948_0,
    i_10_177_2083_0, i_10_177_2154_0, i_10_177_2157_0, i_10_177_2158_0,
    i_10_177_2305_0, i_10_177_2309_0, i_10_177_2353_0, i_10_177_2404_0,
    i_10_177_2407_0, i_10_177_2408_0, i_10_177_2539_0, i_10_177_2633_0,
    i_10_177_2635_0, i_10_177_2705_0, i_10_177_2782_0, i_10_177_2880_0,
    i_10_177_2881_0, i_10_177_2887_0, i_10_177_2953_0, i_10_177_2956_0,
    i_10_177_2983_0, i_10_177_3058_0, i_10_177_3236_0, i_10_177_3316_0,
    i_10_177_3390_0, i_10_177_3494_0, i_10_177_3508_0, i_10_177_3688_0,
    i_10_177_3835_0, i_10_177_3859_0, i_10_177_3860_0, i_10_177_3889_0,
    i_10_177_3890_0, i_10_177_3919_0, i_10_177_3920_0, i_10_177_3928_0,
    i_10_177_3983_0, i_10_177_4087_0, i_10_177_4088_0, i_10_177_4266_0,
    i_10_177_4268_0, i_10_177_4270_0, i_10_177_4271_0, i_10_177_4273_0,
    i_10_177_4274_0, i_10_177_4288_0, i_10_177_4379_0, i_10_177_4460_0,
    i_10_177_4477_0, i_10_177_4569_0, i_10_177_4570_0, i_10_177_4571_0,
    o_10_177_0_0  );
  input  i_10_177_317_0, i_10_177_325_0, i_10_177_372_0, i_10_177_373_0,
    i_10_177_376_0, i_10_177_388_0, i_10_177_405_0, i_10_177_434_0,
    i_10_177_444_0, i_10_177_446_0, i_10_177_447_0, i_10_177_448_0,
    i_10_177_459_0, i_10_177_462_0, i_10_177_466_0, i_10_177_467_0,
    i_10_177_578_0, i_10_177_736_0, i_10_177_737_0, i_10_177_792_0,
    i_10_177_793_0, i_10_177_794_0, i_10_177_799_0, i_10_177_800_0,
    i_10_177_970_0, i_10_177_1002_0, i_10_177_1003_0, i_10_177_1006_0,
    i_10_177_1116_0, i_10_177_1163_0, i_10_177_1183_0, i_10_177_1242_0,
    i_10_177_1305_0, i_10_177_1306_0, i_10_177_1315_0, i_10_177_1344_0,
    i_10_177_1363_0, i_10_177_1441_0, i_10_177_1442_0, i_10_177_1543_0,
    i_10_177_1549_0, i_10_177_1642_0, i_10_177_1729_0, i_10_177_1730_0,
    i_10_177_1823_0, i_10_177_1826_0, i_10_177_1910_0, i_10_177_1948_0,
    i_10_177_2083_0, i_10_177_2154_0, i_10_177_2157_0, i_10_177_2158_0,
    i_10_177_2305_0, i_10_177_2309_0, i_10_177_2353_0, i_10_177_2404_0,
    i_10_177_2407_0, i_10_177_2408_0, i_10_177_2539_0, i_10_177_2633_0,
    i_10_177_2635_0, i_10_177_2705_0, i_10_177_2782_0, i_10_177_2880_0,
    i_10_177_2881_0, i_10_177_2887_0, i_10_177_2953_0, i_10_177_2956_0,
    i_10_177_2983_0, i_10_177_3058_0, i_10_177_3236_0, i_10_177_3316_0,
    i_10_177_3390_0, i_10_177_3494_0, i_10_177_3508_0, i_10_177_3688_0,
    i_10_177_3835_0, i_10_177_3859_0, i_10_177_3860_0, i_10_177_3889_0,
    i_10_177_3890_0, i_10_177_3919_0, i_10_177_3920_0, i_10_177_3928_0,
    i_10_177_3983_0, i_10_177_4087_0, i_10_177_4088_0, i_10_177_4266_0,
    i_10_177_4268_0, i_10_177_4270_0, i_10_177_4271_0, i_10_177_4273_0,
    i_10_177_4274_0, i_10_177_4288_0, i_10_177_4379_0, i_10_177_4460_0,
    i_10_177_4477_0, i_10_177_4569_0, i_10_177_4570_0, i_10_177_4571_0;
  output o_10_177_0_0;
  assign o_10_177_0_0 = 0;
endmodule



// Benchmark "kernel_10_178" written by ABC on Sun Jul 19 10:24:03 2020

module kernel_10_178 ( 
    i_10_178_28_0, i_10_178_82_0, i_10_178_174_0, i_10_178_176_0,
    i_10_178_246_0, i_10_178_289_0, i_10_178_793_0, i_10_178_954_0,
    i_10_178_955_0, i_10_178_961_0, i_10_178_993_0, i_10_178_1272_0,
    i_10_178_1359_0, i_10_178_1378_0, i_10_178_1575_0, i_10_178_1647_0,
    i_10_178_1648_0, i_10_178_1650_0, i_10_178_1683_0, i_10_178_1684_0,
    i_10_178_1686_0, i_10_178_1687_0, i_10_178_1691_0, i_10_178_1818_0,
    i_10_178_1819_0, i_10_178_1820_0, i_10_178_1916_0, i_10_178_1944_0,
    i_10_178_1945_0, i_10_178_1947_0, i_10_178_2178_0, i_10_178_2325_0,
    i_10_178_2361_0, i_10_178_2376_0, i_10_178_2379_0, i_10_178_2404_0,
    i_10_178_2448_0, i_10_178_2449_0, i_10_178_2450_0, i_10_178_2452_0,
    i_10_178_2453_0, i_10_178_2470_0, i_10_178_2502_0, i_10_178_2503_0,
    i_10_178_2505_0, i_10_178_2514_0, i_10_178_2601_0, i_10_178_2602_0,
    i_10_178_2610_0, i_10_178_2628_0, i_10_178_2631_0, i_10_178_2634_0,
    i_10_178_2637_0, i_10_178_2655_0, i_10_178_2663_0, i_10_178_2673_0,
    i_10_178_2674_0, i_10_178_2676_0, i_10_178_2700_0, i_10_178_2701_0,
    i_10_178_2703_0, i_10_178_2712_0, i_10_178_2727_0, i_10_178_2781_0,
    i_10_178_2882_0, i_10_178_2887_0, i_10_178_3033_0, i_10_178_3036_0,
    i_10_178_3042_0, i_10_178_3051_0, i_10_178_3267_0, i_10_178_3277_0,
    i_10_178_3280_0, i_10_178_3385_0, i_10_178_3386_0, i_10_178_3387_0,
    i_10_178_3388_0, i_10_178_3389_0, i_10_178_3447_0, i_10_178_3448_0,
    i_10_178_3611_0, i_10_178_3645_0, i_10_178_3646_0, i_10_178_3648_0,
    i_10_178_3649_0, i_10_178_3681_0, i_10_178_3783_0, i_10_178_3845_0,
    i_10_178_3852_0, i_10_178_3853_0, i_10_178_3854_0, i_10_178_3860_0,
    i_10_178_3894_0, i_10_178_3979_0, i_10_178_3981_0, i_10_178_4050_0,
    i_10_178_4113_0, i_10_178_4287_0, i_10_178_4564_0, i_10_178_4566_0,
    o_10_178_0_0  );
  input  i_10_178_28_0, i_10_178_82_0, i_10_178_174_0, i_10_178_176_0,
    i_10_178_246_0, i_10_178_289_0, i_10_178_793_0, i_10_178_954_0,
    i_10_178_955_0, i_10_178_961_0, i_10_178_993_0, i_10_178_1272_0,
    i_10_178_1359_0, i_10_178_1378_0, i_10_178_1575_0, i_10_178_1647_0,
    i_10_178_1648_0, i_10_178_1650_0, i_10_178_1683_0, i_10_178_1684_0,
    i_10_178_1686_0, i_10_178_1687_0, i_10_178_1691_0, i_10_178_1818_0,
    i_10_178_1819_0, i_10_178_1820_0, i_10_178_1916_0, i_10_178_1944_0,
    i_10_178_1945_0, i_10_178_1947_0, i_10_178_2178_0, i_10_178_2325_0,
    i_10_178_2361_0, i_10_178_2376_0, i_10_178_2379_0, i_10_178_2404_0,
    i_10_178_2448_0, i_10_178_2449_0, i_10_178_2450_0, i_10_178_2452_0,
    i_10_178_2453_0, i_10_178_2470_0, i_10_178_2502_0, i_10_178_2503_0,
    i_10_178_2505_0, i_10_178_2514_0, i_10_178_2601_0, i_10_178_2602_0,
    i_10_178_2610_0, i_10_178_2628_0, i_10_178_2631_0, i_10_178_2634_0,
    i_10_178_2637_0, i_10_178_2655_0, i_10_178_2663_0, i_10_178_2673_0,
    i_10_178_2674_0, i_10_178_2676_0, i_10_178_2700_0, i_10_178_2701_0,
    i_10_178_2703_0, i_10_178_2712_0, i_10_178_2727_0, i_10_178_2781_0,
    i_10_178_2882_0, i_10_178_2887_0, i_10_178_3033_0, i_10_178_3036_0,
    i_10_178_3042_0, i_10_178_3051_0, i_10_178_3267_0, i_10_178_3277_0,
    i_10_178_3280_0, i_10_178_3385_0, i_10_178_3386_0, i_10_178_3387_0,
    i_10_178_3388_0, i_10_178_3389_0, i_10_178_3447_0, i_10_178_3448_0,
    i_10_178_3611_0, i_10_178_3645_0, i_10_178_3646_0, i_10_178_3648_0,
    i_10_178_3649_0, i_10_178_3681_0, i_10_178_3783_0, i_10_178_3845_0,
    i_10_178_3852_0, i_10_178_3853_0, i_10_178_3854_0, i_10_178_3860_0,
    i_10_178_3894_0, i_10_178_3979_0, i_10_178_3981_0, i_10_178_4050_0,
    i_10_178_4113_0, i_10_178_4287_0, i_10_178_4564_0, i_10_178_4566_0;
  output o_10_178_0_0;
  assign o_10_178_0_0 = ~((~i_10_178_2602_0 & ((~i_10_178_28_0 & ((~i_10_178_954_0 & i_10_178_1687_0) | (~i_10_178_1945_0 & ~i_10_178_2502_0 & ~i_10_178_2701_0 & ~i_10_178_2712_0 & i_10_178_3853_0 & ~i_10_178_3860_0 & ~i_10_178_4050_0))) | (~i_10_178_2505_0 & ~i_10_178_3681_0 & ((~i_10_178_1648_0 & ~i_10_178_1947_0 & ~i_10_178_2404_0 & ~i_10_178_2502_0 & ~i_10_178_2503_0) | (~i_10_178_2325_0 & ~i_10_178_2655_0 & ~i_10_178_2781_0 & ~i_10_178_3783_0 & i_10_178_4113_0))) | (i_10_178_2450_0 & ~i_10_178_2628_0) | (~i_10_178_2631_0 & ~i_10_178_2781_0 & ~i_10_178_3267_0 & ~i_10_178_3845_0))) | (~i_10_178_2376_0 & ((~i_10_178_1647_0 & ~i_10_178_1686_0 & ~i_10_178_1687_0 & ~i_10_178_2325_0 & ~i_10_178_2674_0 & ~i_10_178_2781_0) | (~i_10_178_2703_0 & ~i_10_178_3649_0 & i_10_178_3845_0))) | (~i_10_178_3267_0 & ((~i_10_178_1647_0 & ((~i_10_178_2502_0 & ~i_10_178_2781_0 & ~i_10_178_3645_0) | (~i_10_178_289_0 & ~i_10_178_2655_0 & ~i_10_178_3036_0 & ~i_10_178_3042_0 & ~i_10_178_3611_0 & ~i_10_178_3783_0))) | (~i_10_178_3036_0 & ((i_10_178_1683_0 & ~i_10_178_2610_0 & ~i_10_178_2703_0) | (~i_10_178_2470_0 & ~i_10_178_2673_0 & ~i_10_178_2674_0 & ~i_10_178_3648_0 & ~i_10_178_3681_0 & ~i_10_178_3981_0 & ~i_10_178_4287_0 & i_10_178_4564_0))))) | (~i_10_178_2325_0 & ((~i_10_178_1359_0 & ~i_10_178_2404_0 & ~i_10_178_2505_0 & ~i_10_178_2601_0 & ~i_10_178_2674_0 & ~i_10_178_3033_0 & ~i_10_178_3681_0) | (~i_10_178_1944_0 & ~i_10_178_2502_0 & ~i_10_178_2634_0 & i_10_178_2781_0 & i_10_178_3981_0 & ~i_10_178_4113_0))) | (~i_10_178_2404_0 & ~i_10_178_3845_0 & ((~i_10_178_1359_0 & ~i_10_178_2502_0 & i_10_178_3033_0 & i_10_178_3852_0 & ~i_10_178_3979_0) | (~i_10_178_1819_0 & ~i_10_178_2505_0 & ~i_10_178_2781_0 & ~i_10_178_3645_0 & ~i_10_178_3649_0 & ~i_10_178_4050_0))) | (~i_10_178_1359_0 & ((i_10_178_1818_0 & ~i_10_178_2503_0 & ~i_10_178_2610_0 & i_10_178_2634_0 & ~i_10_178_2673_0 & i_10_178_3860_0) | (~i_10_178_1648_0 & ~i_10_178_2448_0 & ~i_10_178_2452_0 & ~i_10_178_2502_0 & ~i_10_178_2505_0 & ~i_10_178_2663_0 & ~i_10_178_4564_0 & ~i_10_178_4566_0))) | (i_10_178_2449_0 & ((~i_10_178_1916_0 & ~i_10_178_3033_0 & i_10_178_3611_0) | (~i_10_178_246_0 & ~i_10_178_2610_0 & ~i_10_178_4564_0))) | (~i_10_178_3681_0 & ((i_10_178_1819_0 & ~i_10_178_2505_0 & i_10_178_3611_0 & ~i_10_178_3979_0) | (i_10_178_954_0 & ~i_10_178_1820_0 & ~i_10_178_2503_0 & ~i_10_178_2673_0 & i_10_178_3385_0 & ~i_10_178_4050_0 & i_10_178_4564_0 & ~i_10_178_4566_0))) | (i_10_178_1820_0 & ~i_10_178_2502_0 & ~i_10_178_2700_0 & ~i_10_178_2781_0 & ~i_10_178_4050_0));
endmodule



// Benchmark "kernel_10_179" written by ABC on Sun Jul 19 10:24:05 2020

module kernel_10_179 ( 
    i_10_179_248_0, i_10_179_250_0, i_10_179_268_0, i_10_179_321_0,
    i_10_179_408_0, i_10_179_409_0, i_10_179_410_0, i_10_179_425_0,
    i_10_179_441_0, i_10_179_444_0, i_10_179_447_0, i_10_179_463_0,
    i_10_179_466_0, i_10_179_566_0, i_10_179_799_0, i_10_179_958_0,
    i_10_179_969_0, i_10_179_990_0, i_10_179_996_0, i_10_179_1031_0,
    i_10_179_1239_0, i_10_179_1250_0, i_10_179_1263_0, i_10_179_1307_0,
    i_10_179_1344_0, i_10_179_1345_0, i_10_179_1348_0, i_10_179_1439_0,
    i_10_179_1546_0, i_10_179_1576_0, i_10_179_1577_0, i_10_179_1686_0,
    i_10_179_1687_0, i_10_179_1818_0, i_10_179_1819_0, i_10_179_1909_0,
    i_10_179_1912_0, i_10_179_2022_0, i_10_179_2023_0, i_10_179_2032_0,
    i_10_179_2200_0, i_10_179_2201_0, i_10_179_2358_0, i_10_179_2359_0,
    i_10_179_2384_0, i_10_179_2456_0, i_10_179_2474_0, i_10_179_2633_0,
    i_10_179_2700_0, i_10_179_2709_0, i_10_179_2710_0, i_10_179_2713_0,
    i_10_179_2727_0, i_10_179_2731_0, i_10_179_2784_0, i_10_179_2785_0,
    i_10_179_2817_0, i_10_179_2818_0, i_10_179_2883_0, i_10_179_2884_0,
    i_10_179_2887_0, i_10_179_3034_0, i_10_179_3037_0, i_10_179_3038_0,
    i_10_179_3040_0, i_10_179_3069_0, i_10_179_3150_0, i_10_179_3151_0,
    i_10_179_3152_0, i_10_179_3155_0, i_10_179_3157_0, i_10_179_3284_0,
    i_10_179_3384_0, i_10_179_3385_0, i_10_179_3403_0, i_10_179_3472_0,
    i_10_179_3520_0, i_10_179_3522_0, i_10_179_3523_0, i_10_179_3525_0,
    i_10_179_3612_0, i_10_179_3613_0, i_10_179_3781_0, i_10_179_3784_0,
    i_10_179_3847_0, i_10_179_3856_0, i_10_179_3859_0, i_10_179_3983_0,
    i_10_179_3990_0, i_10_179_4114_0, i_10_179_4116_0, i_10_179_4119_0,
    i_10_179_4120_0, i_10_179_4121_0, i_10_179_4266_0, i_10_179_4267_0,
    i_10_179_4271_0, i_10_179_4273_0, i_10_179_4288_0, i_10_179_4290_0,
    o_10_179_0_0  );
  input  i_10_179_248_0, i_10_179_250_0, i_10_179_268_0, i_10_179_321_0,
    i_10_179_408_0, i_10_179_409_0, i_10_179_410_0, i_10_179_425_0,
    i_10_179_441_0, i_10_179_444_0, i_10_179_447_0, i_10_179_463_0,
    i_10_179_466_0, i_10_179_566_0, i_10_179_799_0, i_10_179_958_0,
    i_10_179_969_0, i_10_179_990_0, i_10_179_996_0, i_10_179_1031_0,
    i_10_179_1239_0, i_10_179_1250_0, i_10_179_1263_0, i_10_179_1307_0,
    i_10_179_1344_0, i_10_179_1345_0, i_10_179_1348_0, i_10_179_1439_0,
    i_10_179_1546_0, i_10_179_1576_0, i_10_179_1577_0, i_10_179_1686_0,
    i_10_179_1687_0, i_10_179_1818_0, i_10_179_1819_0, i_10_179_1909_0,
    i_10_179_1912_0, i_10_179_2022_0, i_10_179_2023_0, i_10_179_2032_0,
    i_10_179_2200_0, i_10_179_2201_0, i_10_179_2358_0, i_10_179_2359_0,
    i_10_179_2384_0, i_10_179_2456_0, i_10_179_2474_0, i_10_179_2633_0,
    i_10_179_2700_0, i_10_179_2709_0, i_10_179_2710_0, i_10_179_2713_0,
    i_10_179_2727_0, i_10_179_2731_0, i_10_179_2784_0, i_10_179_2785_0,
    i_10_179_2817_0, i_10_179_2818_0, i_10_179_2883_0, i_10_179_2884_0,
    i_10_179_2887_0, i_10_179_3034_0, i_10_179_3037_0, i_10_179_3038_0,
    i_10_179_3040_0, i_10_179_3069_0, i_10_179_3150_0, i_10_179_3151_0,
    i_10_179_3152_0, i_10_179_3155_0, i_10_179_3157_0, i_10_179_3284_0,
    i_10_179_3384_0, i_10_179_3385_0, i_10_179_3403_0, i_10_179_3472_0,
    i_10_179_3520_0, i_10_179_3522_0, i_10_179_3523_0, i_10_179_3525_0,
    i_10_179_3612_0, i_10_179_3613_0, i_10_179_3781_0, i_10_179_3784_0,
    i_10_179_3847_0, i_10_179_3856_0, i_10_179_3859_0, i_10_179_3983_0,
    i_10_179_3990_0, i_10_179_4114_0, i_10_179_4116_0, i_10_179_4119_0,
    i_10_179_4120_0, i_10_179_4121_0, i_10_179_4266_0, i_10_179_4267_0,
    i_10_179_4271_0, i_10_179_4273_0, i_10_179_4288_0, i_10_179_4290_0;
  output o_10_179_0_0;
  assign o_10_179_0_0 = ~((i_10_179_466_0 & ((~i_10_179_2784_0 & ~i_10_179_3403_0 & ~i_10_179_3613_0 & ~i_10_179_3990_0) | (~i_10_179_990_0 & ~i_10_179_1348_0 & ~i_10_179_2817_0 & ~i_10_179_3525_0 & ~i_10_179_3983_0 & ~i_10_179_4116_0))) | (~i_10_179_990_0 & ((~i_10_179_250_0 & ~i_10_179_410_0 & ~i_10_179_996_0 & ~i_10_179_1345_0 & ~i_10_179_2022_0 & ~i_10_179_2709_0 & ~i_10_179_3523_0 & ~i_10_179_3990_0) | (~i_10_179_799_0 & ~i_10_179_958_0 & i_10_179_2359_0 & i_10_179_2727_0 & ~i_10_179_3784_0 & ~i_10_179_4121_0))) | (~i_10_179_1263_0 & ((~i_10_179_250_0 & ~i_10_179_410_0 & ~i_10_179_2384_0 & i_10_179_2633_0 & ~i_10_179_3384_0 & i_10_179_3523_0) | (~i_10_179_408_0 & ~i_10_179_409_0 & ~i_10_179_1348_0 & ~i_10_179_1909_0 & ~i_10_179_2887_0 & ~i_10_179_3403_0 & ~i_10_179_3781_0 & ~i_10_179_3856_0 & ~i_10_179_3990_0))) | (~i_10_179_250_0 & ((~i_10_179_408_0 & ~i_10_179_466_0 & ~i_10_179_1348_0 & ~i_10_179_1686_0 & ~i_10_179_1818_0 & ~i_10_179_2200_0 & ~i_10_179_2384_0 & ~i_10_179_2700_0 & ~i_10_179_2710_0 & ~i_10_179_3284_0 & ~i_10_179_3385_0 & ~i_10_179_4119_0 & ~i_10_179_4273_0) | (~i_10_179_410_0 & ~i_10_179_2713_0 & ~i_10_179_3523_0 & ~i_10_179_3612_0 & i_10_179_3856_0 & ~i_10_179_3990_0 & ~i_10_179_4288_0))) | (~i_10_179_1348_0 & ((~i_10_179_248_0 & ~i_10_179_2785_0 & ~i_10_179_2883_0 & ~i_10_179_3384_0 & ~i_10_179_3522_0 & ~i_10_179_3856_0 & ~i_10_179_4120_0) | (~i_10_179_996_0 & i_10_179_2201_0 & ~i_10_179_3038_0 & ~i_10_179_3784_0 & ~i_10_179_3990_0 & ~i_10_179_4290_0))) | (~i_10_179_996_0 & ((~i_10_179_410_0 & ~i_10_179_1909_0 & ~i_10_179_2023_0 & ~i_10_179_2784_0 & ~i_10_179_3983_0 & ~i_10_179_4116_0 & ~i_10_179_2818_0 & ~i_10_179_3384_0) | (i_10_179_3781_0 & i_10_179_3784_0 & ~i_10_179_4288_0))) | (i_10_179_2633_0 & ((~i_10_179_1344_0 & ~i_10_179_1912_0 & ~i_10_179_2818_0 & ~i_10_179_3523_0 & ~i_10_179_3990_0 & ~i_10_179_4116_0) | (i_10_179_958_0 & ~i_10_179_4121_0))) | (~i_10_179_409_0 & ((~i_10_179_2710_0 & ((~i_10_179_410_0 & ~i_10_179_566_0 & ~i_10_179_1239_0 & ~i_10_179_2359_0 & ~i_10_179_2474_0 & ~i_10_179_2709_0 & ~i_10_179_2887_0 & ~i_10_179_3781_0 & ~i_10_179_4114_0) | (~i_10_179_463_0 & ~i_10_179_2201_0 & ~i_10_179_3520_0 & ~i_10_179_3525_0 & i_10_179_4116_0 & ~i_10_179_4120_0))) | (i_10_179_1819_0 & ~i_10_179_2883_0 & ~i_10_179_3522_0 & ~i_10_179_3525_0))) | (~i_10_179_408_0 & ((~i_10_179_410_0 & ((i_10_179_248_0 & ~i_10_179_441_0 & ~i_10_179_2384_0 & ~i_10_179_2883_0 & ~i_10_179_3612_0) | (~i_10_179_1912_0 & ~i_10_179_3385_0 & ~i_10_179_3403_0 & ~i_10_179_3613_0 & ~i_10_179_4119_0))) | (~i_10_179_4288_0 & ((~i_10_179_1912_0 & i_10_179_2201_0 & ~i_10_179_2883_0 & ~i_10_179_2884_0) | (~i_10_179_1818_0 & ~i_10_179_2713_0 & i_10_179_2731_0 & ~i_10_179_3403_0 & ~i_10_179_3523_0 & ~i_10_179_3612_0 & ~i_10_179_4271_0 & ~i_10_179_4290_0))))) | (~i_10_179_3990_0 & ((~i_10_179_1345_0 & i_10_179_2731_0 & ~i_10_179_2818_0 & i_10_179_3612_0 & ~i_10_179_4119_0) | (i_10_179_3385_0 & i_10_179_3847_0 & ~i_10_179_3856_0 & ~i_10_179_4114_0 & ~i_10_179_4120_0))) | (~i_10_179_3522_0 & ~i_10_179_3525_0 & i_10_179_1239_0 & ~i_10_179_2887_0) | (~i_10_179_1912_0 & ~i_10_179_2884_0 & ~i_10_179_3385_0 & i_10_179_3856_0 & ~i_10_179_4119_0 & ~i_10_179_4121_0));
endmodule



// Benchmark "kernel_10_180" written by ABC on Sun Jul 19 10:24:06 2020

module kernel_10_180 ( 
    i_10_180_22_0, i_10_180_23_0, i_10_180_86_0, i_10_180_245_0,
    i_10_180_248_0, i_10_180_262_0, i_10_180_283_0, i_10_180_284_0,
    i_10_180_317_0, i_10_180_319_0, i_10_180_320_0, i_10_180_391_0,
    i_10_180_439_0, i_10_180_460_0, i_10_180_464_0, i_10_180_479_0,
    i_10_180_496_0, i_10_180_497_0, i_10_180_832_0, i_10_180_932_0,
    i_10_180_947_0, i_10_180_1001_0, i_10_180_1085_0, i_10_180_1223_0,
    i_10_180_1240_0, i_10_180_1243_0, i_10_180_1267_0, i_10_180_1301_0,
    i_10_180_1328_0, i_10_180_1346_0, i_10_180_1433_0, i_10_180_1445_0,
    i_10_180_1487_0, i_10_180_1541_0, i_10_180_1544_0, i_10_180_1577_0,
    i_10_180_1607_0, i_10_180_1622_0, i_10_180_1624_0, i_10_180_1625_0,
    i_10_180_1687_0, i_10_180_1714_0, i_10_180_1741_0, i_10_180_1805_0,
    i_10_180_1821_0, i_10_180_1826_0, i_10_180_1931_0, i_10_180_2017_0,
    i_10_180_2018_0, i_10_180_2026_0, i_10_180_2027_0, i_10_180_2110_0,
    i_10_180_2111_0, i_10_180_2162_0, i_10_180_2198_0, i_10_180_2204_0,
    i_10_180_2359_0, i_10_180_2366_0, i_10_180_2453_0, i_10_180_2567_0,
    i_10_180_2602_0, i_10_180_2605_0, i_10_180_2606_0, i_10_180_2663_0,
    i_10_180_2702_0, i_10_180_2705_0, i_10_180_2719_0, i_10_180_2725_0,
    i_10_180_2732_0, i_10_180_2846_0, i_10_180_2924_0, i_10_180_3025_0,
    i_10_180_3044_0, i_10_180_3070_0, i_10_180_3077_0, i_10_180_3167_0,
    i_10_180_3317_0, i_10_180_3332_0, i_10_180_3377_0, i_10_180_3389_0,
    i_10_180_3523_0, i_10_180_3557_0, i_10_180_3602_0, i_10_180_3613_0,
    i_10_180_3722_0, i_10_180_3725_0, i_10_180_3772_0, i_10_180_3835_0,
    i_10_180_3841_0, i_10_180_3851_0, i_10_180_3856_0, i_10_180_3916_0,
    i_10_180_3989_0, i_10_180_4096_0, i_10_180_4097_0, i_10_180_4114_0,
    i_10_180_4117_0, i_10_180_4123_0, i_10_180_4124_0, i_10_180_4276_0,
    o_10_180_0_0  );
  input  i_10_180_22_0, i_10_180_23_0, i_10_180_86_0, i_10_180_245_0,
    i_10_180_248_0, i_10_180_262_0, i_10_180_283_0, i_10_180_284_0,
    i_10_180_317_0, i_10_180_319_0, i_10_180_320_0, i_10_180_391_0,
    i_10_180_439_0, i_10_180_460_0, i_10_180_464_0, i_10_180_479_0,
    i_10_180_496_0, i_10_180_497_0, i_10_180_832_0, i_10_180_932_0,
    i_10_180_947_0, i_10_180_1001_0, i_10_180_1085_0, i_10_180_1223_0,
    i_10_180_1240_0, i_10_180_1243_0, i_10_180_1267_0, i_10_180_1301_0,
    i_10_180_1328_0, i_10_180_1346_0, i_10_180_1433_0, i_10_180_1445_0,
    i_10_180_1487_0, i_10_180_1541_0, i_10_180_1544_0, i_10_180_1577_0,
    i_10_180_1607_0, i_10_180_1622_0, i_10_180_1624_0, i_10_180_1625_0,
    i_10_180_1687_0, i_10_180_1714_0, i_10_180_1741_0, i_10_180_1805_0,
    i_10_180_1821_0, i_10_180_1826_0, i_10_180_1931_0, i_10_180_2017_0,
    i_10_180_2018_0, i_10_180_2026_0, i_10_180_2027_0, i_10_180_2110_0,
    i_10_180_2111_0, i_10_180_2162_0, i_10_180_2198_0, i_10_180_2204_0,
    i_10_180_2359_0, i_10_180_2366_0, i_10_180_2453_0, i_10_180_2567_0,
    i_10_180_2602_0, i_10_180_2605_0, i_10_180_2606_0, i_10_180_2663_0,
    i_10_180_2702_0, i_10_180_2705_0, i_10_180_2719_0, i_10_180_2725_0,
    i_10_180_2732_0, i_10_180_2846_0, i_10_180_2924_0, i_10_180_3025_0,
    i_10_180_3044_0, i_10_180_3070_0, i_10_180_3077_0, i_10_180_3167_0,
    i_10_180_3317_0, i_10_180_3332_0, i_10_180_3377_0, i_10_180_3389_0,
    i_10_180_3523_0, i_10_180_3557_0, i_10_180_3602_0, i_10_180_3613_0,
    i_10_180_3722_0, i_10_180_3725_0, i_10_180_3772_0, i_10_180_3835_0,
    i_10_180_3841_0, i_10_180_3851_0, i_10_180_3856_0, i_10_180_3916_0,
    i_10_180_3989_0, i_10_180_4096_0, i_10_180_4097_0, i_10_180_4114_0,
    i_10_180_4117_0, i_10_180_4123_0, i_10_180_4124_0, i_10_180_4276_0;
  output o_10_180_0_0;
  assign o_10_180_0_0 = 0;
endmodule



// Benchmark "kernel_10_181" written by ABC on Sun Jul 19 10:24:07 2020

module kernel_10_181 ( 
    i_10_181_85_0, i_10_181_86_0, i_10_181_155_0, i_10_181_158_0,
    i_10_181_243_0, i_10_181_245_0, i_10_181_246_0, i_10_181_287_0,
    i_10_181_319_0, i_10_181_374_0, i_10_181_405_0, i_10_181_423_0,
    i_10_181_436_0, i_10_181_460_0, i_10_181_462_0, i_10_181_463_0,
    i_10_181_466_0, i_10_181_948_0, i_10_181_990_0, i_10_181_991_0,
    i_10_181_992_0, i_10_181_1031_0, i_10_181_1053_0, i_10_181_1173_0,
    i_10_181_1201_0, i_10_181_1202_0, i_10_181_1217_0, i_10_181_1260_0,
    i_10_181_1307_0, i_10_181_1358_0, i_10_181_1443_0, i_10_181_1444_0,
    i_10_181_1543_0, i_10_181_1596_0, i_10_181_1608_0, i_10_181_1622_0,
    i_10_181_1647_0, i_10_181_1648_0, i_10_181_1649_0, i_10_181_1651_0,
    i_10_181_1713_0, i_10_181_1994_0, i_10_181_2000_0, i_10_181_2016_0,
    i_10_181_2018_0, i_10_181_2201_0, i_10_181_2204_0, i_10_181_2324_0,
    i_10_181_2357_0, i_10_181_2459_0, i_10_181_2460_0, i_10_181_2512_0,
    i_10_181_2513_0, i_10_181_2606_0, i_10_181_2641_0, i_10_181_2659_0,
    i_10_181_2660_0, i_10_181_2720_0, i_10_181_2721_0, i_10_181_2725_0,
    i_10_181_2726_0, i_10_181_2782_0, i_10_181_2828_0, i_10_181_2834_0,
    i_10_181_2884_0, i_10_181_2964_0, i_10_181_2965_0, i_10_181_2981_0,
    i_10_181_2984_0, i_10_181_3044_0, i_10_181_3083_0, i_10_181_3201_0,
    i_10_181_3259_0, i_10_181_3272_0, i_10_181_3442_0, i_10_181_3443_0,
    i_10_181_3611_0, i_10_181_3721_0, i_10_181_3722_0, i_10_181_3788_0,
    i_10_181_3807_0, i_10_181_3830_0, i_10_181_3857_0, i_10_181_3860_0,
    i_10_181_3893_0, i_10_181_3910_0, i_10_181_3926_0, i_10_181_3980_0,
    i_10_181_3988_0, i_10_181_4030_0, i_10_181_4031_0, i_10_181_4114_0,
    i_10_181_4115_0, i_10_181_4169_0, i_10_181_4214_0, i_10_181_4277_0,
    i_10_181_4286_0, i_10_181_4317_0, i_10_181_4456_0, i_10_181_4521_0,
    o_10_181_0_0  );
  input  i_10_181_85_0, i_10_181_86_0, i_10_181_155_0, i_10_181_158_0,
    i_10_181_243_0, i_10_181_245_0, i_10_181_246_0, i_10_181_287_0,
    i_10_181_319_0, i_10_181_374_0, i_10_181_405_0, i_10_181_423_0,
    i_10_181_436_0, i_10_181_460_0, i_10_181_462_0, i_10_181_463_0,
    i_10_181_466_0, i_10_181_948_0, i_10_181_990_0, i_10_181_991_0,
    i_10_181_992_0, i_10_181_1031_0, i_10_181_1053_0, i_10_181_1173_0,
    i_10_181_1201_0, i_10_181_1202_0, i_10_181_1217_0, i_10_181_1260_0,
    i_10_181_1307_0, i_10_181_1358_0, i_10_181_1443_0, i_10_181_1444_0,
    i_10_181_1543_0, i_10_181_1596_0, i_10_181_1608_0, i_10_181_1622_0,
    i_10_181_1647_0, i_10_181_1648_0, i_10_181_1649_0, i_10_181_1651_0,
    i_10_181_1713_0, i_10_181_1994_0, i_10_181_2000_0, i_10_181_2016_0,
    i_10_181_2018_0, i_10_181_2201_0, i_10_181_2204_0, i_10_181_2324_0,
    i_10_181_2357_0, i_10_181_2459_0, i_10_181_2460_0, i_10_181_2512_0,
    i_10_181_2513_0, i_10_181_2606_0, i_10_181_2641_0, i_10_181_2659_0,
    i_10_181_2660_0, i_10_181_2720_0, i_10_181_2721_0, i_10_181_2725_0,
    i_10_181_2726_0, i_10_181_2782_0, i_10_181_2828_0, i_10_181_2834_0,
    i_10_181_2884_0, i_10_181_2964_0, i_10_181_2965_0, i_10_181_2981_0,
    i_10_181_2984_0, i_10_181_3044_0, i_10_181_3083_0, i_10_181_3201_0,
    i_10_181_3259_0, i_10_181_3272_0, i_10_181_3442_0, i_10_181_3443_0,
    i_10_181_3611_0, i_10_181_3721_0, i_10_181_3722_0, i_10_181_3788_0,
    i_10_181_3807_0, i_10_181_3830_0, i_10_181_3857_0, i_10_181_3860_0,
    i_10_181_3893_0, i_10_181_3910_0, i_10_181_3926_0, i_10_181_3980_0,
    i_10_181_3988_0, i_10_181_4030_0, i_10_181_4031_0, i_10_181_4114_0,
    i_10_181_4115_0, i_10_181_4169_0, i_10_181_4214_0, i_10_181_4277_0,
    i_10_181_4286_0, i_10_181_4317_0, i_10_181_4456_0, i_10_181_4521_0;
  output o_10_181_0_0;
  assign o_10_181_0_0 = 0;
endmodule



// Benchmark "kernel_10_182" written by ABC on Sun Jul 19 10:24:08 2020

module kernel_10_182 ( 
    i_10_182_172_0, i_10_182_244_0, i_10_182_246_0, i_10_182_247_0,
    i_10_182_253_0, i_10_182_276_0, i_10_182_286_0, i_10_182_405_0,
    i_10_182_426_0, i_10_182_427_0, i_10_182_460_0, i_10_182_467_0,
    i_10_182_747_0, i_10_182_748_0, i_10_182_954_0, i_10_182_955_0,
    i_10_182_956_0, i_10_182_962_0, i_10_182_1026_0, i_10_182_1029_0,
    i_10_182_1234_0, i_10_182_1236_0, i_10_182_1237_0, i_10_182_1241_0,
    i_10_182_1243_0, i_10_182_1308_0, i_10_182_1309_0, i_10_182_1311_0,
    i_10_182_1312_0, i_10_182_1540_0, i_10_182_1542_0, i_10_182_1545_0,
    i_10_182_1650_0, i_10_182_1686_0, i_10_182_1688_0, i_10_182_1818_0,
    i_10_182_1819_0, i_10_182_1820_0, i_10_182_1826_0, i_10_182_1953_0,
    i_10_182_2196_0, i_10_182_2351_0, i_10_182_2354_0, i_10_182_2450_0,
    i_10_182_2452_0, i_10_182_2469_0, i_10_182_2474_0, i_10_182_2601_0,
    i_10_182_2674_0, i_10_182_2677_0, i_10_182_2710_0, i_10_182_2711_0,
    i_10_182_2719_0, i_10_182_2731_0, i_10_182_2917_0, i_10_182_2924_0,
    i_10_182_2980_0, i_10_182_3036_0, i_10_182_3072_0, i_10_182_3075_0,
    i_10_182_3198_0, i_10_182_3199_0, i_10_182_3200_0, i_10_182_3202_0,
    i_10_182_3385_0, i_10_182_3408_0, i_10_182_3522_0, i_10_182_3523_0,
    i_10_182_3582_0, i_10_182_3585_0, i_10_182_3586_0, i_10_182_3612_0,
    i_10_182_3613_0, i_10_182_3615_0, i_10_182_3646_0, i_10_182_3648_0,
    i_10_182_3649_0, i_10_182_3780_0, i_10_182_3781_0, i_10_182_3782_0,
    i_10_182_3783_0, i_10_182_3784_0, i_10_182_3786_0, i_10_182_3787_0,
    i_10_182_3788_0, i_10_182_3835_0, i_10_182_3840_0, i_10_182_3856_0,
    i_10_182_4113_0, i_10_182_4114_0, i_10_182_4116_0, i_10_182_4117_0,
    i_10_182_4216_0, i_10_182_4267_0, i_10_182_4284_0, i_10_182_4288_0,
    i_10_182_4563_0, i_10_182_4564_0, i_10_182_4567_0, i_10_182_4568_0,
    o_10_182_0_0  );
  input  i_10_182_172_0, i_10_182_244_0, i_10_182_246_0, i_10_182_247_0,
    i_10_182_253_0, i_10_182_276_0, i_10_182_286_0, i_10_182_405_0,
    i_10_182_426_0, i_10_182_427_0, i_10_182_460_0, i_10_182_467_0,
    i_10_182_747_0, i_10_182_748_0, i_10_182_954_0, i_10_182_955_0,
    i_10_182_956_0, i_10_182_962_0, i_10_182_1026_0, i_10_182_1029_0,
    i_10_182_1234_0, i_10_182_1236_0, i_10_182_1237_0, i_10_182_1241_0,
    i_10_182_1243_0, i_10_182_1308_0, i_10_182_1309_0, i_10_182_1311_0,
    i_10_182_1312_0, i_10_182_1540_0, i_10_182_1542_0, i_10_182_1545_0,
    i_10_182_1650_0, i_10_182_1686_0, i_10_182_1688_0, i_10_182_1818_0,
    i_10_182_1819_0, i_10_182_1820_0, i_10_182_1826_0, i_10_182_1953_0,
    i_10_182_2196_0, i_10_182_2351_0, i_10_182_2354_0, i_10_182_2450_0,
    i_10_182_2452_0, i_10_182_2469_0, i_10_182_2474_0, i_10_182_2601_0,
    i_10_182_2674_0, i_10_182_2677_0, i_10_182_2710_0, i_10_182_2711_0,
    i_10_182_2719_0, i_10_182_2731_0, i_10_182_2917_0, i_10_182_2924_0,
    i_10_182_2980_0, i_10_182_3036_0, i_10_182_3072_0, i_10_182_3075_0,
    i_10_182_3198_0, i_10_182_3199_0, i_10_182_3200_0, i_10_182_3202_0,
    i_10_182_3385_0, i_10_182_3408_0, i_10_182_3522_0, i_10_182_3523_0,
    i_10_182_3582_0, i_10_182_3585_0, i_10_182_3586_0, i_10_182_3612_0,
    i_10_182_3613_0, i_10_182_3615_0, i_10_182_3646_0, i_10_182_3648_0,
    i_10_182_3649_0, i_10_182_3780_0, i_10_182_3781_0, i_10_182_3782_0,
    i_10_182_3783_0, i_10_182_3784_0, i_10_182_3786_0, i_10_182_3787_0,
    i_10_182_3788_0, i_10_182_3835_0, i_10_182_3840_0, i_10_182_3856_0,
    i_10_182_4113_0, i_10_182_4114_0, i_10_182_4116_0, i_10_182_4117_0,
    i_10_182_4216_0, i_10_182_4267_0, i_10_182_4284_0, i_10_182_4288_0,
    i_10_182_4563_0, i_10_182_4564_0, i_10_182_4567_0, i_10_182_4568_0;
  output o_10_182_0_0;
  assign o_10_182_0_0 = ~((~i_10_182_246_0 & ((i_10_182_286_0 & ~i_10_182_1026_0 & ~i_10_182_1241_0 & ~i_10_182_2469_0 & ~i_10_182_3200_0 & ~i_10_182_3787_0) | (~i_10_182_1243_0 & ~i_10_182_3036_0 & ~i_10_182_3615_0 & ~i_10_182_3783_0 & ~i_10_182_3788_0 & ~i_10_182_4113_0 & ~i_10_182_4216_0))) | (~i_10_182_244_0 & ((~i_10_182_247_0 & ((~i_10_182_747_0 & ~i_10_182_748_0 & ~i_10_182_954_0 & i_10_182_1819_0) | (~i_10_182_962_0 & ~i_10_182_1029_0 & ~i_10_182_2601_0 & ~i_10_182_3198_0 & ~i_10_182_3783_0 & ~i_10_182_4216_0))) | (~i_10_182_3840_0 & ((~i_10_182_2719_0 & ~i_10_182_3198_0 & ~i_10_182_3385_0 & ~i_10_182_3786_0 & ~i_10_182_3856_0) | (~i_10_182_748_0 & ~i_10_182_962_0 & ~i_10_182_1308_0 & ~i_10_182_1542_0 & ~i_10_182_1545_0 & ~i_10_182_2452_0 & ~i_10_182_3072_0 & ~i_10_182_3075_0 & ~i_10_182_4216_0))) | (~i_10_182_1820_0 & ~i_10_182_2196_0 & ~i_10_182_2351_0 & i_10_182_3385_0 & ~i_10_182_4113_0 & ~i_10_182_4284_0))) | (~i_10_182_748_0 & ((~i_10_182_1026_0 & i_10_182_1819_0 & ~i_10_182_2601_0 & ~i_10_182_3582_0 & ~i_10_182_3787_0 & ~i_10_182_3788_0 & ~i_10_182_4216_0) | (~i_10_182_253_0 & ~i_10_182_3036_0 & ~i_10_182_3075_0 & ~i_10_182_3780_0 & i_10_182_4567_0))) | (~i_10_182_2351_0 & ((~i_10_182_1311_0 & ((i_10_182_2354_0 & ~i_10_182_3199_0 & ~i_10_182_3613_0 & ~i_10_182_3786_0) | (~i_10_182_405_0 & ~i_10_182_1029_0 & ~i_10_182_1241_0 & ~i_10_182_1243_0 & ~i_10_182_2450_0 & ~i_10_182_2601_0 & ~i_10_182_2980_0 & ~i_10_182_3072_0 & ~i_10_182_3408_0 & ~i_10_182_3787_0 & ~i_10_182_3788_0 & ~i_10_182_3840_0 & ~i_10_182_4216_0))) | (~i_10_182_1026_0 & ~i_10_182_2469_0 & i_10_182_3523_0 & i_10_182_3615_0 & ~i_10_182_3787_0 & ~i_10_182_4564_0))) | (~i_10_182_1026_0 & ((~i_10_182_747_0 & ~i_10_182_3612_0 & ~i_10_182_3786_0 & i_10_182_3835_0) | (~i_10_182_956_0 & i_10_182_1686_0 & ~i_10_182_3036_0 & ~i_10_182_3835_0 & ~i_10_182_4216_0 & ~i_10_182_4267_0))) | (~i_10_182_3783_0 & ((~i_10_182_747_0 & ~i_10_182_2196_0 & ((~i_10_182_1312_0 & ~i_10_182_3784_0) | (~i_10_182_3202_0 & ~i_10_182_3385_0 & ~i_10_182_3615_0 & ~i_10_182_3788_0 & ~i_10_182_3840_0))) | (~i_10_182_1029_0 & ~i_10_182_2601_0 & ~i_10_182_3200_0 & ~i_10_182_3612_0 & ~i_10_182_3781_0) | (~i_10_182_3408_0 & i_10_182_3615_0 & ~i_10_182_3788_0 & ~i_10_182_3856_0 & ~i_10_182_4116_0))) | (i_10_182_3036_0 & ~i_10_182_3615_0 & ((i_10_182_1236_0 & ~i_10_182_3202_0 & ~i_10_182_3840_0 & ~i_10_182_4114_0) | (~i_10_182_1029_0 & ~i_10_182_1236_0 & i_10_182_3200_0 & i_10_182_3856_0 & ~i_10_182_4117_0))) | (~i_10_182_4117_0 & ((i_10_182_172_0 & i_10_182_2354_0) | i_10_182_4288_0 | (~i_10_182_1650_0 & ~i_10_182_2601_0 & ~i_10_182_3198_0 & ~i_10_182_3199_0))) | (i_10_182_286_0 & ~i_10_182_1826_0 & ~i_10_182_2196_0 & ~i_10_182_3787_0 & ~i_10_182_3840_0) | (~i_10_182_1542_0 & i_10_182_3585_0 & i_10_182_3586_0 & ~i_10_182_4564_0) | (i_10_182_1234_0 & ~i_10_182_1545_0 & ~i_10_182_1820_0 & ~i_10_182_3780_0 & ~i_10_182_4567_0));
endmodule



// Benchmark "kernel_10_183" written by ABC on Sun Jul 19 10:24:09 2020

module kernel_10_183 ( 
    i_10_183_117_0, i_10_183_118_0, i_10_183_136_0, i_10_183_146_0,
    i_10_183_175_0, i_10_183_216_0, i_10_183_220_0, i_10_183_263_0,
    i_10_183_284_0, i_10_183_308_0, i_10_183_347_0, i_10_183_390_0,
    i_10_183_391_0, i_10_183_435_0, i_10_183_508_0, i_10_183_509_0,
    i_10_183_689_0, i_10_183_748_0, i_10_183_892_0, i_10_183_901_0,
    i_10_183_902_0, i_10_183_963_0, i_10_183_1045_0, i_10_183_1046_0,
    i_10_183_1083_0, i_10_183_1234_0, i_10_183_1238_0, i_10_183_1246_0,
    i_10_183_1247_0, i_10_183_1432_0, i_10_183_1433_0, i_10_183_1451_0,
    i_10_183_1534_0, i_10_183_1621_0, i_10_183_1622_0, i_10_183_1683_0,
    i_10_183_1686_0, i_10_183_1689_0, i_10_183_1691_0, i_10_183_1821_0,
    i_10_183_1901_0, i_10_183_1908_0, i_10_183_1909_0, i_10_183_1944_0,
    i_10_183_2035_0, i_10_183_2161_0, i_10_183_2243_0, i_10_183_2246_0,
    i_10_183_2252_0, i_10_183_2326_0, i_10_183_2448_0, i_10_183_2449_0,
    i_10_183_2453_0, i_10_183_2467_0, i_10_183_2468_0, i_10_183_2469_0,
    i_10_183_2512_0, i_10_183_2513_0, i_10_183_2544_0, i_10_183_2565_0,
    i_10_183_2629_0, i_10_183_2630_0, i_10_183_2632_0, i_10_183_2638_0,
    i_10_183_2655_0, i_10_183_2656_0, i_10_183_2663_0, i_10_183_2700_0,
    i_10_183_2718_0, i_10_183_2723_0, i_10_183_2728_0, i_10_183_2911_0,
    i_10_183_3043_0, i_10_183_3069_0, i_10_183_3071_0, i_10_183_3170_0,
    i_10_183_3392_0, i_10_183_3408_0, i_10_183_3409_0, i_10_183_3449_0,
    i_10_183_3465_0, i_10_183_3469_0, i_10_183_3527_0, i_10_183_3538_0,
    i_10_183_3555_0, i_10_183_3562_0, i_10_183_3583_0, i_10_183_3609_0,
    i_10_183_3837_0, i_10_183_3856_0, i_10_183_4121_0, i_10_183_4122_0,
    i_10_183_4278_0, i_10_183_4285_0, i_10_183_4286_0, i_10_183_4288_0,
    i_10_183_4289_0, i_10_183_4428_0, i_10_183_4570_0, i_10_183_4582_0,
    o_10_183_0_0  );
  input  i_10_183_117_0, i_10_183_118_0, i_10_183_136_0, i_10_183_146_0,
    i_10_183_175_0, i_10_183_216_0, i_10_183_220_0, i_10_183_263_0,
    i_10_183_284_0, i_10_183_308_0, i_10_183_347_0, i_10_183_390_0,
    i_10_183_391_0, i_10_183_435_0, i_10_183_508_0, i_10_183_509_0,
    i_10_183_689_0, i_10_183_748_0, i_10_183_892_0, i_10_183_901_0,
    i_10_183_902_0, i_10_183_963_0, i_10_183_1045_0, i_10_183_1046_0,
    i_10_183_1083_0, i_10_183_1234_0, i_10_183_1238_0, i_10_183_1246_0,
    i_10_183_1247_0, i_10_183_1432_0, i_10_183_1433_0, i_10_183_1451_0,
    i_10_183_1534_0, i_10_183_1621_0, i_10_183_1622_0, i_10_183_1683_0,
    i_10_183_1686_0, i_10_183_1689_0, i_10_183_1691_0, i_10_183_1821_0,
    i_10_183_1901_0, i_10_183_1908_0, i_10_183_1909_0, i_10_183_1944_0,
    i_10_183_2035_0, i_10_183_2161_0, i_10_183_2243_0, i_10_183_2246_0,
    i_10_183_2252_0, i_10_183_2326_0, i_10_183_2448_0, i_10_183_2449_0,
    i_10_183_2453_0, i_10_183_2467_0, i_10_183_2468_0, i_10_183_2469_0,
    i_10_183_2512_0, i_10_183_2513_0, i_10_183_2544_0, i_10_183_2565_0,
    i_10_183_2629_0, i_10_183_2630_0, i_10_183_2632_0, i_10_183_2638_0,
    i_10_183_2655_0, i_10_183_2656_0, i_10_183_2663_0, i_10_183_2700_0,
    i_10_183_2718_0, i_10_183_2723_0, i_10_183_2728_0, i_10_183_2911_0,
    i_10_183_3043_0, i_10_183_3069_0, i_10_183_3071_0, i_10_183_3170_0,
    i_10_183_3392_0, i_10_183_3408_0, i_10_183_3409_0, i_10_183_3449_0,
    i_10_183_3465_0, i_10_183_3469_0, i_10_183_3527_0, i_10_183_3538_0,
    i_10_183_3555_0, i_10_183_3562_0, i_10_183_3583_0, i_10_183_3609_0,
    i_10_183_3837_0, i_10_183_3856_0, i_10_183_4121_0, i_10_183_4122_0,
    i_10_183_4278_0, i_10_183_4285_0, i_10_183_4286_0, i_10_183_4288_0,
    i_10_183_4289_0, i_10_183_4428_0, i_10_183_4570_0, i_10_183_4582_0;
  output o_10_183_0_0;
  assign o_10_183_0_0 = 0;
endmodule



// Benchmark "kernel_10_184" written by ABC on Sun Jul 19 10:24:10 2020

module kernel_10_184 ( 
    i_10_184_64_0, i_10_184_180_0, i_10_184_243_0, i_10_184_262_0,
    i_10_184_408_0, i_10_184_424_0, i_10_184_429_0, i_10_184_430_0,
    i_10_184_444_0, i_10_184_445_0, i_10_184_462_0, i_10_184_467_0,
    i_10_184_831_0, i_10_184_921_0, i_10_184_954_0, i_10_184_955_0,
    i_10_184_956_0, i_10_184_957_0, i_10_184_959_0, i_10_184_962_0,
    i_10_184_1002_0, i_10_184_1026_0, i_10_184_1034_0, i_10_184_1080_0,
    i_10_184_1161_0, i_10_184_1162_0, i_10_184_1233_0, i_10_184_1287_0,
    i_10_184_1488_0, i_10_184_1494_0, i_10_184_1533_0, i_10_184_1579_0,
    i_10_184_1614_0, i_10_184_1638_0, i_10_184_1854_0, i_10_184_1872_0,
    i_10_184_1910_0, i_10_184_1914_0, i_10_184_1944_0, i_10_184_1945_0,
    i_10_184_2088_0, i_10_184_2202_0, i_10_184_2304_0, i_10_184_2323_0,
    i_10_184_2349_0, i_10_184_2350_0, i_10_184_2365_0, i_10_184_2376_0,
    i_10_184_2406_0, i_10_184_2409_0, i_10_184_2472_0, i_10_184_2473_0,
    i_10_184_2563_0, i_10_184_2604_0, i_10_184_2629_0, i_10_184_2632_0,
    i_10_184_2657_0, i_10_184_2658_0, i_10_184_2662_0, i_10_184_2676_0,
    i_10_184_2700_0, i_10_184_2705_0, i_10_184_2734_0, i_10_184_2740_0,
    i_10_184_2754_0, i_10_184_2982_0, i_10_184_3034_0, i_10_184_3037_0,
    i_10_184_3070_0, i_10_184_3195_0, i_10_184_3196_0, i_10_184_3283_0,
    i_10_184_3294_0, i_10_184_3312_0, i_10_184_3384_0, i_10_184_3385_0,
    i_10_184_3387_0, i_10_184_3391_0, i_10_184_3432_0, i_10_184_3465_0,
    i_10_184_3469_0, i_10_184_3499_0, i_10_184_3585_0, i_10_184_3609_0,
    i_10_184_3616_0, i_10_184_3645_0, i_10_184_3651_0, i_10_184_3877_0,
    i_10_184_3996_0, i_10_184_4000_0, i_10_184_4113_0, i_10_184_4114_0,
    i_10_184_4115_0, i_10_184_4188_0, i_10_184_4275_0, i_10_184_4287_0,
    i_10_184_4297_0, i_10_184_4369_0, i_10_184_4554_0, i_10_184_4581_0,
    o_10_184_0_0  );
  input  i_10_184_64_0, i_10_184_180_0, i_10_184_243_0, i_10_184_262_0,
    i_10_184_408_0, i_10_184_424_0, i_10_184_429_0, i_10_184_430_0,
    i_10_184_444_0, i_10_184_445_0, i_10_184_462_0, i_10_184_467_0,
    i_10_184_831_0, i_10_184_921_0, i_10_184_954_0, i_10_184_955_0,
    i_10_184_956_0, i_10_184_957_0, i_10_184_959_0, i_10_184_962_0,
    i_10_184_1002_0, i_10_184_1026_0, i_10_184_1034_0, i_10_184_1080_0,
    i_10_184_1161_0, i_10_184_1162_0, i_10_184_1233_0, i_10_184_1287_0,
    i_10_184_1488_0, i_10_184_1494_0, i_10_184_1533_0, i_10_184_1579_0,
    i_10_184_1614_0, i_10_184_1638_0, i_10_184_1854_0, i_10_184_1872_0,
    i_10_184_1910_0, i_10_184_1914_0, i_10_184_1944_0, i_10_184_1945_0,
    i_10_184_2088_0, i_10_184_2202_0, i_10_184_2304_0, i_10_184_2323_0,
    i_10_184_2349_0, i_10_184_2350_0, i_10_184_2365_0, i_10_184_2376_0,
    i_10_184_2406_0, i_10_184_2409_0, i_10_184_2472_0, i_10_184_2473_0,
    i_10_184_2563_0, i_10_184_2604_0, i_10_184_2629_0, i_10_184_2632_0,
    i_10_184_2657_0, i_10_184_2658_0, i_10_184_2662_0, i_10_184_2676_0,
    i_10_184_2700_0, i_10_184_2705_0, i_10_184_2734_0, i_10_184_2740_0,
    i_10_184_2754_0, i_10_184_2982_0, i_10_184_3034_0, i_10_184_3037_0,
    i_10_184_3070_0, i_10_184_3195_0, i_10_184_3196_0, i_10_184_3283_0,
    i_10_184_3294_0, i_10_184_3312_0, i_10_184_3384_0, i_10_184_3385_0,
    i_10_184_3387_0, i_10_184_3391_0, i_10_184_3432_0, i_10_184_3465_0,
    i_10_184_3469_0, i_10_184_3499_0, i_10_184_3585_0, i_10_184_3609_0,
    i_10_184_3616_0, i_10_184_3645_0, i_10_184_3651_0, i_10_184_3877_0,
    i_10_184_3996_0, i_10_184_4000_0, i_10_184_4113_0, i_10_184_4114_0,
    i_10_184_4115_0, i_10_184_4188_0, i_10_184_4275_0, i_10_184_4287_0,
    i_10_184_4297_0, i_10_184_4369_0, i_10_184_4554_0, i_10_184_4581_0;
  output o_10_184_0_0;
  assign o_10_184_0_0 = 0;
endmodule



// Benchmark "kernel_10_185" written by ABC on Sun Jul 19 10:24:11 2020

module kernel_10_185 ( 
    i_10_185_32_0, i_10_185_174_0, i_10_185_223_0, i_10_185_224_0,
    i_10_185_245_0, i_10_185_319_0, i_10_185_320_0, i_10_185_361_0,
    i_10_185_393_0, i_10_185_443_0, i_10_185_460_0, i_10_185_461_0,
    i_10_185_463_0, i_10_185_467_0, i_10_185_499_0, i_10_185_514_0,
    i_10_185_931_0, i_10_185_996_0, i_10_185_999_0, i_10_185_1237_0,
    i_10_185_1245_0, i_10_185_1246_0, i_10_185_1249_0, i_10_185_1297_0,
    i_10_185_1399_0, i_10_185_1432_0, i_10_185_1434_0, i_10_185_1435_0,
    i_10_185_1502_0, i_10_185_1543_0, i_10_185_1580_0, i_10_185_1624_0,
    i_10_185_1625_0, i_10_185_1689_0, i_10_185_1690_0, i_10_185_1807_0,
    i_10_185_1818_0, i_10_185_1819_0, i_10_185_1912_0, i_10_185_1983_0,
    i_10_185_1994_0, i_10_185_1996_0, i_10_185_2003_0, i_10_185_2006_0,
    i_10_185_2337_0, i_10_185_2353_0, i_10_185_2450_0, i_10_185_2474_0,
    i_10_185_2556_0, i_10_185_2629_0, i_10_185_2631_0, i_10_185_2634_0,
    i_10_185_2642_0, i_10_185_2705_0, i_10_185_2731_0, i_10_185_2733_0,
    i_10_185_2734_0, i_10_185_2735_0, i_10_185_2786_0, i_10_185_3041_0,
    i_10_185_3157_0, i_10_185_3284_0, i_10_185_3313_0, i_10_185_3316_0,
    i_10_185_3333_0, i_10_185_3387_0, i_10_185_3434_0, i_10_185_3451_0,
    i_10_185_3470_0, i_10_185_3473_0, i_10_185_3500_0, i_10_185_3525_0,
    i_10_185_3526_0, i_10_185_3543_0, i_10_185_3544_0, i_10_185_3725_0,
    i_10_185_3834_0, i_10_185_3835_0, i_10_185_3838_0, i_10_185_3839_0,
    i_10_185_3841_0, i_10_185_3852_0, i_10_185_3855_0, i_10_185_3883_0,
    i_10_185_3884_0, i_10_185_3895_0, i_10_185_3896_0, i_10_185_3988_0,
    i_10_185_4054_0, i_10_185_4055_0, i_10_185_4115_0, i_10_185_4121_0,
    i_10_185_4207_0, i_10_185_4208_0, i_10_185_4211_0, i_10_185_4282_0,
    i_10_185_4292_0, i_10_185_4588_0, i_10_185_4589_0, i_10_185_4592_0,
    o_10_185_0_0  );
  input  i_10_185_32_0, i_10_185_174_0, i_10_185_223_0, i_10_185_224_0,
    i_10_185_245_0, i_10_185_319_0, i_10_185_320_0, i_10_185_361_0,
    i_10_185_393_0, i_10_185_443_0, i_10_185_460_0, i_10_185_461_0,
    i_10_185_463_0, i_10_185_467_0, i_10_185_499_0, i_10_185_514_0,
    i_10_185_931_0, i_10_185_996_0, i_10_185_999_0, i_10_185_1237_0,
    i_10_185_1245_0, i_10_185_1246_0, i_10_185_1249_0, i_10_185_1297_0,
    i_10_185_1399_0, i_10_185_1432_0, i_10_185_1434_0, i_10_185_1435_0,
    i_10_185_1502_0, i_10_185_1543_0, i_10_185_1580_0, i_10_185_1624_0,
    i_10_185_1625_0, i_10_185_1689_0, i_10_185_1690_0, i_10_185_1807_0,
    i_10_185_1818_0, i_10_185_1819_0, i_10_185_1912_0, i_10_185_1983_0,
    i_10_185_1994_0, i_10_185_1996_0, i_10_185_2003_0, i_10_185_2006_0,
    i_10_185_2337_0, i_10_185_2353_0, i_10_185_2450_0, i_10_185_2474_0,
    i_10_185_2556_0, i_10_185_2629_0, i_10_185_2631_0, i_10_185_2634_0,
    i_10_185_2642_0, i_10_185_2705_0, i_10_185_2731_0, i_10_185_2733_0,
    i_10_185_2734_0, i_10_185_2735_0, i_10_185_2786_0, i_10_185_3041_0,
    i_10_185_3157_0, i_10_185_3284_0, i_10_185_3313_0, i_10_185_3316_0,
    i_10_185_3333_0, i_10_185_3387_0, i_10_185_3434_0, i_10_185_3451_0,
    i_10_185_3470_0, i_10_185_3473_0, i_10_185_3500_0, i_10_185_3525_0,
    i_10_185_3526_0, i_10_185_3543_0, i_10_185_3544_0, i_10_185_3725_0,
    i_10_185_3834_0, i_10_185_3835_0, i_10_185_3838_0, i_10_185_3839_0,
    i_10_185_3841_0, i_10_185_3852_0, i_10_185_3855_0, i_10_185_3883_0,
    i_10_185_3884_0, i_10_185_3895_0, i_10_185_3896_0, i_10_185_3988_0,
    i_10_185_4054_0, i_10_185_4055_0, i_10_185_4115_0, i_10_185_4121_0,
    i_10_185_4207_0, i_10_185_4208_0, i_10_185_4211_0, i_10_185_4282_0,
    i_10_185_4292_0, i_10_185_4588_0, i_10_185_4589_0, i_10_185_4592_0;
  output o_10_185_0_0;
  assign o_10_185_0_0 = 0;
endmodule



// Benchmark "kernel_10_186" written by ABC on Sun Jul 19 10:24:12 2020

module kernel_10_186 ( 
    i_10_186_46_0, i_10_186_47_0, i_10_186_49_0, i_10_186_50_0,
    i_10_186_154_0, i_10_186_179_0, i_10_186_220_0, i_10_186_221_0,
    i_10_186_222_0, i_10_186_280_0, i_10_186_291_0, i_10_186_318_0,
    i_10_186_327_0, i_10_186_328_0, i_10_186_406_0, i_10_186_410_0,
    i_10_186_440_0, i_10_186_445_0, i_10_186_795_0, i_10_186_798_0,
    i_10_186_893_0, i_10_186_1028_0, i_10_186_1037_0, i_10_186_1118_0,
    i_10_186_1121_0, i_10_186_1202_0, i_10_186_1239_0, i_10_186_1242_0,
    i_10_186_1264_0, i_10_186_1266_0, i_10_186_1276_0, i_10_186_1306_0,
    i_10_186_1445_0, i_10_186_1539_0, i_10_186_1653_0, i_10_186_1683_0,
    i_10_186_1685_0, i_10_186_1691_0, i_10_186_1765_0, i_10_186_1767_0,
    i_10_186_1768_0, i_10_186_1769_0, i_10_186_1771_0, i_10_186_1772_0,
    i_10_186_1819_0, i_10_186_1822_0, i_10_186_2201_0, i_10_186_2327_0,
    i_10_186_2361_0, i_10_186_2362_0, i_10_186_2378_0, i_10_186_2381_0,
    i_10_186_2449_0, i_10_186_2460_0, i_10_186_2603_0, i_10_186_2607_0,
    i_10_186_2629_0, i_10_186_2631_0, i_10_186_2635_0, i_10_186_2718_0,
    i_10_186_2723_0, i_10_186_2826_0, i_10_186_2829_0, i_10_186_2831_0,
    i_10_186_2834_0, i_10_186_2917_0, i_10_186_2918_0, i_10_186_2919_0,
    i_10_186_2921_0, i_10_186_2923_0, i_10_186_2924_0, i_10_186_2980_0,
    i_10_186_3048_0, i_10_186_3070_0, i_10_186_3072_0, i_10_186_3091_0,
    i_10_186_3092_0, i_10_186_3283_0, i_10_186_3388_0, i_10_186_3403_0,
    i_10_186_3407_0, i_10_186_3523_0, i_10_186_3551_0, i_10_186_3614_0,
    i_10_186_3809_0, i_10_186_3837_0, i_10_186_3846_0, i_10_186_3850_0,
    i_10_186_3852_0, i_10_186_3853_0, i_10_186_3855_0, i_10_186_3856_0,
    i_10_186_3857_0, i_10_186_4123_0, i_10_186_4284_0, i_10_186_4286_0,
    i_10_186_4288_0, i_10_186_4564_0, i_10_186_4570_0, i_10_186_4571_0,
    o_10_186_0_0  );
  input  i_10_186_46_0, i_10_186_47_0, i_10_186_49_0, i_10_186_50_0,
    i_10_186_154_0, i_10_186_179_0, i_10_186_220_0, i_10_186_221_0,
    i_10_186_222_0, i_10_186_280_0, i_10_186_291_0, i_10_186_318_0,
    i_10_186_327_0, i_10_186_328_0, i_10_186_406_0, i_10_186_410_0,
    i_10_186_440_0, i_10_186_445_0, i_10_186_795_0, i_10_186_798_0,
    i_10_186_893_0, i_10_186_1028_0, i_10_186_1037_0, i_10_186_1118_0,
    i_10_186_1121_0, i_10_186_1202_0, i_10_186_1239_0, i_10_186_1242_0,
    i_10_186_1264_0, i_10_186_1266_0, i_10_186_1276_0, i_10_186_1306_0,
    i_10_186_1445_0, i_10_186_1539_0, i_10_186_1653_0, i_10_186_1683_0,
    i_10_186_1685_0, i_10_186_1691_0, i_10_186_1765_0, i_10_186_1767_0,
    i_10_186_1768_0, i_10_186_1769_0, i_10_186_1771_0, i_10_186_1772_0,
    i_10_186_1819_0, i_10_186_1822_0, i_10_186_2201_0, i_10_186_2327_0,
    i_10_186_2361_0, i_10_186_2362_0, i_10_186_2378_0, i_10_186_2381_0,
    i_10_186_2449_0, i_10_186_2460_0, i_10_186_2603_0, i_10_186_2607_0,
    i_10_186_2629_0, i_10_186_2631_0, i_10_186_2635_0, i_10_186_2718_0,
    i_10_186_2723_0, i_10_186_2826_0, i_10_186_2829_0, i_10_186_2831_0,
    i_10_186_2834_0, i_10_186_2917_0, i_10_186_2918_0, i_10_186_2919_0,
    i_10_186_2921_0, i_10_186_2923_0, i_10_186_2924_0, i_10_186_2980_0,
    i_10_186_3048_0, i_10_186_3070_0, i_10_186_3072_0, i_10_186_3091_0,
    i_10_186_3092_0, i_10_186_3283_0, i_10_186_3388_0, i_10_186_3403_0,
    i_10_186_3407_0, i_10_186_3523_0, i_10_186_3551_0, i_10_186_3614_0,
    i_10_186_3809_0, i_10_186_3837_0, i_10_186_3846_0, i_10_186_3850_0,
    i_10_186_3852_0, i_10_186_3853_0, i_10_186_3855_0, i_10_186_3856_0,
    i_10_186_3857_0, i_10_186_4123_0, i_10_186_4284_0, i_10_186_4286_0,
    i_10_186_4288_0, i_10_186_4564_0, i_10_186_4570_0, i_10_186_4571_0;
  output o_10_186_0_0;
  assign o_10_186_0_0 = 0;
endmodule



// Benchmark "kernel_10_187" written by ABC on Sun Jul 19 10:24:12 2020

module kernel_10_187 ( 
    i_10_187_144_0, i_10_187_147_0, i_10_187_148_0, i_10_187_172_0,
    i_10_187_177_0, i_10_187_222_0, i_10_187_223_0, i_10_187_250_0,
    i_10_187_260_0, i_10_187_266_0, i_10_187_293_0, i_10_187_330_0,
    i_10_187_405_0, i_10_187_408_0, i_10_187_411_0, i_10_187_447_0,
    i_10_187_628_0, i_10_187_629_0, i_10_187_687_0, i_10_187_741_0,
    i_10_187_742_0, i_10_187_745_0, i_10_187_747_0, i_10_187_798_0,
    i_10_187_967_0, i_10_187_970_0, i_10_187_1002_0, i_10_187_1218_0,
    i_10_187_1221_0, i_10_187_1222_0, i_10_187_1236_0, i_10_187_1239_0,
    i_10_187_1240_0, i_10_187_1275_0, i_10_187_1365_0, i_10_187_1434_0,
    i_10_187_1438_0, i_10_187_1444_0, i_10_187_1446_0, i_10_187_1447_0,
    i_10_187_1488_0, i_10_187_1502_0, i_10_187_1821_0, i_10_187_1920_0,
    i_10_187_2001_0, i_10_187_2031_0, i_10_187_2032_0, i_10_187_2037_0,
    i_10_187_2040_0, i_10_187_2110_0, i_10_187_2290_0, i_10_187_2349_0,
    i_10_187_2353_0, i_10_187_2354_0, i_10_187_2383_0, i_10_187_2384_0,
    i_10_187_2406_0, i_10_187_2470_0, i_10_187_2559_0, i_10_187_2608_0,
    i_10_187_2711_0, i_10_187_2715_0, i_10_187_2734_0, i_10_187_2742_0,
    i_10_187_2787_0, i_10_187_2841_0, i_10_187_2847_0, i_10_187_2885_0,
    i_10_187_2960_0, i_10_187_2967_0, i_10_187_3076_0, i_10_187_3077_0,
    i_10_187_3273_0, i_10_187_3283_0, i_10_187_3319_0, i_10_187_3384_0,
    i_10_187_3387_0, i_10_187_3492_0, i_10_187_3504_0, i_10_187_3507_0,
    i_10_187_3508_0, i_10_187_3544_0, i_10_187_3718_0, i_10_187_3721_0,
    i_10_187_3836_0, i_10_187_3840_0, i_10_187_4012_0, i_10_187_4119_0,
    i_10_187_4129_0, i_10_187_4211_0, i_10_187_4220_0, i_10_187_4266_0,
    i_10_187_4269_0, i_10_187_4272_0, i_10_187_4281_0, i_10_187_4292_0,
    i_10_187_4435_0, i_10_187_4564_0, i_10_187_4567_0, i_10_187_4585_0,
    o_10_187_0_0  );
  input  i_10_187_144_0, i_10_187_147_0, i_10_187_148_0, i_10_187_172_0,
    i_10_187_177_0, i_10_187_222_0, i_10_187_223_0, i_10_187_250_0,
    i_10_187_260_0, i_10_187_266_0, i_10_187_293_0, i_10_187_330_0,
    i_10_187_405_0, i_10_187_408_0, i_10_187_411_0, i_10_187_447_0,
    i_10_187_628_0, i_10_187_629_0, i_10_187_687_0, i_10_187_741_0,
    i_10_187_742_0, i_10_187_745_0, i_10_187_747_0, i_10_187_798_0,
    i_10_187_967_0, i_10_187_970_0, i_10_187_1002_0, i_10_187_1218_0,
    i_10_187_1221_0, i_10_187_1222_0, i_10_187_1236_0, i_10_187_1239_0,
    i_10_187_1240_0, i_10_187_1275_0, i_10_187_1365_0, i_10_187_1434_0,
    i_10_187_1438_0, i_10_187_1444_0, i_10_187_1446_0, i_10_187_1447_0,
    i_10_187_1488_0, i_10_187_1502_0, i_10_187_1821_0, i_10_187_1920_0,
    i_10_187_2001_0, i_10_187_2031_0, i_10_187_2032_0, i_10_187_2037_0,
    i_10_187_2040_0, i_10_187_2110_0, i_10_187_2290_0, i_10_187_2349_0,
    i_10_187_2353_0, i_10_187_2354_0, i_10_187_2383_0, i_10_187_2384_0,
    i_10_187_2406_0, i_10_187_2470_0, i_10_187_2559_0, i_10_187_2608_0,
    i_10_187_2711_0, i_10_187_2715_0, i_10_187_2734_0, i_10_187_2742_0,
    i_10_187_2787_0, i_10_187_2841_0, i_10_187_2847_0, i_10_187_2885_0,
    i_10_187_2960_0, i_10_187_2967_0, i_10_187_3076_0, i_10_187_3077_0,
    i_10_187_3273_0, i_10_187_3283_0, i_10_187_3319_0, i_10_187_3384_0,
    i_10_187_3387_0, i_10_187_3492_0, i_10_187_3504_0, i_10_187_3507_0,
    i_10_187_3508_0, i_10_187_3544_0, i_10_187_3718_0, i_10_187_3721_0,
    i_10_187_3836_0, i_10_187_3840_0, i_10_187_4012_0, i_10_187_4119_0,
    i_10_187_4129_0, i_10_187_4211_0, i_10_187_4220_0, i_10_187_4266_0,
    i_10_187_4269_0, i_10_187_4272_0, i_10_187_4281_0, i_10_187_4292_0,
    i_10_187_4435_0, i_10_187_4564_0, i_10_187_4567_0, i_10_187_4585_0;
  output o_10_187_0_0;
  assign o_10_187_0_0 = 0;
endmodule



// Benchmark "kernel_10_188" written by ABC on Sun Jul 19 10:24:14 2020

module kernel_10_188 ( 
    i_10_188_172_0, i_10_188_177_0, i_10_188_183_0, i_10_188_249_0,
    i_10_188_267_0, i_10_188_285_0, i_10_188_286_0, i_10_188_319_0,
    i_10_188_324_0, i_10_188_328_0, i_10_188_408_0, i_10_188_410_0,
    i_10_188_460_0, i_10_188_507_0, i_10_188_753_0, i_10_188_754_0,
    i_10_188_797_0, i_10_188_996_0, i_10_188_1006_0, i_10_188_1041_0,
    i_10_188_1042_0, i_10_188_1309_0, i_10_188_1437_0, i_10_188_1442_0,
    i_10_188_1578_0, i_10_188_1579_0, i_10_188_1654_0, i_10_188_1655_0,
    i_10_188_1684_0, i_10_188_1687_0, i_10_188_1690_0, i_10_188_1815_0,
    i_10_188_1821_0, i_10_188_1823_0, i_10_188_1825_0, i_10_188_1947_0,
    i_10_188_1951_0, i_10_188_1996_0, i_10_188_2019_0, i_10_188_2022_0,
    i_10_188_2349_0, i_10_188_2350_0, i_10_188_2352_0, i_10_188_2353_0,
    i_10_188_2355_0, i_10_188_2451_0, i_10_188_2453_0, i_10_188_2469_0,
    i_10_188_2607_0, i_10_188_2632_0, i_10_188_2633_0, i_10_188_2673_0,
    i_10_188_2703_0, i_10_188_2704_0, i_10_188_2713_0, i_10_188_2715_0,
    i_10_188_2729_0, i_10_188_2734_0, i_10_188_2735_0, i_10_188_2823_0,
    i_10_188_2829_0, i_10_188_2985_0, i_10_188_2986_0, i_10_188_3076_0,
    i_10_188_3270_0, i_10_188_3271_0, i_10_188_3272_0, i_10_188_3274_0,
    i_10_188_3388_0, i_10_188_3391_0, i_10_188_3409_0, i_10_188_3469_0,
    i_10_188_3472_0, i_10_188_3525_0, i_10_188_3582_0, i_10_188_3588_0,
    i_10_188_3589_0, i_10_188_3612_0, i_10_188_3613_0, i_10_188_3780_0,
    i_10_188_3837_0, i_10_188_3841_0, i_10_188_3852_0, i_10_188_3855_0,
    i_10_188_3857_0, i_10_188_3858_0, i_10_188_3894_0, i_10_188_3895_0,
    i_10_188_3990_0, i_10_188_3991_0, i_10_188_4116_0, i_10_188_4127_0,
    i_10_188_4129_0, i_10_188_4267_0, i_10_188_4281_0, i_10_188_4282_0,
    i_10_188_4283_0, i_10_188_4288_0, i_10_188_4290_0, i_10_188_4567_0,
    o_10_188_0_0  );
  input  i_10_188_172_0, i_10_188_177_0, i_10_188_183_0, i_10_188_249_0,
    i_10_188_267_0, i_10_188_285_0, i_10_188_286_0, i_10_188_319_0,
    i_10_188_324_0, i_10_188_328_0, i_10_188_408_0, i_10_188_410_0,
    i_10_188_460_0, i_10_188_507_0, i_10_188_753_0, i_10_188_754_0,
    i_10_188_797_0, i_10_188_996_0, i_10_188_1006_0, i_10_188_1041_0,
    i_10_188_1042_0, i_10_188_1309_0, i_10_188_1437_0, i_10_188_1442_0,
    i_10_188_1578_0, i_10_188_1579_0, i_10_188_1654_0, i_10_188_1655_0,
    i_10_188_1684_0, i_10_188_1687_0, i_10_188_1690_0, i_10_188_1815_0,
    i_10_188_1821_0, i_10_188_1823_0, i_10_188_1825_0, i_10_188_1947_0,
    i_10_188_1951_0, i_10_188_1996_0, i_10_188_2019_0, i_10_188_2022_0,
    i_10_188_2349_0, i_10_188_2350_0, i_10_188_2352_0, i_10_188_2353_0,
    i_10_188_2355_0, i_10_188_2451_0, i_10_188_2453_0, i_10_188_2469_0,
    i_10_188_2607_0, i_10_188_2632_0, i_10_188_2633_0, i_10_188_2673_0,
    i_10_188_2703_0, i_10_188_2704_0, i_10_188_2713_0, i_10_188_2715_0,
    i_10_188_2729_0, i_10_188_2734_0, i_10_188_2735_0, i_10_188_2823_0,
    i_10_188_2829_0, i_10_188_2985_0, i_10_188_2986_0, i_10_188_3076_0,
    i_10_188_3270_0, i_10_188_3271_0, i_10_188_3272_0, i_10_188_3274_0,
    i_10_188_3388_0, i_10_188_3391_0, i_10_188_3409_0, i_10_188_3469_0,
    i_10_188_3472_0, i_10_188_3525_0, i_10_188_3582_0, i_10_188_3588_0,
    i_10_188_3589_0, i_10_188_3612_0, i_10_188_3613_0, i_10_188_3780_0,
    i_10_188_3837_0, i_10_188_3841_0, i_10_188_3852_0, i_10_188_3855_0,
    i_10_188_3857_0, i_10_188_3858_0, i_10_188_3894_0, i_10_188_3895_0,
    i_10_188_3990_0, i_10_188_3991_0, i_10_188_4116_0, i_10_188_4127_0,
    i_10_188_4129_0, i_10_188_4267_0, i_10_188_4281_0, i_10_188_4282_0,
    i_10_188_4283_0, i_10_188_4288_0, i_10_188_4290_0, i_10_188_4567_0;
  output o_10_188_0_0;
  assign o_10_188_0_0 = ~((~i_10_188_1042_0 & ((~i_10_188_797_0 & ~i_10_188_2823_0 & ~i_10_188_3852_0 & ~i_10_188_3895_0 & ~i_10_188_3990_0) | (~i_10_188_172_0 & ~i_10_188_754_0 & ~i_10_188_996_0 & ~i_10_188_1041_0 & ~i_10_188_2607_0 & ~i_10_188_3991_0))) | (~i_10_188_4127_0 & ((~i_10_188_1041_0 & ((~i_10_188_2607_0 & i_10_188_2713_0 & ~i_10_188_2823_0 & ~i_10_188_3271_0 & ~i_10_188_4267_0) | (~i_10_188_285_0 & ~i_10_188_1442_0 & ~i_10_188_2022_0 & i_10_188_2704_0 & ~i_10_188_3589_0 & ~i_10_188_3612_0 & ~i_10_188_3855_0 & ~i_10_188_4283_0))) | (~i_10_188_3895_0 & ((~i_10_188_1309_0 & ~i_10_188_1578_0 & ~i_10_188_2019_0 & ~i_10_188_2453_0 & ~i_10_188_2715_0 & ~i_10_188_3270_0) | (~i_10_188_1815_0 & ~i_10_188_1821_0 & ~i_10_188_4282_0))))) | (~i_10_188_1578_0 & ~i_10_188_3613_0 & ((~i_10_188_319_0 & ~i_10_188_410_0 & ~i_10_188_2633_0 & ~i_10_188_3525_0 & ~i_10_188_4267_0) | (~i_10_188_1821_0 & ~i_10_188_2735_0 & ~i_10_188_4281_0))) | (~i_10_188_410_0 & ((~i_10_188_1815_0 & ~i_10_188_2673_0 & ~i_10_188_2729_0 & ~i_10_188_3894_0 & ~i_10_188_3991_0) | (~i_10_188_1821_0 & ~i_10_188_2703_0 & ~i_10_188_4283_0))) | (~i_10_188_1823_0 & ((~i_10_188_408_0 & ~i_10_188_1947_0 & ~i_10_188_3894_0 & ~i_10_188_3990_0 & ~i_10_188_3991_0 & i_10_188_4116_0) | (~i_10_188_183_0 & ~i_10_188_1687_0 & ~i_10_188_2019_0 & ~i_10_188_2022_0 & ~i_10_188_4282_0))) | (~i_10_188_3895_0 & ((~i_10_188_408_0 & ((~i_10_188_183_0 & ~i_10_188_267_0 & ~i_10_188_1442_0 & ~i_10_188_2022_0 & ~i_10_188_2673_0 & ~i_10_188_2986_0) | (~i_10_188_319_0 & ~i_10_188_460_0 & ~i_10_188_4282_0))) | (i_10_188_1655_0 & i_10_188_4267_0))) | (~i_10_188_183_0 & ((i_10_188_285_0 & ~i_10_188_3894_0 & ~i_10_188_3991_0) | (~i_10_188_319_0 & ~i_10_188_1442_0 & i_10_188_1823_0 & ~i_10_188_3780_0 & ~i_10_188_3990_0 & ~i_10_188_4283_0))) | (i_10_188_328_0 & i_10_188_3841_0) | (~i_10_188_3612_0 & i_10_188_3858_0 & ~i_10_188_3991_0) | (~i_10_188_1442_0 & ~i_10_188_1654_0 & ~i_10_188_1825_0 & ~i_10_188_3852_0 & ~i_10_188_3858_0 & ~i_10_188_3990_0 & ~i_10_188_4129_0) | (~i_10_188_319_0 & ~i_10_188_2673_0 & ~i_10_188_2735_0 & i_10_188_3612_0 & ~i_10_188_3780_0 & ~i_10_188_4116_0 & ~i_10_188_4288_0 & ~i_10_188_4290_0));
endmodule



// Benchmark "kernel_10_189" written by ABC on Sun Jul 19 10:24:15 2020

module kernel_10_189 ( 
    i_10_189_172_0, i_10_189_173_0, i_10_189_219_0, i_10_189_222_0,
    i_10_189_224_0, i_10_189_271_0, i_10_189_279_0, i_10_189_286_0,
    i_10_189_315_0, i_10_189_316_0, i_10_189_318_0, i_10_189_319_0,
    i_10_189_320_0, i_10_189_408_0, i_10_189_442_0, i_10_189_463_0,
    i_10_189_464_0, i_10_189_467_0, i_10_189_716_0, i_10_189_900_0,
    i_10_189_967_0, i_10_189_1084_0, i_10_189_1245_0, i_10_189_1246_0,
    i_10_189_1247_0, i_10_189_1248_0, i_10_189_1249_0, i_10_189_1250_0,
    i_10_189_1305_0, i_10_189_1307_0, i_10_189_1308_0, i_10_189_1311_0,
    i_10_189_1365_0, i_10_189_1651_0, i_10_189_1652_0, i_10_189_1653_0,
    i_10_189_1678_0, i_10_189_1685_0, i_10_189_1687_0, i_10_189_1802_0,
    i_10_189_1822_0, i_10_189_1825_0, i_10_189_1911_0, i_10_189_1912_0,
    i_10_189_1913_0, i_10_189_2198_0, i_10_189_2355_0, i_10_189_2403_0,
    i_10_189_2452_0, i_10_189_2460_0, i_10_189_2506_0, i_10_189_2628_0,
    i_10_189_2629_0, i_10_189_2632_0, i_10_189_2636_0, i_10_189_2701_0,
    i_10_189_2721_0, i_10_189_2722_0, i_10_189_2724_0, i_10_189_2725_0,
    i_10_189_2726_0, i_10_189_2731_0, i_10_189_2782_0, i_10_189_2828_0,
    i_10_189_2829_0, i_10_189_2833_0, i_10_189_2916_0, i_10_189_2919_0,
    i_10_189_2920_0, i_10_189_2922_0, i_10_189_2923_0, i_10_189_3034_0,
    i_10_189_3163_0, i_10_189_3195_0, i_10_189_3284_0, i_10_189_3323_0,
    i_10_189_3325_0, i_10_189_3390_0, i_10_189_3391_0, i_10_189_3402_0,
    i_10_189_3403_0, i_10_189_3586_0, i_10_189_3855_0, i_10_189_3856_0,
    i_10_189_3858_0, i_10_189_3860_0, i_10_189_3979_0, i_10_189_3980_0,
    i_10_189_3982_0, i_10_189_3983_0, i_10_189_3986_0, i_10_189_4117_0,
    i_10_189_4279_0, i_10_189_4285_0, i_10_189_4286_0, i_10_189_4287_0,
    i_10_189_4288_0, i_10_189_4290_0, i_10_189_4291_0, i_10_189_4566_0,
    o_10_189_0_0  );
  input  i_10_189_172_0, i_10_189_173_0, i_10_189_219_0, i_10_189_222_0,
    i_10_189_224_0, i_10_189_271_0, i_10_189_279_0, i_10_189_286_0,
    i_10_189_315_0, i_10_189_316_0, i_10_189_318_0, i_10_189_319_0,
    i_10_189_320_0, i_10_189_408_0, i_10_189_442_0, i_10_189_463_0,
    i_10_189_464_0, i_10_189_467_0, i_10_189_716_0, i_10_189_900_0,
    i_10_189_967_0, i_10_189_1084_0, i_10_189_1245_0, i_10_189_1246_0,
    i_10_189_1247_0, i_10_189_1248_0, i_10_189_1249_0, i_10_189_1250_0,
    i_10_189_1305_0, i_10_189_1307_0, i_10_189_1308_0, i_10_189_1311_0,
    i_10_189_1365_0, i_10_189_1651_0, i_10_189_1652_0, i_10_189_1653_0,
    i_10_189_1678_0, i_10_189_1685_0, i_10_189_1687_0, i_10_189_1802_0,
    i_10_189_1822_0, i_10_189_1825_0, i_10_189_1911_0, i_10_189_1912_0,
    i_10_189_1913_0, i_10_189_2198_0, i_10_189_2355_0, i_10_189_2403_0,
    i_10_189_2452_0, i_10_189_2460_0, i_10_189_2506_0, i_10_189_2628_0,
    i_10_189_2629_0, i_10_189_2632_0, i_10_189_2636_0, i_10_189_2701_0,
    i_10_189_2721_0, i_10_189_2722_0, i_10_189_2724_0, i_10_189_2725_0,
    i_10_189_2726_0, i_10_189_2731_0, i_10_189_2782_0, i_10_189_2828_0,
    i_10_189_2829_0, i_10_189_2833_0, i_10_189_2916_0, i_10_189_2919_0,
    i_10_189_2920_0, i_10_189_2922_0, i_10_189_2923_0, i_10_189_3034_0,
    i_10_189_3163_0, i_10_189_3195_0, i_10_189_3284_0, i_10_189_3323_0,
    i_10_189_3325_0, i_10_189_3390_0, i_10_189_3391_0, i_10_189_3402_0,
    i_10_189_3403_0, i_10_189_3586_0, i_10_189_3855_0, i_10_189_3856_0,
    i_10_189_3858_0, i_10_189_3860_0, i_10_189_3979_0, i_10_189_3980_0,
    i_10_189_3982_0, i_10_189_3983_0, i_10_189_3986_0, i_10_189_4117_0,
    i_10_189_4279_0, i_10_189_4285_0, i_10_189_4286_0, i_10_189_4287_0,
    i_10_189_4288_0, i_10_189_4290_0, i_10_189_4291_0, i_10_189_4566_0;
  output o_10_189_0_0;
  assign o_10_189_0_0 = ~((~i_10_189_4286_0 & ((~i_10_189_408_0 & ((~i_10_189_172_0 & ~i_10_189_224_0 & ~i_10_189_900_0 & ~i_10_189_1685_0 & ~i_10_189_1822_0 & ~i_10_189_2724_0 & ~i_10_189_2725_0 & ~i_10_189_2920_0) | (~i_10_189_467_0 & ~i_10_189_3284_0 & ~i_10_189_3403_0 & ~i_10_189_3586_0 & ~i_10_189_3856_0 & ~i_10_189_4290_0))) | (~i_10_189_1249_0 & ~i_10_189_1911_0 & ((~i_10_189_173_0 & ~i_10_189_1248_0 & ~i_10_189_2922_0 & ~i_10_189_3858_0 & i_10_189_4288_0 & i_10_189_4291_0) | (~i_10_189_1246_0 & ~i_10_189_2724_0 & ~i_10_189_4285_0 & ~i_10_189_4291_0))) | (~i_10_189_4290_0 & ((~i_10_189_219_0 & ~i_10_189_464_0 & ~i_10_189_467_0 & ~i_10_189_2629_0 & ~i_10_189_2632_0 & ~i_10_189_2922_0 & ~i_10_189_3195_0) | (~i_10_189_1250_0 & ~i_10_189_2726_0 & ~i_10_189_2829_0 & ~i_10_189_3586_0 & ~i_10_189_3855_0 & ~i_10_189_4285_0))))) | (~i_10_189_172_0 & ((i_10_189_463_0 & ~i_10_189_1245_0 & ~i_10_189_1250_0 & ~i_10_189_1365_0 & ~i_10_189_2726_0 & i_10_189_2731_0 & ~i_10_189_3860_0 & ~i_10_189_4285_0) | (~i_10_189_716_0 & i_10_189_1913_0 & ~i_10_189_2721_0 & ~i_10_189_2725_0 & ~i_10_189_3855_0 & ~i_10_189_4291_0))) | (~i_10_189_1247_0 & ((~i_10_189_219_0 & ((~i_10_189_900_0 & ~i_10_189_1249_0 & ~i_10_189_1250_0 & ~i_10_189_1307_0 & ~i_10_189_3855_0 & ~i_10_189_3856_0 & ~i_10_189_4285_0) | (~i_10_189_716_0 & ~i_10_189_967_0 & ~i_10_189_1685_0 & ~i_10_189_2460_0 & ~i_10_189_2923_0 & ~i_10_189_3391_0 & ~i_10_189_4287_0))) | (~i_10_189_467_0 & ((~i_10_189_222_0 & ~i_10_189_716_0 & ~i_10_189_2628_0 & ~i_10_189_2724_0 & ~i_10_189_2731_0 & ~i_10_189_2833_0 & ~i_10_189_3403_0) | (~i_10_189_1246_0 & ~i_10_189_1685_0 & i_10_189_1822_0 & ~i_10_189_2452_0 & ~i_10_189_2721_0 & ~i_10_189_4290_0))) | (~i_10_189_1911_0 & ~i_10_189_3860_0 & ((~i_10_189_442_0 & ~i_10_189_1653_0 & i_10_189_1822_0 & ~i_10_189_1913_0 & ~i_10_189_2916_0 & ~i_10_189_3034_0 & ~i_10_189_3390_0 & ~i_10_189_3586_0 & ~i_10_189_3979_0) | (~i_10_189_716_0 & ~i_10_189_1249_0 & ~i_10_189_1307_0 & ~i_10_189_2460_0 & ~i_10_189_2722_0 & ~i_10_189_4288_0))))) | (~i_10_189_1245_0 & ((~i_10_189_224_0 & ~i_10_189_1913_0 & ((~i_10_189_1250_0 & ~i_10_189_1912_0 & ~i_10_189_2452_0 & ~i_10_189_2721_0 & ~i_10_189_2833_0 & ~i_10_189_2916_0) | (~i_10_189_173_0 & ~i_10_189_2922_0 & ~i_10_189_3403_0 & ~i_10_189_3586_0 & ~i_10_189_4285_0 & ~i_10_189_4290_0))) | (~i_10_189_442_0 & ~i_10_189_2829_0 & ~i_10_189_2920_0 & ~i_10_189_2923_0 & ~i_10_189_4288_0))) | (~i_10_189_464_0 & ~i_10_189_4291_0 & (i_10_189_316_0 | (~i_10_189_716_0 & ~i_10_189_2628_0 & ~i_10_189_2636_0 & ~i_10_189_3858_0 & ~i_10_189_4287_0))) | (~i_10_189_173_0 & ((~i_10_189_967_0 & ((~i_10_189_1311_0 & ~i_10_189_1365_0 & ~i_10_189_2198_0 & ~i_10_189_2460_0 & ~i_10_189_3856_0 & ~i_10_189_4285_0 & ~i_10_189_2721_0 & ~i_10_189_2833_0) | (~i_10_189_1246_0 & ~i_10_189_2452_0 & ~i_10_189_2829_0 & ~i_10_189_3391_0 & ~i_10_189_4290_0))) | (~i_10_189_2460_0 & ~i_10_189_2725_0 & ~i_10_189_2920_0 & ~i_10_189_3855_0 & i_10_189_4286_0))) | (~i_10_189_900_0 & ((~i_10_189_1249_0 & ~i_10_189_2833_0 & ((~i_10_189_1687_0 & i_10_189_2828_0 & ~i_10_189_2919_0 & ~i_10_189_3858_0) | (i_10_189_279_0 & ~i_10_189_2460_0 & ~i_10_189_2726_0 & ~i_10_189_3390_0 & ~i_10_189_3856_0 & i_10_189_4287_0))) | (~i_10_189_442_0 & ~i_10_189_1653_0 & ~i_10_189_1685_0 & ~i_10_189_2721_0 & ~i_10_189_2922_0 & ~i_10_189_3856_0 & ~i_10_189_4290_0 & ~i_10_189_4566_0))) | (~i_10_189_1250_0 & ((~i_10_189_1913_0 & ~i_10_189_2629_0 & ~i_10_189_2632_0 & ~i_10_189_2919_0 & ~i_10_189_3391_0 & ~i_10_189_3860_0) | (~i_10_189_1653_0 & ~i_10_189_2628_0 & ~i_10_189_2722_0 & ~i_10_189_4290_0 & ~i_10_189_4566_0))) | (~i_10_189_2923_0 & ((i_10_189_315_0 & ~i_10_189_2916_0) | (~i_10_189_716_0 & i_10_189_1305_0 & ~i_10_189_3403_0 & ~i_10_189_4285_0 & ~i_10_189_4287_0))) | (~i_10_189_4288_0 & ((~i_10_189_1365_0 & ~i_10_189_1912_0 & ~i_10_189_2628_0 & ~i_10_189_2629_0 & ~i_10_189_2725_0 & ~i_10_189_2829_0 & ~i_10_189_3391_0) | (i_10_189_2833_0 & ~i_10_189_3855_0 & i_10_189_4290_0))) | (i_10_189_319_0 & ~i_10_189_463_0));
endmodule



// Benchmark "kernel_10_190" written by ABC on Sun Jul 19 10:24:16 2020

module kernel_10_190 ( 
    i_10_190_14_0, i_10_190_49_0, i_10_190_86_0, i_10_190_176_0,
    i_10_190_179_0, i_10_190_221_0, i_10_190_254_0, i_10_190_283_0,
    i_10_190_287_0, i_10_190_317_0, i_10_190_391_0, i_10_190_464_0,
    i_10_190_509_0, i_10_190_689_0, i_10_190_869_0, i_10_190_1084_0,
    i_10_190_1085_0, i_10_190_1088_0, i_10_190_1103_0, i_10_190_1235_0,
    i_10_190_1237_0, i_10_190_1238_0, i_10_190_1271_0, i_10_190_1298_0,
    i_10_190_1301_0, i_10_190_1439_0, i_10_190_1454_0, i_10_190_1541_0,
    i_10_190_1544_0, i_10_190_1583_0, i_10_190_1622_0, i_10_190_1648_0,
    i_10_190_1651_0, i_10_190_1684_0, i_10_190_1685_0, i_10_190_1687_0,
    i_10_190_1688_0, i_10_190_1981_0, i_10_190_1982_0, i_10_190_1990_0,
    i_10_190_1994_0, i_10_190_2003_0, i_10_190_2020_0, i_10_190_2021_0,
    i_10_190_2030_0, i_10_190_2189_0, i_10_190_2201_0, i_10_190_2204_0,
    i_10_190_2351_0, i_10_190_2356_0, i_10_190_2465_0, i_10_190_2468_0,
    i_10_190_2471_0, i_10_190_2473_0, i_10_190_2479_0, i_10_190_2567_0,
    i_10_190_2629_0, i_10_190_2636_0, i_10_190_2650_0, i_10_190_2651_0,
    i_10_190_2654_0, i_10_190_2660_0, i_10_190_2711_0, i_10_190_2714_0,
    i_10_190_2821_0, i_10_190_2830_0, i_10_190_2831_0, i_10_190_2846_0,
    i_10_190_2917_0, i_10_190_2919_0, i_10_190_2924_0, i_10_190_2966_0,
    i_10_190_2969_0, i_10_190_3043_0, i_10_190_3070_0, i_10_190_3073_0,
    i_10_190_3088_0, i_10_190_3197_0, i_10_190_3323_0, i_10_190_3391_0,
    i_10_190_3503_0, i_10_190_3526_0, i_10_190_3584_0, i_10_190_3733_0,
    i_10_190_3734_0, i_10_190_3786_0, i_10_190_3794_0, i_10_190_3835_0,
    i_10_190_3847_0, i_10_190_3979_0, i_10_190_4028_0, i_10_190_4126_0,
    i_10_190_4127_0, i_10_190_4130_0, i_10_190_4154_0, i_10_190_4172_0,
    i_10_190_4175_0, i_10_190_4279_0, i_10_190_4291_0, i_10_190_4565_0,
    o_10_190_0_0  );
  input  i_10_190_14_0, i_10_190_49_0, i_10_190_86_0, i_10_190_176_0,
    i_10_190_179_0, i_10_190_221_0, i_10_190_254_0, i_10_190_283_0,
    i_10_190_287_0, i_10_190_317_0, i_10_190_391_0, i_10_190_464_0,
    i_10_190_509_0, i_10_190_689_0, i_10_190_869_0, i_10_190_1084_0,
    i_10_190_1085_0, i_10_190_1088_0, i_10_190_1103_0, i_10_190_1235_0,
    i_10_190_1237_0, i_10_190_1238_0, i_10_190_1271_0, i_10_190_1298_0,
    i_10_190_1301_0, i_10_190_1439_0, i_10_190_1454_0, i_10_190_1541_0,
    i_10_190_1544_0, i_10_190_1583_0, i_10_190_1622_0, i_10_190_1648_0,
    i_10_190_1651_0, i_10_190_1684_0, i_10_190_1685_0, i_10_190_1687_0,
    i_10_190_1688_0, i_10_190_1981_0, i_10_190_1982_0, i_10_190_1990_0,
    i_10_190_1994_0, i_10_190_2003_0, i_10_190_2020_0, i_10_190_2021_0,
    i_10_190_2030_0, i_10_190_2189_0, i_10_190_2201_0, i_10_190_2204_0,
    i_10_190_2351_0, i_10_190_2356_0, i_10_190_2465_0, i_10_190_2468_0,
    i_10_190_2471_0, i_10_190_2473_0, i_10_190_2479_0, i_10_190_2567_0,
    i_10_190_2629_0, i_10_190_2636_0, i_10_190_2650_0, i_10_190_2651_0,
    i_10_190_2654_0, i_10_190_2660_0, i_10_190_2711_0, i_10_190_2714_0,
    i_10_190_2821_0, i_10_190_2830_0, i_10_190_2831_0, i_10_190_2846_0,
    i_10_190_2917_0, i_10_190_2919_0, i_10_190_2924_0, i_10_190_2966_0,
    i_10_190_2969_0, i_10_190_3043_0, i_10_190_3070_0, i_10_190_3073_0,
    i_10_190_3088_0, i_10_190_3197_0, i_10_190_3323_0, i_10_190_3391_0,
    i_10_190_3503_0, i_10_190_3526_0, i_10_190_3584_0, i_10_190_3733_0,
    i_10_190_3734_0, i_10_190_3786_0, i_10_190_3794_0, i_10_190_3835_0,
    i_10_190_3847_0, i_10_190_3979_0, i_10_190_4028_0, i_10_190_4126_0,
    i_10_190_4127_0, i_10_190_4130_0, i_10_190_4154_0, i_10_190_4172_0,
    i_10_190_4175_0, i_10_190_4279_0, i_10_190_4291_0, i_10_190_4565_0;
  output o_10_190_0_0;
  assign o_10_190_0_0 = 0;
endmodule



// Benchmark "kernel_10_191" written by ABC on Sun Jul 19 10:24:18 2020

module kernel_10_191 ( 
    i_10_191_87_0, i_10_191_152_0, i_10_191_172_0, i_10_191_176_0,
    i_10_191_221_0, i_10_191_224_0, i_10_191_259_0, i_10_191_260_0,
    i_10_191_325_0, i_10_191_433_0, i_10_191_443_0, i_10_191_445_0,
    i_10_191_446_0, i_10_191_448_0, i_10_191_449_0, i_10_191_454_0,
    i_10_191_461_0, i_10_191_463_0, i_10_191_467_0, i_10_191_716_0,
    i_10_191_794_0, i_10_191_797_0, i_10_191_800_0, i_10_191_899_0,
    i_10_191_904_0, i_10_191_905_0, i_10_191_908_0, i_10_191_965_0,
    i_10_191_971_0, i_10_191_999_0, i_10_191_1000_0, i_10_191_1135_0,
    i_10_191_1165_0, i_10_191_1166_0, i_10_191_1237_0, i_10_191_1240_0,
    i_10_191_1244_0, i_10_191_1245_0, i_10_191_1246_0, i_10_191_1247_0,
    i_10_191_1248_0, i_10_191_1308_0, i_10_191_1311_0, i_10_191_1553_0,
    i_10_191_1818_0, i_10_191_1822_0, i_10_191_1823_0, i_10_191_2181_0,
    i_10_191_2249_0, i_10_191_2309_0, i_10_191_2335_0, i_10_191_2355_0,
    i_10_191_2410_0, i_10_191_2450_0, i_10_191_2453_0, i_10_191_2470_0,
    i_10_191_2630_0, i_10_191_2635_0, i_10_191_2662_0, i_10_191_2663_0,
    i_10_191_2700_0, i_10_191_2713_0, i_10_191_2720_0, i_10_191_2728_0,
    i_10_191_2729_0, i_10_191_2731_0, i_10_191_2735_0, i_10_191_2785_0,
    i_10_191_2824_0, i_10_191_2881_0, i_10_191_2884_0, i_10_191_2917_0,
    i_10_191_2919_0, i_10_191_2920_0, i_10_191_3038_0, i_10_191_3073_0,
    i_10_191_3274_0, i_10_191_3334_0, i_10_191_3387_0, i_10_191_3391_0,
    i_10_191_3493_0, i_10_191_3494_0, i_10_191_3541_0, i_10_191_3649_0,
    i_10_191_3788_0, i_10_191_3836_0, i_10_191_3858_0, i_10_191_3859_0,
    i_10_191_3986_0, i_10_191_4120_0, i_10_191_4121_0, i_10_191_4220_0,
    i_10_191_4270_0, i_10_191_4271_0, i_10_191_4274_0, i_10_191_4291_0,
    i_10_191_4292_0, i_10_191_4564_0, i_10_191_4565_0, i_10_191_4571_0,
    o_10_191_0_0  );
  input  i_10_191_87_0, i_10_191_152_0, i_10_191_172_0, i_10_191_176_0,
    i_10_191_221_0, i_10_191_224_0, i_10_191_259_0, i_10_191_260_0,
    i_10_191_325_0, i_10_191_433_0, i_10_191_443_0, i_10_191_445_0,
    i_10_191_446_0, i_10_191_448_0, i_10_191_449_0, i_10_191_454_0,
    i_10_191_461_0, i_10_191_463_0, i_10_191_467_0, i_10_191_716_0,
    i_10_191_794_0, i_10_191_797_0, i_10_191_800_0, i_10_191_899_0,
    i_10_191_904_0, i_10_191_905_0, i_10_191_908_0, i_10_191_965_0,
    i_10_191_971_0, i_10_191_999_0, i_10_191_1000_0, i_10_191_1135_0,
    i_10_191_1165_0, i_10_191_1166_0, i_10_191_1237_0, i_10_191_1240_0,
    i_10_191_1244_0, i_10_191_1245_0, i_10_191_1246_0, i_10_191_1247_0,
    i_10_191_1248_0, i_10_191_1308_0, i_10_191_1311_0, i_10_191_1553_0,
    i_10_191_1818_0, i_10_191_1822_0, i_10_191_1823_0, i_10_191_2181_0,
    i_10_191_2249_0, i_10_191_2309_0, i_10_191_2335_0, i_10_191_2355_0,
    i_10_191_2410_0, i_10_191_2450_0, i_10_191_2453_0, i_10_191_2470_0,
    i_10_191_2630_0, i_10_191_2635_0, i_10_191_2662_0, i_10_191_2663_0,
    i_10_191_2700_0, i_10_191_2713_0, i_10_191_2720_0, i_10_191_2728_0,
    i_10_191_2729_0, i_10_191_2731_0, i_10_191_2735_0, i_10_191_2785_0,
    i_10_191_2824_0, i_10_191_2881_0, i_10_191_2884_0, i_10_191_2917_0,
    i_10_191_2919_0, i_10_191_2920_0, i_10_191_3038_0, i_10_191_3073_0,
    i_10_191_3274_0, i_10_191_3334_0, i_10_191_3387_0, i_10_191_3391_0,
    i_10_191_3493_0, i_10_191_3494_0, i_10_191_3541_0, i_10_191_3649_0,
    i_10_191_3788_0, i_10_191_3836_0, i_10_191_3858_0, i_10_191_3859_0,
    i_10_191_3986_0, i_10_191_4120_0, i_10_191_4121_0, i_10_191_4220_0,
    i_10_191_4270_0, i_10_191_4271_0, i_10_191_4274_0, i_10_191_4291_0,
    i_10_191_4292_0, i_10_191_4564_0, i_10_191_4565_0, i_10_191_4571_0;
  output o_10_191_0_0;
  assign o_10_191_0_0 = ~((~i_10_191_1247_0 & ((~i_10_191_152_0 & ((~i_10_191_904_0 & ~i_10_191_2635_0 & ~i_10_191_2720_0 & ~i_10_191_3858_0) | (~i_10_191_899_0 & ~i_10_191_1244_0 & ~i_10_191_1308_0 & ~i_10_191_2450_0 & ~i_10_191_3836_0 & ~i_10_191_4271_0 & ~i_10_191_4565_0))) | (~i_10_191_224_0 & ~i_10_191_1240_0 & ~i_10_191_1246_0 & ~i_10_191_3858_0 & ~i_10_191_4121_0) | (~i_10_191_176_0 & ~i_10_191_908_0 & ~i_10_191_1553_0 & ~i_10_191_2335_0 & ~i_10_191_2720_0 & ~i_10_191_2919_0 & i_10_191_4571_0))) | (~i_10_191_176_0 & ((~i_10_191_172_0 & ~i_10_191_1165_0 & ~i_10_191_2720_0 & ~i_10_191_2881_0 & ~i_10_191_3858_0 & ~i_10_191_4271_0) | (~i_10_191_899_0 & ~i_10_191_1166_0 & ~i_10_191_2729_0 & ~i_10_191_3073_0 & ~i_10_191_4571_0))) | (~i_10_191_908_0 & ((~i_10_191_87_0 & ((~i_10_191_446_0 & ~i_10_191_1818_0 & ~i_10_191_2735_0 & ~i_10_191_4120_0) | (~i_10_191_965_0 & ~i_10_191_971_0 & ~i_10_191_1244_0 & ~i_10_191_2713_0 & ~i_10_191_4291_0))) | (~i_10_191_965_0 & ~i_10_191_2728_0 & ~i_10_191_2735_0 & ~i_10_191_2919_0) | (~i_10_191_1165_0 & ~i_10_191_1166_0 & ~i_10_191_2450_0 & ~i_10_191_2662_0 & ~i_10_191_3859_0))) | (~i_10_191_1166_0 & ((~i_10_191_1822_0 & ~i_10_191_4220_0 & ((~i_10_191_87_0 & ~i_10_191_224_0) | (i_10_191_2720_0 & ~i_10_191_3387_0 & ~i_10_191_3649_0 & ~i_10_191_4120_0))) | (~i_10_191_2919_0 & ((~i_10_191_461_0 & ~i_10_191_463_0) | (~i_10_191_1823_0 & i_10_191_2450_0 & ~i_10_191_2720_0 & ~i_10_191_4564_0))))) | (~i_10_191_2663_0 & i_10_191_2881_0) | (~i_10_191_448_0 & ~i_10_191_899_0 & ~i_10_191_904_0 & i_10_191_2635_0 & ~i_10_191_2713_0 & ~i_10_191_3494_0) | (~i_10_191_1248_0 & ~i_10_191_1823_0 & ~i_10_191_2450_0 & i_10_191_2662_0 & ~i_10_191_2735_0 & ~i_10_191_2824_0 & ~i_10_191_4121_0));
endmodule



// Benchmark "kernel_10_192" written by ABC on Sun Jul 19 10:24:19 2020

module kernel_10_192 ( 
    i_10_192_217_0, i_10_192_223_0, i_10_192_224_0, i_10_192_245_0,
    i_10_192_280_0, i_10_192_281_0, i_10_192_283_0, i_10_192_284_0,
    i_10_192_316_0, i_10_192_318_0, i_10_192_319_0, i_10_192_413_0,
    i_10_192_435_0, i_10_192_443_0, i_10_192_460_0, i_10_192_748_0,
    i_10_192_749_0, i_10_192_792_0, i_10_192_793_0, i_10_192_795_0,
    i_10_192_898_0, i_10_192_956_0, i_10_192_1026_0, i_10_192_1027_0,
    i_10_192_1028_0, i_10_192_1033_0, i_10_192_1137_0, i_10_192_1139_0,
    i_10_192_1233_0, i_10_192_1234_0, i_10_192_1243_0, i_10_192_1539_0,
    i_10_192_1541_0, i_10_192_1549_0, i_10_192_1651_0, i_10_192_1654_0,
    i_10_192_1683_0, i_10_192_1684_0, i_10_192_1685_0, i_10_192_1686_0,
    i_10_192_1687_0, i_10_192_1688_0, i_10_192_1689_0, i_10_192_1691_0,
    i_10_192_1818_0, i_10_192_1819_0, i_10_192_1820_0, i_10_192_1821_0,
    i_10_192_1826_0, i_10_192_1913_0, i_10_192_2180_0, i_10_192_2243_0,
    i_10_192_2352_0, i_10_192_2358_0, i_10_192_2452_0, i_10_192_2470_0,
    i_10_192_2628_0, i_10_192_2631_0, i_10_192_2674_0, i_10_192_2675_0,
    i_10_192_2677_0, i_10_192_2701_0, i_10_192_2702_0, i_10_192_2710_0,
    i_10_192_2718_0, i_10_192_2728_0, i_10_192_2983_0, i_10_192_3073_0,
    i_10_192_3195_0, i_10_192_3198_0, i_10_192_3199_0, i_10_192_3203_0,
    i_10_192_3322_0, i_10_192_3407_0, i_10_192_3408_0, i_10_192_3409_0,
    i_10_192_3519_0, i_10_192_3585_0, i_10_192_3588_0, i_10_192_3589_0,
    i_10_192_3609_0, i_10_192_3610_0, i_10_192_3612_0, i_10_192_3614_0,
    i_10_192_3781_0, i_10_192_3784_0, i_10_192_3785_0, i_10_192_3786_0,
    i_10_192_3787_0, i_10_192_3837_0, i_10_192_3855_0, i_10_192_3856_0,
    i_10_192_3857_0, i_10_192_3979_0, i_10_192_3980_0, i_10_192_3987_0,
    i_10_192_4113_0, i_10_192_4287_0, i_10_192_4567_0, i_10_192_4568_0,
    o_10_192_0_0  );
  input  i_10_192_217_0, i_10_192_223_0, i_10_192_224_0, i_10_192_245_0,
    i_10_192_280_0, i_10_192_281_0, i_10_192_283_0, i_10_192_284_0,
    i_10_192_316_0, i_10_192_318_0, i_10_192_319_0, i_10_192_413_0,
    i_10_192_435_0, i_10_192_443_0, i_10_192_460_0, i_10_192_748_0,
    i_10_192_749_0, i_10_192_792_0, i_10_192_793_0, i_10_192_795_0,
    i_10_192_898_0, i_10_192_956_0, i_10_192_1026_0, i_10_192_1027_0,
    i_10_192_1028_0, i_10_192_1033_0, i_10_192_1137_0, i_10_192_1139_0,
    i_10_192_1233_0, i_10_192_1234_0, i_10_192_1243_0, i_10_192_1539_0,
    i_10_192_1541_0, i_10_192_1549_0, i_10_192_1651_0, i_10_192_1654_0,
    i_10_192_1683_0, i_10_192_1684_0, i_10_192_1685_0, i_10_192_1686_0,
    i_10_192_1687_0, i_10_192_1688_0, i_10_192_1689_0, i_10_192_1691_0,
    i_10_192_1818_0, i_10_192_1819_0, i_10_192_1820_0, i_10_192_1821_0,
    i_10_192_1826_0, i_10_192_1913_0, i_10_192_2180_0, i_10_192_2243_0,
    i_10_192_2352_0, i_10_192_2358_0, i_10_192_2452_0, i_10_192_2470_0,
    i_10_192_2628_0, i_10_192_2631_0, i_10_192_2674_0, i_10_192_2675_0,
    i_10_192_2677_0, i_10_192_2701_0, i_10_192_2702_0, i_10_192_2710_0,
    i_10_192_2718_0, i_10_192_2728_0, i_10_192_2983_0, i_10_192_3073_0,
    i_10_192_3195_0, i_10_192_3198_0, i_10_192_3199_0, i_10_192_3203_0,
    i_10_192_3322_0, i_10_192_3407_0, i_10_192_3408_0, i_10_192_3409_0,
    i_10_192_3519_0, i_10_192_3585_0, i_10_192_3588_0, i_10_192_3589_0,
    i_10_192_3609_0, i_10_192_3610_0, i_10_192_3612_0, i_10_192_3614_0,
    i_10_192_3781_0, i_10_192_3784_0, i_10_192_3785_0, i_10_192_3786_0,
    i_10_192_3787_0, i_10_192_3837_0, i_10_192_3855_0, i_10_192_3856_0,
    i_10_192_3857_0, i_10_192_3979_0, i_10_192_3980_0, i_10_192_3987_0,
    i_10_192_4113_0, i_10_192_4287_0, i_10_192_4567_0, i_10_192_4568_0;
  output o_10_192_0_0;
  assign o_10_192_0_0 = ~((~i_10_192_224_0 & ((~i_10_192_245_0 & ~i_10_192_1685_0 & ~i_10_192_3408_0 & ~i_10_192_3786_0 & ~i_10_192_3855_0) | (~i_10_192_413_0 & ~i_10_192_956_0 & ~i_10_192_1243_0 & ~i_10_192_1651_0 & ~i_10_192_3837_0 & ~i_10_192_4567_0))) | (~i_10_192_413_0 & ((~i_10_192_223_0 & ~i_10_192_1539_0 & ~i_10_192_1688_0 & ~i_10_192_1689_0 & ~i_10_192_2452_0 & ~i_10_192_3409_0 & ~i_10_192_3614_0) | (~i_10_192_749_0 & ~i_10_192_898_0 & ~i_10_192_1654_0 & i_10_192_1821_0 & ~i_10_192_1826_0 & ~i_10_192_2628_0 & ~i_10_192_3589_0 & ~i_10_192_3787_0 & ~i_10_192_3980_0 & ~i_10_192_4568_0))) | (~i_10_192_956_0 & ((~i_10_192_898_0 & ~i_10_192_3073_0 & i_10_192_3610_0) | (~i_10_192_795_0 & i_10_192_1243_0 & ~i_10_192_2180_0 & ~i_10_192_2631_0 & ~i_10_192_3610_0 & i_10_192_3857_0))) | (~i_10_192_1539_0 & ((~i_10_192_1028_0 & i_10_192_1684_0 & ~i_10_192_3612_0) | (~i_10_192_795_0 & ~i_10_192_1687_0 & ~i_10_192_1691_0 & ~i_10_192_3857_0 & ~i_10_192_4287_0))) | (~i_10_192_795_0 & ((~i_10_192_2452_0 & ~i_10_192_2631_0 & ~i_10_192_3781_0 & ~i_10_192_3785_0) | (~i_10_192_223_0 & ~i_10_192_748_0 & ~i_10_192_1028_0 & ~i_10_192_1691_0 & ~i_10_192_1826_0 & ~i_10_192_3203_0 & ~i_10_192_3408_0 & ~i_10_192_4568_0))) | (~i_10_192_898_0 & ((~i_10_192_1028_0 & ((~i_10_192_435_0 & ~i_10_192_1027_0 & ~i_10_192_1685_0 & i_10_192_2631_0 & ~i_10_192_2728_0 & ~i_10_192_3588_0 & i_10_192_3785_0) | (~i_10_192_3408_0 & ~i_10_192_3855_0 & ~i_10_192_3857_0))) | (~i_10_192_749_0 & ~i_10_192_3199_0 & ~i_10_192_3614_0) | (~i_10_192_1243_0 & i_10_192_2631_0 & ~i_10_192_2718_0 & ~i_10_192_3195_0 & ~i_10_192_3785_0 & ~i_10_192_3855_0))) | (~i_10_192_1826_0 & ((~i_10_192_223_0 & i_10_192_1651_0 & ~i_10_192_2180_0 & ~i_10_192_3198_0 & ~i_10_192_3407_0) | (~i_10_192_1651_0 & ~i_10_192_1689_0 & ~i_10_192_1821_0 & ~i_10_192_3408_0 & ~i_10_192_3409_0 & i_10_192_3857_0))) | (~i_10_192_223_0 & ((i_10_192_795_0 & ~i_10_192_3203_0 & ~i_10_192_3784_0 & ~i_10_192_3785_0) | (~i_10_192_1687_0 & ~i_10_192_2180_0 & i_10_192_4567_0))) | (~i_10_192_1688_0 & i_10_192_1819_0) | (i_10_192_460_0 & i_10_192_2628_0 & i_10_192_2631_0 & ~i_10_192_3785_0) | (~i_10_192_3199_0 & ~i_10_192_3203_0 & ~i_10_192_3784_0) | (i_10_192_3585_0 & ~i_10_192_3781_0 & ~i_10_192_3786_0) | (i_10_192_1033_0 & ~i_10_192_3409_0 & ~i_10_192_3837_0 & ~i_10_192_4113_0 & ~i_10_192_4567_0) | (i_10_192_2352_0 & ~i_10_192_3408_0 & i_10_192_4568_0));
endmodule



// Benchmark "kernel_10_193" written by ABC on Sun Jul 19 10:24:20 2020

module kernel_10_193 ( 
    i_10_193_89_0, i_10_193_219_0, i_10_193_220_0, i_10_193_224_0,
    i_10_193_286_0, i_10_193_388_0, i_10_193_405_0, i_10_193_410_0,
    i_10_193_445_0, i_10_193_511_0, i_10_193_519_0, i_10_193_628_0,
    i_10_193_696_0, i_10_193_697_0, i_10_193_698_0, i_10_193_797_0,
    i_10_193_799_0, i_10_193_846_0, i_10_193_850_0, i_10_193_853_0,
    i_10_193_949_0, i_10_193_963_0, i_10_193_976_0, i_10_193_1060_0,
    i_10_193_1124_0, i_10_193_1237_0, i_10_193_1247_0, i_10_193_1249_0,
    i_10_193_1250_0, i_10_193_1308_0, i_10_193_1478_0, i_10_193_1651_0,
    i_10_193_1652_0, i_10_193_1688_0, i_10_193_1691_0, i_10_193_1711_0,
    i_10_193_1755_0, i_10_193_1776_0, i_10_193_1819_0, i_10_193_1820_0,
    i_10_193_1821_0, i_10_193_1823_0, i_10_193_1826_0, i_10_193_1913_0,
    i_10_193_1952_0, i_10_193_2020_0, i_10_193_2083_0, i_10_193_2272_0,
    i_10_193_2381_0, i_10_193_2382_0, i_10_193_2514_0, i_10_193_2517_0,
    i_10_193_2518_0, i_10_193_2533_0, i_10_193_2543_0, i_10_193_2563_0,
    i_10_193_2635_0, i_10_193_2653_0, i_10_193_2654_0, i_10_193_2722_0,
    i_10_193_2724_0, i_10_193_2732_0, i_10_193_2758_0, i_10_193_2820_0,
    i_10_193_2830_0, i_10_193_2833_0, i_10_193_2918_0, i_10_193_3049_0,
    i_10_193_3118_0, i_10_193_3165_0, i_10_193_3166_0, i_10_193_3198_0,
    i_10_193_3200_0, i_10_193_3273_0, i_10_193_3275_0, i_10_193_3358_0,
    i_10_193_3388_0, i_10_193_3392_0, i_10_193_3407_0, i_10_193_3409_0,
    i_10_193_3410_0, i_10_193_3544_0, i_10_193_3640_0, i_10_193_3705_0,
    i_10_193_3706_0, i_10_193_3732_0, i_10_193_3832_0, i_10_193_3838_0,
    i_10_193_3840_0, i_10_193_3851_0, i_10_193_3860_0, i_10_193_3905_0,
    i_10_193_3978_0, i_10_193_3979_0, i_10_193_4129_0, i_10_193_4184_0,
    i_10_193_4288_0, i_10_193_4460_0, i_10_193_4480_0, i_10_193_4570_0,
    o_10_193_0_0  );
  input  i_10_193_89_0, i_10_193_219_0, i_10_193_220_0, i_10_193_224_0,
    i_10_193_286_0, i_10_193_388_0, i_10_193_405_0, i_10_193_410_0,
    i_10_193_445_0, i_10_193_511_0, i_10_193_519_0, i_10_193_628_0,
    i_10_193_696_0, i_10_193_697_0, i_10_193_698_0, i_10_193_797_0,
    i_10_193_799_0, i_10_193_846_0, i_10_193_850_0, i_10_193_853_0,
    i_10_193_949_0, i_10_193_963_0, i_10_193_976_0, i_10_193_1060_0,
    i_10_193_1124_0, i_10_193_1237_0, i_10_193_1247_0, i_10_193_1249_0,
    i_10_193_1250_0, i_10_193_1308_0, i_10_193_1478_0, i_10_193_1651_0,
    i_10_193_1652_0, i_10_193_1688_0, i_10_193_1691_0, i_10_193_1711_0,
    i_10_193_1755_0, i_10_193_1776_0, i_10_193_1819_0, i_10_193_1820_0,
    i_10_193_1821_0, i_10_193_1823_0, i_10_193_1826_0, i_10_193_1913_0,
    i_10_193_1952_0, i_10_193_2020_0, i_10_193_2083_0, i_10_193_2272_0,
    i_10_193_2381_0, i_10_193_2382_0, i_10_193_2514_0, i_10_193_2517_0,
    i_10_193_2518_0, i_10_193_2533_0, i_10_193_2543_0, i_10_193_2563_0,
    i_10_193_2635_0, i_10_193_2653_0, i_10_193_2654_0, i_10_193_2722_0,
    i_10_193_2724_0, i_10_193_2732_0, i_10_193_2758_0, i_10_193_2820_0,
    i_10_193_2830_0, i_10_193_2833_0, i_10_193_2918_0, i_10_193_3049_0,
    i_10_193_3118_0, i_10_193_3165_0, i_10_193_3166_0, i_10_193_3198_0,
    i_10_193_3200_0, i_10_193_3273_0, i_10_193_3275_0, i_10_193_3358_0,
    i_10_193_3388_0, i_10_193_3392_0, i_10_193_3407_0, i_10_193_3409_0,
    i_10_193_3410_0, i_10_193_3544_0, i_10_193_3640_0, i_10_193_3705_0,
    i_10_193_3706_0, i_10_193_3732_0, i_10_193_3832_0, i_10_193_3838_0,
    i_10_193_3840_0, i_10_193_3851_0, i_10_193_3860_0, i_10_193_3905_0,
    i_10_193_3978_0, i_10_193_3979_0, i_10_193_4129_0, i_10_193_4184_0,
    i_10_193_4288_0, i_10_193_4460_0, i_10_193_4480_0, i_10_193_4570_0;
  output o_10_193_0_0;
  assign o_10_193_0_0 = 0;
endmodule



// Benchmark "kernel_10_194" written by ABC on Sun Jul 19 10:24:21 2020

module kernel_10_194 ( 
    i_10_194_28_0, i_10_194_118_0, i_10_194_119_0, i_10_194_122_0,
    i_10_194_220_0, i_10_194_221_0, i_10_194_250_0, i_10_194_281_0,
    i_10_194_284_0, i_10_194_316_0, i_10_194_329_0, i_10_194_388_0,
    i_10_194_431_0, i_10_194_433_0, i_10_194_437_0, i_10_194_460_0,
    i_10_194_520_0, i_10_194_749_0, i_10_194_754_0, i_10_194_793_0,
    i_10_194_794_0, i_10_194_797_0, i_10_194_968_0, i_10_194_990_0,
    i_10_194_1000_0, i_10_194_1236_0, i_10_194_1240_0, i_10_194_1241_0,
    i_10_194_1261_0, i_10_194_1308_0, i_10_194_1309_0, i_10_194_1578_0,
    i_10_194_1647_0, i_10_194_1650_0, i_10_194_1651_0, i_10_194_1652_0,
    i_10_194_1686_0, i_10_194_1687_0, i_10_194_1732_0, i_10_194_1821_0,
    i_10_194_1822_0, i_10_194_1912_0, i_10_194_1944_0, i_10_194_2186_0,
    i_10_194_2242_0, i_10_194_2350_0, i_10_194_2352_0, i_10_194_2354_0,
    i_10_194_2355_0, i_10_194_2357_0, i_10_194_2467_0, i_10_194_2473_0,
    i_10_194_2632_0, i_10_194_2633_0, i_10_194_2658_0, i_10_194_2660_0,
    i_10_194_2701_0, i_10_194_2732_0, i_10_194_2788_0, i_10_194_2827_0,
    i_10_194_2832_0, i_10_194_2886_0, i_10_194_2888_0, i_10_194_2922_0,
    i_10_194_3036_0, i_10_194_3037_0, i_10_194_3038_0, i_10_194_3046_0,
    i_10_194_3049_0, i_10_194_3075_0, i_10_194_3076_0, i_10_194_3088_0,
    i_10_194_3198_0, i_10_194_3199_0, i_10_194_3276_0, i_10_194_3390_0,
    i_10_194_3391_0, i_10_194_3406_0, i_10_194_3466_0, i_10_194_3587_0,
    i_10_194_3609_0, i_10_194_3649_0, i_10_194_3650_0, i_10_194_3653_0,
    i_10_194_3782_0, i_10_194_3785_0, i_10_194_3788_0, i_10_194_3855_0,
    i_10_194_3856_0, i_10_194_3893_0, i_10_194_3979_0, i_10_194_3980_0,
    i_10_194_4114_0, i_10_194_4115_0, i_10_194_4117_0, i_10_194_4127_0,
    i_10_194_4270_0, i_10_194_4288_0, i_10_194_4289_0, i_10_194_4567_0,
    o_10_194_0_0  );
  input  i_10_194_28_0, i_10_194_118_0, i_10_194_119_0, i_10_194_122_0,
    i_10_194_220_0, i_10_194_221_0, i_10_194_250_0, i_10_194_281_0,
    i_10_194_284_0, i_10_194_316_0, i_10_194_329_0, i_10_194_388_0,
    i_10_194_431_0, i_10_194_433_0, i_10_194_437_0, i_10_194_460_0,
    i_10_194_520_0, i_10_194_749_0, i_10_194_754_0, i_10_194_793_0,
    i_10_194_794_0, i_10_194_797_0, i_10_194_968_0, i_10_194_990_0,
    i_10_194_1000_0, i_10_194_1236_0, i_10_194_1240_0, i_10_194_1241_0,
    i_10_194_1261_0, i_10_194_1308_0, i_10_194_1309_0, i_10_194_1578_0,
    i_10_194_1647_0, i_10_194_1650_0, i_10_194_1651_0, i_10_194_1652_0,
    i_10_194_1686_0, i_10_194_1687_0, i_10_194_1732_0, i_10_194_1821_0,
    i_10_194_1822_0, i_10_194_1912_0, i_10_194_1944_0, i_10_194_2186_0,
    i_10_194_2242_0, i_10_194_2350_0, i_10_194_2352_0, i_10_194_2354_0,
    i_10_194_2355_0, i_10_194_2357_0, i_10_194_2467_0, i_10_194_2473_0,
    i_10_194_2632_0, i_10_194_2633_0, i_10_194_2658_0, i_10_194_2660_0,
    i_10_194_2701_0, i_10_194_2732_0, i_10_194_2788_0, i_10_194_2827_0,
    i_10_194_2832_0, i_10_194_2886_0, i_10_194_2888_0, i_10_194_2922_0,
    i_10_194_3036_0, i_10_194_3037_0, i_10_194_3038_0, i_10_194_3046_0,
    i_10_194_3049_0, i_10_194_3075_0, i_10_194_3076_0, i_10_194_3088_0,
    i_10_194_3198_0, i_10_194_3199_0, i_10_194_3276_0, i_10_194_3390_0,
    i_10_194_3391_0, i_10_194_3406_0, i_10_194_3466_0, i_10_194_3587_0,
    i_10_194_3609_0, i_10_194_3649_0, i_10_194_3650_0, i_10_194_3653_0,
    i_10_194_3782_0, i_10_194_3785_0, i_10_194_3788_0, i_10_194_3855_0,
    i_10_194_3856_0, i_10_194_3893_0, i_10_194_3979_0, i_10_194_3980_0,
    i_10_194_4114_0, i_10_194_4115_0, i_10_194_4117_0, i_10_194_4127_0,
    i_10_194_4270_0, i_10_194_4288_0, i_10_194_4289_0, i_10_194_4567_0;
  output o_10_194_0_0;
  assign o_10_194_0_0 = ~((~i_10_194_3049_0 & ((~i_10_194_122_0 & ((~i_10_194_431_0 & ~i_10_194_520_0 & ~i_10_194_2186_0 & ~i_10_194_2473_0 & ~i_10_194_3076_0 & ~i_10_194_3088_0 & ~i_10_194_3856_0) | (~i_10_194_433_0 & ~i_10_194_1822_0 & ~i_10_194_1912_0 & ~i_10_194_2660_0 & ~i_10_194_3609_0 & ~i_10_194_4567_0))) | (~i_10_194_1240_0 & ((~i_10_194_1241_0 & i_10_194_1309_0 & ~i_10_194_2352_0 & ~i_10_194_2355_0 & ~i_10_194_2788_0 & i_10_194_3198_0) | (~i_10_194_118_0 & ~i_10_194_431_0 & ~i_10_194_3198_0 & ~i_10_194_3390_0 & ~i_10_194_3587_0 & ~i_10_194_3788_0))) | (~i_10_194_28_0 & ~i_10_194_281_0 & ~i_10_194_437_0 & ~i_10_194_1241_0 & ~i_10_194_1912_0 & ~i_10_194_2186_0 & ~i_10_194_2357_0 & ~i_10_194_2633_0 & ~i_10_194_2788_0 & ~i_10_194_3076_0 & ~i_10_194_3199_0))) | (~i_10_194_2788_0 & ((~i_10_194_118_0 & ((~i_10_194_1308_0 & ~i_10_194_1309_0 & ~i_10_194_2354_0 & ~i_10_194_2357_0) | (~i_10_194_2473_0 & ~i_10_194_3037_0 & ~i_10_194_3038_0))) | (~i_10_194_2467_0 & ~i_10_194_2888_0 & ((~i_10_194_2354_0 & ~i_10_194_3390_0 & ~i_10_194_3466_0 & ~i_10_194_3587_0 & ~i_10_194_3785_0) | (i_10_194_1822_0 & ~i_10_194_2186_0 & i_10_194_2352_0 & ~i_10_194_3391_0 & ~i_10_194_3788_0 & ~i_10_194_3979_0))) | (~i_10_194_2660_0 & ~i_10_194_3076_0 & ~i_10_194_3653_0 & ~i_10_194_3856_0))) | (~i_10_194_122_0 & ((~i_10_194_1000_0 & ~i_10_194_1822_0 & ~i_10_194_2186_0 & ~i_10_194_2886_0 & ~i_10_194_3036_0 & ~i_10_194_3076_0 & ~i_10_194_3390_0 & ~i_10_194_3391_0 & ~i_10_194_3788_0) | (~i_10_194_1821_0 & ~i_10_194_2660_0 & ~i_10_194_2832_0 & ~i_10_194_3037_0 & ~i_10_194_3649_0 & ~i_10_194_3856_0))) | (i_10_194_1236_0 & ~i_10_194_3979_0 & ((~i_10_194_1241_0 & i_10_194_1578_0 & i_10_194_1822_0 & ~i_10_194_3650_0) | (~i_10_194_250_0 & ~i_10_194_3076_0 & ~i_10_194_3587_0 & ~i_10_194_3649_0 & ~i_10_194_3653_0))) | (i_10_194_1912_0 & ((i_10_194_520_0 & ~i_10_194_1308_0 & i_10_194_3785_0) | (~i_10_194_2473_0 & i_10_194_2827_0 & ~i_10_194_3390_0 & ~i_10_194_3391_0 & ~i_10_194_3980_0))) | (i_10_194_1578_0 & ~i_10_194_3036_0 & ~i_10_194_3038_0) | (~i_10_194_2186_0 & ~i_10_194_2658_0 & ~i_10_194_2832_0 & ~i_10_194_3037_0 & ~i_10_194_3587_0) | (~i_10_194_1309_0 & ~i_10_194_1912_0 & ~i_10_194_3856_0 & ~i_10_194_3980_0) | (~i_10_194_1000_0 & ~i_10_194_1241_0 & i_10_194_1652_0 & ~i_10_194_1944_0 & ~i_10_194_4567_0));
endmodule



// Benchmark "kernel_10_195" written by ABC on Sun Jul 19 10:24:22 2020

module kernel_10_195 ( 
    i_10_195_45_0, i_10_195_144_0, i_10_195_219_0, i_10_195_280_0,
    i_10_195_283_0, i_10_195_287_0, i_10_195_316_0, i_10_195_320_0,
    i_10_195_328_0, i_10_195_390_0, i_10_195_392_0, i_10_195_437_0,
    i_10_195_440_0, i_10_195_442_0, i_10_195_463_0, i_10_195_464_0,
    i_10_195_711_0, i_10_195_712_0, i_10_195_821_0, i_10_195_1234_0,
    i_10_195_1240_0, i_10_195_1241_0, i_10_195_1245_0, i_10_195_1246_0,
    i_10_195_1298_0, i_10_195_1363_0, i_10_195_1433_0, i_10_195_1441_0,
    i_10_195_1445_0, i_10_195_1551_0, i_10_195_1552_0, i_10_195_1553_0,
    i_10_195_1580_0, i_10_195_1622_0, i_10_195_1649_0, i_10_195_1655_0,
    i_10_195_1683_0, i_10_195_1684_0, i_10_195_1686_0, i_10_195_1687_0,
    i_10_195_1769_0, i_10_195_1943_0, i_10_195_1952_0, i_10_195_1982_0,
    i_10_195_2003_0, i_10_195_2185_0, i_10_195_2312_0, i_10_195_2349_0,
    i_10_195_2358_0, i_10_195_2361_0, i_10_195_2362_0, i_10_195_2448_0,
    i_10_195_2449_0, i_10_195_2450_0, i_10_195_2456_0, i_10_195_2468_0,
    i_10_195_2473_0, i_10_195_2516_0, i_10_195_2593_0, i_10_195_2629_0,
    i_10_195_2630_0, i_10_195_2631_0, i_10_195_2632_0, i_10_195_2638_0,
    i_10_195_2655_0, i_10_195_2658_0, i_10_195_2660_0, i_10_195_2661_0,
    i_10_195_2718_0, i_10_195_2720_0, i_10_195_2723_0, i_10_195_2728_0,
    i_10_195_2781_0, i_10_195_2818_0, i_10_195_2887_0, i_10_195_2963_0,
    i_10_195_3071_0, i_10_195_3231_0, i_10_195_3388_0, i_10_195_3389_0,
    i_10_195_3469_0, i_10_195_3540_0, i_10_195_3583_0, i_10_195_3586_0,
    i_10_195_3587_0, i_10_195_3650_0, i_10_195_3784_0, i_10_195_3835_0,
    i_10_195_3838_0, i_10_195_3839_0, i_10_195_3884_0, i_10_195_3910_0,
    i_10_195_4028_0, i_10_195_4119_0, i_10_195_4124_0, i_10_195_4127_0,
    i_10_195_4142_0, i_10_195_4145_0, i_10_195_4266_0, i_10_195_4289_0,
    o_10_195_0_0  );
  input  i_10_195_45_0, i_10_195_144_0, i_10_195_219_0, i_10_195_280_0,
    i_10_195_283_0, i_10_195_287_0, i_10_195_316_0, i_10_195_320_0,
    i_10_195_328_0, i_10_195_390_0, i_10_195_392_0, i_10_195_437_0,
    i_10_195_440_0, i_10_195_442_0, i_10_195_463_0, i_10_195_464_0,
    i_10_195_711_0, i_10_195_712_0, i_10_195_821_0, i_10_195_1234_0,
    i_10_195_1240_0, i_10_195_1241_0, i_10_195_1245_0, i_10_195_1246_0,
    i_10_195_1298_0, i_10_195_1363_0, i_10_195_1433_0, i_10_195_1441_0,
    i_10_195_1445_0, i_10_195_1551_0, i_10_195_1552_0, i_10_195_1553_0,
    i_10_195_1580_0, i_10_195_1622_0, i_10_195_1649_0, i_10_195_1655_0,
    i_10_195_1683_0, i_10_195_1684_0, i_10_195_1686_0, i_10_195_1687_0,
    i_10_195_1769_0, i_10_195_1943_0, i_10_195_1952_0, i_10_195_1982_0,
    i_10_195_2003_0, i_10_195_2185_0, i_10_195_2312_0, i_10_195_2349_0,
    i_10_195_2358_0, i_10_195_2361_0, i_10_195_2362_0, i_10_195_2448_0,
    i_10_195_2449_0, i_10_195_2450_0, i_10_195_2456_0, i_10_195_2468_0,
    i_10_195_2473_0, i_10_195_2516_0, i_10_195_2593_0, i_10_195_2629_0,
    i_10_195_2630_0, i_10_195_2631_0, i_10_195_2632_0, i_10_195_2638_0,
    i_10_195_2655_0, i_10_195_2658_0, i_10_195_2660_0, i_10_195_2661_0,
    i_10_195_2718_0, i_10_195_2720_0, i_10_195_2723_0, i_10_195_2728_0,
    i_10_195_2781_0, i_10_195_2818_0, i_10_195_2887_0, i_10_195_2963_0,
    i_10_195_3071_0, i_10_195_3231_0, i_10_195_3388_0, i_10_195_3389_0,
    i_10_195_3469_0, i_10_195_3540_0, i_10_195_3583_0, i_10_195_3586_0,
    i_10_195_3587_0, i_10_195_3650_0, i_10_195_3784_0, i_10_195_3835_0,
    i_10_195_3838_0, i_10_195_3839_0, i_10_195_3884_0, i_10_195_3910_0,
    i_10_195_4028_0, i_10_195_4119_0, i_10_195_4124_0, i_10_195_4127_0,
    i_10_195_4142_0, i_10_195_4145_0, i_10_195_4266_0, i_10_195_4289_0;
  output o_10_195_0_0;
  assign o_10_195_0_0 = 0;
endmodule



// Benchmark "kernel_10_196" written by ABC on Sun Jul 19 10:24:23 2020

module kernel_10_196 ( 
    i_10_196_83_0, i_10_196_283_0, i_10_196_284_0, i_10_196_289_0,
    i_10_196_325_0, i_10_196_442_0, i_10_196_446_0, i_10_196_461_0,
    i_10_196_464_0, i_10_196_504_0, i_10_196_508_0, i_10_196_514_0,
    i_10_196_545_0, i_10_196_892_0, i_10_196_893_0, i_10_196_1027_0,
    i_10_196_1028_0, i_10_196_1135_0, i_10_196_1139_0, i_10_196_1233_0,
    i_10_196_1234_0, i_10_196_1236_0, i_10_196_1238_0, i_10_196_1243_0,
    i_10_196_1244_0, i_10_196_1264_0, i_10_196_1306_0, i_10_196_1313_0,
    i_10_196_1650_0, i_10_196_1652_0, i_10_196_1690_0, i_10_196_1818_0,
    i_10_196_1819_0, i_10_196_1823_0, i_10_196_1909_0, i_10_196_1910_0,
    i_10_196_1912_0, i_10_196_1913_0, i_10_196_1989_0, i_10_196_1990_0,
    i_10_196_1991_0, i_10_196_2017_0, i_10_196_2198_0, i_10_196_2353_0,
    i_10_196_2358_0, i_10_196_2359_0, i_10_196_2360_0, i_10_196_2361_0,
    i_10_196_2362_0, i_10_196_2408_0, i_10_196_2449_0, i_10_196_2457_0,
    i_10_196_2458_0, i_10_196_2459_0, i_10_196_2462_0, i_10_196_2470_0,
    i_10_196_2601_0, i_10_196_2700_0, i_10_196_2709_0, i_10_196_2728_0,
    i_10_196_2818_0, i_10_196_2828_0, i_10_196_2830_0, i_10_196_2882_0,
    i_10_196_2918_0, i_10_196_2920_0, i_10_196_2921_0, i_10_196_3150_0,
    i_10_196_3269_0, i_10_196_3272_0, i_10_196_3277_0, i_10_196_3386_0,
    i_10_196_3388_0, i_10_196_3389_0, i_10_196_3402_0, i_10_196_3406_0,
    i_10_196_3523_0, i_10_196_3587_0, i_10_196_3722_0, i_10_196_3783_0,
    i_10_196_3784_0, i_10_196_3785_0, i_10_196_3787_0, i_10_196_3830_0,
    i_10_196_3834_0, i_10_196_3848_0, i_10_196_3849_0, i_10_196_3850_0,
    i_10_196_3854_0, i_10_196_3855_0, i_10_196_3856_0, i_10_196_3857_0,
    i_10_196_3890_0, i_10_196_3892_0, i_10_196_3982_0, i_10_196_3986_0,
    i_10_196_4024_0, i_10_196_4233_0, i_10_196_4565_0, i_10_196_4567_0,
    o_10_196_0_0  );
  input  i_10_196_83_0, i_10_196_283_0, i_10_196_284_0, i_10_196_289_0,
    i_10_196_325_0, i_10_196_442_0, i_10_196_446_0, i_10_196_461_0,
    i_10_196_464_0, i_10_196_504_0, i_10_196_508_0, i_10_196_514_0,
    i_10_196_545_0, i_10_196_892_0, i_10_196_893_0, i_10_196_1027_0,
    i_10_196_1028_0, i_10_196_1135_0, i_10_196_1139_0, i_10_196_1233_0,
    i_10_196_1234_0, i_10_196_1236_0, i_10_196_1238_0, i_10_196_1243_0,
    i_10_196_1244_0, i_10_196_1264_0, i_10_196_1306_0, i_10_196_1313_0,
    i_10_196_1650_0, i_10_196_1652_0, i_10_196_1690_0, i_10_196_1818_0,
    i_10_196_1819_0, i_10_196_1823_0, i_10_196_1909_0, i_10_196_1910_0,
    i_10_196_1912_0, i_10_196_1913_0, i_10_196_1989_0, i_10_196_1990_0,
    i_10_196_1991_0, i_10_196_2017_0, i_10_196_2198_0, i_10_196_2353_0,
    i_10_196_2358_0, i_10_196_2359_0, i_10_196_2360_0, i_10_196_2361_0,
    i_10_196_2362_0, i_10_196_2408_0, i_10_196_2449_0, i_10_196_2457_0,
    i_10_196_2458_0, i_10_196_2459_0, i_10_196_2462_0, i_10_196_2470_0,
    i_10_196_2601_0, i_10_196_2700_0, i_10_196_2709_0, i_10_196_2728_0,
    i_10_196_2818_0, i_10_196_2828_0, i_10_196_2830_0, i_10_196_2882_0,
    i_10_196_2918_0, i_10_196_2920_0, i_10_196_2921_0, i_10_196_3150_0,
    i_10_196_3269_0, i_10_196_3272_0, i_10_196_3277_0, i_10_196_3386_0,
    i_10_196_3388_0, i_10_196_3389_0, i_10_196_3402_0, i_10_196_3406_0,
    i_10_196_3523_0, i_10_196_3587_0, i_10_196_3722_0, i_10_196_3783_0,
    i_10_196_3784_0, i_10_196_3785_0, i_10_196_3787_0, i_10_196_3830_0,
    i_10_196_3834_0, i_10_196_3848_0, i_10_196_3849_0, i_10_196_3850_0,
    i_10_196_3854_0, i_10_196_3855_0, i_10_196_3856_0, i_10_196_3857_0,
    i_10_196_3890_0, i_10_196_3892_0, i_10_196_3982_0, i_10_196_3986_0,
    i_10_196_4024_0, i_10_196_4233_0, i_10_196_4565_0, i_10_196_4567_0;
  output o_10_196_0_0;
  assign o_10_196_0_0 = ~((~i_10_196_1028_0 & ((~i_10_196_893_0 & ~i_10_196_2601_0 & ~i_10_196_2921_0 & ~i_10_196_3402_0 & ~i_10_196_3783_0 & ~i_10_196_3787_0) | (~i_10_196_283_0 & ~i_10_196_892_0 & ~i_10_196_1313_0 & ~i_10_196_3848_0 & ~i_10_196_3849_0))) | (~i_10_196_892_0 & ((i_10_196_442_0 & ~i_10_196_2457_0 & ~i_10_196_2459_0 & ~i_10_196_3272_0) | (~i_10_196_2458_0 & ~i_10_196_2462_0 & ~i_10_196_2830_0 & ~i_10_196_3386_0))) | (~i_10_196_1238_0 & ((~i_10_196_893_0 & i_10_196_1818_0 & ~i_10_196_2360_0 & ~i_10_196_2458_0 & ~i_10_196_2728_0 & ~i_10_196_3848_0) | (i_10_196_2358_0 & i_10_196_2360_0 & ~i_10_196_2457_0 & ~i_10_196_3269_0 & ~i_10_196_3389_0 & ~i_10_196_3850_0))) | (~i_10_196_893_0 & ~i_10_196_2362_0 & ((~i_10_196_1989_0 & ~i_10_196_2359_0 & ~i_10_196_3784_0) | (~i_10_196_3269_0 & ~i_10_196_3787_0 & ~i_10_196_4024_0))) | (~i_10_196_1313_0 & ~i_10_196_3269_0 & ((~i_10_196_83_0 & ~i_10_196_1989_0 & ~i_10_196_2360_0 & ~i_10_196_2830_0 & ~i_10_196_3389_0) | (i_10_196_283_0 & ~i_10_196_289_0 & ~i_10_196_1690_0 & ~i_10_196_2462_0 & ~i_10_196_3850_0 & ~i_10_196_3855_0 & ~i_10_196_4567_0))) | (~i_10_196_83_0 & ((~i_10_196_1306_0 & ~i_10_196_1690_0 & ~i_10_196_1991_0 & ~i_10_196_2459_0 & ~i_10_196_2728_0 & ~i_10_196_3783_0 & ~i_10_196_3785_0 & ~i_10_196_3855_0) | (i_10_196_2361_0 & ~i_10_196_3386_0 & ~i_10_196_3787_0 & ~i_10_196_3850_0 & ~i_10_196_4024_0))) | (~i_10_196_2360_0 & ~i_10_196_2457_0 & ((~i_10_196_3386_0 & ~i_10_196_3388_0 & ~i_10_196_3857_0) | (~i_10_196_1264_0 & ~i_10_196_2361_0 & ~i_10_196_2601_0 & ~i_10_196_3848_0 & ~i_10_196_4565_0))) | (~i_10_196_2458_0 & ((i_10_196_1306_0 & i_10_196_2449_0 & ~i_10_196_3855_0) | (i_10_196_284_0 & ~i_10_196_1652_0 & ~i_10_196_2470_0 & ~i_10_196_2921_0 & ~i_10_196_3848_0 & ~i_10_196_3857_0))) | (i_10_196_514_0 & i_10_196_2353_0) | (i_10_196_461_0 & ~i_10_196_3388_0) | (~i_10_196_1027_0 & ~i_10_196_1991_0 & ~i_10_196_2459_0 & ~i_10_196_3389_0 & ~i_10_196_3848_0 & ~i_10_196_4024_0) | (i_10_196_1652_0 & ~i_10_196_3787_0 & i_10_196_4024_0 & i_10_196_4567_0));
endmodule



// Benchmark "kernel_10_197" written by ABC on Sun Jul 19 10:24:24 2020

module kernel_10_197 ( 
    i_10_197_89_0, i_10_197_177_0, i_10_197_214_0, i_10_197_259_0,
    i_10_197_325_0, i_10_197_329_0, i_10_197_370_0, i_10_197_446_0,
    i_10_197_518_0, i_10_197_543_0, i_10_197_738_0, i_10_197_793_0,
    i_10_197_797_0, i_10_197_799_0, i_10_197_827_0, i_10_197_963_0,
    i_10_197_967_0, i_10_197_999_0, i_10_197_1083_0, i_10_197_1087_0,
    i_10_197_1120_0, i_10_197_1205_0, i_10_197_1237_0, i_10_197_1245_0,
    i_10_197_1248_0, i_10_197_1306_0, i_10_197_1312_0, i_10_197_1313_0,
    i_10_197_1344_0, i_10_197_1542_0, i_10_197_1553_0, i_10_197_1647_0,
    i_10_197_1650_0, i_10_197_1685_0, i_10_197_1689_0, i_10_197_1690_0,
    i_10_197_1818_0, i_10_197_2019_0, i_10_197_2182_0, i_10_197_2338_0,
    i_10_197_2350_0, i_10_197_2378_0, i_10_197_2404_0, i_10_197_2407_0,
    i_10_197_2451_0, i_10_197_2472_0, i_10_197_2629_0, i_10_197_2631_0,
    i_10_197_2632_0, i_10_197_2636_0, i_10_197_2707_0, i_10_197_2713_0,
    i_10_197_2714_0, i_10_197_2718_0, i_10_197_2727_0, i_10_197_2731_0,
    i_10_197_2781_0, i_10_197_2823_0, i_10_197_2824_0, i_10_197_2828_0,
    i_10_197_2832_0, i_10_197_2850_0, i_10_197_2868_0, i_10_197_2887_0,
    i_10_197_2922_0, i_10_197_2954_0, i_10_197_2957_0, i_10_197_2983_0,
    i_10_197_3037_0, i_10_197_3038_0, i_10_197_3092_0, i_10_197_3268_0,
    i_10_197_3274_0, i_10_197_3280_0, i_10_197_3328_0, i_10_197_3388_0,
    i_10_197_3405_0, i_10_197_3432_0, i_10_197_3444_0, i_10_197_3447_0,
    i_10_197_3526_0, i_10_197_3583_0, i_10_197_3589_0, i_10_197_3612_0,
    i_10_197_3613_0, i_10_197_3616_0, i_10_197_3672_0, i_10_197_3687_0,
    i_10_197_3813_0, i_10_197_3841_0, i_10_197_3843_0, i_10_197_3844_0,
    i_10_197_3946_0, i_10_197_4156_0, i_10_197_4157_0, i_10_197_4175_0,
    i_10_197_4215_0, i_10_197_4272_0, i_10_197_4273_0, i_10_197_4565_0,
    o_10_197_0_0  );
  input  i_10_197_89_0, i_10_197_177_0, i_10_197_214_0, i_10_197_259_0,
    i_10_197_325_0, i_10_197_329_0, i_10_197_370_0, i_10_197_446_0,
    i_10_197_518_0, i_10_197_543_0, i_10_197_738_0, i_10_197_793_0,
    i_10_197_797_0, i_10_197_799_0, i_10_197_827_0, i_10_197_963_0,
    i_10_197_967_0, i_10_197_999_0, i_10_197_1083_0, i_10_197_1087_0,
    i_10_197_1120_0, i_10_197_1205_0, i_10_197_1237_0, i_10_197_1245_0,
    i_10_197_1248_0, i_10_197_1306_0, i_10_197_1312_0, i_10_197_1313_0,
    i_10_197_1344_0, i_10_197_1542_0, i_10_197_1553_0, i_10_197_1647_0,
    i_10_197_1650_0, i_10_197_1685_0, i_10_197_1689_0, i_10_197_1690_0,
    i_10_197_1818_0, i_10_197_2019_0, i_10_197_2182_0, i_10_197_2338_0,
    i_10_197_2350_0, i_10_197_2378_0, i_10_197_2404_0, i_10_197_2407_0,
    i_10_197_2451_0, i_10_197_2472_0, i_10_197_2629_0, i_10_197_2631_0,
    i_10_197_2632_0, i_10_197_2636_0, i_10_197_2707_0, i_10_197_2713_0,
    i_10_197_2714_0, i_10_197_2718_0, i_10_197_2727_0, i_10_197_2731_0,
    i_10_197_2781_0, i_10_197_2823_0, i_10_197_2824_0, i_10_197_2828_0,
    i_10_197_2832_0, i_10_197_2850_0, i_10_197_2868_0, i_10_197_2887_0,
    i_10_197_2922_0, i_10_197_2954_0, i_10_197_2957_0, i_10_197_2983_0,
    i_10_197_3037_0, i_10_197_3038_0, i_10_197_3092_0, i_10_197_3268_0,
    i_10_197_3274_0, i_10_197_3280_0, i_10_197_3328_0, i_10_197_3388_0,
    i_10_197_3405_0, i_10_197_3432_0, i_10_197_3444_0, i_10_197_3447_0,
    i_10_197_3526_0, i_10_197_3583_0, i_10_197_3589_0, i_10_197_3612_0,
    i_10_197_3613_0, i_10_197_3616_0, i_10_197_3672_0, i_10_197_3687_0,
    i_10_197_3813_0, i_10_197_3841_0, i_10_197_3843_0, i_10_197_3844_0,
    i_10_197_3946_0, i_10_197_4156_0, i_10_197_4157_0, i_10_197_4175_0,
    i_10_197_4215_0, i_10_197_4272_0, i_10_197_4273_0, i_10_197_4565_0;
  output o_10_197_0_0;
  assign o_10_197_0_0 = 0;
endmodule



// Benchmark "kernel_10_198" written by ABC on Sun Jul 19 10:24:25 2020

module kernel_10_198 ( 
    i_10_198_24_0, i_10_198_64_0, i_10_198_67_0, i_10_198_70_0,
    i_10_198_175_0, i_10_198_183_0, i_10_198_272_0, i_10_198_283_0,
    i_10_198_319_0, i_10_198_408_0, i_10_198_410_0, i_10_198_434_0,
    i_10_198_458_0, i_10_198_536_0, i_10_198_817_0, i_10_198_905_0,
    i_10_198_906_0, i_10_198_947_0, i_10_198_951_0, i_10_198_956_0,
    i_10_198_1064_0, i_10_198_1119_0, i_10_198_1172_0, i_10_198_1286_0,
    i_10_198_1375_0, i_10_198_1445_0, i_10_198_1482_0, i_10_198_1484_0,
    i_10_198_1551_0, i_10_198_1554_0, i_10_198_1632_0, i_10_198_1641_0,
    i_10_198_1647_0, i_10_198_1684_0, i_10_198_1790_0, i_10_198_1819_0,
    i_10_198_1822_0, i_10_198_1887_0, i_10_198_1911_0, i_10_198_1912_0,
    i_10_198_1915_0, i_10_198_1916_0, i_10_198_1918_0, i_10_198_1919_0,
    i_10_198_1932_0, i_10_198_1933_0, i_10_198_2027_0, i_10_198_2059_0,
    i_10_198_2063_0, i_10_198_2094_0, i_10_198_2095_0, i_10_198_2154_0,
    i_10_198_2157_0, i_10_198_2158_0, i_10_198_2274_0, i_10_198_2275_0,
    i_10_198_2311_0, i_10_198_2312_0, i_10_198_2337_0, i_10_198_2351_0,
    i_10_198_2352_0, i_10_198_2353_0, i_10_198_2354_0, i_10_198_2357_0,
    i_10_198_2452_0, i_10_198_2453_0, i_10_198_2508_0, i_10_198_2509_0,
    i_10_198_2541_0, i_10_198_2557_0, i_10_198_2605_0, i_10_198_2635_0,
    i_10_198_2640_0, i_10_198_2663_0, i_10_198_2698_0, i_10_198_2770_0,
    i_10_198_2820_0, i_10_198_2848_0, i_10_198_2856_0, i_10_198_2857_0,
    i_10_198_2919_0, i_10_198_2922_0, i_10_198_3031_0, i_10_198_3032_0,
    i_10_198_3074_0, i_10_198_3102_0, i_10_198_3103_0, i_10_198_3104_0,
    i_10_198_3229_0, i_10_198_3545_0, i_10_198_3610_0, i_10_198_3647_0,
    i_10_198_3775_0, i_10_198_3805_0, i_10_198_3806_0, i_10_198_3859_0,
    i_10_198_3982_0, i_10_198_4126_0, i_10_198_4364_0, i_10_198_4534_0,
    o_10_198_0_0  );
  input  i_10_198_24_0, i_10_198_64_0, i_10_198_67_0, i_10_198_70_0,
    i_10_198_175_0, i_10_198_183_0, i_10_198_272_0, i_10_198_283_0,
    i_10_198_319_0, i_10_198_408_0, i_10_198_410_0, i_10_198_434_0,
    i_10_198_458_0, i_10_198_536_0, i_10_198_817_0, i_10_198_905_0,
    i_10_198_906_0, i_10_198_947_0, i_10_198_951_0, i_10_198_956_0,
    i_10_198_1064_0, i_10_198_1119_0, i_10_198_1172_0, i_10_198_1286_0,
    i_10_198_1375_0, i_10_198_1445_0, i_10_198_1482_0, i_10_198_1484_0,
    i_10_198_1551_0, i_10_198_1554_0, i_10_198_1632_0, i_10_198_1641_0,
    i_10_198_1647_0, i_10_198_1684_0, i_10_198_1790_0, i_10_198_1819_0,
    i_10_198_1822_0, i_10_198_1887_0, i_10_198_1911_0, i_10_198_1912_0,
    i_10_198_1915_0, i_10_198_1916_0, i_10_198_1918_0, i_10_198_1919_0,
    i_10_198_1932_0, i_10_198_1933_0, i_10_198_2027_0, i_10_198_2059_0,
    i_10_198_2063_0, i_10_198_2094_0, i_10_198_2095_0, i_10_198_2154_0,
    i_10_198_2157_0, i_10_198_2158_0, i_10_198_2274_0, i_10_198_2275_0,
    i_10_198_2311_0, i_10_198_2312_0, i_10_198_2337_0, i_10_198_2351_0,
    i_10_198_2352_0, i_10_198_2353_0, i_10_198_2354_0, i_10_198_2357_0,
    i_10_198_2452_0, i_10_198_2453_0, i_10_198_2508_0, i_10_198_2509_0,
    i_10_198_2541_0, i_10_198_2557_0, i_10_198_2605_0, i_10_198_2635_0,
    i_10_198_2640_0, i_10_198_2663_0, i_10_198_2698_0, i_10_198_2770_0,
    i_10_198_2820_0, i_10_198_2848_0, i_10_198_2856_0, i_10_198_2857_0,
    i_10_198_2919_0, i_10_198_2922_0, i_10_198_3031_0, i_10_198_3032_0,
    i_10_198_3074_0, i_10_198_3102_0, i_10_198_3103_0, i_10_198_3104_0,
    i_10_198_3229_0, i_10_198_3545_0, i_10_198_3610_0, i_10_198_3647_0,
    i_10_198_3775_0, i_10_198_3805_0, i_10_198_3806_0, i_10_198_3859_0,
    i_10_198_3982_0, i_10_198_4126_0, i_10_198_4364_0, i_10_198_4534_0;
  output o_10_198_0_0;
  assign o_10_198_0_0 = 0;
endmodule



// Benchmark "kernel_10_199" written by ABC on Sun Jul 19 10:24:26 2020

module kernel_10_199 ( 
    i_10_199_27_0, i_10_199_124_0, i_10_199_175_0, i_10_199_285_0,
    i_10_199_369_0, i_10_199_433_0, i_10_199_443_0, i_10_199_444_0,
    i_10_199_467_0, i_10_199_501_0, i_10_199_532_0, i_10_199_729_0,
    i_10_199_730_0, i_10_199_732_0, i_10_199_733_0, i_10_199_901_0,
    i_10_199_961_0, i_10_199_999_0, i_10_199_1052_0, i_10_199_1201_0,
    i_10_199_1263_0, i_10_199_1265_0, i_10_199_1270_0, i_10_199_1271_0,
    i_10_199_1308_0, i_10_199_1309_0, i_10_199_1353_0, i_10_199_1361_0,
    i_10_199_1363_0, i_10_199_1638_0, i_10_199_1741_0, i_10_199_1765_0,
    i_10_199_1823_0, i_10_199_1912_0, i_10_199_1947_0, i_10_199_1948_0,
    i_10_199_1957_0, i_10_199_2079_0, i_10_199_2151_0, i_10_199_2166_0,
    i_10_199_2167_0, i_10_199_2304_0, i_10_199_2306_0, i_10_199_2307_0,
    i_10_199_2310_0, i_10_199_2333_0, i_10_199_2335_0, i_10_199_2357_0,
    i_10_199_2436_0, i_10_199_2475_0, i_10_199_2478_0, i_10_199_2511_0,
    i_10_199_2608_0, i_10_199_2614_0, i_10_199_2615_0, i_10_199_2628_0,
    i_10_199_2630_0, i_10_199_2638_0, i_10_199_2655_0, i_10_199_2658_0,
    i_10_199_2659_0, i_10_199_2700_0, i_10_199_2832_0, i_10_199_2871_0,
    i_10_199_2881_0, i_10_199_2916_0, i_10_199_2920_0, i_10_199_2923_0,
    i_10_199_2952_0, i_10_199_2953_0, i_10_199_3037_0, i_10_199_3038_0,
    i_10_199_3040_0, i_10_199_3055_0, i_10_199_3087_0, i_10_199_3204_0,
    i_10_199_3229_0, i_10_199_3356_0, i_10_199_3358_0, i_10_199_3560_0,
    i_10_199_3651_0, i_10_199_3682_0, i_10_199_3683_0, i_10_199_3684_0,
    i_10_199_3685_0, i_10_199_3774_0, i_10_199_3853_0, i_10_199_3889_0,
    i_10_199_3892_0, i_10_199_3894_0, i_10_199_3924_0, i_10_199_3984_0,
    i_10_199_4124_0, i_10_199_4192_0, i_10_199_4230_0, i_10_199_4231_0,
    i_10_199_4374_0, i_10_199_4375_0, i_10_199_4376_0, i_10_199_4580_0,
    o_10_199_0_0  );
  input  i_10_199_27_0, i_10_199_124_0, i_10_199_175_0, i_10_199_285_0,
    i_10_199_369_0, i_10_199_433_0, i_10_199_443_0, i_10_199_444_0,
    i_10_199_467_0, i_10_199_501_0, i_10_199_532_0, i_10_199_729_0,
    i_10_199_730_0, i_10_199_732_0, i_10_199_733_0, i_10_199_901_0,
    i_10_199_961_0, i_10_199_999_0, i_10_199_1052_0, i_10_199_1201_0,
    i_10_199_1263_0, i_10_199_1265_0, i_10_199_1270_0, i_10_199_1271_0,
    i_10_199_1308_0, i_10_199_1309_0, i_10_199_1353_0, i_10_199_1361_0,
    i_10_199_1363_0, i_10_199_1638_0, i_10_199_1741_0, i_10_199_1765_0,
    i_10_199_1823_0, i_10_199_1912_0, i_10_199_1947_0, i_10_199_1948_0,
    i_10_199_1957_0, i_10_199_2079_0, i_10_199_2151_0, i_10_199_2166_0,
    i_10_199_2167_0, i_10_199_2304_0, i_10_199_2306_0, i_10_199_2307_0,
    i_10_199_2310_0, i_10_199_2333_0, i_10_199_2335_0, i_10_199_2357_0,
    i_10_199_2436_0, i_10_199_2475_0, i_10_199_2478_0, i_10_199_2511_0,
    i_10_199_2608_0, i_10_199_2614_0, i_10_199_2615_0, i_10_199_2628_0,
    i_10_199_2630_0, i_10_199_2638_0, i_10_199_2655_0, i_10_199_2658_0,
    i_10_199_2659_0, i_10_199_2700_0, i_10_199_2832_0, i_10_199_2871_0,
    i_10_199_2881_0, i_10_199_2916_0, i_10_199_2920_0, i_10_199_2923_0,
    i_10_199_2952_0, i_10_199_2953_0, i_10_199_3037_0, i_10_199_3038_0,
    i_10_199_3040_0, i_10_199_3055_0, i_10_199_3087_0, i_10_199_3204_0,
    i_10_199_3229_0, i_10_199_3356_0, i_10_199_3358_0, i_10_199_3560_0,
    i_10_199_3651_0, i_10_199_3682_0, i_10_199_3683_0, i_10_199_3684_0,
    i_10_199_3685_0, i_10_199_3774_0, i_10_199_3853_0, i_10_199_3889_0,
    i_10_199_3892_0, i_10_199_3894_0, i_10_199_3924_0, i_10_199_3984_0,
    i_10_199_4124_0, i_10_199_4192_0, i_10_199_4230_0, i_10_199_4231_0,
    i_10_199_4374_0, i_10_199_4375_0, i_10_199_4376_0, i_10_199_4580_0;
  output o_10_199_0_0;
  assign o_10_199_0_0 = 0;
endmodule



// Benchmark "kernel_10_200" written by ABC on Sun Jul 19 10:24:28 2020

module kernel_10_200 ( 
    i_10_200_33_0, i_10_200_123_0, i_10_200_174_0, i_10_200_177_0,
    i_10_200_260_0, i_10_200_286_0, i_10_200_319_0, i_10_200_328_0,
    i_10_200_408_0, i_10_200_412_0, i_10_200_438_0, i_10_200_439_0,
    i_10_200_440_0, i_10_200_511_0, i_10_200_512_0, i_10_200_796_0,
    i_10_200_967_0, i_10_200_1003_0, i_10_200_1236_0, i_10_200_1239_0,
    i_10_200_1311_0, i_10_200_1439_0, i_10_200_1546_0, i_10_200_1619_0,
    i_10_200_1626_0, i_10_200_1627_0, i_10_200_1686_0, i_10_200_1689_0,
    i_10_200_1690_0, i_10_200_1691_0, i_10_200_1821_0, i_10_200_1822_0,
    i_10_200_1823_0, i_10_200_1986_0, i_10_200_1996_0, i_10_200_2031_0,
    i_10_200_2032_0, i_10_200_2361_0, i_10_200_2364_0, i_10_200_2407_0,
    i_10_200_2410_0, i_10_200_2451_0, i_10_200_2452_0, i_10_200_2455_0,
    i_10_200_2472_0, i_10_200_2473_0, i_10_200_2605_0, i_10_200_2634_0,
    i_10_200_2635_0, i_10_200_2636_0, i_10_200_2663_0, i_10_200_2704_0,
    i_10_200_2706_0, i_10_200_2713_0, i_10_200_2716_0, i_10_200_2717_0,
    i_10_200_2722_0, i_10_200_2733_0, i_10_200_2734_0, i_10_200_2788_0,
    i_10_200_2826_0, i_10_200_2827_0, i_10_200_2829_0, i_10_200_2830_0,
    i_10_200_2831_0, i_10_200_2833_0, i_10_200_2883_0, i_10_200_2884_0,
    i_10_200_2885_0, i_10_200_2985_0, i_10_200_2986_0, i_10_200_3049_0,
    i_10_200_3151_0, i_10_200_3202_0, i_10_200_3280_0, i_10_200_3283_0,
    i_10_200_3318_0, i_10_200_3325_0, i_10_200_3328_0, i_10_200_3391_0,
    i_10_200_3403_0, i_10_200_3525_0, i_10_200_3585_0, i_10_200_3615_0,
    i_10_200_3616_0, i_10_200_3617_0, i_10_200_3649_0, i_10_200_3653_0,
    i_10_200_3783_0, i_10_200_3786_0, i_10_200_3834_0, i_10_200_3835_0,
    i_10_200_3856_0, i_10_200_3858_0, i_10_200_3859_0, i_10_200_3912_0,
    i_10_200_3913_0, i_10_200_4281_0, i_10_200_4289_0, i_10_200_4571_0,
    o_10_200_0_0  );
  input  i_10_200_33_0, i_10_200_123_0, i_10_200_174_0, i_10_200_177_0,
    i_10_200_260_0, i_10_200_286_0, i_10_200_319_0, i_10_200_328_0,
    i_10_200_408_0, i_10_200_412_0, i_10_200_438_0, i_10_200_439_0,
    i_10_200_440_0, i_10_200_511_0, i_10_200_512_0, i_10_200_796_0,
    i_10_200_967_0, i_10_200_1003_0, i_10_200_1236_0, i_10_200_1239_0,
    i_10_200_1311_0, i_10_200_1439_0, i_10_200_1546_0, i_10_200_1619_0,
    i_10_200_1626_0, i_10_200_1627_0, i_10_200_1686_0, i_10_200_1689_0,
    i_10_200_1690_0, i_10_200_1691_0, i_10_200_1821_0, i_10_200_1822_0,
    i_10_200_1823_0, i_10_200_1986_0, i_10_200_1996_0, i_10_200_2031_0,
    i_10_200_2032_0, i_10_200_2361_0, i_10_200_2364_0, i_10_200_2407_0,
    i_10_200_2410_0, i_10_200_2451_0, i_10_200_2452_0, i_10_200_2455_0,
    i_10_200_2472_0, i_10_200_2473_0, i_10_200_2605_0, i_10_200_2634_0,
    i_10_200_2635_0, i_10_200_2636_0, i_10_200_2663_0, i_10_200_2704_0,
    i_10_200_2706_0, i_10_200_2713_0, i_10_200_2716_0, i_10_200_2717_0,
    i_10_200_2722_0, i_10_200_2733_0, i_10_200_2734_0, i_10_200_2788_0,
    i_10_200_2826_0, i_10_200_2827_0, i_10_200_2829_0, i_10_200_2830_0,
    i_10_200_2831_0, i_10_200_2833_0, i_10_200_2883_0, i_10_200_2884_0,
    i_10_200_2885_0, i_10_200_2985_0, i_10_200_2986_0, i_10_200_3049_0,
    i_10_200_3151_0, i_10_200_3202_0, i_10_200_3280_0, i_10_200_3283_0,
    i_10_200_3318_0, i_10_200_3325_0, i_10_200_3328_0, i_10_200_3391_0,
    i_10_200_3403_0, i_10_200_3525_0, i_10_200_3585_0, i_10_200_3615_0,
    i_10_200_3616_0, i_10_200_3617_0, i_10_200_3649_0, i_10_200_3653_0,
    i_10_200_3783_0, i_10_200_3786_0, i_10_200_3834_0, i_10_200_3835_0,
    i_10_200_3856_0, i_10_200_3858_0, i_10_200_3859_0, i_10_200_3912_0,
    i_10_200_3913_0, i_10_200_4281_0, i_10_200_4289_0, i_10_200_4571_0;
  output o_10_200_0_0;
  assign o_10_200_0_0 = ~((~i_10_200_177_0 & ((~i_10_200_1689_0 & ~i_10_200_1823_0 & ~i_10_200_2830_0 & ~i_10_200_3403_0 & i_10_200_3649_0) | (~i_10_200_174_0 & ~i_10_200_1691_0 & ~i_10_200_2722_0 & i_10_200_3280_0 & i_10_200_3856_0 & ~i_10_200_3912_0 & ~i_10_200_4289_0))) | (i_10_200_408_0 & ((~i_10_200_1686_0 & ~i_10_200_2722_0 & ~i_10_200_3049_0 & ~i_10_200_3283_0) | (~i_10_200_1823_0 & i_10_200_2713_0 & i_10_200_3856_0))) | (~i_10_200_1236_0 & ((~i_10_200_3283_0 & i_10_200_3617_0) | (~i_10_200_412_0 & ~i_10_200_1822_0 & ~i_10_200_2663_0 & ~i_10_200_2884_0 & ~i_10_200_3912_0 & ~i_10_200_4571_0))) | (~i_10_200_2032_0 & ((~i_10_200_408_0 & ~i_10_200_1626_0 & i_10_200_3653_0) | (~i_10_200_1689_0 & ~i_10_200_1823_0 & ~i_10_200_2451_0 & ~i_10_200_2883_0 & ~i_10_200_3912_0))) | (~i_10_200_1823_0 & ((~i_10_200_2472_0 & i_10_200_2634_0 & i_10_200_3858_0) | (~i_10_200_967_0 & ~i_10_200_2452_0 & ~i_10_200_2733_0 & ~i_10_200_3283_0 & ~i_10_200_3913_0))) | (~i_10_200_3283_0 & ((~i_10_200_967_0 & ~i_10_200_2452_0 & ((~i_10_200_1690_0 & ~i_10_200_3280_0) | (~i_10_200_2722_0 & ~i_10_200_3049_0 & ~i_10_200_3835_0))) | (~i_10_200_1822_0 & i_10_200_3856_0) | (~i_10_200_1546_0 & i_10_200_1691_0 & ~i_10_200_2663_0 & ~i_10_200_2885_0 & ~i_10_200_3783_0 & ~i_10_200_3913_0) | (i_10_200_1003_0 & ~i_10_200_2722_0 & ~i_10_200_2734_0 & ~i_10_200_4281_0))) | (~i_10_200_1821_0 & ((~i_10_200_967_0 & ((~i_10_200_260_0 & ~i_10_200_1003_0 & ~i_10_200_1689_0 & ~i_10_200_2473_0 & ~i_10_200_2716_0 & ~i_10_200_2722_0 & ~i_10_200_3049_0 & ~i_10_200_3403_0) | (i_10_200_2722_0 & ~i_10_200_3913_0 & ~i_10_200_4289_0))) | (~i_10_200_2031_0 & ~i_10_200_2472_0 & ~i_10_200_2716_0 & ~i_10_200_2884_0 & ~i_10_200_3049_0 & ~i_10_200_3403_0 & ~i_10_200_3912_0 & ~i_10_200_3913_0))) | (~i_10_200_2884_0 & ((~i_10_200_1689_0 & i_10_200_2704_0 & ~i_10_200_2986_0) | (~i_10_200_2883_0 & ~i_10_200_3280_0 & i_10_200_3783_0 & ~i_10_200_3913_0 & ~i_10_200_4289_0 & ~i_10_200_4571_0))) | (~i_10_200_4289_0 & ((~i_10_200_3585_0 & (i_10_200_2407_0 | (i_10_200_1823_0 & ~i_10_200_2885_0 & i_10_200_3649_0 & ~i_10_200_3783_0))) | (~i_10_200_796_0 & ~i_10_200_1689_0 & ~i_10_200_2451_0 & ~i_10_200_3391_0 & i_10_200_3649_0 & ~i_10_200_3653_0) | (~i_10_200_123_0 & ~i_10_200_2788_0 & ~i_10_200_3525_0 & i_10_200_3615_0 & ~i_10_200_3913_0))) | (~i_10_200_1689_0 & ((i_10_200_2451_0 & ~i_10_200_2713_0 & i_10_200_3617_0) | (~i_10_200_1439_0 & i_10_200_2635_0 & ~i_10_200_3318_0 & ~i_10_200_3913_0))) | (i_10_200_2827_0 & i_10_200_3403_0 & ~i_10_200_3835_0) | (i_10_200_2831_0 & i_10_200_4289_0));
endmodule



// Benchmark "kernel_10_201" written by ABC on Sun Jul 19 10:24:29 2020

module kernel_10_201 ( 
    i_10_201_24_0, i_10_201_33_0, i_10_201_184_0, i_10_201_283_0,
    i_10_201_320_0, i_10_201_323_0, i_10_201_330_0, i_10_201_332_0,
    i_10_201_393_0, i_10_201_394_0, i_10_201_436_0, i_10_201_440_0,
    i_10_201_444_0, i_10_201_461_0, i_10_201_500_0, i_10_201_503_0,
    i_10_201_696_0, i_10_201_732_0, i_10_201_733_0, i_10_201_734_0,
    i_10_201_931_0, i_10_201_952_0, i_10_201_1002_0, i_10_201_1043_0,
    i_10_201_1047_0, i_10_201_1348_0, i_10_201_1349_0, i_10_201_1482_0,
    i_10_201_1488_0, i_10_201_1528_0, i_10_201_1548_0, i_10_201_1551_0,
    i_10_201_1555_0, i_10_201_1556_0, i_10_201_1655_0, i_10_201_1686_0,
    i_10_201_1767_0, i_10_201_1768_0, i_10_201_1823_0, i_10_201_1869_0,
    i_10_201_1957_0, i_10_201_2003_0, i_10_201_2004_0, i_10_201_2029_0,
    i_10_201_2083_0, i_10_201_2088_0, i_10_201_2156_0, i_10_201_2186_0,
    i_10_201_2204_0, i_10_201_2212_0, i_10_201_2312_0, i_10_201_2382_0,
    i_10_201_2409_0, i_10_201_2453_0, i_10_201_2571_0, i_10_201_2631_0,
    i_10_201_2632_0, i_10_201_2636_0, i_10_201_2659_0, i_10_201_2721_0,
    i_10_201_2722_0, i_10_201_2761_0, i_10_201_2806_0, i_10_201_2917_0,
    i_10_201_2923_0, i_10_201_2956_0, i_10_201_2983_0, i_10_201_2987_0,
    i_10_201_3030_0, i_10_201_3041_0, i_10_201_3131_0, i_10_201_3275_0,
    i_10_201_3361_0, i_10_201_3362_0, i_10_201_3388_0, i_10_201_3537_0,
    i_10_201_3538_0, i_10_201_3554_0, i_10_201_3588_0, i_10_201_3605_0,
    i_10_201_3608_0, i_10_201_3612_0, i_10_201_3615_0, i_10_201_3616_0,
    i_10_201_3837_0, i_10_201_3856_0, i_10_201_3865_0, i_10_201_3981_0,
    i_10_201_3982_0, i_10_201_3984_0, i_10_201_3990_0, i_10_201_3991_0,
    i_10_201_3993_0, i_10_201_4287_0, i_10_201_4288_0, i_10_201_4289_0,
    i_10_201_4292_0, i_10_201_4372_0, i_10_201_4570_0, i_10_201_4571_0,
    o_10_201_0_0  );
  input  i_10_201_24_0, i_10_201_33_0, i_10_201_184_0, i_10_201_283_0,
    i_10_201_320_0, i_10_201_323_0, i_10_201_330_0, i_10_201_332_0,
    i_10_201_393_0, i_10_201_394_0, i_10_201_436_0, i_10_201_440_0,
    i_10_201_444_0, i_10_201_461_0, i_10_201_500_0, i_10_201_503_0,
    i_10_201_696_0, i_10_201_732_0, i_10_201_733_0, i_10_201_734_0,
    i_10_201_931_0, i_10_201_952_0, i_10_201_1002_0, i_10_201_1043_0,
    i_10_201_1047_0, i_10_201_1348_0, i_10_201_1349_0, i_10_201_1482_0,
    i_10_201_1488_0, i_10_201_1528_0, i_10_201_1548_0, i_10_201_1551_0,
    i_10_201_1555_0, i_10_201_1556_0, i_10_201_1655_0, i_10_201_1686_0,
    i_10_201_1767_0, i_10_201_1768_0, i_10_201_1823_0, i_10_201_1869_0,
    i_10_201_1957_0, i_10_201_2003_0, i_10_201_2004_0, i_10_201_2029_0,
    i_10_201_2083_0, i_10_201_2088_0, i_10_201_2156_0, i_10_201_2186_0,
    i_10_201_2204_0, i_10_201_2212_0, i_10_201_2312_0, i_10_201_2382_0,
    i_10_201_2409_0, i_10_201_2453_0, i_10_201_2571_0, i_10_201_2631_0,
    i_10_201_2632_0, i_10_201_2636_0, i_10_201_2659_0, i_10_201_2721_0,
    i_10_201_2722_0, i_10_201_2761_0, i_10_201_2806_0, i_10_201_2917_0,
    i_10_201_2923_0, i_10_201_2956_0, i_10_201_2983_0, i_10_201_2987_0,
    i_10_201_3030_0, i_10_201_3041_0, i_10_201_3131_0, i_10_201_3275_0,
    i_10_201_3361_0, i_10_201_3362_0, i_10_201_3388_0, i_10_201_3537_0,
    i_10_201_3538_0, i_10_201_3554_0, i_10_201_3588_0, i_10_201_3605_0,
    i_10_201_3608_0, i_10_201_3612_0, i_10_201_3615_0, i_10_201_3616_0,
    i_10_201_3837_0, i_10_201_3856_0, i_10_201_3865_0, i_10_201_3981_0,
    i_10_201_3982_0, i_10_201_3984_0, i_10_201_3990_0, i_10_201_3991_0,
    i_10_201_3993_0, i_10_201_4287_0, i_10_201_4288_0, i_10_201_4289_0,
    i_10_201_4292_0, i_10_201_4372_0, i_10_201_4570_0, i_10_201_4571_0;
  output o_10_201_0_0;
  assign o_10_201_0_0 = 0;
endmodule



// Benchmark "kernel_10_202" written by ABC on Sun Jul 19 10:24:30 2020

module kernel_10_202 ( 
    i_10_202_42_0, i_10_202_177_0, i_10_202_220_0, i_10_202_222_0,
    i_10_202_246_0, i_10_202_247_0, i_10_202_249_0, i_10_202_250_0,
    i_10_202_283_0, i_10_202_292_0, i_10_202_442_0, i_10_202_463_0,
    i_10_202_466_0, i_10_202_467_0, i_10_202_566_0, i_10_202_597_0,
    i_10_202_894_0, i_10_202_996_0, i_10_202_1032_0, i_10_202_1033_0,
    i_10_202_1141_0, i_10_202_1239_0, i_10_202_1241_0, i_10_202_1266_0,
    i_10_202_1444_0, i_10_202_1545_0, i_10_202_1578_0, i_10_202_1648_0,
    i_10_202_1653_0, i_10_202_1654_0, i_10_202_1825_0, i_10_202_2004_0,
    i_10_202_2019_0, i_10_202_2022_0, i_10_202_2351_0, i_10_202_2353_0,
    i_10_202_2359_0, i_10_202_2361_0, i_10_202_2364_0, i_10_202_2469_0,
    i_10_202_2470_0, i_10_202_2471_0, i_10_202_2472_0, i_10_202_2473_0,
    i_10_202_2604_0, i_10_202_2607_0, i_10_202_2632_0, i_10_202_2657_0,
    i_10_202_2658_0, i_10_202_2703_0, i_10_202_2704_0, i_10_202_2706_0,
    i_10_202_2721_0, i_10_202_2727_0, i_10_202_2731_0, i_10_202_2781_0,
    i_10_202_2826_0, i_10_202_2833_0, i_10_202_2917_0, i_10_202_3033_0,
    i_10_202_3043_0, i_10_202_3045_0, i_10_202_3072_0, i_10_202_3075_0,
    i_10_202_3158_0, i_10_202_3162_0, i_10_202_3267_0, i_10_202_3270_0,
    i_10_202_3278_0, i_10_202_3279_0, i_10_202_3280_0, i_10_202_3388_0,
    i_10_202_3406_0, i_10_202_3430_0, i_10_202_3493_0, i_10_202_3652_0,
    i_10_202_3684_0, i_10_202_3687_0, i_10_202_3782_0, i_10_202_3787_0,
    i_10_202_3810_0, i_10_202_3811_0, i_10_202_3813_0, i_10_202_3839_0,
    i_10_202_3846_0, i_10_202_3855_0, i_10_202_3858_0, i_10_202_4116_0,
    i_10_202_4117_0, i_10_202_4119_0, i_10_202_4125_0, i_10_202_4128_0,
    i_10_202_4129_0, i_10_202_4215_0, i_10_202_4218_0, i_10_202_4289_0,
    i_10_202_4291_0, i_10_202_4292_0, i_10_202_4564_0, i_10_202_4567_0,
    o_10_202_0_0  );
  input  i_10_202_42_0, i_10_202_177_0, i_10_202_220_0, i_10_202_222_0,
    i_10_202_246_0, i_10_202_247_0, i_10_202_249_0, i_10_202_250_0,
    i_10_202_283_0, i_10_202_292_0, i_10_202_442_0, i_10_202_463_0,
    i_10_202_466_0, i_10_202_467_0, i_10_202_566_0, i_10_202_597_0,
    i_10_202_894_0, i_10_202_996_0, i_10_202_1032_0, i_10_202_1033_0,
    i_10_202_1141_0, i_10_202_1239_0, i_10_202_1241_0, i_10_202_1266_0,
    i_10_202_1444_0, i_10_202_1545_0, i_10_202_1578_0, i_10_202_1648_0,
    i_10_202_1653_0, i_10_202_1654_0, i_10_202_1825_0, i_10_202_2004_0,
    i_10_202_2019_0, i_10_202_2022_0, i_10_202_2351_0, i_10_202_2353_0,
    i_10_202_2359_0, i_10_202_2361_0, i_10_202_2364_0, i_10_202_2469_0,
    i_10_202_2470_0, i_10_202_2471_0, i_10_202_2472_0, i_10_202_2473_0,
    i_10_202_2604_0, i_10_202_2607_0, i_10_202_2632_0, i_10_202_2657_0,
    i_10_202_2658_0, i_10_202_2703_0, i_10_202_2704_0, i_10_202_2706_0,
    i_10_202_2721_0, i_10_202_2727_0, i_10_202_2731_0, i_10_202_2781_0,
    i_10_202_2826_0, i_10_202_2833_0, i_10_202_2917_0, i_10_202_3033_0,
    i_10_202_3043_0, i_10_202_3045_0, i_10_202_3072_0, i_10_202_3075_0,
    i_10_202_3158_0, i_10_202_3162_0, i_10_202_3267_0, i_10_202_3270_0,
    i_10_202_3278_0, i_10_202_3279_0, i_10_202_3280_0, i_10_202_3388_0,
    i_10_202_3406_0, i_10_202_3430_0, i_10_202_3493_0, i_10_202_3652_0,
    i_10_202_3684_0, i_10_202_3687_0, i_10_202_3782_0, i_10_202_3787_0,
    i_10_202_3810_0, i_10_202_3811_0, i_10_202_3813_0, i_10_202_3839_0,
    i_10_202_3846_0, i_10_202_3855_0, i_10_202_3858_0, i_10_202_4116_0,
    i_10_202_4117_0, i_10_202_4119_0, i_10_202_4125_0, i_10_202_4128_0,
    i_10_202_4129_0, i_10_202_4215_0, i_10_202_4218_0, i_10_202_4289_0,
    i_10_202_4291_0, i_10_202_4292_0, i_10_202_4564_0, i_10_202_4567_0;
  output o_10_202_0_0;
  assign o_10_202_0_0 = ~((~i_10_202_3162_0 & ((~i_10_202_246_0 & ((~i_10_202_894_0 & ~i_10_202_996_0 & ~i_10_202_3684_0 & ~i_10_202_3687_0 & ~i_10_202_4119_0) | (~i_10_202_1033_0 & ~i_10_202_1648_0 & ~i_10_202_2351_0 & ~i_10_202_2607_0 & ~i_10_202_3045_0 & ~i_10_202_3267_0 & ~i_10_202_4128_0 & ~i_10_202_4218_0))) | (~i_10_202_250_0 & ~i_10_202_1545_0 & ~i_10_202_2781_0 & ~i_10_202_3075_0 & ~i_10_202_3430_0 & ~i_10_202_3684_0 & i_10_202_4117_0) | (~i_10_202_249_0 & ~i_10_202_2019_0 & ~i_10_202_2607_0 & ~i_10_202_3072_0 & ~i_10_202_4215_0 & ~i_10_202_4218_0) | (~i_10_202_996_0 & ~i_10_202_1032_0 & ~i_10_202_2826_0 & ~i_10_202_3033_0 & i_10_202_3267_0 & ~i_10_202_4129_0 & ~i_10_202_4564_0))) | (~i_10_202_247_0 & ((~i_10_202_442_0 & ~i_10_202_2359_0 & ~i_10_202_2361_0 & ~i_10_202_2607_0 & ~i_10_202_3684_0) | (i_10_202_283_0 & ~i_10_202_292_0 & ~i_10_202_463_0 & ~i_10_202_1654_0 & ~i_10_202_2353_0 & ~i_10_202_3072_0 & ~i_10_202_3687_0 & ~i_10_202_4128_0))) | (~i_10_202_2604_0 & ((~i_10_202_466_0 & ((~i_10_202_566_0 & ~i_10_202_996_0 & ~i_10_202_1654_0 & ~i_10_202_2607_0 & ~i_10_202_2632_0 & ~i_10_202_2833_0 & ~i_10_202_2917_0 & ~i_10_202_3270_0 & ~i_10_202_3279_0 & ~i_10_202_3430_0) | (~i_10_202_463_0 & ~i_10_202_2359_0 & ~i_10_202_2658_0 & ~i_10_202_3787_0 & ~i_10_202_4129_0 & ~i_10_202_4289_0 & ~i_10_202_4564_0))) | (~i_10_202_222_0 & ~i_10_202_2703_0 & ~i_10_202_3270_0 & ~i_10_202_4218_0 & ~i_10_202_4567_0))) | (~i_10_202_2607_0 & ~i_10_202_2706_0 & ((~i_10_202_292_0 & ~i_10_202_1032_0 & ~i_10_202_2359_0 & i_10_202_2632_0 & ~i_10_202_3430_0 & ~i_10_202_3684_0 & ~i_10_202_3782_0) | (~i_10_202_1266_0 & ~i_10_202_1444_0 & ~i_10_202_2361_0 & ~i_10_202_3687_0 & ~i_10_202_3787_0))) | (~i_10_202_3430_0 & ((~i_10_202_1648_0 & ~i_10_202_2658_0 & i_10_202_2731_0 & ~i_10_202_3652_0) | (~i_10_202_4215_0 & ~i_10_202_4218_0 & ~i_10_202_250_0 & ~i_10_202_4116_0))) | (~i_10_202_442_0 & ~i_10_202_2472_0 & ~i_10_202_2727_0 & ~i_10_202_3033_0 & ~i_10_202_3687_0 & ~i_10_202_3846_0 & ~i_10_202_4119_0 & ~i_10_202_4215_0) | (~i_10_202_249_0 & i_10_202_463_0 & ~i_10_202_3045_0 & ~i_10_202_3267_0 & i_10_202_3839_0 & i_10_202_4129_0));
endmodule



// Benchmark "kernel_10_203" written by ABC on Sun Jul 19 10:24:31 2020

module kernel_10_203 ( 
    i_10_203_34_0, i_10_203_176_0, i_10_203_221_0, i_10_203_254_0,
    i_10_203_280_0, i_10_203_328_0, i_10_203_374_0, i_10_203_394_0,
    i_10_203_445_0, i_10_203_446_0, i_10_203_715_0, i_10_203_718_0,
    i_10_203_754_0, i_10_203_792_0, i_10_203_797_0, i_10_203_798_0,
    i_10_203_829_0, i_10_203_830_0, i_10_203_832_0, i_10_203_957_0,
    i_10_203_959_0, i_10_203_1012_0, i_10_203_1031_0, i_10_203_1119_0,
    i_10_203_1234_0, i_10_203_1235_0, i_10_203_1313_0, i_10_203_1544_0,
    i_10_203_1578_0, i_10_203_1579_0, i_10_203_1683_0, i_10_203_1687_0,
    i_10_203_1814_0, i_10_203_1819_0, i_10_203_1820_0, i_10_203_1823_0,
    i_10_203_1919_0, i_10_203_1939_0, i_10_203_2026_0, i_10_203_2178_0,
    i_10_203_2179_0, i_10_203_2309_0, i_10_203_2311_0, i_10_203_2350_0,
    i_10_203_2353_0, i_10_203_2354_0, i_10_203_2365_0, i_10_203_2380_0,
    i_10_203_2404_0, i_10_203_2569_0, i_10_203_2708_0, i_10_203_2721_0,
    i_10_203_2722_0, i_10_203_2731_0, i_10_203_2783_0, i_10_203_2785_0,
    i_10_203_2834_0, i_10_203_3011_0, i_10_203_3099_0, i_10_203_3200_0,
    i_10_203_3202_0, i_10_203_3236_0, i_10_203_3239_0, i_10_203_3275_0,
    i_10_203_3298_0, i_10_203_3352_0, i_10_203_3386_0, i_10_203_3389_0,
    i_10_203_3493_0, i_10_203_3494_0, i_10_203_3542_0, i_10_203_3581_0,
    i_10_203_3583_0, i_10_203_3584_0, i_10_203_3615_0, i_10_203_3616_0,
    i_10_203_3617_0, i_10_203_3636_0, i_10_203_3650_0, i_10_203_3653_0,
    i_10_203_3711_0, i_10_203_3724_0, i_10_203_3781_0, i_10_203_3782_0,
    i_10_203_3783_0, i_10_203_3784_0, i_10_203_3785_0, i_10_203_3786_0,
    i_10_203_3787_0, i_10_203_3788_0, i_10_203_3809_0, i_10_203_3860_0,
    i_10_203_3947_0, i_10_203_4024_0, i_10_203_4118_0, i_10_203_4120_0,
    i_10_203_4121_0, i_10_203_4130_0, i_10_203_4175_0, i_10_203_4214_0,
    o_10_203_0_0  );
  input  i_10_203_34_0, i_10_203_176_0, i_10_203_221_0, i_10_203_254_0,
    i_10_203_280_0, i_10_203_328_0, i_10_203_374_0, i_10_203_394_0,
    i_10_203_445_0, i_10_203_446_0, i_10_203_715_0, i_10_203_718_0,
    i_10_203_754_0, i_10_203_792_0, i_10_203_797_0, i_10_203_798_0,
    i_10_203_829_0, i_10_203_830_0, i_10_203_832_0, i_10_203_957_0,
    i_10_203_959_0, i_10_203_1012_0, i_10_203_1031_0, i_10_203_1119_0,
    i_10_203_1234_0, i_10_203_1235_0, i_10_203_1313_0, i_10_203_1544_0,
    i_10_203_1578_0, i_10_203_1579_0, i_10_203_1683_0, i_10_203_1687_0,
    i_10_203_1814_0, i_10_203_1819_0, i_10_203_1820_0, i_10_203_1823_0,
    i_10_203_1919_0, i_10_203_1939_0, i_10_203_2026_0, i_10_203_2178_0,
    i_10_203_2179_0, i_10_203_2309_0, i_10_203_2311_0, i_10_203_2350_0,
    i_10_203_2353_0, i_10_203_2354_0, i_10_203_2365_0, i_10_203_2380_0,
    i_10_203_2404_0, i_10_203_2569_0, i_10_203_2708_0, i_10_203_2721_0,
    i_10_203_2722_0, i_10_203_2731_0, i_10_203_2783_0, i_10_203_2785_0,
    i_10_203_2834_0, i_10_203_3011_0, i_10_203_3099_0, i_10_203_3200_0,
    i_10_203_3202_0, i_10_203_3236_0, i_10_203_3239_0, i_10_203_3275_0,
    i_10_203_3298_0, i_10_203_3352_0, i_10_203_3386_0, i_10_203_3389_0,
    i_10_203_3493_0, i_10_203_3494_0, i_10_203_3542_0, i_10_203_3581_0,
    i_10_203_3583_0, i_10_203_3584_0, i_10_203_3615_0, i_10_203_3616_0,
    i_10_203_3617_0, i_10_203_3636_0, i_10_203_3650_0, i_10_203_3653_0,
    i_10_203_3711_0, i_10_203_3724_0, i_10_203_3781_0, i_10_203_3782_0,
    i_10_203_3783_0, i_10_203_3784_0, i_10_203_3785_0, i_10_203_3786_0,
    i_10_203_3787_0, i_10_203_3788_0, i_10_203_3809_0, i_10_203_3860_0,
    i_10_203_3947_0, i_10_203_4024_0, i_10_203_4118_0, i_10_203_4120_0,
    i_10_203_4121_0, i_10_203_4130_0, i_10_203_4175_0, i_10_203_4214_0;
  output o_10_203_0_0;
  assign o_10_203_0_0 = 0;
endmodule



// Benchmark "kernel_10_204" written by ABC on Sun Jul 19 10:24:32 2020

module kernel_10_204 ( 
    i_10_204_17_0, i_10_204_68_0, i_10_204_134_0, i_10_204_152_0,
    i_10_204_170_0, i_10_204_223_0, i_10_204_239_0, i_10_204_275_0,
    i_10_204_331_0, i_10_204_373_0, i_10_204_376_0, i_10_204_392_0,
    i_10_204_440_0, i_10_204_445_0, i_10_204_446_0, i_10_204_447_0,
    i_10_204_462_0, i_10_204_518_0, i_10_204_548_0, i_10_204_637_0,
    i_10_204_718_0, i_10_204_719_0, i_10_204_737_0, i_10_204_799_0,
    i_10_204_950_0, i_10_204_989_0, i_10_204_1166_0, i_10_204_1245_0,
    i_10_204_1246_0, i_10_204_1267_0, i_10_204_1312_0, i_10_204_1313_0,
    i_10_204_1438_0, i_10_204_1491_0, i_10_204_1493_0, i_10_204_1538_0,
    i_10_204_1539_0, i_10_204_1583_0, i_10_204_1616_0, i_10_204_1637_0,
    i_10_204_1643_0, i_10_204_1646_0, i_10_204_1651_0, i_10_204_1653_0,
    i_10_204_1691_0, i_10_204_1824_0, i_10_204_1873_0, i_10_204_1940_0,
    i_10_204_1942_0, i_10_204_1951_0, i_10_204_1961_0, i_10_204_2032_0,
    i_10_204_2069_0, i_10_204_2183_0, i_10_204_2231_0, i_10_204_2326_0,
    i_10_204_2330_0, i_10_204_2359_0, i_10_204_2452_0, i_10_204_2474_0,
    i_10_204_2521_0, i_10_204_2535_0, i_10_204_2636_0, i_10_204_2663_0,
    i_10_204_2672_0, i_10_204_2705_0, i_10_204_2865_0, i_10_204_2883_0,
    i_10_204_2884_0, i_10_204_2986_0, i_10_204_2987_0, i_10_204_3072_0,
    i_10_204_3075_0, i_10_204_3122_0, i_10_204_3195_0, i_10_204_3199_0,
    i_10_204_3356_0, i_10_204_3455_0, i_10_204_3469_0, i_10_204_3495_0,
    i_10_204_3509_0, i_10_204_3590_0, i_10_204_3617_0, i_10_204_3650_0,
    i_10_204_3788_0, i_10_204_3801_0, i_10_204_3804_0, i_10_204_3860_0,
    i_10_204_3877_0, i_10_204_3878_0, i_10_204_3910_0, i_10_204_3950_0,
    i_10_204_3991_0, i_10_204_3994_0, i_10_204_3995_0, i_10_204_4138_0,
    i_10_204_4154_0, i_10_204_4183_0, i_10_204_4288_0, i_10_204_4291_0,
    o_10_204_0_0  );
  input  i_10_204_17_0, i_10_204_68_0, i_10_204_134_0, i_10_204_152_0,
    i_10_204_170_0, i_10_204_223_0, i_10_204_239_0, i_10_204_275_0,
    i_10_204_331_0, i_10_204_373_0, i_10_204_376_0, i_10_204_392_0,
    i_10_204_440_0, i_10_204_445_0, i_10_204_446_0, i_10_204_447_0,
    i_10_204_462_0, i_10_204_518_0, i_10_204_548_0, i_10_204_637_0,
    i_10_204_718_0, i_10_204_719_0, i_10_204_737_0, i_10_204_799_0,
    i_10_204_950_0, i_10_204_989_0, i_10_204_1166_0, i_10_204_1245_0,
    i_10_204_1246_0, i_10_204_1267_0, i_10_204_1312_0, i_10_204_1313_0,
    i_10_204_1438_0, i_10_204_1491_0, i_10_204_1493_0, i_10_204_1538_0,
    i_10_204_1539_0, i_10_204_1583_0, i_10_204_1616_0, i_10_204_1637_0,
    i_10_204_1643_0, i_10_204_1646_0, i_10_204_1651_0, i_10_204_1653_0,
    i_10_204_1691_0, i_10_204_1824_0, i_10_204_1873_0, i_10_204_1940_0,
    i_10_204_1942_0, i_10_204_1951_0, i_10_204_1961_0, i_10_204_2032_0,
    i_10_204_2069_0, i_10_204_2183_0, i_10_204_2231_0, i_10_204_2326_0,
    i_10_204_2330_0, i_10_204_2359_0, i_10_204_2452_0, i_10_204_2474_0,
    i_10_204_2521_0, i_10_204_2535_0, i_10_204_2636_0, i_10_204_2663_0,
    i_10_204_2672_0, i_10_204_2705_0, i_10_204_2865_0, i_10_204_2883_0,
    i_10_204_2884_0, i_10_204_2986_0, i_10_204_2987_0, i_10_204_3072_0,
    i_10_204_3075_0, i_10_204_3122_0, i_10_204_3195_0, i_10_204_3199_0,
    i_10_204_3356_0, i_10_204_3455_0, i_10_204_3469_0, i_10_204_3495_0,
    i_10_204_3509_0, i_10_204_3590_0, i_10_204_3617_0, i_10_204_3650_0,
    i_10_204_3788_0, i_10_204_3801_0, i_10_204_3804_0, i_10_204_3860_0,
    i_10_204_3877_0, i_10_204_3878_0, i_10_204_3910_0, i_10_204_3950_0,
    i_10_204_3991_0, i_10_204_3994_0, i_10_204_3995_0, i_10_204_4138_0,
    i_10_204_4154_0, i_10_204_4183_0, i_10_204_4288_0, i_10_204_4291_0;
  output o_10_204_0_0;
  assign o_10_204_0_0 = 0;
endmodule



// Benchmark "kernel_10_205" written by ABC on Sun Jul 19 10:24:33 2020

module kernel_10_205 ( 
    i_10_205_39_0, i_10_205_159_0, i_10_205_251_0, i_10_205_282_0,
    i_10_205_284_0, i_10_205_292_0, i_10_205_296_0, i_10_205_320_0,
    i_10_205_328_0, i_10_205_329_0, i_10_205_368_0, i_10_205_394_0,
    i_10_205_411_0, i_10_205_412_0, i_10_205_413_0, i_10_205_439_0,
    i_10_205_440_0, i_10_205_444_0, i_10_205_447_0, i_10_205_448_0,
    i_10_205_449_0, i_10_205_512_0, i_10_205_800_0, i_10_205_962_0,
    i_10_205_1015_0, i_10_205_1016_0, i_10_205_1034_0, i_10_205_1221_0,
    i_10_205_1222_0, i_10_205_1237_0, i_10_205_1346_0, i_10_205_1348_0,
    i_10_205_1687_0, i_10_205_1688_0, i_10_205_1690_0, i_10_205_1691_0,
    i_10_205_1729_0, i_10_205_1730_0, i_10_205_1733_0, i_10_205_1984_0,
    i_10_205_2003_0, i_10_205_2006_0, i_10_205_2030_0, i_10_205_2357_0,
    i_10_205_2383_0, i_10_205_2384_0, i_10_205_2450_0, i_10_205_2454_0,
    i_10_205_2455_0, i_10_205_2456_0, i_10_205_2464_0, i_10_205_2471_0,
    i_10_205_2512_0, i_10_205_2516_0, i_10_205_2536_0, i_10_205_2537_0,
    i_10_205_2571_0, i_10_205_2601_0, i_10_205_2604_0, i_10_205_2673_0,
    i_10_205_2676_0, i_10_205_2704_0, i_10_205_2714_0, i_10_205_2716_0,
    i_10_205_2717_0, i_10_205_2728_0, i_10_205_2734_0, i_10_205_2743_0,
    i_10_205_2788_0, i_10_205_2831_0, i_10_205_2833_0, i_10_205_2834_0,
    i_10_205_2885_0, i_10_205_2969_0, i_10_205_2980_0, i_10_205_3199_0,
    i_10_205_3278_0, i_10_205_3281_0, i_10_205_3301_0, i_10_205_3506_0,
    i_10_205_3551_0, i_10_205_3561_0, i_10_205_3562_0, i_10_205_3586_0,
    i_10_205_3587_0, i_10_205_3590_0, i_10_205_3613_0, i_10_205_3614_0,
    i_10_205_3616_0, i_10_205_3784_0, i_10_205_3787_0, i_10_205_3840_0,
    i_10_205_3913_0, i_10_205_3983_0, i_10_205_4120_0, i_10_205_4155_0,
    i_10_205_4277_0, i_10_205_4291_0, i_10_205_4292_0, i_10_205_4567_0,
    o_10_205_0_0  );
  input  i_10_205_39_0, i_10_205_159_0, i_10_205_251_0, i_10_205_282_0,
    i_10_205_284_0, i_10_205_292_0, i_10_205_296_0, i_10_205_320_0,
    i_10_205_328_0, i_10_205_329_0, i_10_205_368_0, i_10_205_394_0,
    i_10_205_411_0, i_10_205_412_0, i_10_205_413_0, i_10_205_439_0,
    i_10_205_440_0, i_10_205_444_0, i_10_205_447_0, i_10_205_448_0,
    i_10_205_449_0, i_10_205_512_0, i_10_205_800_0, i_10_205_962_0,
    i_10_205_1015_0, i_10_205_1016_0, i_10_205_1034_0, i_10_205_1221_0,
    i_10_205_1222_0, i_10_205_1237_0, i_10_205_1346_0, i_10_205_1348_0,
    i_10_205_1687_0, i_10_205_1688_0, i_10_205_1690_0, i_10_205_1691_0,
    i_10_205_1729_0, i_10_205_1730_0, i_10_205_1733_0, i_10_205_1984_0,
    i_10_205_2003_0, i_10_205_2006_0, i_10_205_2030_0, i_10_205_2357_0,
    i_10_205_2383_0, i_10_205_2384_0, i_10_205_2450_0, i_10_205_2454_0,
    i_10_205_2455_0, i_10_205_2456_0, i_10_205_2464_0, i_10_205_2471_0,
    i_10_205_2512_0, i_10_205_2516_0, i_10_205_2536_0, i_10_205_2537_0,
    i_10_205_2571_0, i_10_205_2601_0, i_10_205_2604_0, i_10_205_2673_0,
    i_10_205_2676_0, i_10_205_2704_0, i_10_205_2714_0, i_10_205_2716_0,
    i_10_205_2717_0, i_10_205_2728_0, i_10_205_2734_0, i_10_205_2743_0,
    i_10_205_2788_0, i_10_205_2831_0, i_10_205_2833_0, i_10_205_2834_0,
    i_10_205_2885_0, i_10_205_2969_0, i_10_205_2980_0, i_10_205_3199_0,
    i_10_205_3278_0, i_10_205_3281_0, i_10_205_3301_0, i_10_205_3506_0,
    i_10_205_3551_0, i_10_205_3561_0, i_10_205_3562_0, i_10_205_3586_0,
    i_10_205_3587_0, i_10_205_3590_0, i_10_205_3613_0, i_10_205_3614_0,
    i_10_205_3616_0, i_10_205_3784_0, i_10_205_3787_0, i_10_205_3840_0,
    i_10_205_3913_0, i_10_205_3983_0, i_10_205_4120_0, i_10_205_4155_0,
    i_10_205_4277_0, i_10_205_4291_0, i_10_205_4292_0, i_10_205_4567_0;
  output o_10_205_0_0;
  assign o_10_205_0_0 = 0;
endmodule



// Benchmark "kernel_10_206" written by ABC on Sun Jul 19 10:24:33 2020

module kernel_10_206 ( 
    i_10_206_152_0, i_10_206_172_0, i_10_206_222_0, i_10_206_268_0,
    i_10_206_280_0, i_10_206_284_0, i_10_206_285_0, i_10_206_392_0,
    i_10_206_409_0, i_10_206_413_0, i_10_206_431_0, i_10_206_439_0,
    i_10_206_565_0, i_10_206_751_0, i_10_206_754_0, i_10_206_755_0,
    i_10_206_799_0, i_10_206_899_0, i_10_206_954_0, i_10_206_957_0,
    i_10_206_958_0, i_10_206_967_0, i_10_206_1032_0, i_10_206_1033_0,
    i_10_206_1236_0, i_10_206_1238_0, i_10_206_1242_0, i_10_206_1243_0,
    i_10_206_1244_0, i_10_206_1245_0, i_10_206_1249_0, i_10_206_1306_0,
    i_10_206_1345_0, i_10_206_1360_0, i_10_206_1366_0, i_10_206_1549_0,
    i_10_206_1683_0, i_10_206_1823_0, i_10_206_1825_0, i_10_206_1913_0,
    i_10_206_1916_0, i_10_206_1949_0, i_10_206_1952_0, i_10_206_1997_0,
    i_10_206_2311_0, i_10_206_2353_0, i_10_206_2364_0, i_10_206_2410_0,
    i_10_206_2450_0, i_10_206_2457_0, i_10_206_2470_0, i_10_206_2472_0,
    i_10_206_2474_0, i_10_206_2513_0, i_10_206_2705_0, i_10_206_2725_0,
    i_10_206_2735_0, i_10_206_2830_0, i_10_206_2834_0, i_10_206_2917_0,
    i_10_206_2919_0, i_10_206_2923_0, i_10_206_2924_0, i_10_206_2992_0,
    i_10_206_3037_0, i_10_206_3038_0, i_10_206_3039_0, i_10_206_3091_0,
    i_10_206_3199_0, i_10_206_3200_0, i_10_206_3270_0, i_10_206_3283_0,
    i_10_206_3388_0, i_10_206_3525_0, i_10_206_3563_0, i_10_206_3615_0,
    i_10_206_3617_0, i_10_206_3651_0, i_10_206_3780_0, i_10_206_3783_0,
    i_10_206_3784_0, i_10_206_3786_0, i_10_206_3787_0, i_10_206_3788_0,
    i_10_206_3844_0, i_10_206_3847_0, i_10_206_3854_0, i_10_206_3859_0,
    i_10_206_3982_0, i_10_206_3983_0, i_10_206_3986_0, i_10_206_3994_0,
    i_10_206_4116_0, i_10_206_4117_0, i_10_206_4118_0, i_10_206_4267_0,
    i_10_206_4273_0, i_10_206_4564_0, i_10_206_4571_0, i_10_206_4597_0,
    o_10_206_0_0  );
  input  i_10_206_152_0, i_10_206_172_0, i_10_206_222_0, i_10_206_268_0,
    i_10_206_280_0, i_10_206_284_0, i_10_206_285_0, i_10_206_392_0,
    i_10_206_409_0, i_10_206_413_0, i_10_206_431_0, i_10_206_439_0,
    i_10_206_565_0, i_10_206_751_0, i_10_206_754_0, i_10_206_755_0,
    i_10_206_799_0, i_10_206_899_0, i_10_206_954_0, i_10_206_957_0,
    i_10_206_958_0, i_10_206_967_0, i_10_206_1032_0, i_10_206_1033_0,
    i_10_206_1236_0, i_10_206_1238_0, i_10_206_1242_0, i_10_206_1243_0,
    i_10_206_1244_0, i_10_206_1245_0, i_10_206_1249_0, i_10_206_1306_0,
    i_10_206_1345_0, i_10_206_1360_0, i_10_206_1366_0, i_10_206_1549_0,
    i_10_206_1683_0, i_10_206_1823_0, i_10_206_1825_0, i_10_206_1913_0,
    i_10_206_1916_0, i_10_206_1949_0, i_10_206_1952_0, i_10_206_1997_0,
    i_10_206_2311_0, i_10_206_2353_0, i_10_206_2364_0, i_10_206_2410_0,
    i_10_206_2450_0, i_10_206_2457_0, i_10_206_2470_0, i_10_206_2472_0,
    i_10_206_2474_0, i_10_206_2513_0, i_10_206_2705_0, i_10_206_2725_0,
    i_10_206_2735_0, i_10_206_2830_0, i_10_206_2834_0, i_10_206_2917_0,
    i_10_206_2919_0, i_10_206_2923_0, i_10_206_2924_0, i_10_206_2992_0,
    i_10_206_3037_0, i_10_206_3038_0, i_10_206_3039_0, i_10_206_3091_0,
    i_10_206_3199_0, i_10_206_3200_0, i_10_206_3270_0, i_10_206_3283_0,
    i_10_206_3388_0, i_10_206_3525_0, i_10_206_3563_0, i_10_206_3615_0,
    i_10_206_3617_0, i_10_206_3651_0, i_10_206_3780_0, i_10_206_3783_0,
    i_10_206_3784_0, i_10_206_3786_0, i_10_206_3787_0, i_10_206_3788_0,
    i_10_206_3844_0, i_10_206_3847_0, i_10_206_3854_0, i_10_206_3859_0,
    i_10_206_3982_0, i_10_206_3983_0, i_10_206_3986_0, i_10_206_3994_0,
    i_10_206_4116_0, i_10_206_4117_0, i_10_206_4118_0, i_10_206_4267_0,
    i_10_206_4273_0, i_10_206_4564_0, i_10_206_4571_0, i_10_206_4597_0;
  output o_10_206_0_0;
  assign o_10_206_0_0 = 0;
endmodule



// Benchmark "kernel_10_207" written by ABC on Sun Jul 19 10:24:34 2020

module kernel_10_207 ( 
    i_10_207_171_0, i_10_207_178_0, i_10_207_179_0, i_10_207_253_0,
    i_10_207_328_0, i_10_207_329_0, i_10_207_364_0, i_10_207_409_0,
    i_10_207_410_0, i_10_207_443_0, i_10_207_444_0, i_10_207_462_0,
    i_10_207_463_0, i_10_207_466_0, i_10_207_960_0, i_10_207_962_0,
    i_10_207_1032_0, i_10_207_1033_0, i_10_207_1034_0, i_10_207_1165_0,
    i_10_207_1233_0, i_10_207_1242_0, i_10_207_1296_0, i_10_207_1307_0,
    i_10_207_1431_0, i_10_207_1432_0, i_10_207_1443_0, i_10_207_1444_0,
    i_10_207_1539_0, i_10_207_1576_0, i_10_207_1683_0, i_10_207_1686_0,
    i_10_207_1728_0, i_10_207_1818_0, i_10_207_1819_0, i_10_207_2021_0,
    i_10_207_2223_0, i_10_207_2352_0, i_10_207_2359_0, i_10_207_2361_0,
    i_10_207_2364_0, i_10_207_2431_0, i_10_207_2442_0, i_10_207_2449_0,
    i_10_207_2450_0, i_10_207_2451_0, i_10_207_2454_0, i_10_207_2628_0,
    i_10_207_2629_0, i_10_207_2655_0, i_10_207_2658_0, i_10_207_2659_0,
    i_10_207_2661_0, i_10_207_2681_0, i_10_207_2701_0, i_10_207_2714_0,
    i_10_207_2727_0, i_10_207_2784_0, i_10_207_2862_0, i_10_207_2916_0,
    i_10_207_3038_0, i_10_207_3074_0, i_10_207_3267_0, i_10_207_3271_0,
    i_10_207_3277_0, i_10_207_3279_0, i_10_207_3280_0, i_10_207_3282_0,
    i_10_207_3316_0, i_10_207_3331_0, i_10_207_3349_0, i_10_207_3450_0,
    i_10_207_3497_0, i_10_207_3537_0, i_10_207_3538_0, i_10_207_3614_0,
    i_10_207_3617_0, i_10_207_3650_0, i_10_207_3786_0, i_10_207_3787_0,
    i_10_207_3834_0, i_10_207_3846_0, i_10_207_3854_0, i_10_207_4116_0,
    i_10_207_4119_0, i_10_207_4171_0, i_10_207_4172_0, i_10_207_4204_0,
    i_10_207_4219_0, i_10_207_4267_0, i_10_207_4269_0, i_10_207_4270_0,
    i_10_207_4279_0, i_10_207_4284_0, i_10_207_4285_0, i_10_207_4288_0,
    i_10_207_4428_0, i_10_207_4459_0, i_10_207_4582_0, i_10_207_4591_0,
    o_10_207_0_0  );
  input  i_10_207_171_0, i_10_207_178_0, i_10_207_179_0, i_10_207_253_0,
    i_10_207_328_0, i_10_207_329_0, i_10_207_364_0, i_10_207_409_0,
    i_10_207_410_0, i_10_207_443_0, i_10_207_444_0, i_10_207_462_0,
    i_10_207_463_0, i_10_207_466_0, i_10_207_960_0, i_10_207_962_0,
    i_10_207_1032_0, i_10_207_1033_0, i_10_207_1034_0, i_10_207_1165_0,
    i_10_207_1233_0, i_10_207_1242_0, i_10_207_1296_0, i_10_207_1307_0,
    i_10_207_1431_0, i_10_207_1432_0, i_10_207_1443_0, i_10_207_1444_0,
    i_10_207_1539_0, i_10_207_1576_0, i_10_207_1683_0, i_10_207_1686_0,
    i_10_207_1728_0, i_10_207_1818_0, i_10_207_1819_0, i_10_207_2021_0,
    i_10_207_2223_0, i_10_207_2352_0, i_10_207_2359_0, i_10_207_2361_0,
    i_10_207_2364_0, i_10_207_2431_0, i_10_207_2442_0, i_10_207_2449_0,
    i_10_207_2450_0, i_10_207_2451_0, i_10_207_2454_0, i_10_207_2628_0,
    i_10_207_2629_0, i_10_207_2655_0, i_10_207_2658_0, i_10_207_2659_0,
    i_10_207_2661_0, i_10_207_2681_0, i_10_207_2701_0, i_10_207_2714_0,
    i_10_207_2727_0, i_10_207_2784_0, i_10_207_2862_0, i_10_207_2916_0,
    i_10_207_3038_0, i_10_207_3074_0, i_10_207_3267_0, i_10_207_3271_0,
    i_10_207_3277_0, i_10_207_3279_0, i_10_207_3280_0, i_10_207_3282_0,
    i_10_207_3316_0, i_10_207_3331_0, i_10_207_3349_0, i_10_207_3450_0,
    i_10_207_3497_0, i_10_207_3537_0, i_10_207_3538_0, i_10_207_3614_0,
    i_10_207_3617_0, i_10_207_3650_0, i_10_207_3786_0, i_10_207_3787_0,
    i_10_207_3834_0, i_10_207_3846_0, i_10_207_3854_0, i_10_207_4116_0,
    i_10_207_4119_0, i_10_207_4171_0, i_10_207_4172_0, i_10_207_4204_0,
    i_10_207_4219_0, i_10_207_4267_0, i_10_207_4269_0, i_10_207_4270_0,
    i_10_207_4279_0, i_10_207_4284_0, i_10_207_4285_0, i_10_207_4288_0,
    i_10_207_4428_0, i_10_207_4459_0, i_10_207_4582_0, i_10_207_4591_0;
  output o_10_207_0_0;
  assign o_10_207_0_0 = 0;
endmodule



// Benchmark "kernel_10_208" written by ABC on Sun Jul 19 10:24:36 2020

module kernel_10_208 ( 
    i_10_208_28_0, i_10_208_89_0, i_10_208_224_0, i_10_208_247_0,
    i_10_208_283_0, i_10_208_315_0, i_10_208_324_0, i_10_208_325_0,
    i_10_208_408_0, i_10_208_446_0, i_10_208_447_0, i_10_208_463_0,
    i_10_208_464_0, i_10_208_467_0, i_10_208_508_0, i_10_208_510_0,
    i_10_208_737_0, i_10_208_755_0, i_10_208_798_0, i_10_208_800_0,
    i_10_208_966_0, i_10_208_1027_0, i_10_208_1030_0, i_10_208_1034_0,
    i_10_208_1039_0, i_10_208_1140_0, i_10_208_1233_0, i_10_208_1234_0,
    i_10_208_1235_0, i_10_208_1238_0, i_10_208_1241_0, i_10_208_1307_0,
    i_10_208_1313_0, i_10_208_1363_0, i_10_208_1579_0, i_10_208_1650_0,
    i_10_208_1652_0, i_10_208_1820_0, i_10_208_1825_0, i_10_208_1910_0,
    i_10_208_1995_0, i_10_208_1996_0, i_10_208_2179_0, i_10_208_2186_0,
    i_10_208_2338_0, i_10_208_2382_0, i_10_208_2383_0, i_10_208_2384_0,
    i_10_208_2463_0, i_10_208_2464_0, i_10_208_2470_0, i_10_208_2474_0,
    i_10_208_2629_0, i_10_208_2661_0, i_10_208_2680_0, i_10_208_2706_0,
    i_10_208_2707_0, i_10_208_2714_0, i_10_208_2721_0, i_10_208_2730_0,
    i_10_208_2832_0, i_10_208_2833_0, i_10_208_2985_0, i_10_208_3039_0,
    i_10_208_3040_0, i_10_208_3049_0, i_10_208_3162_0, i_10_208_3165_0,
    i_10_208_3196_0, i_10_208_3197_0, i_10_208_3268_0, i_10_208_3270_0,
    i_10_208_3271_0, i_10_208_3321_0, i_10_208_3388_0, i_10_208_3389_0,
    i_10_208_3391_0, i_10_208_3402_0, i_10_208_3406_0, i_10_208_3468_0,
    i_10_208_3582_0, i_10_208_3609_0, i_10_208_3615_0, i_10_208_3785_0,
    i_10_208_3787_0, i_10_208_3834_0, i_10_208_3837_0, i_10_208_3846_0,
    i_10_208_3847_0, i_10_208_3889_0, i_10_208_3984_0, i_10_208_3985_0,
    i_10_208_4030_0, i_10_208_4031_0, i_10_208_4116_0, i_10_208_4128_0,
    i_10_208_4155_0, i_10_208_4217_0, i_10_208_4292_0, i_10_208_4567_0,
    o_10_208_0_0  );
  input  i_10_208_28_0, i_10_208_89_0, i_10_208_224_0, i_10_208_247_0,
    i_10_208_283_0, i_10_208_315_0, i_10_208_324_0, i_10_208_325_0,
    i_10_208_408_0, i_10_208_446_0, i_10_208_447_0, i_10_208_463_0,
    i_10_208_464_0, i_10_208_467_0, i_10_208_508_0, i_10_208_510_0,
    i_10_208_737_0, i_10_208_755_0, i_10_208_798_0, i_10_208_800_0,
    i_10_208_966_0, i_10_208_1027_0, i_10_208_1030_0, i_10_208_1034_0,
    i_10_208_1039_0, i_10_208_1140_0, i_10_208_1233_0, i_10_208_1234_0,
    i_10_208_1235_0, i_10_208_1238_0, i_10_208_1241_0, i_10_208_1307_0,
    i_10_208_1313_0, i_10_208_1363_0, i_10_208_1579_0, i_10_208_1650_0,
    i_10_208_1652_0, i_10_208_1820_0, i_10_208_1825_0, i_10_208_1910_0,
    i_10_208_1995_0, i_10_208_1996_0, i_10_208_2179_0, i_10_208_2186_0,
    i_10_208_2338_0, i_10_208_2382_0, i_10_208_2383_0, i_10_208_2384_0,
    i_10_208_2463_0, i_10_208_2464_0, i_10_208_2470_0, i_10_208_2474_0,
    i_10_208_2629_0, i_10_208_2661_0, i_10_208_2680_0, i_10_208_2706_0,
    i_10_208_2707_0, i_10_208_2714_0, i_10_208_2721_0, i_10_208_2730_0,
    i_10_208_2832_0, i_10_208_2833_0, i_10_208_2985_0, i_10_208_3039_0,
    i_10_208_3040_0, i_10_208_3049_0, i_10_208_3162_0, i_10_208_3165_0,
    i_10_208_3196_0, i_10_208_3197_0, i_10_208_3268_0, i_10_208_3270_0,
    i_10_208_3271_0, i_10_208_3321_0, i_10_208_3388_0, i_10_208_3389_0,
    i_10_208_3391_0, i_10_208_3402_0, i_10_208_3406_0, i_10_208_3468_0,
    i_10_208_3582_0, i_10_208_3609_0, i_10_208_3615_0, i_10_208_3785_0,
    i_10_208_3787_0, i_10_208_3834_0, i_10_208_3837_0, i_10_208_3846_0,
    i_10_208_3847_0, i_10_208_3889_0, i_10_208_3984_0, i_10_208_3985_0,
    i_10_208_4030_0, i_10_208_4031_0, i_10_208_4116_0, i_10_208_4128_0,
    i_10_208_4155_0, i_10_208_4217_0, i_10_208_4292_0, i_10_208_4567_0;
  output o_10_208_0_0;
  assign o_10_208_0_0 = ~((~i_10_208_3785_0 & ((i_10_208_463_0 & ((~i_10_208_283_0 & ~i_10_208_1027_0 & ~i_10_208_2384_0 & i_10_208_2629_0 & ~i_10_208_2833_0 & ~i_10_208_3197_0 & ~i_10_208_3270_0 & ~i_10_208_3271_0 & ~i_10_208_4030_0) | (~i_10_208_89_0 & ~i_10_208_798_0 & ~i_10_208_1307_0 & ~i_10_208_2179_0 & ~i_10_208_3268_0 & ~i_10_208_3834_0 & ~i_10_208_4128_0 & ~i_10_208_4292_0 & ~i_10_208_4567_0))) | (~i_10_208_1996_0 & ((~i_10_208_1363_0 & ~i_10_208_1825_0 & ~i_10_208_2382_0 & i_10_208_2721_0 & i_10_208_3388_0) | (~i_10_208_28_0 & ~i_10_208_2680_0 & ~i_10_208_3039_0 & ~i_10_208_3196_0 & ~i_10_208_3270_0 & ~i_10_208_3406_0 & i_10_208_3834_0 & ~i_10_208_3984_0))) | (~i_10_208_3837_0 & ((~i_10_208_2383_0 & ~i_10_208_2707_0 & ~i_10_208_3270_0 & i_10_208_3846_0) | (~i_10_208_1233_0 & ~i_10_208_2382_0 & i_10_208_2629_0 & ~i_10_208_2706_0 & ~i_10_208_3268_0 & ~i_10_208_3846_0))) | (~i_10_208_447_0 & ~i_10_208_463_0 & ~i_10_208_1652_0 & ~i_10_208_3196_0 & ~i_10_208_3406_0 & i_10_208_3847_0))) | (~i_10_208_3609_0 & ((~i_10_208_28_0 & ((i_10_208_467_0 & ~i_10_208_2707_0 & ~i_10_208_3271_0) | (~i_10_208_446_0 & ~i_10_208_463_0 & ~i_10_208_2383_0 & ~i_10_208_2730_0 & ~i_10_208_3197_0 & ~i_10_208_3837_0 & ~i_10_208_4128_0 & ~i_10_208_4292_0))) | (~i_10_208_447_0 & ~i_10_208_1027_0 & ~i_10_208_1233_0 & ~i_10_208_2179_0 & ~i_10_208_2384_0 & ~i_10_208_2832_0 & ~i_10_208_3406_0 & ~i_10_208_3984_0))) | (~i_10_208_89_0 & ((~i_10_208_1034_0 & ~i_10_208_1235_0 & ~i_10_208_1238_0 & ~i_10_208_2338_0 & ~i_10_208_2384_0 & i_10_208_2730_0 & ~i_10_208_3049_0 & ~i_10_208_3165_0 & ~i_10_208_3270_0 & ~i_10_208_3406_0 & ~i_10_208_3468_0 & ~i_10_208_3615_0) | (i_10_208_1234_0 & i_10_208_1235_0 & i_10_208_1238_0 & ~i_10_208_1995_0 & ~i_10_208_3402_0 & ~i_10_208_4030_0))) | (~i_10_208_3271_0 & ((~i_10_208_463_0 & ((~i_10_208_1652_0 & ~i_10_208_2382_0 & ~i_10_208_3162_0 & ~i_10_208_3582_0 & ~i_10_208_3615_0 & ~i_10_208_3834_0 & ~i_10_208_3837_0) | (~i_10_208_247_0 & ~i_10_208_798_0 & ~i_10_208_1027_0 & ~i_10_208_1307_0 & ~i_10_208_2338_0 & ~i_10_208_3270_0 & ~i_10_208_3846_0 & ~i_10_208_4128_0 & ~i_10_208_4292_0))) | (~i_10_208_2382_0 & ((~i_10_208_1820_0 & ~i_10_208_2179_0 & ~i_10_208_2706_0 & ~i_10_208_2707_0 & ~i_10_208_3196_0 & ~i_10_208_3268_0 & ~i_10_208_3402_0) | (i_10_208_464_0 & ~i_10_208_1650_0 & ~i_10_208_3406_0))))) | (~i_10_208_2179_0 & ((~i_10_208_2985_0 & ((~i_10_208_800_0 & ~i_10_208_2832_0 & ~i_10_208_3889_0 & ((~i_10_208_1027_0 & ~i_10_208_1034_0 & ~i_10_208_1820_0 & i_10_208_2384_0 & ~i_10_208_3582_0) | (~i_10_208_447_0 & ~i_10_208_1650_0 & ~i_10_208_1995_0 & ~i_10_208_3049_0 & ~i_10_208_3406_0 & ~i_10_208_3615_0 & ~i_10_208_3985_0))) | (~i_10_208_1027_0 & ~i_10_208_1030_0 & ~i_10_208_1820_0 & ~i_10_208_2707_0 & ~i_10_208_3049_0 & ~i_10_208_3270_0 & ~i_10_208_3406_0 & ~i_10_208_4567_0))) | (~i_10_208_1241_0 & ~i_10_208_1307_0 & ~i_10_208_2382_0 & ~i_10_208_3049_0 & ~i_10_208_3162_0 & i_10_208_3615_0 & i_10_208_4116_0) | (i_10_208_800_0 & ~i_10_208_1650_0 & i_10_208_3889_0 & i_10_208_4292_0))) | (~i_10_208_1027_0 & ((i_10_208_464_0 & ~i_10_208_1650_0 & ~i_10_208_2383_0 & i_10_208_2629_0) | (~i_10_208_1996_0 & ~i_10_208_2730_0 & i_10_208_3388_0 & ~i_10_208_3846_0 & ~i_10_208_4567_0))) | (i_10_208_1234_0 & ((~i_10_208_1579_0 & ~i_10_208_3270_0 & ~i_10_208_3406_0 & ~i_10_208_3787_0 & ~i_10_208_3834_0) | (~i_10_208_325_0 & ~i_10_208_2629_0 & ~i_10_208_2714_0 & ~i_10_208_2833_0 & ~i_10_208_3837_0 & ~i_10_208_3847_0))) | (~i_10_208_1650_0 & ((~i_10_208_1820_0 & i_10_208_1825_0 & ~i_10_208_2186_0 & ~i_10_208_2464_0 & ~i_10_208_3268_0 & ~i_10_208_3834_0 & ~i_10_208_3984_0) | (~i_10_208_2382_0 & ~i_10_208_2383_0 & ~i_10_208_3165_0 & ~i_10_208_3197_0 & ~i_10_208_3402_0 & ~i_10_208_4128_0 & ~i_10_208_4217_0))) | (~i_10_208_3268_0 & ((~i_10_208_2384_0 & ((~i_10_208_1034_0 & i_10_208_1820_0 & i_10_208_1825_0 & ~i_10_208_2706_0) | (i_10_208_1238_0 & ~i_10_208_2629_0 & ~i_10_208_3040_0 & ~i_10_208_3165_0))) | (i_10_208_283_0 & ~i_10_208_2707_0 & ~i_10_208_3270_0 & ~i_10_208_3582_0 & ~i_10_208_3847_0))) | (~i_10_208_2707_0 & i_10_208_3040_0 & i_10_208_3984_0) | (~i_10_208_224_0 & ~i_10_208_2382_0 & i_10_208_2714_0 & ~i_10_208_2730_0 & ~i_10_208_2832_0 & ~i_10_208_4567_0));
endmodule



// Benchmark "kernel_10_209" written by ABC on Sun Jul 19 10:24:37 2020

module kernel_10_209 ( 
    i_10_209_197_0, i_10_209_202_0, i_10_209_273_0, i_10_209_274_0,
    i_10_209_276_0, i_10_209_277_0, i_10_209_279_0, i_10_209_293_0,
    i_10_209_392_0, i_10_209_408_0, i_10_209_447_0, i_10_209_509_0,
    i_10_209_515_0, i_10_209_792_0, i_10_209_959_0, i_10_209_985_0,
    i_10_209_1256_0, i_10_209_1322_0, i_10_209_1363_0, i_10_209_1394_0,
    i_10_209_1444_0, i_10_209_1462_0, i_10_209_1463_0, i_10_209_1484_0,
    i_10_209_1526_0, i_10_209_1552_0, i_10_209_1570_0, i_10_209_1573_0,
    i_10_209_1610_0, i_10_209_1643_0, i_10_209_1713_0, i_10_209_1716_0,
    i_10_209_1744_0, i_10_209_1764_0, i_10_209_1772_0, i_10_209_1820_0,
    i_10_209_1915_0, i_10_209_2005_0, i_10_209_2011_0, i_10_209_2019_0,
    i_10_209_2020_0, i_10_209_2022_0, i_10_209_2028_0, i_10_209_2182_0,
    i_10_209_2185_0, i_10_209_2186_0, i_10_209_2303_0, i_10_209_2327_0,
    i_10_209_2329_0, i_10_209_2330_0, i_10_209_2359_0, i_10_209_2434_0,
    i_10_209_2482_0, i_10_209_2483_0, i_10_209_2505_0, i_10_209_2506_0,
    i_10_209_2510_0, i_10_209_2634_0, i_10_209_2642_0, i_10_209_2675_0,
    i_10_209_2824_0, i_10_209_2874_0, i_10_209_2884_0, i_10_209_2965_0,
    i_10_209_2986_0, i_10_209_2987_0, i_10_209_3032_0, i_10_209_3039_0,
    i_10_209_3076_0, i_10_209_3320_0, i_10_209_3362_0, i_10_209_3364_0,
    i_10_209_3365_0, i_10_209_3431_0, i_10_209_3437_0, i_10_209_3496_0,
    i_10_209_3521_0, i_10_209_3717_0, i_10_209_3720_0, i_10_209_3806_0,
    i_10_209_3838_0, i_10_209_3841_0, i_10_209_3889_0, i_10_209_3890_0,
    i_10_209_3896_0, i_10_209_3920_0, i_10_209_3965_0, i_10_209_3982_0,
    i_10_209_3989_0, i_10_209_3992_0, i_10_209_4143_0, i_10_209_4144_0,
    i_10_209_4283_0, i_10_209_4360_0, i_10_209_4445_0, i_10_209_4526_0,
    i_10_209_4568_0, i_10_209_4574_0, i_10_209_4577_0, i_10_209_4596_0,
    o_10_209_0_0  );
  input  i_10_209_197_0, i_10_209_202_0, i_10_209_273_0, i_10_209_274_0,
    i_10_209_276_0, i_10_209_277_0, i_10_209_279_0, i_10_209_293_0,
    i_10_209_392_0, i_10_209_408_0, i_10_209_447_0, i_10_209_509_0,
    i_10_209_515_0, i_10_209_792_0, i_10_209_959_0, i_10_209_985_0,
    i_10_209_1256_0, i_10_209_1322_0, i_10_209_1363_0, i_10_209_1394_0,
    i_10_209_1444_0, i_10_209_1462_0, i_10_209_1463_0, i_10_209_1484_0,
    i_10_209_1526_0, i_10_209_1552_0, i_10_209_1570_0, i_10_209_1573_0,
    i_10_209_1610_0, i_10_209_1643_0, i_10_209_1713_0, i_10_209_1716_0,
    i_10_209_1744_0, i_10_209_1764_0, i_10_209_1772_0, i_10_209_1820_0,
    i_10_209_1915_0, i_10_209_2005_0, i_10_209_2011_0, i_10_209_2019_0,
    i_10_209_2020_0, i_10_209_2022_0, i_10_209_2028_0, i_10_209_2182_0,
    i_10_209_2185_0, i_10_209_2186_0, i_10_209_2303_0, i_10_209_2327_0,
    i_10_209_2329_0, i_10_209_2330_0, i_10_209_2359_0, i_10_209_2434_0,
    i_10_209_2482_0, i_10_209_2483_0, i_10_209_2505_0, i_10_209_2506_0,
    i_10_209_2510_0, i_10_209_2634_0, i_10_209_2642_0, i_10_209_2675_0,
    i_10_209_2824_0, i_10_209_2874_0, i_10_209_2884_0, i_10_209_2965_0,
    i_10_209_2986_0, i_10_209_2987_0, i_10_209_3032_0, i_10_209_3039_0,
    i_10_209_3076_0, i_10_209_3320_0, i_10_209_3362_0, i_10_209_3364_0,
    i_10_209_3365_0, i_10_209_3431_0, i_10_209_3437_0, i_10_209_3496_0,
    i_10_209_3521_0, i_10_209_3717_0, i_10_209_3720_0, i_10_209_3806_0,
    i_10_209_3838_0, i_10_209_3841_0, i_10_209_3889_0, i_10_209_3890_0,
    i_10_209_3896_0, i_10_209_3920_0, i_10_209_3965_0, i_10_209_3982_0,
    i_10_209_3989_0, i_10_209_3992_0, i_10_209_4143_0, i_10_209_4144_0,
    i_10_209_4283_0, i_10_209_4360_0, i_10_209_4445_0, i_10_209_4526_0,
    i_10_209_4568_0, i_10_209_4574_0, i_10_209_4577_0, i_10_209_4596_0;
  output o_10_209_0_0;
  assign o_10_209_0_0 = 0;
endmodule



// Benchmark "kernel_10_210" written by ABC on Sun Jul 19 10:24:38 2020

module kernel_10_210 ( 
    i_10_210_175_0, i_10_210_283_0, i_10_210_284_0, i_10_210_285_0,
    i_10_210_286_0, i_10_210_289_0, i_10_210_318_0, i_10_210_325_0,
    i_10_210_390_0, i_10_210_425_0, i_10_210_460_0, i_10_210_463_0,
    i_10_210_464_0, i_10_210_514_0, i_10_210_639_0, i_10_210_752_0,
    i_10_210_892_0, i_10_210_893_0, i_10_210_965_0, i_10_210_967_0,
    i_10_210_990_0, i_10_210_1003_0, i_10_210_1026_0, i_10_210_1235_0,
    i_10_210_1241_0, i_10_210_1296_0, i_10_210_1305_0, i_10_210_1306_0,
    i_10_210_1307_0, i_10_210_1342_0, i_10_210_1542_0, i_10_210_1603_0,
    i_10_210_1629_0, i_10_210_1651_0, i_10_210_1652_0, i_10_210_1653_0,
    i_10_210_1655_0, i_10_210_1720_0, i_10_210_1721_0, i_10_210_1821_0,
    i_10_210_1822_0, i_10_210_1823_0, i_10_210_1909_0, i_10_210_1910_0,
    i_10_210_1916_0, i_10_210_1989_0, i_10_210_1990_0, i_10_210_2026_0,
    i_10_210_2288_0, i_10_210_2359_0, i_10_210_2361_0, i_10_210_2362_0,
    i_10_210_2377_0, i_10_210_2378_0, i_10_210_2566_0, i_10_210_2631_0,
    i_10_210_2656_0, i_10_210_2657_0, i_10_210_2675_0, i_10_210_2702_0,
    i_10_210_2710_0, i_10_210_2725_0, i_10_210_2726_0, i_10_210_2828_0,
    i_10_210_2918_0, i_10_210_2919_0, i_10_210_2980_0, i_10_210_3035_0,
    i_10_210_3069_0, i_10_210_3269_0, i_10_210_3384_0, i_10_210_3389_0,
    i_10_210_3403_0, i_10_210_3405_0, i_10_210_3555_0, i_10_210_3556_0,
    i_10_210_3582_0, i_10_210_3613_0, i_10_210_3615_0, i_10_210_3616_0,
    i_10_210_3617_0, i_10_210_3647_0, i_10_210_3683_0, i_10_210_3846_0,
    i_10_210_3848_0, i_10_210_3856_0, i_10_210_3888_0, i_10_210_3889_0,
    i_10_210_3980_0, i_10_210_4023_0, i_10_210_4096_0, i_10_210_4123_0,
    i_10_210_4125_0, i_10_210_4127_0, i_10_210_4214_0, i_10_210_4287_0,
    i_10_210_4288_0, i_10_210_4565_0, i_10_210_4567_0, i_10_210_4568_0,
    o_10_210_0_0  );
  input  i_10_210_175_0, i_10_210_283_0, i_10_210_284_0, i_10_210_285_0,
    i_10_210_286_0, i_10_210_289_0, i_10_210_318_0, i_10_210_325_0,
    i_10_210_390_0, i_10_210_425_0, i_10_210_460_0, i_10_210_463_0,
    i_10_210_464_0, i_10_210_514_0, i_10_210_639_0, i_10_210_752_0,
    i_10_210_892_0, i_10_210_893_0, i_10_210_965_0, i_10_210_967_0,
    i_10_210_990_0, i_10_210_1003_0, i_10_210_1026_0, i_10_210_1235_0,
    i_10_210_1241_0, i_10_210_1296_0, i_10_210_1305_0, i_10_210_1306_0,
    i_10_210_1307_0, i_10_210_1342_0, i_10_210_1542_0, i_10_210_1603_0,
    i_10_210_1629_0, i_10_210_1651_0, i_10_210_1652_0, i_10_210_1653_0,
    i_10_210_1655_0, i_10_210_1720_0, i_10_210_1721_0, i_10_210_1821_0,
    i_10_210_1822_0, i_10_210_1823_0, i_10_210_1909_0, i_10_210_1910_0,
    i_10_210_1916_0, i_10_210_1989_0, i_10_210_1990_0, i_10_210_2026_0,
    i_10_210_2288_0, i_10_210_2359_0, i_10_210_2361_0, i_10_210_2362_0,
    i_10_210_2377_0, i_10_210_2378_0, i_10_210_2566_0, i_10_210_2631_0,
    i_10_210_2656_0, i_10_210_2657_0, i_10_210_2675_0, i_10_210_2702_0,
    i_10_210_2710_0, i_10_210_2725_0, i_10_210_2726_0, i_10_210_2828_0,
    i_10_210_2918_0, i_10_210_2919_0, i_10_210_2980_0, i_10_210_3035_0,
    i_10_210_3069_0, i_10_210_3269_0, i_10_210_3384_0, i_10_210_3389_0,
    i_10_210_3403_0, i_10_210_3405_0, i_10_210_3555_0, i_10_210_3556_0,
    i_10_210_3582_0, i_10_210_3613_0, i_10_210_3615_0, i_10_210_3616_0,
    i_10_210_3617_0, i_10_210_3647_0, i_10_210_3683_0, i_10_210_3846_0,
    i_10_210_3848_0, i_10_210_3856_0, i_10_210_3888_0, i_10_210_3889_0,
    i_10_210_3980_0, i_10_210_4023_0, i_10_210_4096_0, i_10_210_4123_0,
    i_10_210_4125_0, i_10_210_4127_0, i_10_210_4214_0, i_10_210_4287_0,
    i_10_210_4288_0, i_10_210_4565_0, i_10_210_4567_0, i_10_210_4568_0;
  output o_10_210_0_0;
  assign o_10_210_0_0 = ~((~i_10_210_175_0 & ((~i_10_210_425_0 & ~i_10_210_514_0 & ~i_10_210_892_0 & ~i_10_210_990_0 & ~i_10_210_1823_0 & ~i_10_210_3846_0) | (~i_10_210_325_0 & ~i_10_210_965_0 & i_10_210_1651_0 & ~i_10_210_3683_0 & i_10_210_3848_0 & ~i_10_210_3980_0))) | (~i_10_210_390_0 & ((i_10_210_1821_0 & ~i_10_210_2362_0 & i_10_210_2631_0 & ~i_10_210_2725_0 & ~i_10_210_2980_0 & ~i_10_210_4565_0 & i_10_210_4568_0) | (~i_10_210_2359_0 & ~i_10_210_2377_0 & ~i_10_210_2675_0 & ~i_10_210_2710_0 & ~i_10_210_3035_0 & ~i_10_210_4125_0 & ~i_10_210_4568_0))) | (i_10_210_460_0 & ((~i_10_210_286_0 & ~i_10_210_639_0 & ~i_10_210_1026_0 & ~i_10_210_1342_0 & ~i_10_210_1990_0 & ~i_10_210_2361_0) | (i_10_210_1909_0 & ~i_10_210_4567_0))) | (~i_10_210_460_0 & ((~i_10_210_1542_0 & i_10_210_1655_0 & ~i_10_210_1990_0 & ~i_10_210_3069_0 & ~i_10_210_3582_0 & ~i_10_210_3856_0) | (~i_10_210_892_0 & i_10_210_2919_0 & i_10_210_3889_0 & i_10_210_3980_0 & ~i_10_210_4287_0))) | (i_10_210_463_0 & ((~i_10_210_284_0 & ~i_10_210_639_0 & i_10_210_2631_0 & ~i_10_210_3403_0) | (i_10_210_464_0 & i_10_210_1241_0 & ~i_10_210_4214_0))) | (i_10_210_1909_0 & (i_10_210_464_0 | (i_10_210_325_0 & ~i_10_210_1989_0 & ~i_10_210_3683_0))) | (~i_10_210_2359_0 & ((i_10_210_1655_0 & ~i_10_210_1822_0) | (~i_10_210_2361_0 & ~i_10_210_2631_0 & ~i_10_210_2828_0 & ~i_10_210_3846_0 & ~i_10_210_4123_0 & ~i_10_210_4127_0))) | (~i_10_210_2566_0 & ((i_10_210_3035_0 & i_10_210_3647_0) | (~i_10_210_893_0 & ~i_10_210_1342_0 & ~i_10_210_1989_0 & ~i_10_210_3683_0 & ~i_10_210_3848_0 & ~i_10_210_4287_0))) | (~i_10_210_2919_0 & ((i_10_210_1653_0 & ~i_10_210_1821_0 & ~i_10_210_1989_0) | (~i_10_210_2377_0 & ~i_10_210_2702_0 & i_10_210_3389_0 & ~i_10_210_4565_0 & ~i_10_210_4567_0))) | (~i_10_210_4565_0 & ((~i_10_210_3269_0 & ((~i_10_210_1235_0 & i_10_210_1652_0) | (~i_10_210_639_0 & ~i_10_210_1241_0 & ~i_10_210_2377_0 & ~i_10_210_2378_0 & ~i_10_210_2675_0 & ~i_10_210_2918_0 & ~i_10_210_3582_0 & ~i_10_210_3846_0 & ~i_10_210_4123_0))) | (~i_10_210_284_0 & ~i_10_210_2725_0 & i_10_210_3846_0 & ~i_10_210_4287_0 & i_10_210_4568_0))) | (~i_10_210_2377_0 & ((~i_10_210_284_0 & ((~i_10_210_3846_0 & ~i_10_210_4123_0 & i_10_210_1651_0 & ~i_10_210_1989_0) | (i_10_210_2725_0 & i_10_210_2726_0 & ~i_10_210_3384_0 & i_10_210_3389_0 & ~i_10_210_4214_0))) | (i_10_210_1026_0 & i_10_210_1305_0 & ~i_10_210_3848_0))) | (~i_10_210_1989_0 & ((~i_10_210_1026_0 & i_10_210_1306_0) | (~i_10_210_1651_0 & ~i_10_210_3683_0 & ~i_10_210_3848_0 & ~i_10_210_4288_0))) | (~i_10_210_892_0 & ~i_10_210_3069_0 & ~i_10_210_3384_0 & ~i_10_210_3848_0 & ~i_10_210_4125_0 & ~i_10_210_4127_0) | (i_10_210_285_0 & ~i_10_210_2710_0 & i_10_210_4568_0) | (i_10_210_1910_0 & ~i_10_210_4567_0 & ~i_10_210_4568_0));
endmodule



// Benchmark "kernel_10_211" written by ABC on Sun Jul 19 10:24:39 2020

module kernel_10_211 ( 
    i_10_211_9_0, i_10_211_153_0, i_10_211_174_0, i_10_211_175_0,
    i_10_211_223_0, i_10_211_280_0, i_10_211_284_0, i_10_211_315_0,
    i_10_211_316_0, i_10_211_327_0, i_10_211_390_0, i_10_211_437_0,
    i_10_211_445_0, i_10_211_448_0, i_10_211_459_0, i_10_211_460_0,
    i_10_211_621_0, i_10_211_687_0, i_10_211_688_0, i_10_211_820_0,
    i_10_211_903_0, i_10_211_990_0, i_10_211_1030_0, i_10_211_1080_0,
    i_10_211_1083_0, i_10_211_1107_0, i_10_211_1215_0, i_10_211_1218_0,
    i_10_211_1236_0, i_10_211_1237_0, i_10_211_1239_0, i_10_211_1241_0,
    i_10_211_1264_0, i_10_211_1582_0, i_10_211_1800_0, i_10_211_1818_0,
    i_10_211_1826_0, i_10_211_1945_0, i_10_211_2016_0, i_10_211_2017_0,
    i_10_211_2026_0, i_10_211_2181_0, i_10_211_2199_0, i_10_211_2336_0,
    i_10_211_2352_0, i_10_211_2353_0, i_10_211_2355_0, i_10_211_2377_0,
    i_10_211_2378_0, i_10_211_2379_0, i_10_211_2406_0, i_10_211_2460_0,
    i_10_211_2466_0, i_10_211_2468_0, i_10_211_2471_0, i_10_211_2511_0,
    i_10_211_2514_0, i_10_211_2605_0, i_10_211_2611_0, i_10_211_2657_0,
    i_10_211_2700_0, i_10_211_2709_0, i_10_211_2718_0, i_10_211_2734_0,
    i_10_211_2783_0, i_10_211_2831_0, i_10_211_2881_0, i_10_211_3042_0,
    i_10_211_3069_0, i_10_211_3094_0, i_10_211_3392_0, i_10_211_3409_0,
    i_10_211_3468_0, i_10_211_3493_0, i_10_211_3610_0, i_10_211_3614_0,
    i_10_211_3616_0, i_10_211_3717_0, i_10_211_3720_0, i_10_211_3846_0,
    i_10_211_3855_0, i_10_211_3857_0, i_10_211_3894_0, i_10_211_3905_0,
    i_10_211_3906_0, i_10_211_3907_0, i_10_211_3909_0, i_10_211_4030_0,
    i_10_211_4122_0, i_10_211_4123_0, i_10_211_4168_0, i_10_211_4170_0,
    i_10_211_4176_0, i_10_211_4276_0, i_10_211_4291_0, i_10_211_4410_0,
    i_10_211_4566_0, i_10_211_4567_0, i_10_211_4568_0, i_10_211_4581_0,
    o_10_211_0_0  );
  input  i_10_211_9_0, i_10_211_153_0, i_10_211_174_0, i_10_211_175_0,
    i_10_211_223_0, i_10_211_280_0, i_10_211_284_0, i_10_211_315_0,
    i_10_211_316_0, i_10_211_327_0, i_10_211_390_0, i_10_211_437_0,
    i_10_211_445_0, i_10_211_448_0, i_10_211_459_0, i_10_211_460_0,
    i_10_211_621_0, i_10_211_687_0, i_10_211_688_0, i_10_211_820_0,
    i_10_211_903_0, i_10_211_990_0, i_10_211_1030_0, i_10_211_1080_0,
    i_10_211_1083_0, i_10_211_1107_0, i_10_211_1215_0, i_10_211_1218_0,
    i_10_211_1236_0, i_10_211_1237_0, i_10_211_1239_0, i_10_211_1241_0,
    i_10_211_1264_0, i_10_211_1582_0, i_10_211_1800_0, i_10_211_1818_0,
    i_10_211_1826_0, i_10_211_1945_0, i_10_211_2016_0, i_10_211_2017_0,
    i_10_211_2026_0, i_10_211_2181_0, i_10_211_2199_0, i_10_211_2336_0,
    i_10_211_2352_0, i_10_211_2353_0, i_10_211_2355_0, i_10_211_2377_0,
    i_10_211_2378_0, i_10_211_2379_0, i_10_211_2406_0, i_10_211_2460_0,
    i_10_211_2466_0, i_10_211_2468_0, i_10_211_2471_0, i_10_211_2511_0,
    i_10_211_2514_0, i_10_211_2605_0, i_10_211_2611_0, i_10_211_2657_0,
    i_10_211_2700_0, i_10_211_2709_0, i_10_211_2718_0, i_10_211_2734_0,
    i_10_211_2783_0, i_10_211_2831_0, i_10_211_2881_0, i_10_211_3042_0,
    i_10_211_3069_0, i_10_211_3094_0, i_10_211_3392_0, i_10_211_3409_0,
    i_10_211_3468_0, i_10_211_3493_0, i_10_211_3610_0, i_10_211_3614_0,
    i_10_211_3616_0, i_10_211_3717_0, i_10_211_3720_0, i_10_211_3846_0,
    i_10_211_3855_0, i_10_211_3857_0, i_10_211_3894_0, i_10_211_3905_0,
    i_10_211_3906_0, i_10_211_3907_0, i_10_211_3909_0, i_10_211_4030_0,
    i_10_211_4122_0, i_10_211_4123_0, i_10_211_4168_0, i_10_211_4170_0,
    i_10_211_4176_0, i_10_211_4276_0, i_10_211_4291_0, i_10_211_4410_0,
    i_10_211_4566_0, i_10_211_4567_0, i_10_211_4568_0, i_10_211_4581_0;
  output o_10_211_0_0;
  assign o_10_211_0_0 = 0;
endmodule



// Benchmark "kernel_10_212" written by ABC on Sun Jul 19 10:24:40 2020

module kernel_10_212 ( 
    i_10_212_28_0, i_10_212_175_0, i_10_212_178_0, i_10_212_286_0,
    i_10_212_327_0, i_10_212_444_0, i_10_212_461_0, i_10_212_463_0,
    i_10_212_464_0, i_10_212_514_0, i_10_212_794_0, i_10_212_797_0,
    i_10_212_901_0, i_10_212_956_0, i_10_212_958_0, i_10_212_959_0,
    i_10_212_999_0, i_10_212_1000_0, i_10_212_1009_0, i_10_212_1162_0,
    i_10_212_1241_0, i_10_212_1306_0, i_10_212_1378_0, i_10_212_1379_0,
    i_10_212_1486_0, i_10_212_1576_0, i_10_212_1654_0, i_10_212_1655_0,
    i_10_212_1685_0, i_10_212_1687_0, i_10_212_1688_0, i_10_212_1813_0,
    i_10_212_1821_0, i_10_212_1944_0, i_10_212_1945_0, i_10_212_1946_0,
    i_10_212_2090_0, i_10_212_2183_0, i_10_212_2203_0, i_10_212_2305_0,
    i_10_212_2378_0, i_10_212_2448_0, i_10_212_2449_0, i_10_212_2450_0,
    i_10_212_2455_0, i_10_212_2456_0, i_10_212_2470_0, i_10_212_2471_0,
    i_10_212_2635_0, i_10_212_2636_0, i_10_212_2638_0, i_10_212_2639_0,
    i_10_212_2674_0, i_10_212_2711_0, i_10_212_2717_0, i_10_212_2720_0,
    i_10_212_2727_0, i_10_212_2728_0, i_10_212_3034_0, i_10_212_3035_0,
    i_10_212_3037_0, i_10_212_3042_0, i_10_212_3043_0, i_10_212_3046_0,
    i_10_212_3074_0, i_10_212_3087_0, i_10_212_3203_0, i_10_212_3267_0,
    i_10_212_3271_0, i_10_212_3278_0, i_10_212_3281_0, i_10_212_3384_0,
    i_10_212_3390_0, i_10_212_3392_0, i_10_212_3409_0, i_10_212_3431_0,
    i_10_212_3495_0, i_10_212_3539_0, i_10_212_3725_0, i_10_212_3781_0,
    i_10_212_3786_0, i_10_212_3837_0, i_10_212_3838_0, i_10_212_3857_0,
    i_10_212_3888_0, i_10_212_3890_0, i_10_212_3911_0, i_10_212_3979_0,
    i_10_212_3992_0, i_10_212_4055_0, i_10_212_4117_0, i_10_212_4118_0,
    i_10_212_4119_0, i_10_212_4121_0, i_10_212_4126_0, i_10_212_4280_0,
    i_10_212_4284_0, i_10_212_4370_0, i_10_212_4429_0, i_10_212_4583_0,
    o_10_212_0_0  );
  input  i_10_212_28_0, i_10_212_175_0, i_10_212_178_0, i_10_212_286_0,
    i_10_212_327_0, i_10_212_444_0, i_10_212_461_0, i_10_212_463_0,
    i_10_212_464_0, i_10_212_514_0, i_10_212_794_0, i_10_212_797_0,
    i_10_212_901_0, i_10_212_956_0, i_10_212_958_0, i_10_212_959_0,
    i_10_212_999_0, i_10_212_1000_0, i_10_212_1009_0, i_10_212_1162_0,
    i_10_212_1241_0, i_10_212_1306_0, i_10_212_1378_0, i_10_212_1379_0,
    i_10_212_1486_0, i_10_212_1576_0, i_10_212_1654_0, i_10_212_1655_0,
    i_10_212_1685_0, i_10_212_1687_0, i_10_212_1688_0, i_10_212_1813_0,
    i_10_212_1821_0, i_10_212_1944_0, i_10_212_1945_0, i_10_212_1946_0,
    i_10_212_2090_0, i_10_212_2183_0, i_10_212_2203_0, i_10_212_2305_0,
    i_10_212_2378_0, i_10_212_2448_0, i_10_212_2449_0, i_10_212_2450_0,
    i_10_212_2455_0, i_10_212_2456_0, i_10_212_2470_0, i_10_212_2471_0,
    i_10_212_2635_0, i_10_212_2636_0, i_10_212_2638_0, i_10_212_2639_0,
    i_10_212_2674_0, i_10_212_2711_0, i_10_212_2717_0, i_10_212_2720_0,
    i_10_212_2727_0, i_10_212_2728_0, i_10_212_3034_0, i_10_212_3035_0,
    i_10_212_3037_0, i_10_212_3042_0, i_10_212_3043_0, i_10_212_3046_0,
    i_10_212_3074_0, i_10_212_3087_0, i_10_212_3203_0, i_10_212_3267_0,
    i_10_212_3271_0, i_10_212_3278_0, i_10_212_3281_0, i_10_212_3384_0,
    i_10_212_3390_0, i_10_212_3392_0, i_10_212_3409_0, i_10_212_3431_0,
    i_10_212_3495_0, i_10_212_3539_0, i_10_212_3725_0, i_10_212_3781_0,
    i_10_212_3786_0, i_10_212_3837_0, i_10_212_3838_0, i_10_212_3857_0,
    i_10_212_3888_0, i_10_212_3890_0, i_10_212_3911_0, i_10_212_3979_0,
    i_10_212_3992_0, i_10_212_4055_0, i_10_212_4117_0, i_10_212_4118_0,
    i_10_212_4119_0, i_10_212_4121_0, i_10_212_4126_0, i_10_212_4280_0,
    i_10_212_4284_0, i_10_212_4370_0, i_10_212_4429_0, i_10_212_4583_0;
  output o_10_212_0_0;
  assign o_10_212_0_0 = 0;
endmodule



// Benchmark "kernel_10_213" written by ABC on Sun Jul 19 10:24:40 2020

module kernel_10_213 ( 
    i_10_213_64_0, i_10_213_176_0, i_10_213_177_0, i_10_213_178_0,
    i_10_213_183_0, i_10_213_214_0, i_10_213_262_0, i_10_213_284_0,
    i_10_213_316_0, i_10_213_521_0, i_10_213_757_0, i_10_213_758_0,
    i_10_213_794_0, i_10_213_798_0, i_10_213_799_0, i_10_213_907_0,
    i_10_213_994_0, i_10_213_1000_0, i_10_213_1012_0, i_10_213_1039_0,
    i_10_213_1058_0, i_10_213_1114_0, i_10_213_1300_0, i_10_213_1354_0,
    i_10_213_1355_0, i_10_213_1367_0, i_10_213_1434_0, i_10_213_1577_0,
    i_10_213_1579_0, i_10_213_1622_0, i_10_213_1625_0, i_10_213_1649_0,
    i_10_213_1651_0, i_10_213_1652_0, i_10_213_1684_0, i_10_213_1685_0,
    i_10_213_1689_0, i_10_213_1691_0, i_10_213_1730_0, i_10_213_1822_0,
    i_10_213_1919_0, i_10_213_1982_0, i_10_213_2027_0, i_10_213_2030_0,
    i_10_213_2153_0, i_10_213_2180_0, i_10_213_2201_0, i_10_213_2288_0,
    i_10_213_2360_0, i_10_213_2449_0, i_10_213_2506_0, i_10_213_2533_0,
    i_10_213_2566_0, i_10_213_2567_0, i_10_213_2570_0, i_10_213_2641_0,
    i_10_213_2663_0, i_10_213_2714_0, i_10_213_2719_0, i_10_213_2720_0,
    i_10_213_2728_0, i_10_213_2731_0, i_10_213_2826_0, i_10_213_2829_0,
    i_10_213_2849_0, i_10_213_2924_0, i_10_213_2963_0, i_10_213_3041_0,
    i_10_213_3044_0, i_10_213_3269_0, i_10_213_3280_0, i_10_213_3314_0,
    i_10_213_3316_0, i_10_213_3317_0, i_10_213_3387_0, i_10_213_3406_0,
    i_10_213_3461_0, i_10_213_3539_0, i_10_213_3560_0, i_10_213_3584_0,
    i_10_213_3689_0, i_10_213_3797_0, i_10_213_3834_0, i_10_213_3835_0,
    i_10_213_3839_0, i_10_213_3842_0, i_10_213_3849_0, i_10_213_3852_0,
    i_10_213_3894_0, i_10_213_3895_0, i_10_213_3982_0, i_10_213_4025_0,
    i_10_213_4028_0, i_10_213_4127_0, i_10_213_4172_0, i_10_213_4267_0,
    i_10_213_4283_0, i_10_213_4289_0, i_10_213_4583_0, i_10_213_4596_0,
    o_10_213_0_0  );
  input  i_10_213_64_0, i_10_213_176_0, i_10_213_177_0, i_10_213_178_0,
    i_10_213_183_0, i_10_213_214_0, i_10_213_262_0, i_10_213_284_0,
    i_10_213_316_0, i_10_213_521_0, i_10_213_757_0, i_10_213_758_0,
    i_10_213_794_0, i_10_213_798_0, i_10_213_799_0, i_10_213_907_0,
    i_10_213_994_0, i_10_213_1000_0, i_10_213_1012_0, i_10_213_1039_0,
    i_10_213_1058_0, i_10_213_1114_0, i_10_213_1300_0, i_10_213_1354_0,
    i_10_213_1355_0, i_10_213_1367_0, i_10_213_1434_0, i_10_213_1577_0,
    i_10_213_1579_0, i_10_213_1622_0, i_10_213_1625_0, i_10_213_1649_0,
    i_10_213_1651_0, i_10_213_1652_0, i_10_213_1684_0, i_10_213_1685_0,
    i_10_213_1689_0, i_10_213_1691_0, i_10_213_1730_0, i_10_213_1822_0,
    i_10_213_1919_0, i_10_213_1982_0, i_10_213_2027_0, i_10_213_2030_0,
    i_10_213_2153_0, i_10_213_2180_0, i_10_213_2201_0, i_10_213_2288_0,
    i_10_213_2360_0, i_10_213_2449_0, i_10_213_2506_0, i_10_213_2533_0,
    i_10_213_2566_0, i_10_213_2567_0, i_10_213_2570_0, i_10_213_2641_0,
    i_10_213_2663_0, i_10_213_2714_0, i_10_213_2719_0, i_10_213_2720_0,
    i_10_213_2728_0, i_10_213_2731_0, i_10_213_2826_0, i_10_213_2829_0,
    i_10_213_2849_0, i_10_213_2924_0, i_10_213_2963_0, i_10_213_3041_0,
    i_10_213_3044_0, i_10_213_3269_0, i_10_213_3280_0, i_10_213_3314_0,
    i_10_213_3316_0, i_10_213_3317_0, i_10_213_3387_0, i_10_213_3406_0,
    i_10_213_3461_0, i_10_213_3539_0, i_10_213_3560_0, i_10_213_3584_0,
    i_10_213_3689_0, i_10_213_3797_0, i_10_213_3834_0, i_10_213_3835_0,
    i_10_213_3839_0, i_10_213_3842_0, i_10_213_3849_0, i_10_213_3852_0,
    i_10_213_3894_0, i_10_213_3895_0, i_10_213_3982_0, i_10_213_4025_0,
    i_10_213_4028_0, i_10_213_4127_0, i_10_213_4172_0, i_10_213_4267_0,
    i_10_213_4283_0, i_10_213_4289_0, i_10_213_4583_0, i_10_213_4596_0;
  output o_10_213_0_0;
  assign o_10_213_0_0 = 0;
endmodule



// Benchmark "kernel_10_214" written by ABC on Sun Jul 19 10:24:41 2020

module kernel_10_214 ( 
    i_10_214_42_0, i_10_214_43_0, i_10_214_144_0, i_10_214_145_0,
    i_10_214_159_0, i_10_214_175_0, i_10_214_250_0, i_10_214_287_0,
    i_10_214_293_0, i_10_214_296_0, i_10_214_327_0, i_10_214_328_0,
    i_10_214_391_0, i_10_214_409_0, i_10_214_411_0, i_10_214_430_0,
    i_10_214_539_0, i_10_214_898_0, i_10_214_1084_0, i_10_214_1131_0,
    i_10_214_1132_0, i_10_214_1234_0, i_10_214_1237_0, i_10_214_1239_0,
    i_10_214_1241_0, i_10_214_1269_0, i_10_214_1270_0, i_10_214_1306_0,
    i_10_214_1307_0, i_10_214_1357_0, i_10_214_1362_0, i_10_214_1365_0,
    i_10_214_1444_0, i_10_214_1445_0, i_10_214_1447_0, i_10_214_1448_0,
    i_10_214_1651_0, i_10_214_1654_0, i_10_214_1680_0, i_10_214_1726_0,
    i_10_214_1816_0, i_10_214_1875_0, i_10_214_2019_0, i_10_214_2020_0,
    i_10_214_2022_0, i_10_214_2050_0, i_10_214_2253_0, i_10_214_2256_0,
    i_10_214_2257_0, i_10_214_2258_0, i_10_214_2259_0, i_10_214_2325_0,
    i_10_214_2354_0, i_10_214_2364_0, i_10_214_2454_0, i_10_214_2467_0,
    i_10_214_2514_0, i_10_214_2527_0, i_10_214_2546_0, i_10_214_2571_0,
    i_10_214_2660_0, i_10_214_2675_0, i_10_214_2787_0, i_10_214_2839_0,
    i_10_214_2913_0, i_10_214_2914_0, i_10_214_2979_0, i_10_214_3047_0,
    i_10_214_3237_0, i_10_214_3284_0, i_10_214_3291_0, i_10_214_3389_0,
    i_10_214_3399_0, i_10_214_3433_0, i_10_214_3495_0, i_10_214_3499_0,
    i_10_214_3583_0, i_10_214_3585_0, i_10_214_3586_0, i_10_214_3590_0,
    i_10_214_3687_0, i_10_214_3814_0, i_10_214_3837_0, i_10_214_3846_0,
    i_10_214_3855_0, i_10_214_3856_0, i_10_214_3873_0, i_10_214_3887_0,
    i_10_214_3945_0, i_10_214_3948_0, i_10_214_3973_0, i_10_214_4028_0,
    i_10_214_4055_0, i_10_214_4119_0, i_10_214_4123_0, i_10_214_4128_0,
    i_10_214_4220_0, i_10_214_4236_0, i_10_214_4267_0, i_10_214_4269_0,
    o_10_214_0_0  );
  input  i_10_214_42_0, i_10_214_43_0, i_10_214_144_0, i_10_214_145_0,
    i_10_214_159_0, i_10_214_175_0, i_10_214_250_0, i_10_214_287_0,
    i_10_214_293_0, i_10_214_296_0, i_10_214_327_0, i_10_214_328_0,
    i_10_214_391_0, i_10_214_409_0, i_10_214_411_0, i_10_214_430_0,
    i_10_214_539_0, i_10_214_898_0, i_10_214_1084_0, i_10_214_1131_0,
    i_10_214_1132_0, i_10_214_1234_0, i_10_214_1237_0, i_10_214_1239_0,
    i_10_214_1241_0, i_10_214_1269_0, i_10_214_1270_0, i_10_214_1306_0,
    i_10_214_1307_0, i_10_214_1357_0, i_10_214_1362_0, i_10_214_1365_0,
    i_10_214_1444_0, i_10_214_1445_0, i_10_214_1447_0, i_10_214_1448_0,
    i_10_214_1651_0, i_10_214_1654_0, i_10_214_1680_0, i_10_214_1726_0,
    i_10_214_1816_0, i_10_214_1875_0, i_10_214_2019_0, i_10_214_2020_0,
    i_10_214_2022_0, i_10_214_2050_0, i_10_214_2253_0, i_10_214_2256_0,
    i_10_214_2257_0, i_10_214_2258_0, i_10_214_2259_0, i_10_214_2325_0,
    i_10_214_2354_0, i_10_214_2364_0, i_10_214_2454_0, i_10_214_2467_0,
    i_10_214_2514_0, i_10_214_2527_0, i_10_214_2546_0, i_10_214_2571_0,
    i_10_214_2660_0, i_10_214_2675_0, i_10_214_2787_0, i_10_214_2839_0,
    i_10_214_2913_0, i_10_214_2914_0, i_10_214_2979_0, i_10_214_3047_0,
    i_10_214_3237_0, i_10_214_3284_0, i_10_214_3291_0, i_10_214_3389_0,
    i_10_214_3399_0, i_10_214_3433_0, i_10_214_3495_0, i_10_214_3499_0,
    i_10_214_3583_0, i_10_214_3585_0, i_10_214_3586_0, i_10_214_3590_0,
    i_10_214_3687_0, i_10_214_3814_0, i_10_214_3837_0, i_10_214_3846_0,
    i_10_214_3855_0, i_10_214_3856_0, i_10_214_3873_0, i_10_214_3887_0,
    i_10_214_3945_0, i_10_214_3948_0, i_10_214_3973_0, i_10_214_4028_0,
    i_10_214_4055_0, i_10_214_4119_0, i_10_214_4123_0, i_10_214_4128_0,
    i_10_214_4220_0, i_10_214_4236_0, i_10_214_4267_0, i_10_214_4269_0;
  output o_10_214_0_0;
  assign o_10_214_0_0 = 0;
endmodule



// Benchmark "kernel_10_215" written by ABC on Sun Jul 19 10:24:43 2020

module kernel_10_215 ( 
    i_10_215_144_0, i_10_215_282_0, i_10_215_283_0, i_10_215_284_0,
    i_10_215_288_0, i_10_215_289_0, i_10_215_290_0, i_10_215_316_0,
    i_10_215_423_0, i_10_215_424_0, i_10_215_425_0, i_10_215_446_0,
    i_10_215_449_0, i_10_215_639_0, i_10_215_718_0, i_10_215_793_0,
    i_10_215_794_0, i_10_215_891_0, i_10_215_1003_0, i_10_215_1080_0,
    i_10_215_1083_0, i_10_215_1247_0, i_10_215_1262_0, i_10_215_1360_0,
    i_10_215_1440_0, i_10_215_1441_0, i_10_215_1442_0, i_10_215_1443_0,
    i_10_215_1444_0, i_10_215_1539_0, i_10_215_1543_0, i_10_215_1575_0,
    i_10_215_1576_0, i_10_215_1577_0, i_10_215_1579_0, i_10_215_1581_0,
    i_10_215_1653_0, i_10_215_1654_0, i_10_215_1679_0, i_10_215_1821_0,
    i_10_215_1822_0, i_10_215_1913_0, i_10_215_1945_0, i_10_215_1989_0,
    i_10_215_1990_0, i_10_215_2197_0, i_10_215_2200_0, i_10_215_2349_0,
    i_10_215_2351_0, i_10_215_2355_0, i_10_215_2362_0, i_10_215_2461_0,
    i_10_215_2659_0, i_10_215_2673_0, i_10_215_2674_0, i_10_215_2701_0,
    i_10_215_2709_0, i_10_215_2710_0, i_10_215_2711_0, i_10_215_2826_0,
    i_10_215_2881_0, i_10_215_2918_0, i_10_215_2920_0, i_10_215_3034_0,
    i_10_215_3038_0, i_10_215_3088_0, i_10_215_3196_0, i_10_215_3232_0,
    i_10_215_3267_0, i_10_215_3278_0, i_10_215_3294_0, i_10_215_3384_0,
    i_10_215_3405_0, i_10_215_3430_0, i_10_215_3431_0, i_10_215_3440_0,
    i_10_215_3522_0, i_10_215_3550_0, i_10_215_3584_0, i_10_215_3612_0,
    i_10_215_3614_0, i_10_215_3649_0, i_10_215_3781_0, i_10_215_3788_0,
    i_10_215_3835_0, i_10_215_3839_0, i_10_215_3859_0, i_10_215_3897_0,
    i_10_215_3910_0, i_10_215_3942_0, i_10_215_3990_0, i_10_215_3991_0,
    i_10_215_4051_0, i_10_215_4057_0, i_10_215_4119_0, i_10_215_4168_0,
    i_10_215_4276_0, i_10_215_4279_0, i_10_215_4565_0, i_10_215_4568_0,
    o_10_215_0_0  );
  input  i_10_215_144_0, i_10_215_282_0, i_10_215_283_0, i_10_215_284_0,
    i_10_215_288_0, i_10_215_289_0, i_10_215_290_0, i_10_215_316_0,
    i_10_215_423_0, i_10_215_424_0, i_10_215_425_0, i_10_215_446_0,
    i_10_215_449_0, i_10_215_639_0, i_10_215_718_0, i_10_215_793_0,
    i_10_215_794_0, i_10_215_891_0, i_10_215_1003_0, i_10_215_1080_0,
    i_10_215_1083_0, i_10_215_1247_0, i_10_215_1262_0, i_10_215_1360_0,
    i_10_215_1440_0, i_10_215_1441_0, i_10_215_1442_0, i_10_215_1443_0,
    i_10_215_1444_0, i_10_215_1539_0, i_10_215_1543_0, i_10_215_1575_0,
    i_10_215_1576_0, i_10_215_1577_0, i_10_215_1579_0, i_10_215_1581_0,
    i_10_215_1653_0, i_10_215_1654_0, i_10_215_1679_0, i_10_215_1821_0,
    i_10_215_1822_0, i_10_215_1913_0, i_10_215_1945_0, i_10_215_1989_0,
    i_10_215_1990_0, i_10_215_2197_0, i_10_215_2200_0, i_10_215_2349_0,
    i_10_215_2351_0, i_10_215_2355_0, i_10_215_2362_0, i_10_215_2461_0,
    i_10_215_2659_0, i_10_215_2673_0, i_10_215_2674_0, i_10_215_2701_0,
    i_10_215_2709_0, i_10_215_2710_0, i_10_215_2711_0, i_10_215_2826_0,
    i_10_215_2881_0, i_10_215_2918_0, i_10_215_2920_0, i_10_215_3034_0,
    i_10_215_3038_0, i_10_215_3088_0, i_10_215_3196_0, i_10_215_3232_0,
    i_10_215_3267_0, i_10_215_3278_0, i_10_215_3294_0, i_10_215_3384_0,
    i_10_215_3405_0, i_10_215_3430_0, i_10_215_3431_0, i_10_215_3440_0,
    i_10_215_3522_0, i_10_215_3550_0, i_10_215_3584_0, i_10_215_3612_0,
    i_10_215_3614_0, i_10_215_3649_0, i_10_215_3781_0, i_10_215_3788_0,
    i_10_215_3835_0, i_10_215_3839_0, i_10_215_3859_0, i_10_215_3897_0,
    i_10_215_3910_0, i_10_215_3942_0, i_10_215_3990_0, i_10_215_3991_0,
    i_10_215_4051_0, i_10_215_4057_0, i_10_215_4119_0, i_10_215_4168_0,
    i_10_215_4276_0, i_10_215_4279_0, i_10_215_4565_0, i_10_215_4568_0;
  output o_10_215_0_0;
  assign o_10_215_0_0 = ~((~i_10_215_2674_0 & ((~i_10_215_144_0 & ((~i_10_215_639_0 & ~i_10_215_1440_0 & ~i_10_215_1821_0 & ~i_10_215_1822_0 & ~i_10_215_1989_0 & ~i_10_215_2362_0 & ~i_10_215_2461_0) | (~i_10_215_289_0 & ~i_10_215_424_0 & ~i_10_215_1444_0 & ~i_10_215_1990_0 & ~i_10_215_3038_0 & ~i_10_215_3405_0 & ~i_10_215_3431_0 & ~i_10_215_3614_0))) | (~i_10_215_283_0 & ~i_10_215_425_0 & ~i_10_215_639_0 & ~i_10_215_891_0 & ~i_10_215_1441_0 & ~i_10_215_1443_0 & ~i_10_215_3088_0 & ~i_10_215_3550_0 & ~i_10_215_3584_0 & ~i_10_215_3859_0 & ~i_10_215_3942_0) | (~i_10_215_1654_0 & i_10_215_1821_0 & ~i_10_215_3430_0 & ~i_10_215_4057_0 & i_10_215_4119_0))) | (~i_10_215_284_0 & ((~i_10_215_1440_0 & ~i_10_215_1441_0 & ~i_10_215_1821_0 & ~i_10_215_1989_0 & ~i_10_215_2826_0 & ~i_10_215_2918_0 & ~i_10_215_3034_0 & ~i_10_215_3384_0 & ~i_10_215_3788_0 & ~i_10_215_3942_0 & ~i_10_215_4057_0) | (~i_10_215_423_0 & ~i_10_215_639_0 & ~i_10_215_1247_0 & ~i_10_215_3088_0 & ~i_10_215_3430_0 & ~i_10_215_3522_0 & ~i_10_215_3991_0 & ~i_10_215_4565_0))) | (~i_10_215_1443_0 & ((~i_10_215_282_0 & ~i_10_215_1990_0 & ~i_10_215_3088_0 & ((~i_10_215_289_0 & ~i_10_215_316_0 & ~i_10_215_424_0 & ~i_10_215_2711_0 & ~i_10_215_4057_0) | (~i_10_215_718_0 & ~i_10_215_1822_0 & i_10_215_3584_0 & ~i_10_215_3942_0 & ~i_10_215_4565_0))) | (~i_10_215_289_0 & ~i_10_215_290_0 & ~i_10_215_639_0 & i_10_215_2351_0) | (~i_10_215_1083_0 & ~i_10_215_1360_0 & ~i_10_215_2709_0 & ~i_10_215_2711_0 & ~i_10_215_2881_0 & ~i_10_215_3431_0 & i_10_215_3859_0 & ~i_10_215_4568_0))) | (~i_10_215_282_0 & ((~i_10_215_423_0 & ~i_10_215_639_0 & ~i_10_215_2362_0 & ~i_10_215_2709_0 & ~i_10_215_3584_0 & ~i_10_215_3990_0) | (i_10_215_1913_0 & ~i_10_215_2461_0 & i_10_215_4057_0))) | (~i_10_215_424_0 & ((~i_10_215_793_0 & ~i_10_215_1441_0 & ~i_10_215_1822_0 & ~i_10_215_1990_0 & ~i_10_215_3384_0 & i_10_215_3431_0) | (~i_10_215_3522_0 & ~i_10_215_3612_0 & ~i_10_215_4051_0 & ~i_10_215_4119_0 & ~i_10_215_4568_0))) | (~i_10_215_2362_0 & ((~i_10_215_1360_0 & ((~i_10_215_423_0 & ~i_10_215_425_0 & ~i_10_215_1441_0 & ~i_10_215_3430_0 & ~i_10_215_3550_0) | (~i_10_215_794_0 & ~i_10_215_3088_0 & i_10_215_3835_0 & ~i_10_215_3991_0))) | (i_10_215_1654_0 & ~i_10_215_2709_0 & ~i_10_215_3038_0 & ~i_10_215_3612_0 & ~i_10_215_3788_0 & ~i_10_215_3942_0))) | (~i_10_215_3088_0 & ((~i_10_215_423_0 & ~i_10_215_4057_0 & ((~i_10_215_1441_0 & i_10_215_2826_0 & ~i_10_215_3550_0 & ~i_10_215_3839_0) | (~i_10_215_1440_0 & ~i_10_215_1913_0 & ~i_10_215_2461_0 & ~i_10_215_2918_0 & ~i_10_215_3522_0 & ~i_10_215_3942_0 & ~i_10_215_4051_0))) | (~i_10_215_1247_0 & ~i_10_215_1440_0 & ~i_10_215_1444_0 & ~i_10_215_2709_0 & ~i_10_215_3267_0 & ~i_10_215_3405_0 & ~i_10_215_4051_0 & ~i_10_215_4568_0))) | (i_10_215_2355_0 & (i_10_215_1083_0 | (i_10_215_4057_0 & ~i_10_215_4568_0))) | (~i_10_215_1822_0 & ~i_10_215_2673_0 & i_10_215_3088_0 & ~i_10_215_3431_0 & i_10_215_3835_0) | (i_10_215_1581_0 & i_10_215_3649_0 & i_10_215_4119_0));
endmodule



// Benchmark "kernel_10_216" written by ABC on Sun Jul 19 10:24:43 2020

module kernel_10_216 ( 
    i_10_216_64_0, i_10_216_171_0, i_10_216_175_0, i_10_216_223_0,
    i_10_216_224_0, i_10_216_286_0, i_10_216_290_0, i_10_216_461_0,
    i_10_216_517_0, i_10_216_532_0, i_10_216_533_0, i_10_216_748_0,
    i_10_216_797_0, i_10_216_1026_0, i_10_216_1027_0, i_10_216_1029_0,
    i_10_216_1035_0, i_10_216_1236_0, i_10_216_1242_0, i_10_216_1243_0,
    i_10_216_1315_0, i_10_216_1547_0, i_10_216_1578_0, i_10_216_1579_0,
    i_10_216_1614_0, i_10_216_1687_0, i_10_216_1691_0, i_10_216_1822_0,
    i_10_216_1854_0, i_10_216_1915_0, i_10_216_1916_0, i_10_216_1954_0,
    i_10_216_1989_0, i_10_216_1991_0, i_10_216_1998_0, i_10_216_2151_0,
    i_10_216_2154_0, i_10_216_2179_0, i_10_216_2224_0, i_10_216_2304_0,
    i_10_216_2305_0, i_10_216_2307_0, i_10_216_2358_0, i_10_216_2361_0,
    i_10_216_2362_0, i_10_216_2364_0, i_10_216_2368_0, i_10_216_2448_0,
    i_10_216_2456_0, i_10_216_2457_0, i_10_216_2460_0, i_10_216_2461_0,
    i_10_216_2466_0, i_10_216_2467_0, i_10_216_2629_0, i_10_216_2631_0,
    i_10_216_2632_0, i_10_216_2677_0, i_10_216_2726_0, i_10_216_2730_0,
    i_10_216_2862_0, i_10_216_2983_0, i_10_216_3088_0, i_10_216_3196_0,
    i_10_216_3199_0, i_10_216_3231_0, i_10_216_3283_0, i_10_216_3303_0,
    i_10_216_3330_0, i_10_216_3333_0, i_10_216_3385_0, i_10_216_3442_0,
    i_10_216_3468_0, i_10_216_3520_0, i_10_216_3522_0, i_10_216_3609_0,
    i_10_216_3612_0, i_10_216_3613_0, i_10_216_3614_0, i_10_216_3681_0,
    i_10_216_3682_0, i_10_216_3684_0, i_10_216_3686_0, i_10_216_3840_0,
    i_10_216_3844_0, i_10_216_3856_0, i_10_216_3889_0, i_10_216_3930_0,
    i_10_216_3980_0, i_10_216_4024_0, i_10_216_4113_0, i_10_216_4124_0,
    i_10_216_4143_0, i_10_216_4212_0, i_10_216_4213_0, i_10_216_4216_0,
    i_10_216_4284_0, i_10_216_4350_0, i_10_216_4351_0, i_10_216_4590_0,
    o_10_216_0_0  );
  input  i_10_216_64_0, i_10_216_171_0, i_10_216_175_0, i_10_216_223_0,
    i_10_216_224_0, i_10_216_286_0, i_10_216_290_0, i_10_216_461_0,
    i_10_216_517_0, i_10_216_532_0, i_10_216_533_0, i_10_216_748_0,
    i_10_216_797_0, i_10_216_1026_0, i_10_216_1027_0, i_10_216_1029_0,
    i_10_216_1035_0, i_10_216_1236_0, i_10_216_1242_0, i_10_216_1243_0,
    i_10_216_1315_0, i_10_216_1547_0, i_10_216_1578_0, i_10_216_1579_0,
    i_10_216_1614_0, i_10_216_1687_0, i_10_216_1691_0, i_10_216_1822_0,
    i_10_216_1854_0, i_10_216_1915_0, i_10_216_1916_0, i_10_216_1954_0,
    i_10_216_1989_0, i_10_216_1991_0, i_10_216_1998_0, i_10_216_2151_0,
    i_10_216_2154_0, i_10_216_2179_0, i_10_216_2224_0, i_10_216_2304_0,
    i_10_216_2305_0, i_10_216_2307_0, i_10_216_2358_0, i_10_216_2361_0,
    i_10_216_2362_0, i_10_216_2364_0, i_10_216_2368_0, i_10_216_2448_0,
    i_10_216_2456_0, i_10_216_2457_0, i_10_216_2460_0, i_10_216_2461_0,
    i_10_216_2466_0, i_10_216_2467_0, i_10_216_2629_0, i_10_216_2631_0,
    i_10_216_2632_0, i_10_216_2677_0, i_10_216_2726_0, i_10_216_2730_0,
    i_10_216_2862_0, i_10_216_2983_0, i_10_216_3088_0, i_10_216_3196_0,
    i_10_216_3199_0, i_10_216_3231_0, i_10_216_3283_0, i_10_216_3303_0,
    i_10_216_3330_0, i_10_216_3333_0, i_10_216_3385_0, i_10_216_3442_0,
    i_10_216_3468_0, i_10_216_3520_0, i_10_216_3522_0, i_10_216_3609_0,
    i_10_216_3612_0, i_10_216_3613_0, i_10_216_3614_0, i_10_216_3681_0,
    i_10_216_3682_0, i_10_216_3684_0, i_10_216_3686_0, i_10_216_3840_0,
    i_10_216_3844_0, i_10_216_3856_0, i_10_216_3889_0, i_10_216_3930_0,
    i_10_216_3980_0, i_10_216_4024_0, i_10_216_4113_0, i_10_216_4124_0,
    i_10_216_4143_0, i_10_216_4212_0, i_10_216_4213_0, i_10_216_4216_0,
    i_10_216_4284_0, i_10_216_4350_0, i_10_216_4351_0, i_10_216_4590_0;
  output o_10_216_0_0;
  assign o_10_216_0_0 = 0;
endmodule



// Benchmark "kernel_10_217" written by ABC on Sun Jul 19 10:24:45 2020

module kernel_10_217 ( 
    i_10_217_172_0, i_10_217_177_0, i_10_217_223_0, i_10_217_283_0,
    i_10_217_316_0, i_10_217_318_0, i_10_217_330_0, i_10_217_409_0,
    i_10_217_410_0, i_10_217_411_0, i_10_217_412_0, i_10_217_413_0,
    i_10_217_512_0, i_10_217_993_0, i_10_217_1236_0, i_10_217_1238_0,
    i_10_217_1239_0, i_10_217_1240_0, i_10_217_1241_0, i_10_217_1243_0,
    i_10_217_1310_0, i_10_217_1365_0, i_10_217_1549_0, i_10_217_1552_0,
    i_10_217_1577_0, i_10_217_1581_0, i_10_217_1647_0, i_10_217_1683_0,
    i_10_217_1687_0, i_10_217_1820_0, i_10_217_1821_0, i_10_217_1945_0,
    i_10_217_2244_0, i_10_217_2339_0, i_10_217_2353_0, i_10_217_2381_0,
    i_10_217_2451_0, i_10_217_2453_0, i_10_217_2455_0, i_10_217_2466_0,
    i_10_217_2467_0, i_10_217_2468_0, i_10_217_2469_0, i_10_217_2473_0,
    i_10_217_2629_0, i_10_217_2630_0, i_10_217_2631_0, i_10_217_2632_0,
    i_10_217_2633_0, i_10_217_2635_0, i_10_217_2636_0, i_10_217_2659_0,
    i_10_217_2674_0, i_10_217_2703_0, i_10_217_2706_0, i_10_217_2728_0,
    i_10_217_2731_0, i_10_217_2732_0, i_10_217_2733_0, i_10_217_2781_0,
    i_10_217_2782_0, i_10_217_2785_0, i_10_217_2787_0, i_10_217_2788_0,
    i_10_217_2827_0, i_10_217_2834_0, i_10_217_2886_0, i_10_217_3042_0,
    i_10_217_3043_0, i_10_217_3044_0, i_10_217_3047_0, i_10_217_3151_0,
    i_10_217_3157_0, i_10_217_3158_0, i_10_217_3198_0, i_10_217_3237_0,
    i_10_217_3405_0, i_10_217_3408_0, i_10_217_3468_0, i_10_217_3472_0,
    i_10_217_3582_0, i_10_217_3585_0, i_10_217_3586_0, i_10_217_3588_0,
    i_10_217_3589_0, i_10_217_3617_0, i_10_217_3651_0, i_10_217_3652_0,
    i_10_217_3781_0, i_10_217_3785_0, i_10_217_3847_0, i_10_217_3853_0,
    i_10_217_3907_0, i_10_217_4054_0, i_10_217_4118_0, i_10_217_4119_0,
    i_10_217_4289_0, i_10_217_4292_0, i_10_217_4567_0, i_10_217_4584_0,
    o_10_217_0_0  );
  input  i_10_217_172_0, i_10_217_177_0, i_10_217_223_0, i_10_217_283_0,
    i_10_217_316_0, i_10_217_318_0, i_10_217_330_0, i_10_217_409_0,
    i_10_217_410_0, i_10_217_411_0, i_10_217_412_0, i_10_217_413_0,
    i_10_217_512_0, i_10_217_993_0, i_10_217_1236_0, i_10_217_1238_0,
    i_10_217_1239_0, i_10_217_1240_0, i_10_217_1241_0, i_10_217_1243_0,
    i_10_217_1310_0, i_10_217_1365_0, i_10_217_1549_0, i_10_217_1552_0,
    i_10_217_1577_0, i_10_217_1581_0, i_10_217_1647_0, i_10_217_1683_0,
    i_10_217_1687_0, i_10_217_1820_0, i_10_217_1821_0, i_10_217_1945_0,
    i_10_217_2244_0, i_10_217_2339_0, i_10_217_2353_0, i_10_217_2381_0,
    i_10_217_2451_0, i_10_217_2453_0, i_10_217_2455_0, i_10_217_2466_0,
    i_10_217_2467_0, i_10_217_2468_0, i_10_217_2469_0, i_10_217_2473_0,
    i_10_217_2629_0, i_10_217_2630_0, i_10_217_2631_0, i_10_217_2632_0,
    i_10_217_2633_0, i_10_217_2635_0, i_10_217_2636_0, i_10_217_2659_0,
    i_10_217_2674_0, i_10_217_2703_0, i_10_217_2706_0, i_10_217_2728_0,
    i_10_217_2731_0, i_10_217_2732_0, i_10_217_2733_0, i_10_217_2781_0,
    i_10_217_2782_0, i_10_217_2785_0, i_10_217_2787_0, i_10_217_2788_0,
    i_10_217_2827_0, i_10_217_2834_0, i_10_217_2886_0, i_10_217_3042_0,
    i_10_217_3043_0, i_10_217_3044_0, i_10_217_3047_0, i_10_217_3151_0,
    i_10_217_3157_0, i_10_217_3158_0, i_10_217_3198_0, i_10_217_3237_0,
    i_10_217_3405_0, i_10_217_3408_0, i_10_217_3468_0, i_10_217_3472_0,
    i_10_217_3582_0, i_10_217_3585_0, i_10_217_3586_0, i_10_217_3588_0,
    i_10_217_3589_0, i_10_217_3617_0, i_10_217_3651_0, i_10_217_3652_0,
    i_10_217_3781_0, i_10_217_3785_0, i_10_217_3847_0, i_10_217_3853_0,
    i_10_217_3907_0, i_10_217_4054_0, i_10_217_4118_0, i_10_217_4119_0,
    i_10_217_4289_0, i_10_217_4292_0, i_10_217_4567_0, i_10_217_4584_0;
  output o_10_217_0_0;
  assign o_10_217_0_0 = ~((~i_10_217_3588_0 & ((~i_10_217_283_0 & ((~i_10_217_1241_0 & ~i_10_217_2733_0 & ~i_10_217_3042_0 & ~i_10_217_3585_0 & ~i_10_217_3586_0) | (~i_10_217_412_0 & ~i_10_217_413_0 & ~i_10_217_1365_0 & ~i_10_217_2469_0 & ~i_10_217_2674_0 & ~i_10_217_2785_0 & ~i_10_217_3582_0 & ~i_10_217_4054_0))) | (~i_10_217_2466_0 & ((~i_10_217_318_0 & ~i_10_217_411_0 & ~i_10_217_1241_0 & i_10_217_2728_0) | (~i_10_217_1239_0 & ~i_10_217_2469_0 & ~i_10_217_2473_0 & i_10_217_2731_0 & ~i_10_217_2785_0 & ~i_10_217_3237_0))))) | (~i_10_217_1581_0 & ((~i_10_217_409_0 & ((~i_10_217_318_0 & ~i_10_217_412_0 & ~i_10_217_1236_0 & ~i_10_217_1365_0 & ~i_10_217_2467_0 & ~i_10_217_2787_0 & ~i_10_217_3237_0 & ~i_10_217_3468_0 & ~i_10_217_3781_0) | (~i_10_217_1821_0 & ~i_10_217_2732_0 & ~i_10_217_2781_0 & ~i_10_217_3585_0 & ~i_10_217_4054_0))) | (i_10_217_316_0 & i_10_217_1238_0 & ~i_10_217_2732_0 & ~i_10_217_2781_0 & ~i_10_217_3585_0))) | (~i_10_217_318_0 & ((~i_10_217_1236_0 & ~i_10_217_2473_0 & ~i_10_217_2733_0 & ~i_10_217_2781_0 & ~i_10_217_2782_0 & ~i_10_217_2788_0) | (~i_10_217_993_0 & ~i_10_217_1945_0 & ~i_10_217_2451_0 & ~i_10_217_2468_0 & ~i_10_217_2827_0 & ~i_10_217_3198_0 & ~i_10_217_3237_0 & ~i_10_217_3472_0 & ~i_10_217_3586_0 & ~i_10_217_3853_0 & ~i_10_217_4119_0 & ~i_10_217_4292_0))) | (~i_10_217_1239_0 & ((~i_10_217_412_0 & i_10_217_2732_0 & i_10_217_2733_0 & ~i_10_217_2788_0 & ~i_10_217_3468_0) | (i_10_217_2632_0 & ~i_10_217_2733_0 & ~i_10_217_2782_0 & ~i_10_217_3785_0))) | (~i_10_217_1310_0 & ((i_10_217_993_0 & i_10_217_3198_0) | (~i_10_217_411_0 & ~i_10_217_2469_0 & i_10_217_2732_0 & ~i_10_217_2788_0 & ~i_10_217_3472_0 & ~i_10_217_3582_0))) | (~i_10_217_411_0 & ((i_10_217_2630_0 & ~i_10_217_2787_0 & ~i_10_217_3043_0 & ~i_10_217_3237_0) | (~i_10_217_410_0 & ~i_10_217_1945_0 & i_10_217_2659_0 & ~i_10_217_3472_0 & ~i_10_217_3585_0 & ~i_10_217_4054_0))) | (i_10_217_2632_0 & ((i_10_217_2453_0 & ~i_10_217_3043_0 & ~i_10_217_3468_0) | (~i_10_217_330_0 & ~i_10_217_1365_0 & ~i_10_217_1945_0 & ~i_10_217_2469_0 & ~i_10_217_2787_0 & ~i_10_217_3047_0 & ~i_10_217_3237_0 & ~i_10_217_4054_0))) | (~i_10_217_3585_0 & ((~i_10_217_177_0 & ~i_10_217_2782_0 & ((~i_10_217_1238_0 & ~i_10_217_1365_0 & ~i_10_217_2827_0 & ~i_10_217_3043_0 & ~i_10_217_3047_0 & ~i_10_217_3472_0) | (~i_10_217_2469_0 & i_10_217_4289_0 & ~i_10_217_4567_0))) | (~i_10_217_1365_0 & ~i_10_217_2451_0 & ~i_10_217_2827_0 & ~i_10_217_3472_0 & ~i_10_217_3582_0 & ~i_10_217_3589_0 & ~i_10_217_4054_0 & ~i_10_217_4567_0))) | (~i_10_217_2781_0 & ((~i_10_217_2469_0 & ~i_10_217_2473_0 & ~i_10_217_177_0 & ~i_10_217_413_0 & ~i_10_217_2788_0 & ~i_10_217_2886_0 & ~i_10_217_3042_0 & ~i_10_217_3237_0) | (i_10_217_172_0 & ~i_10_217_1240_0 & i_10_217_2467_0 & i_10_217_3847_0))) | (~i_10_217_172_0 & i_10_217_1687_0 & i_10_217_1821_0 & ~i_10_217_2353_0 & ~i_10_217_2674_0 & ~i_10_217_2703_0 & ~i_10_217_2733_0 & ~i_10_217_3044_0 & ~i_10_217_3047_0 & ~i_10_217_3785_0));
endmodule



// Benchmark "kernel_10_218" written by ABC on Sun Jul 19 10:24:46 2020

module kernel_10_218 ( 
    i_10_218_42_0, i_10_218_89_0, i_10_218_180_0, i_10_218_181_0,
    i_10_218_183_0, i_10_218_184_0, i_10_218_250_0, i_10_218_280_0,
    i_10_218_287_0, i_10_218_292_0, i_10_218_293_0, i_10_218_408_0,
    i_10_218_409_0, i_10_218_412_0, i_10_218_426_0, i_10_218_436_0,
    i_10_218_444_0, i_10_218_795_0, i_10_218_796_0, i_10_218_798_0,
    i_10_218_957_0, i_10_218_958_0, i_10_218_997_0, i_10_218_1119_0,
    i_10_218_1167_0, i_10_218_1168_0, i_10_218_1237_0, i_10_218_1238_0,
    i_10_218_1239_0, i_10_218_1240_0, i_10_218_1247_0, i_10_218_1249_0,
    i_10_218_1250_0, i_10_218_1354_0, i_10_218_1363_0, i_10_218_1543_0,
    i_10_218_1758_0, i_10_218_1763_0, i_10_218_1824_0, i_10_218_1826_0,
    i_10_218_1909_0, i_10_218_1915_0, i_10_218_1995_0, i_10_218_1996_0,
    i_10_218_2005_0, i_10_218_2022_0, i_10_218_2023_0, i_10_218_2334_0,
    i_10_218_2353_0, i_10_218_2474_0, i_10_218_2608_0, i_10_218_2629_0,
    i_10_218_2633_0, i_10_218_2636_0, i_10_218_2677_0, i_10_218_2707_0,
    i_10_218_2719_0, i_10_218_2721_0, i_10_218_2722_0, i_10_218_2723_0,
    i_10_218_2729_0, i_10_218_2785_0, i_10_218_2788_0, i_10_218_2827_0,
    i_10_218_2829_0, i_10_218_2830_0, i_10_218_2923_0, i_10_218_2924_0,
    i_10_218_2983_0, i_10_218_3038_0, i_10_218_3048_0, i_10_218_3076_0,
    i_10_218_3270_0, i_10_218_3271_0, i_10_218_3283_0, i_10_218_3385_0,
    i_10_218_3387_0, i_10_218_3433_0, i_10_218_3612_0, i_10_218_3647_0,
    i_10_218_3649_0, i_10_218_3688_0, i_10_218_3689_0, i_10_218_3720_0,
    i_10_218_3835_0, i_10_218_3836_0, i_10_218_3841_0, i_10_218_3886_0,
    i_10_218_3982_0, i_10_218_3986_0, i_10_218_4027_0, i_10_218_4095_0,
    i_10_218_4120_0, i_10_218_4153_0, i_10_218_4180_0, i_10_218_4188_0,
    i_10_218_4189_0, i_10_218_4191_0, i_10_218_4272_0, i_10_218_4565_0,
    o_10_218_0_0  );
  input  i_10_218_42_0, i_10_218_89_0, i_10_218_180_0, i_10_218_181_0,
    i_10_218_183_0, i_10_218_184_0, i_10_218_250_0, i_10_218_280_0,
    i_10_218_287_0, i_10_218_292_0, i_10_218_293_0, i_10_218_408_0,
    i_10_218_409_0, i_10_218_412_0, i_10_218_426_0, i_10_218_436_0,
    i_10_218_444_0, i_10_218_795_0, i_10_218_796_0, i_10_218_798_0,
    i_10_218_957_0, i_10_218_958_0, i_10_218_997_0, i_10_218_1119_0,
    i_10_218_1167_0, i_10_218_1168_0, i_10_218_1237_0, i_10_218_1238_0,
    i_10_218_1239_0, i_10_218_1240_0, i_10_218_1247_0, i_10_218_1249_0,
    i_10_218_1250_0, i_10_218_1354_0, i_10_218_1363_0, i_10_218_1543_0,
    i_10_218_1758_0, i_10_218_1763_0, i_10_218_1824_0, i_10_218_1826_0,
    i_10_218_1909_0, i_10_218_1915_0, i_10_218_1995_0, i_10_218_1996_0,
    i_10_218_2005_0, i_10_218_2022_0, i_10_218_2023_0, i_10_218_2334_0,
    i_10_218_2353_0, i_10_218_2474_0, i_10_218_2608_0, i_10_218_2629_0,
    i_10_218_2633_0, i_10_218_2636_0, i_10_218_2677_0, i_10_218_2707_0,
    i_10_218_2719_0, i_10_218_2721_0, i_10_218_2722_0, i_10_218_2723_0,
    i_10_218_2729_0, i_10_218_2785_0, i_10_218_2788_0, i_10_218_2827_0,
    i_10_218_2829_0, i_10_218_2830_0, i_10_218_2923_0, i_10_218_2924_0,
    i_10_218_2983_0, i_10_218_3038_0, i_10_218_3048_0, i_10_218_3076_0,
    i_10_218_3270_0, i_10_218_3271_0, i_10_218_3283_0, i_10_218_3385_0,
    i_10_218_3387_0, i_10_218_3433_0, i_10_218_3612_0, i_10_218_3647_0,
    i_10_218_3649_0, i_10_218_3688_0, i_10_218_3689_0, i_10_218_3720_0,
    i_10_218_3835_0, i_10_218_3836_0, i_10_218_3841_0, i_10_218_3886_0,
    i_10_218_3982_0, i_10_218_3986_0, i_10_218_4027_0, i_10_218_4095_0,
    i_10_218_4120_0, i_10_218_4153_0, i_10_218_4180_0, i_10_218_4188_0,
    i_10_218_4189_0, i_10_218_4191_0, i_10_218_4272_0, i_10_218_4565_0;
  output o_10_218_0_0;
  assign o_10_218_0_0 = ~((~i_10_218_183_0 & ((~i_10_218_250_0 & ~i_10_218_795_0 & ~i_10_218_1237_0 & ~i_10_218_1249_0 & ~i_10_218_3048_0 & ~i_10_218_3283_0 & ~i_10_218_3649_0 & ~i_10_218_3689_0 & i_10_218_3835_0) | (~i_10_218_1168_0 & ~i_10_218_1238_0 & ~i_10_218_2005_0 & ~i_10_218_2719_0 & ~i_10_218_2722_0 & ~i_10_218_3271_0 & ~i_10_218_4272_0 & ~i_10_218_4565_0))) | (~i_10_218_287_0 & ((~i_10_218_280_0 & ~i_10_218_426_0 & ~i_10_218_436_0 & i_10_218_444_0 & ~i_10_218_1250_0 & ~i_10_218_2827_0 & ~i_10_218_2830_0 & ~i_10_218_3385_0 & ~i_10_218_3433_0) | (~i_10_218_409_0 & ~i_10_218_1363_0 & ~i_10_218_1996_0 & ~i_10_218_2005_0 & ~i_10_218_2608_0 & ~i_10_218_2707_0 & ~i_10_218_2719_0 & ~i_10_218_2983_0 & ~i_10_218_3841_0))) | (~i_10_218_292_0 & ((~i_10_218_89_0 & ~i_10_218_444_0 & i_10_218_2677_0 & ~i_10_218_3433_0 & i_10_218_3612_0) | (~i_10_218_184_0 & ~i_10_218_293_0 & ~i_10_218_426_0 & ~i_10_218_1363_0 & ~i_10_218_1995_0 & ~i_10_218_1996_0 & ~i_10_218_2023_0 & ~i_10_218_2729_0 & ~i_10_218_2983_0 & ~i_10_218_3038_0 & ~i_10_218_3986_0))) | (~i_10_218_408_0 & ((~i_10_218_280_0 & ~i_10_218_409_0 & ~i_10_218_1995_0 & ~i_10_218_1996_0 & ~i_10_218_2633_0 & ~i_10_218_2924_0) | (~i_10_218_1250_0 & ~i_10_218_2677_0 & ~i_10_218_2830_0 & ~i_10_218_2923_0 & i_10_218_3612_0))) | (~i_10_218_409_0 & ((~i_10_218_180_0 & ~i_10_218_997_0 & ~i_10_218_1247_0 & ~i_10_218_2723_0 & ~i_10_218_3689_0) | (~i_10_218_795_0 & ~i_10_218_1237_0 & ~i_10_218_1249_0 & ~i_10_218_1915_0 & ~i_10_218_3688_0 & ~i_10_218_3835_0 & ~i_10_218_3841_0))) | (~i_10_218_3689_0 & ((~i_10_218_3433_0 & ((~i_10_218_184_0 & ((~i_10_218_1250_0 & ~i_10_218_1824_0 & ~i_10_218_1909_0 & ~i_10_218_2022_0 & ~i_10_218_3076_0 & ~i_10_218_3612_0) | (~i_10_218_426_0 & ~i_10_218_796_0 & i_10_218_2830_0 & ~i_10_218_3688_0))) | (~i_10_218_795_0 & ~i_10_218_997_0 & ~i_10_218_1168_0 & ~i_10_218_1826_0 & ~i_10_218_2722_0 & ~i_10_218_3270_0 & ~i_10_218_3612_0))) | (~i_10_218_250_0 & ~i_10_218_280_0 & ~i_10_218_1168_0 & ~i_10_218_1247_0 & ~i_10_218_1250_0 & ~i_10_218_1996_0 & ~i_10_218_2827_0))) | (~i_10_218_1247_0 & ((~i_10_218_89_0 & ~i_10_218_3433_0 & ((~i_10_218_184_0 & ~i_10_218_293_0 & ~i_10_218_795_0 & ~i_10_218_2474_0 & ~i_10_218_3385_0 & ~i_10_218_3387_0) | (~i_10_218_250_0 & ~i_10_218_1240_0 & ~i_10_218_2005_0 & ~i_10_218_2721_0 & ~i_10_218_2788_0 & ~i_10_218_2829_0 & ~i_10_218_3688_0))) | (~i_10_218_184_0 & i_10_218_796_0 & ~i_10_218_2707_0 & ~i_10_218_2924_0 & ~i_10_218_3076_0 & ~i_10_218_3271_0 & i_10_218_3387_0 & ~i_10_218_3612_0 & ~i_10_218_3982_0))) | (~i_10_218_250_0 & ((~i_10_218_1239_0 & i_10_218_1824_0 & ~i_10_218_2629_0 & ~i_10_218_3270_0 & i_10_218_3387_0 & ~i_10_218_3836_0) | (~i_10_218_798_0 & ~i_10_218_997_0 & ~i_10_218_1995_0 & ~i_10_218_3271_0 & ~i_10_218_3433_0 & i_10_218_4027_0))) | (~i_10_218_280_0 & ((~i_10_218_958_0 & ~i_10_218_1237_0 & ~i_10_218_2636_0 & i_10_218_2719_0) | (~i_10_218_795_0 & ~i_10_218_997_0 & ~i_10_218_2830_0 & i_10_218_2923_0 & ~i_10_218_3433_0 & ~i_10_218_3612_0 & ~i_10_218_4120_0 & ~i_10_218_4565_0))) | (~i_10_218_1915_0 & ((~i_10_218_1237_0 & ~i_10_218_1363_0 & i_10_218_1824_0 & ~i_10_218_1909_0) | (~i_10_218_1239_0 & ~i_10_218_1249_0 & i_10_218_2983_0))) | (~i_10_218_2729_0 & ((~i_10_218_795_0 & i_10_218_1543_0 & ~i_10_218_2707_0) | (i_10_218_436_0 & i_10_218_2830_0 & ~i_10_218_3283_0 & i_10_218_3982_0 & i_10_218_3986_0))) | (~i_10_218_3433_0 & ~i_10_218_3835_0 & ((~i_10_218_1238_0 & ~i_10_218_2636_0 & i_10_218_2830_0) | (~i_10_218_181_0 & i_10_218_1826_0 & ~i_10_218_2785_0 & i_10_218_2827_0 & ~i_10_218_3841_0))) | (~i_10_218_89_0 & i_10_218_2636_0 & ~i_10_218_2829_0 & ~i_10_218_3038_0 & ~i_10_218_3385_0 & ~i_10_218_3841_0 & ~i_10_218_4027_0 & i_10_218_4120_0));
endmodule



// Benchmark "kernel_10_219" written by ABC on Sun Jul 19 10:24:47 2020

module kernel_10_219 ( 
    i_10_219_34_0, i_10_219_66_0, i_10_219_174_0, i_10_219_175_0,
    i_10_219_197_0, i_10_219_260_0, i_10_219_268_0, i_10_219_269_0,
    i_10_219_499_0, i_10_219_538_0, i_10_219_718_0, i_10_219_797_0,
    i_10_219_966_0, i_10_219_967_0, i_10_219_971_0, i_10_219_1030_0,
    i_10_219_1195_0, i_10_219_1196_0, i_10_219_1223_0, i_10_219_1241_0,
    i_10_219_1276_0, i_10_219_1277_0, i_10_219_1285_0, i_10_219_1302_0,
    i_10_219_1545_0, i_10_219_1556_0, i_10_219_1618_0, i_10_219_1641_0,
    i_10_219_1696_0, i_10_219_1697_0, i_10_219_1766_0, i_10_219_1767_0,
    i_10_219_1769_0, i_10_219_1822_0, i_10_219_1908_0, i_10_219_1943_0,
    i_10_219_1949_0, i_10_219_1957_0, i_10_219_2022_0, i_10_219_2023_0,
    i_10_219_2032_0, i_10_219_2033_0, i_10_219_2192_0, i_10_219_2203_0,
    i_10_219_2204_0, i_10_219_2348_0, i_10_219_2355_0, i_10_219_2356_0,
    i_10_219_2357_0, i_10_219_2456_0, i_10_219_2572_0, i_10_219_2580_0,
    i_10_219_2591_0, i_10_219_2599_0, i_10_219_2636_0, i_10_219_2705_0,
    i_10_219_2734_0, i_10_219_2761_0, i_10_219_2784_0, i_10_219_2785_0,
    i_10_219_2869_0, i_10_219_2883_0, i_10_219_2923_0, i_10_219_2959_0,
    i_10_219_2986_0, i_10_219_3026_0, i_10_219_3058_0, i_10_219_3059_0,
    i_10_219_3273_0, i_10_219_3281_0, i_10_219_3329_0, i_10_219_3473_0,
    i_10_219_3506_0, i_10_219_3571_0, i_10_219_3586_0, i_10_219_3605_0,
    i_10_219_3608_0, i_10_219_3616_0, i_10_219_3688_0, i_10_219_3839_0,
    i_10_219_3977_0, i_10_219_3984_0, i_10_219_3985_0, i_10_219_4013_0,
    i_10_219_4094_0, i_10_219_4126_0, i_10_219_4173_0, i_10_219_4183_0,
    i_10_219_4271_0, i_10_219_4272_0, i_10_219_4280_0, i_10_219_4281_0,
    i_10_219_4282_0, i_10_219_4283_0, i_10_219_4360_0, i_10_219_4379_0,
    i_10_219_4381_0, i_10_219_4461_0, i_10_219_4568_0, i_10_219_4569_0,
    o_10_219_0_0  );
  input  i_10_219_34_0, i_10_219_66_0, i_10_219_174_0, i_10_219_175_0,
    i_10_219_197_0, i_10_219_260_0, i_10_219_268_0, i_10_219_269_0,
    i_10_219_499_0, i_10_219_538_0, i_10_219_718_0, i_10_219_797_0,
    i_10_219_966_0, i_10_219_967_0, i_10_219_971_0, i_10_219_1030_0,
    i_10_219_1195_0, i_10_219_1196_0, i_10_219_1223_0, i_10_219_1241_0,
    i_10_219_1276_0, i_10_219_1277_0, i_10_219_1285_0, i_10_219_1302_0,
    i_10_219_1545_0, i_10_219_1556_0, i_10_219_1618_0, i_10_219_1641_0,
    i_10_219_1696_0, i_10_219_1697_0, i_10_219_1766_0, i_10_219_1767_0,
    i_10_219_1769_0, i_10_219_1822_0, i_10_219_1908_0, i_10_219_1943_0,
    i_10_219_1949_0, i_10_219_1957_0, i_10_219_2022_0, i_10_219_2023_0,
    i_10_219_2032_0, i_10_219_2033_0, i_10_219_2192_0, i_10_219_2203_0,
    i_10_219_2204_0, i_10_219_2348_0, i_10_219_2355_0, i_10_219_2356_0,
    i_10_219_2357_0, i_10_219_2456_0, i_10_219_2572_0, i_10_219_2580_0,
    i_10_219_2591_0, i_10_219_2599_0, i_10_219_2636_0, i_10_219_2705_0,
    i_10_219_2734_0, i_10_219_2761_0, i_10_219_2784_0, i_10_219_2785_0,
    i_10_219_2869_0, i_10_219_2883_0, i_10_219_2923_0, i_10_219_2959_0,
    i_10_219_2986_0, i_10_219_3026_0, i_10_219_3058_0, i_10_219_3059_0,
    i_10_219_3273_0, i_10_219_3281_0, i_10_219_3329_0, i_10_219_3473_0,
    i_10_219_3506_0, i_10_219_3571_0, i_10_219_3586_0, i_10_219_3605_0,
    i_10_219_3608_0, i_10_219_3616_0, i_10_219_3688_0, i_10_219_3839_0,
    i_10_219_3977_0, i_10_219_3984_0, i_10_219_3985_0, i_10_219_4013_0,
    i_10_219_4094_0, i_10_219_4126_0, i_10_219_4173_0, i_10_219_4183_0,
    i_10_219_4271_0, i_10_219_4272_0, i_10_219_4280_0, i_10_219_4281_0,
    i_10_219_4282_0, i_10_219_4283_0, i_10_219_4360_0, i_10_219_4379_0,
    i_10_219_4381_0, i_10_219_4461_0, i_10_219_4568_0, i_10_219_4569_0;
  output o_10_219_0_0;
  assign o_10_219_0_0 = 0;
endmodule



// Benchmark "kernel_10_220" written by ABC on Sun Jul 19 10:24:48 2020

module kernel_10_220 ( 
    i_10_220_51_0, i_10_220_88_0, i_10_220_150_0, i_10_220_186_0,
    i_10_220_187_0, i_10_220_258_0, i_10_220_269_0, i_10_220_372_0,
    i_10_220_408_0, i_10_220_464_0, i_10_220_565_0, i_10_220_642_0,
    i_10_220_762_0, i_10_220_793_0, i_10_220_794_0, i_10_220_826_0,
    i_10_220_853_0, i_10_220_854_0, i_10_220_898_0, i_10_220_996_0,
    i_10_220_1083_0, i_10_220_1086_0, i_10_220_1223_0, i_10_220_1305_0,
    i_10_220_1309_0, i_10_220_1396_0, i_10_220_1443_0, i_10_220_1551_0,
    i_10_220_1555_0, i_10_220_1556_0, i_10_220_1635_0, i_10_220_1636_0,
    i_10_220_1650_0, i_10_220_1651_0, i_10_220_1652_0, i_10_220_1653_0,
    i_10_220_1691_0, i_10_220_1713_0, i_10_220_1714_0, i_10_220_1732_0,
    i_10_220_1822_0, i_10_220_1883_0, i_10_220_1984_0, i_10_220_1986_0,
    i_10_220_2014_0, i_10_220_2026_0, i_10_220_2062_0, i_10_220_2157_0,
    i_10_220_2159_0, i_10_220_2227_0, i_10_220_2266_0, i_10_220_2290_0,
    i_10_220_2339_0, i_10_220_2365_0, i_10_220_2446_0, i_10_220_2451_0,
    i_10_220_2465_0, i_10_220_2568_0, i_10_220_2572_0, i_10_220_2634_0,
    i_10_220_2652_0, i_10_220_2661_0, i_10_220_2680_0, i_10_220_2711_0,
    i_10_220_2717_0, i_10_220_2730_0, i_10_220_2731_0, i_10_220_2734_0,
    i_10_220_2806_0, i_10_220_2850_0, i_10_220_3040_0, i_10_220_3091_0,
    i_10_220_3165_0, i_10_220_3166_0, i_10_220_3174_0, i_10_220_3273_0,
    i_10_220_3391_0, i_10_220_3408_0, i_10_220_3409_0, i_10_220_3410_0,
    i_10_220_3561_0, i_10_220_3611_0, i_10_220_3612_0, i_10_220_3613_0,
    i_10_220_3642_0, i_10_220_3803_0, i_10_220_3813_0, i_10_220_3854_0,
    i_10_220_3855_0, i_10_220_3856_0, i_10_220_3905_0, i_10_220_3923_0,
    i_10_220_4102_0, i_10_220_4120_0, i_10_220_4157_0, i_10_220_4174_0,
    i_10_220_4191_0, i_10_220_4269_0, i_10_220_4287_0, i_10_220_4552_0,
    o_10_220_0_0  );
  input  i_10_220_51_0, i_10_220_88_0, i_10_220_150_0, i_10_220_186_0,
    i_10_220_187_0, i_10_220_258_0, i_10_220_269_0, i_10_220_372_0,
    i_10_220_408_0, i_10_220_464_0, i_10_220_565_0, i_10_220_642_0,
    i_10_220_762_0, i_10_220_793_0, i_10_220_794_0, i_10_220_826_0,
    i_10_220_853_0, i_10_220_854_0, i_10_220_898_0, i_10_220_996_0,
    i_10_220_1083_0, i_10_220_1086_0, i_10_220_1223_0, i_10_220_1305_0,
    i_10_220_1309_0, i_10_220_1396_0, i_10_220_1443_0, i_10_220_1551_0,
    i_10_220_1555_0, i_10_220_1556_0, i_10_220_1635_0, i_10_220_1636_0,
    i_10_220_1650_0, i_10_220_1651_0, i_10_220_1652_0, i_10_220_1653_0,
    i_10_220_1691_0, i_10_220_1713_0, i_10_220_1714_0, i_10_220_1732_0,
    i_10_220_1822_0, i_10_220_1883_0, i_10_220_1984_0, i_10_220_1986_0,
    i_10_220_2014_0, i_10_220_2026_0, i_10_220_2062_0, i_10_220_2157_0,
    i_10_220_2159_0, i_10_220_2227_0, i_10_220_2266_0, i_10_220_2290_0,
    i_10_220_2339_0, i_10_220_2365_0, i_10_220_2446_0, i_10_220_2451_0,
    i_10_220_2465_0, i_10_220_2568_0, i_10_220_2572_0, i_10_220_2634_0,
    i_10_220_2652_0, i_10_220_2661_0, i_10_220_2680_0, i_10_220_2711_0,
    i_10_220_2717_0, i_10_220_2730_0, i_10_220_2731_0, i_10_220_2734_0,
    i_10_220_2806_0, i_10_220_2850_0, i_10_220_3040_0, i_10_220_3091_0,
    i_10_220_3165_0, i_10_220_3166_0, i_10_220_3174_0, i_10_220_3273_0,
    i_10_220_3391_0, i_10_220_3408_0, i_10_220_3409_0, i_10_220_3410_0,
    i_10_220_3561_0, i_10_220_3611_0, i_10_220_3612_0, i_10_220_3613_0,
    i_10_220_3642_0, i_10_220_3803_0, i_10_220_3813_0, i_10_220_3854_0,
    i_10_220_3855_0, i_10_220_3856_0, i_10_220_3905_0, i_10_220_3923_0,
    i_10_220_4102_0, i_10_220_4120_0, i_10_220_4157_0, i_10_220_4174_0,
    i_10_220_4191_0, i_10_220_4269_0, i_10_220_4287_0, i_10_220_4552_0;
  output o_10_220_0_0;
  assign o_10_220_0_0 = 0;
endmodule



// Benchmark "kernel_10_221" written by ABC on Sun Jul 19 10:24:49 2020

module kernel_10_221 ( 
    i_10_221_34_0, i_10_221_172_0, i_10_221_224_0, i_10_221_247_0,
    i_10_221_259_0, i_10_221_280_0, i_10_221_283_0, i_10_221_319_0,
    i_10_221_409_0, i_10_221_410_0, i_10_221_447_0, i_10_221_448_0,
    i_10_221_466_0, i_10_221_749_0, i_10_221_752_0, i_10_221_792_0,
    i_10_221_795_0, i_10_221_799_0, i_10_221_955_0, i_10_221_956_0,
    i_10_221_1032_0, i_10_221_1033_0, i_10_221_1034_0, i_10_221_1234_0,
    i_10_221_1235_0, i_10_221_1240_0, i_10_221_1248_0, i_10_221_1305_0,
    i_10_221_1312_0, i_10_221_1432_0, i_10_221_1438_0, i_10_221_1442_0,
    i_10_221_1577_0, i_10_221_1579_0, i_10_221_1647_0, i_10_221_1648_0,
    i_10_221_1650_0, i_10_221_1651_0, i_10_221_1652_0, i_10_221_1687_0,
    i_10_221_1688_0, i_10_221_1689_0, i_10_221_1822_0, i_10_221_1996_0,
    i_10_221_2001_0, i_10_221_2022_0, i_10_221_2025_0, i_10_221_2230_0,
    i_10_221_2324_0, i_10_221_2358_0, i_10_221_2359_0, i_10_221_2361_0,
    i_10_221_2365_0, i_10_221_2455_0, i_10_221_2471_0, i_10_221_2473_0,
    i_10_221_2474_0, i_10_221_2631_0, i_10_221_2655_0, i_10_221_2657_0,
    i_10_221_2661_0, i_10_221_2701_0, i_10_221_2703_0, i_10_221_2713_0,
    i_10_221_2724_0, i_10_221_2923_0, i_10_221_3033_0, i_10_221_3070_0,
    i_10_221_3196_0, i_10_221_3202_0, i_10_221_3203_0, i_10_221_3277_0,
    i_10_221_3279_0, i_10_221_3384_0, i_10_221_3386_0, i_10_221_3391_0,
    i_10_221_3405_0, i_10_221_3406_0, i_10_221_3609_0, i_10_221_3616_0,
    i_10_221_3717_0, i_10_221_3780_0, i_10_221_3782_0, i_10_221_3783_0,
    i_10_221_3785_0, i_10_221_3786_0, i_10_221_3787_0, i_10_221_3808_0,
    i_10_221_3811_0, i_10_221_3839_0, i_10_221_3844_0, i_10_221_3845_0,
    i_10_221_3847_0, i_10_221_3860_0, i_10_221_4114_0, i_10_221_4273_0,
    i_10_221_4278_0, i_10_221_4285_0, i_10_221_4289_0, i_10_221_4291_0,
    o_10_221_0_0  );
  input  i_10_221_34_0, i_10_221_172_0, i_10_221_224_0, i_10_221_247_0,
    i_10_221_259_0, i_10_221_280_0, i_10_221_283_0, i_10_221_319_0,
    i_10_221_409_0, i_10_221_410_0, i_10_221_447_0, i_10_221_448_0,
    i_10_221_466_0, i_10_221_749_0, i_10_221_752_0, i_10_221_792_0,
    i_10_221_795_0, i_10_221_799_0, i_10_221_955_0, i_10_221_956_0,
    i_10_221_1032_0, i_10_221_1033_0, i_10_221_1034_0, i_10_221_1234_0,
    i_10_221_1235_0, i_10_221_1240_0, i_10_221_1248_0, i_10_221_1305_0,
    i_10_221_1312_0, i_10_221_1432_0, i_10_221_1438_0, i_10_221_1442_0,
    i_10_221_1577_0, i_10_221_1579_0, i_10_221_1647_0, i_10_221_1648_0,
    i_10_221_1650_0, i_10_221_1651_0, i_10_221_1652_0, i_10_221_1687_0,
    i_10_221_1688_0, i_10_221_1689_0, i_10_221_1822_0, i_10_221_1996_0,
    i_10_221_2001_0, i_10_221_2022_0, i_10_221_2025_0, i_10_221_2230_0,
    i_10_221_2324_0, i_10_221_2358_0, i_10_221_2359_0, i_10_221_2361_0,
    i_10_221_2365_0, i_10_221_2455_0, i_10_221_2471_0, i_10_221_2473_0,
    i_10_221_2474_0, i_10_221_2631_0, i_10_221_2655_0, i_10_221_2657_0,
    i_10_221_2661_0, i_10_221_2701_0, i_10_221_2703_0, i_10_221_2713_0,
    i_10_221_2724_0, i_10_221_2923_0, i_10_221_3033_0, i_10_221_3070_0,
    i_10_221_3196_0, i_10_221_3202_0, i_10_221_3203_0, i_10_221_3277_0,
    i_10_221_3279_0, i_10_221_3384_0, i_10_221_3386_0, i_10_221_3391_0,
    i_10_221_3405_0, i_10_221_3406_0, i_10_221_3609_0, i_10_221_3616_0,
    i_10_221_3717_0, i_10_221_3780_0, i_10_221_3782_0, i_10_221_3783_0,
    i_10_221_3785_0, i_10_221_3786_0, i_10_221_3787_0, i_10_221_3808_0,
    i_10_221_3811_0, i_10_221_3839_0, i_10_221_3844_0, i_10_221_3845_0,
    i_10_221_3847_0, i_10_221_3860_0, i_10_221_4114_0, i_10_221_4273_0,
    i_10_221_4278_0, i_10_221_4285_0, i_10_221_4289_0, i_10_221_4291_0;
  output o_10_221_0_0;
  assign o_10_221_0_0 = 0;
endmodule



// Benchmark "kernel_10_222" written by ABC on Sun Jul 19 10:24:50 2020

module kernel_10_222 ( 
    i_10_222_218_0, i_10_222_219_0, i_10_222_220_0, i_10_222_221_0,
    i_10_222_279_0, i_10_222_280_0, i_10_222_391_0, i_10_222_424_0,
    i_10_222_425_0, i_10_222_431_0, i_10_222_460_0, i_10_222_461_0,
    i_10_222_462_0, i_10_222_463_0, i_10_222_464_0, i_10_222_712_0,
    i_10_222_713_0, i_10_222_794_0, i_10_222_899_0, i_10_222_990_0,
    i_10_222_999_0, i_10_222_1236_0, i_10_222_1237_0, i_10_222_1243_0,
    i_10_222_1244_0, i_10_222_1247_0, i_10_222_1250_0, i_10_222_1310_0,
    i_10_222_1365_0, i_10_222_1650_0, i_10_222_1652_0, i_10_222_1686_0,
    i_10_222_1688_0, i_10_222_1821_0, i_10_222_1824_0, i_10_222_1825_0,
    i_10_222_1915_0, i_10_222_2022_0, i_10_222_2180_0, i_10_222_2306_0,
    i_10_222_2350_0, i_10_222_2352_0, i_10_222_2353_0, i_10_222_2354_0,
    i_10_222_2359_0, i_10_222_2452_0, i_10_222_2454_0, i_10_222_2455_0,
    i_10_222_2464_0, i_10_222_2468_0, i_10_222_2471_0, i_10_222_2571_0,
    i_10_222_2628_0, i_10_222_2654_0, i_10_222_2660_0, i_10_222_2700_0,
    i_10_222_2701_0, i_10_222_2702_0, i_10_222_2723_0, i_10_222_2726_0,
    i_10_222_2734_0, i_10_222_2880_0, i_10_222_2887_0, i_10_222_2923_0,
    i_10_222_3037_0, i_10_222_3049_0, i_10_222_3050_0, i_10_222_3073_0,
    i_10_222_3165_0, i_10_222_3196_0, i_10_222_3200_0, i_10_222_3271_0,
    i_10_222_3387_0, i_10_222_3406_0, i_10_222_3408_0, i_10_222_3409_0,
    i_10_222_3613_0, i_10_222_3614_0, i_10_222_3645_0, i_10_222_3653_0,
    i_10_222_3732_0, i_10_222_3783_0, i_10_222_3784_0, i_10_222_3785_0,
    i_10_222_3837_0, i_10_222_3848_0, i_10_222_3854_0, i_10_222_3855_0,
    i_10_222_3856_0, i_10_222_3857_0, i_10_222_3991_0, i_10_222_4119_0,
    i_10_222_4120_0, i_10_222_4121_0, i_10_222_4270_0, i_10_222_4288_0,
    i_10_222_4289_0, i_10_222_4564_0, i_10_222_4565_0, i_10_222_4568_0,
    o_10_222_0_0  );
  input  i_10_222_218_0, i_10_222_219_0, i_10_222_220_0, i_10_222_221_0,
    i_10_222_279_0, i_10_222_280_0, i_10_222_391_0, i_10_222_424_0,
    i_10_222_425_0, i_10_222_431_0, i_10_222_460_0, i_10_222_461_0,
    i_10_222_462_0, i_10_222_463_0, i_10_222_464_0, i_10_222_712_0,
    i_10_222_713_0, i_10_222_794_0, i_10_222_899_0, i_10_222_990_0,
    i_10_222_999_0, i_10_222_1236_0, i_10_222_1237_0, i_10_222_1243_0,
    i_10_222_1244_0, i_10_222_1247_0, i_10_222_1250_0, i_10_222_1310_0,
    i_10_222_1365_0, i_10_222_1650_0, i_10_222_1652_0, i_10_222_1686_0,
    i_10_222_1688_0, i_10_222_1821_0, i_10_222_1824_0, i_10_222_1825_0,
    i_10_222_1915_0, i_10_222_2022_0, i_10_222_2180_0, i_10_222_2306_0,
    i_10_222_2350_0, i_10_222_2352_0, i_10_222_2353_0, i_10_222_2354_0,
    i_10_222_2359_0, i_10_222_2452_0, i_10_222_2454_0, i_10_222_2455_0,
    i_10_222_2464_0, i_10_222_2468_0, i_10_222_2471_0, i_10_222_2571_0,
    i_10_222_2628_0, i_10_222_2654_0, i_10_222_2660_0, i_10_222_2700_0,
    i_10_222_2701_0, i_10_222_2702_0, i_10_222_2723_0, i_10_222_2726_0,
    i_10_222_2734_0, i_10_222_2880_0, i_10_222_2887_0, i_10_222_2923_0,
    i_10_222_3037_0, i_10_222_3049_0, i_10_222_3050_0, i_10_222_3073_0,
    i_10_222_3165_0, i_10_222_3196_0, i_10_222_3200_0, i_10_222_3271_0,
    i_10_222_3387_0, i_10_222_3406_0, i_10_222_3408_0, i_10_222_3409_0,
    i_10_222_3613_0, i_10_222_3614_0, i_10_222_3645_0, i_10_222_3653_0,
    i_10_222_3732_0, i_10_222_3783_0, i_10_222_3784_0, i_10_222_3785_0,
    i_10_222_3837_0, i_10_222_3848_0, i_10_222_3854_0, i_10_222_3855_0,
    i_10_222_3856_0, i_10_222_3857_0, i_10_222_3991_0, i_10_222_4119_0,
    i_10_222_4120_0, i_10_222_4121_0, i_10_222_4270_0, i_10_222_4288_0,
    i_10_222_4289_0, i_10_222_4564_0, i_10_222_4565_0, i_10_222_4568_0;
  output o_10_222_0_0;
  assign o_10_222_0_0 = ~((~i_10_222_3857_0 & ((~i_10_222_218_0 & ~i_10_222_3049_0 & ((~i_10_222_712_0 & ~i_10_222_1243_0 & ~i_10_222_1365_0 & ~i_10_222_2571_0 & ~i_10_222_3196_0 & ~i_10_222_3387_0 & ~i_10_222_3614_0) | (~i_10_222_1688_0 & ~i_10_222_2306_0 & ~i_10_222_3856_0))) | (~i_10_222_431_0 & ((~i_10_222_2452_0 & ~i_10_222_2723_0 & ~i_10_222_2734_0 & ~i_10_222_3406_0 & ~i_10_222_3614_0 & ~i_10_222_3645_0 & ~i_10_222_3854_0) | (~i_10_222_713_0 & i_10_222_2350_0 & ~i_10_222_3856_0))) | (~i_10_222_464_0 & ((i_10_222_1237_0 & i_10_222_1825_0 & ~i_10_222_2628_0 & i_10_222_3613_0) | (~i_10_222_460_0 & ~i_10_222_1247_0 & ~i_10_222_1365_0 & ~i_10_222_1650_0 & ~i_10_222_2354_0 & ~i_10_222_2880_0 & ~i_10_222_3645_0))) | (~i_10_222_219_0 & ~i_10_222_899_0 & ~i_10_222_1247_0 & ~i_10_222_1250_0 & i_10_222_2452_0 & ~i_10_222_3784_0 & ~i_10_222_3856_0))) | (~i_10_222_218_0 & ((i_10_222_279_0 & ~i_10_222_1250_0 & ~i_10_222_1650_0 & ~i_10_222_2354_0 & ~i_10_222_2468_0 & ~i_10_222_3037_0 & ~i_10_222_3785_0) | (~i_10_222_2180_0 & i_10_222_4119_0 & i_10_222_4564_0))) | (~i_10_222_463_0 & ((~i_10_222_2571_0 & ((~i_10_222_794_0 & ((~i_10_222_460_0 & ~i_10_222_1310_0 & ~i_10_222_1688_0 & ~i_10_222_3050_0 & ~i_10_222_3408_0) | (~i_10_222_899_0 & ~i_10_222_3613_0 & ~i_10_222_3645_0 & i_10_222_3784_0 & ~i_10_222_3837_0))) | (~i_10_222_221_0 & ~i_10_222_899_0 & ~i_10_222_1824_0 & ~i_10_222_2468_0 & ~i_10_222_3856_0))) | (~i_10_222_2359_0 & ~i_10_222_2923_0 & ~i_10_222_3037_0 & ~i_10_222_3050_0 & ~i_10_222_3196_0 & ~i_10_222_3271_0 & ~i_10_222_3408_0 & ~i_10_222_3783_0) | (i_10_222_1825_0 & i_10_222_3837_0 & ~i_10_222_3855_0))) | (~i_10_222_460_0 & ((~i_10_222_899_0 & ~i_10_222_1237_0 & ~i_10_222_1686_0 & ~i_10_222_1688_0 & ~i_10_222_3049_0 & ~i_10_222_3406_0 & ~i_10_222_3614_0 & ~i_10_222_3653_0) | (~i_10_222_462_0 & ~i_10_222_464_0 & ~i_10_222_1824_0 & ~i_10_222_2660_0 & ~i_10_222_2923_0 & ~i_10_222_3050_0 & ~i_10_222_3785_0))) | (~i_10_222_464_0 & ((~i_10_222_1824_0 & i_10_222_2455_0 & ~i_10_222_3200_0 & ~i_10_222_3645_0 & ~i_10_222_3732_0) | (~i_10_222_461_0 & i_10_222_2350_0 & ~i_10_222_2471_0 & ~i_10_222_3785_0))) | (~i_10_222_712_0 & ((~i_10_222_461_0 & ((~i_10_222_1365_0 & i_10_222_1824_0 & i_10_222_1825_0 & ~i_10_222_2180_0 & ~i_10_222_2464_0 & ~i_10_222_3837_0) | (~i_10_222_221_0 & ~i_10_222_1824_0 & ~i_10_222_2352_0 & ~i_10_222_3049_0 & ~i_10_222_3785_0 & i_10_222_4288_0))) | (~i_10_222_3049_0 & ~i_10_222_3855_0 & i_10_222_4565_0))) | (~i_10_222_221_0 & ((~i_10_222_1310_0 & ((~i_10_222_999_0 & ~i_10_222_3785_0 & i_10_222_4270_0) | (~i_10_222_220_0 & ~i_10_222_1237_0 & ~i_10_222_1365_0 & ~i_10_222_1650_0 & ~i_10_222_1652_0 & ~i_10_222_2352_0 & ~i_10_222_3614_0 & ~i_10_222_4270_0))) | (i_10_222_1688_0 & ~i_10_222_2352_0 & ~i_10_222_2468_0 & ~i_10_222_2726_0 & ~i_10_222_3049_0 & ~i_10_222_3271_0 & i_10_222_3613_0))) | (~i_10_222_1365_0 & ((~i_10_222_425_0 & ~i_10_222_1244_0 & ~i_10_222_2455_0 & ~i_10_222_3196_0 & ~i_10_222_3200_0 & i_10_222_3613_0 & i_10_222_3653_0) | (i_10_222_2352_0 & ~i_10_222_2726_0 & ~i_10_222_3614_0 & ~i_10_222_3837_0 & i_10_222_4120_0))) | (i_10_222_2350_0 & ((i_10_222_2702_0 & i_10_222_3613_0) | (~i_10_222_3614_0 & ~i_10_222_3645_0 & i_10_222_4289_0))) | (~i_10_222_2452_0 & ~i_10_222_2471_0 & ((i_10_222_1237_0 & ~i_10_222_3200_0 & ~i_10_222_3856_0) | (~i_10_222_2734_0 & i_10_222_4270_0))) | (i_10_222_2701_0 & ~i_10_222_3037_0 & i_10_222_3613_0 & ~i_10_222_3855_0));
endmodule



// Benchmark "kernel_10_223" written by ABC on Sun Jul 19 10:24:52 2020

module kernel_10_223 ( 
    i_10_223_174_0, i_10_223_175_0, i_10_223_216_0, i_10_223_268_0,
    i_10_223_279_0, i_10_223_287_0, i_10_223_443_0, i_10_223_466_0,
    i_10_223_508_0, i_10_223_511_0, i_10_223_697_0, i_10_223_797_0,
    i_10_223_798_0, i_10_223_1005_0, i_10_223_1006_0, i_10_223_1234_0,
    i_10_223_1237_0, i_10_223_1240_0, i_10_223_1249_0, i_10_223_1310_0,
    i_10_223_1311_0, i_10_223_1647_0, i_10_223_1648_0, i_10_223_1650_0,
    i_10_223_1651_0, i_10_223_1652_0, i_10_223_1654_0, i_10_223_1684_0,
    i_10_223_1686_0, i_10_223_1820_0, i_10_223_1821_0, i_10_223_1823_0,
    i_10_223_1824_0, i_10_223_1825_0, i_10_223_1910_0, i_10_223_1913_0,
    i_10_223_1952_0, i_10_223_1994_0, i_10_223_1996_0, i_10_223_2179_0,
    i_10_223_2185_0, i_10_223_2203_0, i_10_223_2332_0, i_10_223_2337_0,
    i_10_223_2338_0, i_10_223_2339_0, i_10_223_2353_0, i_10_223_2366_0,
    i_10_223_2377_0, i_10_223_2380_0, i_10_223_2383_0, i_10_223_2384_0,
    i_10_223_2407_0, i_10_223_2408_0, i_10_223_2410_0, i_10_223_2451_0,
    i_10_223_2456_0, i_10_223_2569_0, i_10_223_2571_0, i_10_223_2572_0,
    i_10_223_2711_0, i_10_223_2730_0, i_10_223_2735_0, i_10_223_2883_0,
    i_10_223_3034_0, i_10_223_3037_0, i_10_223_3046_0, i_10_223_3047_0,
    i_10_223_3048_0, i_10_223_3049_0, i_10_223_3050_0, i_10_223_3069_0,
    i_10_223_3072_0, i_10_223_3074_0, i_10_223_3151_0, i_10_223_3153_0,
    i_10_223_3155_0, i_10_223_3158_0, i_10_223_3199_0, i_10_223_3267_0,
    i_10_223_3268_0, i_10_223_3271_0, i_10_223_3327_0, i_10_223_3405_0,
    i_10_223_3469_0, i_10_223_3497_0, i_10_223_3617_0, i_10_223_3650_0,
    i_10_223_3837_0, i_10_223_3838_0, i_10_223_3839_0, i_10_223_3846_0,
    i_10_223_3847_0, i_10_223_4056_0, i_10_223_4117_0, i_10_223_4118_0,
    i_10_223_4119_0, i_10_223_4120_0, i_10_223_4121_0, i_10_223_4285_0,
    o_10_223_0_0  );
  input  i_10_223_174_0, i_10_223_175_0, i_10_223_216_0, i_10_223_268_0,
    i_10_223_279_0, i_10_223_287_0, i_10_223_443_0, i_10_223_466_0,
    i_10_223_508_0, i_10_223_511_0, i_10_223_697_0, i_10_223_797_0,
    i_10_223_798_0, i_10_223_1005_0, i_10_223_1006_0, i_10_223_1234_0,
    i_10_223_1237_0, i_10_223_1240_0, i_10_223_1249_0, i_10_223_1310_0,
    i_10_223_1311_0, i_10_223_1647_0, i_10_223_1648_0, i_10_223_1650_0,
    i_10_223_1651_0, i_10_223_1652_0, i_10_223_1654_0, i_10_223_1684_0,
    i_10_223_1686_0, i_10_223_1820_0, i_10_223_1821_0, i_10_223_1823_0,
    i_10_223_1824_0, i_10_223_1825_0, i_10_223_1910_0, i_10_223_1913_0,
    i_10_223_1952_0, i_10_223_1994_0, i_10_223_1996_0, i_10_223_2179_0,
    i_10_223_2185_0, i_10_223_2203_0, i_10_223_2332_0, i_10_223_2337_0,
    i_10_223_2338_0, i_10_223_2339_0, i_10_223_2353_0, i_10_223_2366_0,
    i_10_223_2377_0, i_10_223_2380_0, i_10_223_2383_0, i_10_223_2384_0,
    i_10_223_2407_0, i_10_223_2408_0, i_10_223_2410_0, i_10_223_2451_0,
    i_10_223_2456_0, i_10_223_2569_0, i_10_223_2571_0, i_10_223_2572_0,
    i_10_223_2711_0, i_10_223_2730_0, i_10_223_2735_0, i_10_223_2883_0,
    i_10_223_3034_0, i_10_223_3037_0, i_10_223_3046_0, i_10_223_3047_0,
    i_10_223_3048_0, i_10_223_3049_0, i_10_223_3050_0, i_10_223_3069_0,
    i_10_223_3072_0, i_10_223_3074_0, i_10_223_3151_0, i_10_223_3153_0,
    i_10_223_3155_0, i_10_223_3158_0, i_10_223_3199_0, i_10_223_3267_0,
    i_10_223_3268_0, i_10_223_3271_0, i_10_223_3327_0, i_10_223_3405_0,
    i_10_223_3469_0, i_10_223_3497_0, i_10_223_3617_0, i_10_223_3650_0,
    i_10_223_3837_0, i_10_223_3838_0, i_10_223_3839_0, i_10_223_3846_0,
    i_10_223_3847_0, i_10_223_4056_0, i_10_223_4117_0, i_10_223_4118_0,
    i_10_223_4119_0, i_10_223_4120_0, i_10_223_4121_0, i_10_223_4285_0;
  output o_10_223_0_0;
  assign o_10_223_0_0 = ~((i_10_223_174_0 & ((~i_10_223_268_0 & ~i_10_223_1310_0 & ~i_10_223_1654_0 & ~i_10_223_2384_0 & ~i_10_223_3267_0 & ~i_10_223_3271_0 & ~i_10_223_3405_0) | (~i_10_223_1821_0 & ~i_10_223_3049_0 & ~i_10_223_3838_0))) | (~i_10_223_174_0 & ((~i_10_223_216_0 & ~i_10_223_268_0 & ~i_10_223_2337_0 & ~i_10_223_2377_0 & ~i_10_223_2380_0 & i_10_223_3037_0 & ~i_10_223_3046_0) | (i_10_223_1654_0 & i_10_223_1823_0 & ~i_10_223_2383_0 & ~i_10_223_2408_0 & ~i_10_223_2735_0 & ~i_10_223_3846_0))) | (i_10_223_279_0 & ((~i_10_223_443_0 & ~i_10_223_797_0 & ~i_10_223_798_0 & ~i_10_223_2451_0 & ~i_10_223_3049_0 & ~i_10_223_3069_0) | (~i_10_223_2332_0 & ~i_10_223_2572_0 & i_10_223_4120_0))) | (i_10_223_287_0 & ((~i_10_223_268_0 & ~i_10_223_279_0 & ~i_10_223_1913_0 & ~i_10_223_2339_0 & ~i_10_223_2383_0 & ~i_10_223_2735_0 & ~i_10_223_3199_0 & ~i_10_223_3497_0 & ~i_10_223_4056_0) | (i_10_223_2353_0 & ~i_10_223_2408_0 & i_10_223_4121_0))) | (~i_10_223_3267_0 & ((~i_10_223_2366_0 & ((~i_10_223_268_0 & ~i_10_223_3069_0 & ((~i_10_223_1647_0 & i_10_223_1824_0 & ~i_10_223_1952_0 & ~i_10_223_2571_0 & ~i_10_223_2572_0 & ~i_10_223_2883_0) | (~i_10_223_798_0 & ~i_10_223_1650_0 & ~i_10_223_2185_0 & ~i_10_223_2332_0 & ~i_10_223_2384_0 & ~i_10_223_3838_0))) | (~i_10_223_2339_0 & ((i_10_223_466_0 & ~i_10_223_1005_0 & ~i_10_223_1821_0 & ~i_10_223_1913_0 & ~i_10_223_2408_0 & ~i_10_223_3047_0) | (~i_10_223_443_0 & ~i_10_223_1310_0 & ~i_10_223_1650_0 & ~i_10_223_1994_0 & ~i_10_223_2179_0 & ~i_10_223_3048_0 & ~i_10_223_3049_0 & ~i_10_223_3271_0))))) | (i_10_223_3847_0 & i_10_223_4117_0) | (~i_10_223_1996_0 & ~i_10_223_3047_0 & ~i_10_223_3268_0 & i_10_223_4120_0))) | (~i_10_223_2407_0 & ((~i_10_223_1005_0 & ((~i_10_223_797_0 & ~i_10_223_1006_0 & ~i_10_223_1311_0 & ~i_10_223_1684_0 & ~i_10_223_1821_0 & ~i_10_223_1996_0 & ~i_10_223_2456_0 & ~i_10_223_2571_0 & ~i_10_223_2711_0 & ~i_10_223_3069_0) | (~i_10_223_1651_0 & ~i_10_223_3072_0 & ~i_10_223_3271_0 & i_10_223_3846_0))) | (~i_10_223_2179_0 & ~i_10_223_3271_0 & ((~i_10_223_216_0 & ~i_10_223_1647_0 & ~i_10_223_1825_0 & ~i_10_223_3048_0 & ~i_10_223_3050_0 & ~i_10_223_3268_0 & i_10_223_3837_0) | (~i_10_223_3405_0 & ~i_10_223_3837_0 & i_10_223_4117_0))) | (~i_10_223_1006_0 & ~i_10_223_1240_0 & ~i_10_223_1651_0 & ~i_10_223_2353_0 & ~i_10_223_2380_0 & ~i_10_223_2384_0 & ~i_10_223_3074_0))) | (~i_10_223_2332_0 & ((~i_10_223_216_0 & ((~i_10_223_1647_0 & ~i_10_223_2179_0 & ~i_10_223_2339_0 & ~i_10_223_2571_0 & i_10_223_3847_0) | (i_10_223_1820_0 & ~i_10_223_2569_0 & ~i_10_223_2572_0 & ~i_10_223_3838_0 & ~i_10_223_4056_0))) | (i_10_223_1652_0 & ~i_10_223_1821_0 & ~i_10_223_2456_0 & i_10_223_4117_0))) | (~i_10_223_1006_0 & ((~i_10_223_1648_0 & ~i_10_223_1996_0 & ~i_10_223_2179_0 & ~i_10_223_2366_0 & ~i_10_223_2384_0 & ~i_10_223_2408_0 & ~i_10_223_2571_0 & ~i_10_223_3047_0 & ~i_10_223_3271_0 & ~i_10_223_3837_0) | (~i_10_223_466_0 & i_10_223_1311_0 & ~i_10_223_3405_0 & i_10_223_3838_0))) | (~i_10_223_1647_0 & ((~i_10_223_2179_0 & ((~i_10_223_1952_0 & ~i_10_223_3037_0 & i_10_223_3650_0 & ~i_10_223_3838_0) | (~i_10_223_2185_0 & ~i_10_223_2572_0 & i_10_223_4118_0))) | (~i_10_223_1654_0 & i_10_223_1684_0 & ~i_10_223_3047_0 & ~i_10_223_3837_0 & ~i_10_223_3839_0) | (~i_10_223_3050_0 & i_10_223_4119_0))) | (~i_10_223_2185_0 & ((~i_10_223_1650_0 & ~i_10_223_1652_0 & ~i_10_223_1684_0 & ~i_10_223_1994_0 & ~i_10_223_2203_0 & ~i_10_223_3049_0 & ~i_10_223_3050_0 & ~i_10_223_3497_0 & ~i_10_223_3847_0) | (~i_10_223_2377_0 & ~i_10_223_3048_0 & ~i_10_223_3839_0 & i_10_223_4119_0))) | (~i_10_223_3199_0 & ((~i_10_223_3271_0 & ~i_10_223_4056_0 & i_10_223_4120_0) | (i_10_223_797_0 & ~i_10_223_1996_0 & ~i_10_223_2377_0 & ~i_10_223_2410_0 & ~i_10_223_2730_0 & ~i_10_223_3049_0 & ~i_10_223_3837_0 & ~i_10_223_4121_0))) | (i_10_223_2730_0 & (i_10_223_697_0 | (~i_10_223_3049_0 & ((~i_10_223_798_0 & ~i_10_223_1821_0 & i_10_223_2410_0) | (~i_10_223_2380_0 & i_10_223_4117_0))))) | (~i_10_223_3839_0 & ((i_10_223_1237_0 & ~i_10_223_1240_0 & i_10_223_1913_0 & i_10_223_2451_0 & ~i_10_223_3650_0 & ~i_10_223_3838_0) | (i_10_223_1821_0 & ~i_10_223_3072_0 & ~i_10_223_3268_0 & i_10_223_4117_0))) | (i_10_223_1651_0 & ~i_10_223_1823_0 & i_10_223_2380_0 & ~i_10_223_2384_0 & i_10_223_3034_0) | (i_10_223_1820_0 & i_10_223_3074_0 & i_10_223_3650_0 & ~i_10_223_3837_0) | (~i_10_223_1686_0 & ~i_10_223_3405_0 & i_10_223_3839_0 & i_10_223_4117_0));
endmodule



// Benchmark "kernel_10_224" written by ABC on Sun Jul 19 10:24:52 2020

module kernel_10_224 ( 
    i_10_224_29_0, i_10_224_216_0, i_10_224_283_0, i_10_224_284_0,
    i_10_224_308_0, i_10_224_374_0, i_10_224_433_0, i_10_224_444_0,
    i_10_224_505_0, i_10_224_558_0, i_10_224_623_0, i_10_224_794_0,
    i_10_224_821_0, i_10_224_847_0, i_10_224_893_0, i_10_224_895_0,
    i_10_224_901_0, i_10_224_1030_0, i_10_224_1031_0, i_10_224_1084_0,
    i_10_224_1085_0, i_10_224_1233_0, i_10_224_1235_0, i_10_224_1243_0,
    i_10_224_1548_0, i_10_224_1575_0, i_10_224_1606_0, i_10_224_1612_0,
    i_10_224_1616_0, i_10_224_1684_0, i_10_224_1825_0, i_10_224_1911_0,
    i_10_224_1956_0, i_10_224_1990_0, i_10_224_1991_0, i_10_224_2090_0,
    i_10_224_2225_0, i_10_224_2242_0, i_10_224_2304_0, i_10_224_2332_0,
    i_10_224_2335_0, i_10_224_2336_0, i_10_224_2361_0, i_10_224_2462_0,
    i_10_224_2556_0, i_10_224_2567_0, i_10_224_2632_0, i_10_224_2638_0,
    i_10_224_2639_0, i_10_224_2660_0, i_10_224_2675_0, i_10_224_2701_0,
    i_10_224_2702_0, i_10_224_2709_0, i_10_224_2728_0, i_10_224_2729_0,
    i_10_224_2783_0, i_10_224_2827_0, i_10_224_2829_0, i_10_224_2830_0,
    i_10_224_2867_0, i_10_224_2880_0, i_10_224_2917_0, i_10_224_2920_0,
    i_10_224_3160_0, i_10_224_3161_0, i_10_224_3315_0, i_10_224_3353_0,
    i_10_224_3385_0, i_10_224_3389_0, i_10_224_3440_0, i_10_224_3448_0,
    i_10_224_3457_0, i_10_224_3458_0, i_10_224_3551_0, i_10_224_3553_0,
    i_10_224_3557_0, i_10_224_3611_0, i_10_224_3614_0, i_10_224_3646_0,
    i_10_224_3784_0, i_10_224_3834_0, i_10_224_3837_0, i_10_224_3848_0,
    i_10_224_3856_0, i_10_224_3857_0, i_10_224_3880_0, i_10_224_3920_0,
    i_10_224_3978_0, i_10_224_4009_0, i_10_224_4010_0, i_10_224_4028_0,
    i_10_224_4051_0, i_10_224_4052_0, i_10_224_4213_0, i_10_224_4214_0,
    i_10_224_4291_0, i_10_224_4302_0, i_10_224_4564_0, i_10_224_4565_0,
    o_10_224_0_0  );
  input  i_10_224_29_0, i_10_224_216_0, i_10_224_283_0, i_10_224_284_0,
    i_10_224_308_0, i_10_224_374_0, i_10_224_433_0, i_10_224_444_0,
    i_10_224_505_0, i_10_224_558_0, i_10_224_623_0, i_10_224_794_0,
    i_10_224_821_0, i_10_224_847_0, i_10_224_893_0, i_10_224_895_0,
    i_10_224_901_0, i_10_224_1030_0, i_10_224_1031_0, i_10_224_1084_0,
    i_10_224_1085_0, i_10_224_1233_0, i_10_224_1235_0, i_10_224_1243_0,
    i_10_224_1548_0, i_10_224_1575_0, i_10_224_1606_0, i_10_224_1612_0,
    i_10_224_1616_0, i_10_224_1684_0, i_10_224_1825_0, i_10_224_1911_0,
    i_10_224_1956_0, i_10_224_1990_0, i_10_224_1991_0, i_10_224_2090_0,
    i_10_224_2225_0, i_10_224_2242_0, i_10_224_2304_0, i_10_224_2332_0,
    i_10_224_2335_0, i_10_224_2336_0, i_10_224_2361_0, i_10_224_2462_0,
    i_10_224_2556_0, i_10_224_2567_0, i_10_224_2632_0, i_10_224_2638_0,
    i_10_224_2639_0, i_10_224_2660_0, i_10_224_2675_0, i_10_224_2701_0,
    i_10_224_2702_0, i_10_224_2709_0, i_10_224_2728_0, i_10_224_2729_0,
    i_10_224_2783_0, i_10_224_2827_0, i_10_224_2829_0, i_10_224_2830_0,
    i_10_224_2867_0, i_10_224_2880_0, i_10_224_2917_0, i_10_224_2920_0,
    i_10_224_3160_0, i_10_224_3161_0, i_10_224_3315_0, i_10_224_3353_0,
    i_10_224_3385_0, i_10_224_3389_0, i_10_224_3440_0, i_10_224_3448_0,
    i_10_224_3457_0, i_10_224_3458_0, i_10_224_3551_0, i_10_224_3553_0,
    i_10_224_3557_0, i_10_224_3611_0, i_10_224_3614_0, i_10_224_3646_0,
    i_10_224_3784_0, i_10_224_3834_0, i_10_224_3837_0, i_10_224_3848_0,
    i_10_224_3856_0, i_10_224_3857_0, i_10_224_3880_0, i_10_224_3920_0,
    i_10_224_3978_0, i_10_224_4009_0, i_10_224_4010_0, i_10_224_4028_0,
    i_10_224_4051_0, i_10_224_4052_0, i_10_224_4213_0, i_10_224_4214_0,
    i_10_224_4291_0, i_10_224_4302_0, i_10_224_4564_0, i_10_224_4565_0;
  output o_10_224_0_0;
  assign o_10_224_0_0 = 0;
endmodule



// Benchmark "kernel_10_225" written by ABC on Sun Jul 19 10:24:53 2020

module kernel_10_225 ( 
    i_10_225_171_0, i_10_225_174_0, i_10_225_185_0, i_10_225_217_0,
    i_10_225_218_0, i_10_225_221_0, i_10_225_223_0, i_10_225_255_0,
    i_10_225_271_0, i_10_225_276_0, i_10_225_315_0, i_10_225_370_0,
    i_10_225_395_0, i_10_225_427_0, i_10_225_433_0, i_10_225_436_0,
    i_10_225_460_0, i_10_225_461_0, i_10_225_712_0, i_10_225_904_0,
    i_10_225_1027_0, i_10_225_1084_0, i_10_225_1120_0, i_10_225_1162_0,
    i_10_225_1237_0, i_10_225_1240_0, i_10_225_1242_0, i_10_225_1243_0,
    i_10_225_1246_0, i_10_225_1264_0, i_10_225_1308_0, i_10_225_1542_0,
    i_10_225_1544_0, i_10_225_1583_0, i_10_225_1650_0, i_10_225_1688_0,
    i_10_225_1908_0, i_10_225_1910_0, i_10_225_2304_0, i_10_225_2310_0,
    i_10_225_2312_0, i_10_225_2356_0, i_10_225_2359_0, i_10_225_2363_0,
    i_10_225_2367_0, i_10_225_2452_0, i_10_225_2458_0, i_10_225_2470_0,
    i_10_225_2471_0, i_10_225_2513_0, i_10_225_2713_0, i_10_225_2714_0,
    i_10_225_2721_0, i_10_225_2727_0, i_10_225_2730_0, i_10_225_2831_0,
    i_10_225_2884_0, i_10_225_2923_0, i_10_225_2982_0, i_10_225_3034_0,
    i_10_225_3036_0, i_10_225_3198_0, i_10_225_3199_0, i_10_225_3280_0,
    i_10_225_3297_0, i_10_225_3335_0, i_10_225_3390_0, i_10_225_3402_0,
    i_10_225_3405_0, i_10_225_3406_0, i_10_225_3410_0, i_10_225_3430_0,
    i_10_225_3586_0, i_10_225_3609_0, i_10_225_3612_0, i_10_225_3616_0,
    i_10_225_3652_0, i_10_225_3689_0, i_10_225_3730_0, i_10_225_3731_0,
    i_10_225_3780_0, i_10_225_3783_0, i_10_225_3784_0, i_10_225_3821_0,
    i_10_225_3840_0, i_10_225_3855_0, i_10_225_3858_0, i_10_225_3892_0,
    i_10_225_3943_0, i_10_225_3991_0, i_10_225_3992_0, i_10_225_3998_0,
    i_10_225_4173_0, i_10_225_4174_0, i_10_225_4213_0, i_10_225_4214_0,
    i_10_225_4274_0, i_10_225_4288_0, i_10_225_4289_0, i_10_225_4567_0,
    o_10_225_0_0  );
  input  i_10_225_171_0, i_10_225_174_0, i_10_225_185_0, i_10_225_217_0,
    i_10_225_218_0, i_10_225_221_0, i_10_225_223_0, i_10_225_255_0,
    i_10_225_271_0, i_10_225_276_0, i_10_225_315_0, i_10_225_370_0,
    i_10_225_395_0, i_10_225_427_0, i_10_225_433_0, i_10_225_436_0,
    i_10_225_460_0, i_10_225_461_0, i_10_225_712_0, i_10_225_904_0,
    i_10_225_1027_0, i_10_225_1084_0, i_10_225_1120_0, i_10_225_1162_0,
    i_10_225_1237_0, i_10_225_1240_0, i_10_225_1242_0, i_10_225_1243_0,
    i_10_225_1246_0, i_10_225_1264_0, i_10_225_1308_0, i_10_225_1542_0,
    i_10_225_1544_0, i_10_225_1583_0, i_10_225_1650_0, i_10_225_1688_0,
    i_10_225_1908_0, i_10_225_1910_0, i_10_225_2304_0, i_10_225_2310_0,
    i_10_225_2312_0, i_10_225_2356_0, i_10_225_2359_0, i_10_225_2363_0,
    i_10_225_2367_0, i_10_225_2452_0, i_10_225_2458_0, i_10_225_2470_0,
    i_10_225_2471_0, i_10_225_2513_0, i_10_225_2713_0, i_10_225_2714_0,
    i_10_225_2721_0, i_10_225_2727_0, i_10_225_2730_0, i_10_225_2831_0,
    i_10_225_2884_0, i_10_225_2923_0, i_10_225_2982_0, i_10_225_3034_0,
    i_10_225_3036_0, i_10_225_3198_0, i_10_225_3199_0, i_10_225_3280_0,
    i_10_225_3297_0, i_10_225_3335_0, i_10_225_3390_0, i_10_225_3402_0,
    i_10_225_3405_0, i_10_225_3406_0, i_10_225_3410_0, i_10_225_3430_0,
    i_10_225_3586_0, i_10_225_3609_0, i_10_225_3612_0, i_10_225_3616_0,
    i_10_225_3652_0, i_10_225_3689_0, i_10_225_3730_0, i_10_225_3731_0,
    i_10_225_3780_0, i_10_225_3783_0, i_10_225_3784_0, i_10_225_3821_0,
    i_10_225_3840_0, i_10_225_3855_0, i_10_225_3858_0, i_10_225_3892_0,
    i_10_225_3943_0, i_10_225_3991_0, i_10_225_3992_0, i_10_225_3998_0,
    i_10_225_4173_0, i_10_225_4174_0, i_10_225_4213_0, i_10_225_4214_0,
    i_10_225_4274_0, i_10_225_4288_0, i_10_225_4289_0, i_10_225_4567_0;
  output o_10_225_0_0;
  assign o_10_225_0_0 = 0;
endmodule



// Benchmark "kernel_10_226" written by ABC on Sun Jul 19 10:24:54 2020

module kernel_10_226 ( 
    i_10_226_223_0, i_10_226_269_0, i_10_226_292_0, i_10_226_320_0,
    i_10_226_323_0, i_10_226_432_0, i_10_226_437_0, i_10_226_446_0,
    i_10_226_448_0, i_10_226_462_0, i_10_226_466_0, i_10_226_503_0,
    i_10_226_509_0, i_10_226_628_0, i_10_226_629_0, i_10_226_711_0,
    i_10_226_716_0, i_10_226_799_0, i_10_226_896_0, i_10_226_968_0,
    i_10_226_1011_0, i_10_226_1034_0, i_10_226_1106_0, i_10_226_1124_0,
    i_10_226_1156_0, i_10_226_1223_0, i_10_226_1270_0, i_10_226_1354_0,
    i_10_226_1439_0, i_10_226_1441_0, i_10_226_1442_0, i_10_226_1448_0,
    i_10_226_1492_0, i_10_226_1545_0, i_10_226_1581_0, i_10_226_1582_0,
    i_10_226_1637_0, i_10_226_1689_0, i_10_226_1690_0, i_10_226_1691_0,
    i_10_226_1736_0, i_10_226_1808_0, i_10_226_1822_0, i_10_226_1984_0,
    i_10_226_1994_0, i_10_226_2005_0, i_10_226_2006_0, i_10_226_2033_0,
    i_10_226_2202_0, i_10_226_2223_0, i_10_226_2347_0, i_10_226_2352_0,
    i_10_226_2365_0, i_10_226_2366_0, i_10_226_2451_0, i_10_226_2474_0,
    i_10_226_2635_0, i_10_226_2659_0, i_10_226_2679_0, i_10_226_2680_0,
    i_10_226_2704_0, i_10_226_2715_0, i_10_226_2722_0, i_10_226_2732_0,
    i_10_226_2762_0, i_10_226_2782_0, i_10_226_2833_0, i_10_226_2919_0,
    i_10_226_2924_0, i_10_226_2969_0, i_10_226_2978_0, i_10_226_3077_0,
    i_10_226_3199_0, i_10_226_3281_0, i_10_226_3389_0, i_10_226_3409_0,
    i_10_226_3465_0, i_10_226_3467_0, i_10_226_3473_0, i_10_226_3494_0,
    i_10_226_3497_0, i_10_226_3538_0, i_10_226_3545_0, i_10_226_3587_0,
    i_10_226_3590_0, i_10_226_3649_0, i_10_226_3853_0, i_10_226_3914_0,
    i_10_226_3923_0, i_10_226_4122_0, i_10_226_4210_0, i_10_226_4211_0,
    i_10_226_4269_0, i_10_226_4271_0, i_10_226_4273_0, i_10_226_4281_0,
    i_10_226_4291_0, i_10_226_4395_0, i_10_226_4584_0, i_10_226_4589_0,
    o_10_226_0_0  );
  input  i_10_226_223_0, i_10_226_269_0, i_10_226_292_0, i_10_226_320_0,
    i_10_226_323_0, i_10_226_432_0, i_10_226_437_0, i_10_226_446_0,
    i_10_226_448_0, i_10_226_462_0, i_10_226_466_0, i_10_226_503_0,
    i_10_226_509_0, i_10_226_628_0, i_10_226_629_0, i_10_226_711_0,
    i_10_226_716_0, i_10_226_799_0, i_10_226_896_0, i_10_226_968_0,
    i_10_226_1011_0, i_10_226_1034_0, i_10_226_1106_0, i_10_226_1124_0,
    i_10_226_1156_0, i_10_226_1223_0, i_10_226_1270_0, i_10_226_1354_0,
    i_10_226_1439_0, i_10_226_1441_0, i_10_226_1442_0, i_10_226_1448_0,
    i_10_226_1492_0, i_10_226_1545_0, i_10_226_1581_0, i_10_226_1582_0,
    i_10_226_1637_0, i_10_226_1689_0, i_10_226_1690_0, i_10_226_1691_0,
    i_10_226_1736_0, i_10_226_1808_0, i_10_226_1822_0, i_10_226_1984_0,
    i_10_226_1994_0, i_10_226_2005_0, i_10_226_2006_0, i_10_226_2033_0,
    i_10_226_2202_0, i_10_226_2223_0, i_10_226_2347_0, i_10_226_2352_0,
    i_10_226_2365_0, i_10_226_2366_0, i_10_226_2451_0, i_10_226_2474_0,
    i_10_226_2635_0, i_10_226_2659_0, i_10_226_2679_0, i_10_226_2680_0,
    i_10_226_2704_0, i_10_226_2715_0, i_10_226_2722_0, i_10_226_2732_0,
    i_10_226_2762_0, i_10_226_2782_0, i_10_226_2833_0, i_10_226_2919_0,
    i_10_226_2924_0, i_10_226_2969_0, i_10_226_2978_0, i_10_226_3077_0,
    i_10_226_3199_0, i_10_226_3281_0, i_10_226_3389_0, i_10_226_3409_0,
    i_10_226_3465_0, i_10_226_3467_0, i_10_226_3473_0, i_10_226_3494_0,
    i_10_226_3497_0, i_10_226_3538_0, i_10_226_3545_0, i_10_226_3587_0,
    i_10_226_3590_0, i_10_226_3649_0, i_10_226_3853_0, i_10_226_3914_0,
    i_10_226_3923_0, i_10_226_4122_0, i_10_226_4210_0, i_10_226_4211_0,
    i_10_226_4269_0, i_10_226_4271_0, i_10_226_4273_0, i_10_226_4281_0,
    i_10_226_4291_0, i_10_226_4395_0, i_10_226_4584_0, i_10_226_4589_0;
  output o_10_226_0_0;
  assign o_10_226_0_0 = 0;
endmodule



// Benchmark "kernel_10_227" written by ABC on Sun Jul 19 10:24:55 2020

module kernel_10_227 ( 
    i_10_227_122_0, i_10_227_171_0, i_10_227_174_0, i_10_227_175_0,
    i_10_227_176_0, i_10_227_282_0, i_10_227_283_0, i_10_227_319_0,
    i_10_227_387_0, i_10_227_409_0, i_10_227_434_0, i_10_227_445_0,
    i_10_227_460_0, i_10_227_461_0, i_10_227_462_0, i_10_227_464_0,
    i_10_227_497_0, i_10_227_713_0, i_10_227_752_0, i_10_227_900_0,
    i_10_227_1048_0, i_10_227_1084_0, i_10_227_1237_0, i_10_227_1238_0,
    i_10_227_1279_0, i_10_227_1310_0, i_10_227_1342_0, i_10_227_1354_0,
    i_10_227_1435_0, i_10_227_1539_0, i_10_227_1540_0, i_10_227_1580_0,
    i_10_227_1651_0, i_10_227_1687_0, i_10_227_1688_0, i_10_227_1690_0,
    i_10_227_1691_0, i_10_227_1909_0, i_10_227_2033_0, i_10_227_2201_0,
    i_10_227_2359_0, i_10_227_2379_0, i_10_227_2452_0, i_10_227_2455_0,
    i_10_227_2468_0, i_10_227_2629_0, i_10_227_2630_0, i_10_227_2644_0,
    i_10_227_2656_0, i_10_227_2657_0, i_10_227_2658_0, i_10_227_2659_0,
    i_10_227_2679_0, i_10_227_2711_0, i_10_227_2720_0, i_10_227_2722_0,
    i_10_227_2789_0, i_10_227_2817_0, i_10_227_3070_0, i_10_227_3071_0,
    i_10_227_3200_0, i_10_227_3276_0, i_10_227_3277_0, i_10_227_3278_0,
    i_10_227_3279_0, i_10_227_3280_0, i_10_227_3281_0, i_10_227_3283_0,
    i_10_227_3316_0, i_10_227_3385_0, i_10_227_3387_0, i_10_227_3392_0,
    i_10_227_3496_0, i_10_227_3538_0, i_10_227_3541_0, i_10_227_3587_0,
    i_10_227_3686_0, i_10_227_3837_0, i_10_227_3838_0, i_10_227_3839_0,
    i_10_227_3849_0, i_10_227_3856_0, i_10_227_3857_0, i_10_227_3859_0,
    i_10_227_3860_0, i_10_227_3888_0, i_10_227_3889_0, i_10_227_3981_0,
    i_10_227_3982_0, i_10_227_4114_0, i_10_227_4118_0, i_10_227_4167_0,
    i_10_227_4170_0, i_10_227_4171_0, i_10_227_4269_0, i_10_227_4270_0,
    i_10_227_4287_0, i_10_227_4288_0, i_10_227_4289_0, i_10_227_4290_0,
    o_10_227_0_0  );
  input  i_10_227_122_0, i_10_227_171_0, i_10_227_174_0, i_10_227_175_0,
    i_10_227_176_0, i_10_227_282_0, i_10_227_283_0, i_10_227_319_0,
    i_10_227_387_0, i_10_227_409_0, i_10_227_434_0, i_10_227_445_0,
    i_10_227_460_0, i_10_227_461_0, i_10_227_462_0, i_10_227_464_0,
    i_10_227_497_0, i_10_227_713_0, i_10_227_752_0, i_10_227_900_0,
    i_10_227_1048_0, i_10_227_1084_0, i_10_227_1237_0, i_10_227_1238_0,
    i_10_227_1279_0, i_10_227_1310_0, i_10_227_1342_0, i_10_227_1354_0,
    i_10_227_1435_0, i_10_227_1539_0, i_10_227_1540_0, i_10_227_1580_0,
    i_10_227_1651_0, i_10_227_1687_0, i_10_227_1688_0, i_10_227_1690_0,
    i_10_227_1691_0, i_10_227_1909_0, i_10_227_2033_0, i_10_227_2201_0,
    i_10_227_2359_0, i_10_227_2379_0, i_10_227_2452_0, i_10_227_2455_0,
    i_10_227_2468_0, i_10_227_2629_0, i_10_227_2630_0, i_10_227_2644_0,
    i_10_227_2656_0, i_10_227_2657_0, i_10_227_2658_0, i_10_227_2659_0,
    i_10_227_2679_0, i_10_227_2711_0, i_10_227_2720_0, i_10_227_2722_0,
    i_10_227_2789_0, i_10_227_2817_0, i_10_227_3070_0, i_10_227_3071_0,
    i_10_227_3200_0, i_10_227_3276_0, i_10_227_3277_0, i_10_227_3278_0,
    i_10_227_3279_0, i_10_227_3280_0, i_10_227_3281_0, i_10_227_3283_0,
    i_10_227_3316_0, i_10_227_3385_0, i_10_227_3387_0, i_10_227_3392_0,
    i_10_227_3496_0, i_10_227_3538_0, i_10_227_3541_0, i_10_227_3587_0,
    i_10_227_3686_0, i_10_227_3837_0, i_10_227_3838_0, i_10_227_3839_0,
    i_10_227_3849_0, i_10_227_3856_0, i_10_227_3857_0, i_10_227_3859_0,
    i_10_227_3860_0, i_10_227_3888_0, i_10_227_3889_0, i_10_227_3981_0,
    i_10_227_3982_0, i_10_227_4114_0, i_10_227_4118_0, i_10_227_4167_0,
    i_10_227_4170_0, i_10_227_4171_0, i_10_227_4269_0, i_10_227_4270_0,
    i_10_227_4287_0, i_10_227_4288_0, i_10_227_4289_0, i_10_227_4290_0;
  output o_10_227_0_0;
  assign o_10_227_0_0 = 0;
endmodule



// Benchmark "kernel_10_228" written by ABC on Sun Jul 19 10:24:56 2020

module kernel_10_228 ( 
    i_10_228_38_0, i_10_228_148_0, i_10_228_286_0, i_10_228_287_0,
    i_10_228_356_0, i_10_228_358_0, i_10_228_359_0, i_10_228_365_0,
    i_10_228_374_0, i_10_228_410_0, i_10_228_428_0, i_10_228_446_0,
    i_10_228_464_0, i_10_228_635_0, i_10_228_719_0, i_10_228_734_0,
    i_10_228_736_0, i_10_228_737_0, i_10_228_755_0, i_10_228_793_0,
    i_10_228_800_0, i_10_228_832_0, i_10_228_905_0, i_10_228_955_0,
    i_10_228_959_0, i_10_228_994_0, i_10_228_1054_0, i_10_228_1088_0,
    i_10_228_1136_0, i_10_228_1162_0, i_10_228_1163_0, i_10_228_1166_0,
    i_10_228_1219_0, i_10_228_1235_0, i_10_228_1238_0, i_10_228_1262_0,
    i_10_228_1289_0, i_10_228_1292_0, i_10_228_1349_0, i_10_228_1355_0,
    i_10_228_1493_0, i_10_228_1535_0, i_10_228_1651_0, i_10_228_1652_0,
    i_10_228_1694_0, i_10_228_1823_0, i_10_228_1847_0, i_10_228_1850_0,
    i_10_228_1913_0, i_10_228_1958_0, i_10_228_2003_0, i_10_228_2207_0,
    i_10_228_2213_0, i_10_228_2249_0, i_10_228_2386_0, i_10_228_2387_0,
    i_10_228_2390_0, i_10_228_2408_0, i_10_228_2452_0, i_10_228_2454_0,
    i_10_228_2455_0, i_10_228_2495_0, i_10_228_2519_0, i_10_228_2543_0,
    i_10_228_2609_0, i_10_228_2611_0, i_10_228_2632_0, i_10_228_2633_0,
    i_10_228_2659_0, i_10_228_2678_0, i_10_228_2833_0, i_10_228_2980_0,
    i_10_228_2984_0, i_10_228_3119_0, i_10_228_3278_0, i_10_228_3283_0,
    i_10_228_3292_0, i_10_228_3293_0, i_10_228_3317_0, i_10_228_3326_0,
    i_10_228_3362_0, i_10_228_3385_0, i_10_228_3386_0, i_10_228_3388_0,
    i_10_228_3526_0, i_10_228_3539_0, i_10_228_3581_0, i_10_228_3584_0,
    i_10_228_3616_0, i_10_228_3638_0, i_10_228_3777_0, i_10_228_3824_0,
    i_10_228_4001_0, i_10_228_4061_0, i_10_228_4064_0, i_10_228_4115_0,
    i_10_228_4306_0, i_10_228_4382_0, i_10_228_4484_0, i_10_228_4571_0,
    o_10_228_0_0  );
  input  i_10_228_38_0, i_10_228_148_0, i_10_228_286_0, i_10_228_287_0,
    i_10_228_356_0, i_10_228_358_0, i_10_228_359_0, i_10_228_365_0,
    i_10_228_374_0, i_10_228_410_0, i_10_228_428_0, i_10_228_446_0,
    i_10_228_464_0, i_10_228_635_0, i_10_228_719_0, i_10_228_734_0,
    i_10_228_736_0, i_10_228_737_0, i_10_228_755_0, i_10_228_793_0,
    i_10_228_800_0, i_10_228_832_0, i_10_228_905_0, i_10_228_955_0,
    i_10_228_959_0, i_10_228_994_0, i_10_228_1054_0, i_10_228_1088_0,
    i_10_228_1136_0, i_10_228_1162_0, i_10_228_1163_0, i_10_228_1166_0,
    i_10_228_1219_0, i_10_228_1235_0, i_10_228_1238_0, i_10_228_1262_0,
    i_10_228_1289_0, i_10_228_1292_0, i_10_228_1349_0, i_10_228_1355_0,
    i_10_228_1493_0, i_10_228_1535_0, i_10_228_1651_0, i_10_228_1652_0,
    i_10_228_1694_0, i_10_228_1823_0, i_10_228_1847_0, i_10_228_1850_0,
    i_10_228_1913_0, i_10_228_1958_0, i_10_228_2003_0, i_10_228_2207_0,
    i_10_228_2213_0, i_10_228_2249_0, i_10_228_2386_0, i_10_228_2387_0,
    i_10_228_2390_0, i_10_228_2408_0, i_10_228_2452_0, i_10_228_2454_0,
    i_10_228_2455_0, i_10_228_2495_0, i_10_228_2519_0, i_10_228_2543_0,
    i_10_228_2609_0, i_10_228_2611_0, i_10_228_2632_0, i_10_228_2633_0,
    i_10_228_2659_0, i_10_228_2678_0, i_10_228_2833_0, i_10_228_2980_0,
    i_10_228_2984_0, i_10_228_3119_0, i_10_228_3278_0, i_10_228_3283_0,
    i_10_228_3292_0, i_10_228_3293_0, i_10_228_3317_0, i_10_228_3326_0,
    i_10_228_3362_0, i_10_228_3385_0, i_10_228_3386_0, i_10_228_3388_0,
    i_10_228_3526_0, i_10_228_3539_0, i_10_228_3581_0, i_10_228_3584_0,
    i_10_228_3616_0, i_10_228_3638_0, i_10_228_3777_0, i_10_228_3824_0,
    i_10_228_4001_0, i_10_228_4061_0, i_10_228_4064_0, i_10_228_4115_0,
    i_10_228_4306_0, i_10_228_4382_0, i_10_228_4484_0, i_10_228_4571_0;
  output o_10_228_0_0;
  assign o_10_228_0_0 = 0;
endmodule



// Benchmark "kernel_10_229" written by ABC on Sun Jul 19 10:24:57 2020

module kernel_10_229 ( 
    i_10_229_174_0, i_10_229_175_0, i_10_229_176_0, i_10_229_184_0,
    i_10_229_270_0, i_10_229_286_0, i_10_229_287_0, i_10_229_319_0,
    i_10_229_409_0, i_10_229_410_0, i_10_229_436_0, i_10_229_438_0,
    i_10_229_440_0, i_10_229_446_0, i_10_229_447_0, i_10_229_448_0,
    i_10_229_449_0, i_10_229_466_0, i_10_229_467_0, i_10_229_518_0,
    i_10_229_717_0, i_10_229_718_0, i_10_229_719_0, i_10_229_755_0,
    i_10_229_793_0, i_10_229_797_0, i_10_229_798_0, i_10_229_799_0,
    i_10_229_958_0, i_10_229_968_0, i_10_229_971_0, i_10_229_1003_0,
    i_10_229_1006_0, i_10_229_1164_0, i_10_229_1165_0, i_10_229_1166_0,
    i_10_229_1169_0, i_10_229_1237_0, i_10_229_1245_0, i_10_229_1247_0,
    i_10_229_1249_0, i_10_229_1250_0, i_10_229_1309_0, i_10_229_1311_0,
    i_10_229_1435_0, i_10_229_1624_0, i_10_229_1654_0, i_10_229_1655_0,
    i_10_229_1765_0, i_10_229_1822_0, i_10_229_1823_0, i_10_229_1909_0,
    i_10_229_2095_0, i_10_229_2179_0, i_10_229_2308_0, i_10_229_2350_0,
    i_10_229_2351_0, i_10_229_2407_0, i_10_229_2634_0, i_10_229_2635_0,
    i_10_229_2636_0, i_10_229_2724_0, i_10_229_2727_0, i_10_229_2728_0,
    i_10_229_2734_0, i_10_229_2783_0, i_10_229_2784_0, i_10_229_2830_0,
    i_10_229_2834_0, i_10_229_2883_0, i_10_229_2920_0, i_10_229_2986_0,
    i_10_229_3038_0, i_10_229_3039_0, i_10_229_3041_0, i_10_229_3048_0,
    i_10_229_3271_0, i_10_229_3273_0, i_10_229_3617_0, i_10_229_3652_0,
    i_10_229_3653_0, i_10_229_3783_0, i_10_229_3839_0, i_10_229_3840_0,
    i_10_229_3846_0, i_10_229_3851_0, i_10_229_3895_0, i_10_229_3982_0,
    i_10_229_3983_0, i_10_229_3985_0, i_10_229_4116_0, i_10_229_4120_0,
    i_10_229_4121_0, i_10_229_4125_0, i_10_229_4188_0, i_10_229_4192_0,
    i_10_229_4270_0, i_10_229_4272_0, i_10_229_4290_0, i_10_229_4291_0,
    o_10_229_0_0  );
  input  i_10_229_174_0, i_10_229_175_0, i_10_229_176_0, i_10_229_184_0,
    i_10_229_270_0, i_10_229_286_0, i_10_229_287_0, i_10_229_319_0,
    i_10_229_409_0, i_10_229_410_0, i_10_229_436_0, i_10_229_438_0,
    i_10_229_440_0, i_10_229_446_0, i_10_229_447_0, i_10_229_448_0,
    i_10_229_449_0, i_10_229_466_0, i_10_229_467_0, i_10_229_518_0,
    i_10_229_717_0, i_10_229_718_0, i_10_229_719_0, i_10_229_755_0,
    i_10_229_793_0, i_10_229_797_0, i_10_229_798_0, i_10_229_799_0,
    i_10_229_958_0, i_10_229_968_0, i_10_229_971_0, i_10_229_1003_0,
    i_10_229_1006_0, i_10_229_1164_0, i_10_229_1165_0, i_10_229_1166_0,
    i_10_229_1169_0, i_10_229_1237_0, i_10_229_1245_0, i_10_229_1247_0,
    i_10_229_1249_0, i_10_229_1250_0, i_10_229_1309_0, i_10_229_1311_0,
    i_10_229_1435_0, i_10_229_1624_0, i_10_229_1654_0, i_10_229_1655_0,
    i_10_229_1765_0, i_10_229_1822_0, i_10_229_1823_0, i_10_229_1909_0,
    i_10_229_2095_0, i_10_229_2179_0, i_10_229_2308_0, i_10_229_2350_0,
    i_10_229_2351_0, i_10_229_2407_0, i_10_229_2634_0, i_10_229_2635_0,
    i_10_229_2636_0, i_10_229_2724_0, i_10_229_2727_0, i_10_229_2728_0,
    i_10_229_2734_0, i_10_229_2783_0, i_10_229_2784_0, i_10_229_2830_0,
    i_10_229_2834_0, i_10_229_2883_0, i_10_229_2920_0, i_10_229_2986_0,
    i_10_229_3038_0, i_10_229_3039_0, i_10_229_3041_0, i_10_229_3048_0,
    i_10_229_3271_0, i_10_229_3273_0, i_10_229_3617_0, i_10_229_3652_0,
    i_10_229_3653_0, i_10_229_3783_0, i_10_229_3839_0, i_10_229_3840_0,
    i_10_229_3846_0, i_10_229_3851_0, i_10_229_3895_0, i_10_229_3982_0,
    i_10_229_3983_0, i_10_229_3985_0, i_10_229_4116_0, i_10_229_4120_0,
    i_10_229_4121_0, i_10_229_4125_0, i_10_229_4188_0, i_10_229_4192_0,
    i_10_229_4270_0, i_10_229_4272_0, i_10_229_4290_0, i_10_229_4291_0;
  output o_10_229_0_0;
  assign o_10_229_0_0 = ~((~i_10_229_448_0 & ((~i_10_229_1249_0 & ~i_10_229_1822_0 & ~i_10_229_3840_0) | (~i_10_229_174_0 & ~i_10_229_184_0 & ~i_10_229_449_0 & ~i_10_229_755_0 & ~i_10_229_3895_0))) | (~i_10_229_174_0 & ((i_10_229_466_0 & ~i_10_229_797_0 & ~i_10_229_1164_0 & ~i_10_229_1166_0 & ~i_10_229_2635_0) | (~i_10_229_718_0 & ~i_10_229_719_0 & ~i_10_229_1165_0 & ~i_10_229_1169_0 & ~i_10_229_1245_0 & ~i_10_229_1247_0 & ~i_10_229_2834_0 & ~i_10_229_3038_0))) | (~i_10_229_1166_0 & ((~i_10_229_449_0 & ~i_10_229_1169_0 & ((~i_10_229_446_0 & ~i_10_229_518_0 & ~i_10_229_718_0 & ~i_10_229_799_0 & ~i_10_229_1165_0) | (~i_10_229_1164_0 & ~i_10_229_1823_0 & ~i_10_229_2727_0 & ~i_10_229_2728_0 & ~i_10_229_2920_0))) | (~i_10_229_1164_0 & ((~i_10_229_175_0 & ~i_10_229_718_0 & ~i_10_229_1311_0 & ~i_10_229_1823_0 & ~i_10_229_4270_0) | (~i_10_229_1247_0 & ~i_10_229_1822_0 & ~i_10_229_2351_0 & ~i_10_229_2734_0 & ~i_10_229_4272_0 & ~i_10_229_4290_0))) | (~i_10_229_1250_0 & ((~i_10_229_447_0 & ~i_10_229_466_0) | (~i_10_229_184_0 & ~i_10_229_717_0 & ~i_10_229_958_0 & ~i_10_229_1245_0 & ~i_10_229_1249_0 & ~i_10_229_3895_0))))) | (~i_10_229_717_0 & ((i_10_229_518_0 & ~i_10_229_718_0 & i_10_229_797_0 & ~i_10_229_1164_0 & ~i_10_229_1247_0 & ~i_10_229_1250_0 & ~i_10_229_2728_0) | (~i_10_229_184_0 & i_10_229_799_0 & ~i_10_229_1822_0 & ~i_10_229_2179_0 & ~i_10_229_4120_0 & ~i_10_229_4291_0))) | (~i_10_229_184_0 & ~i_10_229_1247_0 & ((~i_10_229_971_0 & ~i_10_229_1250_0 & i_10_229_3652_0 & ~i_10_229_3846_0) | (~i_10_229_467_0 & ~i_10_229_718_0 & i_10_229_1823_0 & ~i_10_229_3783_0 & ~i_10_229_4291_0))) | (~i_10_229_718_0 & ((~i_10_229_518_0 & ~i_10_229_798_0 & ~i_10_229_2727_0 & ~i_10_229_3038_0 & ~i_10_229_3895_0) | (i_10_229_1309_0 & ~i_10_229_1823_0 & ~i_10_229_4116_0 & i_10_229_4121_0))) | (~i_10_229_1165_0 & ((i_10_229_1435_0 & ~i_10_229_1822_0 & i_10_229_4121_0) | (~i_10_229_719_0 & ~i_10_229_799_0 & ~i_10_229_1164_0 & ~i_10_229_1169_0 & ~i_10_229_2727_0 & ~i_10_229_2734_0 & i_10_229_4116_0 & ~i_10_229_4270_0))));
endmodule



// Benchmark "kernel_10_230" written by ABC on Sun Jul 19 10:24:58 2020

module kernel_10_230 ( 
    i_10_230_268_0, i_10_230_269_0, i_10_230_282_0, i_10_230_283_0,
    i_10_230_315_0, i_10_230_316_0, i_10_230_321_0, i_10_230_327_0,
    i_10_230_390_0, i_10_230_408_0, i_10_230_412_0, i_10_230_439_0,
    i_10_230_440_0, i_10_230_501_0, i_10_230_516_0, i_10_230_664_0,
    i_10_230_685_0, i_10_230_826_0, i_10_230_960_0, i_10_230_969_0,
    i_10_230_1030_0, i_10_230_1105_0, i_10_230_1113_0, i_10_230_1242_0,
    i_10_230_1248_0, i_10_230_1264_0, i_10_230_1302_0, i_10_230_1303_0,
    i_10_230_1357_0, i_10_230_1447_0, i_10_230_1547_0, i_10_230_1556_0,
    i_10_230_1578_0, i_10_230_1579_0, i_10_230_1580_0, i_10_230_1618_0,
    i_10_230_1627_0, i_10_230_1683_0, i_10_230_1689_0, i_10_230_1734_0,
    i_10_230_1735_0, i_10_230_1806_0, i_10_230_1819_0, i_10_230_1821_0,
    i_10_230_1945_0, i_10_230_1984_0, i_10_230_1986_0, i_10_230_2005_0,
    i_10_230_2035_0, i_10_230_2243_0, i_10_230_2353_0, i_10_230_2355_0,
    i_10_230_2356_0, i_10_230_2383_0, i_10_230_2384_0, i_10_230_2449_0,
    i_10_230_2451_0, i_10_230_2452_0, i_10_230_2472_0, i_10_230_2569_0,
    i_10_230_2572_0, i_10_230_2631_0, i_10_230_2635_0, i_10_230_2662_0,
    i_10_230_2733_0, i_10_230_2734_0, i_10_230_2832_0, i_10_230_2919_0,
    i_10_230_2920_0, i_10_230_3037_0, i_10_230_3069_0, i_10_230_3280_0,
    i_10_230_3281_0, i_10_230_3283_0, i_10_230_3329_0, i_10_230_3390_0,
    i_10_230_3391_0, i_10_230_3472_0, i_10_230_3501_0, i_10_230_3504_0,
    i_10_230_3508_0, i_10_230_3540_0, i_10_230_3541_0, i_10_230_3612_0,
    i_10_230_3613_0, i_10_230_3785_0, i_10_230_3837_0, i_10_230_3839_0,
    i_10_230_3841_0, i_10_230_3850_0, i_10_230_3852_0, i_10_230_3859_0,
    i_10_230_3860_0, i_10_230_3871_0, i_10_230_4030_0, i_10_230_4116_0,
    i_10_230_4117_0, i_10_230_4120_0, i_10_230_4171_0, i_10_230_4173_0,
    o_10_230_0_0  );
  input  i_10_230_268_0, i_10_230_269_0, i_10_230_282_0, i_10_230_283_0,
    i_10_230_315_0, i_10_230_316_0, i_10_230_321_0, i_10_230_327_0,
    i_10_230_390_0, i_10_230_408_0, i_10_230_412_0, i_10_230_439_0,
    i_10_230_440_0, i_10_230_501_0, i_10_230_516_0, i_10_230_664_0,
    i_10_230_685_0, i_10_230_826_0, i_10_230_960_0, i_10_230_969_0,
    i_10_230_1030_0, i_10_230_1105_0, i_10_230_1113_0, i_10_230_1242_0,
    i_10_230_1248_0, i_10_230_1264_0, i_10_230_1302_0, i_10_230_1303_0,
    i_10_230_1357_0, i_10_230_1447_0, i_10_230_1547_0, i_10_230_1556_0,
    i_10_230_1578_0, i_10_230_1579_0, i_10_230_1580_0, i_10_230_1618_0,
    i_10_230_1627_0, i_10_230_1683_0, i_10_230_1689_0, i_10_230_1734_0,
    i_10_230_1735_0, i_10_230_1806_0, i_10_230_1819_0, i_10_230_1821_0,
    i_10_230_1945_0, i_10_230_1984_0, i_10_230_1986_0, i_10_230_2005_0,
    i_10_230_2035_0, i_10_230_2243_0, i_10_230_2353_0, i_10_230_2355_0,
    i_10_230_2356_0, i_10_230_2383_0, i_10_230_2384_0, i_10_230_2449_0,
    i_10_230_2451_0, i_10_230_2452_0, i_10_230_2472_0, i_10_230_2569_0,
    i_10_230_2572_0, i_10_230_2631_0, i_10_230_2635_0, i_10_230_2662_0,
    i_10_230_2733_0, i_10_230_2734_0, i_10_230_2832_0, i_10_230_2919_0,
    i_10_230_2920_0, i_10_230_3037_0, i_10_230_3069_0, i_10_230_3280_0,
    i_10_230_3281_0, i_10_230_3283_0, i_10_230_3329_0, i_10_230_3390_0,
    i_10_230_3391_0, i_10_230_3472_0, i_10_230_3501_0, i_10_230_3504_0,
    i_10_230_3508_0, i_10_230_3540_0, i_10_230_3541_0, i_10_230_3612_0,
    i_10_230_3613_0, i_10_230_3785_0, i_10_230_3837_0, i_10_230_3839_0,
    i_10_230_3841_0, i_10_230_3850_0, i_10_230_3852_0, i_10_230_3859_0,
    i_10_230_3860_0, i_10_230_3871_0, i_10_230_4030_0, i_10_230_4116_0,
    i_10_230_4117_0, i_10_230_4120_0, i_10_230_4171_0, i_10_230_4173_0;
  output o_10_230_0_0;
  assign o_10_230_0_0 = 0;
endmodule



// Benchmark "kernel_10_231" written by ABC on Sun Jul 19 10:24:59 2020

module kernel_10_231 ( 
    i_10_231_28_0, i_10_231_29_0, i_10_231_146_0, i_10_231_172_0,
    i_10_231_220_0, i_10_231_243_0, i_10_231_252_0, i_10_231_387_0,
    i_10_231_433_0, i_10_231_519_0, i_10_231_570_0, i_10_231_687_0,
    i_10_231_711_0, i_10_231_712_0, i_10_231_747_0, i_10_231_748_0,
    i_10_231_752_0, i_10_231_846_0, i_10_231_954_0, i_10_231_1029_0,
    i_10_231_1237_0, i_10_231_1305_0, i_10_231_1309_0, i_10_231_1313_0,
    i_10_231_1377_0, i_10_231_1539_0, i_10_231_1575_0, i_10_231_1614_0,
    i_10_231_1617_0, i_10_231_1683_0, i_10_231_1686_0, i_10_231_1688_0,
    i_10_231_1823_0, i_10_231_1826_0, i_10_231_2178_0, i_10_231_2179_0,
    i_10_231_2308_0, i_10_231_2451_0, i_10_231_2462_0, i_10_231_2463_0,
    i_10_231_2470_0, i_10_231_2471_0, i_10_231_2529_0, i_10_231_2530_0,
    i_10_231_2535_0, i_10_231_2601_0, i_10_231_2602_0, i_10_231_2604_0,
    i_10_231_2628_0, i_10_231_2640_0, i_10_231_2662_0, i_10_231_2728_0,
    i_10_231_2830_0, i_10_231_2831_0, i_10_231_2924_0, i_10_231_2995_0,
    i_10_231_3070_0, i_10_231_3072_0, i_10_231_3156_0, i_10_231_3195_0,
    i_10_231_3196_0, i_10_231_3234_0, i_10_231_3278_0, i_10_231_3385_0,
    i_10_231_3386_0, i_10_231_3389_0, i_10_231_3405_0, i_10_231_3406_0,
    i_10_231_3408_0, i_10_231_3441_0, i_10_231_3444_0, i_10_231_3523_0,
    i_10_231_3525_0, i_10_231_3552_0, i_10_231_3586_0, i_10_231_3609_0,
    i_10_231_3612_0, i_10_231_3616_0, i_10_231_3646_0, i_10_231_3649_0,
    i_10_231_3726_0, i_10_231_3780_0, i_10_231_3781_0, i_10_231_3807_0,
    i_10_231_3808_0, i_10_231_3839_0, i_10_231_3845_0, i_10_231_3849_0,
    i_10_231_3879_0, i_10_231_3880_0, i_10_231_4113_0, i_10_231_4114_0,
    i_10_231_4116_0, i_10_231_4117_0, i_10_231_4118_0, i_10_231_4212_0,
    i_10_231_4216_0, i_10_231_4284_0, i_10_231_4456_0, i_10_231_4582_0,
    o_10_231_0_0  );
  input  i_10_231_28_0, i_10_231_29_0, i_10_231_146_0, i_10_231_172_0,
    i_10_231_220_0, i_10_231_243_0, i_10_231_252_0, i_10_231_387_0,
    i_10_231_433_0, i_10_231_519_0, i_10_231_570_0, i_10_231_687_0,
    i_10_231_711_0, i_10_231_712_0, i_10_231_747_0, i_10_231_748_0,
    i_10_231_752_0, i_10_231_846_0, i_10_231_954_0, i_10_231_1029_0,
    i_10_231_1237_0, i_10_231_1305_0, i_10_231_1309_0, i_10_231_1313_0,
    i_10_231_1377_0, i_10_231_1539_0, i_10_231_1575_0, i_10_231_1614_0,
    i_10_231_1617_0, i_10_231_1683_0, i_10_231_1686_0, i_10_231_1688_0,
    i_10_231_1823_0, i_10_231_1826_0, i_10_231_2178_0, i_10_231_2179_0,
    i_10_231_2308_0, i_10_231_2451_0, i_10_231_2462_0, i_10_231_2463_0,
    i_10_231_2470_0, i_10_231_2471_0, i_10_231_2529_0, i_10_231_2530_0,
    i_10_231_2535_0, i_10_231_2601_0, i_10_231_2602_0, i_10_231_2604_0,
    i_10_231_2628_0, i_10_231_2640_0, i_10_231_2662_0, i_10_231_2728_0,
    i_10_231_2830_0, i_10_231_2831_0, i_10_231_2924_0, i_10_231_2995_0,
    i_10_231_3070_0, i_10_231_3072_0, i_10_231_3156_0, i_10_231_3195_0,
    i_10_231_3196_0, i_10_231_3234_0, i_10_231_3278_0, i_10_231_3385_0,
    i_10_231_3386_0, i_10_231_3389_0, i_10_231_3405_0, i_10_231_3406_0,
    i_10_231_3408_0, i_10_231_3441_0, i_10_231_3444_0, i_10_231_3523_0,
    i_10_231_3525_0, i_10_231_3552_0, i_10_231_3586_0, i_10_231_3609_0,
    i_10_231_3612_0, i_10_231_3616_0, i_10_231_3646_0, i_10_231_3649_0,
    i_10_231_3726_0, i_10_231_3780_0, i_10_231_3781_0, i_10_231_3807_0,
    i_10_231_3808_0, i_10_231_3839_0, i_10_231_3845_0, i_10_231_3849_0,
    i_10_231_3879_0, i_10_231_3880_0, i_10_231_4113_0, i_10_231_4114_0,
    i_10_231_4116_0, i_10_231_4117_0, i_10_231_4118_0, i_10_231_4212_0,
    i_10_231_4216_0, i_10_231_4284_0, i_10_231_4456_0, i_10_231_4582_0;
  output o_10_231_0_0;
  assign o_10_231_0_0 = 0;
endmodule



// Benchmark "kernel_10_232" written by ABC on Sun Jul 19 10:25:00 2020

module kernel_10_232 ( 
    i_10_232_177_0, i_10_232_183_0, i_10_232_184_0, i_10_232_186_0,
    i_10_232_187_0, i_10_232_188_0, i_10_232_220_0, i_10_232_244_0,
    i_10_232_282_0, i_10_232_283_0, i_10_232_284_0, i_10_232_316_0,
    i_10_232_406_0, i_10_232_410_0, i_10_232_429_0, i_10_232_436_0,
    i_10_232_437_0, i_10_232_438_0, i_10_232_439_0, i_10_232_442_0,
    i_10_232_459_0, i_10_232_794_0, i_10_232_996_0, i_10_232_1026_0,
    i_10_232_1027_0, i_10_232_1033_0, i_10_232_1042_0, i_10_232_1043_0,
    i_10_232_1236_0, i_10_232_1247_0, i_10_232_1250_0, i_10_232_1435_0,
    i_10_232_1444_0, i_10_232_1445_0, i_10_232_1447_0, i_10_232_1540_0,
    i_10_232_1543_0, i_10_232_1544_0, i_10_232_1547_0, i_10_232_1575_0,
    i_10_232_1576_0, i_10_232_1579_0, i_10_232_1582_0, i_10_232_1583_0,
    i_10_232_1650_0, i_10_232_1652_0, i_10_232_1653_0, i_10_232_1683_0,
    i_10_232_1684_0, i_10_232_1686_0, i_10_232_1820_0, i_10_232_1821_0,
    i_10_232_1915_0, i_10_232_2183_0, i_10_232_2407_0, i_10_232_2473_0,
    i_10_232_2478_0, i_10_232_2566_0, i_10_232_2628_0, i_10_232_2630_0,
    i_10_232_2633_0, i_10_232_2657_0, i_10_232_2658_0, i_10_232_2659_0,
    i_10_232_2660_0, i_10_232_2662_0, i_10_232_2663_0, i_10_232_2680_0,
    i_10_232_2708_0, i_10_232_2716_0, i_10_232_2728_0, i_10_232_2732_0,
    i_10_232_2883_0, i_10_232_2922_0, i_10_232_3040_0, i_10_232_3069_0,
    i_10_232_3070_0, i_10_232_3152_0, i_10_232_3278_0, i_10_232_3329_0,
    i_10_232_3386_0, i_10_232_3408_0, i_10_232_3465_0, i_10_232_3544_0,
    i_10_232_3783_0, i_10_232_3837_0, i_10_232_3838_0, i_10_232_3839_0,
    i_10_232_3842_0, i_10_232_3846_0, i_10_232_3847_0, i_10_232_3895_0,
    i_10_232_4114_0, i_10_232_4273_0, i_10_232_4278_0, i_10_232_4282_0,
    i_10_232_4286_0, i_10_232_4291_0, i_10_232_4292_0, i_10_232_4563_0,
    o_10_232_0_0  );
  input  i_10_232_177_0, i_10_232_183_0, i_10_232_184_0, i_10_232_186_0,
    i_10_232_187_0, i_10_232_188_0, i_10_232_220_0, i_10_232_244_0,
    i_10_232_282_0, i_10_232_283_0, i_10_232_284_0, i_10_232_316_0,
    i_10_232_406_0, i_10_232_410_0, i_10_232_429_0, i_10_232_436_0,
    i_10_232_437_0, i_10_232_438_0, i_10_232_439_0, i_10_232_442_0,
    i_10_232_459_0, i_10_232_794_0, i_10_232_996_0, i_10_232_1026_0,
    i_10_232_1027_0, i_10_232_1033_0, i_10_232_1042_0, i_10_232_1043_0,
    i_10_232_1236_0, i_10_232_1247_0, i_10_232_1250_0, i_10_232_1435_0,
    i_10_232_1444_0, i_10_232_1445_0, i_10_232_1447_0, i_10_232_1540_0,
    i_10_232_1543_0, i_10_232_1544_0, i_10_232_1547_0, i_10_232_1575_0,
    i_10_232_1576_0, i_10_232_1579_0, i_10_232_1582_0, i_10_232_1583_0,
    i_10_232_1650_0, i_10_232_1652_0, i_10_232_1653_0, i_10_232_1683_0,
    i_10_232_1684_0, i_10_232_1686_0, i_10_232_1820_0, i_10_232_1821_0,
    i_10_232_1915_0, i_10_232_2183_0, i_10_232_2407_0, i_10_232_2473_0,
    i_10_232_2478_0, i_10_232_2566_0, i_10_232_2628_0, i_10_232_2630_0,
    i_10_232_2633_0, i_10_232_2657_0, i_10_232_2658_0, i_10_232_2659_0,
    i_10_232_2660_0, i_10_232_2662_0, i_10_232_2663_0, i_10_232_2680_0,
    i_10_232_2708_0, i_10_232_2716_0, i_10_232_2728_0, i_10_232_2732_0,
    i_10_232_2883_0, i_10_232_2922_0, i_10_232_3040_0, i_10_232_3069_0,
    i_10_232_3070_0, i_10_232_3152_0, i_10_232_3278_0, i_10_232_3329_0,
    i_10_232_3386_0, i_10_232_3408_0, i_10_232_3465_0, i_10_232_3544_0,
    i_10_232_3783_0, i_10_232_3837_0, i_10_232_3838_0, i_10_232_3839_0,
    i_10_232_3842_0, i_10_232_3846_0, i_10_232_3847_0, i_10_232_3895_0,
    i_10_232_4114_0, i_10_232_4273_0, i_10_232_4278_0, i_10_232_4282_0,
    i_10_232_4286_0, i_10_232_4291_0, i_10_232_4292_0, i_10_232_4563_0;
  output o_10_232_0_0;
  assign o_10_232_0_0 = ~((~i_10_232_3846_0 & ((~i_10_232_177_0 & ((~i_10_232_1236_0 & ~i_10_232_1544_0 & ~i_10_232_2708_0) | (~i_10_232_282_0 & i_10_232_1579_0 & ~i_10_232_1583_0 & ~i_10_232_1820_0 & ~i_10_232_2566_0 & ~i_10_232_3465_0))) | (~i_10_232_188_0 & ~i_10_232_1042_0 & ~i_10_232_1247_0 & ~i_10_232_1540_0 & ~i_10_232_1547_0 & ~i_10_232_3070_0))) | (~i_10_232_284_0 & ~i_10_232_3408_0 & ((~i_10_232_1250_0 & ~i_10_232_1543_0 & ~i_10_232_1820_0 & i_10_232_4114_0) | (~i_10_232_1544_0 & i_10_232_1650_0 & ~i_10_232_4291_0))) | (~i_10_232_1540_0 & ((~i_10_232_1042_0 & ((~i_10_232_184_0 & ~i_10_232_1543_0 & ~i_10_232_1544_0 & ~i_10_232_4278_0) | (~i_10_232_186_0 & ~i_10_232_1247_0 & ~i_10_232_1683_0 & ~i_10_232_3783_0 & ~i_10_232_4286_0))) | (~i_10_232_410_0 & ~i_10_232_1652_0 & ~i_10_232_2728_0 & ~i_10_232_3040_0 & ~i_10_232_4273_0))) | (~i_10_232_186_0 & ~i_10_232_3465_0 & ((~i_10_232_282_0 & ~i_10_232_3839_0) | (~i_10_232_459_0 & ~i_10_232_1043_0 & ~i_10_232_2566_0 & ~i_10_232_3070_0 & ~i_10_232_4291_0))) | (~i_10_232_2922_0 & ~i_10_232_3783_0 & ((~i_10_232_283_0 & ~i_10_232_2662_0) | (~i_10_232_1915_0 & ~i_10_232_3069_0 & ~i_10_232_3895_0 & ~i_10_232_4286_0 & ~i_10_232_4291_0))) | (i_10_232_2630_0 & i_10_232_2708_0) | (~i_10_232_187_0 & ~i_10_232_316_0 & ~i_10_232_1683_0 & ~i_10_232_3278_0) | (i_10_232_2883_0 & ~i_10_232_4278_0) | (~i_10_232_188_0 & ~i_10_232_3837_0 & ~i_10_232_4286_0 & ~i_10_232_4292_0));
endmodule



// Benchmark "kernel_10_233" written by ABC on Sun Jul 19 10:25:02 2020

module kernel_10_233 ( 
    i_10_233_153_0, i_10_233_243_0, i_10_233_318_0, i_10_233_442_0,
    i_10_233_460_0, i_10_233_463_0, i_10_233_498_0, i_10_233_513_0,
    i_10_233_516_0, i_10_233_565_0, i_10_233_622_0, i_10_233_864_0,
    i_10_233_865_0, i_10_233_903_0, i_10_233_993_0, i_10_233_1026_0,
    i_10_233_1045_0, i_10_233_1080_0, i_10_233_1235_0, i_10_233_1263_0,
    i_10_233_1264_0, i_10_233_1449_0, i_10_233_1450_0, i_10_233_1551_0,
    i_10_233_1623_0, i_10_233_1683_0, i_10_233_1690_0, i_10_233_1809_0,
    i_10_233_1812_0, i_10_233_1819_0, i_10_233_1825_0, i_10_233_1826_0,
    i_10_233_1878_0, i_10_233_1909_0, i_10_233_1910_0, i_10_233_1913_0,
    i_10_233_1989_0, i_10_233_2002_0, i_10_233_2199_0, i_10_233_2200_0,
    i_10_233_2308_0, i_10_233_2349_0, i_10_233_2353_0, i_10_233_2357_0,
    i_10_233_2376_0, i_10_233_2377_0, i_10_233_2450_0, i_10_233_2451_0,
    i_10_233_2452_0, i_10_233_2453_0, i_10_233_2469_0, i_10_233_2505_0,
    i_10_233_2565_0, i_10_233_2574_0, i_10_233_2657_0, i_10_233_2673_0,
    i_10_233_2700_0, i_10_233_2701_0, i_10_233_2703_0, i_10_233_2723_0,
    i_10_233_2732_0, i_10_233_2735_0, i_10_233_2827_0, i_10_233_2880_0,
    i_10_233_2952_0, i_10_233_2961_0, i_10_233_2983_0, i_10_233_3042_0,
    i_10_233_3159_0, i_10_233_3196_0, i_10_233_3283_0, i_10_233_3284_0,
    i_10_233_3315_0, i_10_233_3388_0, i_10_233_3389_0, i_10_233_3555_0,
    i_10_233_3613_0, i_10_233_3614_0, i_10_233_3649_0, i_10_233_3685_0,
    i_10_233_3780_0, i_10_233_3784_0, i_10_233_3810_0, i_10_233_3839_0,
    i_10_233_3843_0, i_10_233_3858_0, i_10_233_3876_0, i_10_233_3979_0,
    i_10_233_4118_0, i_10_233_4121_0, i_10_233_4122_0, i_10_233_4123_0,
    i_10_233_4126_0, i_10_233_4128_0, i_10_233_4186_0, i_10_233_4266_0,
    i_10_233_4286_0, i_10_233_4289_0, i_10_233_4564_0, i_10_233_4566_0,
    o_10_233_0_0  );
  input  i_10_233_153_0, i_10_233_243_0, i_10_233_318_0, i_10_233_442_0,
    i_10_233_460_0, i_10_233_463_0, i_10_233_498_0, i_10_233_513_0,
    i_10_233_516_0, i_10_233_565_0, i_10_233_622_0, i_10_233_864_0,
    i_10_233_865_0, i_10_233_903_0, i_10_233_993_0, i_10_233_1026_0,
    i_10_233_1045_0, i_10_233_1080_0, i_10_233_1235_0, i_10_233_1263_0,
    i_10_233_1264_0, i_10_233_1449_0, i_10_233_1450_0, i_10_233_1551_0,
    i_10_233_1623_0, i_10_233_1683_0, i_10_233_1690_0, i_10_233_1809_0,
    i_10_233_1812_0, i_10_233_1819_0, i_10_233_1825_0, i_10_233_1826_0,
    i_10_233_1878_0, i_10_233_1909_0, i_10_233_1910_0, i_10_233_1913_0,
    i_10_233_1989_0, i_10_233_2002_0, i_10_233_2199_0, i_10_233_2200_0,
    i_10_233_2308_0, i_10_233_2349_0, i_10_233_2353_0, i_10_233_2357_0,
    i_10_233_2376_0, i_10_233_2377_0, i_10_233_2450_0, i_10_233_2451_0,
    i_10_233_2452_0, i_10_233_2453_0, i_10_233_2469_0, i_10_233_2505_0,
    i_10_233_2565_0, i_10_233_2574_0, i_10_233_2657_0, i_10_233_2673_0,
    i_10_233_2700_0, i_10_233_2701_0, i_10_233_2703_0, i_10_233_2723_0,
    i_10_233_2732_0, i_10_233_2735_0, i_10_233_2827_0, i_10_233_2880_0,
    i_10_233_2952_0, i_10_233_2961_0, i_10_233_2983_0, i_10_233_3042_0,
    i_10_233_3159_0, i_10_233_3196_0, i_10_233_3283_0, i_10_233_3284_0,
    i_10_233_3315_0, i_10_233_3388_0, i_10_233_3389_0, i_10_233_3555_0,
    i_10_233_3613_0, i_10_233_3614_0, i_10_233_3649_0, i_10_233_3685_0,
    i_10_233_3780_0, i_10_233_3784_0, i_10_233_3810_0, i_10_233_3839_0,
    i_10_233_3843_0, i_10_233_3858_0, i_10_233_3876_0, i_10_233_3979_0,
    i_10_233_4118_0, i_10_233_4121_0, i_10_233_4122_0, i_10_233_4123_0,
    i_10_233_4126_0, i_10_233_4128_0, i_10_233_4186_0, i_10_233_4266_0,
    i_10_233_4286_0, i_10_233_4289_0, i_10_233_4564_0, i_10_233_4566_0;
  output o_10_233_0_0;
  assign o_10_233_0_0 = ~((~i_10_233_243_0 & ((~i_10_233_2308_0 & ((~i_10_233_1026_0 & ~i_10_233_3614_0 & ((i_10_233_2357_0 & ~i_10_233_2453_0 & ~i_10_233_2827_0 & ~i_10_233_3389_0 & ~i_10_233_3649_0) | (~i_10_233_565_0 & ~i_10_233_1080_0 & ~i_10_233_1264_0 & ~i_10_233_1551_0 & ~i_10_233_1878_0 & ~i_10_233_1909_0 & ~i_10_233_2199_0 & ~i_10_233_3843_0))) | (~i_10_233_1826_0 & ~i_10_233_2199_0 & ~i_10_233_2353_0 & ~i_10_233_2452_0 & i_10_233_2700_0 & ~i_10_233_2827_0 & ~i_10_233_4128_0))) | (~i_10_233_1878_0 & ((~i_10_233_1989_0 & ~i_10_233_2199_0 & ~i_10_233_2349_0 & ~i_10_233_3159_0) | (~i_10_233_993_0 & ~i_10_233_2200_0 & ~i_10_233_2505_0 & ~i_10_233_4122_0 & ~i_10_233_4266_0))))) | (~i_10_233_993_0 & ~i_10_233_1623_0 & ((~i_10_233_2308_0 & ~i_10_233_2353_0 & ~i_10_233_2505_0 & ~i_10_233_3196_0 & ~i_10_233_4121_0 & ~i_10_233_4123_0) | (~i_10_233_1080_0 & ~i_10_233_1264_0 & ~i_10_233_2377_0 & ~i_10_233_4122_0 & ~i_10_233_4566_0))) | (~i_10_233_1080_0 & ~i_10_233_1812_0 & ((~i_10_233_1263_0 & ~i_10_233_1264_0 & ~i_10_233_2308_0 & ~i_10_233_2376_0 & ~i_10_233_4122_0 & ~i_10_233_4123_0 & ~i_10_233_4128_0) | (~i_10_233_516_0 & ~i_10_233_2505_0 & ~i_10_233_3042_0 & ~i_10_233_4286_0))) | (~i_10_233_1909_0 & ((~i_10_233_1989_0 & ~i_10_233_2353_0 & ~i_10_233_3649_0 & ~i_10_233_3979_0 & ~i_10_233_4122_0) | (~i_10_233_2376_0 & ~i_10_233_2673_0 & ~i_10_233_2701_0 & ~i_10_233_3315_0 & ~i_10_233_4126_0))) | (~i_10_233_2701_0 & ((~i_10_233_2723_0 & ~i_10_233_3784_0 & ~i_10_233_3839_0 & i_10_233_4118_0) | (~i_10_233_1825_0 & ~i_10_233_1878_0 & ~i_10_233_2700_0 & ~i_10_233_3979_0 & ~i_10_233_4566_0))) | (~i_10_233_2827_0 & ((~i_10_233_513_0 & i_10_233_3196_0) | (i_10_233_442_0 & ~i_10_233_2353_0 & ~i_10_233_2377_0 & ~i_10_233_3283_0 & ~i_10_233_4123_0))) | (i_10_233_4289_0 & ((~i_10_233_318_0 & ~i_10_233_1826_0 & ~i_10_233_4126_0 & ~i_10_233_4286_0) | (~i_10_233_3159_0 & i_10_233_4121_0 & i_10_233_4564_0))) | (i_10_233_1819_0 & ~i_10_233_2565_0 & i_10_233_3283_0 & ~i_10_233_3649_0) | (~i_10_233_2002_0 & ~i_10_233_2505_0 & ~i_10_233_3042_0 & ~i_10_233_3613_0 & ~i_10_233_3839_0 & ~i_10_233_3979_0 & ~i_10_233_4123_0 & ~i_10_233_4266_0) | (~i_10_233_903_0 & ~i_10_233_1263_0 & i_10_233_3196_0 & ~i_10_233_4128_0 & ~i_10_233_4289_0));
endmodule



// Benchmark "kernel_10_234" written by ABC on Sun Jul 19 10:25:03 2020

module kernel_10_234 ( 
    i_10_234_31_0, i_10_234_318_0, i_10_234_393_0, i_10_234_444_0,
    i_10_234_447_0, i_10_234_459_0, i_10_234_460_0, i_10_234_463_0,
    i_10_234_467_0, i_10_234_792_0, i_10_234_849_0, i_10_234_970_0,
    i_10_234_1036_0, i_10_234_1039_0, i_10_234_1040_0, i_10_234_1242_0,
    i_10_234_1308_0, i_10_234_1360_0, i_10_234_1382_0, i_10_234_1409_0,
    i_10_234_1444_0, i_10_234_1447_0, i_10_234_1465_0, i_10_234_1552_0,
    i_10_234_1650_0, i_10_234_1757_0, i_10_234_1912_0, i_10_234_1918_0,
    i_10_234_2012_0, i_10_234_2029_0, i_10_234_2096_0, i_10_234_2157_0,
    i_10_234_2332_0, i_10_234_2338_0, i_10_234_2339_0, i_10_234_2434_0,
    i_10_234_2445_0, i_10_234_2461_0, i_10_234_2470_0, i_10_234_2526_0,
    i_10_234_2579_0, i_10_234_2632_0, i_10_234_2659_0, i_10_234_2702_0,
    i_10_234_2705_0, i_10_234_2709_0, i_10_234_2710_0, i_10_234_2711_0,
    i_10_234_2714_0, i_10_234_2887_0, i_10_234_2916_0, i_10_234_2917_0,
    i_10_234_2919_0, i_10_234_2924_0, i_10_234_2954_0, i_10_234_3033_0,
    i_10_234_3057_0, i_10_234_3208_0, i_10_234_3277_0, i_10_234_3279_0,
    i_10_234_3284_0, i_10_234_3297_0, i_10_234_3386_0, i_10_234_3387_0,
    i_10_234_3388_0, i_10_234_3391_0, i_10_234_3403_0, i_10_234_3408_0,
    i_10_234_3409_0, i_10_234_3451_0, i_10_234_3496_0, i_10_234_3497_0,
    i_10_234_3500_0, i_10_234_3550_0, i_10_234_3577_0, i_10_234_3611_0,
    i_10_234_3615_0, i_10_234_3684_0, i_10_234_3717_0, i_10_234_3719_0,
    i_10_234_3720_0, i_10_234_3722_0, i_10_234_3854_0, i_10_234_3860_0,
    i_10_234_3889_0, i_10_234_3965_0, i_10_234_4030_0, i_10_234_4119_0,
    i_10_234_4186_0, i_10_234_4188_0, i_10_234_4189_0, i_10_234_4204_0,
    i_10_234_4270_0, i_10_234_4271_0, i_10_234_4272_0, i_10_234_4273_0,
    i_10_234_4274_0, i_10_234_4290_0, i_10_234_4291_0, i_10_234_4531_0,
    o_10_234_0_0  );
  input  i_10_234_31_0, i_10_234_318_0, i_10_234_393_0, i_10_234_444_0,
    i_10_234_447_0, i_10_234_459_0, i_10_234_460_0, i_10_234_463_0,
    i_10_234_467_0, i_10_234_792_0, i_10_234_849_0, i_10_234_970_0,
    i_10_234_1036_0, i_10_234_1039_0, i_10_234_1040_0, i_10_234_1242_0,
    i_10_234_1308_0, i_10_234_1360_0, i_10_234_1382_0, i_10_234_1409_0,
    i_10_234_1444_0, i_10_234_1447_0, i_10_234_1465_0, i_10_234_1552_0,
    i_10_234_1650_0, i_10_234_1757_0, i_10_234_1912_0, i_10_234_1918_0,
    i_10_234_2012_0, i_10_234_2029_0, i_10_234_2096_0, i_10_234_2157_0,
    i_10_234_2332_0, i_10_234_2338_0, i_10_234_2339_0, i_10_234_2434_0,
    i_10_234_2445_0, i_10_234_2461_0, i_10_234_2470_0, i_10_234_2526_0,
    i_10_234_2579_0, i_10_234_2632_0, i_10_234_2659_0, i_10_234_2702_0,
    i_10_234_2705_0, i_10_234_2709_0, i_10_234_2710_0, i_10_234_2711_0,
    i_10_234_2714_0, i_10_234_2887_0, i_10_234_2916_0, i_10_234_2917_0,
    i_10_234_2919_0, i_10_234_2924_0, i_10_234_2954_0, i_10_234_3033_0,
    i_10_234_3057_0, i_10_234_3208_0, i_10_234_3277_0, i_10_234_3279_0,
    i_10_234_3284_0, i_10_234_3297_0, i_10_234_3386_0, i_10_234_3387_0,
    i_10_234_3388_0, i_10_234_3391_0, i_10_234_3403_0, i_10_234_3408_0,
    i_10_234_3409_0, i_10_234_3451_0, i_10_234_3496_0, i_10_234_3497_0,
    i_10_234_3500_0, i_10_234_3550_0, i_10_234_3577_0, i_10_234_3611_0,
    i_10_234_3615_0, i_10_234_3684_0, i_10_234_3717_0, i_10_234_3719_0,
    i_10_234_3720_0, i_10_234_3722_0, i_10_234_3854_0, i_10_234_3860_0,
    i_10_234_3889_0, i_10_234_3965_0, i_10_234_4030_0, i_10_234_4119_0,
    i_10_234_4186_0, i_10_234_4188_0, i_10_234_4189_0, i_10_234_4204_0,
    i_10_234_4270_0, i_10_234_4271_0, i_10_234_4272_0, i_10_234_4273_0,
    i_10_234_4274_0, i_10_234_4290_0, i_10_234_4291_0, i_10_234_4531_0;
  output o_10_234_0_0;
  assign o_10_234_0_0 = 0;
endmodule



// Benchmark "kernel_10_235" written by ABC on Sun Jul 19 10:25:04 2020

module kernel_10_235 ( 
    i_10_235_49_0, i_10_235_173_0, i_10_235_174_0, i_10_235_175_0,
    i_10_235_176_0, i_10_235_244_0, i_10_235_257_0, i_10_235_315_0,
    i_10_235_371_0, i_10_235_389_0, i_10_235_394_0, i_10_235_395_0,
    i_10_235_407_0, i_10_235_411_0, i_10_235_412_0, i_10_235_427_0,
    i_10_235_435_0, i_10_235_439_0, i_10_235_500_0, i_10_235_503_0,
    i_10_235_520_0, i_10_235_521_0, i_10_235_590_0, i_10_235_716_0,
    i_10_235_792_0, i_10_235_989_0, i_10_235_1031_0, i_10_235_1235_0,
    i_10_235_1244_0, i_10_235_1306_0, i_10_235_1313_0, i_10_235_1362_0,
    i_10_235_1436_0, i_10_235_1583_0, i_10_235_1634_0, i_10_235_1654_0,
    i_10_235_1655_0, i_10_235_1685_0, i_10_235_1686_0, i_10_235_1687_0,
    i_10_235_1688_0, i_10_235_1719_0, i_10_235_1720_0, i_10_235_1824_0,
    i_10_235_1826_0, i_10_235_1909_0, i_10_235_2003_0, i_10_235_2198_0,
    i_10_235_2351_0, i_10_235_2352_0, i_10_235_2380_0, i_10_235_2456_0,
    i_10_235_2468_0, i_10_235_2471_0, i_10_235_2531_0, i_10_235_2634_0,
    i_10_235_2690_0, i_10_235_2719_0, i_10_235_2722_0, i_10_235_2732_0,
    i_10_235_2833_0, i_10_235_2834_0, i_10_235_2923_0, i_10_235_3074_0,
    i_10_235_3200_0, i_10_235_3271_0, i_10_235_3278_0, i_10_235_3332_0,
    i_10_235_3466_0, i_10_235_3506_0, i_10_235_3509_0, i_10_235_3610_0,
    i_10_235_3613_0, i_10_235_3616_0, i_10_235_3646_0, i_10_235_3648_0,
    i_10_235_3649_0, i_10_235_3651_0, i_10_235_3652_0, i_10_235_3653_0,
    i_10_235_3721_0, i_10_235_3780_0, i_10_235_3781_0, i_10_235_3782_0,
    i_10_235_3840_0, i_10_235_3841_0, i_10_235_3842_0, i_10_235_3855_0,
    i_10_235_3856_0, i_10_235_3910_0, i_10_235_3911_0, i_10_235_4029_0,
    i_10_235_4126_0, i_10_235_4171_0, i_10_235_4189_0, i_10_235_4268_0,
    i_10_235_4270_0, i_10_235_4271_0, i_10_235_4288_0, i_10_235_4289_0,
    o_10_235_0_0  );
  input  i_10_235_49_0, i_10_235_173_0, i_10_235_174_0, i_10_235_175_0,
    i_10_235_176_0, i_10_235_244_0, i_10_235_257_0, i_10_235_315_0,
    i_10_235_371_0, i_10_235_389_0, i_10_235_394_0, i_10_235_395_0,
    i_10_235_407_0, i_10_235_411_0, i_10_235_412_0, i_10_235_427_0,
    i_10_235_435_0, i_10_235_439_0, i_10_235_500_0, i_10_235_503_0,
    i_10_235_520_0, i_10_235_521_0, i_10_235_590_0, i_10_235_716_0,
    i_10_235_792_0, i_10_235_989_0, i_10_235_1031_0, i_10_235_1235_0,
    i_10_235_1244_0, i_10_235_1306_0, i_10_235_1313_0, i_10_235_1362_0,
    i_10_235_1436_0, i_10_235_1583_0, i_10_235_1634_0, i_10_235_1654_0,
    i_10_235_1655_0, i_10_235_1685_0, i_10_235_1686_0, i_10_235_1687_0,
    i_10_235_1688_0, i_10_235_1719_0, i_10_235_1720_0, i_10_235_1824_0,
    i_10_235_1826_0, i_10_235_1909_0, i_10_235_2003_0, i_10_235_2198_0,
    i_10_235_2351_0, i_10_235_2352_0, i_10_235_2380_0, i_10_235_2456_0,
    i_10_235_2468_0, i_10_235_2471_0, i_10_235_2531_0, i_10_235_2634_0,
    i_10_235_2690_0, i_10_235_2719_0, i_10_235_2722_0, i_10_235_2732_0,
    i_10_235_2833_0, i_10_235_2834_0, i_10_235_2923_0, i_10_235_3074_0,
    i_10_235_3200_0, i_10_235_3271_0, i_10_235_3278_0, i_10_235_3332_0,
    i_10_235_3466_0, i_10_235_3506_0, i_10_235_3509_0, i_10_235_3610_0,
    i_10_235_3613_0, i_10_235_3616_0, i_10_235_3646_0, i_10_235_3648_0,
    i_10_235_3649_0, i_10_235_3651_0, i_10_235_3652_0, i_10_235_3653_0,
    i_10_235_3721_0, i_10_235_3780_0, i_10_235_3781_0, i_10_235_3782_0,
    i_10_235_3840_0, i_10_235_3841_0, i_10_235_3842_0, i_10_235_3855_0,
    i_10_235_3856_0, i_10_235_3910_0, i_10_235_3911_0, i_10_235_4029_0,
    i_10_235_4126_0, i_10_235_4171_0, i_10_235_4189_0, i_10_235_4268_0,
    i_10_235_4270_0, i_10_235_4271_0, i_10_235_4288_0, i_10_235_4289_0;
  output o_10_235_0_0;
  assign o_10_235_0_0 = 0;
endmodule



// Benchmark "kernel_10_236" written by ABC on Sun Jul 19 10:25:04 2020

module kernel_10_236 ( 
    i_10_236_71_0, i_10_236_89_0, i_10_236_145_0, i_10_236_146_0,
    i_10_236_172_0, i_10_236_174_0, i_10_236_175_0, i_10_236_224_0,
    i_10_236_248_0, i_10_236_286_0, i_10_236_287_0, i_10_236_393_0,
    i_10_236_408_0, i_10_236_439_0, i_10_236_446_0, i_10_236_462_0,
    i_10_236_464_0, i_10_236_466_0, i_10_236_691_0, i_10_236_794_0,
    i_10_236_796_0, i_10_236_800_0, i_10_236_1042_0, i_10_236_1043_0,
    i_10_236_1165_0, i_10_236_1168_0, i_10_236_1237_0, i_10_236_1240_0,
    i_10_236_1241_0, i_10_236_1306_0, i_10_236_1308_0, i_10_236_1364_0,
    i_10_236_1450_0, i_10_236_1540_0, i_10_236_1555_0, i_10_236_1613_0,
    i_10_236_1653_0, i_10_236_1654_0, i_10_236_1735_0, i_10_236_1760_0,
    i_10_236_1821_0, i_10_236_1823_0, i_10_236_1824_0, i_10_236_1915_0,
    i_10_236_2159_0, i_10_236_2246_0, i_10_236_2248_0, i_10_236_2249_0,
    i_10_236_2309_0, i_10_236_2329_0, i_10_236_2350_0, i_10_236_2352_0,
    i_10_236_2361_0, i_10_236_2380_0, i_10_236_2451_0, i_10_236_2456_0,
    i_10_236_2473_0, i_10_236_2581_0, i_10_236_2658_0, i_10_236_2730_0,
    i_10_236_2734_0, i_10_236_2841_0, i_10_236_2881_0, i_10_236_2922_0,
    i_10_236_2923_0, i_10_236_2941_0, i_10_236_2942_0, i_10_236_3036_0,
    i_10_236_3037_0, i_10_236_3073_0, i_10_236_3198_0, i_10_236_3202_0,
    i_10_236_3388_0, i_10_236_3405_0, i_10_236_3470_0, i_10_236_3610_0,
    i_10_236_3613_0, i_10_236_3614_0, i_10_236_3615_0, i_10_236_3649_0,
    i_10_236_3674_0, i_10_236_3686_0, i_10_236_3703_0, i_10_236_3788_0,
    i_10_236_3810_0, i_10_236_3838_0, i_10_236_3853_0, i_10_236_3855_0,
    i_10_236_3856_0, i_10_236_3858_0, i_10_236_3859_0, i_10_236_3860_0,
    i_10_236_3883_0, i_10_236_3967_0, i_10_236_4267_0, i_10_236_4270_0,
    i_10_236_4271_0, i_10_236_4292_0, i_10_236_4463_0, i_10_236_4606_0,
    o_10_236_0_0  );
  input  i_10_236_71_0, i_10_236_89_0, i_10_236_145_0, i_10_236_146_0,
    i_10_236_172_0, i_10_236_174_0, i_10_236_175_0, i_10_236_224_0,
    i_10_236_248_0, i_10_236_286_0, i_10_236_287_0, i_10_236_393_0,
    i_10_236_408_0, i_10_236_439_0, i_10_236_446_0, i_10_236_462_0,
    i_10_236_464_0, i_10_236_466_0, i_10_236_691_0, i_10_236_794_0,
    i_10_236_796_0, i_10_236_800_0, i_10_236_1042_0, i_10_236_1043_0,
    i_10_236_1165_0, i_10_236_1168_0, i_10_236_1237_0, i_10_236_1240_0,
    i_10_236_1241_0, i_10_236_1306_0, i_10_236_1308_0, i_10_236_1364_0,
    i_10_236_1450_0, i_10_236_1540_0, i_10_236_1555_0, i_10_236_1613_0,
    i_10_236_1653_0, i_10_236_1654_0, i_10_236_1735_0, i_10_236_1760_0,
    i_10_236_1821_0, i_10_236_1823_0, i_10_236_1824_0, i_10_236_1915_0,
    i_10_236_2159_0, i_10_236_2246_0, i_10_236_2248_0, i_10_236_2249_0,
    i_10_236_2309_0, i_10_236_2329_0, i_10_236_2350_0, i_10_236_2352_0,
    i_10_236_2361_0, i_10_236_2380_0, i_10_236_2451_0, i_10_236_2456_0,
    i_10_236_2473_0, i_10_236_2581_0, i_10_236_2658_0, i_10_236_2730_0,
    i_10_236_2734_0, i_10_236_2841_0, i_10_236_2881_0, i_10_236_2922_0,
    i_10_236_2923_0, i_10_236_2941_0, i_10_236_2942_0, i_10_236_3036_0,
    i_10_236_3037_0, i_10_236_3073_0, i_10_236_3198_0, i_10_236_3202_0,
    i_10_236_3388_0, i_10_236_3405_0, i_10_236_3470_0, i_10_236_3610_0,
    i_10_236_3613_0, i_10_236_3614_0, i_10_236_3615_0, i_10_236_3649_0,
    i_10_236_3674_0, i_10_236_3686_0, i_10_236_3703_0, i_10_236_3788_0,
    i_10_236_3810_0, i_10_236_3838_0, i_10_236_3853_0, i_10_236_3855_0,
    i_10_236_3856_0, i_10_236_3858_0, i_10_236_3859_0, i_10_236_3860_0,
    i_10_236_3883_0, i_10_236_3967_0, i_10_236_4267_0, i_10_236_4270_0,
    i_10_236_4271_0, i_10_236_4292_0, i_10_236_4463_0, i_10_236_4606_0;
  output o_10_236_0_0;
  assign o_10_236_0_0 = 1;
endmodule



// Benchmark "kernel_10_237" written by ABC on Sun Jul 19 10:25:05 2020

module kernel_10_237 ( 
    i_10_237_66_0, i_10_237_121_0, i_10_237_177_0, i_10_237_193_0,
    i_10_237_252_0, i_10_237_253_0, i_10_237_256_0, i_10_237_262_0,
    i_10_237_393_0, i_10_237_499_0, i_10_237_558_0, i_10_237_561_0,
    i_10_237_562_0, i_10_237_606_0, i_10_237_693_0, i_10_237_694_0,
    i_10_237_696_0, i_10_237_759_0, i_10_237_946_0, i_10_237_1002_0,
    i_10_237_1107_0, i_10_237_1110_0, i_10_237_1129_0, i_10_237_1233_0,
    i_10_237_1236_0, i_10_237_1281_0, i_10_237_1282_0, i_10_237_1296_0,
    i_10_237_1299_0, i_10_237_1432_0, i_10_237_1434_0, i_10_237_1435_0,
    i_10_237_1438_0, i_10_237_1539_0, i_10_237_1540_0, i_10_237_1542_0,
    i_10_237_1549_0, i_10_237_1550_0, i_10_237_1552_0, i_10_237_1553_0,
    i_10_237_1624_0, i_10_237_1625_0, i_10_237_1651_0, i_10_237_1654_0,
    i_10_237_1820_0, i_10_237_2092_0, i_10_237_2155_0, i_10_237_2156_0,
    i_10_237_2235_0, i_10_237_2238_0, i_10_237_2244_0, i_10_237_2289_0,
    i_10_237_2290_0, i_10_237_2350_0, i_10_237_2352_0, i_10_237_2353_0,
    i_10_237_2529_0, i_10_237_2531_0, i_10_237_2556_0, i_10_237_2565_0,
    i_10_237_2566_0, i_10_237_2570_0, i_10_237_2584_0, i_10_237_2587_0,
    i_10_237_2595_0, i_10_237_2694_0, i_10_237_2757_0, i_10_237_2782_0,
    i_10_237_2881_0, i_10_237_2944_0, i_10_237_2957_0, i_10_237_2989_0,
    i_10_237_3055_0, i_10_237_3070_0, i_10_237_3171_0, i_10_237_3198_0,
    i_10_237_3277_0, i_10_237_3279_0, i_10_237_3462_0, i_10_237_3567_0,
    i_10_237_3793_0, i_10_237_3858_0, i_10_237_3979_0, i_10_237_4027_0,
    i_10_237_4053_0, i_10_237_4153_0, i_10_237_4156_0, i_10_237_4167_0,
    i_10_237_4170_0, i_10_237_4171_0, i_10_237_4180_0, i_10_237_4189_0,
    i_10_237_4266_0, i_10_237_4275_0, i_10_237_4279_0, i_10_237_4378_0,
    i_10_237_4545_0, i_10_237_4549_0, i_10_237_4563_0, i_10_237_4564_0,
    o_10_237_0_0  );
  input  i_10_237_66_0, i_10_237_121_0, i_10_237_177_0, i_10_237_193_0,
    i_10_237_252_0, i_10_237_253_0, i_10_237_256_0, i_10_237_262_0,
    i_10_237_393_0, i_10_237_499_0, i_10_237_558_0, i_10_237_561_0,
    i_10_237_562_0, i_10_237_606_0, i_10_237_693_0, i_10_237_694_0,
    i_10_237_696_0, i_10_237_759_0, i_10_237_946_0, i_10_237_1002_0,
    i_10_237_1107_0, i_10_237_1110_0, i_10_237_1129_0, i_10_237_1233_0,
    i_10_237_1236_0, i_10_237_1281_0, i_10_237_1282_0, i_10_237_1296_0,
    i_10_237_1299_0, i_10_237_1432_0, i_10_237_1434_0, i_10_237_1435_0,
    i_10_237_1438_0, i_10_237_1539_0, i_10_237_1540_0, i_10_237_1542_0,
    i_10_237_1549_0, i_10_237_1550_0, i_10_237_1552_0, i_10_237_1553_0,
    i_10_237_1624_0, i_10_237_1625_0, i_10_237_1651_0, i_10_237_1654_0,
    i_10_237_1820_0, i_10_237_2092_0, i_10_237_2155_0, i_10_237_2156_0,
    i_10_237_2235_0, i_10_237_2238_0, i_10_237_2244_0, i_10_237_2289_0,
    i_10_237_2290_0, i_10_237_2350_0, i_10_237_2352_0, i_10_237_2353_0,
    i_10_237_2529_0, i_10_237_2531_0, i_10_237_2556_0, i_10_237_2565_0,
    i_10_237_2566_0, i_10_237_2570_0, i_10_237_2584_0, i_10_237_2587_0,
    i_10_237_2595_0, i_10_237_2694_0, i_10_237_2757_0, i_10_237_2782_0,
    i_10_237_2881_0, i_10_237_2944_0, i_10_237_2957_0, i_10_237_2989_0,
    i_10_237_3055_0, i_10_237_3070_0, i_10_237_3171_0, i_10_237_3198_0,
    i_10_237_3277_0, i_10_237_3279_0, i_10_237_3462_0, i_10_237_3567_0,
    i_10_237_3793_0, i_10_237_3858_0, i_10_237_3979_0, i_10_237_4027_0,
    i_10_237_4053_0, i_10_237_4153_0, i_10_237_4156_0, i_10_237_4167_0,
    i_10_237_4170_0, i_10_237_4171_0, i_10_237_4180_0, i_10_237_4189_0,
    i_10_237_4266_0, i_10_237_4275_0, i_10_237_4279_0, i_10_237_4378_0,
    i_10_237_4545_0, i_10_237_4549_0, i_10_237_4563_0, i_10_237_4564_0;
  output o_10_237_0_0;
  assign o_10_237_0_0 = 0;
endmodule



// Benchmark "kernel_10_238" written by ABC on Sun Jul 19 10:25:06 2020

module kernel_10_238 ( 
    i_10_238_171_0, i_10_238_247_0, i_10_238_282_0, i_10_238_286_0,
    i_10_238_287_0, i_10_238_390_0, i_10_238_406_0, i_10_238_408_0,
    i_10_238_429_0, i_10_238_435_0, i_10_238_444_0, i_10_238_445_0,
    i_10_238_448_0, i_10_238_449_0, i_10_238_521_0, i_10_238_793_0,
    i_10_238_966_0, i_10_238_967_0, i_10_238_992_0, i_10_238_1001_0,
    i_10_238_1007_0, i_10_238_1233_0, i_10_238_1238_0, i_10_238_1241_0,
    i_10_238_1246_0, i_10_238_1311_0, i_10_238_1360_0, i_10_238_1541_0,
    i_10_238_1552_0, i_10_238_1553_0, i_10_238_1555_0, i_10_238_1622_0,
    i_10_238_1655_0, i_10_238_1721_0, i_10_238_1730_0, i_10_238_1820_0,
    i_10_238_1824_0, i_10_238_1825_0, i_10_238_1826_0, i_10_238_1913_0,
    i_10_238_2030_0, i_10_238_2332_0, i_10_238_2333_0, i_10_238_2337_0,
    i_10_238_2338_0, i_10_238_2351_0, i_10_238_2352_0, i_10_238_2353_0,
    i_10_238_2377_0, i_10_238_2379_0, i_10_238_2380_0, i_10_238_2381_0,
    i_10_238_2383_0, i_10_238_2384_0, i_10_238_2405_0, i_10_238_2410_0,
    i_10_238_2570_0, i_10_238_2638_0, i_10_238_2656_0, i_10_238_2658_0,
    i_10_238_2659_0, i_10_238_2660_0, i_10_238_2701_0, i_10_238_2716_0,
    i_10_238_2721_0, i_10_238_2734_0, i_10_238_2917_0, i_10_238_2953_0,
    i_10_238_2963_0, i_10_238_2979_0, i_10_238_2980_0, i_10_238_2985_0,
    i_10_238_3038_0, i_10_238_3045_0, i_10_238_3151_0, i_10_238_3152_0,
    i_10_238_3153_0, i_10_238_3154_0, i_10_238_3155_0, i_10_238_3199_0,
    i_10_238_3268_0, i_10_238_3317_0, i_10_238_3388_0, i_10_238_3389_0,
    i_10_238_3437_0, i_10_238_3495_0, i_10_238_3497_0, i_10_238_3582_0,
    i_10_238_3650_0, i_10_238_3837_0, i_10_238_3842_0, i_10_238_3856_0,
    i_10_238_3857_0, i_10_238_3982_0, i_10_238_4114_0, i_10_238_4267_0,
    i_10_238_4270_0, i_10_238_4271_0, i_10_238_4274_0, i_10_238_4565_0,
    o_10_238_0_0  );
  input  i_10_238_171_0, i_10_238_247_0, i_10_238_282_0, i_10_238_286_0,
    i_10_238_287_0, i_10_238_390_0, i_10_238_406_0, i_10_238_408_0,
    i_10_238_429_0, i_10_238_435_0, i_10_238_444_0, i_10_238_445_0,
    i_10_238_448_0, i_10_238_449_0, i_10_238_521_0, i_10_238_793_0,
    i_10_238_966_0, i_10_238_967_0, i_10_238_992_0, i_10_238_1001_0,
    i_10_238_1007_0, i_10_238_1233_0, i_10_238_1238_0, i_10_238_1241_0,
    i_10_238_1246_0, i_10_238_1311_0, i_10_238_1360_0, i_10_238_1541_0,
    i_10_238_1552_0, i_10_238_1553_0, i_10_238_1555_0, i_10_238_1622_0,
    i_10_238_1655_0, i_10_238_1721_0, i_10_238_1730_0, i_10_238_1820_0,
    i_10_238_1824_0, i_10_238_1825_0, i_10_238_1826_0, i_10_238_1913_0,
    i_10_238_2030_0, i_10_238_2332_0, i_10_238_2333_0, i_10_238_2337_0,
    i_10_238_2338_0, i_10_238_2351_0, i_10_238_2352_0, i_10_238_2353_0,
    i_10_238_2377_0, i_10_238_2379_0, i_10_238_2380_0, i_10_238_2381_0,
    i_10_238_2383_0, i_10_238_2384_0, i_10_238_2405_0, i_10_238_2410_0,
    i_10_238_2570_0, i_10_238_2638_0, i_10_238_2656_0, i_10_238_2658_0,
    i_10_238_2659_0, i_10_238_2660_0, i_10_238_2701_0, i_10_238_2716_0,
    i_10_238_2721_0, i_10_238_2734_0, i_10_238_2917_0, i_10_238_2953_0,
    i_10_238_2963_0, i_10_238_2979_0, i_10_238_2980_0, i_10_238_2985_0,
    i_10_238_3038_0, i_10_238_3045_0, i_10_238_3151_0, i_10_238_3152_0,
    i_10_238_3153_0, i_10_238_3154_0, i_10_238_3155_0, i_10_238_3199_0,
    i_10_238_3268_0, i_10_238_3317_0, i_10_238_3388_0, i_10_238_3389_0,
    i_10_238_3437_0, i_10_238_3495_0, i_10_238_3497_0, i_10_238_3582_0,
    i_10_238_3650_0, i_10_238_3837_0, i_10_238_3842_0, i_10_238_3856_0,
    i_10_238_3857_0, i_10_238_3982_0, i_10_238_4114_0, i_10_238_4267_0,
    i_10_238_4270_0, i_10_238_4271_0, i_10_238_4274_0, i_10_238_4565_0;
  output o_10_238_0_0;
  assign o_10_238_0_0 = ~((~i_10_238_1553_0 & ((i_10_238_287_0 & ((~i_10_238_1001_0 & ~i_10_238_1541_0 & i_10_238_1825_0 & i_10_238_1826_0) | (~i_10_238_1555_0 & ~i_10_238_1730_0 & ~i_10_238_1826_0 & ~i_10_238_2379_0))) | (~i_10_238_2405_0 & ~i_10_238_3317_0 & ((~i_10_238_2030_0 & ~i_10_238_2410_0 & i_10_238_3038_0 & i_10_238_3650_0) | (~i_10_238_992_0 & ~i_10_238_1360_0 & ~i_10_238_1622_0 & ~i_10_238_1730_0 & ~i_10_238_2337_0 & ~i_10_238_2379_0 & ~i_10_238_2570_0 & ~i_10_238_2985_0 & ~i_10_238_3842_0))))) | (~i_10_238_444_0 & ((i_10_238_1241_0 & ~i_10_238_1730_0 & ~i_10_238_2353_0 & ~i_10_238_3199_0 & ~i_10_238_3497_0) | (~i_10_238_992_0 & ~i_10_238_1552_0 & ~i_10_238_1622_0 & ~i_10_238_2332_0 & ~i_10_238_2351_0 & ~i_10_238_3045_0 & ~i_10_238_4271_0))) | (~i_10_238_966_0 & ((~i_10_238_1001_0 & ~i_10_238_1622_0 & ~i_10_238_2377_0 & ~i_10_238_2384_0 & ~i_10_238_2734_0 & i_10_238_3388_0) | (~i_10_238_1552_0 & ~i_10_238_1730_0 & ~i_10_238_2333_0 & ~i_10_238_2337_0 & ~i_10_238_2338_0 & ~i_10_238_4271_0 & ~i_10_238_4274_0))) | (~i_10_238_1622_0 & ((~i_10_238_967_0 & ((~i_10_238_448_0 & ~i_10_238_2332_0 & ~i_10_238_2338_0 & ~i_10_238_2351_0 & ~i_10_238_3317_0 & ~i_10_238_3837_0) | (~i_10_238_449_0 & ~i_10_238_1001_0 & ~i_10_238_1007_0 & ~i_10_238_2030_0 & ~i_10_238_2383_0 & ~i_10_238_2980_0 & ~i_10_238_4267_0))) | (~i_10_238_1555_0 & i_10_238_1825_0 & ~i_10_238_2030_0 & ~i_10_238_2338_0 & ~i_10_238_2353_0 & ~i_10_238_2377_0 & ~i_10_238_3497_0) | (~i_10_238_521_0 & ~i_10_238_2352_0 & i_10_238_4114_0))) | (~i_10_238_2405_0 & ((~i_10_238_1007_0 & ((~i_10_238_1555_0 & i_10_238_1820_0 & ~i_10_238_4271_0) | (~i_10_238_390_0 & ~i_10_238_1001_0 & ~i_10_238_2338_0 & ~i_10_238_2377_0 & ~i_10_238_2660_0 & ~i_10_238_2980_0 & ~i_10_238_2985_0 & ~i_10_238_3317_0 & ~i_10_238_3389_0 & ~i_10_238_3495_0 & ~i_10_238_4274_0))) | (~i_10_238_1360_0 & ~i_10_238_1541_0 & ~i_10_238_2351_0 & ~i_10_238_2383_0 & ~i_10_238_2734_0 & ~i_10_238_3268_0 & ~i_10_238_3389_0 & ~i_10_238_3650_0 & ~i_10_238_4274_0))) | i_10_238_1246_0 | (i_10_238_1825_0 & ~i_10_238_2332_0 & i_10_238_2352_0 & ~i_10_238_2410_0 & ~i_10_238_3495_0 & ~i_10_238_4274_0) | (~i_10_238_1555_0 & i_10_238_2353_0 & ~i_10_238_2716_0 & ~i_10_238_3045_0 & ~i_10_238_3268_0 & i_10_238_3837_0 & ~i_10_238_4271_0));
endmodule



// Benchmark "kernel_10_239" written by ABC on Sun Jul 19 10:25:07 2020

module kernel_10_239 ( 
    i_10_239_30_0, i_10_239_61_0, i_10_239_64_0, i_10_239_249_0,
    i_10_239_250_0, i_10_239_258_0, i_10_239_282_0, i_10_239_292_0,
    i_10_239_318_0, i_10_239_319_0, i_10_239_324_0, i_10_239_327_0,
    i_10_239_361_0, i_10_239_405_0, i_10_239_436_0, i_10_239_438_0,
    i_10_239_444_0, i_10_239_445_0, i_10_239_448_0, i_10_239_627_0,
    i_10_239_663_0, i_10_239_870_0, i_10_239_877_0, i_10_239_954_0,
    i_10_239_959_0, i_10_239_1156_0, i_10_239_1159_0, i_10_239_1234_0,
    i_10_239_1260_0, i_10_239_1308_0, i_10_239_1309_0, i_10_239_1347_0,
    i_10_239_1437_0, i_10_239_1441_0, i_10_239_1542_0, i_10_239_1545_0,
    i_10_239_1546_0, i_10_239_1581_0, i_10_239_1626_0, i_10_239_1641_0,
    i_10_239_1689_0, i_10_239_1690_0, i_10_239_1765_0, i_10_239_1766_0,
    i_10_239_1992_0, i_10_239_2022_0, i_10_239_2031_0, i_10_239_2094_0,
    i_10_239_2199_0, i_10_239_2292_0, i_10_239_2323_0, i_10_239_2346_0,
    i_10_239_2352_0, i_10_239_2355_0, i_10_239_2452_0, i_10_239_2470_0,
    i_10_239_2506_0, i_10_239_2535_0, i_10_239_2634_0, i_10_239_2635_0,
    i_10_239_2712_0, i_10_239_2731_0, i_10_239_2742_0, i_10_239_2850_0,
    i_10_239_2868_0, i_10_239_2888_0, i_10_239_2919_0, i_10_239_2967_0,
    i_10_239_2989_0, i_10_239_3075_0, i_10_239_3076_0, i_10_239_3166_0,
    i_10_239_3279_0, i_10_239_3281_0, i_10_239_3328_0, i_10_239_3336_0,
    i_10_239_3391_0, i_10_239_3431_0, i_10_239_3468_0, i_10_239_3469_0,
    i_10_239_3498_0, i_10_239_3586_0, i_10_239_3588_0, i_10_239_3609_0,
    i_10_239_3616_0, i_10_239_3846_0, i_10_239_3913_0, i_10_239_3984_0,
    i_10_239_4011_0, i_10_239_4113_0, i_10_239_4114_0, i_10_239_4116_0,
    i_10_239_4119_0, i_10_239_4209_0, i_10_239_4216_0, i_10_239_4231_0,
    i_10_239_4272_0, i_10_239_4502_0, i_10_239_4505_0, i_10_239_4568_0,
    o_10_239_0_0  );
  input  i_10_239_30_0, i_10_239_61_0, i_10_239_64_0, i_10_239_249_0,
    i_10_239_250_0, i_10_239_258_0, i_10_239_282_0, i_10_239_292_0,
    i_10_239_318_0, i_10_239_319_0, i_10_239_324_0, i_10_239_327_0,
    i_10_239_361_0, i_10_239_405_0, i_10_239_436_0, i_10_239_438_0,
    i_10_239_444_0, i_10_239_445_0, i_10_239_448_0, i_10_239_627_0,
    i_10_239_663_0, i_10_239_870_0, i_10_239_877_0, i_10_239_954_0,
    i_10_239_959_0, i_10_239_1156_0, i_10_239_1159_0, i_10_239_1234_0,
    i_10_239_1260_0, i_10_239_1308_0, i_10_239_1309_0, i_10_239_1347_0,
    i_10_239_1437_0, i_10_239_1441_0, i_10_239_1542_0, i_10_239_1545_0,
    i_10_239_1546_0, i_10_239_1581_0, i_10_239_1626_0, i_10_239_1641_0,
    i_10_239_1689_0, i_10_239_1690_0, i_10_239_1765_0, i_10_239_1766_0,
    i_10_239_1992_0, i_10_239_2022_0, i_10_239_2031_0, i_10_239_2094_0,
    i_10_239_2199_0, i_10_239_2292_0, i_10_239_2323_0, i_10_239_2346_0,
    i_10_239_2352_0, i_10_239_2355_0, i_10_239_2452_0, i_10_239_2470_0,
    i_10_239_2506_0, i_10_239_2535_0, i_10_239_2634_0, i_10_239_2635_0,
    i_10_239_2712_0, i_10_239_2731_0, i_10_239_2742_0, i_10_239_2850_0,
    i_10_239_2868_0, i_10_239_2888_0, i_10_239_2919_0, i_10_239_2967_0,
    i_10_239_2989_0, i_10_239_3075_0, i_10_239_3076_0, i_10_239_3166_0,
    i_10_239_3279_0, i_10_239_3281_0, i_10_239_3328_0, i_10_239_3336_0,
    i_10_239_3391_0, i_10_239_3431_0, i_10_239_3468_0, i_10_239_3469_0,
    i_10_239_3498_0, i_10_239_3586_0, i_10_239_3588_0, i_10_239_3609_0,
    i_10_239_3616_0, i_10_239_3846_0, i_10_239_3913_0, i_10_239_3984_0,
    i_10_239_4011_0, i_10_239_4113_0, i_10_239_4114_0, i_10_239_4116_0,
    i_10_239_4119_0, i_10_239_4209_0, i_10_239_4216_0, i_10_239_4231_0,
    i_10_239_4272_0, i_10_239_4502_0, i_10_239_4505_0, i_10_239_4568_0;
  output o_10_239_0_0;
  assign o_10_239_0_0 = 0;
endmodule



// Benchmark "kernel_10_240" written by ABC on Sun Jul 19 10:25:08 2020

module kernel_10_240 ( 
    i_10_240_159_0, i_10_240_264_0, i_10_240_265_0, i_10_240_273_0,
    i_10_240_274_0, i_10_240_284_0, i_10_240_286_0, i_10_240_439_0,
    i_10_240_444_0, i_10_240_446_0, i_10_240_447_0, i_10_240_465_0,
    i_10_240_467_0, i_10_240_754_0, i_10_240_755_0, i_10_240_797_0,
    i_10_240_799_0, i_10_240_800_0, i_10_240_898_0, i_10_240_899_0,
    i_10_240_964_0, i_10_240_996_0, i_10_240_1002_0, i_10_240_1027_0,
    i_10_240_1031_0, i_10_240_1032_0, i_10_240_1033_0, i_10_240_1034_0,
    i_10_240_1236_0, i_10_240_1241_0, i_10_240_1245_0, i_10_240_1246_0,
    i_10_240_1306_0, i_10_240_1308_0, i_10_240_1309_0, i_10_240_1312_0,
    i_10_240_1431_0, i_10_240_1576_0, i_10_240_1579_0, i_10_240_1597_0,
    i_10_240_1650_0, i_10_240_1651_0, i_10_240_1652_0, i_10_240_1689_0,
    i_10_240_1813_0, i_10_240_1913_0, i_10_240_1920_0, i_10_240_2202_0,
    i_10_240_2363_0, i_10_240_2383_0, i_10_240_2469_0, i_10_240_2473_0,
    i_10_240_2571_0, i_10_240_2609_0, i_10_240_2635_0, i_10_240_2702_0,
    i_10_240_2717_0, i_10_240_2719_0, i_10_240_2734_0, i_10_240_2829_0,
    i_10_240_2833_0, i_10_240_2880_0, i_10_240_2883_0, i_10_240_2918_0,
    i_10_240_2919_0, i_10_240_2921_0, i_10_240_3074_0, i_10_240_3151_0,
    i_10_240_3163_0, i_10_240_3165_0, i_10_240_3166_0, i_10_240_3196_0,
    i_10_240_3200_0, i_10_240_3274_0, i_10_240_3403_0, i_10_240_3409_0,
    i_10_240_3410_0, i_10_240_3589_0, i_10_240_3610_0, i_10_240_3612_0,
    i_10_240_3616_0, i_10_240_3649_0, i_10_240_3653_0, i_10_240_3781_0,
    i_10_240_3782_0, i_10_240_3855_0, i_10_240_3856_0, i_10_240_3880_0,
    i_10_240_3913_0, i_10_240_4116_0, i_10_240_4117_0, i_10_240_4120_0,
    i_10_240_4126_0, i_10_240_4128_0, i_10_240_4129_0, i_10_240_4130_0,
    i_10_240_4219_0, i_10_240_4273_0, i_10_240_4287_0, i_10_240_4288_0,
    o_10_240_0_0  );
  input  i_10_240_159_0, i_10_240_264_0, i_10_240_265_0, i_10_240_273_0,
    i_10_240_274_0, i_10_240_284_0, i_10_240_286_0, i_10_240_439_0,
    i_10_240_444_0, i_10_240_446_0, i_10_240_447_0, i_10_240_465_0,
    i_10_240_467_0, i_10_240_754_0, i_10_240_755_0, i_10_240_797_0,
    i_10_240_799_0, i_10_240_800_0, i_10_240_898_0, i_10_240_899_0,
    i_10_240_964_0, i_10_240_996_0, i_10_240_1002_0, i_10_240_1027_0,
    i_10_240_1031_0, i_10_240_1032_0, i_10_240_1033_0, i_10_240_1034_0,
    i_10_240_1236_0, i_10_240_1241_0, i_10_240_1245_0, i_10_240_1246_0,
    i_10_240_1306_0, i_10_240_1308_0, i_10_240_1309_0, i_10_240_1312_0,
    i_10_240_1431_0, i_10_240_1576_0, i_10_240_1579_0, i_10_240_1597_0,
    i_10_240_1650_0, i_10_240_1651_0, i_10_240_1652_0, i_10_240_1689_0,
    i_10_240_1813_0, i_10_240_1913_0, i_10_240_1920_0, i_10_240_2202_0,
    i_10_240_2363_0, i_10_240_2383_0, i_10_240_2469_0, i_10_240_2473_0,
    i_10_240_2571_0, i_10_240_2609_0, i_10_240_2635_0, i_10_240_2702_0,
    i_10_240_2717_0, i_10_240_2719_0, i_10_240_2734_0, i_10_240_2829_0,
    i_10_240_2833_0, i_10_240_2880_0, i_10_240_2883_0, i_10_240_2918_0,
    i_10_240_2919_0, i_10_240_2921_0, i_10_240_3074_0, i_10_240_3151_0,
    i_10_240_3163_0, i_10_240_3165_0, i_10_240_3166_0, i_10_240_3196_0,
    i_10_240_3200_0, i_10_240_3274_0, i_10_240_3403_0, i_10_240_3409_0,
    i_10_240_3410_0, i_10_240_3589_0, i_10_240_3610_0, i_10_240_3612_0,
    i_10_240_3616_0, i_10_240_3649_0, i_10_240_3653_0, i_10_240_3781_0,
    i_10_240_3782_0, i_10_240_3855_0, i_10_240_3856_0, i_10_240_3880_0,
    i_10_240_3913_0, i_10_240_4116_0, i_10_240_4117_0, i_10_240_4120_0,
    i_10_240_4126_0, i_10_240_4128_0, i_10_240_4129_0, i_10_240_4130_0,
    i_10_240_4219_0, i_10_240_4273_0, i_10_240_4287_0, i_10_240_4288_0;
  output o_10_240_0_0;
  assign o_10_240_0_0 = ~((~i_10_240_755_0 & ((~i_10_240_1033_0 & ~i_10_240_3200_0 & ~i_10_240_3403_0) | (~i_10_240_3165_0 & ~i_10_240_4219_0))) | (~i_10_240_1027_0 & ~i_10_240_2571_0 & ((~i_10_240_1031_0 & ~i_10_240_2734_0) | (i_10_240_1246_0 & i_10_240_3410_0 & i_10_240_3856_0))) | (~i_10_240_3166_0 & ((~i_10_240_1308_0 & ~i_10_240_3409_0) | (~i_10_240_446_0 & ~i_10_240_2609_0 & ~i_10_240_3410_0 & i_10_240_3616_0))) | (~i_10_240_444_0 & ~i_10_240_1431_0 & ~i_10_240_2635_0 & ~i_10_240_2829_0) | (~i_10_240_1034_0 & ~i_10_240_2880_0 & ~i_10_240_3165_0) | (~i_10_240_899_0 & ~i_10_240_1312_0 & ~i_10_240_2383_0 & ~i_10_240_3781_0) | (i_10_240_2880_0 & i_10_240_3196_0 & ~i_10_240_3410_0 & ~i_10_240_3649_0 & ~i_10_240_3782_0) | (~i_10_240_284_0 & ~i_10_240_2717_0 & ~i_10_240_2883_0 & ~i_10_240_3196_0 & ~i_10_240_4116_0) | (~i_10_240_2363_0 & ~i_10_240_4120_0 & ~i_10_240_4128_0) | (i_10_240_1689_0 & ~i_10_240_4219_0) | (~i_10_240_996_0 & i_10_240_2635_0 & ~i_10_240_3200_0 & ~i_10_240_4287_0));
endmodule



// Benchmark "kernel_10_241" written by ABC on Sun Jul 19 10:25:10 2020

module kernel_10_241 ( 
    i_10_241_171_0, i_10_241_172_0, i_10_241_175_0, i_10_241_176_0,
    i_10_241_220_0, i_10_241_221_0, i_10_241_223_0, i_10_241_250_0,
    i_10_241_282_0, i_10_241_283_0, i_10_241_284_0, i_10_241_432_0,
    i_10_241_433_0, i_10_241_434_0, i_10_241_441_0, i_10_241_463_0,
    i_10_241_794_0, i_10_241_797_0, i_10_241_892_0, i_10_241_968_0,
    i_10_241_1082_0, i_10_241_1236_0, i_10_241_1243_0, i_10_241_1244_0,
    i_10_241_1248_0, i_10_241_1347_0, i_10_241_1348_0, i_10_241_1360_0,
    i_10_241_1365_0, i_10_241_1441_0, i_10_241_1575_0, i_10_241_1652_0,
    i_10_241_1683_0, i_10_241_1687_0, i_10_241_1688_0, i_10_241_1768_0,
    i_10_241_1818_0, i_10_241_1819_0, i_10_241_1824_0, i_10_241_1825_0,
    i_10_241_2186_0, i_10_241_2354_0, i_10_241_2361_0, i_10_241_2382_0,
    i_10_241_2384_0, i_10_241_2448_0, i_10_241_2449_0, i_10_241_2450_0,
    i_10_241_2461_0, i_10_241_2469_0, i_10_241_2629_0, i_10_241_2632_0,
    i_10_241_2633_0, i_10_241_2656_0, i_10_241_2657_0, i_10_241_2658_0,
    i_10_241_2659_0, i_10_241_2721_0, i_10_241_2725_0, i_10_241_2727_0,
    i_10_241_2728_0, i_10_241_2729_0, i_10_241_2787_0, i_10_241_2827_0,
    i_10_241_2829_0, i_10_241_2830_0, i_10_241_2831_0, i_10_241_2883_0,
    i_10_241_2916_0, i_10_241_2983_0, i_10_241_3037_0, i_10_241_3039_0,
    i_10_241_3040_0, i_10_241_3075_0, i_10_241_3151_0, i_10_241_3153_0,
    i_10_241_3156_0, i_10_241_3195_0, i_10_241_3198_0, i_10_241_3238_0,
    i_10_241_3384_0, i_10_241_3387_0, i_10_241_3434_0, i_10_241_3610_0,
    i_10_241_3647_0, i_10_241_3648_0, i_10_241_3649_0, i_10_241_3652_0,
    i_10_241_3653_0, i_10_241_3784_0, i_10_241_3786_0, i_10_241_3835_0,
    i_10_241_3840_0, i_10_241_3855_0, i_10_241_3856_0, i_10_241_3857_0,
    i_10_241_3988_0, i_10_241_4056_0, i_10_241_4266_0, i_10_241_4269_0,
    o_10_241_0_0  );
  input  i_10_241_171_0, i_10_241_172_0, i_10_241_175_0, i_10_241_176_0,
    i_10_241_220_0, i_10_241_221_0, i_10_241_223_0, i_10_241_250_0,
    i_10_241_282_0, i_10_241_283_0, i_10_241_284_0, i_10_241_432_0,
    i_10_241_433_0, i_10_241_434_0, i_10_241_441_0, i_10_241_463_0,
    i_10_241_794_0, i_10_241_797_0, i_10_241_892_0, i_10_241_968_0,
    i_10_241_1082_0, i_10_241_1236_0, i_10_241_1243_0, i_10_241_1244_0,
    i_10_241_1248_0, i_10_241_1347_0, i_10_241_1348_0, i_10_241_1360_0,
    i_10_241_1365_0, i_10_241_1441_0, i_10_241_1575_0, i_10_241_1652_0,
    i_10_241_1683_0, i_10_241_1687_0, i_10_241_1688_0, i_10_241_1768_0,
    i_10_241_1818_0, i_10_241_1819_0, i_10_241_1824_0, i_10_241_1825_0,
    i_10_241_2186_0, i_10_241_2354_0, i_10_241_2361_0, i_10_241_2382_0,
    i_10_241_2384_0, i_10_241_2448_0, i_10_241_2449_0, i_10_241_2450_0,
    i_10_241_2461_0, i_10_241_2469_0, i_10_241_2629_0, i_10_241_2632_0,
    i_10_241_2633_0, i_10_241_2656_0, i_10_241_2657_0, i_10_241_2658_0,
    i_10_241_2659_0, i_10_241_2721_0, i_10_241_2725_0, i_10_241_2727_0,
    i_10_241_2728_0, i_10_241_2729_0, i_10_241_2787_0, i_10_241_2827_0,
    i_10_241_2829_0, i_10_241_2830_0, i_10_241_2831_0, i_10_241_2883_0,
    i_10_241_2916_0, i_10_241_2983_0, i_10_241_3037_0, i_10_241_3039_0,
    i_10_241_3040_0, i_10_241_3075_0, i_10_241_3151_0, i_10_241_3153_0,
    i_10_241_3156_0, i_10_241_3195_0, i_10_241_3198_0, i_10_241_3238_0,
    i_10_241_3384_0, i_10_241_3387_0, i_10_241_3434_0, i_10_241_3610_0,
    i_10_241_3647_0, i_10_241_3648_0, i_10_241_3649_0, i_10_241_3652_0,
    i_10_241_3653_0, i_10_241_3784_0, i_10_241_3786_0, i_10_241_3835_0,
    i_10_241_3840_0, i_10_241_3855_0, i_10_241_3856_0, i_10_241_3857_0,
    i_10_241_3988_0, i_10_241_4056_0, i_10_241_4266_0, i_10_241_4269_0;
  output o_10_241_0_0;
  assign o_10_241_0_0 = ~((~i_10_241_250_0 & ((i_10_241_283_0 & ~i_10_241_1082_0 & ~i_10_241_1243_0 & ~i_10_241_1347_0 & ~i_10_241_2656_0 & ~i_10_241_2727_0 & ~i_10_241_3384_0 & ~i_10_241_3434_0 & ~i_10_241_3784_0) | (i_10_241_797_0 & i_10_241_2354_0 & ~i_10_241_2729_0 & ~i_10_241_3855_0))) | (~i_10_241_2829_0 & ((~i_10_241_283_0 & ((~i_10_241_2659_0 & ~i_10_241_2729_0 & ~i_10_241_2787_0 & i_10_241_3040_0) | (~i_10_241_433_0 & ~i_10_241_2354_0 & ~i_10_241_2469_0 & ~i_10_241_2657_0 & ~i_10_241_2727_0 & ~i_10_241_2728_0 & ~i_10_241_4056_0))) | (~i_10_241_433_0 & ~i_10_241_1244_0 & ~i_10_241_1365_0 & ~i_10_241_1575_0 & ~i_10_241_1652_0 & ~i_10_241_2469_0 & ~i_10_241_2787_0 & ~i_10_241_2827_0 & ~i_10_241_3434_0) | (~i_10_241_432_0 & ~i_10_241_1768_0 & i_10_241_2469_0 & ~i_10_241_3040_0 & ~i_10_241_3784_0))) | (~i_10_241_284_0 & ((~i_10_241_463_0 & ~i_10_241_2658_0 & ~i_10_241_2831_0 & ~i_10_241_3649_0) | (i_10_241_441_0 & ~i_10_241_3855_0 & ~i_10_241_3857_0))) | (~i_10_241_4056_0 & ((~i_10_241_432_0 & ~i_10_241_2361_0 & ~i_10_241_3238_0 & ((~i_10_241_1248_0 & ~i_10_241_2461_0 & ~i_10_241_2469_0 & ~i_10_241_3384_0 & i_10_241_3649_0 & i_10_241_3784_0) | (~i_10_241_433_0 & ~i_10_241_1347_0 & ~i_10_241_2629_0 & ~i_10_241_3040_0 & ~i_10_241_3784_0 & ~i_10_241_3855_0))) | (~i_10_241_892_0 & ((~i_10_241_1082_0 & ~i_10_241_2469_0 & ~i_10_241_2830_0 & ~i_10_241_3649_0) | (~i_10_241_1236_0 & ~i_10_241_2629_0 & ~i_10_241_2729_0 & ~i_10_241_3075_0 & i_10_241_3198_0 & ~i_10_241_3855_0 & ~i_10_241_3857_0 & ~i_10_241_3988_0))))) | (~i_10_241_1082_0 & ((~i_10_241_282_0 & ~i_10_241_1348_0 & ~i_10_241_2729_0 & ~i_10_241_3040_0 & ~i_10_241_3384_0 & ~i_10_241_3648_0) | (~i_10_241_2728_0 & ~i_10_241_2830_0 & ~i_10_241_2831_0 & ~i_10_241_3238_0 & ~i_10_241_3855_0 & ~i_10_241_3857_0))) | (~i_10_241_282_0 & ((~i_10_241_1768_0 & ~i_10_241_2354_0 & ~i_10_241_2361_0 & ~i_10_241_2469_0 & ~i_10_241_2632_0 & ~i_10_241_2659_0 & ~i_10_241_2721_0 & ~i_10_241_2729_0) | (~i_10_241_433_0 & i_10_241_1825_0 & ~i_10_241_2657_0 & i_10_241_3835_0 & ~i_10_241_3988_0))) | (~i_10_241_433_0 & ((~i_10_241_1347_0 & ((i_10_241_2448_0 & ~i_10_241_3784_0) | (~i_10_241_2461_0 & ~i_10_241_2629_0 & ~i_10_241_2728_0 & ~i_10_241_3037_0 & ~i_10_241_3648_0 & ~i_10_241_3855_0))) | (i_10_241_1687_0 & ~i_10_241_2186_0 & ~i_10_241_3039_0))) | (~i_10_241_1365_0 & i_10_241_1825_0 & ((~i_10_241_434_0 & i_10_241_463_0 & ~i_10_241_2469_0 & ~i_10_241_2831_0 & i_10_241_3652_0 & ~i_10_241_3786_0) | (~i_10_241_3855_0 & ~i_10_241_3856_0 & ~i_10_241_3988_0))) | (~i_10_241_2657_0 & ((~i_10_241_1348_0 & ~i_10_241_1768_0 & ~i_10_241_2727_0 & ~i_10_241_2916_0 & ~i_10_241_3075_0 & ~i_10_241_3648_0 & ~i_10_241_3653_0 & ~i_10_241_3786_0) | (~i_10_241_2721_0 & ~i_10_241_3039_0 & ~i_10_241_3387_0 & ~i_10_241_3434_0 & ~i_10_241_3856_0 & ~i_10_241_4269_0))) | (i_10_241_250_0 & i_10_241_2725_0 & ~i_10_241_2787_0 & ~i_10_241_3652_0) | (~i_10_241_1360_0 & i_10_241_1819_0 & ~i_10_241_2186_0 & i_10_241_2633_0 & ~i_10_241_2725_0 & i_10_241_2729_0 & ~i_10_241_2916_0 & ~i_10_241_3784_0 & ~i_10_241_3855_0) | (i_10_241_2449_0 & ~i_10_241_2727_0 & ~i_10_241_3434_0 & ~i_10_241_3857_0));
endmodule



// Benchmark "kernel_10_242" written by ABC on Sun Jul 19 10:25:10 2020

module kernel_10_242 ( 
    i_10_242_22_0, i_10_242_172_0, i_10_242_217_0, i_10_242_273_0,
    i_10_242_274_0, i_10_242_282_0, i_10_242_508_0, i_10_242_531_0,
    i_10_242_586_0, i_10_242_729_0, i_10_242_730_0, i_10_242_733_0,
    i_10_242_792_0, i_10_242_828_0, i_10_242_1120_0, i_10_242_1243_0,
    i_10_242_1245_0, i_10_242_1377_0, i_10_242_1378_0, i_10_242_1386_0,
    i_10_242_1440_0, i_10_242_1521_0, i_10_242_1522_0, i_10_242_1559_0,
    i_10_242_1602_0, i_10_242_1649_0, i_10_242_1651_0, i_10_242_1652_0,
    i_10_242_1684_0, i_10_242_1685_0, i_10_242_1693_0, i_10_242_1767_0,
    i_10_242_1768_0, i_10_242_1824_0, i_10_242_1882_0, i_10_242_1913_0,
    i_10_242_1926_0, i_10_242_1929_0, i_10_242_1944_0, i_10_242_1945_0,
    i_10_242_1947_0, i_10_242_1981_0, i_10_242_2181_0, i_10_242_2331_0,
    i_10_242_2334_0, i_10_242_2376_0, i_10_242_2377_0, i_10_242_2380_0,
    i_10_242_2443_0, i_10_242_2475_0, i_10_242_2542_0, i_10_242_2630_0,
    i_10_242_2640_0, i_10_242_2673_0, i_10_242_2674_0, i_10_242_2689_0,
    i_10_242_2728_0, i_10_242_2729_0, i_10_242_2865_0, i_10_242_2872_0,
    i_10_242_2935_0, i_10_242_2965_0, i_10_242_2990_0, i_10_242_3096_0,
    i_10_242_3224_0, i_10_242_3231_0, i_10_242_3404_0, i_10_242_3519_0,
    i_10_242_3520_0, i_10_242_3521_0, i_10_242_3592_0, i_10_242_3614_0,
    i_10_242_3646_0, i_10_242_3726_0, i_10_242_3846_0, i_10_242_3847_0,
    i_10_242_3849_0, i_10_242_3850_0, i_10_242_3861_0, i_10_242_3889_0,
    i_10_242_3906_0, i_10_242_3961_0, i_10_242_4120_0, i_10_242_4176_0,
    i_10_242_4177_0, i_10_242_4266_0, i_10_242_4267_0, i_10_242_4269_0,
    i_10_242_4275_0, i_10_242_4302_0, i_10_242_4305_0, i_10_242_4306_0,
    i_10_242_4432_0, i_10_242_4437_0, i_10_242_4458_0, i_10_242_4459_0,
    i_10_242_4509_0, i_10_242_4510_0, i_10_242_4519_0, i_10_242_4567_0,
    o_10_242_0_0  );
  input  i_10_242_22_0, i_10_242_172_0, i_10_242_217_0, i_10_242_273_0,
    i_10_242_274_0, i_10_242_282_0, i_10_242_508_0, i_10_242_531_0,
    i_10_242_586_0, i_10_242_729_0, i_10_242_730_0, i_10_242_733_0,
    i_10_242_792_0, i_10_242_828_0, i_10_242_1120_0, i_10_242_1243_0,
    i_10_242_1245_0, i_10_242_1377_0, i_10_242_1378_0, i_10_242_1386_0,
    i_10_242_1440_0, i_10_242_1521_0, i_10_242_1522_0, i_10_242_1559_0,
    i_10_242_1602_0, i_10_242_1649_0, i_10_242_1651_0, i_10_242_1652_0,
    i_10_242_1684_0, i_10_242_1685_0, i_10_242_1693_0, i_10_242_1767_0,
    i_10_242_1768_0, i_10_242_1824_0, i_10_242_1882_0, i_10_242_1913_0,
    i_10_242_1926_0, i_10_242_1929_0, i_10_242_1944_0, i_10_242_1945_0,
    i_10_242_1947_0, i_10_242_1981_0, i_10_242_2181_0, i_10_242_2331_0,
    i_10_242_2334_0, i_10_242_2376_0, i_10_242_2377_0, i_10_242_2380_0,
    i_10_242_2443_0, i_10_242_2475_0, i_10_242_2542_0, i_10_242_2630_0,
    i_10_242_2640_0, i_10_242_2673_0, i_10_242_2674_0, i_10_242_2689_0,
    i_10_242_2728_0, i_10_242_2729_0, i_10_242_2865_0, i_10_242_2872_0,
    i_10_242_2935_0, i_10_242_2965_0, i_10_242_2990_0, i_10_242_3096_0,
    i_10_242_3224_0, i_10_242_3231_0, i_10_242_3404_0, i_10_242_3519_0,
    i_10_242_3520_0, i_10_242_3521_0, i_10_242_3592_0, i_10_242_3614_0,
    i_10_242_3646_0, i_10_242_3726_0, i_10_242_3846_0, i_10_242_3847_0,
    i_10_242_3849_0, i_10_242_3850_0, i_10_242_3861_0, i_10_242_3889_0,
    i_10_242_3906_0, i_10_242_3961_0, i_10_242_4120_0, i_10_242_4176_0,
    i_10_242_4177_0, i_10_242_4266_0, i_10_242_4267_0, i_10_242_4269_0,
    i_10_242_4275_0, i_10_242_4302_0, i_10_242_4305_0, i_10_242_4306_0,
    i_10_242_4432_0, i_10_242_4437_0, i_10_242_4458_0, i_10_242_4459_0,
    i_10_242_4509_0, i_10_242_4510_0, i_10_242_4519_0, i_10_242_4567_0;
  output o_10_242_0_0;
  assign o_10_242_0_0 = 0;
endmodule



// Benchmark "kernel_10_243" written by ABC on Sun Jul 19 10:25:12 2020

module kernel_10_243 ( 
    i_10_243_48_0, i_10_243_49_0, i_10_243_50_0, i_10_243_145_0,
    i_10_243_244_0, i_10_243_253_0, i_10_243_274_0, i_10_243_281_0,
    i_10_243_283_0, i_10_243_284_0, i_10_243_320_0, i_10_243_425_0,
    i_10_243_433_0, i_10_243_450_0, i_10_243_515_0, i_10_243_711_0,
    i_10_243_712_0, i_10_243_796_0, i_10_243_800_0, i_10_243_956_0,
    i_10_243_963_0, i_10_243_1000_0, i_10_243_1237_0, i_10_243_1239_0,
    i_10_243_1241_0, i_10_243_1311_0, i_10_243_1360_0, i_10_243_1433_0,
    i_10_243_1532_0, i_10_243_1539_0, i_10_243_1577_0, i_10_243_1653_0,
    i_10_243_1718_0, i_10_243_1768_0, i_10_243_1769_0, i_10_243_1818_0,
    i_10_243_1819_0, i_10_243_1821_0, i_10_243_1911_0, i_10_243_1912_0,
    i_10_243_1913_0, i_10_243_1916_0, i_10_243_1917_0, i_10_243_2366_0,
    i_10_243_2383_0, i_10_243_2450_0, i_10_243_2452_0, i_10_243_2453_0,
    i_10_243_2459_0, i_10_243_2468_0, i_10_243_2470_0, i_10_243_2543_0,
    i_10_243_2629_0, i_10_243_2630_0, i_10_243_2659_0, i_10_243_2710_0,
    i_10_243_2711_0, i_10_243_2715_0, i_10_243_2717_0, i_10_243_2719_0,
    i_10_243_2721_0, i_10_243_2722_0, i_10_243_2723_0, i_10_243_2728_0,
    i_10_243_2729_0, i_10_243_2781_0, i_10_243_2782_0, i_10_243_2783_0,
    i_10_243_2827_0, i_10_243_2829_0, i_10_243_2830_0, i_10_243_2833_0,
    i_10_243_2916_0, i_10_243_2953_0, i_10_243_3069_0, i_10_243_3155_0,
    i_10_243_3196_0, i_10_243_3278_0, i_10_243_3281_0, i_10_243_3384_0,
    i_10_243_3385_0, i_10_243_3386_0, i_10_243_3405_0, i_10_243_3406_0,
    i_10_243_3466_0, i_10_243_3467_0, i_10_243_3522_0, i_10_243_3523_0,
    i_10_243_3615_0, i_10_243_3616_0, i_10_243_3647_0, i_10_243_3648_0,
    i_10_243_3685_0, i_10_243_3834_0, i_10_243_3848_0, i_10_243_3856_0,
    i_10_243_3857_0, i_10_243_4171_0, i_10_243_4231_0, i_10_243_4279_0,
    o_10_243_0_0  );
  input  i_10_243_48_0, i_10_243_49_0, i_10_243_50_0, i_10_243_145_0,
    i_10_243_244_0, i_10_243_253_0, i_10_243_274_0, i_10_243_281_0,
    i_10_243_283_0, i_10_243_284_0, i_10_243_320_0, i_10_243_425_0,
    i_10_243_433_0, i_10_243_450_0, i_10_243_515_0, i_10_243_711_0,
    i_10_243_712_0, i_10_243_796_0, i_10_243_800_0, i_10_243_956_0,
    i_10_243_963_0, i_10_243_1000_0, i_10_243_1237_0, i_10_243_1239_0,
    i_10_243_1241_0, i_10_243_1311_0, i_10_243_1360_0, i_10_243_1433_0,
    i_10_243_1532_0, i_10_243_1539_0, i_10_243_1577_0, i_10_243_1653_0,
    i_10_243_1718_0, i_10_243_1768_0, i_10_243_1769_0, i_10_243_1818_0,
    i_10_243_1819_0, i_10_243_1821_0, i_10_243_1911_0, i_10_243_1912_0,
    i_10_243_1913_0, i_10_243_1916_0, i_10_243_1917_0, i_10_243_2366_0,
    i_10_243_2383_0, i_10_243_2450_0, i_10_243_2452_0, i_10_243_2453_0,
    i_10_243_2459_0, i_10_243_2468_0, i_10_243_2470_0, i_10_243_2543_0,
    i_10_243_2629_0, i_10_243_2630_0, i_10_243_2659_0, i_10_243_2710_0,
    i_10_243_2711_0, i_10_243_2715_0, i_10_243_2717_0, i_10_243_2719_0,
    i_10_243_2721_0, i_10_243_2722_0, i_10_243_2723_0, i_10_243_2728_0,
    i_10_243_2729_0, i_10_243_2781_0, i_10_243_2782_0, i_10_243_2783_0,
    i_10_243_2827_0, i_10_243_2829_0, i_10_243_2830_0, i_10_243_2833_0,
    i_10_243_2916_0, i_10_243_2953_0, i_10_243_3069_0, i_10_243_3155_0,
    i_10_243_3196_0, i_10_243_3278_0, i_10_243_3281_0, i_10_243_3384_0,
    i_10_243_3385_0, i_10_243_3386_0, i_10_243_3405_0, i_10_243_3406_0,
    i_10_243_3466_0, i_10_243_3467_0, i_10_243_3522_0, i_10_243_3523_0,
    i_10_243_3615_0, i_10_243_3616_0, i_10_243_3647_0, i_10_243_3648_0,
    i_10_243_3685_0, i_10_243_3834_0, i_10_243_3848_0, i_10_243_3856_0,
    i_10_243_3857_0, i_10_243_4171_0, i_10_243_4231_0, i_10_243_4279_0;
  output o_10_243_0_0;
  assign o_10_243_0_0 = ~((~i_10_243_320_0 & ((~i_10_243_1913_0 & i_10_243_2719_0 & ~i_10_243_2722_0 & i_10_243_3278_0 & i_10_243_3405_0) | (~i_10_243_281_0 & ~i_10_243_800_0 & i_10_243_1821_0 & ~i_10_243_2729_0 & ~i_10_243_3281_0 & ~i_10_243_3522_0 & ~i_10_243_3834_0 & ~i_10_243_4231_0))) | (~i_10_243_712_0 & ((i_10_243_1237_0 & ~i_10_243_1768_0 & ~i_10_243_2366_0 & i_10_243_2659_0 & ~i_10_243_2719_0) | (~i_10_243_425_0 & ~i_10_243_1913_0 & ~i_10_243_2459_0 & ~i_10_243_3523_0))) | (~i_10_243_3856_0 & ((~i_10_243_425_0 & ((~i_10_243_433_0 & ~i_10_243_1912_0 & ~i_10_243_3278_0 & ~i_10_243_3467_0) | (~i_10_243_1913_0 & ~i_10_243_2711_0 & ~i_10_243_3848_0))) | (~i_10_243_2453_0 & ~i_10_243_2711_0 & ~i_10_243_3615_0 & ~i_10_243_3857_0 & ~i_10_243_4231_0))) | (~i_10_243_433_0 & ((~i_10_243_515_0 & ~i_10_243_2659_0 & ~i_10_243_2717_0 & ~i_10_243_2723_0 & ~i_10_243_2830_0) | (~i_10_243_1768_0 & ~i_10_243_1769_0 & ~i_10_243_1913_0 & ~i_10_243_2453_0 & ~i_10_243_2459_0 & i_10_243_3857_0))) | (~i_10_243_515_0 & ~i_10_243_3278_0 & ((~i_10_243_284_0 & ~i_10_243_2459_0 & ~i_10_243_2715_0 & ~i_10_243_2728_0) | (~i_10_243_145_0 & ~i_10_243_2470_0 & ~i_10_243_2717_0 & ~i_10_243_3386_0 & ~i_10_243_3405_0 & i_10_243_3522_0))) | (~i_10_243_284_0 & ((~i_10_243_145_0 & i_10_243_450_0 & ~i_10_243_1916_0 & ~i_10_243_2470_0 & i_10_243_2629_0 & ~i_10_243_3386_0) | (i_10_243_1819_0 & ~i_10_243_2450_0 & ~i_10_243_3406_0))) | (~i_10_243_145_0 & ((~i_10_243_796_0 & ~i_10_243_1237_0 & ~i_10_243_2366_0 & ~i_10_243_2717_0 & i_10_243_2722_0 & i_10_243_2723_0 & ~i_10_243_2728_0 & ~i_10_243_3281_0 & ~i_10_243_3384_0 & ~i_10_243_3848_0) | (~i_10_243_283_0 & ~i_10_243_800_0 & ~i_10_243_1769_0 & ~i_10_243_1821_0 & ~i_10_243_3616_0 & ~i_10_243_3857_0))) | (~i_10_243_283_0 & ((~i_10_243_2452_0 & i_10_243_2833_0) | (i_10_243_1577_0 & ~i_10_243_1912_0 & ~i_10_243_3386_0))) | (~i_10_243_2459_0 & ((~i_10_243_1241_0 & ~i_10_243_1769_0 & i_10_243_1821_0 & ~i_10_243_2659_0 & ~i_10_243_2719_0) | (~i_10_243_2829_0 & ~i_10_243_3281_0 & ~i_10_243_3685_0 & i_10_243_4231_0))) | (~i_10_243_1769_0 & ((~i_10_243_2453_0 & ~i_10_243_2719_0 & i_10_243_2833_0) | (~i_10_243_2723_0 & ~i_10_243_3385_0))) | (~i_10_243_2719_0 & ((i_10_243_1239_0 & ~i_10_243_1768_0 & i_10_243_3856_0) | (i_10_243_2459_0 & i_10_243_4231_0))) | (i_10_243_1818_0 & ~i_10_243_2830_0 & ~i_10_243_3281_0) | (i_10_243_320_0 & ~i_10_243_2717_0 & ~i_10_243_2723_0 & ~i_10_243_3405_0) | (~i_10_243_2711_0 & i_10_243_2719_0 & i_10_243_2829_0 & i_10_243_2833_0 & ~i_10_243_3616_0));
endmodule



// Benchmark "kernel_10_244" written by ABC on Sun Jul 19 10:25:13 2020

module kernel_10_244 ( 
    i_10_244_277_0, i_10_244_279_0, i_10_244_282_0, i_10_244_286_0,
    i_10_244_287_0, i_10_244_328_0, i_10_244_329_0, i_10_244_405_0,
    i_10_244_408_0, i_10_244_410_0, i_10_244_413_0, i_10_244_424_0,
    i_10_244_425_0, i_10_244_430_0, i_10_244_436_0, i_10_244_439_0,
    i_10_244_440_0, i_10_244_464_0, i_10_244_518_0, i_10_244_713_0,
    i_10_244_796_0, i_10_244_958_0, i_10_244_959_0, i_10_244_996_0,
    i_10_244_997_0, i_10_244_1138_0, i_10_244_1234_0, i_10_244_1238_0,
    i_10_244_1265_0, i_10_244_1346_0, i_10_244_1546_0, i_10_244_1552_0,
    i_10_244_1555_0, i_10_244_1556_0, i_10_244_1768_0, i_10_244_1818_0,
    i_10_244_1819_0, i_10_244_1823_0, i_10_244_1825_0, i_10_244_1826_0,
    i_10_244_1912_0, i_10_244_1915_0, i_10_244_2021_0, i_10_244_2407_0,
    i_10_244_2408_0, i_10_244_2471_0, i_10_244_2474_0, i_10_244_2508_0,
    i_10_244_2515_0, i_10_244_2542_0, i_10_244_2633_0, i_10_244_2656_0,
    i_10_244_2658_0, i_10_244_2679_0, i_10_244_2680_0, i_10_244_2681_0,
    i_10_244_2705_0, i_10_244_2707_0, i_10_244_2723_0, i_10_244_2726_0,
    i_10_244_2730_0, i_10_244_2732_0, i_10_244_2785_0, i_10_244_2823_0,
    i_10_244_2829_0, i_10_244_2830_0, i_10_244_2831_0, i_10_244_2959_0,
    i_10_244_2979_0, i_10_244_2983_0, i_10_244_2984_0, i_10_244_2986_0,
    i_10_244_3034_0, i_10_244_3039_0, i_10_244_3070_0, i_10_244_3072_0,
    i_10_244_3157_0, i_10_244_3158_0, i_10_244_3387_0, i_10_244_3391_0,
    i_10_244_3496_0, i_10_244_3497_0, i_10_244_3499_0, i_10_244_3519_0,
    i_10_244_3522_0, i_10_244_3523_0, i_10_244_3525_0, i_10_244_3586_0,
    i_10_244_3612_0, i_10_244_3613_0, i_10_244_3614_0, i_10_244_3648_0,
    i_10_244_3784_0, i_10_244_3786_0, i_10_244_3839_0, i_10_244_3847_0,
    i_10_244_3849_0, i_10_244_3855_0, i_10_244_3985_0, i_10_244_3986_0,
    o_10_244_0_0  );
  input  i_10_244_277_0, i_10_244_279_0, i_10_244_282_0, i_10_244_286_0,
    i_10_244_287_0, i_10_244_328_0, i_10_244_329_0, i_10_244_405_0,
    i_10_244_408_0, i_10_244_410_0, i_10_244_413_0, i_10_244_424_0,
    i_10_244_425_0, i_10_244_430_0, i_10_244_436_0, i_10_244_439_0,
    i_10_244_440_0, i_10_244_464_0, i_10_244_518_0, i_10_244_713_0,
    i_10_244_796_0, i_10_244_958_0, i_10_244_959_0, i_10_244_996_0,
    i_10_244_997_0, i_10_244_1138_0, i_10_244_1234_0, i_10_244_1238_0,
    i_10_244_1265_0, i_10_244_1346_0, i_10_244_1546_0, i_10_244_1552_0,
    i_10_244_1555_0, i_10_244_1556_0, i_10_244_1768_0, i_10_244_1818_0,
    i_10_244_1819_0, i_10_244_1823_0, i_10_244_1825_0, i_10_244_1826_0,
    i_10_244_1912_0, i_10_244_1915_0, i_10_244_2021_0, i_10_244_2407_0,
    i_10_244_2408_0, i_10_244_2471_0, i_10_244_2474_0, i_10_244_2508_0,
    i_10_244_2515_0, i_10_244_2542_0, i_10_244_2633_0, i_10_244_2656_0,
    i_10_244_2658_0, i_10_244_2679_0, i_10_244_2680_0, i_10_244_2681_0,
    i_10_244_2705_0, i_10_244_2707_0, i_10_244_2723_0, i_10_244_2726_0,
    i_10_244_2730_0, i_10_244_2732_0, i_10_244_2785_0, i_10_244_2823_0,
    i_10_244_2829_0, i_10_244_2830_0, i_10_244_2831_0, i_10_244_2959_0,
    i_10_244_2979_0, i_10_244_2983_0, i_10_244_2984_0, i_10_244_2986_0,
    i_10_244_3034_0, i_10_244_3039_0, i_10_244_3070_0, i_10_244_3072_0,
    i_10_244_3157_0, i_10_244_3158_0, i_10_244_3387_0, i_10_244_3391_0,
    i_10_244_3496_0, i_10_244_3497_0, i_10_244_3499_0, i_10_244_3519_0,
    i_10_244_3522_0, i_10_244_3523_0, i_10_244_3525_0, i_10_244_3586_0,
    i_10_244_3612_0, i_10_244_3613_0, i_10_244_3614_0, i_10_244_3648_0,
    i_10_244_3784_0, i_10_244_3786_0, i_10_244_3839_0, i_10_244_3847_0,
    i_10_244_3849_0, i_10_244_3855_0, i_10_244_3985_0, i_10_244_3986_0;
  output o_10_244_0_0;
  assign o_10_244_0_0 = ~((~i_10_244_1915_0 & ((~i_10_244_1265_0 & ((~i_10_244_279_0 & ((~i_10_244_410_0 & ~i_10_244_958_0 & ~i_10_244_997_0 & ~i_10_244_1552_0 & ~i_10_244_1825_0 & ~i_10_244_2732_0 & ~i_10_244_2984_0 & ~i_10_244_2986_0 & ~i_10_244_3522_0 & ~i_10_244_3648_0 & ~i_10_244_3839_0) | (~i_10_244_413_0 & ~i_10_244_425_0 & ~i_10_244_1555_0 & ~i_10_244_1556_0 & ~i_10_244_2021_0 & ~i_10_244_2408_0 & ~i_10_244_2508_0 & ~i_10_244_2680_0 & ~i_10_244_2681_0 & ~i_10_244_3612_0 & ~i_10_244_3849_0 & ~i_10_244_3855_0))) | (i_10_244_958_0 & i_10_244_2656_0) | (~i_10_244_328_0 & ~i_10_244_430_0 & ~i_10_244_436_0 & ~i_10_244_440_0 & ~i_10_244_796_0 & ~i_10_244_997_0 & ~i_10_244_1552_0 & ~i_10_244_2707_0 & ~i_10_244_2730_0 & ~i_10_244_3612_0))) | (~i_10_244_436_0 & ((~i_10_244_996_0 & ~i_10_244_3039_0 & ~i_10_244_3523_0 & i_10_244_3612_0 & ~i_10_244_3839_0 & i_10_244_3855_0) | (~i_10_244_329_0 & ~i_10_244_997_0 & ~i_10_244_1238_0 & ~i_10_244_1552_0 & ~i_10_244_1826_0 & ~i_10_244_2407_0 & ~i_10_244_2508_0 & ~i_10_244_2732_0 & ~i_10_244_2983_0 & ~i_10_244_2986_0 & ~i_10_244_3849_0 & ~i_10_244_3985_0))) | (~i_10_244_329_0 & ~i_10_244_439_0 & ~i_10_244_2979_0 & ((~i_10_244_328_0 & ~i_10_244_405_0 & ~i_10_244_410_0 & ~i_10_244_424_0 & ~i_10_244_2984_0 & ~i_10_244_2986_0 & ~i_10_244_430_0 & ~i_10_244_997_0) | (~i_10_244_518_0 & ~i_10_244_1552_0 & ~i_10_244_1823_0 & ~i_10_244_2508_0 & ~i_10_244_2823_0 & ~i_10_244_2983_0 & ~i_10_244_3522_0))))) | (~i_10_244_1555_0 & ((~i_10_244_328_0 & ~i_10_244_2680_0 & ((~i_10_244_424_0 & ~i_10_244_425_0 & ~i_10_244_439_0 & ~i_10_244_440_0 & ~i_10_244_1265_0 & ~i_10_244_2408_0 & ~i_10_244_2679_0 & ~i_10_244_2983_0 & ~i_10_244_2984_0 & ~i_10_244_3497_0) | (i_10_244_282_0 & ~i_10_244_713_0 & ~i_10_244_2407_0 & ~i_10_244_3525_0 & ~i_10_244_3849_0 & i_10_244_3855_0 & ~i_10_244_3986_0))) | (~i_10_244_713_0 & ~i_10_244_2979_0 & ((i_10_244_286_0 & ~i_10_244_436_0 & ~i_10_244_1265_0 & ~i_10_244_2407_0 & ~i_10_244_2508_0 & ~i_10_244_3034_0 & ~i_10_244_3499_0 & ~i_10_244_3519_0 & ~i_10_244_3612_0) | (~i_10_244_439_0 & ~i_10_244_997_0 & ~i_10_244_1556_0 & ~i_10_244_2408_0 & ~i_10_244_2633_0 & ~i_10_244_2785_0 & ~i_10_244_2983_0 & ~i_10_244_2986_0 & ~i_10_244_3497_0 & ~i_10_244_3985_0))) | (~i_10_244_1552_0 & ~i_10_244_2656_0 & ~i_10_244_2679_0 & ((~i_10_244_2407_0 & ~i_10_244_2633_0 & ~i_10_244_2705_0 & ~i_10_244_2726_0 & ~i_10_244_3525_0) | (~i_10_244_425_0 & ~i_10_244_1346_0 & ~i_10_244_2829_0 & ~i_10_244_2983_0 & ~i_10_244_2986_0 & ~i_10_244_3519_0 & ~i_10_244_3614_0 & ~i_10_244_3986_0))))) | (~i_10_244_329_0 & ((~i_10_244_279_0 & ~i_10_244_518_0 & ~i_10_244_996_0 & ~i_10_244_1552_0 & ((~i_10_244_282_0 & ~i_10_244_430_0 & ~i_10_244_1826_0 & ~i_10_244_2508_0 & ~i_10_244_2707_0 & ~i_10_244_2785_0 & ~i_10_244_2979_0) | (~i_10_244_1346_0 & ~i_10_244_2474_0 & ~i_10_244_2681_0 & ~i_10_244_2823_0 & ~i_10_244_3648_0 & ~i_10_244_3839_0 & ~i_10_244_3855_0 & ~i_10_244_3985_0 & ~i_10_244_3986_0))) | (~i_10_244_2408_0 & ~i_10_244_2679_0 & ~i_10_244_430_0 & ~i_10_244_796_0 & ~i_10_244_2829_0 & ~i_10_244_2983_0 & ~i_10_244_3613_0 & ~i_10_244_3986_0))) | (~i_10_244_1552_0 & ((~i_10_244_279_0 & ((i_10_244_464_0 & ~i_10_244_518_0 & ~i_10_244_996_0 & ~i_10_244_997_0 & ~i_10_244_1556_0 & ~i_10_244_1819_0 & ~i_10_244_2681_0 & ~i_10_244_2979_0 & ~i_10_244_3039_0 & i_10_244_3613_0) | (~i_10_244_796_0 & ~i_10_244_2021_0 & ~i_10_244_2656_0 & ~i_10_244_2680_0 & ~i_10_244_2730_0 & ~i_10_244_2823_0 & ~i_10_244_2984_0 & ~i_10_244_3614_0 & ~i_10_244_3849_0))) | (~i_10_244_282_0 & ((~i_10_244_2831_0 & i_10_244_3391_0 & i_10_244_3612_0) | (~i_10_244_424_0 & ~i_10_244_440_0 & ~i_10_244_2471_0 & ~i_10_244_2508_0 & ~i_10_244_2979_0 & ~i_10_244_3525_0 & i_10_244_3855_0))) | (~i_10_244_440_0 & ~i_10_244_518_0 & ~i_10_244_2408_0 & ~i_10_244_2471_0 & i_10_244_2723_0 & ~i_10_244_2979_0 & ~i_10_244_3496_0 & ~i_10_244_3499_0 & ~i_10_244_3612_0))) | (~i_10_244_436_0 & ((i_10_244_1825_0 & ~i_10_244_2633_0 & ~i_10_244_2656_0 & ~i_10_244_2680_0 & ~i_10_244_2707_0 & ~i_10_244_2983_0) | (~i_10_244_440_0 & ~i_10_244_2730_0 & ~i_10_244_3523_0 & ~i_10_244_3612_0 & i_10_244_3613_0 & ~i_10_244_3784_0))) | (~i_10_244_2705_0 & ~i_10_244_2983_0 & i_10_244_3523_0 & i_10_244_3847_0) | (i_10_244_287_0 & ~i_10_244_1912_0 & ~i_10_244_2730_0 & i_10_244_3612_0 & ~i_10_244_3985_0));
endmodule



// Benchmark "kernel_10_245" written by ABC on Sun Jul 19 10:25:14 2020

module kernel_10_245 ( 
    i_10_245_17_0, i_10_245_149_0, i_10_245_187_0, i_10_245_242_0,
    i_10_245_263_0, i_10_245_431_0, i_10_245_448_0, i_10_245_463_0,
    i_10_245_563_0, i_10_245_586_0, i_10_245_587_0, i_10_245_659_0,
    i_10_245_694_0, i_10_245_712_0, i_10_245_824_0, i_10_245_892_0,
    i_10_245_893_0, i_10_245_896_0, i_10_245_899_0, i_10_245_950_0,
    i_10_245_997_0, i_10_245_1000_0, i_10_245_1109_0, i_10_245_1111_0,
    i_10_245_1112_0, i_10_245_1237_0, i_10_245_1270_0, i_10_245_1283_0,
    i_10_245_1300_0, i_10_245_1301_0, i_10_245_1304_0, i_10_245_1345_0,
    i_10_245_1346_0, i_10_245_1388_0, i_10_245_1439_0, i_10_245_1577_0,
    i_10_245_1579_0, i_10_245_1606_0, i_10_245_1732_0, i_10_245_1765_0,
    i_10_245_1799_0, i_10_245_1807_0, i_10_245_1883_0, i_10_245_1913_0,
    i_10_245_1940_0, i_10_245_1985_0, i_10_245_2011_0, i_10_245_2030_0,
    i_10_245_2152_0, i_10_245_2200_0, i_10_245_2210_0, i_10_245_2291_0,
    i_10_245_2350_0, i_10_245_2351_0, i_10_245_2450_0, i_10_245_2453_0,
    i_10_245_2515_0, i_10_245_2533_0, i_10_245_2556_0, i_10_245_2558_0,
    i_10_245_2560_0, i_10_245_2567_0, i_10_245_2570_0, i_10_245_2573_0,
    i_10_245_2660_0, i_10_245_2711_0, i_10_245_2713_0, i_10_245_2833_0,
    i_10_245_2846_0, i_10_245_2876_0, i_10_245_2885_0, i_10_245_2888_0,
    i_10_245_2957_0, i_10_245_3173_0, i_10_245_3277_0, i_10_245_3359_0,
    i_10_245_3395_0, i_10_245_3406_0, i_10_245_3464_0, i_10_245_3470_0,
    i_10_245_3520_0, i_10_245_3521_0, i_10_245_3560_0, i_10_245_3614_0,
    i_10_245_3649_0, i_10_245_3652_0, i_10_245_3841_0, i_10_245_3842_0,
    i_10_245_3920_0, i_10_245_3974_0, i_10_245_3983_0, i_10_245_4031_0,
    i_10_245_4117_0, i_10_245_4145_0, i_10_245_4151_0, i_10_245_4169_0,
    i_10_245_4172_0, i_10_245_4181_0, i_10_245_4268_0, i_10_245_4286_0,
    o_10_245_0_0  );
  input  i_10_245_17_0, i_10_245_149_0, i_10_245_187_0, i_10_245_242_0,
    i_10_245_263_0, i_10_245_431_0, i_10_245_448_0, i_10_245_463_0,
    i_10_245_563_0, i_10_245_586_0, i_10_245_587_0, i_10_245_659_0,
    i_10_245_694_0, i_10_245_712_0, i_10_245_824_0, i_10_245_892_0,
    i_10_245_893_0, i_10_245_896_0, i_10_245_899_0, i_10_245_950_0,
    i_10_245_997_0, i_10_245_1000_0, i_10_245_1109_0, i_10_245_1111_0,
    i_10_245_1112_0, i_10_245_1237_0, i_10_245_1270_0, i_10_245_1283_0,
    i_10_245_1300_0, i_10_245_1301_0, i_10_245_1304_0, i_10_245_1345_0,
    i_10_245_1346_0, i_10_245_1388_0, i_10_245_1439_0, i_10_245_1577_0,
    i_10_245_1579_0, i_10_245_1606_0, i_10_245_1732_0, i_10_245_1765_0,
    i_10_245_1799_0, i_10_245_1807_0, i_10_245_1883_0, i_10_245_1913_0,
    i_10_245_1940_0, i_10_245_1985_0, i_10_245_2011_0, i_10_245_2030_0,
    i_10_245_2152_0, i_10_245_2200_0, i_10_245_2210_0, i_10_245_2291_0,
    i_10_245_2350_0, i_10_245_2351_0, i_10_245_2450_0, i_10_245_2453_0,
    i_10_245_2515_0, i_10_245_2533_0, i_10_245_2556_0, i_10_245_2558_0,
    i_10_245_2560_0, i_10_245_2567_0, i_10_245_2570_0, i_10_245_2573_0,
    i_10_245_2660_0, i_10_245_2711_0, i_10_245_2713_0, i_10_245_2833_0,
    i_10_245_2846_0, i_10_245_2876_0, i_10_245_2885_0, i_10_245_2888_0,
    i_10_245_2957_0, i_10_245_3173_0, i_10_245_3277_0, i_10_245_3359_0,
    i_10_245_3395_0, i_10_245_3406_0, i_10_245_3464_0, i_10_245_3470_0,
    i_10_245_3520_0, i_10_245_3521_0, i_10_245_3560_0, i_10_245_3614_0,
    i_10_245_3649_0, i_10_245_3652_0, i_10_245_3841_0, i_10_245_3842_0,
    i_10_245_3920_0, i_10_245_3974_0, i_10_245_3983_0, i_10_245_4031_0,
    i_10_245_4117_0, i_10_245_4145_0, i_10_245_4151_0, i_10_245_4169_0,
    i_10_245_4172_0, i_10_245_4181_0, i_10_245_4268_0, i_10_245_4286_0;
  output o_10_245_0_0;
  assign o_10_245_0_0 = 0;
endmodule



// Benchmark "kernel_10_246" written by ABC on Sun Jul 19 10:25:15 2020

module kernel_10_246 ( 
    i_10_246_35_0, i_10_246_122_0, i_10_246_161_0, i_10_246_251_0,
    i_10_246_323_0, i_10_246_349_0, i_10_246_390_0, i_10_246_391_0,
    i_10_246_436_0, i_10_246_446_0, i_10_246_448_0, i_10_246_449_0,
    i_10_246_462_0, i_10_246_465_0, i_10_246_601_0, i_10_246_754_0,
    i_10_246_957_0, i_10_246_998_0, i_10_246_1004_0, i_10_246_1033_0,
    i_10_246_1034_0, i_10_246_1052_0, i_10_246_1058_0, i_10_246_1083_0,
    i_10_246_1084_0, i_10_246_1223_0, i_10_246_1291_0, i_10_246_1308_0,
    i_10_246_1382_0, i_10_246_1385_0, i_10_246_1579_0, i_10_246_1580_0,
    i_10_246_1651_0, i_10_246_1655_0, i_10_246_1736_0, i_10_246_1816_0,
    i_10_246_1818_0, i_10_246_1822_0, i_10_246_1823_0, i_10_246_1913_0,
    i_10_246_1961_0, i_10_246_2024_0, i_10_246_2086_0, i_10_246_2264_0,
    i_10_246_2384_0, i_10_246_2452_0, i_10_246_2453_0, i_10_246_2474_0,
    i_10_246_2609_0, i_10_246_2617_0, i_10_246_2657_0, i_10_246_2658_0,
    i_10_246_2700_0, i_10_246_2707_0, i_10_246_2715_0, i_10_246_2786_0,
    i_10_246_2788_0, i_10_246_2789_0, i_10_246_2824_0, i_10_246_2825_0,
    i_10_246_2959_0, i_10_246_2995_0, i_10_246_3094_0, i_10_246_3167_0,
    i_10_246_3238_0, i_10_246_3239_0, i_10_246_3269_0, i_10_246_3280_0,
    i_10_246_3281_0, i_10_246_3419_0, i_10_246_3434_0, i_10_246_3473_0,
    i_10_246_3505_0, i_10_246_3508_0, i_10_246_3526_0, i_10_246_3527_0,
    i_10_246_3587_0, i_10_246_3647_0, i_10_246_3848_0, i_10_246_3883_0,
    i_10_246_3913_0, i_10_246_3914_0, i_10_246_3950_0, i_10_246_3985_0,
    i_10_246_3991_0, i_10_246_3992_0, i_10_246_4004_0, i_10_246_4057_0,
    i_10_246_4113_0, i_10_246_4118_0, i_10_246_4120_0, i_10_246_4130_0,
    i_10_246_4168_0, i_10_246_4172_0, i_10_246_4174_0, i_10_246_4276_0,
    i_10_246_4279_0, i_10_246_4281_0, i_10_246_4454_0, i_10_246_4568_0,
    o_10_246_0_0  );
  input  i_10_246_35_0, i_10_246_122_0, i_10_246_161_0, i_10_246_251_0,
    i_10_246_323_0, i_10_246_349_0, i_10_246_390_0, i_10_246_391_0,
    i_10_246_436_0, i_10_246_446_0, i_10_246_448_0, i_10_246_449_0,
    i_10_246_462_0, i_10_246_465_0, i_10_246_601_0, i_10_246_754_0,
    i_10_246_957_0, i_10_246_998_0, i_10_246_1004_0, i_10_246_1033_0,
    i_10_246_1034_0, i_10_246_1052_0, i_10_246_1058_0, i_10_246_1083_0,
    i_10_246_1084_0, i_10_246_1223_0, i_10_246_1291_0, i_10_246_1308_0,
    i_10_246_1382_0, i_10_246_1385_0, i_10_246_1579_0, i_10_246_1580_0,
    i_10_246_1651_0, i_10_246_1655_0, i_10_246_1736_0, i_10_246_1816_0,
    i_10_246_1818_0, i_10_246_1822_0, i_10_246_1823_0, i_10_246_1913_0,
    i_10_246_1961_0, i_10_246_2024_0, i_10_246_2086_0, i_10_246_2264_0,
    i_10_246_2384_0, i_10_246_2452_0, i_10_246_2453_0, i_10_246_2474_0,
    i_10_246_2609_0, i_10_246_2617_0, i_10_246_2657_0, i_10_246_2658_0,
    i_10_246_2700_0, i_10_246_2707_0, i_10_246_2715_0, i_10_246_2786_0,
    i_10_246_2788_0, i_10_246_2789_0, i_10_246_2824_0, i_10_246_2825_0,
    i_10_246_2959_0, i_10_246_2995_0, i_10_246_3094_0, i_10_246_3167_0,
    i_10_246_3238_0, i_10_246_3239_0, i_10_246_3269_0, i_10_246_3280_0,
    i_10_246_3281_0, i_10_246_3419_0, i_10_246_3434_0, i_10_246_3473_0,
    i_10_246_3505_0, i_10_246_3508_0, i_10_246_3526_0, i_10_246_3527_0,
    i_10_246_3587_0, i_10_246_3647_0, i_10_246_3848_0, i_10_246_3883_0,
    i_10_246_3913_0, i_10_246_3914_0, i_10_246_3950_0, i_10_246_3985_0,
    i_10_246_3991_0, i_10_246_3992_0, i_10_246_4004_0, i_10_246_4057_0,
    i_10_246_4113_0, i_10_246_4118_0, i_10_246_4120_0, i_10_246_4130_0,
    i_10_246_4168_0, i_10_246_4172_0, i_10_246_4174_0, i_10_246_4276_0,
    i_10_246_4279_0, i_10_246_4281_0, i_10_246_4454_0, i_10_246_4568_0;
  output o_10_246_0_0;
  assign o_10_246_0_0 = 0;
endmodule



// Benchmark "kernel_10_247" written by ABC on Sun Jul 19 10:25:16 2020

module kernel_10_247 ( 
    i_10_247_123_0, i_10_247_181_0, i_10_247_183_0, i_10_247_319_0,
    i_10_247_320_0, i_10_247_323_0, i_10_247_328_0, i_10_247_330_0,
    i_10_247_390_0, i_10_247_391_0, i_10_247_408_0, i_10_247_437_0,
    i_10_247_442_0, i_10_247_449_0, i_10_247_755_0, i_10_247_850_0,
    i_10_247_965_0, i_10_247_998_0, i_10_247_1031_0, i_10_247_1048_0,
    i_10_247_1240_0, i_10_247_1241_0, i_10_247_1264_0, i_10_247_1265_0,
    i_10_247_1268_0, i_10_247_1310_0, i_10_247_1345_0, i_10_247_1362_0,
    i_10_247_1363_0, i_10_247_1464_0, i_10_247_1555_0, i_10_247_1651_0,
    i_10_247_1653_0, i_10_247_1684_0, i_10_247_1687_0, i_10_247_1878_0,
    i_10_247_1915_0, i_10_247_1983_0, i_10_247_2056_0, i_10_247_2183_0,
    i_10_247_2200_0, i_10_247_2361_0, i_10_247_2464_0, i_10_247_2466_0,
    i_10_247_2471_0, i_10_247_2474_0, i_10_247_2505_0, i_10_247_2508_0,
    i_10_247_2509_0, i_10_247_2515_0, i_10_247_2632_0, i_10_247_2634_0,
    i_10_247_2635_0, i_10_247_2636_0, i_10_247_2655_0, i_10_247_2661_0,
    i_10_247_2679_0, i_10_247_2681_0, i_10_247_2705_0, i_10_247_2706_0,
    i_10_247_2711_0, i_10_247_2716_0, i_10_247_2718_0, i_10_247_2719_0,
    i_10_247_2728_0, i_10_247_2734_0, i_10_247_2787_0, i_10_247_2826_0,
    i_10_247_2833_0, i_10_247_2886_0, i_10_247_2923_0, i_10_247_3036_0,
    i_10_247_3074_0, i_10_247_3075_0, i_10_247_3076_0, i_10_247_3077_0,
    i_10_247_3165_0, i_10_247_3280_0, i_10_247_3283_0, i_10_247_3315_0,
    i_10_247_3385_0, i_10_247_3388_0, i_10_247_3617_0, i_10_247_3808_0,
    i_10_247_3848_0, i_10_247_3860_0, i_10_247_3892_0, i_10_247_3894_0,
    i_10_247_3982_0, i_10_247_4118_0, i_10_247_4119_0, i_10_247_4130_0,
    i_10_247_4219_0, i_10_247_4261_0, i_10_247_4279_0, i_10_247_4289_0,
    i_10_247_4566_0, i_10_247_4585_0, i_10_247_4586_0, i_10_247_4598_0,
    o_10_247_0_0  );
  input  i_10_247_123_0, i_10_247_181_0, i_10_247_183_0, i_10_247_319_0,
    i_10_247_320_0, i_10_247_323_0, i_10_247_328_0, i_10_247_330_0,
    i_10_247_390_0, i_10_247_391_0, i_10_247_408_0, i_10_247_437_0,
    i_10_247_442_0, i_10_247_449_0, i_10_247_755_0, i_10_247_850_0,
    i_10_247_965_0, i_10_247_998_0, i_10_247_1031_0, i_10_247_1048_0,
    i_10_247_1240_0, i_10_247_1241_0, i_10_247_1264_0, i_10_247_1265_0,
    i_10_247_1268_0, i_10_247_1310_0, i_10_247_1345_0, i_10_247_1362_0,
    i_10_247_1363_0, i_10_247_1464_0, i_10_247_1555_0, i_10_247_1651_0,
    i_10_247_1653_0, i_10_247_1684_0, i_10_247_1687_0, i_10_247_1878_0,
    i_10_247_1915_0, i_10_247_1983_0, i_10_247_2056_0, i_10_247_2183_0,
    i_10_247_2200_0, i_10_247_2361_0, i_10_247_2464_0, i_10_247_2466_0,
    i_10_247_2471_0, i_10_247_2474_0, i_10_247_2505_0, i_10_247_2508_0,
    i_10_247_2509_0, i_10_247_2515_0, i_10_247_2632_0, i_10_247_2634_0,
    i_10_247_2635_0, i_10_247_2636_0, i_10_247_2655_0, i_10_247_2661_0,
    i_10_247_2679_0, i_10_247_2681_0, i_10_247_2705_0, i_10_247_2706_0,
    i_10_247_2711_0, i_10_247_2716_0, i_10_247_2718_0, i_10_247_2719_0,
    i_10_247_2728_0, i_10_247_2734_0, i_10_247_2787_0, i_10_247_2826_0,
    i_10_247_2833_0, i_10_247_2886_0, i_10_247_2923_0, i_10_247_3036_0,
    i_10_247_3074_0, i_10_247_3075_0, i_10_247_3076_0, i_10_247_3077_0,
    i_10_247_3165_0, i_10_247_3280_0, i_10_247_3283_0, i_10_247_3315_0,
    i_10_247_3385_0, i_10_247_3388_0, i_10_247_3617_0, i_10_247_3808_0,
    i_10_247_3848_0, i_10_247_3860_0, i_10_247_3892_0, i_10_247_3894_0,
    i_10_247_3982_0, i_10_247_4118_0, i_10_247_4119_0, i_10_247_4130_0,
    i_10_247_4219_0, i_10_247_4261_0, i_10_247_4279_0, i_10_247_4289_0,
    i_10_247_4566_0, i_10_247_4585_0, i_10_247_4586_0, i_10_247_4598_0;
  output o_10_247_0_0;
  assign o_10_247_0_0 = 0;
endmodule



// Benchmark "kernel_10_248" written by ABC on Sun Jul 19 10:25:16 2020

module kernel_10_248 ( 
    i_10_248_123_0, i_10_248_124_0, i_10_248_149_0, i_10_248_220_0,
    i_10_248_245_0, i_10_248_265_0, i_10_248_282_0, i_10_248_286_0,
    i_10_248_326_0, i_10_248_329_0, i_10_248_447_0, i_10_248_448_0,
    i_10_248_449_0, i_10_248_459_0, i_10_248_467_0, i_10_248_515_0,
    i_10_248_518_0, i_10_248_599_0, i_10_248_713_0, i_10_248_715_0,
    i_10_248_716_0, i_10_248_751_0, i_10_248_755_0, i_10_248_796_0,
    i_10_248_964_0, i_10_248_965_0, i_10_248_1004_0, i_10_248_1239_0,
    i_10_248_1266_0, i_10_248_1384_0, i_10_248_1583_0, i_10_248_1634_0,
    i_10_248_1726_0, i_10_248_1764_0, i_10_248_1822_0, i_10_248_1916_0,
    i_10_248_1945_0, i_10_248_1991_0, i_10_248_2255_0, i_10_248_2349_0,
    i_10_248_2353_0, i_10_248_2354_0, i_10_248_2377_0, i_10_248_2378_0,
    i_10_248_2453_0, i_10_248_2455_0, i_10_248_2469_0, i_10_248_2471_0,
    i_10_248_2504_0, i_10_248_2512_0, i_10_248_2605_0, i_10_248_2606_0,
    i_10_248_2633_0, i_10_248_2657_0, i_10_248_2663_0, i_10_248_2710_0,
    i_10_248_2714_0, i_10_248_2728_0, i_10_248_2729_0, i_10_248_2818_0,
    i_10_248_2918_0, i_10_248_2920_0, i_10_248_2980_0, i_10_248_2982_0,
    i_10_248_3043_0, i_10_248_3044_0, i_10_248_3047_0, i_10_248_3070_0,
    i_10_248_3275_0, i_10_248_3279_0, i_10_248_3391_0, i_10_248_3467_0,
    i_10_248_3473_0, i_10_248_3589_0, i_10_248_3590_0, i_10_248_3609_0,
    i_10_248_3649_0, i_10_248_3650_0, i_10_248_3652_0, i_10_248_3653_0,
    i_10_248_3781_0, i_10_248_3786_0, i_10_248_3809_0, i_10_248_3835_0,
    i_10_248_3842_0, i_10_248_3845_0, i_10_248_3854_0, i_10_248_3875_0,
    i_10_248_3947_0, i_10_248_4115_0, i_10_248_4117_0, i_10_248_4119_0,
    i_10_248_4121_0, i_10_248_4124_0, i_10_248_4214_0, i_10_248_4269_0,
    i_10_248_4285_0, i_10_248_4287_0, i_10_248_4460_0, i_10_248_4569_0,
    o_10_248_0_0  );
  input  i_10_248_123_0, i_10_248_124_0, i_10_248_149_0, i_10_248_220_0,
    i_10_248_245_0, i_10_248_265_0, i_10_248_282_0, i_10_248_286_0,
    i_10_248_326_0, i_10_248_329_0, i_10_248_447_0, i_10_248_448_0,
    i_10_248_449_0, i_10_248_459_0, i_10_248_467_0, i_10_248_515_0,
    i_10_248_518_0, i_10_248_599_0, i_10_248_713_0, i_10_248_715_0,
    i_10_248_716_0, i_10_248_751_0, i_10_248_755_0, i_10_248_796_0,
    i_10_248_964_0, i_10_248_965_0, i_10_248_1004_0, i_10_248_1239_0,
    i_10_248_1266_0, i_10_248_1384_0, i_10_248_1583_0, i_10_248_1634_0,
    i_10_248_1726_0, i_10_248_1764_0, i_10_248_1822_0, i_10_248_1916_0,
    i_10_248_1945_0, i_10_248_1991_0, i_10_248_2255_0, i_10_248_2349_0,
    i_10_248_2353_0, i_10_248_2354_0, i_10_248_2377_0, i_10_248_2378_0,
    i_10_248_2453_0, i_10_248_2455_0, i_10_248_2469_0, i_10_248_2471_0,
    i_10_248_2504_0, i_10_248_2512_0, i_10_248_2605_0, i_10_248_2606_0,
    i_10_248_2633_0, i_10_248_2657_0, i_10_248_2663_0, i_10_248_2710_0,
    i_10_248_2714_0, i_10_248_2728_0, i_10_248_2729_0, i_10_248_2818_0,
    i_10_248_2918_0, i_10_248_2920_0, i_10_248_2980_0, i_10_248_2982_0,
    i_10_248_3043_0, i_10_248_3044_0, i_10_248_3047_0, i_10_248_3070_0,
    i_10_248_3275_0, i_10_248_3279_0, i_10_248_3391_0, i_10_248_3467_0,
    i_10_248_3473_0, i_10_248_3589_0, i_10_248_3590_0, i_10_248_3609_0,
    i_10_248_3649_0, i_10_248_3650_0, i_10_248_3652_0, i_10_248_3653_0,
    i_10_248_3781_0, i_10_248_3786_0, i_10_248_3809_0, i_10_248_3835_0,
    i_10_248_3842_0, i_10_248_3845_0, i_10_248_3854_0, i_10_248_3875_0,
    i_10_248_3947_0, i_10_248_4115_0, i_10_248_4117_0, i_10_248_4119_0,
    i_10_248_4121_0, i_10_248_4124_0, i_10_248_4214_0, i_10_248_4269_0,
    i_10_248_4285_0, i_10_248_4287_0, i_10_248_4460_0, i_10_248_4569_0;
  output o_10_248_0_0;
  assign o_10_248_0_0 = 0;
endmodule



// Benchmark "kernel_10_249" written by ABC on Sun Jul 19 10:25:18 2020

module kernel_10_249 ( 
    i_10_249_221_0, i_10_249_280_0, i_10_249_282_0, i_10_249_283_0,
    i_10_249_284_0, i_10_249_286_0, i_10_249_287_0, i_10_249_433_0,
    i_10_249_435_0, i_10_249_436_0, i_10_249_441_0, i_10_249_442_0,
    i_10_249_445_0, i_10_249_446_0, i_10_249_448_0, i_10_249_466_0,
    i_10_249_507_0, i_10_249_510_0, i_10_249_755_0, i_10_249_793_0,
    i_10_249_794_0, i_10_249_798_0, i_10_249_902_0, i_10_249_957_0,
    i_10_249_958_0, i_10_249_961_0, i_10_249_1032_0, i_10_249_1033_0,
    i_10_249_1237_0, i_10_249_1240_0, i_10_249_1241_0, i_10_249_1365_0,
    i_10_249_1366_0, i_10_249_1545_0, i_10_249_1578_0, i_10_249_1648_0,
    i_10_249_1649_0, i_10_249_1650_0, i_10_249_1651_0, i_10_249_1654_0,
    i_10_249_1686_0, i_10_249_1687_0, i_10_249_1689_0, i_10_249_1819_0,
    i_10_249_1824_0, i_10_249_1825_0, i_10_249_1909_0, i_10_249_1915_0,
    i_10_249_1990_0, i_10_249_2312_0, i_10_249_2338_0, i_10_249_2354_0,
    i_10_249_2366_0, i_10_249_2380_0, i_10_249_2382_0, i_10_249_2454_0,
    i_10_249_2457_0, i_10_249_2460_0, i_10_249_2461_0, i_10_249_2662_0,
    i_10_249_2679_0, i_10_249_2703_0, i_10_249_2704_0, i_10_249_2706_0,
    i_10_249_2707_0, i_10_249_2708_0, i_10_249_2719_0, i_10_249_2731_0,
    i_10_249_2783_0, i_10_249_2827_0, i_10_249_2830_0, i_10_249_2831_0,
    i_10_249_2832_0, i_10_249_2833_0, i_10_249_2919_0, i_10_249_2923_0,
    i_10_249_3038_0, i_10_249_3158_0, i_10_249_3271_0, i_10_249_3387_0,
    i_10_249_3388_0, i_10_249_3389_0, i_10_249_3391_0, i_10_249_3392_0,
    i_10_249_3406_0, i_10_249_3472_0, i_10_249_3588_0, i_10_249_3616_0,
    i_10_249_3783_0, i_10_249_3786_0, i_10_249_3787_0, i_10_249_3838_0,
    i_10_249_3840_0, i_10_249_3841_0, i_10_249_3847_0, i_10_249_3855_0,
    i_10_249_3860_0, i_10_249_4118_0, i_10_249_4121_0, i_10_249_4274_0,
    o_10_249_0_0  );
  input  i_10_249_221_0, i_10_249_280_0, i_10_249_282_0, i_10_249_283_0,
    i_10_249_284_0, i_10_249_286_0, i_10_249_287_0, i_10_249_433_0,
    i_10_249_435_0, i_10_249_436_0, i_10_249_441_0, i_10_249_442_0,
    i_10_249_445_0, i_10_249_446_0, i_10_249_448_0, i_10_249_466_0,
    i_10_249_507_0, i_10_249_510_0, i_10_249_755_0, i_10_249_793_0,
    i_10_249_794_0, i_10_249_798_0, i_10_249_902_0, i_10_249_957_0,
    i_10_249_958_0, i_10_249_961_0, i_10_249_1032_0, i_10_249_1033_0,
    i_10_249_1237_0, i_10_249_1240_0, i_10_249_1241_0, i_10_249_1365_0,
    i_10_249_1366_0, i_10_249_1545_0, i_10_249_1578_0, i_10_249_1648_0,
    i_10_249_1649_0, i_10_249_1650_0, i_10_249_1651_0, i_10_249_1654_0,
    i_10_249_1686_0, i_10_249_1687_0, i_10_249_1689_0, i_10_249_1819_0,
    i_10_249_1824_0, i_10_249_1825_0, i_10_249_1909_0, i_10_249_1915_0,
    i_10_249_1990_0, i_10_249_2312_0, i_10_249_2338_0, i_10_249_2354_0,
    i_10_249_2366_0, i_10_249_2380_0, i_10_249_2382_0, i_10_249_2454_0,
    i_10_249_2457_0, i_10_249_2460_0, i_10_249_2461_0, i_10_249_2662_0,
    i_10_249_2679_0, i_10_249_2703_0, i_10_249_2704_0, i_10_249_2706_0,
    i_10_249_2707_0, i_10_249_2708_0, i_10_249_2719_0, i_10_249_2731_0,
    i_10_249_2783_0, i_10_249_2827_0, i_10_249_2830_0, i_10_249_2831_0,
    i_10_249_2832_0, i_10_249_2833_0, i_10_249_2919_0, i_10_249_2923_0,
    i_10_249_3038_0, i_10_249_3158_0, i_10_249_3271_0, i_10_249_3387_0,
    i_10_249_3388_0, i_10_249_3389_0, i_10_249_3391_0, i_10_249_3392_0,
    i_10_249_3406_0, i_10_249_3472_0, i_10_249_3588_0, i_10_249_3616_0,
    i_10_249_3783_0, i_10_249_3786_0, i_10_249_3787_0, i_10_249_3838_0,
    i_10_249_3840_0, i_10_249_3841_0, i_10_249_3847_0, i_10_249_3855_0,
    i_10_249_3860_0, i_10_249_4118_0, i_10_249_4121_0, i_10_249_4274_0;
  output o_10_249_0_0;
  assign o_10_249_0_0 = ~((~i_10_249_283_0 & ((~i_10_249_282_0 & ~i_10_249_958_0 & ~i_10_249_3389_0 & ~i_10_249_3783_0) | (i_10_249_282_0 & ~i_10_249_2457_0 & ~i_10_249_3786_0))) | (i_10_249_442_0 & ((i_10_249_441_0 & ~i_10_249_957_0 & ~i_10_249_1990_0) | (i_10_249_436_0 & ~i_10_249_958_0 & ~i_10_249_1824_0 & ~i_10_249_3787_0))) | (~i_10_249_436_0 & ((~i_10_249_442_0 & ((~i_10_249_280_0 & ~i_10_249_755_0 & ~i_10_249_958_0 & ~i_10_249_2366_0 & ~i_10_249_2460_0 & ~i_10_249_2832_0 & ~i_10_249_3406_0) | (~i_10_249_448_0 & ~i_10_249_2312_0 & ~i_10_249_2461_0 & ~i_10_249_2831_0 & ~i_10_249_3838_0 & ~i_10_249_3847_0 & ~i_10_249_3855_0))) | (~i_10_249_798_0 & ~i_10_249_961_0 & i_10_249_1687_0 & ~i_10_249_2354_0 & ~i_10_249_2380_0 & ~i_10_249_2827_0))) | (~i_10_249_961_0 & ((i_10_249_1240_0 & i_10_249_3392_0 & i_10_249_3588_0) | (~i_10_249_1032_0 & ~i_10_249_1689_0 & i_10_249_2704_0 & ~i_10_249_3392_0 & ~i_10_249_3787_0))) | (~i_10_249_1237_0 & ((~i_10_249_284_0 & ~i_10_249_1032_0 & ~i_10_249_1686_0 & ~i_10_249_2312_0 & ~i_10_249_2366_0 & ~i_10_249_2380_0 & ~i_10_249_2460_0 & ~i_10_249_2461_0 & ~i_10_249_2708_0 & ~i_10_249_2719_0) | (i_10_249_284_0 & i_10_249_1825_0 & ~i_10_249_2731_0 & ~i_10_249_3387_0 & ~i_10_249_3847_0))) | (i_10_249_1648_0 & (i_10_249_1237_0 | (~i_10_249_435_0 & ~i_10_249_1545_0 & ~i_10_249_1689_0 & ~i_10_249_1990_0 & ~i_10_249_3038_0))) | (~i_10_249_958_0 & ((~i_10_249_435_0 & ((~i_10_249_284_0 & ~i_10_249_2312_0 & ~i_10_249_2457_0 & ~i_10_249_3847_0) | (i_10_249_1237_0 & ~i_10_249_1654_0 & ~i_10_249_2461_0 & ~i_10_249_2827_0 & ~i_10_249_3786_0 & ~i_10_249_4118_0))) | (~i_10_249_2380_0 & ~i_10_249_2461_0 & ~i_10_249_2662_0 & ~i_10_249_2731_0 & ~i_10_249_2783_0 & ~i_10_249_2831_0 & ~i_10_249_2919_0 & ~i_10_249_3038_0 & ~i_10_249_3271_0 & i_10_249_3388_0 & ~i_10_249_3855_0))) | (~i_10_249_2312_0 & ((~i_10_249_284_0 & ((i_10_249_2354_0 & ~i_10_249_2461_0 & ~i_10_249_2831_0) | (i_10_249_286_0 & ~i_10_249_1825_0 & ~i_10_249_3841_0))) | (~i_10_249_2783_0 & ((~i_10_249_282_0 & ~i_10_249_1990_0 & ~i_10_249_2460_0 & ~i_10_249_2833_0 & ~i_10_249_3038_0 & ~i_10_249_3783_0 & ~i_10_249_3838_0 & ~i_10_249_3855_0 & ~i_10_249_4118_0) | (i_10_249_1819_0 & ~i_10_249_3847_0 & ~i_10_249_4121_0))) | (i_10_249_445_0 & ~i_10_249_2719_0 & ~i_10_249_2731_0 & ~i_10_249_3038_0))) | (~i_10_249_3388_0 & ((~i_10_249_282_0 & ((~i_10_249_433_0 & ~i_10_249_1033_0 & ~i_10_249_2461_0 & ~i_10_249_3389_0 & ~i_10_249_3391_0) | (i_10_249_283_0 & i_10_249_3855_0))) | (i_10_249_1687_0 & ~i_10_249_3391_0 & ~i_10_249_3855_0))) | (~i_10_249_1033_0 & ((i_10_249_1240_0 & ~i_10_249_1648_0 & ~i_10_249_3389_0) | (~i_10_249_448_0 & i_10_249_1241_0 & ~i_10_249_2366_0 & ~i_10_249_2783_0 & ~i_10_249_4121_0))) | (~i_10_249_2461_0 & ((i_10_249_1687_0 & ((i_10_249_2731_0 & ~i_10_249_2831_0) | (~i_10_249_1578_0 & ~i_10_249_2380_0 & ~i_10_249_2783_0 & ~i_10_249_4274_0))) | (~i_10_249_433_0 & ~i_10_249_957_0 & ~i_10_249_2783_0 & i_10_249_3841_0) | (i_10_249_2460_0 & i_10_249_2833_0 & ~i_10_249_3847_0))) | (~i_10_249_433_0 & ((i_10_249_793_0 & ~i_10_249_2460_0) | (~i_10_249_957_0 & i_10_249_1237_0 & ~i_10_249_1687_0 & ~i_10_249_3406_0))) | (~i_10_249_4118_0 & ((~i_10_249_957_0 & i_10_249_1650_0 & ~i_10_249_3389_0) | (i_10_249_2366_0 & ~i_10_249_2731_0 & i_10_249_4121_0))) | (~i_10_249_2366_0 & i_10_249_2923_0 & i_10_249_3616_0 & i_10_249_3841_0));
endmodule



// Benchmark "kernel_10_250" written by ABC on Sun Jul 19 10:25:19 2020

module kernel_10_250 ( 
    i_10_250_157_0, i_10_250_174_0, i_10_250_248_0, i_10_250_273_0,
    i_10_250_274_0, i_10_250_277_0, i_10_250_285_0, i_10_250_286_0,
    i_10_250_324_0, i_10_250_428_0, i_10_250_436_0, i_10_250_439_0,
    i_10_250_467_0, i_10_250_793_0, i_10_250_796_0, i_10_250_959_0,
    i_10_250_967_0, i_10_250_968_0, i_10_250_995_0, i_10_250_999_0,
    i_10_250_1027_0, i_10_250_1033_0, i_10_250_1217_0, i_10_250_1241_0,
    i_10_250_1245_0, i_10_250_1250_0, i_10_250_1306_0, i_10_250_1309_0,
    i_10_250_1310_0, i_10_250_1313_0, i_10_250_1432_0, i_10_250_1444_0,
    i_10_250_1647_0, i_10_250_1649_0, i_10_250_1945_0, i_10_250_1949_0,
    i_10_250_1950_0, i_10_250_2019_0, i_10_250_2308_0, i_10_250_2327_0,
    i_10_250_2350_0, i_10_250_2452_0, i_10_250_2471_0, i_10_250_2508_0,
    i_10_250_2509_0, i_10_250_2541_0, i_10_250_2542_0, i_10_250_2628_0,
    i_10_250_2629_0, i_10_250_2630_0, i_10_250_2633_0, i_10_250_2635_0,
    i_10_250_2657_0, i_10_250_2663_0, i_10_250_2713_0, i_10_250_2734_0,
    i_10_250_2735_0, i_10_250_2785_0, i_10_250_2828_0, i_10_250_2830_0,
    i_10_250_2920_0, i_10_250_3033_0, i_10_250_3037_0, i_10_250_3038_0,
    i_10_250_3092_0, i_10_250_3268_0, i_10_250_3271_0, i_10_250_3281_0,
    i_10_250_3384_0, i_10_250_3385_0, i_10_250_3388_0, i_10_250_3433_0,
    i_10_250_3465_0, i_10_250_3472_0, i_10_250_3586_0, i_10_250_3587_0,
    i_10_250_3613_0, i_10_250_3614_0, i_10_250_3616_0, i_10_250_3626_0,
    i_10_250_3646_0, i_10_250_3647_0, i_10_250_3649_0, i_10_250_3650_0,
    i_10_250_3836_0, i_10_250_3838_0, i_10_250_3839_0, i_10_250_3846_0,
    i_10_250_3847_0, i_10_250_3848_0, i_10_250_3857_0, i_10_250_3890_0,
    i_10_250_3980_0, i_10_250_3988_0, i_10_250_3994_0, i_10_250_4055_0,
    i_10_250_4114_0, i_10_250_4116_0, i_10_250_4118_0, i_10_250_4284_0,
    o_10_250_0_0  );
  input  i_10_250_157_0, i_10_250_174_0, i_10_250_248_0, i_10_250_273_0,
    i_10_250_274_0, i_10_250_277_0, i_10_250_285_0, i_10_250_286_0,
    i_10_250_324_0, i_10_250_428_0, i_10_250_436_0, i_10_250_439_0,
    i_10_250_467_0, i_10_250_793_0, i_10_250_796_0, i_10_250_959_0,
    i_10_250_967_0, i_10_250_968_0, i_10_250_995_0, i_10_250_999_0,
    i_10_250_1027_0, i_10_250_1033_0, i_10_250_1217_0, i_10_250_1241_0,
    i_10_250_1245_0, i_10_250_1250_0, i_10_250_1306_0, i_10_250_1309_0,
    i_10_250_1310_0, i_10_250_1313_0, i_10_250_1432_0, i_10_250_1444_0,
    i_10_250_1647_0, i_10_250_1649_0, i_10_250_1945_0, i_10_250_1949_0,
    i_10_250_1950_0, i_10_250_2019_0, i_10_250_2308_0, i_10_250_2327_0,
    i_10_250_2350_0, i_10_250_2452_0, i_10_250_2471_0, i_10_250_2508_0,
    i_10_250_2509_0, i_10_250_2541_0, i_10_250_2542_0, i_10_250_2628_0,
    i_10_250_2629_0, i_10_250_2630_0, i_10_250_2633_0, i_10_250_2635_0,
    i_10_250_2657_0, i_10_250_2663_0, i_10_250_2713_0, i_10_250_2734_0,
    i_10_250_2735_0, i_10_250_2785_0, i_10_250_2828_0, i_10_250_2830_0,
    i_10_250_2920_0, i_10_250_3033_0, i_10_250_3037_0, i_10_250_3038_0,
    i_10_250_3092_0, i_10_250_3268_0, i_10_250_3271_0, i_10_250_3281_0,
    i_10_250_3384_0, i_10_250_3385_0, i_10_250_3388_0, i_10_250_3433_0,
    i_10_250_3465_0, i_10_250_3472_0, i_10_250_3586_0, i_10_250_3587_0,
    i_10_250_3613_0, i_10_250_3614_0, i_10_250_3616_0, i_10_250_3626_0,
    i_10_250_3646_0, i_10_250_3647_0, i_10_250_3649_0, i_10_250_3650_0,
    i_10_250_3836_0, i_10_250_3838_0, i_10_250_3839_0, i_10_250_3846_0,
    i_10_250_3847_0, i_10_250_3848_0, i_10_250_3857_0, i_10_250_3890_0,
    i_10_250_3980_0, i_10_250_3988_0, i_10_250_3994_0, i_10_250_4055_0,
    i_10_250_4114_0, i_10_250_4116_0, i_10_250_4118_0, i_10_250_4284_0;
  output o_10_250_0_0;
  assign o_10_250_0_0 = 0;
endmodule



// Benchmark "kernel_10_251" written by ABC on Sun Jul 19 10:25:20 2020

module kernel_10_251 ( 
    i_10_251_124_0, i_10_251_222_0, i_10_251_246_0, i_10_251_247_0,
    i_10_251_249_0, i_10_251_250_0, i_10_251_280_0, i_10_251_315_0,
    i_10_251_317_0, i_10_251_327_0, i_10_251_329_0, i_10_251_331_0,
    i_10_251_395_0, i_10_251_406_0, i_10_251_409_0, i_10_251_751_0,
    i_10_251_797_0, i_10_251_955_0, i_10_251_956_0, i_10_251_993_0,
    i_10_251_1040_0, i_10_251_1129_0, i_10_251_1234_0, i_10_251_1235_0,
    i_10_251_1238_0, i_10_251_1241_0, i_10_251_1244_0, i_10_251_1246_0,
    i_10_251_1264_0, i_10_251_1309_0, i_10_251_1341_0, i_10_251_1363_0,
    i_10_251_1579_0, i_10_251_1600_0, i_10_251_1651_0, i_10_251_1686_0,
    i_10_251_1689_0, i_10_251_1819_0, i_10_251_1824_0, i_10_251_1950_0,
    i_10_251_2182_0, i_10_251_2203_0, i_10_251_2350_0, i_10_251_2353_0,
    i_10_251_2354_0, i_10_251_2356_0, i_10_251_2357_0, i_10_251_2361_0,
    i_10_251_2364_0, i_10_251_2365_0, i_10_251_2366_0, i_10_251_2454_0,
    i_10_251_2455_0, i_10_251_2456_0, i_10_251_2461_0, i_10_251_2721_0,
    i_10_251_2722_0, i_10_251_2723_0, i_10_251_2725_0, i_10_251_2728_0,
    i_10_251_2885_0, i_10_251_2888_0, i_10_251_2916_0, i_10_251_2922_0,
    i_10_251_2923_0, i_10_251_3034_0, i_10_251_3038_0, i_10_251_3043_0,
    i_10_251_3202_0, i_10_251_3203_0, i_10_251_3275_0, i_10_251_3281_0,
    i_10_251_3284_0, i_10_251_3386_0, i_10_251_3389_0, i_10_251_3392_0,
    i_10_251_3542_0, i_10_251_3586_0, i_10_251_3589_0, i_10_251_3616_0,
    i_10_251_3617_0, i_10_251_3653_0, i_10_251_3780_0, i_10_251_3781_0,
    i_10_251_3785_0, i_10_251_3788_0, i_10_251_3808_0, i_10_251_3814_0,
    i_10_251_3844_0, i_10_251_3845_0, i_10_251_3848_0, i_10_251_3858_0,
    i_10_251_3914_0, i_10_251_3983_0, i_10_251_4117_0, i_10_251_4120_0,
    i_10_251_4286_0, i_10_251_4288_0, i_10_251_4289_0, i_10_251_4563_0,
    o_10_251_0_0  );
  input  i_10_251_124_0, i_10_251_222_0, i_10_251_246_0, i_10_251_247_0,
    i_10_251_249_0, i_10_251_250_0, i_10_251_280_0, i_10_251_315_0,
    i_10_251_317_0, i_10_251_327_0, i_10_251_329_0, i_10_251_331_0,
    i_10_251_395_0, i_10_251_406_0, i_10_251_409_0, i_10_251_751_0,
    i_10_251_797_0, i_10_251_955_0, i_10_251_956_0, i_10_251_993_0,
    i_10_251_1040_0, i_10_251_1129_0, i_10_251_1234_0, i_10_251_1235_0,
    i_10_251_1238_0, i_10_251_1241_0, i_10_251_1244_0, i_10_251_1246_0,
    i_10_251_1264_0, i_10_251_1309_0, i_10_251_1341_0, i_10_251_1363_0,
    i_10_251_1579_0, i_10_251_1600_0, i_10_251_1651_0, i_10_251_1686_0,
    i_10_251_1689_0, i_10_251_1819_0, i_10_251_1824_0, i_10_251_1950_0,
    i_10_251_2182_0, i_10_251_2203_0, i_10_251_2350_0, i_10_251_2353_0,
    i_10_251_2354_0, i_10_251_2356_0, i_10_251_2357_0, i_10_251_2361_0,
    i_10_251_2364_0, i_10_251_2365_0, i_10_251_2366_0, i_10_251_2454_0,
    i_10_251_2455_0, i_10_251_2456_0, i_10_251_2461_0, i_10_251_2721_0,
    i_10_251_2722_0, i_10_251_2723_0, i_10_251_2725_0, i_10_251_2728_0,
    i_10_251_2885_0, i_10_251_2888_0, i_10_251_2916_0, i_10_251_2922_0,
    i_10_251_2923_0, i_10_251_3034_0, i_10_251_3038_0, i_10_251_3043_0,
    i_10_251_3202_0, i_10_251_3203_0, i_10_251_3275_0, i_10_251_3281_0,
    i_10_251_3284_0, i_10_251_3386_0, i_10_251_3389_0, i_10_251_3392_0,
    i_10_251_3542_0, i_10_251_3586_0, i_10_251_3589_0, i_10_251_3616_0,
    i_10_251_3617_0, i_10_251_3653_0, i_10_251_3780_0, i_10_251_3781_0,
    i_10_251_3785_0, i_10_251_3788_0, i_10_251_3808_0, i_10_251_3814_0,
    i_10_251_3844_0, i_10_251_3845_0, i_10_251_3848_0, i_10_251_3858_0,
    i_10_251_3914_0, i_10_251_3983_0, i_10_251_4117_0, i_10_251_4120_0,
    i_10_251_4286_0, i_10_251_4288_0, i_10_251_4289_0, i_10_251_4563_0;
  output o_10_251_0_0;
  assign o_10_251_0_0 = 0;
endmodule



// Benchmark "kernel_10_252" written by ABC on Sun Jul 19 10:25:21 2020

module kernel_10_252 ( 
    i_10_252_150_0, i_10_252_175_0, i_10_252_183_0, i_10_252_219_0,
    i_10_252_220_0, i_10_252_224_0, i_10_252_260_0, i_10_252_281_0,
    i_10_252_286_0, i_10_252_319_0, i_10_252_320_0, i_10_252_409_0,
    i_10_252_432_0, i_10_252_435_0, i_10_252_436_0, i_10_252_441_0,
    i_10_252_444_0, i_10_252_445_0, i_10_252_448_0, i_10_252_461_0,
    i_10_252_462_0, i_10_252_519_0, i_10_252_697_0, i_10_252_795_0,
    i_10_252_796_0, i_10_252_898_0, i_10_252_966_0, i_10_252_967_0,
    i_10_252_1033_0, i_10_252_1237_0, i_10_252_1238_0, i_10_252_1241_0,
    i_10_252_1243_0, i_10_252_1305_0, i_10_252_1308_0, i_10_252_1309_0,
    i_10_252_1437_0, i_10_252_1650_0, i_10_252_1651_0, i_10_252_1681_0,
    i_10_252_1682_0, i_10_252_1819_0, i_10_252_1821_0, i_10_252_1822_0,
    i_10_252_1825_0, i_10_252_2182_0, i_10_252_2331_0, i_10_252_2334_0,
    i_10_252_2382_0, i_10_252_2384_0, i_10_252_2405_0, i_10_252_2452_0,
    i_10_252_2453_0, i_10_252_2455_0, i_10_252_2631_0, i_10_252_2635_0,
    i_10_252_2658_0, i_10_252_2659_0, i_10_252_2660_0, i_10_252_2710_0,
    i_10_252_2733_0, i_10_252_2831_0, i_10_252_2919_0, i_10_252_2920_0,
    i_10_252_3036_0, i_10_252_3037_0, i_10_252_3045_0, i_10_252_3046_0,
    i_10_252_3150_0, i_10_252_3153_0, i_10_252_3165_0, i_10_252_3166_0,
    i_10_252_3270_0, i_10_252_3274_0, i_10_252_3278_0, i_10_252_3280_0,
    i_10_252_3281_0, i_10_252_3326_0, i_10_252_3469_0, i_10_252_3583_0,
    i_10_252_3649_0, i_10_252_3781_0, i_10_252_3846_0, i_10_252_3847_0,
    i_10_252_3853_0, i_10_252_3858_0, i_10_252_3912_0, i_10_252_3915_0,
    i_10_252_3980_0, i_10_252_3985_0, i_10_252_4116_0, i_10_252_4118_0,
    i_10_252_4120_0, i_10_252_4219_0, i_10_252_4269_0, i_10_252_4271_0,
    i_10_252_4283_0, i_10_252_4564_0, i_10_252_4566_0, i_10_252_4567_0,
    o_10_252_0_0  );
  input  i_10_252_150_0, i_10_252_175_0, i_10_252_183_0, i_10_252_219_0,
    i_10_252_220_0, i_10_252_224_0, i_10_252_260_0, i_10_252_281_0,
    i_10_252_286_0, i_10_252_319_0, i_10_252_320_0, i_10_252_409_0,
    i_10_252_432_0, i_10_252_435_0, i_10_252_436_0, i_10_252_441_0,
    i_10_252_444_0, i_10_252_445_0, i_10_252_448_0, i_10_252_461_0,
    i_10_252_462_0, i_10_252_519_0, i_10_252_697_0, i_10_252_795_0,
    i_10_252_796_0, i_10_252_898_0, i_10_252_966_0, i_10_252_967_0,
    i_10_252_1033_0, i_10_252_1237_0, i_10_252_1238_0, i_10_252_1241_0,
    i_10_252_1243_0, i_10_252_1305_0, i_10_252_1308_0, i_10_252_1309_0,
    i_10_252_1437_0, i_10_252_1650_0, i_10_252_1651_0, i_10_252_1681_0,
    i_10_252_1682_0, i_10_252_1819_0, i_10_252_1821_0, i_10_252_1822_0,
    i_10_252_1825_0, i_10_252_2182_0, i_10_252_2331_0, i_10_252_2334_0,
    i_10_252_2382_0, i_10_252_2384_0, i_10_252_2405_0, i_10_252_2452_0,
    i_10_252_2453_0, i_10_252_2455_0, i_10_252_2631_0, i_10_252_2635_0,
    i_10_252_2658_0, i_10_252_2659_0, i_10_252_2660_0, i_10_252_2710_0,
    i_10_252_2733_0, i_10_252_2831_0, i_10_252_2919_0, i_10_252_2920_0,
    i_10_252_3036_0, i_10_252_3037_0, i_10_252_3045_0, i_10_252_3046_0,
    i_10_252_3150_0, i_10_252_3153_0, i_10_252_3165_0, i_10_252_3166_0,
    i_10_252_3270_0, i_10_252_3274_0, i_10_252_3278_0, i_10_252_3280_0,
    i_10_252_3281_0, i_10_252_3326_0, i_10_252_3469_0, i_10_252_3583_0,
    i_10_252_3649_0, i_10_252_3781_0, i_10_252_3846_0, i_10_252_3847_0,
    i_10_252_3853_0, i_10_252_3858_0, i_10_252_3912_0, i_10_252_3915_0,
    i_10_252_3980_0, i_10_252_3985_0, i_10_252_4116_0, i_10_252_4118_0,
    i_10_252_4120_0, i_10_252_4219_0, i_10_252_4269_0, i_10_252_4271_0,
    i_10_252_4283_0, i_10_252_4564_0, i_10_252_4566_0, i_10_252_4567_0;
  output o_10_252_0_0;
  assign o_10_252_0_0 = ~((~i_10_252_432_0 & ((~i_10_252_1243_0 & ~i_10_252_2334_0 & i_10_252_3046_0 & ~i_10_252_3165_0 & i_10_252_3853_0) | (~i_10_252_409_0 & ~i_10_252_444_0 & ~i_10_252_1237_0 & ~i_10_252_1309_0 & ~i_10_252_1650_0 & ~i_10_252_2405_0 & ~i_10_252_2453_0 & ~i_10_252_2455_0 & ~i_10_252_2658_0 & ~i_10_252_3037_0 & ~i_10_252_3045_0 & ~i_10_252_3469_0 & ~i_10_252_3985_0 & ~i_10_252_4116_0 & ~i_10_252_4118_0 & ~i_10_252_4219_0))) | (~i_10_252_4566_0 & ((~i_10_252_3270_0 & ((~i_10_252_220_0 & ~i_10_252_461_0 & ((~i_10_252_2660_0 & ~i_10_252_3036_0 & ~i_10_252_3165_0 & i_10_252_3858_0 & ~i_10_252_3912_0) | (~i_10_252_519_0 & ~i_10_252_966_0 & i_10_252_1819_0 & ~i_10_252_2182_0 & ~i_10_252_4567_0))) | (~i_10_252_4567_0 & ((~i_10_252_441_0 & ~i_10_252_444_0 & ~i_10_252_967_0 & ~i_10_252_1822_0 & i_10_252_1825_0 & ~i_10_252_3165_0 & ~i_10_252_3166_0 & ~i_10_252_3858_0) | (~i_10_252_175_0 & ~i_10_252_796_0 & ~i_10_252_1033_0 & ~i_10_252_1243_0 & ~i_10_252_2453_0 & ~i_10_252_2733_0 & ~i_10_252_2831_0 & ~i_10_252_3846_0 & ~i_10_252_4564_0))))) | (~i_10_252_444_0 & ((~i_10_252_967_0 & ~i_10_252_3037_0 & ((~i_10_252_435_0 & ~i_10_252_441_0 & ~i_10_252_1033_0 & i_10_252_1819_0 & ~i_10_252_2453_0 & ~i_10_252_3846_0) | (~i_10_252_1243_0 & ~i_10_252_1650_0 & ~i_10_252_2384_0 & ~i_10_252_3165_0 & ~i_10_252_3166_0 & ~i_10_252_3847_0 & ~i_10_252_4219_0 & ~i_10_252_4269_0))) | (~i_10_252_150_0 & i_10_252_175_0 & ~i_10_252_448_0 & ~i_10_252_2384_0 & ~i_10_252_2452_0 & ~i_10_252_4219_0 & ~i_10_252_4567_0))) | (i_10_252_281_0 & ~i_10_252_697_0 & ~i_10_252_1437_0 & ~i_10_252_2635_0 & ~i_10_252_3846_0) | (i_10_252_2710_0 & i_10_252_2919_0 & i_10_252_3469_0 & ~i_10_252_3583_0) | (~i_10_252_409_0 & ~i_10_252_966_0 & i_10_252_1241_0 & ~i_10_252_2919_0 & ~i_10_252_3781_0 & ~i_10_252_3847_0))) | (~i_10_252_4120_0 & ((i_10_252_281_0 & ((~i_10_252_220_0 & ~i_10_252_1650_0 & ~i_10_252_2384_0 & ~i_10_252_2631_0 & ~i_10_252_2831_0 & ~i_10_252_3281_0) | (~i_10_252_441_0 & ~i_10_252_1825_0 & ~i_10_252_2405_0 & ~i_10_252_2919_0 & ~i_10_252_3649_0))) | (~i_10_252_1650_0 & ((~i_10_252_462_0 & ~i_10_252_967_0 & ~i_10_252_2831_0 & ~i_10_252_2920_0 & ~i_10_252_3037_0 & ~i_10_252_3274_0 & ~i_10_252_3858_0 & ~i_10_252_3980_0) | (~i_10_252_150_0 & i_10_252_1822_0 & i_10_252_3781_0 & ~i_10_252_4269_0 & ~i_10_252_4271_0 & ~i_10_252_4564_0))) | (i_10_252_1237_0 & i_10_252_1305_0 & ~i_10_252_1825_0 & ~i_10_252_2382_0 & ~i_10_252_2635_0) | (i_10_252_2659_0 & i_10_252_2660_0 & ~i_10_252_3270_0 & ~i_10_252_3469_0 & ~i_10_252_4116_0))) | (~i_10_252_150_0 & ((~i_10_252_220_0 & ((~i_10_252_444_0 & ~i_10_252_1243_0 & i_10_252_2660_0) | (~i_10_252_409_0 & ~i_10_252_519_0 & ~i_10_252_796_0 & ~i_10_252_967_0 & ~i_10_252_2182_0 & ~i_10_252_2384_0 & ~i_10_252_2455_0 & ~i_10_252_2631_0 & ~i_10_252_4269_0 & ~i_10_252_4567_0))) | (~i_10_252_2382_0 & ((~i_10_252_1033_0 & i_10_252_1308_0 & ~i_10_252_2452_0 & ~i_10_252_2635_0 & ~i_10_252_3165_0 & ~i_10_252_3781_0 & ~i_10_252_3912_0 & ~i_10_252_4564_0) | (~i_10_252_409_0 & ~i_10_252_697_0 & ~i_10_252_1308_0 & i_10_252_3278_0 & ~i_10_252_4269_0 & ~i_10_252_4567_0))) | (~i_10_252_175_0 & ~i_10_252_445_0 & ~i_10_252_519_0 & ~i_10_252_898_0 & ~i_10_252_1243_0 & ~i_10_252_1822_0 & ~i_10_252_3037_0 & ~i_10_252_3165_0 & ~i_10_252_4564_0))) | (~i_10_252_175_0 & ((~i_10_252_462_0 & ~i_10_252_519_0 & i_10_252_1305_0 & ~i_10_252_2635_0 & ~i_10_252_3037_0 & ~i_10_252_3846_0) | (~i_10_252_409_0 & ~i_10_252_967_0 & i_10_252_2659_0 & ~i_10_252_2920_0 & ~i_10_252_4269_0))) | (~i_10_252_3847_0 & ((~i_10_252_409_0 & ((i_10_252_448_0 & ~i_10_252_1309_0 & ~i_10_252_1822_0 & ~i_10_252_2182_0 & ~i_10_252_2631_0 & ~i_10_252_2831_0 & i_10_252_4271_0 & ~i_10_252_4564_0) | (~i_10_252_448_0 & ~i_10_252_795_0 & ~i_10_252_966_0 & ~i_10_252_1243_0 & ~i_10_252_2659_0 & ~i_10_252_3165_0 & ~i_10_252_3270_0 & ~i_10_252_3274_0 & ~i_10_252_4219_0 & ~i_10_252_4567_0))) | (~i_10_252_445_0 & ~i_10_252_796_0 & ~i_10_252_1821_0 & i_10_252_2659_0 & ~i_10_252_3165_0 & ~i_10_252_3166_0))) | (~i_10_252_444_0 & ((~i_10_252_519_0 & ~i_10_252_2384_0 & ~i_10_252_2631_0 & i_10_252_2831_0 & ~i_10_252_3165_0 & ~i_10_252_3281_0 & ~i_10_252_3781_0 & ~i_10_252_4219_0) | (i_10_252_2710_0 & ~i_10_252_3166_0 & i_10_252_4118_0 & ~i_10_252_4567_0))) | (~i_10_252_967_0 & ~i_10_252_2919_0 & ((~i_10_252_1243_0 & i_10_252_2710_0 & ~i_10_252_2920_0) | (~i_10_252_795_0 & ~i_10_252_898_0 & ~i_10_252_3036_0 & ~i_10_252_3166_0 & i_10_252_4118_0 & ~i_10_252_4567_0 & ~i_10_252_3469_0 & ~i_10_252_3781_0))) | (~i_10_252_1243_0 & ((~i_10_252_796_0 & ~i_10_252_1033_0 & i_10_252_1822_0 & ~i_10_252_3165_0 & i_10_252_3281_0) | (i_10_252_432_0 & ~i_10_252_445_0 & i_10_252_2710_0 & ~i_10_252_2831_0 & ~i_10_252_3270_0 & ~i_10_252_3649_0))) | (~i_10_252_2635_0 & ((i_10_252_2384_0 & i_10_252_3274_0 & ~i_10_252_3281_0) | (i_10_252_1309_0 & i_10_252_1819_0 & ~i_10_252_2453_0 & i_10_252_4116_0))) | (i_10_252_1309_0 & ((~i_10_252_1308_0 & ~i_10_252_1822_0 & ~i_10_252_2382_0 & i_10_252_2831_0) | (~i_10_252_448_0 & i_10_252_461_0 & ~i_10_252_3649_0))) | (~i_10_252_3270_0 & ((~i_10_252_2331_0 & i_10_252_2659_0 & i_10_252_2660_0 & i_10_252_3853_0) | (~i_10_252_441_0 & ~i_10_252_1651_0 & ~i_10_252_1821_0 & i_10_252_2831_0 & ~i_10_252_3036_0 & ~i_10_252_3165_0 & ~i_10_252_3274_0 & ~i_10_252_3912_0 & ~i_10_252_4271_0))) | (i_10_252_1243_0 & i_10_252_3280_0 & i_10_252_3853_0) | (i_10_252_1822_0 & ~i_10_252_3037_0 & i_10_252_3274_0 & i_10_252_3985_0));
endmodule



// Benchmark "kernel_10_253" written by ABC on Sun Jul 19 10:25:22 2020

module kernel_10_253 ( 
    i_10_253_88_0, i_10_253_148_0, i_10_253_217_0, i_10_253_269_0,
    i_10_253_408_0, i_10_253_424_0, i_10_253_434_0, i_10_253_435_0,
    i_10_253_441_0, i_10_253_442_0, i_10_253_459_0, i_10_253_533_0,
    i_10_253_559_0, i_10_253_733_0, i_10_253_794_0, i_10_253_990_0,
    i_10_253_1036_0, i_10_253_1085_0, i_10_253_1164_0, i_10_253_1222_0,
    i_10_253_1234_0, i_10_253_1241_0, i_10_253_1309_0, i_10_253_1310_0,
    i_10_253_1341_0, i_10_253_1384_0, i_10_253_1552_0, i_10_253_1579_0,
    i_10_253_1580_0, i_10_253_1582_0, i_10_253_1687_0, i_10_253_1688_0,
    i_10_253_1737_0, i_10_253_1806_0, i_10_253_1818_0, i_10_253_1819_0,
    i_10_253_2016_0, i_10_253_2206_0, i_10_253_2250_0, i_10_253_2355_0,
    i_10_253_2356_0, i_10_253_2364_0, i_10_253_2389_0, i_10_253_2451_0,
    i_10_253_2469_0, i_10_253_2470_0, i_10_253_2515_0, i_10_253_2563_0,
    i_10_253_2602_0, i_10_253_2604_0, i_10_253_2606_0, i_10_253_2628_0,
    i_10_253_2629_0, i_10_253_2701_0, i_10_253_2711_0, i_10_253_2725_0,
    i_10_253_2782_0, i_10_253_2789_0, i_10_253_2817_0, i_10_253_2820_0,
    i_10_253_2841_0, i_10_253_2862_0, i_10_253_2863_0, i_10_253_2883_0,
    i_10_253_2884_0, i_10_253_2921_0, i_10_253_3048_0, i_10_253_3124_0,
    i_10_253_3200_0, i_10_253_3268_0, i_10_253_3269_0, i_10_253_3277_0,
    i_10_253_3295_0, i_10_253_3297_0, i_10_253_3357_0, i_10_253_3384_0,
    i_10_253_3387_0, i_10_253_3388_0, i_10_253_3389_0, i_10_253_3408_0,
    i_10_253_3430_0, i_10_253_3520_0, i_10_253_3544_0, i_10_253_3610_0,
    i_10_253_3612_0, i_10_253_3640_0, i_10_253_3649_0, i_10_253_3808_0,
    i_10_253_3835_0, i_10_253_3855_0, i_10_253_3889_0, i_10_253_3920_0,
    i_10_253_3981_0, i_10_253_3991_0, i_10_253_4129_0, i_10_253_4272_0,
    i_10_253_4273_0, i_10_253_4281_0, i_10_253_4290_0, i_10_253_4292_0,
    o_10_253_0_0  );
  input  i_10_253_88_0, i_10_253_148_0, i_10_253_217_0, i_10_253_269_0,
    i_10_253_408_0, i_10_253_424_0, i_10_253_434_0, i_10_253_435_0,
    i_10_253_441_0, i_10_253_442_0, i_10_253_459_0, i_10_253_533_0,
    i_10_253_559_0, i_10_253_733_0, i_10_253_794_0, i_10_253_990_0,
    i_10_253_1036_0, i_10_253_1085_0, i_10_253_1164_0, i_10_253_1222_0,
    i_10_253_1234_0, i_10_253_1241_0, i_10_253_1309_0, i_10_253_1310_0,
    i_10_253_1341_0, i_10_253_1384_0, i_10_253_1552_0, i_10_253_1579_0,
    i_10_253_1580_0, i_10_253_1582_0, i_10_253_1687_0, i_10_253_1688_0,
    i_10_253_1737_0, i_10_253_1806_0, i_10_253_1818_0, i_10_253_1819_0,
    i_10_253_2016_0, i_10_253_2206_0, i_10_253_2250_0, i_10_253_2355_0,
    i_10_253_2356_0, i_10_253_2364_0, i_10_253_2389_0, i_10_253_2451_0,
    i_10_253_2469_0, i_10_253_2470_0, i_10_253_2515_0, i_10_253_2563_0,
    i_10_253_2602_0, i_10_253_2604_0, i_10_253_2606_0, i_10_253_2628_0,
    i_10_253_2629_0, i_10_253_2701_0, i_10_253_2711_0, i_10_253_2725_0,
    i_10_253_2782_0, i_10_253_2789_0, i_10_253_2817_0, i_10_253_2820_0,
    i_10_253_2841_0, i_10_253_2862_0, i_10_253_2863_0, i_10_253_2883_0,
    i_10_253_2884_0, i_10_253_2921_0, i_10_253_3048_0, i_10_253_3124_0,
    i_10_253_3200_0, i_10_253_3268_0, i_10_253_3269_0, i_10_253_3277_0,
    i_10_253_3295_0, i_10_253_3297_0, i_10_253_3357_0, i_10_253_3384_0,
    i_10_253_3387_0, i_10_253_3388_0, i_10_253_3389_0, i_10_253_3408_0,
    i_10_253_3430_0, i_10_253_3520_0, i_10_253_3544_0, i_10_253_3610_0,
    i_10_253_3612_0, i_10_253_3640_0, i_10_253_3649_0, i_10_253_3808_0,
    i_10_253_3835_0, i_10_253_3855_0, i_10_253_3889_0, i_10_253_3920_0,
    i_10_253_3981_0, i_10_253_3991_0, i_10_253_4129_0, i_10_253_4272_0,
    i_10_253_4273_0, i_10_253_4281_0, i_10_253_4290_0, i_10_253_4292_0;
  output o_10_253_0_0;
  assign o_10_253_0_0 = 0;
endmodule



// Benchmark "kernel_10_254" written by ABC on Sun Jul 19 10:25:23 2020

module kernel_10_254 ( 
    i_10_254_40_0, i_10_254_41_0, i_10_254_175_0, i_10_254_185_0,
    i_10_254_197_0, i_10_254_251_0, i_10_254_268_0, i_10_254_269_0,
    i_10_254_280_0, i_10_254_286_0, i_10_254_319_0, i_10_254_320_0,
    i_10_254_410_0, i_10_254_447_0, i_10_254_462_0, i_10_254_463_0,
    i_10_254_533_0, i_10_254_697_0, i_10_254_700_0, i_10_254_701_0,
    i_10_254_737_0, i_10_254_794_0, i_10_254_995_0, i_10_254_997_0,
    i_10_254_998_0, i_10_254_1003_0, i_10_254_1043_0, i_10_254_1088_0,
    i_10_254_1236_0, i_10_254_1237_0, i_10_254_1240_0, i_10_254_1349_0,
    i_10_254_1445_0, i_10_254_1582_0, i_10_254_1601_0, i_10_254_1653_0,
    i_10_254_1654_0, i_10_254_1655_0, i_10_254_1685_0, i_10_254_1817_0,
    i_10_254_1823_0, i_10_254_1946_0, i_10_254_1949_0, i_10_254_2006_0,
    i_10_254_2158_0, i_10_254_2311_0, i_10_254_2334_0, i_10_254_2339_0,
    i_10_254_2355_0, i_10_254_2383_0, i_10_254_2384_0, i_10_254_2453_0,
    i_10_254_2470_0, i_10_254_2471_0, i_10_254_2510_0, i_10_254_2635_0,
    i_10_254_2636_0, i_10_254_2680_0, i_10_254_2681_0, i_10_254_2707_0,
    i_10_254_2729_0, i_10_254_2786_0, i_10_254_2825_0, i_10_254_2828_0,
    i_10_254_2830_0, i_10_254_2883_0, i_10_254_2887_0, i_10_254_2983_0,
    i_10_254_2985_0, i_10_254_3038_0, i_10_254_3073_0, i_10_254_3076_0,
    i_10_254_3196_0, i_10_254_3274_0, i_10_254_3284_0, i_10_254_3290_0,
    i_10_254_3302_0, i_10_254_3409_0, i_10_254_3410_0, i_10_254_3472_0,
    i_10_254_3611_0, i_10_254_3616_0, i_10_254_3649_0, i_10_254_3650_0,
    i_10_254_3688_0, i_10_254_3784_0, i_10_254_3837_0, i_10_254_3853_0,
    i_10_254_3854_0, i_10_254_3857_0, i_10_254_3859_0, i_10_254_3896_0,
    i_10_254_3919_0, i_10_254_3985_0, i_10_254_3986_0, i_10_254_3991_0,
    i_10_254_3994_0, i_10_254_4220_0, i_10_254_4283_0, i_10_254_4289_0,
    o_10_254_0_0  );
  input  i_10_254_40_0, i_10_254_41_0, i_10_254_175_0, i_10_254_185_0,
    i_10_254_197_0, i_10_254_251_0, i_10_254_268_0, i_10_254_269_0,
    i_10_254_280_0, i_10_254_286_0, i_10_254_319_0, i_10_254_320_0,
    i_10_254_410_0, i_10_254_447_0, i_10_254_462_0, i_10_254_463_0,
    i_10_254_533_0, i_10_254_697_0, i_10_254_700_0, i_10_254_701_0,
    i_10_254_737_0, i_10_254_794_0, i_10_254_995_0, i_10_254_997_0,
    i_10_254_998_0, i_10_254_1003_0, i_10_254_1043_0, i_10_254_1088_0,
    i_10_254_1236_0, i_10_254_1237_0, i_10_254_1240_0, i_10_254_1349_0,
    i_10_254_1445_0, i_10_254_1582_0, i_10_254_1601_0, i_10_254_1653_0,
    i_10_254_1654_0, i_10_254_1655_0, i_10_254_1685_0, i_10_254_1817_0,
    i_10_254_1823_0, i_10_254_1946_0, i_10_254_1949_0, i_10_254_2006_0,
    i_10_254_2158_0, i_10_254_2311_0, i_10_254_2334_0, i_10_254_2339_0,
    i_10_254_2355_0, i_10_254_2383_0, i_10_254_2384_0, i_10_254_2453_0,
    i_10_254_2470_0, i_10_254_2471_0, i_10_254_2510_0, i_10_254_2635_0,
    i_10_254_2636_0, i_10_254_2680_0, i_10_254_2681_0, i_10_254_2707_0,
    i_10_254_2729_0, i_10_254_2786_0, i_10_254_2825_0, i_10_254_2828_0,
    i_10_254_2830_0, i_10_254_2883_0, i_10_254_2887_0, i_10_254_2983_0,
    i_10_254_2985_0, i_10_254_3038_0, i_10_254_3073_0, i_10_254_3076_0,
    i_10_254_3196_0, i_10_254_3274_0, i_10_254_3284_0, i_10_254_3290_0,
    i_10_254_3302_0, i_10_254_3409_0, i_10_254_3410_0, i_10_254_3472_0,
    i_10_254_3611_0, i_10_254_3616_0, i_10_254_3649_0, i_10_254_3650_0,
    i_10_254_3688_0, i_10_254_3784_0, i_10_254_3837_0, i_10_254_3853_0,
    i_10_254_3854_0, i_10_254_3857_0, i_10_254_3859_0, i_10_254_3896_0,
    i_10_254_3919_0, i_10_254_3985_0, i_10_254_3986_0, i_10_254_3991_0,
    i_10_254_3994_0, i_10_254_4220_0, i_10_254_4283_0, i_10_254_4289_0;
  output o_10_254_0_0;
  assign o_10_254_0_0 = ~((~i_10_254_2983_0 & ((~i_10_254_320_0 & ((~i_10_254_700_0 & i_10_254_1654_0 & ~i_10_254_1823_0 & ~i_10_254_2681_0 & ~i_10_254_2985_0 & ~i_10_254_3616_0 & ~i_10_254_3784_0) | (~i_10_254_319_0 & ~i_10_254_1043_0 & ~i_10_254_1655_0 & ~i_10_254_2311_0 & ~i_10_254_2825_0 & i_10_254_3616_0 & ~i_10_254_3986_0))) | (~i_10_254_447_0 & ~i_10_254_697_0 & ((~i_10_254_998_0 & ~i_10_254_1685_0 & ~i_10_254_2355_0 & ~i_10_254_2453_0 & ~i_10_254_2680_0 & ~i_10_254_2681_0 & ~i_10_254_2830_0 & ~i_10_254_3076_0 & ~i_10_254_3611_0) | (~i_10_254_997_0 & ~i_10_254_2510_0 & ~i_10_254_2828_0 & ~i_10_254_3649_0 & ~i_10_254_3650_0 & ~i_10_254_3896_0))) | (i_10_254_463_0 & ~i_10_254_995_0 & ~i_10_254_1349_0 & ~i_10_254_1817_0 & ~i_10_254_3985_0))) | (~i_10_254_319_0 & ((~i_10_254_1349_0 & ~i_10_254_1817_0 & ~i_10_254_1949_0 & ~i_10_254_2339_0 & ~i_10_254_2786_0 & ~i_10_254_2887_0 & ~i_10_254_3196_0 & ~i_10_254_3409_0 & ~i_10_254_3611_0) | (i_10_254_3859_0 & ~i_10_254_3896_0 & ~i_10_254_3994_0))) | (i_10_254_463_0 & ((i_10_254_286_0 & i_10_254_998_0 & i_10_254_3284_0) | (~i_10_254_320_0 & ~i_10_254_997_0 & ~i_10_254_998_0 & ~i_10_254_2681_0 & ~i_10_254_3688_0))) | (i_10_254_286_0 & ((~i_10_254_1655_0 & i_10_254_2680_0 & ~i_10_254_3688_0 & ~i_10_254_3837_0) | (~i_10_254_995_0 & ~i_10_254_998_0 & ~i_10_254_1349_0 & ~i_10_254_2339_0 & ~i_10_254_3616_0 & ~i_10_254_3991_0 & ~i_10_254_4289_0))) | (~i_10_254_2729_0 & ((~i_10_254_410_0 & ((~i_10_254_700_0 & ~i_10_254_1445_0 & ~i_10_254_1817_0 & ~i_10_254_1949_0 & ~i_10_254_2510_0 & ~i_10_254_2828_0 & ~i_10_254_3896_0 & ~i_10_254_3991_0) | (~i_10_254_175_0 & ~i_10_254_1043_0 & ~i_10_254_2339_0 & ~i_10_254_2355_0 & ~i_10_254_2471_0 & ~i_10_254_2887_0 & ~i_10_254_3854_0 & ~i_10_254_4283_0))) | (~i_10_254_1349_0 & ~i_10_254_2339_0 & ((~i_10_254_320_0 & ~i_10_254_700_0 & ~i_10_254_995_0 & ~i_10_254_1949_0 & ~i_10_254_2887_0 & ~i_10_254_3409_0 & ~i_10_254_3985_0) | (~i_10_254_462_0 & i_10_254_1655_0 & ~i_10_254_1817_0 & ~i_10_254_3038_0 & ~i_10_254_3196_0 & ~i_10_254_3649_0 & ~i_10_254_3853_0 & i_10_254_3986_0 & ~i_10_254_4289_0))) | (i_10_254_995_0 & ~i_10_254_1655_0 & i_10_254_2680_0 & i_10_254_3854_0))) | (~i_10_254_997_0 & ((~i_10_254_320_0 & ~i_10_254_2339_0 & ((~i_10_254_251_0 & ~i_10_254_701_0 & ~i_10_254_2355_0 & ~i_10_254_2883_0 & ~i_10_254_3274_0) | (~i_10_254_286_0 & i_10_254_2983_0 & ~i_10_254_3650_0 & ~i_10_254_3853_0 & ~i_10_254_3986_0))) | (i_10_254_462_0 & ~i_10_254_2510_0 & ~i_10_254_3616_0 & ~i_10_254_3649_0))) | (~i_10_254_2830_0 & ((~i_10_254_1349_0 & ((~i_10_254_995_0 & i_10_254_1823_0 & ~i_10_254_2883_0 & ~i_10_254_3611_0 & ~i_10_254_3896_0) | (~i_10_254_697_0 & ~i_10_254_701_0 & ~i_10_254_1817_0 & ~i_10_254_2311_0 & ~i_10_254_2510_0 & i_10_254_3854_0 & ~i_10_254_3985_0 & ~i_10_254_3991_0))) | (i_10_254_1653_0 & i_10_254_3038_0 & ~i_10_254_3985_0) | (~i_10_254_410_0 & ~i_10_254_2825_0 & ~i_10_254_3616_0 & ~i_10_254_3688_0 & i_10_254_3985_0))) | (~i_10_254_3991_0 & ((~i_10_254_3274_0 & ((~i_10_254_998_0 & ~i_10_254_2510_0 & ~i_10_254_3611_0 & ~i_10_254_3649_0 & ~i_10_254_3650_0 & ~i_10_254_3985_0) | (i_10_254_1240_0 & ~i_10_254_2470_0 & ~i_10_254_2471_0 & ~i_10_254_3994_0 & ~i_10_254_4220_0))) | (i_10_254_3649_0 & i_10_254_3857_0 & i_10_254_4220_0))) | (~i_10_254_1582_0 & i_10_254_1654_0 & i_10_254_2680_0 & ~i_10_254_3616_0 & ~i_10_254_3986_0));
endmodule



// Benchmark "kernel_10_255" written by ABC on Sun Jul 19 10:25:25 2020

module kernel_10_255 ( 
    i_10_255_35_0, i_10_255_175_0, i_10_255_176_0, i_10_255_218_0,
    i_10_255_223_0, i_10_255_282_0, i_10_255_410_0, i_10_255_444_0,
    i_10_255_460_0, i_10_255_462_0, i_10_255_463_0, i_10_255_464_0,
    i_10_255_798_0, i_10_255_799_0, i_10_255_969_0, i_10_255_970_0,
    i_10_255_994_0, i_10_255_1005_0, i_10_255_1030_0, i_10_255_1138_0,
    i_10_255_1236_0, i_10_255_1237_0, i_10_255_1238_0, i_10_255_1260_0,
    i_10_255_1305_0, i_10_255_1309_0, i_10_255_1310_0, i_10_255_1362_0,
    i_10_255_1654_0, i_10_255_1686_0, i_10_255_1687_0, i_10_255_1819_0,
    i_10_255_1820_0, i_10_255_1823_0, i_10_255_1909_0, i_10_255_1911_0,
    i_10_255_1944_0, i_10_255_1989_0, i_10_255_1990_0, i_10_255_2180_0,
    i_10_255_2183_0, i_10_255_2305_0, i_10_255_2310_0, i_10_255_2409_0,
    i_10_255_2450_0, i_10_255_2472_0, i_10_255_2632_0, i_10_255_2657_0,
    i_10_255_2659_0, i_10_255_2701_0, i_10_255_2711_0, i_10_255_2713_0,
    i_10_255_2727_0, i_10_255_2785_0, i_10_255_2830_0, i_10_255_2833_0,
    i_10_255_2881_0, i_10_255_2883_0, i_10_255_2885_0, i_10_255_2920_0,
    i_10_255_3034_0, i_10_255_3036_0, i_10_255_3037_0, i_10_255_3038_0,
    i_10_255_3039_0, i_10_255_3040_0, i_10_255_3069_0, i_10_255_3199_0,
    i_10_255_3200_0, i_10_255_3323_0, i_10_255_3386_0, i_10_255_3389_0,
    i_10_255_3403_0, i_10_255_3405_0, i_10_255_3406_0, i_10_255_3585_0,
    i_10_255_3588_0, i_10_255_3590_0, i_10_255_3649_0, i_10_255_3652_0,
    i_10_255_3653_0, i_10_255_3835_0, i_10_255_3842_0, i_10_255_3846_0,
    i_10_255_3848_0, i_10_255_3857_0, i_10_255_3882_0, i_10_255_3981_0,
    i_10_255_3982_0, i_10_255_3985_0, i_10_255_4116_0, i_10_255_4118_0,
    i_10_255_4125_0, i_10_255_4126_0, i_10_255_4127_0, i_10_255_4218_0,
    i_10_255_4269_0, i_10_255_4273_0, i_10_255_4289_0, i_10_255_4566_0,
    o_10_255_0_0  );
  input  i_10_255_35_0, i_10_255_175_0, i_10_255_176_0, i_10_255_218_0,
    i_10_255_223_0, i_10_255_282_0, i_10_255_410_0, i_10_255_444_0,
    i_10_255_460_0, i_10_255_462_0, i_10_255_463_0, i_10_255_464_0,
    i_10_255_798_0, i_10_255_799_0, i_10_255_969_0, i_10_255_970_0,
    i_10_255_994_0, i_10_255_1005_0, i_10_255_1030_0, i_10_255_1138_0,
    i_10_255_1236_0, i_10_255_1237_0, i_10_255_1238_0, i_10_255_1260_0,
    i_10_255_1305_0, i_10_255_1309_0, i_10_255_1310_0, i_10_255_1362_0,
    i_10_255_1654_0, i_10_255_1686_0, i_10_255_1687_0, i_10_255_1819_0,
    i_10_255_1820_0, i_10_255_1823_0, i_10_255_1909_0, i_10_255_1911_0,
    i_10_255_1944_0, i_10_255_1989_0, i_10_255_1990_0, i_10_255_2180_0,
    i_10_255_2183_0, i_10_255_2305_0, i_10_255_2310_0, i_10_255_2409_0,
    i_10_255_2450_0, i_10_255_2472_0, i_10_255_2632_0, i_10_255_2657_0,
    i_10_255_2659_0, i_10_255_2701_0, i_10_255_2711_0, i_10_255_2713_0,
    i_10_255_2727_0, i_10_255_2785_0, i_10_255_2830_0, i_10_255_2833_0,
    i_10_255_2881_0, i_10_255_2883_0, i_10_255_2885_0, i_10_255_2920_0,
    i_10_255_3034_0, i_10_255_3036_0, i_10_255_3037_0, i_10_255_3038_0,
    i_10_255_3039_0, i_10_255_3040_0, i_10_255_3069_0, i_10_255_3199_0,
    i_10_255_3200_0, i_10_255_3323_0, i_10_255_3386_0, i_10_255_3389_0,
    i_10_255_3403_0, i_10_255_3405_0, i_10_255_3406_0, i_10_255_3585_0,
    i_10_255_3588_0, i_10_255_3590_0, i_10_255_3649_0, i_10_255_3652_0,
    i_10_255_3653_0, i_10_255_3835_0, i_10_255_3842_0, i_10_255_3846_0,
    i_10_255_3848_0, i_10_255_3857_0, i_10_255_3882_0, i_10_255_3981_0,
    i_10_255_3982_0, i_10_255_3985_0, i_10_255_4116_0, i_10_255_4118_0,
    i_10_255_4125_0, i_10_255_4126_0, i_10_255_4127_0, i_10_255_4218_0,
    i_10_255_4269_0, i_10_255_4273_0, i_10_255_4289_0, i_10_255_4566_0;
  output o_10_255_0_0;
  assign o_10_255_0_0 = ~((i_10_255_175_0 & ((~i_10_255_460_0 & i_10_255_1237_0 & ~i_10_255_1944_0 & ~i_10_255_2310_0 & ~i_10_255_2632_0 & ~i_10_255_2830_0 & ~i_10_255_3649_0 & ~i_10_255_3857_0) | (~i_10_255_463_0 & i_10_255_798_0 & ~i_10_255_3036_0 & i_10_255_3389_0 & ~i_10_255_4273_0))) | (i_10_255_176_0 & ((i_10_255_464_0 & ~i_10_255_1260_0 & ~i_10_255_1654_0 & ~i_10_255_2472_0 & ~i_10_255_3036_0 & ~i_10_255_3039_0) | (~i_10_255_969_0 & i_10_255_2632_0 & ~i_10_255_3037_0 & ~i_10_255_3649_0))) | (~i_10_255_970_0 & ((~i_10_255_35_0 & ~i_10_255_444_0 & ~i_10_255_798_0 & ~i_10_255_1236_0 & ((i_10_255_3200_0 & ~i_10_255_3590_0 & i_10_255_3652_0) | (~i_10_255_1823_0 & ~i_10_255_2180_0 & ~i_10_255_2659_0 & ~i_10_255_3039_0 & ~i_10_255_3985_0))) | (~i_10_255_282_0 & ~i_10_255_3406_0 & ((~i_10_255_969_0 & ~i_10_255_1030_0 & ~i_10_255_1305_0 & ~i_10_255_2183_0 & ~i_10_255_2310_0 & ~i_10_255_2659_0 & ~i_10_255_2883_0 & ~i_10_255_2920_0 & ~i_10_255_3040_0 & ~i_10_255_3405_0 & ~i_10_255_3835_0 & ~i_10_255_3857_0) | (~i_10_255_2180_0 & i_10_255_2920_0 & ~i_10_255_3649_0 & ~i_10_255_4566_0))) | (~i_10_255_462_0 & ((~i_10_255_3037_0 & ~i_10_255_3649_0 & ~i_10_255_799_0 & ~i_10_255_1911_0) | (~i_10_255_464_0 & i_10_255_1819_0 & i_10_255_3835_0))) | (~i_10_255_2727_0 & ((~i_10_255_2310_0 & i_10_255_2701_0 & ~i_10_255_2830_0 & ~i_10_255_3034_0 & ~i_10_255_3037_0) | (~i_10_255_3038_0 & i_10_255_3848_0))) | (~i_10_255_460_0 & ~i_10_255_464_0 & ~i_10_255_1005_0 & ~i_10_255_1260_0 & ~i_10_255_1911_0 & ~i_10_255_1944_0 & ~i_10_255_3038_0 & ~i_10_255_3652_0 & ~i_10_255_3835_0 & ~i_10_255_4566_0))) | (~i_10_255_282_0 & ((i_10_255_1687_0 & ~i_10_255_2183_0 & ~i_10_255_2659_0 & ~i_10_255_3585_0 & i_10_255_3653_0) | (~i_10_255_1260_0 & i_10_255_2632_0 & ~i_10_255_3036_0 & ~i_10_255_3037_0 & ~i_10_255_3653_0 & ~i_10_255_3982_0 & i_10_255_4118_0 & ~i_10_255_4273_0))) | (~i_10_255_463_0 & ((~i_10_255_3588_0 & ((~i_10_255_460_0 & ((~i_10_255_35_0 & ~i_10_255_969_0 & ~i_10_255_1237_0 & ~i_10_255_2409_0 & ~i_10_255_2659_0 & ~i_10_255_2833_0 & ~i_10_255_3200_0 & ~i_10_255_3405_0) | (~i_10_255_464_0 & ~i_10_255_1944_0 & ~i_10_255_2310_0 & ~i_10_255_3040_0 & ~i_10_255_4273_0 & ~i_10_255_4566_0))) | (~i_10_255_1310_0 & i_10_255_2833_0 & ~i_10_255_3199_0))) | (~i_10_255_464_0 & ~i_10_255_1236_0 & ~i_10_255_1238_0 & ~i_10_255_2409_0 & ~i_10_255_2701_0 & ~i_10_255_2920_0 & ~i_10_255_3037_0))) | (~i_10_255_2727_0 & ((~i_10_255_35_0 & ~i_10_255_2409_0 & ~i_10_255_2701_0 & ~i_10_255_3039_0 & ~i_10_255_4566_0 & ((i_10_255_464_0 & ~i_10_255_3034_0 & ~i_10_255_3036_0 & ~i_10_255_3590_0) | (~i_10_255_969_0 & ~i_10_255_2885_0 & ~i_10_255_3585_0 & ~i_10_255_3857_0))) | (i_10_255_1819_0 & ~i_10_255_3037_0 & i_10_255_3846_0) | (i_10_255_3406_0 & ~i_10_255_3585_0 & ~i_10_255_3590_0 & ~i_10_255_4269_0))) | (~i_10_255_799_0 & ((i_10_255_1819_0 & ~i_10_255_3649_0 & i_10_255_3848_0) | (~i_10_255_798_0 & ~i_10_255_969_0 & ~i_10_255_1236_0 & ~i_10_255_1823_0 & ~i_10_255_3038_0 & ~i_10_255_3039_0 & ~i_10_255_3857_0 & i_10_255_3982_0))) | (~i_10_255_3588_0 & ((~i_10_255_798_0 & ~i_10_255_3590_0 & i_10_255_3652_0 & ((~i_10_255_410_0 & ~i_10_255_1005_0 & ~i_10_255_2310_0 & ~i_10_255_2885_0 & i_10_255_3199_0) | (~i_10_255_460_0 & ~i_10_255_1305_0 & ~i_10_255_1944_0 & ~i_10_255_4273_0 & ~i_10_255_4566_0 & i_10_255_3649_0 & ~i_10_255_3985_0))) | (~i_10_255_1309_0 & ~i_10_255_1909_0 & ~i_10_255_2657_0 & i_10_255_2659_0 & ~i_10_255_3835_0))) | (~i_10_255_1005_0 & ((~i_10_255_460_0 & ((~i_10_255_969_0 & ~i_10_255_2472_0 & ~i_10_255_3038_0 & ~i_10_255_3848_0 & i_10_255_3981_0) | (~i_10_255_1260_0 & i_10_255_1654_0 & ~i_10_255_3585_0 & i_10_255_4118_0 & ~i_10_255_4273_0))) | (~i_10_255_410_0 & i_10_255_2713_0 & ~i_10_255_2830_0 & ~i_10_255_3405_0 & ~i_10_255_3406_0 & i_10_255_3590_0))) | (~i_10_255_4269_0 & ((~i_10_255_410_0 & ((~i_10_255_2632_0 & i_10_255_2713_0 & ~i_10_255_2830_0 & ~i_10_255_2920_0 & ~i_10_255_3038_0 & ~i_10_255_3389_0) | (~i_10_255_175_0 & ~i_10_255_1030_0 & i_10_255_1687_0 & ~i_10_255_2711_0 & i_10_255_3649_0 & ~i_10_255_3652_0 & ~i_10_255_4289_0))) | (i_10_255_799_0 & ~i_10_255_1686_0 & ~i_10_255_3037_0 & ~i_10_255_3038_0 & ~i_10_255_3585_0 & ~i_10_255_3848_0 & ~i_10_255_4118_0))) | (~i_10_255_969_0 & ~i_10_255_1944_0 & ~i_10_255_2881_0 & ((i_10_255_1819_0 & ~i_10_255_2920_0 & i_10_255_4116_0) | (~i_10_255_1911_0 & ~i_10_255_2409_0 & ~i_10_255_2657_0 & ~i_10_255_3038_0 & ~i_10_255_3039_0 & ~i_10_255_3040_0 & ~i_10_255_3585_0 & ~i_10_255_3857_0 & ~i_10_255_3982_0 & ~i_10_255_4116_0))) | (i_10_255_1909_0 & i_10_255_3034_0 & ~i_10_255_3040_0) | (~i_10_255_462_0 & ~i_10_255_3038_0 & i_10_255_3386_0) | (~i_10_255_2310_0 & i_10_255_4218_0 & i_10_255_4566_0) | (~i_10_255_1236_0 & ~i_10_255_2830_0 & ~i_10_255_3037_0 & i_10_255_4269_0 & ~i_10_255_4566_0));
endmodule



// Benchmark "kernel_10_256" written by ABC on Sun Jul 19 10:25:26 2020

module kernel_10_256 ( 
    i_10_256_41_0, i_10_256_255_0, i_10_256_282_0, i_10_256_409_0,
    i_10_256_423_0, i_10_256_430_0, i_10_256_431_0, i_10_256_436_0,
    i_10_256_444_0, i_10_256_445_0, i_10_256_446_0, i_10_256_447_0,
    i_10_256_448_0, i_10_256_466_0, i_10_256_716_0, i_10_256_794_0,
    i_10_256_796_0, i_10_256_800_0, i_10_256_967_0, i_10_256_968_0,
    i_10_256_969_0, i_10_256_970_0, i_10_256_1240_0, i_10_256_1241_0,
    i_10_256_1243_0, i_10_256_1266_0, i_10_256_1365_0, i_10_256_1452_0,
    i_10_256_1453_0, i_10_256_1548_0, i_10_256_1580_0, i_10_256_1582_0,
    i_10_256_1583_0, i_10_256_1629_0, i_10_256_1650_0, i_10_256_1651_0,
    i_10_256_1655_0, i_10_256_1683_0, i_10_256_1690_0, i_10_256_1691_0,
    i_10_256_2203_0, i_10_256_2352_0, i_10_256_2362_0, i_10_256_2363_0,
    i_10_256_2364_0, i_10_256_2365_0, i_10_256_2366_0, i_10_256_2376_0,
    i_10_256_2410_0, i_10_256_2411_0, i_10_256_2469_0, i_10_256_2470_0,
    i_10_256_2472_0, i_10_256_2473_0, i_10_256_2474_0, i_10_256_2631_0,
    i_10_256_2632_0, i_10_256_2659_0, i_10_256_2660_0, i_10_256_2661_0,
    i_10_256_2662_0, i_10_256_2663_0, i_10_256_2702_0, i_10_256_2716_0,
    i_10_256_2734_0, i_10_256_2735_0, i_10_256_2831_0, i_10_256_2832_0,
    i_10_256_2982_0, i_10_256_3049_0, i_10_256_3087_0, i_10_256_3165_0,
    i_10_256_3385_0, i_10_256_3386_0, i_10_256_3388_0, i_10_256_3389_0,
    i_10_256_3390_0, i_10_256_3391_0, i_10_256_3392_0, i_10_256_3468_0,
    i_10_256_3469_0, i_10_256_3470_0, i_10_256_3586_0, i_10_256_3587_0,
    i_10_256_3588_0, i_10_256_3589_0, i_10_256_3590_0, i_10_256_3783_0,
    i_10_256_3784_0, i_10_256_3787_0, i_10_256_3834_0, i_10_256_3843_0,
    i_10_256_4058_0, i_10_256_4116_0, i_10_256_4117_0, i_10_256_4119_0,
    i_10_256_4165_0, i_10_256_4270_0, i_10_256_4365_0, i_10_256_4585_0,
    o_10_256_0_0  );
  input  i_10_256_41_0, i_10_256_255_0, i_10_256_282_0, i_10_256_409_0,
    i_10_256_423_0, i_10_256_430_0, i_10_256_431_0, i_10_256_436_0,
    i_10_256_444_0, i_10_256_445_0, i_10_256_446_0, i_10_256_447_0,
    i_10_256_448_0, i_10_256_466_0, i_10_256_716_0, i_10_256_794_0,
    i_10_256_796_0, i_10_256_800_0, i_10_256_967_0, i_10_256_968_0,
    i_10_256_969_0, i_10_256_970_0, i_10_256_1240_0, i_10_256_1241_0,
    i_10_256_1243_0, i_10_256_1266_0, i_10_256_1365_0, i_10_256_1452_0,
    i_10_256_1453_0, i_10_256_1548_0, i_10_256_1580_0, i_10_256_1582_0,
    i_10_256_1583_0, i_10_256_1629_0, i_10_256_1650_0, i_10_256_1651_0,
    i_10_256_1655_0, i_10_256_1683_0, i_10_256_1690_0, i_10_256_1691_0,
    i_10_256_2203_0, i_10_256_2352_0, i_10_256_2362_0, i_10_256_2363_0,
    i_10_256_2364_0, i_10_256_2365_0, i_10_256_2366_0, i_10_256_2376_0,
    i_10_256_2410_0, i_10_256_2411_0, i_10_256_2469_0, i_10_256_2470_0,
    i_10_256_2472_0, i_10_256_2473_0, i_10_256_2474_0, i_10_256_2631_0,
    i_10_256_2632_0, i_10_256_2659_0, i_10_256_2660_0, i_10_256_2661_0,
    i_10_256_2662_0, i_10_256_2663_0, i_10_256_2702_0, i_10_256_2716_0,
    i_10_256_2734_0, i_10_256_2735_0, i_10_256_2831_0, i_10_256_2832_0,
    i_10_256_2982_0, i_10_256_3049_0, i_10_256_3087_0, i_10_256_3165_0,
    i_10_256_3385_0, i_10_256_3386_0, i_10_256_3388_0, i_10_256_3389_0,
    i_10_256_3390_0, i_10_256_3391_0, i_10_256_3392_0, i_10_256_3468_0,
    i_10_256_3469_0, i_10_256_3470_0, i_10_256_3586_0, i_10_256_3587_0,
    i_10_256_3588_0, i_10_256_3589_0, i_10_256_3590_0, i_10_256_3783_0,
    i_10_256_3784_0, i_10_256_3787_0, i_10_256_3834_0, i_10_256_3843_0,
    i_10_256_4058_0, i_10_256_4116_0, i_10_256_4117_0, i_10_256_4119_0,
    i_10_256_4165_0, i_10_256_4270_0, i_10_256_4365_0, i_10_256_4585_0;
  output o_10_256_0_0;
  assign o_10_256_0_0 = 0;
endmodule



// Benchmark "kernel_10_257" written by ABC on Sun Jul 19 10:25:27 2020

module kernel_10_257 ( 
    i_10_257_149_0, i_10_257_174_0, i_10_257_175_0, i_10_257_177_0,
    i_10_257_178_0, i_10_257_183_0, i_10_257_184_0, i_10_257_185_0,
    i_10_257_187_0, i_10_257_286_0, i_10_257_319_0, i_10_257_328_0,
    i_10_257_329_0, i_10_257_408_0, i_10_257_409_0, i_10_257_410_0,
    i_10_257_442_0, i_10_257_463_0, i_10_257_510_0, i_10_257_753_0,
    i_10_257_754_0, i_10_257_796_0, i_10_257_967_0, i_10_257_1032_0,
    i_10_257_1042_0, i_10_257_1043_0, i_10_257_1169_0, i_10_257_1250_0,
    i_10_257_1263_0, i_10_257_1582_0, i_10_257_1651_0, i_10_257_1652_0,
    i_10_257_1653_0, i_10_257_1654_0, i_10_257_1655_0, i_10_257_1684_0,
    i_10_257_1821_0, i_10_257_1822_0, i_10_257_1824_0, i_10_257_1825_0,
    i_10_257_1826_0, i_10_257_1910_0, i_10_257_1952_0, i_10_257_2185_0,
    i_10_257_2307_0, i_10_257_2352_0, i_10_257_2353_0, i_10_257_2354_0,
    i_10_257_2355_0, i_10_257_2410_0, i_10_257_2452_0, i_10_257_2454_0,
    i_10_257_2470_0, i_10_257_2473_0, i_10_257_2474_0, i_10_257_2608_0,
    i_10_257_2701_0, i_10_257_2704_0, i_10_257_2713_0, i_10_257_2716_0,
    i_10_257_2735_0, i_10_257_2833_0, i_10_257_2916_0, i_10_257_2919_0,
    i_10_257_2920_0, i_10_257_2921_0, i_10_257_2980_0, i_10_257_2985_0,
    i_10_257_3035_0, i_10_257_3050_0, i_10_257_3152_0, i_10_257_3162_0,
    i_10_257_3271_0, i_10_257_3279_0, i_10_257_3280_0, i_10_257_3387_0,
    i_10_257_3388_0, i_10_257_3390_0, i_10_257_3391_0, i_10_257_3405_0,
    i_10_257_3472_0, i_10_257_3611_0, i_10_257_3613_0, i_10_257_3614_0,
    i_10_257_3615_0, i_10_257_3646_0, i_10_257_3647_0, i_10_257_3653_0,
    i_10_257_3725_0, i_10_257_3834_0, i_10_257_3837_0, i_10_257_3840_0,
    i_10_257_3857_0, i_10_257_3895_0, i_10_257_3990_0, i_10_257_3991_0,
    i_10_257_4115_0, i_10_257_4182_0, i_10_257_4189_0, i_10_257_4282_0,
    o_10_257_0_0  );
  input  i_10_257_149_0, i_10_257_174_0, i_10_257_175_0, i_10_257_177_0,
    i_10_257_178_0, i_10_257_183_0, i_10_257_184_0, i_10_257_185_0,
    i_10_257_187_0, i_10_257_286_0, i_10_257_319_0, i_10_257_328_0,
    i_10_257_329_0, i_10_257_408_0, i_10_257_409_0, i_10_257_410_0,
    i_10_257_442_0, i_10_257_463_0, i_10_257_510_0, i_10_257_753_0,
    i_10_257_754_0, i_10_257_796_0, i_10_257_967_0, i_10_257_1032_0,
    i_10_257_1042_0, i_10_257_1043_0, i_10_257_1169_0, i_10_257_1250_0,
    i_10_257_1263_0, i_10_257_1582_0, i_10_257_1651_0, i_10_257_1652_0,
    i_10_257_1653_0, i_10_257_1654_0, i_10_257_1655_0, i_10_257_1684_0,
    i_10_257_1821_0, i_10_257_1822_0, i_10_257_1824_0, i_10_257_1825_0,
    i_10_257_1826_0, i_10_257_1910_0, i_10_257_1952_0, i_10_257_2185_0,
    i_10_257_2307_0, i_10_257_2352_0, i_10_257_2353_0, i_10_257_2354_0,
    i_10_257_2355_0, i_10_257_2410_0, i_10_257_2452_0, i_10_257_2454_0,
    i_10_257_2470_0, i_10_257_2473_0, i_10_257_2474_0, i_10_257_2608_0,
    i_10_257_2701_0, i_10_257_2704_0, i_10_257_2713_0, i_10_257_2716_0,
    i_10_257_2735_0, i_10_257_2833_0, i_10_257_2916_0, i_10_257_2919_0,
    i_10_257_2920_0, i_10_257_2921_0, i_10_257_2980_0, i_10_257_2985_0,
    i_10_257_3035_0, i_10_257_3050_0, i_10_257_3152_0, i_10_257_3162_0,
    i_10_257_3271_0, i_10_257_3279_0, i_10_257_3280_0, i_10_257_3387_0,
    i_10_257_3388_0, i_10_257_3390_0, i_10_257_3391_0, i_10_257_3405_0,
    i_10_257_3472_0, i_10_257_3611_0, i_10_257_3613_0, i_10_257_3614_0,
    i_10_257_3615_0, i_10_257_3646_0, i_10_257_3647_0, i_10_257_3653_0,
    i_10_257_3725_0, i_10_257_3834_0, i_10_257_3837_0, i_10_257_3840_0,
    i_10_257_3857_0, i_10_257_3895_0, i_10_257_3990_0, i_10_257_3991_0,
    i_10_257_4115_0, i_10_257_4182_0, i_10_257_4189_0, i_10_257_4282_0;
  output o_10_257_0_0;
  assign o_10_257_0_0 = ~((i_10_257_174_0 & ((i_10_257_1655_0 & ~i_10_257_2916_0 & i_10_257_2921_0 & ~i_10_257_3895_0 & ~i_10_257_3991_0) | (~i_10_257_184_0 & ~i_10_257_2354_0 & ~i_10_257_2473_0 & ~i_10_257_2919_0 & ~i_10_257_2920_0 & ~i_10_257_2921_0 & ~i_10_257_3405_0 & ~i_10_257_3611_0 & ~i_10_257_4282_0))) | (~i_10_257_2735_0 & ((~i_10_257_174_0 & ((~i_10_257_175_0 & ~i_10_257_442_0 & ~i_10_257_1822_0) | (~i_10_257_1910_0 & ~i_10_257_3035_0 & ~i_10_257_3405_0 & i_10_257_3646_0))) | (i_10_257_319_0 & ~i_10_257_408_0 & ~i_10_257_753_0 & ~i_10_257_754_0 & ~i_10_257_1825_0 & ~i_10_257_2307_0 & ~i_10_257_2713_0) | (~i_10_257_1821_0 & i_10_257_1825_0 & ~i_10_257_3653_0) | (~i_10_257_1042_0 & ~i_10_257_1043_0 & ~i_10_257_1652_0 & i_10_257_2704_0 & ~i_10_257_3990_0))) | (~i_10_257_184_0 & ((~i_10_257_175_0 & ~i_10_257_2921_0 & ~i_10_257_3647_0 & ~i_10_257_3990_0) | (~i_10_257_408_0 & ~i_10_257_410_0 & ~i_10_257_3837_0 & ~i_10_257_3991_0))) | (~i_10_257_175_0 & ~i_10_257_753_0 & ((~i_10_257_329_0 & ~i_10_257_1263_0 & ~i_10_257_1822_0 & i_10_257_3611_0 & i_10_257_3991_0) | (~i_10_257_185_0 & ~i_10_257_409_0 & ~i_10_257_410_0 & ~i_10_257_1653_0 & ~i_10_257_2410_0 & ~i_10_257_2452_0 & ~i_10_257_4282_0))) | (~i_10_257_187_0 & ((i_10_257_1824_0 & ~i_10_257_2701_0 & ~i_10_257_3162_0 & ~i_10_257_3834_0) | (~i_10_257_442_0 & ~i_10_257_1042_0 & ~i_10_257_1169_0 & ~i_10_257_2608_0 & ~i_10_257_2916_0 & ~i_10_257_3614_0 & ~i_10_257_3653_0 & ~i_10_257_3991_0))) | (~i_10_257_2919_0 & ((~i_10_257_410_0 & ((~i_10_257_408_0 & ~i_10_257_2704_0 & ~i_10_257_2920_0) | (~i_10_257_1043_0 & ~i_10_257_2452_0 & ~i_10_257_3990_0 & ~i_10_257_4115_0))) | (i_10_257_1825_0 & ~i_10_257_1952_0 & ~i_10_257_3614_0 & i_10_257_3653_0) | (~i_10_257_185_0 & ~i_10_257_1651_0 & ~i_10_257_1910_0 & ~i_10_257_2701_0 & ~i_10_257_3895_0 & ~i_10_257_4115_0 & ~i_10_257_4282_0))) | (i_10_257_2713_0 & ((~i_10_257_408_0 & i_10_257_3857_0 & i_10_257_4115_0) | (~i_10_257_183_0 & ~i_10_257_3614_0 & ~i_10_257_4115_0))) | (i_10_257_2980_0 & (i_10_257_2307_0 | (~i_10_257_1250_0 & ~i_10_257_3405_0 & ~i_10_257_3895_0))) | (~i_10_257_408_0 & ((~i_10_257_409_0 & i_10_257_3647_0 & ~i_10_257_3990_0 & (~i_10_257_3611_0 | (~i_10_257_1032_0 & ~i_10_257_1042_0 & ~i_10_257_1043_0 & i_10_257_3035_0))) | (~i_10_257_1169_0 & ~i_10_257_1684_0 & ~i_10_257_2704_0 & ~i_10_257_3834_0 & ~i_10_257_3991_0))) | (i_10_257_328_0 & ~i_10_257_442_0 & i_10_257_1263_0 & ~i_10_257_1822_0) | (~i_10_257_1821_0 & ~i_10_257_2608_0 & i_10_257_3405_0) | (i_10_257_1825_0 & i_10_257_1826_0 & ~i_10_257_2452_0 & ~i_10_257_3405_0 & i_10_257_3991_0) | (~i_10_257_409_0 & i_10_257_796_0 & ~i_10_257_1653_0 & ~i_10_257_3990_0 & ~i_10_257_4115_0 & ~i_10_257_4282_0));
endmodule



// Benchmark "kernel_10_258" written by ABC on Sun Jul 19 10:25:28 2020

module kernel_10_258 ( 
    i_10_258_177_0, i_10_258_252_0, i_10_258_282_0, i_10_258_284_0,
    i_10_258_290_0, i_10_258_324_0, i_10_258_370_0, i_10_258_430_0,
    i_10_258_438_0, i_10_258_442_0, i_10_258_464_0, i_10_258_504_0,
    i_10_258_595_0, i_10_258_717_0, i_10_258_793_0, i_10_258_891_0,
    i_10_258_999_0, i_10_258_1000_0, i_10_258_1053_0, i_10_258_1245_0,
    i_10_258_1313_0, i_10_258_1443_0, i_10_258_1445_0, i_10_258_1654_0,
    i_10_258_1655_0, i_10_258_1719_0, i_10_258_1809_0, i_10_258_1819_0,
    i_10_258_1824_0, i_10_258_1825_0, i_10_258_1948_0, i_10_258_1990_0,
    i_10_258_1991_0, i_10_258_2181_0, i_10_258_2184_0, i_10_258_2245_0,
    i_10_258_2322_0, i_10_258_2331_0, i_10_258_2353_0, i_10_258_2356_0,
    i_10_258_2361_0, i_10_258_2379_0, i_10_258_2380_0, i_10_258_2453_0,
    i_10_258_2461_0, i_10_258_2566_0, i_10_258_2638_0, i_10_258_2680_0,
    i_10_258_2700_0, i_10_258_2704_0, i_10_258_2709_0, i_10_258_2881_0,
    i_10_258_2882_0, i_10_258_2885_0, i_10_258_2953_0, i_10_258_3033_0,
    i_10_258_3042_0, i_10_258_3043_0, i_10_258_3044_0, i_10_258_3045_0,
    i_10_258_3156_0, i_10_258_3196_0, i_10_258_3200_0, i_10_258_3267_0,
    i_10_258_3268_0, i_10_258_3277_0, i_10_258_3280_0, i_10_258_3288_0,
    i_10_258_3385_0, i_10_258_3386_0, i_10_258_3406_0, i_10_258_3465_0,
    i_10_258_3468_0, i_10_258_3495_0, i_10_258_3496_0, i_10_258_3525_0,
    i_10_258_3609_0, i_10_258_3610_0, i_10_258_3617_0, i_10_258_3647_0,
    i_10_258_3651_0, i_10_258_3780_0, i_10_258_3785_0, i_10_258_3836_0,
    i_10_258_3837_0, i_10_258_3851_0, i_10_258_3856_0, i_10_258_3859_0,
    i_10_258_4113_0, i_10_258_4122_0, i_10_258_4123_0, i_10_258_4126_0,
    i_10_258_4213_0, i_10_258_4231_0, i_10_258_4269_0, i_10_258_4290_0,
    i_10_258_4564_0, i_10_258_4566_0, i_10_258_4567_0, i_10_258_4568_0,
    o_10_258_0_0  );
  input  i_10_258_177_0, i_10_258_252_0, i_10_258_282_0, i_10_258_284_0,
    i_10_258_290_0, i_10_258_324_0, i_10_258_370_0, i_10_258_430_0,
    i_10_258_438_0, i_10_258_442_0, i_10_258_464_0, i_10_258_504_0,
    i_10_258_595_0, i_10_258_717_0, i_10_258_793_0, i_10_258_891_0,
    i_10_258_999_0, i_10_258_1000_0, i_10_258_1053_0, i_10_258_1245_0,
    i_10_258_1313_0, i_10_258_1443_0, i_10_258_1445_0, i_10_258_1654_0,
    i_10_258_1655_0, i_10_258_1719_0, i_10_258_1809_0, i_10_258_1819_0,
    i_10_258_1824_0, i_10_258_1825_0, i_10_258_1948_0, i_10_258_1990_0,
    i_10_258_1991_0, i_10_258_2181_0, i_10_258_2184_0, i_10_258_2245_0,
    i_10_258_2322_0, i_10_258_2331_0, i_10_258_2353_0, i_10_258_2356_0,
    i_10_258_2361_0, i_10_258_2379_0, i_10_258_2380_0, i_10_258_2453_0,
    i_10_258_2461_0, i_10_258_2566_0, i_10_258_2638_0, i_10_258_2680_0,
    i_10_258_2700_0, i_10_258_2704_0, i_10_258_2709_0, i_10_258_2881_0,
    i_10_258_2882_0, i_10_258_2885_0, i_10_258_2953_0, i_10_258_3033_0,
    i_10_258_3042_0, i_10_258_3043_0, i_10_258_3044_0, i_10_258_3045_0,
    i_10_258_3156_0, i_10_258_3196_0, i_10_258_3200_0, i_10_258_3267_0,
    i_10_258_3268_0, i_10_258_3277_0, i_10_258_3280_0, i_10_258_3288_0,
    i_10_258_3385_0, i_10_258_3386_0, i_10_258_3406_0, i_10_258_3465_0,
    i_10_258_3468_0, i_10_258_3495_0, i_10_258_3496_0, i_10_258_3525_0,
    i_10_258_3609_0, i_10_258_3610_0, i_10_258_3617_0, i_10_258_3647_0,
    i_10_258_3651_0, i_10_258_3780_0, i_10_258_3785_0, i_10_258_3836_0,
    i_10_258_3837_0, i_10_258_3851_0, i_10_258_3856_0, i_10_258_3859_0,
    i_10_258_4113_0, i_10_258_4122_0, i_10_258_4123_0, i_10_258_4126_0,
    i_10_258_4213_0, i_10_258_4231_0, i_10_258_4269_0, i_10_258_4290_0,
    i_10_258_4564_0, i_10_258_4566_0, i_10_258_4567_0, i_10_258_4568_0;
  output o_10_258_0_0;
  assign o_10_258_0_0 = ~((~i_10_258_3042_0 & ((~i_10_258_177_0 & ~i_10_258_3267_0 & ((~i_10_258_290_0 & ~i_10_258_1443_0 & ~i_10_258_2566_0 & ~i_10_258_4269_0) | (~i_10_258_2680_0 & ~i_10_258_4126_0 & ~i_10_258_4568_0))) | (~i_10_258_1443_0 & ~i_10_258_1824_0 & ~i_10_258_2353_0 & ~i_10_258_2380_0 & ~i_10_258_3033_0 & i_10_258_3385_0 & ~i_10_258_3785_0 & ~i_10_258_4126_0))) | (~i_10_258_2322_0 & ((~i_10_258_252_0 & ~i_10_258_3268_0 & ((~i_10_258_430_0 & ~i_10_258_1991_0 & ~i_10_258_2361_0 & ~i_10_258_3277_0 & ~i_10_258_3468_0 & ~i_10_258_3495_0 & ~i_10_258_4122_0) | (~i_10_258_717_0 & ~i_10_258_2638_0 & ~i_10_258_2680_0 & ~i_10_258_2700_0 & ~i_10_258_3044_0 & ~i_10_258_3785_0 & ~i_10_258_3836_0 & ~i_10_258_4123_0 & ~i_10_258_4126_0))) | (~i_10_258_2379_0 & ((~i_10_258_793_0 & ~i_10_258_891_0 & ~i_10_258_2461_0 & ~i_10_258_2709_0 & ~i_10_258_3495_0 & ~i_10_258_3496_0 & ~i_10_258_4231_0 & ~i_10_258_4269_0) | (~i_10_258_430_0 & ~i_10_258_1655_0 & ~i_10_258_2680_0 & ~i_10_258_3647_0 & ~i_10_258_3785_0 & ~i_10_258_3837_0 & ~i_10_258_3851_0 & ~i_10_258_4123_0 & ~i_10_258_4566_0))) | (~i_10_258_3045_0 & i_10_258_3856_0 & ~i_10_258_4123_0 & ~i_10_258_4564_0) | (~i_10_258_2700_0 & i_10_258_3609_0 & ~i_10_258_4568_0))) | (~i_10_258_4231_0 & ((~i_10_258_282_0 & ((~i_10_258_717_0 & ~i_10_258_1819_0 & ~i_10_258_3043_0 & ~i_10_258_3196_0 & ~i_10_258_3268_0) | (~i_10_258_430_0 & i_10_258_1655_0 & ~i_10_258_2356_0 & ~i_10_258_3837_0 & ~i_10_258_4213_0))) | (~i_10_258_284_0 & ~i_10_258_999_0 & ~i_10_258_1443_0 & i_10_258_1819_0 & ~i_10_258_1991_0 & ~i_10_258_2181_0 & ~i_10_258_2331_0 & ~i_10_258_2709_0 & ~i_10_258_3496_0))) | (~i_10_258_1445_0 & ~i_10_258_2181_0 & ((~i_10_258_1000_0 & ~i_10_258_1824_0 & ~i_10_258_2379_0 & ~i_10_258_3268_0 & ~i_10_258_3525_0 & ~i_10_258_3851_0 & ~i_10_258_4122_0 & ~i_10_258_4213_0 & ~i_10_258_4566_0) | (~i_10_258_324_0 & ~i_10_258_3043_0 & ~i_10_258_3495_0 & ~i_10_258_4123_0 & ~i_10_258_4567_0))) | (~i_10_258_1825_0 & ~i_10_258_3465_0 & ((~i_10_258_793_0 & ~i_10_258_2184_0 & i_10_258_2356_0 & ~i_10_258_2885_0 & ~i_10_258_3385_0 & i_10_258_3837_0) | (~i_10_258_290_0 & ~i_10_258_430_0 & ~i_10_258_1443_0 & ~i_10_258_4123_0 & ~i_10_258_4126_0 & ~i_10_258_2379_0 & ~i_10_258_2380_0))) | (~i_10_258_2353_0 & ((~i_10_258_2331_0 & ~i_10_258_2700_0 & ~i_10_258_3043_0 & ~i_10_258_3468_0 & ~i_10_258_3495_0 & ~i_10_258_4123_0) | (i_10_258_1655_0 & ~i_10_258_4126_0 & ~i_10_258_4564_0))) | (i_10_258_2322_0 & i_10_258_3610_0 & ~i_10_258_4126_0) | (~i_10_258_2638_0 & i_10_258_3836_0 & i_10_258_3856_0) | (i_10_258_2356_0 & i_10_258_2461_0 & ~i_10_258_4566_0) | (i_10_258_1654_0 & ~i_10_258_2700_0 & ~i_10_258_3651_0 & ~i_10_258_4269_0 & ~i_10_258_4568_0));
endmodule



// Benchmark "kernel_10_259" written by ABC on Sun Jul 19 10:25:29 2020

module kernel_10_259 ( 
    i_10_259_119_0, i_10_259_174_0, i_10_259_331_0, i_10_259_332_0,
    i_10_259_361_0, i_10_259_409_0, i_10_259_446_0, i_10_259_519_0,
    i_10_259_895_0, i_10_259_906_0, i_10_259_951_0, i_10_259_1039_0,
    i_10_259_1041_0, i_10_259_1042_0, i_10_259_1122_0, i_10_259_1204_0,
    i_10_259_1241_0, i_10_259_1266_0, i_10_259_1267_0, i_10_259_1271_0,
    i_10_259_1308_0, i_10_259_1309_0, i_10_259_1311_0, i_10_259_1312_0,
    i_10_259_1353_0, i_10_259_1354_0, i_10_259_1546_0, i_10_259_1647_0,
    i_10_259_1651_0, i_10_259_1654_0, i_10_259_1824_0, i_10_259_1911_0,
    i_10_259_1912_0, i_10_259_1950_0, i_10_259_2002_0, i_10_259_2326_0,
    i_10_259_2355_0, i_10_259_2356_0, i_10_259_2357_0, i_10_259_2454_0,
    i_10_259_2467_0, i_10_259_2515_0, i_10_259_2607_0, i_10_259_2630_0,
    i_10_259_2632_0, i_10_259_2655_0, i_10_259_2656_0, i_10_259_2676_0,
    i_10_259_2679_0, i_10_259_2703_0, i_10_259_2704_0, i_10_259_2722_0,
    i_10_259_2733_0, i_10_259_2784_0, i_10_259_2788_0, i_10_259_2820_0,
    i_10_259_2823_0, i_10_259_2833_0, i_10_259_2834_0, i_10_259_2883_0,
    i_10_259_2919_0, i_10_259_2955_0, i_10_259_2985_0, i_10_259_2986_0,
    i_10_259_3088_0, i_10_259_3163_0, i_10_259_3272_0, i_10_259_3297_0,
    i_10_259_3388_0, i_10_259_3406_0, i_10_259_3407_0, i_10_259_3433_0,
    i_10_259_3434_0, i_10_259_3450_0, i_10_259_3496_0, i_10_259_3614_0,
    i_10_259_3700_0, i_10_259_3723_0, i_10_259_3834_0, i_10_259_3852_0,
    i_10_259_3859_0, i_10_259_3860_0, i_10_259_3894_0, i_10_259_3895_0,
    i_10_259_3896_0, i_10_259_3964_0, i_10_259_3980_0, i_10_259_3981_0,
    i_10_259_3982_0, i_10_259_3987_0, i_10_259_4116_0, i_10_259_4129_0,
    i_10_259_4130_0, i_10_259_4281_0, i_10_259_4282_0, i_10_259_4285_0,
    i_10_259_4288_0, i_10_259_4291_0, i_10_259_4292_0, i_10_259_4579_0,
    o_10_259_0_0  );
  input  i_10_259_119_0, i_10_259_174_0, i_10_259_331_0, i_10_259_332_0,
    i_10_259_361_0, i_10_259_409_0, i_10_259_446_0, i_10_259_519_0,
    i_10_259_895_0, i_10_259_906_0, i_10_259_951_0, i_10_259_1039_0,
    i_10_259_1041_0, i_10_259_1042_0, i_10_259_1122_0, i_10_259_1204_0,
    i_10_259_1241_0, i_10_259_1266_0, i_10_259_1267_0, i_10_259_1271_0,
    i_10_259_1308_0, i_10_259_1309_0, i_10_259_1311_0, i_10_259_1312_0,
    i_10_259_1353_0, i_10_259_1354_0, i_10_259_1546_0, i_10_259_1647_0,
    i_10_259_1651_0, i_10_259_1654_0, i_10_259_1824_0, i_10_259_1911_0,
    i_10_259_1912_0, i_10_259_1950_0, i_10_259_2002_0, i_10_259_2326_0,
    i_10_259_2355_0, i_10_259_2356_0, i_10_259_2357_0, i_10_259_2454_0,
    i_10_259_2467_0, i_10_259_2515_0, i_10_259_2607_0, i_10_259_2630_0,
    i_10_259_2632_0, i_10_259_2655_0, i_10_259_2656_0, i_10_259_2676_0,
    i_10_259_2679_0, i_10_259_2703_0, i_10_259_2704_0, i_10_259_2722_0,
    i_10_259_2733_0, i_10_259_2784_0, i_10_259_2788_0, i_10_259_2820_0,
    i_10_259_2823_0, i_10_259_2833_0, i_10_259_2834_0, i_10_259_2883_0,
    i_10_259_2919_0, i_10_259_2955_0, i_10_259_2985_0, i_10_259_2986_0,
    i_10_259_3088_0, i_10_259_3163_0, i_10_259_3272_0, i_10_259_3297_0,
    i_10_259_3388_0, i_10_259_3406_0, i_10_259_3407_0, i_10_259_3433_0,
    i_10_259_3434_0, i_10_259_3450_0, i_10_259_3496_0, i_10_259_3614_0,
    i_10_259_3700_0, i_10_259_3723_0, i_10_259_3834_0, i_10_259_3852_0,
    i_10_259_3859_0, i_10_259_3860_0, i_10_259_3894_0, i_10_259_3895_0,
    i_10_259_3896_0, i_10_259_3964_0, i_10_259_3980_0, i_10_259_3981_0,
    i_10_259_3982_0, i_10_259_3987_0, i_10_259_4116_0, i_10_259_4129_0,
    i_10_259_4130_0, i_10_259_4281_0, i_10_259_4282_0, i_10_259_4285_0,
    i_10_259_4288_0, i_10_259_4291_0, i_10_259_4292_0, i_10_259_4579_0;
  output o_10_259_0_0;
  assign o_10_259_0_0 = 0;
endmodule



// Benchmark "kernel_10_260" written by ABC on Sun Jul 19 10:25:30 2020

module kernel_10_260 ( 
    i_10_260_28_0, i_10_260_55_0, i_10_260_56_0, i_10_260_250_0,
    i_10_260_251_0, i_10_260_282_0, i_10_260_294_0, i_10_260_321_0,
    i_10_260_322_0, i_10_260_430_0, i_10_260_431_0, i_10_260_463_0,
    i_10_260_517_0, i_10_260_593_0, i_10_260_706_0, i_10_260_797_0,
    i_10_260_799_0, i_10_260_876_0, i_10_260_898_0, i_10_260_906_0,
    i_10_260_921_0, i_10_260_930_0, i_10_260_945_0, i_10_260_969_0,
    i_10_260_1029_0, i_10_260_1165_0, i_10_260_1237_0, i_10_260_1238_0,
    i_10_260_1239_0, i_10_260_1347_0, i_10_260_1364_0, i_10_260_1369_0,
    i_10_260_1385_0, i_10_260_1489_0, i_10_260_1543_0, i_10_260_1546_0,
    i_10_260_1547_0, i_10_260_1628_0, i_10_260_1630_0, i_10_260_1695_0,
    i_10_260_1718_0, i_10_260_1908_0, i_10_260_1996_0, i_10_260_2023_0,
    i_10_260_2326_0, i_10_260_2353_0, i_10_260_2356_0, i_10_260_2357_0,
    i_10_260_2568_0, i_10_260_2571_0, i_10_260_2608_0, i_10_260_2609_0,
    i_10_260_2632_0, i_10_260_2679_0, i_10_260_2691_0, i_10_260_2694_0,
    i_10_260_2695_0, i_10_260_2710_0, i_10_260_2716_0, i_10_260_2782_0,
    i_10_260_2788_0, i_10_260_2789_0, i_10_260_2828_0, i_10_260_2830_0,
    i_10_260_2850_0, i_10_260_2851_0, i_10_260_2921_0, i_10_260_2982_0,
    i_10_260_3072_0, i_10_260_3073_0, i_10_260_3076_0, i_10_260_3093_0,
    i_10_260_3271_0, i_10_260_3293_0, i_10_260_3301_0, i_10_260_3359_0,
    i_10_260_3390_0, i_10_260_3391_0, i_10_260_3434_0, i_10_260_3561_0,
    i_10_260_3582_0, i_10_260_3583_0, i_10_260_3590_0, i_10_260_3784_0,
    i_10_260_3813_0, i_10_260_3815_0, i_10_260_3855_0, i_10_260_3856_0,
    i_10_260_3877_0, i_10_260_3889_0, i_10_260_3945_0, i_10_260_4031_0,
    i_10_260_4119_0, i_10_260_4173_0, i_10_260_4236_0, i_10_260_4266_0,
    i_10_260_4278_0, i_10_260_4281_0, i_10_260_4461_0, i_10_260_4566_0,
    o_10_260_0_0  );
  input  i_10_260_28_0, i_10_260_55_0, i_10_260_56_0, i_10_260_250_0,
    i_10_260_251_0, i_10_260_282_0, i_10_260_294_0, i_10_260_321_0,
    i_10_260_322_0, i_10_260_430_0, i_10_260_431_0, i_10_260_463_0,
    i_10_260_517_0, i_10_260_593_0, i_10_260_706_0, i_10_260_797_0,
    i_10_260_799_0, i_10_260_876_0, i_10_260_898_0, i_10_260_906_0,
    i_10_260_921_0, i_10_260_930_0, i_10_260_945_0, i_10_260_969_0,
    i_10_260_1029_0, i_10_260_1165_0, i_10_260_1237_0, i_10_260_1238_0,
    i_10_260_1239_0, i_10_260_1347_0, i_10_260_1364_0, i_10_260_1369_0,
    i_10_260_1385_0, i_10_260_1489_0, i_10_260_1543_0, i_10_260_1546_0,
    i_10_260_1547_0, i_10_260_1628_0, i_10_260_1630_0, i_10_260_1695_0,
    i_10_260_1718_0, i_10_260_1908_0, i_10_260_1996_0, i_10_260_2023_0,
    i_10_260_2326_0, i_10_260_2353_0, i_10_260_2356_0, i_10_260_2357_0,
    i_10_260_2568_0, i_10_260_2571_0, i_10_260_2608_0, i_10_260_2609_0,
    i_10_260_2632_0, i_10_260_2679_0, i_10_260_2691_0, i_10_260_2694_0,
    i_10_260_2695_0, i_10_260_2710_0, i_10_260_2716_0, i_10_260_2782_0,
    i_10_260_2788_0, i_10_260_2789_0, i_10_260_2828_0, i_10_260_2830_0,
    i_10_260_2850_0, i_10_260_2851_0, i_10_260_2921_0, i_10_260_2982_0,
    i_10_260_3072_0, i_10_260_3073_0, i_10_260_3076_0, i_10_260_3093_0,
    i_10_260_3271_0, i_10_260_3293_0, i_10_260_3301_0, i_10_260_3359_0,
    i_10_260_3390_0, i_10_260_3391_0, i_10_260_3434_0, i_10_260_3561_0,
    i_10_260_3582_0, i_10_260_3583_0, i_10_260_3590_0, i_10_260_3784_0,
    i_10_260_3813_0, i_10_260_3815_0, i_10_260_3855_0, i_10_260_3856_0,
    i_10_260_3877_0, i_10_260_3889_0, i_10_260_3945_0, i_10_260_4031_0,
    i_10_260_4119_0, i_10_260_4173_0, i_10_260_4236_0, i_10_260_4266_0,
    i_10_260_4278_0, i_10_260_4281_0, i_10_260_4461_0, i_10_260_4566_0;
  output o_10_260_0_0;
  assign o_10_260_0_0 = 0;
endmodule



// Benchmark "kernel_10_261" written by ABC on Sun Jul 19 10:25:31 2020

module kernel_10_261 ( 
    i_10_261_123_0, i_10_261_148_0, i_10_261_178_0, i_10_261_267_0,
    i_10_261_277_0, i_10_261_282_0, i_10_261_283_0, i_10_261_292_0,
    i_10_261_408_0, i_10_261_510_0, i_10_261_520_0, i_10_261_663_0,
    i_10_261_1005_0, i_10_261_1006_0, i_10_261_1236_0, i_10_261_1266_0,
    i_10_261_1309_0, i_10_261_1312_0, i_10_261_1437_0, i_10_261_1438_0,
    i_10_261_1546_0, i_10_261_1552_0, i_10_261_1555_0, i_10_261_1579_0,
    i_10_261_1626_0, i_10_261_1689_0, i_10_261_1716_0, i_10_261_1734_0,
    i_10_261_1735_0, i_10_261_1806_0, i_10_261_1951_0, i_10_261_1992_0,
    i_10_261_2031_0, i_10_261_2311_0, i_10_261_2353_0, i_10_261_2355_0,
    i_10_261_2356_0, i_10_261_2408_0, i_10_261_2453_0, i_10_261_2469_0,
    i_10_261_2472_0, i_10_261_2571_0, i_10_261_2632_0, i_10_261_2662_0,
    i_10_261_2663_0, i_10_261_2715_0, i_10_261_2716_0, i_10_261_2730_0,
    i_10_261_2731_0, i_10_261_2734_0, i_10_261_2785_0, i_10_261_2827_0,
    i_10_261_2850_0, i_10_261_2884_0, i_10_261_2887_0, i_10_261_2922_0,
    i_10_261_2967_0, i_10_261_2985_0, i_10_261_3045_0, i_10_261_3072_0,
    i_10_261_3075_0, i_10_261_3196_0, i_10_261_3199_0, i_10_261_3201_0,
    i_10_261_3278_0, i_10_261_3279_0, i_10_261_3283_0, i_10_261_3318_0,
    i_10_261_3386_0, i_10_261_3391_0, i_10_261_3471_0, i_10_261_3507_0,
    i_10_261_3525_0, i_10_261_3540_0, i_10_261_3585_0, i_10_261_3613_0,
    i_10_261_3616_0, i_10_261_3688_0, i_10_261_3782_0, i_10_261_3783_0,
    i_10_261_3784_0, i_10_261_3787_0, i_10_261_3811_0, i_10_261_3837_0,
    i_10_261_3838_0, i_10_261_3846_0, i_10_261_3859_0, i_10_261_3909_0,
    i_10_261_3985_0, i_10_261_4056_0, i_10_261_4116_0, i_10_261_4117_0,
    i_10_261_4120_0, i_10_261_4121_0, i_10_261_4173_0, i_10_261_4272_0,
    i_10_261_4273_0, i_10_261_4281_0, i_10_261_4282_0, i_10_261_4290_0,
    o_10_261_0_0  );
  input  i_10_261_123_0, i_10_261_148_0, i_10_261_178_0, i_10_261_267_0,
    i_10_261_277_0, i_10_261_282_0, i_10_261_283_0, i_10_261_292_0,
    i_10_261_408_0, i_10_261_510_0, i_10_261_520_0, i_10_261_663_0,
    i_10_261_1005_0, i_10_261_1006_0, i_10_261_1236_0, i_10_261_1266_0,
    i_10_261_1309_0, i_10_261_1312_0, i_10_261_1437_0, i_10_261_1438_0,
    i_10_261_1546_0, i_10_261_1552_0, i_10_261_1555_0, i_10_261_1579_0,
    i_10_261_1626_0, i_10_261_1689_0, i_10_261_1716_0, i_10_261_1734_0,
    i_10_261_1735_0, i_10_261_1806_0, i_10_261_1951_0, i_10_261_1992_0,
    i_10_261_2031_0, i_10_261_2311_0, i_10_261_2353_0, i_10_261_2355_0,
    i_10_261_2356_0, i_10_261_2408_0, i_10_261_2453_0, i_10_261_2469_0,
    i_10_261_2472_0, i_10_261_2571_0, i_10_261_2632_0, i_10_261_2662_0,
    i_10_261_2663_0, i_10_261_2715_0, i_10_261_2716_0, i_10_261_2730_0,
    i_10_261_2731_0, i_10_261_2734_0, i_10_261_2785_0, i_10_261_2827_0,
    i_10_261_2850_0, i_10_261_2884_0, i_10_261_2887_0, i_10_261_2922_0,
    i_10_261_2967_0, i_10_261_2985_0, i_10_261_3045_0, i_10_261_3072_0,
    i_10_261_3075_0, i_10_261_3196_0, i_10_261_3199_0, i_10_261_3201_0,
    i_10_261_3278_0, i_10_261_3279_0, i_10_261_3283_0, i_10_261_3318_0,
    i_10_261_3386_0, i_10_261_3391_0, i_10_261_3471_0, i_10_261_3507_0,
    i_10_261_3525_0, i_10_261_3540_0, i_10_261_3585_0, i_10_261_3613_0,
    i_10_261_3616_0, i_10_261_3688_0, i_10_261_3782_0, i_10_261_3783_0,
    i_10_261_3784_0, i_10_261_3787_0, i_10_261_3811_0, i_10_261_3837_0,
    i_10_261_3838_0, i_10_261_3846_0, i_10_261_3859_0, i_10_261_3909_0,
    i_10_261_3985_0, i_10_261_4056_0, i_10_261_4116_0, i_10_261_4117_0,
    i_10_261_4120_0, i_10_261_4121_0, i_10_261_4173_0, i_10_261_4272_0,
    i_10_261_4273_0, i_10_261_4281_0, i_10_261_4282_0, i_10_261_4290_0;
  output o_10_261_0_0;
  assign o_10_261_0_0 = ~((~i_10_261_282_0 & i_10_261_3985_0 & ((~i_10_261_1236_0 & ~i_10_261_2355_0 & ~i_10_261_2408_0 & ~i_10_261_2734_0) | (~i_10_261_283_0 & ~i_10_261_1689_0 & ~i_10_261_2715_0 & ~i_10_261_2827_0 & ~i_10_261_3507_0))) | (~i_10_261_1005_0 & ((~i_10_261_1437_0 & ~i_10_261_1626_0 & ~i_10_261_2715_0) | (~i_10_261_267_0 & ~i_10_261_1546_0 & ~i_10_261_3199_0 & ~i_10_261_4272_0 & ~i_10_261_4282_0))) | (~i_10_261_2571_0 & ((~i_10_261_267_0 & ((~i_10_261_148_0 & ~i_10_261_408_0 & ~i_10_261_1552_0 & ~i_10_261_1555_0 & ~i_10_261_2031_0 & i_10_261_2734_0) | (~i_10_261_2408_0 & ~i_10_261_3283_0 & ~i_10_261_3507_0 & ~i_10_261_3985_0))) | (i_10_261_2353_0 & i_10_261_2731_0 & ~i_10_261_2922_0 & ~i_10_261_3075_0 & ~i_10_261_3782_0))) | (i_10_261_3199_0 & ((~i_10_261_3283_0 & ~i_10_261_3540_0) | (~i_10_261_2469_0 & ~i_10_261_3782_0))) | (~i_10_261_3837_0 & ((~i_10_261_1006_0 & ~i_10_261_2356_0 & i_10_261_2827_0 & ~i_10_261_3283_0) | (~i_10_261_1735_0 & ~i_10_261_2311_0 & i_10_261_3688_0))) | (~i_10_261_4281_0 & ((~i_10_261_1555_0 & ~i_10_261_2884_0 & ~i_10_261_3279_0) | (~i_10_261_520_0 & ~i_10_261_2355_0 & i_10_261_3283_0 & ~i_10_261_3318_0 & ~i_10_261_3616_0 & i_10_261_3838_0))) | (i_10_261_3196_0 & i_10_261_3616_0));
endmodule



// Benchmark "kernel_10_262" written by ABC on Sun Jul 19 10:25:32 2020

module kernel_10_262 ( 
    i_10_262_319_0, i_10_262_390_0, i_10_262_408_0, i_10_262_409_0,
    i_10_262_410_0, i_10_262_411_0, i_10_262_413_0, i_10_262_441_0,
    i_10_262_444_0, i_10_262_499_0, i_10_262_586_0, i_10_262_736_0,
    i_10_262_737_0, i_10_262_797_0, i_10_262_853_0, i_10_262_931_0,
    i_10_262_1034_0, i_10_262_1119_0, i_10_262_1181_0, i_10_262_1239_0,
    i_10_262_1240_0, i_10_262_1241_0, i_10_262_1276_0, i_10_262_1308_0,
    i_10_262_1347_0, i_10_262_1438_0, i_10_262_1439_0, i_10_262_1545_0,
    i_10_262_1552_0, i_10_262_1579_0, i_10_262_1583_0, i_10_262_1650_0,
    i_10_262_1651_0, i_10_262_1766_0, i_10_262_1804_0, i_10_262_1807_0,
    i_10_262_1819_0, i_10_262_1821_0, i_10_262_1822_0, i_10_262_2200_0,
    i_10_262_2223_0, i_10_262_2355_0, i_10_262_2356_0, i_10_262_2380_0,
    i_10_262_2389_0, i_10_262_2391_0, i_10_262_2392_0, i_10_262_2410_0,
    i_10_262_2435_0, i_10_262_2441_0, i_10_262_2443_0, i_10_262_2444_0,
    i_10_262_2450_0, i_10_262_2452_0, i_10_262_2459_0, i_10_262_2635_0,
    i_10_262_2650_0, i_10_262_2658_0, i_10_262_2660_0, i_10_262_2679_0,
    i_10_262_2695_0, i_10_262_2704_0, i_10_262_2716_0, i_10_262_2733_0,
    i_10_262_2734_0, i_10_262_2784_0, i_10_262_2821_0, i_10_262_2884_0,
    i_10_262_2888_0, i_10_262_2983_0, i_10_262_3072_0, i_10_262_3075_0,
    i_10_262_3076_0, i_10_262_3117_0, i_10_262_3166_0, i_10_262_3202_0,
    i_10_262_3468_0, i_10_262_3471_0, i_10_262_3539_0, i_10_262_3541_0,
    i_10_262_3544_0, i_10_262_3609_0, i_10_262_3684_0, i_10_262_3775_0,
    i_10_262_3805_0, i_10_262_3840_0, i_10_262_3846_0, i_10_262_3857_0,
    i_10_262_3893_0, i_10_262_4013_0, i_10_262_4173_0, i_10_262_4175_0,
    i_10_262_4182_0, i_10_262_4475_0, i_10_262_4524_0, i_10_262_4563_0,
    i_10_262_4564_0, i_10_262_4568_0, i_10_262_4588_0, i_10_262_4598_0,
    o_10_262_0_0  );
  input  i_10_262_319_0, i_10_262_390_0, i_10_262_408_0, i_10_262_409_0,
    i_10_262_410_0, i_10_262_411_0, i_10_262_413_0, i_10_262_441_0,
    i_10_262_444_0, i_10_262_499_0, i_10_262_586_0, i_10_262_736_0,
    i_10_262_737_0, i_10_262_797_0, i_10_262_853_0, i_10_262_931_0,
    i_10_262_1034_0, i_10_262_1119_0, i_10_262_1181_0, i_10_262_1239_0,
    i_10_262_1240_0, i_10_262_1241_0, i_10_262_1276_0, i_10_262_1308_0,
    i_10_262_1347_0, i_10_262_1438_0, i_10_262_1439_0, i_10_262_1545_0,
    i_10_262_1552_0, i_10_262_1579_0, i_10_262_1583_0, i_10_262_1650_0,
    i_10_262_1651_0, i_10_262_1766_0, i_10_262_1804_0, i_10_262_1807_0,
    i_10_262_1819_0, i_10_262_1821_0, i_10_262_1822_0, i_10_262_2200_0,
    i_10_262_2223_0, i_10_262_2355_0, i_10_262_2356_0, i_10_262_2380_0,
    i_10_262_2389_0, i_10_262_2391_0, i_10_262_2392_0, i_10_262_2410_0,
    i_10_262_2435_0, i_10_262_2441_0, i_10_262_2443_0, i_10_262_2444_0,
    i_10_262_2450_0, i_10_262_2452_0, i_10_262_2459_0, i_10_262_2635_0,
    i_10_262_2650_0, i_10_262_2658_0, i_10_262_2660_0, i_10_262_2679_0,
    i_10_262_2695_0, i_10_262_2704_0, i_10_262_2716_0, i_10_262_2733_0,
    i_10_262_2734_0, i_10_262_2784_0, i_10_262_2821_0, i_10_262_2884_0,
    i_10_262_2888_0, i_10_262_2983_0, i_10_262_3072_0, i_10_262_3075_0,
    i_10_262_3076_0, i_10_262_3117_0, i_10_262_3166_0, i_10_262_3202_0,
    i_10_262_3468_0, i_10_262_3471_0, i_10_262_3539_0, i_10_262_3541_0,
    i_10_262_3544_0, i_10_262_3609_0, i_10_262_3684_0, i_10_262_3775_0,
    i_10_262_3805_0, i_10_262_3840_0, i_10_262_3846_0, i_10_262_3857_0,
    i_10_262_3893_0, i_10_262_4013_0, i_10_262_4173_0, i_10_262_4175_0,
    i_10_262_4182_0, i_10_262_4475_0, i_10_262_4524_0, i_10_262_4563_0,
    i_10_262_4564_0, i_10_262_4568_0, i_10_262_4588_0, i_10_262_4598_0;
  output o_10_262_0_0;
  assign o_10_262_0_0 = 0;
endmodule



// Benchmark "kernel_10_263" written by ABC on Sun Jul 19 10:25:33 2020

module kernel_10_263 ( 
    i_10_263_243_0, i_10_263_283_0, i_10_263_444_0, i_10_263_459_0,
    i_10_263_460_0, i_10_263_464_0, i_10_263_751_0, i_10_263_793_0,
    i_10_263_795_0, i_10_263_966_0, i_10_263_968_0, i_10_263_999_0,
    i_10_263_1000_0, i_10_263_1041_0, i_10_263_1235_0, i_10_263_1236_0,
    i_10_263_1243_0, i_10_263_1246_0, i_10_263_1247_0, i_10_263_1249_0,
    i_10_263_1445_0, i_10_263_1539_0, i_10_263_1541_0, i_10_263_1819_0,
    i_10_263_1821_0, i_10_263_1823_0, i_10_263_1911_0, i_10_263_1912_0,
    i_10_263_1913_0, i_10_263_2004_0, i_10_263_2179_0, i_10_263_2180_0,
    i_10_263_2354_0, i_10_263_2377_0, i_10_263_2467_0, i_10_263_2473_0,
    i_10_263_2628_0, i_10_263_2630_0, i_10_263_2631_0, i_10_263_2634_0,
    i_10_263_2655_0, i_10_263_2657_0, i_10_263_2658_0, i_10_263_2660_0,
    i_10_263_2680_0, i_10_263_2681_0, i_10_263_2700_0, i_10_263_2701_0,
    i_10_263_2720_0, i_10_263_2721_0, i_10_263_2722_0, i_10_263_2727_0,
    i_10_263_2728_0, i_10_263_2732_0, i_10_263_2733_0, i_10_263_2735_0,
    i_10_263_2818_0, i_10_263_2827_0, i_10_263_2829_0, i_10_263_2830_0,
    i_10_263_2833_0, i_10_263_2883_0, i_10_263_2884_0, i_10_263_2919_0,
    i_10_263_2920_0, i_10_263_3034_0, i_10_263_3038_0, i_10_263_3069_0,
    i_10_263_3070_0, i_10_263_3071_0, i_10_263_3087_0, i_10_263_3198_0,
    i_10_263_3268_0, i_10_263_3270_0, i_10_263_3385_0, i_10_263_3388_0,
    i_10_263_3389_0, i_10_263_3469_0, i_10_263_3537_0, i_10_263_3589_0,
    i_10_263_3612_0, i_10_263_3681_0, i_10_263_3687_0, i_10_263_3781_0,
    i_10_263_3787_0, i_10_263_3852_0, i_10_263_3853_0, i_10_263_3854_0,
    i_10_263_3860_0, i_10_263_3888_0, i_10_263_3889_0, i_10_263_3912_0,
    i_10_263_3978_0, i_10_263_3990_0, i_10_263_3991_0, i_10_263_4266_0,
    i_10_263_4267_0, i_10_263_4290_0, i_10_263_4429_0, i_10_263_4571_0,
    o_10_263_0_0  );
  input  i_10_263_243_0, i_10_263_283_0, i_10_263_444_0, i_10_263_459_0,
    i_10_263_460_0, i_10_263_464_0, i_10_263_751_0, i_10_263_793_0,
    i_10_263_795_0, i_10_263_966_0, i_10_263_968_0, i_10_263_999_0,
    i_10_263_1000_0, i_10_263_1041_0, i_10_263_1235_0, i_10_263_1236_0,
    i_10_263_1243_0, i_10_263_1246_0, i_10_263_1247_0, i_10_263_1249_0,
    i_10_263_1445_0, i_10_263_1539_0, i_10_263_1541_0, i_10_263_1819_0,
    i_10_263_1821_0, i_10_263_1823_0, i_10_263_1911_0, i_10_263_1912_0,
    i_10_263_1913_0, i_10_263_2004_0, i_10_263_2179_0, i_10_263_2180_0,
    i_10_263_2354_0, i_10_263_2377_0, i_10_263_2467_0, i_10_263_2473_0,
    i_10_263_2628_0, i_10_263_2630_0, i_10_263_2631_0, i_10_263_2634_0,
    i_10_263_2655_0, i_10_263_2657_0, i_10_263_2658_0, i_10_263_2660_0,
    i_10_263_2680_0, i_10_263_2681_0, i_10_263_2700_0, i_10_263_2701_0,
    i_10_263_2720_0, i_10_263_2721_0, i_10_263_2722_0, i_10_263_2727_0,
    i_10_263_2728_0, i_10_263_2732_0, i_10_263_2733_0, i_10_263_2735_0,
    i_10_263_2818_0, i_10_263_2827_0, i_10_263_2829_0, i_10_263_2830_0,
    i_10_263_2833_0, i_10_263_2883_0, i_10_263_2884_0, i_10_263_2919_0,
    i_10_263_2920_0, i_10_263_3034_0, i_10_263_3038_0, i_10_263_3069_0,
    i_10_263_3070_0, i_10_263_3071_0, i_10_263_3087_0, i_10_263_3198_0,
    i_10_263_3268_0, i_10_263_3270_0, i_10_263_3385_0, i_10_263_3388_0,
    i_10_263_3389_0, i_10_263_3469_0, i_10_263_3537_0, i_10_263_3589_0,
    i_10_263_3612_0, i_10_263_3681_0, i_10_263_3687_0, i_10_263_3781_0,
    i_10_263_3787_0, i_10_263_3852_0, i_10_263_3853_0, i_10_263_3854_0,
    i_10_263_3860_0, i_10_263_3888_0, i_10_263_3889_0, i_10_263_3912_0,
    i_10_263_3978_0, i_10_263_3990_0, i_10_263_3991_0, i_10_263_4266_0,
    i_10_263_4267_0, i_10_263_4290_0, i_10_263_4429_0, i_10_263_4571_0;
  output o_10_263_0_0;
  assign o_10_263_0_0 = ~((~i_10_263_3069_0 & ((i_10_263_283_0 & ((~i_10_263_968_0 & ~i_10_263_1445_0 & ~i_10_263_2377_0 & ~i_10_263_2733_0 & ~i_10_263_2884_0 & ~i_10_263_3537_0 & ~i_10_263_3889_0) | (~i_10_263_2473_0 & ~i_10_263_2829_0 & ~i_10_263_3469_0 & ~i_10_263_3991_0))) | (~i_10_263_966_0 & ((~i_10_263_968_0 & ~i_10_263_3888_0 & ~i_10_263_3991_0 & ((~i_10_263_444_0 & ~i_10_263_999_0 & ~i_10_263_2004_0 & ~i_10_263_2179_0 & ~i_10_263_2473_0 & ~i_10_263_3589_0 & ~i_10_263_3612_0) | (~i_10_263_1821_0 & ~i_10_263_2377_0 & ~i_10_263_2660_0 & ~i_10_263_2680_0 & ~i_10_263_2728_0 & ~i_10_263_3852_0 & ~i_10_263_3912_0))) | (~i_10_263_2377_0 & ~i_10_263_2680_0 & ~i_10_263_2681_0 & ~i_10_263_2833_0 & ~i_10_263_2883_0 & ~i_10_263_2884_0 & ~i_10_263_3070_0 & ~i_10_263_3071_0 & ~i_10_263_3589_0 & ~i_10_263_3681_0 & ~i_10_263_3860_0 & ~i_10_263_3889_0 & ~i_10_263_3912_0 & ~i_10_263_3978_0))) | (~i_10_263_999_0 & ((i_10_263_1819_0 & ~i_10_263_2354_0 & ~i_10_263_2630_0 & ~i_10_263_2655_0 & ~i_10_263_2884_0 & ~i_10_263_3469_0 & ~i_10_263_3681_0 & ~i_10_263_3888_0) | (~i_10_263_1246_0 & ~i_10_263_2004_0 & ~i_10_263_2681_0 & ~i_10_263_3268_0 & i_10_263_3852_0 & ~i_10_263_3912_0 & ~i_10_263_3991_0))) | (i_10_263_1235_0 & ~i_10_263_1821_0 & ~i_10_263_3268_0 & ~i_10_263_3681_0 & ~i_10_263_4290_0))) | (~i_10_263_283_0 & ((~i_10_263_464_0 & ~i_10_263_2631_0 & ~i_10_263_2733_0 & ~i_10_263_2883_0 & i_10_263_3389_0) | (~i_10_263_444_0 & ~i_10_263_1912_0 & i_10_263_2658_0 & ~i_10_263_2735_0 & ~i_10_263_2884_0 & i_10_263_3612_0))) | (~i_10_263_2004_0 & ((~i_10_263_2919_0 & ((~i_10_263_459_0 & ~i_10_263_3537_0 & ((~i_10_263_795_0 & ~i_10_263_1821_0 & ~i_10_263_1823_0 & ~i_10_263_2179_0 & ~i_10_263_2680_0 & ~i_10_263_2829_0 & ~i_10_263_3198_0 & ~i_10_263_3853_0 & ~i_10_263_3888_0) | (i_10_263_2728_0 & ~i_10_263_3385_0 & ~i_10_263_3612_0 & ~i_10_263_3990_0))) | (~i_10_263_464_0 & ~i_10_263_2473_0 & ~i_10_263_2701_0 & ~i_10_263_3038_0 & ~i_10_263_3469_0 & ~i_10_263_3681_0 & ~i_10_263_3889_0 & ~i_10_263_3978_0 & ~i_10_263_3990_0 & ~i_10_263_3991_0))) | (~i_10_263_999_0 & ~i_10_263_3991_0 & ((~i_10_263_3198_0 & ~i_10_263_3681_0 & i_10_263_3853_0) | (~i_10_263_966_0 & ~i_10_263_1235_0 & ~i_10_263_1539_0 & ~i_10_263_2884_0 & ~i_10_263_2920_0 & ~i_10_263_3589_0 & ~i_10_263_3889_0 & ~i_10_263_3990_0))) | (~i_10_263_3681_0 & ((~i_10_263_1000_0 & ~i_10_263_1823_0 & ~i_10_263_2883_0 & ~i_10_263_3537_0 & ~i_10_263_3612_0 & i_10_263_3853_0 & ~i_10_263_3888_0) | (~i_10_263_968_0 & ~i_10_263_1539_0 & ~i_10_263_1821_0 & ~i_10_263_2721_0 & ~i_10_263_2884_0 & ~i_10_263_3087_0 & ~i_10_263_3198_0 & ~i_10_263_3889_0 & ~i_10_263_4267_0))))) | (~i_10_263_2919_0 & ((i_10_263_460_0 & ((~i_10_263_966_0 & ~i_10_263_968_0 & ~i_10_263_2727_0 & ~i_10_263_2818_0 & ~i_10_263_3038_0 & ~i_10_263_3912_0 & ~i_10_263_3978_0 & ~i_10_263_3990_0) | (~i_10_263_1539_0 & ~i_10_263_2354_0 & ~i_10_263_2680_0 & ~i_10_263_3681_0 & ~i_10_263_3889_0 & ~i_10_263_3991_0))) | (i_10_263_793_0 & ~i_10_263_1235_0 & ~i_10_263_2180_0 & ~i_10_263_2634_0 & ~i_10_263_2884_0 & ~i_10_263_3270_0 & ~i_10_263_3537_0 & ~i_10_263_3681_0 & ~i_10_263_3888_0))) | (~i_10_263_3990_0 & ((~i_10_263_999_0 & ((~i_10_263_1236_0 & ~i_10_263_1821_0 & i_10_263_2827_0 & ~i_10_263_3537_0) | (~i_10_263_966_0 & ~i_10_263_968_0 & ~i_10_263_1243_0 & ~i_10_263_2700_0 & ~i_10_263_2735_0 & ~i_10_263_2818_0 & ~i_10_263_2883_0 & ~i_10_263_3198_0 & ~i_10_263_3853_0 & ~i_10_263_3978_0))) | (~i_10_263_3681_0 & ~i_10_263_3889_0 & ((~i_10_263_1236_0 & ~i_10_263_2180_0 & ~i_10_263_2680_0 & ~i_10_263_2720_0 & ~i_10_263_2735_0 & ~i_10_263_3034_0 & ~i_10_263_3071_0 & ~i_10_263_3198_0 & ~i_10_263_3469_0 & ~i_10_263_3860_0 & ~i_10_263_3888_0 & ~i_10_263_3978_0) | (~i_10_263_2179_0 & ~i_10_263_2631_0 & ~i_10_263_2700_0 & ~i_10_263_2721_0 & ~i_10_263_2884_0 & i_10_263_2920_0 & ~i_10_263_3070_0 & ~i_10_263_3385_0 & ~i_10_263_4571_0))))) | (~i_10_263_2884_0 & ((~i_10_263_1000_0 & ((i_10_263_2630_0 & ~i_10_263_3198_0 & i_10_263_3860_0) | (~i_10_263_444_0 & ~i_10_263_1541_0 & ~i_10_263_2681_0 & ~i_10_263_2701_0 & ~i_10_263_2883_0 & ~i_10_263_2920_0 & i_10_263_3852_0 & ~i_10_263_4266_0))) | (~i_10_263_2701_0 & i_10_263_2722_0 & ~i_10_263_2735_0 & ~i_10_263_2883_0 & ~i_10_263_3070_0 & ~i_10_263_3589_0))) | (i_10_263_2722_0 & ((~i_10_263_1243_0 & ~i_10_263_2680_0 & i_10_263_2728_0 & ~i_10_263_3270_0) | (i_10_263_2634_0 & i_10_263_2829_0 & ~i_10_263_3991_0))) | (~i_10_263_2680_0 & ~i_10_263_3681_0 & ~i_10_263_3860_0 & ~i_10_263_3991_0 & ~i_10_263_4266_0 & ((~i_10_263_2354_0 & i_10_263_2728_0 & ~i_10_263_3087_0) | (~i_10_263_1235_0 & ~i_10_263_2179_0 & ~i_10_263_2473_0 & ~i_10_263_2631_0 & ~i_10_263_2830_0 & ~i_10_263_2833_0 & ~i_10_263_3034_0 & ~i_10_263_3385_0 & ~i_10_263_3912_0 & ~i_10_263_4571_0))) | (i_10_263_2377_0 & ~i_10_263_2628_0 & i_10_263_3038_0 & ~i_10_263_3268_0) | (i_10_263_999_0 & ~i_10_263_1821_0 & i_10_263_2728_0 & ~i_10_263_2733_0 & ~i_10_263_3388_0));
endmodule



// Benchmark "kernel_10_264" written by ABC on Sun Jul 19 10:25:34 2020

module kernel_10_264 ( 
    i_10_264_155_0, i_10_264_177_0, i_10_264_220_0, i_10_264_223_0,
    i_10_264_224_0, i_10_264_247_0, i_10_264_249_0, i_10_264_272_0,
    i_10_264_281_0, i_10_264_290_0, i_10_264_291_0, i_10_264_292_0,
    i_10_264_318_0, i_10_264_326_0, i_10_264_329_0, i_10_264_406_0,
    i_10_264_407_0, i_10_264_408_0, i_10_264_497_0, i_10_264_593_0,
    i_10_264_797_0, i_10_264_830_0, i_10_264_832_0, i_10_264_833_0,
    i_10_264_896_0, i_10_264_899_0, i_10_264_931_0, i_10_264_954_0,
    i_10_264_955_0, i_10_264_957_0, i_10_264_1057_0, i_10_264_1121_0,
    i_10_264_1264_0, i_10_264_1273_0, i_10_264_1305_0, i_10_264_1308_0,
    i_10_264_1345_0, i_10_264_1363_0, i_10_264_1364_0, i_10_264_1367_0,
    i_10_264_1444_0, i_10_264_1648_0, i_10_264_1651_0, i_10_264_1688_0,
    i_10_264_1724_0, i_10_264_1765_0, i_10_264_1913_0, i_10_264_1921_0,
    i_10_264_1996_0, i_10_264_1997_0, i_10_264_2023_0, i_10_264_2255_0,
    i_10_264_2310_0, i_10_264_2351_0, i_10_264_2362_0, i_10_264_2365_0,
    i_10_264_2452_0, i_10_264_2516_0, i_10_264_2518_0, i_10_264_2655_0,
    i_10_264_2656_0, i_10_264_2657_0, i_10_264_2714_0, i_10_264_2718_0,
    i_10_264_2719_0, i_10_264_2720_0, i_10_264_2731_0, i_10_264_2782_0,
    i_10_264_2784_0, i_10_264_2787_0, i_10_264_2884_0, i_10_264_2984_0,
    i_10_264_3047_0, i_10_264_3050_0, i_10_264_3077_0, i_10_264_3092_0,
    i_10_264_3281_0, i_10_264_3290_0, i_10_264_3302_0, i_10_264_3356_0,
    i_10_264_3406_0, i_10_264_3407_0, i_10_264_3494_0, i_10_264_3497_0,
    i_10_264_3526_0, i_10_264_3527_0, i_10_264_3542_0, i_10_264_3641_0,
    i_10_264_3688_0, i_10_264_3780_0, i_10_264_3852_0, i_10_264_3854_0,
    i_10_264_3984_0, i_10_264_3995_0, i_10_264_4054_0, i_10_264_4055_0,
    i_10_264_4121_0, i_10_264_4171_0, i_10_264_4237_0, i_10_264_4268_0,
    o_10_264_0_0  );
  input  i_10_264_155_0, i_10_264_177_0, i_10_264_220_0, i_10_264_223_0,
    i_10_264_224_0, i_10_264_247_0, i_10_264_249_0, i_10_264_272_0,
    i_10_264_281_0, i_10_264_290_0, i_10_264_291_0, i_10_264_292_0,
    i_10_264_318_0, i_10_264_326_0, i_10_264_329_0, i_10_264_406_0,
    i_10_264_407_0, i_10_264_408_0, i_10_264_497_0, i_10_264_593_0,
    i_10_264_797_0, i_10_264_830_0, i_10_264_832_0, i_10_264_833_0,
    i_10_264_896_0, i_10_264_899_0, i_10_264_931_0, i_10_264_954_0,
    i_10_264_955_0, i_10_264_957_0, i_10_264_1057_0, i_10_264_1121_0,
    i_10_264_1264_0, i_10_264_1273_0, i_10_264_1305_0, i_10_264_1308_0,
    i_10_264_1345_0, i_10_264_1363_0, i_10_264_1364_0, i_10_264_1367_0,
    i_10_264_1444_0, i_10_264_1648_0, i_10_264_1651_0, i_10_264_1688_0,
    i_10_264_1724_0, i_10_264_1765_0, i_10_264_1913_0, i_10_264_1921_0,
    i_10_264_1996_0, i_10_264_1997_0, i_10_264_2023_0, i_10_264_2255_0,
    i_10_264_2310_0, i_10_264_2351_0, i_10_264_2362_0, i_10_264_2365_0,
    i_10_264_2452_0, i_10_264_2516_0, i_10_264_2518_0, i_10_264_2655_0,
    i_10_264_2656_0, i_10_264_2657_0, i_10_264_2714_0, i_10_264_2718_0,
    i_10_264_2719_0, i_10_264_2720_0, i_10_264_2731_0, i_10_264_2782_0,
    i_10_264_2784_0, i_10_264_2787_0, i_10_264_2884_0, i_10_264_2984_0,
    i_10_264_3047_0, i_10_264_3050_0, i_10_264_3077_0, i_10_264_3092_0,
    i_10_264_3281_0, i_10_264_3290_0, i_10_264_3302_0, i_10_264_3356_0,
    i_10_264_3406_0, i_10_264_3407_0, i_10_264_3494_0, i_10_264_3497_0,
    i_10_264_3526_0, i_10_264_3527_0, i_10_264_3542_0, i_10_264_3641_0,
    i_10_264_3688_0, i_10_264_3780_0, i_10_264_3852_0, i_10_264_3854_0,
    i_10_264_3984_0, i_10_264_3995_0, i_10_264_4054_0, i_10_264_4055_0,
    i_10_264_4121_0, i_10_264_4171_0, i_10_264_4237_0, i_10_264_4268_0;
  output o_10_264_0_0;
  assign o_10_264_0_0 = 0;
endmodule



// Benchmark "kernel_10_265" written by ABC on Sun Jul 19 10:25:35 2020

module kernel_10_265 ( 
    i_10_265_210_0, i_10_265_277_0, i_10_265_279_0, i_10_265_280_0,
    i_10_265_287_0, i_10_265_444_0, i_10_265_447_0, i_10_265_499_0,
    i_10_265_517_0, i_10_265_586_0, i_10_265_587_0, i_10_265_607_0,
    i_10_265_792_0, i_10_265_793_0, i_10_265_796_0, i_10_265_798_0,
    i_10_265_799_0, i_10_265_904_0, i_10_265_1049_0, i_10_265_1123_0,
    i_10_265_1164_0, i_10_265_1171_0, i_10_265_1200_0, i_10_265_1201_0,
    i_10_265_1234_0, i_10_265_1305_0, i_10_265_1362_0, i_10_265_1444_0,
    i_10_265_1447_0, i_10_265_1448_0, i_10_265_1602_0, i_10_265_1651_0,
    i_10_265_1652_0, i_10_265_1732_0, i_10_265_1818_0, i_10_265_1822_0,
    i_10_265_1881_0, i_10_265_1882_0, i_10_265_2155_0, i_10_265_2329_0,
    i_10_265_2338_0, i_10_265_2362_0, i_10_265_2382_0, i_10_265_2448_0,
    i_10_265_2449_0, i_10_265_2451_0, i_10_265_2475_0, i_10_265_2543_0,
    i_10_265_2659_0, i_10_265_2660_0, i_10_265_2662_0, i_10_265_2663_0,
    i_10_265_2728_0, i_10_265_2731_0, i_10_265_2814_0, i_10_265_2888_0,
    i_10_265_2916_0, i_10_265_2917_0, i_10_265_2919_0, i_10_265_2922_0,
    i_10_265_2979_0, i_10_265_3039_0, i_10_265_3047_0, i_10_265_3049_0,
    i_10_265_3050_0, i_10_265_3092_0, i_10_265_3109_0, i_10_265_3169_0,
    i_10_265_3172_0, i_10_265_3282_0, i_10_265_3294_0, i_10_265_3388_0,
    i_10_265_3496_0, i_10_265_3615_0, i_10_265_3684_0, i_10_265_3720_0,
    i_10_265_3721_0, i_10_265_3729_0, i_10_265_3787_0, i_10_265_3851_0,
    i_10_265_3854_0, i_10_265_3859_0, i_10_265_3892_0, i_10_265_3919_0,
    i_10_265_3950_0, i_10_265_4024_0, i_10_265_4117_0, i_10_265_4170_0,
    i_10_265_4189_0, i_10_265_4277_0, i_10_265_4290_0, i_10_265_4326_0,
    i_10_265_4354_0, i_10_265_4371_0, i_10_265_4449_0, i_10_265_4476_0,
    i_10_265_4477_0, i_10_265_4539_0, i_10_265_4575_0, i_10_265_4593_0,
    o_10_265_0_0  );
  input  i_10_265_210_0, i_10_265_277_0, i_10_265_279_0, i_10_265_280_0,
    i_10_265_287_0, i_10_265_444_0, i_10_265_447_0, i_10_265_499_0,
    i_10_265_517_0, i_10_265_586_0, i_10_265_587_0, i_10_265_607_0,
    i_10_265_792_0, i_10_265_793_0, i_10_265_796_0, i_10_265_798_0,
    i_10_265_799_0, i_10_265_904_0, i_10_265_1049_0, i_10_265_1123_0,
    i_10_265_1164_0, i_10_265_1171_0, i_10_265_1200_0, i_10_265_1201_0,
    i_10_265_1234_0, i_10_265_1305_0, i_10_265_1362_0, i_10_265_1444_0,
    i_10_265_1447_0, i_10_265_1448_0, i_10_265_1602_0, i_10_265_1651_0,
    i_10_265_1652_0, i_10_265_1732_0, i_10_265_1818_0, i_10_265_1822_0,
    i_10_265_1881_0, i_10_265_1882_0, i_10_265_2155_0, i_10_265_2329_0,
    i_10_265_2338_0, i_10_265_2362_0, i_10_265_2382_0, i_10_265_2448_0,
    i_10_265_2449_0, i_10_265_2451_0, i_10_265_2475_0, i_10_265_2543_0,
    i_10_265_2659_0, i_10_265_2660_0, i_10_265_2662_0, i_10_265_2663_0,
    i_10_265_2728_0, i_10_265_2731_0, i_10_265_2814_0, i_10_265_2888_0,
    i_10_265_2916_0, i_10_265_2917_0, i_10_265_2919_0, i_10_265_2922_0,
    i_10_265_2979_0, i_10_265_3039_0, i_10_265_3047_0, i_10_265_3049_0,
    i_10_265_3050_0, i_10_265_3092_0, i_10_265_3109_0, i_10_265_3169_0,
    i_10_265_3172_0, i_10_265_3282_0, i_10_265_3294_0, i_10_265_3388_0,
    i_10_265_3496_0, i_10_265_3615_0, i_10_265_3684_0, i_10_265_3720_0,
    i_10_265_3721_0, i_10_265_3729_0, i_10_265_3787_0, i_10_265_3851_0,
    i_10_265_3854_0, i_10_265_3859_0, i_10_265_3892_0, i_10_265_3919_0,
    i_10_265_3950_0, i_10_265_4024_0, i_10_265_4117_0, i_10_265_4170_0,
    i_10_265_4189_0, i_10_265_4277_0, i_10_265_4290_0, i_10_265_4326_0,
    i_10_265_4354_0, i_10_265_4371_0, i_10_265_4449_0, i_10_265_4476_0,
    i_10_265_4477_0, i_10_265_4539_0, i_10_265_4575_0, i_10_265_4593_0;
  output o_10_265_0_0;
  assign o_10_265_0_0 = 0;
endmodule



// Benchmark "kernel_10_266" written by ABC on Sun Jul 19 10:25:36 2020

module kernel_10_266 ( 
    i_10_266_33_0, i_10_266_39_0, i_10_266_69_0, i_10_266_144_0,
    i_10_266_146_0, i_10_266_178_0, i_10_266_248_0, i_10_266_257_0,
    i_10_266_271_0, i_10_266_282_0, i_10_266_406_0, i_10_266_429_0,
    i_10_266_445_0, i_10_266_502_0, i_10_266_520_0, i_10_266_561_0,
    i_10_266_585_0, i_10_266_598_0, i_10_266_642_0, i_10_266_730_0,
    i_10_266_731_0, i_10_266_733_0, i_10_266_734_0, i_10_266_737_0,
    i_10_266_832_0, i_10_266_847_0, i_10_266_848_0, i_10_266_1003_0,
    i_10_266_1039_0, i_10_266_1233_0, i_10_266_1234_0, i_10_266_1239_0,
    i_10_266_1268_0, i_10_266_1307_0, i_10_266_1347_0, i_10_266_1353_0,
    i_10_266_1365_0, i_10_266_1441_0, i_10_266_1442_0, i_10_266_1611_0,
    i_10_266_1650_0, i_10_266_1697_0, i_10_266_1717_0, i_10_266_1824_0,
    i_10_266_1825_0, i_10_266_1872_0, i_10_266_1942_0, i_10_266_2079_0,
    i_10_266_2179_0, i_10_266_2206_0, i_10_266_2376_0, i_10_266_2379_0,
    i_10_266_2434_0, i_10_266_2452_0, i_10_266_2457_0, i_10_266_2463_0,
    i_10_266_2471_0, i_10_266_2504_0, i_10_266_2602_0, i_10_266_2617_0,
    i_10_266_2632_0, i_10_266_2658_0, i_10_266_2724_0, i_10_266_2730_0,
    i_10_266_2789_0, i_10_266_2829_0, i_10_266_2869_0, i_10_266_2920_0,
    i_10_266_2922_0, i_10_266_3038_0, i_10_266_3076_0, i_10_266_3097_0,
    i_10_266_3098_0, i_10_266_3101_0, i_10_266_3198_0, i_10_266_3201_0,
    i_10_266_3203_0, i_10_266_3282_0, i_10_266_3351_0, i_10_266_3469_0,
    i_10_266_3472_0, i_10_266_3473_0, i_10_266_3496_0, i_10_266_3525_0,
    i_10_266_3612_0, i_10_266_3650_0, i_10_266_3685_0, i_10_266_3717_0,
    i_10_266_3783_0, i_10_266_3786_0, i_10_266_3787_0, i_10_266_3788_0,
    i_10_266_3810_0, i_10_266_3834_0, i_10_266_3835_0, i_10_266_3857_0,
    i_10_266_4054_0, i_10_266_4101_0, i_10_266_4279_0, i_10_266_4563_0,
    o_10_266_0_0  );
  input  i_10_266_33_0, i_10_266_39_0, i_10_266_69_0, i_10_266_144_0,
    i_10_266_146_0, i_10_266_178_0, i_10_266_248_0, i_10_266_257_0,
    i_10_266_271_0, i_10_266_282_0, i_10_266_406_0, i_10_266_429_0,
    i_10_266_445_0, i_10_266_502_0, i_10_266_520_0, i_10_266_561_0,
    i_10_266_585_0, i_10_266_598_0, i_10_266_642_0, i_10_266_730_0,
    i_10_266_731_0, i_10_266_733_0, i_10_266_734_0, i_10_266_737_0,
    i_10_266_832_0, i_10_266_847_0, i_10_266_848_0, i_10_266_1003_0,
    i_10_266_1039_0, i_10_266_1233_0, i_10_266_1234_0, i_10_266_1239_0,
    i_10_266_1268_0, i_10_266_1307_0, i_10_266_1347_0, i_10_266_1353_0,
    i_10_266_1365_0, i_10_266_1441_0, i_10_266_1442_0, i_10_266_1611_0,
    i_10_266_1650_0, i_10_266_1697_0, i_10_266_1717_0, i_10_266_1824_0,
    i_10_266_1825_0, i_10_266_1872_0, i_10_266_1942_0, i_10_266_2079_0,
    i_10_266_2179_0, i_10_266_2206_0, i_10_266_2376_0, i_10_266_2379_0,
    i_10_266_2434_0, i_10_266_2452_0, i_10_266_2457_0, i_10_266_2463_0,
    i_10_266_2471_0, i_10_266_2504_0, i_10_266_2602_0, i_10_266_2617_0,
    i_10_266_2632_0, i_10_266_2658_0, i_10_266_2724_0, i_10_266_2730_0,
    i_10_266_2789_0, i_10_266_2829_0, i_10_266_2869_0, i_10_266_2920_0,
    i_10_266_2922_0, i_10_266_3038_0, i_10_266_3076_0, i_10_266_3097_0,
    i_10_266_3098_0, i_10_266_3101_0, i_10_266_3198_0, i_10_266_3201_0,
    i_10_266_3203_0, i_10_266_3282_0, i_10_266_3351_0, i_10_266_3469_0,
    i_10_266_3472_0, i_10_266_3473_0, i_10_266_3496_0, i_10_266_3525_0,
    i_10_266_3612_0, i_10_266_3650_0, i_10_266_3685_0, i_10_266_3717_0,
    i_10_266_3783_0, i_10_266_3786_0, i_10_266_3787_0, i_10_266_3788_0,
    i_10_266_3810_0, i_10_266_3834_0, i_10_266_3835_0, i_10_266_3857_0,
    i_10_266_4054_0, i_10_266_4101_0, i_10_266_4279_0, i_10_266_4563_0;
  output o_10_266_0_0;
  assign o_10_266_0_0 = 0;
endmodule



// Benchmark "kernel_10_267" written by ABC on Sun Jul 19 10:25:37 2020

module kernel_10_267 ( 
    i_10_267_34_0, i_10_267_85_0, i_10_267_86_0, i_10_267_89_0,
    i_10_267_121_0, i_10_267_151_0, i_10_267_172_0, i_10_267_249_0,
    i_10_267_283_0, i_10_267_330_0, i_10_267_427_0, i_10_267_431_0,
    i_10_267_438_0, i_10_267_445_0, i_10_267_465_0, i_10_267_520_0,
    i_10_267_565_0, i_10_267_898_0, i_10_267_996_0, i_10_267_1003_0,
    i_10_267_1032_0, i_10_267_1033_0, i_10_267_1165_0, i_10_267_1166_0,
    i_10_267_1168_0, i_10_267_1173_0, i_10_267_1174_0, i_10_267_1233_0,
    i_10_267_1237_0, i_10_267_1239_0, i_10_267_1293_0, i_10_267_1365_0,
    i_10_267_1381_0, i_10_267_1488_0, i_10_267_1491_0, i_10_267_1536_0,
    i_10_267_1537_0, i_10_267_1583_0, i_10_267_1691_0, i_10_267_1821_0,
    i_10_267_1824_0, i_10_267_1997_0, i_10_267_2004_0, i_10_267_2352_0,
    i_10_267_2382_0, i_10_267_2391_0, i_10_267_2392_0, i_10_267_2463_0,
    i_10_267_2508_0, i_10_267_2542_0, i_10_267_2607_0, i_10_267_2634_0,
    i_10_267_2635_0, i_10_267_2653_0, i_10_267_2654_0, i_10_267_2660_0,
    i_10_267_2680_0, i_10_267_2703_0, i_10_267_2705_0, i_10_267_2724_0,
    i_10_267_2725_0, i_10_267_2729_0, i_10_267_2730_0, i_10_267_2731_0,
    i_10_267_2733_0, i_10_267_2734_0, i_10_267_2787_0, i_10_267_2828_0,
    i_10_267_2834_0, i_10_267_2920_0, i_10_267_2986_0, i_10_267_3120_0,
    i_10_267_3150_0, i_10_267_3151_0, i_10_267_3152_0, i_10_267_3162_0,
    i_10_267_3163_0, i_10_267_3165_0, i_10_267_3195_0, i_10_267_3202_0,
    i_10_267_3300_0, i_10_267_3496_0, i_10_267_3522_0, i_10_267_3616_0,
    i_10_267_3617_0, i_10_267_3688_0, i_10_267_3689_0, i_10_267_3733_0,
    i_10_267_3839_0, i_10_267_3846_0, i_10_267_3847_0, i_10_267_3856_0,
    i_10_267_4116_0, i_10_267_4117_0, i_10_267_4120_0, i_10_267_4128_0,
    i_10_267_4288_0, i_10_267_4290_0, i_10_267_4566_0, i_10_267_4567_0,
    o_10_267_0_0  );
  input  i_10_267_34_0, i_10_267_85_0, i_10_267_86_0, i_10_267_89_0,
    i_10_267_121_0, i_10_267_151_0, i_10_267_172_0, i_10_267_249_0,
    i_10_267_283_0, i_10_267_330_0, i_10_267_427_0, i_10_267_431_0,
    i_10_267_438_0, i_10_267_445_0, i_10_267_465_0, i_10_267_520_0,
    i_10_267_565_0, i_10_267_898_0, i_10_267_996_0, i_10_267_1003_0,
    i_10_267_1032_0, i_10_267_1033_0, i_10_267_1165_0, i_10_267_1166_0,
    i_10_267_1168_0, i_10_267_1173_0, i_10_267_1174_0, i_10_267_1233_0,
    i_10_267_1237_0, i_10_267_1239_0, i_10_267_1293_0, i_10_267_1365_0,
    i_10_267_1381_0, i_10_267_1488_0, i_10_267_1491_0, i_10_267_1536_0,
    i_10_267_1537_0, i_10_267_1583_0, i_10_267_1691_0, i_10_267_1821_0,
    i_10_267_1824_0, i_10_267_1997_0, i_10_267_2004_0, i_10_267_2352_0,
    i_10_267_2382_0, i_10_267_2391_0, i_10_267_2392_0, i_10_267_2463_0,
    i_10_267_2508_0, i_10_267_2542_0, i_10_267_2607_0, i_10_267_2634_0,
    i_10_267_2635_0, i_10_267_2653_0, i_10_267_2654_0, i_10_267_2660_0,
    i_10_267_2680_0, i_10_267_2703_0, i_10_267_2705_0, i_10_267_2724_0,
    i_10_267_2725_0, i_10_267_2729_0, i_10_267_2730_0, i_10_267_2731_0,
    i_10_267_2733_0, i_10_267_2734_0, i_10_267_2787_0, i_10_267_2828_0,
    i_10_267_2834_0, i_10_267_2920_0, i_10_267_2986_0, i_10_267_3120_0,
    i_10_267_3150_0, i_10_267_3151_0, i_10_267_3152_0, i_10_267_3162_0,
    i_10_267_3163_0, i_10_267_3165_0, i_10_267_3195_0, i_10_267_3202_0,
    i_10_267_3300_0, i_10_267_3496_0, i_10_267_3522_0, i_10_267_3616_0,
    i_10_267_3617_0, i_10_267_3688_0, i_10_267_3689_0, i_10_267_3733_0,
    i_10_267_3839_0, i_10_267_3846_0, i_10_267_3847_0, i_10_267_3856_0,
    i_10_267_4116_0, i_10_267_4117_0, i_10_267_4120_0, i_10_267_4128_0,
    i_10_267_4288_0, i_10_267_4290_0, i_10_267_4566_0, i_10_267_4567_0;
  output o_10_267_0_0;
  assign o_10_267_0_0 = ~((~i_10_267_89_0 & ((~i_10_267_431_0 & ~i_10_267_1365_0 & ~i_10_267_2463_0 & ~i_10_267_2634_0 & ~i_10_267_3162_0) | (~i_10_267_898_0 & ~i_10_267_1165_0 & i_10_267_1824_0 & ~i_10_267_3846_0 & ~i_10_267_3847_0 & ~i_10_267_4128_0))) | (~i_10_267_3162_0 & ((~i_10_267_445_0 & ((~i_10_267_1168_0 & ~i_10_267_1821_0 & ~i_10_267_2382_0 & ~i_10_267_2734_0) | (~i_10_267_465_0 & i_10_267_2635_0 & ~i_10_267_2730_0 & ~i_10_267_3733_0 & ~i_10_267_4567_0))) | (~i_10_267_172_0 & ~i_10_267_520_0 & ~i_10_267_1032_0 & ~i_10_267_1033_0 & ~i_10_267_1165_0 & ~i_10_267_1166_0 & ~i_10_267_3847_0))) | (~i_10_267_3165_0 & ((~i_10_267_85_0 & ~i_10_267_172_0 & ~i_10_267_1168_0 & ((~i_10_267_151_0 & ~i_10_267_1233_0 & ~i_10_267_1365_0 & ~i_10_267_2725_0 & ~i_10_267_4116_0) | (~i_10_267_996_0 & ~i_10_267_1491_0 & ~i_10_267_2729_0 & ~i_10_267_3163_0 & ~i_10_267_3195_0 & ~i_10_267_3202_0 & ~i_10_267_4567_0))) | (~i_10_267_898_0 & ~i_10_267_1033_0 & ~i_10_267_1166_0 & ~i_10_267_2607_0 & i_10_267_2660_0 & ~i_10_267_4128_0) | (~i_10_267_1237_0 & ~i_10_267_2382_0 & ~i_10_267_2733_0 & ~i_10_267_3846_0 & ~i_10_267_4290_0))) | (~i_10_267_1165_0 & ((i_10_267_2352_0 & ~i_10_267_2680_0 & ~i_10_267_2986_0) | (~i_10_267_996_0 & i_10_267_1239_0 & ~i_10_267_4288_0 & ~i_10_267_4566_0))) | (~i_10_267_1166_0 & ((~i_10_267_2635_0 & ~i_10_267_2920_0 & ~i_10_267_4120_0) | (~i_10_267_85_0 & ~i_10_267_1233_0 & ~i_10_267_1239_0 & ~i_10_267_2725_0 & ~i_10_267_2734_0 & i_10_267_4566_0))) | (~i_10_267_2680_0 & ((~i_10_267_1233_0 & i_10_267_2635_0 & ~i_10_267_2828_0 & ~i_10_267_2986_0 & i_10_267_3522_0 & ~i_10_267_3847_0) | (~i_10_267_427_0 & ~i_10_267_1491_0 & ~i_10_267_2352_0 & ~i_10_267_2463_0 & i_10_267_2731_0 & i_10_267_4116_0 & ~i_10_267_4128_0))) | (~i_10_267_2730_0 & ((i_10_267_172_0 & ~i_10_267_1033_0 & i_10_267_2834_0) | (i_10_267_445_0 & ~i_10_267_1239_0 & ~i_10_267_3847_0 & ~i_10_267_3856_0 & ~i_10_267_4120_0))) | (~i_10_267_4290_0 & ((~i_10_267_1488_0 & ~i_10_267_2634_0) | (i_10_267_2920_0 & i_10_267_3856_0) | (~i_10_267_2607_0 & ~i_10_267_2660_0 & i_10_267_3616_0 & ~i_10_267_3846_0 & ~i_10_267_4128_0))) | (~i_10_267_249_0 & i_10_267_465_0 & ~i_10_267_2731_0 & ~i_10_267_3163_0 & ~i_10_267_3847_0 & ~i_10_267_4566_0 & ~i_10_267_4567_0));
endmodule



// Benchmark "kernel_10_268" written by ABC on Sun Jul 19 10:25:38 2020

module kernel_10_268 ( 
    i_10_268_34_0, i_10_268_42_0, i_10_268_51_0, i_10_268_52_0,
    i_10_268_53_0, i_10_268_142_0, i_10_268_151_0, i_10_268_177_0,
    i_10_268_184_0, i_10_268_287_0, i_10_268_294_0, i_10_268_321_0,
    i_10_268_430_0, i_10_268_431_0, i_10_268_445_0, i_10_268_447_0,
    i_10_268_464_0, i_10_268_465_0, i_10_268_637_0, i_10_268_699_0,
    i_10_268_834_0, i_10_268_897_0, i_10_268_934_0, i_10_268_957_0,
    i_10_268_961_0, i_10_268_966_0, i_10_268_971_0, i_10_268_1087_0,
    i_10_268_1236_0, i_10_268_1239_0, i_10_268_1241_0, i_10_268_1311_0,
    i_10_268_1543_0, i_10_268_1582_0, i_10_268_1583_0, i_10_268_1636_0,
    i_10_268_1645_0, i_10_268_1687_0, i_10_268_1688_0, i_10_268_1696_0,
    i_10_268_1725_0, i_10_268_1816_0, i_10_268_1823_0, i_10_268_1957_0,
    i_10_268_2040_0, i_10_268_2391_0, i_10_268_2471_0, i_10_268_2472_0,
    i_10_268_2535_0, i_10_268_2545_0, i_10_268_2632_0, i_10_268_2633_0,
    i_10_268_2679_0, i_10_268_2706_0, i_10_268_2707_0, i_10_268_2708_0,
    i_10_268_2716_0, i_10_268_2717_0, i_10_268_2730_0, i_10_268_2830_0,
    i_10_268_2913_0, i_10_268_3198_0, i_10_268_3238_0, i_10_268_3390_0,
    i_10_268_3468_0, i_10_268_3469_0, i_10_268_3495_0, i_10_268_3496_0,
    i_10_268_3497_0, i_10_268_3498_0, i_10_268_3500_0, i_10_268_3509_0,
    i_10_268_3541_0, i_10_268_3588_0, i_10_268_3648_0, i_10_268_3651_0,
    i_10_268_3783_0, i_10_268_3784_0, i_10_268_3785_0, i_10_268_3787_0,
    i_10_268_3846_0, i_10_268_3849_0, i_10_268_3851_0, i_10_268_3859_0,
    i_10_268_3886_0, i_10_268_3949_0, i_10_268_3999_0, i_10_268_4119_0,
    i_10_268_4121_0, i_10_268_4165_0, i_10_268_4242_0, i_10_268_4269_0,
    i_10_268_4270_0, i_10_268_4287_0, i_10_268_4462_0, i_10_268_4463_0,
    i_10_268_4566_0, i_10_268_4567_0, i_10_268_4570_0, i_10_268_4588_0,
    o_10_268_0_0  );
  input  i_10_268_34_0, i_10_268_42_0, i_10_268_51_0, i_10_268_52_0,
    i_10_268_53_0, i_10_268_142_0, i_10_268_151_0, i_10_268_177_0,
    i_10_268_184_0, i_10_268_287_0, i_10_268_294_0, i_10_268_321_0,
    i_10_268_430_0, i_10_268_431_0, i_10_268_445_0, i_10_268_447_0,
    i_10_268_464_0, i_10_268_465_0, i_10_268_637_0, i_10_268_699_0,
    i_10_268_834_0, i_10_268_897_0, i_10_268_934_0, i_10_268_957_0,
    i_10_268_961_0, i_10_268_966_0, i_10_268_971_0, i_10_268_1087_0,
    i_10_268_1236_0, i_10_268_1239_0, i_10_268_1241_0, i_10_268_1311_0,
    i_10_268_1543_0, i_10_268_1582_0, i_10_268_1583_0, i_10_268_1636_0,
    i_10_268_1645_0, i_10_268_1687_0, i_10_268_1688_0, i_10_268_1696_0,
    i_10_268_1725_0, i_10_268_1816_0, i_10_268_1823_0, i_10_268_1957_0,
    i_10_268_2040_0, i_10_268_2391_0, i_10_268_2471_0, i_10_268_2472_0,
    i_10_268_2535_0, i_10_268_2545_0, i_10_268_2632_0, i_10_268_2633_0,
    i_10_268_2679_0, i_10_268_2706_0, i_10_268_2707_0, i_10_268_2708_0,
    i_10_268_2716_0, i_10_268_2717_0, i_10_268_2730_0, i_10_268_2830_0,
    i_10_268_2913_0, i_10_268_3198_0, i_10_268_3238_0, i_10_268_3390_0,
    i_10_268_3468_0, i_10_268_3469_0, i_10_268_3495_0, i_10_268_3496_0,
    i_10_268_3497_0, i_10_268_3498_0, i_10_268_3500_0, i_10_268_3509_0,
    i_10_268_3541_0, i_10_268_3588_0, i_10_268_3648_0, i_10_268_3651_0,
    i_10_268_3783_0, i_10_268_3784_0, i_10_268_3785_0, i_10_268_3787_0,
    i_10_268_3846_0, i_10_268_3849_0, i_10_268_3851_0, i_10_268_3859_0,
    i_10_268_3886_0, i_10_268_3949_0, i_10_268_3999_0, i_10_268_4119_0,
    i_10_268_4121_0, i_10_268_4165_0, i_10_268_4242_0, i_10_268_4269_0,
    i_10_268_4270_0, i_10_268_4287_0, i_10_268_4462_0, i_10_268_4463_0,
    i_10_268_4566_0, i_10_268_4567_0, i_10_268_4570_0, i_10_268_4588_0;
  output o_10_268_0_0;
  assign o_10_268_0_0 = 0;
endmodule



// Benchmark "kernel_10_269" written by ABC on Sun Jul 19 10:25:39 2020

module kernel_10_269 ( 
    i_10_269_25_0, i_10_269_187_0, i_10_269_249_0, i_10_269_258_0,
    i_10_269_259_0, i_10_269_260_0, i_10_269_276_0, i_10_269_277_0,
    i_10_269_282_0, i_10_269_283_0, i_10_269_321_0, i_10_269_426_0,
    i_10_269_517_0, i_10_269_600_0, i_10_269_717_0, i_10_269_728_0,
    i_10_269_754_0, i_10_269_800_0, i_10_269_850_0, i_10_269_853_0,
    i_10_269_997_0, i_10_269_998_0, i_10_269_1033_0, i_10_269_1034_0,
    i_10_269_1124_0, i_10_269_1194_0, i_10_269_1195_0, i_10_269_1239_0,
    i_10_269_1240_0, i_10_269_1249_0, i_10_269_1250_0, i_10_269_1356_0,
    i_10_269_1515_0, i_10_269_1579_0, i_10_269_1583_0, i_10_269_1618_0,
    i_10_269_1619_0, i_10_269_1653_0, i_10_269_1654_0, i_10_269_1687_0,
    i_10_269_1688_0, i_10_269_1819_0, i_10_269_1820_0, i_10_269_1821_0,
    i_10_269_1823_0, i_10_269_1826_0, i_10_269_1833_0, i_10_269_1960_0,
    i_10_269_2352_0, i_10_269_2355_0, i_10_269_2356_0, i_10_269_2357_0,
    i_10_269_2436_0, i_10_269_2457_0, i_10_269_2458_0, i_10_269_2460_0,
    i_10_269_2509_0, i_10_269_2563_0, i_10_269_2634_0, i_10_269_2716_0,
    i_10_269_2823_0, i_10_269_2868_0, i_10_269_2887_0, i_10_269_2895_0,
    i_10_269_3192_0, i_10_269_3195_0, i_10_269_3273_0, i_10_269_3319_0,
    i_10_269_3391_0, i_10_269_3401_0, i_10_269_3434_0, i_10_269_3508_0,
    i_10_269_3562_0, i_10_269_3610_0, i_10_269_3651_0, i_10_269_3687_0,
    i_10_269_3775_0, i_10_269_3783_0, i_10_269_3787_0, i_10_269_3813_0,
    i_10_269_3814_0, i_10_269_3815_0, i_10_269_3846_0, i_10_269_3910_0,
    i_10_269_3946_0, i_10_269_3947_0, i_10_269_3948_0, i_10_269_4012_0,
    i_10_269_4013_0, i_10_269_4055_0, i_10_269_4117_0, i_10_269_4118_0,
    i_10_269_4171_0, i_10_269_4279_0, i_10_269_4280_0, i_10_269_4290_0,
    i_10_269_4291_0, i_10_269_4369_0, i_10_269_4461_0, i_10_269_4462_0,
    o_10_269_0_0  );
  input  i_10_269_25_0, i_10_269_187_0, i_10_269_249_0, i_10_269_258_0,
    i_10_269_259_0, i_10_269_260_0, i_10_269_276_0, i_10_269_277_0,
    i_10_269_282_0, i_10_269_283_0, i_10_269_321_0, i_10_269_426_0,
    i_10_269_517_0, i_10_269_600_0, i_10_269_717_0, i_10_269_728_0,
    i_10_269_754_0, i_10_269_800_0, i_10_269_850_0, i_10_269_853_0,
    i_10_269_997_0, i_10_269_998_0, i_10_269_1033_0, i_10_269_1034_0,
    i_10_269_1124_0, i_10_269_1194_0, i_10_269_1195_0, i_10_269_1239_0,
    i_10_269_1240_0, i_10_269_1249_0, i_10_269_1250_0, i_10_269_1356_0,
    i_10_269_1515_0, i_10_269_1579_0, i_10_269_1583_0, i_10_269_1618_0,
    i_10_269_1619_0, i_10_269_1653_0, i_10_269_1654_0, i_10_269_1687_0,
    i_10_269_1688_0, i_10_269_1819_0, i_10_269_1820_0, i_10_269_1821_0,
    i_10_269_1823_0, i_10_269_1826_0, i_10_269_1833_0, i_10_269_1960_0,
    i_10_269_2352_0, i_10_269_2355_0, i_10_269_2356_0, i_10_269_2357_0,
    i_10_269_2436_0, i_10_269_2457_0, i_10_269_2458_0, i_10_269_2460_0,
    i_10_269_2509_0, i_10_269_2563_0, i_10_269_2634_0, i_10_269_2716_0,
    i_10_269_2823_0, i_10_269_2868_0, i_10_269_2887_0, i_10_269_2895_0,
    i_10_269_3192_0, i_10_269_3195_0, i_10_269_3273_0, i_10_269_3319_0,
    i_10_269_3391_0, i_10_269_3401_0, i_10_269_3434_0, i_10_269_3508_0,
    i_10_269_3562_0, i_10_269_3610_0, i_10_269_3651_0, i_10_269_3687_0,
    i_10_269_3775_0, i_10_269_3783_0, i_10_269_3787_0, i_10_269_3813_0,
    i_10_269_3814_0, i_10_269_3815_0, i_10_269_3846_0, i_10_269_3910_0,
    i_10_269_3946_0, i_10_269_3947_0, i_10_269_3948_0, i_10_269_4012_0,
    i_10_269_4013_0, i_10_269_4055_0, i_10_269_4117_0, i_10_269_4118_0,
    i_10_269_4171_0, i_10_269_4279_0, i_10_269_4280_0, i_10_269_4290_0,
    i_10_269_4291_0, i_10_269_4369_0, i_10_269_4461_0, i_10_269_4462_0;
  output o_10_269_0_0;
  assign o_10_269_0_0 = 0;
endmodule



// Benchmark "kernel_10_270" written by ABC on Sun Jul 19 10:25:40 2020

module kernel_10_270 ( 
    i_10_270_29_0, i_10_270_145_0, i_10_270_146_0, i_10_270_176_0,
    i_10_270_221_0, i_10_270_247_0, i_10_270_254_0, i_10_270_281_0,
    i_10_270_318_0, i_10_270_319_0, i_10_270_391_0, i_10_270_434_0,
    i_10_270_461_0, i_10_270_462_0, i_10_270_463_0, i_10_270_464_0,
    i_10_270_513_0, i_10_270_711_0, i_10_270_713_0, i_10_270_749_0,
    i_10_270_800_0, i_10_270_954_0, i_10_270_992_0, i_10_270_1027_0,
    i_10_270_1046_0, i_10_270_1049_0, i_10_270_1083_0, i_10_270_1220_0,
    i_10_270_1349_0, i_10_270_1361_0, i_10_270_1396_0, i_10_270_1397_0,
    i_10_270_1451_0, i_10_270_1539_0, i_10_270_1616_0, i_10_270_1622_0,
    i_10_270_1685_0, i_10_270_1821_0, i_10_270_1822_0, i_10_270_1954_0,
    i_10_270_1981_0, i_10_270_2066_0, i_10_270_2201_0, i_10_270_2349_0,
    i_10_270_2351_0, i_10_270_2353_0, i_10_270_2453_0, i_10_270_2471_0,
    i_10_270_2601_0, i_10_270_2612_0, i_10_270_2660_0, i_10_270_2701_0,
    i_10_270_2702_0, i_10_270_2704_0, i_10_270_2711_0, i_10_270_2722_0,
    i_10_270_2723_0, i_10_270_2783_0, i_10_270_2920_0, i_10_270_3038_0,
    i_10_270_3044_0, i_10_270_3196_0, i_10_270_3198_0, i_10_270_3199_0,
    i_10_270_3232_0, i_10_270_3278_0, i_10_270_3314_0, i_10_270_3388_0,
    i_10_270_3407_0, i_10_270_3503_0, i_10_270_3519_0, i_10_270_3520_0,
    i_10_270_3584_0, i_10_270_3586_0, i_10_270_3620_0, i_10_270_3645_0,
    i_10_270_3646_0, i_10_270_3683_0, i_10_270_3728_0, i_10_270_3783_0,
    i_10_270_3785_0, i_10_270_3837_0, i_10_270_3838_0, i_10_270_3839_0,
    i_10_270_3852_0, i_10_270_3859_0, i_10_270_3980_0, i_10_270_4115_0,
    i_10_270_4117_0, i_10_270_4126_0, i_10_270_4153_0, i_10_270_4171_0,
    i_10_270_4172_0, i_10_270_4275_0, i_10_270_4279_0, i_10_270_4280_0,
    i_10_270_4288_0, i_10_270_4289_0, i_10_270_4566_0, i_10_270_4568_0,
    o_10_270_0_0  );
  input  i_10_270_29_0, i_10_270_145_0, i_10_270_146_0, i_10_270_176_0,
    i_10_270_221_0, i_10_270_247_0, i_10_270_254_0, i_10_270_281_0,
    i_10_270_318_0, i_10_270_319_0, i_10_270_391_0, i_10_270_434_0,
    i_10_270_461_0, i_10_270_462_0, i_10_270_463_0, i_10_270_464_0,
    i_10_270_513_0, i_10_270_711_0, i_10_270_713_0, i_10_270_749_0,
    i_10_270_800_0, i_10_270_954_0, i_10_270_992_0, i_10_270_1027_0,
    i_10_270_1046_0, i_10_270_1049_0, i_10_270_1083_0, i_10_270_1220_0,
    i_10_270_1349_0, i_10_270_1361_0, i_10_270_1396_0, i_10_270_1397_0,
    i_10_270_1451_0, i_10_270_1539_0, i_10_270_1616_0, i_10_270_1622_0,
    i_10_270_1685_0, i_10_270_1821_0, i_10_270_1822_0, i_10_270_1954_0,
    i_10_270_1981_0, i_10_270_2066_0, i_10_270_2201_0, i_10_270_2349_0,
    i_10_270_2351_0, i_10_270_2353_0, i_10_270_2453_0, i_10_270_2471_0,
    i_10_270_2601_0, i_10_270_2612_0, i_10_270_2660_0, i_10_270_2701_0,
    i_10_270_2702_0, i_10_270_2704_0, i_10_270_2711_0, i_10_270_2722_0,
    i_10_270_2723_0, i_10_270_2783_0, i_10_270_2920_0, i_10_270_3038_0,
    i_10_270_3044_0, i_10_270_3196_0, i_10_270_3198_0, i_10_270_3199_0,
    i_10_270_3232_0, i_10_270_3278_0, i_10_270_3314_0, i_10_270_3388_0,
    i_10_270_3407_0, i_10_270_3503_0, i_10_270_3519_0, i_10_270_3520_0,
    i_10_270_3584_0, i_10_270_3586_0, i_10_270_3620_0, i_10_270_3645_0,
    i_10_270_3646_0, i_10_270_3683_0, i_10_270_3728_0, i_10_270_3783_0,
    i_10_270_3785_0, i_10_270_3837_0, i_10_270_3838_0, i_10_270_3839_0,
    i_10_270_3852_0, i_10_270_3859_0, i_10_270_3980_0, i_10_270_4115_0,
    i_10_270_4117_0, i_10_270_4126_0, i_10_270_4153_0, i_10_270_4171_0,
    i_10_270_4172_0, i_10_270_4275_0, i_10_270_4279_0, i_10_270_4280_0,
    i_10_270_4288_0, i_10_270_4289_0, i_10_270_4566_0, i_10_270_4568_0;
  output o_10_270_0_0;
  assign o_10_270_0_0 = 0;
endmodule



// Benchmark "kernel_10_271" written by ABC on Sun Jul 19 10:25:41 2020

module kernel_10_271 ( 
    i_10_271_161_0, i_10_271_175_0, i_10_271_183_0, i_10_271_187_0,
    i_10_271_220_0, i_10_271_246_0, i_10_271_248_0, i_10_271_251_0,
    i_10_271_268_0, i_10_271_279_0, i_10_271_285_0, i_10_271_410_0,
    i_10_271_431_0, i_10_271_446_0, i_10_271_462_0, i_10_271_463_0,
    i_10_271_464_0, i_10_271_465_0, i_10_271_466_0, i_10_271_467_0,
    i_10_271_754_0, i_10_271_755_0, i_10_271_799_0, i_10_271_995_0,
    i_10_271_997_0, i_10_271_1237_0, i_10_271_1238_0, i_10_271_1239_0,
    i_10_271_1240_0, i_10_271_1241_0, i_10_271_1312_0, i_10_271_1362_0,
    i_10_271_1363_0, i_10_271_1434_0, i_10_271_1436_0, i_10_271_1438_0,
    i_10_271_1439_0, i_10_271_1545_0, i_10_271_1654_0, i_10_271_1655_0,
    i_10_271_1685_0, i_10_271_1821_0, i_10_271_1825_0, i_10_271_1911_0,
    i_10_271_1912_0, i_10_271_2338_0, i_10_271_2339_0, i_10_271_2349_0,
    i_10_271_2350_0, i_10_271_2351_0, i_10_271_2356_0, i_10_271_2357_0,
    i_10_271_2361_0, i_10_271_2364_0, i_10_271_2383_0, i_10_271_2384_0,
    i_10_271_2455_0, i_10_271_2463_0, i_10_271_2464_0, i_10_271_2470_0,
    i_10_271_2609_0, i_10_271_2635_0, i_10_271_2636_0, i_10_271_2658_0,
    i_10_271_2662_0, i_10_271_2713_0, i_10_271_2732_0, i_10_271_2735_0,
    i_10_271_2916_0, i_10_271_2921_0, i_10_271_2985_0, i_10_271_2986_0,
    i_10_271_2987_0, i_10_271_3070_0, i_10_271_3151_0, i_10_271_3163_0,
    i_10_271_3195_0, i_10_271_3237_0, i_10_271_3238_0, i_10_271_3271_0,
    i_10_271_3275_0, i_10_271_3278_0, i_10_271_3390_0, i_10_271_3686_0,
    i_10_271_3837_0, i_10_271_3839_0, i_10_271_3840_0, i_10_271_3841_0,
    i_10_271_3852_0, i_10_271_3860_0, i_10_271_3892_0, i_10_271_4116_0,
    i_10_271_4117_0, i_10_271_4118_0, i_10_271_4121_0, i_10_271_4130_0,
    i_10_271_4269_0, i_10_271_4270_0, i_10_271_4288_0, i_10_271_4289_0,
    o_10_271_0_0  );
  input  i_10_271_161_0, i_10_271_175_0, i_10_271_183_0, i_10_271_187_0,
    i_10_271_220_0, i_10_271_246_0, i_10_271_248_0, i_10_271_251_0,
    i_10_271_268_0, i_10_271_279_0, i_10_271_285_0, i_10_271_410_0,
    i_10_271_431_0, i_10_271_446_0, i_10_271_462_0, i_10_271_463_0,
    i_10_271_464_0, i_10_271_465_0, i_10_271_466_0, i_10_271_467_0,
    i_10_271_754_0, i_10_271_755_0, i_10_271_799_0, i_10_271_995_0,
    i_10_271_997_0, i_10_271_1237_0, i_10_271_1238_0, i_10_271_1239_0,
    i_10_271_1240_0, i_10_271_1241_0, i_10_271_1312_0, i_10_271_1362_0,
    i_10_271_1363_0, i_10_271_1434_0, i_10_271_1436_0, i_10_271_1438_0,
    i_10_271_1439_0, i_10_271_1545_0, i_10_271_1654_0, i_10_271_1655_0,
    i_10_271_1685_0, i_10_271_1821_0, i_10_271_1825_0, i_10_271_1911_0,
    i_10_271_1912_0, i_10_271_2338_0, i_10_271_2339_0, i_10_271_2349_0,
    i_10_271_2350_0, i_10_271_2351_0, i_10_271_2356_0, i_10_271_2357_0,
    i_10_271_2361_0, i_10_271_2364_0, i_10_271_2383_0, i_10_271_2384_0,
    i_10_271_2455_0, i_10_271_2463_0, i_10_271_2464_0, i_10_271_2470_0,
    i_10_271_2609_0, i_10_271_2635_0, i_10_271_2636_0, i_10_271_2658_0,
    i_10_271_2662_0, i_10_271_2713_0, i_10_271_2732_0, i_10_271_2735_0,
    i_10_271_2916_0, i_10_271_2921_0, i_10_271_2985_0, i_10_271_2986_0,
    i_10_271_2987_0, i_10_271_3070_0, i_10_271_3151_0, i_10_271_3163_0,
    i_10_271_3195_0, i_10_271_3237_0, i_10_271_3238_0, i_10_271_3271_0,
    i_10_271_3275_0, i_10_271_3278_0, i_10_271_3390_0, i_10_271_3686_0,
    i_10_271_3837_0, i_10_271_3839_0, i_10_271_3840_0, i_10_271_3841_0,
    i_10_271_3852_0, i_10_271_3860_0, i_10_271_3892_0, i_10_271_4116_0,
    i_10_271_4117_0, i_10_271_4118_0, i_10_271_4121_0, i_10_271_4130_0,
    i_10_271_4269_0, i_10_271_4270_0, i_10_271_4288_0, i_10_271_4289_0;
  output o_10_271_0_0;
  assign o_10_271_0_0 = ~((~i_10_271_246_0 & ((i_10_271_462_0 & ~i_10_271_2383_0 & ~i_10_271_2985_0 & ~i_10_271_3839_0 & ~i_10_271_4118_0) | (~i_10_271_220_0 & ~i_10_271_248_0 & i_10_271_1821_0 & ~i_10_271_2916_0 & i_10_271_3070_0 & ~i_10_271_4269_0))) | (i_10_271_279_0 & ((~i_10_271_220_0 & ~i_10_271_410_0 & ~i_10_271_1545_0 & ~i_10_271_2338_0 & ~i_10_271_2361_0 & ~i_10_271_2732_0 & ~i_10_271_2916_0 & ~i_10_271_3237_0 & ~i_10_271_4121_0) | (~i_10_271_755_0 & ~i_10_271_1821_0 & ~i_10_271_2364_0 & ~i_10_271_2986_0 & ~i_10_271_3839_0 & ~i_10_271_3860_0 & ~i_10_271_4270_0))) | (~i_10_271_2635_0 & ((~i_10_271_220_0 & ((~i_10_271_995_0 & ~i_10_271_2339_0 & ~i_10_271_2916_0 & ~i_10_271_2921_0 & ~i_10_271_4116_0 & ~i_10_271_4118_0) | (i_10_271_464_0 & ~i_10_271_4288_0))) | (~i_10_271_446_0 & ((~i_10_271_2349_0 & ~i_10_271_2361_0 & ~i_10_271_2636_0 & ~i_10_271_4116_0 & ~i_10_271_4118_0 & ~i_10_271_4121_0 & ~i_10_271_4269_0) | (~i_10_271_2658_0 & i_10_271_2916_0 & i_10_271_4117_0 & i_10_271_4289_0))) | i_10_271_3237_0 | (~i_10_271_279_0 & ~i_10_271_754_0 & ~i_10_271_2361_0 & ~i_10_271_2609_0 & ~i_10_271_2636_0 & ~i_10_271_2916_0 & ~i_10_271_3070_0 & ~i_10_271_4270_0))) | (~i_10_271_248_0 & ((~i_10_271_431_0 & ((~i_10_271_755_0 & ~i_10_271_2364_0 & ~i_10_271_2986_0 & ~i_10_271_3163_0 & i_10_271_3841_0) | (i_10_271_466_0 & ~i_10_271_2356_0 & ~i_10_271_2921_0 & ~i_10_271_2987_0 & i_10_271_4288_0))) | (~i_10_271_754_0 & ~i_10_271_3163_0 & ((~i_10_271_997_0 & ~i_10_271_1821_0 & ~i_10_271_3275_0 & i_10_271_3892_0 & ~i_10_271_4121_0) | (~i_10_271_251_0 & i_10_271_466_0 & i_10_271_467_0 & ~i_10_271_2364_0 & ~i_10_271_2987_0 & ~i_10_271_3237_0 & ~i_10_271_4116_0 & ~i_10_271_4130_0))) | (~i_10_271_279_0 & ~i_10_271_1654_0 & ~i_10_271_2361_0 & ~i_10_271_2383_0 & ~i_10_271_2455_0 & ~i_10_271_2609_0 & ~i_10_271_2916_0 & ~i_10_271_3271_0 & ~i_10_271_4117_0) | (~i_10_271_410_0 & ~i_10_271_755_0 & ~i_10_271_995_0 & ~i_10_271_1545_0 & i_10_271_1654_0 & ~i_10_271_2463_0 & ~i_10_271_2985_0 & ~i_10_271_3275_0 & ~i_10_271_3390_0 & ~i_10_271_4270_0))) | (i_10_271_462_0 & (i_10_271_1237_0 | (~i_10_271_175_0 & i_10_271_799_0 & ~i_10_271_2356_0 & ~i_10_271_2361_0 & ~i_10_271_2986_0))) | (i_10_271_464_0 & ~i_10_271_1655_0 & (i_10_271_3892_0 | (~i_10_271_251_0 & ~i_10_271_2351_0 & ~i_10_271_2356_0 & ~i_10_271_2364_0 & ~i_10_271_2455_0 & ~i_10_271_2609_0 & ~i_10_271_3070_0 & ~i_10_271_3275_0 & ~i_10_271_3840_0 & ~i_10_271_4116_0))) | (~i_10_271_464_0 & i_10_271_466_0 & ((~i_10_271_1821_0 & ~i_10_271_2986_0 & ~i_10_271_3271_0 & ~i_10_271_4118_0) | (~i_10_271_251_0 & ~i_10_271_463_0 & ~i_10_271_1241_0 & ~i_10_271_2357_0 & ~i_10_271_2463_0 & ~i_10_271_3837_0 & ~i_10_271_3841_0 & ~i_10_271_3852_0 & i_10_271_4117_0 & ~i_10_271_4288_0))) | (~i_10_271_3390_0 & ((~i_10_271_251_0 & ((~i_10_271_997_0 & i_10_271_1240_0 & ~i_10_271_2609_0 & ~i_10_271_3238_0) | (~i_10_271_1237_0 & ~i_10_271_1434_0 & i_10_271_1825_0 & ~i_10_271_2349_0 & ~i_10_271_2356_0 & ~i_10_271_2383_0 & ~i_10_271_2662_0 & ~i_10_271_2916_0 & ~i_10_271_3275_0))) | (~i_10_271_1654_0 & ~i_10_271_4116_0 & ~i_10_271_4118_0 & ~i_10_271_4121_0 & ~i_10_271_4130_0 & i_10_271_4288_0))) | (~i_10_271_754_0 & ((~i_10_271_410_0 & ~i_10_271_2636_0 & ((~i_10_271_1438_0 & i_10_271_2350_0 & ~i_10_271_2609_0 & ~i_10_271_2916_0 & ~i_10_271_3837_0) | (~i_10_271_995_0 & ~i_10_271_1436_0 & i_10_271_1825_0 & ~i_10_271_2735_0 & ~i_10_271_3275_0 & ~i_10_271_3852_0 & ~i_10_271_4289_0))) | (~i_10_271_1821_0 & i_10_271_1825_0 & ~i_10_271_2349_0 & ~i_10_271_2384_0 & i_10_271_3195_0) | (~i_10_271_183_0 & i_10_271_463_0 & ~i_10_271_799_0 & ~i_10_271_2364_0 & ~i_10_271_2735_0 & ~i_10_271_2921_0 & ~i_10_271_3070_0 & ~i_10_271_3238_0 & ~i_10_271_3839_0))) | (i_10_271_463_0 & ((~i_10_271_997_0 & i_10_271_1238_0 & ~i_10_271_4269_0) | (~i_10_271_2350_0 & ~i_10_271_2384_0 & i_10_271_2455_0 & ~i_10_271_2463_0 & ~i_10_271_2916_0 & ~i_10_271_3686_0 & ~i_10_271_4270_0))) | (~i_10_271_1654_0 & ((~i_10_271_995_0 & ((i_10_271_3686_0 & ~i_10_271_3839_0 & ~i_10_271_4116_0) | (~i_10_271_446_0 & ~i_10_271_1237_0 & ~i_10_271_2364_0 & ~i_10_271_2383_0 & ~i_10_271_2609_0 & ~i_10_271_3070_0 & ~i_10_271_3163_0 & ~i_10_271_3195_0 & ~i_10_271_4117_0))) | (i_10_271_3271_0 & i_10_271_3841_0))) | (~i_10_271_1821_0 & ((~i_10_271_755_0 & ~i_10_271_2384_0 & ~i_10_271_2609_0 & ~i_10_271_3070_0 & ~i_10_271_3271_0 & i_10_271_3841_0 & ~i_10_271_4269_0) | (i_10_271_1237_0 & ~i_10_271_1545_0 & ~i_10_271_2357_0 & ~i_10_271_4270_0))) | (~i_10_271_2916_0 & ((~i_10_271_1363_0 & i_10_271_2351_0 & i_10_271_2713_0 & ~i_10_271_2921_0) | (i_10_271_2658_0 & ~i_10_271_2662_0 & ~i_10_271_4118_0))) | (i_10_271_1239_0 & i_10_271_1240_0 & i_10_271_2455_0 & ~i_10_271_2713_0) | (i_10_271_1685_0 & ~i_10_271_2349_0 & ~i_10_271_2350_0 & ~i_10_271_2658_0 & i_10_271_3070_0 & i_10_271_3852_0 & ~i_10_271_4117_0) | (i_10_271_1821_0 & ~i_10_271_3195_0 & i_10_271_4117_0 & ~i_10_271_4269_0 & ~i_10_271_4270_0 & i_10_271_4288_0) | (i_10_271_175_0 & ~i_10_271_410_0 & i_10_271_2350_0 & i_10_271_4289_0));
endmodule



// Benchmark "kernel_10_272" written by ABC on Sun Jul 19 10:25:42 2020

module kernel_10_272 ( 
    i_10_272_22_0, i_10_272_135_0, i_10_272_144_0, i_10_272_193_0,
    i_10_272_218_0, i_10_272_274_0, i_10_272_284_0, i_10_272_289_0,
    i_10_272_371_0, i_10_272_460_0, i_10_272_461_0, i_10_272_694_0,
    i_10_272_792_0, i_10_272_846_0, i_10_272_900_0, i_10_272_901_0,
    i_10_272_949_0, i_10_272_1280_0, i_10_272_1315_0, i_10_272_1360_0,
    i_10_272_1369_0, i_10_272_1370_0, i_10_272_1391_0, i_10_272_1441_0,
    i_10_272_1442_0, i_10_272_1479_0, i_10_272_1566_0, i_10_272_1567_0,
    i_10_272_1568_0, i_10_272_1651_0, i_10_272_1714_0, i_10_272_1818_0,
    i_10_272_1911_0, i_10_272_1924_0, i_10_272_1927_0, i_10_272_1930_0,
    i_10_272_1979_0, i_10_272_1984_0, i_10_272_2080_0, i_10_272_2089_0,
    i_10_272_2125_0, i_10_272_2151_0, i_10_272_2155_0, i_10_272_2269_0,
    i_10_272_2305_0, i_10_272_2306_0, i_10_272_2324_0, i_10_272_2350_0,
    i_10_272_2460_0, i_10_272_2475_0, i_10_272_2502_0, i_10_272_2503_0,
    i_10_272_2504_0, i_10_272_2506_0, i_10_272_2550_0, i_10_272_2629_0,
    i_10_272_2630_0, i_10_272_2677_0, i_10_272_2692_0, i_10_272_2729_0,
    i_10_272_2767_0, i_10_272_2803_0, i_10_272_2804_0, i_10_272_2953_0,
    i_10_272_2957_0, i_10_272_2959_0, i_10_272_3025_0, i_10_272_3026_0,
    i_10_272_3029_0, i_10_272_3096_0, i_10_272_3097_0, i_10_272_3214_0,
    i_10_272_3258_0, i_10_272_3298_0, i_10_272_3321_0, i_10_272_3357_0,
    i_10_272_3358_0, i_10_272_3540_0, i_10_272_3602_0, i_10_272_3651_0,
    i_10_272_3802_0, i_10_272_3838_0, i_10_272_3848_0, i_10_272_3979_0,
    i_10_272_3980_0, i_10_272_3994_0, i_10_272_4068_0, i_10_272_4089_0,
    i_10_272_4090_0, i_10_272_4114_0, i_10_272_4230_0, i_10_272_4266_0,
    i_10_272_4270_0, i_10_272_4279_0, i_10_272_4280_0, i_10_272_4357_0,
    i_10_272_4358_0, i_10_272_4403_0, i_10_272_4433_0, i_10_272_4440_0,
    o_10_272_0_0  );
  input  i_10_272_22_0, i_10_272_135_0, i_10_272_144_0, i_10_272_193_0,
    i_10_272_218_0, i_10_272_274_0, i_10_272_284_0, i_10_272_289_0,
    i_10_272_371_0, i_10_272_460_0, i_10_272_461_0, i_10_272_694_0,
    i_10_272_792_0, i_10_272_846_0, i_10_272_900_0, i_10_272_901_0,
    i_10_272_949_0, i_10_272_1280_0, i_10_272_1315_0, i_10_272_1360_0,
    i_10_272_1369_0, i_10_272_1370_0, i_10_272_1391_0, i_10_272_1441_0,
    i_10_272_1442_0, i_10_272_1479_0, i_10_272_1566_0, i_10_272_1567_0,
    i_10_272_1568_0, i_10_272_1651_0, i_10_272_1714_0, i_10_272_1818_0,
    i_10_272_1911_0, i_10_272_1924_0, i_10_272_1927_0, i_10_272_1930_0,
    i_10_272_1979_0, i_10_272_1984_0, i_10_272_2080_0, i_10_272_2089_0,
    i_10_272_2125_0, i_10_272_2151_0, i_10_272_2155_0, i_10_272_2269_0,
    i_10_272_2305_0, i_10_272_2306_0, i_10_272_2324_0, i_10_272_2350_0,
    i_10_272_2460_0, i_10_272_2475_0, i_10_272_2502_0, i_10_272_2503_0,
    i_10_272_2504_0, i_10_272_2506_0, i_10_272_2550_0, i_10_272_2629_0,
    i_10_272_2630_0, i_10_272_2677_0, i_10_272_2692_0, i_10_272_2729_0,
    i_10_272_2767_0, i_10_272_2803_0, i_10_272_2804_0, i_10_272_2953_0,
    i_10_272_2957_0, i_10_272_2959_0, i_10_272_3025_0, i_10_272_3026_0,
    i_10_272_3029_0, i_10_272_3096_0, i_10_272_3097_0, i_10_272_3214_0,
    i_10_272_3258_0, i_10_272_3298_0, i_10_272_3321_0, i_10_272_3357_0,
    i_10_272_3358_0, i_10_272_3540_0, i_10_272_3602_0, i_10_272_3651_0,
    i_10_272_3802_0, i_10_272_3838_0, i_10_272_3848_0, i_10_272_3979_0,
    i_10_272_3980_0, i_10_272_3994_0, i_10_272_4068_0, i_10_272_4089_0,
    i_10_272_4090_0, i_10_272_4114_0, i_10_272_4230_0, i_10_272_4266_0,
    i_10_272_4270_0, i_10_272_4279_0, i_10_272_4280_0, i_10_272_4357_0,
    i_10_272_4358_0, i_10_272_4403_0, i_10_272_4433_0, i_10_272_4440_0;
  output o_10_272_0_0;
  assign o_10_272_0_0 = 0;
endmodule



// Benchmark "kernel_10_273" written by ABC on Sun Jul 19 10:25:43 2020

module kernel_10_273 ( 
    i_10_273_281_0, i_10_273_282_0, i_10_273_283_0, i_10_273_296_0,
    i_10_273_327_0, i_10_273_328_0, i_10_273_408_0, i_10_273_411_0,
    i_10_273_413_0, i_10_273_425_0, i_10_273_443_0, i_10_273_712_0,
    i_10_273_748_0, i_10_273_800_0, i_10_273_1134_0, i_10_273_1235_0,
    i_10_273_1240_0, i_10_273_1248_0, i_10_273_1263_0, i_10_273_1264_0,
    i_10_273_1309_0, i_10_273_1366_0, i_10_273_1445_0, i_10_273_1580_0,
    i_10_273_1649_0, i_10_273_1819_0, i_10_273_1821_0, i_10_273_1823_0,
    i_10_273_1824_0, i_10_273_1876_0, i_10_273_1910_0, i_10_273_1911_0,
    i_10_273_1912_0, i_10_273_1913_0, i_10_273_1948_0, i_10_273_1989_0,
    i_10_273_2180_0, i_10_273_2186_0, i_10_273_2353_0, i_10_273_2354_0,
    i_10_273_2362_0, i_10_273_2380_0, i_10_273_2453_0, i_10_273_2468_0,
    i_10_273_2632_0, i_10_273_2634_0, i_10_273_2635_0, i_10_273_2636_0,
    i_10_273_2659_0, i_10_273_2660_0, i_10_273_2677_0, i_10_273_2711_0,
    i_10_273_2718_0, i_10_273_2719_0, i_10_273_2721_0, i_10_273_2722_0,
    i_10_273_2731_0, i_10_273_2781_0, i_10_273_2916_0, i_10_273_2921_0,
    i_10_273_2979_0, i_10_273_2980_0, i_10_273_2981_0, i_10_273_3033_0,
    i_10_273_3034_0, i_10_273_3035_0, i_10_273_3039_0, i_10_273_3040_0,
    i_10_273_3069_0, i_10_273_3196_0, i_10_273_3281_0, i_10_273_3283_0,
    i_10_273_3284_0, i_10_273_3324_0, i_10_273_3384_0, i_10_273_3388_0,
    i_10_273_3389_0, i_10_273_3392_0, i_10_273_3406_0, i_10_273_3437_0,
    i_10_273_3519_0, i_10_273_3520_0, i_10_273_3523_0, i_10_273_3613_0,
    i_10_273_3649_0, i_10_273_3650_0, i_10_273_3835_0, i_10_273_3849_0,
    i_10_273_3850_0, i_10_273_3855_0, i_10_273_3856_0, i_10_273_3857_0,
    i_10_273_3859_0, i_10_273_3906_0, i_10_273_3991_0, i_10_273_4114_0,
    i_10_273_4121_0, i_10_273_4563_0, i_10_273_4566_0, i_10_273_4568_0,
    o_10_273_0_0  );
  input  i_10_273_281_0, i_10_273_282_0, i_10_273_283_0, i_10_273_296_0,
    i_10_273_327_0, i_10_273_328_0, i_10_273_408_0, i_10_273_411_0,
    i_10_273_413_0, i_10_273_425_0, i_10_273_443_0, i_10_273_712_0,
    i_10_273_748_0, i_10_273_800_0, i_10_273_1134_0, i_10_273_1235_0,
    i_10_273_1240_0, i_10_273_1248_0, i_10_273_1263_0, i_10_273_1264_0,
    i_10_273_1309_0, i_10_273_1366_0, i_10_273_1445_0, i_10_273_1580_0,
    i_10_273_1649_0, i_10_273_1819_0, i_10_273_1821_0, i_10_273_1823_0,
    i_10_273_1824_0, i_10_273_1876_0, i_10_273_1910_0, i_10_273_1911_0,
    i_10_273_1912_0, i_10_273_1913_0, i_10_273_1948_0, i_10_273_1989_0,
    i_10_273_2180_0, i_10_273_2186_0, i_10_273_2353_0, i_10_273_2354_0,
    i_10_273_2362_0, i_10_273_2380_0, i_10_273_2453_0, i_10_273_2468_0,
    i_10_273_2632_0, i_10_273_2634_0, i_10_273_2635_0, i_10_273_2636_0,
    i_10_273_2659_0, i_10_273_2660_0, i_10_273_2677_0, i_10_273_2711_0,
    i_10_273_2718_0, i_10_273_2719_0, i_10_273_2721_0, i_10_273_2722_0,
    i_10_273_2731_0, i_10_273_2781_0, i_10_273_2916_0, i_10_273_2921_0,
    i_10_273_2979_0, i_10_273_2980_0, i_10_273_2981_0, i_10_273_3033_0,
    i_10_273_3034_0, i_10_273_3035_0, i_10_273_3039_0, i_10_273_3040_0,
    i_10_273_3069_0, i_10_273_3196_0, i_10_273_3281_0, i_10_273_3283_0,
    i_10_273_3284_0, i_10_273_3324_0, i_10_273_3384_0, i_10_273_3388_0,
    i_10_273_3389_0, i_10_273_3392_0, i_10_273_3406_0, i_10_273_3437_0,
    i_10_273_3519_0, i_10_273_3520_0, i_10_273_3523_0, i_10_273_3613_0,
    i_10_273_3649_0, i_10_273_3650_0, i_10_273_3835_0, i_10_273_3849_0,
    i_10_273_3850_0, i_10_273_3855_0, i_10_273_3856_0, i_10_273_3857_0,
    i_10_273_3859_0, i_10_273_3906_0, i_10_273_3991_0, i_10_273_4114_0,
    i_10_273_4121_0, i_10_273_4563_0, i_10_273_4566_0, i_10_273_4568_0;
  output o_10_273_0_0;
  assign o_10_273_0_0 = ~((~i_10_273_296_0 & ~i_10_273_2980_0 & ((~i_10_273_1911_0 & ~i_10_273_2635_0 & ~i_10_273_2711_0 & ~i_10_273_3649_0) | (~i_10_273_1248_0 & ~i_10_273_1263_0 & ~i_10_273_2636_0 & ~i_10_273_3281_0 & ~i_10_273_3906_0 & ~i_10_273_4114_0))) | (~i_10_273_413_0 & ((~i_10_273_327_0 & ~i_10_273_1912_0 & ~i_10_273_2981_0) | (~i_10_273_408_0 & ~i_10_273_748_0 & ~i_10_273_1445_0 & ~i_10_273_1649_0 & ~i_10_273_1876_0 & ~i_10_273_2731_0 & ~i_10_273_2921_0 & ~i_10_273_3284_0 & ~i_10_273_3519_0))) | (~i_10_273_3437_0 & ((~i_10_273_327_0 & ((~i_10_273_408_0 & ~i_10_273_1264_0 & i_10_273_2722_0 & ~i_10_273_3519_0 & ~i_10_273_3857_0) | (~i_10_273_1912_0 & ~i_10_273_2719_0 & ~i_10_273_3039_0 & i_10_273_4114_0))) | (~i_10_273_1263_0 & i_10_273_2634_0 & ~i_10_273_3856_0) | (~i_10_273_408_0 & ~i_10_273_411_0 & ~i_10_273_1876_0 & ~i_10_273_2711_0 & ~i_10_273_2718_0 & ~i_10_273_3283_0 & ~i_10_273_3392_0 & ~i_10_273_3520_0 & ~i_10_273_3906_0))) | (~i_10_273_1264_0 & ((~i_10_273_327_0 & ~i_10_273_748_0 & ~i_10_273_2659_0 & ~i_10_273_3040_0 & ~i_10_273_3855_0) | (~i_10_273_1821_0 & ~i_10_273_1912_0 & ~i_10_273_2718_0 & ~i_10_273_3039_0 & ~i_10_273_3281_0 & ~i_10_273_3650_0 & ~i_10_273_4566_0))) | (~i_10_273_748_0 & (i_10_273_3850_0 | (~i_10_273_800_0 & ~i_10_273_1240_0 & ~i_10_273_1876_0 & i_10_273_2731_0 & i_10_273_3859_0))) | (~i_10_273_2659_0 & ((i_10_273_3283_0 & i_10_273_3859_0) | (~i_10_273_1913_0 & ~i_10_273_2353_0 & ~i_10_273_2634_0 & ~i_10_273_3859_0 & ~i_10_273_4114_0))) | (~i_10_273_2722_0 & ((i_10_273_2635_0 & i_10_273_2721_0 & i_10_273_2731_0) | (~i_10_273_1445_0 & ~i_10_273_3519_0 & ~i_10_273_3855_0 & ~i_10_273_3857_0))) | (i_10_273_1819_0 & i_10_273_2453_0 & ~i_10_273_3033_0 & ~i_10_273_3406_0) | (~i_10_273_1309_0 & ~i_10_273_1821_0 & ~i_10_273_2354_0 & ~i_10_273_2468_0 & ~i_10_273_3649_0 & ~i_10_273_3855_0) | (~i_10_273_281_0 & ~i_10_273_283_0 & ~i_10_273_3281_0 & i_10_273_3835_0) | (~i_10_273_712_0 & ~i_10_273_1263_0 & i_10_273_3406_0 & ~i_10_273_3857_0 & ~i_10_273_3859_0));
endmodule



// Benchmark "kernel_10_274" written by ABC on Sun Jul 19 10:25:44 2020

module kernel_10_274 ( 
    i_10_274_27_0, i_10_274_28_0, i_10_274_29_0, i_10_274_117_0,
    i_10_274_118_0, i_10_274_119_0, i_10_274_122_0, i_10_274_153_0,
    i_10_274_174_0, i_10_274_279_0, i_10_274_280_0, i_10_274_286_0,
    i_10_274_316_0, i_10_274_462_0, i_10_274_464_0, i_10_274_514_0,
    i_10_274_559_0, i_10_274_793_0, i_10_274_958_0, i_10_274_1235_0,
    i_10_274_1240_0, i_10_274_1242_0, i_10_274_1309_0, i_10_274_1310_0,
    i_10_274_1549_0, i_10_274_1652_0, i_10_274_1686_0, i_10_274_1687_0,
    i_10_274_1820_0, i_10_274_1822_0, i_10_274_2018_0, i_10_274_2026_0,
    i_10_274_2029_0, i_10_274_2179_0, i_10_274_2180_0, i_10_274_2200_0,
    i_10_274_2350_0, i_10_274_2352_0, i_10_274_2380_0, i_10_274_2449_0,
    i_10_274_2452_0, i_10_274_2453_0, i_10_274_2466_0, i_10_274_2467_0,
    i_10_274_2470_0, i_10_274_2471_0, i_10_274_2502_0, i_10_274_2610_0,
    i_10_274_2628_0, i_10_274_2631_0, i_10_274_2659_0, i_10_274_2663_0,
    i_10_274_2700_0, i_10_274_2701_0, i_10_274_2719_0, i_10_274_2782_0,
    i_10_274_2827_0, i_10_274_2919_0, i_10_274_3036_0, i_10_274_3037_0,
    i_10_274_3088_0, i_10_274_3089_0, i_10_274_3155_0, i_10_274_3200_0,
    i_10_274_3385_0, i_10_274_3390_0, i_10_274_3519_0, i_10_274_3520_0,
    i_10_274_3525_0, i_10_274_3583_0, i_10_274_3586_0, i_10_274_3587_0,
    i_10_274_3613_0, i_10_274_3646_0, i_10_274_3649_0, i_10_274_3785_0,
    i_10_274_3837_0, i_10_274_3842_0, i_10_274_3847_0, i_10_274_3851_0,
    i_10_274_3854_0, i_10_274_3855_0, i_10_274_3856_0, i_10_274_3857_0,
    i_10_274_3860_0, i_10_274_3907_0, i_10_274_3978_0, i_10_274_4051_0,
    i_10_274_4052_0, i_10_274_4113_0, i_10_274_4114_0, i_10_274_4120_0,
    i_10_274_4168_0, i_10_274_4276_0, i_10_274_4288_0, i_10_274_4289_0,
    i_10_274_4564_0, i_10_274_4565_0, i_10_274_4568_0, i_10_274_4570_0,
    o_10_274_0_0  );
  input  i_10_274_27_0, i_10_274_28_0, i_10_274_29_0, i_10_274_117_0,
    i_10_274_118_0, i_10_274_119_0, i_10_274_122_0, i_10_274_153_0,
    i_10_274_174_0, i_10_274_279_0, i_10_274_280_0, i_10_274_286_0,
    i_10_274_316_0, i_10_274_462_0, i_10_274_464_0, i_10_274_514_0,
    i_10_274_559_0, i_10_274_793_0, i_10_274_958_0, i_10_274_1235_0,
    i_10_274_1240_0, i_10_274_1242_0, i_10_274_1309_0, i_10_274_1310_0,
    i_10_274_1549_0, i_10_274_1652_0, i_10_274_1686_0, i_10_274_1687_0,
    i_10_274_1820_0, i_10_274_1822_0, i_10_274_2018_0, i_10_274_2026_0,
    i_10_274_2029_0, i_10_274_2179_0, i_10_274_2180_0, i_10_274_2200_0,
    i_10_274_2350_0, i_10_274_2352_0, i_10_274_2380_0, i_10_274_2449_0,
    i_10_274_2452_0, i_10_274_2453_0, i_10_274_2466_0, i_10_274_2467_0,
    i_10_274_2470_0, i_10_274_2471_0, i_10_274_2502_0, i_10_274_2610_0,
    i_10_274_2628_0, i_10_274_2631_0, i_10_274_2659_0, i_10_274_2663_0,
    i_10_274_2700_0, i_10_274_2701_0, i_10_274_2719_0, i_10_274_2782_0,
    i_10_274_2827_0, i_10_274_2919_0, i_10_274_3036_0, i_10_274_3037_0,
    i_10_274_3088_0, i_10_274_3089_0, i_10_274_3155_0, i_10_274_3200_0,
    i_10_274_3385_0, i_10_274_3390_0, i_10_274_3519_0, i_10_274_3520_0,
    i_10_274_3525_0, i_10_274_3583_0, i_10_274_3586_0, i_10_274_3587_0,
    i_10_274_3613_0, i_10_274_3646_0, i_10_274_3649_0, i_10_274_3785_0,
    i_10_274_3837_0, i_10_274_3842_0, i_10_274_3847_0, i_10_274_3851_0,
    i_10_274_3854_0, i_10_274_3855_0, i_10_274_3856_0, i_10_274_3857_0,
    i_10_274_3860_0, i_10_274_3907_0, i_10_274_3978_0, i_10_274_4051_0,
    i_10_274_4052_0, i_10_274_4113_0, i_10_274_4114_0, i_10_274_4120_0,
    i_10_274_4168_0, i_10_274_4276_0, i_10_274_4288_0, i_10_274_4289_0,
    i_10_274_4564_0, i_10_274_4565_0, i_10_274_4568_0, i_10_274_4570_0;
  output o_10_274_0_0;
  assign o_10_274_0_0 = ~((~i_10_274_28_0 & ((~i_10_274_29_0 & ((~i_10_274_27_0 & ~i_10_274_122_0 & ~i_10_274_174_0 & i_10_274_464_0 & ~i_10_274_1240_0 & ~i_10_274_3037_0 & i_10_274_3649_0 & ~i_10_274_3842_0 & ~i_10_274_3860_0) | (~i_10_274_286_0 & i_10_274_1652_0 & ~i_10_274_2179_0 & i_10_274_3856_0 & ~i_10_274_4570_0))) | (~i_10_274_117_0 & ~i_10_274_464_0 & ~i_10_274_2663_0 & ~i_10_274_3586_0 & i_10_274_4114_0))) | (~i_10_274_286_0 & ~i_10_274_3200_0 & ((i_10_274_2200_0 & ~i_10_274_2453_0 & ~i_10_274_2470_0 & ~i_10_274_2610_0 & ~i_10_274_3036_0 & ~i_10_274_3390_0 & ~i_10_274_3854_0) | (~i_10_274_27_0 & ~i_10_274_174_0 & ~i_10_274_3089_0 & ~i_10_274_3586_0 & ~i_10_274_3842_0 & ~i_10_274_3860_0 & ~i_10_274_4120_0))) | (~i_10_274_27_0 & ((i_10_274_2467_0 & ~i_10_274_2827_0 & ~i_10_274_3583_0) | (i_10_274_2200_0 & ~i_10_274_3842_0 & i_10_274_4113_0))) | (~i_10_274_1310_0 & (~i_10_274_3856_0 | (i_10_274_3847_0 & i_10_274_3857_0))) | (~i_10_274_2919_0 & ((i_10_274_1686_0 & ((~i_10_274_122_0 & ~i_10_274_3036_0 & ~i_10_274_3856_0) | (~i_10_274_174_0 & i_10_274_2452_0 & ~i_10_274_2663_0 & i_10_274_3385_0 & ~i_10_274_4120_0))) | (~i_10_274_2663_0 & ~i_10_274_3037_0 & i_10_274_3837_0 & ~i_10_274_3856_0 & ~i_10_274_3860_0))) | (~i_10_274_174_0 & ((i_10_274_3390_0 & ~i_10_274_3586_0 & ~i_10_274_3587_0) | (~i_10_274_464_0 & ~i_10_274_3613_0 & ~i_10_274_3856_0 & i_10_274_3857_0))) | (~i_10_274_1822_0 & ((i_10_274_464_0 & ~i_10_274_958_0 & ~i_10_274_2663_0 & ~i_10_274_3855_0) | (~i_10_274_3036_0 & ~i_10_274_3857_0 & ~i_10_274_3860_0))) | (i_10_274_2352_0 & ((~i_10_274_464_0 & ~i_10_274_2467_0 & ~i_10_274_2471_0 & ~i_10_274_2663_0 & ~i_10_274_3842_0 & ~i_10_274_3851_0) | (~i_10_274_2470_0 & i_10_274_3525_0 & ~i_10_274_3860_0))) | (~i_10_274_464_0 & ((i_10_274_2663_0 & ~i_10_274_3037_0 & ~i_10_274_3587_0 & ~i_10_274_3649_0 & ~i_10_274_3837_0) | (~i_10_274_2352_0 & ~i_10_274_2452_0 & ~i_10_274_2659_0 & i_10_274_3860_0 & ~i_10_274_4051_0))) | (~i_10_274_2471_0 & ((~i_10_274_3037_0 & ~i_10_274_3649_0 & ~i_10_274_3842_0 & ~i_10_274_3857_0 & ~i_10_274_3860_0) | (~i_10_274_2452_0 & ~i_10_274_2659_0 & ~i_10_274_3613_0 & i_10_274_3842_0 & ~i_10_274_3855_0 & ~i_10_274_4113_0))) | (~i_10_274_2452_0 & ~i_10_274_3649_0 & ((~i_10_274_2663_0 & i_10_274_3390_0) | (~i_10_274_1240_0 & ~i_10_274_3857_0 & ~i_10_274_3860_0))) | (~i_10_274_1309_0 & ~i_10_274_2502_0) | (i_10_274_1652_0 & i_10_274_2701_0) | (i_10_274_514_0 & ~i_10_274_2827_0 & ~i_10_274_3037_0) | (i_10_274_2200_0 & ~i_10_274_3613_0 & i_10_274_3851_0 & ~i_10_274_3855_0) | (~i_10_274_2470_0 & i_10_274_2631_0 & ~i_10_274_3586_0 & ~i_10_274_3856_0) | (i_10_274_2466_0 & ~i_10_274_3583_0 & i_10_274_3837_0 & i_10_274_3978_0) | (i_10_274_2719_0 & ~i_10_274_4052_0) | (~i_10_274_2179_0 & i_10_274_2449_0 & ~i_10_274_4114_0) | (~i_10_274_1235_0 & ~i_10_274_3036_0 & ~i_10_274_3842_0 & i_10_274_3847_0 & ~i_10_274_4568_0));
endmodule



// Benchmark "kernel_10_275" written by ABC on Sun Jul 19 10:25:46 2020

module kernel_10_275 ( 
    i_10_275_69_0, i_10_275_176_0, i_10_275_178_0, i_10_275_283_0,
    i_10_275_284_0, i_10_275_328_0, i_10_275_329_0, i_10_275_406_0,
    i_10_275_409_0, i_10_275_410_0, i_10_275_412_0, i_10_275_458_0,
    i_10_275_462_0, i_10_275_463_0, i_10_275_464_0, i_10_275_466_0,
    i_10_275_467_0, i_10_275_511_0, i_10_275_799_0, i_10_275_800_0,
    i_10_275_959_0, i_10_275_962_0, i_10_275_1002_0, i_10_275_1233_0,
    i_10_275_1307_0, i_10_275_1312_0, i_10_275_1547_0, i_10_275_1552_0,
    i_10_275_1553_0, i_10_275_1555_0, i_10_275_1556_0, i_10_275_1626_0,
    i_10_275_1652_0, i_10_275_1691_0, i_10_275_1716_0, i_10_275_1717_0,
    i_10_275_1726_0, i_10_275_1821_0, i_10_275_1822_0, i_10_275_1825_0,
    i_10_275_1949_0, i_10_275_2005_0, i_10_275_2159_0, i_10_275_2199_0,
    i_10_275_2311_0, i_10_275_2312_0, i_10_275_2352_0, i_10_275_2353_0,
    i_10_275_2354_0, i_10_275_2355_0, i_10_275_2407_0, i_10_275_2473_0,
    i_10_275_2631_0, i_10_275_2632_0, i_10_275_2635_0, i_10_275_2656_0,
    i_10_275_2661_0, i_10_275_2663_0, i_10_275_2725_0, i_10_275_2730_0,
    i_10_275_2731_0, i_10_275_2827_0, i_10_275_2832_0, i_10_275_2834_0,
    i_10_275_2880_0, i_10_275_2881_0, i_10_275_2921_0, i_10_275_2923_0,
    i_10_275_2924_0, i_10_275_3075_0, i_10_275_3076_0, i_10_275_3094_0,
    i_10_275_3155_0, i_10_275_3385_0, i_10_275_3388_0, i_10_275_3389_0,
    i_10_275_3391_0, i_10_275_3392_0, i_10_275_3497_0, i_10_275_3541_0,
    i_10_275_3545_0, i_10_275_3551_0, i_10_275_3614_0, i_10_275_3783_0,
    i_10_275_3788_0, i_10_275_3835_0, i_10_275_3854_0, i_10_275_3856_0,
    i_10_275_3859_0, i_10_275_3860_0, i_10_275_3894_0, i_10_275_3982_0,
    i_10_275_3994_0, i_10_275_4050_0, i_10_275_4124_0, i_10_275_4220_0,
    i_10_275_4237_0, i_10_275_4270_0, i_10_275_4273_0, i_10_275_4564_0,
    o_10_275_0_0  );
  input  i_10_275_69_0, i_10_275_176_0, i_10_275_178_0, i_10_275_283_0,
    i_10_275_284_0, i_10_275_328_0, i_10_275_329_0, i_10_275_406_0,
    i_10_275_409_0, i_10_275_410_0, i_10_275_412_0, i_10_275_458_0,
    i_10_275_462_0, i_10_275_463_0, i_10_275_464_0, i_10_275_466_0,
    i_10_275_467_0, i_10_275_511_0, i_10_275_799_0, i_10_275_800_0,
    i_10_275_959_0, i_10_275_962_0, i_10_275_1002_0, i_10_275_1233_0,
    i_10_275_1307_0, i_10_275_1312_0, i_10_275_1547_0, i_10_275_1552_0,
    i_10_275_1553_0, i_10_275_1555_0, i_10_275_1556_0, i_10_275_1626_0,
    i_10_275_1652_0, i_10_275_1691_0, i_10_275_1716_0, i_10_275_1717_0,
    i_10_275_1726_0, i_10_275_1821_0, i_10_275_1822_0, i_10_275_1825_0,
    i_10_275_1949_0, i_10_275_2005_0, i_10_275_2159_0, i_10_275_2199_0,
    i_10_275_2311_0, i_10_275_2312_0, i_10_275_2352_0, i_10_275_2353_0,
    i_10_275_2354_0, i_10_275_2355_0, i_10_275_2407_0, i_10_275_2473_0,
    i_10_275_2631_0, i_10_275_2632_0, i_10_275_2635_0, i_10_275_2656_0,
    i_10_275_2661_0, i_10_275_2663_0, i_10_275_2725_0, i_10_275_2730_0,
    i_10_275_2731_0, i_10_275_2827_0, i_10_275_2832_0, i_10_275_2834_0,
    i_10_275_2880_0, i_10_275_2881_0, i_10_275_2921_0, i_10_275_2923_0,
    i_10_275_2924_0, i_10_275_3075_0, i_10_275_3076_0, i_10_275_3094_0,
    i_10_275_3155_0, i_10_275_3385_0, i_10_275_3388_0, i_10_275_3389_0,
    i_10_275_3391_0, i_10_275_3392_0, i_10_275_3497_0, i_10_275_3541_0,
    i_10_275_3545_0, i_10_275_3551_0, i_10_275_3614_0, i_10_275_3783_0,
    i_10_275_3788_0, i_10_275_3835_0, i_10_275_3854_0, i_10_275_3856_0,
    i_10_275_3859_0, i_10_275_3860_0, i_10_275_3894_0, i_10_275_3982_0,
    i_10_275_3994_0, i_10_275_4050_0, i_10_275_4124_0, i_10_275_4220_0,
    i_10_275_4237_0, i_10_275_4270_0, i_10_275_4273_0, i_10_275_4564_0;
  output o_10_275_0_0;
  assign o_10_275_0_0 = ~((~i_10_275_283_0 & ((~i_10_275_1553_0 & ~i_10_275_2353_0 & ~i_10_275_3094_0 & ~i_10_275_3392_0 & ~i_10_275_3541_0) | (i_10_275_1652_0 & i_10_275_3614_0))) | (~i_10_275_328_0 & ~i_10_275_3385_0 & ((~i_10_275_1552_0 & ~i_10_275_1626_0 & ~i_10_275_2354_0 & ~i_10_275_2881_0) | (~i_10_275_799_0 & ~i_10_275_1556_0 & ~i_10_275_3075_0 & ~i_10_275_3545_0 & ~i_10_275_3783_0 & ~i_10_275_4220_0 & ~i_10_275_4270_0))) | (~i_10_275_4220_0 & ((~i_10_275_458_0 & ((i_10_275_176_0 & ~i_10_275_1553_0 & ~i_10_275_2355_0 & ~i_10_275_2656_0 & ~i_10_275_2881_0 & ~i_10_275_3541_0 & ~i_10_275_3545_0 & ~i_10_275_3788_0) | (~i_10_275_1547_0 & ~i_10_275_2005_0 & ~i_10_275_2827_0 & ~i_10_275_3076_0 & ~i_10_275_3391_0 & ~i_10_275_4237_0))) | (~i_10_275_1552_0 & ((~i_10_275_329_0 & ~i_10_275_1821_0 & ~i_10_275_2311_0 & ~i_10_275_2473_0 & ~i_10_275_3392_0 & ~i_10_275_3545_0 & ~i_10_275_3835_0 & ~i_10_275_4124_0 & ~i_10_275_4270_0) | (~i_10_275_1553_0 & ~i_10_275_1691_0 & i_10_275_2725_0 & ~i_10_275_3075_0 & ~i_10_275_3076_0 & ~i_10_275_4273_0))))) | (~i_10_275_3835_0 & ((i_10_275_464_0 & (~i_10_275_2352_0 | i_10_275_3614_0)) | (i_10_275_463_0 & ~i_10_275_1825_0 & ~i_10_275_2312_0 & ~i_10_275_2355_0 & ~i_10_275_2407_0))) | (i_10_275_466_0 & ((~i_10_275_1312_0 & ~i_10_275_1556_0 & ~i_10_275_2311_0 & ~i_10_275_3075_0 & ~i_10_275_3389_0) | (i_10_275_1825_0 & ~i_10_275_2355_0 & i_10_275_2635_0 & ~i_10_275_2924_0 & ~i_10_275_3497_0 & ~i_10_275_3614_0))) | (~i_10_275_1547_0 & ((~i_10_275_178_0 & ((i_10_275_2731_0 & ~i_10_275_3392_0 & i_10_275_3856_0) | (~i_10_275_176_0 & ~i_10_275_959_0 & ~i_10_275_1002_0 & ~i_10_275_1652_0 & ~i_10_275_2312_0 & ~i_10_275_3076_0 & ~i_10_275_3854_0 & ~i_10_275_3982_0))) | (~i_10_275_329_0 & ~i_10_275_1556_0 & ~i_10_275_2352_0 & ~i_10_275_3389_0 & ~i_10_275_3391_0) | (~i_10_275_1002_0 & ~i_10_275_1307_0 & ~i_10_275_1555_0 & ~i_10_275_2311_0 & ~i_10_275_3076_0 & ~i_10_275_3392_0 & ~i_10_275_3551_0 & ~i_10_275_4237_0))) | (~i_10_275_329_0 & ((~i_10_275_2312_0 & ~i_10_275_2355_0 & i_10_275_2661_0) | (~i_10_275_1626_0 & ~i_10_275_2352_0 & ~i_10_275_2354_0 & i_10_275_2923_0))) | (~i_10_275_1556_0 & ((~i_10_275_1652_0 & ~i_10_275_1822_0 & ~i_10_275_2312_0 & i_10_275_3859_0) | (~i_10_275_412_0 & ~i_10_275_1691_0 & ~i_10_275_2631_0 & ~i_10_275_2632_0 & ~i_10_275_3075_0 & i_10_275_3391_0 & ~i_10_275_3497_0 & ~i_10_275_3545_0 & ~i_10_275_3860_0 & ~i_10_275_4124_0))) | (~i_10_275_3854_0 & ((~i_10_275_2631_0 & i_10_275_2827_0 & ((i_10_275_329_0 & ~i_10_275_463_0 & ~i_10_275_467_0 & i_10_275_1307_0 & i_10_275_2407_0) | (i_10_275_2352_0 & i_10_275_4124_0))) | (~i_10_275_466_0 & ~i_10_275_1233_0 & i_10_275_1825_0 & ~i_10_275_2005_0 & ~i_10_275_2354_0))) | (~i_10_275_2312_0 & ((~i_10_275_2354_0 & (i_10_275_3860_0 | (~i_10_275_178_0 & ~i_10_275_1626_0 & ~i_10_275_2407_0 & ~i_10_275_2632_0 & ~i_10_275_3788_0))) | (~i_10_275_3075_0 & ((i_10_275_799_0 & ~i_10_275_2311_0 & ~i_10_275_2632_0 & ~i_10_275_3392_0 & ~i_10_275_3497_0 & ~i_10_275_3856_0) | (i_10_275_962_0 & ~i_10_275_1552_0 & ~i_10_275_3545_0 & ~i_10_275_3859_0 & ~i_10_275_4564_0))) | (~i_10_275_284_0 & ~i_10_275_2473_0 & ~i_10_275_2656_0 & i_10_275_2881_0 & ~i_10_275_3545_0))) | (i_10_275_2924_0 & i_10_275_3094_0 & i_10_275_3389_0) | (i_10_275_1652_0 & ~i_10_275_3783_0 & i_10_275_3859_0));
endmodule



// Benchmark "kernel_10_276" written by ABC on Sun Jul 19 10:25:47 2020

module kernel_10_276 ( 
    i_10_276_160_0, i_10_276_259_0, i_10_276_282_0, i_10_276_283_0,
    i_10_276_315_0, i_10_276_320_0, i_10_276_328_0, i_10_276_367_0,
    i_10_276_393_0, i_10_276_425_0, i_10_276_436_0, i_10_276_445_0,
    i_10_276_446_0, i_10_276_447_0, i_10_276_463_0, i_10_276_464_0,
    i_10_276_715_0, i_10_276_750_0, i_10_276_864_0, i_10_276_1005_0,
    i_10_276_1104_0, i_10_276_1237_0, i_10_276_1296_0, i_10_276_1308_0,
    i_10_276_1309_0, i_10_276_1341_0, i_10_276_1365_0, i_10_276_1432_0,
    i_10_276_1575_0, i_10_276_1576_0, i_10_276_1626_0, i_10_276_1648_0,
    i_10_276_1651_0, i_10_276_1653_0, i_10_276_1683_0, i_10_276_1684_0,
    i_10_276_1687_0, i_10_276_1688_0, i_10_276_1689_0, i_10_276_1690_0,
    i_10_276_1710_0, i_10_276_1711_0, i_10_276_1821_0, i_10_276_1824_0,
    i_10_276_1826_0, i_10_276_1995_0, i_10_276_2349_0, i_10_276_2362_0,
    i_10_276_2364_0, i_10_276_2365_0, i_10_276_2453_0, i_10_276_2456_0,
    i_10_276_2460_0, i_10_276_2463_0, i_10_276_2468_0, i_10_276_2479_0,
    i_10_276_2511_0, i_10_276_2513_0, i_10_276_2565_0, i_10_276_2628_0,
    i_10_276_2631_0, i_10_276_2633_0, i_10_276_2657_0, i_10_276_2658_0,
    i_10_276_2660_0, i_10_276_2728_0, i_10_276_2731_0, i_10_276_2742_0,
    i_10_276_2754_0, i_10_276_2830_0, i_10_276_2831_0, i_10_276_2834_0,
    i_10_276_2869_0, i_10_276_2924_0, i_10_276_2953_0, i_10_276_2976_0,
    i_10_276_3036_0, i_10_276_3038_0, i_10_276_3075_0, i_10_276_3268_0,
    i_10_276_3280_0, i_10_276_3281_0, i_10_276_3501_0, i_10_276_3537_0,
    i_10_276_3582_0, i_10_276_3610_0, i_10_276_3611_0, i_10_276_3855_0,
    i_10_276_3856_0, i_10_276_3858_0, i_10_276_3860_0, i_10_276_3893_0,
    i_10_276_3919_0, i_10_276_4114_0, i_10_276_4116_0, i_10_276_4123_0,
    i_10_276_4156_0, i_10_276_4167_0, i_10_276_4275_0, i_10_276_4582_0,
    o_10_276_0_0  );
  input  i_10_276_160_0, i_10_276_259_0, i_10_276_282_0, i_10_276_283_0,
    i_10_276_315_0, i_10_276_320_0, i_10_276_328_0, i_10_276_367_0,
    i_10_276_393_0, i_10_276_425_0, i_10_276_436_0, i_10_276_445_0,
    i_10_276_446_0, i_10_276_447_0, i_10_276_463_0, i_10_276_464_0,
    i_10_276_715_0, i_10_276_750_0, i_10_276_864_0, i_10_276_1005_0,
    i_10_276_1104_0, i_10_276_1237_0, i_10_276_1296_0, i_10_276_1308_0,
    i_10_276_1309_0, i_10_276_1341_0, i_10_276_1365_0, i_10_276_1432_0,
    i_10_276_1575_0, i_10_276_1576_0, i_10_276_1626_0, i_10_276_1648_0,
    i_10_276_1651_0, i_10_276_1653_0, i_10_276_1683_0, i_10_276_1684_0,
    i_10_276_1687_0, i_10_276_1688_0, i_10_276_1689_0, i_10_276_1690_0,
    i_10_276_1710_0, i_10_276_1711_0, i_10_276_1821_0, i_10_276_1824_0,
    i_10_276_1826_0, i_10_276_1995_0, i_10_276_2349_0, i_10_276_2362_0,
    i_10_276_2364_0, i_10_276_2365_0, i_10_276_2453_0, i_10_276_2456_0,
    i_10_276_2460_0, i_10_276_2463_0, i_10_276_2468_0, i_10_276_2479_0,
    i_10_276_2511_0, i_10_276_2513_0, i_10_276_2565_0, i_10_276_2628_0,
    i_10_276_2631_0, i_10_276_2633_0, i_10_276_2657_0, i_10_276_2658_0,
    i_10_276_2660_0, i_10_276_2728_0, i_10_276_2731_0, i_10_276_2742_0,
    i_10_276_2754_0, i_10_276_2830_0, i_10_276_2831_0, i_10_276_2834_0,
    i_10_276_2869_0, i_10_276_2924_0, i_10_276_2953_0, i_10_276_2976_0,
    i_10_276_3036_0, i_10_276_3038_0, i_10_276_3075_0, i_10_276_3268_0,
    i_10_276_3280_0, i_10_276_3281_0, i_10_276_3501_0, i_10_276_3537_0,
    i_10_276_3582_0, i_10_276_3610_0, i_10_276_3611_0, i_10_276_3855_0,
    i_10_276_3856_0, i_10_276_3858_0, i_10_276_3860_0, i_10_276_3893_0,
    i_10_276_3919_0, i_10_276_4114_0, i_10_276_4116_0, i_10_276_4123_0,
    i_10_276_4156_0, i_10_276_4167_0, i_10_276_4275_0, i_10_276_4582_0;
  output o_10_276_0_0;
  assign o_10_276_0_0 = 0;
endmodule



// Benchmark "kernel_10_277" written by ABC on Sun Jul 19 10:25:47 2020

module kernel_10_277 ( 
    i_10_277_47_0, i_10_277_179_0, i_10_277_254_0, i_10_277_281_0,
    i_10_277_285_0, i_10_277_388_0, i_10_277_391_0, i_10_277_406_0,
    i_10_277_506_0, i_10_277_542_0, i_10_277_560_0, i_10_277_623_0,
    i_10_277_712_0, i_10_277_983_0, i_10_277_1000_0, i_10_277_1001_0,
    i_10_277_1003_0, i_10_277_1028_0, i_10_277_1100_0, i_10_277_1190_0,
    i_10_277_1207_0, i_10_277_1243_0, i_10_277_1280_0, i_10_277_1362_0,
    i_10_277_1363_0, i_10_277_1366_0, i_10_277_1397_0, i_10_277_1436_0,
    i_10_277_1541_0, i_10_277_1568_0, i_10_277_1577_0, i_10_277_1582_0,
    i_10_277_1613_0, i_10_277_1654_0, i_10_277_1655_0, i_10_277_1687_0,
    i_10_277_1688_0, i_10_277_1693_0, i_10_277_1730_0, i_10_277_1819_0,
    i_10_277_1820_0, i_10_277_1826_0, i_10_277_1828_0, i_10_277_1955_0,
    i_10_277_2020_0, i_10_277_2027_0, i_10_277_2350_0, i_10_277_2362_0,
    i_10_277_2365_0, i_10_277_2377_0, i_10_277_2435_0, i_10_277_2467_0,
    i_10_277_2470_0, i_10_277_2476_0, i_10_277_2531_0, i_10_277_2533_0,
    i_10_277_2534_0, i_10_277_2567_0, i_10_277_2661_0, i_10_277_2702_0,
    i_10_277_2705_0, i_10_277_2711_0, i_10_277_2713_0, i_10_277_2719_0,
    i_10_277_2755_0, i_10_277_2836_0, i_10_277_2846_0, i_10_277_2863_0,
    i_10_277_2867_0, i_10_277_3041_0, i_10_277_3042_0, i_10_277_3045_0,
    i_10_277_3074_0, i_10_277_3196_0, i_10_277_3232_0, i_10_277_3332_0,
    i_10_277_3350_0, i_10_277_3387_0, i_10_277_3388_0, i_10_277_3407_0,
    i_10_277_3439_0, i_10_277_3440_0, i_10_277_3449_0, i_10_277_3484_0,
    i_10_277_3503_0, i_10_277_3519_0, i_10_277_3609_0, i_10_277_3808_0,
    i_10_277_3837_0, i_10_277_3842_0, i_10_277_3908_0, i_10_277_3911_0,
    i_10_277_3982_0, i_10_277_4113_0, i_10_277_4114_0, i_10_277_4124_0,
    i_10_277_4145_0, i_10_277_4151_0, i_10_277_4268_0, i_10_277_4286_0,
    o_10_277_0_0  );
  input  i_10_277_47_0, i_10_277_179_0, i_10_277_254_0, i_10_277_281_0,
    i_10_277_285_0, i_10_277_388_0, i_10_277_391_0, i_10_277_406_0,
    i_10_277_506_0, i_10_277_542_0, i_10_277_560_0, i_10_277_623_0,
    i_10_277_712_0, i_10_277_983_0, i_10_277_1000_0, i_10_277_1001_0,
    i_10_277_1003_0, i_10_277_1028_0, i_10_277_1100_0, i_10_277_1190_0,
    i_10_277_1207_0, i_10_277_1243_0, i_10_277_1280_0, i_10_277_1362_0,
    i_10_277_1363_0, i_10_277_1366_0, i_10_277_1397_0, i_10_277_1436_0,
    i_10_277_1541_0, i_10_277_1568_0, i_10_277_1577_0, i_10_277_1582_0,
    i_10_277_1613_0, i_10_277_1654_0, i_10_277_1655_0, i_10_277_1687_0,
    i_10_277_1688_0, i_10_277_1693_0, i_10_277_1730_0, i_10_277_1819_0,
    i_10_277_1820_0, i_10_277_1826_0, i_10_277_1828_0, i_10_277_1955_0,
    i_10_277_2020_0, i_10_277_2027_0, i_10_277_2350_0, i_10_277_2362_0,
    i_10_277_2365_0, i_10_277_2377_0, i_10_277_2435_0, i_10_277_2467_0,
    i_10_277_2470_0, i_10_277_2476_0, i_10_277_2531_0, i_10_277_2533_0,
    i_10_277_2534_0, i_10_277_2567_0, i_10_277_2661_0, i_10_277_2702_0,
    i_10_277_2705_0, i_10_277_2711_0, i_10_277_2713_0, i_10_277_2719_0,
    i_10_277_2755_0, i_10_277_2836_0, i_10_277_2846_0, i_10_277_2863_0,
    i_10_277_2867_0, i_10_277_3041_0, i_10_277_3042_0, i_10_277_3045_0,
    i_10_277_3074_0, i_10_277_3196_0, i_10_277_3232_0, i_10_277_3332_0,
    i_10_277_3350_0, i_10_277_3387_0, i_10_277_3388_0, i_10_277_3407_0,
    i_10_277_3439_0, i_10_277_3440_0, i_10_277_3449_0, i_10_277_3484_0,
    i_10_277_3503_0, i_10_277_3519_0, i_10_277_3609_0, i_10_277_3808_0,
    i_10_277_3837_0, i_10_277_3842_0, i_10_277_3908_0, i_10_277_3911_0,
    i_10_277_3982_0, i_10_277_4113_0, i_10_277_4114_0, i_10_277_4124_0,
    i_10_277_4145_0, i_10_277_4151_0, i_10_277_4268_0, i_10_277_4286_0;
  output o_10_277_0_0;
  assign o_10_277_0_0 = 0;
endmodule



// Benchmark "kernel_10_278" written by ABC on Sun Jul 19 10:25:48 2020

module kernel_10_278 ( 
    i_10_278_21_0, i_10_278_22_0, i_10_278_23_0, i_10_278_27_0,
    i_10_278_55_0, i_10_278_82_0, i_10_278_171_0, i_10_278_270_0,
    i_10_278_373_0, i_10_278_460_0, i_10_278_461_0, i_10_278_468_0,
    i_10_278_469_0, i_10_278_477_0, i_10_278_478_0, i_10_278_495_0,
    i_10_278_498_0, i_10_278_567_0, i_10_278_568_0, i_10_278_569_0,
    i_10_278_675_0, i_10_278_676_0, i_10_278_730_0, i_10_278_901_0,
    i_10_278_945_0, i_10_278_999_0, i_10_278_1171_0, i_10_278_1235_0,
    i_10_278_1280_0, i_10_278_1368_0, i_10_278_1521_0, i_10_278_1522_0,
    i_10_278_1566_0, i_10_278_1569_0, i_10_278_1570_0, i_10_278_1690_0,
    i_10_278_1691_0, i_10_278_1728_0, i_10_278_1729_0, i_10_278_1737_0,
    i_10_278_1768_0, i_10_278_1845_0, i_10_278_1927_0, i_10_278_1944_0,
    i_10_278_1945_0, i_10_278_2025_0, i_10_278_2180_0, i_10_278_2244_0,
    i_10_278_2322_0, i_10_278_2325_0, i_10_278_2333_0, i_10_278_2334_0,
    i_10_278_2358_0, i_10_278_2538_0, i_10_278_2569_0, i_10_278_2602_0,
    i_10_278_2610_0, i_10_278_2709_0, i_10_278_2764_0, i_10_278_2817_0,
    i_10_278_2839_0, i_10_278_2919_0, i_10_278_2981_0, i_10_278_3025_0,
    i_10_278_3096_0, i_10_278_3186_0, i_10_278_3258_0, i_10_278_3268_0,
    i_10_278_3288_0, i_10_278_3357_0, i_10_278_3358_0, i_10_278_3359_0,
    i_10_278_3474_0, i_10_278_3583_0, i_10_278_3600_0, i_10_278_3601_0,
    i_10_278_3615_0, i_10_278_3651_0, i_10_278_3727_0, i_10_278_3799_0,
    i_10_278_3802_0, i_10_278_3850_0, i_10_278_3860_0, i_10_278_3861_0,
    i_10_278_3870_0, i_10_278_3892_0, i_10_278_3927_0, i_10_278_3942_0,
    i_10_278_4068_0, i_10_278_4069_0, i_10_278_4086_0, i_10_278_4095_0,
    i_10_278_4116_0, i_10_278_4185_0, i_10_278_4231_0, i_10_278_4430_0,
    i_10_278_4432_0, i_10_278_4433_0, i_10_278_4437_0, i_10_278_4446_0,
    o_10_278_0_0  );
  input  i_10_278_21_0, i_10_278_22_0, i_10_278_23_0, i_10_278_27_0,
    i_10_278_55_0, i_10_278_82_0, i_10_278_171_0, i_10_278_270_0,
    i_10_278_373_0, i_10_278_460_0, i_10_278_461_0, i_10_278_468_0,
    i_10_278_469_0, i_10_278_477_0, i_10_278_478_0, i_10_278_495_0,
    i_10_278_498_0, i_10_278_567_0, i_10_278_568_0, i_10_278_569_0,
    i_10_278_675_0, i_10_278_676_0, i_10_278_730_0, i_10_278_901_0,
    i_10_278_945_0, i_10_278_999_0, i_10_278_1171_0, i_10_278_1235_0,
    i_10_278_1280_0, i_10_278_1368_0, i_10_278_1521_0, i_10_278_1522_0,
    i_10_278_1566_0, i_10_278_1569_0, i_10_278_1570_0, i_10_278_1690_0,
    i_10_278_1691_0, i_10_278_1728_0, i_10_278_1729_0, i_10_278_1737_0,
    i_10_278_1768_0, i_10_278_1845_0, i_10_278_1927_0, i_10_278_1944_0,
    i_10_278_1945_0, i_10_278_2025_0, i_10_278_2180_0, i_10_278_2244_0,
    i_10_278_2322_0, i_10_278_2325_0, i_10_278_2333_0, i_10_278_2334_0,
    i_10_278_2358_0, i_10_278_2538_0, i_10_278_2569_0, i_10_278_2602_0,
    i_10_278_2610_0, i_10_278_2709_0, i_10_278_2764_0, i_10_278_2817_0,
    i_10_278_2839_0, i_10_278_2919_0, i_10_278_2981_0, i_10_278_3025_0,
    i_10_278_3096_0, i_10_278_3186_0, i_10_278_3258_0, i_10_278_3268_0,
    i_10_278_3288_0, i_10_278_3357_0, i_10_278_3358_0, i_10_278_3359_0,
    i_10_278_3474_0, i_10_278_3583_0, i_10_278_3600_0, i_10_278_3601_0,
    i_10_278_3615_0, i_10_278_3651_0, i_10_278_3727_0, i_10_278_3799_0,
    i_10_278_3802_0, i_10_278_3850_0, i_10_278_3860_0, i_10_278_3861_0,
    i_10_278_3870_0, i_10_278_3892_0, i_10_278_3927_0, i_10_278_3942_0,
    i_10_278_4068_0, i_10_278_4069_0, i_10_278_4086_0, i_10_278_4095_0,
    i_10_278_4116_0, i_10_278_4185_0, i_10_278_4231_0, i_10_278_4430_0,
    i_10_278_4432_0, i_10_278_4433_0, i_10_278_4437_0, i_10_278_4446_0;
  output o_10_278_0_0;
  assign o_10_278_0_0 = 0;
endmodule



// Benchmark "kernel_10_279" written by ABC on Sun Jul 19 10:25:49 2020

module kernel_10_279 ( 
    i_10_279_33_0, i_10_279_34_0, i_10_279_40_0, i_10_279_82_0,
    i_10_279_124_0, i_10_279_185_0, i_10_279_187_0, i_10_279_196_0,
    i_10_279_272_0, i_10_279_275_0, i_10_279_282_0, i_10_279_321_0,
    i_10_279_374_0, i_10_279_390_0, i_10_279_393_0, i_10_279_394_0,
    i_10_279_465_0, i_10_279_499_0, i_10_279_564_0, i_10_279_629_0,
    i_10_279_700_0, i_10_279_906_0, i_10_279_988_0, i_10_279_1048_0,
    i_10_279_1201_0, i_10_279_1234_0, i_10_279_1241_0, i_10_279_1249_0,
    i_10_279_1312_0, i_10_279_1365_0, i_10_279_1366_0, i_10_279_1543_0,
    i_10_279_1547_0, i_10_279_1641_0, i_10_279_1646_0, i_10_279_1651_0,
    i_10_279_1756_0, i_10_279_1905_0, i_10_279_1906_0, i_10_279_1930_0,
    i_10_279_1931_0, i_10_279_1933_0, i_10_279_1934_0, i_10_279_1941_0,
    i_10_279_1942_0, i_10_279_1951_0, i_10_279_1952_0, i_10_279_2094_0,
    i_10_279_2095_0, i_10_279_2245_0, i_10_279_2275_0, i_10_279_2276_0,
    i_10_279_2330_0, i_10_279_2380_0, i_10_279_2464_0, i_10_279_2515_0,
    i_10_279_2518_0, i_10_279_2632_0, i_10_279_2678_0, i_10_279_2726_0,
    i_10_279_2823_0, i_10_279_2851_0, i_10_279_2947_0, i_10_279_2982_0,
    i_10_279_2986_0, i_10_279_3050_0, i_10_279_3076_0, i_10_279_3093_0,
    i_10_279_3100_0, i_10_279_3208_0, i_10_279_3315_0, i_10_279_3316_0,
    i_10_279_3356_0, i_10_279_3392_0, i_10_279_3466_0, i_10_279_3471_0,
    i_10_279_3472_0, i_10_279_3495_0, i_10_279_3544_0, i_10_279_3585_0,
    i_10_279_3588_0, i_10_279_3589_0, i_10_279_3613_0, i_10_279_3624_0,
    i_10_279_3625_0, i_10_279_3649_0, i_10_279_3653_0, i_10_279_3751_0,
    i_10_279_3805_0, i_10_279_3931_0, i_10_279_3985_0, i_10_279_4189_0,
    i_10_279_4237_0, i_10_279_4287_0, i_10_279_4292_0, i_10_279_4524_0,
    i_10_279_4525_0, i_10_279_4526_0, i_10_279_4533_0, i_10_279_4534_0,
    o_10_279_0_0  );
  input  i_10_279_33_0, i_10_279_34_0, i_10_279_40_0, i_10_279_82_0,
    i_10_279_124_0, i_10_279_185_0, i_10_279_187_0, i_10_279_196_0,
    i_10_279_272_0, i_10_279_275_0, i_10_279_282_0, i_10_279_321_0,
    i_10_279_374_0, i_10_279_390_0, i_10_279_393_0, i_10_279_394_0,
    i_10_279_465_0, i_10_279_499_0, i_10_279_564_0, i_10_279_629_0,
    i_10_279_700_0, i_10_279_906_0, i_10_279_988_0, i_10_279_1048_0,
    i_10_279_1201_0, i_10_279_1234_0, i_10_279_1241_0, i_10_279_1249_0,
    i_10_279_1312_0, i_10_279_1365_0, i_10_279_1366_0, i_10_279_1543_0,
    i_10_279_1547_0, i_10_279_1641_0, i_10_279_1646_0, i_10_279_1651_0,
    i_10_279_1756_0, i_10_279_1905_0, i_10_279_1906_0, i_10_279_1930_0,
    i_10_279_1931_0, i_10_279_1933_0, i_10_279_1934_0, i_10_279_1941_0,
    i_10_279_1942_0, i_10_279_1951_0, i_10_279_1952_0, i_10_279_2094_0,
    i_10_279_2095_0, i_10_279_2245_0, i_10_279_2275_0, i_10_279_2276_0,
    i_10_279_2330_0, i_10_279_2380_0, i_10_279_2464_0, i_10_279_2515_0,
    i_10_279_2518_0, i_10_279_2632_0, i_10_279_2678_0, i_10_279_2726_0,
    i_10_279_2823_0, i_10_279_2851_0, i_10_279_2947_0, i_10_279_2982_0,
    i_10_279_2986_0, i_10_279_3050_0, i_10_279_3076_0, i_10_279_3093_0,
    i_10_279_3100_0, i_10_279_3208_0, i_10_279_3315_0, i_10_279_3316_0,
    i_10_279_3356_0, i_10_279_3392_0, i_10_279_3466_0, i_10_279_3471_0,
    i_10_279_3472_0, i_10_279_3495_0, i_10_279_3544_0, i_10_279_3585_0,
    i_10_279_3588_0, i_10_279_3589_0, i_10_279_3613_0, i_10_279_3624_0,
    i_10_279_3625_0, i_10_279_3649_0, i_10_279_3653_0, i_10_279_3751_0,
    i_10_279_3805_0, i_10_279_3931_0, i_10_279_3985_0, i_10_279_4189_0,
    i_10_279_4237_0, i_10_279_4287_0, i_10_279_4292_0, i_10_279_4524_0,
    i_10_279_4525_0, i_10_279_4526_0, i_10_279_4533_0, i_10_279_4534_0;
  output o_10_279_0_0;
  assign o_10_279_0_0 = 0;
endmodule



// Benchmark "kernel_10_280" written by ABC on Sun Jul 19 10:25:50 2020

module kernel_10_280 ( 
    i_10_280_27_0, i_10_280_117_0, i_10_280_207_0, i_10_280_262_0,
    i_10_280_282_0, i_10_280_283_0, i_10_280_284_0, i_10_280_287_0,
    i_10_280_325_0, i_10_280_369_0, i_10_280_390_0, i_10_280_423_0,
    i_10_280_426_0, i_10_280_433_0, i_10_280_434_0, i_10_280_558_0,
    i_10_280_730_0, i_10_280_793_0, i_10_280_797_0, i_10_280_945_0,
    i_10_280_958_0, i_10_280_969_0, i_10_280_996_0, i_10_280_1044_0,
    i_10_280_1163_0, i_10_280_1236_0, i_10_280_1341_0, i_10_280_1359_0,
    i_10_280_1377_0, i_10_280_1449_0, i_10_280_1450_0, i_10_280_1494_0,
    i_10_280_1611_0, i_10_280_1620_0, i_10_280_1630_0, i_10_280_1651_0,
    i_10_280_1684_0, i_10_280_1686_0, i_10_280_1689_0, i_10_280_1768_0,
    i_10_280_1818_0, i_10_280_1820_0, i_10_280_1822_0, i_10_280_1823_0,
    i_10_280_1825_0, i_10_280_1899_0, i_10_280_1944_0, i_10_280_2019_0,
    i_10_280_2089_0, i_10_280_2091_0, i_10_280_2178_0, i_10_280_2350_0,
    i_10_280_2403_0, i_10_280_2502_0, i_10_280_2505_0, i_10_280_2514_0,
    i_10_280_2601_0, i_10_280_2610_0, i_10_280_2611_0, i_10_280_2655_0,
    i_10_280_2661_0, i_10_280_2673_0, i_10_280_2700_0, i_10_280_2721_0,
    i_10_280_2729_0, i_10_280_2784_0, i_10_280_2817_0, i_10_280_2880_0,
    i_10_280_2907_0, i_10_280_2919_0, i_10_280_3036_0, i_10_280_3198_0,
    i_10_280_3231_0, i_10_280_3384_0, i_10_280_3385_0, i_10_280_3387_0,
    i_10_280_3402_0, i_10_280_3409_0, i_10_280_3468_0, i_10_280_3496_0,
    i_10_280_3555_0, i_10_280_3590_0, i_10_280_3618_0, i_10_280_3646_0,
    i_10_280_3786_0, i_10_280_3787_0, i_10_280_3837_0, i_10_280_3851_0,
    i_10_280_3895_0, i_10_280_3942_0, i_10_280_3978_0, i_10_280_3979_0,
    i_10_280_4053_0, i_10_280_4125_0, i_10_280_4176_0, i_10_280_4230_0,
    i_10_280_4419_0, i_10_280_4527_0, i_10_280_4567_0, i_10_280_4581_0,
    o_10_280_0_0  );
  input  i_10_280_27_0, i_10_280_117_0, i_10_280_207_0, i_10_280_262_0,
    i_10_280_282_0, i_10_280_283_0, i_10_280_284_0, i_10_280_287_0,
    i_10_280_325_0, i_10_280_369_0, i_10_280_390_0, i_10_280_423_0,
    i_10_280_426_0, i_10_280_433_0, i_10_280_434_0, i_10_280_558_0,
    i_10_280_730_0, i_10_280_793_0, i_10_280_797_0, i_10_280_945_0,
    i_10_280_958_0, i_10_280_969_0, i_10_280_996_0, i_10_280_1044_0,
    i_10_280_1163_0, i_10_280_1236_0, i_10_280_1341_0, i_10_280_1359_0,
    i_10_280_1377_0, i_10_280_1449_0, i_10_280_1450_0, i_10_280_1494_0,
    i_10_280_1611_0, i_10_280_1620_0, i_10_280_1630_0, i_10_280_1651_0,
    i_10_280_1684_0, i_10_280_1686_0, i_10_280_1689_0, i_10_280_1768_0,
    i_10_280_1818_0, i_10_280_1820_0, i_10_280_1822_0, i_10_280_1823_0,
    i_10_280_1825_0, i_10_280_1899_0, i_10_280_1944_0, i_10_280_2019_0,
    i_10_280_2089_0, i_10_280_2091_0, i_10_280_2178_0, i_10_280_2350_0,
    i_10_280_2403_0, i_10_280_2502_0, i_10_280_2505_0, i_10_280_2514_0,
    i_10_280_2601_0, i_10_280_2610_0, i_10_280_2611_0, i_10_280_2655_0,
    i_10_280_2661_0, i_10_280_2673_0, i_10_280_2700_0, i_10_280_2721_0,
    i_10_280_2729_0, i_10_280_2784_0, i_10_280_2817_0, i_10_280_2880_0,
    i_10_280_2907_0, i_10_280_2919_0, i_10_280_3036_0, i_10_280_3198_0,
    i_10_280_3231_0, i_10_280_3384_0, i_10_280_3385_0, i_10_280_3387_0,
    i_10_280_3402_0, i_10_280_3409_0, i_10_280_3468_0, i_10_280_3496_0,
    i_10_280_3555_0, i_10_280_3590_0, i_10_280_3618_0, i_10_280_3646_0,
    i_10_280_3786_0, i_10_280_3787_0, i_10_280_3837_0, i_10_280_3851_0,
    i_10_280_3895_0, i_10_280_3942_0, i_10_280_3978_0, i_10_280_3979_0,
    i_10_280_4053_0, i_10_280_4125_0, i_10_280_4176_0, i_10_280_4230_0,
    i_10_280_4419_0, i_10_280_4527_0, i_10_280_4567_0, i_10_280_4581_0;
  output o_10_280_0_0;
  assign o_10_280_0_0 = ~((~i_10_280_797_0 & ((~i_10_280_426_0 & ~i_10_280_1359_0 & ~i_10_280_2505_0 & ~i_10_280_2919_0 & ~i_10_280_3468_0 & ~i_10_280_3942_0) | (i_10_280_1825_0 & i_10_280_2610_0 & ~i_10_280_2611_0 & i_10_280_4567_0))) | (~i_10_280_958_0 & ((~i_10_280_1823_0 & ~i_10_280_2610_0 & ~i_10_280_2611_0 & i_10_280_3646_0 & ~i_10_280_4125_0) | (~i_10_280_2502_0 & i_10_280_2729_0 & ~i_10_280_3231_0 & ~i_10_280_4230_0))) | (~i_10_280_2502_0 & ((~i_10_280_1163_0 & ((~i_10_280_558_0 & ~i_10_280_1359_0 & ~i_10_280_1818_0 & ~i_10_280_1820_0 & ~i_10_280_2178_0) | (~i_10_280_2019_0 & ~i_10_280_2505_0 & ~i_10_280_2700_0))) | (~i_10_280_1823_0 & ~i_10_280_1825_0 & ~i_10_280_2610_0 & ~i_10_280_2673_0))) | (~i_10_280_1341_0 & ((~i_10_280_27_0 & ~i_10_280_1651_0 & ~i_10_280_1689_0 & i_10_280_1825_0 & i_10_280_2403_0) | (~i_10_280_996_0 & ~i_10_280_1359_0 & ~i_10_280_1620_0 & ~i_10_280_2601_0 & ~i_10_280_2655_0 & ~i_10_280_4230_0))) | (~i_10_280_1359_0 & ((~i_10_280_2403_0 & ~i_10_280_2505_0 & ~i_10_280_2673_0 & ~i_10_280_3646_0) | (~i_10_280_2721_0 & i_10_280_2729_0 & ~i_10_280_3786_0 & ~i_10_280_3851_0 & i_10_280_3978_0 & ~i_10_280_4053_0))) | (~i_10_280_1611_0 & ~i_10_280_4125_0 & (i_10_280_2655_0 | (~i_10_280_1822_0 & ~i_10_280_3036_0 & ~i_10_280_3851_0 & ~i_10_280_3942_0))) | (i_10_280_434_0 & ~i_10_280_2611_0) | (~i_10_280_2610_0 & ~i_10_280_4230_0 & ~i_10_280_4567_0));
endmodule



// Benchmark "kernel_10_281" written by ABC on Sun Jul 19 10:25:51 2020

module kernel_10_281 ( 
    i_10_281_40_0, i_10_281_171_0, i_10_281_174_0, i_10_281_253_0,
    i_10_281_280_0, i_10_281_282_0, i_10_281_283_0, i_10_281_424_0,
    i_10_281_444_0, i_10_281_463_0, i_10_281_464_0, i_10_281_713_0,
    i_10_281_749_0, i_10_281_820_0, i_10_281_967_0, i_10_281_1027_0,
    i_10_281_1028_0, i_10_281_1040_0, i_10_281_1235_0, i_10_281_1236_0,
    i_10_281_1237_0, i_10_281_1243_0, i_10_281_1296_0, i_10_281_1305_0,
    i_10_281_1359_0, i_10_281_1444_0, i_10_281_1540_0, i_10_281_1541_0,
    i_10_281_1650_0, i_10_281_1683_0, i_10_281_1684_0, i_10_281_1686_0,
    i_10_281_1687_0, i_10_281_1691_0, i_10_281_1730_0, i_10_281_1765_0,
    i_10_281_1801_0, i_10_281_1821_0, i_10_281_1824_0, i_10_281_1954_0,
    i_10_281_2027_0, i_10_281_2199_0, i_10_281_2350_0, i_10_281_2467_0,
    i_10_281_2470_0, i_10_281_2557_0, i_10_281_2566_0, i_10_281_2602_0,
    i_10_281_2628_0, i_10_281_2631_0, i_10_281_2632_0, i_10_281_2633_0,
    i_10_281_2659_0, i_10_281_2728_0, i_10_281_2731_0, i_10_281_2818_0,
    i_10_281_2828_0, i_10_281_2920_0, i_10_281_2921_0, i_10_281_3037_0,
    i_10_281_3070_0, i_10_281_3198_0, i_10_281_3199_0, i_10_281_3200_0,
    i_10_281_3277_0, i_10_281_3278_0, i_10_281_3281_0, i_10_281_3386_0,
    i_10_281_3389_0, i_10_281_3406_0, i_10_281_3407_0, i_10_281_3522_0,
    i_10_281_3523_0, i_10_281_3538_0, i_10_281_3541_0, i_10_281_3584_0,
    i_10_281_3613_0, i_10_281_3615_0, i_10_281_3646_0, i_10_281_3650_0,
    i_10_281_3781_0, i_10_281_3782_0, i_10_281_3784_0, i_10_281_3837_0,
    i_10_281_3846_0, i_10_281_3853_0, i_10_281_3854_0, i_10_281_3856_0,
    i_10_281_3857_0, i_10_281_4115_0, i_10_281_4121_0, i_10_281_4171_0,
    i_10_281_4204_0, i_10_281_4267_0, i_10_281_4275_0, i_10_281_4276_0,
    i_10_281_4285_0, i_10_281_4286_0, i_10_281_4567_0, i_10_281_4582_0,
    o_10_281_0_0  );
  input  i_10_281_40_0, i_10_281_171_0, i_10_281_174_0, i_10_281_253_0,
    i_10_281_280_0, i_10_281_282_0, i_10_281_283_0, i_10_281_424_0,
    i_10_281_444_0, i_10_281_463_0, i_10_281_464_0, i_10_281_713_0,
    i_10_281_749_0, i_10_281_820_0, i_10_281_967_0, i_10_281_1027_0,
    i_10_281_1028_0, i_10_281_1040_0, i_10_281_1235_0, i_10_281_1236_0,
    i_10_281_1237_0, i_10_281_1243_0, i_10_281_1296_0, i_10_281_1305_0,
    i_10_281_1359_0, i_10_281_1444_0, i_10_281_1540_0, i_10_281_1541_0,
    i_10_281_1650_0, i_10_281_1683_0, i_10_281_1684_0, i_10_281_1686_0,
    i_10_281_1687_0, i_10_281_1691_0, i_10_281_1730_0, i_10_281_1765_0,
    i_10_281_1801_0, i_10_281_1821_0, i_10_281_1824_0, i_10_281_1954_0,
    i_10_281_2027_0, i_10_281_2199_0, i_10_281_2350_0, i_10_281_2467_0,
    i_10_281_2470_0, i_10_281_2557_0, i_10_281_2566_0, i_10_281_2602_0,
    i_10_281_2628_0, i_10_281_2631_0, i_10_281_2632_0, i_10_281_2633_0,
    i_10_281_2659_0, i_10_281_2728_0, i_10_281_2731_0, i_10_281_2818_0,
    i_10_281_2828_0, i_10_281_2920_0, i_10_281_2921_0, i_10_281_3037_0,
    i_10_281_3070_0, i_10_281_3198_0, i_10_281_3199_0, i_10_281_3200_0,
    i_10_281_3277_0, i_10_281_3278_0, i_10_281_3281_0, i_10_281_3386_0,
    i_10_281_3389_0, i_10_281_3406_0, i_10_281_3407_0, i_10_281_3522_0,
    i_10_281_3523_0, i_10_281_3538_0, i_10_281_3541_0, i_10_281_3584_0,
    i_10_281_3613_0, i_10_281_3615_0, i_10_281_3646_0, i_10_281_3650_0,
    i_10_281_3781_0, i_10_281_3782_0, i_10_281_3784_0, i_10_281_3837_0,
    i_10_281_3846_0, i_10_281_3853_0, i_10_281_3854_0, i_10_281_3856_0,
    i_10_281_3857_0, i_10_281_4115_0, i_10_281_4121_0, i_10_281_4171_0,
    i_10_281_4204_0, i_10_281_4267_0, i_10_281_4275_0, i_10_281_4276_0,
    i_10_281_4285_0, i_10_281_4286_0, i_10_281_4567_0, i_10_281_4582_0;
  output o_10_281_0_0;
  assign o_10_281_0_0 = 0;
endmodule



// Benchmark "kernel_10_282" written by ABC on Sun Jul 19 10:25:52 2020

module kernel_10_282 ( 
    i_10_282_64_0, i_10_282_144_0, i_10_282_177_0, i_10_282_189_0,
    i_10_282_190_0, i_10_282_275_0, i_10_282_315_0, i_10_282_369_0,
    i_10_282_388_0, i_10_282_391_0, i_10_282_443_0, i_10_282_447_0,
    i_10_282_459_0, i_10_282_460_0, i_10_282_463_0, i_10_282_465_0,
    i_10_282_535_0, i_10_282_536_0, i_10_282_585_0, i_10_282_588_0,
    i_10_282_698_0, i_10_282_700_0, i_10_282_800_0, i_10_282_967_0,
    i_10_282_994_0, i_10_282_1233_0, i_10_282_1290_0, i_10_282_1307_0,
    i_10_282_1312_0, i_10_282_1343_0, i_10_282_1417_0, i_10_282_1444_0,
    i_10_282_1447_0, i_10_282_1476_0, i_10_282_1551_0, i_10_282_1552_0,
    i_10_282_1556_0, i_10_282_1618_0, i_10_282_1648_0, i_10_282_1651_0,
    i_10_282_1801_0, i_10_282_1820_0, i_10_282_1826_0, i_10_282_1980_0,
    i_10_282_1982_0, i_10_282_2304_0, i_10_282_2305_0, i_10_282_2352_0,
    i_10_282_2430_0, i_10_282_2451_0, i_10_282_2514_0, i_10_282_2607_0,
    i_10_282_2608_0, i_10_282_2609_0, i_10_282_2629_0, i_10_282_2630_0,
    i_10_282_2641_0, i_10_282_2655_0, i_10_282_2660_0, i_10_282_2679_0,
    i_10_282_2722_0, i_10_282_2726_0, i_10_282_2734_0, i_10_282_2829_0,
    i_10_282_2830_0, i_10_282_2832_0, i_10_282_2923_0, i_10_282_3034_0,
    i_10_282_3036_0, i_10_282_3199_0, i_10_282_3271_0, i_10_282_3317_0,
    i_10_282_3402_0, i_10_282_3403_0, i_10_282_3405_0, i_10_282_3408_0,
    i_10_282_3469_0, i_10_282_3492_0, i_10_282_3493_0, i_10_282_3495_0,
    i_10_282_3523_0, i_10_282_3540_0, i_10_282_3639_0, i_10_282_3649_0,
    i_10_282_3682_0, i_10_282_3706_0, i_10_282_3846_0, i_10_282_3855_0,
    i_10_282_3857_0, i_10_282_3978_0, i_10_282_3979_0, i_10_282_3986_0,
    i_10_282_4030_0, i_10_282_4171_0, i_10_282_4266_0, i_10_282_4352_0,
    i_10_282_4354_0, i_10_282_4567_0, i_10_282_4582_0, i_10_282_4595_0,
    o_10_282_0_0  );
  input  i_10_282_64_0, i_10_282_144_0, i_10_282_177_0, i_10_282_189_0,
    i_10_282_190_0, i_10_282_275_0, i_10_282_315_0, i_10_282_369_0,
    i_10_282_388_0, i_10_282_391_0, i_10_282_443_0, i_10_282_447_0,
    i_10_282_459_0, i_10_282_460_0, i_10_282_463_0, i_10_282_465_0,
    i_10_282_535_0, i_10_282_536_0, i_10_282_585_0, i_10_282_588_0,
    i_10_282_698_0, i_10_282_700_0, i_10_282_800_0, i_10_282_967_0,
    i_10_282_994_0, i_10_282_1233_0, i_10_282_1290_0, i_10_282_1307_0,
    i_10_282_1312_0, i_10_282_1343_0, i_10_282_1417_0, i_10_282_1444_0,
    i_10_282_1447_0, i_10_282_1476_0, i_10_282_1551_0, i_10_282_1552_0,
    i_10_282_1556_0, i_10_282_1618_0, i_10_282_1648_0, i_10_282_1651_0,
    i_10_282_1801_0, i_10_282_1820_0, i_10_282_1826_0, i_10_282_1980_0,
    i_10_282_1982_0, i_10_282_2304_0, i_10_282_2305_0, i_10_282_2352_0,
    i_10_282_2430_0, i_10_282_2451_0, i_10_282_2514_0, i_10_282_2607_0,
    i_10_282_2608_0, i_10_282_2609_0, i_10_282_2629_0, i_10_282_2630_0,
    i_10_282_2641_0, i_10_282_2655_0, i_10_282_2660_0, i_10_282_2679_0,
    i_10_282_2722_0, i_10_282_2726_0, i_10_282_2734_0, i_10_282_2829_0,
    i_10_282_2830_0, i_10_282_2832_0, i_10_282_2923_0, i_10_282_3034_0,
    i_10_282_3036_0, i_10_282_3199_0, i_10_282_3271_0, i_10_282_3317_0,
    i_10_282_3402_0, i_10_282_3403_0, i_10_282_3405_0, i_10_282_3408_0,
    i_10_282_3469_0, i_10_282_3492_0, i_10_282_3493_0, i_10_282_3495_0,
    i_10_282_3523_0, i_10_282_3540_0, i_10_282_3639_0, i_10_282_3649_0,
    i_10_282_3682_0, i_10_282_3706_0, i_10_282_3846_0, i_10_282_3855_0,
    i_10_282_3857_0, i_10_282_3978_0, i_10_282_3979_0, i_10_282_3986_0,
    i_10_282_4030_0, i_10_282_4171_0, i_10_282_4266_0, i_10_282_4352_0,
    i_10_282_4354_0, i_10_282_4567_0, i_10_282_4582_0, i_10_282_4595_0;
  output o_10_282_0_0;
  assign o_10_282_0_0 = 0;
endmodule



// Benchmark "kernel_10_283" written by ABC on Sun Jul 19 10:25:53 2020

module kernel_10_283 ( 
    i_10_283_222_0, i_10_283_324_0, i_10_283_433_0, i_10_283_442_0,
    i_10_283_444_0, i_10_283_463_0, i_10_283_513_0, i_10_283_516_0,
    i_10_283_793_0, i_10_283_794_0, i_10_283_796_0, i_10_283_900_0,
    i_10_283_954_0, i_10_283_959_0, i_10_283_966_0, i_10_283_967_0,
    i_10_283_968_0, i_10_283_990_0, i_10_283_1027_0, i_10_283_1028_0,
    i_10_283_1031_0, i_10_283_1036_0, i_10_283_1235_0, i_10_283_1263_0,
    i_10_283_1359_0, i_10_283_1444_0, i_10_283_1651_0, i_10_283_1654_0,
    i_10_283_1683_0, i_10_283_1684_0, i_10_283_1689_0, i_10_283_1812_0,
    i_10_283_1818_0, i_10_283_1819_0, i_10_283_1823_0, i_10_283_1825_0,
    i_10_283_1872_0, i_10_283_2322_0, i_10_283_2325_0, i_10_283_2351_0,
    i_10_283_2356_0, i_10_283_2461_0, i_10_283_2502_0, i_10_283_2604_0,
    i_10_283_2635_0, i_10_283_2673_0, i_10_283_2674_0, i_10_283_2700_0,
    i_10_283_2701_0, i_10_283_2723_0, i_10_283_2781_0, i_10_283_2782_0,
    i_10_283_2817_0, i_10_283_2828_0, i_10_283_2919_0, i_10_283_2921_0,
    i_10_283_2979_0, i_10_283_2980_0, i_10_283_3043_0, i_10_283_3071_0,
    i_10_283_3073_0, i_10_283_3200_0, i_10_283_3201_0, i_10_283_3387_0,
    i_10_283_3389_0, i_10_283_3391_0, i_10_283_3405_0, i_10_283_3406_0,
    i_10_283_3519_0, i_10_283_3522_0, i_10_283_3582_0, i_10_283_3585_0,
    i_10_283_3684_0, i_10_283_3780_0, i_10_283_3781_0, i_10_283_3783_0,
    i_10_283_3784_0, i_10_283_3788_0, i_10_283_3838_0, i_10_283_3839_0,
    i_10_283_3841_0, i_10_283_3854_0, i_10_283_3855_0, i_10_283_3889_0,
    i_10_283_3979_0, i_10_283_3980_0, i_10_283_3991_0, i_10_283_4027_0,
    i_10_283_4030_0, i_10_283_4116_0, i_10_283_4117_0, i_10_283_4230_0,
    i_10_283_4266_0, i_10_283_4267_0, i_10_283_4285_0, i_10_283_4292_0,
    i_10_283_4458_0, i_10_283_4461_0, i_10_283_4564_0, i_10_283_4566_0,
    o_10_283_0_0  );
  input  i_10_283_222_0, i_10_283_324_0, i_10_283_433_0, i_10_283_442_0,
    i_10_283_444_0, i_10_283_463_0, i_10_283_513_0, i_10_283_516_0,
    i_10_283_793_0, i_10_283_794_0, i_10_283_796_0, i_10_283_900_0,
    i_10_283_954_0, i_10_283_959_0, i_10_283_966_0, i_10_283_967_0,
    i_10_283_968_0, i_10_283_990_0, i_10_283_1027_0, i_10_283_1028_0,
    i_10_283_1031_0, i_10_283_1036_0, i_10_283_1235_0, i_10_283_1263_0,
    i_10_283_1359_0, i_10_283_1444_0, i_10_283_1651_0, i_10_283_1654_0,
    i_10_283_1683_0, i_10_283_1684_0, i_10_283_1689_0, i_10_283_1812_0,
    i_10_283_1818_0, i_10_283_1819_0, i_10_283_1823_0, i_10_283_1825_0,
    i_10_283_1872_0, i_10_283_2322_0, i_10_283_2325_0, i_10_283_2351_0,
    i_10_283_2356_0, i_10_283_2461_0, i_10_283_2502_0, i_10_283_2604_0,
    i_10_283_2635_0, i_10_283_2673_0, i_10_283_2674_0, i_10_283_2700_0,
    i_10_283_2701_0, i_10_283_2723_0, i_10_283_2781_0, i_10_283_2782_0,
    i_10_283_2817_0, i_10_283_2828_0, i_10_283_2919_0, i_10_283_2921_0,
    i_10_283_2979_0, i_10_283_2980_0, i_10_283_3043_0, i_10_283_3071_0,
    i_10_283_3073_0, i_10_283_3200_0, i_10_283_3201_0, i_10_283_3387_0,
    i_10_283_3389_0, i_10_283_3391_0, i_10_283_3405_0, i_10_283_3406_0,
    i_10_283_3519_0, i_10_283_3522_0, i_10_283_3582_0, i_10_283_3585_0,
    i_10_283_3684_0, i_10_283_3780_0, i_10_283_3781_0, i_10_283_3783_0,
    i_10_283_3784_0, i_10_283_3788_0, i_10_283_3838_0, i_10_283_3839_0,
    i_10_283_3841_0, i_10_283_3854_0, i_10_283_3855_0, i_10_283_3889_0,
    i_10_283_3979_0, i_10_283_3980_0, i_10_283_3991_0, i_10_283_4027_0,
    i_10_283_4030_0, i_10_283_4116_0, i_10_283_4117_0, i_10_283_4230_0,
    i_10_283_4266_0, i_10_283_4267_0, i_10_283_4285_0, i_10_283_4292_0,
    i_10_283_4458_0, i_10_283_4461_0, i_10_283_4564_0, i_10_283_4566_0;
  output o_10_283_0_0;
  assign o_10_283_0_0 = ~((~i_10_283_4230_0 & ((~i_10_283_444_0 & ((~i_10_283_796_0 & ~i_10_283_990_0 & ~i_10_283_1036_0 & ~i_10_283_1444_0 & ~i_10_283_1812_0 & ~i_10_283_1872_0 & ~i_10_283_3387_0 & ~i_10_283_3781_0 & ~i_10_283_3854_0) | (~i_10_283_900_0 & ~i_10_283_966_0 & ~i_10_283_2674_0 & ~i_10_283_3522_0 & ~i_10_283_3788_0 & ~i_10_283_3889_0 & ~i_10_283_4030_0))) | (~i_10_283_900_0 & ((~i_10_283_1689_0 & ~i_10_283_1812_0 & i_10_283_1825_0 & ~i_10_283_1872_0 & ~i_10_283_2322_0 & ~i_10_283_2325_0 & ~i_10_283_2351_0 & ~i_10_283_2723_0 & ~i_10_283_3522_0) | (~i_10_283_954_0 & ~i_10_283_2356_0 & ~i_10_283_2674_0 & ~i_10_283_2979_0 & ~i_10_283_3841_0 & ~i_10_283_4117_0 & ~i_10_283_4266_0 & ~i_10_283_4564_0))) | (~i_10_283_966_0 & ((~i_10_283_513_0 & ~i_10_283_1359_0 & i_10_283_2635_0 & ~i_10_283_2980_0 & ~i_10_283_3522_0 & ~i_10_283_3841_0 & ~i_10_283_3854_0) | (~i_10_283_324_0 & ~i_10_283_1036_0 & ~i_10_283_1263_0 & ~i_10_283_1689_0 & ~i_10_283_1812_0 & ~i_10_283_2604_0 & ~i_10_283_2673_0 & ~i_10_283_2828_0 & ~i_10_283_3387_0 & ~i_10_283_3788_0 & ~i_10_283_3839_0 & ~i_10_283_4564_0))) | (~i_10_283_516_0 & ~i_10_283_1359_0 & ~i_10_283_2325_0 & ~i_10_283_2817_0 & ~i_10_283_3519_0 & ~i_10_283_4267_0))) | (~i_10_283_796_0 & ((~i_10_283_516_0 & ~i_10_283_1825_0 & ~i_10_283_2322_0 & ~i_10_283_2817_0 & ~i_10_283_3522_0 & ~i_10_283_4564_0) | (~i_10_283_900_0 & ~i_10_283_967_0 & ~i_10_283_2325_0 & ~i_10_283_2673_0 & ~i_10_283_2723_0 & ~i_10_283_3043_0 & ~i_10_283_3519_0 & ~i_10_283_3784_0 & ~i_10_283_4566_0))) | (~i_10_283_2322_0 & ((~i_10_283_4267_0 & ((~i_10_283_900_0 & ~i_10_283_2325_0 & ((~i_10_283_222_0 & ~i_10_283_1654_0 & ~i_10_283_1825_0 & ~i_10_283_2700_0 & ~i_10_283_3043_0 & ~i_10_283_3389_0 & ~i_10_283_3522_0 & ~i_10_283_3838_0) | (~i_10_283_968_0 & ~i_10_283_1263_0 & ~i_10_283_1651_0 & ~i_10_283_2502_0 & ~i_10_283_3991_0 & ~i_10_283_4117_0))) | (~i_10_283_513_0 & i_10_283_793_0 & i_10_283_1819_0 & ~i_10_283_2604_0 & ~i_10_283_2980_0 & ~i_10_283_3582_0 & ~i_10_283_3839_0))) | (~i_10_283_2700_0 & ((i_10_283_1036_0 & ~i_10_283_2635_0 & ~i_10_283_3980_0 & ~i_10_283_4564_0) | (~i_10_283_442_0 & ~i_10_283_1654_0 & ~i_10_283_3585_0 & i_10_283_4566_0))) | (~i_10_283_954_0 & ~i_10_283_966_0 & ~i_10_283_968_0 & ~i_10_283_1359_0 & ~i_10_283_1825_0 & ~i_10_283_1872_0 & ~i_10_283_2979_0 & ~i_10_283_2980_0 & ~i_10_283_3200_0 & ~i_10_283_3519_0 & ~i_10_283_3522_0))) | (~i_10_283_324_0 & ((~i_10_283_222_0 & ((~i_10_283_900_0 & ~i_10_283_966_0 & ~i_10_283_1651_0 & ~i_10_283_2673_0 & ~i_10_283_2980_0 & ~i_10_283_3889_0) | (~i_10_283_463_0 & ~i_10_283_513_0 & ~i_10_283_1444_0 & ~i_10_283_1818_0 & ~i_10_283_2351_0 & ~i_10_283_2782_0 & ~i_10_283_3200_0 & ~i_10_283_3519_0 & ~i_10_283_4266_0))) | (~i_10_283_513_0 & ~i_10_283_966_0 & ~i_10_283_1444_0 & ~i_10_283_2502_0 & ~i_10_283_2701_0 & ~i_10_283_3979_0 & ~i_10_283_3991_0))) | (i_10_283_4292_0 & ((i_10_283_2356_0 & ~i_10_283_2700_0) | (i_10_283_1825_0 & i_10_283_3389_0 & i_10_283_3585_0 & ~i_10_283_4267_0))) | (i_10_283_1036_0 & i_10_283_1819_0 & ~i_10_283_2919_0 & i_10_283_2921_0) | (i_10_283_794_0 & ~i_10_283_966_0 & ~i_10_283_1263_0 & ~i_10_283_1823_0 & i_10_283_2635_0 & ~i_10_283_2674_0 & ~i_10_283_3684_0 & ~i_10_283_3788_0 & ~i_10_283_3839_0 & ~i_10_283_4266_0));
endmodule



// Benchmark "kernel_10_284" written by ABC on Sun Jul 19 10:25:54 2020

module kernel_10_284 ( 
    i_10_284_65_0, i_10_284_178_0, i_10_284_181_0, i_10_284_220_0,
    i_10_284_280_0, i_10_284_425_0, i_10_284_434_0, i_10_284_448_0,
    i_10_284_460_0, i_10_284_796_0, i_10_284_1036_0, i_10_284_1200_0,
    i_10_284_1233_0, i_10_284_1234_0, i_10_284_1240_0, i_10_284_1242_0,
    i_10_284_1342_0, i_10_284_1359_0, i_10_284_1550_0, i_10_284_1576_0,
    i_10_284_1651_0, i_10_284_1819_0, i_10_284_1913_0, i_10_284_1945_0,
    i_10_284_1946_0, i_10_284_1949_0, i_10_284_1991_0, i_10_284_2178_0,
    i_10_284_2179_0, i_10_284_2305_0, i_10_284_2306_0, i_10_284_2324_0,
    i_10_284_2333_0, i_10_284_2354_0, i_10_284_2358_0, i_10_284_2359_0,
    i_10_284_2362_0, i_10_284_2363_0, i_10_284_2378_0, i_10_284_2381_0,
    i_10_284_2404_0, i_10_284_2451_0, i_10_284_2453_0, i_10_284_2463_0,
    i_10_284_2467_0, i_10_284_2475_0, i_10_284_2476_0, i_10_284_2503_0,
    i_10_284_2628_0, i_10_284_2634_0, i_10_284_2635_0, i_10_284_2659_0,
    i_10_284_2660_0, i_10_284_2674_0, i_10_284_2704_0, i_10_284_2709_0,
    i_10_284_2710_0, i_10_284_2711_0, i_10_284_2721_0, i_10_284_2727_0,
    i_10_284_2730_0, i_10_284_2731_0, i_10_284_2732_0, i_10_284_2828_0,
    i_10_284_2886_0, i_10_284_2916_0, i_10_284_2924_0, i_10_284_3034_0,
    i_10_284_3035_0, i_10_284_3040_0, i_10_284_3087_0, i_10_284_3088_0,
    i_10_284_3203_0, i_10_284_3268_0, i_10_284_3269_0, i_10_284_3384_0,
    i_10_284_3403_0, i_10_284_3404_0, i_10_284_3405_0, i_10_284_3406_0,
    i_10_284_3407_0, i_10_284_3648_0, i_10_284_3682_0, i_10_284_3838_0,
    i_10_284_3848_0, i_10_284_3858_0, i_10_284_3893_0, i_10_284_3908_0,
    i_10_284_3978_0, i_10_284_3991_0, i_10_284_4051_0, i_10_284_4052_0,
    i_10_284_4116_0, i_10_284_4121_0, i_10_284_4129_0, i_10_284_4214_0,
    i_10_284_4231_0, i_10_284_4232_0, i_10_284_4270_0, i_10_284_4528_0,
    o_10_284_0_0  );
  input  i_10_284_65_0, i_10_284_178_0, i_10_284_181_0, i_10_284_220_0,
    i_10_284_280_0, i_10_284_425_0, i_10_284_434_0, i_10_284_448_0,
    i_10_284_460_0, i_10_284_796_0, i_10_284_1036_0, i_10_284_1200_0,
    i_10_284_1233_0, i_10_284_1234_0, i_10_284_1240_0, i_10_284_1242_0,
    i_10_284_1342_0, i_10_284_1359_0, i_10_284_1550_0, i_10_284_1576_0,
    i_10_284_1651_0, i_10_284_1819_0, i_10_284_1913_0, i_10_284_1945_0,
    i_10_284_1946_0, i_10_284_1949_0, i_10_284_1991_0, i_10_284_2178_0,
    i_10_284_2179_0, i_10_284_2305_0, i_10_284_2306_0, i_10_284_2324_0,
    i_10_284_2333_0, i_10_284_2354_0, i_10_284_2358_0, i_10_284_2359_0,
    i_10_284_2362_0, i_10_284_2363_0, i_10_284_2378_0, i_10_284_2381_0,
    i_10_284_2404_0, i_10_284_2451_0, i_10_284_2453_0, i_10_284_2463_0,
    i_10_284_2467_0, i_10_284_2475_0, i_10_284_2476_0, i_10_284_2503_0,
    i_10_284_2628_0, i_10_284_2634_0, i_10_284_2635_0, i_10_284_2659_0,
    i_10_284_2660_0, i_10_284_2674_0, i_10_284_2704_0, i_10_284_2709_0,
    i_10_284_2710_0, i_10_284_2711_0, i_10_284_2721_0, i_10_284_2727_0,
    i_10_284_2730_0, i_10_284_2731_0, i_10_284_2732_0, i_10_284_2828_0,
    i_10_284_2886_0, i_10_284_2916_0, i_10_284_2924_0, i_10_284_3034_0,
    i_10_284_3035_0, i_10_284_3040_0, i_10_284_3087_0, i_10_284_3088_0,
    i_10_284_3203_0, i_10_284_3268_0, i_10_284_3269_0, i_10_284_3384_0,
    i_10_284_3403_0, i_10_284_3404_0, i_10_284_3405_0, i_10_284_3406_0,
    i_10_284_3407_0, i_10_284_3648_0, i_10_284_3682_0, i_10_284_3838_0,
    i_10_284_3848_0, i_10_284_3858_0, i_10_284_3893_0, i_10_284_3908_0,
    i_10_284_3978_0, i_10_284_3991_0, i_10_284_4051_0, i_10_284_4052_0,
    i_10_284_4116_0, i_10_284_4121_0, i_10_284_4129_0, i_10_284_4214_0,
    i_10_284_4231_0, i_10_284_4232_0, i_10_284_4270_0, i_10_284_4528_0;
  output o_10_284_0_0;
  assign o_10_284_0_0 = ~((~i_10_284_434_0 & ((~i_10_284_280_0 & ~i_10_284_2178_0 & ~i_10_284_2363_0 & ~i_10_284_2451_0 & ~i_10_284_2709_0 & ~i_10_284_2886_0 & ~i_10_284_3269_0 & ~i_10_284_3404_0 & ~i_10_284_3682_0 & ~i_10_284_3908_0) | (~i_10_284_1240_0 & ~i_10_284_1342_0 & ~i_10_284_2660_0 & ~i_10_284_2674_0 & i_10_284_2709_0 & ~i_10_284_3268_0 & ~i_10_284_3838_0 & ~i_10_284_4121_0))) | (i_10_284_1234_0 & ((i_10_284_425_0 & ~i_10_284_796_0 & i_10_284_2710_0) | (i_10_284_796_0 & ~i_10_284_1342_0 & ~i_10_284_1359_0 & ~i_10_284_2306_0 & ~i_10_284_4231_0 & ~i_10_284_4232_0))) | (i_10_284_796_0 & ((~i_10_284_1550_0 & ~i_10_284_2179_0 & ~i_10_284_2305_0 & ~i_10_284_2363_0 & ~i_10_284_2463_0 & ~i_10_284_2467_0 & ~i_10_284_2886_0 & ~i_10_284_4116_0) | (~i_10_284_178_0 & ~i_10_284_2306_0 & ~i_10_284_2359_0 & ~i_10_284_2635_0 & i_10_284_3405_0 & ~i_10_284_3991_0 & ~i_10_284_4231_0))) | (~i_10_284_1550_0 & ((i_10_284_280_0 & ~i_10_284_1949_0 & ~i_10_284_2178_0 & ~i_10_284_2324_0 & ~i_10_284_2381_0 & ~i_10_284_2709_0 & ~i_10_284_2710_0 & ~i_10_284_2732_0 & ~i_10_284_2886_0 & ~i_10_284_4214_0 & ~i_10_284_4231_0) | (~i_10_284_448_0 & ~i_10_284_2628_0 & i_10_284_2828_0 & ~i_10_284_2924_0 & ~i_10_284_3088_0 & ~i_10_284_3269_0 & ~i_10_284_3405_0 & ~i_10_284_4232_0))) | (i_10_284_1819_0 & ((i_10_284_181_0 & i_10_284_3838_0) | (~i_10_284_1342_0 & ~i_10_284_1991_0 & ~i_10_284_2305_0 & ~i_10_284_2453_0 & ~i_10_284_3268_0 & ~i_10_284_3269_0 & ~i_10_284_4232_0))) | (~i_10_284_4232_0 & ((~i_10_284_425_0 & ~i_10_284_2305_0 & ~i_10_284_4214_0 & ((~i_10_284_460_0 & ~i_10_284_1240_0 & ~i_10_284_1991_0 & ~i_10_284_2358_0 & ~i_10_284_2381_0 & ~i_10_284_2634_0 & ~i_10_284_2924_0) | (~i_10_284_220_0 & ~i_10_284_1342_0 & ~i_10_284_2178_0 & ~i_10_284_2362_0 & ~i_10_284_2378_0 & ~i_10_284_2476_0 & ~i_10_284_2886_0 & ~i_10_284_3404_0))) | (~i_10_284_3682_0 & ((~i_10_284_2704_0 & ~i_10_284_3268_0 & ~i_10_284_3403_0 & i_10_284_3848_0) | (~i_10_284_1342_0 & ~i_10_284_1945_0 & ~i_10_284_2324_0 & ~i_10_284_2363_0 & ~i_10_284_2674_0 & ~i_10_284_2721_0 & ~i_10_284_2924_0 & ~i_10_284_3269_0 & ~i_10_284_3404_0 & ~i_10_284_4129_0))))) | (~i_10_284_2475_0 & ((~i_10_284_2359_0 & ((~i_10_284_425_0 & ~i_10_284_4214_0 & ((i_10_284_460_0 & ~i_10_284_2362_0 & ~i_10_284_2476_0 & ~i_10_284_2674_0 & ~i_10_284_3203_0) | (~i_10_284_1991_0 & ~i_10_284_2333_0 & ~i_10_284_2828_0 & ~i_10_284_3406_0 & ~i_10_284_3407_0 & ~i_10_284_3682_0 & ~i_10_284_4231_0))) | (~i_10_284_2324_0 & ~i_10_284_2333_0 & ~i_10_284_2362_0 & ~i_10_284_2453_0 & ~i_10_284_2660_0 & ~i_10_284_2710_0 & ~i_10_284_2924_0 & ~i_10_284_4231_0))) | (~i_10_284_1240_0 & ~i_10_284_2306_0 & ~i_10_284_2358_0 & ~i_10_284_2453_0 & ~i_10_284_2463_0 & ~i_10_284_2476_0 & ~i_10_284_2660_0 & ~i_10_284_3407_0 & ~i_10_284_3682_0 & ~i_10_284_3848_0 & ~i_10_284_3978_0 & ~i_10_284_4052_0))) | (~i_10_284_2306_0 & ((i_10_284_1240_0 & ~i_10_284_2362_0 & ~i_10_284_3407_0 & ~i_10_284_3682_0 & ~i_10_284_3978_0) | (~i_10_284_2324_0 & ~i_10_284_2358_0 & ~i_10_284_2453_0 & ~i_10_284_2659_0 & ~i_10_284_3087_0 & ~i_10_284_3403_0 & ~i_10_284_3858_0 & ~i_10_284_4270_0))) | (~i_10_284_3087_0 & ~i_10_284_3407_0 & ((i_10_284_1036_0 & ~i_10_284_2463_0 & i_10_284_3978_0) | (~i_10_284_2674_0 & ~i_10_284_3203_0 & i_10_284_3406_0 & ~i_10_284_3682_0 & i_10_284_3838_0 & ~i_10_284_4129_0 & ~i_10_284_4214_0))) | (~i_10_284_3406_0 & ((~i_10_284_3384_0 & ~i_10_284_3848_0 & i_10_284_4121_0 & i_10_284_4214_0) | (~i_10_284_1946_0 & ~i_10_284_2305_0 & ~i_10_284_2363_0 & ~i_10_284_4214_0 & ~i_10_284_4231_0 & ~i_10_284_3268_0 & ~i_10_284_4129_0))) | (i_10_284_3838_0 & ((~i_10_284_1240_0 & ~i_10_284_2451_0 & ~i_10_284_2711_0 & ~i_10_284_2924_0 & ~i_10_284_3269_0) | (i_10_284_2731_0 & ~i_10_284_3203_0 & i_10_284_4129_0))));
endmodule



// Benchmark "kernel_10_285" written by ABC on Sun Jul 19 10:25:56 2020

module kernel_10_285 ( 
    i_10_285_121_0, i_10_285_148_0, i_10_285_171_0, i_10_285_174_0,
    i_10_285_175_0, i_10_285_219_0, i_10_285_220_0, i_10_285_244_0,
    i_10_285_271_0, i_10_285_279_0, i_10_285_280_0, i_10_285_281_0,
    i_10_285_328_0, i_10_285_390_0, i_10_285_435_0, i_10_285_439_0,
    i_10_285_447_0, i_10_285_507_0, i_10_285_747_0, i_10_285_748_0,
    i_10_285_750_0, i_10_285_793_0, i_10_285_891_0, i_10_285_1000_0,
    i_10_285_1026_0, i_10_285_1027_0, i_10_285_1028_0, i_10_285_1029_0,
    i_10_285_1233_0, i_10_285_1242_0, i_10_285_1306_0, i_10_285_1307_0,
    i_10_285_1308_0, i_10_285_1309_0, i_10_285_1311_0, i_10_285_1312_0,
    i_10_285_1539_0, i_10_285_1540_0, i_10_285_1575_0, i_10_285_1576_0,
    i_10_285_1647_0, i_10_285_1648_0, i_10_285_1651_0, i_10_285_1655_0,
    i_10_285_1711_0, i_10_285_1818_0, i_10_285_1822_0, i_10_285_2196_0,
    i_10_285_2199_0, i_10_285_2202_0, i_10_285_2349_0, i_10_285_2350_0,
    i_10_285_2364_0, i_10_285_2406_0, i_10_285_2463_0, i_10_285_2466_0,
    i_10_285_2467_0, i_10_285_2468_0, i_10_285_2470_0, i_10_285_2512_0,
    i_10_285_2530_0, i_10_285_2604_0, i_10_285_2628_0, i_10_285_2629_0,
    i_10_285_2674_0, i_10_285_2710_0, i_10_285_2711_0, i_10_285_2720_0,
    i_10_285_2722_0, i_10_285_2727_0, i_10_285_2732_0, i_10_285_2829_0,
    i_10_285_2830_0, i_10_285_2981_0, i_10_285_3038_0, i_10_285_3154_0,
    i_10_285_3159_0, i_10_285_3198_0, i_10_285_3270_0, i_10_285_3271_0,
    i_10_285_3322_0, i_10_285_3408_0, i_10_285_3409_0, i_10_285_3465_0,
    i_10_285_3466_0, i_10_285_3582_0, i_10_285_3586_0, i_10_285_3785_0,
    i_10_285_3807_0, i_10_285_3808_0, i_10_285_3841_0, i_10_285_3842_0,
    i_10_285_3853_0, i_10_285_3855_0, i_10_285_3857_0, i_10_285_4113_0,
    i_10_285_4114_0, i_10_285_4119_0, i_10_285_4269_0, i_10_285_4288_0,
    o_10_285_0_0  );
  input  i_10_285_121_0, i_10_285_148_0, i_10_285_171_0, i_10_285_174_0,
    i_10_285_175_0, i_10_285_219_0, i_10_285_220_0, i_10_285_244_0,
    i_10_285_271_0, i_10_285_279_0, i_10_285_280_0, i_10_285_281_0,
    i_10_285_328_0, i_10_285_390_0, i_10_285_435_0, i_10_285_439_0,
    i_10_285_447_0, i_10_285_507_0, i_10_285_747_0, i_10_285_748_0,
    i_10_285_750_0, i_10_285_793_0, i_10_285_891_0, i_10_285_1000_0,
    i_10_285_1026_0, i_10_285_1027_0, i_10_285_1028_0, i_10_285_1029_0,
    i_10_285_1233_0, i_10_285_1242_0, i_10_285_1306_0, i_10_285_1307_0,
    i_10_285_1308_0, i_10_285_1309_0, i_10_285_1311_0, i_10_285_1312_0,
    i_10_285_1539_0, i_10_285_1540_0, i_10_285_1575_0, i_10_285_1576_0,
    i_10_285_1647_0, i_10_285_1648_0, i_10_285_1651_0, i_10_285_1655_0,
    i_10_285_1711_0, i_10_285_1818_0, i_10_285_1822_0, i_10_285_2196_0,
    i_10_285_2199_0, i_10_285_2202_0, i_10_285_2349_0, i_10_285_2350_0,
    i_10_285_2364_0, i_10_285_2406_0, i_10_285_2463_0, i_10_285_2466_0,
    i_10_285_2467_0, i_10_285_2468_0, i_10_285_2470_0, i_10_285_2512_0,
    i_10_285_2530_0, i_10_285_2604_0, i_10_285_2628_0, i_10_285_2629_0,
    i_10_285_2674_0, i_10_285_2710_0, i_10_285_2711_0, i_10_285_2720_0,
    i_10_285_2722_0, i_10_285_2727_0, i_10_285_2732_0, i_10_285_2829_0,
    i_10_285_2830_0, i_10_285_2981_0, i_10_285_3038_0, i_10_285_3154_0,
    i_10_285_3159_0, i_10_285_3198_0, i_10_285_3270_0, i_10_285_3271_0,
    i_10_285_3322_0, i_10_285_3408_0, i_10_285_3409_0, i_10_285_3465_0,
    i_10_285_3466_0, i_10_285_3582_0, i_10_285_3586_0, i_10_285_3785_0,
    i_10_285_3807_0, i_10_285_3808_0, i_10_285_3841_0, i_10_285_3842_0,
    i_10_285_3853_0, i_10_285_3855_0, i_10_285_3857_0, i_10_285_4113_0,
    i_10_285_4114_0, i_10_285_4119_0, i_10_285_4269_0, i_10_285_4288_0;
  output o_10_285_0_0;
  assign o_10_285_0_0 = ~((i_10_285_148_0 & ((~i_10_285_1026_0 & ~i_10_285_3785_0) | (~i_10_285_1029_0 & i_10_285_1822_0 & ~i_10_285_2628_0 & ~i_10_285_3586_0 & ~i_10_285_3842_0))) | (~i_10_285_175_0 & ((~i_10_285_1309_0 & ~i_10_285_2199_0 & i_10_285_3271_0 & ~i_10_285_3785_0 & ~i_10_285_3855_0) | (~i_10_285_148_0 & ~i_10_285_1648_0 & ~i_10_285_2830_0 & ~i_10_285_3270_0 & ~i_10_285_3408_0 & ~i_10_285_3842_0 & i_10_285_4119_0))) | (~i_10_285_2199_0 & ((~i_10_285_220_0 & ((~i_10_285_390_0 & ~i_10_285_1306_0 & ~i_10_285_1311_0 & ~i_10_285_1540_0 & ~i_10_285_1647_0 & ~i_10_285_2406_0 & ~i_10_285_2722_0 & ~i_10_285_2829_0 & ~i_10_285_3853_0) | (~i_10_285_174_0 & ~i_10_285_2364_0 & ~i_10_285_2720_0 & ~i_10_285_3159_0 & ~i_10_285_3198_0 & ~i_10_285_3270_0 & ~i_10_285_3409_0 & ~i_10_285_3842_0 & ~i_10_285_3855_0))) | (~i_10_285_2406_0 & ((~i_10_285_435_0 & ~i_10_285_3409_0 & ((i_10_285_439_0 & ~i_10_285_1647_0 & i_10_285_1822_0 & ~i_10_285_2829_0) | (~i_10_285_1307_0 & ~i_10_285_2364_0 & ~i_10_285_3198_0 & ~i_10_285_3586_0 & ~i_10_285_3857_0 & ~i_10_285_4113_0))) | (~i_10_285_1027_0 & ~i_10_285_1242_0 & ~i_10_285_1311_0 & ~i_10_285_1651_0 & ~i_10_285_3198_0 & ~i_10_285_3785_0 & i_10_285_3857_0 & ~i_10_285_4119_0))) | (~i_10_285_748_0 & ((~i_10_285_439_0 & ~i_10_285_3198_0 & ((~i_10_285_328_0 & ~i_10_285_891_0 & ~i_10_285_1026_0 & ~i_10_285_1311_0 & ~i_10_285_2350_0 & ~i_10_285_3408_0) | (~i_10_285_1822_0 & ~i_10_285_2829_0 & ~i_10_285_3271_0 & ~i_10_285_4113_0))) | (i_10_285_281_0 & ~i_10_285_1539_0 & ~i_10_285_3408_0))) | (~i_10_285_3842_0 & ~i_10_285_3855_0 & i_10_285_3038_0 & ~i_10_285_3198_0) | (i_10_285_2470_0 & i_10_285_2829_0 & ~i_10_285_3270_0 & i_10_285_3855_0 & i_10_285_3857_0))) | (i_10_285_279_0 & ((~i_10_285_244_0 & ~i_10_285_390_0 & ~i_10_285_747_0 & ~i_10_285_1029_0 & ~i_10_285_1647_0 & ~i_10_285_3842_0) | (i_10_285_793_0 & ~i_10_285_2463_0 & i_10_285_3841_0 & i_10_285_3853_0))) | (i_10_285_793_0 & ((~i_10_285_439_0 & ~i_10_285_447_0 & ~i_10_285_747_0 & ~i_10_285_1028_0 & ~i_10_285_1540_0 & ~i_10_285_2202_0 & ~i_10_285_2463_0) | (~i_10_285_1648_0 & ~i_10_285_2829_0 & ~i_10_285_2981_0 & ~i_10_285_3841_0 & ~i_10_285_4114_0))) | (~i_10_285_1311_0 & ((~i_10_285_748_0 & ~i_10_285_3409_0 & ((~i_10_285_1242_0 & ~i_10_285_1307_0 & ~i_10_285_2196_0 & ~i_10_285_2364_0 & ~i_10_285_2406_0 & i_10_285_2830_0 & ~i_10_285_3038_0 & ~i_10_285_3408_0) | (~i_10_285_121_0 & ~i_10_285_747_0 & ~i_10_285_750_0 & ~i_10_285_1028_0 & ~i_10_285_1312_0 & ~i_10_285_2829_0 & ~i_10_285_3198_0 & ~i_10_285_3855_0))) | (~i_10_285_279_0 & ~i_10_285_328_0 & ~i_10_285_439_0 & ~i_10_285_1575_0 & ~i_10_285_2202_0 & ~i_10_285_2629_0 & ~i_10_285_3270_0 & ~i_10_285_3271_0) | (~i_10_285_1028_0 & ~i_10_285_1308_0 & ~i_10_285_3408_0 & i_10_285_3857_0 & ~i_10_285_4113_0))) | (~i_10_285_3198_0 & ((~i_10_285_328_0 & ((~i_10_285_2350_0 & i_10_285_2467_0 & ~i_10_285_2711_0 & ~i_10_285_3409_0) | (~i_10_285_219_0 & ~i_10_285_439_0 & ~i_10_285_748_0 & i_10_285_3857_0 & ~i_10_285_4113_0 & ~i_10_285_793_0 & ~i_10_285_1312_0))) | (~i_10_285_1309_0 & i_10_285_1822_0 & i_10_285_2830_0) | (i_10_285_2710_0 & ~i_10_285_2829_0 & ~i_10_285_3582_0) | (i_10_285_175_0 & ~i_10_285_2604_0 & ~i_10_285_2732_0 & ~i_10_285_3842_0 & ~i_10_285_4113_0))) | (~i_10_285_747_0 & ((~i_10_285_219_0 & ~i_10_285_435_0 & ~i_10_285_1308_0 & ~i_10_285_1309_0 & ~i_10_285_1312_0 & ~i_10_285_2364_0 & ~i_10_285_2629_0) | (~i_10_285_244_0 & ~i_10_285_439_0 & ~i_10_285_1029_0 & ~i_10_285_1648_0 & ~i_10_285_1655_0 & ~i_10_285_2829_0 & ~i_10_285_3270_0 & ~i_10_285_3841_0 & ~i_10_285_3842_0))) | (~i_10_285_219_0 & ((~i_10_285_244_0 & i_10_285_1655_0 & ~i_10_285_2202_0 & i_10_285_3038_0) | (~i_10_285_171_0 & i_10_285_280_0 & ~i_10_285_390_0 & ~i_10_285_748_0 & ~i_10_285_1026_0 & ~i_10_285_2727_0 & ~i_10_285_3841_0))) | (~i_10_285_4113_0 & ((~i_10_285_439_0 & ~i_10_285_4114_0 & ((~i_10_285_1026_0 & ~i_10_285_1312_0 & ~i_10_285_2830_0 & ~i_10_285_3270_0 & ~i_10_285_3842_0) | (~i_10_285_1308_0 & ~i_10_285_2364_0 & ~i_10_285_3855_0 & ~i_10_285_4269_0))) | i_10_285_2468_0 | (i_10_285_174_0 & ~i_10_285_2202_0 & ~i_10_285_3409_0 & ~i_10_285_3855_0))) | (~i_10_285_1026_0 & ((~i_10_285_2406_0 & i_10_285_2470_0 & ~i_10_285_2732_0 & ~i_10_285_3785_0) | (~i_10_285_1309_0 & ~i_10_285_1575_0 & ~i_10_285_2364_0 & ~i_10_285_2463_0 & ~i_10_285_2720_0 & ~i_10_285_3270_0 & ~i_10_285_3841_0))) | (i_10_285_3586_0 & ((i_10_285_2364_0 & (~i_10_285_1309_0 | (i_10_285_2199_0 & i_10_285_2732_0) | (~i_10_285_2406_0 & i_10_285_4119_0))) | (~i_10_285_1539_0 & i_10_285_2467_0 & ~i_10_285_2830_0))) | (~i_10_285_244_0 & ~i_10_285_1575_0 & ~i_10_285_1647_0 & i_10_285_1818_0 & ~i_10_285_3785_0) | (~i_10_285_2364_0 & i_10_285_2711_0 & i_10_285_3409_0 & ~i_10_285_3841_0));
endmodule



// Benchmark "kernel_10_286" written by ABC on Sun Jul 19 10:25:57 2020

module kernel_10_286 ( 
    i_10_286_208_0, i_10_286_209_0, i_10_286_218_0, i_10_286_270_0,
    i_10_286_271_0, i_10_286_272_0, i_10_286_281_0, i_10_286_283_0,
    i_10_286_407_0, i_10_286_424_0, i_10_286_425_0, i_10_286_433_0,
    i_10_286_437_0, i_10_286_445_0, i_10_286_465_0, i_10_286_508_0,
    i_10_286_902_0, i_10_286_986_0, i_10_286_1036_0, i_10_286_1117_0,
    i_10_286_1118_0, i_10_286_1217_0, i_10_286_1235_0, i_10_286_1243_0,
    i_10_286_1244_0, i_10_286_1361_0, i_10_286_1444_0, i_10_286_1445_0,
    i_10_286_1822_0, i_10_286_1823_0, i_10_286_1882_0, i_10_286_1883_0,
    i_10_286_1990_0, i_10_286_2089_0, i_10_286_2323_0, i_10_286_2327_0,
    i_10_286_2333_0, i_10_286_2351_0, i_10_286_2368_0, i_10_286_2369_0,
    i_10_286_2432_0, i_10_286_2441_0, i_10_286_2462_0, i_10_286_2606_0,
    i_10_286_2630_0, i_10_286_2634_0, i_10_286_2639_0, i_10_286_2674_0,
    i_10_286_2675_0, i_10_286_2701_0, i_10_286_2702_0, i_10_286_2705_0,
    i_10_286_2728_0, i_10_286_2819_0, i_10_286_2831_0, i_10_286_2863_0,
    i_10_286_2864_0, i_10_286_2917_0, i_10_286_2920_0, i_10_286_2921_0,
    i_10_286_3034_0, i_10_286_3224_0, i_10_286_3281_0, i_10_286_3298_0,
    i_10_286_3349_0, i_10_286_3406_0, i_10_286_3466_0, i_10_286_3647_0,
    i_10_286_3682_0, i_10_286_3782_0, i_10_286_3785_0, i_10_286_3847_0,
    i_10_286_3848_0, i_10_286_3849_0, i_10_286_3857_0, i_10_286_3889_0,
    i_10_286_3890_0, i_10_286_3893_0, i_10_286_3980_0, i_10_286_4028_0,
    i_10_286_4118_0, i_10_286_4142_0, i_10_286_4185_0, i_10_286_4186_0,
    i_10_286_4187_0, i_10_286_4276_0, i_10_286_4277_0, i_10_286_4285_0,
    i_10_286_4286_0, i_10_286_4288_0, i_10_286_4289_0, i_10_286_4290_0,
    i_10_286_4291_0, i_10_286_4510_0, i_10_286_4511_0, i_10_286_4563_0,
    i_10_286_4564_0, i_10_286_4571_0, i_10_286_4583_0, i_10_286_4601_0,
    o_10_286_0_0  );
  input  i_10_286_208_0, i_10_286_209_0, i_10_286_218_0, i_10_286_270_0,
    i_10_286_271_0, i_10_286_272_0, i_10_286_281_0, i_10_286_283_0,
    i_10_286_407_0, i_10_286_424_0, i_10_286_425_0, i_10_286_433_0,
    i_10_286_437_0, i_10_286_445_0, i_10_286_465_0, i_10_286_508_0,
    i_10_286_902_0, i_10_286_986_0, i_10_286_1036_0, i_10_286_1117_0,
    i_10_286_1118_0, i_10_286_1217_0, i_10_286_1235_0, i_10_286_1243_0,
    i_10_286_1244_0, i_10_286_1361_0, i_10_286_1444_0, i_10_286_1445_0,
    i_10_286_1822_0, i_10_286_1823_0, i_10_286_1882_0, i_10_286_1883_0,
    i_10_286_1990_0, i_10_286_2089_0, i_10_286_2323_0, i_10_286_2327_0,
    i_10_286_2333_0, i_10_286_2351_0, i_10_286_2368_0, i_10_286_2369_0,
    i_10_286_2432_0, i_10_286_2441_0, i_10_286_2462_0, i_10_286_2606_0,
    i_10_286_2630_0, i_10_286_2634_0, i_10_286_2639_0, i_10_286_2674_0,
    i_10_286_2675_0, i_10_286_2701_0, i_10_286_2702_0, i_10_286_2705_0,
    i_10_286_2728_0, i_10_286_2819_0, i_10_286_2831_0, i_10_286_2863_0,
    i_10_286_2864_0, i_10_286_2917_0, i_10_286_2920_0, i_10_286_2921_0,
    i_10_286_3034_0, i_10_286_3224_0, i_10_286_3281_0, i_10_286_3298_0,
    i_10_286_3349_0, i_10_286_3406_0, i_10_286_3466_0, i_10_286_3647_0,
    i_10_286_3682_0, i_10_286_3782_0, i_10_286_3785_0, i_10_286_3847_0,
    i_10_286_3848_0, i_10_286_3849_0, i_10_286_3857_0, i_10_286_3889_0,
    i_10_286_3890_0, i_10_286_3893_0, i_10_286_3980_0, i_10_286_4028_0,
    i_10_286_4118_0, i_10_286_4142_0, i_10_286_4185_0, i_10_286_4186_0,
    i_10_286_4187_0, i_10_286_4276_0, i_10_286_4277_0, i_10_286_4285_0,
    i_10_286_4286_0, i_10_286_4288_0, i_10_286_4289_0, i_10_286_4290_0,
    i_10_286_4291_0, i_10_286_4510_0, i_10_286_4511_0, i_10_286_4563_0,
    i_10_286_4564_0, i_10_286_4571_0, i_10_286_4583_0, i_10_286_4601_0;
  output o_10_286_0_0;
  assign o_10_286_0_0 = 0;
endmodule



// Benchmark "kernel_10_287" written by ABC on Sun Jul 19 10:25:58 2020

module kernel_10_287 ( 
    i_10_287_34_0, i_10_287_89_0, i_10_287_174_0, i_10_287_175_0,
    i_10_287_176_0, i_10_287_177_0, i_10_287_178_0, i_10_287_249_0,
    i_10_287_267_0, i_10_287_277_0, i_10_287_283_0, i_10_287_284_0,
    i_10_287_412_0, i_10_287_440_0, i_10_287_509_0, i_10_287_796_0,
    i_10_287_898_0, i_10_287_963_0, i_10_287_1033_0, i_10_287_1034_0,
    i_10_287_1165_0, i_10_287_1237_0, i_10_287_1311_0, i_10_287_1362_0,
    i_10_287_1440_0, i_10_287_1491_0, i_10_287_1549_0, i_10_287_1550_0,
    i_10_287_1651_0, i_10_287_1654_0, i_10_287_1655_0, i_10_287_1821_0,
    i_10_287_1822_0, i_10_287_1823_0, i_10_287_2026_0, i_10_287_2334_0,
    i_10_287_2350_0, i_10_287_2351_0, i_10_287_2353_0, i_10_287_2354_0,
    i_10_287_2407_0, i_10_287_2408_0, i_10_287_2449_0, i_10_287_2452_0,
    i_10_287_2453_0, i_10_287_2465_0, i_10_287_2608_0, i_10_287_2609_0,
    i_10_287_2631_0, i_10_287_2635_0, i_10_287_2636_0, i_10_287_2644_0,
    i_10_287_2678_0, i_10_287_2725_0, i_10_287_2733_0, i_10_287_2735_0,
    i_10_287_2829_0, i_10_287_2919_0, i_10_287_3076_0, i_10_287_3154_0,
    i_10_287_3155_0, i_10_287_3156_0, i_10_287_3162_0, i_10_287_3165_0,
    i_10_287_3166_0, i_10_287_3167_0, i_10_287_3201_0, i_10_287_3237_0,
    i_10_287_3279_0, i_10_287_3280_0, i_10_287_3282_0, i_10_287_3385_0,
    i_10_287_3386_0, i_10_287_3388_0, i_10_287_3389_0, i_10_287_3390_0,
    i_10_287_3525_0, i_10_287_3586_0, i_10_287_3587_0, i_10_287_3613_0,
    i_10_287_3614_0, i_10_287_3853_0, i_10_287_3855_0, i_10_287_3891_0,
    i_10_287_3912_0, i_10_287_3991_0, i_10_287_4113_0, i_10_287_4117_0,
    i_10_287_4118_0, i_10_287_4119_0, i_10_287_4121_0, i_10_287_4125_0,
    i_10_287_4126_0, i_10_287_4128_0, i_10_287_4129_0, i_10_287_4130_0,
    i_10_287_4174_0, i_10_287_4219_0, i_10_287_4272_0, i_10_287_4292_0,
    o_10_287_0_0  );
  input  i_10_287_34_0, i_10_287_89_0, i_10_287_174_0, i_10_287_175_0,
    i_10_287_176_0, i_10_287_177_0, i_10_287_178_0, i_10_287_249_0,
    i_10_287_267_0, i_10_287_277_0, i_10_287_283_0, i_10_287_284_0,
    i_10_287_412_0, i_10_287_440_0, i_10_287_509_0, i_10_287_796_0,
    i_10_287_898_0, i_10_287_963_0, i_10_287_1033_0, i_10_287_1034_0,
    i_10_287_1165_0, i_10_287_1237_0, i_10_287_1311_0, i_10_287_1362_0,
    i_10_287_1440_0, i_10_287_1491_0, i_10_287_1549_0, i_10_287_1550_0,
    i_10_287_1651_0, i_10_287_1654_0, i_10_287_1655_0, i_10_287_1821_0,
    i_10_287_1822_0, i_10_287_1823_0, i_10_287_2026_0, i_10_287_2334_0,
    i_10_287_2350_0, i_10_287_2351_0, i_10_287_2353_0, i_10_287_2354_0,
    i_10_287_2407_0, i_10_287_2408_0, i_10_287_2449_0, i_10_287_2452_0,
    i_10_287_2453_0, i_10_287_2465_0, i_10_287_2608_0, i_10_287_2609_0,
    i_10_287_2631_0, i_10_287_2635_0, i_10_287_2636_0, i_10_287_2644_0,
    i_10_287_2678_0, i_10_287_2725_0, i_10_287_2733_0, i_10_287_2735_0,
    i_10_287_2829_0, i_10_287_2919_0, i_10_287_3076_0, i_10_287_3154_0,
    i_10_287_3155_0, i_10_287_3156_0, i_10_287_3162_0, i_10_287_3165_0,
    i_10_287_3166_0, i_10_287_3167_0, i_10_287_3201_0, i_10_287_3237_0,
    i_10_287_3279_0, i_10_287_3280_0, i_10_287_3282_0, i_10_287_3385_0,
    i_10_287_3386_0, i_10_287_3388_0, i_10_287_3389_0, i_10_287_3390_0,
    i_10_287_3525_0, i_10_287_3586_0, i_10_287_3587_0, i_10_287_3613_0,
    i_10_287_3614_0, i_10_287_3853_0, i_10_287_3855_0, i_10_287_3891_0,
    i_10_287_3912_0, i_10_287_3991_0, i_10_287_4113_0, i_10_287_4117_0,
    i_10_287_4118_0, i_10_287_4119_0, i_10_287_4121_0, i_10_287_4125_0,
    i_10_287_4126_0, i_10_287_4128_0, i_10_287_4129_0, i_10_287_4130_0,
    i_10_287_4174_0, i_10_287_4219_0, i_10_287_4272_0, i_10_287_4292_0;
  output o_10_287_0_0;
  assign o_10_287_0_0 = ~((~i_10_287_174_0 & ((~i_10_287_440_0 & ~i_10_287_1165_0 & ~i_10_287_2449_0 & ~i_10_287_2644_0 & ~i_10_287_2733_0 & ~i_10_287_3167_0) | (~i_10_287_1651_0 & ~i_10_287_2351_0 & ~i_10_287_2465_0 & ~i_10_287_3386_0 & ~i_10_287_3525_0 & ~i_10_287_3614_0 & ~i_10_287_4130_0))) | (~i_10_287_1655_0 & ((i_10_287_178_0 & ((~i_10_287_2350_0 & ~i_10_287_2353_0 & i_10_287_3237_0 & ~i_10_287_4118_0) | (~i_10_287_3279_0 & ~i_10_287_3853_0 & ~i_10_287_3891_0 & ~i_10_287_4121_0 & ~i_10_287_4129_0 & ~i_10_287_4272_0))) | (~i_10_287_1237_0 & ~i_10_287_1651_0 & ~i_10_287_1821_0 & ~i_10_287_2354_0 & i_10_287_4117_0))) | (~i_10_287_178_0 & ((i_10_287_2353_0 & i_10_287_3282_0) | (~i_10_287_89_0 & ~i_10_287_249_0 & ~i_10_287_440_0 & ~i_10_287_1033_0 & ~i_10_287_1034_0 & ~i_10_287_1165_0 & ~i_10_287_4128_0))) | (i_10_287_283_0 & ((~i_10_287_1237_0 & ~i_10_287_2919_0 & ~i_10_287_3282_0) | (~i_10_287_89_0 & ~i_10_287_2635_0 & ~i_10_287_4117_0))) | (~i_10_287_4292_0 & ((~i_10_287_898_0 & ~i_10_287_1440_0 & ((~i_10_287_89_0 & ~i_10_287_2026_0 & ~i_10_287_2919_0 & ~i_10_287_3279_0 & ~i_10_287_3912_0 & ~i_10_287_3991_0) | (~i_10_287_1491_0 & i_10_287_1651_0 & ~i_10_287_2449_0 & ~i_10_287_3165_0 & ~i_10_287_4121_0 & ~i_10_287_4130_0))) | (~i_10_287_1362_0 & ~i_10_287_2635_0 & ~i_10_287_2733_0 & i_10_287_3388_0) | (i_10_287_175_0 & i_10_287_796_0 & ~i_10_287_1491_0 & ~i_10_287_3237_0 & ~i_10_287_3385_0 & i_10_287_4117_0 & ~i_10_287_4130_0 & ~i_10_287_4272_0))) | (~i_10_287_1033_0 & ((i_10_287_1237_0 & i_10_287_1823_0 & i_10_287_2452_0 & ~i_10_287_3853_0 & ~i_10_287_3891_0 & ~i_10_287_2678_0 & ~i_10_287_2829_0) | (~i_10_287_249_0 & ~i_10_287_1165_0 & ~i_10_287_2452_0 & ~i_10_287_2644_0 & ~i_10_287_3166_0 & ~i_10_287_3991_0))) | (~i_10_287_249_0 & ((~i_10_287_89_0 & ~i_10_287_284_0 & ~i_10_287_796_0 & ~i_10_287_2465_0 & ~i_10_287_2678_0 & ~i_10_287_3165_0 & ~i_10_287_3201_0 & ~i_10_287_3855_0 & ~i_10_287_4174_0) | (~i_10_287_963_0 & ~i_10_287_2351_0 & ~i_10_287_2608_0 & i_10_287_2631_0 & ~i_10_287_2735_0 & ~i_10_287_2919_0 & i_10_287_4117_0 & ~i_10_287_4272_0))) | (~i_10_287_3167_0 & ((~i_10_287_89_0 & ((~i_10_287_1165_0 & ~i_10_287_1491_0 & ~i_10_287_2609_0 & ((~i_10_287_176_0 & ~i_10_287_3162_0 & ~i_10_287_3165_0 & ~i_10_287_3525_0) | (~i_10_287_1440_0 & ~i_10_287_2449_0 & ~i_10_287_3237_0 & ~i_10_287_3280_0 & ~i_10_287_4128_0))) | (~i_10_287_175_0 & ~i_10_287_1654_0 & ~i_10_287_2644_0 & ~i_10_287_3613_0 & ~i_10_287_4219_0))) | (~i_10_287_1311_0 & ~i_10_287_2408_0 & i_10_287_2452_0 & ~i_10_287_2733_0 & ~i_10_287_3165_0 & ~i_10_287_3891_0 & ~i_10_287_4119_0 & ~i_10_287_4121_0 & ~i_10_287_4219_0))) | (~i_10_287_176_0 & ((i_10_287_2407_0 & ~i_10_287_2919_0 & ~i_10_287_3165_0 & ~i_10_287_3280_0) | (~i_10_287_440_0 & ~i_10_287_1362_0 & i_10_287_2635_0 & ~i_10_287_3237_0 & ~i_10_287_3891_0 & ~i_10_287_3991_0 & ~i_10_287_4121_0 & ~i_10_287_4128_0 & ~i_10_287_4129_0))) | (i_10_287_284_0 & ~i_10_287_2644_0 & ~i_10_287_2919_0 & ~i_10_287_4121_0) | (i_10_287_2354_0 & ~i_10_287_2453_0 & ~i_10_287_2636_0 & ~i_10_287_3162_0) | (~i_10_287_1362_0 & i_10_287_2350_0 & ~i_10_287_2725_0 & ~i_10_287_3912_0 & ~i_10_287_4126_0));
endmodule



// Benchmark "kernel_10_288" written by ABC on Sun Jul 19 10:25:59 2020

module kernel_10_288 ( 
    i_10_288_48_0, i_10_288_63_0, i_10_288_81_0, i_10_288_117_0,
    i_10_288_174_0, i_10_288_178_0, i_10_288_219_0, i_10_288_220_0,
    i_10_288_222_0, i_10_288_223_0, i_10_288_224_0, i_10_288_261_0,
    i_10_288_285_0, i_10_288_286_0, i_10_288_367_0, i_10_288_406_0,
    i_10_288_427_0, i_10_288_439_0, i_10_288_531_0, i_10_288_534_0,
    i_10_288_736_0, i_10_288_901_0, i_10_288_957_0, i_10_288_999_0,
    i_10_288_1041_0, i_10_288_1156_0, i_10_288_1233_0, i_10_288_1236_0,
    i_10_288_1296_0, i_10_288_1310_0, i_10_288_1341_0, i_10_288_1359_0,
    i_10_288_1440_0, i_10_288_1441_0, i_10_288_1476_0, i_10_288_1540_0,
    i_10_288_1614_0, i_10_288_1653_0, i_10_288_1655_0, i_10_288_1711_0,
    i_10_288_1719_0, i_10_288_1764_0, i_10_288_1765_0, i_10_288_1821_0,
    i_10_288_1890_0, i_10_288_1909_0, i_10_288_1912_0, i_10_288_1916_0,
    i_10_288_1945_0, i_10_288_2019_0, i_10_288_2109_0, i_10_288_2160_0,
    i_10_288_2178_0, i_10_288_2236_0, i_10_288_2254_0, i_10_288_2350_0,
    i_10_288_2361_0, i_10_288_2377_0, i_10_288_2466_0, i_10_288_2469_0,
    i_10_288_2515_0, i_10_288_2541_0, i_10_288_2655_0, i_10_288_2676_0,
    i_10_288_2704_0, i_10_288_2709_0, i_10_288_2742_0, i_10_288_2844_0,
    i_10_288_2923_0, i_10_288_3033_0, i_10_288_3040_0, i_10_288_3095_0,
    i_10_288_3114_0, i_10_288_3231_0, i_10_288_3270_0, i_10_288_3277_0,
    i_10_288_3289_0, i_10_288_3331_0, i_10_288_3434_0, i_10_288_3465_0,
    i_10_288_3492_0, i_10_288_3523_0, i_10_288_3526_0, i_10_288_3538_0,
    i_10_288_3561_0, i_10_288_3582_0, i_10_288_3837_0, i_10_288_3852_0,
    i_10_288_3853_0, i_10_288_3859_0, i_10_288_3901_0, i_10_288_4114_0,
    i_10_288_4161_0, i_10_288_4218_0, i_10_288_4219_0, i_10_288_4222_0,
    i_10_288_4234_0, i_10_288_4311_0, i_10_288_4554_0, i_10_288_4580_0,
    o_10_288_0_0  );
  input  i_10_288_48_0, i_10_288_63_0, i_10_288_81_0, i_10_288_117_0,
    i_10_288_174_0, i_10_288_178_0, i_10_288_219_0, i_10_288_220_0,
    i_10_288_222_0, i_10_288_223_0, i_10_288_224_0, i_10_288_261_0,
    i_10_288_285_0, i_10_288_286_0, i_10_288_367_0, i_10_288_406_0,
    i_10_288_427_0, i_10_288_439_0, i_10_288_531_0, i_10_288_534_0,
    i_10_288_736_0, i_10_288_901_0, i_10_288_957_0, i_10_288_999_0,
    i_10_288_1041_0, i_10_288_1156_0, i_10_288_1233_0, i_10_288_1236_0,
    i_10_288_1296_0, i_10_288_1310_0, i_10_288_1341_0, i_10_288_1359_0,
    i_10_288_1440_0, i_10_288_1441_0, i_10_288_1476_0, i_10_288_1540_0,
    i_10_288_1614_0, i_10_288_1653_0, i_10_288_1655_0, i_10_288_1711_0,
    i_10_288_1719_0, i_10_288_1764_0, i_10_288_1765_0, i_10_288_1821_0,
    i_10_288_1890_0, i_10_288_1909_0, i_10_288_1912_0, i_10_288_1916_0,
    i_10_288_1945_0, i_10_288_2019_0, i_10_288_2109_0, i_10_288_2160_0,
    i_10_288_2178_0, i_10_288_2236_0, i_10_288_2254_0, i_10_288_2350_0,
    i_10_288_2361_0, i_10_288_2377_0, i_10_288_2466_0, i_10_288_2469_0,
    i_10_288_2515_0, i_10_288_2541_0, i_10_288_2655_0, i_10_288_2676_0,
    i_10_288_2704_0, i_10_288_2709_0, i_10_288_2742_0, i_10_288_2844_0,
    i_10_288_2923_0, i_10_288_3033_0, i_10_288_3040_0, i_10_288_3095_0,
    i_10_288_3114_0, i_10_288_3231_0, i_10_288_3270_0, i_10_288_3277_0,
    i_10_288_3289_0, i_10_288_3331_0, i_10_288_3434_0, i_10_288_3465_0,
    i_10_288_3492_0, i_10_288_3523_0, i_10_288_3526_0, i_10_288_3538_0,
    i_10_288_3561_0, i_10_288_3582_0, i_10_288_3837_0, i_10_288_3852_0,
    i_10_288_3853_0, i_10_288_3859_0, i_10_288_3901_0, i_10_288_4114_0,
    i_10_288_4161_0, i_10_288_4218_0, i_10_288_4219_0, i_10_288_4222_0,
    i_10_288_4234_0, i_10_288_4311_0, i_10_288_4554_0, i_10_288_4580_0;
  output o_10_288_0_0;
  assign o_10_288_0_0 = 0;
endmodule



// Benchmark "kernel_10_289" written by ABC on Sun Jul 19 10:26:01 2020

module kernel_10_289 ( 
    i_10_289_124_0, i_10_289_125_0, i_10_289_174_0, i_10_289_177_0,
    i_10_289_183_0, i_10_289_184_0, i_10_289_280_0, i_10_289_285_0,
    i_10_289_286_0, i_10_289_287_0, i_10_289_317_0, i_10_289_318_0,
    i_10_289_319_0, i_10_289_446_0, i_10_289_449_0, i_10_289_460_0,
    i_10_289_462_0, i_10_289_463_0, i_10_289_464_0, i_10_289_510_0,
    i_10_289_511_0, i_10_289_514_0, i_10_289_749_0, i_10_289_955_0,
    i_10_289_993_0, i_10_289_1006_0, i_10_289_1034_0, i_10_289_1037_0,
    i_10_289_1244_0, i_10_289_1247_0, i_10_289_1308_0, i_10_289_1310_0,
    i_10_289_1363_0, i_10_289_1380_0, i_10_289_1552_0, i_10_289_1653_0,
    i_10_289_1685_0, i_10_289_1819_0, i_10_289_1820_0, i_10_289_1822_0,
    i_10_289_1823_0, i_10_289_1825_0, i_10_289_1826_0, i_10_289_1950_0,
    i_10_289_1995_0, i_10_289_2095_0, i_10_289_2351_0, i_10_289_2354_0,
    i_10_289_2356_0, i_10_289_2361_0, i_10_289_2362_0, i_10_289_2455_0,
    i_10_289_2469_0, i_10_289_2632_0, i_10_289_2702_0, i_10_289_2713_0,
    i_10_289_2715_0, i_10_289_2722_0, i_10_289_2724_0, i_10_289_2725_0,
    i_10_289_2731_0, i_10_289_2734_0, i_10_289_2829_0, i_10_289_2830_0,
    i_10_289_2834_0, i_10_289_2920_0, i_10_289_3040_0, i_10_289_3041_0,
    i_10_289_3151_0, i_10_289_3195_0, i_10_289_3196_0, i_10_289_3197_0,
    i_10_289_3198_0, i_10_289_3199_0, i_10_289_3270_0, i_10_289_3271_0,
    i_10_289_3328_0, i_10_289_3387_0, i_10_289_3388_0, i_10_289_3389_0,
    i_10_289_3391_0, i_10_289_3392_0, i_10_289_3610_0, i_10_289_3613_0,
    i_10_289_3647_0, i_10_289_3649_0, i_10_289_3653_0, i_10_289_3780_0,
    i_10_289_3781_0, i_10_289_3782_0, i_10_289_3837_0, i_10_289_3838_0,
    i_10_289_3839_0, i_10_289_3842_0, i_10_289_3856_0, i_10_289_3967_0,
    i_10_289_3985_0, i_10_289_4114_0, i_10_289_4291_0, i_10_289_4427_0,
    o_10_289_0_0  );
  input  i_10_289_124_0, i_10_289_125_0, i_10_289_174_0, i_10_289_177_0,
    i_10_289_183_0, i_10_289_184_0, i_10_289_280_0, i_10_289_285_0,
    i_10_289_286_0, i_10_289_287_0, i_10_289_317_0, i_10_289_318_0,
    i_10_289_319_0, i_10_289_446_0, i_10_289_449_0, i_10_289_460_0,
    i_10_289_462_0, i_10_289_463_0, i_10_289_464_0, i_10_289_510_0,
    i_10_289_511_0, i_10_289_514_0, i_10_289_749_0, i_10_289_955_0,
    i_10_289_993_0, i_10_289_1006_0, i_10_289_1034_0, i_10_289_1037_0,
    i_10_289_1244_0, i_10_289_1247_0, i_10_289_1308_0, i_10_289_1310_0,
    i_10_289_1363_0, i_10_289_1380_0, i_10_289_1552_0, i_10_289_1653_0,
    i_10_289_1685_0, i_10_289_1819_0, i_10_289_1820_0, i_10_289_1822_0,
    i_10_289_1823_0, i_10_289_1825_0, i_10_289_1826_0, i_10_289_1950_0,
    i_10_289_1995_0, i_10_289_2095_0, i_10_289_2351_0, i_10_289_2354_0,
    i_10_289_2356_0, i_10_289_2361_0, i_10_289_2362_0, i_10_289_2455_0,
    i_10_289_2469_0, i_10_289_2632_0, i_10_289_2702_0, i_10_289_2713_0,
    i_10_289_2715_0, i_10_289_2722_0, i_10_289_2724_0, i_10_289_2725_0,
    i_10_289_2731_0, i_10_289_2734_0, i_10_289_2829_0, i_10_289_2830_0,
    i_10_289_2834_0, i_10_289_2920_0, i_10_289_3040_0, i_10_289_3041_0,
    i_10_289_3151_0, i_10_289_3195_0, i_10_289_3196_0, i_10_289_3197_0,
    i_10_289_3198_0, i_10_289_3199_0, i_10_289_3270_0, i_10_289_3271_0,
    i_10_289_3328_0, i_10_289_3387_0, i_10_289_3388_0, i_10_289_3389_0,
    i_10_289_3391_0, i_10_289_3392_0, i_10_289_3610_0, i_10_289_3613_0,
    i_10_289_3647_0, i_10_289_3649_0, i_10_289_3653_0, i_10_289_3780_0,
    i_10_289_3781_0, i_10_289_3782_0, i_10_289_3837_0, i_10_289_3838_0,
    i_10_289_3839_0, i_10_289_3842_0, i_10_289_3856_0, i_10_289_3967_0,
    i_10_289_3985_0, i_10_289_4114_0, i_10_289_4291_0, i_10_289_4427_0;
  output o_10_289_0_0;
  assign o_10_289_0_0 = ~((~i_10_289_460_0 & ((~i_10_289_183_0 & ~i_10_289_184_0 & i_10_289_993_0) | (~i_10_289_174_0 & ~i_10_289_464_0 & ~i_10_289_514_0 & ~i_10_289_1006_0 & ~i_10_289_2469_0 & ~i_10_289_2722_0 & ~i_10_289_2731_0 & ~i_10_289_3195_0))) | (~i_10_289_464_0 & ((~i_10_289_174_0 & ~i_10_289_462_0 & ~i_10_289_1685_0 & ~i_10_289_3040_0) | (~i_10_289_749_0 & ~i_10_289_1244_0 & ~i_10_289_1950_0 & ~i_10_289_3199_0 & i_10_289_3838_0))) | (~i_10_289_174_0 & ((~i_10_289_1244_0 & i_10_289_1825_0 & i_10_289_1826_0 & ~i_10_289_2722_0 & ~i_10_289_3199_0 & ~i_10_289_3613_0) | (~i_10_289_124_0 & ~i_10_289_1820_0 & ~i_10_289_2469_0 & ~i_10_289_2734_0 & ~i_10_289_3196_0 & ~i_10_289_3780_0 & ~i_10_289_4114_0 & ~i_10_289_4291_0))) | (~i_10_289_124_0 & ((~i_10_289_446_0 & ~i_10_289_1363_0 & i_10_289_1825_0 & ~i_10_289_2731_0 & i_10_289_3199_0 & ~i_10_289_3838_0) | (~i_10_289_514_0 & ~i_10_289_2469_0 & ~i_10_289_3199_0 & ~i_10_289_3780_0 & i_10_289_3856_0 & ~i_10_289_4291_0))) | (~i_10_289_183_0 & ((~i_10_289_2734_0 & ((~i_10_289_280_0 & ~i_10_289_3198_0 & ~i_10_289_3837_0 & ((i_10_289_2632_0 & ~i_10_289_2702_0 & i_10_289_3196_0 & i_10_289_3649_0) | (~i_10_289_446_0 & ~i_10_289_955_0 & ~i_10_289_1037_0 & i_10_289_3610_0 & ~i_10_289_3780_0))) | (~i_10_289_1006_0 & ~i_10_289_2920_0 & ~i_10_289_3780_0 & ~i_10_289_3782_0))) | (~i_10_289_446_0 & ~i_10_289_1244_0 & ~i_10_289_1363_0 & i_10_289_1825_0 & ~i_10_289_1950_0 & ~i_10_289_2362_0) | (~i_10_289_993_0 & ~i_10_289_1037_0 & i_10_289_2632_0 & ~i_10_289_3649_0 & ~i_10_289_3837_0) | (~i_10_289_3041_0 & ~i_10_289_3195_0 & ~i_10_289_3197_0 & ~i_10_289_3199_0 & ~i_10_289_3838_0) | (~i_10_289_125_0 & ~i_10_289_184_0 & ~i_10_289_1823_0 & ~i_10_289_3613_0 & ~i_10_289_3839_0 & ~i_10_289_3985_0))) | (~i_10_289_3985_0 & ((~i_10_289_125_0 & ((~i_10_289_184_0 & ~i_10_289_462_0 & ~i_10_289_514_0 & ~i_10_289_1037_0 & ~i_10_289_1244_0 & ~i_10_289_1247_0 & i_10_289_1822_0 & ~i_10_289_1826_0 & ~i_10_289_2469_0) | (~i_10_289_280_0 & i_10_289_1310_0 & ~i_10_289_2920_0 & i_10_289_3653_0))) | (~i_10_289_514_0 & ~i_10_289_1037_0 & ~i_10_289_1823_0 & i_10_289_1826_0 & ~i_10_289_2734_0 & ~i_10_289_3782_0))) | (~i_10_289_462_0 & ((i_10_289_514_0 & i_10_289_1037_0) | (i_10_289_2455_0 & i_10_289_2830_0))) | (~i_10_289_1819_0 & ~i_10_289_3041_0 & ((~i_10_289_749_0 & ~i_10_289_1244_0 & ~i_10_289_1820_0 & ~i_10_289_3195_0 & ~i_10_289_3649_0 & ~i_10_289_3653_0) | (~i_10_289_184_0 & ~i_10_289_1950_0 & ~i_10_289_2920_0 & ~i_10_289_3782_0 & ~i_10_289_4114_0))) | (~i_10_289_3198_0 & ((~i_10_289_1820_0 & (i_10_289_317_0 | (~i_10_289_1653_0 & i_10_289_1826_0 & ~i_10_289_2830_0 & i_10_289_3653_0))) | (~i_10_289_280_0 & ~i_10_289_3195_0 & ~i_10_289_3196_0 & ~i_10_289_3197_0 & ~i_10_289_3839_0))) | (~i_10_289_3781_0 & ((i_10_289_286_0 & ~i_10_289_1363_0 & ~i_10_289_2362_0 & ~i_10_289_2829_0 & ~i_10_289_2920_0) | (~i_10_289_463_0 & ~i_10_289_1006_0 & ~i_10_289_3197_0))) | (~i_10_289_1247_0 & i_10_289_1825_0 & ~i_10_289_2361_0 & ~i_10_289_3610_0 & ~i_10_289_3613_0) | (i_10_289_2724_0 & ~i_10_289_3040_0 & ~i_10_289_3780_0));
endmodule



// Benchmark "kernel_10_290" written by ABC on Sun Jul 19 10:26:02 2020

module kernel_10_290 ( 
    i_10_290_36_0, i_10_290_64_0, i_10_290_68_0, i_10_290_119_0,
    i_10_290_191_0, i_10_290_254_0, i_10_290_262_0, i_10_290_316_0,
    i_10_290_319_0, i_10_290_411_0, i_10_290_433_0, i_10_290_443_0,
    i_10_290_448_0, i_10_290_497_0, i_10_290_514_0, i_10_290_515_0,
    i_10_290_695_0, i_10_290_712_0, i_10_290_829_0, i_10_290_830_0,
    i_10_290_1036_0, i_10_290_1037_0, i_10_290_1082_0, i_10_290_1099_0,
    i_10_290_1108_0, i_10_290_1109_0, i_10_290_1235_0, i_10_290_1265_0,
    i_10_290_1273_0, i_10_290_1301_0, i_10_290_1360_0, i_10_290_1361_0,
    i_10_290_1433_0, i_10_290_1451_0, i_10_290_1540_0, i_10_290_1541_0,
    i_10_290_1544_0, i_10_290_1621_0, i_10_290_1622_0, i_10_290_1739_0,
    i_10_290_1801_0, i_10_290_1802_0, i_10_290_1804_0, i_10_290_1874_0,
    i_10_290_1981_0, i_10_290_1996_0, i_10_290_1997_0, i_10_290_2018_0,
    i_10_290_2111_0, i_10_290_2153_0, i_10_290_2198_0, i_10_290_2201_0,
    i_10_290_2305_0, i_10_290_2306_0, i_10_290_2350_0, i_10_290_2351_0,
    i_10_290_2365_0, i_10_290_2376_0, i_10_290_2377_0, i_10_290_2467_0,
    i_10_290_2531_0, i_10_290_2558_0, i_10_290_2567_0, i_10_290_2585_0,
    i_10_290_2594_0, i_10_290_2609_0, i_10_290_2612_0, i_10_290_2615_0,
    i_10_290_2629_0, i_10_290_2653_0, i_10_290_2654_0, i_10_290_2675_0,
    i_10_290_2714_0, i_10_290_2830_0, i_10_290_2935_0, i_10_290_3092_0,
    i_10_290_3199_0, i_10_290_3280_0, i_10_290_3404_0, i_10_290_3410_0,
    i_10_290_3467_0, i_10_290_3494_0, i_10_290_3538_0, i_10_290_3584_0,
    i_10_290_3686_0, i_10_290_3692_0, i_10_290_3699_0, i_10_290_3794_0,
    i_10_290_3836_0, i_10_290_3839_0, i_10_290_3851_0, i_10_290_4115_0,
    i_10_290_4151_0, i_10_290_4154_0, i_10_290_4275_0, i_10_290_4278_0,
    i_10_290_4291_0, i_10_290_4547_0, i_10_290_4569_0, i_10_290_4571_0,
    o_10_290_0_0  );
  input  i_10_290_36_0, i_10_290_64_0, i_10_290_68_0, i_10_290_119_0,
    i_10_290_191_0, i_10_290_254_0, i_10_290_262_0, i_10_290_316_0,
    i_10_290_319_0, i_10_290_411_0, i_10_290_433_0, i_10_290_443_0,
    i_10_290_448_0, i_10_290_497_0, i_10_290_514_0, i_10_290_515_0,
    i_10_290_695_0, i_10_290_712_0, i_10_290_829_0, i_10_290_830_0,
    i_10_290_1036_0, i_10_290_1037_0, i_10_290_1082_0, i_10_290_1099_0,
    i_10_290_1108_0, i_10_290_1109_0, i_10_290_1235_0, i_10_290_1265_0,
    i_10_290_1273_0, i_10_290_1301_0, i_10_290_1360_0, i_10_290_1361_0,
    i_10_290_1433_0, i_10_290_1451_0, i_10_290_1540_0, i_10_290_1541_0,
    i_10_290_1544_0, i_10_290_1621_0, i_10_290_1622_0, i_10_290_1739_0,
    i_10_290_1801_0, i_10_290_1802_0, i_10_290_1804_0, i_10_290_1874_0,
    i_10_290_1981_0, i_10_290_1996_0, i_10_290_1997_0, i_10_290_2018_0,
    i_10_290_2111_0, i_10_290_2153_0, i_10_290_2198_0, i_10_290_2201_0,
    i_10_290_2305_0, i_10_290_2306_0, i_10_290_2350_0, i_10_290_2351_0,
    i_10_290_2365_0, i_10_290_2376_0, i_10_290_2377_0, i_10_290_2467_0,
    i_10_290_2531_0, i_10_290_2558_0, i_10_290_2567_0, i_10_290_2585_0,
    i_10_290_2594_0, i_10_290_2609_0, i_10_290_2612_0, i_10_290_2615_0,
    i_10_290_2629_0, i_10_290_2653_0, i_10_290_2654_0, i_10_290_2675_0,
    i_10_290_2714_0, i_10_290_2830_0, i_10_290_2935_0, i_10_290_3092_0,
    i_10_290_3199_0, i_10_290_3280_0, i_10_290_3404_0, i_10_290_3410_0,
    i_10_290_3467_0, i_10_290_3494_0, i_10_290_3538_0, i_10_290_3584_0,
    i_10_290_3686_0, i_10_290_3692_0, i_10_290_3699_0, i_10_290_3794_0,
    i_10_290_3836_0, i_10_290_3839_0, i_10_290_3851_0, i_10_290_4115_0,
    i_10_290_4151_0, i_10_290_4154_0, i_10_290_4275_0, i_10_290_4278_0,
    i_10_290_4291_0, i_10_290_4547_0, i_10_290_4569_0, i_10_290_4571_0;
  output o_10_290_0_0;
  assign o_10_290_0_0 = 0;
endmodule



// Benchmark "kernel_10_291" written by ABC on Sun Jul 19 10:26:03 2020

module kernel_10_291 ( 
    i_10_291_41_0, i_10_291_43_0, i_10_291_46_0, i_10_291_63_0,
    i_10_291_65_0, i_10_291_155_0, i_10_291_246_0, i_10_291_248_0,
    i_10_291_249_0, i_10_291_289_0, i_10_291_409_0, i_10_291_595_0,
    i_10_291_608_0, i_10_291_712_0, i_10_291_713_0, i_10_291_756_0,
    i_10_291_875_0, i_10_291_901_0, i_10_291_947_0, i_10_291_993_0,
    i_10_291_1010_0, i_10_291_1120_0, i_10_291_1157_0, i_10_291_1433_0,
    i_10_291_1488_0, i_10_291_1540_0, i_10_291_1614_0, i_10_291_1649_0,
    i_10_291_1703_0, i_10_291_1710_0, i_10_291_1802_0, i_10_291_1873_0,
    i_10_291_1915_0, i_10_291_1916_0, i_10_291_1947_0, i_10_291_2021_0,
    i_10_291_2030_0, i_10_291_2054_0, i_10_291_2109_0, i_10_291_2162_0,
    i_10_291_2180_0, i_10_291_2218_0, i_10_291_2304_0, i_10_291_2333_0,
    i_10_291_2336_0, i_10_291_2351_0, i_10_291_2359_0, i_10_291_2366_0,
    i_10_291_2431_0, i_10_291_2450_0, i_10_291_2451_0, i_10_291_2529_0,
    i_10_291_2602_0, i_10_291_2702_0, i_10_291_2705_0, i_10_291_2709_0,
    i_10_291_2713_0, i_10_291_2720_0, i_10_291_2863_0, i_10_291_2864_0,
    i_10_291_2923_0, i_10_291_3024_0, i_10_291_3071_0, i_10_291_3073_0,
    i_10_291_3074_0, i_10_291_3223_0, i_10_291_3227_0, i_10_291_3269_0,
    i_10_291_3278_0, i_10_291_3280_0, i_10_291_3287_0, i_10_291_3304_0,
    i_10_291_3330_0, i_10_291_3331_0, i_10_291_3385_0, i_10_291_3387_0,
    i_10_291_3403_0, i_10_291_3431_0, i_10_291_3523_0, i_10_291_3619_0,
    i_10_291_3647_0, i_10_291_3651_0, i_10_291_3730_0, i_10_291_3771_0,
    i_10_291_3774_0, i_10_291_3807_0, i_10_291_3834_0, i_10_291_3838_0,
    i_10_291_3839_0, i_10_291_3840_0, i_10_291_3849_0, i_10_291_3893_0,
    i_10_291_3902_0, i_10_291_3989_0, i_10_291_3993_0, i_10_291_4118_0,
    i_10_291_4188_0, i_10_291_4217_0, i_10_291_4302_0, i_10_291_4430_0,
    o_10_291_0_0  );
  input  i_10_291_41_0, i_10_291_43_0, i_10_291_46_0, i_10_291_63_0,
    i_10_291_65_0, i_10_291_155_0, i_10_291_246_0, i_10_291_248_0,
    i_10_291_249_0, i_10_291_289_0, i_10_291_409_0, i_10_291_595_0,
    i_10_291_608_0, i_10_291_712_0, i_10_291_713_0, i_10_291_756_0,
    i_10_291_875_0, i_10_291_901_0, i_10_291_947_0, i_10_291_993_0,
    i_10_291_1010_0, i_10_291_1120_0, i_10_291_1157_0, i_10_291_1433_0,
    i_10_291_1488_0, i_10_291_1540_0, i_10_291_1614_0, i_10_291_1649_0,
    i_10_291_1703_0, i_10_291_1710_0, i_10_291_1802_0, i_10_291_1873_0,
    i_10_291_1915_0, i_10_291_1916_0, i_10_291_1947_0, i_10_291_2021_0,
    i_10_291_2030_0, i_10_291_2054_0, i_10_291_2109_0, i_10_291_2162_0,
    i_10_291_2180_0, i_10_291_2218_0, i_10_291_2304_0, i_10_291_2333_0,
    i_10_291_2336_0, i_10_291_2351_0, i_10_291_2359_0, i_10_291_2366_0,
    i_10_291_2431_0, i_10_291_2450_0, i_10_291_2451_0, i_10_291_2529_0,
    i_10_291_2602_0, i_10_291_2702_0, i_10_291_2705_0, i_10_291_2709_0,
    i_10_291_2713_0, i_10_291_2720_0, i_10_291_2863_0, i_10_291_2864_0,
    i_10_291_2923_0, i_10_291_3024_0, i_10_291_3071_0, i_10_291_3073_0,
    i_10_291_3074_0, i_10_291_3223_0, i_10_291_3227_0, i_10_291_3269_0,
    i_10_291_3278_0, i_10_291_3280_0, i_10_291_3287_0, i_10_291_3304_0,
    i_10_291_3330_0, i_10_291_3331_0, i_10_291_3385_0, i_10_291_3387_0,
    i_10_291_3403_0, i_10_291_3431_0, i_10_291_3523_0, i_10_291_3619_0,
    i_10_291_3647_0, i_10_291_3651_0, i_10_291_3730_0, i_10_291_3771_0,
    i_10_291_3774_0, i_10_291_3807_0, i_10_291_3834_0, i_10_291_3838_0,
    i_10_291_3839_0, i_10_291_3840_0, i_10_291_3849_0, i_10_291_3893_0,
    i_10_291_3902_0, i_10_291_3989_0, i_10_291_3993_0, i_10_291_4118_0,
    i_10_291_4188_0, i_10_291_4217_0, i_10_291_4302_0, i_10_291_4430_0;
  output o_10_291_0_0;
  assign o_10_291_0_0 = 0;
endmodule



// Benchmark "kernel_10_292" written by ABC on Sun Jul 19 10:26:04 2020

module kernel_10_292 ( 
    i_10_292_68_0, i_10_292_175_0, i_10_292_247_0, i_10_292_273_0,
    i_10_292_319_0, i_10_292_328_0, i_10_292_355_0, i_10_292_363_0,
    i_10_292_390_0, i_10_292_425_0, i_10_292_435_0, i_10_292_442_0,
    i_10_292_443_0, i_10_292_465_0, i_10_292_518_0, i_10_292_608_0,
    i_10_292_631_0, i_10_292_734_0, i_10_292_736_0, i_10_292_793_0,
    i_10_292_794_0, i_10_292_796_0, i_10_292_799_0, i_10_292_908_0,
    i_10_292_956_0, i_10_292_977_0, i_10_292_993_0, i_10_292_1041_0,
    i_10_292_1163_0, i_10_292_1184_0, i_10_292_1194_0, i_10_292_1195_0,
    i_10_292_1220_0, i_10_292_1276_0, i_10_292_1360_0, i_10_292_1583_0,
    i_10_292_1683_0, i_10_292_1790_0, i_10_292_1894_0, i_10_292_1900_0,
    i_10_292_1911_0, i_10_292_1912_0, i_10_292_2003_0, i_10_292_2027_0,
    i_10_292_2030_0, i_10_292_2083_0, i_10_292_2158_0, i_10_292_2308_0,
    i_10_292_2309_0, i_10_292_2336_0, i_10_292_2359_0, i_10_292_2379_0,
    i_10_292_2381_0, i_10_292_2389_0, i_10_292_2480_0, i_10_292_2498_0,
    i_10_292_2542_0, i_10_292_2543_0, i_10_292_2603_0, i_10_292_2606_0,
    i_10_292_2629_0, i_10_292_2662_0, i_10_292_2727_0, i_10_292_2859_0,
    i_10_292_2923_0, i_10_292_2952_0, i_10_292_2983_0, i_10_292_2984_0,
    i_10_292_3044_0, i_10_292_3047_0, i_10_292_3056_0, i_10_292_3195_0,
    i_10_292_3196_0, i_10_292_3231_0, i_10_292_3273_0, i_10_292_3275_0,
    i_10_292_3300_0, i_10_292_3302_0, i_10_292_3325_0, i_10_292_3362_0,
    i_10_292_3363_0, i_10_292_3541_0, i_10_292_3647_0, i_10_292_3653_0,
    i_10_292_3684_0, i_10_292_3857_0, i_10_292_3875_0, i_10_292_3893_0,
    i_10_292_3945_0, i_10_292_3995_0, i_10_292_4113_0, i_10_292_4122_0,
    i_10_292_4220_0, i_10_292_4237_0, i_10_292_4275_0, i_10_292_4278_0,
    i_10_292_4295_0, i_10_292_4378_0, i_10_292_4381_0, i_10_292_4478_0,
    o_10_292_0_0  );
  input  i_10_292_68_0, i_10_292_175_0, i_10_292_247_0, i_10_292_273_0,
    i_10_292_319_0, i_10_292_328_0, i_10_292_355_0, i_10_292_363_0,
    i_10_292_390_0, i_10_292_425_0, i_10_292_435_0, i_10_292_442_0,
    i_10_292_443_0, i_10_292_465_0, i_10_292_518_0, i_10_292_608_0,
    i_10_292_631_0, i_10_292_734_0, i_10_292_736_0, i_10_292_793_0,
    i_10_292_794_0, i_10_292_796_0, i_10_292_799_0, i_10_292_908_0,
    i_10_292_956_0, i_10_292_977_0, i_10_292_993_0, i_10_292_1041_0,
    i_10_292_1163_0, i_10_292_1184_0, i_10_292_1194_0, i_10_292_1195_0,
    i_10_292_1220_0, i_10_292_1276_0, i_10_292_1360_0, i_10_292_1583_0,
    i_10_292_1683_0, i_10_292_1790_0, i_10_292_1894_0, i_10_292_1900_0,
    i_10_292_1911_0, i_10_292_1912_0, i_10_292_2003_0, i_10_292_2027_0,
    i_10_292_2030_0, i_10_292_2083_0, i_10_292_2158_0, i_10_292_2308_0,
    i_10_292_2309_0, i_10_292_2336_0, i_10_292_2359_0, i_10_292_2379_0,
    i_10_292_2381_0, i_10_292_2389_0, i_10_292_2480_0, i_10_292_2498_0,
    i_10_292_2542_0, i_10_292_2543_0, i_10_292_2603_0, i_10_292_2606_0,
    i_10_292_2629_0, i_10_292_2662_0, i_10_292_2727_0, i_10_292_2859_0,
    i_10_292_2923_0, i_10_292_2952_0, i_10_292_2983_0, i_10_292_2984_0,
    i_10_292_3044_0, i_10_292_3047_0, i_10_292_3056_0, i_10_292_3195_0,
    i_10_292_3196_0, i_10_292_3231_0, i_10_292_3273_0, i_10_292_3275_0,
    i_10_292_3300_0, i_10_292_3302_0, i_10_292_3325_0, i_10_292_3362_0,
    i_10_292_3363_0, i_10_292_3541_0, i_10_292_3647_0, i_10_292_3653_0,
    i_10_292_3684_0, i_10_292_3857_0, i_10_292_3875_0, i_10_292_3893_0,
    i_10_292_3945_0, i_10_292_3995_0, i_10_292_4113_0, i_10_292_4122_0,
    i_10_292_4220_0, i_10_292_4237_0, i_10_292_4275_0, i_10_292_4278_0,
    i_10_292_4295_0, i_10_292_4378_0, i_10_292_4381_0, i_10_292_4478_0;
  output o_10_292_0_0;
  assign o_10_292_0_0 = 0;
endmodule



// Benchmark "kernel_10_293" written by ABC on Sun Jul 19 10:26:05 2020

module kernel_10_293 ( 
    i_10_293_28_0, i_10_293_29_0, i_10_293_31_0, i_10_293_32_0,
    i_10_293_45_0, i_10_293_46_0, i_10_293_124_0, i_10_293_224_0,
    i_10_293_408_0, i_10_293_437_0, i_10_293_443_0, i_10_293_444_0,
    i_10_293_461_0, i_10_293_465_0, i_10_293_466_0, i_10_293_516_0,
    i_10_293_517_0, i_10_293_732_0, i_10_293_733_0, i_10_293_753_0,
    i_10_293_754_0, i_10_293_755_0, i_10_293_928_0, i_10_293_961_0,
    i_10_293_1032_0, i_10_293_1305_0, i_10_293_1306_0, i_10_293_1310_0,
    i_10_293_1312_0, i_10_293_1313_0, i_10_293_1546_0, i_10_293_1559_0,
    i_10_293_1616_0, i_10_293_1648_0, i_10_293_1800_0, i_10_293_1818_0,
    i_10_293_1948_0, i_10_293_1949_0, i_10_293_1951_0, i_10_293_1952_0,
    i_10_293_2006_0, i_10_293_2366_0, i_10_293_2407_0, i_10_293_2473_0,
    i_10_293_2603_0, i_10_293_2632_0, i_10_293_2633_0, i_10_293_2635_0,
    i_10_293_2655_0, i_10_293_2656_0, i_10_293_2657_0, i_10_293_2660_0,
    i_10_293_2718_0, i_10_293_2719_0, i_10_293_2722_0, i_10_293_2723_0,
    i_10_293_2724_0, i_10_293_2726_0, i_10_293_2735_0, i_10_293_2826_0,
    i_10_293_2827_0, i_10_293_2828_0, i_10_293_2887_0, i_10_293_2924_0,
    i_10_293_2986_0, i_10_293_3036_0, i_10_293_3039_0, i_10_293_3040_0,
    i_10_293_3041_0, i_10_293_3045_0, i_10_293_3046_0, i_10_293_3196_0,
    i_10_293_3276_0, i_10_293_3278_0, i_10_293_3279_0, i_10_293_3349_0,
    i_10_293_3390_0, i_10_293_3391_0, i_10_293_3392_0, i_10_293_3494_0,
    i_10_293_3522_0, i_10_293_3587_0, i_10_293_3610_0, i_10_293_3611_0,
    i_10_293_3646_0, i_10_293_3649_0, i_10_293_3651_0, i_10_293_3653_0,
    i_10_293_3688_0, i_10_293_3689_0, i_10_293_3727_0, i_10_293_3728_0,
    i_10_293_3780_0, i_10_293_3781_0, i_10_293_3852_0, i_10_293_3853_0,
    i_10_293_3856_0, i_10_293_3859_0, i_10_293_4025_0, i_10_293_4127_0,
    o_10_293_0_0  );
  input  i_10_293_28_0, i_10_293_29_0, i_10_293_31_0, i_10_293_32_0,
    i_10_293_45_0, i_10_293_46_0, i_10_293_124_0, i_10_293_224_0,
    i_10_293_408_0, i_10_293_437_0, i_10_293_443_0, i_10_293_444_0,
    i_10_293_461_0, i_10_293_465_0, i_10_293_466_0, i_10_293_516_0,
    i_10_293_517_0, i_10_293_732_0, i_10_293_733_0, i_10_293_753_0,
    i_10_293_754_0, i_10_293_755_0, i_10_293_928_0, i_10_293_961_0,
    i_10_293_1032_0, i_10_293_1305_0, i_10_293_1306_0, i_10_293_1310_0,
    i_10_293_1312_0, i_10_293_1313_0, i_10_293_1546_0, i_10_293_1559_0,
    i_10_293_1616_0, i_10_293_1648_0, i_10_293_1800_0, i_10_293_1818_0,
    i_10_293_1948_0, i_10_293_1949_0, i_10_293_1951_0, i_10_293_1952_0,
    i_10_293_2006_0, i_10_293_2366_0, i_10_293_2407_0, i_10_293_2473_0,
    i_10_293_2603_0, i_10_293_2632_0, i_10_293_2633_0, i_10_293_2635_0,
    i_10_293_2655_0, i_10_293_2656_0, i_10_293_2657_0, i_10_293_2660_0,
    i_10_293_2718_0, i_10_293_2719_0, i_10_293_2722_0, i_10_293_2723_0,
    i_10_293_2724_0, i_10_293_2726_0, i_10_293_2735_0, i_10_293_2826_0,
    i_10_293_2827_0, i_10_293_2828_0, i_10_293_2887_0, i_10_293_2924_0,
    i_10_293_2986_0, i_10_293_3036_0, i_10_293_3039_0, i_10_293_3040_0,
    i_10_293_3041_0, i_10_293_3045_0, i_10_293_3046_0, i_10_293_3196_0,
    i_10_293_3276_0, i_10_293_3278_0, i_10_293_3279_0, i_10_293_3349_0,
    i_10_293_3390_0, i_10_293_3391_0, i_10_293_3392_0, i_10_293_3494_0,
    i_10_293_3522_0, i_10_293_3587_0, i_10_293_3610_0, i_10_293_3611_0,
    i_10_293_3646_0, i_10_293_3649_0, i_10_293_3651_0, i_10_293_3653_0,
    i_10_293_3688_0, i_10_293_3689_0, i_10_293_3727_0, i_10_293_3728_0,
    i_10_293_3780_0, i_10_293_3781_0, i_10_293_3852_0, i_10_293_3853_0,
    i_10_293_3856_0, i_10_293_3859_0, i_10_293_4025_0, i_10_293_4127_0;
  output o_10_293_0_0;
  assign o_10_293_0_0 = 0;
endmodule



// Benchmark "kernel_10_294" written by ABC on Sun Jul 19 10:26:06 2020

module kernel_10_294 ( 
    i_10_294_118_0, i_10_294_175_0, i_10_294_186_0, i_10_294_243_0,
    i_10_294_282_0, i_10_294_283_0, i_10_294_284_0, i_10_294_285_0,
    i_10_294_318_0, i_10_294_319_0, i_10_294_408_0, i_10_294_409_0,
    i_10_294_410_0, i_10_294_412_0, i_10_294_430_0, i_10_294_431_0,
    i_10_294_460_0, i_10_294_461_0, i_10_294_508_0, i_10_294_511_0,
    i_10_294_737_0, i_10_294_1002_0, i_10_294_1135_0, i_10_294_1168_0,
    i_10_294_1234_0, i_10_294_1235_0, i_10_294_1237_0, i_10_294_1238_0,
    i_10_294_1307_0, i_10_294_1309_0, i_10_294_1310_0, i_10_294_1552_0,
    i_10_294_1555_0, i_10_294_1575_0, i_10_294_1582_0, i_10_294_1615_0,
    i_10_294_1647_0, i_10_294_1652_0, i_10_294_1653_0, i_10_294_1681_0,
    i_10_294_1687_0, i_10_294_1821_0, i_10_294_1822_0, i_10_294_1823_0,
    i_10_294_1825_0, i_10_294_1826_0, i_10_294_1914_0, i_10_294_1915_0,
    i_10_294_1916_0, i_10_294_2022_0, i_10_294_2311_0, i_10_294_2355_0,
    i_10_294_2362_0, i_10_294_2383_0, i_10_294_2453_0, i_10_294_2456_0,
    i_10_294_2473_0, i_10_294_2631_0, i_10_294_2634_0, i_10_294_2655_0,
    i_10_294_2656_0, i_10_294_2658_0, i_10_294_2659_0, i_10_294_2679_0,
    i_10_294_2704_0, i_10_294_2706_0, i_10_294_2707_0, i_10_294_2715_0,
    i_10_294_2716_0, i_10_294_2719_0, i_10_294_2735_0, i_10_294_2788_0,
    i_10_294_2831_0, i_10_294_2888_0, i_10_294_2983_0, i_10_294_3034_0,
    i_10_294_3040_0, i_10_294_3044_0, i_10_294_3046_0, i_10_294_3196_0,
    i_10_294_3197_0, i_10_294_3279_0, i_10_294_3319_0, i_10_294_3387_0,
    i_10_294_3392_0, i_10_294_3405_0, i_10_294_3409_0, i_10_294_3613_0,
    i_10_294_3783_0, i_10_294_3835_0, i_10_294_3840_0, i_10_294_3842_0,
    i_10_294_3847_0, i_10_294_3854_0, i_10_294_3981_0, i_10_294_4050_0,
    i_10_294_4119_0, i_10_294_4130_0, i_10_294_4191_0, i_10_294_4289_0,
    o_10_294_0_0  );
  input  i_10_294_118_0, i_10_294_175_0, i_10_294_186_0, i_10_294_243_0,
    i_10_294_282_0, i_10_294_283_0, i_10_294_284_0, i_10_294_285_0,
    i_10_294_318_0, i_10_294_319_0, i_10_294_408_0, i_10_294_409_0,
    i_10_294_410_0, i_10_294_412_0, i_10_294_430_0, i_10_294_431_0,
    i_10_294_460_0, i_10_294_461_0, i_10_294_508_0, i_10_294_511_0,
    i_10_294_737_0, i_10_294_1002_0, i_10_294_1135_0, i_10_294_1168_0,
    i_10_294_1234_0, i_10_294_1235_0, i_10_294_1237_0, i_10_294_1238_0,
    i_10_294_1307_0, i_10_294_1309_0, i_10_294_1310_0, i_10_294_1552_0,
    i_10_294_1555_0, i_10_294_1575_0, i_10_294_1582_0, i_10_294_1615_0,
    i_10_294_1647_0, i_10_294_1652_0, i_10_294_1653_0, i_10_294_1681_0,
    i_10_294_1687_0, i_10_294_1821_0, i_10_294_1822_0, i_10_294_1823_0,
    i_10_294_1825_0, i_10_294_1826_0, i_10_294_1914_0, i_10_294_1915_0,
    i_10_294_1916_0, i_10_294_2022_0, i_10_294_2311_0, i_10_294_2355_0,
    i_10_294_2362_0, i_10_294_2383_0, i_10_294_2453_0, i_10_294_2456_0,
    i_10_294_2473_0, i_10_294_2631_0, i_10_294_2634_0, i_10_294_2655_0,
    i_10_294_2656_0, i_10_294_2658_0, i_10_294_2659_0, i_10_294_2679_0,
    i_10_294_2704_0, i_10_294_2706_0, i_10_294_2707_0, i_10_294_2715_0,
    i_10_294_2716_0, i_10_294_2719_0, i_10_294_2735_0, i_10_294_2788_0,
    i_10_294_2831_0, i_10_294_2888_0, i_10_294_2983_0, i_10_294_3034_0,
    i_10_294_3040_0, i_10_294_3044_0, i_10_294_3046_0, i_10_294_3196_0,
    i_10_294_3197_0, i_10_294_3279_0, i_10_294_3319_0, i_10_294_3387_0,
    i_10_294_3392_0, i_10_294_3405_0, i_10_294_3409_0, i_10_294_3613_0,
    i_10_294_3783_0, i_10_294_3835_0, i_10_294_3840_0, i_10_294_3842_0,
    i_10_294_3847_0, i_10_294_3854_0, i_10_294_3981_0, i_10_294_4050_0,
    i_10_294_4119_0, i_10_294_4130_0, i_10_294_4191_0, i_10_294_4289_0;
  output o_10_294_0_0;
  assign o_10_294_0_0 = ~((~i_10_294_282_0 & ((~i_10_294_118_0 & ~i_10_294_319_0 & ~i_10_294_408_0 & ~i_10_294_412_0 & ~i_10_294_1310_0 & ~i_10_294_3405_0) | (~i_10_294_284_0 & ~i_10_294_1307_0 & i_10_294_1309_0 & i_10_294_1821_0 & ~i_10_294_3034_0 & ~i_10_294_4119_0))) | (~i_10_294_283_0 & ((~i_10_294_318_0 & ((~i_10_294_409_0 & ~i_10_294_1822_0) | (~i_10_294_284_0 & ~i_10_294_319_0 & ~i_10_294_2655_0 & ~i_10_294_2706_0 & i_10_294_3847_0))) | (~i_10_294_1168_0 & ~i_10_294_1234_0 & ~i_10_294_2679_0 & ~i_10_294_2716_0 & i_10_294_3613_0 & ~i_10_294_3854_0 & ~i_10_294_4050_0 & ~i_10_294_4130_0))) | (~i_10_294_408_0 & ((~i_10_294_409_0 & ~i_10_294_2656_0 & ((~i_10_294_2735_0 & ~i_10_294_2831_0 & ~i_10_294_3387_0) | (~i_10_294_186_0 & ~i_10_294_412_0 & ~i_10_294_3613_0))) | (~i_10_294_412_0 & ~i_10_294_461_0 & i_10_294_1825_0 & ~i_10_294_2362_0 & ~i_10_294_2634_0) | (~i_10_294_118_0 & ~i_10_294_410_0 & ~i_10_294_1238_0 & ~i_10_294_2022_0 & ~i_10_294_4050_0))) | (~i_10_294_186_0 & ~i_10_294_1234_0 & ((~i_10_294_1237_0 & ~i_10_294_1582_0 & ~i_10_294_1821_0 & ~i_10_294_2453_0 & ~i_10_294_2788_0) | (~i_10_294_118_0 & ~i_10_294_243_0 & ~i_10_294_409_0 & ~i_10_294_2704_0 & ~i_10_294_3044_0 & ~i_10_294_3854_0))) | (~i_10_294_243_0 & ((~i_10_294_1652_0 & ~i_10_294_1653_0 & ~i_10_294_1821_0 & ~i_10_294_1823_0 & ~i_10_294_2456_0 & ~i_10_294_3387_0 & ~i_10_294_4130_0) | (~i_10_294_409_0 & ~i_10_294_1307_0 & ~i_10_294_3783_0 & i_10_294_4289_0))) | (~i_10_294_409_0 & ((~i_10_294_1821_0 & ~i_10_294_1823_0 & i_10_294_2355_0 & ~i_10_294_2715_0) | (i_10_294_1825_0 & ~i_10_294_4050_0))) | (~i_10_294_118_0 & ((~i_10_294_410_0 & ((~i_10_294_1822_0 & ~i_10_294_1823_0 & ~i_10_294_2022_0 & ~i_10_294_3044_0 & ~i_10_294_3279_0 & ~i_10_294_3392_0 & ~i_10_294_3847_0) | (~i_10_294_2355_0 & ~i_10_294_2658_0 & ~i_10_294_2706_0 & ~i_10_294_4050_0))) | (i_10_294_175_0 & i_10_294_1307_0 & ~i_10_294_3040_0 & i_10_294_3196_0))) | (~i_10_294_2362_0 & ((i_10_294_1309_0 & ~i_10_294_2658_0 & ~i_10_294_2659_0 & ~i_10_294_2707_0 & ~i_10_294_2983_0 & i_10_294_3613_0 & ~i_10_294_3783_0 & ~i_10_294_4050_0) | (~i_10_294_1237_0 & i_10_294_1310_0 & ~i_10_294_1652_0 & ~i_10_294_2634_0 & ~i_10_294_3854_0 & ~i_10_294_4130_0))) | (~i_10_294_4119_0 & ((~i_10_294_175_0 & ~i_10_294_1653_0 & ~i_10_294_2831_0 & i_10_294_3040_0) | (~i_10_294_319_0 & i_10_294_1652_0 & ~i_10_294_1821_0 & ~i_10_294_3405_0 & ~i_10_294_3847_0 & ~i_10_294_3854_0))) | (i_10_294_1687_0 & ~i_10_294_3613_0));
endmodule



// Benchmark "kernel_10_295" written by ABC on Sun Jul 19 10:26:08 2020

module kernel_10_295 ( 
    i_10_295_28_0, i_10_295_171_0, i_10_295_174_0, i_10_295_178_0,
    i_10_295_183_0, i_10_295_185_0, i_10_295_317_0, i_10_295_390_0,
    i_10_295_410_0, i_10_295_427_0, i_10_295_442_0, i_10_295_443_0,
    i_10_295_459_0, i_10_295_566_0, i_10_295_748_0, i_10_295_792_0,
    i_10_295_798_0, i_10_295_1027_0, i_10_295_1033_0, i_10_295_1034_0,
    i_10_295_1042_0, i_10_295_1043_0, i_10_295_1236_0, i_10_295_1245_0,
    i_10_295_1246_0, i_10_295_1247_0, i_10_295_1539_0, i_10_295_1542_0,
    i_10_295_1543_0, i_10_295_1575_0, i_10_295_1576_0, i_10_295_1650_0,
    i_10_295_1655_0, i_10_295_1683_0, i_10_295_1684_0, i_10_295_1686_0,
    i_10_295_1688_0, i_10_295_1769_0, i_10_295_1911_0, i_10_295_1912_0,
    i_10_295_1913_0, i_10_295_1915_0, i_10_295_1948_0, i_10_295_1949_0,
    i_10_295_1997_0, i_10_295_2201_0, i_10_295_2353_0, i_10_295_2380_0,
    i_10_295_2448_0, i_10_295_2470_0, i_10_295_2632_0, i_10_295_2636_0,
    i_10_295_2659_0, i_10_295_2661_0, i_10_295_2662_0, i_10_295_2701_0,
    i_10_295_2706_0, i_10_295_2709_0, i_10_295_2721_0, i_10_295_2723_0,
    i_10_295_2728_0, i_10_295_2729_0, i_10_295_2827_0, i_10_295_2828_0,
    i_10_295_2831_0, i_10_295_3035_0, i_10_295_3040_0, i_10_295_3041_0,
    i_10_295_3043_0, i_10_295_3152_0, i_10_295_3198_0, i_10_295_3199_0,
    i_10_295_3277_0, i_10_295_3329_0, i_10_295_3388_0, i_10_295_3497_0,
    i_10_295_3525_0, i_10_295_3583_0, i_10_295_3586_0, i_10_295_3614_0,
    i_10_295_3649_0, i_10_295_3653_0, i_10_295_3780_0, i_10_295_3783_0,
    i_10_295_3837_0, i_10_295_3839_0, i_10_295_3855_0, i_10_295_3858_0,
    i_10_295_3894_0, i_10_295_3895_0, i_10_295_3896_0, i_10_295_3985_0,
    i_10_295_4116_0, i_10_295_4128_0, i_10_295_4129_0, i_10_295_4169_0,
    i_10_295_4276_0, i_10_295_4290_0, i_10_295_4291_0, i_10_295_4535_0,
    o_10_295_0_0  );
  input  i_10_295_28_0, i_10_295_171_0, i_10_295_174_0, i_10_295_178_0,
    i_10_295_183_0, i_10_295_185_0, i_10_295_317_0, i_10_295_390_0,
    i_10_295_410_0, i_10_295_427_0, i_10_295_442_0, i_10_295_443_0,
    i_10_295_459_0, i_10_295_566_0, i_10_295_748_0, i_10_295_792_0,
    i_10_295_798_0, i_10_295_1027_0, i_10_295_1033_0, i_10_295_1034_0,
    i_10_295_1042_0, i_10_295_1043_0, i_10_295_1236_0, i_10_295_1245_0,
    i_10_295_1246_0, i_10_295_1247_0, i_10_295_1539_0, i_10_295_1542_0,
    i_10_295_1543_0, i_10_295_1575_0, i_10_295_1576_0, i_10_295_1650_0,
    i_10_295_1655_0, i_10_295_1683_0, i_10_295_1684_0, i_10_295_1686_0,
    i_10_295_1688_0, i_10_295_1769_0, i_10_295_1911_0, i_10_295_1912_0,
    i_10_295_1913_0, i_10_295_1915_0, i_10_295_1948_0, i_10_295_1949_0,
    i_10_295_1997_0, i_10_295_2201_0, i_10_295_2353_0, i_10_295_2380_0,
    i_10_295_2448_0, i_10_295_2470_0, i_10_295_2632_0, i_10_295_2636_0,
    i_10_295_2659_0, i_10_295_2661_0, i_10_295_2662_0, i_10_295_2701_0,
    i_10_295_2706_0, i_10_295_2709_0, i_10_295_2721_0, i_10_295_2723_0,
    i_10_295_2728_0, i_10_295_2729_0, i_10_295_2827_0, i_10_295_2828_0,
    i_10_295_2831_0, i_10_295_3035_0, i_10_295_3040_0, i_10_295_3041_0,
    i_10_295_3043_0, i_10_295_3152_0, i_10_295_3198_0, i_10_295_3199_0,
    i_10_295_3277_0, i_10_295_3329_0, i_10_295_3388_0, i_10_295_3497_0,
    i_10_295_3525_0, i_10_295_3583_0, i_10_295_3586_0, i_10_295_3614_0,
    i_10_295_3649_0, i_10_295_3653_0, i_10_295_3780_0, i_10_295_3783_0,
    i_10_295_3837_0, i_10_295_3839_0, i_10_295_3855_0, i_10_295_3858_0,
    i_10_295_3894_0, i_10_295_3895_0, i_10_295_3896_0, i_10_295_3985_0,
    i_10_295_4116_0, i_10_295_4128_0, i_10_295_4129_0, i_10_295_4169_0,
    i_10_295_4276_0, i_10_295_4290_0, i_10_295_4291_0, i_10_295_4535_0;
  output o_10_295_0_0;
  assign o_10_295_0_0 = ~((~i_10_295_28_0 & ((~i_10_295_317_0 & i_10_295_1033_0 & ~i_10_295_2448_0 & ~i_10_295_2632_0 & ~i_10_295_3614_0) | (~i_10_295_183_0 & ~i_10_295_185_0 & ~i_10_295_390_0 & ~i_10_295_1043_0 & ~i_10_295_1542_0 & ~i_10_295_1575_0 & ~i_10_295_2201_0 & ~i_10_295_3653_0 & ~i_10_295_3985_0))) | (~i_10_295_798_0 & ((i_10_295_171_0 & i_10_295_2659_0 & ~i_10_295_2661_0 & ~i_10_295_3614_0) | (~i_10_295_1539_0 & ~i_10_295_1576_0 & ~i_10_295_2828_0 & ~i_10_295_2831_0 & ~i_10_295_3896_0))) | (~i_10_295_2709_0 & ((~i_10_295_1246_0 & ((~i_10_295_1769_0 & ~i_10_295_2448_0 & ~i_10_295_3198_0 & ~i_10_295_3839_0 & ~i_10_295_4276_0) | (~i_10_295_317_0 & ~i_10_295_1684_0 & ~i_10_295_1686_0 & ~i_10_295_1911_0 & ~i_10_295_2636_0 & ~i_10_295_3043_0 & ~i_10_295_3388_0 & ~i_10_295_3896_0 & ~i_10_295_4291_0))) | (~i_10_295_174_0 & ~i_10_295_1042_0 & ~i_10_295_1575_0 & ~i_10_295_1686_0 & ~i_10_295_1769_0 & ~i_10_295_2659_0 & ~i_10_295_2721_0 & ~i_10_295_3041_0 & ~i_10_295_3837_0))) | (~i_10_295_1042_0 & ((~i_10_295_390_0 & ((~i_10_295_185_0 & ~i_10_295_1236_0 & ~i_10_295_1575_0 & ~i_10_295_1683_0 & ~i_10_295_1769_0 & ~i_10_295_2659_0 & ~i_10_295_2827_0 & ~i_10_295_3277_0) | (~i_10_295_171_0 & ~i_10_295_1650_0 & ~i_10_295_1912_0 & ~i_10_295_2729_0 & ~i_10_295_3041_0 & i_10_295_3388_0 & ~i_10_295_3894_0))) | (~i_10_295_748_0 & ~i_10_295_1043_0 & ~i_10_295_1575_0 & ~i_10_295_3040_0 & ~i_10_295_3198_0 & ~i_10_295_4169_0))) | (~i_10_295_171_0 & ~i_10_295_3614_0 & ((~i_10_295_1913_0 & i_10_295_2659_0 & i_10_295_2721_0 & ~i_10_295_3277_0 & ~i_10_295_3780_0 & ~i_10_295_3837_0) | (~i_10_295_1245_0 & ~i_10_295_1539_0 & i_10_295_2353_0 & ~i_10_295_2721_0 & ~i_10_295_3855_0 & ~i_10_295_3896_0))) | (~i_10_295_1911_0 & ((~i_10_295_185_0 & ~i_10_295_1236_0 & ((~i_10_295_748_0 & ~i_10_295_1027_0 & ~i_10_295_1539_0 & ~i_10_295_1769_0 & ~i_10_295_2729_0 & ~i_10_295_3035_0 & ~i_10_295_3198_0) | (~i_10_295_1245_0 & ~i_10_295_1542_0 & ~i_10_295_1576_0 & ~i_10_295_1915_0 & ~i_10_295_2828_0 & ~i_10_295_3043_0 & ~i_10_295_3895_0))) | (~i_10_295_178_0 & ~i_10_295_390_0 & ~i_10_295_748_0 & ~i_10_295_1043_0 & ~i_10_295_1683_0 & ~i_10_295_1912_0 & ~i_10_295_1915_0 & ~i_10_295_2448_0 & ~i_10_295_3199_0 & ~i_10_295_4290_0))) | (~i_10_295_1539_0 & ((~i_10_295_410_0 & ~i_10_295_1245_0 & ~i_10_295_1769_0 & ~i_10_295_2201_0 & ~i_10_295_3277_0 & ~i_10_295_3855_0 & ~i_10_295_3895_0 & ~i_10_295_3896_0) | (~i_10_295_183_0 & i_10_295_442_0 & ~i_10_295_1688_0 & ~i_10_295_4169_0))) | (~i_10_295_2721_0 & ((~i_10_295_443_0 & ~i_10_295_1043_0 & ~i_10_295_1684_0 & ~i_10_295_2728_0 & ~i_10_295_3388_0 & ~i_10_295_3780_0 & ~i_10_295_3783_0 & ~i_10_295_3894_0) | (~i_10_295_748_0 & ~i_10_295_792_0 & ~i_10_295_3041_0 & i_10_295_3586_0 & ~i_10_295_4276_0))) | (i_10_295_317_0 & ~i_10_295_2632_0 & ~i_10_295_3839_0) | (i_10_295_174_0 & i_10_295_178_0 & ~i_10_295_1033_0 & i_10_295_2706_0 & ~i_10_295_3040_0 & ~i_10_295_3858_0) | (i_10_295_1769_0 & i_10_295_2662_0 & ~i_10_295_3985_0) | (~i_10_295_390_0 & ~i_10_295_566_0 & ~i_10_295_1912_0 & ~i_10_295_1913_0 & i_10_295_2448_0 & ~i_10_295_3783_0 & ~i_10_295_3894_0 & ~i_10_295_4128_0) | (i_10_295_443_0 & i_10_295_1043_0 & ~i_10_295_4291_0));
endmodule



// Benchmark "kernel_10_296" written by ABC on Sun Jul 19 10:26:09 2020

module kernel_10_296 ( 
    i_10_296_9_0, i_10_296_223_0, i_10_296_270_0, i_10_296_272_0,
    i_10_296_279_0, i_10_296_285_0, i_10_296_447_0, i_10_296_462_0,
    i_10_296_464_0, i_10_296_505_0, i_10_296_506_0, i_10_296_507_0,
    i_10_296_508_0, i_10_296_513_0, i_10_296_516_0, i_10_296_711_0,
    i_10_296_712_0, i_10_296_749_0, i_10_296_957_0, i_10_296_967_0,
    i_10_296_999_0, i_10_296_1080_0, i_10_296_1083_0, i_10_296_1098_0,
    i_10_296_1215_0, i_10_296_1239_0, i_10_296_1263_0, i_10_296_1306_0,
    i_10_296_1539_0, i_10_296_1549_0, i_10_296_1578_0, i_10_296_1653_0,
    i_10_296_1686_0, i_10_296_1782_0, i_10_296_1821_0, i_10_296_1822_0,
    i_10_296_1990_0, i_10_296_2016_0, i_10_296_2088_0, i_10_296_2179_0,
    i_10_296_2196_0, i_10_296_2197_0, i_10_296_2199_0, i_10_296_2352_0,
    i_10_296_2376_0, i_10_296_2448_0, i_10_296_2502_0, i_10_296_2574_0,
    i_10_296_2604_0, i_10_296_2610_0, i_10_296_2629_0, i_10_296_2630_0,
    i_10_296_2631_0, i_10_296_2655_0, i_10_296_2659_0, i_10_296_2662_0,
    i_10_296_2673_0, i_10_296_2700_0, i_10_296_2701_0, i_10_296_2703_0,
    i_10_296_2713_0, i_10_296_2882_0, i_10_296_2917_0, i_10_296_2979_0,
    i_10_296_3046_0, i_10_296_3054_0, i_10_296_3055_0, i_10_296_3088_0,
    i_10_296_3158_0, i_10_296_3328_0, i_10_296_3329_0, i_10_296_3385_0,
    i_10_296_3387_0, i_10_296_3538_0, i_10_296_3616_0, i_10_296_3681_0,
    i_10_296_3781_0, i_10_296_3785_0, i_10_296_3844_0, i_10_296_3852_0,
    i_10_296_3853_0, i_10_296_3854_0, i_10_296_3855_0, i_10_296_3858_0,
    i_10_296_3859_0, i_10_296_3860_0, i_10_296_3978_0, i_10_296_3979_0,
    i_10_296_4122_0, i_10_296_4123_0, i_10_296_4126_0, i_10_296_4167_0,
    i_10_296_4168_0, i_10_296_4170_0, i_10_296_4266_0, i_10_296_4267_0,
    i_10_296_4269_0, i_10_296_4275_0, i_10_296_4278_0, i_10_296_4567_0,
    o_10_296_0_0  );
  input  i_10_296_9_0, i_10_296_223_0, i_10_296_270_0, i_10_296_272_0,
    i_10_296_279_0, i_10_296_285_0, i_10_296_447_0, i_10_296_462_0,
    i_10_296_464_0, i_10_296_505_0, i_10_296_506_0, i_10_296_507_0,
    i_10_296_508_0, i_10_296_513_0, i_10_296_516_0, i_10_296_711_0,
    i_10_296_712_0, i_10_296_749_0, i_10_296_957_0, i_10_296_967_0,
    i_10_296_999_0, i_10_296_1080_0, i_10_296_1083_0, i_10_296_1098_0,
    i_10_296_1215_0, i_10_296_1239_0, i_10_296_1263_0, i_10_296_1306_0,
    i_10_296_1539_0, i_10_296_1549_0, i_10_296_1578_0, i_10_296_1653_0,
    i_10_296_1686_0, i_10_296_1782_0, i_10_296_1821_0, i_10_296_1822_0,
    i_10_296_1990_0, i_10_296_2016_0, i_10_296_2088_0, i_10_296_2179_0,
    i_10_296_2196_0, i_10_296_2197_0, i_10_296_2199_0, i_10_296_2352_0,
    i_10_296_2376_0, i_10_296_2448_0, i_10_296_2502_0, i_10_296_2574_0,
    i_10_296_2604_0, i_10_296_2610_0, i_10_296_2629_0, i_10_296_2630_0,
    i_10_296_2631_0, i_10_296_2655_0, i_10_296_2659_0, i_10_296_2662_0,
    i_10_296_2673_0, i_10_296_2700_0, i_10_296_2701_0, i_10_296_2703_0,
    i_10_296_2713_0, i_10_296_2882_0, i_10_296_2917_0, i_10_296_2979_0,
    i_10_296_3046_0, i_10_296_3054_0, i_10_296_3055_0, i_10_296_3088_0,
    i_10_296_3158_0, i_10_296_3328_0, i_10_296_3329_0, i_10_296_3385_0,
    i_10_296_3387_0, i_10_296_3538_0, i_10_296_3616_0, i_10_296_3681_0,
    i_10_296_3781_0, i_10_296_3785_0, i_10_296_3844_0, i_10_296_3852_0,
    i_10_296_3853_0, i_10_296_3854_0, i_10_296_3855_0, i_10_296_3858_0,
    i_10_296_3859_0, i_10_296_3860_0, i_10_296_3978_0, i_10_296_3979_0,
    i_10_296_4122_0, i_10_296_4123_0, i_10_296_4126_0, i_10_296_4167_0,
    i_10_296_4168_0, i_10_296_4170_0, i_10_296_4266_0, i_10_296_4267_0,
    i_10_296_4269_0, i_10_296_4275_0, i_10_296_4278_0, i_10_296_4567_0;
  output o_10_296_0_0;
  assign o_10_296_0_0 = ~((~i_10_296_516_0 & ((~i_10_296_749_0 & ~i_10_296_1539_0 & ~i_10_296_1549_0 & ~i_10_296_1578_0 & ~i_10_296_3681_0) | (~i_10_296_1822_0 & ~i_10_296_2604_0 & i_10_296_3853_0))) | (~i_10_296_2196_0 & ((~i_10_296_957_0 & ((~i_10_296_1263_0 & ~i_10_296_1539_0 & ~i_10_296_2197_0 & ~i_10_296_2199_0 & ~i_10_296_2376_0 & ~i_10_296_2630_0 & ~i_10_296_2673_0 & ~i_10_296_3046_0) | (i_10_296_2917_0 & ~i_10_296_3681_0 & ~i_10_296_4123_0))) | (i_10_296_1306_0 & ~i_10_296_2199_0) | (~i_10_296_999_0 & ~i_10_296_1083_0 & ~i_10_296_1578_0 & ~i_10_296_2502_0 & ~i_10_296_2629_0 & ~i_10_296_3978_0 & ~i_10_296_4275_0))) | (~i_10_296_4122_0 & ((~i_10_296_1822_0 & ((~i_10_296_1549_0 & ~i_10_296_2662_0 & ~i_10_296_4123_0) | (~i_10_296_2376_0 & i_10_296_2630_0 & ~i_10_296_4275_0))) | (i_10_296_516_0 & ~i_10_296_1080_0 & ~i_10_296_2376_0 & ~i_10_296_4167_0 & ~i_10_296_4269_0 & ~i_10_296_4275_0))) | (~i_10_296_2701_0 & ((~i_10_296_1549_0 & ~i_10_296_3844_0 & ~i_10_296_3978_0 & ~i_10_296_4167_0) | (~i_10_296_2700_0 & ~i_10_296_4168_0))) | (~i_10_296_1549_0 & ((i_10_296_285_0 & ~i_10_296_999_0 & ~i_10_296_2376_0 & ~i_10_296_2502_0 & i_10_296_2882_0) | (~i_10_296_2882_0 & i_10_296_3046_0 & ~i_10_296_3785_0 & ~i_10_296_4167_0 & ~i_10_296_4275_0))) | (i_10_296_967_0 & ~i_10_296_3681_0 & i_10_296_3844_0) | (i_10_296_1653_0 & i_10_296_2629_0 & i_10_296_2979_0 & ~i_10_296_3978_0 & ~i_10_296_3979_0) | (i_10_296_3616_0 & ~i_10_296_3781_0 & ~i_10_296_4168_0) | (~i_10_296_1083_0 & ~i_10_296_2016_0 & ~i_10_296_4266_0 & ~i_10_296_4275_0));
endmodule



// Benchmark "kernel_10_297" written by ABC on Sun Jul 19 10:26:10 2020

module kernel_10_297 ( 
    i_10_297_175_0, i_10_297_283_0, i_10_297_287_0, i_10_297_390_0,
    i_10_297_426_0, i_10_297_429_0, i_10_297_430_0, i_10_297_467_0,
    i_10_297_506_0, i_10_297_516_0, i_10_297_518_0, i_10_297_519_0,
    i_10_297_714_0, i_10_297_735_0, i_10_297_799_0, i_10_297_958_0,
    i_10_297_967_0, i_10_297_1000_0, i_10_297_1002_0, i_10_297_1263_0,
    i_10_297_1264_0, i_10_297_1309_0, i_10_297_1492_0, i_10_297_1552_0,
    i_10_297_1554_0, i_10_297_1578_0, i_10_297_1635_0, i_10_297_1651_0,
    i_10_297_1690_0, i_10_297_1695_0, i_10_297_1820_0, i_10_297_1823_0,
    i_10_297_1824_0, i_10_297_1875_0, i_10_297_1913_0, i_10_297_1938_0,
    i_10_297_1995_0, i_10_297_2184_0, i_10_297_2253_0, i_10_297_2310_0,
    i_10_297_2311_0, i_10_297_2329_0, i_10_297_2352_0, i_10_297_2452_0,
    i_10_297_2453_0, i_10_297_2467_0, i_10_297_2481_0, i_10_297_2508_0,
    i_10_297_2541_0, i_10_297_2628_0, i_10_297_2629_0, i_10_297_2630_0,
    i_10_297_2676_0, i_10_297_2679_0, i_10_297_2680_0, i_10_297_2708_0,
    i_10_297_2710_0, i_10_297_2715_0, i_10_297_2716_0, i_10_297_2824_0,
    i_10_297_2833_0, i_10_297_2919_0, i_10_297_3038_0, i_10_297_3041_0,
    i_10_297_3237_0, i_10_297_3315_0, i_10_297_3318_0, i_10_297_3321_0,
    i_10_297_3322_0, i_10_297_3325_0, i_10_297_3326_0, i_10_297_3388_0,
    i_10_297_3471_0, i_10_297_3495_0, i_10_297_3496_0, i_10_297_3504_0,
    i_10_297_3525_0, i_10_297_3541_0, i_10_297_3586_0, i_10_297_3588_0,
    i_10_297_3611_0, i_10_297_3648_0, i_10_297_3652_0, i_10_297_3782_0,
    i_10_297_3783_0, i_10_297_3784_0, i_10_297_3786_0, i_10_297_3836_0,
    i_10_297_3840_0, i_10_297_3848_0, i_10_297_3853_0, i_10_297_3859_0,
    i_10_297_3948_0, i_10_297_3949_0, i_10_297_3985_0, i_10_297_4057_0,
    i_10_297_4270_0, i_10_297_4272_0, i_10_297_4287_0, i_10_297_4291_0,
    o_10_297_0_0  );
  input  i_10_297_175_0, i_10_297_283_0, i_10_297_287_0, i_10_297_390_0,
    i_10_297_426_0, i_10_297_429_0, i_10_297_430_0, i_10_297_467_0,
    i_10_297_506_0, i_10_297_516_0, i_10_297_518_0, i_10_297_519_0,
    i_10_297_714_0, i_10_297_735_0, i_10_297_799_0, i_10_297_958_0,
    i_10_297_967_0, i_10_297_1000_0, i_10_297_1002_0, i_10_297_1263_0,
    i_10_297_1264_0, i_10_297_1309_0, i_10_297_1492_0, i_10_297_1552_0,
    i_10_297_1554_0, i_10_297_1578_0, i_10_297_1635_0, i_10_297_1651_0,
    i_10_297_1690_0, i_10_297_1695_0, i_10_297_1820_0, i_10_297_1823_0,
    i_10_297_1824_0, i_10_297_1875_0, i_10_297_1913_0, i_10_297_1938_0,
    i_10_297_1995_0, i_10_297_2184_0, i_10_297_2253_0, i_10_297_2310_0,
    i_10_297_2311_0, i_10_297_2329_0, i_10_297_2352_0, i_10_297_2452_0,
    i_10_297_2453_0, i_10_297_2467_0, i_10_297_2481_0, i_10_297_2508_0,
    i_10_297_2541_0, i_10_297_2628_0, i_10_297_2629_0, i_10_297_2630_0,
    i_10_297_2676_0, i_10_297_2679_0, i_10_297_2680_0, i_10_297_2708_0,
    i_10_297_2710_0, i_10_297_2715_0, i_10_297_2716_0, i_10_297_2824_0,
    i_10_297_2833_0, i_10_297_2919_0, i_10_297_3038_0, i_10_297_3041_0,
    i_10_297_3237_0, i_10_297_3315_0, i_10_297_3318_0, i_10_297_3321_0,
    i_10_297_3322_0, i_10_297_3325_0, i_10_297_3326_0, i_10_297_3388_0,
    i_10_297_3471_0, i_10_297_3495_0, i_10_297_3496_0, i_10_297_3504_0,
    i_10_297_3525_0, i_10_297_3541_0, i_10_297_3586_0, i_10_297_3588_0,
    i_10_297_3611_0, i_10_297_3648_0, i_10_297_3652_0, i_10_297_3782_0,
    i_10_297_3783_0, i_10_297_3784_0, i_10_297_3786_0, i_10_297_3836_0,
    i_10_297_3840_0, i_10_297_3848_0, i_10_297_3853_0, i_10_297_3859_0,
    i_10_297_3948_0, i_10_297_3949_0, i_10_297_3985_0, i_10_297_4057_0,
    i_10_297_4270_0, i_10_297_4272_0, i_10_297_4287_0, i_10_297_4291_0;
  output o_10_297_0_0;
  assign o_10_297_0_0 = ~((~i_10_297_426_0 & ((~i_10_297_2481_0 & ~i_10_297_2680_0 & ~i_10_297_3495_0 & ~i_10_297_3504_0) | (~i_10_297_519_0 & ~i_10_297_1264_0 & ~i_10_297_2508_0 & i_10_297_2715_0 & ~i_10_297_3315_0 & ~i_10_297_3948_0))) | (i_10_297_1820_0 & ((~i_10_297_516_0 & ~i_10_297_2716_0) | (~i_10_297_3237_0 & i_10_297_3504_0 & i_10_297_3588_0 & ~i_10_297_3848_0 & ~i_10_297_3949_0))) | (i_10_297_1824_0 & ((~i_10_297_390_0 & ~i_10_297_2679_0 & ~i_10_297_3948_0) | (i_10_297_3388_0 & i_10_297_3853_0 & i_10_297_4287_0))) | (~i_10_297_1824_0 & ((~i_10_297_1000_0 & i_10_297_3541_0 & ~i_10_297_3985_0) | (~i_10_297_2311_0 & ~i_10_297_2676_0 & ~i_10_297_3318_0 & ~i_10_297_3948_0 & ~i_10_297_4287_0))) | (~i_10_297_2481_0 & ((~i_10_297_714_0 & ~i_10_297_2467_0 & ~i_10_297_3237_0 & ~i_10_297_3496_0 & ~i_10_297_3541_0) | (~i_10_297_2329_0 & ~i_10_297_3495_0 & ~i_10_297_3948_0 & ~i_10_297_4272_0))) | (~i_10_297_2329_0 & (~i_10_297_4287_0 | (~i_10_297_2710_0 & i_10_297_3541_0))) | (~i_10_297_2508_0 & ((~i_10_297_2716_0 & ~i_10_297_3496_0 & ~i_10_297_3504_0 & ~i_10_297_3948_0) | (~i_10_297_1578_0 & ~i_10_297_1823_0 & ~i_10_297_2715_0 & ~i_10_297_3495_0 & ~i_10_297_3949_0))) | (~i_10_297_1651_0 & ~i_10_297_2310_0 & ~i_10_297_2352_0 & ~i_10_297_3496_0 & ~i_10_297_3586_0) | (~i_10_297_1264_0 & ~i_10_297_2708_0 & i_10_297_2710_0 & ~i_10_297_2833_0 & ~i_10_297_3948_0 & ~i_10_297_4270_0));
endmodule



// Benchmark "kernel_10_298" written by ABC on Sun Jul 19 10:26:11 2020

module kernel_10_298 ( 
    i_10_298_118_0, i_10_298_217_0, i_10_298_221_0, i_10_298_279_0,
    i_10_298_280_0, i_10_298_281_0, i_10_298_284_0, i_10_298_329_0,
    i_10_298_389_0, i_10_298_410_0, i_10_298_463_0, i_10_298_711_0,
    i_10_298_712_0, i_10_298_748_0, i_10_298_749_0, i_10_298_794_0,
    i_10_298_796_0, i_10_298_990_0, i_10_298_999_0, i_10_298_1000_0,
    i_10_298_1086_0, i_10_298_1234_0, i_10_298_1237_0, i_10_298_1246_0,
    i_10_298_1308_0, i_10_298_1309_0, i_10_298_1310_0, i_10_298_1359_0,
    i_10_298_1541_0, i_10_298_1577_0, i_10_298_1613_0, i_10_298_1647_0,
    i_10_298_1648_0, i_10_298_1649_0, i_10_298_1651_0, i_10_298_1654_0,
    i_10_298_1655_0, i_10_298_1684_0, i_10_298_1687_0, i_10_298_1820_0,
    i_10_298_1911_0, i_10_298_1912_0, i_10_298_1913_0, i_10_298_1916_0,
    i_10_298_1949_0, i_10_298_2352_0, i_10_298_2353_0, i_10_298_2354_0,
    i_10_298_2358_0, i_10_298_2359_0, i_10_298_2361_0, i_10_298_2449_0,
    i_10_298_2455_0, i_10_298_2630_0, i_10_298_2633_0, i_10_298_2635_0,
    i_10_298_2659_0, i_10_298_2660_0, i_10_298_2718_0, i_10_298_2721_0,
    i_10_298_2722_0, i_10_298_2723_0, i_10_298_2727_0, i_10_298_2729_0,
    i_10_298_2817_0, i_10_298_2818_0, i_10_298_2919_0, i_10_298_2920_0,
    i_10_298_2921_0, i_10_298_2980_0, i_10_298_3034_0, i_10_298_3035_0,
    i_10_298_3038_0, i_10_298_3042_0, i_10_298_3043_0, i_10_298_3157_0,
    i_10_298_3277_0, i_10_298_3278_0, i_10_298_3279_0, i_10_298_3388_0,
    i_10_298_3466_0, i_10_298_3523_0, i_10_298_3556_0, i_10_298_3613_0,
    i_10_298_3645_0, i_10_298_3834_0, i_10_298_3840_0, i_10_298_3846_0,
    i_10_298_3857_0, i_10_298_3906_0, i_10_298_3907_0, i_10_298_3908_0,
    i_10_298_3979_0, i_10_298_4051_0, i_10_298_4113_0, i_10_298_4114_0,
    i_10_298_4118_0, i_10_298_4271_0, i_10_298_4288_0, i_10_298_4289_0,
    o_10_298_0_0  );
  input  i_10_298_118_0, i_10_298_217_0, i_10_298_221_0, i_10_298_279_0,
    i_10_298_280_0, i_10_298_281_0, i_10_298_284_0, i_10_298_329_0,
    i_10_298_389_0, i_10_298_410_0, i_10_298_463_0, i_10_298_711_0,
    i_10_298_712_0, i_10_298_748_0, i_10_298_749_0, i_10_298_794_0,
    i_10_298_796_0, i_10_298_990_0, i_10_298_999_0, i_10_298_1000_0,
    i_10_298_1086_0, i_10_298_1234_0, i_10_298_1237_0, i_10_298_1246_0,
    i_10_298_1308_0, i_10_298_1309_0, i_10_298_1310_0, i_10_298_1359_0,
    i_10_298_1541_0, i_10_298_1577_0, i_10_298_1613_0, i_10_298_1647_0,
    i_10_298_1648_0, i_10_298_1649_0, i_10_298_1651_0, i_10_298_1654_0,
    i_10_298_1655_0, i_10_298_1684_0, i_10_298_1687_0, i_10_298_1820_0,
    i_10_298_1911_0, i_10_298_1912_0, i_10_298_1913_0, i_10_298_1916_0,
    i_10_298_1949_0, i_10_298_2352_0, i_10_298_2353_0, i_10_298_2354_0,
    i_10_298_2358_0, i_10_298_2359_0, i_10_298_2361_0, i_10_298_2449_0,
    i_10_298_2455_0, i_10_298_2630_0, i_10_298_2633_0, i_10_298_2635_0,
    i_10_298_2659_0, i_10_298_2660_0, i_10_298_2718_0, i_10_298_2721_0,
    i_10_298_2722_0, i_10_298_2723_0, i_10_298_2727_0, i_10_298_2729_0,
    i_10_298_2817_0, i_10_298_2818_0, i_10_298_2919_0, i_10_298_2920_0,
    i_10_298_2921_0, i_10_298_2980_0, i_10_298_3034_0, i_10_298_3035_0,
    i_10_298_3038_0, i_10_298_3042_0, i_10_298_3043_0, i_10_298_3157_0,
    i_10_298_3277_0, i_10_298_3278_0, i_10_298_3279_0, i_10_298_3388_0,
    i_10_298_3466_0, i_10_298_3523_0, i_10_298_3556_0, i_10_298_3613_0,
    i_10_298_3645_0, i_10_298_3834_0, i_10_298_3840_0, i_10_298_3846_0,
    i_10_298_3857_0, i_10_298_3906_0, i_10_298_3907_0, i_10_298_3908_0,
    i_10_298_3979_0, i_10_298_4051_0, i_10_298_4113_0, i_10_298_4114_0,
    i_10_298_4118_0, i_10_298_4271_0, i_10_298_4288_0, i_10_298_4289_0;
  output o_10_298_0_0;
  assign o_10_298_0_0 = ~((~i_10_298_796_0 & ((~i_10_298_1647_0 & ~i_10_298_1911_0 & ~i_10_298_2721_0 & ~i_10_298_2723_0 & ~i_10_298_2980_0) | (~i_10_298_410_0 & ~i_10_298_748_0 & ~i_10_298_1916_0 & ~i_10_298_2352_0 & ~i_10_298_2729_0 & ~i_10_298_3523_0 & ~i_10_298_3840_0 & ~i_10_298_3908_0 & ~i_10_298_4289_0))) | (~i_10_298_1912_0 & ((~i_10_298_749_0 & ((~i_10_298_711_0 & ~i_10_298_990_0 & ~i_10_298_1913_0 & ~i_10_298_1916_0 & ~i_10_298_2354_0) | (~i_10_298_1237_0 & ~i_10_298_2660_0 & ~i_10_298_2721_0 & ~i_10_298_3034_0 & i_10_298_3613_0 & ~i_10_298_4271_0))) | (i_10_298_4118_0 & ((~i_10_298_217_0 & ~i_10_298_794_0 & ~i_10_298_990_0 & ~i_10_298_1911_0 & ~i_10_298_2718_0 & ~i_10_298_2818_0) | (i_10_298_281_0 & ~i_10_298_748_0 & ~i_10_298_2455_0 & i_10_298_2660_0 & ~i_10_298_2920_0))))) | (~i_10_298_711_0 & ((~i_10_298_1911_0 & ~i_10_298_2718_0 & i_10_298_3035_0) | (~i_10_298_712_0 & ~i_10_298_749_0 & ~i_10_298_1309_0 & ~i_10_298_1310_0 & ~i_10_298_3906_0))) | (i_10_298_1654_0 & ((~i_10_298_1310_0 & ~i_10_298_2718_0 & ~i_10_298_2722_0 & ~i_10_298_2817_0 & ~i_10_298_3034_0) | (~i_10_298_329_0 & ~i_10_298_1684_0 & i_10_298_2723_0 & ~i_10_298_3613_0 & ~i_10_298_3906_0))) | (i_10_298_1687_0 & ((~i_10_298_284_0 & ~i_10_298_463_0 & ~i_10_298_2723_0) | (~i_10_298_410_0 & ~i_10_298_748_0 & ~i_10_298_1916_0 & ~i_10_298_2817_0 & i_10_298_2919_0 & ~i_10_298_3834_0))) | (~i_10_298_410_0 & ((~i_10_298_748_0 & ~i_10_298_1916_0 & ~i_10_298_1949_0 & ~i_10_298_2354_0 & ~i_10_298_2455_0 & i_10_298_2635_0) | (i_10_298_280_0 & i_10_298_2659_0 & ~i_10_298_3279_0 & i_10_298_3388_0))) | (~i_10_298_748_0 & ((~i_10_298_1246_0 & ~i_10_298_2455_0 & ~i_10_298_2659_0 & ~i_10_298_2818_0 & ~i_10_298_3388_0 & ~i_10_298_3857_0) | (~i_10_298_749_0 & ~i_10_298_1086_0 & ~i_10_298_1308_0 & ~i_10_298_2919_0 & ~i_10_298_4051_0 & i_10_298_4288_0))) | (~i_10_298_1246_0 & ~i_10_298_3388_0 & ((~i_10_298_1916_0 & i_10_298_2635_0 & ~i_10_298_2659_0 & i_10_298_2723_0 & ~i_10_298_2919_0) | (~i_10_298_2723_0 & ~i_10_298_3278_0 & ~i_10_298_3279_0 & i_10_298_3613_0 & ~i_10_298_3834_0 & ~i_10_298_3840_0 & ~i_10_298_3906_0 & ~i_10_298_4271_0))) | (~i_10_298_2659_0 & ((i_10_298_796_0 & i_10_298_2635_0 & ~i_10_298_3840_0 & ~i_10_298_3857_0) | (i_10_298_794_0 & ~i_10_298_4114_0))) | (~i_10_298_2722_0 & ((~i_10_298_1913_0 & ~i_10_298_2718_0 & ~i_10_298_2980_0 & i_10_298_3038_0) | (i_10_298_329_0 & ~i_10_298_4114_0))) | (~i_10_298_1655_0 & i_10_298_2359_0 & ~i_10_298_2729_0) | (i_10_298_1577_0 & ~i_10_298_2353_0 & i_10_298_3613_0 & i_10_298_3834_0));
endmodule



// Benchmark "kernel_10_299" written by ABC on Sun Jul 19 10:26:13 2020

module kernel_10_299 ( 
    i_10_299_175_0, i_10_299_221_0, i_10_299_280_0, i_10_299_285_0,
    i_10_299_286_0, i_10_299_390_0, i_10_299_465_0, i_10_299_466_0,
    i_10_299_753_0, i_10_299_796_0, i_10_299_957_0, i_10_299_967_0,
    i_10_299_1032_0, i_10_299_1035_0, i_10_299_1236_0, i_10_299_1237_0,
    i_10_299_1239_0, i_10_299_1240_0, i_10_299_1242_0, i_10_299_1243_0,
    i_10_299_1248_0, i_10_299_1249_0, i_10_299_1263_0, i_10_299_1341_0,
    i_10_299_1359_0, i_10_299_1444_0, i_10_299_1545_0, i_10_299_1555_0,
    i_10_299_1576_0, i_10_299_1647_0, i_10_299_1650_0, i_10_299_1651_0,
    i_10_299_1683_0, i_10_299_1812_0, i_10_299_1819_0, i_10_299_1913_0,
    i_10_299_1915_0, i_10_299_1945_0, i_10_299_2185_0, i_10_299_2197_0,
    i_10_299_2199_0, i_10_299_2352_0, i_10_299_2353_0, i_10_299_2361_0,
    i_10_299_2449_0, i_10_299_2456_0, i_10_299_2467_0, i_10_299_2471_0,
    i_10_299_2601_0, i_10_299_2602_0, i_10_299_2604_0, i_10_299_2607_0,
    i_10_299_2628_0, i_10_299_2629_0, i_10_299_2634_0, i_10_299_2636_0,
    i_10_299_2659_0, i_10_299_2662_0, i_10_299_2700_0, i_10_299_2709_0,
    i_10_299_2731_0, i_10_299_2827_0, i_10_299_2830_0, i_10_299_2833_0,
    i_10_299_2981_0, i_10_299_3033_0, i_10_299_3034_0, i_10_299_3036_0,
    i_10_299_3037_0, i_10_299_3329_0, i_10_299_3389_0, i_10_299_3466_0,
    i_10_299_3549_0, i_10_299_3583_0, i_10_299_3586_0, i_10_299_3624_0,
    i_10_299_3645_0, i_10_299_3646_0, i_10_299_3647_0, i_10_299_3648_0,
    i_10_299_3649_0, i_10_299_3717_0, i_10_299_3718_0, i_10_299_3840_0,
    i_10_299_3843_0, i_10_299_3847_0, i_10_299_3848_0, i_10_299_3850_0,
    i_10_299_3852_0, i_10_299_3860_0, i_10_299_3870_0, i_10_299_3888_0,
    i_10_299_3982_0, i_10_299_4116_0, i_10_299_4117_0, i_10_299_4217_0,
    i_10_299_4275_0, i_10_299_4276_0, i_10_299_4564_0, i_10_299_4566_0,
    o_10_299_0_0  );
  input  i_10_299_175_0, i_10_299_221_0, i_10_299_280_0, i_10_299_285_0,
    i_10_299_286_0, i_10_299_390_0, i_10_299_465_0, i_10_299_466_0,
    i_10_299_753_0, i_10_299_796_0, i_10_299_957_0, i_10_299_967_0,
    i_10_299_1032_0, i_10_299_1035_0, i_10_299_1236_0, i_10_299_1237_0,
    i_10_299_1239_0, i_10_299_1240_0, i_10_299_1242_0, i_10_299_1243_0,
    i_10_299_1248_0, i_10_299_1249_0, i_10_299_1263_0, i_10_299_1341_0,
    i_10_299_1359_0, i_10_299_1444_0, i_10_299_1545_0, i_10_299_1555_0,
    i_10_299_1576_0, i_10_299_1647_0, i_10_299_1650_0, i_10_299_1651_0,
    i_10_299_1683_0, i_10_299_1812_0, i_10_299_1819_0, i_10_299_1913_0,
    i_10_299_1915_0, i_10_299_1945_0, i_10_299_2185_0, i_10_299_2197_0,
    i_10_299_2199_0, i_10_299_2352_0, i_10_299_2353_0, i_10_299_2361_0,
    i_10_299_2449_0, i_10_299_2456_0, i_10_299_2467_0, i_10_299_2471_0,
    i_10_299_2601_0, i_10_299_2602_0, i_10_299_2604_0, i_10_299_2607_0,
    i_10_299_2628_0, i_10_299_2629_0, i_10_299_2634_0, i_10_299_2636_0,
    i_10_299_2659_0, i_10_299_2662_0, i_10_299_2700_0, i_10_299_2709_0,
    i_10_299_2731_0, i_10_299_2827_0, i_10_299_2830_0, i_10_299_2833_0,
    i_10_299_2981_0, i_10_299_3033_0, i_10_299_3034_0, i_10_299_3036_0,
    i_10_299_3037_0, i_10_299_3329_0, i_10_299_3389_0, i_10_299_3466_0,
    i_10_299_3549_0, i_10_299_3583_0, i_10_299_3586_0, i_10_299_3624_0,
    i_10_299_3645_0, i_10_299_3646_0, i_10_299_3647_0, i_10_299_3648_0,
    i_10_299_3649_0, i_10_299_3717_0, i_10_299_3718_0, i_10_299_3840_0,
    i_10_299_3843_0, i_10_299_3847_0, i_10_299_3848_0, i_10_299_3850_0,
    i_10_299_3852_0, i_10_299_3860_0, i_10_299_3870_0, i_10_299_3888_0,
    i_10_299_3982_0, i_10_299_4116_0, i_10_299_4117_0, i_10_299_4217_0,
    i_10_299_4275_0, i_10_299_4276_0, i_10_299_4564_0, i_10_299_4566_0;
  output o_10_299_0_0;
  assign o_10_299_0_0 = ~((~i_10_299_286_0 & ((i_10_299_2361_0 & ~i_10_299_2601_0 & ~i_10_299_2607_0 & ~i_10_299_2659_0 & ~i_10_299_3036_0) | (~i_10_299_957_0 & ~i_10_299_967_0 & ~i_10_299_1545_0 & ~i_10_299_1683_0 & ~i_10_299_2602_0 & ~i_10_299_3888_0))) | (~i_10_299_2601_0 & ((~i_10_299_1263_0 & ((~i_10_299_957_0 & ~i_10_299_1035_0 & ~i_10_299_2602_0 & ~i_10_299_3036_0) | (~i_10_299_796_0 & ~i_10_299_967_0 & ~i_10_299_1242_0 & ~i_10_299_2361_0 & ~i_10_299_4566_0))) | (~i_10_299_1236_0 & ~i_10_299_1647_0 & i_10_299_1819_0 & ~i_10_299_2456_0 & ~i_10_299_2830_0) | (~i_10_299_1576_0 & ~i_10_299_3847_0 & ~i_10_299_3888_0))) | (~i_10_299_796_0 & ((~i_10_299_1035_0 & ~i_10_299_1243_0 & ~i_10_299_1248_0 & ~i_10_299_1819_0 & ~i_10_299_2353_0) | (~i_10_299_465_0 & ~i_10_299_1545_0 & i_10_299_3850_0 & ~i_10_299_3888_0))) | (~i_10_299_1035_0 & ((~i_10_299_1243_0 & i_10_299_2629_0 & ~i_10_299_3648_0) | (~i_10_299_221_0 & ~i_10_299_2197_0 & ~i_10_299_2352_0 & ~i_10_299_3037_0 & ~i_10_299_3843_0))) | (~i_10_299_1243_0 & ((~i_10_299_1647_0 & ~i_10_299_1650_0 & ~i_10_299_3852_0 & ~i_10_299_3888_0) | (~i_10_299_2361_0 & ~i_10_299_2602_0 & ~i_10_299_3847_0 & ~i_10_299_4275_0))) | (~i_10_299_2197_0 & ((~i_10_299_1545_0 & ~i_10_299_1812_0 & ~i_10_299_1915_0 & ~i_10_299_3033_0 & ~i_10_299_3645_0) | (~i_10_299_1032_0 & i_10_299_3982_0))) | (~i_10_299_3033_0 & ((i_10_299_2449_0 & ~i_10_299_2602_0 & ~i_10_299_3847_0 & ~i_10_299_3848_0) | (~i_10_299_1576_0 & ~i_10_299_2700_0 & ~i_10_299_3850_0 & i_10_299_4117_0))) | (i_10_299_2731_0 & ~i_10_299_3888_0 & ~i_10_299_4117_0));
endmodule



// Benchmark "kernel_10_300" written by ABC on Sun Jul 19 10:26:14 2020

module kernel_10_300 ( 
    i_10_300_171_0, i_10_300_172_0, i_10_300_175_0, i_10_300_222_0,
    i_10_300_244_0, i_10_300_279_0, i_10_300_283_0, i_10_300_328_0,
    i_10_300_409_0, i_10_300_436_0, i_10_300_441_0, i_10_300_442_0,
    i_10_300_443_0, i_10_300_462_0, i_10_300_696_0, i_10_300_748_0,
    i_10_300_990_0, i_10_300_991_0, i_10_300_1026_0, i_10_300_1029_0,
    i_10_300_1233_0, i_10_300_1234_0, i_10_300_1238_0, i_10_300_1262_0,
    i_10_300_1265_0, i_10_300_1308_0, i_10_300_1309_0, i_10_300_1310_0,
    i_10_300_1445_0, i_10_300_1539_0, i_10_300_1540_0, i_10_300_1541_0,
    i_10_300_1575_0, i_10_300_1576_0, i_10_300_1651_0, i_10_300_1819_0,
    i_10_300_1822_0, i_10_300_1911_0, i_10_300_1912_0, i_10_300_1944_0,
    i_10_300_2179_0, i_10_300_2180_0, i_10_300_2197_0, i_10_300_2198_0,
    i_10_300_2201_0, i_10_300_2351_0, i_10_300_2450_0, i_10_300_2453_0,
    i_10_300_2468_0, i_10_300_2469_0, i_10_300_2470_0, i_10_300_2471_0,
    i_10_300_2629_0, i_10_300_2630_0, i_10_300_2633_0, i_10_300_2636_0,
    i_10_300_2661_0, i_10_300_2702_0, i_10_300_2817_0, i_10_300_2820_0,
    i_10_300_2827_0, i_10_300_2830_0, i_10_300_2881_0, i_10_300_2882_0,
    i_10_300_2884_0, i_10_300_2885_0, i_10_300_2888_0, i_10_300_3071_0,
    i_10_300_3078_0, i_10_300_3196_0, i_10_300_3198_0, i_10_300_3199_0,
    i_10_300_3200_0, i_10_300_3202_0, i_10_300_3203_0, i_10_300_3391_0,
    i_10_300_3403_0, i_10_300_3583_0, i_10_300_3586_0, i_10_300_3611_0,
    i_10_300_3613_0, i_10_300_3614_0, i_10_300_3645_0, i_10_300_3788_0,
    i_10_300_3834_0, i_10_300_3839_0, i_10_300_3846_0, i_10_300_3851_0,
    i_10_300_3853_0, i_10_300_3854_0, i_10_300_3888_0, i_10_300_3994_0,
    i_10_300_4113_0, i_10_300_4114_0, i_10_300_4116_0, i_10_300_4129_0,
    i_10_300_4278_0, i_10_300_4291_0, i_10_300_4292_0, i_10_300_4457_0,
    o_10_300_0_0  );
  input  i_10_300_171_0, i_10_300_172_0, i_10_300_175_0, i_10_300_222_0,
    i_10_300_244_0, i_10_300_279_0, i_10_300_283_0, i_10_300_328_0,
    i_10_300_409_0, i_10_300_436_0, i_10_300_441_0, i_10_300_442_0,
    i_10_300_443_0, i_10_300_462_0, i_10_300_696_0, i_10_300_748_0,
    i_10_300_990_0, i_10_300_991_0, i_10_300_1026_0, i_10_300_1029_0,
    i_10_300_1233_0, i_10_300_1234_0, i_10_300_1238_0, i_10_300_1262_0,
    i_10_300_1265_0, i_10_300_1308_0, i_10_300_1309_0, i_10_300_1310_0,
    i_10_300_1445_0, i_10_300_1539_0, i_10_300_1540_0, i_10_300_1541_0,
    i_10_300_1575_0, i_10_300_1576_0, i_10_300_1651_0, i_10_300_1819_0,
    i_10_300_1822_0, i_10_300_1911_0, i_10_300_1912_0, i_10_300_1944_0,
    i_10_300_2179_0, i_10_300_2180_0, i_10_300_2197_0, i_10_300_2198_0,
    i_10_300_2201_0, i_10_300_2351_0, i_10_300_2450_0, i_10_300_2453_0,
    i_10_300_2468_0, i_10_300_2469_0, i_10_300_2470_0, i_10_300_2471_0,
    i_10_300_2629_0, i_10_300_2630_0, i_10_300_2633_0, i_10_300_2636_0,
    i_10_300_2661_0, i_10_300_2702_0, i_10_300_2817_0, i_10_300_2820_0,
    i_10_300_2827_0, i_10_300_2830_0, i_10_300_2881_0, i_10_300_2882_0,
    i_10_300_2884_0, i_10_300_2885_0, i_10_300_2888_0, i_10_300_3071_0,
    i_10_300_3078_0, i_10_300_3196_0, i_10_300_3198_0, i_10_300_3199_0,
    i_10_300_3200_0, i_10_300_3202_0, i_10_300_3203_0, i_10_300_3391_0,
    i_10_300_3403_0, i_10_300_3583_0, i_10_300_3586_0, i_10_300_3611_0,
    i_10_300_3613_0, i_10_300_3614_0, i_10_300_3645_0, i_10_300_3788_0,
    i_10_300_3834_0, i_10_300_3839_0, i_10_300_3846_0, i_10_300_3851_0,
    i_10_300_3853_0, i_10_300_3854_0, i_10_300_3888_0, i_10_300_3994_0,
    i_10_300_4113_0, i_10_300_4114_0, i_10_300_4116_0, i_10_300_4129_0,
    i_10_300_4278_0, i_10_300_4291_0, i_10_300_4292_0, i_10_300_4457_0;
  output o_10_300_0_0;
  assign o_10_300_0_0 = ~((i_10_300_442_0 & ((~i_10_300_748_0 & ~i_10_300_991_0 & ~i_10_300_3614_0) | (~i_10_300_244_0 & ~i_10_300_696_0 & ~i_10_300_1029_0 & ~i_10_300_2884_0 & ~i_10_300_2888_0 & ~i_10_300_3851_0))) | (~i_10_300_2888_0 & ((~i_10_300_696_0 & ~i_10_300_4129_0 & ((~i_10_300_1234_0 & ~i_10_300_1309_0 & ~i_10_300_1310_0 & ~i_10_300_1541_0 & ~i_10_300_1575_0 & ~i_10_300_3203_0 & ~i_10_300_3391_0 & ~i_10_300_3403_0) | (~i_10_300_328_0 & ~i_10_300_991_0 & ~i_10_300_1539_0 & ~i_10_300_1576_0 & ~i_10_300_2201_0 & ~i_10_300_2827_0 & ~i_10_300_3839_0 & ~i_10_300_3994_0))) | (~i_10_300_1576_0 & ~i_10_300_3614_0 & ((~i_10_300_462_0 & ~i_10_300_748_0 & ~i_10_300_1540_0 & ~i_10_300_1911_0 & ~i_10_300_2197_0 & ~i_10_300_2468_0 & ~i_10_300_2820_0 & ~i_10_300_2882_0 & ~i_10_300_3888_0) | (~i_10_300_409_0 & ~i_10_300_990_0 & ~i_10_300_1541_0 & ~i_10_300_2630_0 & ~i_10_300_3611_0 & ~i_10_300_3613_0 & ~i_10_300_4278_0))) | (~i_10_300_3199_0 & ~i_10_300_3203_0 & i_10_300_3583_0 & i_10_300_3586_0 & ~i_10_300_3613_0))) | (~i_10_300_3203_0 & ((~i_10_300_328_0 & ((~i_10_300_171_0 & ~i_10_300_1540_0 & i_10_300_1819_0 & ~i_10_300_1822_0 & ~i_10_300_2453_0 & ~i_10_300_2884_0 & ~i_10_300_3613_0) | (~i_10_300_283_0 & ~i_10_300_409_0 & ~i_10_300_748_0 & ~i_10_300_1262_0 & ~i_10_300_1310_0 & ~i_10_300_2636_0 & ~i_10_300_2817_0 & ~i_10_300_3071_0 & ~i_10_300_3200_0 & ~i_10_300_3614_0 & ~i_10_300_3888_0))) | (~i_10_300_2885_0 & ((~i_10_300_409_0 & ~i_10_300_462_0 & i_10_300_1822_0 & ~i_10_300_2197_0 & ~i_10_300_2453_0 & ~i_10_300_3196_0 & ~i_10_300_3202_0 & ~i_10_300_3391_0) | (~i_10_300_2201_0 & i_10_300_2636_0 & ~i_10_300_2830_0 & ~i_10_300_2884_0 & i_10_300_3586_0))) | (~i_10_300_4291_0 & ((~i_10_300_244_0 & i_10_300_283_0 & ~i_10_300_436_0 & ~i_10_300_1262_0 & ~i_10_300_2180_0 & ~i_10_300_2450_0 & ~i_10_300_3196_0 & ~i_10_300_3200_0 & ~i_10_300_3611_0 & ~i_10_300_3888_0) | (~i_10_300_748_0 & ~i_10_300_1575_0 & i_10_300_1651_0 & ~i_10_300_2661_0 & ~i_10_300_2827_0 & ~i_10_300_3071_0 & ~i_10_300_3198_0 & ~i_10_300_3391_0 & ~i_10_300_3994_0 & ~i_10_300_4278_0))))) | (~i_10_300_462_0 & ((~i_10_300_1262_0 & ~i_10_300_1310_0 & ~i_10_300_1540_0 & i_10_300_2827_0 & ~i_10_300_2881_0 & ~i_10_300_3391_0 & ~i_10_300_3851_0 & ~i_10_300_3888_0) | (~i_10_300_244_0 & ~i_10_300_1911_0 & ~i_10_300_2201_0 & ~i_10_300_2629_0 & ~i_10_300_2633_0 & ~i_10_300_2817_0 & ~i_10_300_3200_0 & ~i_10_300_3994_0 & ~i_10_300_4129_0 & ~i_10_300_4291_0))) | (~i_10_300_244_0 & ~i_10_300_2885_0 & ((i_10_300_1234_0 & ~i_10_300_1911_0 & ~i_10_300_2820_0 & ~i_10_300_3613_0 & ~i_10_300_3888_0 & ~i_10_300_4113_0) | (i_10_300_1238_0 & ~i_10_300_1575_0 & ~i_10_300_1912_0 & ~i_10_300_2636_0 & ~i_10_300_3198_0 & ~i_10_300_3403_0 & ~i_10_300_4292_0))) | (~i_10_300_1576_0 & ((~i_10_300_1029_0 & i_10_300_1539_0 & i_10_300_3853_0) | (~i_10_300_436_0 & ~i_10_300_1238_0 & i_10_300_1309_0 & ~i_10_300_1575_0 & ~i_10_300_2198_0 & ~i_10_300_2351_0 & ~i_10_300_2471_0 & ~i_10_300_2636_0 & ~i_10_300_3202_0 & ~i_10_300_3403_0 & i_10_300_3613_0 & ~i_10_300_4278_0))) | (~i_10_300_3994_0 & ((~i_10_300_1911_0 & ((~i_10_300_409_0 & ~i_10_300_436_0 & ~i_10_300_991_0 & ~i_10_300_1262_0 & ~i_10_300_1541_0 & ~i_10_300_2179_0 & ~i_10_300_2661_0 & ~i_10_300_2817_0 & ~i_10_300_3199_0) | (i_10_300_172_0 & i_10_300_175_0 & ~i_10_300_1265_0 & ~i_10_300_1445_0 & ~i_10_300_2197_0 & ~i_10_300_3788_0 & ~i_10_300_4129_0))) | (~i_10_300_2197_0 & ~i_10_300_2201_0 & ~i_10_300_2453_0 & ~i_10_300_3199_0 & ~i_10_300_4114_0 & ~i_10_300_4291_0))) | (~i_10_300_436_0 & ~i_10_300_2197_0 & ((~i_10_300_1539_0 & ~i_10_300_1540_0 & ~i_10_300_2198_0 & ~i_10_300_2830_0 & ~i_10_300_2884_0 & ~i_10_300_3196_0 & ~i_10_300_3200_0) | (~i_10_300_328_0 & ~i_10_300_990_0 & ~i_10_300_3071_0 & ~i_10_300_3202_0 & ~i_10_300_3614_0 & ~i_10_300_4113_0 & ~i_10_300_4292_0))) | (~i_10_300_2820_0 & i_10_300_2884_0 & ~i_10_300_3199_0 & i_10_300_3391_0 & ~i_10_300_4292_0));
endmodule



// Benchmark "kernel_10_301" written by ABC on Sun Jul 19 10:26:15 2020

module kernel_10_301 ( 
    i_10_301_44_0, i_10_301_152_0, i_10_301_171_0, i_10_301_179_0,
    i_10_301_187_0, i_10_301_188_0, i_10_301_251_0, i_10_301_327_0,
    i_10_301_329_0, i_10_301_332_0, i_10_301_394_0, i_10_301_463_0,
    i_10_301_465_0, i_10_301_518_0, i_10_301_520_0, i_10_301_521_0,
    i_10_301_565_0, i_10_301_566_0, i_10_301_638_0, i_10_301_796_0,
    i_10_301_799_0, i_10_301_800_0, i_10_301_899_0, i_10_301_908_0,
    i_10_301_959_0, i_10_301_995_0, i_10_301_998_0, i_10_301_1166_0,
    i_10_301_1204_0, i_10_301_1235_0, i_10_301_1241_0, i_10_301_1264_0,
    i_10_301_1276_0, i_10_301_1313_0, i_10_301_1653_0, i_10_301_1817_0,
    i_10_301_1826_0, i_10_301_1889_0, i_10_301_1913_0, i_10_301_1997_0,
    i_10_301_2006_0, i_10_301_2024_0, i_10_301_2032_0, i_10_301_2033_0,
    i_10_301_2041_0, i_10_301_2353_0, i_10_301_2365_0, i_10_301_2450_0,
    i_10_301_2452_0, i_10_301_2464_0, i_10_301_2468_0, i_10_301_2510_0,
    i_10_301_2515_0, i_10_301_2568_0, i_10_301_2609_0, i_10_301_2681_0,
    i_10_301_2717_0, i_10_301_2734_0, i_10_301_2830_0, i_10_301_2882_0,
    i_10_301_2885_0, i_10_301_2888_0, i_10_301_2986_0, i_10_301_3033_0,
    i_10_301_3059_0, i_10_301_3200_0, i_10_301_3239_0, i_10_301_3270_0,
    i_10_301_3280_0, i_10_301_3283_0, i_10_301_3302_0, i_10_301_3409_0,
    i_10_301_3473_0, i_10_301_3497_0, i_10_301_3509_0, i_10_301_3526_0,
    i_10_301_3552_0, i_10_301_3613_0, i_10_301_3689_0, i_10_301_3783_0,
    i_10_301_3851_0, i_10_301_3852_0, i_10_301_3859_0, i_10_301_3878_0,
    i_10_301_3913_0, i_10_301_3914_0, i_10_301_3923_0, i_10_301_3983_0,
    i_10_301_3995_0, i_10_301_4023_0, i_10_301_4168_0, i_10_301_4237_0,
    i_10_301_4271_0, i_10_301_4272_0, i_10_301_4274_0, i_10_301_4287_0,
    i_10_301_4463_0, i_10_301_4568_0, i_10_301_4569_0, i_10_301_4571_0,
    o_10_301_0_0  );
  input  i_10_301_44_0, i_10_301_152_0, i_10_301_171_0, i_10_301_179_0,
    i_10_301_187_0, i_10_301_188_0, i_10_301_251_0, i_10_301_327_0,
    i_10_301_329_0, i_10_301_332_0, i_10_301_394_0, i_10_301_463_0,
    i_10_301_465_0, i_10_301_518_0, i_10_301_520_0, i_10_301_521_0,
    i_10_301_565_0, i_10_301_566_0, i_10_301_638_0, i_10_301_796_0,
    i_10_301_799_0, i_10_301_800_0, i_10_301_899_0, i_10_301_908_0,
    i_10_301_959_0, i_10_301_995_0, i_10_301_998_0, i_10_301_1166_0,
    i_10_301_1204_0, i_10_301_1235_0, i_10_301_1241_0, i_10_301_1264_0,
    i_10_301_1276_0, i_10_301_1313_0, i_10_301_1653_0, i_10_301_1817_0,
    i_10_301_1826_0, i_10_301_1889_0, i_10_301_1913_0, i_10_301_1997_0,
    i_10_301_2006_0, i_10_301_2024_0, i_10_301_2032_0, i_10_301_2033_0,
    i_10_301_2041_0, i_10_301_2353_0, i_10_301_2365_0, i_10_301_2450_0,
    i_10_301_2452_0, i_10_301_2464_0, i_10_301_2468_0, i_10_301_2510_0,
    i_10_301_2515_0, i_10_301_2568_0, i_10_301_2609_0, i_10_301_2681_0,
    i_10_301_2717_0, i_10_301_2734_0, i_10_301_2830_0, i_10_301_2882_0,
    i_10_301_2885_0, i_10_301_2888_0, i_10_301_2986_0, i_10_301_3033_0,
    i_10_301_3059_0, i_10_301_3200_0, i_10_301_3239_0, i_10_301_3270_0,
    i_10_301_3280_0, i_10_301_3283_0, i_10_301_3302_0, i_10_301_3409_0,
    i_10_301_3473_0, i_10_301_3497_0, i_10_301_3509_0, i_10_301_3526_0,
    i_10_301_3552_0, i_10_301_3613_0, i_10_301_3689_0, i_10_301_3783_0,
    i_10_301_3851_0, i_10_301_3852_0, i_10_301_3859_0, i_10_301_3878_0,
    i_10_301_3913_0, i_10_301_3914_0, i_10_301_3923_0, i_10_301_3983_0,
    i_10_301_3995_0, i_10_301_4023_0, i_10_301_4168_0, i_10_301_4237_0,
    i_10_301_4271_0, i_10_301_4272_0, i_10_301_4274_0, i_10_301_4287_0,
    i_10_301_4463_0, i_10_301_4568_0, i_10_301_4569_0, i_10_301_4571_0;
  output o_10_301_0_0;
  assign o_10_301_0_0 = ~((~i_10_301_179_0 & ((~i_10_301_2830_0 & ~i_10_301_3509_0 & i_10_301_3995_0 & ~i_10_301_4237_0) | (~i_10_301_188_0 & ~i_10_301_899_0 & ~i_10_301_2032_0 & ~i_10_301_2681_0 & ~i_10_301_3033_0 & ~i_10_301_3270_0 & ~i_10_301_4569_0))) | (~i_10_301_332_0 & ((~i_10_301_463_0 & i_10_301_520_0 & ~i_10_301_796_0 & ~i_10_301_2033_0 & ~i_10_301_2830_0 & ~i_10_301_3851_0 & ~i_10_301_4271_0) | (~i_10_301_908_0 & ~i_10_301_2353_0 & i_10_301_2681_0 & ~i_10_301_3509_0 & ~i_10_301_4571_0))) | (~i_10_301_4237_0 & ((~i_10_301_188_0 & ((~i_10_301_908_0 & i_10_301_1826_0 & ~i_10_301_2033_0 & ~i_10_301_2681_0 & ~i_10_301_2882_0) | (~i_10_301_3851_0 & ~i_10_301_4271_0 & ~i_10_301_2024_0 & ~i_10_301_3239_0))) | (~i_10_301_1997_0 & ~i_10_301_2006_0 & ((~i_10_301_1166_0 & ~i_10_301_1264_0 & ~i_10_301_3852_0 & ~i_10_301_4271_0 & ~i_10_301_4274_0) | (~i_10_301_2033_0 & ~i_10_301_2365_0 & ~i_10_301_3200_0 & ~i_10_301_4568_0))) | (~i_10_301_908_0 & i_10_301_1826_0 & ~i_10_301_2365_0 & ~i_10_301_2717_0 & ~i_10_301_3852_0) | (~i_10_301_152_0 & ~i_10_301_899_0 & ~i_10_301_1913_0 & ~i_10_301_2024_0 & ~i_10_301_2032_0 & ~i_10_301_2450_0 & ~i_10_301_2885_0 & ~i_10_301_3689_0))) | (~i_10_301_899_0 & ((~i_10_301_187_0 & ~i_10_301_2006_0 & ~i_10_301_2986_0 & ~i_10_301_3239_0 & ~i_10_301_3283_0 & ~i_10_301_3613_0 & ~i_10_301_3689_0 & ~i_10_301_3852_0 & ~i_10_301_3995_0) | (~i_10_301_518_0 & ~i_10_301_521_0 & ~i_10_301_998_0 & ~i_10_301_2510_0 & ~i_10_301_2681_0 & ~i_10_301_3497_0 & ~i_10_301_3509_0 & ~i_10_301_4023_0 & ~i_10_301_4272_0))) | (~i_10_301_521_0 & ((~i_10_301_520_0 & ~i_10_301_1241_0 & ~i_10_301_3689_0) | (i_10_301_188_0 & ~i_10_301_1166_0 & ~i_10_301_3239_0 & i_10_301_4274_0))) | (~i_10_301_3689_0 & ~i_10_301_3914_0 & ((~i_10_301_329_0 & ~i_10_301_465_0 & i_10_301_520_0 & ~i_10_301_2885_0 & ~i_10_301_3613_0 & i_10_301_4274_0 & ~i_10_301_4287_0) | (~i_10_301_188_0 & ~i_10_301_2024_0 & ~i_10_301_3497_0 & ~i_10_301_3913_0 & ~i_10_301_4571_0))) | (~i_10_301_565_0 & i_10_301_2450_0 & i_10_301_2609_0) | (~i_10_301_799_0 & i_10_301_3200_0 & i_10_301_3239_0) | (i_10_301_1653_0 & ~i_10_301_2830_0 & ~i_10_301_3239_0 & ~i_10_301_3783_0 & ~i_10_301_4571_0) | (i_10_301_796_0 & i_10_301_1826_0 & i_10_301_3613_0 & ~i_10_301_4271_0 & ~i_10_301_4272_0) | (i_10_301_2986_0 & i_10_301_3270_0 & ~i_10_301_4568_0));
endmodule



// Benchmark "kernel_10_302" written by ABC on Sun Jul 19 10:26:17 2020

module kernel_10_302 ( 
    i_10_302_118_0, i_10_302_171_0, i_10_302_172_0, i_10_302_244_0,
    i_10_302_249_0, i_10_302_282_0, i_10_302_285_0, i_10_302_410_0,
    i_10_302_431_0, i_10_302_462_0, i_10_302_467_0, i_10_302_800_0,
    i_10_302_957_0, i_10_302_958_0, i_10_302_959_0, i_10_302_1236_0,
    i_10_302_1237_0, i_10_302_1238_0, i_10_302_1240_0, i_10_302_1241_0,
    i_10_302_1246_0, i_10_302_1308_0, i_10_302_1309_0, i_10_302_1581_0,
    i_10_302_1582_0, i_10_302_1648_0, i_10_302_1649_0, i_10_302_1687_0,
    i_10_302_1819_0, i_10_302_1820_0, i_10_302_1821_0, i_10_302_1911_0,
    i_10_302_1916_0, i_10_302_1944_0, i_10_302_1945_0, i_10_302_1946_0,
    i_10_302_2027_0, i_10_302_2178_0, i_10_302_2179_0, i_10_302_2181_0,
    i_10_302_2184_0, i_10_302_2185_0, i_10_302_2186_0, i_10_302_2333_0,
    i_10_302_2364_0, i_10_302_2404_0, i_10_302_2407_0, i_10_302_2448_0,
    i_10_302_2503_0, i_10_302_2629_0, i_10_302_2630_0, i_10_302_2632_0,
    i_10_302_2658_0, i_10_302_2673_0, i_10_302_2700_0, i_10_302_2710_0,
    i_10_302_2712_0, i_10_302_2713_0, i_10_302_2722_0, i_10_302_2724_0,
    i_10_302_2731_0, i_10_302_2733_0, i_10_302_2882_0, i_10_302_2920_0,
    i_10_302_2923_0, i_10_302_2986_0, i_10_302_3034_0, i_10_302_3036_0,
    i_10_302_3037_0, i_10_302_3150_0, i_10_302_3156_0, i_10_302_3160_0,
    i_10_302_3195_0, i_10_302_3231_0, i_10_302_3276_0, i_10_302_3277_0,
    i_10_302_3278_0, i_10_302_3282_0, i_10_302_3409_0, i_10_302_3586_0,
    i_10_302_3611_0, i_10_302_3612_0, i_10_302_3613_0, i_10_302_3646_0,
    i_10_302_3648_0, i_10_302_3649_0, i_10_302_3784_0, i_10_302_3786_0,
    i_10_302_3787_0, i_10_302_3834_0, i_10_302_3835_0, i_10_302_3838_0,
    i_10_302_3849_0, i_10_302_4052_0, i_10_302_4267_0, i_10_302_4563_0,
    i_10_302_4566_0, i_10_302_4567_0, i_10_302_4568_0, i_10_302_4593_0,
    o_10_302_0_0  );
  input  i_10_302_118_0, i_10_302_171_0, i_10_302_172_0, i_10_302_244_0,
    i_10_302_249_0, i_10_302_282_0, i_10_302_285_0, i_10_302_410_0,
    i_10_302_431_0, i_10_302_462_0, i_10_302_467_0, i_10_302_800_0,
    i_10_302_957_0, i_10_302_958_0, i_10_302_959_0, i_10_302_1236_0,
    i_10_302_1237_0, i_10_302_1238_0, i_10_302_1240_0, i_10_302_1241_0,
    i_10_302_1246_0, i_10_302_1308_0, i_10_302_1309_0, i_10_302_1581_0,
    i_10_302_1582_0, i_10_302_1648_0, i_10_302_1649_0, i_10_302_1687_0,
    i_10_302_1819_0, i_10_302_1820_0, i_10_302_1821_0, i_10_302_1911_0,
    i_10_302_1916_0, i_10_302_1944_0, i_10_302_1945_0, i_10_302_1946_0,
    i_10_302_2027_0, i_10_302_2178_0, i_10_302_2179_0, i_10_302_2181_0,
    i_10_302_2184_0, i_10_302_2185_0, i_10_302_2186_0, i_10_302_2333_0,
    i_10_302_2364_0, i_10_302_2404_0, i_10_302_2407_0, i_10_302_2448_0,
    i_10_302_2503_0, i_10_302_2629_0, i_10_302_2630_0, i_10_302_2632_0,
    i_10_302_2658_0, i_10_302_2673_0, i_10_302_2700_0, i_10_302_2710_0,
    i_10_302_2712_0, i_10_302_2713_0, i_10_302_2722_0, i_10_302_2724_0,
    i_10_302_2731_0, i_10_302_2733_0, i_10_302_2882_0, i_10_302_2920_0,
    i_10_302_2923_0, i_10_302_2986_0, i_10_302_3034_0, i_10_302_3036_0,
    i_10_302_3037_0, i_10_302_3150_0, i_10_302_3156_0, i_10_302_3160_0,
    i_10_302_3195_0, i_10_302_3231_0, i_10_302_3276_0, i_10_302_3277_0,
    i_10_302_3278_0, i_10_302_3282_0, i_10_302_3409_0, i_10_302_3586_0,
    i_10_302_3611_0, i_10_302_3612_0, i_10_302_3613_0, i_10_302_3646_0,
    i_10_302_3648_0, i_10_302_3649_0, i_10_302_3784_0, i_10_302_3786_0,
    i_10_302_3787_0, i_10_302_3834_0, i_10_302_3835_0, i_10_302_3838_0,
    i_10_302_3849_0, i_10_302_4052_0, i_10_302_4267_0, i_10_302_4563_0,
    i_10_302_4566_0, i_10_302_4567_0, i_10_302_4568_0, i_10_302_4593_0;
  output o_10_302_0_0;
  assign o_10_302_0_0 = ~((~i_10_302_171_0 & ((~i_10_302_285_0 & ~i_10_302_1649_0 & ~i_10_302_1944_0 & ~i_10_302_2186_0 & ~i_10_302_2731_0 & ~i_10_302_3278_0 & i_10_302_3835_0 & i_10_302_3838_0) | (~i_10_302_249_0 & ~i_10_302_1582_0 & ~i_10_302_1648_0 & ~i_10_302_1945_0 & ~i_10_302_2184_0 & ~i_10_302_2333_0 & ~i_10_302_2407_0 & ~i_10_302_2503_0 & ~i_10_302_2724_0 & ~i_10_302_3612_0 & ~i_10_302_3646_0 & ~i_10_302_3784_0 & ~i_10_302_3786_0 & ~i_10_302_3787_0 & ~i_10_302_4267_0))) | (~i_10_302_958_0 & ((~i_10_302_249_0 & ~i_10_302_1944_0 & ((~i_10_302_959_0 & ~i_10_302_2184_0 & ~i_10_302_2186_0 & ~i_10_302_2629_0 & ~i_10_302_3786_0 & i_10_302_3835_0) | (~i_10_302_1236_0 & i_10_302_1821_0 & ~i_10_302_2407_0 & ~i_10_302_2630_0 & ~i_10_302_2710_0 & ~i_10_302_3036_0 & ~i_10_302_3646_0 & ~i_10_302_3787_0 & ~i_10_302_3849_0))) | (i_10_302_1819_0 & ((~i_10_302_959_0 & ~i_10_302_2700_0 & ~i_10_302_2722_0 & ~i_10_302_3586_0 & i_10_302_3611_0) | (~i_10_302_2181_0 & ~i_10_302_2503_0 & i_10_302_2733_0 & ~i_10_302_3784_0))) | (~i_10_302_2185_0 & ((~i_10_302_1649_0 & ~i_10_302_1945_0 & ~i_10_302_2700_0 & i_10_302_3277_0) | (i_10_302_1241_0 & ~i_10_302_2181_0 & ~i_10_302_2186_0 & ~i_10_302_2503_0 & ~i_10_302_2920_0 & ~i_10_302_4052_0))) | (i_10_302_1649_0 & ~i_10_302_2178_0 & ~i_10_302_2404_0 & ~i_10_302_2407_0 & ~i_10_302_2630_0 & ~i_10_302_2724_0 & ~i_10_302_3231_0 & ~i_10_302_3786_0 & ~i_10_302_4052_0) | (~i_10_302_244_0 & ~i_10_302_800_0 & ~i_10_302_1238_0 & ~i_10_302_1946_0 & i_10_302_2920_0 & i_10_302_2923_0 & ~i_10_302_3160_0 & ~i_10_302_3611_0 & ~i_10_302_3646_0 & ~i_10_302_4267_0))) | (~i_10_302_467_0 & ((~i_10_302_172_0 & ~i_10_302_282_0 & ~i_10_302_1581_0 & ~i_10_302_1582_0 & ~i_10_302_2184_0 & ~i_10_302_2185_0 & ~i_10_302_2630_0 & ~i_10_302_2700_0 & ~i_10_302_2724_0 & ~i_10_302_3646_0 & ~i_10_302_3787_0) | (i_10_302_1240_0 & ~i_10_302_2658_0 & ~i_10_302_3649_0 & ~i_10_302_4563_0))) | (~i_10_302_1946_0 & ((~i_10_302_959_0 & ~i_10_302_2184_0 & ~i_10_302_2503_0 & ((~i_10_302_244_0 & ~i_10_302_1581_0 & ~i_10_302_1649_0 & ~i_10_302_1821_0 & ~i_10_302_2179_0 & ~i_10_302_2185_0 & ~i_10_302_2629_0 & ~i_10_302_3036_0 & ~i_10_302_3277_0 & ~i_10_302_3586_0) | (~i_10_302_1236_0 & ~i_10_302_2178_0 & ~i_10_302_2404_0 & ~i_10_302_2407_0 & ~i_10_302_3034_0 & ~i_10_302_3037_0 & ~i_10_302_3649_0 & ~i_10_302_3784_0 & ~i_10_302_3849_0 & ~i_10_302_4563_0))) | (~i_10_302_1309_0 & ((~i_10_302_1916_0 & i_10_302_2724_0 & ~i_10_302_3277_0 & ~i_10_302_3649_0 & ~i_10_302_4267_0 & ~i_10_302_4563_0) | (~i_10_302_3612_0 & ~i_10_302_3646_0 & ~i_10_302_2185_0 & ~i_10_302_2920_0 & ~i_10_302_3786_0 & ~i_10_302_3787_0 & ~i_10_302_3849_0 & ~i_10_302_4566_0))) | (i_10_302_462_0 & ~i_10_302_957_0 & ~i_10_302_1648_0 & ~i_10_302_1821_0 & i_10_302_2632_0 & ~i_10_302_2673_0 & ~i_10_302_3276_0 & ~i_10_302_3409_0 & ~i_10_302_3838_0))) | (~i_10_302_244_0 & ((i_10_302_1819_0 & ~i_10_302_1945_0 & ~i_10_302_2185_0 & ~i_10_302_2503_0 & ~i_10_302_2673_0 & i_10_302_2731_0 & ~i_10_302_3276_0 & ~i_10_302_3786_0 & ~i_10_302_3838_0) | (i_10_302_467_0 & ~i_10_302_1687_0 & ~i_10_302_2186_0 & ~i_10_302_2658_0 & ~i_10_302_3036_0 & ~i_10_302_3646_0 & i_10_302_3784_0 & ~i_10_302_4563_0))) | (i_10_302_462_0 & ~i_10_302_2658_0 & ((i_10_302_2731_0 & ~i_10_302_3037_0 & i_10_302_3838_0) | (~i_10_302_1241_0 & ~i_10_302_1581_0 & ~i_10_302_1582_0 & ~i_10_302_2179_0 & ~i_10_302_2404_0 & ~i_10_302_2407_0 & ~i_10_302_3034_0 & ~i_10_302_3786_0 & ~i_10_302_4563_0 & ~i_10_302_4566_0))) | (~i_10_302_2179_0 & ((i_10_302_467_0 & i_10_302_3646_0 & ((i_10_302_1820_0 & ~i_10_302_2185_0 & i_10_302_2629_0 & ~i_10_302_2700_0 & ~i_10_302_3787_0 & ~i_10_302_4052_0) | (~i_10_302_1582_0 & ~i_10_302_1648_0 & ~i_10_302_2404_0 & i_10_302_2632_0 & ~i_10_302_2882_0 & ~i_10_302_3612_0 & ~i_10_302_4568_0))) | (i_10_302_285_0 & ~i_10_302_800_0 & ~i_10_302_1648_0 & ~i_10_302_1944_0 & ~i_10_302_2184_0 & i_10_302_2731_0 & ~i_10_302_3787_0 & ~i_10_302_3835_0))) | (~i_10_302_3786_0 & ((~i_10_302_959_0 & ((~i_10_302_1944_0 & ~i_10_302_1945_0 & ~i_10_302_2184_0 & ~i_10_302_2333_0 & ~i_10_302_2503_0 & ~i_10_302_2700_0 & i_10_302_2722_0 & ~i_10_302_3160_0 & ~i_10_302_3649_0) | (~i_10_302_957_0 & i_10_302_1237_0 & ~i_10_302_1582_0 & ~i_10_302_2407_0 & ~i_10_302_2632_0 & ~i_10_302_2673_0 & ~i_10_302_4052_0 & ~i_10_302_4566_0))) | (~i_10_302_1649_0 & i_10_302_1820_0 & ~i_10_302_2404_0 & ~i_10_302_3409_0 & ~i_10_302_3787_0 & ~i_10_302_4267_0))) | (~i_10_302_1582_0 & ((~i_10_302_957_0 & ~i_10_302_2333_0 & ~i_10_302_2407_0 & ~i_10_302_3648_0 & i_10_302_3835_0) | (~i_10_302_1649_0 & ~i_10_302_2404_0 & i_10_302_3611_0 & ~i_10_302_4052_0))) | (~i_10_302_957_0 & ~i_10_302_2185_0 & ((i_10_302_1236_0 & ~i_10_302_1648_0 & ~i_10_302_1944_0 & ~i_10_302_2733_0 & ~i_10_302_2920_0 & ~i_10_302_3160_0 & ~i_10_302_3277_0 & ~i_10_302_3784_0 & ~i_10_302_3787_0) | (i_10_302_1820_0 & ~i_10_302_2178_0 & ~i_10_302_2186_0 & ~i_10_302_2503_0 & i_10_302_3834_0))) | (~i_10_302_3037_0 & ((i_10_302_410_0 & ~i_10_302_2632_0 & ~i_10_302_3036_0 & i_10_302_3648_0 & ~i_10_302_3787_0) | (i_10_302_1238_0 & ~i_10_302_1246_0 & ~i_10_302_2364_0 & ~i_10_302_2404_0 & ~i_10_302_2986_0 & ~i_10_302_3034_0 & ~i_10_302_4052_0 & ~i_10_302_4567_0))) | (i_10_302_3195_0 & i_10_302_3278_0 & i_10_302_3611_0) | (~i_10_302_1581_0 & i_10_302_1687_0 & ~i_10_302_2629_0 & ~i_10_302_3646_0 & ~i_10_302_3784_0) | (~i_10_302_3787_0 & ~i_10_302_4267_0 & ~i_10_302_2333_0 & i_10_302_2712_0) | (i_10_302_2724_0 & i_10_302_3282_0 & ~i_10_302_3648_0 & ~i_10_302_4563_0));
endmodule



// Benchmark "kernel_10_303" written by ABC on Sun Jul 19 10:26:18 2020

module kernel_10_303 ( 
    i_10_303_175_0, i_10_303_217_0, i_10_303_221_0, i_10_303_262_0,
    i_10_303_282_0, i_10_303_283_0, i_10_303_315_0, i_10_303_320_0,
    i_10_303_426_0, i_10_303_432_0, i_10_303_466_0, i_10_303_510_0,
    i_10_303_626_0, i_10_303_631_0, i_10_303_830_0, i_10_303_954_0,
    i_10_303_990_0, i_10_303_991_0, i_10_303_1026_0, i_10_303_1027_0,
    i_10_303_1030_0, i_10_303_1117_0, i_10_303_1236_0, i_10_303_1264_0,
    i_10_303_1300_0, i_10_303_1307_0, i_10_303_1341_0, i_10_303_1431_0,
    i_10_303_1432_0, i_10_303_1539_0, i_10_303_1578_0, i_10_303_1579_0,
    i_10_303_1620_0, i_10_303_1683_0, i_10_303_1684_0, i_10_303_1818_0,
    i_10_303_2197_0, i_10_303_2359_0, i_10_303_2361_0, i_10_303_2362_0,
    i_10_303_2376_0, i_10_303_2377_0, i_10_303_2408_0, i_10_303_2565_0,
    i_10_303_2566_0, i_10_303_2638_0, i_10_303_2659_0, i_10_303_2704_0,
    i_10_303_2729_0, i_10_303_2740_0, i_10_303_2743_0, i_10_303_2844_0,
    i_10_303_2845_0, i_10_303_2885_0, i_10_303_2918_0, i_10_303_2919_0,
    i_10_303_2921_0, i_10_303_3042_0, i_10_303_3196_0, i_10_303_3223_0,
    i_10_303_3268_0, i_10_303_3384_0, i_10_303_3386_0, i_10_303_3387_0,
    i_10_303_3402_0, i_10_303_3403_0, i_10_303_3431_0, i_10_303_3452_0,
    i_10_303_3469_0, i_10_303_3485_0, i_10_303_3538_0, i_10_303_3649_0,
    i_10_303_3650_0, i_10_303_3652_0, i_10_303_3682_0, i_10_303_3781_0,
    i_10_303_3782_0, i_10_303_3783_0, i_10_303_3784_0, i_10_303_3785_0,
    i_10_303_3838_0, i_10_303_3844_0, i_10_303_3852_0, i_10_303_3853_0,
    i_10_303_3854_0, i_10_303_3961_0, i_10_303_3980_0, i_10_303_4023_0,
    i_10_303_4052_0, i_10_303_4143_0, i_10_303_4168_0, i_10_303_4173_0,
    i_10_303_4175_0, i_10_303_4213_0, i_10_303_4214_0, i_10_303_4270_0,
    i_10_303_4420_0, i_10_303_4511_0, i_10_303_4581_0, i_10_303_4600_0,
    o_10_303_0_0  );
  input  i_10_303_175_0, i_10_303_217_0, i_10_303_221_0, i_10_303_262_0,
    i_10_303_282_0, i_10_303_283_0, i_10_303_315_0, i_10_303_320_0,
    i_10_303_426_0, i_10_303_432_0, i_10_303_466_0, i_10_303_510_0,
    i_10_303_626_0, i_10_303_631_0, i_10_303_830_0, i_10_303_954_0,
    i_10_303_990_0, i_10_303_991_0, i_10_303_1026_0, i_10_303_1027_0,
    i_10_303_1030_0, i_10_303_1117_0, i_10_303_1236_0, i_10_303_1264_0,
    i_10_303_1300_0, i_10_303_1307_0, i_10_303_1341_0, i_10_303_1431_0,
    i_10_303_1432_0, i_10_303_1539_0, i_10_303_1578_0, i_10_303_1579_0,
    i_10_303_1620_0, i_10_303_1683_0, i_10_303_1684_0, i_10_303_1818_0,
    i_10_303_2197_0, i_10_303_2359_0, i_10_303_2361_0, i_10_303_2362_0,
    i_10_303_2376_0, i_10_303_2377_0, i_10_303_2408_0, i_10_303_2565_0,
    i_10_303_2566_0, i_10_303_2638_0, i_10_303_2659_0, i_10_303_2704_0,
    i_10_303_2729_0, i_10_303_2740_0, i_10_303_2743_0, i_10_303_2844_0,
    i_10_303_2845_0, i_10_303_2885_0, i_10_303_2918_0, i_10_303_2919_0,
    i_10_303_2921_0, i_10_303_3042_0, i_10_303_3196_0, i_10_303_3223_0,
    i_10_303_3268_0, i_10_303_3384_0, i_10_303_3386_0, i_10_303_3387_0,
    i_10_303_3402_0, i_10_303_3403_0, i_10_303_3431_0, i_10_303_3452_0,
    i_10_303_3469_0, i_10_303_3485_0, i_10_303_3538_0, i_10_303_3649_0,
    i_10_303_3650_0, i_10_303_3652_0, i_10_303_3682_0, i_10_303_3781_0,
    i_10_303_3782_0, i_10_303_3783_0, i_10_303_3784_0, i_10_303_3785_0,
    i_10_303_3838_0, i_10_303_3844_0, i_10_303_3852_0, i_10_303_3853_0,
    i_10_303_3854_0, i_10_303_3961_0, i_10_303_3980_0, i_10_303_4023_0,
    i_10_303_4052_0, i_10_303_4143_0, i_10_303_4168_0, i_10_303_4173_0,
    i_10_303_4175_0, i_10_303_4213_0, i_10_303_4214_0, i_10_303_4270_0,
    i_10_303_4420_0, i_10_303_4511_0, i_10_303_4581_0, i_10_303_4600_0;
  output o_10_303_0_0;
  assign o_10_303_0_0 = 0;
endmodule



// Benchmark "kernel_10_304" written by ABC on Sun Jul 19 10:26:18 2020

module kernel_10_304 ( 
    i_10_304_29_0, i_10_304_154_0, i_10_304_181_0, i_10_304_282_0,
    i_10_304_315_0, i_10_304_316_0, i_10_304_319_0, i_10_304_390_0,
    i_10_304_436_0, i_10_304_464_0, i_10_304_465_0, i_10_304_467_0,
    i_10_304_505_0, i_10_304_820_0, i_10_304_829_0, i_10_304_999_0,
    i_10_304_1053_0, i_10_304_1081_0, i_10_304_1083_0, i_10_304_1084_0,
    i_10_304_1154_0, i_10_304_1239_0, i_10_304_1240_0, i_10_304_1241_0,
    i_10_304_1265_0, i_10_304_1360_0, i_10_304_1539_0, i_10_304_1540_0,
    i_10_304_1542_0, i_10_304_1575_0, i_10_304_1579_0, i_10_304_1620_0,
    i_10_304_1621_0, i_10_304_1622_0, i_10_304_1650_0, i_10_304_1686_0,
    i_10_304_1687_0, i_10_304_1688_0, i_10_304_1909_0, i_10_304_1999_0,
    i_10_304_2008_0, i_10_304_2025_0, i_10_304_2183_0, i_10_304_2196_0,
    i_10_304_2197_0, i_10_304_2198_0, i_10_304_2199_0, i_10_304_2236_0,
    i_10_304_2350_0, i_10_304_2352_0, i_10_304_2353_0, i_10_304_2364_0,
    i_10_304_2406_0, i_10_304_2407_0, i_10_304_2572_0, i_10_304_2636_0,
    i_10_304_2659_0, i_10_304_2674_0, i_10_304_2675_0, i_10_304_2700_0,
    i_10_304_2701_0, i_10_304_2831_0, i_10_304_2882_0, i_10_304_2884_0,
    i_10_304_2922_0, i_10_304_2923_0, i_10_304_3276_0, i_10_304_3277_0,
    i_10_304_3278_0, i_10_304_3279_0, i_10_304_3280_0, i_10_304_3281_0,
    i_10_304_3316_0, i_10_304_3429_0, i_10_304_3448_0, i_10_304_3468_0,
    i_10_304_3469_0, i_10_304_3538_0, i_10_304_3541_0, i_10_304_3542_0,
    i_10_304_3555_0, i_10_304_3558_0, i_10_304_3559_0, i_10_304_3586_0,
    i_10_304_3836_0, i_10_304_3979_0, i_10_304_3980_0, i_10_304_4050_0,
    i_10_304_4113_0, i_10_304_4119_0, i_10_304_4125_0, i_10_304_4126_0,
    i_10_304_4127_0, i_10_304_4167_0, i_10_304_4170_0, i_10_304_4172_0,
    i_10_304_4276_0, i_10_304_4282_0, i_10_304_4546_0, i_10_304_4565_0,
    o_10_304_0_0  );
  input  i_10_304_29_0, i_10_304_154_0, i_10_304_181_0, i_10_304_282_0,
    i_10_304_315_0, i_10_304_316_0, i_10_304_319_0, i_10_304_390_0,
    i_10_304_436_0, i_10_304_464_0, i_10_304_465_0, i_10_304_467_0,
    i_10_304_505_0, i_10_304_820_0, i_10_304_829_0, i_10_304_999_0,
    i_10_304_1053_0, i_10_304_1081_0, i_10_304_1083_0, i_10_304_1084_0,
    i_10_304_1154_0, i_10_304_1239_0, i_10_304_1240_0, i_10_304_1241_0,
    i_10_304_1265_0, i_10_304_1360_0, i_10_304_1539_0, i_10_304_1540_0,
    i_10_304_1542_0, i_10_304_1575_0, i_10_304_1579_0, i_10_304_1620_0,
    i_10_304_1621_0, i_10_304_1622_0, i_10_304_1650_0, i_10_304_1686_0,
    i_10_304_1687_0, i_10_304_1688_0, i_10_304_1909_0, i_10_304_1999_0,
    i_10_304_2008_0, i_10_304_2025_0, i_10_304_2183_0, i_10_304_2196_0,
    i_10_304_2197_0, i_10_304_2198_0, i_10_304_2199_0, i_10_304_2236_0,
    i_10_304_2350_0, i_10_304_2352_0, i_10_304_2353_0, i_10_304_2364_0,
    i_10_304_2406_0, i_10_304_2407_0, i_10_304_2572_0, i_10_304_2636_0,
    i_10_304_2659_0, i_10_304_2674_0, i_10_304_2675_0, i_10_304_2700_0,
    i_10_304_2701_0, i_10_304_2831_0, i_10_304_2882_0, i_10_304_2884_0,
    i_10_304_2922_0, i_10_304_2923_0, i_10_304_3276_0, i_10_304_3277_0,
    i_10_304_3278_0, i_10_304_3279_0, i_10_304_3280_0, i_10_304_3281_0,
    i_10_304_3316_0, i_10_304_3429_0, i_10_304_3448_0, i_10_304_3468_0,
    i_10_304_3469_0, i_10_304_3538_0, i_10_304_3541_0, i_10_304_3542_0,
    i_10_304_3555_0, i_10_304_3558_0, i_10_304_3559_0, i_10_304_3586_0,
    i_10_304_3836_0, i_10_304_3979_0, i_10_304_3980_0, i_10_304_4050_0,
    i_10_304_4113_0, i_10_304_4119_0, i_10_304_4125_0, i_10_304_4126_0,
    i_10_304_4127_0, i_10_304_4167_0, i_10_304_4170_0, i_10_304_4172_0,
    i_10_304_4276_0, i_10_304_4282_0, i_10_304_4546_0, i_10_304_4565_0;
  output o_10_304_0_0;
  assign o_10_304_0_0 = 0;
endmodule



// Benchmark "kernel_10_305" written by ABC on Sun Jul 19 10:26:19 2020

module kernel_10_305 ( 
    i_10_305_32_0, i_10_305_152_0, i_10_305_157_0, i_10_305_174_0,
    i_10_305_179_0, i_10_305_256_0, i_10_305_257_0, i_10_305_262_0,
    i_10_305_266_0, i_10_305_281_0, i_10_305_394_0, i_10_305_410_0,
    i_10_305_430_0, i_10_305_440_0, i_10_305_441_0, i_10_305_464_0,
    i_10_305_548_0, i_10_305_796_0, i_10_305_800_0, i_10_305_962_0,
    i_10_305_1003_0, i_10_305_1004_0, i_10_305_1031_0, i_10_305_1039_0,
    i_10_305_1084_0, i_10_305_1234_0, i_10_305_1236_0, i_10_305_1250_0,
    i_10_305_1344_0, i_10_305_1432_0, i_10_305_1433_0, i_10_305_1546_0,
    i_10_305_1555_0, i_10_305_1556_0, i_10_305_1655_0, i_10_305_1687_0,
    i_10_305_1689_0, i_10_305_1690_0, i_10_305_1813_0, i_10_305_1826_0,
    i_10_305_1915_0, i_10_305_1945_0, i_10_305_1946_0, i_10_305_1948_0,
    i_10_305_2332_0, i_10_305_2356_0, i_10_305_2382_0, i_10_305_2448_0,
    i_10_305_2452_0, i_10_305_2456_0, i_10_305_2468_0, i_10_305_2516_0,
    i_10_305_2519_0, i_10_305_2628_0, i_10_305_2632_0, i_10_305_2633_0,
    i_10_305_2636_0, i_10_305_2657_0, i_10_305_2660_0, i_10_305_2707_0,
    i_10_305_2719_0, i_10_305_2721_0, i_10_305_2727_0, i_10_305_2730_0,
    i_10_305_2731_0, i_10_305_2781_0, i_10_305_2785_0, i_10_305_2829_0,
    i_10_305_2830_0, i_10_305_2832_0, i_10_305_2833_0, i_10_305_3013_0,
    i_10_305_3033_0, i_10_305_3034_0, i_10_305_3076_0, i_10_305_3199_0,
    i_10_305_3200_0, i_10_305_3201_0, i_10_305_3316_0, i_10_305_3386_0,
    i_10_305_3469_0, i_10_305_3473_0, i_10_305_3493_0, i_10_305_3541_0,
    i_10_305_3587_0, i_10_305_3615_0, i_10_305_3626_0, i_10_305_3646_0,
    i_10_305_3841_0, i_10_305_3849_0, i_10_305_3850_0, i_10_305_3853_0,
    i_10_305_3859_0, i_10_305_3990_0, i_10_305_4052_0, i_10_305_4114_0,
    i_10_305_4115_0, i_10_305_4117_0, i_10_305_4121_0, i_10_305_4288_0,
    o_10_305_0_0  );
  input  i_10_305_32_0, i_10_305_152_0, i_10_305_157_0, i_10_305_174_0,
    i_10_305_179_0, i_10_305_256_0, i_10_305_257_0, i_10_305_262_0,
    i_10_305_266_0, i_10_305_281_0, i_10_305_394_0, i_10_305_410_0,
    i_10_305_430_0, i_10_305_440_0, i_10_305_441_0, i_10_305_464_0,
    i_10_305_548_0, i_10_305_796_0, i_10_305_800_0, i_10_305_962_0,
    i_10_305_1003_0, i_10_305_1004_0, i_10_305_1031_0, i_10_305_1039_0,
    i_10_305_1084_0, i_10_305_1234_0, i_10_305_1236_0, i_10_305_1250_0,
    i_10_305_1344_0, i_10_305_1432_0, i_10_305_1433_0, i_10_305_1546_0,
    i_10_305_1555_0, i_10_305_1556_0, i_10_305_1655_0, i_10_305_1687_0,
    i_10_305_1689_0, i_10_305_1690_0, i_10_305_1813_0, i_10_305_1826_0,
    i_10_305_1915_0, i_10_305_1945_0, i_10_305_1946_0, i_10_305_1948_0,
    i_10_305_2332_0, i_10_305_2356_0, i_10_305_2382_0, i_10_305_2448_0,
    i_10_305_2452_0, i_10_305_2456_0, i_10_305_2468_0, i_10_305_2516_0,
    i_10_305_2519_0, i_10_305_2628_0, i_10_305_2632_0, i_10_305_2633_0,
    i_10_305_2636_0, i_10_305_2657_0, i_10_305_2660_0, i_10_305_2707_0,
    i_10_305_2719_0, i_10_305_2721_0, i_10_305_2727_0, i_10_305_2730_0,
    i_10_305_2731_0, i_10_305_2781_0, i_10_305_2785_0, i_10_305_2829_0,
    i_10_305_2830_0, i_10_305_2832_0, i_10_305_2833_0, i_10_305_3013_0,
    i_10_305_3033_0, i_10_305_3034_0, i_10_305_3076_0, i_10_305_3199_0,
    i_10_305_3200_0, i_10_305_3201_0, i_10_305_3316_0, i_10_305_3386_0,
    i_10_305_3469_0, i_10_305_3473_0, i_10_305_3493_0, i_10_305_3541_0,
    i_10_305_3587_0, i_10_305_3615_0, i_10_305_3626_0, i_10_305_3646_0,
    i_10_305_3841_0, i_10_305_3849_0, i_10_305_3850_0, i_10_305_3853_0,
    i_10_305_3859_0, i_10_305_3990_0, i_10_305_4052_0, i_10_305_4114_0,
    i_10_305_4115_0, i_10_305_4117_0, i_10_305_4121_0, i_10_305_4288_0;
  output o_10_305_0_0;
  assign o_10_305_0_0 = 0;
endmodule



// Benchmark "kernel_10_306" written by ABC on Sun Jul 19 10:26:21 2020

module kernel_10_306 ( 
    i_10_306_118_0, i_10_306_153_0, i_10_306_243_0, i_10_306_244_0,
    i_10_306_253_0, i_10_306_284_0, i_10_306_388_0, i_10_306_390_0,
    i_10_306_460_0, i_10_306_462_0, i_10_306_513_0, i_10_306_687_0,
    i_10_306_711_0, i_10_306_747_0, i_10_306_748_0, i_10_306_794_0,
    i_10_306_1000_0, i_10_306_1035_0, i_10_306_1242_0, i_10_306_1246_0,
    i_10_306_1261_0, i_10_306_1263_0, i_10_306_1307_0, i_10_306_1308_0,
    i_10_306_1359_0, i_10_306_1360_0, i_10_306_1530_0, i_10_306_1612_0,
    i_10_306_1647_0, i_10_306_1648_0, i_10_306_1650_0, i_10_306_1651_0,
    i_10_306_1652_0, i_10_306_1654_0, i_10_306_1674_0, i_10_306_1683_0,
    i_10_306_1711_0, i_10_306_1809_0, i_10_306_1810_0, i_10_306_1819_0,
    i_10_306_1822_0, i_10_306_1911_0, i_10_306_1913_0, i_10_306_2178_0,
    i_10_306_2179_0, i_10_306_2199_0, i_10_306_2202_0, i_10_306_2308_0,
    i_10_306_2349_0, i_10_306_2350_0, i_10_306_2355_0, i_10_306_2380_0,
    i_10_306_2406_0, i_10_306_2451_0, i_10_306_2452_0, i_10_306_2467_0,
    i_10_306_2513_0, i_10_306_2601_0, i_10_306_2628_0, i_10_306_2631_0,
    i_10_306_2658_0, i_10_306_2659_0, i_10_306_2660_0, i_10_306_2718_0,
    i_10_306_2721_0, i_10_306_2722_0, i_10_306_2727_0, i_10_306_2740_0,
    i_10_306_2817_0, i_10_306_2818_0, i_10_306_2820_0, i_10_306_2829_0,
    i_10_306_2834_0, i_10_306_2881_0, i_10_306_3088_0, i_10_306_3231_0,
    i_10_306_3386_0, i_10_306_3466_0, i_10_306_3519_0, i_10_306_3522_0,
    i_10_306_3583_0, i_10_306_3646_0, i_10_306_3647_0, i_10_306_3788_0,
    i_10_306_3834_0, i_10_306_3847_0, i_10_306_3848_0, i_10_306_3856_0,
    i_10_306_3889_0, i_10_306_3906_0, i_10_306_3980_0, i_10_306_4023_0,
    i_10_306_4113_0, i_10_306_4122_0, i_10_306_4267_0, i_10_306_4269_0,
    i_10_306_4273_0, i_10_306_4284_0, i_10_306_4287_0, i_10_306_4571_0,
    o_10_306_0_0  );
  input  i_10_306_118_0, i_10_306_153_0, i_10_306_243_0, i_10_306_244_0,
    i_10_306_253_0, i_10_306_284_0, i_10_306_388_0, i_10_306_390_0,
    i_10_306_460_0, i_10_306_462_0, i_10_306_513_0, i_10_306_687_0,
    i_10_306_711_0, i_10_306_747_0, i_10_306_748_0, i_10_306_794_0,
    i_10_306_1000_0, i_10_306_1035_0, i_10_306_1242_0, i_10_306_1246_0,
    i_10_306_1261_0, i_10_306_1263_0, i_10_306_1307_0, i_10_306_1308_0,
    i_10_306_1359_0, i_10_306_1360_0, i_10_306_1530_0, i_10_306_1612_0,
    i_10_306_1647_0, i_10_306_1648_0, i_10_306_1650_0, i_10_306_1651_0,
    i_10_306_1652_0, i_10_306_1654_0, i_10_306_1674_0, i_10_306_1683_0,
    i_10_306_1711_0, i_10_306_1809_0, i_10_306_1810_0, i_10_306_1819_0,
    i_10_306_1822_0, i_10_306_1911_0, i_10_306_1913_0, i_10_306_2178_0,
    i_10_306_2179_0, i_10_306_2199_0, i_10_306_2202_0, i_10_306_2308_0,
    i_10_306_2349_0, i_10_306_2350_0, i_10_306_2355_0, i_10_306_2380_0,
    i_10_306_2406_0, i_10_306_2451_0, i_10_306_2452_0, i_10_306_2467_0,
    i_10_306_2513_0, i_10_306_2601_0, i_10_306_2628_0, i_10_306_2631_0,
    i_10_306_2658_0, i_10_306_2659_0, i_10_306_2660_0, i_10_306_2718_0,
    i_10_306_2721_0, i_10_306_2722_0, i_10_306_2727_0, i_10_306_2740_0,
    i_10_306_2817_0, i_10_306_2818_0, i_10_306_2820_0, i_10_306_2829_0,
    i_10_306_2834_0, i_10_306_2881_0, i_10_306_3088_0, i_10_306_3231_0,
    i_10_306_3386_0, i_10_306_3466_0, i_10_306_3519_0, i_10_306_3522_0,
    i_10_306_3583_0, i_10_306_3646_0, i_10_306_3647_0, i_10_306_3788_0,
    i_10_306_3834_0, i_10_306_3847_0, i_10_306_3848_0, i_10_306_3856_0,
    i_10_306_3889_0, i_10_306_3906_0, i_10_306_3980_0, i_10_306_4023_0,
    i_10_306_4113_0, i_10_306_4122_0, i_10_306_4267_0, i_10_306_4269_0,
    i_10_306_4273_0, i_10_306_4284_0, i_10_306_4287_0, i_10_306_4571_0;
  output o_10_306_0_0;
  assign o_10_306_0_0 = ~((~i_10_306_747_0 & ((~i_10_306_253_0 & ((~i_10_306_1246_0 & ~i_10_306_1648_0 & ~i_10_306_2406_0) | (~i_10_306_462_0 & ~i_10_306_748_0 & i_10_306_794_0 & ~i_10_306_1035_0 & ~i_10_306_1263_0 & ~i_10_306_2349_0 & ~i_10_306_3519_0 & ~i_10_306_4269_0))) | (~i_10_306_513_0 & ((~i_10_306_748_0 & i_10_306_1654_0 & ~i_10_306_2601_0 & ~i_10_306_3583_0 & ~i_10_306_3847_0 & ~i_10_306_4269_0) | (~i_10_306_2406_0 & ~i_10_306_2658_0 & ~i_10_306_2829_0 & ~i_10_306_3386_0 & ~i_10_306_3647_0 & ~i_10_306_4287_0))) | (~i_10_306_462_0 & ~i_10_306_1035_0 & ~i_10_306_1652_0 & i_10_306_2628_0 & ~i_10_306_2721_0 & ~i_10_306_3848_0))) | (~i_10_306_748_0 & ((~i_10_306_513_0 & ((~i_10_306_1035_0 & ~i_10_306_1242_0 & ~i_10_306_1647_0 & ~i_10_306_2601_0 & ~i_10_306_3788_0) | (~i_10_306_243_0 & ~i_10_306_1359_0 & ~i_10_306_1652_0 & ~i_10_306_4267_0 & ~i_10_306_4273_0))) | (~i_10_306_3231_0 & ((~i_10_306_1650_0 & ~i_10_306_1809_0 & ~i_10_306_2601_0) | (~i_10_306_1242_0 & ~i_10_306_1648_0 & ~i_10_306_3647_0))) | (~i_10_306_1035_0 & ~i_10_306_1647_0 & ~i_10_306_2349_0 & ~i_10_306_2628_0 & ~i_10_306_3847_0))) | (~i_10_306_711_0 & ((~i_10_306_1308_0 & ~i_10_306_1359_0 & ~i_10_306_1647_0 & ~i_10_306_1809_0 & ~i_10_306_2601_0 & ~i_10_306_2727_0 & ~i_10_306_4267_0) | (i_10_306_460_0 & ~i_10_306_1035_0 & ~i_10_306_1648_0 & ~i_10_306_3906_0 & ~i_10_306_4273_0))) | (~i_10_306_244_0 & ((~i_10_306_1035_0 & ((~i_10_306_1242_0 & ~i_10_306_1263_0 & ~i_10_306_1307_0 & ~i_10_306_1913_0 & ~i_10_306_2406_0 & ~i_10_306_2601_0 & ~i_10_306_2817_0 & ~i_10_306_3386_0 & ~i_10_306_3889_0 & ~i_10_306_3980_0) | (~i_10_306_462_0 & ~i_10_306_1000_0 & ~i_10_306_1359_0 & ~i_10_306_2178_0 & ~i_10_306_2718_0 & ~i_10_306_3834_0 & i_10_306_4267_0))) | (i_10_306_1651_0 & ~i_10_306_1652_0 & ~i_10_306_2718_0 & ~i_10_306_2721_0 & ~i_10_306_2727_0 & ~i_10_306_3856_0 & ~i_10_306_3889_0))) | (~i_10_306_462_0 & ((~i_10_306_1652_0 & i_10_306_2178_0 & i_10_306_3980_0) | (i_10_306_2349_0 & ~i_10_306_2350_0 & ~i_10_306_4113_0))) | (~i_10_306_2628_0 & ((~i_10_306_1648_0 & ~i_10_306_1652_0) | (~i_10_306_1308_0 & ~i_10_306_2355_0 & i_10_306_3834_0 & ~i_10_306_3889_0 & ~i_10_306_4113_0 & ~i_10_306_4287_0))) | (~i_10_306_2355_0 & ((i_10_306_2179_0 & i_10_306_2308_0 & i_10_306_3980_0) | (~i_10_306_794_0 & ~i_10_306_1242_0 & ~i_10_306_2452_0 & ~i_10_306_2718_0 & ~i_10_306_2727_0 & ~i_10_306_2818_0 & ~i_10_306_2829_0 & ~i_10_306_3231_0 & ~i_10_306_3834_0 & ~i_10_306_4284_0))) | (i_10_306_1612_0 & ~i_10_306_3646_0 & ~i_10_306_3848_0));
endmodule



// Benchmark "kernel_10_307" written by ABC on Sun Jul 19 10:26:22 2020

module kernel_10_307 ( 
    i_10_307_177_0, i_10_307_266_0, i_10_307_268_0, i_10_307_269_0,
    i_10_307_276_0, i_10_307_282_0, i_10_307_319_0, i_10_307_323_0,
    i_10_307_388_0, i_10_307_391_0, i_10_307_393_0, i_10_307_431_0,
    i_10_307_439_0, i_10_307_464_0, i_10_307_560_0, i_10_307_798_0,
    i_10_307_799_0, i_10_307_800_0, i_10_307_1026_0, i_10_307_1136_0,
    i_10_307_1233_0, i_10_307_1241_0, i_10_307_1246_0, i_10_307_1267_0,
    i_10_307_1308_0, i_10_307_1309_0, i_10_307_1310_0, i_10_307_1312_0,
    i_10_307_1582_0, i_10_307_1583_0, i_10_307_1655_0, i_10_307_1821_0,
    i_10_307_1822_0, i_10_307_1823_0, i_10_307_1912_0, i_10_307_1915_0,
    i_10_307_2006_0, i_10_307_2179_0, i_10_307_2354_0, i_10_307_2356_0,
    i_10_307_2357_0, i_10_307_2365_0, i_10_307_2452_0, i_10_307_2453_0,
    i_10_307_2471_0, i_10_307_2472_0, i_10_307_2473_0, i_10_307_2516_0,
    i_10_307_2611_0, i_10_307_2631_0, i_10_307_2632_0, i_10_307_2635_0,
    i_10_307_2663_0, i_10_307_2721_0, i_10_307_2722_0, i_10_307_2723_0,
    i_10_307_2731_0, i_10_307_2732_0, i_10_307_2733_0, i_10_307_2734_0,
    i_10_307_2735_0, i_10_307_2834_0, i_10_307_2883_0, i_10_307_2884_0,
    i_10_307_2923_0, i_10_307_3035_0, i_10_307_3037_0, i_10_307_3045_0,
    i_10_307_3048_0, i_10_307_3049_0, i_10_307_3151_0, i_10_307_3154_0,
    i_10_307_3155_0, i_10_307_3201_0, i_10_307_3388_0, i_10_307_3389_0,
    i_10_307_3472_0, i_10_307_3523_0, i_10_307_3613_0, i_10_307_3688_0,
    i_10_307_3780_0, i_10_307_3783_0, i_10_307_3785_0, i_10_307_3837_0,
    i_10_307_3847_0, i_10_307_3850_0, i_10_307_3851_0, i_10_307_3855_0,
    i_10_307_3984_0, i_10_307_3985_0, i_10_307_3986_0, i_10_307_4128_0,
    i_10_307_4129_0, i_10_307_4130_0, i_10_307_4271_0, i_10_307_4282_0,
    i_10_307_4290_0, i_10_307_4291_0, i_10_307_4568_0, i_10_307_4571_0,
    o_10_307_0_0  );
  input  i_10_307_177_0, i_10_307_266_0, i_10_307_268_0, i_10_307_269_0,
    i_10_307_276_0, i_10_307_282_0, i_10_307_319_0, i_10_307_323_0,
    i_10_307_388_0, i_10_307_391_0, i_10_307_393_0, i_10_307_431_0,
    i_10_307_439_0, i_10_307_464_0, i_10_307_560_0, i_10_307_798_0,
    i_10_307_799_0, i_10_307_800_0, i_10_307_1026_0, i_10_307_1136_0,
    i_10_307_1233_0, i_10_307_1241_0, i_10_307_1246_0, i_10_307_1267_0,
    i_10_307_1308_0, i_10_307_1309_0, i_10_307_1310_0, i_10_307_1312_0,
    i_10_307_1582_0, i_10_307_1583_0, i_10_307_1655_0, i_10_307_1821_0,
    i_10_307_1822_0, i_10_307_1823_0, i_10_307_1912_0, i_10_307_1915_0,
    i_10_307_2006_0, i_10_307_2179_0, i_10_307_2354_0, i_10_307_2356_0,
    i_10_307_2357_0, i_10_307_2365_0, i_10_307_2452_0, i_10_307_2453_0,
    i_10_307_2471_0, i_10_307_2472_0, i_10_307_2473_0, i_10_307_2516_0,
    i_10_307_2611_0, i_10_307_2631_0, i_10_307_2632_0, i_10_307_2635_0,
    i_10_307_2663_0, i_10_307_2721_0, i_10_307_2722_0, i_10_307_2723_0,
    i_10_307_2731_0, i_10_307_2732_0, i_10_307_2733_0, i_10_307_2734_0,
    i_10_307_2735_0, i_10_307_2834_0, i_10_307_2883_0, i_10_307_2884_0,
    i_10_307_2923_0, i_10_307_3035_0, i_10_307_3037_0, i_10_307_3045_0,
    i_10_307_3048_0, i_10_307_3049_0, i_10_307_3151_0, i_10_307_3154_0,
    i_10_307_3155_0, i_10_307_3201_0, i_10_307_3388_0, i_10_307_3389_0,
    i_10_307_3472_0, i_10_307_3523_0, i_10_307_3613_0, i_10_307_3688_0,
    i_10_307_3780_0, i_10_307_3783_0, i_10_307_3785_0, i_10_307_3837_0,
    i_10_307_3847_0, i_10_307_3850_0, i_10_307_3851_0, i_10_307_3855_0,
    i_10_307_3984_0, i_10_307_3985_0, i_10_307_3986_0, i_10_307_4128_0,
    i_10_307_4129_0, i_10_307_4130_0, i_10_307_4271_0, i_10_307_4282_0,
    i_10_307_4290_0, i_10_307_4291_0, i_10_307_4568_0, i_10_307_4571_0;
  output o_10_307_0_0;
  assign o_10_307_0_0 = ~((~i_10_307_268_0 & ~i_10_307_3780_0 & ((~i_10_307_1583_0 & ~i_10_307_1915_0 & ~i_10_307_2179_0 & ~i_10_307_2357_0 & ~i_10_307_2734_0 & ~i_10_307_3037_0 & ~i_10_307_3984_0) | (~i_10_307_319_0 & ~i_10_307_2356_0 & ~i_10_307_2611_0 & ~i_10_307_2663_0 & ~i_10_307_2733_0 & ~i_10_307_2834_0 & ~i_10_307_2883_0 & ~i_10_307_4282_0))) | (~i_10_307_2834_0 & ((~i_10_307_319_0 & ((i_10_307_2723_0 & ~i_10_307_2733_0 & ~i_10_307_3785_0) | (~i_10_307_560_0 & ~i_10_307_1821_0 & i_10_307_3037_0 & ~i_10_307_3049_0 & ~i_10_307_3472_0 & ~i_10_307_3847_0 & ~i_10_307_4282_0))) | (~i_10_307_269_0 & ~i_10_307_282_0 & ~i_10_307_388_0 & ~i_10_307_560_0 & ~i_10_307_1583_0 & ~i_10_307_2733_0 & ~i_10_307_2735_0 & ~i_10_307_3049_0 & ~i_10_307_3201_0 & ~i_10_307_3783_0))) | (~i_10_307_323_0 & ((~i_10_307_266_0 & ~i_10_307_269_0 & ~i_10_307_1308_0 & ~i_10_307_2611_0 & ~i_10_307_4129_0 & ~i_10_307_4282_0) | (~i_10_307_1583_0 & ~i_10_307_1655_0 & ~i_10_307_2453_0 & ~i_10_307_2472_0 & i_10_307_4291_0))) | (~i_10_307_266_0 & ((~i_10_307_269_0 & ~i_10_307_393_0 & ~i_10_307_1026_0 & i_10_307_1308_0 & ~i_10_307_1583_0 & ~i_10_307_2179_0 & ~i_10_307_2734_0 & ~i_10_307_2884_0) | (~i_10_307_1582_0 & ~i_10_307_1822_0 & ~i_10_307_2006_0 & ~i_10_307_2735_0 & ~i_10_307_3855_0 & ~i_10_307_4282_0))) | (i_10_307_2632_0 & ((~i_10_307_388_0 & ((~i_10_307_439_0 & ~i_10_307_1823_0 & ~i_10_307_2635_0 & i_10_307_3035_0 & ~i_10_307_3472_0) | (~i_10_307_2471_0 & ~i_10_307_2735_0 & ~i_10_307_2884_0 & ~i_10_307_3045_0 & ~i_10_307_3389_0 & ~i_10_307_3783_0 & ~i_10_307_3851_0 & ~i_10_307_3986_0))) | (~i_10_307_1582_0 & i_10_307_2721_0 & ~i_10_307_3045_0) | (i_10_307_2631_0 & i_10_307_2635_0 & i_10_307_2834_0 & ~i_10_307_3472_0 & ~i_10_307_4282_0))) | (~i_10_307_439_0 & ((~i_10_307_464_0 & i_10_307_1582_0 & ~i_10_307_2453_0 & ~i_10_307_2734_0 & ~i_10_307_3049_0 & ~i_10_307_3613_0 & ~i_10_307_3986_0) | (~i_10_307_391_0 & ~i_10_307_2179_0 & ~i_10_307_2884_0 & i_10_307_2923_0 & ~i_10_307_4282_0))) | (~i_10_307_1267_0 & ~i_10_307_3855_0 & ((~i_10_307_1309_0 & ~i_10_307_1310_0 & ~i_10_307_2723_0 & ~i_10_307_3045_0 & ~i_10_307_3049_0 & ~i_10_307_3783_0 & i_10_307_3837_0) | (~i_10_307_269_0 & ~i_10_307_560_0 & ~i_10_307_2006_0 & ~i_10_307_2452_0 & ~i_10_307_2472_0 & ~i_10_307_2883_0 & ~i_10_307_3035_0 & ~i_10_307_3847_0 & ~i_10_307_3985_0 & ~i_10_307_3986_0))) | (~i_10_307_1821_0 & ((~i_10_307_1655_0 & ~i_10_307_1822_0 & ~i_10_307_2357_0 & ~i_10_307_2611_0 & ~i_10_307_3035_0 & ~i_10_307_3049_0) | (~i_10_307_1582_0 & ~i_10_307_3037_0 & i_10_307_3837_0))) | (i_10_307_2722_0 & ((~i_10_307_2723_0 & i_10_307_3780_0) | (~i_10_307_2006_0 & ~i_10_307_2611_0 & ~i_10_307_3035_0 & ~i_10_307_3613_0 & ~i_10_307_3837_0 & ~i_10_307_3984_0))) | (~i_10_307_3472_0 & ((i_10_307_2354_0 & ~i_10_307_2453_0 & i_10_307_3389_0) | (~i_10_307_2179_0 & ~i_10_307_2356_0 & ~i_10_307_2357_0 & i_10_307_2453_0 & ~i_10_307_3785_0 & ~i_10_307_3986_0 & ~i_10_307_4128_0 & ~i_10_307_4282_0))) | (~i_10_307_1310_0 & i_10_307_2452_0 & i_10_307_2611_0 & ~i_10_307_3045_0 & ~i_10_307_3837_0) | (~i_10_307_3613_0 & i_10_307_3780_0 & i_10_307_3847_0) | (i_10_307_1026_0 & i_10_307_3388_0 & ~i_10_307_3688_0 & ~i_10_307_4282_0 & ~i_10_307_4291_0));
endmodule



// Benchmark "kernel_10_308" written by ABC on Sun Jul 19 10:26:23 2020

module kernel_10_308 ( 
    i_10_308_89_0, i_10_308_146_0, i_10_308_221_0, i_10_308_284_0,
    i_10_308_286_0, i_10_308_320_0, i_10_308_327_0, i_10_308_329_0,
    i_10_308_330_0, i_10_308_331_0, i_10_308_437_0, i_10_308_443_0,
    i_10_308_462_0, i_10_308_463_0, i_10_308_464_0, i_10_308_467_0,
    i_10_308_514_0, i_10_308_711_0, i_10_308_719_0, i_10_308_748_0,
    i_10_308_749_0, i_10_308_797_0, i_10_308_800_0, i_10_308_990_0,
    i_10_308_991_0, i_10_308_1036_0, i_10_308_1174_0, i_10_308_1235_0,
    i_10_308_1239_0, i_10_308_1240_0, i_10_308_1241_0, i_10_308_1263_0,
    i_10_308_1265_0, i_10_308_1310_0, i_10_308_1342_0, i_10_308_1397_0,
    i_10_308_1610_0, i_10_308_1685_0, i_10_308_1826_0, i_10_308_1908_0,
    i_10_308_1911_0, i_10_308_1916_0, i_10_308_1990_0, i_10_308_1998_0,
    i_10_308_2200_0, i_10_308_2201_0, i_10_308_2335_0, i_10_308_2354_0,
    i_10_308_2407_0, i_10_308_2454_0, i_10_308_2456_0, i_10_308_2470_0,
    i_10_308_2503_0, i_10_308_2516_0, i_10_308_2567_0, i_10_308_2602_0,
    i_10_308_2605_0, i_10_308_2606_0, i_10_308_2629_0, i_10_308_2630_0,
    i_10_308_2661_0, i_10_308_2716_0, i_10_308_2720_0, i_10_308_2722_0,
    i_10_308_2724_0, i_10_308_2729_0, i_10_308_2782_0, i_10_308_2817_0,
    i_10_308_2829_0, i_10_308_2883_0, i_10_308_2953_0, i_10_308_3087_0,
    i_10_308_3088_0, i_10_308_3128_0, i_10_308_3199_0, i_10_308_3201_0,
    i_10_308_3202_0, i_10_308_3267_0, i_10_308_3385_0, i_10_308_3404_0,
    i_10_308_3523_0, i_10_308_3544_0, i_10_308_3557_0, i_10_308_3613_0,
    i_10_308_3614_0, i_10_308_3720_0, i_10_308_3733_0, i_10_308_3837_0,
    i_10_308_3847_0, i_10_308_3856_0, i_10_308_3881_0, i_10_308_4115_0,
    i_10_308_4277_0, i_10_308_4280_0, i_10_308_4284_0, i_10_308_4289_0,
    i_10_308_4351_0, i_10_308_4432_0, i_10_308_4569_0, i_10_308_4570_0,
    o_10_308_0_0  );
  input  i_10_308_89_0, i_10_308_146_0, i_10_308_221_0, i_10_308_284_0,
    i_10_308_286_0, i_10_308_320_0, i_10_308_327_0, i_10_308_329_0,
    i_10_308_330_0, i_10_308_331_0, i_10_308_437_0, i_10_308_443_0,
    i_10_308_462_0, i_10_308_463_0, i_10_308_464_0, i_10_308_467_0,
    i_10_308_514_0, i_10_308_711_0, i_10_308_719_0, i_10_308_748_0,
    i_10_308_749_0, i_10_308_797_0, i_10_308_800_0, i_10_308_990_0,
    i_10_308_991_0, i_10_308_1036_0, i_10_308_1174_0, i_10_308_1235_0,
    i_10_308_1239_0, i_10_308_1240_0, i_10_308_1241_0, i_10_308_1263_0,
    i_10_308_1265_0, i_10_308_1310_0, i_10_308_1342_0, i_10_308_1397_0,
    i_10_308_1610_0, i_10_308_1685_0, i_10_308_1826_0, i_10_308_1908_0,
    i_10_308_1911_0, i_10_308_1916_0, i_10_308_1990_0, i_10_308_1998_0,
    i_10_308_2200_0, i_10_308_2201_0, i_10_308_2335_0, i_10_308_2354_0,
    i_10_308_2407_0, i_10_308_2454_0, i_10_308_2456_0, i_10_308_2470_0,
    i_10_308_2503_0, i_10_308_2516_0, i_10_308_2567_0, i_10_308_2602_0,
    i_10_308_2605_0, i_10_308_2606_0, i_10_308_2629_0, i_10_308_2630_0,
    i_10_308_2661_0, i_10_308_2716_0, i_10_308_2720_0, i_10_308_2722_0,
    i_10_308_2724_0, i_10_308_2729_0, i_10_308_2782_0, i_10_308_2817_0,
    i_10_308_2829_0, i_10_308_2883_0, i_10_308_2953_0, i_10_308_3087_0,
    i_10_308_3088_0, i_10_308_3128_0, i_10_308_3199_0, i_10_308_3201_0,
    i_10_308_3202_0, i_10_308_3267_0, i_10_308_3385_0, i_10_308_3404_0,
    i_10_308_3523_0, i_10_308_3544_0, i_10_308_3557_0, i_10_308_3613_0,
    i_10_308_3614_0, i_10_308_3720_0, i_10_308_3733_0, i_10_308_3837_0,
    i_10_308_3847_0, i_10_308_3856_0, i_10_308_3881_0, i_10_308_4115_0,
    i_10_308_4277_0, i_10_308_4280_0, i_10_308_4284_0, i_10_308_4289_0,
    i_10_308_4351_0, i_10_308_4432_0, i_10_308_4569_0, i_10_308_4570_0;
  output o_10_308_0_0;
  assign o_10_308_0_0 = 0;
endmodule



// Benchmark "kernel_10_309" written by ABC on Sun Jul 19 10:26:25 2020

module kernel_10_309 ( 
    i_10_309_175_0, i_10_309_218_0, i_10_309_244_0, i_10_309_245_0,
    i_10_309_409_0, i_10_309_410_0, i_10_309_436_0, i_10_309_439_0,
    i_10_309_445_0, i_10_309_459_0, i_10_309_467_0, i_10_309_507_0,
    i_10_309_796_0, i_10_309_896_0, i_10_309_990_0, i_10_309_991_0,
    i_10_309_992_0, i_10_309_997_0, i_10_309_1000_0, i_10_309_1003_0,
    i_10_309_1006_0, i_10_309_1042_0, i_10_309_1043_0, i_10_309_1234_0,
    i_10_309_1236_0, i_10_309_1308_0, i_10_309_1309_0, i_10_309_1310_0,
    i_10_309_1312_0, i_10_309_1487_0, i_10_309_1649_0, i_10_309_1652_0,
    i_10_309_1654_0, i_10_309_1690_0, i_10_309_1769_0, i_10_309_1819_0,
    i_10_309_1820_0, i_10_309_1821_0, i_10_309_1824_0, i_10_309_1909_0,
    i_10_309_1916_0, i_10_309_1951_0, i_10_309_1952_0, i_10_309_2185_0,
    i_10_309_2452_0, i_10_309_2453_0, i_10_309_2473_0, i_10_309_2566_0,
    i_10_309_2628_0, i_10_309_2629_0, i_10_309_2704_0, i_10_309_2723_0,
    i_10_309_2724_0, i_10_309_2782_0, i_10_309_2817_0, i_10_309_2829_0,
    i_10_309_2831_0, i_10_309_2832_0, i_10_309_2833_0, i_10_309_2884_0,
    i_10_309_2885_0, i_10_309_2917_0, i_10_309_3034_0, i_10_309_3070_0,
    i_10_309_3151_0, i_10_309_3197_0, i_10_309_3198_0, i_10_309_3200_0,
    i_10_309_3272_0, i_10_309_3326_0, i_10_309_3385_0, i_10_309_3407_0,
    i_10_309_3466_0, i_10_309_3467_0, i_10_309_3499_0, i_10_309_3523_0,
    i_10_309_3585_0, i_10_309_3589_0, i_10_309_3610_0, i_10_309_3613_0,
    i_10_309_3614_0, i_10_309_3616_0, i_10_309_3617_0, i_10_309_3689_0,
    i_10_309_3785_0, i_10_309_3788_0, i_10_309_3835_0, i_10_309_3843_0,
    i_10_309_3986_0, i_10_309_3991_0, i_10_309_3992_0, i_10_309_4113_0,
    i_10_309_4114_0, i_10_309_4115_0, i_10_309_4122_0, i_10_309_4123_0,
    i_10_309_4284_0, i_10_309_4287_0, i_10_309_4563_0, i_10_309_4564_0,
    o_10_309_0_0  );
  input  i_10_309_175_0, i_10_309_218_0, i_10_309_244_0, i_10_309_245_0,
    i_10_309_409_0, i_10_309_410_0, i_10_309_436_0, i_10_309_439_0,
    i_10_309_445_0, i_10_309_459_0, i_10_309_467_0, i_10_309_507_0,
    i_10_309_796_0, i_10_309_896_0, i_10_309_990_0, i_10_309_991_0,
    i_10_309_992_0, i_10_309_997_0, i_10_309_1000_0, i_10_309_1003_0,
    i_10_309_1006_0, i_10_309_1042_0, i_10_309_1043_0, i_10_309_1234_0,
    i_10_309_1236_0, i_10_309_1308_0, i_10_309_1309_0, i_10_309_1310_0,
    i_10_309_1312_0, i_10_309_1487_0, i_10_309_1649_0, i_10_309_1652_0,
    i_10_309_1654_0, i_10_309_1690_0, i_10_309_1769_0, i_10_309_1819_0,
    i_10_309_1820_0, i_10_309_1821_0, i_10_309_1824_0, i_10_309_1909_0,
    i_10_309_1916_0, i_10_309_1951_0, i_10_309_1952_0, i_10_309_2185_0,
    i_10_309_2452_0, i_10_309_2453_0, i_10_309_2473_0, i_10_309_2566_0,
    i_10_309_2628_0, i_10_309_2629_0, i_10_309_2704_0, i_10_309_2723_0,
    i_10_309_2724_0, i_10_309_2782_0, i_10_309_2817_0, i_10_309_2829_0,
    i_10_309_2831_0, i_10_309_2832_0, i_10_309_2833_0, i_10_309_2884_0,
    i_10_309_2885_0, i_10_309_2917_0, i_10_309_3034_0, i_10_309_3070_0,
    i_10_309_3151_0, i_10_309_3197_0, i_10_309_3198_0, i_10_309_3200_0,
    i_10_309_3272_0, i_10_309_3326_0, i_10_309_3385_0, i_10_309_3407_0,
    i_10_309_3466_0, i_10_309_3467_0, i_10_309_3499_0, i_10_309_3523_0,
    i_10_309_3585_0, i_10_309_3589_0, i_10_309_3610_0, i_10_309_3613_0,
    i_10_309_3614_0, i_10_309_3616_0, i_10_309_3617_0, i_10_309_3689_0,
    i_10_309_3785_0, i_10_309_3788_0, i_10_309_3835_0, i_10_309_3843_0,
    i_10_309_3986_0, i_10_309_3991_0, i_10_309_3992_0, i_10_309_4113_0,
    i_10_309_4114_0, i_10_309_4115_0, i_10_309_4122_0, i_10_309_4123_0,
    i_10_309_4284_0, i_10_309_4287_0, i_10_309_4563_0, i_10_309_4564_0;
  output o_10_309_0_0;
  assign o_10_309_0_0 = ~((~i_10_309_1916_0 & ((~i_10_309_175_0 & ((~i_10_309_410_0 & ~i_10_309_796_0 & ~i_10_309_896_0 & ~i_10_309_990_0 & ~i_10_309_1487_0 & ~i_10_309_1649_0 & ~i_10_309_1821_0 & ~i_10_309_2885_0 & ~i_10_309_3070_0 & ~i_10_309_3407_0 & ~i_10_309_3523_0 & ~i_10_309_3613_0) | (~i_10_309_2829_0 & i_10_309_3589_0 & i_10_309_3689_0))) | (~i_10_309_4115_0 & ((~i_10_309_436_0 & ~i_10_309_3197_0 & ~i_10_309_3523_0 & ((~i_10_309_439_0 & ~i_10_309_1042_0 & ~i_10_309_1043_0 & ~i_10_309_1769_0 & ~i_10_309_1821_0 & ~i_10_309_2453_0 & ~i_10_309_2817_0 & ~i_10_309_3617_0) | (~i_10_309_796_0 & ~i_10_309_997_0 & ~i_10_309_1690_0 & ~i_10_309_2829_0 & ~i_10_309_3198_0 & ~i_10_309_3272_0 & ~i_10_309_3785_0))) | (~i_10_309_991_0 & ~i_10_309_1043_0 & ~i_10_309_1236_0 & ~i_10_309_2452_0 & ~i_10_309_2817_0 & ~i_10_309_3385_0 & ~i_10_309_3613_0 & ~i_10_309_3689_0))) | (~i_10_309_991_0 & ~i_10_309_3785_0 & ((~i_10_309_1042_0 & ~i_10_309_1309_0 & ~i_10_309_1312_0 & ~i_10_309_2885_0 & i_10_309_3610_0) | (~i_10_309_992_0 & ~i_10_309_1909_0 & i_10_309_3272_0 & ~i_10_309_3614_0))))) | (~i_10_309_175_0 & ((i_10_309_1006_0 & ~i_10_309_2831_0 & ~i_10_309_3614_0) | (~i_10_309_244_0 & ~i_10_309_245_0 & ~i_10_309_990_0 & ~i_10_309_991_0 & ~i_10_309_1042_0 & ~i_10_309_1043_0 & ~i_10_309_1312_0 & ~i_10_309_1654_0 & ~i_10_309_2833_0 & ~i_10_309_3407_0 & ~i_10_309_3788_0 & ~i_10_309_3986_0 & ~i_10_309_4284_0))) | (~i_10_309_244_0 & ((i_10_309_445_0 & i_10_309_796_0 & ~i_10_309_992_0 & ~i_10_309_1308_0 & ~i_10_309_2723_0 & ~i_10_309_2817_0 & ~i_10_309_2885_0) | (~i_10_309_1310_0 & ~i_10_309_3407_0 & i_10_309_3585_0 & ~i_10_309_3992_0))) | (i_10_309_445_0 & ((~i_10_309_410_0 & ~i_10_309_467_0 & ~i_10_309_1951_0 & ~i_10_309_2884_0 & ~i_10_309_3197_0 & ~i_10_309_3272_0 & ~i_10_309_3385_0) | (~i_10_309_992_0 & ~i_10_309_1649_0 & i_10_309_3589_0))) | (i_10_309_459_0 & ((~i_10_309_245_0 & ~i_10_309_409_0 & ~i_10_309_1310_0 & ~i_10_309_2884_0 & ~i_10_309_3385_0 & ~i_10_309_4115_0) | (~i_10_309_218_0 & ~i_10_309_410_0 & ~i_10_309_990_0 & ~i_10_309_992_0 & ~i_10_309_2885_0 & ~i_10_309_3070_0 & ~i_10_309_3407_0 & ~i_10_309_3785_0 & ~i_10_309_3992_0 & ~i_10_309_4287_0))) | (~i_10_309_991_0 & ((~i_10_309_409_0 & ~i_10_309_3992_0 & ((~i_10_309_997_0 & ~i_10_309_1310_0 & ~i_10_309_2724_0 & ~i_10_309_2833_0 & ~i_10_309_3272_0 & ~i_10_309_3986_0 & ~i_10_309_3991_0 & ~i_10_309_4114_0) | (~i_10_309_896_0 & ~i_10_309_992_0 & ~i_10_309_1309_0 & ~i_10_309_2885_0 & ~i_10_309_3197_0 & ~i_10_309_3614_0 & ~i_10_309_4284_0))) | (~i_10_309_1309_0 & ((~i_10_309_992_0 & ~i_10_309_3614_0 & ((~i_10_309_1043_0 & ~i_10_309_1308_0 & ~i_10_309_1649_0 & ~i_10_309_2629_0 & ~i_10_309_2917_0) | (~i_10_309_1821_0 & ~i_10_309_2452_0 & ~i_10_309_2884_0 & ~i_10_309_3070_0 & ~i_10_309_3272_0))) | (~i_10_309_997_0 & i_10_309_4563_0))) | (i_10_309_2473_0 & ~i_10_309_3617_0 & ~i_10_309_3991_0))) | (~i_10_309_245_0 & ((~i_10_309_992_0 & ((~i_10_309_410_0 & ~i_10_309_1042_0 & ((~i_10_309_997_0 & ~i_10_309_1769_0 & ~i_10_309_1824_0 & ~i_10_309_2628_0 & ~i_10_309_2724_0 & ~i_10_309_2885_0 & ~i_10_309_3788_0 & ~i_10_309_4114_0) | (~i_10_309_459_0 & ~i_10_309_1909_0 & ~i_10_309_2452_0 & ~i_10_309_2453_0 & ~i_10_309_2833_0 & ~i_10_309_3585_0 & ~i_10_309_3614_0 & ~i_10_309_4113_0 & ~i_10_309_4122_0))) | (i_10_309_2782_0 & ~i_10_309_3613_0 & ~i_10_309_4115_0))) | (~i_10_309_2704_0 & i_10_309_3034_0 & ~i_10_309_3197_0) | (~i_10_309_2452_0 & ~i_10_309_2628_0 & ~i_10_309_2723_0 & ~i_10_309_2829_0 & ~i_10_309_3614_0 & ~i_10_309_3992_0))) | (~i_10_309_990_0 & ((i_10_309_1824_0 & ~i_10_309_2832_0 & ~i_10_309_3070_0 & i_10_309_3613_0 & ~i_10_309_3614_0 & ~i_10_309_3617_0) | (~i_10_309_997_0 & i_10_309_1654_0 & ~i_10_309_1824_0 & ~i_10_309_2723_0 & ~i_10_309_3385_0 & ~i_10_309_3610_0 & ~i_10_309_3785_0 & ~i_10_309_3986_0))) | (~i_10_309_992_0 & ((~i_10_309_467_0 & ~i_10_309_796_0 & ~i_10_309_1312_0 & ~i_10_309_2723_0 & ~i_10_309_2832_0 & ~i_10_309_2917_0 & ~i_10_309_3986_0 & ~i_10_309_4114_0) | (~i_10_309_445_0 & ~i_10_309_1308_0 & ~i_10_309_2884_0 & ~i_10_309_2885_0 & ~i_10_309_3523_0 & i_10_309_4284_0))) | (~i_10_309_3992_0 & ((i_10_309_1821_0 & i_10_309_1952_0) | (i_10_309_796_0 & ~i_10_309_896_0 & ~i_10_309_1310_0 & ~i_10_309_2704_0 & ~i_10_309_2829_0 & i_10_309_2833_0 & ~i_10_309_3617_0))) | (i_10_309_2628_0 & ~i_10_309_2629_0 & ~i_10_309_3070_0 & i_10_309_3843_0 & ~i_10_309_4115_0));
endmodule



// Benchmark "kernel_10_310" written by ABC on Sun Jul 19 10:26:26 2020

module kernel_10_310 ( 
    i_10_310_33_0, i_10_310_247_0, i_10_310_248_0, i_10_310_249_0,
    i_10_310_282_0, i_10_310_283_0, i_10_310_287_0, i_10_310_430_0,
    i_10_310_435_0, i_10_310_436_0, i_10_310_438_0, i_10_310_444_0,
    i_10_310_445_0, i_10_310_449_0, i_10_310_462_0, i_10_310_465_0,
    i_10_310_466_0, i_10_310_517_0, i_10_310_747_0, i_10_310_748_0,
    i_10_310_754_0, i_10_310_795_0, i_10_310_796_0, i_10_310_956_0,
    i_10_310_959_0, i_10_310_1233_0, i_10_310_1243_0, i_10_310_1246_0,
    i_10_310_1267_0, i_10_310_1306_0, i_10_310_1311_0, i_10_310_1360_0,
    i_10_310_1442_0, i_10_310_1578_0, i_10_310_1651_0, i_10_310_1654_0,
    i_10_310_1684_0, i_10_310_1689_0, i_10_310_1823_0, i_10_310_2254_0,
    i_10_310_2304_0, i_10_310_2310_0, i_10_310_2311_0, i_10_310_2312_0,
    i_10_310_2350_0, i_10_310_2454_0, i_10_310_2473_0, i_10_310_2474_0,
    i_10_310_2628_0, i_10_310_2631_0, i_10_310_2632_0, i_10_310_2634_0,
    i_10_310_2705_0, i_10_310_2727_0, i_10_310_2728_0, i_10_310_2821_0,
    i_10_310_2881_0, i_10_310_2887_0, i_10_310_2888_0, i_10_310_2913_0,
    i_10_310_2916_0, i_10_310_2923_0, i_10_310_3033_0, i_10_310_3034_0,
    i_10_310_3036_0, i_10_310_3037_0, i_10_310_3038_0, i_10_310_3040_0,
    i_10_310_3041_0, i_10_310_3074_0, i_10_310_3196_0, i_10_310_3197_0,
    i_10_310_3198_0, i_10_310_3202_0, i_10_310_3280_0, i_10_310_3387_0,
    i_10_310_3390_0, i_10_310_3392_0, i_10_310_3402_0, i_10_310_3403_0,
    i_10_310_3469_0, i_10_310_3493_0, i_10_310_3497_0, i_10_310_3614_0,
    i_10_310_3615_0, i_10_310_3649_0, i_10_310_3727_0, i_10_310_3780_0,
    i_10_310_3781_0, i_10_310_3837_0, i_10_310_3860_0, i_10_310_3906_0,
    i_10_310_3907_0, i_10_310_3972_0, i_10_310_3994_0, i_10_310_4113_0,
    i_10_310_4278_0, i_10_310_4279_0, i_10_310_4462_0, i_10_310_4525_0,
    o_10_310_0_0  );
  input  i_10_310_33_0, i_10_310_247_0, i_10_310_248_0, i_10_310_249_0,
    i_10_310_282_0, i_10_310_283_0, i_10_310_287_0, i_10_310_430_0,
    i_10_310_435_0, i_10_310_436_0, i_10_310_438_0, i_10_310_444_0,
    i_10_310_445_0, i_10_310_449_0, i_10_310_462_0, i_10_310_465_0,
    i_10_310_466_0, i_10_310_517_0, i_10_310_747_0, i_10_310_748_0,
    i_10_310_754_0, i_10_310_795_0, i_10_310_796_0, i_10_310_956_0,
    i_10_310_959_0, i_10_310_1233_0, i_10_310_1243_0, i_10_310_1246_0,
    i_10_310_1267_0, i_10_310_1306_0, i_10_310_1311_0, i_10_310_1360_0,
    i_10_310_1442_0, i_10_310_1578_0, i_10_310_1651_0, i_10_310_1654_0,
    i_10_310_1684_0, i_10_310_1689_0, i_10_310_1823_0, i_10_310_2254_0,
    i_10_310_2304_0, i_10_310_2310_0, i_10_310_2311_0, i_10_310_2312_0,
    i_10_310_2350_0, i_10_310_2454_0, i_10_310_2473_0, i_10_310_2474_0,
    i_10_310_2628_0, i_10_310_2631_0, i_10_310_2632_0, i_10_310_2634_0,
    i_10_310_2705_0, i_10_310_2727_0, i_10_310_2728_0, i_10_310_2821_0,
    i_10_310_2881_0, i_10_310_2887_0, i_10_310_2888_0, i_10_310_2913_0,
    i_10_310_2916_0, i_10_310_2923_0, i_10_310_3033_0, i_10_310_3034_0,
    i_10_310_3036_0, i_10_310_3037_0, i_10_310_3038_0, i_10_310_3040_0,
    i_10_310_3041_0, i_10_310_3074_0, i_10_310_3196_0, i_10_310_3197_0,
    i_10_310_3198_0, i_10_310_3202_0, i_10_310_3280_0, i_10_310_3387_0,
    i_10_310_3390_0, i_10_310_3392_0, i_10_310_3402_0, i_10_310_3403_0,
    i_10_310_3469_0, i_10_310_3493_0, i_10_310_3497_0, i_10_310_3614_0,
    i_10_310_3615_0, i_10_310_3649_0, i_10_310_3727_0, i_10_310_3780_0,
    i_10_310_3781_0, i_10_310_3837_0, i_10_310_3860_0, i_10_310_3906_0,
    i_10_310_3907_0, i_10_310_3972_0, i_10_310_3994_0, i_10_310_4113_0,
    i_10_310_4278_0, i_10_310_4279_0, i_10_310_4462_0, i_10_310_4525_0;
  output o_10_310_0_0;
  assign o_10_310_0_0 = 0;
endmodule



// Benchmark "kernel_10_311" written by ABC on Sun Jul 19 10:26:27 2020

module kernel_10_311 ( 
    i_10_311_86_0, i_10_311_387_0, i_10_311_388_0, i_10_311_409_0,
    i_10_311_423_0, i_10_311_433_0, i_10_311_461_0, i_10_311_496_0,
    i_10_311_514_0, i_10_311_693_0, i_10_311_694_0, i_10_311_714_0,
    i_10_311_733_0, i_10_311_734_0, i_10_311_735_0, i_10_311_796_0,
    i_10_311_799_0, i_10_311_800_0, i_10_311_901_0, i_10_311_993_0,
    i_10_311_999_0, i_10_311_1037_0, i_10_311_1237_0, i_10_311_1238_0,
    i_10_311_1239_0, i_10_311_1278_0, i_10_311_1307_0, i_10_311_1341_0,
    i_10_311_1342_0, i_10_311_1343_0, i_10_311_1354_0, i_10_311_1549_0,
    i_10_311_1576_0, i_10_311_1621_0, i_10_311_1650_0, i_10_311_1651_0,
    i_10_311_1685_0, i_10_311_1714_0, i_10_311_1818_0, i_10_311_1825_0,
    i_10_311_1826_0, i_10_311_1908_0, i_10_311_1909_0, i_10_311_1910_0,
    i_10_311_1944_0, i_10_311_2080_0, i_10_311_2263_0, i_10_311_2312_0,
    i_10_311_2327_0, i_10_311_2349_0, i_10_311_2350_0, i_10_311_2351_0,
    i_10_311_2383_0, i_10_311_2448_0, i_10_311_2454_0, i_10_311_2458_0,
    i_10_311_2566_0, i_10_311_2632_0, i_10_311_2635_0, i_10_311_2636_0,
    i_10_311_2720_0, i_10_311_2721_0, i_10_311_2820_0, i_10_311_2821_0,
    i_10_311_2882_0, i_10_311_2884_0, i_10_311_2885_0, i_10_311_2983_0,
    i_10_311_3197_0, i_10_311_3276_0, i_10_311_3277_0, i_10_311_3385_0,
    i_10_311_3613_0, i_10_311_3614_0, i_10_311_3615_0, i_10_311_3616_0,
    i_10_311_3650_0, i_10_311_3837_0, i_10_311_3840_0, i_10_311_3842_0,
    i_10_311_3853_0, i_10_311_3856_0, i_10_311_3859_0, i_10_311_3888_0,
    i_10_311_3889_0, i_10_311_3891_0, i_10_311_3979_0, i_10_311_3988_0,
    i_10_311_4027_0, i_10_311_4113_0, i_10_311_4154_0, i_10_311_4176_0,
    i_10_311_4177_0, i_10_311_4216_0, i_10_311_4275_0, i_10_311_4288_0,
    i_10_311_4291_0, i_10_311_4568_0, i_10_311_4587_0, i_10_311_4592_0,
    o_10_311_0_0  );
  input  i_10_311_86_0, i_10_311_387_0, i_10_311_388_0, i_10_311_409_0,
    i_10_311_423_0, i_10_311_433_0, i_10_311_461_0, i_10_311_496_0,
    i_10_311_514_0, i_10_311_693_0, i_10_311_694_0, i_10_311_714_0,
    i_10_311_733_0, i_10_311_734_0, i_10_311_735_0, i_10_311_796_0,
    i_10_311_799_0, i_10_311_800_0, i_10_311_901_0, i_10_311_993_0,
    i_10_311_999_0, i_10_311_1037_0, i_10_311_1237_0, i_10_311_1238_0,
    i_10_311_1239_0, i_10_311_1278_0, i_10_311_1307_0, i_10_311_1341_0,
    i_10_311_1342_0, i_10_311_1343_0, i_10_311_1354_0, i_10_311_1549_0,
    i_10_311_1576_0, i_10_311_1621_0, i_10_311_1650_0, i_10_311_1651_0,
    i_10_311_1685_0, i_10_311_1714_0, i_10_311_1818_0, i_10_311_1825_0,
    i_10_311_1826_0, i_10_311_1908_0, i_10_311_1909_0, i_10_311_1910_0,
    i_10_311_1944_0, i_10_311_2080_0, i_10_311_2263_0, i_10_311_2312_0,
    i_10_311_2327_0, i_10_311_2349_0, i_10_311_2350_0, i_10_311_2351_0,
    i_10_311_2383_0, i_10_311_2448_0, i_10_311_2454_0, i_10_311_2458_0,
    i_10_311_2566_0, i_10_311_2632_0, i_10_311_2635_0, i_10_311_2636_0,
    i_10_311_2720_0, i_10_311_2721_0, i_10_311_2820_0, i_10_311_2821_0,
    i_10_311_2882_0, i_10_311_2884_0, i_10_311_2885_0, i_10_311_2983_0,
    i_10_311_3197_0, i_10_311_3276_0, i_10_311_3277_0, i_10_311_3385_0,
    i_10_311_3613_0, i_10_311_3614_0, i_10_311_3615_0, i_10_311_3616_0,
    i_10_311_3650_0, i_10_311_3837_0, i_10_311_3840_0, i_10_311_3842_0,
    i_10_311_3853_0, i_10_311_3856_0, i_10_311_3859_0, i_10_311_3888_0,
    i_10_311_3889_0, i_10_311_3891_0, i_10_311_3979_0, i_10_311_3988_0,
    i_10_311_4027_0, i_10_311_4113_0, i_10_311_4154_0, i_10_311_4176_0,
    i_10_311_4177_0, i_10_311_4216_0, i_10_311_4275_0, i_10_311_4288_0,
    i_10_311_4291_0, i_10_311_4568_0, i_10_311_4587_0, i_10_311_4592_0;
  output o_10_311_0_0;
  assign o_10_311_0_0 = 0;
endmodule



// Benchmark "kernel_10_312" written by ABC on Sun Jul 19 10:26:27 2020

module kernel_10_312 ( 
    i_10_312_118_0, i_10_312_218_0, i_10_312_282_0, i_10_312_283_0,
    i_10_312_287_0, i_10_312_316_0, i_10_312_407_0, i_10_312_409_0,
    i_10_312_432_0, i_10_312_433_0, i_10_312_434_0, i_10_312_435_0,
    i_10_312_437_0, i_10_312_448_0, i_10_312_799_0, i_10_312_800_0,
    i_10_312_962_0, i_10_312_1029_0, i_10_312_1030_0, i_10_312_1033_0,
    i_10_312_1241_0, i_10_312_1309_0, i_10_312_1310_0, i_10_312_1365_0,
    i_10_312_1556_0, i_10_312_1650_0, i_10_312_1651_0, i_10_312_1654_0,
    i_10_312_1684_0, i_10_312_1685_0, i_10_312_1821_0, i_10_312_1825_0,
    i_10_312_1996_0, i_10_312_2179_0, i_10_312_2349_0, i_10_312_2350_0,
    i_10_312_2351_0, i_10_312_2361_0, i_10_312_2364_0, i_10_312_2365_0,
    i_10_312_2407_0, i_10_312_2453_0, i_10_312_2458_0, i_10_312_2461_0,
    i_10_312_2463_0, i_10_312_2467_0, i_10_312_2474_0, i_10_312_2571_0,
    i_10_312_2611_0, i_10_312_2634_0, i_10_312_2657_0, i_10_312_2661_0,
    i_10_312_2701_0, i_10_312_2704_0, i_10_312_2707_0, i_10_312_2714_0,
    i_10_312_2721_0, i_10_312_2731_0, i_10_312_2733_0, i_10_312_2788_0,
    i_10_312_2821_0, i_10_312_2824_0, i_10_312_2825_0, i_10_312_2831_0,
    i_10_312_2881_0, i_10_312_2882_0, i_10_312_2919_0, i_10_312_3036_0,
    i_10_312_3037_0, i_10_312_3038_0, i_10_312_3041_0, i_10_312_3050_0,
    i_10_312_3088_0, i_10_312_3196_0, i_10_312_3199_0, i_10_312_3391_0,
    i_10_312_3403_0, i_10_312_3404_0, i_10_312_3583_0, i_10_312_3613_0,
    i_10_312_3614_0, i_10_312_3648_0, i_10_312_3786_0, i_10_312_3839_0,
    i_10_312_3840_0, i_10_312_3843_0, i_10_312_3855_0, i_10_312_3856_0,
    i_10_312_3857_0, i_10_312_3858_0, i_10_312_3859_0, i_10_312_3994_0,
    i_10_312_4128_0, i_10_312_4168_0, i_10_312_4170_0, i_10_312_4172_0,
    i_10_312_4267_0, i_10_312_4273_0, i_10_312_4565_0, i_10_312_4570_0,
    o_10_312_0_0  );
  input  i_10_312_118_0, i_10_312_218_0, i_10_312_282_0, i_10_312_283_0,
    i_10_312_287_0, i_10_312_316_0, i_10_312_407_0, i_10_312_409_0,
    i_10_312_432_0, i_10_312_433_0, i_10_312_434_0, i_10_312_435_0,
    i_10_312_437_0, i_10_312_448_0, i_10_312_799_0, i_10_312_800_0,
    i_10_312_962_0, i_10_312_1029_0, i_10_312_1030_0, i_10_312_1033_0,
    i_10_312_1241_0, i_10_312_1309_0, i_10_312_1310_0, i_10_312_1365_0,
    i_10_312_1556_0, i_10_312_1650_0, i_10_312_1651_0, i_10_312_1654_0,
    i_10_312_1684_0, i_10_312_1685_0, i_10_312_1821_0, i_10_312_1825_0,
    i_10_312_1996_0, i_10_312_2179_0, i_10_312_2349_0, i_10_312_2350_0,
    i_10_312_2351_0, i_10_312_2361_0, i_10_312_2364_0, i_10_312_2365_0,
    i_10_312_2407_0, i_10_312_2453_0, i_10_312_2458_0, i_10_312_2461_0,
    i_10_312_2463_0, i_10_312_2467_0, i_10_312_2474_0, i_10_312_2571_0,
    i_10_312_2611_0, i_10_312_2634_0, i_10_312_2657_0, i_10_312_2661_0,
    i_10_312_2701_0, i_10_312_2704_0, i_10_312_2707_0, i_10_312_2714_0,
    i_10_312_2721_0, i_10_312_2731_0, i_10_312_2733_0, i_10_312_2788_0,
    i_10_312_2821_0, i_10_312_2824_0, i_10_312_2825_0, i_10_312_2831_0,
    i_10_312_2881_0, i_10_312_2882_0, i_10_312_2919_0, i_10_312_3036_0,
    i_10_312_3037_0, i_10_312_3038_0, i_10_312_3041_0, i_10_312_3050_0,
    i_10_312_3088_0, i_10_312_3196_0, i_10_312_3199_0, i_10_312_3391_0,
    i_10_312_3403_0, i_10_312_3404_0, i_10_312_3583_0, i_10_312_3613_0,
    i_10_312_3614_0, i_10_312_3648_0, i_10_312_3786_0, i_10_312_3839_0,
    i_10_312_3840_0, i_10_312_3843_0, i_10_312_3855_0, i_10_312_3856_0,
    i_10_312_3857_0, i_10_312_3858_0, i_10_312_3859_0, i_10_312_3994_0,
    i_10_312_4128_0, i_10_312_4168_0, i_10_312_4170_0, i_10_312_4172_0,
    i_10_312_4267_0, i_10_312_4273_0, i_10_312_4565_0, i_10_312_4570_0;
  output o_10_312_0_0;
  assign o_10_312_0_0 = 0;
endmodule



// Benchmark "kernel_10_313" written by ABC on Sun Jul 19 10:26:28 2020

module kernel_10_313 ( 
    i_10_313_48_0, i_10_313_156_0, i_10_313_216_0, i_10_313_223_0,
    i_10_313_252_0, i_10_313_327_0, i_10_313_387_0, i_10_313_408_0,
    i_10_313_409_0, i_10_313_410_0, i_10_313_445_0, i_10_313_463_0,
    i_10_313_498_0, i_10_313_504_0, i_10_313_516_0, i_10_313_531_0,
    i_10_313_532_0, i_10_313_748_0, i_10_313_750_0, i_10_313_753_0,
    i_10_313_867_0, i_10_313_906_0, i_10_313_957_0, i_10_313_958_0,
    i_10_313_990_0, i_10_313_1084_0, i_10_313_1134_0, i_10_313_1162_0,
    i_10_313_1218_0, i_10_313_1221_0, i_10_313_1236_0, i_10_313_1238_0,
    i_10_313_1262_0, i_10_313_1263_0, i_10_313_1266_0, i_10_313_1290_0,
    i_10_313_1310_0, i_10_313_1312_0, i_10_313_1347_0, i_10_313_1348_0,
    i_10_313_1398_0, i_10_313_1485_0, i_10_313_1545_0, i_10_313_1655_0,
    i_10_313_1683_0, i_10_313_1690_0, i_10_313_1822_0, i_10_313_1848_0,
    i_10_313_1947_0, i_10_313_1999_0, i_10_313_2361_0, i_10_313_2380_0,
    i_10_313_2452_0, i_10_313_2541_0, i_10_313_2577_0, i_10_313_2632_0,
    i_10_313_2634_0, i_10_313_2657_0, i_10_313_2660_0, i_10_313_2661_0,
    i_10_313_2677_0, i_10_313_2723_0, i_10_313_2728_0, i_10_313_2817_0,
    i_10_313_2881_0, i_10_313_2979_0, i_10_313_2983_0, i_10_313_3038_0,
    i_10_313_3040_0, i_10_313_3231_0, i_10_313_3232_0, i_10_313_3276_0,
    i_10_313_3277_0, i_10_313_3279_0, i_10_313_3281_0, i_10_313_3283_0,
    i_10_313_3388_0, i_10_313_3391_0, i_10_313_3466_0, i_10_313_3467_0,
    i_10_313_3496_0, i_10_313_3522_0, i_10_313_3613_0, i_10_313_3614_0,
    i_10_313_3648_0, i_10_313_3684_0, i_10_313_3782_0, i_10_313_3785_0,
    i_10_313_3786_0, i_10_313_3852_0, i_10_313_3910_0, i_10_313_3979_0,
    i_10_313_4113_0, i_10_313_4114_0, i_10_313_4266_0, i_10_313_4270_0,
    i_10_313_4275_0, i_10_313_4290_0, i_10_313_4291_0, i_10_313_4584_0,
    o_10_313_0_0  );
  input  i_10_313_48_0, i_10_313_156_0, i_10_313_216_0, i_10_313_223_0,
    i_10_313_252_0, i_10_313_327_0, i_10_313_387_0, i_10_313_408_0,
    i_10_313_409_0, i_10_313_410_0, i_10_313_445_0, i_10_313_463_0,
    i_10_313_498_0, i_10_313_504_0, i_10_313_516_0, i_10_313_531_0,
    i_10_313_532_0, i_10_313_748_0, i_10_313_750_0, i_10_313_753_0,
    i_10_313_867_0, i_10_313_906_0, i_10_313_957_0, i_10_313_958_0,
    i_10_313_990_0, i_10_313_1084_0, i_10_313_1134_0, i_10_313_1162_0,
    i_10_313_1218_0, i_10_313_1221_0, i_10_313_1236_0, i_10_313_1238_0,
    i_10_313_1262_0, i_10_313_1263_0, i_10_313_1266_0, i_10_313_1290_0,
    i_10_313_1310_0, i_10_313_1312_0, i_10_313_1347_0, i_10_313_1348_0,
    i_10_313_1398_0, i_10_313_1485_0, i_10_313_1545_0, i_10_313_1655_0,
    i_10_313_1683_0, i_10_313_1690_0, i_10_313_1822_0, i_10_313_1848_0,
    i_10_313_1947_0, i_10_313_1999_0, i_10_313_2361_0, i_10_313_2380_0,
    i_10_313_2452_0, i_10_313_2541_0, i_10_313_2577_0, i_10_313_2632_0,
    i_10_313_2634_0, i_10_313_2657_0, i_10_313_2660_0, i_10_313_2661_0,
    i_10_313_2677_0, i_10_313_2723_0, i_10_313_2728_0, i_10_313_2817_0,
    i_10_313_2881_0, i_10_313_2979_0, i_10_313_2983_0, i_10_313_3038_0,
    i_10_313_3040_0, i_10_313_3231_0, i_10_313_3232_0, i_10_313_3276_0,
    i_10_313_3277_0, i_10_313_3279_0, i_10_313_3281_0, i_10_313_3283_0,
    i_10_313_3388_0, i_10_313_3391_0, i_10_313_3466_0, i_10_313_3467_0,
    i_10_313_3496_0, i_10_313_3522_0, i_10_313_3613_0, i_10_313_3614_0,
    i_10_313_3648_0, i_10_313_3684_0, i_10_313_3782_0, i_10_313_3785_0,
    i_10_313_3786_0, i_10_313_3852_0, i_10_313_3910_0, i_10_313_3979_0,
    i_10_313_4113_0, i_10_313_4114_0, i_10_313_4266_0, i_10_313_4270_0,
    i_10_313_4275_0, i_10_313_4290_0, i_10_313_4291_0, i_10_313_4584_0;
  output o_10_313_0_0;
  assign o_10_313_0_0 = 0;
endmodule



// Benchmark "kernel_10_314" written by ABC on Sun Jul 19 10:26:29 2020

module kernel_10_314 ( 
    i_10_314_174_0, i_10_314_179_0, i_10_314_220_0, i_10_314_221_0,
    i_10_314_224_0, i_10_314_283_0, i_10_314_321_0, i_10_314_371_0,
    i_10_314_501_0, i_10_314_734_0, i_10_314_799_0, i_10_314_957_0,
    i_10_314_958_0, i_10_314_1054_0, i_10_314_1234_0, i_10_314_1236_0,
    i_10_314_1237_0, i_10_314_1431_0, i_10_314_1432_0, i_10_314_1541_0,
    i_10_314_1544_0, i_10_314_1578_0, i_10_314_1626_0, i_10_314_1635_0,
    i_10_314_1651_0, i_10_314_1655_0, i_10_314_1683_0, i_10_314_1684_0,
    i_10_314_1689_0, i_10_314_1690_0, i_10_314_1714_0, i_10_314_1735_0,
    i_10_314_1804_0, i_10_314_1805_0, i_10_314_1807_0, i_10_314_2003_0,
    i_10_314_2019_0, i_10_314_2029_0, i_10_314_2200_0, i_10_314_2201_0,
    i_10_314_2330_0, i_10_314_2353_0, i_10_314_2365_0, i_10_314_2366_0,
    i_10_314_2452_0, i_10_314_2481_0, i_10_314_2599_0, i_10_314_2605_0,
    i_10_314_2628_0, i_10_314_2631_0, i_10_314_2716_0, i_10_314_2718_0,
    i_10_314_2730_0, i_10_314_2731_0, i_10_314_2732_0, i_10_314_2733_0,
    i_10_314_2734_0, i_10_314_2757_0, i_10_314_2886_0, i_10_314_2966_0,
    i_10_314_2968_0, i_10_314_3162_0, i_10_314_3269_0, i_10_314_3278_0,
    i_10_314_3280_0, i_10_314_3282_0, i_10_314_3283_0, i_10_314_3284_0,
    i_10_314_3315_0, i_10_314_3387_0, i_10_314_3410_0, i_10_314_3430_0,
    i_10_314_3468_0, i_10_314_3469_0, i_10_314_3525_0, i_10_314_3545_0,
    i_10_314_3583_0, i_10_314_3612_0, i_10_314_3646_0, i_10_314_3648_0,
    i_10_314_3649_0, i_10_314_3811_0, i_10_314_3841_0, i_10_314_3855_0,
    i_10_314_3913_0, i_10_314_3988_0, i_10_314_4051_0, i_10_314_4099_0,
    i_10_314_4113_0, i_10_314_4114_0, i_10_314_4121_0, i_10_314_4129_0,
    i_10_314_4130_0, i_10_314_4215_0, i_10_314_4276_0, i_10_314_4291_0,
    i_10_314_4306_0, i_10_314_4565_0, i_10_314_4567_0, i_10_314_4568_0,
    o_10_314_0_0  );
  input  i_10_314_174_0, i_10_314_179_0, i_10_314_220_0, i_10_314_221_0,
    i_10_314_224_0, i_10_314_283_0, i_10_314_321_0, i_10_314_371_0,
    i_10_314_501_0, i_10_314_734_0, i_10_314_799_0, i_10_314_957_0,
    i_10_314_958_0, i_10_314_1054_0, i_10_314_1234_0, i_10_314_1236_0,
    i_10_314_1237_0, i_10_314_1431_0, i_10_314_1432_0, i_10_314_1541_0,
    i_10_314_1544_0, i_10_314_1578_0, i_10_314_1626_0, i_10_314_1635_0,
    i_10_314_1651_0, i_10_314_1655_0, i_10_314_1683_0, i_10_314_1684_0,
    i_10_314_1689_0, i_10_314_1690_0, i_10_314_1714_0, i_10_314_1735_0,
    i_10_314_1804_0, i_10_314_1805_0, i_10_314_1807_0, i_10_314_2003_0,
    i_10_314_2019_0, i_10_314_2029_0, i_10_314_2200_0, i_10_314_2201_0,
    i_10_314_2330_0, i_10_314_2353_0, i_10_314_2365_0, i_10_314_2366_0,
    i_10_314_2452_0, i_10_314_2481_0, i_10_314_2599_0, i_10_314_2605_0,
    i_10_314_2628_0, i_10_314_2631_0, i_10_314_2716_0, i_10_314_2718_0,
    i_10_314_2730_0, i_10_314_2731_0, i_10_314_2732_0, i_10_314_2733_0,
    i_10_314_2734_0, i_10_314_2757_0, i_10_314_2886_0, i_10_314_2966_0,
    i_10_314_2968_0, i_10_314_3162_0, i_10_314_3269_0, i_10_314_3278_0,
    i_10_314_3280_0, i_10_314_3282_0, i_10_314_3283_0, i_10_314_3284_0,
    i_10_314_3315_0, i_10_314_3387_0, i_10_314_3410_0, i_10_314_3430_0,
    i_10_314_3468_0, i_10_314_3469_0, i_10_314_3525_0, i_10_314_3545_0,
    i_10_314_3583_0, i_10_314_3612_0, i_10_314_3646_0, i_10_314_3648_0,
    i_10_314_3649_0, i_10_314_3811_0, i_10_314_3841_0, i_10_314_3855_0,
    i_10_314_3913_0, i_10_314_3988_0, i_10_314_4051_0, i_10_314_4099_0,
    i_10_314_4113_0, i_10_314_4114_0, i_10_314_4121_0, i_10_314_4129_0,
    i_10_314_4130_0, i_10_314_4215_0, i_10_314_4276_0, i_10_314_4291_0,
    i_10_314_4306_0, i_10_314_4565_0, i_10_314_4567_0, i_10_314_4568_0;
  output o_10_314_0_0;
  assign o_10_314_0_0 = 0;
endmodule



// Benchmark "kernel_10_315" written by ABC on Sun Jul 19 10:26:31 2020

module kernel_10_315 ( 
    i_10_315_173_0, i_10_315_328_0, i_10_315_410_0, i_10_315_427_0,
    i_10_315_443_0, i_10_315_445_0, i_10_315_463_0, i_10_315_466_0,
    i_10_315_515_0, i_10_315_716_0, i_10_315_892_0, i_10_315_958_0,
    i_10_315_1027_0, i_10_315_1028_0, i_10_315_1237_0, i_10_315_1244_0,
    i_10_315_1246_0, i_10_315_1249_0, i_10_315_1308_0, i_10_315_1310_0,
    i_10_315_1312_0, i_10_315_1313_0, i_10_315_1541_0, i_10_315_1631_0,
    i_10_315_1652_0, i_10_315_1675_0, i_10_315_1676_0, i_10_315_1685_0,
    i_10_315_1687_0, i_10_315_1691_0, i_10_315_1820_0, i_10_315_1825_0,
    i_10_315_1910_0, i_10_315_1916_0, i_10_315_2026_0, i_10_315_2027_0,
    i_10_315_2243_0, i_10_315_2378_0, i_10_315_2468_0, i_10_315_2566_0,
    i_10_315_2567_0, i_10_315_2608_0, i_10_315_2635_0, i_10_315_2701_0,
    i_10_315_2711_0, i_10_315_2719_0, i_10_315_2720_0, i_10_315_2722_0,
    i_10_315_2723_0, i_10_315_2727_0, i_10_315_2728_0, i_10_315_2729_0,
    i_10_315_2731_0, i_10_315_2786_0, i_10_315_2829_0, i_10_315_2917_0,
    i_10_315_2919_0, i_10_315_2920_0, i_10_315_2924_0, i_10_315_2980_0,
    i_10_315_3042_0, i_10_315_3044_0, i_10_315_3277_0, i_10_315_3281_0,
    i_10_315_3385_0, i_10_315_3387_0, i_10_315_3389_0, i_10_315_3392_0,
    i_10_315_3539_0, i_10_315_3542_0, i_10_315_3586_0, i_10_315_3611_0,
    i_10_315_3646_0, i_10_315_3727_0, i_10_315_3787_0, i_10_315_3839_0,
    i_10_315_3843_0, i_10_315_3844_0, i_10_315_3846_0, i_10_315_3848_0,
    i_10_315_3851_0, i_10_315_3852_0, i_10_315_3855_0, i_10_315_3857_0,
    i_10_315_3906_0, i_10_315_3908_0, i_10_315_3979_0, i_10_315_4213_0,
    i_10_315_4216_0, i_10_315_4268_0, i_10_315_4271_0, i_10_315_4284_0,
    i_10_315_4285_0, i_10_315_4286_0, i_10_315_4288_0, i_10_315_4289_0,
    i_10_315_4290_0, i_10_315_4563_0, i_10_315_4564_0, i_10_315_4566_0,
    o_10_315_0_0  );
  input  i_10_315_173_0, i_10_315_328_0, i_10_315_410_0, i_10_315_427_0,
    i_10_315_443_0, i_10_315_445_0, i_10_315_463_0, i_10_315_466_0,
    i_10_315_515_0, i_10_315_716_0, i_10_315_892_0, i_10_315_958_0,
    i_10_315_1027_0, i_10_315_1028_0, i_10_315_1237_0, i_10_315_1244_0,
    i_10_315_1246_0, i_10_315_1249_0, i_10_315_1308_0, i_10_315_1310_0,
    i_10_315_1312_0, i_10_315_1313_0, i_10_315_1541_0, i_10_315_1631_0,
    i_10_315_1652_0, i_10_315_1675_0, i_10_315_1676_0, i_10_315_1685_0,
    i_10_315_1687_0, i_10_315_1691_0, i_10_315_1820_0, i_10_315_1825_0,
    i_10_315_1910_0, i_10_315_1916_0, i_10_315_2026_0, i_10_315_2027_0,
    i_10_315_2243_0, i_10_315_2378_0, i_10_315_2468_0, i_10_315_2566_0,
    i_10_315_2567_0, i_10_315_2608_0, i_10_315_2635_0, i_10_315_2701_0,
    i_10_315_2711_0, i_10_315_2719_0, i_10_315_2720_0, i_10_315_2722_0,
    i_10_315_2723_0, i_10_315_2727_0, i_10_315_2728_0, i_10_315_2729_0,
    i_10_315_2731_0, i_10_315_2786_0, i_10_315_2829_0, i_10_315_2917_0,
    i_10_315_2919_0, i_10_315_2920_0, i_10_315_2924_0, i_10_315_2980_0,
    i_10_315_3042_0, i_10_315_3044_0, i_10_315_3277_0, i_10_315_3281_0,
    i_10_315_3385_0, i_10_315_3387_0, i_10_315_3389_0, i_10_315_3392_0,
    i_10_315_3539_0, i_10_315_3542_0, i_10_315_3586_0, i_10_315_3611_0,
    i_10_315_3646_0, i_10_315_3727_0, i_10_315_3787_0, i_10_315_3839_0,
    i_10_315_3843_0, i_10_315_3844_0, i_10_315_3846_0, i_10_315_3848_0,
    i_10_315_3851_0, i_10_315_3852_0, i_10_315_3855_0, i_10_315_3857_0,
    i_10_315_3906_0, i_10_315_3908_0, i_10_315_3979_0, i_10_315_4213_0,
    i_10_315_4216_0, i_10_315_4268_0, i_10_315_4271_0, i_10_315_4284_0,
    i_10_315_4285_0, i_10_315_4286_0, i_10_315_4288_0, i_10_315_4289_0,
    i_10_315_4290_0, i_10_315_4563_0, i_10_315_4564_0, i_10_315_4566_0;
  output o_10_315_0_0;
  assign o_10_315_0_0 = ~((~i_10_315_173_0 & ~i_10_315_1027_0 & ~i_10_315_1685_0 & ((~i_10_315_1244_0 & ~i_10_315_2723_0 & ~i_10_315_3281_0 & ~i_10_315_3844_0) | (~i_10_315_2468_0 & ~i_10_315_2731_0 & ~i_10_315_3044_0 & ~i_10_315_3611_0 & ~i_10_315_3851_0 & ~i_10_315_3906_0 & ~i_10_315_4566_0))) | (~i_10_315_3846_0 & ((~i_10_315_515_0 & ((~i_10_315_716_0 & ~i_10_315_1028_0 & ~i_10_315_1687_0 & ~i_10_315_1820_0 & ~i_10_315_1916_0 & ~i_10_315_2468_0 & ~i_10_315_2727_0) | (~i_10_315_328_0 & ~i_10_315_892_0 & ~i_10_315_3389_0 & ~i_10_315_3908_0 & ~i_10_315_4216_0 & ~i_10_315_4285_0))) | (~i_10_315_1916_0 & ~i_10_315_2468_0 & ~i_10_315_2719_0 & ~i_10_315_2980_0 & ~i_10_315_3044_0 & ~i_10_315_3839_0 & ~i_10_315_4271_0))) | (~i_10_315_716_0 & ((~i_10_315_1028_0 & ~i_10_315_1249_0 & ~i_10_315_2027_0 & ((~i_10_315_892_0 & ~i_10_315_2378_0 & ~i_10_315_2566_0 & ~i_10_315_2720_0 & i_10_315_2731_0 & ~i_10_315_3848_0 & ~i_10_315_3908_0) | (~i_10_315_1246_0 & ~i_10_315_1308_0 & ~i_10_315_1313_0 & ~i_10_315_2026_0 & ~i_10_315_3906_0 & ~i_10_315_4566_0 & ~i_10_315_2468_0 & ~i_10_315_2567_0))) | (~i_10_315_3539_0 & ((~i_10_315_1244_0 & ~i_10_315_1310_0 & ~i_10_315_2378_0 & ~i_10_315_2727_0 & ~i_10_315_2731_0 & ~i_10_315_3855_0 & ~i_10_315_3906_0 & ~i_10_315_3908_0) | (~i_10_315_2567_0 & ~i_10_315_2728_0 & ~i_10_315_4288_0 & ~i_10_315_4563_0))))) | (~i_10_315_892_0 & ((~i_10_315_1244_0 & ~i_10_315_2727_0 & ~i_10_315_3389_0 & ~i_10_315_3539_0 & ~i_10_315_3908_0 & i_10_315_4288_0) | (~i_10_315_427_0 & ~i_10_315_1691_0 & ~i_10_315_2378_0 & ~i_10_315_2711_0 & ~i_10_315_3586_0 & ~i_10_315_3848_0 & ~i_10_315_4289_0))) | (~i_10_315_3389_0 & ((~i_10_315_1687_0 & ((i_10_315_463_0 & ~i_10_315_1246_0 & ~i_10_315_2566_0 & ~i_10_315_2980_0 & ~i_10_315_3852_0 & ~i_10_315_4268_0) | (~i_10_315_1691_0 & ~i_10_315_2026_0 & ~i_10_315_2567_0 & ~i_10_315_2608_0 & ~i_10_315_3281_0 & ~i_10_315_4563_0 & ~i_10_315_4566_0))) | (~i_10_315_2729_0 & ~i_10_315_3843_0 & ~i_10_315_3855_0 & i_10_315_4566_0))) | (~i_10_315_2567_0 & ((i_10_315_1825_0 & ~i_10_315_2701_0 & ~i_10_315_2719_0 & ~i_10_315_2722_0 & ~i_10_315_2723_0 & ~i_10_315_3727_0 & ~i_10_315_3906_0) | (~i_10_315_2566_0 & ~i_10_315_2728_0 & ~i_10_315_3787_0 & ~i_10_315_3839_0 & ~i_10_315_4213_0 & ~i_10_315_4268_0))) | (i_10_315_1308_0 & i_10_315_3277_0 & ~i_10_315_3855_0) | (i_10_315_1249_0 & ~i_10_315_2635_0 & ~i_10_315_3042_0 & ~i_10_315_3281_0 & ~i_10_315_3857_0) | (~i_10_315_2608_0 & ~i_10_315_2920_0 & ~i_10_315_3392_0 & ~i_10_315_4284_0 & ~i_10_315_4285_0 & ~i_10_315_4286_0 & ~i_10_315_4566_0));
endmodule



// Benchmark "kernel_10_316" written by ABC on Sun Jul 19 10:26:32 2020

module kernel_10_316 ( 
    i_10_316_81_0, i_10_316_224_0, i_10_316_280_0, i_10_316_284_0,
    i_10_316_286_0, i_10_316_316_0, i_10_316_317_0, i_10_316_328_0,
    i_10_316_390_0, i_10_316_464_0, i_10_316_796_0, i_10_316_799_0,
    i_10_316_800_0, i_10_316_957_0, i_10_316_1000_0, i_10_316_1153_0,
    i_10_316_1236_0, i_10_316_1241_0, i_10_316_1248_0, i_10_316_1263_0,
    i_10_316_1267_0, i_10_316_1307_0, i_10_316_1308_0, i_10_316_1309_0,
    i_10_316_1310_0, i_10_316_1544_0, i_10_316_1575_0, i_10_316_1579_0,
    i_10_316_1655_0, i_10_316_1810_0, i_10_316_1821_0, i_10_316_2017_0,
    i_10_316_2197_0, i_10_316_2312_0, i_10_316_2349_0, i_10_316_2350_0,
    i_10_316_2351_0, i_10_316_2352_0, i_10_316_2353_0, i_10_316_2354_0,
    i_10_316_2355_0, i_10_316_2359_0, i_10_316_2377_0, i_10_316_2378_0,
    i_10_316_2379_0, i_10_316_2380_0, i_10_316_2381_0, i_10_316_2383_0,
    i_10_316_2407_0, i_10_316_2409_0, i_10_316_2448_0, i_10_316_2449_0,
    i_10_316_2452_0, i_10_316_2453_0, i_10_316_2454_0, i_10_316_2471_0,
    i_10_316_2503_0, i_10_316_2506_0, i_10_316_2507_0, i_10_316_2604_0,
    i_10_316_2605_0, i_10_316_2657_0, i_10_316_2659_0, i_10_316_2700_0,
    i_10_316_2701_0, i_10_316_2727_0, i_10_316_2880_0, i_10_316_2882_0,
    i_10_316_2919_0, i_10_316_2965_0, i_10_316_3280_0, i_10_316_3283_0,
    i_10_316_3384_0, i_10_316_3385_0, i_10_316_3403_0, i_10_316_3537_0,
    i_10_316_3586_0, i_10_316_3587_0, i_10_316_3610_0, i_10_316_3613_0,
    i_10_316_3616_0, i_10_316_3836_0, i_10_316_3841_0, i_10_316_3853_0,
    i_10_316_3854_0, i_10_316_3856_0, i_10_316_3890_0, i_10_316_3982_0,
    i_10_316_4113_0, i_10_316_4115_0, i_10_316_4119_0, i_10_316_4127_0,
    i_10_316_4168_0, i_10_316_4271_0, i_10_316_4276_0, i_10_316_4277_0,
    i_10_316_4288_0, i_10_316_4566_0, i_10_316_4567_0, i_10_316_4568_0,
    o_10_316_0_0  );
  input  i_10_316_81_0, i_10_316_224_0, i_10_316_280_0, i_10_316_284_0,
    i_10_316_286_0, i_10_316_316_0, i_10_316_317_0, i_10_316_328_0,
    i_10_316_390_0, i_10_316_464_0, i_10_316_796_0, i_10_316_799_0,
    i_10_316_800_0, i_10_316_957_0, i_10_316_1000_0, i_10_316_1153_0,
    i_10_316_1236_0, i_10_316_1241_0, i_10_316_1248_0, i_10_316_1263_0,
    i_10_316_1267_0, i_10_316_1307_0, i_10_316_1308_0, i_10_316_1309_0,
    i_10_316_1310_0, i_10_316_1544_0, i_10_316_1575_0, i_10_316_1579_0,
    i_10_316_1655_0, i_10_316_1810_0, i_10_316_1821_0, i_10_316_2017_0,
    i_10_316_2197_0, i_10_316_2312_0, i_10_316_2349_0, i_10_316_2350_0,
    i_10_316_2351_0, i_10_316_2352_0, i_10_316_2353_0, i_10_316_2354_0,
    i_10_316_2355_0, i_10_316_2359_0, i_10_316_2377_0, i_10_316_2378_0,
    i_10_316_2379_0, i_10_316_2380_0, i_10_316_2381_0, i_10_316_2383_0,
    i_10_316_2407_0, i_10_316_2409_0, i_10_316_2448_0, i_10_316_2449_0,
    i_10_316_2452_0, i_10_316_2453_0, i_10_316_2454_0, i_10_316_2471_0,
    i_10_316_2503_0, i_10_316_2506_0, i_10_316_2507_0, i_10_316_2604_0,
    i_10_316_2605_0, i_10_316_2657_0, i_10_316_2659_0, i_10_316_2700_0,
    i_10_316_2701_0, i_10_316_2727_0, i_10_316_2880_0, i_10_316_2882_0,
    i_10_316_2919_0, i_10_316_2965_0, i_10_316_3280_0, i_10_316_3283_0,
    i_10_316_3384_0, i_10_316_3385_0, i_10_316_3403_0, i_10_316_3537_0,
    i_10_316_3586_0, i_10_316_3587_0, i_10_316_3610_0, i_10_316_3613_0,
    i_10_316_3616_0, i_10_316_3836_0, i_10_316_3841_0, i_10_316_3853_0,
    i_10_316_3854_0, i_10_316_3856_0, i_10_316_3890_0, i_10_316_3982_0,
    i_10_316_4113_0, i_10_316_4115_0, i_10_316_4119_0, i_10_316_4127_0,
    i_10_316_4168_0, i_10_316_4271_0, i_10_316_4276_0, i_10_316_4277_0,
    i_10_316_4288_0, i_10_316_4566_0, i_10_316_4567_0, i_10_316_4568_0;
  output o_10_316_0_0;
  assign o_10_316_0_0 = ~((~i_10_316_2378_0 & ((~i_10_316_4276_0 & ((~i_10_316_316_0 & ((~i_10_316_1000_0 & ~i_10_316_2312_0 & ~i_10_316_2355_0 & ~i_10_316_2377_0 & ~i_10_316_2381_0 & ~i_10_316_2506_0) | (~i_10_316_390_0 & ~i_10_316_957_0 & ~i_10_316_2352_0 & ~i_10_316_2383_0 & ~i_10_316_3610_0 & ~i_10_316_3890_0 & ~i_10_316_4127_0))) | (~i_10_316_317_0 & ~i_10_316_328_0 & ~i_10_316_1544_0 & ~i_10_316_2353_0 & ~i_10_316_2407_0 & ~i_10_316_4271_0))) | (~i_10_316_1000_0 & ((~i_10_316_1575_0 & ((~i_10_316_1263_0 & ~i_10_316_1309_0 & ~i_10_316_2605_0 & ~i_10_316_4113_0 & i_10_316_4119_0) | (~i_10_316_1655_0 & ~i_10_316_2354_0 & ~i_10_316_2727_0 & ~i_10_316_3890_0 & ~i_10_316_3982_0 & ~i_10_316_4119_0 & ~i_10_316_4271_0))) | (~i_10_316_317_0 & ~i_10_316_796_0 & ~i_10_316_2407_0 & ~i_10_316_2604_0 & ~i_10_316_4119_0) | (i_10_316_796_0 & ~i_10_316_2312_0 & ~i_10_316_2503_0 & ~i_10_316_2727_0 & i_10_316_4271_0))) | (~i_10_316_2379_0 & ((~i_10_316_1810_0 & ~i_10_316_2354_0 & ~i_10_316_2409_0 & ~i_10_316_3613_0 & ~i_10_316_4113_0 & ~i_10_316_4277_0 & ~i_10_316_4288_0) | (~i_10_316_328_0 & i_10_316_1579_0 & ~i_10_316_2507_0 & ~i_10_316_2604_0 & ~i_10_316_2919_0 & ~i_10_316_3537_0 & ~i_10_316_3890_0 & ~i_10_316_4168_0 & ~i_10_316_4566_0))) | (~i_10_316_280_0 & ~i_10_316_1248_0 & ~i_10_316_2377_0 & ~i_10_316_2409_0 & ~i_10_316_2604_0 & ~i_10_316_2657_0 & ~i_10_316_2659_0 & ~i_10_316_3610_0 & ~i_10_316_3890_0 & ~i_10_316_4119_0))) | (~i_10_316_1248_0 & ((~i_10_316_81_0 & ~i_10_316_1000_0 & ~i_10_316_1263_0 & ~i_10_316_1821_0 & ~i_10_316_2017_0 & ~i_10_316_2197_0 & ~i_10_316_2351_0 & ~i_10_316_2503_0 & ~i_10_316_3982_0) | (i_10_316_286_0 & ~i_10_316_2355_0 & ~i_10_316_2409_0 & ~i_10_316_2657_0 & ~i_10_316_4271_0 & ~i_10_316_4277_0))) | (i_10_316_286_0 & ~i_10_316_2351_0 & ((~i_10_316_1263_0 & ~i_10_316_2312_0 & ~i_10_316_2503_0 & ~i_10_316_4271_0 & ~i_10_316_4277_0 & ~i_10_316_2727_0 & ~i_10_316_4119_0) | (~i_10_316_1267_0 & ~i_10_316_2507_0 & ~i_10_316_2701_0 & ~i_10_316_3613_0 & ~i_10_316_4566_0))) | (~i_10_316_4276_0 & ((~i_10_316_1000_0 & ~i_10_316_2507_0 & ~i_10_316_4566_0 & ((~i_10_316_1579_0 & ~i_10_316_2350_0 & ~i_10_316_2355_0) | (~i_10_316_1810_0 & ~i_10_316_2377_0 & ~i_10_316_2407_0 & ~i_10_316_2503_0 & ~i_10_316_2605_0 & ~i_10_316_2659_0))) | (i_10_316_1655_0 & ~i_10_316_2312_0 & ~i_10_316_2359_0 & ~i_10_316_2380_0 & ~i_10_316_2409_0 & i_10_316_2605_0))) | (~i_10_316_1310_0 & ((~i_10_316_2381_0 & i_10_316_3587_0) | (~i_10_316_2409_0 & ~i_10_316_3537_0 & i_10_316_3854_0 & ~i_10_316_3890_0 & ~i_10_316_4277_0 & ~i_10_316_4566_0))) | (~i_10_316_4277_0 & ((~i_10_316_1810_0 & ((~i_10_316_286_0 & ~i_10_316_1263_0 & ~i_10_316_1308_0 & ~i_10_316_2017_0 & ~i_10_316_2700_0 & ~i_10_316_4271_0) | (~i_10_316_1307_0 & ~i_10_316_2349_0 & ~i_10_316_4115_0 & ~i_10_316_4168_0 & ~i_10_316_4567_0))) | (~i_10_316_2700_0 & ~i_10_316_2727_0 & i_10_316_3613_0 & ~i_10_316_3841_0))) | (~i_10_316_2354_0 & ((~i_10_316_2379_0 & i_10_316_2381_0 & ~i_10_316_2407_0 & ~i_10_316_2659_0) | (i_10_316_1000_0 & ~i_10_316_2352_0 & ~i_10_316_2353_0 & ~i_10_316_2355_0 & ~i_10_316_2503_0 & ~i_10_316_2657_0 & ~i_10_316_2882_0 & ~i_10_316_2919_0 & ~i_10_316_3385_0))) | (~i_10_316_2377_0 & ((i_10_316_464_0 & i_10_316_799_0 & ~i_10_316_2700_0) | (~i_10_316_957_0 & ~i_10_316_1579_0 & ~i_10_316_2312_0 & ~i_10_316_2383_0 & ~i_10_316_2409_0 & ~i_10_316_3841_0 & ~i_10_316_3854_0 & ~i_10_316_4115_0 & ~i_10_316_4127_0 & ~i_10_316_4168_0))) | (~i_10_316_2701_0 & ((i_10_316_2919_0 & i_10_316_3384_0) | (i_10_316_2659_0 & i_10_316_3587_0 & ~i_10_316_3982_0))) | (i_10_316_224_0 & ~i_10_316_2355_0 & i_10_316_4119_0) | (i_10_316_2452_0 & ~i_10_316_4127_0) | (i_10_316_957_0 & ~i_10_316_1821_0 & ~i_10_316_2407_0 & ~i_10_316_4119_0 & i_10_316_4568_0));
endmodule



// Benchmark "kernel_10_317" written by ABC on Sun Jul 19 10:26:33 2020

module kernel_10_317 ( 
    i_10_317_88_0, i_10_317_89_0, i_10_317_117_0, i_10_317_149_0,
    i_10_317_178_0, i_10_317_182_0, i_10_317_276_0, i_10_317_277_0,
    i_10_317_282_0, i_10_317_375_0, i_10_317_409_0, i_10_317_410_0,
    i_10_317_436_0, i_10_317_449_0, i_10_317_459_0, i_10_317_460_0,
    i_10_317_461_0, i_10_317_467_0, i_10_317_473_0, i_10_317_515_0,
    i_10_317_578_0, i_10_317_581_0, i_10_317_800_0, i_10_317_906_0,
    i_10_317_1010_0, i_10_317_1040_0, i_10_317_1041_0, i_10_317_1168_0,
    i_10_317_1233_0, i_10_317_1240_0, i_10_317_1241_0, i_10_317_1292_0,
    i_10_317_1310_0, i_10_317_1348_0, i_10_317_1634_0, i_10_317_1650_0,
    i_10_317_1724_0, i_10_317_1767_0, i_10_317_1773_0, i_10_317_1822_0,
    i_10_317_1823_0, i_10_317_1912_0, i_10_317_1950_0, i_10_317_1951_0,
    i_10_317_2038_0, i_10_317_2183_0, i_10_317_2308_0, i_10_317_2337_0,
    i_10_317_2351_0, i_10_317_2352_0, i_10_317_2353_0, i_10_317_2378_0,
    i_10_317_2408_0, i_10_317_2451_0, i_10_317_2470_0, i_10_317_2474_0,
    i_10_317_2509_0, i_10_317_2606_0, i_10_317_2638_0, i_10_317_2711_0,
    i_10_317_2715_0, i_10_317_2741_0, i_10_317_2788_0, i_10_317_2865_0,
    i_10_317_2914_0, i_10_317_2915_0, i_10_317_2924_0, i_10_317_2957_0,
    i_10_317_2983_0, i_10_317_3001_0, i_10_317_3041_0, i_10_317_3046_0,
    i_10_317_3208_0, i_10_317_3209_0, i_10_317_3272_0, i_10_317_3329_0,
    i_10_317_3432_0, i_10_317_3494_0, i_10_317_3500_0, i_10_317_3585_0,
    i_10_317_3588_0, i_10_317_3589_0, i_10_317_3617_0, i_10_317_3733_0,
    i_10_317_3785_0, i_10_317_3806_0, i_10_317_3855_0, i_10_317_3886_0,
    i_10_317_3895_0, i_10_317_3946_0, i_10_317_3967_0, i_10_317_4054_0,
    i_10_317_4182_0, i_10_317_4183_0, i_10_317_4270_0, i_10_317_4273_0,
    i_10_317_4274_0, i_10_317_4463_0, i_10_317_4477_0, i_10_317_4478_0,
    o_10_317_0_0  );
  input  i_10_317_88_0, i_10_317_89_0, i_10_317_117_0, i_10_317_149_0,
    i_10_317_178_0, i_10_317_182_0, i_10_317_276_0, i_10_317_277_0,
    i_10_317_282_0, i_10_317_375_0, i_10_317_409_0, i_10_317_410_0,
    i_10_317_436_0, i_10_317_449_0, i_10_317_459_0, i_10_317_460_0,
    i_10_317_461_0, i_10_317_467_0, i_10_317_473_0, i_10_317_515_0,
    i_10_317_578_0, i_10_317_581_0, i_10_317_800_0, i_10_317_906_0,
    i_10_317_1010_0, i_10_317_1040_0, i_10_317_1041_0, i_10_317_1168_0,
    i_10_317_1233_0, i_10_317_1240_0, i_10_317_1241_0, i_10_317_1292_0,
    i_10_317_1310_0, i_10_317_1348_0, i_10_317_1634_0, i_10_317_1650_0,
    i_10_317_1724_0, i_10_317_1767_0, i_10_317_1773_0, i_10_317_1822_0,
    i_10_317_1823_0, i_10_317_1912_0, i_10_317_1950_0, i_10_317_1951_0,
    i_10_317_2038_0, i_10_317_2183_0, i_10_317_2308_0, i_10_317_2337_0,
    i_10_317_2351_0, i_10_317_2352_0, i_10_317_2353_0, i_10_317_2378_0,
    i_10_317_2408_0, i_10_317_2451_0, i_10_317_2470_0, i_10_317_2474_0,
    i_10_317_2509_0, i_10_317_2606_0, i_10_317_2638_0, i_10_317_2711_0,
    i_10_317_2715_0, i_10_317_2741_0, i_10_317_2788_0, i_10_317_2865_0,
    i_10_317_2914_0, i_10_317_2915_0, i_10_317_2924_0, i_10_317_2957_0,
    i_10_317_2983_0, i_10_317_3001_0, i_10_317_3041_0, i_10_317_3046_0,
    i_10_317_3208_0, i_10_317_3209_0, i_10_317_3272_0, i_10_317_3329_0,
    i_10_317_3432_0, i_10_317_3494_0, i_10_317_3500_0, i_10_317_3585_0,
    i_10_317_3588_0, i_10_317_3589_0, i_10_317_3617_0, i_10_317_3733_0,
    i_10_317_3785_0, i_10_317_3806_0, i_10_317_3855_0, i_10_317_3886_0,
    i_10_317_3895_0, i_10_317_3946_0, i_10_317_3967_0, i_10_317_4054_0,
    i_10_317_4182_0, i_10_317_4183_0, i_10_317_4270_0, i_10_317_4273_0,
    i_10_317_4274_0, i_10_317_4463_0, i_10_317_4477_0, i_10_317_4478_0;
  output o_10_317_0_0;
  assign o_10_317_0_0 = 0;
endmodule



// Benchmark "kernel_10_318" written by ABC on Sun Jul 19 10:26:34 2020

module kernel_10_318 ( 
    i_10_318_28_0, i_10_318_37_0, i_10_318_155_0, i_10_318_193_0,
    i_10_318_273_0, i_10_318_280_0, i_10_318_282_0, i_10_318_332_0,
    i_10_318_424_0, i_10_318_432_0, i_10_318_435_0, i_10_318_436_0,
    i_10_318_437_0, i_10_318_521_0, i_10_318_629_0, i_10_318_752_0,
    i_10_318_779_0, i_10_318_847_0, i_10_318_929_0, i_10_318_1095_0,
    i_10_318_1121_0, i_10_318_1129_0, i_10_318_1239_0, i_10_318_1266_0,
    i_10_318_1268_0, i_10_318_1315_0, i_10_318_1343_0, i_10_318_1355_0,
    i_10_318_1441_0, i_10_318_1548_0, i_10_318_1549_0, i_10_318_1552_0,
    i_10_318_1555_0, i_10_318_1766_0, i_10_318_1797_0, i_10_318_1813_0,
    i_10_318_1814_0, i_10_318_1817_0, i_10_318_1880_0, i_10_318_1992_0,
    i_10_318_2007_0, i_10_318_2206_0, i_10_318_2242_0, i_10_318_2243_0,
    i_10_318_2349_0, i_10_318_2351_0, i_10_318_2353_0, i_10_318_2355_0,
    i_10_318_2356_0, i_10_318_2432_0, i_10_318_2476_0, i_10_318_2541_0,
    i_10_318_2556_0, i_10_318_2565_0, i_10_318_2583_0, i_10_318_2606_0,
    i_10_318_2701_0, i_10_318_2720_0, i_10_318_2727_0, i_10_318_2728_0,
    i_10_318_2756_0, i_10_318_2803_0, i_10_318_2804_0, i_10_318_2844_0,
    i_10_318_2864_0, i_10_318_2883_0, i_10_318_2920_0, i_10_318_2954_0,
    i_10_318_3033_0, i_10_318_3089_0, i_10_318_3238_0, i_10_318_3276_0,
    i_10_318_3277_0, i_10_318_3312_0, i_10_318_3521_0, i_10_318_3523_0,
    i_10_318_3602_0, i_10_318_3700_0, i_10_318_3746_0, i_10_318_3748_0,
    i_10_318_3812_0, i_10_318_3854_0, i_10_318_3855_0, i_10_318_3882_0,
    i_10_318_3989_0, i_10_318_4007_0, i_10_318_4114_0, i_10_318_4115_0,
    i_10_318_4125_0, i_10_318_4147_0, i_10_318_4171_0, i_10_318_4304_0,
    i_10_318_4439_0, i_10_318_4457_0, i_10_318_4522_0, i_10_318_4525_0,
    i_10_318_4532_0, i_10_318_4573_0, i_10_318_4574_0, i_10_318_4591_0,
    o_10_318_0_0  );
  input  i_10_318_28_0, i_10_318_37_0, i_10_318_155_0, i_10_318_193_0,
    i_10_318_273_0, i_10_318_280_0, i_10_318_282_0, i_10_318_332_0,
    i_10_318_424_0, i_10_318_432_0, i_10_318_435_0, i_10_318_436_0,
    i_10_318_437_0, i_10_318_521_0, i_10_318_629_0, i_10_318_752_0,
    i_10_318_779_0, i_10_318_847_0, i_10_318_929_0, i_10_318_1095_0,
    i_10_318_1121_0, i_10_318_1129_0, i_10_318_1239_0, i_10_318_1266_0,
    i_10_318_1268_0, i_10_318_1315_0, i_10_318_1343_0, i_10_318_1355_0,
    i_10_318_1441_0, i_10_318_1548_0, i_10_318_1549_0, i_10_318_1552_0,
    i_10_318_1555_0, i_10_318_1766_0, i_10_318_1797_0, i_10_318_1813_0,
    i_10_318_1814_0, i_10_318_1817_0, i_10_318_1880_0, i_10_318_1992_0,
    i_10_318_2007_0, i_10_318_2206_0, i_10_318_2242_0, i_10_318_2243_0,
    i_10_318_2349_0, i_10_318_2351_0, i_10_318_2353_0, i_10_318_2355_0,
    i_10_318_2356_0, i_10_318_2432_0, i_10_318_2476_0, i_10_318_2541_0,
    i_10_318_2556_0, i_10_318_2565_0, i_10_318_2583_0, i_10_318_2606_0,
    i_10_318_2701_0, i_10_318_2720_0, i_10_318_2727_0, i_10_318_2728_0,
    i_10_318_2756_0, i_10_318_2803_0, i_10_318_2804_0, i_10_318_2844_0,
    i_10_318_2864_0, i_10_318_2883_0, i_10_318_2920_0, i_10_318_2954_0,
    i_10_318_3033_0, i_10_318_3089_0, i_10_318_3238_0, i_10_318_3276_0,
    i_10_318_3277_0, i_10_318_3312_0, i_10_318_3521_0, i_10_318_3523_0,
    i_10_318_3602_0, i_10_318_3700_0, i_10_318_3746_0, i_10_318_3748_0,
    i_10_318_3812_0, i_10_318_3854_0, i_10_318_3855_0, i_10_318_3882_0,
    i_10_318_3989_0, i_10_318_4007_0, i_10_318_4114_0, i_10_318_4115_0,
    i_10_318_4125_0, i_10_318_4147_0, i_10_318_4171_0, i_10_318_4304_0,
    i_10_318_4439_0, i_10_318_4457_0, i_10_318_4522_0, i_10_318_4525_0,
    i_10_318_4532_0, i_10_318_4573_0, i_10_318_4574_0, i_10_318_4591_0;
  output o_10_318_0_0;
  assign o_10_318_0_0 = 0;
endmodule



// Benchmark "kernel_10_319" written by ABC on Sun Jul 19 10:26:35 2020

module kernel_10_319 ( 
    i_10_319_28_0, i_10_319_30_0, i_10_319_147_0, i_10_319_259_0,
    i_10_319_292_0, i_10_319_387_0, i_10_319_390_0, i_10_319_391_0,
    i_10_319_462_0, i_10_319_501_0, i_10_319_633_0, i_10_319_642_0,
    i_10_319_961_0, i_10_319_999_0, i_10_319_1002_0, i_10_319_1056_0,
    i_10_319_1236_0, i_10_319_1237_0, i_10_319_1239_0, i_10_319_1365_0,
    i_10_319_1391_0, i_10_319_1431_0, i_10_319_1434_0, i_10_319_1578_0,
    i_10_319_1579_0, i_10_319_1614_0, i_10_319_1623_0, i_10_319_1650_0,
    i_10_319_1696_0, i_10_319_1731_0, i_10_319_1821_0, i_10_319_1915_0,
    i_10_319_1920_0, i_10_319_1923_0, i_10_319_1938_0, i_10_319_1951_0,
    i_10_319_1992_0, i_10_319_2204_0, i_10_319_2235_0, i_10_319_2267_0,
    i_10_319_2291_0, i_10_319_2325_0, i_10_319_2355_0, i_10_319_2365_0,
    i_10_319_2448_0, i_10_319_2454_0, i_10_319_2466_0, i_10_319_2469_0,
    i_10_319_2470_0, i_10_319_2478_0, i_10_319_2514_0, i_10_319_2565_0,
    i_10_319_2571_0, i_10_319_2590_0, i_10_319_2607_0, i_10_319_2679_0,
    i_10_319_2709_0, i_10_319_2733_0, i_10_319_2742_0, i_10_319_2781_0,
    i_10_319_2784_0, i_10_319_2833_0, i_10_319_2994_0, i_10_319_2995_0,
    i_10_319_3040_0, i_10_319_3042_0, i_10_319_3045_0, i_10_319_3235_0,
    i_10_319_3280_0, i_10_319_3283_0, i_10_319_3318_0, i_10_319_3384_0,
    i_10_319_3387_0, i_10_319_3450_0, i_10_319_3469_0, i_10_319_3471_0,
    i_10_319_3472_0, i_10_319_3500_0, i_10_319_3504_0, i_10_319_3562_0,
    i_10_319_3610_0, i_10_319_3616_0, i_10_319_3625_0, i_10_319_3774_0,
    i_10_319_3807_0, i_10_319_3876_0, i_10_319_3882_0, i_10_319_3942_0,
    i_10_319_3981_0, i_10_319_3982_0, i_10_319_4053_0, i_10_319_4098_0,
    i_10_319_4102_0, i_10_319_4113_0, i_10_319_4189_0, i_10_319_4219_0,
    i_10_319_4226_0, i_10_319_4289_0, i_10_319_4372_0, i_10_319_4585_0,
    o_10_319_0_0  );
  input  i_10_319_28_0, i_10_319_30_0, i_10_319_147_0, i_10_319_259_0,
    i_10_319_292_0, i_10_319_387_0, i_10_319_390_0, i_10_319_391_0,
    i_10_319_462_0, i_10_319_501_0, i_10_319_633_0, i_10_319_642_0,
    i_10_319_961_0, i_10_319_999_0, i_10_319_1002_0, i_10_319_1056_0,
    i_10_319_1236_0, i_10_319_1237_0, i_10_319_1239_0, i_10_319_1365_0,
    i_10_319_1391_0, i_10_319_1431_0, i_10_319_1434_0, i_10_319_1578_0,
    i_10_319_1579_0, i_10_319_1614_0, i_10_319_1623_0, i_10_319_1650_0,
    i_10_319_1696_0, i_10_319_1731_0, i_10_319_1821_0, i_10_319_1915_0,
    i_10_319_1920_0, i_10_319_1923_0, i_10_319_1938_0, i_10_319_1951_0,
    i_10_319_1992_0, i_10_319_2204_0, i_10_319_2235_0, i_10_319_2267_0,
    i_10_319_2291_0, i_10_319_2325_0, i_10_319_2355_0, i_10_319_2365_0,
    i_10_319_2448_0, i_10_319_2454_0, i_10_319_2466_0, i_10_319_2469_0,
    i_10_319_2470_0, i_10_319_2478_0, i_10_319_2514_0, i_10_319_2565_0,
    i_10_319_2571_0, i_10_319_2590_0, i_10_319_2607_0, i_10_319_2679_0,
    i_10_319_2709_0, i_10_319_2733_0, i_10_319_2742_0, i_10_319_2781_0,
    i_10_319_2784_0, i_10_319_2833_0, i_10_319_2994_0, i_10_319_2995_0,
    i_10_319_3040_0, i_10_319_3042_0, i_10_319_3045_0, i_10_319_3235_0,
    i_10_319_3280_0, i_10_319_3283_0, i_10_319_3318_0, i_10_319_3384_0,
    i_10_319_3387_0, i_10_319_3450_0, i_10_319_3469_0, i_10_319_3471_0,
    i_10_319_3472_0, i_10_319_3500_0, i_10_319_3504_0, i_10_319_3562_0,
    i_10_319_3610_0, i_10_319_3616_0, i_10_319_3625_0, i_10_319_3774_0,
    i_10_319_3807_0, i_10_319_3876_0, i_10_319_3882_0, i_10_319_3942_0,
    i_10_319_3981_0, i_10_319_3982_0, i_10_319_4053_0, i_10_319_4098_0,
    i_10_319_4102_0, i_10_319_4113_0, i_10_319_4189_0, i_10_319_4219_0,
    i_10_319_4226_0, i_10_319_4289_0, i_10_319_4372_0, i_10_319_4585_0;
  output o_10_319_0_0;
  assign o_10_319_0_0 = 0;
endmodule



// Benchmark "kernel_10_320" written by ABC on Sun Jul 19 10:26:36 2020

module kernel_10_320 ( 
    i_10_320_223_0, i_10_320_224_0, i_10_320_269_0, i_10_320_281_0,
    i_10_320_316_0, i_10_320_319_0, i_10_320_323_0, i_10_320_328_0,
    i_10_320_410_0, i_10_320_433_0, i_10_320_435_0, i_10_320_444_0,
    i_10_320_445_0, i_10_320_447_0, i_10_320_464_0, i_10_320_465_0,
    i_10_320_518_0, i_10_320_749_0, i_10_320_993_0, i_10_320_1006_0,
    i_10_320_1042_0, i_10_320_1043_0, i_10_320_1081_0, i_10_320_1237_0,
    i_10_320_1238_0, i_10_320_1241_0, i_10_320_1246_0, i_10_320_1296_0,
    i_10_320_1308_0, i_10_320_1309_0, i_10_320_1310_0, i_10_320_1348_0,
    i_10_320_1363_0, i_10_320_1543_0, i_10_320_1579_0, i_10_320_1582_0,
    i_10_320_1628_0, i_10_320_1653_0, i_10_320_1821_0, i_10_320_1824_0,
    i_10_320_1825_0, i_10_320_1911_0, i_10_320_1912_0, i_10_320_1913_0,
    i_10_320_1990_0, i_10_320_2186_0, i_10_320_2358_0, i_10_320_2380_0,
    i_10_320_2383_0, i_10_320_2633_0, i_10_320_2635_0, i_10_320_2657_0,
    i_10_320_2659_0, i_10_320_2660_0, i_10_320_2707_0, i_10_320_2708_0,
    i_10_320_2710_0, i_10_320_2718_0, i_10_320_2732_0, i_10_320_2789_0,
    i_10_320_2817_0, i_10_320_2818_0, i_10_320_2819_0, i_10_320_2828_0,
    i_10_320_2882_0, i_10_320_2920_0, i_10_320_2921_0, i_10_320_2924_0,
    i_10_320_3033_0, i_10_320_3076_0, i_10_320_3155_0, i_10_320_3199_0,
    i_10_320_3276_0, i_10_320_3338_0, i_10_320_3386_0, i_10_320_3389_0,
    i_10_320_3407_0, i_10_320_3523_0, i_10_320_3544_0, i_10_320_3584_0,
    i_10_320_3612_0, i_10_320_3613_0, i_10_320_3614_0, i_10_320_3649_0,
    i_10_320_3785_0, i_10_320_3834_0, i_10_320_3847_0, i_10_320_3848_0,
    i_10_320_3850_0, i_10_320_3857_0, i_10_320_3907_0, i_10_320_3986_0,
    i_10_320_4116_0, i_10_320_4117_0, i_10_320_4118_0, i_10_320_4119_0,
    i_10_320_4120_0, i_10_320_4125_0, i_10_320_4564_0, i_10_320_4565_0,
    o_10_320_0_0  );
  input  i_10_320_223_0, i_10_320_224_0, i_10_320_269_0, i_10_320_281_0,
    i_10_320_316_0, i_10_320_319_0, i_10_320_323_0, i_10_320_328_0,
    i_10_320_410_0, i_10_320_433_0, i_10_320_435_0, i_10_320_444_0,
    i_10_320_445_0, i_10_320_447_0, i_10_320_464_0, i_10_320_465_0,
    i_10_320_518_0, i_10_320_749_0, i_10_320_993_0, i_10_320_1006_0,
    i_10_320_1042_0, i_10_320_1043_0, i_10_320_1081_0, i_10_320_1237_0,
    i_10_320_1238_0, i_10_320_1241_0, i_10_320_1246_0, i_10_320_1296_0,
    i_10_320_1308_0, i_10_320_1309_0, i_10_320_1310_0, i_10_320_1348_0,
    i_10_320_1363_0, i_10_320_1543_0, i_10_320_1579_0, i_10_320_1582_0,
    i_10_320_1628_0, i_10_320_1653_0, i_10_320_1821_0, i_10_320_1824_0,
    i_10_320_1825_0, i_10_320_1911_0, i_10_320_1912_0, i_10_320_1913_0,
    i_10_320_1990_0, i_10_320_2186_0, i_10_320_2358_0, i_10_320_2380_0,
    i_10_320_2383_0, i_10_320_2633_0, i_10_320_2635_0, i_10_320_2657_0,
    i_10_320_2659_0, i_10_320_2660_0, i_10_320_2707_0, i_10_320_2708_0,
    i_10_320_2710_0, i_10_320_2718_0, i_10_320_2732_0, i_10_320_2789_0,
    i_10_320_2817_0, i_10_320_2818_0, i_10_320_2819_0, i_10_320_2828_0,
    i_10_320_2882_0, i_10_320_2920_0, i_10_320_2921_0, i_10_320_2924_0,
    i_10_320_3033_0, i_10_320_3076_0, i_10_320_3155_0, i_10_320_3199_0,
    i_10_320_3276_0, i_10_320_3338_0, i_10_320_3386_0, i_10_320_3389_0,
    i_10_320_3407_0, i_10_320_3523_0, i_10_320_3544_0, i_10_320_3584_0,
    i_10_320_3612_0, i_10_320_3613_0, i_10_320_3614_0, i_10_320_3649_0,
    i_10_320_3785_0, i_10_320_3834_0, i_10_320_3847_0, i_10_320_3848_0,
    i_10_320_3850_0, i_10_320_3857_0, i_10_320_3907_0, i_10_320_3986_0,
    i_10_320_4116_0, i_10_320_4117_0, i_10_320_4118_0, i_10_320_4119_0,
    i_10_320_4120_0, i_10_320_4125_0, i_10_320_4564_0, i_10_320_4565_0;
  output o_10_320_0_0;
  assign o_10_320_0_0 = ~((~i_10_320_1913_0 & ((~i_10_320_269_0 & ((~i_10_320_1238_0 & ((~i_10_320_281_0 & ((~i_10_320_319_0 & ~i_10_320_1363_0 & ~i_10_320_1653_0 & ~i_10_320_1821_0 & ~i_10_320_1911_0 & ~i_10_320_2633_0) | (~i_10_320_328_0 & ~i_10_320_444_0 & ~i_10_320_1912_0 & ~i_10_320_2383_0 & ~i_10_320_2659_0 & ~i_10_320_2732_0 & ~i_10_320_3276_0))) | (~i_10_320_1081_0 & ~i_10_320_1912_0 & i_10_320_3649_0 & ~i_10_320_3907_0 & i_10_320_4117_0))) | (~i_10_320_749_0 & ~i_10_320_1912_0 & ~i_10_320_2789_0 & ~i_10_320_2818_0 & ~i_10_320_3033_0 & i_10_320_4117_0))) | (~i_10_320_1042_0 & ((~i_10_320_410_0 & ~i_10_320_433_0 & ~i_10_320_444_0 & ~i_10_320_1081_0 & ~i_10_320_1309_0 & ~i_10_320_2921_0 & ~i_10_320_3386_0 & ~i_10_320_3407_0 & ~i_10_320_3857_0 & ~i_10_320_3986_0) | (~i_10_320_1990_0 & i_10_320_2358_0 & ~i_10_320_2707_0 & ~i_10_320_2708_0 & ~i_10_320_2789_0 & ~i_10_320_4564_0))) | (~i_10_320_1821_0 & ~i_10_320_3584_0 & ((~i_10_320_464_0 & ~i_10_320_749_0 & ~i_10_320_1238_0 & ~i_10_320_1241_0 & ~i_10_320_1911_0 & ~i_10_320_1912_0 & ~i_10_320_2635_0 & ~i_10_320_3612_0) | (~i_10_320_1237_0 & ~i_10_320_1309_0 & ~i_10_320_3523_0 & ~i_10_320_3544_0 & ~i_10_320_3785_0))) | (i_10_320_445_0 & ~i_10_320_1006_0 & i_10_320_1825_0 & ~i_10_320_2817_0 & ~i_10_320_3649_0) | (~i_10_320_1310_0 & ~i_10_320_1348_0 & ~i_10_320_1911_0 & i_10_320_4119_0))) | (~i_10_320_1043_0 & ((~i_10_320_269_0 & ((~i_10_320_1238_0 & i_10_320_1309_0 & ~i_10_320_1911_0 & ~i_10_320_2718_0 & ~i_10_320_2789_0 & ~i_10_320_2819_0 & ~i_10_320_3033_0 & ~i_10_320_3544_0 & ~i_10_320_3857_0) | (~i_10_320_1308_0 & ~i_10_320_1310_0 & ~i_10_320_1348_0 & ~i_10_320_1363_0 & ~i_10_320_1628_0 & ~i_10_320_2657_0 & ~i_10_320_2659_0 & ~i_10_320_2817_0 & ~i_10_320_3986_0))) | (~i_10_320_1310_0 & ~i_10_320_1348_0 & ~i_10_320_433_0 & i_10_320_444_0 & ~i_10_320_1911_0 & ~i_10_320_1912_0 & ~i_10_320_3612_0 & ~i_10_320_3986_0) | (~i_10_320_281_0 & ~i_10_320_328_0 & ~i_10_320_1238_0 & ~i_10_320_2789_0 & i_10_320_2882_0 & i_10_320_3614_0))) | (~i_10_320_1237_0 & ((~i_10_320_1912_0 & i_10_320_2921_0 & ~i_10_320_3613_0) | (~i_10_320_1238_0 & ~i_10_320_1348_0 & ~i_10_320_2383_0 & i_10_320_2635_0 & ~i_10_320_2660_0 & ~i_10_320_2708_0 & ~i_10_320_2710_0 & ~i_10_320_2732_0 & ~i_10_320_3544_0 & ~i_10_320_3847_0))) | (~i_10_320_1309_0 & ((~i_10_320_410_0 & ~i_10_320_518_0 & ~i_10_320_1310_0 & ~i_10_320_1653_0 & i_10_320_1825_0 & ~i_10_320_2789_0 & ~i_10_320_2817_0 & ~i_10_320_3076_0 & ~i_10_320_3986_0) | (~i_10_320_2818_0 & i_10_320_2924_0 & i_10_320_4120_0))) | (~i_10_320_2708_0 & ((~i_10_320_410_0 & ((~i_10_320_323_0 & ~i_10_320_328_0 & ~i_10_320_1081_0 & ~i_10_320_1348_0 & ~i_10_320_1653_0 & ~i_10_320_2186_0 & ~i_10_320_2659_0 & ~i_10_320_2660_0 & ~i_10_320_2819_0 & ~i_10_320_3544_0 & ~i_10_320_3785_0 & ~i_10_320_3907_0 & ~i_10_320_4116_0) | (i_10_320_2920_0 & i_10_320_2924_0 & ~i_10_320_4120_0))) | (~i_10_320_433_0 & ~i_10_320_518_0 & ~i_10_320_1911_0 & ~i_10_320_2657_0 & ~i_10_320_2789_0 & ~i_10_320_2819_0 & ~i_10_320_2924_0 & ~i_10_320_3076_0 & ~i_10_320_3386_0 & ~i_10_320_3614_0 & ~i_10_320_3785_0) | (i_10_320_2718_0 & ~i_10_320_2818_0 & i_10_320_4119_0 & i_10_320_4120_0))) | (~i_10_320_518_0 & ((~i_10_320_1042_0 & ~i_10_320_1310_0 & i_10_320_1824_0 & ~i_10_320_2358_0 & ~i_10_320_2659_0 & ~i_10_320_2660_0 & ~i_10_320_3857_0) | (~i_10_320_464_0 & ~i_10_320_1308_0 & i_10_320_1653_0 & ~i_10_320_3649_0 & ~i_10_320_4119_0))) | (~i_10_320_2660_0 & ((~i_10_320_1310_0 & ~i_10_320_1821_0 & ((~i_10_320_224_0 & i_10_320_323_0 & ~i_10_320_1363_0 & ~i_10_320_1912_0 & i_10_320_3386_0) | (~i_10_320_2657_0 & ~i_10_320_2718_0 & ~i_10_320_3076_0 & ~i_10_320_3199_0 & ~i_10_320_3613_0 & ~i_10_320_3614_0 & i_10_320_3649_0))) | (~i_10_320_2718_0 & ~i_10_320_2732_0 & ~i_10_320_2882_0 & ~i_10_320_3389_0 & ~i_10_320_3584_0 & ~i_10_320_3649_0 & i_10_320_3857_0 & ~i_10_320_3986_0))) | (~i_10_320_3523_0 & ((i_10_320_2710_0 & i_10_320_2732_0 & i_10_320_3389_0) | (i_10_320_2707_0 & ~i_10_320_3986_0 & i_10_320_4119_0))));
endmodule



// Benchmark "kernel_10_321" written by ABC on Sun Jul 19 10:26:37 2020

module kernel_10_321 ( 
    i_10_321_117_0, i_10_321_175_0, i_10_321_180_0, i_10_321_268_0,
    i_10_321_279_0, i_10_321_319_0, i_10_321_407_0, i_10_321_408_0,
    i_10_321_427_0, i_10_321_428_0, i_10_321_440_0, i_10_321_444_0,
    i_10_321_445_0, i_10_321_461_0, i_10_321_462_0, i_10_321_712_0,
    i_10_321_748_0, i_10_321_796_0, i_10_321_897_0, i_10_321_958_0,
    i_10_321_1005_0, i_10_321_1166_0, i_10_321_1233_0, i_10_321_1238_0,
    i_10_321_1242_0, i_10_321_1366_0, i_10_321_1367_0, i_10_321_1385_0,
    i_10_321_1444_0, i_10_321_1612_0, i_10_321_1654_0, i_10_321_1655_0,
    i_10_321_1683_0, i_10_321_1821_0, i_10_321_1822_0, i_10_321_1823_0,
    i_10_321_1824_0, i_10_321_1911_0, i_10_321_1946_0, i_10_321_2001_0,
    i_10_321_2004_0, i_10_321_2020_0, i_10_321_2199_0, i_10_321_2311_0,
    i_10_321_2355_0, i_10_321_2451_0, i_10_321_2452_0, i_10_321_2460_0,
    i_10_321_2629_0, i_10_321_2631_0, i_10_321_2633_0, i_10_321_2643_0,
    i_10_321_2662_0, i_10_321_2721_0, i_10_321_2730_0, i_10_321_2733_0,
    i_10_321_2830_0, i_10_321_2882_0, i_10_321_2885_0, i_10_321_2916_0,
    i_10_321_2917_0, i_10_321_2985_0, i_10_321_2986_0, i_10_321_3035_0,
    i_10_321_3036_0, i_10_321_3040_0, i_10_321_3087_0, i_10_321_3094_0,
    i_10_321_3195_0, i_10_321_3196_0, i_10_321_3280_0, i_10_321_3284_0,
    i_10_321_3403_0, i_10_321_3469_0, i_10_321_3497_0, i_10_321_3541_0,
    i_10_321_3590_0, i_10_321_3609_0, i_10_321_3614_0, i_10_321_3682_0,
    i_10_321_3683_0, i_10_321_3721_0, i_10_321_3843_0, i_10_321_3847_0,
    i_10_321_3855_0, i_10_321_3858_0, i_10_321_3859_0, i_10_321_3918_0,
    i_10_321_3980_0, i_10_321_3983_0, i_10_321_4113_0, i_10_321_4119_0,
    i_10_321_4120_0, i_10_321_4122_0, i_10_321_4183_0, i_10_321_4189_0,
    i_10_321_4275_0, i_10_321_4288_0, i_10_321_4517_0, i_10_321_4566_0,
    o_10_321_0_0  );
  input  i_10_321_117_0, i_10_321_175_0, i_10_321_180_0, i_10_321_268_0,
    i_10_321_279_0, i_10_321_319_0, i_10_321_407_0, i_10_321_408_0,
    i_10_321_427_0, i_10_321_428_0, i_10_321_440_0, i_10_321_444_0,
    i_10_321_445_0, i_10_321_461_0, i_10_321_462_0, i_10_321_712_0,
    i_10_321_748_0, i_10_321_796_0, i_10_321_897_0, i_10_321_958_0,
    i_10_321_1005_0, i_10_321_1166_0, i_10_321_1233_0, i_10_321_1238_0,
    i_10_321_1242_0, i_10_321_1366_0, i_10_321_1367_0, i_10_321_1385_0,
    i_10_321_1444_0, i_10_321_1612_0, i_10_321_1654_0, i_10_321_1655_0,
    i_10_321_1683_0, i_10_321_1821_0, i_10_321_1822_0, i_10_321_1823_0,
    i_10_321_1824_0, i_10_321_1911_0, i_10_321_1946_0, i_10_321_2001_0,
    i_10_321_2004_0, i_10_321_2020_0, i_10_321_2199_0, i_10_321_2311_0,
    i_10_321_2355_0, i_10_321_2451_0, i_10_321_2452_0, i_10_321_2460_0,
    i_10_321_2629_0, i_10_321_2631_0, i_10_321_2633_0, i_10_321_2643_0,
    i_10_321_2662_0, i_10_321_2721_0, i_10_321_2730_0, i_10_321_2733_0,
    i_10_321_2830_0, i_10_321_2882_0, i_10_321_2885_0, i_10_321_2916_0,
    i_10_321_2917_0, i_10_321_2985_0, i_10_321_2986_0, i_10_321_3035_0,
    i_10_321_3036_0, i_10_321_3040_0, i_10_321_3087_0, i_10_321_3094_0,
    i_10_321_3195_0, i_10_321_3196_0, i_10_321_3280_0, i_10_321_3284_0,
    i_10_321_3403_0, i_10_321_3469_0, i_10_321_3497_0, i_10_321_3541_0,
    i_10_321_3590_0, i_10_321_3609_0, i_10_321_3614_0, i_10_321_3682_0,
    i_10_321_3683_0, i_10_321_3721_0, i_10_321_3843_0, i_10_321_3847_0,
    i_10_321_3855_0, i_10_321_3858_0, i_10_321_3859_0, i_10_321_3918_0,
    i_10_321_3980_0, i_10_321_3983_0, i_10_321_4113_0, i_10_321_4119_0,
    i_10_321_4120_0, i_10_321_4122_0, i_10_321_4183_0, i_10_321_4189_0,
    i_10_321_4275_0, i_10_321_4288_0, i_10_321_4517_0, i_10_321_4566_0;
  output o_10_321_0_0;
  assign o_10_321_0_0 = 0;
endmodule



// Benchmark "kernel_10_322" written by ABC on Sun Jul 19 10:26:38 2020

module kernel_10_322 ( 
    i_10_322_40_0, i_10_322_41_0, i_10_322_43_0, i_10_322_120_0,
    i_10_322_124_0, i_10_322_172_0, i_10_322_179_0, i_10_322_224_0,
    i_10_322_293_0, i_10_322_315_0, i_10_322_324_0, i_10_322_325_0,
    i_10_322_328_0, i_10_322_390_0, i_10_322_391_0, i_10_322_407_0,
    i_10_322_410_0, i_10_322_413_0, i_10_322_446_0, i_10_322_539_0,
    i_10_322_561_0, i_10_322_796_0, i_10_322_800_0, i_10_322_826_0,
    i_10_322_905_0, i_10_322_961_0, i_10_322_998_0, i_10_322_1006_0,
    i_10_322_1087_0, i_10_322_1157_0, i_10_322_1160_0, i_10_322_1239_0,
    i_10_322_1241_0, i_10_322_1307_0, i_10_322_1309_0, i_10_322_1310_0,
    i_10_322_1349_0, i_10_322_1364_0, i_10_322_1432_0, i_10_322_1448_0,
    i_10_322_1451_0, i_10_322_1649_0, i_10_322_1715_0, i_10_322_1874_0,
    i_10_322_1903_0, i_10_322_1921_0, i_10_322_1947_0, i_10_322_2267_0,
    i_10_322_2363_0, i_10_322_2365_0, i_10_322_2366_0, i_10_322_2411_0,
    i_10_322_2471_0, i_10_322_2510_0, i_10_322_2557_0, i_10_322_2561_0,
    i_10_322_2606_0, i_10_322_2609_0, i_10_322_2611_0, i_10_322_2616_0,
    i_10_322_2617_0, i_10_322_2629_0, i_10_322_2632_0, i_10_322_2702_0,
    i_10_322_2704_0, i_10_322_2705_0, i_10_322_2710_0, i_10_322_2735_0,
    i_10_322_2786_0, i_10_322_2823_0, i_10_322_2882_0, i_10_322_2920_0,
    i_10_322_2957_0, i_10_322_3047_0, i_10_322_3049_0, i_10_322_3090_0,
    i_10_322_3093_0, i_10_322_3236_0, i_10_322_3239_0, i_10_322_3292_0,
    i_10_322_3401_0, i_10_322_3473_0, i_10_322_3527_0, i_10_322_3563_0,
    i_10_322_3781_0, i_10_322_3793_0, i_10_322_3811_0, i_10_322_3812_0,
    i_10_322_3835_0, i_10_322_3836_0, i_10_322_4052_0, i_10_322_4055_0,
    i_10_322_4121_0, i_10_322_4130_0, i_10_322_4171_0, i_10_322_4175_0,
    i_10_322_4281_0, i_10_322_4372_0, i_10_322_4571_0, i_10_322_4586_0,
    o_10_322_0_0  );
  input  i_10_322_40_0, i_10_322_41_0, i_10_322_43_0, i_10_322_120_0,
    i_10_322_124_0, i_10_322_172_0, i_10_322_179_0, i_10_322_224_0,
    i_10_322_293_0, i_10_322_315_0, i_10_322_324_0, i_10_322_325_0,
    i_10_322_328_0, i_10_322_390_0, i_10_322_391_0, i_10_322_407_0,
    i_10_322_410_0, i_10_322_413_0, i_10_322_446_0, i_10_322_539_0,
    i_10_322_561_0, i_10_322_796_0, i_10_322_800_0, i_10_322_826_0,
    i_10_322_905_0, i_10_322_961_0, i_10_322_998_0, i_10_322_1006_0,
    i_10_322_1087_0, i_10_322_1157_0, i_10_322_1160_0, i_10_322_1239_0,
    i_10_322_1241_0, i_10_322_1307_0, i_10_322_1309_0, i_10_322_1310_0,
    i_10_322_1349_0, i_10_322_1364_0, i_10_322_1432_0, i_10_322_1448_0,
    i_10_322_1451_0, i_10_322_1649_0, i_10_322_1715_0, i_10_322_1874_0,
    i_10_322_1903_0, i_10_322_1921_0, i_10_322_1947_0, i_10_322_2267_0,
    i_10_322_2363_0, i_10_322_2365_0, i_10_322_2366_0, i_10_322_2411_0,
    i_10_322_2471_0, i_10_322_2510_0, i_10_322_2557_0, i_10_322_2561_0,
    i_10_322_2606_0, i_10_322_2609_0, i_10_322_2611_0, i_10_322_2616_0,
    i_10_322_2617_0, i_10_322_2629_0, i_10_322_2632_0, i_10_322_2702_0,
    i_10_322_2704_0, i_10_322_2705_0, i_10_322_2710_0, i_10_322_2735_0,
    i_10_322_2786_0, i_10_322_2823_0, i_10_322_2882_0, i_10_322_2920_0,
    i_10_322_2957_0, i_10_322_3047_0, i_10_322_3049_0, i_10_322_3090_0,
    i_10_322_3093_0, i_10_322_3236_0, i_10_322_3239_0, i_10_322_3292_0,
    i_10_322_3401_0, i_10_322_3473_0, i_10_322_3527_0, i_10_322_3563_0,
    i_10_322_3781_0, i_10_322_3793_0, i_10_322_3811_0, i_10_322_3812_0,
    i_10_322_3835_0, i_10_322_3836_0, i_10_322_4052_0, i_10_322_4055_0,
    i_10_322_4121_0, i_10_322_4130_0, i_10_322_4171_0, i_10_322_4175_0,
    i_10_322_4281_0, i_10_322_4372_0, i_10_322_4571_0, i_10_322_4586_0;
  output o_10_322_0_0;
  assign o_10_322_0_0 = 0;
endmodule



// Benchmark "kernel_10_323" written by ABC on Sun Jul 19 10:26:39 2020

module kernel_10_323 ( 
    i_10_323_175_0, i_10_323_178_0, i_10_323_287_0, i_10_323_315_0,
    i_10_323_405_0, i_10_323_496_0, i_10_323_506_0, i_10_323_638_0,
    i_10_323_766_0, i_10_323_796_0, i_10_323_797_0, i_10_323_821_0,
    i_10_323_874_0, i_10_323_899_0, i_10_323_1000_0, i_10_323_1001_0,
    i_10_323_1103_0, i_10_323_1112_0, i_10_323_1207_0, i_10_323_1211_0,
    i_10_323_1235_0, i_10_323_1240_0, i_10_323_1274_0, i_10_323_1283_0,
    i_10_323_1301_0, i_10_323_1306_0, i_10_323_1363_0, i_10_323_1400_0,
    i_10_323_1541_0, i_10_323_1562_0, i_10_323_1565_0, i_10_323_1634_0,
    i_10_323_1688_0, i_10_323_1724_0, i_10_323_1729_0, i_10_323_1733_0,
    i_10_323_1799_0, i_10_323_1802_0, i_10_323_1804_0, i_10_323_1805_0,
    i_10_323_1916_0, i_10_323_1981_0, i_10_323_1984_0, i_10_323_2006_0,
    i_10_323_2186_0, i_10_323_2198_0, i_10_323_2201_0, i_10_323_2237_0,
    i_10_323_2249_0, i_10_323_2258_0, i_10_323_2566_0, i_10_323_2714_0,
    i_10_323_2717_0, i_10_323_2722_0, i_10_323_2728_0, i_10_323_2729_0,
    i_10_323_2747_0, i_10_323_2848_0, i_10_323_2890_0, i_10_323_2915_0,
    i_10_323_2965_0, i_10_323_2966_0, i_10_323_2975_0, i_10_323_3025_0,
    i_10_323_3053_0, i_10_323_3233_0, i_10_323_3281_0, i_10_323_3293_0,
    i_10_323_3296_0, i_10_323_3384_0, i_10_323_3433_0, i_10_323_3436_0,
    i_10_323_3470_0, i_10_323_3503_0, i_10_323_3539_0, i_10_323_3542_0,
    i_10_323_3566_0, i_10_323_3569_0, i_10_323_3586_0, i_10_323_3587_0,
    i_10_323_3620_0, i_10_323_3646_0, i_10_323_3682_0, i_10_323_3715_0,
    i_10_323_3787_0, i_10_323_3793_0, i_10_323_3796_0, i_10_323_3803_0,
    i_10_323_3839_0, i_10_323_3844_0, i_10_323_4007_0, i_10_323_4028_0,
    i_10_323_4150_0, i_10_323_4168_0, i_10_323_4169_0, i_10_323_4277_0,
    i_10_323_4547_0, i_10_323_4570_0, i_10_323_4571_0, i_10_323_4586_0,
    o_10_323_0_0  );
  input  i_10_323_175_0, i_10_323_178_0, i_10_323_287_0, i_10_323_315_0,
    i_10_323_405_0, i_10_323_496_0, i_10_323_506_0, i_10_323_638_0,
    i_10_323_766_0, i_10_323_796_0, i_10_323_797_0, i_10_323_821_0,
    i_10_323_874_0, i_10_323_899_0, i_10_323_1000_0, i_10_323_1001_0,
    i_10_323_1103_0, i_10_323_1112_0, i_10_323_1207_0, i_10_323_1211_0,
    i_10_323_1235_0, i_10_323_1240_0, i_10_323_1274_0, i_10_323_1283_0,
    i_10_323_1301_0, i_10_323_1306_0, i_10_323_1363_0, i_10_323_1400_0,
    i_10_323_1541_0, i_10_323_1562_0, i_10_323_1565_0, i_10_323_1634_0,
    i_10_323_1688_0, i_10_323_1724_0, i_10_323_1729_0, i_10_323_1733_0,
    i_10_323_1799_0, i_10_323_1802_0, i_10_323_1804_0, i_10_323_1805_0,
    i_10_323_1916_0, i_10_323_1981_0, i_10_323_1984_0, i_10_323_2006_0,
    i_10_323_2186_0, i_10_323_2198_0, i_10_323_2201_0, i_10_323_2237_0,
    i_10_323_2249_0, i_10_323_2258_0, i_10_323_2566_0, i_10_323_2714_0,
    i_10_323_2717_0, i_10_323_2722_0, i_10_323_2728_0, i_10_323_2729_0,
    i_10_323_2747_0, i_10_323_2848_0, i_10_323_2890_0, i_10_323_2915_0,
    i_10_323_2965_0, i_10_323_2966_0, i_10_323_2975_0, i_10_323_3025_0,
    i_10_323_3053_0, i_10_323_3233_0, i_10_323_3281_0, i_10_323_3293_0,
    i_10_323_3296_0, i_10_323_3384_0, i_10_323_3433_0, i_10_323_3436_0,
    i_10_323_3470_0, i_10_323_3503_0, i_10_323_3539_0, i_10_323_3542_0,
    i_10_323_3566_0, i_10_323_3569_0, i_10_323_3586_0, i_10_323_3587_0,
    i_10_323_3620_0, i_10_323_3646_0, i_10_323_3682_0, i_10_323_3715_0,
    i_10_323_3787_0, i_10_323_3793_0, i_10_323_3796_0, i_10_323_3803_0,
    i_10_323_3839_0, i_10_323_3844_0, i_10_323_4007_0, i_10_323_4028_0,
    i_10_323_4150_0, i_10_323_4168_0, i_10_323_4169_0, i_10_323_4277_0,
    i_10_323_4547_0, i_10_323_4570_0, i_10_323_4571_0, i_10_323_4586_0;
  output o_10_323_0_0;
  assign o_10_323_0_0 = 0;
endmodule



// Benchmark "kernel_10_324" written by ABC on Sun Jul 19 10:26:40 2020

module kernel_10_324 ( 
    i_10_324_220_0, i_10_324_223_0, i_10_324_247_0, i_10_324_248_0,
    i_10_324_446_0, i_10_324_462_0, i_10_324_520_0, i_10_324_733_0,
    i_10_324_736_0, i_10_324_797_0, i_10_324_927_0, i_10_324_928_0,
    i_10_324_929_0, i_10_324_971_0, i_10_324_1028_0, i_10_324_1040_0,
    i_10_324_1083_0, i_10_324_1117_0, i_10_324_1233_0, i_10_324_1236_0,
    i_10_324_1237_0, i_10_324_1239_0, i_10_324_1243_0, i_10_324_1305_0,
    i_10_324_1306_0, i_10_324_1342_0, i_10_324_1446_0, i_10_324_1546_0,
    i_10_324_1547_0, i_10_324_1549_0, i_10_324_1551_0, i_10_324_1552_0,
    i_10_324_1648_0, i_10_324_1649_0, i_10_324_1683_0, i_10_324_1684_0,
    i_10_324_1685_0, i_10_324_1688_0, i_10_324_1691_0, i_10_324_1818_0,
    i_10_324_1819_0, i_10_324_1823_0, i_10_324_1826_0, i_10_324_1910_0,
    i_10_324_1915_0, i_10_324_1916_0, i_10_324_1991_0, i_10_324_2006_0,
    i_10_324_2309_0, i_10_324_2353_0, i_10_324_2357_0, i_10_324_2362_0,
    i_10_324_2379_0, i_10_324_2380_0, i_10_324_2430_0, i_10_324_2450_0,
    i_10_324_2451_0, i_10_324_2452_0, i_10_324_2569_0, i_10_324_2573_0,
    i_10_324_2725_0, i_10_324_2727_0, i_10_324_2832_0, i_10_324_2923_0,
    i_10_324_3072_0, i_10_324_3073_0, i_10_324_3087_0, i_10_324_3195_0,
    i_10_324_3196_0, i_10_324_3278_0, i_10_324_3385_0, i_10_324_3388_0,
    i_10_324_3391_0, i_10_324_3407_0, i_10_324_3433_0, i_10_324_3538_0,
    i_10_324_3550_0, i_10_324_3551_0, i_10_324_3586_0, i_10_324_3612_0,
    i_10_324_3648_0, i_10_324_3649_0, i_10_324_3650_0, i_10_324_3787_0,
    i_10_324_3838_0, i_10_324_3839_0, i_10_324_3847_0, i_10_324_3848_0,
    i_10_324_3855_0, i_10_324_3856_0, i_10_324_4009_0, i_10_324_4027_0,
    i_10_324_4057_0, i_10_324_4153_0, i_10_324_4175_0, i_10_324_4286_0,
    i_10_324_4375_0, i_10_324_4376_0, i_10_324_4564_0, i_10_324_4568_0,
    o_10_324_0_0  );
  input  i_10_324_220_0, i_10_324_223_0, i_10_324_247_0, i_10_324_248_0,
    i_10_324_446_0, i_10_324_462_0, i_10_324_520_0, i_10_324_733_0,
    i_10_324_736_0, i_10_324_797_0, i_10_324_927_0, i_10_324_928_0,
    i_10_324_929_0, i_10_324_971_0, i_10_324_1028_0, i_10_324_1040_0,
    i_10_324_1083_0, i_10_324_1117_0, i_10_324_1233_0, i_10_324_1236_0,
    i_10_324_1237_0, i_10_324_1239_0, i_10_324_1243_0, i_10_324_1305_0,
    i_10_324_1306_0, i_10_324_1342_0, i_10_324_1446_0, i_10_324_1546_0,
    i_10_324_1547_0, i_10_324_1549_0, i_10_324_1551_0, i_10_324_1552_0,
    i_10_324_1648_0, i_10_324_1649_0, i_10_324_1683_0, i_10_324_1684_0,
    i_10_324_1685_0, i_10_324_1688_0, i_10_324_1691_0, i_10_324_1818_0,
    i_10_324_1819_0, i_10_324_1823_0, i_10_324_1826_0, i_10_324_1910_0,
    i_10_324_1915_0, i_10_324_1916_0, i_10_324_1991_0, i_10_324_2006_0,
    i_10_324_2309_0, i_10_324_2353_0, i_10_324_2357_0, i_10_324_2362_0,
    i_10_324_2379_0, i_10_324_2380_0, i_10_324_2430_0, i_10_324_2450_0,
    i_10_324_2451_0, i_10_324_2452_0, i_10_324_2569_0, i_10_324_2573_0,
    i_10_324_2725_0, i_10_324_2727_0, i_10_324_2832_0, i_10_324_2923_0,
    i_10_324_3072_0, i_10_324_3073_0, i_10_324_3087_0, i_10_324_3195_0,
    i_10_324_3196_0, i_10_324_3278_0, i_10_324_3385_0, i_10_324_3388_0,
    i_10_324_3391_0, i_10_324_3407_0, i_10_324_3433_0, i_10_324_3538_0,
    i_10_324_3550_0, i_10_324_3551_0, i_10_324_3586_0, i_10_324_3612_0,
    i_10_324_3648_0, i_10_324_3649_0, i_10_324_3650_0, i_10_324_3787_0,
    i_10_324_3838_0, i_10_324_3839_0, i_10_324_3847_0, i_10_324_3848_0,
    i_10_324_3855_0, i_10_324_3856_0, i_10_324_4009_0, i_10_324_4027_0,
    i_10_324_4057_0, i_10_324_4153_0, i_10_324_4175_0, i_10_324_4286_0,
    i_10_324_4375_0, i_10_324_4376_0, i_10_324_4564_0, i_10_324_4568_0;
  output o_10_324_0_0;
  assign o_10_324_0_0 = 0;
endmodule



// Benchmark "kernel_10_325" written by ABC on Sun Jul 19 10:26:41 2020

module kernel_10_325 ( 
    i_10_325_31_0, i_10_325_33_0, i_10_325_40_0, i_10_325_43_0,
    i_10_325_151_0, i_10_325_222_0, i_10_325_248_0, i_10_325_251_0,
    i_10_325_285_0, i_10_325_286_0, i_10_325_287_0, i_10_325_318_0,
    i_10_325_319_0, i_10_325_409_0, i_10_325_410_0, i_10_325_412_0,
    i_10_325_413_0, i_10_325_428_0, i_10_325_434_0, i_10_325_436_0,
    i_10_325_437_0, i_10_325_439_0, i_10_325_520_0, i_10_325_964_0,
    i_10_325_996_0, i_10_325_997_0, i_10_325_1004_0, i_10_325_1030_0,
    i_10_325_1041_0, i_10_325_1042_0, i_10_325_1043_0, i_10_325_1169_0,
    i_10_325_1236_0, i_10_325_1294_0, i_10_325_1311_0, i_10_325_1343_0,
    i_10_325_1344_0, i_10_325_1346_0, i_10_325_1546_0, i_10_325_1653_0,
    i_10_325_1655_0, i_10_325_1735_0, i_10_325_1815_0, i_10_325_1880_0,
    i_10_325_1908_0, i_10_325_1909_0, i_10_325_1913_0, i_10_325_2023_0,
    i_10_325_2245_0, i_10_325_2352_0, i_10_325_2353_0, i_10_325_2354_0,
    i_10_325_2355_0, i_10_325_2365_0, i_10_325_2452_0, i_10_325_2453_0,
    i_10_325_2455_0, i_10_325_2469_0, i_10_325_2471_0, i_10_325_2705_0,
    i_10_325_2724_0, i_10_325_2731_0, i_10_325_2832_0, i_10_325_2833_0,
    i_10_325_2869_0, i_10_325_2886_0, i_10_325_2887_0, i_10_325_3036_0,
    i_10_325_3037_0, i_10_325_3039_0, i_10_325_3045_0, i_10_325_3164_0,
    i_10_325_3166_0, i_10_325_3272_0, i_10_325_3280_0, i_10_325_3301_0,
    i_10_325_3433_0, i_10_325_3523_0, i_10_325_3526_0, i_10_325_3527_0,
    i_10_325_3585_0, i_10_325_3586_0, i_10_325_3611_0, i_10_325_3613_0,
    i_10_325_3616_0, i_10_325_3650_0, i_10_325_3784_0, i_10_325_3838_0,
    i_10_325_3893_0, i_10_325_3994_0, i_10_325_3995_0, i_10_325_4030_0,
    i_10_325_4116_0, i_10_325_4117_0, i_10_325_4172_0, i_10_325_4220_0,
    i_10_325_4273_0, i_10_325_4274_0, i_10_325_4282_0, i_10_325_4283_0,
    o_10_325_0_0  );
  input  i_10_325_31_0, i_10_325_33_0, i_10_325_40_0, i_10_325_43_0,
    i_10_325_151_0, i_10_325_222_0, i_10_325_248_0, i_10_325_251_0,
    i_10_325_285_0, i_10_325_286_0, i_10_325_287_0, i_10_325_318_0,
    i_10_325_319_0, i_10_325_409_0, i_10_325_410_0, i_10_325_412_0,
    i_10_325_413_0, i_10_325_428_0, i_10_325_434_0, i_10_325_436_0,
    i_10_325_437_0, i_10_325_439_0, i_10_325_520_0, i_10_325_964_0,
    i_10_325_996_0, i_10_325_997_0, i_10_325_1004_0, i_10_325_1030_0,
    i_10_325_1041_0, i_10_325_1042_0, i_10_325_1043_0, i_10_325_1169_0,
    i_10_325_1236_0, i_10_325_1294_0, i_10_325_1311_0, i_10_325_1343_0,
    i_10_325_1344_0, i_10_325_1346_0, i_10_325_1546_0, i_10_325_1653_0,
    i_10_325_1655_0, i_10_325_1735_0, i_10_325_1815_0, i_10_325_1880_0,
    i_10_325_1908_0, i_10_325_1909_0, i_10_325_1913_0, i_10_325_2023_0,
    i_10_325_2245_0, i_10_325_2352_0, i_10_325_2353_0, i_10_325_2354_0,
    i_10_325_2355_0, i_10_325_2365_0, i_10_325_2452_0, i_10_325_2453_0,
    i_10_325_2455_0, i_10_325_2469_0, i_10_325_2471_0, i_10_325_2705_0,
    i_10_325_2724_0, i_10_325_2731_0, i_10_325_2832_0, i_10_325_2833_0,
    i_10_325_2869_0, i_10_325_2886_0, i_10_325_2887_0, i_10_325_3036_0,
    i_10_325_3037_0, i_10_325_3039_0, i_10_325_3045_0, i_10_325_3164_0,
    i_10_325_3166_0, i_10_325_3272_0, i_10_325_3280_0, i_10_325_3301_0,
    i_10_325_3433_0, i_10_325_3523_0, i_10_325_3526_0, i_10_325_3527_0,
    i_10_325_3585_0, i_10_325_3586_0, i_10_325_3611_0, i_10_325_3613_0,
    i_10_325_3616_0, i_10_325_3650_0, i_10_325_3784_0, i_10_325_3838_0,
    i_10_325_3893_0, i_10_325_3994_0, i_10_325_3995_0, i_10_325_4030_0,
    i_10_325_4116_0, i_10_325_4117_0, i_10_325_4172_0, i_10_325_4220_0,
    i_10_325_4273_0, i_10_325_4274_0, i_10_325_4282_0, i_10_325_4283_0;
  output o_10_325_0_0;
  assign o_10_325_0_0 = ~((i_10_325_287_0 & ((~i_10_325_251_0 & ~i_10_325_1043_0 & ~i_10_325_1908_0 & ~i_10_325_2471_0 & ~i_10_325_3164_0) | (i_10_325_410_0 & ~i_10_325_997_0 & i_10_325_2455_0 & ~i_10_325_3272_0 & i_10_325_3616_0))) | (~i_10_325_409_0 & ((~i_10_325_439_0 & ~i_10_325_1042_0 & ~i_10_325_1913_0 & ~i_10_325_2887_0 & ~i_10_325_3166_0 & ~i_10_325_3523_0) | (~i_10_325_287_0 & ~i_10_325_437_0 & ~i_10_325_1344_0 & ~i_10_325_1346_0 & ~i_10_325_1655_0 & ~i_10_325_3994_0))) | (~i_10_325_413_0 & ((~i_10_325_318_0 & ~i_10_325_520_0 & ~i_10_325_1042_0 & ~i_10_325_1343_0 & ~i_10_325_1346_0 & ~i_10_325_3586_0) | (~i_10_325_251_0 & i_10_325_1653_0 & ~i_10_325_2455_0 & ~i_10_325_3280_0 & ~i_10_325_3611_0 & ~i_10_325_3616_0 & ~i_10_325_4283_0))) | (~i_10_325_997_0 & ((~i_10_325_437_0 & ~i_10_325_996_0 & ((~i_10_325_410_0 & ~i_10_325_412_0 & ~i_10_325_1042_0 & ~i_10_325_2469_0 & ~i_10_325_3838_0) | (~i_10_325_1041_0 & ~i_10_325_1343_0 & ~i_10_325_4117_0 & ~i_10_325_4273_0))) | (~i_10_325_1344_0 & ~i_10_325_2365_0 & ~i_10_325_2453_0 & ~i_10_325_3280_0 & ~i_10_325_3838_0) | (~i_10_325_251_0 & ~i_10_325_1043_0 & ~i_10_325_1343_0 & ~i_10_325_1908_0 & ~i_10_325_3523_0 & ~i_10_325_4116_0))) | (~i_10_325_251_0 & ((i_10_325_2353_0 & i_10_325_2354_0) | (i_10_325_285_0 & ~i_10_325_1030_0 & ~i_10_325_1909_0 & i_10_325_2705_0 & ~i_10_325_2887_0 & ~i_10_325_4283_0))) | (~i_10_325_410_0 & ((~i_10_325_1346_0 & ~i_10_325_2705_0 & ~i_10_325_2887_0 & ~i_10_325_3527_0 & ~i_10_325_3995_0 & ~i_10_325_4282_0) | (~i_10_325_437_0 & ~i_10_325_1041_0 & ~i_10_325_2471_0 & ~i_10_325_3166_0 & ~i_10_325_3280_0 & ~i_10_325_4283_0))) | (~i_10_325_1042_0 & ~i_10_325_1908_0 & ((~i_10_325_1043_0 & ~i_10_325_1346_0 & ~i_10_325_2023_0 & ~i_10_325_3526_0) | (~i_10_325_319_0 & i_10_325_1653_0 & ~i_10_325_1913_0 & ~i_10_325_3613_0 & ~i_10_325_3650_0))) | (i_10_325_1236_0 & ((i_10_325_3280_0 & ~i_10_325_3527_0 & i_10_325_3616_0) | (i_10_325_1041_0 & ~i_10_325_4273_0))) | (~i_10_325_3995_0 & ((~i_10_325_1909_0 & ((~i_10_325_520_0 & ~i_10_325_2023_0 & i_10_325_2705_0) | (~i_10_325_439_0 & ~i_10_325_1346_0 & ~i_10_325_2453_0 & ~i_10_325_3994_0))) | (~i_10_325_2832_0 & ~i_10_325_2887_0 & ~i_10_325_3036_0 & i_10_325_3433_0 & ~i_10_325_3611_0 & ~i_10_325_4117_0))) | (i_10_325_410_0 & ~i_10_325_3611_0 & ~i_10_325_3838_0 & ~i_10_325_3994_0 & ~i_10_325_4117_0 & ~i_10_325_4220_0) | (~i_10_325_1169_0 & ~i_10_325_1913_0 & i_10_325_2469_0 & ~i_10_325_4283_0));
endmodule



// Benchmark "kernel_10_326" written by ABC on Sun Jul 19 10:26:43 2020

module kernel_10_326 ( 
    i_10_326_171_0, i_10_326_174_0, i_10_326_221_0, i_10_326_244_0,
    i_10_326_263_0, i_10_326_280_0, i_10_326_282_0, i_10_326_283_0,
    i_10_326_320_0, i_10_326_390_0, i_10_326_393_0, i_10_326_406_0,
    i_10_326_409_0, i_10_326_445_0, i_10_326_446_0, i_10_326_448_0,
    i_10_326_451_0, i_10_326_460_0, i_10_326_466_0, i_10_326_560_0,
    i_10_326_589_0, i_10_326_699_0, i_10_326_748_0, i_10_326_797_0,
    i_10_326_906_0, i_10_326_954_0, i_10_326_1002_0, i_10_326_1005_0,
    i_10_326_1027_0, i_10_326_1032_0, i_10_326_1238_0, i_10_326_1305_0,
    i_10_326_1307_0, i_10_326_1348_0, i_10_326_1447_0, i_10_326_1626_0,
    i_10_326_1651_0, i_10_326_1652_0, i_10_326_1655_0, i_10_326_1767_0,
    i_10_326_1768_0, i_10_326_1769_0, i_10_326_1818_0, i_10_326_1819_0,
    i_10_326_1821_0, i_10_326_1824_0, i_10_326_1910_0, i_10_326_1911_0,
    i_10_326_1949_0, i_10_326_1995_0, i_10_326_2310_0, i_10_326_2334_0,
    i_10_326_2376_0, i_10_326_2384_0, i_10_326_2460_0, i_10_326_2461_0,
    i_10_326_2565_0, i_10_326_2647_0, i_10_326_2658_0, i_10_326_2679_0,
    i_10_326_2704_0, i_10_326_2718_0, i_10_326_2721_0, i_10_326_2728_0,
    i_10_326_2826_0, i_10_326_2829_0, i_10_326_2830_0, i_10_326_2831_0,
    i_10_326_2921_0, i_10_326_2924_0, i_10_326_3157_0, i_10_326_3280_0,
    i_10_326_3386_0, i_10_326_3387_0, i_10_326_3388_0, i_10_326_3403_0,
    i_10_326_3436_0, i_10_326_3437_0, i_10_326_3540_0, i_10_326_3541_0,
    i_10_326_3550_0, i_10_326_3610_0, i_10_326_3835_0, i_10_326_3853_0,
    i_10_326_3854_0, i_10_326_3855_0, i_10_326_3856_0, i_10_326_3860_0,
    i_10_326_3984_0, i_10_326_4025_0, i_10_326_4026_0, i_10_326_4027_0,
    i_10_326_4117_0, i_10_326_4118_0, i_10_326_4120_0, i_10_326_4122_0,
    i_10_326_4128_0, i_10_326_4174_0, i_10_326_4548_0, i_10_326_4571_0,
    o_10_326_0_0  );
  input  i_10_326_171_0, i_10_326_174_0, i_10_326_221_0, i_10_326_244_0,
    i_10_326_263_0, i_10_326_280_0, i_10_326_282_0, i_10_326_283_0,
    i_10_326_320_0, i_10_326_390_0, i_10_326_393_0, i_10_326_406_0,
    i_10_326_409_0, i_10_326_445_0, i_10_326_446_0, i_10_326_448_0,
    i_10_326_451_0, i_10_326_460_0, i_10_326_466_0, i_10_326_560_0,
    i_10_326_589_0, i_10_326_699_0, i_10_326_748_0, i_10_326_797_0,
    i_10_326_906_0, i_10_326_954_0, i_10_326_1002_0, i_10_326_1005_0,
    i_10_326_1027_0, i_10_326_1032_0, i_10_326_1238_0, i_10_326_1305_0,
    i_10_326_1307_0, i_10_326_1348_0, i_10_326_1447_0, i_10_326_1626_0,
    i_10_326_1651_0, i_10_326_1652_0, i_10_326_1655_0, i_10_326_1767_0,
    i_10_326_1768_0, i_10_326_1769_0, i_10_326_1818_0, i_10_326_1819_0,
    i_10_326_1821_0, i_10_326_1824_0, i_10_326_1910_0, i_10_326_1911_0,
    i_10_326_1949_0, i_10_326_1995_0, i_10_326_2310_0, i_10_326_2334_0,
    i_10_326_2376_0, i_10_326_2384_0, i_10_326_2460_0, i_10_326_2461_0,
    i_10_326_2565_0, i_10_326_2647_0, i_10_326_2658_0, i_10_326_2679_0,
    i_10_326_2704_0, i_10_326_2718_0, i_10_326_2721_0, i_10_326_2728_0,
    i_10_326_2826_0, i_10_326_2829_0, i_10_326_2830_0, i_10_326_2831_0,
    i_10_326_2921_0, i_10_326_2924_0, i_10_326_3157_0, i_10_326_3280_0,
    i_10_326_3386_0, i_10_326_3387_0, i_10_326_3388_0, i_10_326_3403_0,
    i_10_326_3436_0, i_10_326_3437_0, i_10_326_3540_0, i_10_326_3541_0,
    i_10_326_3550_0, i_10_326_3610_0, i_10_326_3835_0, i_10_326_3853_0,
    i_10_326_3854_0, i_10_326_3855_0, i_10_326_3856_0, i_10_326_3860_0,
    i_10_326_3984_0, i_10_326_4025_0, i_10_326_4026_0, i_10_326_4027_0,
    i_10_326_4117_0, i_10_326_4118_0, i_10_326_4120_0, i_10_326_4122_0,
    i_10_326_4128_0, i_10_326_4174_0, i_10_326_4548_0, i_10_326_4571_0;
  output o_10_326_0_0;
  assign o_10_326_0_0 = ~((~i_10_326_171_0 & ((~i_10_326_699_0 & ~i_10_326_1305_0 & ~i_10_326_1911_0 & ~i_10_326_3280_0 & ~i_10_326_3436_0 & ~i_10_326_3550_0 & ~i_10_326_3860_0 & ~i_10_326_4026_0 & ~i_10_326_4128_0) | (~i_10_326_390_0 & ~i_10_326_1002_0 & ~i_10_326_1767_0 & ~i_10_326_1995_0 & ~i_10_326_2310_0 & ~i_10_326_2679_0 & ~i_10_326_2831_0 & i_10_326_3387_0 & ~i_10_326_3853_0 & ~i_10_326_4571_0))) | (~i_10_326_1002_0 & ((~i_10_326_283_0 & ((~i_10_326_460_0 & ~i_10_326_1027_0 & ~i_10_326_1238_0 & ~i_10_326_2460_0 & ~i_10_326_3835_0) | (~i_10_326_1768_0 & ~i_10_326_3280_0 & ~i_10_326_3550_0 & ~i_10_326_4026_0))) | (~i_10_326_3984_0 & ((~i_10_326_699_0 & ((~i_10_326_221_0 & ~i_10_326_1032_0 & ~i_10_326_1767_0 & ~i_10_326_1768_0 & ~i_10_326_2310_0 & ~i_10_326_2565_0 & ~i_10_326_2721_0 & ~i_10_326_3550_0) | (~i_10_326_390_0 & ~i_10_326_2728_0 & ~i_10_326_2829_0 & ~i_10_326_3437_0 & ~i_10_326_3610_0 & ~i_10_326_4571_0))) | (~i_10_326_393_0 & i_10_326_1238_0 & ~i_10_326_1995_0 & ~i_10_326_2461_0 & ~i_10_326_4118_0))) | (~i_10_326_320_0 & ~i_10_326_1769_0 & ~i_10_326_2310_0 & ~i_10_326_2334_0 & ~i_10_326_2565_0 & ~i_10_326_3387_0) | (~i_10_326_2461_0 & ~i_10_326_2679_0 & ~i_10_326_3437_0 & ~i_10_326_3550_0 & i_10_326_4118_0 & ~i_10_326_4128_0))) | (~i_10_326_446_0 & ((i_10_326_1238_0 & ~i_10_326_1305_0 & ~i_10_326_1307_0 & ~i_10_326_2376_0 & ~i_10_326_3856_0) | (~i_10_326_393_0 & ~i_10_326_2310_0 & i_10_326_3984_0 & i_10_326_4025_0))) | (~i_10_326_2310_0 & ((~i_10_326_1027_0 & ~i_10_326_2728_0 & i_10_326_4026_0 & ((~i_10_326_174_0 & ~i_10_326_797_0 & i_10_326_1032_0 & ~i_10_326_1824_0 & i_10_326_3860_0) | (~i_10_326_282_0 & ~i_10_326_1652_0 & ~i_10_326_2679_0 & ~i_10_326_2830_0 & ~i_10_326_4122_0 & ~i_10_326_4174_0))) | (~i_10_326_1032_0 & ~i_10_326_1769_0 & ~i_10_326_2658_0 & ~i_10_326_3437_0 & ~i_10_326_4026_0 & ~i_10_326_4122_0) | (~i_10_326_320_0 & ~i_10_326_451_0 & ~i_10_326_699_0 & ~i_10_326_1307_0 & ~i_10_326_1821_0 & ~i_10_326_1995_0 & ~i_10_326_3403_0 & ~i_10_326_3436_0 & ~i_10_326_3550_0 & ~i_10_326_4120_0 & ~i_10_326_4128_0 & ~i_10_326_4571_0))) | (~i_10_326_393_0 & ((~i_10_326_699_0 & ((~i_10_326_906_0 & ~i_10_326_1626_0 & ~i_10_326_1911_0 & ~i_10_326_2565_0 & ~i_10_326_3550_0 & ~i_10_326_3856_0 & i_10_326_4026_0) | (~i_10_326_390_0 & ~i_10_326_1767_0 & ~i_10_326_1769_0 & ~i_10_326_2460_0 & ~i_10_326_4026_0))) | (~i_10_326_2460_0 & ~i_10_326_2704_0 & ~i_10_326_2718_0 & ~i_10_326_3856_0 & ~i_10_326_4120_0 & ~i_10_326_4122_0))) | (~i_10_326_390_0 & ((i_10_326_446_0 & ~i_10_326_3280_0 & ~i_10_326_4026_0) | (~i_10_326_2728_0 & ~i_10_326_3387_0 & ~i_10_326_3388_0 & i_10_326_3835_0 & ~i_10_326_4174_0))) | (i_10_326_1655_0 & (i_10_326_1819_0 | (~i_10_326_448_0 & ~i_10_326_1767_0 & ~i_10_326_2721_0 & ~i_10_326_3280_0))) | (~i_10_326_3853_0 & ((i_10_326_283_0 & ~i_10_326_445_0 & ~i_10_326_1005_0 & ~i_10_326_1767_0 & ~i_10_326_2721_0 & ~i_10_326_2831_0 & ~i_10_326_4122_0) | (~i_10_326_954_0 & i_10_326_1819_0 & ~i_10_326_1824_0 & i_10_326_4174_0))) | (~i_10_326_3984_0 & ((~i_10_326_3388_0 & ~i_10_326_4026_0) | (~i_10_326_460_0 & ~i_10_326_1447_0 & ~i_10_326_2376_0 & ~i_10_326_2461_0 & ~i_10_326_3280_0 & ~i_10_326_3436_0 & ~i_10_326_4128_0))) | (~i_10_326_466_0 & ~i_10_326_2830_0 & i_10_326_4117_0));
endmodule



// Benchmark "kernel_10_327" written by ABC on Sun Jul 19 10:26:43 2020

module kernel_10_327 ( 
    i_10_327_32_0, i_10_327_158_0, i_10_327_185_0, i_10_327_284_0,
    i_10_327_390_0, i_10_327_391_0, i_10_327_392_0, i_10_327_436_0,
    i_10_327_437_0, i_10_327_443_0, i_10_327_464_0, i_10_327_718_0,
    i_10_327_854_0, i_10_327_955_0, i_10_327_961_0, i_10_327_964_0,
    i_10_327_992_0, i_10_327_1003_0, i_10_327_1036_0, i_10_327_1043_0,
    i_10_327_1045_0, i_10_327_1058_0, i_10_327_1082_0, i_10_327_1083_0,
    i_10_327_1120_0, i_10_327_1240_0, i_10_327_1247_0, i_10_327_1268_0,
    i_10_327_1365_0, i_10_327_1366_0, i_10_327_1367_0, i_10_327_1380_0,
    i_10_327_1436_0, i_10_327_1443_0, i_10_327_1448_0, i_10_327_1489_0,
    i_10_327_1597_0, i_10_327_1651_0, i_10_327_1772_0, i_10_327_1797_0,
    i_10_327_1806_0, i_10_327_1919_0, i_10_327_1954_0, i_10_327_2018_0,
    i_10_327_2095_0, i_10_327_2096_0, i_10_327_2349_0, i_10_327_2357_0,
    i_10_327_2362_0, i_10_327_2366_0, i_10_327_2381_0, i_10_327_2465_0,
    i_10_327_2492_0, i_10_327_2511_0, i_10_327_2514_0, i_10_327_2560_0,
    i_10_327_2565_0, i_10_327_2603_0, i_10_327_2659_0, i_10_327_2660_0,
    i_10_327_2702_0, i_10_327_2743_0, i_10_327_2744_0, i_10_327_2781_0,
    i_10_327_2782_0, i_10_327_2831_0, i_10_327_2834_0, i_10_327_3159_0,
    i_10_327_3162_0, i_10_327_3283_0, i_10_327_3284_0, i_10_327_3450_0,
    i_10_327_3452_0, i_10_327_3470_0, i_10_327_3703_0, i_10_327_3704_0,
    i_10_327_3747_0, i_10_327_3835_0, i_10_327_3853_0, i_10_327_3879_0,
    i_10_327_3923_0, i_10_327_4056_0, i_10_327_4057_0, i_10_327_4114_0,
    i_10_327_4144_0, i_10_327_4220_0, i_10_327_4237_0, i_10_327_4238_0,
    i_10_327_4268_0, i_10_327_4275_0, i_10_327_4278_0, i_10_327_4280_0,
    i_10_327_4282_0, i_10_327_4342_0, i_10_327_4436_0, i_10_327_4521_0,
    i_10_327_4522_0, i_10_327_4523_0, i_10_327_4565_0, i_10_327_4571_0,
    o_10_327_0_0  );
  input  i_10_327_32_0, i_10_327_158_0, i_10_327_185_0, i_10_327_284_0,
    i_10_327_390_0, i_10_327_391_0, i_10_327_392_0, i_10_327_436_0,
    i_10_327_437_0, i_10_327_443_0, i_10_327_464_0, i_10_327_718_0,
    i_10_327_854_0, i_10_327_955_0, i_10_327_961_0, i_10_327_964_0,
    i_10_327_992_0, i_10_327_1003_0, i_10_327_1036_0, i_10_327_1043_0,
    i_10_327_1045_0, i_10_327_1058_0, i_10_327_1082_0, i_10_327_1083_0,
    i_10_327_1120_0, i_10_327_1240_0, i_10_327_1247_0, i_10_327_1268_0,
    i_10_327_1365_0, i_10_327_1366_0, i_10_327_1367_0, i_10_327_1380_0,
    i_10_327_1436_0, i_10_327_1443_0, i_10_327_1448_0, i_10_327_1489_0,
    i_10_327_1597_0, i_10_327_1651_0, i_10_327_1772_0, i_10_327_1797_0,
    i_10_327_1806_0, i_10_327_1919_0, i_10_327_1954_0, i_10_327_2018_0,
    i_10_327_2095_0, i_10_327_2096_0, i_10_327_2349_0, i_10_327_2357_0,
    i_10_327_2362_0, i_10_327_2366_0, i_10_327_2381_0, i_10_327_2465_0,
    i_10_327_2492_0, i_10_327_2511_0, i_10_327_2514_0, i_10_327_2560_0,
    i_10_327_2565_0, i_10_327_2603_0, i_10_327_2659_0, i_10_327_2660_0,
    i_10_327_2702_0, i_10_327_2743_0, i_10_327_2744_0, i_10_327_2781_0,
    i_10_327_2782_0, i_10_327_2831_0, i_10_327_2834_0, i_10_327_3159_0,
    i_10_327_3162_0, i_10_327_3283_0, i_10_327_3284_0, i_10_327_3450_0,
    i_10_327_3452_0, i_10_327_3470_0, i_10_327_3703_0, i_10_327_3704_0,
    i_10_327_3747_0, i_10_327_3835_0, i_10_327_3853_0, i_10_327_3879_0,
    i_10_327_3923_0, i_10_327_4056_0, i_10_327_4057_0, i_10_327_4114_0,
    i_10_327_4144_0, i_10_327_4220_0, i_10_327_4237_0, i_10_327_4238_0,
    i_10_327_4268_0, i_10_327_4275_0, i_10_327_4278_0, i_10_327_4280_0,
    i_10_327_4282_0, i_10_327_4342_0, i_10_327_4436_0, i_10_327_4521_0,
    i_10_327_4522_0, i_10_327_4523_0, i_10_327_4565_0, i_10_327_4571_0;
  output o_10_327_0_0;
  assign o_10_327_0_0 = 0;
endmodule



// Benchmark "kernel_10_328" written by ABC on Sun Jul 19 10:26:44 2020

module kernel_10_328 ( 
    i_10_328_48_0, i_10_328_174_0, i_10_328_175_0, i_10_328_220_0,
    i_10_328_279_0, i_10_328_282_0, i_10_328_283_0, i_10_328_329_0,
    i_10_328_445_0, i_10_328_446_0, i_10_328_459_0, i_10_328_460_0,
    i_10_328_462_0, i_10_328_463_0, i_10_328_685_0, i_10_328_686_0,
    i_10_328_748_0, i_10_328_828_0, i_10_328_963_0, i_10_328_990_0,
    i_10_328_997_0, i_10_328_1026_0, i_10_328_1035_0, i_10_328_1036_0,
    i_10_328_1161_0, i_10_328_1162_0, i_10_328_1266_0, i_10_328_1268_0,
    i_10_328_1288_0, i_10_328_1306_0, i_10_328_1307_0, i_10_328_1486_0,
    i_10_328_1532_0, i_10_328_1551_0, i_10_328_1562_0, i_10_328_1647_0,
    i_10_328_1648_0, i_10_328_1649_0, i_10_328_1683_0, i_10_328_1766_0,
    i_10_328_1823_0, i_10_328_1825_0, i_10_328_1917_0, i_10_328_1946_0,
    i_10_328_2353_0, i_10_328_2448_0, i_10_328_2451_0, i_10_328_2452_0,
    i_10_328_2454_0, i_10_328_2472_0, i_10_328_2473_0, i_10_328_2503_0,
    i_10_328_2539_0, i_10_328_2603_0, i_10_328_2605_0, i_10_328_2629_0,
    i_10_328_2630_0, i_10_328_2632_0, i_10_328_2657_0, i_10_328_2658_0,
    i_10_328_2661_0, i_10_328_2726_0, i_10_328_2727_0, i_10_328_2787_0,
    i_10_328_2817_0, i_10_328_2820_0, i_10_328_2822_0, i_10_328_2826_0,
    i_10_328_2827_0, i_10_328_2828_0, i_10_328_2880_0, i_10_328_2881_0,
    i_10_328_3034_0, i_10_328_3035_0, i_10_328_3282_0, i_10_328_3312_0,
    i_10_328_3313_0, i_10_328_3384_0, i_10_328_3388_0, i_10_328_3522_0,
    i_10_328_3523_0, i_10_328_3525_0, i_10_328_3526_0, i_10_328_3646_0,
    i_10_328_3840_0, i_10_328_3980_0, i_10_328_3987_0, i_10_328_3998_0,
    i_10_328_4113_0, i_10_328_4115_0, i_10_328_4117_0, i_10_328_4168_0,
    i_10_328_4275_0, i_10_328_4284_0, i_10_328_4285_0, i_10_328_4287_0,
    i_10_328_4288_0, i_10_328_4456_0, i_10_328_4563_0, i_10_328_4564_0,
    o_10_328_0_0  );
  input  i_10_328_48_0, i_10_328_174_0, i_10_328_175_0, i_10_328_220_0,
    i_10_328_279_0, i_10_328_282_0, i_10_328_283_0, i_10_328_329_0,
    i_10_328_445_0, i_10_328_446_0, i_10_328_459_0, i_10_328_460_0,
    i_10_328_462_0, i_10_328_463_0, i_10_328_685_0, i_10_328_686_0,
    i_10_328_748_0, i_10_328_828_0, i_10_328_963_0, i_10_328_990_0,
    i_10_328_997_0, i_10_328_1026_0, i_10_328_1035_0, i_10_328_1036_0,
    i_10_328_1161_0, i_10_328_1162_0, i_10_328_1266_0, i_10_328_1268_0,
    i_10_328_1288_0, i_10_328_1306_0, i_10_328_1307_0, i_10_328_1486_0,
    i_10_328_1532_0, i_10_328_1551_0, i_10_328_1562_0, i_10_328_1647_0,
    i_10_328_1648_0, i_10_328_1649_0, i_10_328_1683_0, i_10_328_1766_0,
    i_10_328_1823_0, i_10_328_1825_0, i_10_328_1917_0, i_10_328_1946_0,
    i_10_328_2353_0, i_10_328_2448_0, i_10_328_2451_0, i_10_328_2452_0,
    i_10_328_2454_0, i_10_328_2472_0, i_10_328_2473_0, i_10_328_2503_0,
    i_10_328_2539_0, i_10_328_2603_0, i_10_328_2605_0, i_10_328_2629_0,
    i_10_328_2630_0, i_10_328_2632_0, i_10_328_2657_0, i_10_328_2658_0,
    i_10_328_2661_0, i_10_328_2726_0, i_10_328_2727_0, i_10_328_2787_0,
    i_10_328_2817_0, i_10_328_2820_0, i_10_328_2822_0, i_10_328_2826_0,
    i_10_328_2827_0, i_10_328_2828_0, i_10_328_2880_0, i_10_328_2881_0,
    i_10_328_3034_0, i_10_328_3035_0, i_10_328_3282_0, i_10_328_3312_0,
    i_10_328_3313_0, i_10_328_3384_0, i_10_328_3388_0, i_10_328_3522_0,
    i_10_328_3523_0, i_10_328_3525_0, i_10_328_3526_0, i_10_328_3646_0,
    i_10_328_3840_0, i_10_328_3980_0, i_10_328_3987_0, i_10_328_3998_0,
    i_10_328_4113_0, i_10_328_4115_0, i_10_328_4117_0, i_10_328_4168_0,
    i_10_328_4275_0, i_10_328_4284_0, i_10_328_4285_0, i_10_328_4287_0,
    i_10_328_4288_0, i_10_328_4456_0, i_10_328_4563_0, i_10_328_4564_0;
  output o_10_328_0_0;
  assign o_10_328_0_0 = 0;
endmodule



// Benchmark "kernel_10_329" written by ABC on Sun Jul 19 10:26:45 2020

module kernel_10_329 ( 
    i_10_329_175_0, i_10_329_267_0, i_10_329_281_0, i_10_329_284_0,
    i_10_329_286_0, i_10_329_393_0, i_10_329_405_0, i_10_329_406_0,
    i_10_329_408_0, i_10_329_409_0, i_10_329_412_0, i_10_329_439_0,
    i_10_329_444_0, i_10_329_447_0, i_10_329_448_0, i_10_329_462_0,
    i_10_329_467_0, i_10_329_713_0, i_10_329_793_0, i_10_329_798_0,
    i_10_329_1002_0, i_10_329_1005_0, i_10_329_1054_0, i_10_329_1061_0,
    i_10_329_1122_0, i_10_329_1215_0, i_10_329_1239_0, i_10_329_1247_0,
    i_10_329_1249_0, i_10_329_1296_0, i_10_329_1313_0, i_10_329_1437_0,
    i_10_329_1542_0, i_10_329_1626_0, i_10_329_1650_0, i_10_329_1684_0,
    i_10_329_1685_0, i_10_329_1686_0, i_10_329_1728_0, i_10_329_1730_0,
    i_10_329_1768_0, i_10_329_1821_0, i_10_329_1914_0, i_10_329_1915_0,
    i_10_329_1952_0, i_10_329_2025_0, i_10_329_2029_0, i_10_329_2324_0,
    i_10_329_2327_0, i_10_329_2355_0, i_10_329_2453_0, i_10_329_2454_0,
    i_10_329_2455_0, i_10_329_2469_0, i_10_329_2517_0, i_10_329_2565_0,
    i_10_329_2628_0, i_10_329_2632_0, i_10_329_2634_0, i_10_329_2636_0,
    i_10_329_2655_0, i_10_329_2658_0, i_10_329_2659_0, i_10_329_2662_0,
    i_10_329_2663_0, i_10_329_2678_0, i_10_329_2702_0, i_10_329_2704_0,
    i_10_329_2706_0, i_10_329_2711_0, i_10_329_2725_0, i_10_329_2730_0,
    i_10_329_2732_0, i_10_329_2737_0, i_10_329_2784_0, i_10_329_2785_0,
    i_10_329_2804_0, i_10_329_2954_0, i_10_329_2979_0, i_10_329_2996_0,
    i_10_329_3033_0, i_10_329_3071_0, i_10_329_3279_0, i_10_329_3284_0,
    i_10_329_3320_0, i_10_329_3388_0, i_10_329_3389_0, i_10_329_3471_0,
    i_10_329_3525_0, i_10_329_3545_0, i_10_329_3561_0, i_10_329_3586_0,
    i_10_329_3613_0, i_10_329_3780_0, i_10_329_3784_0, i_10_329_3837_0,
    i_10_329_3859_0, i_10_329_4117_0, i_10_329_4124_0, i_10_329_4272_0,
    o_10_329_0_0  );
  input  i_10_329_175_0, i_10_329_267_0, i_10_329_281_0, i_10_329_284_0,
    i_10_329_286_0, i_10_329_393_0, i_10_329_405_0, i_10_329_406_0,
    i_10_329_408_0, i_10_329_409_0, i_10_329_412_0, i_10_329_439_0,
    i_10_329_444_0, i_10_329_447_0, i_10_329_448_0, i_10_329_462_0,
    i_10_329_467_0, i_10_329_713_0, i_10_329_793_0, i_10_329_798_0,
    i_10_329_1002_0, i_10_329_1005_0, i_10_329_1054_0, i_10_329_1061_0,
    i_10_329_1122_0, i_10_329_1215_0, i_10_329_1239_0, i_10_329_1247_0,
    i_10_329_1249_0, i_10_329_1296_0, i_10_329_1313_0, i_10_329_1437_0,
    i_10_329_1542_0, i_10_329_1626_0, i_10_329_1650_0, i_10_329_1684_0,
    i_10_329_1685_0, i_10_329_1686_0, i_10_329_1728_0, i_10_329_1730_0,
    i_10_329_1768_0, i_10_329_1821_0, i_10_329_1914_0, i_10_329_1915_0,
    i_10_329_1952_0, i_10_329_2025_0, i_10_329_2029_0, i_10_329_2324_0,
    i_10_329_2327_0, i_10_329_2355_0, i_10_329_2453_0, i_10_329_2454_0,
    i_10_329_2455_0, i_10_329_2469_0, i_10_329_2517_0, i_10_329_2565_0,
    i_10_329_2628_0, i_10_329_2632_0, i_10_329_2634_0, i_10_329_2636_0,
    i_10_329_2655_0, i_10_329_2658_0, i_10_329_2659_0, i_10_329_2662_0,
    i_10_329_2663_0, i_10_329_2678_0, i_10_329_2702_0, i_10_329_2704_0,
    i_10_329_2706_0, i_10_329_2711_0, i_10_329_2725_0, i_10_329_2730_0,
    i_10_329_2732_0, i_10_329_2737_0, i_10_329_2784_0, i_10_329_2785_0,
    i_10_329_2804_0, i_10_329_2954_0, i_10_329_2979_0, i_10_329_2996_0,
    i_10_329_3033_0, i_10_329_3071_0, i_10_329_3279_0, i_10_329_3284_0,
    i_10_329_3320_0, i_10_329_3388_0, i_10_329_3389_0, i_10_329_3471_0,
    i_10_329_3525_0, i_10_329_3545_0, i_10_329_3561_0, i_10_329_3586_0,
    i_10_329_3613_0, i_10_329_3780_0, i_10_329_3784_0, i_10_329_3837_0,
    i_10_329_3859_0, i_10_329_4117_0, i_10_329_4124_0, i_10_329_4272_0;
  output o_10_329_0_0;
  assign o_10_329_0_0 = 0;
endmodule



// Benchmark "kernel_10_330" written by ABC on Sun Jul 19 10:26:46 2020

module kernel_10_330 ( 
    i_10_330_33_0, i_10_330_34_0, i_10_330_123_0, i_10_330_143_0,
    i_10_330_256_0, i_10_330_265_0, i_10_330_266_0, i_10_330_272_0,
    i_10_330_274_0, i_10_330_275_0, i_10_330_283_0, i_10_330_432_0,
    i_10_330_448_0, i_10_330_449_0, i_10_330_498_0, i_10_330_501_0,
    i_10_330_502_0, i_10_330_506_0, i_10_330_564_0, i_10_330_565_0,
    i_10_330_628_0, i_10_330_719_0, i_10_330_745_0, i_10_330_753_0,
    i_10_330_1005_0, i_10_330_1030_0, i_10_330_1034_0, i_10_330_1111_0,
    i_10_330_1115_0, i_10_330_1165_0, i_10_330_1213_0, i_10_330_1240_0,
    i_10_330_1243_0, i_10_330_1261_0, i_10_330_1302_0, i_10_330_1303_0,
    i_10_330_1326_0, i_10_330_1348_0, i_10_330_1435_0, i_10_330_1439_0,
    i_10_330_1542_0, i_10_330_1583_0, i_10_330_1732_0, i_10_330_1820_0,
    i_10_330_1821_0, i_10_330_1950_0, i_10_330_1959_0, i_10_330_2035_0,
    i_10_330_2204_0, i_10_330_2294_0, i_10_330_2350_0, i_10_330_2351_0,
    i_10_330_2354_0, i_10_330_2355_0, i_10_330_2408_0, i_10_330_2515_0,
    i_10_330_2533_0, i_10_330_2560_0, i_10_330_2714_0, i_10_330_2744_0,
    i_10_330_2760_0, i_10_330_2761_0, i_10_330_2785_0, i_10_330_2839_0,
    i_10_330_2840_0, i_10_330_2851_0, i_10_330_2869_0, i_10_330_2870_0,
    i_10_330_2885_0, i_10_330_2968_0, i_10_330_2969_0, i_10_330_3048_0,
    i_10_330_3049_0, i_10_330_3195_0, i_10_330_3200_0, i_10_330_3337_0,
    i_10_330_3388_0, i_10_330_3435_0, i_10_330_3504_0, i_10_330_3543_0,
    i_10_330_3544_0, i_10_330_3649_0, i_10_330_3651_0, i_10_330_3747_0,
    i_10_330_3797_0, i_10_330_3804_0, i_10_330_3853_0, i_10_330_3857_0,
    i_10_330_3984_0, i_10_330_4000_0, i_10_330_4117_0, i_10_330_4210_0,
    i_10_330_4211_0, i_10_330_4269_0, i_10_330_4272_0, i_10_330_4273_0,
    i_10_330_4291_0, i_10_330_4392_0, i_10_330_4564_0, i_10_330_4589_0,
    o_10_330_0_0  );
  input  i_10_330_33_0, i_10_330_34_0, i_10_330_123_0, i_10_330_143_0,
    i_10_330_256_0, i_10_330_265_0, i_10_330_266_0, i_10_330_272_0,
    i_10_330_274_0, i_10_330_275_0, i_10_330_283_0, i_10_330_432_0,
    i_10_330_448_0, i_10_330_449_0, i_10_330_498_0, i_10_330_501_0,
    i_10_330_502_0, i_10_330_506_0, i_10_330_564_0, i_10_330_565_0,
    i_10_330_628_0, i_10_330_719_0, i_10_330_745_0, i_10_330_753_0,
    i_10_330_1005_0, i_10_330_1030_0, i_10_330_1034_0, i_10_330_1111_0,
    i_10_330_1115_0, i_10_330_1165_0, i_10_330_1213_0, i_10_330_1240_0,
    i_10_330_1243_0, i_10_330_1261_0, i_10_330_1302_0, i_10_330_1303_0,
    i_10_330_1326_0, i_10_330_1348_0, i_10_330_1435_0, i_10_330_1439_0,
    i_10_330_1542_0, i_10_330_1583_0, i_10_330_1732_0, i_10_330_1820_0,
    i_10_330_1821_0, i_10_330_1950_0, i_10_330_1959_0, i_10_330_2035_0,
    i_10_330_2204_0, i_10_330_2294_0, i_10_330_2350_0, i_10_330_2351_0,
    i_10_330_2354_0, i_10_330_2355_0, i_10_330_2408_0, i_10_330_2515_0,
    i_10_330_2533_0, i_10_330_2560_0, i_10_330_2714_0, i_10_330_2744_0,
    i_10_330_2760_0, i_10_330_2761_0, i_10_330_2785_0, i_10_330_2839_0,
    i_10_330_2840_0, i_10_330_2851_0, i_10_330_2869_0, i_10_330_2870_0,
    i_10_330_2885_0, i_10_330_2968_0, i_10_330_2969_0, i_10_330_3048_0,
    i_10_330_3049_0, i_10_330_3195_0, i_10_330_3200_0, i_10_330_3337_0,
    i_10_330_3388_0, i_10_330_3435_0, i_10_330_3504_0, i_10_330_3543_0,
    i_10_330_3544_0, i_10_330_3649_0, i_10_330_3651_0, i_10_330_3747_0,
    i_10_330_3797_0, i_10_330_3804_0, i_10_330_3853_0, i_10_330_3857_0,
    i_10_330_3984_0, i_10_330_4000_0, i_10_330_4117_0, i_10_330_4210_0,
    i_10_330_4211_0, i_10_330_4269_0, i_10_330_4272_0, i_10_330_4273_0,
    i_10_330_4291_0, i_10_330_4392_0, i_10_330_4564_0, i_10_330_4589_0;
  output o_10_330_0_0;
  assign o_10_330_0_0 = 0;
endmodule



// Benchmark "kernel_10_331" written by ABC on Sun Jul 19 10:26:47 2020

module kernel_10_331 ( 
    i_10_331_49_0, i_10_331_173_0, i_10_331_409_0, i_10_331_460_0,
    i_10_331_464_0, i_10_331_496_0, i_10_331_700_0, i_10_331_712_0,
    i_10_331_713_0, i_10_331_718_0, i_10_331_748_0, i_10_331_749_0,
    i_10_331_752_0, i_10_331_893_0, i_10_331_949_0, i_10_331_1028_0,
    i_10_331_1163_0, i_10_331_1235_0, i_10_331_1236_0, i_10_331_1237_0,
    i_10_331_1264_0, i_10_331_1306_0, i_10_331_1307_0, i_10_331_1308_0,
    i_10_331_1309_0, i_10_331_1310_0, i_10_331_1313_0, i_10_331_1577_0,
    i_10_331_1612_0, i_10_331_1684_0, i_10_331_1685_0, i_10_331_1688_0,
    i_10_331_1766_0, i_10_331_1812_0, i_10_331_1813_0, i_10_331_1821_0,
    i_10_331_2180_0, i_10_331_2359_0, i_10_331_2448_0, i_10_331_2467_0,
    i_10_331_2526_0, i_10_331_2606_0, i_10_331_2631_0, i_10_331_2641_0,
    i_10_331_2657_0, i_10_331_2660_0, i_10_331_2701_0, i_10_331_2702_0,
    i_10_331_2711_0, i_10_331_2719_0, i_10_331_2720_0, i_10_331_2728_0,
    i_10_331_2733_0, i_10_331_2818_0, i_10_331_2830_0, i_10_331_2831_0,
    i_10_331_2833_0, i_10_331_2884_0, i_10_331_2885_0, i_10_331_2921_0,
    i_10_331_2923_0, i_10_331_3070_0, i_10_331_3233_0, i_10_331_3268_0,
    i_10_331_3269_0, i_10_331_3280_0, i_10_331_3297_0, i_10_331_3385_0,
    i_10_331_3386_0, i_10_331_3390_0, i_10_331_3391_0, i_10_331_3392_0,
    i_10_331_3406_0, i_10_331_3462_0, i_10_331_3523_0, i_10_331_3585_0,
    i_10_331_3613_0, i_10_331_3614_0, i_10_331_3647_0, i_10_331_3649_0,
    i_10_331_3650_0, i_10_331_3727_0, i_10_331_3732_0, i_10_331_3781_0,
    i_10_331_3782_0, i_10_331_3783_0, i_10_331_3784_0, i_10_331_3787_0,
    i_10_331_3835_0, i_10_331_3837_0, i_10_331_3888_0, i_10_331_3909_0,
    i_10_331_4115_0, i_10_331_4125_0, i_10_331_4169_0, i_10_331_4212_0,
    i_10_331_4285_0, i_10_331_4286_0, i_10_331_4518_0, i_10_331_4565_0,
    o_10_331_0_0  );
  input  i_10_331_49_0, i_10_331_173_0, i_10_331_409_0, i_10_331_460_0,
    i_10_331_464_0, i_10_331_496_0, i_10_331_700_0, i_10_331_712_0,
    i_10_331_713_0, i_10_331_718_0, i_10_331_748_0, i_10_331_749_0,
    i_10_331_752_0, i_10_331_893_0, i_10_331_949_0, i_10_331_1028_0,
    i_10_331_1163_0, i_10_331_1235_0, i_10_331_1236_0, i_10_331_1237_0,
    i_10_331_1264_0, i_10_331_1306_0, i_10_331_1307_0, i_10_331_1308_0,
    i_10_331_1309_0, i_10_331_1310_0, i_10_331_1313_0, i_10_331_1577_0,
    i_10_331_1612_0, i_10_331_1684_0, i_10_331_1685_0, i_10_331_1688_0,
    i_10_331_1766_0, i_10_331_1812_0, i_10_331_1813_0, i_10_331_1821_0,
    i_10_331_2180_0, i_10_331_2359_0, i_10_331_2448_0, i_10_331_2467_0,
    i_10_331_2526_0, i_10_331_2606_0, i_10_331_2631_0, i_10_331_2641_0,
    i_10_331_2657_0, i_10_331_2660_0, i_10_331_2701_0, i_10_331_2702_0,
    i_10_331_2711_0, i_10_331_2719_0, i_10_331_2720_0, i_10_331_2728_0,
    i_10_331_2733_0, i_10_331_2818_0, i_10_331_2830_0, i_10_331_2831_0,
    i_10_331_2833_0, i_10_331_2884_0, i_10_331_2885_0, i_10_331_2921_0,
    i_10_331_2923_0, i_10_331_3070_0, i_10_331_3233_0, i_10_331_3268_0,
    i_10_331_3269_0, i_10_331_3280_0, i_10_331_3297_0, i_10_331_3385_0,
    i_10_331_3386_0, i_10_331_3390_0, i_10_331_3391_0, i_10_331_3392_0,
    i_10_331_3406_0, i_10_331_3462_0, i_10_331_3523_0, i_10_331_3585_0,
    i_10_331_3613_0, i_10_331_3614_0, i_10_331_3647_0, i_10_331_3649_0,
    i_10_331_3650_0, i_10_331_3727_0, i_10_331_3732_0, i_10_331_3781_0,
    i_10_331_3782_0, i_10_331_3783_0, i_10_331_3784_0, i_10_331_3787_0,
    i_10_331_3835_0, i_10_331_3837_0, i_10_331_3888_0, i_10_331_3909_0,
    i_10_331_4115_0, i_10_331_4125_0, i_10_331_4169_0, i_10_331_4212_0,
    i_10_331_4285_0, i_10_331_4286_0, i_10_331_4518_0, i_10_331_4565_0;
  output o_10_331_0_0;
  assign o_10_331_0_0 = 0;
endmodule



// Benchmark "kernel_10_332" written by ABC on Sun Jul 19 10:26:48 2020

module kernel_10_332 ( 
    i_10_332_11_0, i_10_332_254_0, i_10_332_320_0, i_10_332_344_0,
    i_10_332_392_0, i_10_332_394_0, i_10_332_433_0, i_10_332_464_0,
    i_10_332_497_0, i_10_332_821_0, i_10_332_824_0, i_10_332_931_0,
    i_10_332_1100_0, i_10_332_1210_0, i_10_332_1220_0, i_10_332_1235_0,
    i_10_332_1238_0, i_10_332_1297_0, i_10_332_1298_0, i_10_332_1300_0,
    i_10_332_1307_0, i_10_332_1433_0, i_10_332_1540_0, i_10_332_1541_0,
    i_10_332_1622_0, i_10_332_1625_0, i_10_332_1684_0, i_10_332_1685_0,
    i_10_332_1688_0, i_10_332_1730_0, i_10_332_1733_0, i_10_332_1805_0,
    i_10_332_1822_0, i_10_332_1825_0, i_10_332_1985_0, i_10_332_1990_0,
    i_10_332_2108_0, i_10_332_2162_0, i_10_332_2201_0, i_10_332_2288_0,
    i_10_332_2345_0, i_10_332_2351_0, i_10_332_2358_0, i_10_332_2359_0,
    i_10_332_2360_0, i_10_332_2408_0, i_10_332_2466_0, i_10_332_2467_0,
    i_10_332_2470_0, i_10_332_2507_0, i_10_332_2530_0, i_10_332_2558_0,
    i_10_332_2561_0, i_10_332_2566_0, i_10_332_2567_0, i_10_332_2570_0,
    i_10_332_2606_0, i_10_332_2632_0, i_10_332_2638_0, i_10_332_2641_0,
    i_10_332_2702_0, i_10_332_2705_0, i_10_332_2710_0, i_10_332_2722_0,
    i_10_332_2729_0, i_10_332_2755_0, i_10_332_2852_0, i_10_332_2963_0,
    i_10_332_3043_0, i_10_332_3070_0, i_10_332_3290_0, i_10_332_3317_0,
    i_10_332_3332_0, i_10_332_3461_0, i_10_332_3503_0, i_10_332_3539_0,
    i_10_332_3545_0, i_10_332_3548_0, i_10_332_3556_0, i_10_332_3557_0,
    i_10_332_3584_0, i_10_332_3586_0, i_10_332_3835_0, i_10_332_3836_0,
    i_10_332_3839_0, i_10_332_3847_0, i_10_332_3848_0, i_10_332_3854_0,
    i_10_332_3908_0, i_10_332_4007_0, i_10_332_4060_0, i_10_332_4123_0,
    i_10_332_4154_0, i_10_332_4169_0, i_10_332_4172_0, i_10_332_4267_0,
    i_10_332_4277_0, i_10_332_4429_0, i_10_332_4433_0, i_10_332_4566_0,
    o_10_332_0_0  );
  input  i_10_332_11_0, i_10_332_254_0, i_10_332_320_0, i_10_332_344_0,
    i_10_332_392_0, i_10_332_394_0, i_10_332_433_0, i_10_332_464_0,
    i_10_332_497_0, i_10_332_821_0, i_10_332_824_0, i_10_332_931_0,
    i_10_332_1100_0, i_10_332_1210_0, i_10_332_1220_0, i_10_332_1235_0,
    i_10_332_1238_0, i_10_332_1297_0, i_10_332_1298_0, i_10_332_1300_0,
    i_10_332_1307_0, i_10_332_1433_0, i_10_332_1540_0, i_10_332_1541_0,
    i_10_332_1622_0, i_10_332_1625_0, i_10_332_1684_0, i_10_332_1685_0,
    i_10_332_1688_0, i_10_332_1730_0, i_10_332_1733_0, i_10_332_1805_0,
    i_10_332_1822_0, i_10_332_1825_0, i_10_332_1985_0, i_10_332_1990_0,
    i_10_332_2108_0, i_10_332_2162_0, i_10_332_2201_0, i_10_332_2288_0,
    i_10_332_2345_0, i_10_332_2351_0, i_10_332_2358_0, i_10_332_2359_0,
    i_10_332_2360_0, i_10_332_2408_0, i_10_332_2466_0, i_10_332_2467_0,
    i_10_332_2470_0, i_10_332_2507_0, i_10_332_2530_0, i_10_332_2558_0,
    i_10_332_2561_0, i_10_332_2566_0, i_10_332_2567_0, i_10_332_2570_0,
    i_10_332_2606_0, i_10_332_2632_0, i_10_332_2638_0, i_10_332_2641_0,
    i_10_332_2702_0, i_10_332_2705_0, i_10_332_2710_0, i_10_332_2722_0,
    i_10_332_2729_0, i_10_332_2755_0, i_10_332_2852_0, i_10_332_2963_0,
    i_10_332_3043_0, i_10_332_3070_0, i_10_332_3290_0, i_10_332_3317_0,
    i_10_332_3332_0, i_10_332_3461_0, i_10_332_3503_0, i_10_332_3539_0,
    i_10_332_3545_0, i_10_332_3548_0, i_10_332_3556_0, i_10_332_3557_0,
    i_10_332_3584_0, i_10_332_3586_0, i_10_332_3835_0, i_10_332_3836_0,
    i_10_332_3839_0, i_10_332_3847_0, i_10_332_3848_0, i_10_332_3854_0,
    i_10_332_3908_0, i_10_332_4007_0, i_10_332_4060_0, i_10_332_4123_0,
    i_10_332_4154_0, i_10_332_4169_0, i_10_332_4172_0, i_10_332_4267_0,
    i_10_332_4277_0, i_10_332_4429_0, i_10_332_4433_0, i_10_332_4566_0;
  output o_10_332_0_0;
  assign o_10_332_0_0 = 0;
endmodule



// Benchmark "kernel_10_333" written by ABC on Sun Jul 19 10:26:48 2020

module kernel_10_333 ( 
    i_10_333_14_0, i_10_333_35_0, i_10_333_80_0, i_10_333_160_0,
    i_10_333_223_0, i_10_333_268_0, i_10_333_269_0, i_10_333_296_0,
    i_10_333_410_0, i_10_333_413_0, i_10_333_439_0, i_10_333_440_0,
    i_10_333_463_0, i_10_333_511_0, i_10_333_512_0, i_10_333_692_0,
    i_10_333_755_0, i_10_333_872_0, i_10_333_1033_0, i_10_333_1034_0,
    i_10_333_1041_0, i_10_333_1042_0, i_10_333_1043_0, i_10_333_1052_0,
    i_10_333_1059_0, i_10_333_1139_0, i_10_333_1157_0, i_10_333_1160_0,
    i_10_333_1175_0, i_10_333_1205_0, i_10_333_1241_0, i_10_333_1249_0,
    i_10_333_1294_0, i_10_333_1303_0, i_10_333_1312_0, i_10_333_1348_0,
    i_10_333_1356_0, i_10_333_1362_0, i_10_333_1366_0, i_10_333_1367_0,
    i_10_333_1439_0, i_10_333_1457_0, i_10_333_1545_0, i_10_333_1546_0,
    i_10_333_1547_0, i_10_333_1582_0, i_10_333_1583_0, i_10_333_1627_0,
    i_10_333_1651_0, i_10_333_1655_0, i_10_333_1690_0, i_10_333_1733_0,
    i_10_333_1735_0, i_10_333_1736_0, i_10_333_1772_0, i_10_333_1781_0,
    i_10_333_1817_0, i_10_333_1850_0, i_10_333_1913_0, i_10_333_1915_0,
    i_10_333_1984_0, i_10_333_1987_0, i_10_333_1988_0, i_10_333_2356_0,
    i_10_333_2453_0, i_10_333_2467_0, i_10_333_2560_0, i_10_333_2609_0,
    i_10_333_2660_0, i_10_333_2702_0, i_10_333_2723_0, i_10_333_2743_0,
    i_10_333_2816_0, i_10_333_2829_0, i_10_333_2830_0, i_10_333_2839_0,
    i_10_333_2851_0, i_10_333_2965_0, i_10_333_2968_0, i_10_333_2969_0,
    i_10_333_2987_0, i_10_333_3049_0, i_10_333_3274_0, i_10_333_3392_0,
    i_10_333_3409_0, i_10_333_3437_0, i_10_333_3508_0, i_10_333_3544_0,
    i_10_333_3614_0, i_10_333_3859_0, i_10_333_3984_0, i_10_333_3985_0,
    i_10_333_4117_0, i_10_333_4118_0, i_10_333_4119_0, i_10_333_4238_0,
    i_10_333_4288_0, i_10_333_4462_0, i_10_333_4570_0, i_10_333_4571_0,
    o_10_333_0_0  );
  input  i_10_333_14_0, i_10_333_35_0, i_10_333_80_0, i_10_333_160_0,
    i_10_333_223_0, i_10_333_268_0, i_10_333_269_0, i_10_333_296_0,
    i_10_333_410_0, i_10_333_413_0, i_10_333_439_0, i_10_333_440_0,
    i_10_333_463_0, i_10_333_511_0, i_10_333_512_0, i_10_333_692_0,
    i_10_333_755_0, i_10_333_872_0, i_10_333_1033_0, i_10_333_1034_0,
    i_10_333_1041_0, i_10_333_1042_0, i_10_333_1043_0, i_10_333_1052_0,
    i_10_333_1059_0, i_10_333_1139_0, i_10_333_1157_0, i_10_333_1160_0,
    i_10_333_1175_0, i_10_333_1205_0, i_10_333_1241_0, i_10_333_1249_0,
    i_10_333_1294_0, i_10_333_1303_0, i_10_333_1312_0, i_10_333_1348_0,
    i_10_333_1356_0, i_10_333_1362_0, i_10_333_1366_0, i_10_333_1367_0,
    i_10_333_1439_0, i_10_333_1457_0, i_10_333_1545_0, i_10_333_1546_0,
    i_10_333_1547_0, i_10_333_1582_0, i_10_333_1583_0, i_10_333_1627_0,
    i_10_333_1651_0, i_10_333_1655_0, i_10_333_1690_0, i_10_333_1733_0,
    i_10_333_1735_0, i_10_333_1736_0, i_10_333_1772_0, i_10_333_1781_0,
    i_10_333_1817_0, i_10_333_1850_0, i_10_333_1913_0, i_10_333_1915_0,
    i_10_333_1984_0, i_10_333_1987_0, i_10_333_1988_0, i_10_333_2356_0,
    i_10_333_2453_0, i_10_333_2467_0, i_10_333_2560_0, i_10_333_2609_0,
    i_10_333_2660_0, i_10_333_2702_0, i_10_333_2723_0, i_10_333_2743_0,
    i_10_333_2816_0, i_10_333_2829_0, i_10_333_2830_0, i_10_333_2839_0,
    i_10_333_2851_0, i_10_333_2965_0, i_10_333_2968_0, i_10_333_2969_0,
    i_10_333_2987_0, i_10_333_3049_0, i_10_333_3274_0, i_10_333_3392_0,
    i_10_333_3409_0, i_10_333_3437_0, i_10_333_3508_0, i_10_333_3544_0,
    i_10_333_3614_0, i_10_333_3859_0, i_10_333_3984_0, i_10_333_3985_0,
    i_10_333_4117_0, i_10_333_4118_0, i_10_333_4119_0, i_10_333_4238_0,
    i_10_333_4288_0, i_10_333_4462_0, i_10_333_4570_0, i_10_333_4571_0;
  output o_10_333_0_0;
  assign o_10_333_0_0 = 0;
endmodule



// Benchmark "kernel_10_334" written by ABC on Sun Jul 19 10:26:49 2020

module kernel_10_334 ( 
    i_10_334_13_0, i_10_334_15_0, i_10_334_16_0, i_10_334_22_0,
    i_10_334_39_0, i_10_334_40_0, i_10_334_121_0, i_10_334_160_0,
    i_10_334_281_0, i_10_334_286_0, i_10_334_433_0, i_10_334_434_0,
    i_10_334_513_0, i_10_334_514_0, i_10_334_595_0, i_10_334_598_0,
    i_10_334_635_0, i_10_334_661_0, i_10_334_691_0, i_10_334_800_0,
    i_10_334_872_0, i_10_334_907_0, i_10_334_1060_0, i_10_334_1159_0,
    i_10_334_1169_0, i_10_334_1175_0, i_10_334_1399_0, i_10_334_1439_0,
    i_10_334_1487_0, i_10_334_1542_0, i_10_334_1545_0, i_10_334_1713_0,
    i_10_334_1850_0, i_10_334_1877_0, i_10_334_1879_0, i_10_334_1880_0,
    i_10_334_2020_0, i_10_334_2023_0, i_10_334_2024_0, i_10_334_2029_0,
    i_10_334_2030_0, i_10_334_2037_0, i_10_334_2112_0, i_10_334_2203_0,
    i_10_334_2204_0, i_10_334_2222_0, i_10_334_2243_0, i_10_334_2245_0,
    i_10_334_2380_0, i_10_334_2410_0, i_10_334_2411_0, i_10_334_2467_0,
    i_10_334_2468_0, i_10_334_2472_0, i_10_334_2598_0, i_10_334_2599_0,
    i_10_334_2608_0, i_10_334_2616_0, i_10_334_2660_0, i_10_334_2663_0,
    i_10_334_2678_0, i_10_334_2707_0, i_10_334_2708_0, i_10_334_2711_0,
    i_10_334_2714_0, i_10_334_2722_0, i_10_334_2733_0, i_10_334_2735_0,
    i_10_334_2789_0, i_10_334_2821_0, i_10_334_2824_0, i_10_334_2884_0,
    i_10_334_2885_0, i_10_334_2987_0, i_10_334_3046_0, i_10_334_3072_0,
    i_10_334_3075_0, i_10_334_3076_0, i_10_334_3077_0, i_10_334_3109_0,
    i_10_334_3163_0, i_10_334_3199_0, i_10_334_3407_0, i_10_334_3469_0,
    i_10_334_3472_0, i_10_334_3473_0, i_10_334_3522_0, i_10_334_3586_0,
    i_10_334_3589_0, i_10_334_3590_0, i_10_334_3622_0, i_10_334_3653_0,
    i_10_334_3683_0, i_10_334_3724_0, i_10_334_3839_0, i_10_334_3909_0,
    i_10_334_3910_0, i_10_334_4121_0, i_10_334_4124_0, i_10_334_4526_0,
    o_10_334_0_0  );
  input  i_10_334_13_0, i_10_334_15_0, i_10_334_16_0, i_10_334_22_0,
    i_10_334_39_0, i_10_334_40_0, i_10_334_121_0, i_10_334_160_0,
    i_10_334_281_0, i_10_334_286_0, i_10_334_433_0, i_10_334_434_0,
    i_10_334_513_0, i_10_334_514_0, i_10_334_595_0, i_10_334_598_0,
    i_10_334_635_0, i_10_334_661_0, i_10_334_691_0, i_10_334_800_0,
    i_10_334_872_0, i_10_334_907_0, i_10_334_1060_0, i_10_334_1159_0,
    i_10_334_1169_0, i_10_334_1175_0, i_10_334_1399_0, i_10_334_1439_0,
    i_10_334_1487_0, i_10_334_1542_0, i_10_334_1545_0, i_10_334_1713_0,
    i_10_334_1850_0, i_10_334_1877_0, i_10_334_1879_0, i_10_334_1880_0,
    i_10_334_2020_0, i_10_334_2023_0, i_10_334_2024_0, i_10_334_2029_0,
    i_10_334_2030_0, i_10_334_2037_0, i_10_334_2112_0, i_10_334_2203_0,
    i_10_334_2204_0, i_10_334_2222_0, i_10_334_2243_0, i_10_334_2245_0,
    i_10_334_2380_0, i_10_334_2410_0, i_10_334_2411_0, i_10_334_2467_0,
    i_10_334_2468_0, i_10_334_2472_0, i_10_334_2598_0, i_10_334_2599_0,
    i_10_334_2608_0, i_10_334_2616_0, i_10_334_2660_0, i_10_334_2663_0,
    i_10_334_2678_0, i_10_334_2707_0, i_10_334_2708_0, i_10_334_2711_0,
    i_10_334_2714_0, i_10_334_2722_0, i_10_334_2733_0, i_10_334_2735_0,
    i_10_334_2789_0, i_10_334_2821_0, i_10_334_2824_0, i_10_334_2884_0,
    i_10_334_2885_0, i_10_334_2987_0, i_10_334_3046_0, i_10_334_3072_0,
    i_10_334_3075_0, i_10_334_3076_0, i_10_334_3077_0, i_10_334_3109_0,
    i_10_334_3163_0, i_10_334_3199_0, i_10_334_3407_0, i_10_334_3469_0,
    i_10_334_3472_0, i_10_334_3473_0, i_10_334_3522_0, i_10_334_3586_0,
    i_10_334_3589_0, i_10_334_3590_0, i_10_334_3622_0, i_10_334_3653_0,
    i_10_334_3683_0, i_10_334_3724_0, i_10_334_3839_0, i_10_334_3909_0,
    i_10_334_3910_0, i_10_334_4121_0, i_10_334_4124_0, i_10_334_4526_0;
  output o_10_334_0_0;
  assign o_10_334_0_0 = 0;
endmodule



// Benchmark "kernel_10_335" written by ABC on Sun Jul 19 10:26:50 2020

module kernel_10_335 ( 
    i_10_335_146_0, i_10_335_175_0, i_10_335_284_0, i_10_335_407_0,
    i_10_335_441_0, i_10_335_442_0, i_10_335_443_0, i_10_335_444_0,
    i_10_335_793_0, i_10_335_794_0, i_10_335_800_0, i_10_335_964_0,
    i_10_335_966_0, i_10_335_1117_0, i_10_335_1205_0, i_10_335_1264_0,
    i_10_335_1307_0, i_10_335_1308_0, i_10_335_1346_0, i_10_335_1575_0,
    i_10_335_1620_0, i_10_335_1636_0, i_10_335_1647_0, i_10_335_1651_0,
    i_10_335_1652_0, i_10_335_1683_0, i_10_335_1684_0, i_10_335_1685_0,
    i_10_335_1820_0, i_10_335_1826_0, i_10_335_1915_0, i_10_335_1947_0,
    i_10_335_2000_0, i_10_335_2158_0, i_10_335_2159_0, i_10_335_2333_0,
    i_10_335_2350_0, i_10_335_2352_0, i_10_335_2454_0, i_10_335_2470_0,
    i_10_335_2514_0, i_10_335_2556_0, i_10_335_2631_0, i_10_335_2632_0,
    i_10_335_2701_0, i_10_335_2711_0, i_10_335_2719_0, i_10_335_2789_0,
    i_10_335_2831_0, i_10_335_2850_0, i_10_335_2884_0, i_10_335_2888_0,
    i_10_335_2920_0, i_10_335_2921_0, i_10_335_2923_0, i_10_335_2924_0,
    i_10_335_2952_0, i_10_335_2979_0, i_10_335_3090_0, i_10_335_3239_0,
    i_10_335_3270_0, i_10_335_3387_0, i_10_335_3388_0, i_10_335_3391_0,
    i_10_335_3406_0, i_10_335_3434_0, i_10_335_3522_0, i_10_335_3523_0,
    i_10_335_3524_0, i_10_335_3525_0, i_10_335_3526_0, i_10_335_3527_0,
    i_10_335_3590_0, i_10_335_3610_0, i_10_335_3611_0, i_10_335_3613_0,
    i_10_335_3614_0, i_10_335_3682_0, i_10_335_3683_0, i_10_335_3704_0,
    i_10_335_3730_0, i_10_335_3783_0, i_10_335_3835_0, i_10_335_3844_0,
    i_10_335_3854_0, i_10_335_3860_0, i_10_335_3995_0, i_10_335_4191_0,
    i_10_335_4192_0, i_10_335_4215_0, i_10_335_4216_0, i_10_335_4218_0,
    i_10_335_4269_0, i_10_335_4290_0, i_10_335_4291_0, i_10_335_4459_0,
    i_10_335_4460_0, i_10_335_4462_0, i_10_335_4560_0, i_10_335_4570_0,
    o_10_335_0_0  );
  input  i_10_335_146_0, i_10_335_175_0, i_10_335_284_0, i_10_335_407_0,
    i_10_335_441_0, i_10_335_442_0, i_10_335_443_0, i_10_335_444_0,
    i_10_335_793_0, i_10_335_794_0, i_10_335_800_0, i_10_335_964_0,
    i_10_335_966_0, i_10_335_1117_0, i_10_335_1205_0, i_10_335_1264_0,
    i_10_335_1307_0, i_10_335_1308_0, i_10_335_1346_0, i_10_335_1575_0,
    i_10_335_1620_0, i_10_335_1636_0, i_10_335_1647_0, i_10_335_1651_0,
    i_10_335_1652_0, i_10_335_1683_0, i_10_335_1684_0, i_10_335_1685_0,
    i_10_335_1820_0, i_10_335_1826_0, i_10_335_1915_0, i_10_335_1947_0,
    i_10_335_2000_0, i_10_335_2158_0, i_10_335_2159_0, i_10_335_2333_0,
    i_10_335_2350_0, i_10_335_2352_0, i_10_335_2454_0, i_10_335_2470_0,
    i_10_335_2514_0, i_10_335_2556_0, i_10_335_2631_0, i_10_335_2632_0,
    i_10_335_2701_0, i_10_335_2711_0, i_10_335_2719_0, i_10_335_2789_0,
    i_10_335_2831_0, i_10_335_2850_0, i_10_335_2884_0, i_10_335_2888_0,
    i_10_335_2920_0, i_10_335_2921_0, i_10_335_2923_0, i_10_335_2924_0,
    i_10_335_2952_0, i_10_335_2979_0, i_10_335_3090_0, i_10_335_3239_0,
    i_10_335_3270_0, i_10_335_3387_0, i_10_335_3388_0, i_10_335_3391_0,
    i_10_335_3406_0, i_10_335_3434_0, i_10_335_3522_0, i_10_335_3523_0,
    i_10_335_3524_0, i_10_335_3525_0, i_10_335_3526_0, i_10_335_3527_0,
    i_10_335_3590_0, i_10_335_3610_0, i_10_335_3611_0, i_10_335_3613_0,
    i_10_335_3614_0, i_10_335_3682_0, i_10_335_3683_0, i_10_335_3704_0,
    i_10_335_3730_0, i_10_335_3783_0, i_10_335_3835_0, i_10_335_3844_0,
    i_10_335_3854_0, i_10_335_3860_0, i_10_335_3995_0, i_10_335_4191_0,
    i_10_335_4192_0, i_10_335_4215_0, i_10_335_4216_0, i_10_335_4218_0,
    i_10_335_4269_0, i_10_335_4290_0, i_10_335_4291_0, i_10_335_4459_0,
    i_10_335_4460_0, i_10_335_4462_0, i_10_335_4560_0, i_10_335_4570_0;
  output o_10_335_0_0;
  assign o_10_335_0_0 = 0;
endmodule



// Benchmark "kernel_10_336" written by ABC on Sun Jul 19 10:26:52 2020

module kernel_10_336 ( 
    i_10_336_70_0, i_10_336_71_0, i_10_336_174_0, i_10_336_175_0,
    i_10_336_278_0, i_10_336_286_0, i_10_336_328_0, i_10_336_329_0,
    i_10_336_442_0, i_10_336_445_0, i_10_336_446_0, i_10_336_448_0,
    i_10_336_449_0, i_10_336_466_0, i_10_336_505_0, i_10_336_623_0,
    i_10_336_700_0, i_10_336_794_0, i_10_336_958_0, i_10_336_960_0,
    i_10_336_961_0, i_10_336_1031_0, i_10_336_1043_0, i_10_336_1233_0,
    i_10_336_1239_0, i_10_336_1308_0, i_10_336_1312_0, i_10_336_1313_0,
    i_10_336_1347_0, i_10_336_1348_0, i_10_336_1349_0, i_10_336_1547_0,
    i_10_336_1556_0, i_10_336_1653_0, i_10_336_1684_0, i_10_336_1717_0,
    i_10_336_1718_0, i_10_336_1768_0, i_10_336_1822_0, i_10_336_1823_0,
    i_10_336_1824_0, i_10_336_1825_0, i_10_336_1877_0, i_10_336_1991_0,
    i_10_336_2021_0, i_10_336_2166_0, i_10_336_2167_0, i_10_336_2198_0,
    i_10_336_2200_0, i_10_336_2363_0, i_10_336_2382_0, i_10_336_2449_0,
    i_10_336_2450_0, i_10_336_2452_0, i_10_336_2460_0, i_10_336_2461_0,
    i_10_336_2631_0, i_10_336_2634_0, i_10_336_2661_0, i_10_336_2663_0,
    i_10_336_2703_0, i_10_336_2704_0, i_10_336_2716_0, i_10_336_2717_0,
    i_10_336_2722_0, i_10_336_2723_0, i_10_336_2733_0, i_10_336_2734_0,
    i_10_336_2825_0, i_10_336_2829_0, i_10_336_2887_0, i_10_336_2923_0,
    i_10_336_2924_0, i_10_336_3046_0, i_10_336_3047_0, i_10_336_3076_0,
    i_10_336_3077_0, i_10_336_3151_0, i_10_336_3153_0, i_10_336_3284_0,
    i_10_336_3388_0, i_10_336_3389_0, i_10_336_3390_0, i_10_336_3391_0,
    i_10_336_3392_0, i_10_336_3434_0, i_10_336_3472_0, i_10_336_3616_0,
    i_10_336_3617_0, i_10_336_3650_0, i_10_336_3653_0, i_10_336_3775_0,
    i_10_336_3786_0, i_10_336_3835_0, i_10_336_3841_0, i_10_336_3851_0,
    i_10_336_3856_0, i_10_336_4117_0, i_10_336_4287_0, i_10_336_4571_0,
    o_10_336_0_0  );
  input  i_10_336_70_0, i_10_336_71_0, i_10_336_174_0, i_10_336_175_0,
    i_10_336_278_0, i_10_336_286_0, i_10_336_328_0, i_10_336_329_0,
    i_10_336_442_0, i_10_336_445_0, i_10_336_446_0, i_10_336_448_0,
    i_10_336_449_0, i_10_336_466_0, i_10_336_505_0, i_10_336_623_0,
    i_10_336_700_0, i_10_336_794_0, i_10_336_958_0, i_10_336_960_0,
    i_10_336_961_0, i_10_336_1031_0, i_10_336_1043_0, i_10_336_1233_0,
    i_10_336_1239_0, i_10_336_1308_0, i_10_336_1312_0, i_10_336_1313_0,
    i_10_336_1347_0, i_10_336_1348_0, i_10_336_1349_0, i_10_336_1547_0,
    i_10_336_1556_0, i_10_336_1653_0, i_10_336_1684_0, i_10_336_1717_0,
    i_10_336_1718_0, i_10_336_1768_0, i_10_336_1822_0, i_10_336_1823_0,
    i_10_336_1824_0, i_10_336_1825_0, i_10_336_1877_0, i_10_336_1991_0,
    i_10_336_2021_0, i_10_336_2166_0, i_10_336_2167_0, i_10_336_2198_0,
    i_10_336_2200_0, i_10_336_2363_0, i_10_336_2382_0, i_10_336_2449_0,
    i_10_336_2450_0, i_10_336_2452_0, i_10_336_2460_0, i_10_336_2461_0,
    i_10_336_2631_0, i_10_336_2634_0, i_10_336_2661_0, i_10_336_2663_0,
    i_10_336_2703_0, i_10_336_2704_0, i_10_336_2716_0, i_10_336_2717_0,
    i_10_336_2722_0, i_10_336_2723_0, i_10_336_2733_0, i_10_336_2734_0,
    i_10_336_2825_0, i_10_336_2829_0, i_10_336_2887_0, i_10_336_2923_0,
    i_10_336_2924_0, i_10_336_3046_0, i_10_336_3047_0, i_10_336_3076_0,
    i_10_336_3077_0, i_10_336_3151_0, i_10_336_3153_0, i_10_336_3284_0,
    i_10_336_3388_0, i_10_336_3389_0, i_10_336_3390_0, i_10_336_3391_0,
    i_10_336_3392_0, i_10_336_3434_0, i_10_336_3472_0, i_10_336_3616_0,
    i_10_336_3617_0, i_10_336_3650_0, i_10_336_3653_0, i_10_336_3775_0,
    i_10_336_3786_0, i_10_336_3835_0, i_10_336_3841_0, i_10_336_3851_0,
    i_10_336_3856_0, i_10_336_4117_0, i_10_336_4287_0, i_10_336_4571_0;
  output o_10_336_0_0;
  assign o_10_336_0_0 = ~((~i_10_336_3077_0 & ((i_10_336_466_0 & ((~i_10_336_960_0 & ~i_10_336_1349_0 & i_10_336_1825_0 & ~i_10_336_2198_0 & ~i_10_336_2716_0 & ~i_10_336_3047_0) | (i_10_336_1308_0 & ~i_10_336_2460_0 & ~i_10_336_3076_0 & ~i_10_336_3388_0 & ~i_10_336_3390_0 & ~i_10_336_3851_0))) | (~i_10_336_1031_0 & ~i_10_336_1347_0 & ~i_10_336_2198_0 & ~i_10_336_2631_0 & ((~i_10_336_329_0 & ~i_10_336_958_0 & ~i_10_336_961_0 & ~i_10_336_1822_0 & ~i_10_336_1991_0 & ~i_10_336_2021_0 & ~i_10_336_2460_0 & ~i_10_336_3434_0 & ~i_10_336_3616_0) | (~i_10_336_1239_0 & ~i_10_336_1556_0 & ~i_10_336_1877_0 & ~i_10_336_2663_0 & ~i_10_336_3650_0 & i_10_336_3856_0 & ~i_10_336_4117_0))) | (~i_10_336_329_0 & ((i_10_336_286_0 & ~i_10_336_1877_0 & ~i_10_336_2461_0 & ~i_10_336_2717_0 & ~i_10_336_3390_0 & ~i_10_336_3472_0) | (i_10_336_449_0 & ~i_10_336_1547_0 & ~i_10_336_3851_0))) | (~i_10_336_1308_0 & ((i_10_336_2450_0 & ~i_10_336_2452_0 & ~i_10_336_2722_0 & ~i_10_336_3391_0 & ~i_10_336_3786_0) | (i_10_336_1684_0 & ~i_10_336_1825_0 & i_10_336_2198_0 & ~i_10_336_2734_0 & ~i_10_336_3650_0 & ~i_10_336_4117_0))) | (~i_10_336_1349_0 & i_10_336_1825_0 & i_10_336_2663_0) | (~i_10_336_1547_0 & ~i_10_336_1768_0 & ~i_10_336_1823_0 & ~i_10_336_3390_0 & i_10_336_3616_0 & ~i_10_336_3617_0))) | (i_10_336_1233_0 & (i_10_336_446_0 | (~i_10_336_2200_0 & ~i_10_336_2452_0 & ~i_10_336_2723_0 & ~i_10_336_3835_0 & i_10_336_3856_0))) | (i_10_336_446_0 & (i_10_336_3835_0 | (i_10_336_448_0 & ~i_10_336_1547_0))) | (~i_10_336_1308_0 & ((~i_10_336_958_0 & i_10_336_1031_0 & ~i_10_336_2200_0 & i_10_336_2449_0 & ~i_10_336_3392_0) | (~i_10_336_1031_0 & ~i_10_336_2452_0 & ~i_10_336_2722_0 & ~i_10_336_3388_0 & i_10_336_3835_0 & ~i_10_336_4117_0))) | (i_10_336_1312_0 & ((~i_10_336_329_0 & ~i_10_336_958_0 & ~i_10_336_1239_0 & ~i_10_336_2452_0 & ~i_10_336_2634_0 & ~i_10_336_3389_0) | (~i_10_336_328_0 & ~i_10_336_1547_0 & ~i_10_336_2198_0 & ~i_10_336_3390_0 & ~i_10_336_3841_0))) | (~i_10_336_3653_0 & ((~i_10_336_329_0 & ((i_10_336_794_0 & ~i_10_336_1031_0 & ~i_10_336_1233_0 & ~i_10_336_2829_0 & ~i_10_336_3616_0) | (~i_10_336_448_0 & ~i_10_336_960_0 & ~i_10_336_961_0 & ~i_10_336_1348_0 & ~i_10_336_1768_0 & ~i_10_336_2198_0 & ~i_10_336_2460_0 & ~i_10_336_3047_0 & i_10_336_3388_0 & ~i_10_336_3434_0 & ~i_10_336_3786_0))) | (i_10_336_174_0 & ~i_10_336_2461_0 & ~i_10_336_2717_0 & ~i_10_336_3392_0))) | (~i_10_336_2452_0 & ((~i_10_336_1031_0 & ((~i_10_336_2716_0 & ~i_10_336_2722_0 & ~i_10_336_3392_0 & ~i_10_336_3434_0 & ~i_10_336_3650_0 & ~i_10_336_4117_0) | (~i_10_336_328_0 & ~i_10_336_794_0 & ~i_10_336_958_0 & ~i_10_336_1768_0 & ~i_10_336_1825_0 & ~i_10_336_2021_0 & ~i_10_336_2198_0 & ~i_10_336_3391_0 & ~i_10_336_4287_0))) | (~i_10_336_1547_0 & i_10_336_3046_0 & ~i_10_336_3388_0))) | (~i_10_336_2200_0 & ((~i_10_336_328_0 & ((~i_10_336_958_0 & ~i_10_336_1312_0 & ~i_10_336_1313_0 & ~i_10_336_1347_0 & ~i_10_336_1556_0 & ~i_10_336_2198_0 & i_10_336_2631_0) | (~i_10_336_961_0 & ~i_10_336_1349_0 & ~i_10_336_1547_0 & ~i_10_336_1768_0 & ~i_10_336_2461_0 & ~i_10_336_2634_0 & ~i_10_336_2829_0 & ~i_10_336_2887_0 & ~i_10_336_3650_0 & ~i_10_336_3835_0))) | (~i_10_336_958_0 & ~i_10_336_1824_0 & ~i_10_336_2021_0 & ~i_10_336_2198_0 & ~i_10_336_2363_0 & ~i_10_336_2461_0 & ~i_10_336_2634_0 & ~i_10_336_2661_0 & ~i_10_336_2704_0 & ~i_10_336_2717_0) | (i_10_336_1822_0 & i_10_336_2923_0) | (~i_10_336_960_0 & ~i_10_336_1348_0 & ~i_10_336_1877_0 & i_10_336_4571_0))) | (~i_10_336_1877_0 & ((~i_10_336_960_0 & ~i_10_336_3851_0 & ((~i_10_336_466_0 & i_10_336_2734_0 & ~i_10_336_3388_0 & ~i_10_336_3390_0) | (~i_10_336_961_0 & ~i_10_336_1556_0 & ~i_10_336_2363_0 & ~i_10_336_2722_0 & ~i_10_336_3392_0 & ~i_10_336_3786_0 & ~i_10_336_3835_0 & i_10_336_3841_0))) | (i_10_336_174_0 & i_10_336_175_0 & ~i_10_336_442_0 & ~i_10_336_3472_0))) | (i_10_336_174_0 & ((i_10_336_1239_0 & ~i_10_336_1768_0) | (i_10_336_1825_0 & ~i_10_336_3786_0))) | (~i_10_336_961_0 & ~i_10_336_3389_0 & ((~i_10_336_1556_0 & ~i_10_336_1653_0 & ~i_10_336_2450_0 & i_10_336_2733_0 & ~i_10_336_2825_0) | (~i_10_336_958_0 & ~i_10_336_1348_0 & i_10_336_1825_0 & ~i_10_336_3284_0 & ~i_10_336_3617_0))) | (~i_10_336_1348_0 & ((~i_10_336_700_0 & ~i_10_336_1653_0 & ~i_10_336_2021_0 & ~i_10_336_2461_0 & i_10_336_2661_0) | (~i_10_336_1768_0 & i_10_336_2450_0 & ~i_10_336_3392_0 & i_10_336_3617_0))) | (~i_10_336_3392_0 & ((i_10_336_445_0 & ~i_10_336_2363_0 & ~i_10_336_2722_0) | (~i_10_336_958_0 & i_10_336_1653_0 & ~i_10_336_2825_0 & ~i_10_336_3076_0 & i_10_336_3617_0))) | (~i_10_336_958_0 & ~i_10_336_2363_0 & ((i_10_336_1823_0 & ~i_10_336_2198_0 & ~i_10_336_2717_0 & ~i_10_336_2829_0) | (~i_10_336_1556_0 & ~i_10_336_3616_0 & ~i_10_336_3650_0 & i_10_336_4287_0))) | (i_10_336_1991_0 & ~i_10_336_2631_0 & i_10_336_4287_0) | (i_10_336_442_0 & i_10_336_3046_0));
endmodule



// Benchmark "kernel_10_337" written by ABC on Sun Jul 19 10:26:53 2020

module kernel_10_337 ( 
    i_10_337_276_0, i_10_337_282_0, i_10_337_320_0, i_10_337_321_0,
    i_10_337_328_0, i_10_337_442_0, i_10_337_443_0, i_10_337_447_0,
    i_10_337_448_0, i_10_337_462_0, i_10_337_514_0, i_10_337_516_0,
    i_10_337_519_0, i_10_337_561_0, i_10_337_718_0, i_10_337_795_0,
    i_10_337_798_0, i_10_337_969_0, i_10_337_970_0, i_10_337_993_0,
    i_10_337_1164_0, i_10_337_1234_0, i_10_337_1438_0, i_10_337_1445_0,
    i_10_337_1492_0, i_10_337_1578_0, i_10_337_1581_0, i_10_337_1641_0,
    i_10_337_1652_0, i_10_337_1653_0, i_10_337_1807_0, i_10_337_1815_0,
    i_10_337_1822_0, i_10_337_1946_0, i_10_337_2030_0, i_10_337_2182_0,
    i_10_337_2251_0, i_10_337_2308_0, i_10_337_2310_0, i_10_337_2311_0,
    i_10_337_2349_0, i_10_337_2350_0, i_10_337_2351_0, i_10_337_2352_0,
    i_10_337_2353_0, i_10_337_2356_0, i_10_337_2383_0, i_10_337_2410_0,
    i_10_337_2450_0, i_10_337_2454_0, i_10_337_2544_0, i_10_337_2634_0,
    i_10_337_2676_0, i_10_337_2717_0, i_10_337_2724_0, i_10_337_2727_0,
    i_10_337_2730_0, i_10_337_2743_0, i_10_337_2784_0, i_10_337_2785_0,
    i_10_337_2955_0, i_10_337_2982_0, i_10_337_2985_0, i_10_337_2986_0,
    i_10_337_3040_0, i_10_337_3091_0, i_10_337_3102_0, i_10_337_3103_0,
    i_10_337_3120_0, i_10_337_3156_0, i_10_337_3198_0, i_10_337_3232_0,
    i_10_337_3283_0, i_10_337_3298_0, i_10_337_3468_0, i_10_337_3493_0,
    i_10_337_3494_0, i_10_337_3496_0, i_10_337_3525_0, i_10_337_3588_0,
    i_10_337_3611_0, i_10_337_3649_0, i_10_337_3653_0, i_10_337_3786_0,
    i_10_337_3805_0, i_10_337_3857_0, i_10_337_3874_0, i_10_337_3896_0,
    i_10_337_3949_0, i_10_337_3979_0, i_10_337_4113_0, i_10_337_4117_0,
    i_10_337_4119_0, i_10_337_4146_0, i_10_337_4266_0, i_10_337_4270_0,
    i_10_337_4271_0, i_10_337_4281_0, i_10_337_4285_0, i_10_337_4288_0,
    o_10_337_0_0  );
  input  i_10_337_276_0, i_10_337_282_0, i_10_337_320_0, i_10_337_321_0,
    i_10_337_328_0, i_10_337_442_0, i_10_337_443_0, i_10_337_447_0,
    i_10_337_448_0, i_10_337_462_0, i_10_337_514_0, i_10_337_516_0,
    i_10_337_519_0, i_10_337_561_0, i_10_337_718_0, i_10_337_795_0,
    i_10_337_798_0, i_10_337_969_0, i_10_337_970_0, i_10_337_993_0,
    i_10_337_1164_0, i_10_337_1234_0, i_10_337_1438_0, i_10_337_1445_0,
    i_10_337_1492_0, i_10_337_1578_0, i_10_337_1581_0, i_10_337_1641_0,
    i_10_337_1652_0, i_10_337_1653_0, i_10_337_1807_0, i_10_337_1815_0,
    i_10_337_1822_0, i_10_337_1946_0, i_10_337_2030_0, i_10_337_2182_0,
    i_10_337_2251_0, i_10_337_2308_0, i_10_337_2310_0, i_10_337_2311_0,
    i_10_337_2349_0, i_10_337_2350_0, i_10_337_2351_0, i_10_337_2352_0,
    i_10_337_2353_0, i_10_337_2356_0, i_10_337_2383_0, i_10_337_2410_0,
    i_10_337_2450_0, i_10_337_2454_0, i_10_337_2544_0, i_10_337_2634_0,
    i_10_337_2676_0, i_10_337_2717_0, i_10_337_2724_0, i_10_337_2727_0,
    i_10_337_2730_0, i_10_337_2743_0, i_10_337_2784_0, i_10_337_2785_0,
    i_10_337_2955_0, i_10_337_2982_0, i_10_337_2985_0, i_10_337_2986_0,
    i_10_337_3040_0, i_10_337_3091_0, i_10_337_3102_0, i_10_337_3103_0,
    i_10_337_3120_0, i_10_337_3156_0, i_10_337_3198_0, i_10_337_3232_0,
    i_10_337_3283_0, i_10_337_3298_0, i_10_337_3468_0, i_10_337_3493_0,
    i_10_337_3494_0, i_10_337_3496_0, i_10_337_3525_0, i_10_337_3588_0,
    i_10_337_3611_0, i_10_337_3649_0, i_10_337_3653_0, i_10_337_3786_0,
    i_10_337_3805_0, i_10_337_3857_0, i_10_337_3874_0, i_10_337_3896_0,
    i_10_337_3949_0, i_10_337_3979_0, i_10_337_4113_0, i_10_337_4117_0,
    i_10_337_4119_0, i_10_337_4146_0, i_10_337_4266_0, i_10_337_4270_0,
    i_10_337_4271_0, i_10_337_4281_0, i_10_337_4285_0, i_10_337_4288_0;
  output o_10_337_0_0;
  assign o_10_337_0_0 = ~((~i_10_337_718_0 & ((~i_10_337_519_0 & ((~i_10_337_993_0 & ~i_10_337_2383_0 & ~i_10_337_2784_0) | (~i_10_337_4271_0 & i_10_337_4288_0))) | (~i_10_337_321_0 & ~i_10_337_795_0 & ~i_10_337_1445_0 & ~i_10_337_2982_0 & ~i_10_337_4266_0) | (~i_10_337_2349_0 & ~i_10_337_3232_0 & ~i_10_337_3979_0 & ~i_10_337_4270_0) | (~i_10_337_969_0 & ~i_10_337_1652_0 & ~i_10_337_2454_0 & ~i_10_337_3496_0 & ~i_10_337_3525_0 & ~i_10_337_4271_0 & ~i_10_337_4285_0 & ~i_10_337_4288_0))) | (~i_10_337_3949_0 & ((~i_10_337_1164_0 & ~i_10_337_2311_0 & ((~i_10_337_1492_0 & ~i_10_337_1822_0 & ~i_10_337_2676_0 & ~i_10_337_2784_0 & ~i_10_337_3493_0 & ~i_10_337_3979_0) | (~i_10_337_516_0 & ~i_10_337_2730_0 & ~i_10_337_2982_0 & ~i_10_337_3232_0 & ~i_10_337_3496_0 & ~i_10_337_4281_0))) | (~i_10_337_448_0 & ~i_10_337_514_0 & ~i_10_337_2450_0 & ~i_10_337_2454_0 & ~i_10_337_3198_0 & ~i_10_337_3494_0 & ~i_10_337_3653_0))) | (~i_10_337_2351_0 & ((~i_10_337_447_0 & ~i_10_337_798_0 & ~i_10_337_969_0 & ~i_10_337_1581_0 & ~i_10_337_3493_0) | (~i_10_337_795_0 & i_10_337_1652_0 & ~i_10_337_3496_0 & ~i_10_337_4119_0))) | (~i_10_337_969_0 & ((i_10_337_1822_0 & ~i_10_337_2676_0 & ~i_10_337_2982_0 & ~i_10_337_2985_0 & ~i_10_337_3496_0 & ~i_10_337_3857_0 & ~i_10_337_4281_0) | (~i_10_337_1815_0 & ~i_10_337_2410_0 & ~i_10_337_2450_0 & ~i_10_337_2724_0 & ~i_10_337_2986_0 & ~i_10_337_3493_0 & ~i_10_337_3494_0 & ~i_10_337_4285_0))) | (~i_10_337_2982_0 & ((~i_10_337_2350_0 & ~i_10_337_2717_0 & ~i_10_337_3232_0 & ~i_10_337_3468_0) | (~i_10_337_282_0 & ~i_10_337_1492_0 & ~i_10_337_2986_0 & i_10_337_3232_0 & ~i_10_337_3493_0))) | (i_10_337_3611_0 & (~i_10_337_2352_0 | (~i_10_337_2986_0 & ~i_10_337_3857_0))) | (i_10_337_328_0 & ~i_10_337_442_0 & ~i_10_337_2308_0 & ~i_10_337_2349_0 & i_10_337_2353_0 & i_10_337_2986_0 & i_10_337_3649_0 & ~i_10_337_3653_0) | (~i_10_337_1653_0 & ~i_10_337_1822_0 & ~i_10_337_2030_0 & ~i_10_337_3494_0 & ~i_10_337_4119_0 & ~i_10_337_4266_0) | (i_10_337_2410_0 & ~i_10_337_2676_0 & ~i_10_337_4270_0) | (i_10_337_3896_0 & ~i_10_337_4271_0));
endmodule



// Benchmark "kernel_10_338" written by ABC on Sun Jul 19 10:26:54 2020

module kernel_10_338 ( 
    i_10_338_171_0, i_10_338_172_0, i_10_338_177_0, i_10_338_220_0,
    i_10_338_223_0, i_10_338_271_0, i_10_338_272_0, i_10_338_274_0,
    i_10_338_282_0, i_10_338_318_0, i_10_338_427_0, i_10_338_430_0,
    i_10_338_435_0, i_10_338_438_0, i_10_338_442_0, i_10_338_446_0,
    i_10_338_463_0, i_10_338_711_0, i_10_338_712_0, i_10_338_1030_0,
    i_10_338_1037_0, i_10_338_1238_0, i_10_338_1305_0, i_10_338_1311_0,
    i_10_338_1343_0, i_10_338_1346_0, i_10_338_1548_0, i_10_338_1549_0,
    i_10_338_1551_0, i_10_338_1552_0, i_10_338_1651_0, i_10_338_1652_0,
    i_10_338_1654_0, i_10_338_1655_0, i_10_338_1683_0, i_10_338_1764_0,
    i_10_338_1765_0, i_10_338_1819_0, i_10_338_1822_0, i_10_338_1824_0,
    i_10_338_1910_0, i_10_338_2197_0, i_10_338_2358_0, i_10_338_2381_0,
    i_10_338_2382_0, i_10_338_2383_0, i_10_338_2410_0, i_10_338_2635_0,
    i_10_338_2636_0, i_10_338_2662_0, i_10_338_2704_0, i_10_338_2707_0,
    i_10_338_2710_0, i_10_338_2712_0, i_10_338_2728_0, i_10_338_2731_0,
    i_10_338_2732_0, i_10_338_2783_0, i_10_338_2821_0, i_10_338_2832_0,
    i_10_338_2880_0, i_10_338_2883_0, i_10_338_2884_0, i_10_338_2885_0,
    i_10_338_2886_0, i_10_338_2887_0, i_10_338_2888_0, i_10_338_3040_0,
    i_10_338_3070_0, i_10_338_3151_0, i_10_338_3198_0, i_10_338_3277_0,
    i_10_338_3326_0, i_10_338_3384_0, i_10_338_3385_0, i_10_338_3386_0,
    i_10_338_3387_0, i_10_338_3405_0, i_10_338_3406_0, i_10_338_3409_0,
    i_10_338_3410_0, i_10_338_3588_0, i_10_338_3614_0, i_10_338_3684_0,
    i_10_338_3842_0, i_10_338_3856_0, i_10_338_3857_0, i_10_338_3859_0,
    i_10_338_3860_0, i_10_338_3891_0, i_10_338_3983_0, i_10_338_3994_0,
    i_10_338_3995_0, i_10_338_4118_0, i_10_338_4126_0, i_10_338_4287_0,
    i_10_338_4288_0, i_10_338_4290_0, i_10_338_4292_0, i_10_338_4594_0,
    o_10_338_0_0  );
  input  i_10_338_171_0, i_10_338_172_0, i_10_338_177_0, i_10_338_220_0,
    i_10_338_223_0, i_10_338_271_0, i_10_338_272_0, i_10_338_274_0,
    i_10_338_282_0, i_10_338_318_0, i_10_338_427_0, i_10_338_430_0,
    i_10_338_435_0, i_10_338_438_0, i_10_338_442_0, i_10_338_446_0,
    i_10_338_463_0, i_10_338_711_0, i_10_338_712_0, i_10_338_1030_0,
    i_10_338_1037_0, i_10_338_1238_0, i_10_338_1305_0, i_10_338_1311_0,
    i_10_338_1343_0, i_10_338_1346_0, i_10_338_1548_0, i_10_338_1549_0,
    i_10_338_1551_0, i_10_338_1552_0, i_10_338_1651_0, i_10_338_1652_0,
    i_10_338_1654_0, i_10_338_1655_0, i_10_338_1683_0, i_10_338_1764_0,
    i_10_338_1765_0, i_10_338_1819_0, i_10_338_1822_0, i_10_338_1824_0,
    i_10_338_1910_0, i_10_338_2197_0, i_10_338_2358_0, i_10_338_2381_0,
    i_10_338_2382_0, i_10_338_2383_0, i_10_338_2410_0, i_10_338_2635_0,
    i_10_338_2636_0, i_10_338_2662_0, i_10_338_2704_0, i_10_338_2707_0,
    i_10_338_2710_0, i_10_338_2712_0, i_10_338_2728_0, i_10_338_2731_0,
    i_10_338_2732_0, i_10_338_2783_0, i_10_338_2821_0, i_10_338_2832_0,
    i_10_338_2880_0, i_10_338_2883_0, i_10_338_2884_0, i_10_338_2885_0,
    i_10_338_2886_0, i_10_338_2887_0, i_10_338_2888_0, i_10_338_3040_0,
    i_10_338_3070_0, i_10_338_3151_0, i_10_338_3198_0, i_10_338_3277_0,
    i_10_338_3326_0, i_10_338_3384_0, i_10_338_3385_0, i_10_338_3386_0,
    i_10_338_3387_0, i_10_338_3405_0, i_10_338_3406_0, i_10_338_3409_0,
    i_10_338_3410_0, i_10_338_3588_0, i_10_338_3614_0, i_10_338_3684_0,
    i_10_338_3842_0, i_10_338_3856_0, i_10_338_3857_0, i_10_338_3859_0,
    i_10_338_3860_0, i_10_338_3891_0, i_10_338_3983_0, i_10_338_3994_0,
    i_10_338_3995_0, i_10_338_4118_0, i_10_338_4126_0, i_10_338_4287_0,
    i_10_338_4288_0, i_10_338_4290_0, i_10_338_4292_0, i_10_338_4594_0;
  output o_10_338_0_0;
  assign o_10_338_0_0 = ~((i_10_338_177_0 & ((~i_10_338_2884_0 & ~i_10_338_4290_0) | (~i_10_338_282_0 & ~i_10_338_1305_0 & i_10_338_1822_0 & ~i_10_338_2886_0 & ~i_10_338_3387_0 & ~i_10_338_3983_0 & ~i_10_338_4292_0))) | (~i_10_338_282_0 & ((i_10_338_1824_0 & i_10_338_2636_0 & ~i_10_338_2704_0 & ~i_10_338_3387_0 & i_10_338_4118_0) | (~i_10_338_1549_0 & i_10_338_1652_0 & i_10_338_2635_0 & ~i_10_338_3995_0 & ~i_10_338_4290_0))) | (~i_10_338_427_0 & ((~i_10_338_463_0 & i_10_338_1683_0 & ~i_10_338_2886_0 & i_10_338_4287_0) | (~i_10_338_430_0 & i_10_338_435_0 & ~i_10_338_4288_0 & ~i_10_338_4290_0))) | (~i_10_338_446_0 & ((~i_10_338_430_0 & ((~i_10_338_2885_0 & ~i_10_338_2886_0 & ~i_10_338_2888_0 & ~i_10_338_3588_0 & ~i_10_338_4287_0) | (~i_10_338_1551_0 & ~i_10_338_2382_0 & ~i_10_338_2884_0 & ~i_10_338_3406_0 & ~i_10_338_4290_0))) | (~i_10_338_1551_0 & ~i_10_338_1552_0 & i_10_338_1822_0 & i_10_338_2707_0 & ~i_10_338_2887_0 & ~i_10_338_3277_0))) | (~i_10_338_438_0 & ((~i_10_338_1552_0 & ~i_10_338_1819_0 & ~i_10_338_1824_0 & ~i_10_338_2635_0 & ~i_10_338_2636_0 & ~i_10_338_2704_0 & ~i_10_338_2887_0 & ~i_10_338_2888_0 & ~i_10_338_3384_0 & ~i_10_338_3385_0 & ~i_10_338_3387_0) | (i_10_338_1651_0 & ~i_10_338_3405_0 & ~i_10_338_3842_0))) | (i_10_338_446_0 & ((i_10_338_463_0 & ~i_10_338_1822_0 & i_10_338_3588_0) | (~i_10_338_2884_0 & ~i_10_338_2887_0 & ~i_10_338_3385_0 & ~i_10_338_3588_0 & ~i_10_338_3860_0))) | (~i_10_338_1037_0 & ((~i_10_338_1548_0 & i_10_338_1819_0 & ~i_10_338_2888_0 & ~i_10_338_3384_0) | (~i_10_338_318_0 & ~i_10_338_2636_0 & ~i_10_338_2731_0 & ~i_10_338_2884_0 & ~i_10_338_2886_0 & ~i_10_338_4288_0))) | (~i_10_338_2884_0 & ((~i_10_338_1549_0 & ((~i_10_338_1683_0 & ~i_10_338_1764_0 & ~i_10_338_1824_0 & ~i_10_338_2636_0 & ~i_10_338_2883_0 & ~i_10_338_3856_0 & ~i_10_338_3891_0) | (~i_10_338_435_0 & i_10_338_1822_0 & i_10_338_4288_0 & ~i_10_338_4290_0))) | (~i_10_338_1551_0 & i_10_338_2635_0 & ~i_10_338_2887_0 & i_10_338_3406_0 & i_10_338_3856_0) | (~i_10_338_2662_0 & ~i_10_338_3385_0 & i_10_338_3588_0 & ~i_10_338_4287_0 & i_10_338_4292_0))) | (~i_10_338_1551_0 & ((~i_10_338_1343_0 & ~i_10_338_2887_0 & i_10_338_3983_0) | (i_10_338_2731_0 & ~i_10_338_2886_0 & ~i_10_338_4292_0))) | (i_10_338_463_0 & ((~i_10_338_2883_0 & ~i_10_338_2888_0 & ((i_10_338_427_0 & ~i_10_338_1305_0 & i_10_338_4290_0) | (~i_10_338_2885_0 & ~i_10_338_3995_0 & ~i_10_338_4290_0))) | (~i_10_338_177_0 & ~i_10_338_2731_0 & ~i_10_338_2886_0 & ~i_10_338_2887_0 & ~i_10_338_3387_0 & ~i_10_338_3406_0))) | (~i_10_338_2887_0 & (i_10_338_4126_0 | (~i_10_338_1552_0 & i_10_338_2832_0 & ~i_10_338_4118_0))) | (i_10_338_318_0 & ~i_10_338_1238_0 & i_10_338_1311_0 & ~i_10_338_2382_0 & ~i_10_338_2383_0 & ~i_10_338_3405_0 & ~i_10_338_3856_0) | (i_10_338_282_0 & ~i_10_338_1824_0 & ~i_10_338_2712_0 & ~i_10_338_3857_0 & i_10_338_4118_0));
endmodule



// Benchmark "kernel_10_339" written by ABC on Sun Jul 19 10:26:55 2020

module kernel_10_339 ( 
    i_10_339_255_0, i_10_339_277_0, i_10_339_280_0, i_10_339_281_0,
    i_10_339_315_0, i_10_339_318_0, i_10_339_322_0, i_10_339_387_0,
    i_10_339_393_0, i_10_339_406_0, i_10_339_408_0, i_10_339_441_0,
    i_10_339_442_0, i_10_339_462_0, i_10_339_465_0, i_10_339_519_0,
    i_10_339_747_0, i_10_339_795_0, i_10_339_798_0, i_10_339_963_0,
    i_10_339_1026_0, i_10_339_1029_0, i_10_339_1241_0, i_10_339_1308_0,
    i_10_339_1362_0, i_10_339_1431_0, i_10_339_1434_0, i_10_339_1435_0,
    i_10_339_1444_0, i_10_339_1539_0, i_10_339_1540_0, i_10_339_1542_0,
    i_10_339_1545_0, i_10_339_1578_0, i_10_339_1626_0, i_10_339_1648_0,
    i_10_339_1683_0, i_10_339_1684_0, i_10_339_1686_0, i_10_339_1689_0,
    i_10_339_1719_0, i_10_339_1806_0, i_10_339_1819_0, i_10_339_1821_0,
    i_10_339_1823_0, i_10_339_1826_0, i_10_339_2028_0, i_10_339_2179_0,
    i_10_339_2180_0, i_10_339_2349_0, i_10_339_2350_0, i_10_339_2407_0,
    i_10_339_2451_0, i_10_339_2469_0, i_10_339_2628_0, i_10_339_2631_0,
    i_10_339_2632_0, i_10_339_2636_0, i_10_339_2656_0, i_10_339_2659_0,
    i_10_339_2660_0, i_10_339_2661_0, i_10_339_2728_0, i_10_339_2731_0,
    i_10_339_2733_0, i_10_339_2785_0, i_10_339_2829_0, i_10_339_2880_0,
    i_10_339_2921_0, i_10_339_2967_0, i_10_339_3034_0, i_10_339_3069_0,
    i_10_339_3072_0, i_10_339_3151_0, i_10_339_3153_0, i_10_339_3154_0,
    i_10_339_3270_0, i_10_339_3271_0, i_10_339_3280_0, i_10_339_3318_0,
    i_10_339_3325_0, i_10_339_3336_0, i_10_339_3468_0, i_10_339_3523_0,
    i_10_339_3543_0, i_10_339_3615_0, i_10_339_3648_0, i_10_339_3835_0,
    i_10_339_3837_0, i_10_339_3847_0, i_10_339_3909_0, i_10_339_3910_0,
    i_10_339_3993_0, i_10_339_3994_0, i_10_339_4118_0, i_10_339_4170_0,
    i_10_339_4270_0, i_10_339_4272_0, i_10_339_4275_0, i_10_339_4566_0,
    o_10_339_0_0  );
  input  i_10_339_255_0, i_10_339_277_0, i_10_339_280_0, i_10_339_281_0,
    i_10_339_315_0, i_10_339_318_0, i_10_339_322_0, i_10_339_387_0,
    i_10_339_393_0, i_10_339_406_0, i_10_339_408_0, i_10_339_441_0,
    i_10_339_442_0, i_10_339_462_0, i_10_339_465_0, i_10_339_519_0,
    i_10_339_747_0, i_10_339_795_0, i_10_339_798_0, i_10_339_963_0,
    i_10_339_1026_0, i_10_339_1029_0, i_10_339_1241_0, i_10_339_1308_0,
    i_10_339_1362_0, i_10_339_1431_0, i_10_339_1434_0, i_10_339_1435_0,
    i_10_339_1444_0, i_10_339_1539_0, i_10_339_1540_0, i_10_339_1542_0,
    i_10_339_1545_0, i_10_339_1578_0, i_10_339_1626_0, i_10_339_1648_0,
    i_10_339_1683_0, i_10_339_1684_0, i_10_339_1686_0, i_10_339_1689_0,
    i_10_339_1719_0, i_10_339_1806_0, i_10_339_1819_0, i_10_339_1821_0,
    i_10_339_1823_0, i_10_339_1826_0, i_10_339_2028_0, i_10_339_2179_0,
    i_10_339_2180_0, i_10_339_2349_0, i_10_339_2350_0, i_10_339_2407_0,
    i_10_339_2451_0, i_10_339_2469_0, i_10_339_2628_0, i_10_339_2631_0,
    i_10_339_2632_0, i_10_339_2636_0, i_10_339_2656_0, i_10_339_2659_0,
    i_10_339_2660_0, i_10_339_2661_0, i_10_339_2728_0, i_10_339_2731_0,
    i_10_339_2733_0, i_10_339_2785_0, i_10_339_2829_0, i_10_339_2880_0,
    i_10_339_2921_0, i_10_339_2967_0, i_10_339_3034_0, i_10_339_3069_0,
    i_10_339_3072_0, i_10_339_3151_0, i_10_339_3153_0, i_10_339_3154_0,
    i_10_339_3270_0, i_10_339_3271_0, i_10_339_3280_0, i_10_339_3318_0,
    i_10_339_3325_0, i_10_339_3336_0, i_10_339_3468_0, i_10_339_3523_0,
    i_10_339_3543_0, i_10_339_3615_0, i_10_339_3648_0, i_10_339_3835_0,
    i_10_339_3837_0, i_10_339_3847_0, i_10_339_3909_0, i_10_339_3910_0,
    i_10_339_3993_0, i_10_339_3994_0, i_10_339_4118_0, i_10_339_4170_0,
    i_10_339_4270_0, i_10_339_4272_0, i_10_339_4275_0, i_10_339_4566_0;
  output o_10_339_0_0;
  assign o_10_339_0_0 = ~((~i_10_339_1431_0 & ((~i_10_339_255_0 & ((~i_10_339_1434_0 & ~i_10_339_1539_0 & ~i_10_339_1542_0 & ~i_10_339_1545_0) | (~i_10_339_393_0 & ~i_10_339_406_0 & ~i_10_339_747_0 & ~i_10_339_1626_0 & ~i_10_339_1823_0 & ~i_10_339_2451_0 & ~i_10_339_2469_0 & ~i_10_339_2880_0 & ~i_10_339_3271_0))) | (~i_10_339_1241_0 & ~i_10_339_1539_0 & ~i_10_339_1545_0 & ~i_10_339_3069_0 & ~i_10_339_3468_0) | (~i_10_339_1540_0 & ~i_10_339_1686_0 & ~i_10_339_2733_0 & i_10_339_4118_0))) | (~i_10_339_1026_0 & ~i_10_339_1626_0 & ~i_10_339_2636_0 & ((~i_10_339_519_0 & ~i_10_339_2469_0 & ~i_10_339_2733_0 & ~i_10_339_2785_0 & ~i_10_339_2880_0 & ~i_10_339_2921_0 & ~i_10_339_3072_0 & ~i_10_339_3543_0 & ~i_10_339_3615_0) | (~i_10_339_322_0 & ~i_10_339_798_0 & ~i_10_339_1683_0 & ~i_10_339_3648_0 & ~i_10_339_3909_0 & ~i_10_339_4118_0))) | (~i_10_339_1542_0 & ((~i_10_339_1029_0 & ~i_10_339_2659_0 & ((~i_10_339_747_0 & ~i_10_339_1578_0 & ~i_10_339_2180_0 & ~i_10_339_2733_0 & ~i_10_339_2880_0 & ~i_10_339_3543_0) | (i_10_339_1026_0 & ~i_10_339_2179_0 & i_10_339_2728_0 & ~i_10_339_3280_0 & ~i_10_339_3468_0 & ~i_10_339_4566_0))) | (~i_10_339_1683_0 & i_10_339_2659_0 & ~i_10_339_3069_0))) | (~i_10_339_3072_0 & ((~i_10_339_442_0 & ~i_10_339_1578_0 & ~i_10_339_3280_0 & i_10_339_3835_0 & ~i_10_339_3847_0) | (~i_10_339_1689_0 & ~i_10_339_2349_0 & ~i_10_339_3069_0 & ~i_10_339_3468_0 & ~i_10_339_3543_0 & ~i_10_339_3994_0 & ~i_10_339_4275_0))) | (i_10_339_2636_0 & i_10_339_2921_0));
endmodule



// Benchmark "kernel_10_340" written by ABC on Sun Jul 19 10:26:56 2020

module kernel_10_340 ( 
    i_10_340_34_0, i_10_340_61_0, i_10_340_259_0, i_10_340_273_0,
    i_10_340_282_0, i_10_340_283_0, i_10_340_284_0, i_10_340_301_0,
    i_10_340_444_0, i_10_340_637_0, i_10_340_642_0, i_10_340_717_0,
    i_10_340_718_0, i_10_340_755_0, i_10_340_958_0, i_10_340_962_0,
    i_10_340_1030_0, i_10_340_1034_0, i_10_340_1243_0, i_10_340_1248_0,
    i_10_340_1249_0, i_10_340_1250_0, i_10_340_1265_0, i_10_340_1309_0,
    i_10_340_1385_0, i_10_340_1448_0, i_10_340_1546_0, i_10_340_1547_0,
    i_10_340_1582_0, i_10_340_1619_0, i_10_340_1689_0, i_10_340_1690_0,
    i_10_340_1691_0, i_10_340_1760_0, i_10_340_1824_0, i_10_340_1825_0,
    i_10_340_1961_0, i_10_340_2167_0, i_10_340_2168_0, i_10_340_2185_0,
    i_10_340_2186_0, i_10_340_2199_0, i_10_340_2203_0, i_10_340_2204_0,
    i_10_340_2273_0, i_10_340_2338_0, i_10_340_2352_0, i_10_340_2355_0,
    i_10_340_2356_0, i_10_340_2357_0, i_10_340_2472_0, i_10_340_2536_0,
    i_10_340_2609_0, i_10_340_2632_0, i_10_340_2662_0, i_10_340_2694_0,
    i_10_340_2955_0, i_10_340_3038_0, i_10_340_3075_0, i_10_340_3076_0,
    i_10_340_3177_0, i_10_340_3199_0, i_10_340_3202_0, i_10_340_3239_0,
    i_10_340_3268_0, i_10_340_3274_0, i_10_340_3275_0, i_10_340_3306_0,
    i_10_340_3337_0, i_10_340_3389_0, i_10_340_3390_0, i_10_340_3434_0,
    i_10_340_3468_0, i_10_340_3551_0, i_10_340_3613_0, i_10_340_3626_0,
    i_10_340_3650_0, i_10_340_3734_0, i_10_340_3786_0, i_10_340_3795_0,
    i_10_340_3810_0, i_10_340_3814_0, i_10_340_3815_0, i_10_340_3846_0,
    i_10_340_3847_0, i_10_340_3848_0, i_10_340_3850_0, i_10_340_3851_0,
    i_10_340_3856_0, i_10_340_3877_0, i_10_340_4000_0, i_10_340_4013_0,
    i_10_340_4116_0, i_10_340_4119_0, i_10_340_4120_0, i_10_340_4174_0,
    i_10_340_4220_0, i_10_340_4264_0, i_10_340_4292_0, i_10_340_4585_0,
    o_10_340_0_0  );
  input  i_10_340_34_0, i_10_340_61_0, i_10_340_259_0, i_10_340_273_0,
    i_10_340_282_0, i_10_340_283_0, i_10_340_284_0, i_10_340_301_0,
    i_10_340_444_0, i_10_340_637_0, i_10_340_642_0, i_10_340_717_0,
    i_10_340_718_0, i_10_340_755_0, i_10_340_958_0, i_10_340_962_0,
    i_10_340_1030_0, i_10_340_1034_0, i_10_340_1243_0, i_10_340_1248_0,
    i_10_340_1249_0, i_10_340_1250_0, i_10_340_1265_0, i_10_340_1309_0,
    i_10_340_1385_0, i_10_340_1448_0, i_10_340_1546_0, i_10_340_1547_0,
    i_10_340_1582_0, i_10_340_1619_0, i_10_340_1689_0, i_10_340_1690_0,
    i_10_340_1691_0, i_10_340_1760_0, i_10_340_1824_0, i_10_340_1825_0,
    i_10_340_1961_0, i_10_340_2167_0, i_10_340_2168_0, i_10_340_2185_0,
    i_10_340_2186_0, i_10_340_2199_0, i_10_340_2203_0, i_10_340_2204_0,
    i_10_340_2273_0, i_10_340_2338_0, i_10_340_2352_0, i_10_340_2355_0,
    i_10_340_2356_0, i_10_340_2357_0, i_10_340_2472_0, i_10_340_2536_0,
    i_10_340_2609_0, i_10_340_2632_0, i_10_340_2662_0, i_10_340_2694_0,
    i_10_340_2955_0, i_10_340_3038_0, i_10_340_3075_0, i_10_340_3076_0,
    i_10_340_3177_0, i_10_340_3199_0, i_10_340_3202_0, i_10_340_3239_0,
    i_10_340_3268_0, i_10_340_3274_0, i_10_340_3275_0, i_10_340_3306_0,
    i_10_340_3337_0, i_10_340_3389_0, i_10_340_3390_0, i_10_340_3434_0,
    i_10_340_3468_0, i_10_340_3551_0, i_10_340_3613_0, i_10_340_3626_0,
    i_10_340_3650_0, i_10_340_3734_0, i_10_340_3786_0, i_10_340_3795_0,
    i_10_340_3810_0, i_10_340_3814_0, i_10_340_3815_0, i_10_340_3846_0,
    i_10_340_3847_0, i_10_340_3848_0, i_10_340_3850_0, i_10_340_3851_0,
    i_10_340_3856_0, i_10_340_3877_0, i_10_340_4000_0, i_10_340_4013_0,
    i_10_340_4116_0, i_10_340_4119_0, i_10_340_4120_0, i_10_340_4174_0,
    i_10_340_4220_0, i_10_340_4264_0, i_10_340_4292_0, i_10_340_4585_0;
  output o_10_340_0_0;
  assign o_10_340_0_0 = 0;
endmodule



// Benchmark "kernel_10_341" written by ABC on Sun Jul 19 10:26:57 2020

module kernel_10_341 ( 
    i_10_341_30_0, i_10_341_34_0, i_10_341_175_0, i_10_341_282_0,
    i_10_341_283_0, i_10_341_319_0, i_10_341_390_0, i_10_341_410_0,
    i_10_341_412_0, i_10_341_445_0, i_10_341_466_0, i_10_341_542_0,
    i_10_341_714_0, i_10_341_798_0, i_10_341_799_0, i_10_341_954_0,
    i_10_341_958_0, i_10_341_968_0, i_10_341_1026_0, i_10_341_1027_0,
    i_10_341_1028_0, i_10_341_1029_0, i_10_341_1233_0, i_10_341_1234_0,
    i_10_341_1264_0, i_10_341_1265_0, i_10_341_1305_0, i_10_341_1306_0,
    i_10_341_1313_0, i_10_341_1542_0, i_10_341_1596_0, i_10_341_1653_0,
    i_10_341_1655_0, i_10_341_1691_0, i_10_341_1824_0, i_10_341_1825_0,
    i_10_341_2006_0, i_10_341_2016_0, i_10_341_2081_0, i_10_341_2185_0,
    i_10_341_2198_0, i_10_341_2307_0, i_10_341_2310_0, i_10_341_2350_0,
    i_10_341_2352_0, i_10_341_2353_0, i_10_341_2361_0, i_10_341_2471_0,
    i_10_341_2629_0, i_10_341_2635_0, i_10_341_2657_0, i_10_341_2677_0,
    i_10_341_2713_0, i_10_341_2714_0, i_10_341_2718_0, i_10_341_2726_0,
    i_10_341_2739_0, i_10_341_2824_0, i_10_341_2829_0, i_10_341_2922_0,
    i_10_341_2952_0, i_10_341_3033_0, i_10_341_3034_0, i_10_341_3076_0,
    i_10_341_3231_0, i_10_341_3232_0, i_10_341_3270_0, i_10_341_3331_0,
    i_10_341_3333_0, i_10_341_3429_0, i_10_341_3546_0, i_10_341_3616_0,
    i_10_341_3617_0, i_10_341_3626_0, i_10_341_3649_0, i_10_341_3650_0,
    i_10_341_3689_0, i_10_341_3718_0, i_10_341_3780_0, i_10_341_3783_0,
    i_10_341_3784_0, i_10_341_3786_0, i_10_341_3787_0, i_10_341_3788_0,
    i_10_341_3808_0, i_10_341_3810_0, i_10_341_3811_0, i_10_341_3843_0,
    i_10_341_3844_0, i_10_341_3846_0, i_10_341_3854_0, i_10_341_4115_0,
    i_10_341_4116_0, i_10_341_4119_0, i_10_341_4121_0, i_10_341_4122_0,
    i_10_341_4123_0, i_10_341_4126_0, i_10_341_4167_0, i_10_341_4275_0,
    o_10_341_0_0  );
  input  i_10_341_30_0, i_10_341_34_0, i_10_341_175_0, i_10_341_282_0,
    i_10_341_283_0, i_10_341_319_0, i_10_341_390_0, i_10_341_410_0,
    i_10_341_412_0, i_10_341_445_0, i_10_341_466_0, i_10_341_542_0,
    i_10_341_714_0, i_10_341_798_0, i_10_341_799_0, i_10_341_954_0,
    i_10_341_958_0, i_10_341_968_0, i_10_341_1026_0, i_10_341_1027_0,
    i_10_341_1028_0, i_10_341_1029_0, i_10_341_1233_0, i_10_341_1234_0,
    i_10_341_1264_0, i_10_341_1265_0, i_10_341_1305_0, i_10_341_1306_0,
    i_10_341_1313_0, i_10_341_1542_0, i_10_341_1596_0, i_10_341_1653_0,
    i_10_341_1655_0, i_10_341_1691_0, i_10_341_1824_0, i_10_341_1825_0,
    i_10_341_2006_0, i_10_341_2016_0, i_10_341_2081_0, i_10_341_2185_0,
    i_10_341_2198_0, i_10_341_2307_0, i_10_341_2310_0, i_10_341_2350_0,
    i_10_341_2352_0, i_10_341_2353_0, i_10_341_2361_0, i_10_341_2471_0,
    i_10_341_2629_0, i_10_341_2635_0, i_10_341_2657_0, i_10_341_2677_0,
    i_10_341_2713_0, i_10_341_2714_0, i_10_341_2718_0, i_10_341_2726_0,
    i_10_341_2739_0, i_10_341_2824_0, i_10_341_2829_0, i_10_341_2922_0,
    i_10_341_2952_0, i_10_341_3033_0, i_10_341_3034_0, i_10_341_3076_0,
    i_10_341_3231_0, i_10_341_3232_0, i_10_341_3270_0, i_10_341_3331_0,
    i_10_341_3333_0, i_10_341_3429_0, i_10_341_3546_0, i_10_341_3616_0,
    i_10_341_3617_0, i_10_341_3626_0, i_10_341_3649_0, i_10_341_3650_0,
    i_10_341_3689_0, i_10_341_3718_0, i_10_341_3780_0, i_10_341_3783_0,
    i_10_341_3784_0, i_10_341_3786_0, i_10_341_3787_0, i_10_341_3788_0,
    i_10_341_3808_0, i_10_341_3810_0, i_10_341_3811_0, i_10_341_3843_0,
    i_10_341_3844_0, i_10_341_3846_0, i_10_341_3854_0, i_10_341_4115_0,
    i_10_341_4116_0, i_10_341_4119_0, i_10_341_4121_0, i_10_341_4122_0,
    i_10_341_4123_0, i_10_341_4126_0, i_10_341_4167_0, i_10_341_4275_0;
  output o_10_341_0_0;
  assign o_10_341_0_0 = 0;
endmodule



// Benchmark "kernel_10_342" written by ABC on Sun Jul 19 10:26:58 2020

module kernel_10_342 ( 
    i_10_342_48_0, i_10_342_51_0, i_10_342_52_0, i_10_342_219_0,
    i_10_342_221_0, i_10_342_223_0, i_10_342_267_0, i_10_342_284_0,
    i_10_342_286_0, i_10_342_295_0, i_10_342_461_0, i_10_342_462_0,
    i_10_342_463_0, i_10_342_699_0, i_10_342_796_0, i_10_342_852_0,
    i_10_342_897_0, i_10_342_898_0, i_10_342_1037_0, i_10_342_1050_0,
    i_10_342_1113_0, i_10_342_1195_0, i_10_342_1250_0, i_10_342_1346_0,
    i_10_342_1435_0, i_10_342_1575_0, i_10_342_1616_0, i_10_342_1623_0,
    i_10_342_1685_0, i_10_342_1688_0, i_10_342_1771_0, i_10_342_1821_0,
    i_10_342_1824_0, i_10_342_2211_0, i_10_342_2263_0, i_10_342_2357_0,
    i_10_342_2365_0, i_10_342_2438_0, i_10_342_2454_0, i_10_342_2455_0,
    i_10_342_2465_0, i_10_342_2474_0, i_10_342_2514_0, i_10_342_2515_0,
    i_10_342_2568_0, i_10_342_2631_0, i_10_342_2632_0, i_10_342_2641_0,
    i_10_342_2652_0, i_10_342_2653_0, i_10_342_2705_0, i_10_342_2712_0,
    i_10_342_2715_0, i_10_342_2723_0, i_10_342_2828_0, i_10_342_2832_0,
    i_10_342_2885_0, i_10_342_2888_0, i_10_342_2923_0, i_10_342_2924_0,
    i_10_342_2982_0, i_10_342_2986_0, i_10_342_3093_0, i_10_342_3094_0,
    i_10_342_3270_0, i_10_342_3273_0, i_10_342_3275_0, i_10_342_3276_0,
    i_10_342_3277_0, i_10_342_3390_0, i_10_342_3391_0, i_10_342_3392_0,
    i_10_342_3407_0, i_10_342_3561_0, i_10_342_3612_0, i_10_342_3613_0,
    i_10_342_3617_0, i_10_342_3732_0, i_10_342_3839_0, i_10_342_3841_0,
    i_10_342_3847_0, i_10_342_3855_0, i_10_342_3856_0, i_10_342_3858_0,
    i_10_342_3892_0, i_10_342_3893_0, i_10_342_3894_0, i_10_342_3982_0,
    i_10_342_3983_0, i_10_342_3985_0, i_10_342_3992_0, i_10_342_4027_0,
    i_10_342_4029_0, i_10_342_4031_0, i_10_342_4120_0, i_10_342_4154_0,
    i_10_342_4156_0, i_10_342_4218_0, i_10_342_4219_0, i_10_342_4506_0,
    o_10_342_0_0  );
  input  i_10_342_48_0, i_10_342_51_0, i_10_342_52_0, i_10_342_219_0,
    i_10_342_221_0, i_10_342_223_0, i_10_342_267_0, i_10_342_284_0,
    i_10_342_286_0, i_10_342_295_0, i_10_342_461_0, i_10_342_462_0,
    i_10_342_463_0, i_10_342_699_0, i_10_342_796_0, i_10_342_852_0,
    i_10_342_897_0, i_10_342_898_0, i_10_342_1037_0, i_10_342_1050_0,
    i_10_342_1113_0, i_10_342_1195_0, i_10_342_1250_0, i_10_342_1346_0,
    i_10_342_1435_0, i_10_342_1575_0, i_10_342_1616_0, i_10_342_1623_0,
    i_10_342_1685_0, i_10_342_1688_0, i_10_342_1771_0, i_10_342_1821_0,
    i_10_342_1824_0, i_10_342_2211_0, i_10_342_2263_0, i_10_342_2357_0,
    i_10_342_2365_0, i_10_342_2438_0, i_10_342_2454_0, i_10_342_2455_0,
    i_10_342_2465_0, i_10_342_2474_0, i_10_342_2514_0, i_10_342_2515_0,
    i_10_342_2568_0, i_10_342_2631_0, i_10_342_2632_0, i_10_342_2641_0,
    i_10_342_2652_0, i_10_342_2653_0, i_10_342_2705_0, i_10_342_2712_0,
    i_10_342_2715_0, i_10_342_2723_0, i_10_342_2828_0, i_10_342_2832_0,
    i_10_342_2885_0, i_10_342_2888_0, i_10_342_2923_0, i_10_342_2924_0,
    i_10_342_2982_0, i_10_342_2986_0, i_10_342_3093_0, i_10_342_3094_0,
    i_10_342_3270_0, i_10_342_3273_0, i_10_342_3275_0, i_10_342_3276_0,
    i_10_342_3277_0, i_10_342_3390_0, i_10_342_3391_0, i_10_342_3392_0,
    i_10_342_3407_0, i_10_342_3561_0, i_10_342_3612_0, i_10_342_3613_0,
    i_10_342_3617_0, i_10_342_3732_0, i_10_342_3839_0, i_10_342_3841_0,
    i_10_342_3847_0, i_10_342_3855_0, i_10_342_3856_0, i_10_342_3858_0,
    i_10_342_3892_0, i_10_342_3893_0, i_10_342_3894_0, i_10_342_3982_0,
    i_10_342_3983_0, i_10_342_3985_0, i_10_342_3992_0, i_10_342_4027_0,
    i_10_342_4029_0, i_10_342_4031_0, i_10_342_4120_0, i_10_342_4154_0,
    i_10_342_4156_0, i_10_342_4218_0, i_10_342_4219_0, i_10_342_4506_0;
  output o_10_342_0_0;
  assign o_10_342_0_0 = 0;
endmodule



// Benchmark "kernel_10_343" written by ABC on Sun Jul 19 10:26:59 2020

module kernel_10_343 ( 
    i_10_343_37_0, i_10_343_63_0, i_10_343_91_0, i_10_343_221_0,
    i_10_343_261_0, i_10_343_292_0, i_10_343_327_0, i_10_343_413_0,
    i_10_343_440_0, i_10_343_464_0, i_10_343_585_0, i_10_343_589_0,
    i_10_343_632_0, i_10_343_697_0, i_10_343_725_0, i_10_343_733_0,
    i_10_343_792_0, i_10_343_793_0, i_10_343_832_0, i_10_343_833_0,
    i_10_343_877_0, i_10_343_891_0, i_10_343_892_0, i_10_343_920_0,
    i_10_343_931_0, i_10_343_964_0, i_10_343_967_0, i_10_343_968_0,
    i_10_343_970_0, i_10_343_1008_0, i_10_343_1029_0, i_10_343_1031_0,
    i_10_343_1117_0, i_10_343_1163_0, i_10_343_1216_0, i_10_343_1270_0,
    i_10_343_1288_0, i_10_343_1291_0, i_10_343_1310_0, i_10_343_1311_0,
    i_10_343_1363_0, i_10_343_1687_0, i_10_343_1766_0, i_10_343_1801_0,
    i_10_343_1810_0, i_10_343_1819_0, i_10_343_1823_0, i_10_343_1980_0,
    i_10_343_1999_0, i_10_343_2002_0, i_10_343_2224_0, i_10_343_2308_0,
    i_10_343_2351_0, i_10_343_2407_0, i_10_343_2449_0, i_10_343_2489_0,
    i_10_343_2517_0, i_10_343_2518_0, i_10_343_2539_0, i_10_343_2565_0,
    i_10_343_2678_0, i_10_343_2710_0, i_10_343_2721_0, i_10_343_2722_0,
    i_10_343_2821_0, i_10_343_2822_0, i_10_343_2980_0, i_10_343_2984_0,
    i_10_343_3010_0, i_10_343_3013_0, i_10_343_3274_0, i_10_343_3298_0,
    i_10_343_3331_0, i_10_343_3332_0, i_10_343_3349_0, i_10_343_3470_0,
    i_10_343_3539_0, i_10_343_3587_0, i_10_343_3610_0, i_10_343_3622_0,
    i_10_343_3623_0, i_10_343_3651_0, i_10_343_3685_0, i_10_343_3820_0,
    i_10_343_3970_0, i_10_343_3992_0, i_10_343_3997_0, i_10_343_4009_0,
    i_10_343_4060_0, i_10_343_4061_0, i_10_343_4118_0, i_10_343_4226_0,
    i_10_343_4387_0, i_10_343_4429_0, i_10_343_4522_0, i_10_343_4525_0,
    i_10_343_4571_0, i_10_343_4582_0, i_10_343_4583_0, i_10_343_4588_0,
    o_10_343_0_0  );
  input  i_10_343_37_0, i_10_343_63_0, i_10_343_91_0, i_10_343_221_0,
    i_10_343_261_0, i_10_343_292_0, i_10_343_327_0, i_10_343_413_0,
    i_10_343_440_0, i_10_343_464_0, i_10_343_585_0, i_10_343_589_0,
    i_10_343_632_0, i_10_343_697_0, i_10_343_725_0, i_10_343_733_0,
    i_10_343_792_0, i_10_343_793_0, i_10_343_832_0, i_10_343_833_0,
    i_10_343_877_0, i_10_343_891_0, i_10_343_892_0, i_10_343_920_0,
    i_10_343_931_0, i_10_343_964_0, i_10_343_967_0, i_10_343_968_0,
    i_10_343_970_0, i_10_343_1008_0, i_10_343_1029_0, i_10_343_1031_0,
    i_10_343_1117_0, i_10_343_1163_0, i_10_343_1216_0, i_10_343_1270_0,
    i_10_343_1288_0, i_10_343_1291_0, i_10_343_1310_0, i_10_343_1311_0,
    i_10_343_1363_0, i_10_343_1687_0, i_10_343_1766_0, i_10_343_1801_0,
    i_10_343_1810_0, i_10_343_1819_0, i_10_343_1823_0, i_10_343_1980_0,
    i_10_343_1999_0, i_10_343_2002_0, i_10_343_2224_0, i_10_343_2308_0,
    i_10_343_2351_0, i_10_343_2407_0, i_10_343_2449_0, i_10_343_2489_0,
    i_10_343_2517_0, i_10_343_2518_0, i_10_343_2539_0, i_10_343_2565_0,
    i_10_343_2678_0, i_10_343_2710_0, i_10_343_2721_0, i_10_343_2722_0,
    i_10_343_2821_0, i_10_343_2822_0, i_10_343_2980_0, i_10_343_2984_0,
    i_10_343_3010_0, i_10_343_3013_0, i_10_343_3274_0, i_10_343_3298_0,
    i_10_343_3331_0, i_10_343_3332_0, i_10_343_3349_0, i_10_343_3470_0,
    i_10_343_3539_0, i_10_343_3587_0, i_10_343_3610_0, i_10_343_3622_0,
    i_10_343_3623_0, i_10_343_3651_0, i_10_343_3685_0, i_10_343_3820_0,
    i_10_343_3970_0, i_10_343_3992_0, i_10_343_3997_0, i_10_343_4009_0,
    i_10_343_4060_0, i_10_343_4061_0, i_10_343_4118_0, i_10_343_4226_0,
    i_10_343_4387_0, i_10_343_4429_0, i_10_343_4522_0, i_10_343_4525_0,
    i_10_343_4571_0, i_10_343_4582_0, i_10_343_4583_0, i_10_343_4588_0;
  output o_10_343_0_0;
  assign o_10_343_0_0 = 0;
endmodule



// Benchmark "kernel_10_344" written by ABC on Sun Jul 19 10:26:59 2020

module kernel_10_344 ( 
    i_10_344_86_0, i_10_344_144_0, i_10_344_149_0, i_10_344_172_0,
    i_10_344_173_0, i_10_344_184_0, i_10_344_185_0, i_10_344_253_0,
    i_10_344_254_0, i_10_344_311_0, i_10_344_374_0, i_10_344_423_0,
    i_10_344_424_0, i_10_344_428_0, i_10_344_465_0, i_10_344_560_0,
    i_10_344_692_0, i_10_344_734_0, i_10_344_779_0, i_10_344_792_0,
    i_10_344_900_0, i_10_344_901_0, i_10_344_923_0, i_10_344_963_0,
    i_10_344_997_0, i_10_344_1003_0, i_10_344_1030_0, i_10_344_1053_0,
    i_10_344_1123_0, i_10_344_1162_0, i_10_344_1205_0, i_10_344_1328_0,
    i_10_344_1486_0, i_10_344_1654_0, i_10_344_1683_0, i_10_344_1685_0,
    i_10_344_1768_0, i_10_344_1792_0, i_10_344_1801_0, i_10_344_1854_0,
    i_10_344_1864_0, i_10_344_1905_0, i_10_344_1942_0, i_10_344_1949_0,
    i_10_344_2002_0, i_10_344_2090_0, i_10_344_2255_0, i_10_344_2356_0,
    i_10_344_2383_0, i_10_344_2450_0, i_10_344_2453_0, i_10_344_2461_0,
    i_10_344_2479_0, i_10_344_2513_0, i_10_344_2531_0, i_10_344_2578_0,
    i_10_344_2663_0, i_10_344_2709_0, i_10_344_2713_0, i_10_344_2722_0,
    i_10_344_2727_0, i_10_344_2740_0, i_10_344_2783_0, i_10_344_2804_0,
    i_10_344_2823_0, i_10_344_2827_0, i_10_344_2880_0, i_10_344_2887_0,
    i_10_344_2998_0, i_10_344_3007_0, i_10_344_3119_0, i_10_344_3197_0,
    i_10_344_3231_0, i_10_344_3290_0, i_10_344_3386_0, i_10_344_3451_0,
    i_10_344_3452_0, i_10_344_3466_0, i_10_344_3493_0, i_10_344_3501_0,
    i_10_344_3552_0, i_10_344_3589_0, i_10_344_3590_0, i_10_344_3616_0,
    i_10_344_3702_0, i_10_344_3788_0, i_10_344_3838_0, i_10_344_3858_0,
    i_10_344_3880_0, i_10_344_3883_0, i_10_344_3943_0, i_10_344_4055_0,
    i_10_344_4114_0, i_10_344_4115_0, i_10_344_4213_0, i_10_344_4217_0,
    i_10_344_4220_0, i_10_344_4281_0, i_10_344_4340_0, i_10_344_4451_0,
    o_10_344_0_0  );
  input  i_10_344_86_0, i_10_344_144_0, i_10_344_149_0, i_10_344_172_0,
    i_10_344_173_0, i_10_344_184_0, i_10_344_185_0, i_10_344_253_0,
    i_10_344_254_0, i_10_344_311_0, i_10_344_374_0, i_10_344_423_0,
    i_10_344_424_0, i_10_344_428_0, i_10_344_465_0, i_10_344_560_0,
    i_10_344_692_0, i_10_344_734_0, i_10_344_779_0, i_10_344_792_0,
    i_10_344_900_0, i_10_344_901_0, i_10_344_923_0, i_10_344_963_0,
    i_10_344_997_0, i_10_344_1003_0, i_10_344_1030_0, i_10_344_1053_0,
    i_10_344_1123_0, i_10_344_1162_0, i_10_344_1205_0, i_10_344_1328_0,
    i_10_344_1486_0, i_10_344_1654_0, i_10_344_1683_0, i_10_344_1685_0,
    i_10_344_1768_0, i_10_344_1792_0, i_10_344_1801_0, i_10_344_1854_0,
    i_10_344_1864_0, i_10_344_1905_0, i_10_344_1942_0, i_10_344_1949_0,
    i_10_344_2002_0, i_10_344_2090_0, i_10_344_2255_0, i_10_344_2356_0,
    i_10_344_2383_0, i_10_344_2450_0, i_10_344_2453_0, i_10_344_2461_0,
    i_10_344_2479_0, i_10_344_2513_0, i_10_344_2531_0, i_10_344_2578_0,
    i_10_344_2663_0, i_10_344_2709_0, i_10_344_2713_0, i_10_344_2722_0,
    i_10_344_2727_0, i_10_344_2740_0, i_10_344_2783_0, i_10_344_2804_0,
    i_10_344_2823_0, i_10_344_2827_0, i_10_344_2880_0, i_10_344_2887_0,
    i_10_344_2998_0, i_10_344_3007_0, i_10_344_3119_0, i_10_344_3197_0,
    i_10_344_3231_0, i_10_344_3290_0, i_10_344_3386_0, i_10_344_3451_0,
    i_10_344_3452_0, i_10_344_3466_0, i_10_344_3493_0, i_10_344_3501_0,
    i_10_344_3552_0, i_10_344_3589_0, i_10_344_3590_0, i_10_344_3616_0,
    i_10_344_3702_0, i_10_344_3788_0, i_10_344_3838_0, i_10_344_3858_0,
    i_10_344_3880_0, i_10_344_3883_0, i_10_344_3943_0, i_10_344_4055_0,
    i_10_344_4114_0, i_10_344_4115_0, i_10_344_4213_0, i_10_344_4217_0,
    i_10_344_4220_0, i_10_344_4281_0, i_10_344_4340_0, i_10_344_4451_0;
  output o_10_344_0_0;
  assign o_10_344_0_0 = 0;
endmodule



// Benchmark "kernel_10_345" written by ABC on Sun Jul 19 10:27:01 2020

module kernel_10_345 ( 
    i_10_345_269_0, i_10_345_283_0, i_10_345_284_0, i_10_345_286_0,
    i_10_345_327_0, i_10_345_408_0, i_10_345_409_0, i_10_345_410_0,
    i_10_345_413_0, i_10_345_441_0, i_10_345_444_0, i_10_345_520_0,
    i_10_345_521_0, i_10_345_718_0, i_10_345_793_0, i_10_345_797_0,
    i_10_345_1237_0, i_10_345_1238_0, i_10_345_1299_0, i_10_345_1310_0,
    i_10_345_1312_0, i_10_345_1313_0, i_10_345_1552_0, i_10_345_1555_0,
    i_10_345_1652_0, i_10_345_1819_0, i_10_345_1824_0, i_10_345_1826_0,
    i_10_345_1995_0, i_10_345_1996_0, i_10_345_2022_0, i_10_345_2185_0,
    i_10_345_2197_0, i_10_345_2200_0, i_10_345_2311_0, i_10_345_2312_0,
    i_10_345_2332_0, i_10_345_2352_0, i_10_345_2353_0, i_10_345_2354_0,
    i_10_345_2361_0, i_10_345_2376_0, i_10_345_2377_0, i_10_345_2378_0,
    i_10_345_2382_0, i_10_345_2383_0, i_10_345_2407_0, i_10_345_2410_0,
    i_10_345_2411_0, i_10_345_2462_0, i_10_345_2628_0, i_10_345_2632_0,
    i_10_345_2633_0, i_10_345_2658_0, i_10_345_2661_0, i_10_345_2718_0,
    i_10_345_2735_0, i_10_345_2782_0, i_10_345_2785_0, i_10_345_2788_0,
    i_10_345_2827_0, i_10_345_2828_0, i_10_345_2831_0, i_10_345_2922_0,
    i_10_345_2923_0, i_10_345_2924_0, i_10_345_2983_0, i_10_345_2986_0,
    i_10_345_3049_0, i_10_345_3050_0, i_10_345_3203_0, i_10_345_3271_0,
    i_10_345_3272_0, i_10_345_3282_0, i_10_345_3387_0, i_10_345_3389_0,
    i_10_345_3391_0, i_10_345_3392_0, i_10_345_3405_0, i_10_345_3408_0,
    i_10_345_3497_0, i_10_345_3652_0, i_10_345_3846_0, i_10_345_3847_0,
    i_10_345_3848_0, i_10_345_3851_0, i_10_345_3857_0, i_10_345_3858_0,
    i_10_345_3859_0, i_10_345_3895_0, i_10_345_3986_0, i_10_345_4129_0,
    i_10_345_4269_0, i_10_345_4270_0, i_10_345_4271_0, i_10_345_4277_0,
    i_10_345_4292_0, i_10_345_4567_0, i_10_345_4568_0, i_10_345_4569_0,
    o_10_345_0_0  );
  input  i_10_345_269_0, i_10_345_283_0, i_10_345_284_0, i_10_345_286_0,
    i_10_345_327_0, i_10_345_408_0, i_10_345_409_0, i_10_345_410_0,
    i_10_345_413_0, i_10_345_441_0, i_10_345_444_0, i_10_345_520_0,
    i_10_345_521_0, i_10_345_718_0, i_10_345_793_0, i_10_345_797_0,
    i_10_345_1237_0, i_10_345_1238_0, i_10_345_1299_0, i_10_345_1310_0,
    i_10_345_1312_0, i_10_345_1313_0, i_10_345_1552_0, i_10_345_1555_0,
    i_10_345_1652_0, i_10_345_1819_0, i_10_345_1824_0, i_10_345_1826_0,
    i_10_345_1995_0, i_10_345_1996_0, i_10_345_2022_0, i_10_345_2185_0,
    i_10_345_2197_0, i_10_345_2200_0, i_10_345_2311_0, i_10_345_2312_0,
    i_10_345_2332_0, i_10_345_2352_0, i_10_345_2353_0, i_10_345_2354_0,
    i_10_345_2361_0, i_10_345_2376_0, i_10_345_2377_0, i_10_345_2378_0,
    i_10_345_2382_0, i_10_345_2383_0, i_10_345_2407_0, i_10_345_2410_0,
    i_10_345_2411_0, i_10_345_2462_0, i_10_345_2628_0, i_10_345_2632_0,
    i_10_345_2633_0, i_10_345_2658_0, i_10_345_2661_0, i_10_345_2718_0,
    i_10_345_2735_0, i_10_345_2782_0, i_10_345_2785_0, i_10_345_2788_0,
    i_10_345_2827_0, i_10_345_2828_0, i_10_345_2831_0, i_10_345_2922_0,
    i_10_345_2923_0, i_10_345_2924_0, i_10_345_2983_0, i_10_345_2986_0,
    i_10_345_3049_0, i_10_345_3050_0, i_10_345_3203_0, i_10_345_3271_0,
    i_10_345_3272_0, i_10_345_3282_0, i_10_345_3387_0, i_10_345_3389_0,
    i_10_345_3391_0, i_10_345_3392_0, i_10_345_3405_0, i_10_345_3408_0,
    i_10_345_3497_0, i_10_345_3652_0, i_10_345_3846_0, i_10_345_3847_0,
    i_10_345_3848_0, i_10_345_3851_0, i_10_345_3857_0, i_10_345_3858_0,
    i_10_345_3859_0, i_10_345_3895_0, i_10_345_3986_0, i_10_345_4129_0,
    i_10_345_4269_0, i_10_345_4270_0, i_10_345_4271_0, i_10_345_4277_0,
    i_10_345_4292_0, i_10_345_4567_0, i_10_345_4568_0, i_10_345_4569_0;
  output o_10_345_0_0;
  assign o_10_345_0_0 = ~((~i_10_345_2828_0 & ((~i_10_345_520_0 & ((~i_10_345_521_0 & ~i_10_345_1552_0 & ~i_10_345_1995_0 & ~i_10_345_2200_0 & ~i_10_345_2377_0 & ~i_10_345_2378_0 & ~i_10_345_2462_0 & ~i_10_345_2735_0 & ~i_10_345_3857_0) | (~i_10_345_284_0 & i_10_345_2658_0 & i_10_345_3859_0))) | (~i_10_345_2353_0 & ((~i_10_345_2983_0 & ~i_10_345_3391_0 & ~i_10_345_3846_0 & ~i_10_345_3848_0 & ~i_10_345_3986_0 & ~i_10_345_4270_0) | (~i_10_345_410_0 & ~i_10_345_2312_0 & ~i_10_345_2376_0 & ~i_10_345_2986_0 & ~i_10_345_3895_0 & ~i_10_345_4277_0 & ~i_10_345_4567_0 & ~i_10_345_4568_0))) | (~i_10_345_283_0 & ~i_10_345_521_0 & ~i_10_345_2352_0 & ~i_10_345_2378_0 & ~i_10_345_2407_0 & ~i_10_345_2410_0 & ~i_10_345_2827_0 & ~i_10_345_3392_0))) | (~i_10_345_284_0 & ((i_10_345_286_0 & ~i_10_345_2312_0 & ~i_10_345_2376_0 & ~i_10_345_2382_0 & ~i_10_345_2411_0) | (~i_10_345_2377_0 & ~i_10_345_2378_0 & i_10_345_520_0 & ~i_10_345_1555_0 & ~i_10_345_2718_0 & ~i_10_345_2831_0 & ~i_10_345_3391_0 & ~i_10_345_3497_0 & ~i_10_345_3846_0))) | (~i_10_345_521_0 & ((i_10_345_1312_0 & ~i_10_345_2312_0 & ~i_10_345_2376_0 & ~i_10_345_2410_0 & ~i_10_345_2831_0) | (~i_10_345_327_0 & ~i_10_345_797_0 & ~i_10_345_1819_0 & ~i_10_345_2200_0 & ~i_10_345_2377_0 & ~i_10_345_2378_0 & ~i_10_345_3652_0 & ~i_10_345_3847_0 & ~i_10_345_3986_0))) | (~i_10_345_3282_0 & ((~i_10_345_1310_0 & ((~i_10_345_283_0 & ~i_10_345_327_0 & ~i_10_345_2185_0 & ~i_10_345_2377_0 & ~i_10_345_2378_0 & ~i_10_345_2382_0 & ~i_10_345_2462_0 & ~i_10_345_3272_0 & ~i_10_345_3497_0 & ~i_10_345_4292_0) | (~i_10_345_718_0 & ~i_10_345_797_0 & ~i_10_345_2332_0 & ~i_10_345_2361_0 & ~i_10_345_2628_0 & ~i_10_345_2658_0 & ~i_10_345_3846_0 & ~i_10_345_3857_0 & ~i_10_345_4271_0 & ~i_10_345_4568_0 & ~i_10_345_4569_0))) | (i_10_345_409_0 & ~i_10_345_1555_0 & ~i_10_345_2383_0 & ~i_10_345_2462_0 & ~i_10_345_2628_0 & ~i_10_345_2632_0 & ~i_10_345_2633_0))) | (~i_10_345_2352_0 & ((~i_10_345_283_0 & ((~i_10_345_2632_0 & ~i_10_345_2658_0 & i_10_345_2827_0 & ~i_10_345_3848_0) | (~i_10_345_2378_0 & ~i_10_345_3272_0 & ~i_10_345_3846_0 & ~i_10_345_3851_0 & i_10_345_3859_0))) | (~i_10_345_2983_0 & ((~i_10_345_327_0 & ~i_10_345_718_0 & ~i_10_345_2312_0 & ~i_10_345_2354_0 & ~i_10_345_2377_0 & ~i_10_345_2378_0 & ~i_10_345_2831_0 & ~i_10_345_3851_0) | (~i_10_345_3847_0 & ~i_10_345_4568_0 & i_10_345_4569_0))) | (i_10_345_2632_0 & i_10_345_2782_0))) | (i_10_345_1819_0 & ((~i_10_345_2633_0 & i_10_345_2658_0 & i_10_345_4567_0) | (~i_10_345_2377_0 & i_10_345_2782_0 & ~i_10_345_4568_0))) | (~i_10_345_2312_0 & ((~i_10_345_2332_0 & ~i_10_345_2827_0 & ~i_10_345_3846_0 & i_10_345_4129_0 & ~i_10_345_4277_0) | (~i_10_345_327_0 & i_10_345_1826_0 & ~i_10_345_2378_0 & ~i_10_345_3895_0 & ~i_10_345_4567_0 & ~i_10_345_4568_0))) | (~i_10_345_4292_0 & ((~i_10_345_327_0 & ~i_10_345_4277_0 & ((~i_10_345_2462_0 & i_10_345_2632_0 & ~i_10_345_3857_0 & i_10_345_3858_0) | (~i_10_345_718_0 & ~i_10_345_1555_0 & ~i_10_345_2197_0 & ~i_10_345_2361_0 & ~i_10_345_4271_0 & ~i_10_345_4568_0 & ~i_10_345_4569_0 & ~i_10_345_2376_0 & ~i_10_345_2377_0))) | (~i_10_345_2197_0 & ((~i_10_345_444_0 & ~i_10_345_2377_0 & ~i_10_345_2378_0 & ~i_10_345_2633_0 & ~i_10_345_2986_0 & ~i_10_345_3203_0 & ~i_10_345_3408_0 & ~i_10_345_3847_0) | (~i_10_345_718_0 & ~i_10_345_2411_0 & ~i_10_345_3389_0 & i_10_345_3652_0 & ~i_10_345_4569_0))))) | (~i_10_345_2378_0 & ((~i_10_345_1555_0 & ((i_10_345_441_0 & ~i_10_345_2332_0 & ~i_10_345_2353_0 & ~i_10_345_3848_0) | (~i_10_345_718_0 & ~i_10_345_2376_0 & i_10_345_2735_0 & ~i_10_345_2827_0 & ~i_10_345_2831_0 & ~i_10_345_3895_0))) | (~i_10_345_2332_0 & i_10_345_2382_0 & ~i_10_345_2827_0 & ~i_10_345_2983_0 & ~i_10_345_2986_0 & ~i_10_345_3652_0))) | (~i_10_345_2353_0 & ~i_10_345_2377_0 & i_10_345_2924_0 & ~i_10_345_3391_0 & ~i_10_345_3392_0) | (i_10_345_327_0 & i_10_345_1824_0 & ~i_10_345_2983_0 & ~i_10_345_4567_0));
endmodule



// Benchmark "kernel_10_346" written by ABC on Sun Jul 19 10:27:02 2020

module kernel_10_346 ( 
    i_10_346_86_0, i_10_346_172_0, i_10_346_173_0, i_10_346_181_0,
    i_10_346_185_0, i_10_346_326_0, i_10_346_446_0, i_10_346_449_0,
    i_10_346_499_0, i_10_346_588_0, i_10_346_591_0, i_10_346_800_0,
    i_10_346_971_0, i_10_346_1234_0, i_10_346_1238_0, i_10_346_1246_0,
    i_10_346_1273_0, i_10_346_1363_0, i_10_346_1367_0, i_10_346_1412_0,
    i_10_346_1543_0, i_10_346_1553_0, i_10_346_1648_0, i_10_346_1651_0,
    i_10_346_1655_0, i_10_346_1760_0, i_10_346_1765_0, i_10_346_1777_0,
    i_10_346_1819_0, i_10_346_1820_0, i_10_346_1822_0, i_10_346_1825_0,
    i_10_346_1886_0, i_10_346_1888_0, i_10_346_1909_0, i_10_346_1949_0,
    i_10_346_2093_0, i_10_346_2096_0, i_10_346_2311_0, i_10_346_2336_0,
    i_10_346_2339_0, i_10_346_2448_0, i_10_346_2449_0, i_10_346_2450_0,
    i_10_346_2456_0, i_10_346_2543_0, i_10_346_2606_0, i_10_346_2638_0,
    i_10_346_2642_0, i_10_346_2702_0, i_10_346_2703_0, i_10_346_2725_0,
    i_10_346_2731_0, i_10_346_2788_0, i_10_346_2833_0, i_10_346_2866_0,
    i_10_346_2867_0, i_10_346_2869_0, i_10_346_2870_0, i_10_346_2917_0,
    i_10_346_2920_0, i_10_346_2923_0, i_10_346_3033_0, i_10_346_3037_0,
    i_10_346_3040_0, i_10_346_3092_0, i_10_346_3196_0, i_10_346_3197_0,
    i_10_346_3199_0, i_10_346_3202_0, i_10_346_3203_0, i_10_346_3386_0,
    i_10_346_3390_0, i_10_346_3392_0, i_10_346_3471_0, i_10_346_3586_0,
    i_10_346_3587_0, i_10_346_3588_0, i_10_346_3589_0, i_10_346_3611_0,
    i_10_346_3683_0, i_10_346_3731_0, i_10_346_3734_0, i_10_346_3884_0,
    i_10_346_3923_0, i_10_346_3964_0, i_10_346_3965_0, i_10_346_4117_0,
    i_10_346_4118_0, i_10_346_4120_0, i_10_346_4180_0, i_10_346_4267_0,
    i_10_346_4274_0, i_10_346_4283_0, i_10_346_4310_0, i_10_346_4561_0,
    i_10_346_4588_0, i_10_346_4592_0, i_10_346_4603_0, i_10_346_4604_0,
    o_10_346_0_0  );
  input  i_10_346_86_0, i_10_346_172_0, i_10_346_173_0, i_10_346_181_0,
    i_10_346_185_0, i_10_346_326_0, i_10_346_446_0, i_10_346_449_0,
    i_10_346_499_0, i_10_346_588_0, i_10_346_591_0, i_10_346_800_0,
    i_10_346_971_0, i_10_346_1234_0, i_10_346_1238_0, i_10_346_1246_0,
    i_10_346_1273_0, i_10_346_1363_0, i_10_346_1367_0, i_10_346_1412_0,
    i_10_346_1543_0, i_10_346_1553_0, i_10_346_1648_0, i_10_346_1651_0,
    i_10_346_1655_0, i_10_346_1760_0, i_10_346_1765_0, i_10_346_1777_0,
    i_10_346_1819_0, i_10_346_1820_0, i_10_346_1822_0, i_10_346_1825_0,
    i_10_346_1886_0, i_10_346_1888_0, i_10_346_1909_0, i_10_346_1949_0,
    i_10_346_2093_0, i_10_346_2096_0, i_10_346_2311_0, i_10_346_2336_0,
    i_10_346_2339_0, i_10_346_2448_0, i_10_346_2449_0, i_10_346_2450_0,
    i_10_346_2456_0, i_10_346_2543_0, i_10_346_2606_0, i_10_346_2638_0,
    i_10_346_2642_0, i_10_346_2702_0, i_10_346_2703_0, i_10_346_2725_0,
    i_10_346_2731_0, i_10_346_2788_0, i_10_346_2833_0, i_10_346_2866_0,
    i_10_346_2867_0, i_10_346_2869_0, i_10_346_2870_0, i_10_346_2917_0,
    i_10_346_2920_0, i_10_346_2923_0, i_10_346_3033_0, i_10_346_3037_0,
    i_10_346_3040_0, i_10_346_3092_0, i_10_346_3196_0, i_10_346_3197_0,
    i_10_346_3199_0, i_10_346_3202_0, i_10_346_3203_0, i_10_346_3386_0,
    i_10_346_3390_0, i_10_346_3392_0, i_10_346_3471_0, i_10_346_3586_0,
    i_10_346_3587_0, i_10_346_3588_0, i_10_346_3589_0, i_10_346_3611_0,
    i_10_346_3683_0, i_10_346_3731_0, i_10_346_3734_0, i_10_346_3884_0,
    i_10_346_3923_0, i_10_346_3964_0, i_10_346_3965_0, i_10_346_4117_0,
    i_10_346_4118_0, i_10_346_4120_0, i_10_346_4180_0, i_10_346_4267_0,
    i_10_346_4274_0, i_10_346_4283_0, i_10_346_4310_0, i_10_346_4561_0,
    i_10_346_4588_0, i_10_346_4592_0, i_10_346_4603_0, i_10_346_4604_0;
  output o_10_346_0_0;
  assign o_10_346_0_0 = 0;
endmodule



// Benchmark "kernel_10_347" written by ABC on Sun Jul 19 10:27:04 2020

module kernel_10_347 ( 
    i_10_347_247_0, i_10_347_330_0, i_10_347_393_0, i_10_347_405_0,
    i_10_347_423_0, i_10_347_424_0, i_10_347_438_0, i_10_347_442_0,
    i_10_347_444_0, i_10_347_459_0, i_10_347_463_0, i_10_347_464_0,
    i_10_347_467_0, i_10_347_507_0, i_10_347_562_0, i_10_347_711_0,
    i_10_347_792_0, i_10_347_956_0, i_10_347_1026_0, i_10_347_1305_0,
    i_10_347_1438_0, i_10_347_1548_0, i_10_347_1579_0, i_10_347_1654_0,
    i_10_347_1655_0, i_10_347_1683_0, i_10_347_1819_0, i_10_347_1821_0,
    i_10_347_1913_0, i_10_347_2202_0, i_10_347_2337_0, i_10_347_2350_0,
    i_10_347_2351_0, i_10_347_2352_0, i_10_347_2353_0, i_10_347_2354_0,
    i_10_347_2355_0, i_10_347_2365_0, i_10_347_2379_0, i_10_347_2451_0,
    i_10_347_2452_0, i_10_347_2571_0, i_10_347_2633_0, i_10_347_2634_0,
    i_10_347_2658_0, i_10_347_2701_0, i_10_347_2710_0, i_10_347_2732_0,
    i_10_347_2733_0, i_10_347_2781_0, i_10_347_2830_0, i_10_347_2883_0,
    i_10_347_2884_0, i_10_347_2888_0, i_10_347_2922_0, i_10_347_2985_0,
    i_10_347_3038_0, i_10_347_3048_0, i_10_347_3087_0, i_10_347_3152_0,
    i_10_347_3154_0, i_10_347_3165_0, i_10_347_3198_0, i_10_347_3199_0,
    i_10_347_3277_0, i_10_347_3280_0, i_10_347_3283_0, i_10_347_3385_0,
    i_10_347_3386_0, i_10_347_3405_0, i_10_347_3406_0, i_10_347_3408_0,
    i_10_347_3471_0, i_10_347_3610_0, i_10_347_3612_0, i_10_347_3613_0,
    i_10_347_3616_0, i_10_347_3702_0, i_10_347_3834_0, i_10_347_3837_0,
    i_10_347_3847_0, i_10_347_3850_0, i_10_347_3851_0, i_10_347_3855_0,
    i_10_347_3894_0, i_10_347_3982_0, i_10_347_4027_0, i_10_347_4116_0,
    i_10_347_4117_0, i_10_347_4120_0, i_10_347_4125_0, i_10_347_4126_0,
    i_10_347_4127_0, i_10_347_4285_0, i_10_347_4292_0, i_10_347_4563_0,
    i_10_347_4564_0, i_10_347_4566_0, i_10_347_4567_0, i_10_347_4568_0,
    o_10_347_0_0  );
  input  i_10_347_247_0, i_10_347_330_0, i_10_347_393_0, i_10_347_405_0,
    i_10_347_423_0, i_10_347_424_0, i_10_347_438_0, i_10_347_442_0,
    i_10_347_444_0, i_10_347_459_0, i_10_347_463_0, i_10_347_464_0,
    i_10_347_467_0, i_10_347_507_0, i_10_347_562_0, i_10_347_711_0,
    i_10_347_792_0, i_10_347_956_0, i_10_347_1026_0, i_10_347_1305_0,
    i_10_347_1438_0, i_10_347_1548_0, i_10_347_1579_0, i_10_347_1654_0,
    i_10_347_1655_0, i_10_347_1683_0, i_10_347_1819_0, i_10_347_1821_0,
    i_10_347_1913_0, i_10_347_2202_0, i_10_347_2337_0, i_10_347_2350_0,
    i_10_347_2351_0, i_10_347_2352_0, i_10_347_2353_0, i_10_347_2354_0,
    i_10_347_2355_0, i_10_347_2365_0, i_10_347_2379_0, i_10_347_2451_0,
    i_10_347_2452_0, i_10_347_2571_0, i_10_347_2633_0, i_10_347_2634_0,
    i_10_347_2658_0, i_10_347_2701_0, i_10_347_2710_0, i_10_347_2732_0,
    i_10_347_2733_0, i_10_347_2781_0, i_10_347_2830_0, i_10_347_2883_0,
    i_10_347_2884_0, i_10_347_2888_0, i_10_347_2922_0, i_10_347_2985_0,
    i_10_347_3038_0, i_10_347_3048_0, i_10_347_3087_0, i_10_347_3152_0,
    i_10_347_3154_0, i_10_347_3165_0, i_10_347_3198_0, i_10_347_3199_0,
    i_10_347_3277_0, i_10_347_3280_0, i_10_347_3283_0, i_10_347_3385_0,
    i_10_347_3386_0, i_10_347_3405_0, i_10_347_3406_0, i_10_347_3408_0,
    i_10_347_3471_0, i_10_347_3610_0, i_10_347_3612_0, i_10_347_3613_0,
    i_10_347_3616_0, i_10_347_3702_0, i_10_347_3834_0, i_10_347_3837_0,
    i_10_347_3847_0, i_10_347_3850_0, i_10_347_3851_0, i_10_347_3855_0,
    i_10_347_3894_0, i_10_347_3982_0, i_10_347_4027_0, i_10_347_4116_0,
    i_10_347_4117_0, i_10_347_4120_0, i_10_347_4125_0, i_10_347_4126_0,
    i_10_347_4127_0, i_10_347_4285_0, i_10_347_4292_0, i_10_347_4563_0,
    i_10_347_4564_0, i_10_347_4566_0, i_10_347_4567_0, i_10_347_4568_0;
  output o_10_347_0_0;
  assign o_10_347_0_0 = ~((~i_10_347_423_0 & ((~i_10_347_711_0 & i_10_347_1819_0 & i_10_347_2732_0 & ~i_10_347_3408_0 & ~i_10_347_3471_0) | (~i_10_347_424_0 & ~i_10_347_438_0 & ~i_10_347_1026_0 & ~i_10_347_1305_0 & ~i_10_347_2658_0 & ~i_10_347_2884_0 & i_10_347_4120_0))) | (~i_10_347_442_0 & ((~i_10_347_424_0 & ~i_10_347_438_0 & ~i_10_347_464_0 & ~i_10_347_2202_0 & ~i_10_347_2451_0 & ~i_10_347_2733_0 & ~i_10_347_3280_0 & ~i_10_347_3405_0) | (~i_10_347_459_0 & i_10_347_1819_0 & ~i_10_347_3612_0 & ~i_10_347_3613_0 & ~i_10_347_4120_0 & ~i_10_347_4127_0))) | (i_10_347_464_0 & ((~i_10_347_1548_0 & ~i_10_347_1579_0 & ~i_10_347_2884_0 & ~i_10_347_3280_0 & ~i_10_347_3610_0 & ~i_10_347_3612_0 & ~i_10_347_3837_0) | (~i_10_347_438_0 & ~i_10_347_1026_0 & ~i_10_347_1683_0 & ~i_10_347_1913_0 & ~i_10_347_2633_0 & ~i_10_347_2883_0 & ~i_10_347_3087_0 & ~i_10_347_3834_0 & ~i_10_347_3855_0))) | (~i_10_347_2451_0 & ((~i_10_347_438_0 & ((~i_10_347_711_0 & ~i_10_347_2452_0 & ~i_10_347_3048_0 & i_10_347_3198_0 & ~i_10_347_3386_0 & ~i_10_347_3612_0) | (i_10_347_1579_0 & ~i_10_347_2883_0 & ~i_10_347_3405_0 & ~i_10_347_3616_0))) | (i_10_347_467_0 & ((~i_10_347_562_0 & ~i_10_347_2634_0 & ~i_10_347_2733_0 & ~i_10_347_2888_0 & ~i_10_347_3408_0 & ~i_10_347_3471_0) | (i_10_347_2658_0 & ~i_10_347_3048_0 & i_10_347_4027_0 & ~i_10_347_4117_0))) | (~i_10_347_3087_0 & ~i_10_347_3280_0 & ((i_10_347_459_0 & ~i_10_347_467_0 & ~i_10_347_792_0 & ~i_10_347_1438_0 & ~i_10_347_3038_0 & ~i_10_347_3385_0) | (~i_10_347_2634_0 & ~i_10_347_3616_0 & ~i_10_347_3837_0 & ~i_10_347_4285_0 & ~i_10_347_4566_0))) | (~i_10_347_424_0 & ~i_10_347_711_0 & ~i_10_347_2888_0 & ~i_10_347_3048_0 & ~i_10_347_3198_0 & ~i_10_347_4292_0))) | (~i_10_347_3610_0 & ((~i_10_347_393_0 & ~i_10_347_3165_0 & ~i_10_347_3613_0 & ((~i_10_347_424_0 & ~i_10_347_2571_0 & ~i_10_347_2633_0 & ~i_10_347_2710_0 & ~i_10_347_2883_0 & ~i_10_347_3471_0 & ~i_10_347_3850_0) | (~i_10_347_1683_0 & ~i_10_347_2733_0 & ~i_10_347_2884_0 & ~i_10_347_3277_0 & ~i_10_347_4292_0))) | (~i_10_347_424_0 & ~i_10_347_1683_0 & ~i_10_347_2353_0 & ~i_10_347_2354_0 & ~i_10_347_2634_0 & ~i_10_347_2883_0 & ~i_10_347_2922_0 & ~i_10_347_3405_0 & ~i_10_347_3612_0) | (~i_10_347_2733_0 & ~i_10_347_3038_0 & ~i_10_347_3087_0 & ~i_10_347_3198_0 & ~i_10_347_3277_0 & ~i_10_347_3283_0 & ~i_10_347_3406_0 & ~i_10_347_4567_0))) | (~i_10_347_393_0 & ~i_10_347_1026_0 & ~i_10_347_2710_0 & ((~i_10_347_247_0 & ~i_10_347_467_0 & ~i_10_347_1683_0 & ~i_10_347_2354_0 & ~i_10_347_2781_0 & ~i_10_347_3199_0 & ~i_10_347_3837_0 & ~i_10_347_3855_0) | (i_10_347_1819_0 & ~i_10_347_3087_0 & ~i_10_347_3405_0 & ~i_10_347_3616_0 & ~i_10_347_4120_0))) | (~i_10_347_438_0 & ~i_10_347_2884_0 & ~i_10_347_3855_0 & ((~i_10_347_1821_0 & ~i_10_347_1913_0 & i_10_347_2633_0 & ~i_10_347_3087_0) | (~i_10_347_956_0 & ~i_10_347_1819_0 & i_10_347_2452_0 & ~i_10_347_2658_0 & ~i_10_347_3850_0))) | (~i_10_347_1438_0 & ((~i_10_347_711_0 & ~i_10_347_3198_0 & ((~i_10_347_2337_0 & ~i_10_347_3612_0 & i_10_347_4027_0) | (~i_10_347_2379_0 & ~i_10_347_3613_0 & i_10_347_4285_0))) | (~i_10_347_1305_0 & ~i_10_347_2452_0 & ~i_10_347_2633_0 & ~i_10_347_2883_0 & ~i_10_347_3277_0 & ~i_10_347_3385_0 & ~i_10_347_3408_0 & ~i_10_347_3616_0 & ~i_10_347_3834_0 & ~i_10_347_4566_0))) | (i_10_347_4126_0 & (i_10_347_2732_0 | (i_10_347_2351_0 & ~i_10_347_2634_0 & ~i_10_347_2888_0))) | (i_10_347_792_0 & i_10_347_2781_0 & ~i_10_347_3087_0 & ~i_10_347_3280_0) | (i_10_347_2830_0 & i_10_347_3087_0 & ~i_10_347_3894_0) | (~i_10_347_444_0 & ~i_10_347_464_0 & ~i_10_347_792_0 & ~i_10_347_1683_0 & i_10_347_2633_0 & i_10_347_4117_0) | (~i_10_347_3198_0 & ~i_10_347_3405_0 & i_10_347_4568_0));
endmodule



// Benchmark "kernel_10_348" written by ABC on Sun Jul 19 10:27:05 2020

module kernel_10_348 ( 
    i_10_348_171_0, i_10_348_174_0, i_10_348_175_0, i_10_348_184_0,
    i_10_348_220_0, i_10_348_223_0, i_10_348_247_0, i_10_348_265_0,
    i_10_348_269_0, i_10_348_270_0, i_10_348_271_0, i_10_348_273_0,
    i_10_348_283_0, i_10_348_284_0, i_10_348_287_0, i_10_348_395_0,
    i_10_348_405_0, i_10_348_408_0, i_10_348_412_0, i_10_348_436_0,
    i_10_348_798_0, i_10_348_958_0, i_10_348_1004_0, i_10_348_1006_0,
    i_10_348_1085_0, i_10_348_1310_0, i_10_348_1434_0, i_10_348_1435_0,
    i_10_348_1438_0, i_10_348_1451_0, i_10_348_1547_0, i_10_348_1554_0,
    i_10_348_1555_0, i_10_348_1619_0, i_10_348_1877_0, i_10_348_1945_0,
    i_10_348_1947_0, i_10_348_1948_0, i_10_348_1949_0, i_10_348_1951_0,
    i_10_348_1952_0, i_10_348_2185_0, i_10_348_2310_0, i_10_348_2312_0,
    i_10_348_2350_0, i_10_348_2353_0, i_10_348_2354_0, i_10_348_2356_0,
    i_10_348_2357_0, i_10_348_2407_0, i_10_348_2408_0, i_10_348_2411_0,
    i_10_348_2449_0, i_10_348_2470_0, i_10_348_2471_0, i_10_348_2510_0,
    i_10_348_2663_0, i_10_348_2681_0, i_10_348_2730_0, i_10_348_2781_0,
    i_10_348_2821_0, i_10_348_2920_0, i_10_348_2921_0, i_10_348_2923_0,
    i_10_348_2924_0, i_10_348_3034_0, i_10_348_3047_0, i_10_348_3050_0,
    i_10_348_3077_0, i_10_348_3090_0, i_10_348_3151_0, i_10_348_3157_0,
    i_10_348_3199_0, i_10_348_3272_0, i_10_348_3275_0, i_10_348_3281_0,
    i_10_348_3301_0, i_10_348_3384_0, i_10_348_3385_0, i_10_348_3392_0,
    i_10_348_3472_0, i_10_348_3473_0, i_10_348_3545_0, i_10_348_3560_0,
    i_10_348_3586_0, i_10_348_3588_0, i_10_348_3590_0, i_10_348_3784_0,
    i_10_348_3859_0, i_10_348_3895_0, i_10_348_3986_0, i_10_348_4054_0,
    i_10_348_4115_0, i_10_348_4116_0, i_10_348_4117_0, i_10_348_4118_0,
    i_10_348_4273_0, i_10_348_4283_0, i_10_348_4285_0, i_10_348_4567_0,
    o_10_348_0_0  );
  input  i_10_348_171_0, i_10_348_174_0, i_10_348_175_0, i_10_348_184_0,
    i_10_348_220_0, i_10_348_223_0, i_10_348_247_0, i_10_348_265_0,
    i_10_348_269_0, i_10_348_270_0, i_10_348_271_0, i_10_348_273_0,
    i_10_348_283_0, i_10_348_284_0, i_10_348_287_0, i_10_348_395_0,
    i_10_348_405_0, i_10_348_408_0, i_10_348_412_0, i_10_348_436_0,
    i_10_348_798_0, i_10_348_958_0, i_10_348_1004_0, i_10_348_1006_0,
    i_10_348_1085_0, i_10_348_1310_0, i_10_348_1434_0, i_10_348_1435_0,
    i_10_348_1438_0, i_10_348_1451_0, i_10_348_1547_0, i_10_348_1554_0,
    i_10_348_1555_0, i_10_348_1619_0, i_10_348_1877_0, i_10_348_1945_0,
    i_10_348_1947_0, i_10_348_1948_0, i_10_348_1949_0, i_10_348_1951_0,
    i_10_348_1952_0, i_10_348_2185_0, i_10_348_2310_0, i_10_348_2312_0,
    i_10_348_2350_0, i_10_348_2353_0, i_10_348_2354_0, i_10_348_2356_0,
    i_10_348_2357_0, i_10_348_2407_0, i_10_348_2408_0, i_10_348_2411_0,
    i_10_348_2449_0, i_10_348_2470_0, i_10_348_2471_0, i_10_348_2510_0,
    i_10_348_2663_0, i_10_348_2681_0, i_10_348_2730_0, i_10_348_2781_0,
    i_10_348_2821_0, i_10_348_2920_0, i_10_348_2921_0, i_10_348_2923_0,
    i_10_348_2924_0, i_10_348_3034_0, i_10_348_3047_0, i_10_348_3050_0,
    i_10_348_3077_0, i_10_348_3090_0, i_10_348_3151_0, i_10_348_3157_0,
    i_10_348_3199_0, i_10_348_3272_0, i_10_348_3275_0, i_10_348_3281_0,
    i_10_348_3301_0, i_10_348_3384_0, i_10_348_3385_0, i_10_348_3392_0,
    i_10_348_3472_0, i_10_348_3473_0, i_10_348_3545_0, i_10_348_3560_0,
    i_10_348_3586_0, i_10_348_3588_0, i_10_348_3590_0, i_10_348_3784_0,
    i_10_348_3859_0, i_10_348_3895_0, i_10_348_3986_0, i_10_348_4054_0,
    i_10_348_4115_0, i_10_348_4116_0, i_10_348_4117_0, i_10_348_4118_0,
    i_10_348_4273_0, i_10_348_4283_0, i_10_348_4285_0, i_10_348_4567_0;
  output o_10_348_0_0;
  assign o_10_348_0_0 = ~((~i_10_348_269_0 & ((~i_10_348_1004_0 & ~i_10_348_1006_0 & ~i_10_348_1555_0 & ~i_10_348_2185_0 & ~i_10_348_3090_0) | (~i_10_348_1948_0 & ~i_10_348_2312_0 & ~i_10_348_3545_0))) | (~i_10_348_1004_0 & ((~i_10_348_265_0 & ~i_10_348_2312_0 & ~i_10_348_2357_0) | (~i_10_348_395_0 & ~i_10_348_958_0 & ~i_10_348_1877_0 & ~i_10_348_1947_0 & ~i_10_348_1948_0 & ~i_10_348_3392_0))) | (~i_10_348_395_0 & ((~i_10_348_1435_0 & i_10_348_2354_0 & i_10_348_3472_0) | (~i_10_348_2408_0 & ~i_10_348_3077_0 & ~i_10_348_3588_0 & i_10_348_3986_0 & ~i_10_348_4054_0))) | (~i_10_348_2312_0 & ((~i_10_348_1438_0 & ((i_10_348_1434_0 & i_10_348_2730_0 & ~i_10_348_3473_0) | (i_10_348_2923_0 & ~i_10_348_3986_0))) | (i_10_348_1952_0 & i_10_348_2924_0 & ~i_10_348_3895_0))) | (~i_10_348_1952_0 & ((~i_10_348_1555_0 & ((~i_10_348_1949_0 & ~i_10_348_3392_0 & ~i_10_348_3545_0) | (i_10_348_287_0 & ~i_10_348_1554_0 & ~i_10_348_2449_0 & i_10_348_2470_0 & ~i_10_348_4116_0 & i_10_348_4273_0))) | (~i_10_348_2681_0 & i_10_348_3050_0 & ~i_10_348_3473_0))) | (~i_10_348_1947_0 & ((i_10_348_1310_0 & ~i_10_348_1619_0 & ~i_10_348_2357_0 & ~i_10_348_3034_0 & ~i_10_348_3281_0) | (~i_10_348_175_0 & ~i_10_348_436_0 & ~i_10_348_798_0 & ~i_10_348_1951_0 & ~i_10_348_2510_0 & ~i_10_348_3545_0))) | (~i_10_348_3473_0 & ((~i_10_348_1434_0 & ~i_10_348_2411_0 & ~i_10_348_2510_0) | (~i_10_348_283_0 & ~i_10_348_4054_0 & ~i_10_348_4567_0))) | (~i_10_348_284_0 & ~i_10_348_1085_0 & ~i_10_348_1951_0 & ~i_10_348_2681_0 & ~i_10_348_3986_0 & ~i_10_348_4116_0));
endmodule



// Benchmark "kernel_10_349" written by ABC on Sun Jul 19 10:27:06 2020

module kernel_10_349 ( 
    i_10_349_17_0, i_10_349_67_0, i_10_349_118_0, i_10_349_245_0,
    i_10_349_252_0, i_10_349_279_0, i_10_349_281_0, i_10_349_317_0,
    i_10_349_320_0, i_10_349_325_0, i_10_349_326_0, i_10_349_389_0,
    i_10_349_395_0, i_10_349_410_0, i_10_349_428_0, i_10_349_434_0,
    i_10_349_442_0, i_10_349_464_0, i_10_349_506_0, i_10_349_792_0,
    i_10_349_968_0, i_10_349_994_0, i_10_349_1098_0, i_10_349_1235_0,
    i_10_349_1307_0, i_10_349_1311_0, i_10_349_1313_0, i_10_349_1343_0,
    i_10_349_1379_0, i_10_349_1454_0, i_10_349_1456_0, i_10_349_1544_0,
    i_10_349_1547_0, i_10_349_1576_0, i_10_349_1625_0, i_10_349_1655_0,
    i_10_349_1985_0, i_10_349_1993_0, i_10_349_1994_0, i_10_349_1997_0,
    i_10_349_2201_0, i_10_349_2203_0, i_10_349_2443_0, i_10_349_2444_0,
    i_10_349_2448_0, i_10_349_2450_0, i_10_349_2455_0, i_10_349_2456_0,
    i_10_349_2471_0, i_10_349_2529_0, i_10_349_2534_0, i_10_349_2584_0,
    i_10_349_2592_0, i_10_349_2639_0, i_10_349_2703_0, i_10_349_2705_0,
    i_10_349_2713_0, i_10_349_2716_0, i_10_349_2717_0, i_10_349_2828_0,
    i_10_349_2830_0, i_10_349_2834_0, i_10_349_2867_0, i_10_349_2870_0,
    i_10_349_2881_0, i_10_349_2882_0, i_10_349_2884_0, i_10_349_2885_0,
    i_10_349_2984_0, i_10_349_3041_0, i_10_349_3277_0, i_10_349_3278_0,
    i_10_349_3317_0, i_10_349_3384_0, i_10_349_3388_0, i_10_349_3409_0,
    i_10_349_3452_0, i_10_349_3523_0, i_10_349_3610_0, i_10_349_3611_0,
    i_10_349_3615_0, i_10_349_3653_0, i_10_349_3700_0, i_10_349_3703_0,
    i_10_349_3775_0, i_10_349_3836_0, i_10_349_3837_0, i_10_349_3857_0,
    i_10_349_3860_0, i_10_349_3912_0, i_10_349_3914_0, i_10_349_3983_0,
    i_10_349_4163_0, i_10_349_4175_0, i_10_349_4214_0, i_10_349_4273_0,
    i_10_349_4283_0, i_10_349_4288_0, i_10_349_4588_0, i_10_349_4592_0,
    o_10_349_0_0  );
  input  i_10_349_17_0, i_10_349_67_0, i_10_349_118_0, i_10_349_245_0,
    i_10_349_252_0, i_10_349_279_0, i_10_349_281_0, i_10_349_317_0,
    i_10_349_320_0, i_10_349_325_0, i_10_349_326_0, i_10_349_389_0,
    i_10_349_395_0, i_10_349_410_0, i_10_349_428_0, i_10_349_434_0,
    i_10_349_442_0, i_10_349_464_0, i_10_349_506_0, i_10_349_792_0,
    i_10_349_968_0, i_10_349_994_0, i_10_349_1098_0, i_10_349_1235_0,
    i_10_349_1307_0, i_10_349_1311_0, i_10_349_1313_0, i_10_349_1343_0,
    i_10_349_1379_0, i_10_349_1454_0, i_10_349_1456_0, i_10_349_1544_0,
    i_10_349_1547_0, i_10_349_1576_0, i_10_349_1625_0, i_10_349_1655_0,
    i_10_349_1985_0, i_10_349_1993_0, i_10_349_1994_0, i_10_349_1997_0,
    i_10_349_2201_0, i_10_349_2203_0, i_10_349_2443_0, i_10_349_2444_0,
    i_10_349_2448_0, i_10_349_2450_0, i_10_349_2455_0, i_10_349_2456_0,
    i_10_349_2471_0, i_10_349_2529_0, i_10_349_2534_0, i_10_349_2584_0,
    i_10_349_2592_0, i_10_349_2639_0, i_10_349_2703_0, i_10_349_2705_0,
    i_10_349_2713_0, i_10_349_2716_0, i_10_349_2717_0, i_10_349_2828_0,
    i_10_349_2830_0, i_10_349_2834_0, i_10_349_2867_0, i_10_349_2870_0,
    i_10_349_2881_0, i_10_349_2882_0, i_10_349_2884_0, i_10_349_2885_0,
    i_10_349_2984_0, i_10_349_3041_0, i_10_349_3277_0, i_10_349_3278_0,
    i_10_349_3317_0, i_10_349_3384_0, i_10_349_3388_0, i_10_349_3409_0,
    i_10_349_3452_0, i_10_349_3523_0, i_10_349_3610_0, i_10_349_3611_0,
    i_10_349_3615_0, i_10_349_3653_0, i_10_349_3700_0, i_10_349_3703_0,
    i_10_349_3775_0, i_10_349_3836_0, i_10_349_3837_0, i_10_349_3857_0,
    i_10_349_3860_0, i_10_349_3912_0, i_10_349_3914_0, i_10_349_3983_0,
    i_10_349_4163_0, i_10_349_4175_0, i_10_349_4214_0, i_10_349_4273_0,
    i_10_349_4283_0, i_10_349_4288_0, i_10_349_4588_0, i_10_349_4592_0;
  output o_10_349_0_0;
  assign o_10_349_0_0 = 0;
endmodule



// Benchmark "kernel_10_350" written by ABC on Sun Jul 19 10:27:06 2020

module kernel_10_350 ( 
    i_10_350_27_0, i_10_350_220_0, i_10_350_249_0, i_10_350_282_0,
    i_10_350_284_0, i_10_350_293_0, i_10_350_327_0, i_10_350_412_0,
    i_10_350_428_0, i_10_350_517_0, i_10_350_518_0, i_10_350_520_0,
    i_10_350_798_0, i_10_350_800_0, i_10_350_955_0, i_10_350_957_0,
    i_10_350_961_0, i_10_350_1033_0, i_10_350_1035_0, i_10_350_1152_0,
    i_10_350_1243_0, i_10_350_1245_0, i_10_350_1246_0, i_10_350_1247_0,
    i_10_350_1310_0, i_10_350_1311_0, i_10_350_1384_0, i_10_350_1539_0,
    i_10_350_1617_0, i_10_350_1683_0, i_10_350_1686_0, i_10_350_1690_0,
    i_10_350_1691_0, i_10_350_1820_0, i_10_350_1822_0, i_10_350_1825_0,
    i_10_350_1908_0, i_10_350_1911_0, i_10_350_1912_0, i_10_350_2186_0,
    i_10_350_2349_0, i_10_350_2350_0, i_10_350_2360_0, i_10_350_2361_0,
    i_10_350_2406_0, i_10_350_2452_0, i_10_350_2467_0, i_10_350_2468_0,
    i_10_350_2470_0, i_10_350_2473_0, i_10_350_2655_0, i_10_350_2679_0,
    i_10_350_2719_0, i_10_350_2725_0, i_10_350_2726_0, i_10_350_2740_0,
    i_10_350_2827_0, i_10_350_3036_0, i_10_350_3048_0, i_10_350_3074_0,
    i_10_350_3075_0, i_10_350_3201_0, i_10_350_3269_0, i_10_350_3387_0,
    i_10_350_3391_0, i_10_350_3392_0, i_10_350_3453_0, i_10_350_3520_0,
    i_10_350_3523_0, i_10_350_3609_0, i_10_350_3612_0, i_10_350_3613_0,
    i_10_350_3614_0, i_10_350_3617_0, i_10_350_3624_0, i_10_350_3648_0,
    i_10_350_3651_0, i_10_350_3652_0, i_10_350_3706_0, i_10_350_3723_0,
    i_10_350_3730_0, i_10_350_3780_0, i_10_350_3834_0, i_10_350_3835_0,
    i_10_350_3839_0, i_10_350_3840_0, i_10_350_3860_0, i_10_350_3993_0,
    i_10_350_4114_0, i_10_350_4120_0, i_10_350_4126_0, i_10_350_4215_0,
    i_10_350_4216_0, i_10_350_4219_0, i_10_350_4236_0, i_10_350_4273_0,
    i_10_350_4291_0, i_10_350_4563_0, i_10_350_4566_0, i_10_350_4568_0,
    o_10_350_0_0  );
  input  i_10_350_27_0, i_10_350_220_0, i_10_350_249_0, i_10_350_282_0,
    i_10_350_284_0, i_10_350_293_0, i_10_350_327_0, i_10_350_412_0,
    i_10_350_428_0, i_10_350_517_0, i_10_350_518_0, i_10_350_520_0,
    i_10_350_798_0, i_10_350_800_0, i_10_350_955_0, i_10_350_957_0,
    i_10_350_961_0, i_10_350_1033_0, i_10_350_1035_0, i_10_350_1152_0,
    i_10_350_1243_0, i_10_350_1245_0, i_10_350_1246_0, i_10_350_1247_0,
    i_10_350_1310_0, i_10_350_1311_0, i_10_350_1384_0, i_10_350_1539_0,
    i_10_350_1617_0, i_10_350_1683_0, i_10_350_1686_0, i_10_350_1690_0,
    i_10_350_1691_0, i_10_350_1820_0, i_10_350_1822_0, i_10_350_1825_0,
    i_10_350_1908_0, i_10_350_1911_0, i_10_350_1912_0, i_10_350_2186_0,
    i_10_350_2349_0, i_10_350_2350_0, i_10_350_2360_0, i_10_350_2361_0,
    i_10_350_2406_0, i_10_350_2452_0, i_10_350_2467_0, i_10_350_2468_0,
    i_10_350_2470_0, i_10_350_2473_0, i_10_350_2655_0, i_10_350_2679_0,
    i_10_350_2719_0, i_10_350_2725_0, i_10_350_2726_0, i_10_350_2740_0,
    i_10_350_2827_0, i_10_350_3036_0, i_10_350_3048_0, i_10_350_3074_0,
    i_10_350_3075_0, i_10_350_3201_0, i_10_350_3269_0, i_10_350_3387_0,
    i_10_350_3391_0, i_10_350_3392_0, i_10_350_3453_0, i_10_350_3520_0,
    i_10_350_3523_0, i_10_350_3609_0, i_10_350_3612_0, i_10_350_3613_0,
    i_10_350_3614_0, i_10_350_3617_0, i_10_350_3624_0, i_10_350_3648_0,
    i_10_350_3651_0, i_10_350_3652_0, i_10_350_3706_0, i_10_350_3723_0,
    i_10_350_3730_0, i_10_350_3780_0, i_10_350_3834_0, i_10_350_3835_0,
    i_10_350_3839_0, i_10_350_3840_0, i_10_350_3860_0, i_10_350_3993_0,
    i_10_350_4114_0, i_10_350_4120_0, i_10_350_4126_0, i_10_350_4215_0,
    i_10_350_4216_0, i_10_350_4219_0, i_10_350_4236_0, i_10_350_4273_0,
    i_10_350_4291_0, i_10_350_4563_0, i_10_350_4566_0, i_10_350_4568_0;
  output o_10_350_0_0;
  assign o_10_350_0_0 = 0;
endmodule



// Benchmark "kernel_10_351" written by ABC on Sun Jul 19 10:27:08 2020

module kernel_10_351 ( 
    i_10_351_131_0, i_10_351_182_0, i_10_351_220_0, i_10_351_307_0,
    i_10_351_350_0, i_10_351_361_0, i_10_351_374_0, i_10_351_388_0,
    i_10_351_433_0, i_10_351_560_0, i_10_351_563_0, i_10_351_566_0,
    i_10_351_716_0, i_10_351_751_0, i_10_351_819_0, i_10_351_907_0,
    i_10_351_931_0, i_10_351_955_0, i_10_351_1046_0, i_10_351_1049_0,
    i_10_351_1084_0, i_10_351_1237_0, i_10_351_1247_0, i_10_351_1305_0,
    i_10_351_1308_0, i_10_351_1309_0, i_10_351_1310_0, i_10_351_1454_0,
    i_10_351_1488_0, i_10_351_1489_0, i_10_351_1543_0, i_10_351_1616_0,
    i_10_351_1648_0, i_10_351_1649_0, i_10_351_1652_0, i_10_351_1654_0,
    i_10_351_1688_0, i_10_351_1689_0, i_10_351_1864_0, i_10_351_2026_0,
    i_10_351_2038_0, i_10_351_2061_0, i_10_351_2080_0, i_10_351_2081_0,
    i_10_351_2201_0, i_10_351_2254_0, i_10_351_2514_0, i_10_351_2515_0,
    i_10_351_2533_0, i_10_351_2610_0, i_10_351_2657_0, i_10_351_2660_0,
    i_10_351_2729_0, i_10_351_2731_0, i_10_351_2740_0, i_10_351_2741_0,
    i_10_351_2830_0, i_10_351_2999_0, i_10_351_3039_0, i_10_351_3070_0,
    i_10_351_3292_0, i_10_351_3388_0, i_10_351_3389_0, i_10_351_3492_0,
    i_10_351_3542_0, i_10_351_3583_0, i_10_351_3587_0, i_10_351_3618_0,
    i_10_351_3646_0, i_10_351_3647_0, i_10_351_3649_0, i_10_351_3650_0,
    i_10_351_3682_0, i_10_351_3788_0, i_10_351_3807_0, i_10_351_3853_0,
    i_10_351_3854_0, i_10_351_3856_0, i_10_351_3857_0, i_10_351_3910_0,
    i_10_351_3911_0, i_10_351_3978_0, i_10_351_3979_0, i_10_351_4051_0,
    i_10_351_4052_0, i_10_351_4054_0, i_10_351_4055_0, i_10_351_4113_0,
    i_10_351_4114_0, i_10_351_4117_0, i_10_351_4191_0, i_10_351_4216_0,
    i_10_351_4311_0, i_10_351_4394_0, i_10_351_4400_0, i_10_351_4451_0,
    i_10_351_4528_0, i_10_351_4529_0, i_10_351_4531_0, i_10_351_4567_0,
    o_10_351_0_0  );
  input  i_10_351_131_0, i_10_351_182_0, i_10_351_220_0, i_10_351_307_0,
    i_10_351_350_0, i_10_351_361_0, i_10_351_374_0, i_10_351_388_0,
    i_10_351_433_0, i_10_351_560_0, i_10_351_563_0, i_10_351_566_0,
    i_10_351_716_0, i_10_351_751_0, i_10_351_819_0, i_10_351_907_0,
    i_10_351_931_0, i_10_351_955_0, i_10_351_1046_0, i_10_351_1049_0,
    i_10_351_1084_0, i_10_351_1237_0, i_10_351_1247_0, i_10_351_1305_0,
    i_10_351_1308_0, i_10_351_1309_0, i_10_351_1310_0, i_10_351_1454_0,
    i_10_351_1488_0, i_10_351_1489_0, i_10_351_1543_0, i_10_351_1616_0,
    i_10_351_1648_0, i_10_351_1649_0, i_10_351_1652_0, i_10_351_1654_0,
    i_10_351_1688_0, i_10_351_1689_0, i_10_351_1864_0, i_10_351_2026_0,
    i_10_351_2038_0, i_10_351_2061_0, i_10_351_2080_0, i_10_351_2081_0,
    i_10_351_2201_0, i_10_351_2254_0, i_10_351_2514_0, i_10_351_2515_0,
    i_10_351_2533_0, i_10_351_2610_0, i_10_351_2657_0, i_10_351_2660_0,
    i_10_351_2729_0, i_10_351_2731_0, i_10_351_2740_0, i_10_351_2741_0,
    i_10_351_2830_0, i_10_351_2999_0, i_10_351_3039_0, i_10_351_3070_0,
    i_10_351_3292_0, i_10_351_3388_0, i_10_351_3389_0, i_10_351_3492_0,
    i_10_351_3542_0, i_10_351_3583_0, i_10_351_3587_0, i_10_351_3618_0,
    i_10_351_3646_0, i_10_351_3647_0, i_10_351_3649_0, i_10_351_3650_0,
    i_10_351_3682_0, i_10_351_3788_0, i_10_351_3807_0, i_10_351_3853_0,
    i_10_351_3854_0, i_10_351_3856_0, i_10_351_3857_0, i_10_351_3910_0,
    i_10_351_3911_0, i_10_351_3978_0, i_10_351_3979_0, i_10_351_4051_0,
    i_10_351_4052_0, i_10_351_4054_0, i_10_351_4055_0, i_10_351_4113_0,
    i_10_351_4114_0, i_10_351_4117_0, i_10_351_4191_0, i_10_351_4216_0,
    i_10_351_4311_0, i_10_351_4394_0, i_10_351_4400_0, i_10_351_4451_0,
    i_10_351_4528_0, i_10_351_4529_0, i_10_351_4531_0, i_10_351_4567_0;
  output o_10_351_0_0;
  assign o_10_351_0_0 = 0;
endmodule



// Benchmark "kernel_10_352" written by ABC on Sun Jul 19 10:27:09 2020

module kernel_10_352 ( 
    i_10_352_281_0, i_10_352_282_0, i_10_352_284_0, i_10_352_293_0,
    i_10_352_320_0, i_10_352_322_0, i_10_352_328_0, i_10_352_329_0,
    i_10_352_405_0, i_10_352_409_0, i_10_352_410_0, i_10_352_412_0,
    i_10_352_436_0, i_10_352_445_0, i_10_352_446_0, i_10_352_448_0,
    i_10_352_466_0, i_10_352_467_0, i_10_352_796_0, i_10_352_959_0,
    i_10_352_960_0, i_10_352_961_0, i_10_352_991_0, i_10_352_992_0,
    i_10_352_994_0, i_10_352_996_0, i_10_352_1233_0, i_10_352_1237_0,
    i_10_352_1263_0, i_10_352_1264_0, i_10_352_1309_0, i_10_352_1348_0,
    i_10_352_1653_0, i_10_352_1769_0, i_10_352_1819_0, i_10_352_1820_0,
    i_10_352_1821_0, i_10_352_1822_0, i_10_352_1876_0, i_10_352_1877_0,
    i_10_352_1912_0, i_10_352_1913_0, i_10_352_1989_0, i_10_352_1990_0,
    i_10_352_2351_0, i_10_352_2352_0, i_10_352_2357_0, i_10_352_2362_0,
    i_10_352_2382_0, i_10_352_2383_0, i_10_352_2456_0, i_10_352_2603_0,
    i_10_352_2634_0, i_10_352_2655_0, i_10_352_2656_0, i_10_352_2657_0,
    i_10_352_2659_0, i_10_352_2663_0, i_10_352_2713_0, i_10_352_2714_0,
    i_10_352_2715_0, i_10_352_2716_0, i_10_352_2717_0, i_10_352_2718_0,
    i_10_352_2719_0, i_10_352_2722_0, i_10_352_2730_0, i_10_352_2819_0,
    i_10_352_2826_0, i_10_352_2827_0, i_10_352_2829_0, i_10_352_2830_0,
    i_10_352_2883_0, i_10_352_2919_0, i_10_352_2923_0, i_10_352_2981_0,
    i_10_352_3034_0, i_10_352_3035_0, i_10_352_3037_0, i_10_352_3070_0,
    i_10_352_3076_0, i_10_352_3094_0, i_10_352_3385_0, i_10_352_3388_0,
    i_10_352_3390_0, i_10_352_3406_0, i_10_352_3407_0, i_10_352_3434_0,
    i_10_352_3520_0, i_10_352_3521_0, i_10_352_3523_0, i_10_352_3610_0,
    i_10_352_3834_0, i_10_352_3835_0, i_10_352_3855_0, i_10_352_3859_0,
    i_10_352_4268_0, i_10_352_4271_0, i_10_352_4277_0, i_10_352_4570_0,
    o_10_352_0_0  );
  input  i_10_352_281_0, i_10_352_282_0, i_10_352_284_0, i_10_352_293_0,
    i_10_352_320_0, i_10_352_322_0, i_10_352_328_0, i_10_352_329_0,
    i_10_352_405_0, i_10_352_409_0, i_10_352_410_0, i_10_352_412_0,
    i_10_352_436_0, i_10_352_445_0, i_10_352_446_0, i_10_352_448_0,
    i_10_352_466_0, i_10_352_467_0, i_10_352_796_0, i_10_352_959_0,
    i_10_352_960_0, i_10_352_961_0, i_10_352_991_0, i_10_352_992_0,
    i_10_352_994_0, i_10_352_996_0, i_10_352_1233_0, i_10_352_1237_0,
    i_10_352_1263_0, i_10_352_1264_0, i_10_352_1309_0, i_10_352_1348_0,
    i_10_352_1653_0, i_10_352_1769_0, i_10_352_1819_0, i_10_352_1820_0,
    i_10_352_1821_0, i_10_352_1822_0, i_10_352_1876_0, i_10_352_1877_0,
    i_10_352_1912_0, i_10_352_1913_0, i_10_352_1989_0, i_10_352_1990_0,
    i_10_352_2351_0, i_10_352_2352_0, i_10_352_2357_0, i_10_352_2362_0,
    i_10_352_2382_0, i_10_352_2383_0, i_10_352_2456_0, i_10_352_2603_0,
    i_10_352_2634_0, i_10_352_2655_0, i_10_352_2656_0, i_10_352_2657_0,
    i_10_352_2659_0, i_10_352_2663_0, i_10_352_2713_0, i_10_352_2714_0,
    i_10_352_2715_0, i_10_352_2716_0, i_10_352_2717_0, i_10_352_2718_0,
    i_10_352_2719_0, i_10_352_2722_0, i_10_352_2730_0, i_10_352_2819_0,
    i_10_352_2826_0, i_10_352_2827_0, i_10_352_2829_0, i_10_352_2830_0,
    i_10_352_2883_0, i_10_352_2919_0, i_10_352_2923_0, i_10_352_2981_0,
    i_10_352_3034_0, i_10_352_3035_0, i_10_352_3037_0, i_10_352_3070_0,
    i_10_352_3076_0, i_10_352_3094_0, i_10_352_3385_0, i_10_352_3388_0,
    i_10_352_3390_0, i_10_352_3406_0, i_10_352_3407_0, i_10_352_3434_0,
    i_10_352_3520_0, i_10_352_3521_0, i_10_352_3523_0, i_10_352_3610_0,
    i_10_352_3834_0, i_10_352_3835_0, i_10_352_3855_0, i_10_352_3859_0,
    i_10_352_4268_0, i_10_352_4271_0, i_10_352_4277_0, i_10_352_4570_0;
  output o_10_352_0_0;
  assign o_10_352_0_0 = ~((~i_10_352_2656_0 & ((~i_10_352_282_0 & ((~i_10_352_293_0 & ~i_10_352_1348_0 & ~i_10_352_2819_0 & ~i_10_352_3834_0 & i_10_352_3859_0) | (~i_10_352_320_0 & ~i_10_352_1912_0 & ~i_10_352_2715_0 & i_10_352_2923_0 & ~i_10_352_2981_0 & ~i_10_352_3523_0 & ~i_10_352_3859_0))) | (~i_10_352_329_0 & ~i_10_352_436_0 & i_10_352_796_0 & ~i_10_352_1348_0 & ~i_10_352_2362_0 & ~i_10_352_2717_0 & ~i_10_352_3407_0) | (~i_10_352_293_0 & ~i_10_352_328_0 & ~i_10_352_991_0 & ~i_10_352_2657_0 & ~i_10_352_2716_0 & ~i_10_352_3520_0))) | (~i_10_352_328_0 & ((~i_10_352_409_0 & ~i_10_352_1348_0 & ~i_10_352_1912_0 & ~i_10_352_1990_0 & i_10_352_2634_0 & ~i_10_352_2819_0 & ~i_10_352_3094_0) | (i_10_352_466_0 & ~i_10_352_991_0 & ~i_10_352_992_0 & ~i_10_352_2716_0 & ~i_10_352_3610_0))) | (~i_10_352_960_0 & ((~i_10_352_796_0 & i_10_352_1309_0 & ~i_10_352_1876_0 & ~i_10_352_2657_0 & ~i_10_352_2830_0 & ~i_10_352_3035_0 & ~i_10_352_3406_0) | (~i_10_352_992_0 & ~i_10_352_996_0 & ~i_10_352_1912_0 & ~i_10_352_1989_0 & ~i_10_352_2362_0 & ~i_10_352_2603_0 & ~i_10_352_2714_0 & ~i_10_352_3076_0 & ~i_10_352_3385_0 & ~i_10_352_3434_0 & ~i_10_352_3521_0))) | (~i_10_352_3390_0 & ((~i_10_352_320_0 & ((~i_10_352_991_0 & ~i_10_352_994_0 & i_10_352_1653_0 & ~i_10_352_3076_0 & ~i_10_352_3407_0) | (~i_10_352_996_0 & ~i_10_352_1769_0 & ~i_10_352_2351_0 & ~i_10_352_2352_0 & ~i_10_352_2659_0 & ~i_10_352_2819_0 & ~i_10_352_3434_0 & ~i_10_352_3521_0 & ~i_10_352_3835_0 & ~i_10_352_3855_0))) | (~i_10_352_992_0 & ((~i_10_352_1263_0 & ~i_10_352_1913_0 & ~i_10_352_2657_0 & ~i_10_352_2659_0 & ~i_10_352_2715_0 & ~i_10_352_2830_0 & ~i_10_352_3076_0) | (~i_10_352_1348_0 & ~i_10_352_2362_0 & ~i_10_352_2717_0 & ~i_10_352_2827_0 & ~i_10_352_3520_0 & ~i_10_352_3521_0))) | (~i_10_352_1989_0 & ~i_10_352_2657_0 & ~i_10_352_2717_0 & i_10_352_2719_0 & ~i_10_352_2883_0 & i_10_352_2923_0))) | (~i_10_352_3523_0 & ((~i_10_352_994_0 & ((i_10_352_991_0 & i_10_352_1819_0) | (~i_10_352_2603_0 & ~i_10_352_2719_0 & ~i_10_352_2829_0 & ~i_10_352_2919_0 & ~i_10_352_3076_0 & ~i_10_352_3388_0 & ~i_10_352_3434_0 & ~i_10_352_3855_0))) | (~i_10_352_2827_0 & i_10_352_3385_0 & ~i_10_352_3388_0 & i_10_352_3855_0))) | (~i_10_352_1348_0 & ~i_10_352_2819_0 & ((~i_10_352_410_0 & ~i_10_352_1769_0 & i_10_352_1819_0 & ~i_10_352_3520_0) | (~i_10_352_281_0 & ~i_10_352_412_0 & ~i_10_352_991_0 & ~i_10_352_1821_0 & ~i_10_352_1990_0 & ~i_10_352_2655_0 & ~i_10_352_2714_0 & ~i_10_352_4271_0))) | (i_10_352_1819_0 & ((i_10_352_1820_0 & ~i_10_352_1821_0 & ~i_10_352_1822_0 & ~i_10_352_1876_0 & ~i_10_352_1912_0 & ~i_10_352_2981_0 & ~i_10_352_3521_0) | (i_10_352_2919_0 & i_10_352_3407_0 & ~i_10_352_3855_0))) | (~i_10_352_1912_0 & ((i_10_352_994_0 & i_10_352_2718_0 & ~i_10_352_2719_0 & i_10_352_2919_0 & i_10_352_3407_0) | (~i_10_352_320_0 & ~i_10_352_991_0 & ~i_10_352_1263_0 & ~i_10_352_1769_0 & ~i_10_352_1877_0 & ~i_10_352_1913_0 & ~i_10_352_2382_0 & ~i_10_352_2826_0 & ~i_10_352_3434_0))) | (~i_10_352_991_0 & ((i_10_352_1822_0 & i_10_352_3385_0 & ~i_10_352_3388_0 & ~i_10_352_3406_0) | (~i_10_352_329_0 & ~i_10_352_405_0 & ~i_10_352_2659_0 & ~i_10_352_2830_0 & ~i_10_352_3070_0 & ~i_10_352_3094_0 & ~i_10_352_3407_0 & i_10_352_3835_0))) | (~i_10_352_284_0 & i_10_352_446_0 & ~i_10_352_1820_0 & ~i_10_352_1876_0 & ~i_10_352_3521_0 & ~i_10_352_4268_0));
endmodule



// Benchmark "kernel_10_353" written by ABC on Sun Jul 19 10:27:10 2020

module kernel_10_353 ( 
    i_10_353_43_0, i_10_353_44_0, i_10_353_49_0, i_10_353_89_0,
    i_10_353_176_0, i_10_353_179_0, i_10_353_224_0, i_10_353_248_0,
    i_10_353_279_0, i_10_353_281_0, i_10_353_282_0, i_10_353_295_0,
    i_10_353_316_0, i_10_353_317_0, i_10_353_319_0, i_10_353_320_0,
    i_10_353_328_0, i_10_353_412_0, i_10_353_413_0, i_10_353_434_0,
    i_10_353_441_0, i_10_353_467_0, i_10_353_643_0, i_10_353_715_0,
    i_10_353_716_0, i_10_353_795_0, i_10_353_796_0, i_10_353_896_0,
    i_10_353_898_0, i_10_353_958_0, i_10_353_997_0, i_10_353_1004_0,
    i_10_353_1236_0, i_10_353_1238_0, i_10_353_1241_0, i_10_353_1244_0,
    i_10_353_1247_0, i_10_353_1261_0, i_10_353_1262_0, i_10_353_1313_0,
    i_10_353_1365_0, i_10_353_1366_0, i_10_353_1645_0, i_10_353_1654_0,
    i_10_353_1687_0, i_10_353_1732_0, i_10_353_1824_0, i_10_353_1994_0,
    i_10_353_1999_0, i_10_353_2002_0, i_10_353_2005_0, i_10_353_2024_0,
    i_10_353_2057_0, i_10_353_2165_0, i_10_353_2351_0, i_10_353_2362_0,
    i_10_353_2363_0, i_10_353_2365_0, i_10_353_2366_0, i_10_353_2377_0,
    i_10_353_2449_0, i_10_353_2467_0, i_10_353_2470_0, i_10_353_2471_0,
    i_10_353_2603_0, i_10_353_2630_0, i_10_353_2675_0, i_10_353_2678_0,
    i_10_353_2680_0, i_10_353_2723_0, i_10_353_2725_0, i_10_353_2785_0,
    i_10_353_2786_0, i_10_353_2884_0, i_10_353_2981_0, i_10_353_3074_0,
    i_10_353_3077_0, i_10_353_3272_0, i_10_353_3613_0, i_10_353_3616_0,
    i_10_353_3617_0, i_10_353_3721_0, i_10_353_3722_0, i_10_353_3809_0,
    i_10_353_3841_0, i_10_353_3853_0, i_10_353_3875_0, i_10_353_3911_0,
    i_10_353_3949_0, i_10_353_3993_0, i_10_353_3994_0, i_10_353_3995_0,
    i_10_353_4115_0, i_10_353_4117_0, i_10_353_4120_0, i_10_353_4121_0,
    i_10_353_4130_0, i_10_353_4175_0, i_10_353_4220_0, i_10_353_4276_0,
    o_10_353_0_0  );
  input  i_10_353_43_0, i_10_353_44_0, i_10_353_49_0, i_10_353_89_0,
    i_10_353_176_0, i_10_353_179_0, i_10_353_224_0, i_10_353_248_0,
    i_10_353_279_0, i_10_353_281_0, i_10_353_282_0, i_10_353_295_0,
    i_10_353_316_0, i_10_353_317_0, i_10_353_319_0, i_10_353_320_0,
    i_10_353_328_0, i_10_353_412_0, i_10_353_413_0, i_10_353_434_0,
    i_10_353_441_0, i_10_353_467_0, i_10_353_643_0, i_10_353_715_0,
    i_10_353_716_0, i_10_353_795_0, i_10_353_796_0, i_10_353_896_0,
    i_10_353_898_0, i_10_353_958_0, i_10_353_997_0, i_10_353_1004_0,
    i_10_353_1236_0, i_10_353_1238_0, i_10_353_1241_0, i_10_353_1244_0,
    i_10_353_1247_0, i_10_353_1261_0, i_10_353_1262_0, i_10_353_1313_0,
    i_10_353_1365_0, i_10_353_1366_0, i_10_353_1645_0, i_10_353_1654_0,
    i_10_353_1687_0, i_10_353_1732_0, i_10_353_1824_0, i_10_353_1994_0,
    i_10_353_1999_0, i_10_353_2002_0, i_10_353_2005_0, i_10_353_2024_0,
    i_10_353_2057_0, i_10_353_2165_0, i_10_353_2351_0, i_10_353_2362_0,
    i_10_353_2363_0, i_10_353_2365_0, i_10_353_2366_0, i_10_353_2377_0,
    i_10_353_2449_0, i_10_353_2467_0, i_10_353_2470_0, i_10_353_2471_0,
    i_10_353_2603_0, i_10_353_2630_0, i_10_353_2675_0, i_10_353_2678_0,
    i_10_353_2680_0, i_10_353_2723_0, i_10_353_2725_0, i_10_353_2785_0,
    i_10_353_2786_0, i_10_353_2884_0, i_10_353_2981_0, i_10_353_3074_0,
    i_10_353_3077_0, i_10_353_3272_0, i_10_353_3613_0, i_10_353_3616_0,
    i_10_353_3617_0, i_10_353_3721_0, i_10_353_3722_0, i_10_353_3809_0,
    i_10_353_3841_0, i_10_353_3853_0, i_10_353_3875_0, i_10_353_3911_0,
    i_10_353_3949_0, i_10_353_3993_0, i_10_353_3994_0, i_10_353_3995_0,
    i_10_353_4115_0, i_10_353_4117_0, i_10_353_4120_0, i_10_353_4121_0,
    i_10_353_4130_0, i_10_353_4175_0, i_10_353_4220_0, i_10_353_4276_0;
  output o_10_353_0_0;
  assign o_10_353_0_0 = 0;
endmodule



// Benchmark "kernel_10_354" written by ABC on Sun Jul 19 10:27:11 2020

module kernel_10_354 ( 
    i_10_354_83_0, i_10_354_89_0, i_10_354_172_0, i_10_354_177_0,
    i_10_354_187_0, i_10_354_188_0, i_10_354_214_0, i_10_354_224_0,
    i_10_354_283_0, i_10_354_284_0, i_10_354_318_0, i_10_354_371_0,
    i_10_354_406_0, i_10_354_410_0, i_10_354_413_0, i_10_354_446_0,
    i_10_354_799_0, i_10_354_800_0, i_10_354_906_0, i_10_354_907_0,
    i_10_354_908_0, i_10_354_919_0, i_10_354_920_0, i_10_354_1237_0,
    i_10_354_1238_0, i_10_354_1239_0, i_10_354_1240_0, i_10_354_1245_0,
    i_10_354_1249_0, i_10_354_1250_0, i_10_354_1367_0, i_10_354_1618_0,
    i_10_354_1651_0, i_10_354_1686_0, i_10_354_1687_0, i_10_354_1688_0,
    i_10_354_1767_0, i_10_354_1768_0, i_10_354_1802_0, i_10_354_1888_0,
    i_10_354_1907_0, i_10_354_1909_0, i_10_354_1912_0, i_10_354_1914_0,
    i_10_354_1940_0, i_10_354_1951_0, i_10_354_1952_0, i_10_354_1960_0,
    i_10_354_2020_0, i_10_354_2312_0, i_10_354_2452_0, i_10_354_2455_0,
    i_10_354_2462_0, i_10_354_2463_0, i_10_354_2464_0, i_10_354_2509_0,
    i_10_354_2629_0, i_10_354_2632_0, i_10_354_2634_0, i_10_354_2707_0,
    i_10_354_2708_0, i_10_354_2730_0, i_10_354_2732_0, i_10_354_2758_0,
    i_10_354_2783_0, i_10_354_2922_0, i_10_354_2924_0, i_10_354_3011_0,
    i_10_354_3014_0, i_10_354_3038_0, i_10_354_3185_0, i_10_354_3198_0,
    i_10_354_3199_0, i_10_354_3320_0, i_10_354_3387_0, i_10_354_3613_0,
    i_10_354_3614_0, i_10_354_3689_0, i_10_354_3707_0, i_10_354_3839_0,
    i_10_354_3857_0, i_10_354_3884_0, i_10_354_3887_0, i_10_354_3895_0,
    i_10_354_3967_0, i_10_354_3982_0, i_10_354_4183_0, i_10_354_4184_0,
    i_10_354_4193_0, i_10_354_4270_0, i_10_354_4272_0, i_10_354_4273_0,
    i_10_354_4274_0, i_10_354_4279_0, i_10_354_4298_0, i_10_354_4534_0,
    i_10_354_4567_0, i_10_354_4568_0, i_10_354_4606_0, i_10_354_4607_0,
    o_10_354_0_0  );
  input  i_10_354_83_0, i_10_354_89_0, i_10_354_172_0, i_10_354_177_0,
    i_10_354_187_0, i_10_354_188_0, i_10_354_214_0, i_10_354_224_0,
    i_10_354_283_0, i_10_354_284_0, i_10_354_318_0, i_10_354_371_0,
    i_10_354_406_0, i_10_354_410_0, i_10_354_413_0, i_10_354_446_0,
    i_10_354_799_0, i_10_354_800_0, i_10_354_906_0, i_10_354_907_0,
    i_10_354_908_0, i_10_354_919_0, i_10_354_920_0, i_10_354_1237_0,
    i_10_354_1238_0, i_10_354_1239_0, i_10_354_1240_0, i_10_354_1245_0,
    i_10_354_1249_0, i_10_354_1250_0, i_10_354_1367_0, i_10_354_1618_0,
    i_10_354_1651_0, i_10_354_1686_0, i_10_354_1687_0, i_10_354_1688_0,
    i_10_354_1767_0, i_10_354_1768_0, i_10_354_1802_0, i_10_354_1888_0,
    i_10_354_1907_0, i_10_354_1909_0, i_10_354_1912_0, i_10_354_1914_0,
    i_10_354_1940_0, i_10_354_1951_0, i_10_354_1952_0, i_10_354_1960_0,
    i_10_354_2020_0, i_10_354_2312_0, i_10_354_2452_0, i_10_354_2455_0,
    i_10_354_2462_0, i_10_354_2463_0, i_10_354_2464_0, i_10_354_2509_0,
    i_10_354_2629_0, i_10_354_2632_0, i_10_354_2634_0, i_10_354_2707_0,
    i_10_354_2708_0, i_10_354_2730_0, i_10_354_2732_0, i_10_354_2758_0,
    i_10_354_2783_0, i_10_354_2922_0, i_10_354_2924_0, i_10_354_3011_0,
    i_10_354_3014_0, i_10_354_3038_0, i_10_354_3185_0, i_10_354_3198_0,
    i_10_354_3199_0, i_10_354_3320_0, i_10_354_3387_0, i_10_354_3613_0,
    i_10_354_3614_0, i_10_354_3689_0, i_10_354_3707_0, i_10_354_3839_0,
    i_10_354_3857_0, i_10_354_3884_0, i_10_354_3887_0, i_10_354_3895_0,
    i_10_354_3967_0, i_10_354_3982_0, i_10_354_4183_0, i_10_354_4184_0,
    i_10_354_4193_0, i_10_354_4270_0, i_10_354_4272_0, i_10_354_4273_0,
    i_10_354_4274_0, i_10_354_4279_0, i_10_354_4298_0, i_10_354_4534_0,
    i_10_354_4567_0, i_10_354_4568_0, i_10_354_4606_0, i_10_354_4607_0;
  output o_10_354_0_0;
  assign o_10_354_0_0 = 0;
endmodule



// Benchmark "kernel_10_355" written by ABC on Sun Jul 19 10:27:12 2020

module kernel_10_355 ( 
    i_10_355_27_0, i_10_355_48_0, i_10_355_49_0, i_10_355_130_0,
    i_10_355_144_0, i_10_355_145_0, i_10_355_172_0, i_10_355_176_0,
    i_10_355_283_0, i_10_355_324_0, i_10_355_495_0, i_10_355_513_0,
    i_10_355_586_0, i_10_355_587_0, i_10_355_623_0, i_10_355_711_0,
    i_10_355_733_0, i_10_355_792_0, i_10_355_795_0, i_10_355_821_0,
    i_10_355_918_0, i_10_355_963_0, i_10_355_981_0, i_10_355_999_0,
    i_10_355_1027_0, i_10_355_1044_0, i_10_355_1081_0, i_10_355_1161_0,
    i_10_355_1215_0, i_10_355_1216_0, i_10_355_1218_0, i_10_355_1236_0,
    i_10_355_1237_0, i_10_355_1280_0, i_10_355_1446_0, i_10_355_1476_0,
    i_10_355_1477_0, i_10_355_1478_0, i_10_355_1548_0, i_10_355_1617_0,
    i_10_355_1639_0, i_10_355_1764_0, i_10_355_1812_0, i_10_355_1822_0,
    i_10_355_1911_0, i_10_355_1915_0, i_10_355_1953_0, i_10_355_1956_0,
    i_10_355_1990_0, i_10_355_1998_0, i_10_355_2089_0, i_10_355_2179_0,
    i_10_355_2180_0, i_10_355_2199_0, i_10_355_2201_0, i_10_355_2304_0,
    i_10_355_2410_0, i_10_355_2485_0, i_10_355_2493_0, i_10_355_2631_0,
    i_10_355_2659_0, i_10_355_2662_0, i_10_355_2688_0, i_10_355_2922_0,
    i_10_355_2955_0, i_10_355_2981_0, i_10_355_3070_0, i_10_355_3097_0,
    i_10_355_3114_0, i_10_355_3115_0, i_10_355_3277_0, i_10_355_3278_0,
    i_10_355_3312_0, i_10_355_3331_0, i_10_355_3348_0, i_10_355_3439_0,
    i_10_355_3492_0, i_10_355_3493_0, i_10_355_3539_0, i_10_355_3589_0,
    i_10_355_3645_0, i_10_355_3646_0, i_10_355_3794_0, i_10_355_3871_0,
    i_10_355_3879_0, i_10_355_3997_0, i_10_355_4007_0, i_10_355_4059_0,
    i_10_355_4060_0, i_10_355_4063_0, i_10_355_4114_0, i_10_355_4126_0,
    i_10_355_4267_0, i_10_355_4286_0, i_10_355_4293_0, i_10_355_4294_0,
    i_10_355_4311_0, i_10_355_4314_0, i_10_355_4581_0, i_10_355_4582_0,
    o_10_355_0_0  );
  input  i_10_355_27_0, i_10_355_48_0, i_10_355_49_0, i_10_355_130_0,
    i_10_355_144_0, i_10_355_145_0, i_10_355_172_0, i_10_355_176_0,
    i_10_355_283_0, i_10_355_324_0, i_10_355_495_0, i_10_355_513_0,
    i_10_355_586_0, i_10_355_587_0, i_10_355_623_0, i_10_355_711_0,
    i_10_355_733_0, i_10_355_792_0, i_10_355_795_0, i_10_355_821_0,
    i_10_355_918_0, i_10_355_963_0, i_10_355_981_0, i_10_355_999_0,
    i_10_355_1027_0, i_10_355_1044_0, i_10_355_1081_0, i_10_355_1161_0,
    i_10_355_1215_0, i_10_355_1216_0, i_10_355_1218_0, i_10_355_1236_0,
    i_10_355_1237_0, i_10_355_1280_0, i_10_355_1446_0, i_10_355_1476_0,
    i_10_355_1477_0, i_10_355_1478_0, i_10_355_1548_0, i_10_355_1617_0,
    i_10_355_1639_0, i_10_355_1764_0, i_10_355_1812_0, i_10_355_1822_0,
    i_10_355_1911_0, i_10_355_1915_0, i_10_355_1953_0, i_10_355_1956_0,
    i_10_355_1990_0, i_10_355_1998_0, i_10_355_2089_0, i_10_355_2179_0,
    i_10_355_2180_0, i_10_355_2199_0, i_10_355_2201_0, i_10_355_2304_0,
    i_10_355_2410_0, i_10_355_2485_0, i_10_355_2493_0, i_10_355_2631_0,
    i_10_355_2659_0, i_10_355_2662_0, i_10_355_2688_0, i_10_355_2922_0,
    i_10_355_2955_0, i_10_355_2981_0, i_10_355_3070_0, i_10_355_3097_0,
    i_10_355_3114_0, i_10_355_3115_0, i_10_355_3277_0, i_10_355_3278_0,
    i_10_355_3312_0, i_10_355_3331_0, i_10_355_3348_0, i_10_355_3439_0,
    i_10_355_3492_0, i_10_355_3493_0, i_10_355_3539_0, i_10_355_3589_0,
    i_10_355_3645_0, i_10_355_3646_0, i_10_355_3794_0, i_10_355_3871_0,
    i_10_355_3879_0, i_10_355_3997_0, i_10_355_4007_0, i_10_355_4059_0,
    i_10_355_4060_0, i_10_355_4063_0, i_10_355_4114_0, i_10_355_4126_0,
    i_10_355_4267_0, i_10_355_4286_0, i_10_355_4293_0, i_10_355_4294_0,
    i_10_355_4311_0, i_10_355_4314_0, i_10_355_4581_0, i_10_355_4582_0;
  output o_10_355_0_0;
  assign o_10_355_0_0 = 0;
endmodule



// Benchmark "kernel_10_356" written by ABC on Sun Jul 19 10:27:13 2020

module kernel_10_356 ( 
    i_10_356_122_0, i_10_356_124_0, i_10_356_175_0, i_10_356_220_0,
    i_10_356_246_0, i_10_356_248_0, i_10_356_319_0, i_10_356_423_0,
    i_10_356_426_0, i_10_356_427_0, i_10_356_442_0, i_10_356_445_0,
    i_10_356_459_0, i_10_356_460_0, i_10_356_461_0, i_10_356_463_0,
    i_10_356_464_0, i_10_356_466_0, i_10_356_795_0, i_10_356_800_0,
    i_10_356_896_0, i_10_356_956_0, i_10_356_959_0, i_10_356_1030_0,
    i_10_356_1233_0, i_10_356_1234_0, i_10_356_1241_0, i_10_356_1312_0,
    i_10_356_1362_0, i_10_356_1379_0, i_10_356_1381_0, i_10_356_1445_0,
    i_10_356_1541_0, i_10_356_1551_0, i_10_356_1552_0, i_10_356_1579_0,
    i_10_356_1583_0, i_10_356_1654_0, i_10_356_1690_0, i_10_356_1825_0,
    i_10_356_1826_0, i_10_356_1909_0, i_10_356_1948_0, i_10_356_2203_0,
    i_10_356_2350_0, i_10_356_2351_0, i_10_356_2353_0, i_10_356_2360_0,
    i_10_356_2377_0, i_10_356_2452_0, i_10_356_2459_0, i_10_356_2467_0,
    i_10_356_2471_0, i_10_356_2629_0, i_10_356_2660_0, i_10_356_2661_0,
    i_10_356_2710_0, i_10_356_2713_0, i_10_356_2721_0, i_10_356_2725_0,
    i_10_356_2728_0, i_10_356_2731_0, i_10_356_2830_0, i_10_356_2831_0,
    i_10_356_2917_0, i_10_356_3037_0, i_10_356_3038_0, i_10_356_3046_0,
    i_10_356_3075_0, i_10_356_3196_0, i_10_356_3199_0, i_10_356_3202_0,
    i_10_356_3270_0, i_10_356_3271_0, i_10_356_3272_0, i_10_356_3281_0,
    i_10_356_3387_0, i_10_356_3388_0, i_10_356_3467_0, i_10_356_3493_0,
    i_10_356_3611_0, i_10_356_3613_0, i_10_356_3647_0, i_10_356_3650_0,
    i_10_356_3781_0, i_10_356_3785_0, i_10_356_3835_0, i_10_356_3837_0,
    i_10_356_3838_0, i_10_356_3844_0, i_10_356_3845_0, i_10_356_3846_0,
    i_10_356_3853_0, i_10_356_3855_0, i_10_356_3880_0, i_10_356_4121_0,
    i_10_356_4267_0, i_10_356_4269_0, i_10_356_4279_0, i_10_356_4286_0,
    o_10_356_0_0  );
  input  i_10_356_122_0, i_10_356_124_0, i_10_356_175_0, i_10_356_220_0,
    i_10_356_246_0, i_10_356_248_0, i_10_356_319_0, i_10_356_423_0,
    i_10_356_426_0, i_10_356_427_0, i_10_356_442_0, i_10_356_445_0,
    i_10_356_459_0, i_10_356_460_0, i_10_356_461_0, i_10_356_463_0,
    i_10_356_464_0, i_10_356_466_0, i_10_356_795_0, i_10_356_800_0,
    i_10_356_896_0, i_10_356_956_0, i_10_356_959_0, i_10_356_1030_0,
    i_10_356_1233_0, i_10_356_1234_0, i_10_356_1241_0, i_10_356_1312_0,
    i_10_356_1362_0, i_10_356_1379_0, i_10_356_1381_0, i_10_356_1445_0,
    i_10_356_1541_0, i_10_356_1551_0, i_10_356_1552_0, i_10_356_1579_0,
    i_10_356_1583_0, i_10_356_1654_0, i_10_356_1690_0, i_10_356_1825_0,
    i_10_356_1826_0, i_10_356_1909_0, i_10_356_1948_0, i_10_356_2203_0,
    i_10_356_2350_0, i_10_356_2351_0, i_10_356_2353_0, i_10_356_2360_0,
    i_10_356_2377_0, i_10_356_2452_0, i_10_356_2459_0, i_10_356_2467_0,
    i_10_356_2471_0, i_10_356_2629_0, i_10_356_2660_0, i_10_356_2661_0,
    i_10_356_2710_0, i_10_356_2713_0, i_10_356_2721_0, i_10_356_2725_0,
    i_10_356_2728_0, i_10_356_2731_0, i_10_356_2830_0, i_10_356_2831_0,
    i_10_356_2917_0, i_10_356_3037_0, i_10_356_3038_0, i_10_356_3046_0,
    i_10_356_3075_0, i_10_356_3196_0, i_10_356_3199_0, i_10_356_3202_0,
    i_10_356_3270_0, i_10_356_3271_0, i_10_356_3272_0, i_10_356_3281_0,
    i_10_356_3387_0, i_10_356_3388_0, i_10_356_3467_0, i_10_356_3493_0,
    i_10_356_3611_0, i_10_356_3613_0, i_10_356_3647_0, i_10_356_3650_0,
    i_10_356_3781_0, i_10_356_3785_0, i_10_356_3835_0, i_10_356_3837_0,
    i_10_356_3838_0, i_10_356_3844_0, i_10_356_3845_0, i_10_356_3846_0,
    i_10_356_3853_0, i_10_356_3855_0, i_10_356_3880_0, i_10_356_4121_0,
    i_10_356_4267_0, i_10_356_4269_0, i_10_356_4279_0, i_10_356_4286_0;
  output o_10_356_0_0;
  assign o_10_356_0_0 = 0;
endmodule



// Benchmark "kernel_10_357" written by ABC on Sun Jul 19 10:27:14 2020

module kernel_10_357 ( 
    i_10_357_145_0, i_10_357_151_0, i_10_357_178_0, i_10_357_179_0,
    i_10_357_186_0, i_10_357_284_0, i_10_357_285_0, i_10_357_443_0,
    i_10_357_445_0, i_10_357_446_0, i_10_357_449_0, i_10_357_465_0,
    i_10_357_466_0, i_10_357_519_0, i_10_357_520_0, i_10_357_719_0,
    i_10_357_755_0, i_10_357_793_0, i_10_357_798_0, i_10_357_799_0,
    i_10_357_966_0, i_10_357_967_0, i_10_357_971_0, i_10_357_997_0,
    i_10_357_1026_0, i_10_357_1166_0, i_10_357_1242_0, i_10_357_1246_0,
    i_10_357_1247_0, i_10_357_1250_0, i_10_357_1308_0, i_10_357_1309_0,
    i_10_357_1363_0, i_10_357_1537_0, i_10_357_1543_0, i_10_357_1580_0,
    i_10_357_1582_0, i_10_357_1583_0, i_10_357_1613_0, i_10_357_1616_0,
    i_10_357_1617_0, i_10_357_1686_0, i_10_357_1819_0, i_10_357_2004_0,
    i_10_357_2005_0, i_10_357_2248_0, i_10_357_2359_0, i_10_357_2361_0,
    i_10_357_2456_0, i_10_357_2607_0, i_10_357_2634_0, i_10_357_2635_0,
    i_10_357_2637_0, i_10_357_2638_0, i_10_357_2660_0, i_10_357_2701_0,
    i_10_357_2703_0, i_10_357_2704_0, i_10_357_2705_0, i_10_357_2718_0,
    i_10_357_2719_0, i_10_357_2725_0, i_10_357_2727_0, i_10_357_2729_0,
    i_10_357_2923_0, i_10_357_3039_0, i_10_357_3041_0, i_10_357_3198_0,
    i_10_357_3199_0, i_10_357_3200_0, i_10_357_3276_0, i_10_357_3277_0,
    i_10_357_3278_0, i_10_357_3392_0, i_10_357_3410_0, i_10_357_3493_0,
    i_10_357_3617_0, i_10_357_3721_0, i_10_357_3783_0, i_10_357_3785_0,
    i_10_357_3788_0, i_10_357_3848_0, i_10_357_3856_0, i_10_357_3857_0,
    i_10_357_3899_0, i_10_357_3913_0, i_10_357_3914_0, i_10_357_4027_0,
    i_10_357_4087_0, i_10_357_4117_0, i_10_357_4118_0, i_10_357_4119_0,
    i_10_357_4121_0, i_10_357_4150_0, i_10_357_4267_0, i_10_357_4269_0,
    i_10_357_4273_0, i_10_357_4289_0, i_10_357_4462_0, i_10_357_4527_0,
    o_10_357_0_0  );
  input  i_10_357_145_0, i_10_357_151_0, i_10_357_178_0, i_10_357_179_0,
    i_10_357_186_0, i_10_357_284_0, i_10_357_285_0, i_10_357_443_0,
    i_10_357_445_0, i_10_357_446_0, i_10_357_449_0, i_10_357_465_0,
    i_10_357_466_0, i_10_357_519_0, i_10_357_520_0, i_10_357_719_0,
    i_10_357_755_0, i_10_357_793_0, i_10_357_798_0, i_10_357_799_0,
    i_10_357_966_0, i_10_357_967_0, i_10_357_971_0, i_10_357_997_0,
    i_10_357_1026_0, i_10_357_1166_0, i_10_357_1242_0, i_10_357_1246_0,
    i_10_357_1247_0, i_10_357_1250_0, i_10_357_1308_0, i_10_357_1309_0,
    i_10_357_1363_0, i_10_357_1537_0, i_10_357_1543_0, i_10_357_1580_0,
    i_10_357_1582_0, i_10_357_1583_0, i_10_357_1613_0, i_10_357_1616_0,
    i_10_357_1617_0, i_10_357_1686_0, i_10_357_1819_0, i_10_357_2004_0,
    i_10_357_2005_0, i_10_357_2248_0, i_10_357_2359_0, i_10_357_2361_0,
    i_10_357_2456_0, i_10_357_2607_0, i_10_357_2634_0, i_10_357_2635_0,
    i_10_357_2637_0, i_10_357_2638_0, i_10_357_2660_0, i_10_357_2701_0,
    i_10_357_2703_0, i_10_357_2704_0, i_10_357_2705_0, i_10_357_2718_0,
    i_10_357_2719_0, i_10_357_2725_0, i_10_357_2727_0, i_10_357_2729_0,
    i_10_357_2923_0, i_10_357_3039_0, i_10_357_3041_0, i_10_357_3198_0,
    i_10_357_3199_0, i_10_357_3200_0, i_10_357_3276_0, i_10_357_3277_0,
    i_10_357_3278_0, i_10_357_3392_0, i_10_357_3410_0, i_10_357_3493_0,
    i_10_357_3617_0, i_10_357_3721_0, i_10_357_3783_0, i_10_357_3785_0,
    i_10_357_3788_0, i_10_357_3848_0, i_10_357_3856_0, i_10_357_3857_0,
    i_10_357_3899_0, i_10_357_3913_0, i_10_357_3914_0, i_10_357_4027_0,
    i_10_357_4087_0, i_10_357_4117_0, i_10_357_4118_0, i_10_357_4119_0,
    i_10_357_4121_0, i_10_357_4150_0, i_10_357_4267_0, i_10_357_4269_0,
    i_10_357_4273_0, i_10_357_4289_0, i_10_357_4462_0, i_10_357_4527_0;
  output o_10_357_0_0;
  assign o_10_357_0_0 = 0;
endmodule



// Benchmark "kernel_10_358" written by ABC on Sun Jul 19 10:27:15 2020

module kernel_10_358 ( 
    i_10_358_66_0, i_10_358_119_0, i_10_358_121_0, i_10_358_175_0,
    i_10_358_181_0, i_10_358_287_0, i_10_358_316_0, i_10_358_346_0,
    i_10_358_432_0, i_10_358_433_0, i_10_358_443_0, i_10_358_446_0,
    i_10_358_515_0, i_10_358_535_0, i_10_358_800_0, i_10_358_909_0,
    i_10_358_957_0, i_10_358_959_0, i_10_358_1008_0, i_10_358_1048_0,
    i_10_358_1055_0, i_10_358_1119_0, i_10_358_1187_0, i_10_358_1234_0,
    i_10_358_1288_0, i_10_358_1305_0, i_10_358_1361_0, i_10_358_1363_0,
    i_10_358_1364_0, i_10_358_1371_0, i_10_358_1447_0, i_10_358_1495_0,
    i_10_358_1581_0, i_10_358_1607_0, i_10_358_1746_0, i_10_358_1882_0,
    i_10_358_1949_0, i_10_358_1955_0, i_10_358_1979_0, i_10_358_2200_0,
    i_10_358_2308_0, i_10_358_2309_0, i_10_358_2354_0, i_10_358_2365_0,
    i_10_358_2458_0, i_10_358_2464_0, i_10_358_2476_0, i_10_358_2565_0,
    i_10_358_2566_0, i_10_358_2610_0, i_10_358_2641_0, i_10_358_2673_0,
    i_10_358_2677_0, i_10_358_2710_0, i_10_358_2711_0, i_10_358_2729_0,
    i_10_358_2731_0, i_10_358_2782_0, i_10_358_3008_0, i_10_358_3037_0,
    i_10_358_3043_0, i_10_358_3088_0, i_10_358_3202_0, i_10_358_3211_0,
    i_10_358_3222_0, i_10_358_3226_0, i_10_358_3238_0, i_10_358_3239_0,
    i_10_358_3267_0, i_10_358_3268_0, i_10_358_3291_0, i_10_358_3319_0,
    i_10_358_3350_0, i_10_358_3384_0, i_10_358_3447_0, i_10_358_3448_0,
    i_10_358_3549_0, i_10_358_3550_0, i_10_358_3551_0, i_10_358_3681_0,
    i_10_358_3686_0, i_10_358_3775_0, i_10_358_3835_0, i_10_358_3837_0,
    i_10_358_3879_0, i_10_358_3919_0, i_10_358_3980_0, i_10_358_3987_0,
    i_10_358_4052_0, i_10_358_4213_0, i_10_358_4232_0, i_10_358_4286_0,
    i_10_358_4306_0, i_10_358_4366_0, i_10_358_4369_0, i_10_358_4370_0,
    i_10_358_4455_0, i_10_358_4460_0, i_10_358_4563_0, i_10_358_4564_0,
    o_10_358_0_0  );
  input  i_10_358_66_0, i_10_358_119_0, i_10_358_121_0, i_10_358_175_0,
    i_10_358_181_0, i_10_358_287_0, i_10_358_316_0, i_10_358_346_0,
    i_10_358_432_0, i_10_358_433_0, i_10_358_443_0, i_10_358_446_0,
    i_10_358_515_0, i_10_358_535_0, i_10_358_800_0, i_10_358_909_0,
    i_10_358_957_0, i_10_358_959_0, i_10_358_1008_0, i_10_358_1048_0,
    i_10_358_1055_0, i_10_358_1119_0, i_10_358_1187_0, i_10_358_1234_0,
    i_10_358_1288_0, i_10_358_1305_0, i_10_358_1361_0, i_10_358_1363_0,
    i_10_358_1364_0, i_10_358_1371_0, i_10_358_1447_0, i_10_358_1495_0,
    i_10_358_1581_0, i_10_358_1607_0, i_10_358_1746_0, i_10_358_1882_0,
    i_10_358_1949_0, i_10_358_1955_0, i_10_358_1979_0, i_10_358_2200_0,
    i_10_358_2308_0, i_10_358_2309_0, i_10_358_2354_0, i_10_358_2365_0,
    i_10_358_2458_0, i_10_358_2464_0, i_10_358_2476_0, i_10_358_2565_0,
    i_10_358_2566_0, i_10_358_2610_0, i_10_358_2641_0, i_10_358_2673_0,
    i_10_358_2677_0, i_10_358_2710_0, i_10_358_2711_0, i_10_358_2729_0,
    i_10_358_2731_0, i_10_358_2782_0, i_10_358_3008_0, i_10_358_3037_0,
    i_10_358_3043_0, i_10_358_3088_0, i_10_358_3202_0, i_10_358_3211_0,
    i_10_358_3222_0, i_10_358_3226_0, i_10_358_3238_0, i_10_358_3239_0,
    i_10_358_3267_0, i_10_358_3268_0, i_10_358_3291_0, i_10_358_3319_0,
    i_10_358_3350_0, i_10_358_3384_0, i_10_358_3447_0, i_10_358_3448_0,
    i_10_358_3549_0, i_10_358_3550_0, i_10_358_3551_0, i_10_358_3681_0,
    i_10_358_3686_0, i_10_358_3775_0, i_10_358_3835_0, i_10_358_3837_0,
    i_10_358_3879_0, i_10_358_3919_0, i_10_358_3980_0, i_10_358_3987_0,
    i_10_358_4052_0, i_10_358_4213_0, i_10_358_4232_0, i_10_358_4286_0,
    i_10_358_4306_0, i_10_358_4366_0, i_10_358_4369_0, i_10_358_4370_0,
    i_10_358_4455_0, i_10_358_4460_0, i_10_358_4563_0, i_10_358_4564_0;
  output o_10_358_0_0;
  assign o_10_358_0_0 = 0;
endmodule



// Benchmark "kernel_10_359" written by ABC on Sun Jul 19 10:27:16 2020

module kernel_10_359 ( 
    i_10_359_173_0, i_10_359_196_0, i_10_359_280_0, i_10_359_315_0,
    i_10_359_388_0, i_10_359_394_0, i_10_359_395_0, i_10_359_437_0,
    i_10_359_513_0, i_10_359_722_0, i_10_359_854_0, i_10_359_948_0,
    i_10_359_949_0, i_10_359_964_0, i_10_359_965_0, i_10_359_1035_0,
    i_10_359_1036_0, i_10_359_1112_0, i_10_359_1121_0, i_10_359_1131_0,
    i_10_359_1237_0, i_10_359_1308_0, i_10_359_1309_0, i_10_359_1353_0,
    i_10_359_1354_0, i_10_359_1357_0, i_10_359_1363_0, i_10_359_1435_0,
    i_10_359_1438_0, i_10_359_1579_0, i_10_359_1650_0, i_10_359_1652_0,
    i_10_359_1653_0, i_10_359_1820_0, i_10_359_1909_0, i_10_359_1912_0,
    i_10_359_1929_0, i_10_359_1947_0, i_10_359_1950_0, i_10_359_1984_0,
    i_10_359_1985_0, i_10_359_2016_0, i_10_359_2209_0, i_10_359_2351_0,
    i_10_359_2512_0, i_10_359_2651_0, i_10_359_2656_0, i_10_359_2657_0,
    i_10_359_2659_0, i_10_359_2695_0, i_10_359_2709_0, i_10_359_2710_0,
    i_10_359_2732_0, i_10_359_2754_0, i_10_359_2826_0, i_10_359_2828_0,
    i_10_359_2831_0, i_10_359_2832_0, i_10_359_2840_0, i_10_359_2880_0,
    i_10_359_2916_0, i_10_359_2918_0, i_10_359_2919_0, i_10_359_2920_0,
    i_10_359_2921_0, i_10_359_2922_0, i_10_359_3046_0, i_10_359_3087_0,
    i_10_359_3090_0, i_10_359_3235_0, i_10_359_3269_0, i_10_359_3272_0,
    i_10_359_3313_0, i_10_359_3315_0, i_10_359_3321_0, i_10_359_3356_0,
    i_10_359_3432_0, i_10_359_3538_0, i_10_359_3585_0, i_10_359_3610_0,
    i_10_359_3651_0, i_10_359_3652_0, i_10_359_3664_0, i_10_359_3699_0,
    i_10_359_3718_0, i_10_359_3775_0, i_10_359_3786_0, i_10_359_3811_0,
    i_10_359_3901_0, i_10_359_3981_0, i_10_359_3982_0, i_10_359_3984_0,
    i_10_359_4091_0, i_10_359_4118_0, i_10_359_4268_0, i_10_359_4285_0,
    i_10_359_4288_0, i_10_359_4290_0, i_10_359_4291_0, i_10_359_4593_0,
    o_10_359_0_0  );
  input  i_10_359_173_0, i_10_359_196_0, i_10_359_280_0, i_10_359_315_0,
    i_10_359_388_0, i_10_359_394_0, i_10_359_395_0, i_10_359_437_0,
    i_10_359_513_0, i_10_359_722_0, i_10_359_854_0, i_10_359_948_0,
    i_10_359_949_0, i_10_359_964_0, i_10_359_965_0, i_10_359_1035_0,
    i_10_359_1036_0, i_10_359_1112_0, i_10_359_1121_0, i_10_359_1131_0,
    i_10_359_1237_0, i_10_359_1308_0, i_10_359_1309_0, i_10_359_1353_0,
    i_10_359_1354_0, i_10_359_1357_0, i_10_359_1363_0, i_10_359_1435_0,
    i_10_359_1438_0, i_10_359_1579_0, i_10_359_1650_0, i_10_359_1652_0,
    i_10_359_1653_0, i_10_359_1820_0, i_10_359_1909_0, i_10_359_1912_0,
    i_10_359_1929_0, i_10_359_1947_0, i_10_359_1950_0, i_10_359_1984_0,
    i_10_359_1985_0, i_10_359_2016_0, i_10_359_2209_0, i_10_359_2351_0,
    i_10_359_2512_0, i_10_359_2651_0, i_10_359_2656_0, i_10_359_2657_0,
    i_10_359_2659_0, i_10_359_2695_0, i_10_359_2709_0, i_10_359_2710_0,
    i_10_359_2732_0, i_10_359_2754_0, i_10_359_2826_0, i_10_359_2828_0,
    i_10_359_2831_0, i_10_359_2832_0, i_10_359_2840_0, i_10_359_2880_0,
    i_10_359_2916_0, i_10_359_2918_0, i_10_359_2919_0, i_10_359_2920_0,
    i_10_359_2921_0, i_10_359_2922_0, i_10_359_3046_0, i_10_359_3087_0,
    i_10_359_3090_0, i_10_359_3235_0, i_10_359_3269_0, i_10_359_3272_0,
    i_10_359_3313_0, i_10_359_3315_0, i_10_359_3321_0, i_10_359_3356_0,
    i_10_359_3432_0, i_10_359_3538_0, i_10_359_3585_0, i_10_359_3610_0,
    i_10_359_3651_0, i_10_359_3652_0, i_10_359_3664_0, i_10_359_3699_0,
    i_10_359_3718_0, i_10_359_3775_0, i_10_359_3786_0, i_10_359_3811_0,
    i_10_359_3901_0, i_10_359_3981_0, i_10_359_3982_0, i_10_359_3984_0,
    i_10_359_4091_0, i_10_359_4118_0, i_10_359_4268_0, i_10_359_4285_0,
    i_10_359_4288_0, i_10_359_4290_0, i_10_359_4291_0, i_10_359_4593_0;
  output o_10_359_0_0;
  assign o_10_359_0_0 = 0;
endmodule



// Benchmark "kernel_10_360" written by ABC on Sun Jul 19 10:27:17 2020

module kernel_10_360 ( 
    i_10_360_177_0, i_10_360_178_0, i_10_360_279_0, i_10_360_282_0,
    i_10_360_283_0, i_10_360_296_0, i_10_360_328_0, i_10_360_329_0,
    i_10_360_410_0, i_10_360_438_0, i_10_360_459_0, i_10_360_466_0,
    i_10_360_467_0, i_10_360_506_0, i_10_360_509_0, i_10_360_799_0,
    i_10_360_955_0, i_10_360_1005_0, i_10_360_1006_0, i_10_360_1007_0,
    i_10_360_1236_0, i_10_360_1239_0, i_10_360_1248_0, i_10_360_1249_0,
    i_10_360_1263_0, i_10_360_1264_0, i_10_360_1305_0, i_10_360_1448_0,
    i_10_360_1551_0, i_10_360_1552_0, i_10_360_1554_0, i_10_360_1556_0,
    i_10_360_1582_0, i_10_360_1626_0, i_10_360_1651_0, i_10_360_1678_0,
    i_10_360_1683_0, i_10_360_1689_0, i_10_360_1691_0, i_10_360_1716_0,
    i_10_360_1822_0, i_10_360_1823_0, i_10_360_1825_0, i_10_360_1912_0,
    i_10_360_2204_0, i_10_360_2310_0, i_10_360_2311_0, i_10_360_2312_0,
    i_10_360_2352_0, i_10_360_2354_0, i_10_360_2357_0, i_10_360_2364_0,
    i_10_360_2408_0, i_10_360_2469_0, i_10_360_2470_0, i_10_360_2481_0,
    i_10_360_2633_0, i_10_360_2635_0, i_10_360_2661_0, i_10_360_2663_0,
    i_10_360_2704_0, i_10_360_2708_0, i_10_360_2715_0, i_10_360_2716_0,
    i_10_360_2717_0, i_10_360_2727_0, i_10_360_2731_0, i_10_360_2732_0,
    i_10_360_2735_0, i_10_360_2832_0, i_10_360_2923_0, i_10_360_3072_0,
    i_10_360_3157_0, i_10_360_3158_0, i_10_360_3279_0, i_10_360_3280_0,
    i_10_360_3386_0, i_10_360_3497_0, i_10_360_3501_0, i_10_360_3540_0,
    i_10_360_3543_0, i_10_360_3585_0, i_10_360_3586_0, i_10_360_3649_0,
    i_10_360_3650_0, i_10_360_3653_0, i_10_360_3784_0, i_10_360_3788_0,
    i_10_360_3847_0, i_10_360_3859_0, i_10_360_3895_0, i_10_360_3896_0,
    i_10_360_3906_0, i_10_360_3985_0, i_10_360_4116_0, i_10_360_4117_0,
    i_10_360_4118_0, i_10_360_4121_0, i_10_360_4236_0, i_10_360_4237_0,
    o_10_360_0_0  );
  input  i_10_360_177_0, i_10_360_178_0, i_10_360_279_0, i_10_360_282_0,
    i_10_360_283_0, i_10_360_296_0, i_10_360_328_0, i_10_360_329_0,
    i_10_360_410_0, i_10_360_438_0, i_10_360_459_0, i_10_360_466_0,
    i_10_360_467_0, i_10_360_506_0, i_10_360_509_0, i_10_360_799_0,
    i_10_360_955_0, i_10_360_1005_0, i_10_360_1006_0, i_10_360_1007_0,
    i_10_360_1236_0, i_10_360_1239_0, i_10_360_1248_0, i_10_360_1249_0,
    i_10_360_1263_0, i_10_360_1264_0, i_10_360_1305_0, i_10_360_1448_0,
    i_10_360_1551_0, i_10_360_1552_0, i_10_360_1554_0, i_10_360_1556_0,
    i_10_360_1582_0, i_10_360_1626_0, i_10_360_1651_0, i_10_360_1678_0,
    i_10_360_1683_0, i_10_360_1689_0, i_10_360_1691_0, i_10_360_1716_0,
    i_10_360_1822_0, i_10_360_1823_0, i_10_360_1825_0, i_10_360_1912_0,
    i_10_360_2204_0, i_10_360_2310_0, i_10_360_2311_0, i_10_360_2312_0,
    i_10_360_2352_0, i_10_360_2354_0, i_10_360_2357_0, i_10_360_2364_0,
    i_10_360_2408_0, i_10_360_2469_0, i_10_360_2470_0, i_10_360_2481_0,
    i_10_360_2633_0, i_10_360_2635_0, i_10_360_2661_0, i_10_360_2663_0,
    i_10_360_2704_0, i_10_360_2708_0, i_10_360_2715_0, i_10_360_2716_0,
    i_10_360_2717_0, i_10_360_2727_0, i_10_360_2731_0, i_10_360_2732_0,
    i_10_360_2735_0, i_10_360_2832_0, i_10_360_2923_0, i_10_360_3072_0,
    i_10_360_3157_0, i_10_360_3158_0, i_10_360_3279_0, i_10_360_3280_0,
    i_10_360_3386_0, i_10_360_3497_0, i_10_360_3501_0, i_10_360_3540_0,
    i_10_360_3543_0, i_10_360_3585_0, i_10_360_3586_0, i_10_360_3649_0,
    i_10_360_3650_0, i_10_360_3653_0, i_10_360_3784_0, i_10_360_3788_0,
    i_10_360_3847_0, i_10_360_3859_0, i_10_360_3895_0, i_10_360_3896_0,
    i_10_360_3906_0, i_10_360_3985_0, i_10_360_4116_0, i_10_360_4117_0,
    i_10_360_4118_0, i_10_360_4121_0, i_10_360_4236_0, i_10_360_4237_0;
  output o_10_360_0_0;
  assign o_10_360_0_0 = ~((~i_10_360_2312_0 & ((~i_10_360_282_0 & ((~i_10_360_296_0 & ~i_10_360_1556_0 & ~i_10_360_1626_0 & ~i_10_360_2310_0 & ~i_10_360_2311_0 & ~i_10_360_2481_0 & ~i_10_360_3072_0 & ~i_10_360_3906_0 & ~i_10_360_3985_0) | (~i_10_360_178_0 & ~i_10_360_1448_0 & ~i_10_360_1554_0 & ~i_10_360_3585_0 & ~i_10_360_4237_0))) | (~i_10_360_3543_0 & ((~i_10_360_1006_0 & ((~i_10_360_410_0 & ~i_10_360_2311_0 & ~i_10_360_2408_0 & i_10_360_2727_0 & ~i_10_360_2832_0 & ~i_10_360_3501_0 & ~i_10_360_3985_0 & ~i_10_360_4236_0) | (~i_10_360_1007_0 & i_10_360_1691_0 & ~i_10_360_2704_0 & ~i_10_360_3649_0 & ~i_10_360_4237_0))) | (~i_10_360_177_0 & ~i_10_360_1005_0 & ~i_10_360_1683_0 & ~i_10_360_1823_0 & ~i_10_360_2704_0 & ~i_10_360_3279_0 & ~i_10_360_3650_0 & ~i_10_360_3847_0 & ~i_10_360_3859_0))) | (~i_10_360_1448_0 & i_10_360_2661_0 & i_10_360_3653_0))) | (~i_10_360_1551_0 & ((~i_10_360_177_0 & ((~i_10_360_1007_0 & ~i_10_360_1264_0 & ~i_10_360_2364_0 & ~i_10_360_2633_0 & ~i_10_360_2715_0 & i_10_360_2732_0 & ~i_10_360_3788_0) | (~i_10_360_1626_0 & ~i_10_360_2635_0 & ~i_10_360_3543_0 & i_10_360_3649_0 & ~i_10_360_3906_0))) | (~i_10_360_283_0 & i_10_360_1236_0 & i_10_360_1239_0 & ~i_10_360_2715_0 & ~i_10_360_2717_0 & ~i_10_360_3540_0 & ~i_10_360_4237_0))) | (~i_10_360_1005_0 & ~i_10_360_3585_0 & ((~i_10_360_1236_0 & ~i_10_360_2704_0 & ~i_10_360_2716_0 & ~i_10_360_3586_0 & ~i_10_360_3650_0) | (~i_10_360_329_0 & ~i_10_360_1007_0 & ~i_10_360_2311_0 & ~i_10_360_2470_0 & ~i_10_360_2481_0 & ~i_10_360_2727_0 & ~i_10_360_3543_0 & ~i_10_360_3906_0))) | (~i_10_360_1552_0 & ((i_10_360_1683_0 & ~i_10_360_1912_0 & ~i_10_360_2352_0 & ~i_10_360_2715_0 & ~i_10_360_2717_0 & ~i_10_360_2732_0 & ~i_10_360_3072_0) | (~i_10_360_296_0 & ~i_10_360_328_0 & ~i_10_360_1689_0 & ~i_10_360_2716_0 & ~i_10_360_3280_0 & ~i_10_360_3497_0 & ~i_10_360_3501_0 & ~i_10_360_3543_0))) | (~i_10_360_328_0 & ~i_10_360_2715_0 & ((~i_10_360_1263_0 & ~i_10_360_2352_0 & i_10_360_2633_0 & i_10_360_2635_0 & ~i_10_360_3497_0 & ~i_10_360_3540_0) | (~i_10_360_283_0 & ~i_10_360_1006_0 & ~i_10_360_1554_0 & ~i_10_360_1626_0 & ~i_10_360_2481_0 & ~i_10_360_3501_0 & ~i_10_360_3543_0 & ~i_10_360_4236_0))) | (~i_10_360_1006_0 & ((i_10_360_178_0 & ~i_10_360_1264_0 & i_10_360_2708_0 & ~i_10_360_2732_0 & ~i_10_360_3280_0 & ~i_10_360_4236_0) | (i_10_360_2633_0 & ~i_10_360_3501_0 & ~i_10_360_3895_0 & ~i_10_360_4237_0))) | (~i_10_360_4236_0 & ((~i_10_360_1305_0 & ~i_10_360_1582_0 & i_10_360_2731_0 & ~i_10_360_2732_0 & ~i_10_360_3386_0 & ~i_10_360_3540_0 & ~i_10_360_3650_0) | (~i_10_360_3279_0 & ~i_10_360_3280_0 & i_10_360_4116_0 & ~i_10_360_4237_0))) | (~i_10_360_1239_0 & i_10_360_1689_0 & i_10_360_1912_0) | (~i_10_360_459_0 & ~i_10_360_1007_0 & ~i_10_360_1448_0 & ~i_10_360_1683_0 & ~i_10_360_2310_0 & ~i_10_360_2311_0 & ~i_10_360_2408_0 & ~i_10_360_2469_0 & ~i_10_360_2716_0 & ~i_10_360_3906_0 & ~i_10_360_3985_0) | (i_10_360_3649_0 & i_10_360_4117_0 & ~i_10_360_4118_0));
endmodule



// Benchmark "kernel_10_361" written by ABC on Sun Jul 19 10:27:18 2020

module kernel_10_361 ( 
    i_10_361_172_0, i_10_361_244_0, i_10_361_430_0, i_10_361_431_0,
    i_10_361_444_0, i_10_361_447_0, i_10_361_466_0, i_10_361_467_0,
    i_10_361_589_0, i_10_361_744_0, i_10_361_798_0, i_10_361_820_0,
    i_10_361_1007_0, i_10_361_1032_0, i_10_361_1043_0, i_10_361_1060_0,
    i_10_361_1061_0, i_10_361_1083_0, i_10_361_1132_0, i_10_361_1215_0,
    i_10_361_1233_0, i_10_361_1237_0, i_10_361_1241_0, i_10_361_1349_0,
    i_10_361_1580_0, i_10_361_1582_0, i_10_361_1648_0, i_10_361_1649_0,
    i_10_361_1652_0, i_10_361_1654_0, i_10_361_1684_0, i_10_361_1687_0,
    i_10_361_1690_0, i_10_361_1736_0, i_10_361_1772_0, i_10_361_1821_0,
    i_10_361_1822_0, i_10_361_2023_0, i_10_361_2201_0, i_10_361_2349_0,
    i_10_361_2352_0, i_10_361_2355_0, i_10_361_2374_0, i_10_361_2450_0,
    i_10_361_2468_0, i_10_361_2516_0, i_10_361_2584_0, i_10_361_2632_0,
    i_10_361_2634_0, i_10_361_2659_0, i_10_361_2701_0, i_10_361_2707_0,
    i_10_361_2727_0, i_10_361_2729_0, i_10_361_2741_0, i_10_361_2743_0,
    i_10_361_2829_0, i_10_361_2831_0, i_10_361_2919_0, i_10_361_2921_0,
    i_10_361_2923_0, i_10_361_3073_0, i_10_361_3075_0, i_10_361_3199_0,
    i_10_361_3271_0, i_10_361_3283_0, i_10_361_3326_0, i_10_361_3384_0,
    i_10_361_3387_0, i_10_361_3388_0, i_10_361_3390_0, i_10_361_3391_0,
    i_10_361_3468_0, i_10_361_3470_0, i_10_361_3522_0, i_10_361_3523_0,
    i_10_361_3544_0, i_10_361_3613_0, i_10_361_3615_0, i_10_361_3616_0,
    i_10_361_3617_0, i_10_361_3649_0, i_10_361_3668_0, i_10_361_3726_0,
    i_10_361_3784_0, i_10_361_3838_0, i_10_361_3848_0, i_10_361_3853_0,
    i_10_361_3855_0, i_10_361_3857_0, i_10_361_3990_0, i_10_361_4173_0,
    i_10_361_4174_0, i_10_361_4208_0, i_10_361_4238_0, i_10_361_4281_0,
    i_10_361_4287_0, i_10_361_4288_0, i_10_361_4289_0, i_10_361_4571_0,
    o_10_361_0_0  );
  input  i_10_361_172_0, i_10_361_244_0, i_10_361_430_0, i_10_361_431_0,
    i_10_361_444_0, i_10_361_447_0, i_10_361_466_0, i_10_361_467_0,
    i_10_361_589_0, i_10_361_744_0, i_10_361_798_0, i_10_361_820_0,
    i_10_361_1007_0, i_10_361_1032_0, i_10_361_1043_0, i_10_361_1060_0,
    i_10_361_1061_0, i_10_361_1083_0, i_10_361_1132_0, i_10_361_1215_0,
    i_10_361_1233_0, i_10_361_1237_0, i_10_361_1241_0, i_10_361_1349_0,
    i_10_361_1580_0, i_10_361_1582_0, i_10_361_1648_0, i_10_361_1649_0,
    i_10_361_1652_0, i_10_361_1654_0, i_10_361_1684_0, i_10_361_1687_0,
    i_10_361_1690_0, i_10_361_1736_0, i_10_361_1772_0, i_10_361_1821_0,
    i_10_361_1822_0, i_10_361_2023_0, i_10_361_2201_0, i_10_361_2349_0,
    i_10_361_2352_0, i_10_361_2355_0, i_10_361_2374_0, i_10_361_2450_0,
    i_10_361_2468_0, i_10_361_2516_0, i_10_361_2584_0, i_10_361_2632_0,
    i_10_361_2634_0, i_10_361_2659_0, i_10_361_2701_0, i_10_361_2707_0,
    i_10_361_2727_0, i_10_361_2729_0, i_10_361_2741_0, i_10_361_2743_0,
    i_10_361_2829_0, i_10_361_2831_0, i_10_361_2919_0, i_10_361_2921_0,
    i_10_361_2923_0, i_10_361_3073_0, i_10_361_3075_0, i_10_361_3199_0,
    i_10_361_3271_0, i_10_361_3283_0, i_10_361_3326_0, i_10_361_3384_0,
    i_10_361_3387_0, i_10_361_3388_0, i_10_361_3390_0, i_10_361_3391_0,
    i_10_361_3468_0, i_10_361_3470_0, i_10_361_3522_0, i_10_361_3523_0,
    i_10_361_3544_0, i_10_361_3613_0, i_10_361_3615_0, i_10_361_3616_0,
    i_10_361_3617_0, i_10_361_3649_0, i_10_361_3668_0, i_10_361_3726_0,
    i_10_361_3784_0, i_10_361_3838_0, i_10_361_3848_0, i_10_361_3853_0,
    i_10_361_3855_0, i_10_361_3857_0, i_10_361_3990_0, i_10_361_4173_0,
    i_10_361_4174_0, i_10_361_4208_0, i_10_361_4238_0, i_10_361_4281_0,
    i_10_361_4287_0, i_10_361_4288_0, i_10_361_4289_0, i_10_361_4571_0;
  output o_10_361_0_0;
  assign o_10_361_0_0 = 0;
endmodule



// Benchmark "kernel_10_362" written by ABC on Sun Jul 19 10:27:19 2020

module kernel_10_362 ( 
    i_10_362_85_0, i_10_362_261_0, i_10_362_279_0, i_10_362_281_0,
    i_10_362_284_0, i_10_362_285_0, i_10_362_393_0, i_10_362_436_0,
    i_10_362_498_0, i_10_362_502_0, i_10_362_558_0, i_10_362_600_0,
    i_10_362_643_0, i_10_362_698_0, i_10_362_711_0, i_10_362_724_0,
    i_10_362_727_0, i_10_362_822_0, i_10_362_852_0, i_10_362_876_0,
    i_10_362_1029_0, i_10_362_1086_0, i_10_362_1133_0, i_10_362_1222_0,
    i_10_362_1239_0, i_10_362_1299_0, i_10_362_1332_0, i_10_362_1348_0,
    i_10_362_1434_0, i_10_362_1449_0, i_10_362_1542_0, i_10_362_1551_0,
    i_10_362_1579_0, i_10_362_1605_0, i_10_362_1623_0, i_10_362_1624_0,
    i_10_362_1711_0, i_10_362_1803_0, i_10_362_1804_0, i_10_362_1954_0,
    i_10_362_1956_0, i_10_362_2001_0, i_10_362_2002_0, i_10_362_2010_0,
    i_10_362_2028_0, i_10_362_2091_0, i_10_362_2109_0, i_10_362_2155_0,
    i_10_362_2162_0, i_10_362_2202_0, i_10_362_2349_0, i_10_362_2356_0,
    i_10_362_2451_0, i_10_362_2452_0, i_10_362_2515_0, i_10_362_2599_0,
    i_10_362_2730_0, i_10_362_2731_0, i_10_362_2732_0, i_10_362_2737_0,
    i_10_362_2742_0, i_10_362_2743_0, i_10_362_2744_0, i_10_362_2832_0,
    i_10_362_2880_0, i_10_362_2884_0, i_10_362_2955_0, i_10_362_2958_0,
    i_10_362_2974_0, i_10_362_3048_0, i_10_362_3109_0, i_10_362_3162_0,
    i_10_362_3272_0, i_10_362_3392_0, i_10_362_3472_0, i_10_362_3492_0,
    i_10_362_3504_0, i_10_362_3544_0, i_10_362_3546_0, i_10_362_3729_0,
    i_10_362_3777_0, i_10_362_3840_0, i_10_362_3851_0, i_10_362_3859_0,
    i_10_362_3860_0, i_10_362_3922_0, i_10_362_3978_0, i_10_362_4126_0,
    i_10_362_4216_0, i_10_362_4218_0, i_10_362_4269_0, i_10_362_4270_0,
    i_10_362_4278_0, i_10_362_4287_0, i_10_362_4392_0, i_10_362_4563_0,
    i_10_362_4571_0, i_10_362_4582_0, i_10_362_4585_0, i_10_362_4588_0,
    o_10_362_0_0  );
  input  i_10_362_85_0, i_10_362_261_0, i_10_362_279_0, i_10_362_281_0,
    i_10_362_284_0, i_10_362_285_0, i_10_362_393_0, i_10_362_436_0,
    i_10_362_498_0, i_10_362_502_0, i_10_362_558_0, i_10_362_600_0,
    i_10_362_643_0, i_10_362_698_0, i_10_362_711_0, i_10_362_724_0,
    i_10_362_727_0, i_10_362_822_0, i_10_362_852_0, i_10_362_876_0,
    i_10_362_1029_0, i_10_362_1086_0, i_10_362_1133_0, i_10_362_1222_0,
    i_10_362_1239_0, i_10_362_1299_0, i_10_362_1332_0, i_10_362_1348_0,
    i_10_362_1434_0, i_10_362_1449_0, i_10_362_1542_0, i_10_362_1551_0,
    i_10_362_1579_0, i_10_362_1605_0, i_10_362_1623_0, i_10_362_1624_0,
    i_10_362_1711_0, i_10_362_1803_0, i_10_362_1804_0, i_10_362_1954_0,
    i_10_362_1956_0, i_10_362_2001_0, i_10_362_2002_0, i_10_362_2010_0,
    i_10_362_2028_0, i_10_362_2091_0, i_10_362_2109_0, i_10_362_2155_0,
    i_10_362_2162_0, i_10_362_2202_0, i_10_362_2349_0, i_10_362_2356_0,
    i_10_362_2451_0, i_10_362_2452_0, i_10_362_2515_0, i_10_362_2599_0,
    i_10_362_2730_0, i_10_362_2731_0, i_10_362_2732_0, i_10_362_2737_0,
    i_10_362_2742_0, i_10_362_2743_0, i_10_362_2744_0, i_10_362_2832_0,
    i_10_362_2880_0, i_10_362_2884_0, i_10_362_2955_0, i_10_362_2958_0,
    i_10_362_2974_0, i_10_362_3048_0, i_10_362_3109_0, i_10_362_3162_0,
    i_10_362_3272_0, i_10_362_3392_0, i_10_362_3472_0, i_10_362_3492_0,
    i_10_362_3504_0, i_10_362_3544_0, i_10_362_3546_0, i_10_362_3729_0,
    i_10_362_3777_0, i_10_362_3840_0, i_10_362_3851_0, i_10_362_3859_0,
    i_10_362_3860_0, i_10_362_3922_0, i_10_362_3978_0, i_10_362_4126_0,
    i_10_362_4216_0, i_10_362_4218_0, i_10_362_4269_0, i_10_362_4270_0,
    i_10_362_4278_0, i_10_362_4287_0, i_10_362_4392_0, i_10_362_4563_0,
    i_10_362_4571_0, i_10_362_4582_0, i_10_362_4585_0, i_10_362_4588_0;
  output o_10_362_0_0;
  assign o_10_362_0_0 = 0;
endmodule



// Benchmark "kernel_10_363" written by ABC on Sun Jul 19 10:27:20 2020

module kernel_10_363 ( 
    i_10_363_52_0, i_10_363_160_0, i_10_363_276_0, i_10_363_319_0,
    i_10_363_328_0, i_10_363_388_0, i_10_363_393_0, i_10_363_439_0,
    i_10_363_446_0, i_10_363_463_0, i_10_363_466_0, i_10_363_634_0,
    i_10_363_635_0, i_10_363_718_0, i_10_363_793_0, i_10_363_795_0,
    i_10_363_796_0, i_10_363_797_0, i_10_363_799_0, i_10_363_830_0,
    i_10_363_832_0, i_10_363_919_0, i_10_363_996_0, i_10_363_1116_0,
    i_10_363_1209_0, i_10_363_1210_0, i_10_363_1270_0, i_10_363_1295_0,
    i_10_363_1305_0, i_10_363_1477_0, i_10_363_1492_0, i_10_363_1493_0,
    i_10_363_1580_0, i_10_363_1655_0, i_10_363_1690_0, i_10_363_1821_0,
    i_10_363_1822_0, i_10_363_1823_0, i_10_363_1885_0, i_10_363_1889_0,
    i_10_363_1937_0, i_10_363_1939_0, i_10_363_1940_0, i_10_363_1957_0,
    i_10_363_2002_0, i_10_363_2004_0, i_10_363_2006_0, i_10_363_2086_0,
    i_10_363_2245_0, i_10_363_2386_0, i_10_363_2453_0, i_10_363_2455_0,
    i_10_363_2467_0, i_10_363_2474_0, i_10_363_2516_0, i_10_363_2582_0,
    i_10_363_2681_0, i_10_363_2701_0, i_10_363_2715_0, i_10_363_2716_0,
    i_10_363_2740_0, i_10_363_2825_0, i_10_363_2923_0, i_10_363_2983_0,
    i_10_363_2987_0, i_10_363_3119_0, i_10_363_3122_0, i_10_363_3270_0,
    i_10_363_3274_0, i_10_363_3387_0, i_10_363_3392_0, i_10_363_3466_0,
    i_10_363_3467_0, i_10_363_3496_0, i_10_363_3497_0, i_10_363_3538_0,
    i_10_363_3539_0, i_10_363_3541_0, i_10_363_3586_0, i_10_363_3622_0,
    i_10_363_3644_0, i_10_363_3645_0, i_10_363_3786_0, i_10_363_3878_0,
    i_10_363_3879_0, i_10_363_3946_0, i_10_363_4061_0, i_10_363_4116_0,
    i_10_363_4118_0, i_10_363_4119_0, i_10_363_4120_0, i_10_363_4121_0,
    i_10_363_4125_0, i_10_363_4155_0, i_10_363_4156_0, i_10_363_4269_0,
    i_10_363_4270_0, i_10_363_4273_0, i_10_363_4566_0, i_10_363_4569_0,
    o_10_363_0_0  );
  input  i_10_363_52_0, i_10_363_160_0, i_10_363_276_0, i_10_363_319_0,
    i_10_363_328_0, i_10_363_388_0, i_10_363_393_0, i_10_363_439_0,
    i_10_363_446_0, i_10_363_463_0, i_10_363_466_0, i_10_363_634_0,
    i_10_363_635_0, i_10_363_718_0, i_10_363_793_0, i_10_363_795_0,
    i_10_363_796_0, i_10_363_797_0, i_10_363_799_0, i_10_363_830_0,
    i_10_363_832_0, i_10_363_919_0, i_10_363_996_0, i_10_363_1116_0,
    i_10_363_1209_0, i_10_363_1210_0, i_10_363_1270_0, i_10_363_1295_0,
    i_10_363_1305_0, i_10_363_1477_0, i_10_363_1492_0, i_10_363_1493_0,
    i_10_363_1580_0, i_10_363_1655_0, i_10_363_1690_0, i_10_363_1821_0,
    i_10_363_1822_0, i_10_363_1823_0, i_10_363_1885_0, i_10_363_1889_0,
    i_10_363_1937_0, i_10_363_1939_0, i_10_363_1940_0, i_10_363_1957_0,
    i_10_363_2002_0, i_10_363_2004_0, i_10_363_2006_0, i_10_363_2086_0,
    i_10_363_2245_0, i_10_363_2386_0, i_10_363_2453_0, i_10_363_2455_0,
    i_10_363_2467_0, i_10_363_2474_0, i_10_363_2516_0, i_10_363_2582_0,
    i_10_363_2681_0, i_10_363_2701_0, i_10_363_2715_0, i_10_363_2716_0,
    i_10_363_2740_0, i_10_363_2825_0, i_10_363_2923_0, i_10_363_2983_0,
    i_10_363_2987_0, i_10_363_3119_0, i_10_363_3122_0, i_10_363_3270_0,
    i_10_363_3274_0, i_10_363_3387_0, i_10_363_3392_0, i_10_363_3466_0,
    i_10_363_3467_0, i_10_363_3496_0, i_10_363_3497_0, i_10_363_3538_0,
    i_10_363_3539_0, i_10_363_3541_0, i_10_363_3586_0, i_10_363_3622_0,
    i_10_363_3644_0, i_10_363_3645_0, i_10_363_3786_0, i_10_363_3878_0,
    i_10_363_3879_0, i_10_363_3946_0, i_10_363_4061_0, i_10_363_4116_0,
    i_10_363_4118_0, i_10_363_4119_0, i_10_363_4120_0, i_10_363_4121_0,
    i_10_363_4125_0, i_10_363_4155_0, i_10_363_4156_0, i_10_363_4269_0,
    i_10_363_4270_0, i_10_363_4273_0, i_10_363_4566_0, i_10_363_4569_0;
  output o_10_363_0_0;
  assign o_10_363_0_0 = 0;
endmodule



// Benchmark "kernel_10_364" written by ABC on Sun Jul 19 10:27:21 2020

module kernel_10_364 ( 
    i_10_364_38_0, i_10_364_43_0, i_10_364_47_0, i_10_364_118_0,
    i_10_364_127_0, i_10_364_130_0, i_10_364_131_0, i_10_364_171_0,
    i_10_364_181_0, i_10_364_244_0, i_10_364_349_0, i_10_364_361_0,
    i_10_364_391_0, i_10_364_424_0, i_10_364_427_0, i_10_364_437_0,
    i_10_364_439_0, i_10_364_442_0, i_10_364_459_0, i_10_364_560_0,
    i_10_364_740_0, i_10_364_794_0, i_10_364_820_0, i_10_364_956_0,
    i_10_364_982_0, i_10_364_999_0, i_10_364_1000_0, i_10_364_1084_0,
    i_10_364_1088_0, i_10_364_1215_0, i_10_364_1234_0, i_10_364_1235_0,
    i_10_364_1236_0, i_10_364_1237_0, i_10_364_1296_0, i_10_364_1345_0,
    i_10_364_1378_0, i_10_364_1546_0, i_10_364_1579_0, i_10_364_1693_0,
    i_10_364_1909_0, i_10_364_1944_0, i_10_364_1947_0, i_10_364_2025_0,
    i_10_364_2037_0, i_10_364_2089_0, i_10_364_2113_0, i_10_364_2204_0,
    i_10_364_2270_0, i_10_364_2272_0, i_10_364_2305_0, i_10_364_2341_0,
    i_10_364_2351_0, i_10_364_2354_0, i_10_364_2361_0, i_10_364_2453_0,
    i_10_364_2455_0, i_10_364_2459_0, i_10_364_2468_0, i_10_364_2606_0,
    i_10_364_2631_0, i_10_364_2634_0, i_10_364_2700_0, i_10_364_2703_0,
    i_10_364_2725_0, i_10_364_2783_0, i_10_364_2863_0, i_10_364_2910_0,
    i_10_364_2961_0, i_10_364_3036_0, i_10_364_3037_0, i_10_364_3038_0,
    i_10_364_3042_0, i_10_364_3154_0, i_10_364_3163_0, i_10_364_3232_0,
    i_10_364_3352_0, i_10_364_3356_0, i_10_364_3466_0, i_10_364_3523_0,
    i_10_364_3541_0, i_10_364_3553_0, i_10_364_3556_0, i_10_364_3582_0,
    i_10_364_3584_0, i_10_364_3617_0, i_10_364_3686_0, i_10_364_3838_0,
    i_10_364_3860_0, i_10_364_4023_0, i_10_364_4053_0, i_10_364_4118_0,
    i_10_364_4154_0, i_10_364_4169_0, i_10_364_4204_0, i_10_364_4367_0,
    i_10_364_4394_0, i_10_364_4395_0, i_10_364_4432_0, i_10_364_4593_0,
    o_10_364_0_0  );
  input  i_10_364_38_0, i_10_364_43_0, i_10_364_47_0, i_10_364_118_0,
    i_10_364_127_0, i_10_364_130_0, i_10_364_131_0, i_10_364_171_0,
    i_10_364_181_0, i_10_364_244_0, i_10_364_349_0, i_10_364_361_0,
    i_10_364_391_0, i_10_364_424_0, i_10_364_427_0, i_10_364_437_0,
    i_10_364_439_0, i_10_364_442_0, i_10_364_459_0, i_10_364_560_0,
    i_10_364_740_0, i_10_364_794_0, i_10_364_820_0, i_10_364_956_0,
    i_10_364_982_0, i_10_364_999_0, i_10_364_1000_0, i_10_364_1084_0,
    i_10_364_1088_0, i_10_364_1215_0, i_10_364_1234_0, i_10_364_1235_0,
    i_10_364_1236_0, i_10_364_1237_0, i_10_364_1296_0, i_10_364_1345_0,
    i_10_364_1378_0, i_10_364_1546_0, i_10_364_1579_0, i_10_364_1693_0,
    i_10_364_1909_0, i_10_364_1944_0, i_10_364_1947_0, i_10_364_2025_0,
    i_10_364_2037_0, i_10_364_2089_0, i_10_364_2113_0, i_10_364_2204_0,
    i_10_364_2270_0, i_10_364_2272_0, i_10_364_2305_0, i_10_364_2341_0,
    i_10_364_2351_0, i_10_364_2354_0, i_10_364_2361_0, i_10_364_2453_0,
    i_10_364_2455_0, i_10_364_2459_0, i_10_364_2468_0, i_10_364_2606_0,
    i_10_364_2631_0, i_10_364_2634_0, i_10_364_2700_0, i_10_364_2703_0,
    i_10_364_2725_0, i_10_364_2783_0, i_10_364_2863_0, i_10_364_2910_0,
    i_10_364_2961_0, i_10_364_3036_0, i_10_364_3037_0, i_10_364_3038_0,
    i_10_364_3042_0, i_10_364_3154_0, i_10_364_3163_0, i_10_364_3232_0,
    i_10_364_3352_0, i_10_364_3356_0, i_10_364_3466_0, i_10_364_3523_0,
    i_10_364_3541_0, i_10_364_3553_0, i_10_364_3556_0, i_10_364_3582_0,
    i_10_364_3584_0, i_10_364_3617_0, i_10_364_3686_0, i_10_364_3838_0,
    i_10_364_3860_0, i_10_364_4023_0, i_10_364_4053_0, i_10_364_4118_0,
    i_10_364_4154_0, i_10_364_4169_0, i_10_364_4204_0, i_10_364_4367_0,
    i_10_364_4394_0, i_10_364_4395_0, i_10_364_4432_0, i_10_364_4593_0;
  output o_10_364_0_0;
  assign o_10_364_0_0 = 0;
endmodule



// Benchmark "kernel_10_365" written by ABC on Sun Jul 19 10:27:22 2020

module kernel_10_365 ( 
    i_10_365_216_0, i_10_365_246_0, i_10_365_249_0, i_10_365_275_0,
    i_10_365_278_0, i_10_365_282_0, i_10_365_283_0, i_10_365_287_0,
    i_10_365_324_0, i_10_365_329_0, i_10_365_465_0, i_10_365_508_0,
    i_10_365_750_0, i_10_365_751_0, i_10_365_799_0, i_10_365_898_0,
    i_10_365_957_0, i_10_365_1002_0, i_10_365_1029_0, i_10_365_1032_0,
    i_10_365_1128_0, i_10_365_1138_0, i_10_365_1139_0, i_10_365_1162_0,
    i_10_365_1239_0, i_10_365_1240_0, i_10_365_1241_0, i_10_365_1242_0,
    i_10_365_1243_0, i_10_365_1244_0, i_10_365_1245_0, i_10_365_1265_0,
    i_10_365_1308_0, i_10_365_1345_0, i_10_365_1575_0, i_10_365_1578_0,
    i_10_365_1579_0, i_10_365_1581_0, i_10_365_1614_0, i_10_365_1647_0,
    i_10_365_1650_0, i_10_365_1651_0, i_10_365_1655_0, i_10_365_1687_0,
    i_10_365_1764_0, i_10_365_1819_0, i_10_365_1826_0, i_10_365_2355_0,
    i_10_365_2449_0, i_10_365_2456_0, i_10_365_2463_0, i_10_365_2604_0,
    i_10_365_2628_0, i_10_365_2631_0, i_10_365_2632_0, i_10_365_2643_0,
    i_10_365_2718_0, i_10_365_2724_0, i_10_365_2832_0, i_10_365_2833_0,
    i_10_365_2916_0, i_10_365_2917_0, i_10_365_2919_0, i_10_365_2922_0,
    i_10_365_2979_0, i_10_365_3034_0, i_10_365_3037_0, i_10_365_3162_0,
    i_10_365_3203_0, i_10_365_3277_0, i_10_365_3280_0, i_10_365_3325_0,
    i_10_365_3386_0, i_10_365_3402_0, i_10_365_3409_0, i_10_365_3588_0,
    i_10_365_3645_0, i_10_365_3648_0, i_10_365_3653_0, i_10_365_3729_0,
    i_10_365_3781_0, i_10_365_3783_0, i_10_365_3785_0, i_10_365_3786_0,
    i_10_365_3841_0, i_10_365_3844_0, i_10_365_3852_0, i_10_365_3855_0,
    i_10_365_4115_0, i_10_365_4116_0, i_10_365_4117_0, i_10_365_4118_0,
    i_10_365_4119_0, i_10_365_4120_0, i_10_365_4129_0, i_10_365_4278_0,
    i_10_365_4290_0, i_10_365_4564_0, i_10_365_4565_0, i_10_365_4566_0,
    o_10_365_0_0  );
  input  i_10_365_216_0, i_10_365_246_0, i_10_365_249_0, i_10_365_275_0,
    i_10_365_278_0, i_10_365_282_0, i_10_365_283_0, i_10_365_287_0,
    i_10_365_324_0, i_10_365_329_0, i_10_365_465_0, i_10_365_508_0,
    i_10_365_750_0, i_10_365_751_0, i_10_365_799_0, i_10_365_898_0,
    i_10_365_957_0, i_10_365_1002_0, i_10_365_1029_0, i_10_365_1032_0,
    i_10_365_1128_0, i_10_365_1138_0, i_10_365_1139_0, i_10_365_1162_0,
    i_10_365_1239_0, i_10_365_1240_0, i_10_365_1241_0, i_10_365_1242_0,
    i_10_365_1243_0, i_10_365_1244_0, i_10_365_1245_0, i_10_365_1265_0,
    i_10_365_1308_0, i_10_365_1345_0, i_10_365_1575_0, i_10_365_1578_0,
    i_10_365_1579_0, i_10_365_1581_0, i_10_365_1614_0, i_10_365_1647_0,
    i_10_365_1650_0, i_10_365_1651_0, i_10_365_1655_0, i_10_365_1687_0,
    i_10_365_1764_0, i_10_365_1819_0, i_10_365_1826_0, i_10_365_2355_0,
    i_10_365_2449_0, i_10_365_2456_0, i_10_365_2463_0, i_10_365_2604_0,
    i_10_365_2628_0, i_10_365_2631_0, i_10_365_2632_0, i_10_365_2643_0,
    i_10_365_2718_0, i_10_365_2724_0, i_10_365_2832_0, i_10_365_2833_0,
    i_10_365_2916_0, i_10_365_2917_0, i_10_365_2919_0, i_10_365_2922_0,
    i_10_365_2979_0, i_10_365_3034_0, i_10_365_3037_0, i_10_365_3162_0,
    i_10_365_3203_0, i_10_365_3277_0, i_10_365_3280_0, i_10_365_3325_0,
    i_10_365_3386_0, i_10_365_3402_0, i_10_365_3409_0, i_10_365_3588_0,
    i_10_365_3645_0, i_10_365_3648_0, i_10_365_3653_0, i_10_365_3729_0,
    i_10_365_3781_0, i_10_365_3783_0, i_10_365_3785_0, i_10_365_3786_0,
    i_10_365_3841_0, i_10_365_3844_0, i_10_365_3852_0, i_10_365_3855_0,
    i_10_365_4115_0, i_10_365_4116_0, i_10_365_4117_0, i_10_365_4118_0,
    i_10_365_4119_0, i_10_365_4120_0, i_10_365_4129_0, i_10_365_4278_0,
    i_10_365_4290_0, i_10_365_4564_0, i_10_365_4565_0, i_10_365_4566_0;
  output o_10_365_0_0;
  assign o_10_365_0_0 = ~((~i_10_365_751_0 & ((~i_10_365_2463_0 & ~i_10_365_2832_0 & ~i_10_365_2922_0 & i_10_365_4118_0 & i_10_365_4120_0) | (i_10_365_1655_0 & ~i_10_365_2355_0 & ~i_10_365_4115_0 & ~i_10_365_4565_0 & i_10_365_4566_0))) | (~i_10_365_1575_0 & ((~i_10_365_1581_0 & ~i_10_365_2463_0 & ~i_10_365_3037_0 & ~i_10_365_3409_0) | (i_10_365_799_0 & ~i_10_365_957_0 & ~i_10_365_3402_0 & ~i_10_365_3781_0))) | (~i_10_365_4565_0 & ((~i_10_365_957_0 & ((~i_10_365_2604_0 & i_10_365_2628_0 & ~i_10_365_3781_0 & ~i_10_365_3855_0 & ~i_10_365_4119_0) | (~i_10_365_1029_0 & ~i_10_365_2449_0 & ~i_10_365_2832_0 & ~i_10_365_3386_0 & ~i_10_365_3786_0 & ~i_10_365_3852_0 & ~i_10_365_4120_0))) | (~i_10_365_287_0 & ~i_10_365_750_0 & ~i_10_365_1029_0 & ~i_10_365_1162_0 & ~i_10_365_1826_0 & ~i_10_365_3402_0 & ~i_10_365_4278_0))) | (~i_10_365_2643_0 & ((~i_10_365_750_0 & ((~i_10_365_1242_0 & ~i_10_365_2604_0 & ~i_10_365_3162_0 & ~i_10_365_3729_0) | (~i_10_365_1029_0 & ~i_10_365_1032_0 & ~i_10_365_3280_0 & i_10_365_3781_0))) | (~i_10_365_1245_0 & ((i_10_365_1647_0 & ~i_10_365_2449_0 & ~i_10_365_2604_0 & ~i_10_365_3203_0 & ~i_10_365_4116_0) | (i_10_365_1819_0 & ~i_10_365_3162_0 & ~i_10_365_4119_0))) | (~i_10_365_2604_0 & ((~i_10_365_216_0 & ~i_10_365_3648_0 & ~i_10_365_3781_0 & i_10_365_4117_0) | (~i_10_365_1029_0 & ~i_10_365_1647_0 & ~i_10_365_4566_0))))) | (~i_10_365_750_0 & ((~i_10_365_465_0 & ~i_10_365_1243_0 & ~i_10_365_1579_0 & ~i_10_365_1819_0 & ~i_10_365_3162_0) | (~i_10_365_1265_0 & ~i_10_365_3034_0 & i_10_365_3648_0 & i_10_365_3653_0 & ~i_10_365_4129_0 & ~i_10_365_4566_0))) | (~i_10_365_1242_0 & ((~i_10_365_898_0 & ~i_10_365_1578_0 & ~i_10_365_2604_0 & ~i_10_365_3729_0) | (~i_10_365_249_0 & i_10_365_465_0 & ~i_10_365_1647_0 & ~i_10_365_2449_0 & ~i_10_365_2718_0 & ~i_10_365_4566_0))) | (~i_10_365_1245_0 & ~i_10_365_1650_0 & ~i_10_365_2832_0 & ~i_10_365_2833_0) | (~i_10_365_1647_0 & i_10_365_3588_0) | (~i_10_365_2724_0 & ~i_10_365_2922_0 & ~i_10_365_3783_0 & i_10_365_4118_0 & i_10_365_4120_0) | (i_10_365_3037_0 & ~i_10_365_4116_0 & i_10_365_4565_0));
endmodule



// Benchmark "kernel_10_366" written by ABC on Sun Jul 19 10:27:23 2020

module kernel_10_366 ( 
    i_10_366_28_0, i_10_366_70_0, i_10_366_102_0, i_10_366_103_0,
    i_10_366_120_0, i_10_366_214_0, i_10_366_220_0, i_10_366_223_0,
    i_10_366_279_0, i_10_366_280_0, i_10_366_372_0, i_10_366_373_0,
    i_10_366_375_0, i_10_366_408_0, i_10_366_424_0, i_10_366_459_0,
    i_10_366_461_0, i_10_366_463_0, i_10_366_499_0, i_10_366_586_0,
    i_10_366_588_0, i_10_366_724_0, i_10_366_792_0, i_10_366_795_0,
    i_10_366_798_0, i_10_366_919_0, i_10_366_922_0, i_10_366_957_0,
    i_10_366_960_0, i_10_366_999_0, i_10_366_1002_0, i_10_366_1039_0,
    i_10_366_1045_0, i_10_366_1164_0, i_10_366_1201_0, i_10_366_1233_0,
    i_10_366_1237_0, i_10_366_1240_0, i_10_366_1263_0, i_10_366_1380_0,
    i_10_366_1429_0, i_10_366_1648_0, i_10_366_1653_0, i_10_366_1785_0,
    i_10_366_1821_0, i_10_366_1866_0, i_10_366_1940_0, i_10_366_2004_0,
    i_10_366_2032_0, i_10_366_2094_0, i_10_366_2248_0, i_10_366_2329_0,
    i_10_366_2337_0, i_10_366_2450_0, i_10_366_2452_0, i_10_366_2470_0,
    i_10_366_2509_0, i_10_366_2510_0, i_10_366_2673_0, i_10_366_2676_0,
    i_10_366_2713_0, i_10_366_2782_0, i_10_366_2783_0, i_10_366_2839_0,
    i_10_366_2865_0, i_10_366_2869_0, i_10_366_2874_0, i_10_366_2881_0,
    i_10_366_2919_0, i_10_366_2923_0, i_10_366_2992_0, i_10_366_3070_0,
    i_10_366_3210_0, i_10_366_3238_0, i_10_366_3336_0, i_10_366_3433_0,
    i_10_366_3450_0, i_10_366_3470_0, i_10_366_3480_0, i_10_366_3496_0,
    i_10_366_3497_0, i_10_366_3559_0, i_10_366_3562_0, i_10_366_3645_0,
    i_10_366_3687_0, i_10_366_3837_0, i_10_366_3838_0, i_10_366_3841_0,
    i_10_366_3874_0, i_10_366_4055_0, i_10_366_4152_0, i_10_366_4234_0,
    i_10_366_4422_0, i_10_366_4423_0, i_10_366_4426_0, i_10_366_4434_0,
    i_10_366_4446_0, i_10_366_4447_0, i_10_366_4578_0, i_10_366_4579_0,
    o_10_366_0_0  );
  input  i_10_366_28_0, i_10_366_70_0, i_10_366_102_0, i_10_366_103_0,
    i_10_366_120_0, i_10_366_214_0, i_10_366_220_0, i_10_366_223_0,
    i_10_366_279_0, i_10_366_280_0, i_10_366_372_0, i_10_366_373_0,
    i_10_366_375_0, i_10_366_408_0, i_10_366_424_0, i_10_366_459_0,
    i_10_366_461_0, i_10_366_463_0, i_10_366_499_0, i_10_366_586_0,
    i_10_366_588_0, i_10_366_724_0, i_10_366_792_0, i_10_366_795_0,
    i_10_366_798_0, i_10_366_919_0, i_10_366_922_0, i_10_366_957_0,
    i_10_366_960_0, i_10_366_999_0, i_10_366_1002_0, i_10_366_1039_0,
    i_10_366_1045_0, i_10_366_1164_0, i_10_366_1201_0, i_10_366_1233_0,
    i_10_366_1237_0, i_10_366_1240_0, i_10_366_1263_0, i_10_366_1380_0,
    i_10_366_1429_0, i_10_366_1648_0, i_10_366_1653_0, i_10_366_1785_0,
    i_10_366_1821_0, i_10_366_1866_0, i_10_366_1940_0, i_10_366_2004_0,
    i_10_366_2032_0, i_10_366_2094_0, i_10_366_2248_0, i_10_366_2329_0,
    i_10_366_2337_0, i_10_366_2450_0, i_10_366_2452_0, i_10_366_2470_0,
    i_10_366_2509_0, i_10_366_2510_0, i_10_366_2673_0, i_10_366_2676_0,
    i_10_366_2713_0, i_10_366_2782_0, i_10_366_2783_0, i_10_366_2839_0,
    i_10_366_2865_0, i_10_366_2869_0, i_10_366_2874_0, i_10_366_2881_0,
    i_10_366_2919_0, i_10_366_2923_0, i_10_366_2992_0, i_10_366_3070_0,
    i_10_366_3210_0, i_10_366_3238_0, i_10_366_3336_0, i_10_366_3433_0,
    i_10_366_3450_0, i_10_366_3470_0, i_10_366_3480_0, i_10_366_3496_0,
    i_10_366_3497_0, i_10_366_3559_0, i_10_366_3562_0, i_10_366_3645_0,
    i_10_366_3687_0, i_10_366_3837_0, i_10_366_3838_0, i_10_366_3841_0,
    i_10_366_3874_0, i_10_366_4055_0, i_10_366_4152_0, i_10_366_4234_0,
    i_10_366_4422_0, i_10_366_4423_0, i_10_366_4426_0, i_10_366_4434_0,
    i_10_366_4446_0, i_10_366_4447_0, i_10_366_4578_0, i_10_366_4579_0;
  output o_10_366_0_0;
  assign o_10_366_0_0 = 0;
endmodule



// Benchmark "kernel_10_367" written by ABC on Sun Jul 19 10:27:25 2020

module kernel_10_367 ( 
    i_10_367_150_0, i_10_367_181_0, i_10_367_201_0, i_10_367_291_0,
    i_10_367_427_0, i_10_367_434_0, i_10_367_463_0, i_10_367_465_0,
    i_10_367_496_0, i_10_367_507_0, i_10_367_558_0, i_10_367_589_0,
    i_10_367_604_0, i_10_367_607_0, i_10_367_792_0, i_10_367_819_0,
    i_10_367_839_0, i_10_367_903_0, i_10_367_928_0, i_10_367_945_0,
    i_10_367_981_0, i_10_367_1080_0, i_10_367_1092_0, i_10_367_1120_0,
    i_10_367_1279_0, i_10_367_1353_0, i_10_367_1397_0, i_10_367_1440_0,
    i_10_367_1452_0, i_10_367_1548_0, i_10_367_1566_0, i_10_367_1652_0,
    i_10_367_1796_0, i_10_367_1819_0, i_10_367_1820_0, i_10_367_1825_0,
    i_10_367_1875_0, i_10_367_1999_0, i_10_367_2016_0, i_10_367_2018_0,
    i_10_367_2025_0, i_10_367_2107_0, i_10_367_2178_0, i_10_367_2180_0,
    i_10_367_2334_0, i_10_367_2341_0, i_10_367_2450_0, i_10_367_2502_0,
    i_10_367_2511_0, i_10_367_2556_0, i_10_367_2595_0, i_10_367_2596_0,
    i_10_367_2614_0, i_10_367_2629_0, i_10_367_2632_0, i_10_367_2635_0,
    i_10_367_2638_0, i_10_367_2664_0, i_10_367_2700_0, i_10_367_2707_0,
    i_10_367_2714_0, i_10_367_2718_0, i_10_367_2821_0, i_10_367_2831_0,
    i_10_367_2866_0, i_10_367_2881_0, i_10_367_2917_0, i_10_367_2918_0,
    i_10_367_2944_0, i_10_367_2947_0, i_10_367_2952_0, i_10_367_2953_0,
    i_10_367_3106_0, i_10_367_3235_0, i_10_367_3238_0, i_10_367_3267_0,
    i_10_367_3279_0, i_10_367_3465_0, i_10_367_3493_0, i_10_367_3520_0,
    i_10_367_3540_0, i_10_367_3541_0, i_10_367_3612_0, i_10_367_3619_0,
    i_10_367_3684_0, i_10_367_3685_0, i_10_367_3838_0, i_10_367_3855_0,
    i_10_367_3856_0, i_10_367_3883_0, i_10_367_3943_0, i_10_367_3988_0,
    i_10_367_3993_0, i_10_367_4113_0, i_10_367_4122_0, i_10_367_4194_0,
    i_10_367_4213_0, i_10_367_4268_0, i_10_367_4393_0, i_10_367_4594_0,
    o_10_367_0_0  );
  input  i_10_367_150_0, i_10_367_181_0, i_10_367_201_0, i_10_367_291_0,
    i_10_367_427_0, i_10_367_434_0, i_10_367_463_0, i_10_367_465_0,
    i_10_367_496_0, i_10_367_507_0, i_10_367_558_0, i_10_367_589_0,
    i_10_367_604_0, i_10_367_607_0, i_10_367_792_0, i_10_367_819_0,
    i_10_367_839_0, i_10_367_903_0, i_10_367_928_0, i_10_367_945_0,
    i_10_367_981_0, i_10_367_1080_0, i_10_367_1092_0, i_10_367_1120_0,
    i_10_367_1279_0, i_10_367_1353_0, i_10_367_1397_0, i_10_367_1440_0,
    i_10_367_1452_0, i_10_367_1548_0, i_10_367_1566_0, i_10_367_1652_0,
    i_10_367_1796_0, i_10_367_1819_0, i_10_367_1820_0, i_10_367_1825_0,
    i_10_367_1875_0, i_10_367_1999_0, i_10_367_2016_0, i_10_367_2018_0,
    i_10_367_2025_0, i_10_367_2107_0, i_10_367_2178_0, i_10_367_2180_0,
    i_10_367_2334_0, i_10_367_2341_0, i_10_367_2450_0, i_10_367_2502_0,
    i_10_367_2511_0, i_10_367_2556_0, i_10_367_2595_0, i_10_367_2596_0,
    i_10_367_2614_0, i_10_367_2629_0, i_10_367_2632_0, i_10_367_2635_0,
    i_10_367_2638_0, i_10_367_2664_0, i_10_367_2700_0, i_10_367_2707_0,
    i_10_367_2714_0, i_10_367_2718_0, i_10_367_2821_0, i_10_367_2831_0,
    i_10_367_2866_0, i_10_367_2881_0, i_10_367_2917_0, i_10_367_2918_0,
    i_10_367_2944_0, i_10_367_2947_0, i_10_367_2952_0, i_10_367_2953_0,
    i_10_367_3106_0, i_10_367_3235_0, i_10_367_3238_0, i_10_367_3267_0,
    i_10_367_3279_0, i_10_367_3465_0, i_10_367_3493_0, i_10_367_3520_0,
    i_10_367_3540_0, i_10_367_3541_0, i_10_367_3612_0, i_10_367_3619_0,
    i_10_367_3684_0, i_10_367_3685_0, i_10_367_3838_0, i_10_367_3855_0,
    i_10_367_3856_0, i_10_367_3883_0, i_10_367_3943_0, i_10_367_3988_0,
    i_10_367_3993_0, i_10_367_4113_0, i_10_367_4122_0, i_10_367_4194_0,
    i_10_367_4213_0, i_10_367_4268_0, i_10_367_4393_0, i_10_367_4594_0;
  output o_10_367_0_0;
  assign o_10_367_0_0 = 0;
endmodule



// Benchmark "kernel_10_368" written by ABC on Sun Jul 19 10:27:25 2020

module kernel_10_368 ( 
    i_10_368_29_0, i_10_368_253_0, i_10_368_270_0, i_10_368_271_0,
    i_10_368_284_0, i_10_368_287_0, i_10_368_390_0, i_10_368_391_0,
    i_10_368_392_0, i_10_368_495_0, i_10_368_558_0, i_10_368_694_0,
    i_10_368_963_0, i_10_368_1002_0, i_10_368_1029_0, i_10_368_1045_0,
    i_10_368_1107_0, i_10_368_1108_0, i_10_368_1206_0, i_10_368_1235_0,
    i_10_368_1238_0, i_10_368_1243_0, i_10_368_1244_0, i_10_368_1296_0,
    i_10_368_1297_0, i_10_368_1310_0, i_10_368_1528_0, i_10_368_1550_0,
    i_10_368_1575_0, i_10_368_1576_0, i_10_368_1621_0, i_10_368_1630_0,
    i_10_368_1683_0, i_10_368_1685_0, i_10_368_1686_0, i_10_368_1687_0,
    i_10_368_1688_0, i_10_368_1735_0, i_10_368_1794_0, i_10_368_1798_0,
    i_10_368_1800_0, i_10_368_1801_0, i_10_368_1820_0, i_10_368_1911_0,
    i_10_368_1912_0, i_10_368_1981_0, i_10_368_1999_0, i_10_368_2107_0,
    i_10_368_2349_0, i_10_368_2351_0, i_10_368_2380_0, i_10_368_2439_0,
    i_10_368_2440_0, i_10_368_2443_0, i_10_368_2467_0, i_10_368_2542_0,
    i_10_368_2548_0, i_10_368_2556_0, i_10_368_2566_0, i_10_368_2621_0,
    i_10_368_2701_0, i_10_368_2702_0, i_10_368_2719_0, i_10_368_2720_0,
    i_10_368_2730_0, i_10_368_2755_0, i_10_368_2817_0, i_10_368_2882_0,
    i_10_368_2969_0, i_10_368_3070_0, i_10_368_3171_0, i_10_368_3278_0,
    i_10_368_3321_0, i_10_368_3323_0, i_10_368_3355_0, i_10_368_3386_0,
    i_10_368_3407_0, i_10_368_3463_0, i_10_368_3525_0, i_10_368_3555_0,
    i_10_368_3574_0, i_10_368_3583_0, i_10_368_3647_0, i_10_368_3703_0,
    i_10_368_3704_0, i_10_368_3707_0, i_10_368_3783_0, i_10_368_3785_0,
    i_10_368_3817_0, i_10_368_3857_0, i_10_368_3871_0, i_10_368_3909_0,
    i_10_368_3910_0, i_10_368_4140_0, i_10_368_4177_0, i_10_368_4270_0,
    i_10_368_4284_0, i_10_368_4307_0, i_10_368_4431_0, i_10_368_4582_0,
    o_10_368_0_0  );
  input  i_10_368_29_0, i_10_368_253_0, i_10_368_270_0, i_10_368_271_0,
    i_10_368_284_0, i_10_368_287_0, i_10_368_390_0, i_10_368_391_0,
    i_10_368_392_0, i_10_368_495_0, i_10_368_558_0, i_10_368_694_0,
    i_10_368_963_0, i_10_368_1002_0, i_10_368_1029_0, i_10_368_1045_0,
    i_10_368_1107_0, i_10_368_1108_0, i_10_368_1206_0, i_10_368_1235_0,
    i_10_368_1238_0, i_10_368_1243_0, i_10_368_1244_0, i_10_368_1296_0,
    i_10_368_1297_0, i_10_368_1310_0, i_10_368_1528_0, i_10_368_1550_0,
    i_10_368_1575_0, i_10_368_1576_0, i_10_368_1621_0, i_10_368_1630_0,
    i_10_368_1683_0, i_10_368_1685_0, i_10_368_1686_0, i_10_368_1687_0,
    i_10_368_1688_0, i_10_368_1735_0, i_10_368_1794_0, i_10_368_1798_0,
    i_10_368_1800_0, i_10_368_1801_0, i_10_368_1820_0, i_10_368_1911_0,
    i_10_368_1912_0, i_10_368_1981_0, i_10_368_1999_0, i_10_368_2107_0,
    i_10_368_2349_0, i_10_368_2351_0, i_10_368_2380_0, i_10_368_2439_0,
    i_10_368_2440_0, i_10_368_2443_0, i_10_368_2467_0, i_10_368_2542_0,
    i_10_368_2548_0, i_10_368_2556_0, i_10_368_2566_0, i_10_368_2621_0,
    i_10_368_2701_0, i_10_368_2702_0, i_10_368_2719_0, i_10_368_2720_0,
    i_10_368_2730_0, i_10_368_2755_0, i_10_368_2817_0, i_10_368_2882_0,
    i_10_368_2969_0, i_10_368_3070_0, i_10_368_3171_0, i_10_368_3278_0,
    i_10_368_3321_0, i_10_368_3323_0, i_10_368_3355_0, i_10_368_3386_0,
    i_10_368_3407_0, i_10_368_3463_0, i_10_368_3525_0, i_10_368_3555_0,
    i_10_368_3574_0, i_10_368_3583_0, i_10_368_3647_0, i_10_368_3703_0,
    i_10_368_3704_0, i_10_368_3707_0, i_10_368_3783_0, i_10_368_3785_0,
    i_10_368_3817_0, i_10_368_3857_0, i_10_368_3871_0, i_10_368_3909_0,
    i_10_368_3910_0, i_10_368_4140_0, i_10_368_4177_0, i_10_368_4270_0,
    i_10_368_4284_0, i_10_368_4307_0, i_10_368_4431_0, i_10_368_4582_0;
  output o_10_368_0_0;
  assign o_10_368_0_0 = 0;
endmodule



// Benchmark "kernel_10_369" written by ABC on Sun Jul 19 10:27:27 2020

module kernel_10_369 ( 
    i_10_369_263_0, i_10_369_271_0, i_10_369_286_0, i_10_369_326_0,
    i_10_369_412_0, i_10_369_424_0, i_10_369_425_0, i_10_369_427_0,
    i_10_369_464_0, i_10_369_640_0, i_10_369_712_0, i_10_369_1082_0,
    i_10_369_1084_0, i_10_369_1136_0, i_10_369_1238_0, i_10_369_1241_0,
    i_10_369_1305_0, i_10_369_1306_0, i_10_369_1309_0, i_10_369_1310_0,
    i_10_369_1313_0, i_10_369_1445_0, i_10_369_1543_0, i_10_369_1549_0,
    i_10_369_1550_0, i_10_369_1603_0, i_10_369_1648_0, i_10_369_1650_0,
    i_10_369_1651_0, i_10_369_1654_0, i_10_369_1685_0, i_10_369_1687_0,
    i_10_369_1690_0, i_10_369_1818_0, i_10_369_1819_0, i_10_369_1825_0,
    i_10_369_1994_0, i_10_369_2306_0, i_10_369_2349_0, i_10_369_2350_0,
    i_10_369_2362_0, i_10_369_2363_0, i_10_369_2377_0, i_10_369_2407_0,
    i_10_369_2448_0, i_10_369_2629_0, i_10_369_2630_0, i_10_369_2705_0,
    i_10_369_2710_0, i_10_369_2711_0, i_10_369_2827_0, i_10_369_2828_0,
    i_10_369_2832_0, i_10_369_2884_0, i_10_369_2888_0, i_10_369_2919_0,
    i_10_369_2920_0, i_10_369_2921_0, i_10_369_2922_0, i_10_369_2980_0,
    i_10_369_3033_0, i_10_369_3092_0, i_10_369_3152_0, i_10_369_3277_0,
    i_10_369_3386_0, i_10_369_3388_0, i_10_369_3403_0, i_10_369_3404_0,
    i_10_369_3523_0, i_10_369_3547_0, i_10_369_3613_0, i_10_369_3617_0,
    i_10_369_3646_0, i_10_369_3649_0, i_10_369_3787_0, i_10_369_3834_0,
    i_10_369_3841_0, i_10_369_3847_0, i_10_369_3851_0, i_10_369_3852_0,
    i_10_369_3853_0, i_10_369_3854_0, i_10_369_3857_0, i_10_369_3890_0,
    i_10_369_3982_0, i_10_369_3990_0, i_10_369_4121_0, i_10_369_4122_0,
    i_10_369_4123_0, i_10_369_4189_0, i_10_369_4231_0, i_10_369_4270_0,
    i_10_369_4271_0, i_10_369_4285_0, i_10_369_4286_0, i_10_369_4287_0,
    i_10_369_4288_0, i_10_369_4567_0, i_10_369_4568_0, i_10_369_4592_0,
    o_10_369_0_0  );
  input  i_10_369_263_0, i_10_369_271_0, i_10_369_286_0, i_10_369_326_0,
    i_10_369_412_0, i_10_369_424_0, i_10_369_425_0, i_10_369_427_0,
    i_10_369_464_0, i_10_369_640_0, i_10_369_712_0, i_10_369_1082_0,
    i_10_369_1084_0, i_10_369_1136_0, i_10_369_1238_0, i_10_369_1241_0,
    i_10_369_1305_0, i_10_369_1306_0, i_10_369_1309_0, i_10_369_1310_0,
    i_10_369_1313_0, i_10_369_1445_0, i_10_369_1543_0, i_10_369_1549_0,
    i_10_369_1550_0, i_10_369_1603_0, i_10_369_1648_0, i_10_369_1650_0,
    i_10_369_1651_0, i_10_369_1654_0, i_10_369_1685_0, i_10_369_1687_0,
    i_10_369_1690_0, i_10_369_1818_0, i_10_369_1819_0, i_10_369_1825_0,
    i_10_369_1994_0, i_10_369_2306_0, i_10_369_2349_0, i_10_369_2350_0,
    i_10_369_2362_0, i_10_369_2363_0, i_10_369_2377_0, i_10_369_2407_0,
    i_10_369_2448_0, i_10_369_2629_0, i_10_369_2630_0, i_10_369_2705_0,
    i_10_369_2710_0, i_10_369_2711_0, i_10_369_2827_0, i_10_369_2828_0,
    i_10_369_2832_0, i_10_369_2884_0, i_10_369_2888_0, i_10_369_2919_0,
    i_10_369_2920_0, i_10_369_2921_0, i_10_369_2922_0, i_10_369_2980_0,
    i_10_369_3033_0, i_10_369_3092_0, i_10_369_3152_0, i_10_369_3277_0,
    i_10_369_3386_0, i_10_369_3388_0, i_10_369_3403_0, i_10_369_3404_0,
    i_10_369_3523_0, i_10_369_3547_0, i_10_369_3613_0, i_10_369_3617_0,
    i_10_369_3646_0, i_10_369_3649_0, i_10_369_3787_0, i_10_369_3834_0,
    i_10_369_3841_0, i_10_369_3847_0, i_10_369_3851_0, i_10_369_3852_0,
    i_10_369_3853_0, i_10_369_3854_0, i_10_369_3857_0, i_10_369_3890_0,
    i_10_369_3982_0, i_10_369_3990_0, i_10_369_4121_0, i_10_369_4122_0,
    i_10_369_4123_0, i_10_369_4189_0, i_10_369_4231_0, i_10_369_4270_0,
    i_10_369_4271_0, i_10_369_4285_0, i_10_369_4286_0, i_10_369_4287_0,
    i_10_369_4288_0, i_10_369_4567_0, i_10_369_4568_0, i_10_369_4592_0;
  output o_10_369_0_0;
  assign o_10_369_0_0 = ~((~i_10_369_4287_0 & ((~i_10_369_326_0 & ((~i_10_369_427_0 & ~i_10_369_1238_0 & i_10_369_2350_0 & ~i_10_369_2710_0 & ~i_10_369_3523_0 & ~i_10_369_3834_0) | (i_10_369_1651_0 & i_10_369_1654_0 & ~i_10_369_2349_0 & ~i_10_369_2888_0 & ~i_10_369_3982_0 & ~i_10_369_4123_0 & ~i_10_369_4288_0))) | (~i_10_369_425_0 & ~i_10_369_2710_0 & ((~i_10_369_427_0 & ~i_10_369_1543_0 & ~i_10_369_2921_0 & ~i_10_369_3523_0 & ~i_10_369_4270_0) | (~i_10_369_1994_0 & ~i_10_369_3404_0 & ~i_10_369_3847_0 & ~i_10_369_3851_0 & ~i_10_369_4288_0))) | (~i_10_369_3851_0 & ((i_10_369_1651_0 & ~i_10_369_2362_0 & ~i_10_369_2921_0 & ~i_10_369_3033_0 & ~i_10_369_4285_0) | (i_10_369_1241_0 & ~i_10_369_2711_0 & ~i_10_369_4286_0))))) | (~i_10_369_640_0 & ((i_10_369_1651_0 & ~i_10_369_1818_0 & ~i_10_369_2705_0 & i_10_369_2921_0 & i_10_369_4271_0) | (~i_10_369_427_0 & ~i_10_369_712_0 & ~i_10_369_2629_0 & ~i_10_369_2919_0 & ~i_10_369_3404_0 & ~i_10_369_4285_0 & ~i_10_369_4567_0))) | (~i_10_369_1238_0 & ((~i_10_369_424_0 & ~i_10_369_464_0 & ~i_10_369_1445_0 & ~i_10_369_1543_0 & i_10_369_1651_0 & ~i_10_369_1687_0 & ~i_10_369_1690_0 & ~i_10_369_2362_0 & ~i_10_369_3890_0) | (i_10_369_1241_0 & ~i_10_369_4288_0))) | (~i_10_369_425_0 & ((~i_10_369_424_0 & ((i_10_369_1306_0 & ~i_10_369_2921_0 & ~i_10_369_3092_0) | (~i_10_369_286_0 & ~i_10_369_1445_0 & i_10_369_1818_0 & ~i_10_369_2884_0 & ~i_10_369_3403_0 & ~i_10_369_3834_0 & ~i_10_369_3854_0))) | (~i_10_369_1445_0 & ((~i_10_369_427_0 & ~i_10_369_2363_0 & ~i_10_369_2711_0 & ~i_10_369_2919_0 & ~i_10_369_4288_0) | (~i_10_369_2306_0 & ~i_10_369_3092_0 & i_10_369_3386_0 & ~i_10_369_4122_0 & ~i_10_369_4286_0 & ~i_10_369_4567_0 & ~i_10_369_4568_0))))) | (~i_10_369_464_0 & ((~i_10_369_1241_0 & ~i_10_369_1654_0 & ~i_10_369_1685_0 & ~i_10_369_2362_0 & ~i_10_369_2711_0 & ~i_10_369_2980_0 & ~i_10_369_3388_0 & ~i_10_369_4122_0 & ~i_10_369_4285_0) | (~i_10_369_1550_0 & ~i_10_369_2710_0 & ~i_10_369_2832_0 & ~i_10_369_3386_0 & ~i_10_369_3403_0 & ~i_10_369_3841_0 & ~i_10_369_4567_0))) | (~i_10_369_4285_0 & ((~i_10_369_1654_0 & ~i_10_369_2629_0 & ((~i_10_369_1690_0 & i_10_369_1825_0 & ~i_10_369_2711_0 & ~i_10_369_3388_0) | (i_10_369_427_0 & ~i_10_369_3404_0 & ~i_10_369_3852_0 & i_10_369_4288_0 & ~i_10_369_4568_0))) | (~i_10_369_2350_0 & ~i_10_369_2705_0 & i_10_369_2710_0 & ~i_10_369_3386_0 & ~i_10_369_3403_0 & ~i_10_369_4567_0))) | (~i_10_369_1687_0 & ((~i_10_369_427_0 & i_10_369_464_0 & ~i_10_369_2919_0 & ~i_10_369_2920_0 & ~i_10_369_3388_0) | (~i_10_369_1549_0 & ~i_10_369_2363_0 & ~i_10_369_2710_0 & i_10_369_2920_0 & ~i_10_369_3404_0 & ~i_10_369_3547_0 & ~i_10_369_3787_0 & ~i_10_369_3834_0 & i_10_369_3847_0))) | (i_10_369_464_0 & ((~i_10_369_1445_0 & i_10_369_2705_0 & ~i_10_369_3403_0 & ~i_10_369_3613_0 & ~i_10_369_3787_0) | (~i_10_369_712_0 & ~i_10_369_1549_0 & ~i_10_369_1550_0 & ~i_10_369_2448_0 & ~i_10_369_2919_0 & ~i_10_369_4121_0 & ~i_10_369_4122_0 & ~i_10_369_4567_0))) | (~i_10_369_2377_0 & ((~i_10_369_1549_0 & ((i_10_369_1818_0 & i_10_369_2448_0 & ~i_10_369_2980_0 & ~i_10_369_3403_0 & ~i_10_369_3523_0) | (~i_10_369_427_0 & i_10_369_1819_0 & ~i_10_369_2630_0 & ~i_10_369_2919_0 & ~i_10_369_2921_0 & ~i_10_369_3857_0))) | (~i_10_369_1685_0 & ~i_10_369_2711_0 & i_10_369_3854_0) | (i_10_369_1310_0 & ~i_10_369_3277_0 & ~i_10_369_4231_0))) | (~i_10_369_3386_0 & ((i_10_369_2349_0 & ~i_10_369_2922_0 & i_10_369_3033_0) | (~i_10_369_427_0 & ~i_10_369_1543_0 & ~i_10_369_1550_0 & ~i_10_369_2363_0 & ~i_10_369_2920_0 & ~i_10_369_2921_0 & ~i_10_369_3033_0 & ~i_10_369_3847_0 & ~i_10_369_3890_0))) | (~i_10_369_427_0 & ((i_10_369_3649_0 & i_10_369_3847_0) | (~i_10_369_1550_0 & i_10_369_2350_0 & ~i_10_369_3523_0 & ~i_10_369_3982_0 & ~i_10_369_4123_0 & ~i_10_369_4568_0))) | (i_10_369_1650_0 & ~i_10_369_1690_0 & ~i_10_369_3404_0 & i_10_369_3852_0) | (~i_10_369_1550_0 & i_10_369_1648_0 & ~i_10_369_2710_0 & ~i_10_369_2711_0 & ~i_10_369_2884_0 & ~i_10_369_3851_0 & ~i_10_369_4231_0) | (i_10_369_1309_0 & ~i_10_369_1994_0 & ~i_10_369_2832_0 & ~i_10_369_2980_0 & ~i_10_369_4123_0 & ~i_10_369_4288_0));
endmodule



// Benchmark "kernel_10_370" written by ABC on Sun Jul 19 10:27:28 2020

module kernel_10_370 ( 
    i_10_370_39_0, i_10_370_48_0, i_10_370_171_0, i_10_370_174_0,
    i_10_370_175_0, i_10_370_193_0, i_10_370_247_0, i_10_370_249_0,
    i_10_370_289_0, i_10_370_318_0, i_10_370_327_0, i_10_370_330_0,
    i_10_370_364_0, i_10_370_405_0, i_10_370_406_0, i_10_370_412_0,
    i_10_370_435_0, i_10_370_520_0, i_10_370_594_0, i_10_370_633_0,
    i_10_370_793_0, i_10_370_832_0, i_10_370_877_0, i_10_370_1002_0,
    i_10_370_1155_0, i_10_370_1266_0, i_10_370_1270_0, i_10_370_1293_0,
    i_10_370_1306_0, i_10_370_1327_0, i_10_370_1329_0, i_10_370_1341_0,
    i_10_370_1344_0, i_10_370_1365_0, i_10_370_1366_0, i_10_370_1441_0,
    i_10_370_1576_0, i_10_370_1714_0, i_10_370_1825_0, i_10_370_1873_0,
    i_10_370_1878_0, i_10_370_1992_0, i_10_370_1996_0, i_10_370_2016_0,
    i_10_370_2020_0, i_10_370_2202_0, i_10_370_2241_0, i_10_370_2250_0,
    i_10_370_2317_0, i_10_370_2326_0, i_10_370_2352_0, i_10_370_2359_0,
    i_10_370_2364_0, i_10_370_2380_0, i_10_370_2406_0, i_10_370_2449_0,
    i_10_370_2473_0, i_10_370_2586_0, i_10_370_2604_0, i_10_370_2605_0,
    i_10_370_2608_0, i_10_370_2643_0, i_10_370_2676_0, i_10_370_2701_0,
    i_10_370_2704_0, i_10_370_2720_0, i_10_370_2721_0, i_10_370_2724_0,
    i_10_370_2782_0, i_10_370_2785_0, i_10_370_2786_0, i_10_370_2834_0,
    i_10_370_2881_0, i_10_370_2882_0, i_10_370_2994_0, i_10_370_3030_0,
    i_10_370_3075_0, i_10_370_3165_0, i_10_370_3198_0, i_10_370_3199_0,
    i_10_370_3273_0, i_10_370_3297_0, i_10_370_3300_0, i_10_370_3588_0,
    i_10_370_3589_0, i_10_370_3703_0, i_10_370_3714_0, i_10_370_3975_0,
    i_10_370_4126_0, i_10_370_4156_0, i_10_370_4233_0, i_10_370_4260_0,
    i_10_370_4273_0, i_10_370_4276_0, i_10_370_4378_0, i_10_370_4505_0,
    i_10_370_4522_0, i_10_370_4524_0, i_10_370_4581_0, i_10_370_4585_0,
    o_10_370_0_0  );
  input  i_10_370_39_0, i_10_370_48_0, i_10_370_171_0, i_10_370_174_0,
    i_10_370_175_0, i_10_370_193_0, i_10_370_247_0, i_10_370_249_0,
    i_10_370_289_0, i_10_370_318_0, i_10_370_327_0, i_10_370_330_0,
    i_10_370_364_0, i_10_370_405_0, i_10_370_406_0, i_10_370_412_0,
    i_10_370_435_0, i_10_370_520_0, i_10_370_594_0, i_10_370_633_0,
    i_10_370_793_0, i_10_370_832_0, i_10_370_877_0, i_10_370_1002_0,
    i_10_370_1155_0, i_10_370_1266_0, i_10_370_1270_0, i_10_370_1293_0,
    i_10_370_1306_0, i_10_370_1327_0, i_10_370_1329_0, i_10_370_1341_0,
    i_10_370_1344_0, i_10_370_1365_0, i_10_370_1366_0, i_10_370_1441_0,
    i_10_370_1576_0, i_10_370_1714_0, i_10_370_1825_0, i_10_370_1873_0,
    i_10_370_1878_0, i_10_370_1992_0, i_10_370_1996_0, i_10_370_2016_0,
    i_10_370_2020_0, i_10_370_2202_0, i_10_370_2241_0, i_10_370_2250_0,
    i_10_370_2317_0, i_10_370_2326_0, i_10_370_2352_0, i_10_370_2359_0,
    i_10_370_2364_0, i_10_370_2380_0, i_10_370_2406_0, i_10_370_2449_0,
    i_10_370_2473_0, i_10_370_2586_0, i_10_370_2604_0, i_10_370_2605_0,
    i_10_370_2608_0, i_10_370_2643_0, i_10_370_2676_0, i_10_370_2701_0,
    i_10_370_2704_0, i_10_370_2720_0, i_10_370_2721_0, i_10_370_2724_0,
    i_10_370_2782_0, i_10_370_2785_0, i_10_370_2786_0, i_10_370_2834_0,
    i_10_370_2881_0, i_10_370_2882_0, i_10_370_2994_0, i_10_370_3030_0,
    i_10_370_3075_0, i_10_370_3165_0, i_10_370_3198_0, i_10_370_3199_0,
    i_10_370_3273_0, i_10_370_3297_0, i_10_370_3300_0, i_10_370_3588_0,
    i_10_370_3589_0, i_10_370_3703_0, i_10_370_3714_0, i_10_370_3975_0,
    i_10_370_4126_0, i_10_370_4156_0, i_10_370_4233_0, i_10_370_4260_0,
    i_10_370_4273_0, i_10_370_4276_0, i_10_370_4378_0, i_10_370_4505_0,
    i_10_370_4522_0, i_10_370_4524_0, i_10_370_4581_0, i_10_370_4585_0;
  output o_10_370_0_0;
  assign o_10_370_0_0 = 0;
endmodule



// Benchmark "kernel_10_371" written by ABC on Sun Jul 19 10:27:29 2020

module kernel_10_371 ( 
    i_10_371_156_0, i_10_371_220_0, i_10_371_249_0, i_10_371_279_0,
    i_10_371_390_0, i_10_371_391_0, i_10_371_423_0, i_10_371_441_0,
    i_10_371_447_0, i_10_371_459_0, i_10_371_513_0, i_10_371_516_0,
    i_10_371_519_0, i_10_371_600_0, i_10_371_636_0, i_10_371_637_0,
    i_10_371_718_0, i_10_371_795_0, i_10_371_796_0, i_10_371_898_0,
    i_10_371_1087_0, i_10_371_1122_0, i_10_371_1248_0, i_10_371_1306_0,
    i_10_371_1307_0, i_10_371_1308_0, i_10_371_1339_0, i_10_371_1359_0,
    i_10_371_1377_0, i_10_371_1485_0, i_10_371_1486_0, i_10_371_1541_0,
    i_10_371_1642_0, i_10_371_1683_0, i_10_371_1684_0, i_10_371_1685_0,
    i_10_371_1824_0, i_10_371_1915_0, i_10_371_1950_0, i_10_371_2061_0,
    i_10_371_2185_0, i_10_371_2247_0, i_10_371_2384_0, i_10_371_2391_0,
    i_10_371_2451_0, i_10_371_2452_0, i_10_371_2468_0, i_10_371_2562_0,
    i_10_371_2634_0, i_10_371_2679_0, i_10_371_2715_0, i_10_371_2718_0,
    i_10_371_2719_0, i_10_371_2721_0, i_10_371_2727_0, i_10_371_2742_0,
    i_10_371_2743_0, i_10_371_2781_0, i_10_371_2785_0, i_10_371_2786_0,
    i_10_371_2832_0, i_10_371_2833_0, i_10_371_2916_0, i_10_371_2919_0,
    i_10_371_2982_0, i_10_371_3047_0, i_10_371_3201_0, i_10_371_3234_0,
    i_10_371_3237_0, i_10_371_3276_0, i_10_371_3279_0, i_10_371_3312_0,
    i_10_371_3390_0, i_10_371_3468_0, i_10_371_3471_0, i_10_371_3472_0,
    i_10_371_3495_0, i_10_371_3519_0, i_10_371_3522_0, i_10_371_3525_0,
    i_10_371_3586_0, i_10_371_3589_0, i_10_371_3590_0, i_10_371_3834_0,
    i_10_371_3841_0, i_10_371_3844_0, i_10_371_3853_0, i_10_371_3858_0,
    i_10_371_3877_0, i_10_371_3906_0, i_10_371_3949_0, i_10_371_3985_0,
    i_10_371_4114_0, i_10_371_4228_0, i_10_371_4229_0, i_10_371_4271_0,
    i_10_371_4287_0, i_10_371_4317_0, i_10_371_4318_0, i_10_371_4588_0,
    o_10_371_0_0  );
  input  i_10_371_156_0, i_10_371_220_0, i_10_371_249_0, i_10_371_279_0,
    i_10_371_390_0, i_10_371_391_0, i_10_371_423_0, i_10_371_441_0,
    i_10_371_447_0, i_10_371_459_0, i_10_371_513_0, i_10_371_516_0,
    i_10_371_519_0, i_10_371_600_0, i_10_371_636_0, i_10_371_637_0,
    i_10_371_718_0, i_10_371_795_0, i_10_371_796_0, i_10_371_898_0,
    i_10_371_1087_0, i_10_371_1122_0, i_10_371_1248_0, i_10_371_1306_0,
    i_10_371_1307_0, i_10_371_1308_0, i_10_371_1339_0, i_10_371_1359_0,
    i_10_371_1377_0, i_10_371_1485_0, i_10_371_1486_0, i_10_371_1541_0,
    i_10_371_1642_0, i_10_371_1683_0, i_10_371_1684_0, i_10_371_1685_0,
    i_10_371_1824_0, i_10_371_1915_0, i_10_371_1950_0, i_10_371_2061_0,
    i_10_371_2185_0, i_10_371_2247_0, i_10_371_2384_0, i_10_371_2391_0,
    i_10_371_2451_0, i_10_371_2452_0, i_10_371_2468_0, i_10_371_2562_0,
    i_10_371_2634_0, i_10_371_2679_0, i_10_371_2715_0, i_10_371_2718_0,
    i_10_371_2719_0, i_10_371_2721_0, i_10_371_2727_0, i_10_371_2742_0,
    i_10_371_2743_0, i_10_371_2781_0, i_10_371_2785_0, i_10_371_2786_0,
    i_10_371_2832_0, i_10_371_2833_0, i_10_371_2916_0, i_10_371_2919_0,
    i_10_371_2982_0, i_10_371_3047_0, i_10_371_3201_0, i_10_371_3234_0,
    i_10_371_3237_0, i_10_371_3276_0, i_10_371_3279_0, i_10_371_3312_0,
    i_10_371_3390_0, i_10_371_3468_0, i_10_371_3471_0, i_10_371_3472_0,
    i_10_371_3495_0, i_10_371_3519_0, i_10_371_3522_0, i_10_371_3525_0,
    i_10_371_3586_0, i_10_371_3589_0, i_10_371_3590_0, i_10_371_3834_0,
    i_10_371_3841_0, i_10_371_3844_0, i_10_371_3853_0, i_10_371_3858_0,
    i_10_371_3877_0, i_10_371_3906_0, i_10_371_3949_0, i_10_371_3985_0,
    i_10_371_4114_0, i_10_371_4228_0, i_10_371_4229_0, i_10_371_4271_0,
    i_10_371_4287_0, i_10_371_4317_0, i_10_371_4318_0, i_10_371_4588_0;
  output o_10_371_0_0;
  assign o_10_371_0_0 = ~((~i_10_371_279_0 & ((i_10_371_3276_0 & ~i_10_371_3312_0 & ~i_10_371_3906_0 & ~i_10_371_4114_0) | (~i_10_371_447_0 & ~i_10_371_1486_0 & ~i_10_371_2468_0 & ~i_10_371_2715_0 & ~i_10_371_2727_0 & ~i_10_371_3841_0 & i_10_371_4287_0))) | (~i_10_371_513_0 & ((~i_10_371_2452_0 & ~i_10_371_2719_0 & ~i_10_371_3234_0 & ~i_10_371_3495_0 & ~i_10_371_3844_0 & i_10_371_4271_0) | (~i_10_371_447_0 & ~i_10_371_1359_0 & ~i_10_371_3841_0 & ~i_10_371_3853_0 & i_10_371_4287_0))) | (~i_10_371_447_0 & ((~i_10_371_423_0 & i_10_371_1308_0 & ~i_10_371_2468_0) | (~i_10_371_1485_0 & ~i_10_371_2719_0 & ~i_10_371_3390_0 & ~i_10_371_4287_0))) | (~i_10_371_423_0 & ((~i_10_371_1248_0 & ~i_10_371_1684_0 & ~i_10_371_2727_0 & i_10_371_2832_0 & i_10_371_2833_0) | (~i_10_371_441_0 & ~i_10_371_1824_0 & ~i_10_371_2634_0 & ~i_10_371_4287_0))) | (~i_10_371_795_0 & ((~i_10_371_898_0 & ~i_10_371_2452_0) | (~i_10_371_796_0 & i_10_371_1950_0 & ~i_10_371_2727_0))) | (~i_10_371_898_0 & ~i_10_371_2384_0 & ((~i_10_371_516_0 & ~i_10_371_1359_0 & ~i_10_371_2451_0 & ~i_10_371_3906_0) | (~i_10_371_1684_0 & ~i_10_371_2781_0 & ~i_10_371_3237_0 & ~i_10_371_3841_0 & ~i_10_371_4287_0))) | (~i_10_371_516_0 & ((~i_10_371_718_0 & ~i_10_371_1683_0 & ~i_10_371_2451_0 & ~i_10_371_3237_0 & ~i_10_371_3279_0 & ~i_10_371_3589_0) | (i_10_371_3201_0 & ~i_10_371_4287_0))) | (~i_10_371_1248_0 & ((i_10_371_459_0 & i_10_371_1307_0 & ~i_10_371_1485_0 & ~i_10_371_1824_0) | (i_10_371_279_0 & ~i_10_371_1359_0 & ~i_10_371_1684_0 & ~i_10_371_1685_0 & ~i_10_371_2833_0 & ~i_10_371_3906_0 & ~i_10_371_3949_0))) | (~i_10_371_2721_0 & ((~i_10_371_1359_0 & ((~i_10_371_2727_0 & ~i_10_371_3234_0 & ~i_10_371_3237_0 & ~i_10_371_3586_0 & ~i_10_371_3589_0) | (~i_10_371_3312_0 & ~i_10_371_3468_0 & ~i_10_371_3590_0 & ~i_10_371_4287_0))) | (~i_10_371_1684_0 & ~i_10_371_2715_0 & ~i_10_371_2916_0 & ~i_10_371_2919_0))) | (~i_10_371_2916_0 & ~i_10_371_3237_0 & ((~i_10_371_220_0 & ~i_10_371_1685_0 & ~i_10_371_2919_0 & ~i_10_371_3312_0 & ~i_10_371_3495_0 & ~i_10_371_3525_0) | (~i_10_371_1308_0 & ~i_10_371_1485_0 & ~i_10_371_2833_0 & ~i_10_371_3234_0 & ~i_10_371_3390_0 & ~i_10_371_3519_0 & ~i_10_371_4271_0))) | (i_10_371_3853_0 & ((~i_10_371_1950_0 & ~i_10_371_2718_0 & i_10_371_2919_0 & i_10_371_3858_0) | (~i_10_371_2452_0 & i_10_371_4271_0))) | (i_10_371_1950_0 & i_10_371_2384_0 & ~i_10_371_3834_0) | (~i_10_371_2715_0 & ~i_10_371_2727_0 & ~i_10_371_3276_0 & ~i_10_371_4287_0));
endmodule



// Benchmark "kernel_10_372" written by ABC on Sun Jul 19 10:27:30 2020

module kernel_10_372 ( 
    i_10_372_40_0, i_10_372_43_0, i_10_372_176_0, i_10_372_257_0,
    i_10_372_266_0, i_10_372_269_0, i_10_372_323_0, i_10_372_374_0,
    i_10_372_394_0, i_10_372_395_0, i_10_372_410_0, i_10_372_413_0,
    i_10_372_439_0, i_10_372_440_0, i_10_372_449_0, i_10_372_640_0,
    i_10_372_743_0, i_10_372_797_0, i_10_372_1004_0, i_10_372_1007_0,
    i_10_372_1034_0, i_10_372_1042_0, i_10_372_1222_0, i_10_372_1223_0,
    i_10_372_1235_0, i_10_372_1237_0, i_10_372_1238_0, i_10_372_1240_0,
    i_10_372_1303_0, i_10_372_1308_0, i_10_372_1310_0, i_10_372_1366_0,
    i_10_372_1385_0, i_10_372_1435_0, i_10_372_1436_0, i_10_372_1439_0,
    i_10_372_1544_0, i_10_372_1552_0, i_10_372_1612_0, i_10_372_1717_0,
    i_10_372_1736_0, i_10_372_1823_0, i_10_372_1916_0, i_10_372_1919_0,
    i_10_372_1956_0, i_10_372_1988_0, i_10_372_2006_0, i_10_372_2023_0,
    i_10_372_2029_0, i_10_372_2033_0, i_10_372_2204_0, i_10_372_2312_0,
    i_10_372_2348_0, i_10_372_2354_0, i_10_372_2608_0, i_10_372_2633_0,
    i_10_372_2635_0, i_10_372_2636_0, i_10_372_2735_0, i_10_372_2761_0,
    i_10_372_2786_0, i_10_372_2789_0, i_10_372_2830_0, i_10_372_2843_0,
    i_10_372_2870_0, i_10_372_2966_0, i_10_372_3024_0, i_10_372_3040_0,
    i_10_372_3049_0, i_10_372_3050_0, i_10_372_3074_0, i_10_372_3077_0,
    i_10_372_3391_0, i_10_372_3392_0, i_10_372_3473_0, i_10_372_3506_0,
    i_10_372_3563_0, i_10_372_3584_0, i_10_372_3586_0, i_10_372_3587_0,
    i_10_372_3589_0, i_10_372_3590_0, i_10_372_3612_0, i_10_372_3721_0,
    i_10_372_3722_0, i_10_372_3734_0, i_10_372_3854_0, i_10_372_3860_0,
    i_10_372_3986_0, i_10_372_4004_0, i_10_372_4161_0, i_10_372_4175_0,
    i_10_372_4210_0, i_10_372_4211_0, i_10_372_4217_0, i_10_372_4268_0,
    i_10_372_4271_0, i_10_372_4273_0, i_10_372_4489_0, i_10_372_4535_0,
    o_10_372_0_0  );
  input  i_10_372_40_0, i_10_372_43_0, i_10_372_176_0, i_10_372_257_0,
    i_10_372_266_0, i_10_372_269_0, i_10_372_323_0, i_10_372_374_0,
    i_10_372_394_0, i_10_372_395_0, i_10_372_410_0, i_10_372_413_0,
    i_10_372_439_0, i_10_372_440_0, i_10_372_449_0, i_10_372_640_0,
    i_10_372_743_0, i_10_372_797_0, i_10_372_1004_0, i_10_372_1007_0,
    i_10_372_1034_0, i_10_372_1042_0, i_10_372_1222_0, i_10_372_1223_0,
    i_10_372_1235_0, i_10_372_1237_0, i_10_372_1238_0, i_10_372_1240_0,
    i_10_372_1303_0, i_10_372_1308_0, i_10_372_1310_0, i_10_372_1366_0,
    i_10_372_1385_0, i_10_372_1435_0, i_10_372_1436_0, i_10_372_1439_0,
    i_10_372_1544_0, i_10_372_1552_0, i_10_372_1612_0, i_10_372_1717_0,
    i_10_372_1736_0, i_10_372_1823_0, i_10_372_1916_0, i_10_372_1919_0,
    i_10_372_1956_0, i_10_372_1988_0, i_10_372_2006_0, i_10_372_2023_0,
    i_10_372_2029_0, i_10_372_2033_0, i_10_372_2204_0, i_10_372_2312_0,
    i_10_372_2348_0, i_10_372_2354_0, i_10_372_2608_0, i_10_372_2633_0,
    i_10_372_2635_0, i_10_372_2636_0, i_10_372_2735_0, i_10_372_2761_0,
    i_10_372_2786_0, i_10_372_2789_0, i_10_372_2830_0, i_10_372_2843_0,
    i_10_372_2870_0, i_10_372_2966_0, i_10_372_3024_0, i_10_372_3040_0,
    i_10_372_3049_0, i_10_372_3050_0, i_10_372_3074_0, i_10_372_3077_0,
    i_10_372_3391_0, i_10_372_3392_0, i_10_372_3473_0, i_10_372_3506_0,
    i_10_372_3563_0, i_10_372_3584_0, i_10_372_3586_0, i_10_372_3587_0,
    i_10_372_3589_0, i_10_372_3590_0, i_10_372_3612_0, i_10_372_3721_0,
    i_10_372_3722_0, i_10_372_3734_0, i_10_372_3854_0, i_10_372_3860_0,
    i_10_372_3986_0, i_10_372_4004_0, i_10_372_4161_0, i_10_372_4175_0,
    i_10_372_4210_0, i_10_372_4211_0, i_10_372_4217_0, i_10_372_4268_0,
    i_10_372_4271_0, i_10_372_4273_0, i_10_372_4489_0, i_10_372_4535_0;
  output o_10_372_0_0;
  assign o_10_372_0_0 = 0;
endmodule



// Benchmark "kernel_10_373" written by ABC on Sun Jul 19 10:27:31 2020

module kernel_10_373 ( 
    i_10_373_150_0, i_10_373_176_0, i_10_373_390_0, i_10_373_394_0,
    i_10_373_395_0, i_10_373_409_0, i_10_373_412_0, i_10_373_429_0,
    i_10_373_430_0, i_10_373_431_0, i_10_373_445_0, i_10_373_448_0,
    i_10_373_457_0, i_10_373_460_0, i_10_373_505_0, i_10_373_508_0,
    i_10_373_717_0, i_10_373_796_0, i_10_373_799_0, i_10_373_907_0,
    i_10_373_908_0, i_10_373_957_0, i_10_373_966_0, i_10_373_967_0,
    i_10_373_1005_0, i_10_373_1307_0, i_10_373_1312_0, i_10_373_1313_0,
    i_10_373_1583_0, i_10_373_1652_0, i_10_373_1653_0, i_10_373_1655_0,
    i_10_373_1689_0, i_10_373_1690_0, i_10_373_1823_0, i_10_373_1826_0,
    i_10_373_1995_0, i_10_373_2033_0, i_10_373_2351_0, i_10_373_2365_0,
    i_10_373_2407_0, i_10_373_2451_0, i_10_373_2452_0, i_10_373_2453_0,
    i_10_373_2455_0, i_10_373_2469_0, i_10_373_2472_0, i_10_373_2473_0,
    i_10_373_2636_0, i_10_373_2659_0, i_10_373_2660_0, i_10_373_2703_0,
    i_10_373_2704_0, i_10_373_2706_0, i_10_373_2707_0, i_10_373_2708_0,
    i_10_373_2786_0, i_10_373_2788_0, i_10_373_2789_0, i_10_373_2824_0,
    i_10_373_2830_0, i_10_373_2833_0, i_10_373_2922_0, i_10_373_2923_0,
    i_10_373_3071_0, i_10_373_3157_0, i_10_373_3158_0, i_10_373_3196_0,
    i_10_373_3197_0, i_10_373_3272_0, i_10_373_3283_0, i_10_373_3284_0,
    i_10_373_3315_0, i_10_373_3328_0, i_10_373_3329_0, i_10_373_3388_0,
    i_10_373_3391_0, i_10_373_3392_0, i_10_373_3468_0, i_10_373_3469_0,
    i_10_373_3470_0, i_10_373_3542_0, i_10_373_3544_0, i_10_373_3545_0,
    i_10_373_3589_0, i_10_373_3613_0, i_10_373_3787_0, i_10_373_3837_0,
    i_10_373_3840_0, i_10_373_3846_0, i_10_373_3847_0, i_10_373_3859_0,
    i_10_373_3860_0, i_10_373_4057_0, i_10_373_4121_0, i_10_373_4129_0,
    i_10_373_4270_0, i_10_373_4274_0, i_10_373_4287_0, i_10_373_4292_0,
    o_10_373_0_0  );
  input  i_10_373_150_0, i_10_373_176_0, i_10_373_390_0, i_10_373_394_0,
    i_10_373_395_0, i_10_373_409_0, i_10_373_412_0, i_10_373_429_0,
    i_10_373_430_0, i_10_373_431_0, i_10_373_445_0, i_10_373_448_0,
    i_10_373_457_0, i_10_373_460_0, i_10_373_505_0, i_10_373_508_0,
    i_10_373_717_0, i_10_373_796_0, i_10_373_799_0, i_10_373_907_0,
    i_10_373_908_0, i_10_373_957_0, i_10_373_966_0, i_10_373_967_0,
    i_10_373_1005_0, i_10_373_1307_0, i_10_373_1312_0, i_10_373_1313_0,
    i_10_373_1583_0, i_10_373_1652_0, i_10_373_1653_0, i_10_373_1655_0,
    i_10_373_1689_0, i_10_373_1690_0, i_10_373_1823_0, i_10_373_1826_0,
    i_10_373_1995_0, i_10_373_2033_0, i_10_373_2351_0, i_10_373_2365_0,
    i_10_373_2407_0, i_10_373_2451_0, i_10_373_2452_0, i_10_373_2453_0,
    i_10_373_2455_0, i_10_373_2469_0, i_10_373_2472_0, i_10_373_2473_0,
    i_10_373_2636_0, i_10_373_2659_0, i_10_373_2660_0, i_10_373_2703_0,
    i_10_373_2704_0, i_10_373_2706_0, i_10_373_2707_0, i_10_373_2708_0,
    i_10_373_2786_0, i_10_373_2788_0, i_10_373_2789_0, i_10_373_2824_0,
    i_10_373_2830_0, i_10_373_2833_0, i_10_373_2922_0, i_10_373_2923_0,
    i_10_373_3071_0, i_10_373_3157_0, i_10_373_3158_0, i_10_373_3196_0,
    i_10_373_3197_0, i_10_373_3272_0, i_10_373_3283_0, i_10_373_3284_0,
    i_10_373_3315_0, i_10_373_3328_0, i_10_373_3329_0, i_10_373_3388_0,
    i_10_373_3391_0, i_10_373_3392_0, i_10_373_3468_0, i_10_373_3469_0,
    i_10_373_3470_0, i_10_373_3542_0, i_10_373_3544_0, i_10_373_3545_0,
    i_10_373_3589_0, i_10_373_3613_0, i_10_373_3787_0, i_10_373_3837_0,
    i_10_373_3840_0, i_10_373_3846_0, i_10_373_3847_0, i_10_373_3859_0,
    i_10_373_3860_0, i_10_373_4057_0, i_10_373_4121_0, i_10_373_4129_0,
    i_10_373_4270_0, i_10_373_4274_0, i_10_373_4287_0, i_10_373_4292_0;
  output o_10_373_0_0;
  assign o_10_373_0_0 = ~((~i_10_373_445_0 & ((~i_10_373_429_0 & i_10_373_796_0 & ~i_10_373_3284_0 & ~i_10_373_3315_0 & ~i_10_373_3470_0 & ~i_10_373_3542_0 & ~i_10_373_4270_0) | (~i_10_373_799_0 & ~i_10_373_1312_0 & ~i_10_373_1583_0 & ~i_10_373_1689_0 & ~i_10_373_1823_0 & ~i_10_373_2472_0 & ~i_10_373_2833_0 & ~i_10_373_3469_0 & ~i_10_373_4287_0 & ~i_10_373_4292_0))) | (~i_10_373_430_0 & ((~i_10_373_966_0 & ((~i_10_373_390_0 & ~i_10_373_431_0 & ((~i_10_373_429_0 & ~i_10_373_1652_0 & ~i_10_373_1689_0 & ~i_10_373_1690_0 & ~i_10_373_2451_0 & ~i_10_373_2452_0 & ~i_10_373_3283_0 & ~i_10_373_3542_0 & ~i_10_373_3544_0 & ~i_10_373_3846_0) | (~i_10_373_150_0 & ~i_10_373_394_0 & ~i_10_373_460_0 & ~i_10_373_967_0 & ~i_10_373_1005_0 & ~i_10_373_1313_0 & ~i_10_373_1995_0 & ~i_10_373_2833_0 & ~i_10_373_3315_0 & ~i_10_373_3469_0 & ~i_10_373_3470_0 & ~i_10_373_3859_0 & ~i_10_373_4274_0))) | (~i_10_373_3468_0 & ((~i_10_373_717_0 & ~i_10_373_908_0 & ~i_10_373_1583_0 & ~i_10_373_2452_0 & i_10_373_3859_0) | (~i_10_373_395_0 & ~i_10_373_457_0 & ~i_10_373_1690_0 & ~i_10_373_2407_0 & ~i_10_373_2455_0 & ~i_10_373_3071_0 & ~i_10_373_3388_0 & ~i_10_373_3392_0 & ~i_10_373_3787_0 & ~i_10_373_3846_0 & ~i_10_373_4287_0))))) | (~i_10_373_460_0 & ~i_10_373_957_0 & ~i_10_373_1312_0 & ~i_10_373_1823_0 & i_10_373_2452_0 & ~i_10_373_3284_0 & ~i_10_373_3392_0 & ~i_10_373_3544_0) | (~i_10_373_717_0 & ~i_10_373_1307_0 & ~i_10_373_2473_0 & i_10_373_2636_0 & ~i_10_373_3470_0 & ~i_10_373_3545_0 & ~i_10_373_3589_0))) | (~i_10_373_429_0 & ((~i_10_373_390_0 & ~i_10_373_394_0 & ~i_10_373_395_0 & ~i_10_373_957_0 & ~i_10_373_2033_0 & ~i_10_373_2351_0 & i_10_373_2452_0 & i_10_373_2453_0 & ~i_10_373_3388_0) | (~i_10_373_448_0 & ~i_10_373_967_0 & i_10_373_1312_0 & ~i_10_373_2469_0 & ~i_10_373_3391_0 & ~i_10_373_3469_0 & ~i_10_373_3470_0 & ~i_10_373_3542_0 & ~i_10_373_4292_0))) | (~i_10_373_431_0 & ((~i_10_373_390_0 & ~i_10_373_2469_0 & ~i_10_373_2786_0 & ~i_10_373_2824_0 & i_10_373_2922_0 & ~i_10_373_3589_0 & ~i_10_373_3846_0 & ~i_10_373_4121_0) | (i_10_373_1655_0 & ~i_10_373_2472_0 & ~i_10_373_3283_0 & ~i_10_373_3542_0 & ~i_10_373_4057_0 & ~i_10_373_4274_0))) | (~i_10_373_796_0 & ((~i_10_373_390_0 & ~i_10_373_966_0 & i_10_373_1823_0 & ~i_10_373_3284_0 & ~i_10_373_3392_0 & ~i_10_373_3542_0 & ~i_10_373_3589_0 & ~i_10_373_3613_0) | (~i_10_373_799_0 & ~i_10_373_1690_0 & ~i_10_373_2473_0 & i_10_373_3197_0 & ~i_10_373_3545_0 & ~i_10_373_3787_0))) | (~i_10_373_150_0 & ((~i_10_373_2469_0 & ((~i_10_373_395_0 & ~i_10_373_3468_0 & ((~i_10_373_907_0 & ~i_10_373_967_0 & ~i_10_373_3196_0 & ~i_10_373_3283_0 & ~i_10_373_3469_0 & ~i_10_373_3470_0 & ~i_10_373_3613_0) | (~i_10_373_966_0 & ~i_10_373_2472_0 & ~i_10_373_2824_0 & ~i_10_373_3284_0 & ~i_10_373_3388_0 & ~i_10_373_4121_0 & ~i_10_373_4270_0))) | (~i_10_373_390_0 & ~i_10_373_2033_0 & ~i_10_373_2472_0 & ~i_10_373_3388_0 & ~i_10_373_3470_0 & i_10_373_3837_0 & ~i_10_373_3840_0))) | (~i_10_373_907_0 & ~i_10_373_967_0 & i_10_373_1655_0 & ~i_10_373_3315_0 & ~i_10_373_3468_0 & ~i_10_373_3542_0 & ~i_10_373_3545_0) | (~i_10_373_966_0 & ~i_10_373_1690_0 & i_10_373_2703_0 & ~i_10_373_3388_0 & ~i_10_373_3787_0 & ~i_10_373_3847_0 & ~i_10_373_4057_0) | (~i_10_373_394_0 & ~i_10_373_1689_0 & i_10_373_1826_0 & ~i_10_373_2351_0 & ~i_10_373_3469_0 & ~i_10_373_4129_0 & ~i_10_373_4292_0))) | (~i_10_373_460_0 & ((~i_10_373_394_0 & ((~i_10_373_2472_0 & i_10_373_2703_0 & i_10_373_2704_0 & ~i_10_373_3391_0) | (i_10_373_390_0 & ~i_10_373_957_0 & ~i_10_373_2455_0 & ~i_10_373_2469_0 & ~i_10_373_3846_0))) | (i_10_373_1312_0 & i_10_373_2469_0 & ~i_10_373_2472_0 & ~i_10_373_3589_0))) | (~i_10_373_3837_0 & ((i_10_373_1823_0 & ~i_10_373_2469_0 & ~i_10_373_4287_0 & ((i_10_373_1826_0 & ~i_10_373_2033_0 & ~i_10_373_3284_0) | (~i_10_373_2351_0 & ~i_10_373_3470_0 & ~i_10_373_3589_0 & ~i_10_373_3846_0 & ~i_10_373_3847_0))) | (i_10_373_3272_0 & ~i_10_373_3392_0 & ~i_10_373_3847_0) | (~i_10_373_967_0 & ~i_10_373_3196_0 & ~i_10_373_3283_0 & ~i_10_373_3388_0 & ~i_10_373_3859_0 & i_10_373_4287_0))) | (~i_10_373_390_0 & ~i_10_373_3542_0 & ((~i_10_373_967_0 & ~i_10_373_3315_0 & ((~i_10_373_395_0 & ~i_10_373_412_0 & ~i_10_373_957_0 & ~i_10_373_2452_0 & ~i_10_373_2453_0 & ~i_10_373_2455_0 & ~i_10_373_2472_0 & ~i_10_373_2473_0 & ~i_10_373_2786_0 & ~i_10_373_2830_0) | (i_10_373_2922_0 & ~i_10_373_3840_0))) | (~i_10_373_966_0 & ~i_10_373_2472_0 & ~i_10_373_2659_0 & ~i_10_373_3283_0 & ~i_10_373_3284_0 & ~i_10_373_3469_0 & ~i_10_373_3470_0 & ~i_10_373_3787_0 & ~i_10_373_3847_0))) | (i_10_373_2704_0 & ((i_10_373_1652_0 & i_10_373_2703_0) | (~i_10_373_2451_0 & i_10_373_2923_0 & ~i_10_373_3283_0 & ~i_10_373_4292_0))) | (~i_10_373_1823_0 & i_10_373_2365_0) | (i_10_373_2833_0 & ~i_10_373_3613_0 & i_10_373_4287_0) | (i_10_373_3272_0 & i_10_373_3847_0 & ~i_10_373_4287_0));
endmodule



// Benchmark "kernel_10_374" written by ABC on Sun Jul 19 10:27:32 2020

module kernel_10_374 ( 
    i_10_374_117_0, i_10_374_171_0, i_10_374_173_0, i_10_374_222_0,
    i_10_374_249_0, i_10_374_250_0, i_10_374_282_0, i_10_374_283_0,
    i_10_374_295_0, i_10_374_316_0, i_10_374_423_0, i_10_374_425_0,
    i_10_374_431_0, i_10_374_433_0, i_10_374_449_0, i_10_374_467_0,
    i_10_374_748_0, i_10_374_795_0, i_10_374_799_0, i_10_374_892_0,
    i_10_374_893_0, i_10_374_957_0, i_10_374_958_0, i_10_374_959_0,
    i_10_374_960_0, i_10_374_1239_0, i_10_374_1309_0, i_10_374_1360_0,
    i_10_374_1578_0, i_10_374_1619_0, i_10_374_1648_0, i_10_374_1650_0,
    i_10_374_1652_0, i_10_374_1822_0, i_10_374_1913_0, i_10_374_1944_0,
    i_10_374_2178_0, i_10_374_2358_0, i_10_374_2361_0, i_10_374_2382_0,
    i_10_374_2409_0, i_10_374_2452_0, i_10_374_2454_0, i_10_374_2456_0,
    i_10_374_2632_0, i_10_374_2658_0, i_10_374_2661_0, i_10_374_2663_0,
    i_10_374_2702_0, i_10_374_2721_0, i_10_374_2725_0, i_10_374_2729_0,
    i_10_374_2731_0, i_10_374_2732_0, i_10_374_2734_0, i_10_374_2827_0,
    i_10_374_2884_0, i_10_374_3033_0, i_10_374_3036_0, i_10_374_3037_0,
    i_10_374_3042_0, i_10_374_3075_0, i_10_374_3085_0, i_10_374_3087_0,
    i_10_374_3150_0, i_10_374_3152_0, i_10_374_3154_0, i_10_374_3195_0,
    i_10_374_3196_0, i_10_374_3276_0, i_10_374_3279_0, i_10_374_3388_0,
    i_10_374_3583_0, i_10_374_3589_0, i_10_374_3612_0, i_10_374_3617_0,
    i_10_374_3645_0, i_10_374_3646_0, i_10_374_3647_0, i_10_374_3653_0,
    i_10_374_3783_0, i_10_374_3785_0, i_10_374_3835_0, i_10_374_3837_0,
    i_10_374_3838_0, i_10_374_3839_0, i_10_374_3848_0, i_10_374_3854_0,
    i_10_374_3855_0, i_10_374_3856_0, i_10_374_3857_0, i_10_374_3889_0,
    i_10_374_4024_0, i_10_374_4051_0, i_10_374_4120_0, i_10_374_4168_0,
    i_10_374_4212_0, i_10_374_4288_0, i_10_374_4291_0, i_10_374_4566_0,
    o_10_374_0_0  );
  input  i_10_374_117_0, i_10_374_171_0, i_10_374_173_0, i_10_374_222_0,
    i_10_374_249_0, i_10_374_250_0, i_10_374_282_0, i_10_374_283_0,
    i_10_374_295_0, i_10_374_316_0, i_10_374_423_0, i_10_374_425_0,
    i_10_374_431_0, i_10_374_433_0, i_10_374_449_0, i_10_374_467_0,
    i_10_374_748_0, i_10_374_795_0, i_10_374_799_0, i_10_374_892_0,
    i_10_374_893_0, i_10_374_957_0, i_10_374_958_0, i_10_374_959_0,
    i_10_374_960_0, i_10_374_1239_0, i_10_374_1309_0, i_10_374_1360_0,
    i_10_374_1578_0, i_10_374_1619_0, i_10_374_1648_0, i_10_374_1650_0,
    i_10_374_1652_0, i_10_374_1822_0, i_10_374_1913_0, i_10_374_1944_0,
    i_10_374_2178_0, i_10_374_2358_0, i_10_374_2361_0, i_10_374_2382_0,
    i_10_374_2409_0, i_10_374_2452_0, i_10_374_2454_0, i_10_374_2456_0,
    i_10_374_2632_0, i_10_374_2658_0, i_10_374_2661_0, i_10_374_2663_0,
    i_10_374_2702_0, i_10_374_2721_0, i_10_374_2725_0, i_10_374_2729_0,
    i_10_374_2731_0, i_10_374_2732_0, i_10_374_2734_0, i_10_374_2827_0,
    i_10_374_2884_0, i_10_374_3033_0, i_10_374_3036_0, i_10_374_3037_0,
    i_10_374_3042_0, i_10_374_3075_0, i_10_374_3085_0, i_10_374_3087_0,
    i_10_374_3150_0, i_10_374_3152_0, i_10_374_3154_0, i_10_374_3195_0,
    i_10_374_3196_0, i_10_374_3276_0, i_10_374_3279_0, i_10_374_3388_0,
    i_10_374_3583_0, i_10_374_3589_0, i_10_374_3612_0, i_10_374_3617_0,
    i_10_374_3645_0, i_10_374_3646_0, i_10_374_3647_0, i_10_374_3653_0,
    i_10_374_3783_0, i_10_374_3785_0, i_10_374_3835_0, i_10_374_3837_0,
    i_10_374_3838_0, i_10_374_3839_0, i_10_374_3848_0, i_10_374_3854_0,
    i_10_374_3855_0, i_10_374_3856_0, i_10_374_3857_0, i_10_374_3889_0,
    i_10_374_4024_0, i_10_374_4051_0, i_10_374_4120_0, i_10_374_4168_0,
    i_10_374_4212_0, i_10_374_4288_0, i_10_374_4291_0, i_10_374_4566_0;
  output o_10_374_0_0;
  assign o_10_374_0_0 = ~((~i_10_374_957_0 & ((~i_10_374_295_0 & ((~i_10_374_892_0 & ~i_10_374_893_0 & ~i_10_374_1239_0 & ~i_10_374_1360_0 & ~i_10_374_3036_0 & ~i_10_374_3037_0 & ~i_10_374_3783_0 & ~i_10_374_3848_0) | (~i_10_374_958_0 & ~i_10_374_1944_0 & ~i_10_374_2178_0 & ~i_10_374_2827_0 & ~i_10_374_3087_0 & ~i_10_374_4051_0))) | (~i_10_374_1360_0 & i_10_374_2663_0 & ~i_10_374_3075_0 & ~i_10_374_3087_0))) | (~i_10_374_249_0 & ((~i_10_374_1944_0 & ((~i_10_374_250_0 & ((~i_10_374_425_0 & ~i_10_374_958_0 & ~i_10_374_1360_0 & ~i_10_374_3042_0) | (~i_10_374_117_0 & ~i_10_374_959_0 & ~i_10_374_960_0 & ~i_10_374_3087_0 & ~i_10_374_3783_0 & ~i_10_374_4212_0))) | (~i_10_374_425_0 & ~i_10_374_893_0 & ~i_10_374_2661_0 & ~i_10_374_2884_0 & ~i_10_374_3033_0 & ~i_10_374_3839_0 & ~i_10_374_3848_0 & ~i_10_374_4120_0))) | (~i_10_374_250_0 & ((~i_10_374_283_0 & ~i_10_374_423_0 & ~i_10_374_960_0 & ~i_10_374_1913_0 & ~i_10_374_3087_0) | (~i_10_374_3583_0 & ~i_10_374_3855_0 & ~i_10_374_4212_0))) | (i_10_374_2725_0 & ~i_10_374_3612_0 & i_10_374_4120_0 & ~i_10_374_4566_0))) | (~i_10_374_960_0 & ((~i_10_374_431_0 & ((~i_10_374_958_0 & ~i_10_374_959_0 & ~i_10_374_2178_0 & ~i_10_374_2358_0 & ~i_10_374_3075_0) | (~i_10_374_433_0 & ~i_10_374_1239_0 & ~i_10_374_1360_0 & ~i_10_374_1648_0 & i_10_374_2827_0 & ~i_10_374_3036_0 & ~i_10_374_3087_0 & ~i_10_374_3837_0 & ~i_10_374_4051_0))) | (~i_10_374_449_0 & ((~i_10_374_117_0 & ~i_10_374_2661_0 & ~i_10_374_3589_0 & ~i_10_374_3653_0 & ~i_10_374_3854_0 & ~i_10_374_3855_0 & ~i_10_374_4024_0) | (~i_10_374_893_0 & ~i_10_374_959_0 & ~i_10_374_1822_0 & ~i_10_374_2452_0 & i_10_374_2731_0 & ~i_10_374_4291_0))) | (~i_10_374_2456_0 & ~i_10_374_2702_0 & i_10_374_3854_0 & ~i_10_374_3855_0 & i_10_374_4120_0 & ~i_10_374_4566_0))) | (~i_10_374_892_0 & ((~i_10_374_958_0 & ~i_10_374_2178_0 & i_10_374_3195_0) | (~i_10_374_117_0 & ~i_10_374_1360_0 & ~i_10_374_2456_0 & ~i_10_374_2729_0 & ~i_10_374_3589_0 & ~i_10_374_3848_0 & ~i_10_374_3855_0 & ~i_10_374_4566_0))) | (~i_10_374_117_0 & ((~i_10_374_449_0 & ~i_10_374_3195_0 & ~i_10_374_3583_0 & ~i_10_374_3612_0 & ~i_10_374_3854_0 & ~i_10_374_3855_0 & ~i_10_374_3856_0) | (~i_10_374_958_0 & ~i_10_374_1239_0 & ~i_10_374_2827_0 & i_10_374_3856_0 & ~i_10_374_4291_0))) | (i_10_374_3196_0 & ((i_10_374_467_0 & i_10_374_1650_0) | (~i_10_374_2827_0 & i_10_374_3195_0 & i_10_374_4291_0))) | (i_10_374_295_0 & i_10_374_3617_0) | (~i_10_374_3036_0 & i_10_374_3835_0 & ~i_10_374_3857_0) | (~i_10_374_3612_0 & ~i_10_374_3856_0 & ~i_10_374_4024_0 & ~i_10_374_4120_0));
endmodule



// Benchmark "kernel_10_375" written by ABC on Sun Jul 19 10:27:33 2020

module kernel_10_375 ( 
    i_10_375_189_0, i_10_375_220_0, i_10_375_283_0, i_10_375_284_0,
    i_10_375_318_0, i_10_375_361_0, i_10_375_364_0, i_10_375_390_0,
    i_10_375_433_0, i_10_375_444_0, i_10_375_467_0, i_10_375_505_0,
    i_10_375_639_0, i_10_375_739_0, i_10_375_750_0, i_10_375_945_0,
    i_10_375_946_0, i_10_375_948_0, i_10_375_949_0, i_10_375_1000_0,
    i_10_375_1002_0, i_10_375_1027_0, i_10_375_1028_0, i_10_375_1030_0,
    i_10_375_1056_0, i_10_375_1152_0, i_10_375_1153_0, i_10_375_1236_0,
    i_10_375_1237_0, i_10_375_1238_0, i_10_375_1244_0, i_10_375_1270_0,
    i_10_375_1311_0, i_10_375_1312_0, i_10_375_1315_0, i_10_375_1360_0,
    i_10_375_1362_0, i_10_375_1395_0, i_10_375_1440_0, i_10_375_1620_0,
    i_10_375_1650_0, i_10_375_1651_0, i_10_375_1713_0, i_10_375_1737_0,
    i_10_375_1740_0, i_10_375_1981_0, i_10_375_1990_0, i_10_375_2019_0,
    i_10_375_2028_0, i_10_375_2152_0, i_10_375_2153_0, i_10_375_2233_0,
    i_10_375_2359_0, i_10_375_2364_0, i_10_375_2430_0, i_10_375_2456_0,
    i_10_375_2473_0, i_10_375_2556_0, i_10_375_2567_0, i_10_375_2632_0,
    i_10_375_2754_0, i_10_375_2784_0, i_10_375_2817_0, i_10_375_2844_0,
    i_10_375_2863_0, i_10_375_2961_0, i_10_375_3070_0, i_10_375_3071_0,
    i_10_375_3087_0, i_10_375_3088_0, i_10_375_3127_0, i_10_375_3196_0,
    i_10_375_3312_0, i_10_375_3313_0, i_10_375_3472_0, i_10_375_3541_0,
    i_10_375_3583_0, i_10_375_3653_0, i_10_375_3682_0, i_10_375_3683_0,
    i_10_375_3700_0, i_10_375_3784_0, i_10_375_3838_0, i_10_375_3846_0,
    i_10_375_3889_0, i_10_375_3979_0, i_10_375_3991_0, i_10_375_4123_0,
    i_10_375_4126_0, i_10_375_4169_0, i_10_375_4214_0, i_10_375_4230_0,
    i_10_375_4258_0, i_10_375_4269_0, i_10_375_4292_0, i_10_375_4350_0,
    i_10_375_4370_0, i_10_375_4375_0, i_10_375_4437_0, i_10_375_4456_0,
    o_10_375_0_0  );
  input  i_10_375_189_0, i_10_375_220_0, i_10_375_283_0, i_10_375_284_0,
    i_10_375_318_0, i_10_375_361_0, i_10_375_364_0, i_10_375_390_0,
    i_10_375_433_0, i_10_375_444_0, i_10_375_467_0, i_10_375_505_0,
    i_10_375_639_0, i_10_375_739_0, i_10_375_750_0, i_10_375_945_0,
    i_10_375_946_0, i_10_375_948_0, i_10_375_949_0, i_10_375_1000_0,
    i_10_375_1002_0, i_10_375_1027_0, i_10_375_1028_0, i_10_375_1030_0,
    i_10_375_1056_0, i_10_375_1152_0, i_10_375_1153_0, i_10_375_1236_0,
    i_10_375_1237_0, i_10_375_1238_0, i_10_375_1244_0, i_10_375_1270_0,
    i_10_375_1311_0, i_10_375_1312_0, i_10_375_1315_0, i_10_375_1360_0,
    i_10_375_1362_0, i_10_375_1395_0, i_10_375_1440_0, i_10_375_1620_0,
    i_10_375_1650_0, i_10_375_1651_0, i_10_375_1713_0, i_10_375_1737_0,
    i_10_375_1740_0, i_10_375_1981_0, i_10_375_1990_0, i_10_375_2019_0,
    i_10_375_2028_0, i_10_375_2152_0, i_10_375_2153_0, i_10_375_2233_0,
    i_10_375_2359_0, i_10_375_2364_0, i_10_375_2430_0, i_10_375_2456_0,
    i_10_375_2473_0, i_10_375_2556_0, i_10_375_2567_0, i_10_375_2632_0,
    i_10_375_2754_0, i_10_375_2784_0, i_10_375_2817_0, i_10_375_2844_0,
    i_10_375_2863_0, i_10_375_2961_0, i_10_375_3070_0, i_10_375_3071_0,
    i_10_375_3087_0, i_10_375_3088_0, i_10_375_3127_0, i_10_375_3196_0,
    i_10_375_3312_0, i_10_375_3313_0, i_10_375_3472_0, i_10_375_3541_0,
    i_10_375_3583_0, i_10_375_3653_0, i_10_375_3682_0, i_10_375_3683_0,
    i_10_375_3700_0, i_10_375_3784_0, i_10_375_3838_0, i_10_375_3846_0,
    i_10_375_3889_0, i_10_375_3979_0, i_10_375_3991_0, i_10_375_4123_0,
    i_10_375_4126_0, i_10_375_4169_0, i_10_375_4214_0, i_10_375_4230_0,
    i_10_375_4258_0, i_10_375_4269_0, i_10_375_4292_0, i_10_375_4350_0,
    i_10_375_4370_0, i_10_375_4375_0, i_10_375_4437_0, i_10_375_4456_0;
  output o_10_375_0_0;
  assign o_10_375_0_0 = 0;
endmodule



// Benchmark "kernel_10_376" written by ABC on Sun Jul 19 10:27:35 2020

module kernel_10_376 ( 
    i_10_376_178_0, i_10_376_184_0, i_10_376_220_0, i_10_376_221_0,
    i_10_376_282_0, i_10_376_283_0, i_10_376_284_0, i_10_376_287_0,
    i_10_376_317_0, i_10_376_319_0, i_10_376_393_0, i_10_376_430_0,
    i_10_376_441_0, i_10_376_445_0, i_10_376_463_0, i_10_376_466_0,
    i_10_376_504_0, i_10_376_511_0, i_10_376_512_0, i_10_376_520_0,
    i_10_376_755_0, i_10_376_797_0, i_10_376_964_0, i_10_376_1033_0,
    i_10_376_1124_0, i_10_376_1136_0, i_10_376_1138_0, i_10_376_1236_0,
    i_10_376_1237_0, i_10_376_1249_0, i_10_376_1260_0, i_10_376_1365_0,
    i_10_376_1366_0, i_10_376_1555_0, i_10_376_1556_0, i_10_376_1575_0,
    i_10_376_1684_0, i_10_376_1689_0, i_10_376_1821_0, i_10_376_1824_0,
    i_10_376_1825_0, i_10_376_1826_0, i_10_376_1912_0, i_10_376_1914_0,
    i_10_376_1915_0, i_10_376_2017_0, i_10_376_2357_0, i_10_376_2451_0,
    i_10_376_2454_0, i_10_376_2455_0, i_10_376_2456_0, i_10_376_2466_0,
    i_10_376_2467_0, i_10_376_2635_0, i_10_376_2658_0, i_10_376_2659_0,
    i_10_376_2660_0, i_10_376_2680_0, i_10_376_2701_0, i_10_376_2721_0,
    i_10_376_2723_0, i_10_376_2731_0, i_10_376_2787_0, i_10_376_2818_0,
    i_10_376_2824_0, i_10_376_2826_0, i_10_376_2827_0, i_10_376_2830_0,
    i_10_376_2883_0, i_10_376_2884_0, i_10_376_2885_0, i_10_376_2982_0,
    i_10_376_3035_0, i_10_376_3039_0, i_10_376_3041_0, i_10_376_3069_0,
    i_10_376_3150_0, i_10_376_3151_0, i_10_376_3158_0, i_10_376_3267_0,
    i_10_376_3271_0, i_10_376_3328_0, i_10_376_3391_0, i_10_376_3409_0,
    i_10_376_3586_0, i_10_376_3587_0, i_10_376_3612_0, i_10_376_3613_0,
    i_10_376_3615_0, i_10_376_3783_0, i_10_376_3847_0, i_10_376_3850_0,
    i_10_376_3855_0, i_10_376_3856_0, i_10_376_3858_0, i_10_376_3982_0,
    i_10_376_4117_0, i_10_376_4118_0, i_10_376_4119_0, i_10_376_4270_0,
    o_10_376_0_0  );
  input  i_10_376_178_0, i_10_376_184_0, i_10_376_220_0, i_10_376_221_0,
    i_10_376_282_0, i_10_376_283_0, i_10_376_284_0, i_10_376_287_0,
    i_10_376_317_0, i_10_376_319_0, i_10_376_393_0, i_10_376_430_0,
    i_10_376_441_0, i_10_376_445_0, i_10_376_463_0, i_10_376_466_0,
    i_10_376_504_0, i_10_376_511_0, i_10_376_512_0, i_10_376_520_0,
    i_10_376_755_0, i_10_376_797_0, i_10_376_964_0, i_10_376_1033_0,
    i_10_376_1124_0, i_10_376_1136_0, i_10_376_1138_0, i_10_376_1236_0,
    i_10_376_1237_0, i_10_376_1249_0, i_10_376_1260_0, i_10_376_1365_0,
    i_10_376_1366_0, i_10_376_1555_0, i_10_376_1556_0, i_10_376_1575_0,
    i_10_376_1684_0, i_10_376_1689_0, i_10_376_1821_0, i_10_376_1824_0,
    i_10_376_1825_0, i_10_376_1826_0, i_10_376_1912_0, i_10_376_1914_0,
    i_10_376_1915_0, i_10_376_2017_0, i_10_376_2357_0, i_10_376_2451_0,
    i_10_376_2454_0, i_10_376_2455_0, i_10_376_2456_0, i_10_376_2466_0,
    i_10_376_2467_0, i_10_376_2635_0, i_10_376_2658_0, i_10_376_2659_0,
    i_10_376_2660_0, i_10_376_2680_0, i_10_376_2701_0, i_10_376_2721_0,
    i_10_376_2723_0, i_10_376_2731_0, i_10_376_2787_0, i_10_376_2818_0,
    i_10_376_2824_0, i_10_376_2826_0, i_10_376_2827_0, i_10_376_2830_0,
    i_10_376_2883_0, i_10_376_2884_0, i_10_376_2885_0, i_10_376_2982_0,
    i_10_376_3035_0, i_10_376_3039_0, i_10_376_3041_0, i_10_376_3069_0,
    i_10_376_3150_0, i_10_376_3151_0, i_10_376_3158_0, i_10_376_3267_0,
    i_10_376_3271_0, i_10_376_3328_0, i_10_376_3391_0, i_10_376_3409_0,
    i_10_376_3586_0, i_10_376_3587_0, i_10_376_3612_0, i_10_376_3613_0,
    i_10_376_3615_0, i_10_376_3783_0, i_10_376_3847_0, i_10_376_3850_0,
    i_10_376_3855_0, i_10_376_3856_0, i_10_376_3858_0, i_10_376_3982_0,
    i_10_376_4117_0, i_10_376_4118_0, i_10_376_4119_0, i_10_376_4270_0;
  output o_10_376_0_0;
  assign o_10_376_0_0 = ~((~i_10_376_178_0 & ((i_10_376_466_0 & ~i_10_376_2451_0 & i_10_376_2701_0 & ~i_10_376_3069_0 & ~i_10_376_3586_0) | (i_10_376_520_0 & ~i_10_376_2884_0 & ~i_10_376_2982_0 & i_10_376_3041_0 & i_10_376_3613_0 & ~i_10_376_3615_0 & ~i_10_376_3855_0))) | (~i_10_376_2787_0 & ((~i_10_376_184_0 & ((~i_10_376_220_0 & ~i_10_376_1236_0 & ~i_10_376_2723_0 & ~i_10_376_2826_0 & ~i_10_376_3035_0 & ~i_10_376_3267_0 & ~i_10_376_3586_0 & i_10_376_3856_0) | (~i_10_376_221_0 & i_10_376_283_0 & i_10_376_1915_0 & i_10_376_2455_0 & ~i_10_376_4119_0))) | (~i_10_376_1366_0 & ~i_10_376_3612_0 & ((~i_10_376_220_0 & ~i_10_376_221_0 & ~i_10_376_2467_0 & ~i_10_376_2660_0 & ~i_10_376_3035_0 & ~i_10_376_3855_0) | (~i_10_376_1915_0 & i_10_376_2731_0 & ~i_10_376_3613_0 & ~i_10_376_3847_0 & ~i_10_376_4270_0))) | (~i_10_376_1684_0 & ((~i_10_376_1821_0 & i_10_376_2827_0 & i_10_376_3391_0) | (~i_10_376_1236_0 & ~i_10_376_2721_0 & ~i_10_376_2827_0 & ~i_10_376_3035_0 & ~i_10_376_3069_0 & i_10_376_3612_0))) | (~i_10_376_1365_0 & i_10_376_2455_0 & i_10_376_2456_0 & ~i_10_376_2818_0) | (~i_10_376_284_0 & i_10_376_1689_0 & ~i_10_376_1825_0 & ~i_10_376_1826_0 & ~i_10_376_1912_0 & ~i_10_376_3850_0))) | (~i_10_376_221_0 & ~i_10_376_2818_0 & ((i_10_376_284_0 & ~i_10_376_520_0 & ~i_10_376_1365_0 & ~i_10_376_1912_0 & i_10_376_2635_0 & ~i_10_376_3271_0) | (~i_10_376_2658_0 & ~i_10_376_3391_0 & i_10_376_4118_0))) | (~i_10_376_1684_0 & ((~i_10_376_393_0 & ~i_10_376_2826_0 & ((~i_10_376_1237_0 & ~i_10_376_2721_0 & ~i_10_376_3587_0 & ~i_10_376_3612_0 & i_10_376_3856_0) | (~i_10_376_1555_0 & ~i_10_376_1912_0 & ~i_10_376_2466_0 & ~i_10_376_2660_0 & ~i_10_376_3856_0 & ~i_10_376_3982_0 & ~i_10_376_4118_0))) | (~i_10_376_184_0 & ~i_10_376_445_0 & ~i_10_376_1365_0 & ~i_10_376_1555_0 & ~i_10_376_1912_0 & ~i_10_376_3035_0 & ~i_10_376_3069_0 & ~i_10_376_3267_0 & ~i_10_376_3850_0 & ~i_10_376_3856_0 & ~i_10_376_3982_0))) | (~i_10_376_184_0 & ((~i_10_376_441_0 & i_10_376_1249_0 & ~i_10_376_1912_0 & ~i_10_376_2660_0) | (~i_10_376_463_0 & ~i_10_376_1249_0 & ~i_10_376_1365_0 & ~i_10_376_1366_0 & i_10_376_2701_0))) | (~i_10_376_441_0 & i_10_376_1826_0 & ((~i_10_376_282_0 & ~i_10_376_283_0 & ~i_10_376_1365_0 & ~i_10_376_1575_0) | (i_10_376_1825_0 & i_10_376_2456_0 & ~i_10_376_2466_0))) | (~i_10_376_1236_0 & ((~i_10_376_463_0 & ~i_10_376_1821_0 & ~i_10_376_1912_0 & ~i_10_376_3267_0) | (i_10_376_2659_0 & i_10_376_2731_0 & ~i_10_376_3615_0 & ~i_10_376_3855_0 & ~i_10_376_3982_0))) | (~i_10_376_463_0 & ((i_10_376_284_0 & ~i_10_376_2659_0) | (~i_10_376_1912_0 & ~i_10_376_2660_0 & i_10_376_2731_0 & ~i_10_376_3586_0 & ~i_10_376_3783_0))) | (~i_10_376_1249_0 & ((~i_10_376_1366_0 & i_10_376_1824_0 & ~i_10_376_2658_0) | (i_10_376_3409_0 & ~i_10_376_3586_0 & ~i_10_376_3783_0))) | (i_10_376_1825_0 & ((i_10_376_220_0 & i_10_376_1684_0) | (~i_10_376_3039_0 & i_10_376_3409_0))) | (~i_10_376_1365_0 & ((~i_10_376_1237_0 & ((~i_10_376_284_0 & ~i_10_376_2723_0 & ~i_10_376_3783_0 & ~i_10_376_3856_0) | (i_10_376_1033_0 & ~i_10_376_4117_0))) | (~i_10_376_1912_0 & ~i_10_376_3613_0 & ((~i_10_376_2466_0 & ~i_10_376_2659_0 & ~i_10_376_3855_0) | (~i_10_376_1366_0 & ~i_10_376_1821_0 & ~i_10_376_3267_0 & ~i_10_376_3612_0 & i_10_376_4117_0))))) | (~i_10_376_1237_0 & ((i_10_376_2017_0 & ~i_10_376_2467_0) | (~i_10_376_2658_0 & ~i_10_376_2659_0 & ~i_10_376_3587_0 & ~i_10_376_3855_0))) | (~i_10_376_1366_0 & ~i_10_376_2830_0 & ((i_10_376_178_0 & i_10_376_1821_0 & ~i_10_376_2466_0 & ~i_10_376_3039_0) | (i_10_376_2824_0 & ~i_10_376_3855_0))) | (i_10_376_2884_0 & ~i_10_376_3612_0 & ~i_10_376_3858_0));
endmodule



// Benchmark "kernel_10_377" written by ABC on Sun Jul 19 10:27:36 2020

module kernel_10_377 ( 
    i_10_377_180_0, i_10_377_222_0, i_10_377_276_0, i_10_377_283_0,
    i_10_377_284_0, i_10_377_324_0, i_10_377_325_0, i_10_377_388_0,
    i_10_377_426_0, i_10_377_435_0, i_10_377_436_0, i_10_377_442_0,
    i_10_377_443_0, i_10_377_459_0, i_10_377_465_0, i_10_377_466_0,
    i_10_377_514_0, i_10_377_958_0, i_10_377_959_0, i_10_377_960_0,
    i_10_377_961_0, i_10_377_962_0, i_10_377_1163_0, i_10_377_1164_0,
    i_10_377_1233_0, i_10_377_1236_0, i_10_377_1245_0, i_10_377_1248_0,
    i_10_377_1432_0, i_10_377_1546_0, i_10_377_1582_0, i_10_377_1652_0,
    i_10_377_1690_0, i_10_377_1720_0, i_10_377_1759_0, i_10_377_1760_0,
    i_10_377_1820_0, i_10_377_1822_0, i_10_377_1823_0, i_10_377_1824_0,
    i_10_377_1826_0, i_10_377_2029_0, i_10_377_2352_0, i_10_377_2380_0,
    i_10_377_2452_0, i_10_377_2453_0, i_10_377_2630_0, i_10_377_2658_0,
    i_10_377_2659_0, i_10_377_2660_0, i_10_377_2702_0, i_10_377_2708_0,
    i_10_377_2713_0, i_10_377_2721_0, i_10_377_2722_0, i_10_377_2724_0,
    i_10_377_2727_0, i_10_377_2728_0, i_10_377_2730_0, i_10_377_2731_0,
    i_10_377_2735_0, i_10_377_2982_0, i_10_377_3033_0, i_10_377_3034_0,
    i_10_377_3035_0, i_10_377_3036_0, i_10_377_3037_0, i_10_377_3069_0,
    i_10_377_3150_0, i_10_377_3231_0, i_10_377_3268_0, i_10_377_3271_0,
    i_10_377_3316_0, i_10_377_3332_0, i_10_377_3388_0, i_10_377_3389_0,
    i_10_377_3391_0, i_10_377_3469_0, i_10_377_3494_0, i_10_377_3537_0,
    i_10_377_3616_0, i_10_377_3649_0, i_10_377_3783_0, i_10_377_3837_0,
    i_10_377_3847_0, i_10_377_3848_0, i_10_377_3849_0, i_10_377_3850_0,
    i_10_377_3857_0, i_10_377_3983_0, i_10_377_4113_0, i_10_377_4120_0,
    i_10_377_4121_0, i_10_377_4185_0, i_10_377_4269_0, i_10_377_4279_0,
    i_10_377_4285_0, i_10_377_4286_0, i_10_377_4289_0, i_10_377_4563_0,
    o_10_377_0_0  );
  input  i_10_377_180_0, i_10_377_222_0, i_10_377_276_0, i_10_377_283_0,
    i_10_377_284_0, i_10_377_324_0, i_10_377_325_0, i_10_377_388_0,
    i_10_377_426_0, i_10_377_435_0, i_10_377_436_0, i_10_377_442_0,
    i_10_377_443_0, i_10_377_459_0, i_10_377_465_0, i_10_377_466_0,
    i_10_377_514_0, i_10_377_958_0, i_10_377_959_0, i_10_377_960_0,
    i_10_377_961_0, i_10_377_962_0, i_10_377_1163_0, i_10_377_1164_0,
    i_10_377_1233_0, i_10_377_1236_0, i_10_377_1245_0, i_10_377_1248_0,
    i_10_377_1432_0, i_10_377_1546_0, i_10_377_1582_0, i_10_377_1652_0,
    i_10_377_1690_0, i_10_377_1720_0, i_10_377_1759_0, i_10_377_1760_0,
    i_10_377_1820_0, i_10_377_1822_0, i_10_377_1823_0, i_10_377_1824_0,
    i_10_377_1826_0, i_10_377_2029_0, i_10_377_2352_0, i_10_377_2380_0,
    i_10_377_2452_0, i_10_377_2453_0, i_10_377_2630_0, i_10_377_2658_0,
    i_10_377_2659_0, i_10_377_2660_0, i_10_377_2702_0, i_10_377_2708_0,
    i_10_377_2713_0, i_10_377_2721_0, i_10_377_2722_0, i_10_377_2724_0,
    i_10_377_2727_0, i_10_377_2728_0, i_10_377_2730_0, i_10_377_2731_0,
    i_10_377_2735_0, i_10_377_2982_0, i_10_377_3033_0, i_10_377_3034_0,
    i_10_377_3035_0, i_10_377_3036_0, i_10_377_3037_0, i_10_377_3069_0,
    i_10_377_3150_0, i_10_377_3231_0, i_10_377_3268_0, i_10_377_3271_0,
    i_10_377_3316_0, i_10_377_3332_0, i_10_377_3388_0, i_10_377_3389_0,
    i_10_377_3391_0, i_10_377_3469_0, i_10_377_3494_0, i_10_377_3537_0,
    i_10_377_3616_0, i_10_377_3649_0, i_10_377_3783_0, i_10_377_3837_0,
    i_10_377_3847_0, i_10_377_3848_0, i_10_377_3849_0, i_10_377_3850_0,
    i_10_377_3857_0, i_10_377_3983_0, i_10_377_4113_0, i_10_377_4120_0,
    i_10_377_4121_0, i_10_377_4185_0, i_10_377_4269_0, i_10_377_4279_0,
    i_10_377_4285_0, i_10_377_4286_0, i_10_377_4289_0, i_10_377_4563_0;
  output o_10_377_0_0;
  assign o_10_377_0_0 = ~((~i_10_377_180_0 & ((~i_10_377_283_0 & ((i_10_377_443_0 & ~i_10_377_958_0 & ~i_10_377_3391_0 & ~i_10_377_3537_0 & ~i_10_377_3847_0 & ~i_10_377_3850_0) | (~i_10_377_961_0 & ~i_10_377_1233_0 & ~i_10_377_2029_0 & ~i_10_377_2352_0 & ~i_10_377_2660_0 & ~i_10_377_2735_0 & ~i_10_377_3848_0 & ~i_10_377_3849_0 & ~i_10_377_4120_0 & ~i_10_377_4563_0))) | (~i_10_377_959_0 & ~i_10_377_3033_0 & ((~i_10_377_962_0 & i_10_377_2630_0 & ~i_10_377_2724_0 & ~i_10_377_3649_0) | (~i_10_377_960_0 & ~i_10_377_2352_0 & ~i_10_377_2630_0 & ~i_10_377_3036_0 & ~i_10_377_3231_0 & ~i_10_377_3391_0 & ~i_10_377_3848_0 & ~i_10_377_4285_0 & ~i_10_377_4563_0))) | (~i_10_377_961_0 & ((i_10_377_1823_0 & ~i_10_377_2352_0 & ~i_10_377_2702_0 & i_10_377_2728_0 & ~i_10_377_2730_0 & ~i_10_377_3034_0 & ~i_10_377_3849_0) | (~i_10_377_958_0 & ~i_10_377_1546_0 & ~i_10_377_2728_0 & ~i_10_377_2735_0 & i_10_377_3033_0 & ~i_10_377_3847_0 & ~i_10_377_4269_0))) | (~i_10_377_958_0 & ~i_10_377_2730_0 & ~i_10_377_4279_0 & ((~i_10_377_962_0 & ~i_10_377_2380_0 & ~i_10_377_2731_0 & ~i_10_377_3035_0 & ~i_10_377_3036_0 & ~i_10_377_3069_0 & ~i_10_377_3537_0) | (~i_10_377_443_0 & i_10_377_465_0 & ~i_10_377_1546_0 & ~i_10_377_2708_0 & ~i_10_377_3389_0 & ~i_10_377_3847_0))) | (~i_10_377_1432_0 & ((~i_10_377_1248_0 & ~i_10_377_2029_0 & i_10_377_2380_0 & ~i_10_377_3037_0) | (~i_10_377_466_0 & ~i_10_377_962_0 & ~i_10_377_1164_0 & ~i_10_377_1823_0 & ~i_10_377_3035_0 & ~i_10_377_3036_0 & ~i_10_377_3316_0 & ~i_10_377_3783_0 & ~i_10_377_3848_0))))) | (~i_10_377_284_0 & ((~i_10_377_961_0 & ~i_10_377_1432_0 & ~i_10_377_1822_0 & ~i_10_377_2722_0 & ~i_10_377_2735_0 & ~i_10_377_3036_0 & ~i_10_377_3037_0 & ~i_10_377_3316_0) | (i_10_377_283_0 & ~i_10_377_459_0 & ~i_10_377_958_0 & ~i_10_377_2452_0 & ~i_10_377_2730_0 & ~i_10_377_3469_0 & ~i_10_377_3850_0))) | (~i_10_377_459_0 & ((i_10_377_514_0 & i_10_377_1820_0 & i_10_377_2630_0) | (~i_10_377_1236_0 & ~i_10_377_1582_0 & i_10_377_1823_0 & ~i_10_377_3848_0 & ~i_10_377_3857_0 & ~i_10_377_3983_0))) | (~i_10_377_3849_0 & ((~i_10_377_3847_0 & ((~i_10_377_960_0 & ((~i_10_377_465_0 & ~i_10_377_959_0 & ~i_10_377_1164_0 & ~i_10_377_2708_0 & ~i_10_377_3033_0 & ~i_10_377_3388_0 & ~i_10_377_3391_0) | (~i_10_377_1233_0 & ~i_10_377_1248_0 & ~i_10_377_1582_0 & i_10_377_3857_0 & ~i_10_377_4121_0))) | (~i_10_377_388_0 & i_10_377_514_0 & i_10_377_2728_0))) | (i_10_377_2722_0 & ~i_10_377_3850_0 & ((~i_10_377_961_0 & ~i_10_377_3035_0 & ~i_10_377_3037_0 & ~i_10_377_3469_0) | (~i_10_377_1164_0 & i_10_377_4113_0))) | (~i_10_377_958_0 & i_10_377_1432_0 & ~i_10_377_1690_0 & ~i_10_377_2380_0 & ~i_10_377_2452_0 & ~i_10_377_3069_0 & ~i_10_377_3271_0 & ~i_10_377_3316_0 & ~i_10_377_3469_0) | (~i_10_377_962_0 & ~i_10_377_1163_0 & ~i_10_377_1546_0 & i_10_377_1820_0 & ~i_10_377_2727_0 & ~i_10_377_3537_0 & ~i_10_377_3783_0 & ~i_10_377_4120_0))) | (~i_10_377_958_0 & ((~i_10_377_1164_0 & ~i_10_377_1245_0 & ~i_10_377_1432_0 & ~i_10_377_2735_0 & ~i_10_377_3391_0 & ~i_10_377_3848_0 & ~i_10_377_4120_0) | (~i_10_377_388_0 & ~i_10_377_2029_0 & ~i_10_377_2730_0 & ~i_10_377_3033_0 & ~i_10_377_3037_0 & ~i_10_377_3316_0 & ~i_10_377_3537_0 & ~i_10_377_4121_0))) | (~i_10_377_2727_0 & ((~i_10_377_959_0 & ~i_10_377_2352_0 & ((~i_10_377_1822_0 & ~i_10_377_3037_0 & ~i_10_377_3271_0 & ~i_10_377_4269_0) | (~i_10_377_436_0 & ~i_10_377_1163_0 & ~i_10_377_1582_0 & ~i_10_377_2452_0 & ~i_10_377_2728_0 & ~i_10_377_2730_0 & ~i_10_377_3469_0 & ~i_10_377_4289_0))) | (~i_10_377_388_0 & ~i_10_377_1163_0 & ~i_10_377_2029_0 & ~i_10_377_3036_0 & ~i_10_377_3316_0 & ~i_10_377_3537_0 & ~i_10_377_4121_0 & ~i_10_377_4285_0 & i_10_377_4289_0))) | (~i_10_377_388_0 & ((i_10_377_435_0 & i_10_377_1652_0 & ~i_10_377_2730_0) | (~i_10_377_962_0 & ~i_10_377_1248_0 & ~i_10_377_1546_0 & ~i_10_377_3037_0 & ~i_10_377_3316_0 & ~i_10_377_3391_0 & ~i_10_377_3850_0 & ~i_10_377_3983_0 & ~i_10_377_4269_0))) | (~i_10_377_3033_0 & ~i_10_377_4120_0 & ((i_10_377_465_0 & ~i_10_377_1233_0 & ~i_10_377_1245_0 & ~i_10_377_2659_0 & i_10_377_2731_0) | (~i_10_377_1164_0 & ~i_10_377_1690_0 & ~i_10_377_2728_0 & i_10_377_3037_0 & ~i_10_377_3316_0 & ~i_10_377_3391_0 & ~i_10_377_3850_0 & ~i_10_377_3983_0 & ~i_10_377_4121_0 & ~i_10_377_4269_0))) | (~i_10_377_3783_0 & ((~i_10_377_959_0 & ~i_10_377_1546_0 & ~i_10_377_1822_0 & ~i_10_377_3037_0 & i_10_377_3616_0 & ~i_10_377_3850_0) | (~i_10_377_3316_0 & ~i_10_377_3391_0 & ~i_10_377_2731_0 & ~i_10_377_3069_0 & ~i_10_377_4285_0 & ~i_10_377_4563_0 & ~i_10_377_3469_0 & ~i_10_377_3649_0))) | (i_10_377_2713_0 & ~i_10_377_3388_0 & ~i_10_377_3389_0 & i_10_377_3391_0 & ~i_10_377_4269_0));
endmodule



// Benchmark "kernel_10_378" written by ABC on Sun Jul 19 10:27:37 2020

module kernel_10_378 ( 
    i_10_378_145_0, i_10_378_171_0, i_10_378_173_0, i_10_378_223_0,
    i_10_378_247_0, i_10_378_261_0, i_10_378_262_0, i_10_378_263_0,
    i_10_378_270_0, i_10_378_273_0, i_10_378_282_0, i_10_378_315_0,
    i_10_378_316_0, i_10_378_317_0, i_10_378_319_0, i_10_378_320_0,
    i_10_378_388_0, i_10_378_389_0, i_10_378_391_0, i_10_378_392_0,
    i_10_378_406_0, i_10_378_407_0, i_10_378_428_0, i_10_378_433_0,
    i_10_378_434_0, i_10_378_437_0, i_10_378_442_0, i_10_378_445_0,
    i_10_378_623_0, i_10_378_792_0, i_10_378_892_0, i_10_378_994_0,
    i_10_378_1000_0, i_10_378_1001_0, i_10_378_1081_0, i_10_378_1082_0,
    i_10_378_1100_0, i_10_378_1103_0, i_10_378_1138_0, i_10_378_1217_0,
    i_10_378_1219_0, i_10_378_1233_0, i_10_378_1296_0, i_10_378_1299_0,
    i_10_378_1307_0, i_10_378_1343_0, i_10_378_1433_0, i_10_378_1544_0,
    i_10_378_1553_0, i_10_378_1580_0, i_10_378_1650_0, i_10_378_1652_0,
    i_10_378_1655_0, i_10_378_1765_0, i_10_378_1823_0, i_10_378_1825_0,
    i_10_378_1826_0, i_10_378_1910_0, i_10_378_2000_0, i_10_378_2198_0,
    i_10_378_2200_0, i_10_378_2362_0, i_10_378_2448_0, i_10_378_2518_0,
    i_10_378_2602_0, i_10_378_2657_0, i_10_378_2660_0, i_10_378_2721_0,
    i_10_378_2781_0, i_10_378_2830_0, i_10_378_2832_0, i_10_378_2918_0,
    i_10_378_3038_0, i_10_378_3072_0, i_10_378_3151_0, i_10_378_3196_0,
    i_10_378_3197_0, i_10_378_3200_0, i_10_378_3202_0, i_10_378_3203_0,
    i_10_378_3323_0, i_10_378_3405_0, i_10_378_3431_0, i_10_378_3470_0,
    i_10_378_3538_0, i_10_378_3539_0, i_10_378_3610_0, i_10_378_3647_0,
    i_10_378_3793_0, i_10_378_3834_0, i_10_378_3836_0, i_10_378_3838_0,
    i_10_378_3844_0, i_10_378_3880_0, i_10_378_3979_0, i_10_378_3980_0,
    i_10_378_4117_0, i_10_378_4169_0, i_10_378_4277_0, i_10_378_4283_0,
    o_10_378_0_0  );
  input  i_10_378_145_0, i_10_378_171_0, i_10_378_173_0, i_10_378_223_0,
    i_10_378_247_0, i_10_378_261_0, i_10_378_262_0, i_10_378_263_0,
    i_10_378_270_0, i_10_378_273_0, i_10_378_282_0, i_10_378_315_0,
    i_10_378_316_0, i_10_378_317_0, i_10_378_319_0, i_10_378_320_0,
    i_10_378_388_0, i_10_378_389_0, i_10_378_391_0, i_10_378_392_0,
    i_10_378_406_0, i_10_378_407_0, i_10_378_428_0, i_10_378_433_0,
    i_10_378_434_0, i_10_378_437_0, i_10_378_442_0, i_10_378_445_0,
    i_10_378_623_0, i_10_378_792_0, i_10_378_892_0, i_10_378_994_0,
    i_10_378_1000_0, i_10_378_1001_0, i_10_378_1081_0, i_10_378_1082_0,
    i_10_378_1100_0, i_10_378_1103_0, i_10_378_1138_0, i_10_378_1217_0,
    i_10_378_1219_0, i_10_378_1233_0, i_10_378_1296_0, i_10_378_1299_0,
    i_10_378_1307_0, i_10_378_1343_0, i_10_378_1433_0, i_10_378_1544_0,
    i_10_378_1553_0, i_10_378_1580_0, i_10_378_1650_0, i_10_378_1652_0,
    i_10_378_1655_0, i_10_378_1765_0, i_10_378_1823_0, i_10_378_1825_0,
    i_10_378_1826_0, i_10_378_1910_0, i_10_378_2000_0, i_10_378_2198_0,
    i_10_378_2200_0, i_10_378_2362_0, i_10_378_2448_0, i_10_378_2518_0,
    i_10_378_2602_0, i_10_378_2657_0, i_10_378_2660_0, i_10_378_2721_0,
    i_10_378_2781_0, i_10_378_2830_0, i_10_378_2832_0, i_10_378_2918_0,
    i_10_378_3038_0, i_10_378_3072_0, i_10_378_3151_0, i_10_378_3196_0,
    i_10_378_3197_0, i_10_378_3200_0, i_10_378_3202_0, i_10_378_3203_0,
    i_10_378_3323_0, i_10_378_3405_0, i_10_378_3431_0, i_10_378_3470_0,
    i_10_378_3538_0, i_10_378_3539_0, i_10_378_3610_0, i_10_378_3647_0,
    i_10_378_3793_0, i_10_378_3834_0, i_10_378_3836_0, i_10_378_3838_0,
    i_10_378_3844_0, i_10_378_3880_0, i_10_378_3979_0, i_10_378_3980_0,
    i_10_378_4117_0, i_10_378_4169_0, i_10_378_4277_0, i_10_378_4283_0;
  output o_10_378_0_0;
  assign o_10_378_0_0 = ~((~i_10_378_263_0 & ((~i_10_378_389_0 & ~i_10_378_434_0 & ~i_10_378_437_0) | (~i_10_378_433_0 & ~i_10_378_1001_0 & ~i_10_378_1233_0 & ~i_10_378_1544_0 & ~i_10_378_3202_0 & ~i_10_378_3431_0))) | (~i_10_378_388_0 & ((~i_10_378_261_0 & ~i_10_378_1081_0 & ~i_10_378_1343_0 & ~i_10_378_3470_0 & ~i_10_378_3538_0 & ~i_10_378_3539_0) | (~i_10_378_392_0 & ~i_10_378_1001_0 & ~i_10_378_3196_0 & ~i_10_378_4277_0))) | (~i_10_378_389_0 & ~i_10_378_1826_0 & ((~i_10_378_320_0 & ~i_10_378_994_0 & ~i_10_378_1000_0 & ~i_10_378_1001_0 & ~i_10_378_4117_0) | (~i_10_378_262_0 & ~i_10_378_391_0 & ~i_10_378_3538_0 & ~i_10_378_4277_0))) | (~i_10_378_392_0 & ((~i_10_378_391_0 & ~i_10_378_437_0 & ~i_10_378_994_0 & ~i_10_378_3038_0 & ~i_10_378_3539_0) | (~i_10_378_145_0 & ~i_10_378_1082_0 & ~i_10_378_2000_0 & ~i_10_378_2448_0 & ~i_10_378_3197_0 & ~i_10_378_3200_0 & ~i_10_378_3844_0 & ~i_10_378_4283_0))) | (~i_10_378_1001_0 & ((i_10_378_173_0 & ~i_10_378_1307_0 & ~i_10_378_3538_0) | (~i_10_378_433_0 & ~i_10_378_3200_0 & ~i_10_378_3610_0 & ~i_10_378_3980_0 & ~i_10_378_4277_0))) | (i_10_378_171_0 & i_10_378_1655_0 & ~i_10_378_2000_0 & ~i_10_378_3038_0));
endmodule



// Benchmark "kernel_10_379" written by ABC on Sun Jul 19 10:27:38 2020

module kernel_10_379 ( 
    i_10_379_31_0, i_10_379_247_0, i_10_379_346_0, i_10_379_391_0,
    i_10_379_394_0, i_10_379_435_0, i_10_379_438_0, i_10_379_443_0,
    i_10_379_518_0, i_10_379_560_0, i_10_379_563_0, i_10_379_597_0,
    i_10_379_623_0, i_10_379_714_0, i_10_379_798_0, i_10_379_968_0,
    i_10_379_1010_0, i_10_379_1051_0, i_10_379_1236_0, i_10_379_1238_0,
    i_10_379_1240_0, i_10_379_1241_0, i_10_379_1269_0, i_10_379_1310_0,
    i_10_379_1359_0, i_10_379_1362_0, i_10_379_1364_0, i_10_379_1498_0,
    i_10_379_1543_0, i_10_379_1550_0, i_10_379_1632_0, i_10_379_1652_0,
    i_10_379_1684_0, i_10_379_1807_0, i_10_379_1822_0, i_10_379_1874_0,
    i_10_379_2021_0, i_10_379_2329_0, i_10_379_2354_0, i_10_379_2454_0,
    i_10_379_2468_0, i_10_379_2507_0, i_10_379_2513_0, i_10_379_2531_0,
    i_10_379_2566_0, i_10_379_2569_0, i_10_379_2612_0, i_10_379_2621_0,
    i_10_379_2635_0, i_10_379_2659_0, i_10_379_2660_0, i_10_379_2674_0,
    i_10_379_2707_0, i_10_379_2718_0, i_10_379_2719_0, i_10_379_2720_0,
    i_10_379_2722_0, i_10_379_2729_0, i_10_379_2821_0, i_10_379_2827_0,
    i_10_379_2830_0, i_10_379_2918_0, i_10_379_2919_0, i_10_379_2920_0,
    i_10_379_2921_0, i_10_379_3034_0, i_10_379_3072_0, i_10_379_3233_0,
    i_10_379_3285_0, i_10_379_3286_0, i_10_379_3355_0, i_10_379_3402_0,
    i_10_379_3434_0, i_10_379_3436_0, i_10_379_3437_0, i_10_379_3493_0,
    i_10_379_3505_0, i_10_379_3544_0, i_10_379_3613_0, i_10_379_3625_0,
    i_10_379_3653_0, i_10_379_3683_0, i_10_379_3688_0, i_10_379_3728_0,
    i_10_379_3827_0, i_10_379_3837_0, i_10_379_3846_0, i_10_379_3857_0,
    i_10_379_3890_0, i_10_379_4025_0, i_10_379_4122_0, i_10_379_4123_0,
    i_10_379_4124_0, i_10_379_4279_0, i_10_379_4288_0, i_10_379_4289_0,
    i_10_379_4307_0, i_10_379_4564_0, i_10_379_4582_0, i_10_379_4590_0,
    o_10_379_0_0  );
  input  i_10_379_31_0, i_10_379_247_0, i_10_379_346_0, i_10_379_391_0,
    i_10_379_394_0, i_10_379_435_0, i_10_379_438_0, i_10_379_443_0,
    i_10_379_518_0, i_10_379_560_0, i_10_379_563_0, i_10_379_597_0,
    i_10_379_623_0, i_10_379_714_0, i_10_379_798_0, i_10_379_968_0,
    i_10_379_1010_0, i_10_379_1051_0, i_10_379_1236_0, i_10_379_1238_0,
    i_10_379_1240_0, i_10_379_1241_0, i_10_379_1269_0, i_10_379_1310_0,
    i_10_379_1359_0, i_10_379_1362_0, i_10_379_1364_0, i_10_379_1498_0,
    i_10_379_1543_0, i_10_379_1550_0, i_10_379_1632_0, i_10_379_1652_0,
    i_10_379_1684_0, i_10_379_1807_0, i_10_379_1822_0, i_10_379_1874_0,
    i_10_379_2021_0, i_10_379_2329_0, i_10_379_2354_0, i_10_379_2454_0,
    i_10_379_2468_0, i_10_379_2507_0, i_10_379_2513_0, i_10_379_2531_0,
    i_10_379_2566_0, i_10_379_2569_0, i_10_379_2612_0, i_10_379_2621_0,
    i_10_379_2635_0, i_10_379_2659_0, i_10_379_2660_0, i_10_379_2674_0,
    i_10_379_2707_0, i_10_379_2718_0, i_10_379_2719_0, i_10_379_2720_0,
    i_10_379_2722_0, i_10_379_2729_0, i_10_379_2821_0, i_10_379_2827_0,
    i_10_379_2830_0, i_10_379_2918_0, i_10_379_2919_0, i_10_379_2920_0,
    i_10_379_2921_0, i_10_379_3034_0, i_10_379_3072_0, i_10_379_3233_0,
    i_10_379_3285_0, i_10_379_3286_0, i_10_379_3355_0, i_10_379_3402_0,
    i_10_379_3434_0, i_10_379_3436_0, i_10_379_3437_0, i_10_379_3493_0,
    i_10_379_3505_0, i_10_379_3544_0, i_10_379_3613_0, i_10_379_3625_0,
    i_10_379_3653_0, i_10_379_3683_0, i_10_379_3688_0, i_10_379_3728_0,
    i_10_379_3827_0, i_10_379_3837_0, i_10_379_3846_0, i_10_379_3857_0,
    i_10_379_3890_0, i_10_379_4025_0, i_10_379_4122_0, i_10_379_4123_0,
    i_10_379_4124_0, i_10_379_4279_0, i_10_379_4288_0, i_10_379_4289_0,
    i_10_379_4307_0, i_10_379_4564_0, i_10_379_4582_0, i_10_379_4590_0;
  output o_10_379_0_0;
  assign o_10_379_0_0 = 0;
endmodule



// Benchmark "kernel_10_380" written by ABC on Sun Jul 19 10:27:39 2020

module kernel_10_380 ( 
    i_10_380_174_0, i_10_380_175_0, i_10_380_178_0, i_10_380_264_0,
    i_10_380_265_0, i_10_380_268_0, i_10_380_284_0, i_10_380_289_0,
    i_10_380_315_0, i_10_380_316_0, i_10_380_324_0, i_10_380_446_0,
    i_10_380_464_0, i_10_380_503_0, i_10_380_629_0, i_10_380_718_0,
    i_10_380_748_0, i_10_380_754_0, i_10_380_931_0, i_10_380_997_0,
    i_10_380_1121_0, i_10_380_1221_0, i_10_380_1237_0, i_10_380_1239_0,
    i_10_380_1361_0, i_10_380_1432_0, i_10_380_1435_0, i_10_380_1438_0,
    i_10_380_1539_0, i_10_380_1581_0, i_10_380_1627_0, i_10_380_1650_0,
    i_10_380_1651_0, i_10_380_1652_0, i_10_380_1683_0, i_10_380_1686_0,
    i_10_380_1687_0, i_10_380_1689_0, i_10_380_1713_0, i_10_380_1717_0,
    i_10_380_1769_0, i_10_380_1819_0, i_10_380_1821_0, i_10_380_1823_0,
    i_10_380_1948_0, i_10_380_2032_0, i_10_380_2346_0, i_10_380_2347_0,
    i_10_380_2352_0, i_10_380_2362_0, i_10_380_2363_0, i_10_380_2451_0,
    i_10_380_2452_0, i_10_380_2471_0, i_10_380_2631_0, i_10_380_2632_0,
    i_10_380_2659_0, i_10_380_2709_0, i_10_380_2710_0, i_10_380_2727_0,
    i_10_380_2734_0, i_10_380_2735_0, i_10_380_2823_0, i_10_380_2850_0,
    i_10_380_2888_0, i_10_380_2919_0, i_10_380_2965_0, i_10_380_2967_0,
    i_10_380_2968_0, i_10_380_2980_0, i_10_380_3043_0, i_10_380_3049_0,
    i_10_380_3070_0, i_10_380_3199_0, i_10_380_3281_0, i_10_380_3283_0,
    i_10_380_3284_0, i_10_380_3380_0, i_10_380_3392_0, i_10_380_3504_0,
    i_10_380_3612_0, i_10_380_3781_0, i_10_380_3784_0, i_10_380_3840_0,
    i_10_380_3985_0, i_10_380_3993_0, i_10_380_4026_0, i_10_380_4113_0,
    i_10_380_4115_0, i_10_380_4119_0, i_10_380_4149_0, i_10_380_4173_0,
    i_10_380_4174_0, i_10_380_4212_0, i_10_380_4219_0, i_10_380_4269_0,
    i_10_380_4272_0, i_10_380_4276_0, i_10_380_4288_0, i_10_380_4571_0,
    o_10_380_0_0  );
  input  i_10_380_174_0, i_10_380_175_0, i_10_380_178_0, i_10_380_264_0,
    i_10_380_265_0, i_10_380_268_0, i_10_380_284_0, i_10_380_289_0,
    i_10_380_315_0, i_10_380_316_0, i_10_380_324_0, i_10_380_446_0,
    i_10_380_464_0, i_10_380_503_0, i_10_380_629_0, i_10_380_718_0,
    i_10_380_748_0, i_10_380_754_0, i_10_380_931_0, i_10_380_997_0,
    i_10_380_1121_0, i_10_380_1221_0, i_10_380_1237_0, i_10_380_1239_0,
    i_10_380_1361_0, i_10_380_1432_0, i_10_380_1435_0, i_10_380_1438_0,
    i_10_380_1539_0, i_10_380_1581_0, i_10_380_1627_0, i_10_380_1650_0,
    i_10_380_1651_0, i_10_380_1652_0, i_10_380_1683_0, i_10_380_1686_0,
    i_10_380_1687_0, i_10_380_1689_0, i_10_380_1713_0, i_10_380_1717_0,
    i_10_380_1769_0, i_10_380_1819_0, i_10_380_1821_0, i_10_380_1823_0,
    i_10_380_1948_0, i_10_380_2032_0, i_10_380_2346_0, i_10_380_2347_0,
    i_10_380_2352_0, i_10_380_2362_0, i_10_380_2363_0, i_10_380_2451_0,
    i_10_380_2452_0, i_10_380_2471_0, i_10_380_2631_0, i_10_380_2632_0,
    i_10_380_2659_0, i_10_380_2709_0, i_10_380_2710_0, i_10_380_2727_0,
    i_10_380_2734_0, i_10_380_2735_0, i_10_380_2823_0, i_10_380_2850_0,
    i_10_380_2888_0, i_10_380_2919_0, i_10_380_2965_0, i_10_380_2967_0,
    i_10_380_2968_0, i_10_380_2980_0, i_10_380_3043_0, i_10_380_3049_0,
    i_10_380_3070_0, i_10_380_3199_0, i_10_380_3281_0, i_10_380_3283_0,
    i_10_380_3284_0, i_10_380_3380_0, i_10_380_3392_0, i_10_380_3504_0,
    i_10_380_3612_0, i_10_380_3781_0, i_10_380_3784_0, i_10_380_3840_0,
    i_10_380_3985_0, i_10_380_3993_0, i_10_380_4026_0, i_10_380_4113_0,
    i_10_380_4115_0, i_10_380_4119_0, i_10_380_4149_0, i_10_380_4173_0,
    i_10_380_4174_0, i_10_380_4212_0, i_10_380_4219_0, i_10_380_4269_0,
    i_10_380_4272_0, i_10_380_4276_0, i_10_380_4288_0, i_10_380_4571_0;
  output o_10_380_0_0;
  assign o_10_380_0_0 = 0;
endmodule



// Benchmark "kernel_10_381" written by ABC on Sun Jul 19 10:27:40 2020

module kernel_10_381 ( 
    i_10_381_176_0, i_10_381_178_0, i_10_381_185_0, i_10_381_187_0,
    i_10_381_188_0, i_10_381_213_0, i_10_381_390_0, i_10_381_408_0,
    i_10_381_410_0, i_10_381_430_0, i_10_381_431_0, i_10_381_508_0,
    i_10_381_511_0, i_10_381_512_0, i_10_381_795_0, i_10_381_796_0,
    i_10_381_957_0, i_10_381_997_0, i_10_381_1028_0, i_10_381_1032_0,
    i_10_381_1042_0, i_10_381_1043_0, i_10_381_1141_0, i_10_381_1142_0,
    i_10_381_1237_0, i_10_381_1238_0, i_10_381_1261_0, i_10_381_1305_0,
    i_10_381_1308_0, i_10_381_1310_0, i_10_381_1365_0, i_10_381_1366_0,
    i_10_381_1367_0, i_10_381_1487_0, i_10_381_1580_0, i_10_381_1582_0,
    i_10_381_1583_0, i_10_381_1653_0, i_10_381_1683_0, i_10_381_1823_0,
    i_10_381_1824_0, i_10_381_1825_0, i_10_381_1913_0, i_10_381_2021_0,
    i_10_381_2185_0, i_10_381_2186_0, i_10_381_2309_0, i_10_381_2355_0,
    i_10_381_2453_0, i_10_381_2703_0, i_10_381_2705_0, i_10_381_2706_0,
    i_10_381_2707_0, i_10_381_2708_0, i_10_381_2716_0, i_10_381_2717_0,
    i_10_381_2730_0, i_10_381_2732_0, i_10_381_2734_0, i_10_381_2830_0,
    i_10_381_2831_0, i_10_381_2833_0, i_10_381_2870_0, i_10_381_2919_0,
    i_10_381_3037_0, i_10_381_3041_0, i_10_381_3151_0, i_10_381_3152_0,
    i_10_381_3199_0, i_10_381_3200_0, i_10_381_3270_0, i_10_381_3271_0,
    i_10_381_3284_0, i_10_381_3387_0, i_10_381_3388_0, i_10_381_3389_0,
    i_10_381_3390_0, i_10_381_3406_0, i_10_381_3523_0, i_10_381_3611_0,
    i_10_381_3614_0, i_10_381_3617_0, i_10_381_3651_0, i_10_381_3788_0,
    i_10_381_3895_0, i_10_381_3896_0, i_10_381_3991_0, i_10_381_4031_0,
    i_10_381_4119_0, i_10_381_4171_0, i_10_381_4172_0, i_10_381_4175_0,
    i_10_381_4182_0, i_10_381_4183_0, i_10_381_4192_0, i_10_381_4272_0,
    i_10_381_4273_0, i_10_381_4280_0, i_10_381_4282_0, i_10_381_4283_0,
    o_10_381_0_0  );
  input  i_10_381_176_0, i_10_381_178_0, i_10_381_185_0, i_10_381_187_0,
    i_10_381_188_0, i_10_381_213_0, i_10_381_390_0, i_10_381_408_0,
    i_10_381_410_0, i_10_381_430_0, i_10_381_431_0, i_10_381_508_0,
    i_10_381_511_0, i_10_381_512_0, i_10_381_795_0, i_10_381_796_0,
    i_10_381_957_0, i_10_381_997_0, i_10_381_1028_0, i_10_381_1032_0,
    i_10_381_1042_0, i_10_381_1043_0, i_10_381_1141_0, i_10_381_1142_0,
    i_10_381_1237_0, i_10_381_1238_0, i_10_381_1261_0, i_10_381_1305_0,
    i_10_381_1308_0, i_10_381_1310_0, i_10_381_1365_0, i_10_381_1366_0,
    i_10_381_1367_0, i_10_381_1487_0, i_10_381_1580_0, i_10_381_1582_0,
    i_10_381_1583_0, i_10_381_1653_0, i_10_381_1683_0, i_10_381_1823_0,
    i_10_381_1824_0, i_10_381_1825_0, i_10_381_1913_0, i_10_381_2021_0,
    i_10_381_2185_0, i_10_381_2186_0, i_10_381_2309_0, i_10_381_2355_0,
    i_10_381_2453_0, i_10_381_2703_0, i_10_381_2705_0, i_10_381_2706_0,
    i_10_381_2707_0, i_10_381_2708_0, i_10_381_2716_0, i_10_381_2717_0,
    i_10_381_2730_0, i_10_381_2732_0, i_10_381_2734_0, i_10_381_2830_0,
    i_10_381_2831_0, i_10_381_2833_0, i_10_381_2870_0, i_10_381_2919_0,
    i_10_381_3037_0, i_10_381_3041_0, i_10_381_3151_0, i_10_381_3152_0,
    i_10_381_3199_0, i_10_381_3200_0, i_10_381_3270_0, i_10_381_3271_0,
    i_10_381_3284_0, i_10_381_3387_0, i_10_381_3388_0, i_10_381_3389_0,
    i_10_381_3390_0, i_10_381_3406_0, i_10_381_3523_0, i_10_381_3611_0,
    i_10_381_3614_0, i_10_381_3617_0, i_10_381_3651_0, i_10_381_3788_0,
    i_10_381_3895_0, i_10_381_3896_0, i_10_381_3991_0, i_10_381_4031_0,
    i_10_381_4119_0, i_10_381_4171_0, i_10_381_4172_0, i_10_381_4175_0,
    i_10_381_4182_0, i_10_381_4183_0, i_10_381_4192_0, i_10_381_4272_0,
    i_10_381_4273_0, i_10_381_4280_0, i_10_381_4282_0, i_10_381_4283_0;
  output o_10_381_0_0;
  assign o_10_381_0_0 = ~((~i_10_381_2833_0 & ((~i_10_381_408_0 & ((~i_10_381_1043_0 & ~i_10_381_2453_0 & ~i_10_381_2716_0 & ~i_10_381_2734_0 & ~i_10_381_2830_0) | (~i_10_381_997_0 & ~i_10_381_1028_0 & ~i_10_381_1042_0 & ~i_10_381_1305_0 & ~i_10_381_2919_0 & ~i_10_381_3200_0 & ~i_10_381_4175_0))) | (~i_10_381_2703_0 & i_10_381_3284_0 & ~i_10_381_3611_0 & ~i_10_381_4172_0 & ~i_10_381_4280_0))) | (~i_10_381_1032_0 & ((~i_10_381_410_0 & ~i_10_381_1028_0 & ~i_10_381_1653_0 & ~i_10_381_2705_0) | (~i_10_381_188_0 & ~i_10_381_1683_0 & ~i_10_381_2919_0 & ~i_10_381_3991_0 & ~i_10_381_4171_0 & ~i_10_381_4280_0))) | (~i_10_381_1366_0 & ((~i_10_381_1028_0 & ~i_10_381_1261_0 & ~i_10_381_1487_0 & ~i_10_381_2021_0 & ~i_10_381_3284_0 & ~i_10_381_3617_0 & ~i_10_381_3896_0) | (~i_10_381_176_0 & ~i_10_381_1043_0 & ~i_10_381_2717_0 & ~i_10_381_2831_0 & ~i_10_381_3200_0 & ~i_10_381_4175_0))) | (~i_10_381_1367_0 & ~i_10_381_1823_0 & ((~i_10_381_997_0 & ~i_10_381_1028_0 & ~i_10_381_1042_0 & ~i_10_381_1487_0 & ~i_10_381_3284_0 & ~i_10_381_4171_0) | (~i_10_381_795_0 & i_10_381_1237_0 & ~i_10_381_2831_0 & ~i_10_381_4175_0))) | (~i_10_381_1028_0 & ((~i_10_381_1653_0 & i_10_381_1683_0 & ~i_10_381_2708_0 & ~i_10_381_3406_0) | (i_10_381_1825_0 & ~i_10_381_2453_0 & ~i_10_381_3614_0 & i_10_381_4272_0))) | (~i_10_381_1487_0 & ((~i_10_381_2705_0 & ~i_10_381_3896_0 & ~i_10_381_4119_0 & ~i_10_381_4272_0 & ~i_10_381_4282_0) | (~i_10_381_1308_0 & ~i_10_381_2732_0 & ~i_10_381_2919_0 & ~i_10_381_3895_0 & ~i_10_381_4172_0 & ~i_10_381_4283_0))) | (i_10_381_3388_0 & (~i_10_381_4172_0 | ~i_10_381_4283_0)) | (~i_10_381_3896_0 & ((i_10_381_796_0 & ~i_10_381_2453_0 & ~i_10_381_4119_0) | (i_10_381_2703_0 & ~i_10_381_2732_0 & ~i_10_381_3199_0 & ~i_10_381_3895_0 & ~i_10_381_4172_0))) | (~i_10_381_1238_0 & ~i_10_381_2707_0 & ~i_10_381_2708_0 & ~i_10_381_4280_0));
endmodule



// Benchmark "kernel_10_382" written by ABC on Sun Jul 19 10:27:41 2020

module kernel_10_382 ( 
    i_10_382_15_0, i_10_382_48_0, i_10_382_219_0, i_10_382_222_0,
    i_10_382_264_0, i_10_382_285_0, i_10_382_286_0, i_10_382_316_0,
    i_10_382_321_0, i_10_382_374_0, i_10_382_387_0, i_10_382_390_0,
    i_10_382_408_0, i_10_382_623_0, i_10_382_626_0, i_10_382_750_0,
    i_10_382_800_0, i_10_382_961_0, i_10_382_1049_0, i_10_382_1233_0,
    i_10_382_1234_0, i_10_382_1240_0, i_10_382_1296_0, i_10_382_1312_0,
    i_10_382_1346_0, i_10_382_1544_0, i_10_382_1549_0, i_10_382_1550_0,
    i_10_382_1686_0, i_10_382_1731_0, i_10_382_1732_0, i_10_382_1764_0,
    i_10_382_1810_0, i_10_382_1980_0, i_10_382_1990_0, i_10_382_2028_0,
    i_10_382_2031_0, i_10_382_2198_0, i_10_382_2199_0, i_10_382_2201_0,
    i_10_382_2349_0, i_10_382_2350_0, i_10_382_2352_0, i_10_382_2353_0,
    i_10_382_2364_0, i_10_382_2448_0, i_10_382_2458_0, i_10_382_2466_0,
    i_10_382_2469_0, i_10_382_2470_0, i_10_382_2472_0, i_10_382_2514_0,
    i_10_382_2565_0, i_10_382_2568_0, i_10_382_2570_0, i_10_382_2571_0,
    i_10_382_2628_0, i_10_382_2730_0, i_10_382_2781_0, i_10_382_2819_0,
    i_10_382_2822_0, i_10_382_2839_0, i_10_382_2880_0, i_10_382_2881_0,
    i_10_382_2982_0, i_10_382_3039_0, i_10_382_3087_0, i_10_382_3277_0,
    i_10_382_3283_0, i_10_382_3315_0, i_10_382_3318_0, i_10_382_3353_0,
    i_10_382_3392_0, i_10_382_3465_0, i_10_382_3468_0, i_10_382_3471_0,
    i_10_382_3507_0, i_10_382_3519_0, i_10_382_3543_0, i_10_382_3555_0,
    i_10_382_3582_0, i_10_382_3583_0, i_10_382_3585_0, i_10_382_3616_0,
    i_10_382_3838_0, i_10_382_3840_0, i_10_382_3980_0, i_10_382_4113_0,
    i_10_382_4115_0, i_10_382_4123_0, i_10_382_4168_0, i_10_382_4170_0,
    i_10_382_4266_0, i_10_382_4276_0, i_10_382_4285_0, i_10_382_4289_0,
    i_10_382_4290_0, i_10_382_4374_0, i_10_382_4461_0, i_10_382_4585_0,
    o_10_382_0_0  );
  input  i_10_382_15_0, i_10_382_48_0, i_10_382_219_0, i_10_382_222_0,
    i_10_382_264_0, i_10_382_285_0, i_10_382_286_0, i_10_382_316_0,
    i_10_382_321_0, i_10_382_374_0, i_10_382_387_0, i_10_382_390_0,
    i_10_382_408_0, i_10_382_623_0, i_10_382_626_0, i_10_382_750_0,
    i_10_382_800_0, i_10_382_961_0, i_10_382_1049_0, i_10_382_1233_0,
    i_10_382_1234_0, i_10_382_1240_0, i_10_382_1296_0, i_10_382_1312_0,
    i_10_382_1346_0, i_10_382_1544_0, i_10_382_1549_0, i_10_382_1550_0,
    i_10_382_1686_0, i_10_382_1731_0, i_10_382_1732_0, i_10_382_1764_0,
    i_10_382_1810_0, i_10_382_1980_0, i_10_382_1990_0, i_10_382_2028_0,
    i_10_382_2031_0, i_10_382_2198_0, i_10_382_2199_0, i_10_382_2201_0,
    i_10_382_2349_0, i_10_382_2350_0, i_10_382_2352_0, i_10_382_2353_0,
    i_10_382_2364_0, i_10_382_2448_0, i_10_382_2458_0, i_10_382_2466_0,
    i_10_382_2469_0, i_10_382_2470_0, i_10_382_2472_0, i_10_382_2514_0,
    i_10_382_2565_0, i_10_382_2568_0, i_10_382_2570_0, i_10_382_2571_0,
    i_10_382_2628_0, i_10_382_2730_0, i_10_382_2781_0, i_10_382_2819_0,
    i_10_382_2822_0, i_10_382_2839_0, i_10_382_2880_0, i_10_382_2881_0,
    i_10_382_2982_0, i_10_382_3039_0, i_10_382_3087_0, i_10_382_3277_0,
    i_10_382_3283_0, i_10_382_3315_0, i_10_382_3318_0, i_10_382_3353_0,
    i_10_382_3392_0, i_10_382_3465_0, i_10_382_3468_0, i_10_382_3471_0,
    i_10_382_3507_0, i_10_382_3519_0, i_10_382_3543_0, i_10_382_3555_0,
    i_10_382_3582_0, i_10_382_3583_0, i_10_382_3585_0, i_10_382_3616_0,
    i_10_382_3838_0, i_10_382_3840_0, i_10_382_3980_0, i_10_382_4113_0,
    i_10_382_4115_0, i_10_382_4123_0, i_10_382_4168_0, i_10_382_4170_0,
    i_10_382_4266_0, i_10_382_4276_0, i_10_382_4285_0, i_10_382_4289_0,
    i_10_382_4290_0, i_10_382_4374_0, i_10_382_4461_0, i_10_382_4585_0;
  output o_10_382_0_0;
  assign o_10_382_0_0 = 0;
endmodule



// Benchmark "kernel_10_383" written by ABC on Sun Jul 19 10:27:42 2020

module kernel_10_383 ( 
    i_10_383_9_0, i_10_383_16_0, i_10_383_66_0, i_10_383_67_0,
    i_10_383_69_0, i_10_383_148_0, i_10_383_159_0, i_10_383_160_0,
    i_10_383_224_0, i_10_383_237_0, i_10_383_245_0, i_10_383_251_0,
    i_10_383_253_0, i_10_383_256_0, i_10_383_261_0, i_10_383_270_0,
    i_10_383_290_0, i_10_383_293_0, i_10_383_318_0, i_10_383_321_0,
    i_10_383_331_0, i_10_383_368_0, i_10_383_373_0, i_10_383_393_0,
    i_10_383_519_0, i_10_383_541_0, i_10_383_627_0, i_10_383_688_0,
    i_10_383_721_0, i_10_383_823_0, i_10_383_1029_0, i_10_383_1030_0,
    i_10_383_1042_0, i_10_383_1110_0, i_10_383_1221_0, i_10_383_1239_0,
    i_10_383_1296_0, i_10_383_1299_0, i_10_383_1306_0, i_10_383_1359_0,
    i_10_383_1362_0, i_10_383_1431_0, i_10_383_1435_0, i_10_383_1438_0,
    i_10_383_1445_0, i_10_383_1513_0, i_10_383_1540_0, i_10_383_1553_0,
    i_10_383_1612_0, i_10_383_1798_0, i_10_383_1876_0, i_10_383_1879_0,
    i_10_383_1956_0, i_10_383_1966_0, i_10_383_2019_0, i_10_383_2022_0,
    i_10_383_2023_0, i_10_383_2196_0, i_10_383_2202_0, i_10_383_2203_0,
    i_10_383_2207_0, i_10_383_2326_0, i_10_383_2533_0, i_10_383_2535_0,
    i_10_383_2554_0, i_10_383_2565_0, i_10_383_2569_0, i_10_383_2587_0,
    i_10_383_2676_0, i_10_383_2709_0, i_10_383_2713_0, i_10_383_2724_0,
    i_10_383_2806_0, i_10_383_2913_0, i_10_383_2914_0, i_10_383_2989_0,
    i_10_383_2992_0, i_10_383_3072_0, i_10_383_3073_0, i_10_383_3177_0,
    i_10_383_3201_0, i_10_383_3268_0, i_10_383_3297_0, i_10_383_3469_0,
    i_10_383_3470_0, i_10_383_3472_0, i_10_383_3473_0, i_10_383_3504_0,
    i_10_383_3615_0, i_10_383_3777_0, i_10_383_3793_0, i_10_383_3814_0,
    i_10_383_3815_0, i_10_383_3840_0, i_10_383_3850_0, i_10_383_4120_0,
    i_10_383_4171_0, i_10_383_4174_0, i_10_383_4400_0, i_10_383_4587_0,
    o_10_383_0_0  );
  input  i_10_383_9_0, i_10_383_16_0, i_10_383_66_0, i_10_383_67_0,
    i_10_383_69_0, i_10_383_148_0, i_10_383_159_0, i_10_383_160_0,
    i_10_383_224_0, i_10_383_237_0, i_10_383_245_0, i_10_383_251_0,
    i_10_383_253_0, i_10_383_256_0, i_10_383_261_0, i_10_383_270_0,
    i_10_383_290_0, i_10_383_293_0, i_10_383_318_0, i_10_383_321_0,
    i_10_383_331_0, i_10_383_368_0, i_10_383_373_0, i_10_383_393_0,
    i_10_383_519_0, i_10_383_541_0, i_10_383_627_0, i_10_383_688_0,
    i_10_383_721_0, i_10_383_823_0, i_10_383_1029_0, i_10_383_1030_0,
    i_10_383_1042_0, i_10_383_1110_0, i_10_383_1221_0, i_10_383_1239_0,
    i_10_383_1296_0, i_10_383_1299_0, i_10_383_1306_0, i_10_383_1359_0,
    i_10_383_1362_0, i_10_383_1431_0, i_10_383_1435_0, i_10_383_1438_0,
    i_10_383_1445_0, i_10_383_1513_0, i_10_383_1540_0, i_10_383_1553_0,
    i_10_383_1612_0, i_10_383_1798_0, i_10_383_1876_0, i_10_383_1879_0,
    i_10_383_1956_0, i_10_383_1966_0, i_10_383_2019_0, i_10_383_2022_0,
    i_10_383_2023_0, i_10_383_2196_0, i_10_383_2202_0, i_10_383_2203_0,
    i_10_383_2207_0, i_10_383_2326_0, i_10_383_2533_0, i_10_383_2535_0,
    i_10_383_2554_0, i_10_383_2565_0, i_10_383_2569_0, i_10_383_2587_0,
    i_10_383_2676_0, i_10_383_2709_0, i_10_383_2713_0, i_10_383_2724_0,
    i_10_383_2806_0, i_10_383_2913_0, i_10_383_2914_0, i_10_383_2989_0,
    i_10_383_2992_0, i_10_383_3072_0, i_10_383_3073_0, i_10_383_3177_0,
    i_10_383_3201_0, i_10_383_3268_0, i_10_383_3297_0, i_10_383_3469_0,
    i_10_383_3470_0, i_10_383_3472_0, i_10_383_3473_0, i_10_383_3504_0,
    i_10_383_3615_0, i_10_383_3777_0, i_10_383_3793_0, i_10_383_3814_0,
    i_10_383_3815_0, i_10_383_3840_0, i_10_383_3850_0, i_10_383_4120_0,
    i_10_383_4171_0, i_10_383_4174_0, i_10_383_4400_0, i_10_383_4587_0;
  output o_10_383_0_0;
  assign o_10_383_0_0 = 0;
endmodule



// Benchmark "kernel_10_384" written by ABC on Sun Jul 19 10:27:43 2020

module kernel_10_384 ( 
    i_10_384_118_0, i_10_384_124_0, i_10_384_247_0, i_10_384_280_0,
    i_10_384_321_0, i_10_384_322_0, i_10_384_323_0, i_10_384_388_0,
    i_10_384_389_0, i_10_384_424_0, i_10_384_433_0, i_10_384_436_0,
    i_10_384_445_0, i_10_384_446_0, i_10_384_506_0, i_10_384_507_0,
    i_10_384_508_0, i_10_384_509_0, i_10_384_565_0, i_10_384_713_0,
    i_10_384_755_0, i_10_384_797_0, i_10_384_893_0, i_10_384_954_0,
    i_10_384_990_0, i_10_384_1027_0, i_10_384_1031_0, i_10_384_1043_0,
    i_10_384_1237_0, i_10_384_1309_0, i_10_384_1310_0, i_10_384_1575_0,
    i_10_384_1647_0, i_10_384_1648_0, i_10_384_1650_0, i_10_384_1691_0,
    i_10_384_1818_0, i_10_384_1819_0, i_10_384_1821_0, i_10_384_1822_0,
    i_10_384_2002_0, i_10_384_2197_0, i_10_384_2199_0, i_10_384_2357_0,
    i_10_384_2361_0, i_10_384_2410_0, i_10_384_2451_0, i_10_384_2452_0,
    i_10_384_2453_0, i_10_384_2467_0, i_10_384_2468_0, i_10_384_2700_0,
    i_10_384_2701_0, i_10_384_2702_0, i_10_384_2707_0, i_10_384_2709_0,
    i_10_384_2716_0, i_10_384_2817_0, i_10_384_2818_0, i_10_384_2826_0,
    i_10_384_2830_0, i_10_384_2883_0, i_10_384_2884_0, i_10_384_3037_0,
    i_10_384_3069_0, i_10_384_3088_0, i_10_384_3152_0, i_10_384_3278_0,
    i_10_384_3280_0, i_10_384_3281_0, i_10_384_3385_0, i_10_384_3386_0,
    i_10_384_3389_0, i_10_384_3390_0, i_10_384_3403_0, i_10_384_3404_0,
    i_10_384_3409_0, i_10_384_3583_0, i_10_384_3613_0, i_10_384_3614_0,
    i_10_384_3648_0, i_10_384_3650_0, i_10_384_3682_0, i_10_384_3835_0,
    i_10_384_3839_0, i_10_384_3847_0, i_10_384_3848_0, i_10_384_3851_0,
    i_10_384_3856_0, i_10_384_3860_0, i_10_384_3983_0, i_10_384_3992_0,
    i_10_384_4126_0, i_10_384_4127_0, i_10_384_4277_0, i_10_384_4292_0,
    i_10_384_4564_0, i_10_384_4565_0, i_10_384_4567_0, i_10_384_4568_0,
    o_10_384_0_0  );
  input  i_10_384_118_0, i_10_384_124_0, i_10_384_247_0, i_10_384_280_0,
    i_10_384_321_0, i_10_384_322_0, i_10_384_323_0, i_10_384_388_0,
    i_10_384_389_0, i_10_384_424_0, i_10_384_433_0, i_10_384_436_0,
    i_10_384_445_0, i_10_384_446_0, i_10_384_506_0, i_10_384_507_0,
    i_10_384_508_0, i_10_384_509_0, i_10_384_565_0, i_10_384_713_0,
    i_10_384_755_0, i_10_384_797_0, i_10_384_893_0, i_10_384_954_0,
    i_10_384_990_0, i_10_384_1027_0, i_10_384_1031_0, i_10_384_1043_0,
    i_10_384_1237_0, i_10_384_1309_0, i_10_384_1310_0, i_10_384_1575_0,
    i_10_384_1647_0, i_10_384_1648_0, i_10_384_1650_0, i_10_384_1691_0,
    i_10_384_1818_0, i_10_384_1819_0, i_10_384_1821_0, i_10_384_1822_0,
    i_10_384_2002_0, i_10_384_2197_0, i_10_384_2199_0, i_10_384_2357_0,
    i_10_384_2361_0, i_10_384_2410_0, i_10_384_2451_0, i_10_384_2452_0,
    i_10_384_2453_0, i_10_384_2467_0, i_10_384_2468_0, i_10_384_2700_0,
    i_10_384_2701_0, i_10_384_2702_0, i_10_384_2707_0, i_10_384_2709_0,
    i_10_384_2716_0, i_10_384_2817_0, i_10_384_2818_0, i_10_384_2826_0,
    i_10_384_2830_0, i_10_384_2883_0, i_10_384_2884_0, i_10_384_3037_0,
    i_10_384_3069_0, i_10_384_3088_0, i_10_384_3152_0, i_10_384_3278_0,
    i_10_384_3280_0, i_10_384_3281_0, i_10_384_3385_0, i_10_384_3386_0,
    i_10_384_3389_0, i_10_384_3390_0, i_10_384_3403_0, i_10_384_3404_0,
    i_10_384_3409_0, i_10_384_3583_0, i_10_384_3613_0, i_10_384_3614_0,
    i_10_384_3648_0, i_10_384_3650_0, i_10_384_3682_0, i_10_384_3835_0,
    i_10_384_3839_0, i_10_384_3847_0, i_10_384_3848_0, i_10_384_3851_0,
    i_10_384_3856_0, i_10_384_3860_0, i_10_384_3983_0, i_10_384_3992_0,
    i_10_384_4126_0, i_10_384_4127_0, i_10_384_4277_0, i_10_384_4292_0,
    i_10_384_4564_0, i_10_384_4565_0, i_10_384_4567_0, i_10_384_4568_0;
  output o_10_384_0_0;
  assign o_10_384_0_0 = ~((~i_10_384_323_0 & ((~i_10_384_322_0 & ((~i_10_384_389_0 & i_10_384_1027_0 & ~i_10_384_2818_0) | (~i_10_384_2453_0 & ~i_10_384_2467_0 & ~i_10_384_2817_0 & ~i_10_384_2883_0 & ~i_10_384_3088_0 & ~i_10_384_3281_0))) | (~i_10_384_1691_0 & ~i_10_384_2451_0 & ~i_10_384_2468_0 & ~i_10_384_3088_0 & ~i_10_384_3389_0 & i_10_384_3860_0))) | (i_10_384_445_0 & ((i_10_384_2709_0 & ~i_10_384_3281_0 & ~i_10_384_3613_0) | (i_10_384_446_0 & ~i_10_384_2467_0 & ~i_10_384_2818_0 & ~i_10_384_2883_0 & ~i_10_384_3280_0 & ~i_10_384_3648_0 & i_10_384_3856_0))) | (~i_10_384_565_0 & ((~i_10_384_436_0 & ~i_10_384_445_0 & i_10_384_1818_0 & ~i_10_384_2818_0 & ~i_10_384_3088_0) | (~i_10_384_424_0 & ~i_10_384_2884_0 & i_10_384_3847_0))) | (~i_10_384_3281_0 & ((~i_10_384_436_0 & ((~i_10_384_1237_0 & ~i_10_384_1650_0 & i_10_384_1821_0 & i_10_384_3613_0) | (~i_10_384_2199_0 & ~i_10_384_2451_0 & ~i_10_384_2452_0 & ~i_10_384_2716_0 & ~i_10_384_3390_0 & ~i_10_384_3583_0 & ~i_10_384_3847_0 & ~i_10_384_3860_0))) | (~i_10_384_2817_0 & ((~i_10_384_118_0 & ~i_10_384_797_0 & ~i_10_384_2707_0 & ~i_10_384_2826_0 & ~i_10_384_3278_0 & ~i_10_384_3280_0 & ~i_10_384_3835_0 & ~i_10_384_3847_0) | (~i_10_384_1819_0 & ~i_10_384_2467_0 & ~i_10_384_2818_0 & i_10_384_3385_0 & ~i_10_384_3390_0 & ~i_10_384_3404_0 & ~i_10_384_3992_0))))) | (~i_10_384_3409_0 & ((~i_10_384_118_0 & ((i_10_384_1237_0 & ~i_10_384_1822_0 & ~i_10_384_2357_0 & ~i_10_384_2451_0 & ~i_10_384_3278_0) | (~i_10_384_713_0 & ~i_10_384_1031_0 & ~i_10_384_1310_0 & ~i_10_384_1650_0 & ~i_10_384_1821_0 & ~i_10_384_2361_0 & ~i_10_384_2883_0 & ~i_10_384_3404_0 & ~i_10_384_4126_0))) | (~i_10_384_1821_0 & i_10_384_2451_0 & i_10_384_2817_0 & ~i_10_384_3278_0 & i_10_384_3856_0))) | (~i_10_384_1031_0 & ((~i_10_384_424_0 & ~i_10_384_1309_0 & i_10_384_1819_0 & ~i_10_384_3278_0) | (~i_10_384_446_0 & ~i_10_384_1043_0 & i_10_384_3037_0 & ~i_10_384_3280_0 & ~i_10_384_3386_0 & ~i_10_384_3390_0 & ~i_10_384_3583_0 & i_10_384_3650_0 & ~i_10_384_3860_0 & ~i_10_384_4565_0))) | (~i_10_384_424_0 & ((~i_10_384_713_0 & ~i_10_384_755_0 & ~i_10_384_1043_0 & ~i_10_384_2357_0 & ~i_10_384_2716_0 & ~i_10_384_2818_0 & ~i_10_384_2883_0 & ~i_10_384_2884_0 & ~i_10_384_3037_0) | (~i_10_384_1237_0 & ~i_10_384_3403_0 & ~i_10_384_3583_0 & i_10_384_3835_0 & ~i_10_384_3856_0))) | (i_10_384_1650_0 & ((~i_10_384_1309_0 & ~i_10_384_2884_0 & ~i_10_384_3278_0 & i_10_384_3409_0) | (i_10_384_2709_0 & ~i_10_384_2817_0 & ~i_10_384_3614_0))) | (~i_10_384_2451_0 & ((i_10_384_2701_0 & ~i_10_384_3037_0) | (i_10_384_1237_0 & i_10_384_1310_0 & ~i_10_384_1691_0 & ~i_10_384_2361_0 & ~i_10_384_2818_0 & ~i_10_384_2830_0 & ~i_10_384_2884_0 & ~i_10_384_3088_0))) | (~i_10_384_2467_0 & ((~i_10_384_1237_0 & ~i_10_384_1310_0 & i_10_384_1648_0) | (~i_10_384_2707_0 & i_10_384_3278_0 & ~i_10_384_3390_0 & ~i_10_384_3614_0 & ~i_10_384_3856_0))) | (~i_10_384_2818_0 & ~i_10_384_2883_0 & ~i_10_384_2884_0 & ((i_10_384_1819_0 & ~i_10_384_3088_0 & ~i_10_384_3613_0 & i_10_384_3835_0) | (~i_10_384_433_0 & ~i_10_384_2357_0 & ~i_10_384_2707_0 & ~i_10_384_2817_0 & ~i_10_384_2830_0 & ~i_10_384_3278_0 & ~i_10_384_3385_0 & ~i_10_384_3386_0 & ~i_10_384_3848_0))));
endmodule



// Benchmark "kernel_10_385" written by ABC on Sun Jul 19 10:27:44 2020

module kernel_10_385 ( 
    i_10_385_125_0, i_10_385_132_0, i_10_385_174_0, i_10_385_178_0,
    i_10_385_250_0, i_10_385_251_0, i_10_385_268_0, i_10_385_282_0,
    i_10_385_318_0, i_10_385_391_0, i_10_385_393_0, i_10_385_394_0,
    i_10_385_395_0, i_10_385_409_0, i_10_385_436_0, i_10_385_441_0,
    i_10_385_442_0, i_10_385_448_0, i_10_385_561_0, i_10_385_564_0,
    i_10_385_733_0, i_10_385_734_0, i_10_385_736_0, i_10_385_795_0,
    i_10_385_798_0, i_10_385_800_0, i_10_385_825_0, i_10_385_967_0,
    i_10_385_970_0, i_10_385_1002_0, i_10_385_1005_0, i_10_385_1006_0,
    i_10_385_1033_0, i_10_385_1113_0, i_10_385_1164_0, i_10_385_1233_0,
    i_10_385_1247_0, i_10_385_1306_0, i_10_385_1500_0, i_10_385_1689_0,
    i_10_385_1767_0, i_10_385_1821_0, i_10_385_1822_0, i_10_385_1920_0,
    i_10_385_2004_0, i_10_385_2351_0, i_10_385_2354_0, i_10_385_2361_0,
    i_10_385_2362_0, i_10_385_2381_0, i_10_385_2407_0, i_10_385_2448_0,
    i_10_385_2449_0, i_10_385_2453_0, i_10_385_2455_0, i_10_385_2518_0,
    i_10_385_2562_0, i_10_385_2630_0, i_10_385_2636_0, i_10_385_2662_0,
    i_10_385_2711_0, i_10_385_2725_0, i_10_385_2730_0, i_10_385_2732_0,
    i_10_385_2734_0, i_10_385_2833_0, i_10_385_2888_0, i_10_385_2955_0,
    i_10_385_2983_0, i_10_385_3042_0, i_10_385_3043_0, i_10_385_3049_0,
    i_10_385_3074_0, i_10_385_3283_0, i_10_385_3390_0, i_10_385_3437_0,
    i_10_385_3471_0, i_10_385_3472_0, i_10_385_3541_0, i_10_385_3542_0,
    i_10_385_3586_0, i_10_385_3588_0, i_10_385_3589_0, i_10_385_3612_0,
    i_10_385_3814_0, i_10_385_3850_0, i_10_385_3930_0, i_10_385_3985_0,
    i_10_385_3990_0, i_10_385_4024_0, i_10_385_4056_0, i_10_385_4057_0,
    i_10_385_4116_0, i_10_385_4117_0, i_10_385_4272_0, i_10_385_4292_0,
    i_10_385_4374_0, i_10_385_4570_0, i_10_385_4597_0, i_10_385_4598_0,
    o_10_385_0_0  );
  input  i_10_385_125_0, i_10_385_132_0, i_10_385_174_0, i_10_385_178_0,
    i_10_385_250_0, i_10_385_251_0, i_10_385_268_0, i_10_385_282_0,
    i_10_385_318_0, i_10_385_391_0, i_10_385_393_0, i_10_385_394_0,
    i_10_385_395_0, i_10_385_409_0, i_10_385_436_0, i_10_385_441_0,
    i_10_385_442_0, i_10_385_448_0, i_10_385_561_0, i_10_385_564_0,
    i_10_385_733_0, i_10_385_734_0, i_10_385_736_0, i_10_385_795_0,
    i_10_385_798_0, i_10_385_800_0, i_10_385_825_0, i_10_385_967_0,
    i_10_385_970_0, i_10_385_1002_0, i_10_385_1005_0, i_10_385_1006_0,
    i_10_385_1033_0, i_10_385_1113_0, i_10_385_1164_0, i_10_385_1233_0,
    i_10_385_1247_0, i_10_385_1306_0, i_10_385_1500_0, i_10_385_1689_0,
    i_10_385_1767_0, i_10_385_1821_0, i_10_385_1822_0, i_10_385_1920_0,
    i_10_385_2004_0, i_10_385_2351_0, i_10_385_2354_0, i_10_385_2361_0,
    i_10_385_2362_0, i_10_385_2381_0, i_10_385_2407_0, i_10_385_2448_0,
    i_10_385_2449_0, i_10_385_2453_0, i_10_385_2455_0, i_10_385_2518_0,
    i_10_385_2562_0, i_10_385_2630_0, i_10_385_2636_0, i_10_385_2662_0,
    i_10_385_2711_0, i_10_385_2725_0, i_10_385_2730_0, i_10_385_2732_0,
    i_10_385_2734_0, i_10_385_2833_0, i_10_385_2888_0, i_10_385_2955_0,
    i_10_385_2983_0, i_10_385_3042_0, i_10_385_3043_0, i_10_385_3049_0,
    i_10_385_3074_0, i_10_385_3283_0, i_10_385_3390_0, i_10_385_3437_0,
    i_10_385_3471_0, i_10_385_3472_0, i_10_385_3541_0, i_10_385_3542_0,
    i_10_385_3586_0, i_10_385_3588_0, i_10_385_3589_0, i_10_385_3612_0,
    i_10_385_3814_0, i_10_385_3850_0, i_10_385_3930_0, i_10_385_3985_0,
    i_10_385_3990_0, i_10_385_4024_0, i_10_385_4056_0, i_10_385_4057_0,
    i_10_385_4116_0, i_10_385_4117_0, i_10_385_4272_0, i_10_385_4292_0,
    i_10_385_4374_0, i_10_385_4570_0, i_10_385_4597_0, i_10_385_4598_0;
  output o_10_385_0_0;
  assign o_10_385_0_0 = 0;
endmodule



// Benchmark "kernel_10_386" written by ABC on Sun Jul 19 10:27:46 2020

module kernel_10_386 ( 
    i_10_386_172_0, i_10_386_183_0, i_10_386_265_0, i_10_386_275_0,
    i_10_386_327_0, i_10_386_328_0, i_10_386_390_0, i_10_386_393_0,
    i_10_386_394_0, i_10_386_408_0, i_10_386_427_0, i_10_386_429_0,
    i_10_386_437_0, i_10_386_440_0, i_10_386_538_0, i_10_386_539_0,
    i_10_386_701_0, i_10_386_735_0, i_10_386_755_0, i_10_386_996_0,
    i_10_386_997_0, i_10_386_1002_0, i_10_386_1003_0, i_10_386_1087_0,
    i_10_386_1138_0, i_10_386_1141_0, i_10_386_1168_0, i_10_386_1233_0,
    i_10_386_1264_0, i_10_386_1348_0, i_10_386_1349_0, i_10_386_1434_0,
    i_10_386_1435_0, i_10_386_1445_0, i_10_386_1555_0, i_10_386_1652_0,
    i_10_386_1655_0, i_10_386_1717_0, i_10_386_1769_0, i_10_386_1772_0,
    i_10_386_1818_0, i_10_386_1822_0, i_10_386_1823_0, i_10_386_1912_0,
    i_10_386_1913_0, i_10_386_1948_0, i_10_386_1949_0, i_10_386_2181_0,
    i_10_386_2184_0, i_10_386_2185_0, i_10_386_2199_0, i_10_386_2204_0,
    i_10_386_2311_0, i_10_386_2312_0, i_10_386_2329_0, i_10_386_2406_0,
    i_10_386_2407_0, i_10_386_2408_0, i_10_386_2455_0, i_10_386_2469_0,
    i_10_386_2481_0, i_10_386_2629_0, i_10_386_2631_0, i_10_386_2657_0,
    i_10_386_2679_0, i_10_386_2713_0, i_10_386_2716_0, i_10_386_2833_0,
    i_10_386_2919_0, i_10_386_2921_0, i_10_386_2922_0, i_10_386_2923_0,
    i_10_386_2982_0, i_10_386_2983_0, i_10_386_3041_0, i_10_386_3047_0,
    i_10_386_3093_0, i_10_386_3094_0, i_10_386_3152_0, i_10_386_3154_0,
    i_10_386_3155_0, i_10_386_3210_0, i_10_386_3472_0, i_10_386_3473_0,
    i_10_386_3497_0, i_10_386_3543_0, i_10_386_3544_0, i_10_386_3588_0,
    i_10_386_3855_0, i_10_386_3856_0, i_10_386_3859_0, i_10_386_4057_0,
    i_10_386_4114_0, i_10_386_4117_0, i_10_386_4175_0, i_10_386_4236_0,
    i_10_386_4238_0, i_10_386_4290_0, i_10_386_4291_0, i_10_386_4533_0,
    o_10_386_0_0  );
  input  i_10_386_172_0, i_10_386_183_0, i_10_386_265_0, i_10_386_275_0,
    i_10_386_327_0, i_10_386_328_0, i_10_386_390_0, i_10_386_393_0,
    i_10_386_394_0, i_10_386_408_0, i_10_386_427_0, i_10_386_429_0,
    i_10_386_437_0, i_10_386_440_0, i_10_386_538_0, i_10_386_539_0,
    i_10_386_701_0, i_10_386_735_0, i_10_386_755_0, i_10_386_996_0,
    i_10_386_997_0, i_10_386_1002_0, i_10_386_1003_0, i_10_386_1087_0,
    i_10_386_1138_0, i_10_386_1141_0, i_10_386_1168_0, i_10_386_1233_0,
    i_10_386_1264_0, i_10_386_1348_0, i_10_386_1349_0, i_10_386_1434_0,
    i_10_386_1435_0, i_10_386_1445_0, i_10_386_1555_0, i_10_386_1652_0,
    i_10_386_1655_0, i_10_386_1717_0, i_10_386_1769_0, i_10_386_1772_0,
    i_10_386_1818_0, i_10_386_1822_0, i_10_386_1823_0, i_10_386_1912_0,
    i_10_386_1913_0, i_10_386_1948_0, i_10_386_1949_0, i_10_386_2181_0,
    i_10_386_2184_0, i_10_386_2185_0, i_10_386_2199_0, i_10_386_2204_0,
    i_10_386_2311_0, i_10_386_2312_0, i_10_386_2329_0, i_10_386_2406_0,
    i_10_386_2407_0, i_10_386_2408_0, i_10_386_2455_0, i_10_386_2469_0,
    i_10_386_2481_0, i_10_386_2629_0, i_10_386_2631_0, i_10_386_2657_0,
    i_10_386_2679_0, i_10_386_2713_0, i_10_386_2716_0, i_10_386_2833_0,
    i_10_386_2919_0, i_10_386_2921_0, i_10_386_2922_0, i_10_386_2923_0,
    i_10_386_2982_0, i_10_386_2983_0, i_10_386_3041_0, i_10_386_3047_0,
    i_10_386_3093_0, i_10_386_3094_0, i_10_386_3152_0, i_10_386_3154_0,
    i_10_386_3155_0, i_10_386_3210_0, i_10_386_3472_0, i_10_386_3473_0,
    i_10_386_3497_0, i_10_386_3543_0, i_10_386_3544_0, i_10_386_3588_0,
    i_10_386_3855_0, i_10_386_3856_0, i_10_386_3859_0, i_10_386_4057_0,
    i_10_386_4114_0, i_10_386_4117_0, i_10_386_4175_0, i_10_386_4236_0,
    i_10_386_4238_0, i_10_386_4290_0, i_10_386_4291_0, i_10_386_4533_0;
  output o_10_386_0_0;
  assign o_10_386_0_0 = ~((~i_10_386_4236_0 & ((~i_10_386_3497_0 & ((~i_10_386_390_0 & ((~i_10_386_437_0 & ~i_10_386_3093_0) | (~i_10_386_1349_0 & ~i_10_386_3588_0))) | (~i_10_386_1913_0 & ~i_10_386_2716_0 & ~i_10_386_3093_0))) | (~i_10_386_427_0 & i_10_386_1435_0 & ~i_10_386_4175_0 & ~i_10_386_4238_0))) | (~i_10_386_1445_0 & ((~i_10_386_265_0 & ~i_10_386_394_0 & ~i_10_386_1349_0 & ~i_10_386_2406_0) | (~i_10_386_701_0 & ~i_10_386_2408_0 & ~i_10_386_2469_0 & ~i_10_386_3543_0 & i_10_386_3856_0))) | (~i_10_386_394_0 & ~i_10_386_4290_0 & ((~i_10_386_1264_0 & ~i_10_386_1822_0 & ~i_10_386_2982_0) | (~i_10_386_427_0 & ~i_10_386_1348_0 & ~i_10_386_2312_0 & ~i_10_386_3041_0 & ~i_10_386_4238_0))) | (~i_10_386_2312_0 & i_10_386_2923_0) | (~i_10_386_2408_0 & i_10_386_2629_0 & ~i_10_386_3093_0) | (~i_10_386_1003_0 & ~i_10_386_1435_0 & ~i_10_386_1772_0 & ~i_10_386_2713_0 & ~i_10_386_3473_0 & ~i_10_386_4238_0) | (~i_10_386_327_0 & ~i_10_386_2311_0 & ~i_10_386_3544_0 & ~i_10_386_4057_0) | (~i_10_386_429_0 & ~i_10_386_1002_0 & ~i_10_386_3047_0 & ~i_10_386_3094_0 & ~i_10_386_3856_0 & ~i_10_386_4114_0) | (~i_10_386_997_0 & ~i_10_386_1769_0 & ~i_10_386_2204_0 & ~i_10_386_2407_0 & ~i_10_386_2481_0 & ~i_10_386_4117_0) | (~i_10_386_1912_0 & ~i_10_386_3588_0 & i_10_386_4291_0));
endmodule



// Benchmark "kernel_10_387" written by ABC on Sun Jul 19 10:27:46 2020

module kernel_10_387 ( 
    i_10_387_45_0, i_10_387_48_0, i_10_387_120_0, i_10_387_144_0,
    i_10_387_145_0, i_10_387_177_0, i_10_387_219_0, i_10_387_246_0,
    i_10_387_280_0, i_10_387_285_0, i_10_387_286_0, i_10_387_315_0,
    i_10_387_373_0, i_10_387_448_0, i_10_387_449_0, i_10_387_461_0,
    i_10_387_462_0, i_10_387_467_0, i_10_387_747_0, i_10_387_796_0,
    i_10_387_797_0, i_10_387_798_0, i_10_387_799_0, i_10_387_967_0,
    i_10_387_981_0, i_10_387_1030_0, i_10_387_1242_0, i_10_387_1266_0,
    i_10_387_1305_0, i_10_387_1309_0, i_10_387_1342_0, i_10_387_1446_0,
    i_10_387_1482_0, i_10_387_1578_0, i_10_387_1629_0, i_10_387_1632_0,
    i_10_387_1638_0, i_10_387_1686_0, i_10_387_1689_0, i_10_387_1791_0,
    i_10_387_1916_0, i_10_387_1925_0, i_10_387_1951_0, i_10_387_1952_0,
    i_10_387_2025_0, i_10_387_2311_0, i_10_387_2312_0, i_10_387_2349_0,
    i_10_387_2350_0, i_10_387_2469_0, i_10_387_2565_0, i_10_387_2628_0,
    i_10_387_2638_0, i_10_387_2658_0, i_10_387_2659_0, i_10_387_2673_0,
    i_10_387_2700_0, i_10_387_2721_0, i_10_387_2727_0, i_10_387_2728_0,
    i_10_387_2817_0, i_10_387_2969_0, i_10_387_3043_0, i_10_387_3114_0,
    i_10_387_3277_0, i_10_387_3283_0, i_10_387_3312_0, i_10_387_3348_0,
    i_10_387_3360_0, i_10_387_3384_0, i_10_387_3387_0, i_10_387_3388_0,
    i_10_387_3393_0, i_10_387_3468_0, i_10_387_3471_0, i_10_387_3504_0,
    i_10_387_3585_0, i_10_387_3619_0, i_10_387_3652_0, i_10_387_3784_0,
    i_10_387_3843_0, i_10_387_3844_0, i_10_387_3845_0, i_10_387_3847_0,
    i_10_387_3856_0, i_10_387_3870_0, i_10_387_3913_0, i_10_387_4030_0,
    i_10_387_4116_0, i_10_387_4117_0, i_10_387_4125_0, i_10_387_4129_0,
    i_10_387_4152_0, i_10_387_4153_0, i_10_387_4170_0, i_10_387_4267_0,
    i_10_387_4275_0, i_10_387_4284_0, i_10_387_4290_0, i_10_387_4565_0,
    o_10_387_0_0  );
  input  i_10_387_45_0, i_10_387_48_0, i_10_387_120_0, i_10_387_144_0,
    i_10_387_145_0, i_10_387_177_0, i_10_387_219_0, i_10_387_246_0,
    i_10_387_280_0, i_10_387_285_0, i_10_387_286_0, i_10_387_315_0,
    i_10_387_373_0, i_10_387_448_0, i_10_387_449_0, i_10_387_461_0,
    i_10_387_462_0, i_10_387_467_0, i_10_387_747_0, i_10_387_796_0,
    i_10_387_797_0, i_10_387_798_0, i_10_387_799_0, i_10_387_967_0,
    i_10_387_981_0, i_10_387_1030_0, i_10_387_1242_0, i_10_387_1266_0,
    i_10_387_1305_0, i_10_387_1309_0, i_10_387_1342_0, i_10_387_1446_0,
    i_10_387_1482_0, i_10_387_1578_0, i_10_387_1629_0, i_10_387_1632_0,
    i_10_387_1638_0, i_10_387_1686_0, i_10_387_1689_0, i_10_387_1791_0,
    i_10_387_1916_0, i_10_387_1925_0, i_10_387_1951_0, i_10_387_1952_0,
    i_10_387_2025_0, i_10_387_2311_0, i_10_387_2312_0, i_10_387_2349_0,
    i_10_387_2350_0, i_10_387_2469_0, i_10_387_2565_0, i_10_387_2628_0,
    i_10_387_2638_0, i_10_387_2658_0, i_10_387_2659_0, i_10_387_2673_0,
    i_10_387_2700_0, i_10_387_2721_0, i_10_387_2727_0, i_10_387_2728_0,
    i_10_387_2817_0, i_10_387_2969_0, i_10_387_3043_0, i_10_387_3114_0,
    i_10_387_3277_0, i_10_387_3283_0, i_10_387_3312_0, i_10_387_3348_0,
    i_10_387_3360_0, i_10_387_3384_0, i_10_387_3387_0, i_10_387_3388_0,
    i_10_387_3393_0, i_10_387_3468_0, i_10_387_3471_0, i_10_387_3504_0,
    i_10_387_3585_0, i_10_387_3619_0, i_10_387_3652_0, i_10_387_3784_0,
    i_10_387_3843_0, i_10_387_3844_0, i_10_387_3845_0, i_10_387_3847_0,
    i_10_387_3856_0, i_10_387_3870_0, i_10_387_3913_0, i_10_387_4030_0,
    i_10_387_4116_0, i_10_387_4117_0, i_10_387_4125_0, i_10_387_4129_0,
    i_10_387_4152_0, i_10_387_4153_0, i_10_387_4170_0, i_10_387_4267_0,
    i_10_387_4275_0, i_10_387_4284_0, i_10_387_4290_0, i_10_387_4565_0;
  output o_10_387_0_0;
  assign o_10_387_0_0 = 0;
endmodule



// Benchmark "kernel_10_388" written by ABC on Sun Jul 19 10:27:47 2020

module kernel_10_388 ( 
    i_10_388_150_0, i_10_388_256_0, i_10_388_294_0, i_10_388_409_0,
    i_10_388_410_0, i_10_388_429_0, i_10_388_430_0, i_10_388_438_0,
    i_10_388_439_0, i_10_388_447_0, i_10_388_627_0, i_10_388_645_0,
    i_10_388_796_0, i_10_388_798_0, i_10_388_799_0, i_10_388_897_0,
    i_10_388_1033_0, i_10_388_1051_0, i_10_388_1203_0, i_10_388_1245_0,
    i_10_388_1249_0, i_10_388_1364_0, i_10_388_1367_0, i_10_388_1384_0,
    i_10_388_1444_0, i_10_388_1552_0, i_10_388_1608_0, i_10_388_1618_0,
    i_10_388_1650_0, i_10_388_1653_0, i_10_388_1808_0, i_10_388_1822_0,
    i_10_388_1915_0, i_10_388_1951_0, i_10_388_1995_0, i_10_388_1996_0,
    i_10_388_2265_0, i_10_388_2338_0, i_10_388_2350_0, i_10_388_2351_0,
    i_10_388_2352_0, i_10_388_2355_0, i_10_388_2356_0, i_10_388_2364_0,
    i_10_388_2446_0, i_10_388_2447_0, i_10_388_2451_0, i_10_388_2463_0,
    i_10_388_2481_0, i_10_388_2482_0, i_10_388_2514_0, i_10_388_2515_0,
    i_10_388_2543_0, i_10_388_2607_0, i_10_388_2634_0, i_10_388_2643_0,
    i_10_388_2644_0, i_10_388_2716_0, i_10_388_2717_0, i_10_388_2718_0,
    i_10_388_2720_0, i_10_388_2726_0, i_10_388_2731_0, i_10_388_2735_0,
    i_10_388_2866_0, i_10_388_2919_0, i_10_388_2920_0, i_10_388_2922_0,
    i_10_388_3165_0, i_10_388_3166_0, i_10_388_3175_0, i_10_388_3196_0,
    i_10_388_3228_0, i_10_388_3270_0, i_10_388_3276_0, i_10_388_3280_0,
    i_10_388_3281_0, i_10_388_3283_0, i_10_388_3544_0, i_10_388_3561_0,
    i_10_388_3610_0, i_10_388_3612_0, i_10_388_3613_0, i_10_388_3706_0,
    i_10_388_3785_0, i_10_388_3838_0, i_10_388_3855_0, i_10_388_3904_0,
    i_10_388_3991_0, i_10_388_3992_0, i_10_388_4026_0, i_10_388_4027_0,
    i_10_388_4028_0, i_10_388_4029_0, i_10_388_4215_0, i_10_388_4219_0,
    i_10_388_4236_0, i_10_388_4276_0, i_10_388_4291_0, i_10_388_4480_0,
    o_10_388_0_0  );
  input  i_10_388_150_0, i_10_388_256_0, i_10_388_294_0, i_10_388_409_0,
    i_10_388_410_0, i_10_388_429_0, i_10_388_430_0, i_10_388_438_0,
    i_10_388_439_0, i_10_388_447_0, i_10_388_627_0, i_10_388_645_0,
    i_10_388_796_0, i_10_388_798_0, i_10_388_799_0, i_10_388_897_0,
    i_10_388_1033_0, i_10_388_1051_0, i_10_388_1203_0, i_10_388_1245_0,
    i_10_388_1249_0, i_10_388_1364_0, i_10_388_1367_0, i_10_388_1384_0,
    i_10_388_1444_0, i_10_388_1552_0, i_10_388_1608_0, i_10_388_1618_0,
    i_10_388_1650_0, i_10_388_1653_0, i_10_388_1808_0, i_10_388_1822_0,
    i_10_388_1915_0, i_10_388_1951_0, i_10_388_1995_0, i_10_388_1996_0,
    i_10_388_2265_0, i_10_388_2338_0, i_10_388_2350_0, i_10_388_2351_0,
    i_10_388_2352_0, i_10_388_2355_0, i_10_388_2356_0, i_10_388_2364_0,
    i_10_388_2446_0, i_10_388_2447_0, i_10_388_2451_0, i_10_388_2463_0,
    i_10_388_2481_0, i_10_388_2482_0, i_10_388_2514_0, i_10_388_2515_0,
    i_10_388_2543_0, i_10_388_2607_0, i_10_388_2634_0, i_10_388_2643_0,
    i_10_388_2644_0, i_10_388_2716_0, i_10_388_2717_0, i_10_388_2718_0,
    i_10_388_2720_0, i_10_388_2726_0, i_10_388_2731_0, i_10_388_2735_0,
    i_10_388_2866_0, i_10_388_2919_0, i_10_388_2920_0, i_10_388_2922_0,
    i_10_388_3165_0, i_10_388_3166_0, i_10_388_3175_0, i_10_388_3196_0,
    i_10_388_3228_0, i_10_388_3270_0, i_10_388_3276_0, i_10_388_3280_0,
    i_10_388_3281_0, i_10_388_3283_0, i_10_388_3544_0, i_10_388_3561_0,
    i_10_388_3610_0, i_10_388_3612_0, i_10_388_3613_0, i_10_388_3706_0,
    i_10_388_3785_0, i_10_388_3838_0, i_10_388_3855_0, i_10_388_3904_0,
    i_10_388_3991_0, i_10_388_3992_0, i_10_388_4026_0, i_10_388_4027_0,
    i_10_388_4028_0, i_10_388_4029_0, i_10_388_4215_0, i_10_388_4219_0,
    i_10_388_4236_0, i_10_388_4276_0, i_10_388_4291_0, i_10_388_4480_0;
  output o_10_388_0_0;
  assign o_10_388_0_0 = 0;
endmodule



// Benchmark "kernel_10_389" written by ABC on Sun Jul 19 10:27:48 2020

module kernel_10_389 ( 
    i_10_389_35_0, i_10_389_71_0, i_10_389_242_0, i_10_389_251_0,
    i_10_389_275_0, i_10_389_283_0, i_10_389_284_0, i_10_389_285_0,
    i_10_389_368_0, i_10_389_448_0, i_10_389_466_0, i_10_389_467_0,
    i_10_389_545_0, i_10_389_719_0, i_10_389_752_0, i_10_389_800_0,
    i_10_389_954_0, i_10_389_959_0, i_10_389_1031_0, i_10_389_1032_0,
    i_10_389_1033_0, i_10_389_1034_0, i_10_389_1244_0, i_10_389_1248_0,
    i_10_389_1250_0, i_10_389_1345_0, i_10_389_1439_0, i_10_389_1448_0,
    i_10_389_1619_0, i_10_389_1687_0, i_10_389_1819_0, i_10_389_1822_0,
    i_10_389_1823_0, i_10_389_1825_0, i_10_389_1958_0, i_10_389_1961_0,
    i_10_389_1995_0, i_10_389_1996_0, i_10_389_2185_0, i_10_389_2186_0,
    i_10_389_2311_0, i_10_389_2312_0, i_10_389_2361_0, i_10_389_2363_0,
    i_10_389_2365_0, i_10_389_2470_0, i_10_389_2573_0, i_10_389_2609_0,
    i_10_389_2632_0, i_10_389_2658_0, i_10_389_2663_0, i_10_389_2704_0,
    i_10_389_2705_0, i_10_389_2708_0, i_10_389_2711_0, i_10_389_2714_0,
    i_10_389_2717_0, i_10_389_2732_0, i_10_389_2735_0, i_10_389_2744_0,
    i_10_389_2830_0, i_10_389_2831_0, i_10_389_3034_0, i_10_389_3037_0,
    i_10_389_3038_0, i_10_389_3077_0, i_10_389_3198_0, i_10_389_3199_0,
    i_10_389_3272_0, i_10_389_3275_0, i_10_389_3384_0, i_10_389_3389_0,
    i_10_389_3443_0, i_10_389_3446_0, i_10_389_3472_0, i_10_389_3525_0,
    i_10_389_3584_0, i_10_389_3613_0, i_10_389_3614_0, i_10_389_3784_0,
    i_10_389_3785_0, i_10_389_3787_0, i_10_389_3788_0, i_10_389_3840_0,
    i_10_389_3842_0, i_10_389_3848_0, i_10_389_3849_0, i_10_389_3855_0,
    i_10_389_3949_0, i_10_389_3991_0, i_10_389_4113_0, i_10_389_4114_0,
    i_10_389_4118_0, i_10_389_4121_0, i_10_389_4127_0, i_10_389_4170_0,
    i_10_389_4220_0, i_10_389_4280_0, i_10_389_4291_0, i_10_389_4571_0,
    o_10_389_0_0  );
  input  i_10_389_35_0, i_10_389_71_0, i_10_389_242_0, i_10_389_251_0,
    i_10_389_275_0, i_10_389_283_0, i_10_389_284_0, i_10_389_285_0,
    i_10_389_368_0, i_10_389_448_0, i_10_389_466_0, i_10_389_467_0,
    i_10_389_545_0, i_10_389_719_0, i_10_389_752_0, i_10_389_800_0,
    i_10_389_954_0, i_10_389_959_0, i_10_389_1031_0, i_10_389_1032_0,
    i_10_389_1033_0, i_10_389_1034_0, i_10_389_1244_0, i_10_389_1248_0,
    i_10_389_1250_0, i_10_389_1345_0, i_10_389_1439_0, i_10_389_1448_0,
    i_10_389_1619_0, i_10_389_1687_0, i_10_389_1819_0, i_10_389_1822_0,
    i_10_389_1823_0, i_10_389_1825_0, i_10_389_1958_0, i_10_389_1961_0,
    i_10_389_1995_0, i_10_389_1996_0, i_10_389_2185_0, i_10_389_2186_0,
    i_10_389_2311_0, i_10_389_2312_0, i_10_389_2361_0, i_10_389_2363_0,
    i_10_389_2365_0, i_10_389_2470_0, i_10_389_2573_0, i_10_389_2609_0,
    i_10_389_2632_0, i_10_389_2658_0, i_10_389_2663_0, i_10_389_2704_0,
    i_10_389_2705_0, i_10_389_2708_0, i_10_389_2711_0, i_10_389_2714_0,
    i_10_389_2717_0, i_10_389_2732_0, i_10_389_2735_0, i_10_389_2744_0,
    i_10_389_2830_0, i_10_389_2831_0, i_10_389_3034_0, i_10_389_3037_0,
    i_10_389_3038_0, i_10_389_3077_0, i_10_389_3198_0, i_10_389_3199_0,
    i_10_389_3272_0, i_10_389_3275_0, i_10_389_3384_0, i_10_389_3389_0,
    i_10_389_3443_0, i_10_389_3446_0, i_10_389_3472_0, i_10_389_3525_0,
    i_10_389_3584_0, i_10_389_3613_0, i_10_389_3614_0, i_10_389_3784_0,
    i_10_389_3785_0, i_10_389_3787_0, i_10_389_3788_0, i_10_389_3840_0,
    i_10_389_3842_0, i_10_389_3848_0, i_10_389_3849_0, i_10_389_3855_0,
    i_10_389_3949_0, i_10_389_3991_0, i_10_389_4113_0, i_10_389_4114_0,
    i_10_389_4118_0, i_10_389_4121_0, i_10_389_4127_0, i_10_389_4170_0,
    i_10_389_4220_0, i_10_389_4280_0, i_10_389_4291_0, i_10_389_4571_0;
  output o_10_389_0_0;
  assign o_10_389_0_0 = 0;
endmodule



// Benchmark "kernel_10_390" written by ABC on Sun Jul 19 10:27:49 2020

module kernel_10_390 ( 
    i_10_390_47_0, i_10_390_49_0, i_10_390_50_0, i_10_390_137_0,
    i_10_390_171_0, i_10_390_172_0, i_10_390_178_0, i_10_390_216_0,
    i_10_390_221_0, i_10_390_245_0, i_10_390_248_0, i_10_390_287_0,
    i_10_390_515_0, i_10_390_544_0, i_10_390_545_0, i_10_390_662_0,
    i_10_390_689_0, i_10_390_716_0, i_10_390_748_0, i_10_390_749_0,
    i_10_390_796_0, i_10_390_954_0, i_10_390_964_0, i_10_390_965_0,
    i_10_390_983_0, i_10_390_1028_0, i_10_390_1031_0, i_10_390_1181_0,
    i_10_390_1184_0, i_10_390_1217_0, i_10_390_1242_0, i_10_390_1244_0,
    i_10_390_1310_0, i_10_390_1355_0, i_10_390_1487_0, i_10_390_1531_0,
    i_10_390_1532_0, i_10_390_1541_0, i_10_390_1559_0, i_10_390_1580_0,
    i_10_390_1616_0, i_10_390_1653_0, i_10_390_1685_0, i_10_390_2003_0,
    i_10_390_2035_0, i_10_390_2081_0, i_10_390_2161_0, i_10_390_2305_0,
    i_10_390_2306_0, i_10_390_2308_0, i_10_390_2327_0, i_10_390_2330_0,
    i_10_390_2363_0, i_10_390_2458_0, i_10_390_2459_0, i_10_390_2463_0,
    i_10_390_2471_0, i_10_390_2473_0, i_10_390_2567_0, i_10_390_2602_0,
    i_10_390_2603_0, i_10_390_2630_0, i_10_390_2659_0, i_10_390_2660_0,
    i_10_390_2737_0, i_10_390_2738_0, i_10_390_3074_0, i_10_390_3199_0,
    i_10_390_3200_0, i_10_390_3233_0, i_10_390_3281_0, i_10_390_3290_0,
    i_10_390_3388_0, i_10_390_3406_0, i_10_390_3407_0, i_10_390_3445_0,
    i_10_390_3550_0, i_10_390_3584_0, i_10_390_3587_0, i_10_390_3610_0,
    i_10_390_3613_0, i_10_390_3614_0, i_10_390_3619_0, i_10_390_3620_0,
    i_10_390_3647_0, i_10_390_3800_0, i_10_390_3871_0, i_10_390_3908_0,
    i_10_390_3998_0, i_10_390_4064_0, i_10_390_4115_0, i_10_390_4126_0,
    i_10_390_4217_0, i_10_390_4220_0, i_10_390_4268_0, i_10_390_4276_0,
    i_10_390_4285_0, i_10_390_4287_0, i_10_390_4288_0, i_10_390_4289_0,
    o_10_390_0_0  );
  input  i_10_390_47_0, i_10_390_49_0, i_10_390_50_0, i_10_390_137_0,
    i_10_390_171_0, i_10_390_172_0, i_10_390_178_0, i_10_390_216_0,
    i_10_390_221_0, i_10_390_245_0, i_10_390_248_0, i_10_390_287_0,
    i_10_390_515_0, i_10_390_544_0, i_10_390_545_0, i_10_390_662_0,
    i_10_390_689_0, i_10_390_716_0, i_10_390_748_0, i_10_390_749_0,
    i_10_390_796_0, i_10_390_954_0, i_10_390_964_0, i_10_390_965_0,
    i_10_390_983_0, i_10_390_1028_0, i_10_390_1031_0, i_10_390_1181_0,
    i_10_390_1184_0, i_10_390_1217_0, i_10_390_1242_0, i_10_390_1244_0,
    i_10_390_1310_0, i_10_390_1355_0, i_10_390_1487_0, i_10_390_1531_0,
    i_10_390_1532_0, i_10_390_1541_0, i_10_390_1559_0, i_10_390_1580_0,
    i_10_390_1616_0, i_10_390_1653_0, i_10_390_1685_0, i_10_390_2003_0,
    i_10_390_2035_0, i_10_390_2081_0, i_10_390_2161_0, i_10_390_2305_0,
    i_10_390_2306_0, i_10_390_2308_0, i_10_390_2327_0, i_10_390_2330_0,
    i_10_390_2363_0, i_10_390_2458_0, i_10_390_2459_0, i_10_390_2463_0,
    i_10_390_2471_0, i_10_390_2473_0, i_10_390_2567_0, i_10_390_2602_0,
    i_10_390_2603_0, i_10_390_2630_0, i_10_390_2659_0, i_10_390_2660_0,
    i_10_390_2737_0, i_10_390_2738_0, i_10_390_3074_0, i_10_390_3199_0,
    i_10_390_3200_0, i_10_390_3233_0, i_10_390_3281_0, i_10_390_3290_0,
    i_10_390_3388_0, i_10_390_3406_0, i_10_390_3407_0, i_10_390_3445_0,
    i_10_390_3550_0, i_10_390_3584_0, i_10_390_3587_0, i_10_390_3610_0,
    i_10_390_3613_0, i_10_390_3614_0, i_10_390_3619_0, i_10_390_3620_0,
    i_10_390_3647_0, i_10_390_3800_0, i_10_390_3871_0, i_10_390_3908_0,
    i_10_390_3998_0, i_10_390_4064_0, i_10_390_4115_0, i_10_390_4126_0,
    i_10_390_4217_0, i_10_390_4220_0, i_10_390_4268_0, i_10_390_4276_0,
    i_10_390_4285_0, i_10_390_4287_0, i_10_390_4288_0, i_10_390_4289_0;
  output o_10_390_0_0;
  assign o_10_390_0_0 = 0;
endmodule



// Benchmark "kernel_10_391" written by ABC on Sun Jul 19 10:27:50 2020

module kernel_10_391 ( 
    i_10_391_47_0, i_10_391_51_0, i_10_391_83_0, i_10_391_155_0,
    i_10_391_217_0, i_10_391_220_0, i_10_391_245_0, i_10_391_281_0,
    i_10_391_283_0, i_10_391_286_0, i_10_391_319_0, i_10_391_329_0,
    i_10_391_389_0, i_10_391_409_0, i_10_391_434_0, i_10_391_436_0,
    i_10_391_441_0, i_10_391_442_0, i_10_391_462_0, i_10_391_465_0,
    i_10_391_639_0, i_10_391_640_0, i_10_391_643_0, i_10_391_985_0,
    i_10_391_1026_0, i_10_391_1029_0, i_10_391_1046_0, i_10_391_1059_0,
    i_10_391_1207_0, i_10_391_1237_0, i_10_391_1250_0, i_10_391_1264_0,
    i_10_391_1492_0, i_10_391_1543_0, i_10_391_1683_0, i_10_391_1689_0,
    i_10_391_1824_0, i_10_391_1825_0, i_10_391_1826_0, i_10_391_1915_0,
    i_10_391_1992_0, i_10_391_1999_0, i_10_391_2000_0, i_10_391_2016_0,
    i_10_391_2352_0, i_10_391_2436_0, i_10_391_2448_0, i_10_391_2449_0,
    i_10_391_2452_0, i_10_391_2464_0, i_10_391_2465_0, i_10_391_2628_0,
    i_10_391_2631_0, i_10_391_2642_0, i_10_391_2656_0, i_10_391_2659_0,
    i_10_391_2660_0, i_10_391_2674_0, i_10_391_2727_0, i_10_391_2728_0,
    i_10_391_2729_0, i_10_391_2819_0, i_10_391_2829_0, i_10_391_2830_0,
    i_10_391_2833_0, i_10_391_2963_0, i_10_391_2964_0, i_10_391_2982_0,
    i_10_391_2986_0, i_10_391_3045_0, i_10_391_3087_0, i_10_391_3088_0,
    i_10_391_3089_0, i_10_391_3094_0, i_10_391_3161_0, i_10_391_3233_0,
    i_10_391_3289_0, i_10_391_3388_0, i_10_391_3391_0, i_10_391_3434_0,
    i_10_391_3504_0, i_10_391_3522_0, i_10_391_3523_0, i_10_391_3524_0,
    i_10_391_3682_0, i_10_391_3700_0, i_10_391_3783_0, i_10_391_3809_0,
    i_10_391_3838_0, i_10_391_3856_0, i_10_391_3857_0, i_10_391_4029_0,
    i_10_391_4054_0, i_10_391_4127_0, i_10_391_4153_0, i_10_391_4172_0,
    i_10_391_4275_0, i_10_391_4280_0, i_10_391_4282_0, i_10_391_4292_0,
    o_10_391_0_0  );
  input  i_10_391_47_0, i_10_391_51_0, i_10_391_83_0, i_10_391_155_0,
    i_10_391_217_0, i_10_391_220_0, i_10_391_245_0, i_10_391_281_0,
    i_10_391_283_0, i_10_391_286_0, i_10_391_319_0, i_10_391_329_0,
    i_10_391_389_0, i_10_391_409_0, i_10_391_434_0, i_10_391_436_0,
    i_10_391_441_0, i_10_391_442_0, i_10_391_462_0, i_10_391_465_0,
    i_10_391_639_0, i_10_391_640_0, i_10_391_643_0, i_10_391_985_0,
    i_10_391_1026_0, i_10_391_1029_0, i_10_391_1046_0, i_10_391_1059_0,
    i_10_391_1207_0, i_10_391_1237_0, i_10_391_1250_0, i_10_391_1264_0,
    i_10_391_1492_0, i_10_391_1543_0, i_10_391_1683_0, i_10_391_1689_0,
    i_10_391_1824_0, i_10_391_1825_0, i_10_391_1826_0, i_10_391_1915_0,
    i_10_391_1992_0, i_10_391_1999_0, i_10_391_2000_0, i_10_391_2016_0,
    i_10_391_2352_0, i_10_391_2436_0, i_10_391_2448_0, i_10_391_2449_0,
    i_10_391_2452_0, i_10_391_2464_0, i_10_391_2465_0, i_10_391_2628_0,
    i_10_391_2631_0, i_10_391_2642_0, i_10_391_2656_0, i_10_391_2659_0,
    i_10_391_2660_0, i_10_391_2674_0, i_10_391_2727_0, i_10_391_2728_0,
    i_10_391_2729_0, i_10_391_2819_0, i_10_391_2829_0, i_10_391_2830_0,
    i_10_391_2833_0, i_10_391_2963_0, i_10_391_2964_0, i_10_391_2982_0,
    i_10_391_2986_0, i_10_391_3045_0, i_10_391_3087_0, i_10_391_3088_0,
    i_10_391_3089_0, i_10_391_3094_0, i_10_391_3161_0, i_10_391_3233_0,
    i_10_391_3289_0, i_10_391_3388_0, i_10_391_3391_0, i_10_391_3434_0,
    i_10_391_3504_0, i_10_391_3522_0, i_10_391_3523_0, i_10_391_3524_0,
    i_10_391_3682_0, i_10_391_3700_0, i_10_391_3783_0, i_10_391_3809_0,
    i_10_391_3838_0, i_10_391_3856_0, i_10_391_3857_0, i_10_391_4029_0,
    i_10_391_4054_0, i_10_391_4127_0, i_10_391_4153_0, i_10_391_4172_0,
    i_10_391_4275_0, i_10_391_4280_0, i_10_391_4282_0, i_10_391_4292_0;
  output o_10_391_0_0;
  assign o_10_391_0_0 = 0;
endmodule



// Benchmark "kernel_10_392" written by ABC on Sun Jul 19 10:27:51 2020

module kernel_10_392 ( 
    i_10_392_281_0, i_10_392_282_0, i_10_392_295_0, i_10_392_296_0,
    i_10_392_327_0, i_10_392_328_0, i_10_392_329_0, i_10_392_407_0,
    i_10_392_433_0, i_10_392_434_0, i_10_392_441_0, i_10_392_442_0,
    i_10_392_443_0, i_10_392_444_0, i_10_392_445_0, i_10_392_749_0,
    i_10_392_796_0, i_10_392_960_0, i_10_392_1233_0, i_10_392_1234_0,
    i_10_392_1235_0, i_10_392_1239_0, i_10_392_1263_0, i_10_392_1311_0,
    i_10_392_1312_0, i_10_392_1348_0, i_10_392_1431_0, i_10_392_1432_0,
    i_10_392_1447_0, i_10_392_1654_0, i_10_392_1767_0, i_10_392_1768_0,
    i_10_392_1819_0, i_10_392_1822_0, i_10_392_1823_0, i_10_392_1824_0,
    i_10_392_1825_0, i_10_392_1911_0, i_10_392_1912_0, i_10_392_1913_0,
    i_10_392_1946_0, i_10_392_2180_0, i_10_392_2457_0, i_10_392_2458_0,
    i_10_392_2470_0, i_10_392_2629_0, i_10_392_2630_0, i_10_392_2656_0,
    i_10_392_2658_0, i_10_392_2659_0, i_10_392_2663_0, i_10_392_2711_0,
    i_10_392_2716_0, i_10_392_2718_0, i_10_392_2719_0, i_10_392_2722_0,
    i_10_392_2723_0, i_10_392_2781_0, i_10_392_2782_0, i_10_392_2783_0,
    i_10_392_2817_0, i_10_392_2819_0, i_10_392_2826_0, i_10_392_2827_0,
    i_10_392_2830_0, i_10_392_2831_0, i_10_392_2923_0, i_10_392_2981_0,
    i_10_392_3033_0, i_10_392_3034_0, i_10_392_3035_0, i_10_392_3047_0,
    i_10_392_3196_0, i_10_392_3323_0, i_10_392_3392_0, i_10_392_3403_0,
    i_10_392_3409_0, i_10_392_3523_0, i_10_392_3583_0, i_10_392_3609_0,
    i_10_392_3612_0, i_10_392_3613_0, i_10_392_3682_0, i_10_392_3783_0,
    i_10_392_3785_0, i_10_392_3838_0, i_10_392_3839_0, i_10_392_3852_0,
    i_10_392_3853_0, i_10_392_3857_0, i_10_392_3906_0, i_10_392_3907_0,
    i_10_392_3991_0, i_10_392_4113_0, i_10_392_4116_0, i_10_392_4118_0,
    i_10_392_4267_0, i_10_392_4285_0, i_10_392_4288_0, i_10_392_4566_0,
    o_10_392_0_0  );
  input  i_10_392_281_0, i_10_392_282_0, i_10_392_295_0, i_10_392_296_0,
    i_10_392_327_0, i_10_392_328_0, i_10_392_329_0, i_10_392_407_0,
    i_10_392_433_0, i_10_392_434_0, i_10_392_441_0, i_10_392_442_0,
    i_10_392_443_0, i_10_392_444_0, i_10_392_445_0, i_10_392_749_0,
    i_10_392_796_0, i_10_392_960_0, i_10_392_1233_0, i_10_392_1234_0,
    i_10_392_1235_0, i_10_392_1239_0, i_10_392_1263_0, i_10_392_1311_0,
    i_10_392_1312_0, i_10_392_1348_0, i_10_392_1431_0, i_10_392_1432_0,
    i_10_392_1447_0, i_10_392_1654_0, i_10_392_1767_0, i_10_392_1768_0,
    i_10_392_1819_0, i_10_392_1822_0, i_10_392_1823_0, i_10_392_1824_0,
    i_10_392_1825_0, i_10_392_1911_0, i_10_392_1912_0, i_10_392_1913_0,
    i_10_392_1946_0, i_10_392_2180_0, i_10_392_2457_0, i_10_392_2458_0,
    i_10_392_2470_0, i_10_392_2629_0, i_10_392_2630_0, i_10_392_2656_0,
    i_10_392_2658_0, i_10_392_2659_0, i_10_392_2663_0, i_10_392_2711_0,
    i_10_392_2716_0, i_10_392_2718_0, i_10_392_2719_0, i_10_392_2722_0,
    i_10_392_2723_0, i_10_392_2781_0, i_10_392_2782_0, i_10_392_2783_0,
    i_10_392_2817_0, i_10_392_2819_0, i_10_392_2826_0, i_10_392_2827_0,
    i_10_392_2830_0, i_10_392_2831_0, i_10_392_2923_0, i_10_392_2981_0,
    i_10_392_3033_0, i_10_392_3034_0, i_10_392_3035_0, i_10_392_3047_0,
    i_10_392_3196_0, i_10_392_3323_0, i_10_392_3392_0, i_10_392_3403_0,
    i_10_392_3409_0, i_10_392_3523_0, i_10_392_3583_0, i_10_392_3609_0,
    i_10_392_3612_0, i_10_392_3613_0, i_10_392_3682_0, i_10_392_3783_0,
    i_10_392_3785_0, i_10_392_3838_0, i_10_392_3839_0, i_10_392_3852_0,
    i_10_392_3853_0, i_10_392_3857_0, i_10_392_3906_0, i_10_392_3907_0,
    i_10_392_3991_0, i_10_392_4113_0, i_10_392_4116_0, i_10_392_4118_0,
    i_10_392_4267_0, i_10_392_4285_0, i_10_392_4288_0, i_10_392_4566_0;
  output o_10_392_0_0;
  assign o_10_392_0_0 = ~((~i_10_392_3907_0 & ((~i_10_392_281_0 & ((~i_10_392_442_0 & ~i_10_392_445_0 & ~i_10_392_1234_0 & ~i_10_392_1767_0 & ~i_10_392_1822_0 & ~i_10_392_1946_0 & i_10_392_2830_0 & ~i_10_392_3392_0 & ~i_10_392_3409_0 & ~i_10_392_3523_0 & ~i_10_392_3612_0 & ~i_10_392_3906_0) | (~i_10_392_282_0 & i_10_392_1819_0 & ~i_10_392_3613_0 & ~i_10_392_4113_0))) | (~i_10_392_282_0 & ~i_10_392_1768_0 & ~i_10_392_3785_0 & ((~i_10_392_295_0 & ~i_10_392_327_0 & ~i_10_392_1312_0 & ~i_10_392_2629_0 & ~i_10_392_2630_0 & ~i_10_392_2817_0 & ~i_10_392_3047_0) | (~i_10_392_433_0 & ~i_10_392_434_0 & ~i_10_392_1233_0 & ~i_10_392_2830_0 & ~i_10_392_3392_0 & ~i_10_392_3783_0 & ~i_10_392_3838_0))) | (~i_10_392_296_0 & ~i_10_392_1911_0 & ~i_10_392_2458_0 & ~i_10_392_2656_0 & ~i_10_392_2718_0 & ~i_10_392_3613_0 & ~i_10_392_3838_0 & ~i_10_392_3857_0))) | (~i_10_392_282_0 & ~i_10_392_4116_0 & ((~i_10_392_1912_0 & ~i_10_392_2630_0 & ~i_10_392_3403_0 & ~i_10_392_3857_0 & ~i_10_392_4118_0) | (~i_10_392_1911_0 & ~i_10_392_2719_0 & ~i_10_392_3991_0 & i_10_392_4288_0))) | (~i_10_392_1767_0 & ((~i_10_392_327_0 & ((~i_10_392_434_0 & ~i_10_392_1654_0 & i_10_392_1825_0 & ~i_10_392_2718_0) | (~i_10_392_329_0 & ~i_10_392_749_0 & ~i_10_392_1348_0 & ~i_10_392_2457_0 & ~i_10_392_2711_0 & ~i_10_392_2719_0 & ~i_10_392_2923_0))) | (~i_10_392_433_0 & ~i_10_392_1912_0 & ~i_10_392_2719_0 & ~i_10_392_2830_0 & ~i_10_392_2981_0) | (~i_10_392_328_0 & ~i_10_392_1913_0 & ~i_10_392_2457_0 & ~i_10_392_2630_0 & ~i_10_392_2819_0 & ~i_10_392_3409_0 & ~i_10_392_3785_0 & ~i_10_392_3906_0))) | (~i_10_392_433_0 & ((~i_10_392_434_0 & ~i_10_392_1263_0 & ~i_10_392_3852_0 & ((~i_10_392_296_0 & ~i_10_392_1348_0 & ~i_10_392_1768_0 & ~i_10_392_2629_0 & ~i_10_392_2656_0 & ~i_10_392_2819_0 & ~i_10_392_3609_0 & ~i_10_392_3839_0) | (~i_10_392_1822_0 & ~i_10_392_3857_0 & i_10_392_4116_0))) | (~i_10_392_1912_0 & ~i_10_392_2457_0 & ~i_10_392_2658_0 & ~i_10_392_2819_0 & i_10_392_2827_0 & ~i_10_392_3047_0) | (~i_10_392_1911_0 & ~i_10_392_2817_0 & i_10_392_3852_0 & ~i_10_392_3857_0 & ~i_10_392_4285_0))) | (~i_10_392_2819_0 & ((~i_10_392_434_0 & ((~i_10_392_1768_0 & i_10_392_1819_0 & ~i_10_392_1823_0 & i_10_392_3853_0) | (~i_10_392_1912_0 & ~i_10_392_1913_0 & ~i_10_392_2716_0 & ~i_10_392_3609_0 & ~i_10_392_3853_0 & ~i_10_392_4113_0 & ~i_10_392_4566_0))) | (~i_10_392_328_0 & ~i_10_392_2457_0 & ~i_10_392_2711_0 & ~i_10_392_2723_0 & i_10_392_3853_0))) | (~i_10_392_4288_0 & ((~i_10_392_328_0 & ((i_10_392_1825_0 & ~i_10_392_3857_0) | (~i_10_392_445_0 & ~i_10_392_1768_0 & ~i_10_392_2711_0 & ~i_10_392_2981_0 & i_10_392_3852_0 & ~i_10_392_4566_0))) | (i_10_392_1825_0 & i_10_392_1913_0 & ~i_10_392_2723_0))) | (~i_10_392_1768_0 & ~i_10_392_3612_0 & ((i_10_392_1825_0 & i_10_392_3839_0) | (~i_10_392_1348_0 & ~i_10_392_1911_0 & ~i_10_392_2718_0 & ~i_10_392_2981_0 & ~i_10_392_3403_0 & ~i_10_392_3857_0 & ~i_10_392_4285_0 & ~i_10_392_4566_0))) | (~i_10_392_444_0 & i_10_392_1654_0 & ~i_10_392_1822_0 & ~i_10_392_2629_0 & ~i_10_392_2716_0) | (i_10_392_445_0 & ~i_10_392_1239_0 & ~i_10_392_1823_0 & ~i_10_392_2817_0 & ~i_10_392_2831_0 & ~i_10_392_2981_0) | (i_10_392_3196_0 & ~i_10_392_3609_0 & i_10_392_3991_0 & i_10_392_4118_0) | (~i_10_392_1912_0 & ~i_10_392_2711_0 & i_10_392_2719_0 & ~i_10_392_3783_0 & ~i_10_392_4113_0 & i_10_392_4288_0 & ~i_10_392_4566_0) | (i_10_392_444_0 & i_10_392_3838_0 & ~i_10_392_3839_0 & i_10_392_4566_0));
endmodule



// Benchmark "kernel_10_393" written by ABC on Sun Jul 19 10:27:52 2020

module kernel_10_393 ( 
    i_10_393_100_0, i_10_393_133_0, i_10_393_134_0, i_10_393_174_0,
    i_10_393_175_0, i_10_393_190_0, i_10_393_282_0, i_10_393_432_0,
    i_10_393_444_0, i_10_393_446_0, i_10_393_514_0, i_10_393_643_0,
    i_10_393_715_0, i_10_393_796_0, i_10_393_829_0, i_10_393_830_0,
    i_10_393_836_0, i_10_393_853_0, i_10_393_896_0, i_10_393_905_0,
    i_10_393_965_0, i_10_393_990_0, i_10_393_991_0, i_10_393_1051_0,
    i_10_393_1233_0, i_10_393_1289_0, i_10_393_1305_0, i_10_393_1306_0,
    i_10_393_1342_0, i_10_393_1366_0, i_10_393_1434_0, i_10_393_1478_0,
    i_10_393_1558_0, i_10_393_1640_0, i_10_393_1913_0, i_10_393_1949_0,
    i_10_393_1991_0, i_10_393_2020_0, i_10_393_2349_0, i_10_393_2351_0,
    i_10_393_2352_0, i_10_393_2353_0, i_10_393_2354_0, i_10_393_2363_0,
    i_10_393_2365_0, i_10_393_2366_0, i_10_393_2470_0, i_10_393_2515_0,
    i_10_393_2527_0, i_10_393_2539_0, i_10_393_2629_0, i_10_393_2675_0,
    i_10_393_2744_0, i_10_393_2817_0, i_10_393_2818_0, i_10_393_2855_0,
    i_10_393_2881_0, i_10_393_2917_0, i_10_393_2918_0, i_10_393_2921_0,
    i_10_393_2980_0, i_10_393_3083_0, i_10_393_3107_0, i_10_393_3114_0,
    i_10_393_3197_0, i_10_393_3269_0, i_10_393_3298_0, i_10_393_3352_0,
    i_10_393_3391_0, i_10_393_3392_0, i_10_393_3403_0, i_10_393_3443_0,
    i_10_393_3460_0, i_10_393_3471_0, i_10_393_3497_0, i_10_393_3502_0,
    i_10_393_3503_0, i_10_393_3539_0, i_10_393_3609_0, i_10_393_3612_0,
    i_10_393_3615_0, i_10_393_3617_0, i_10_393_3625_0, i_10_393_3626_0,
    i_10_393_3683_0, i_10_393_3729_0, i_10_393_3730_0, i_10_393_3731_0,
    i_10_393_3776_0, i_10_393_3833_0, i_10_393_3858_0, i_10_393_3899_0,
    i_10_393_4118_0, i_10_393_4185_0, i_10_393_4276_0, i_10_393_4277_0,
    i_10_393_4403_0, i_10_393_4457_0, i_10_393_4573_0, i_10_393_4583_0,
    o_10_393_0_0  );
  input  i_10_393_100_0, i_10_393_133_0, i_10_393_134_0, i_10_393_174_0,
    i_10_393_175_0, i_10_393_190_0, i_10_393_282_0, i_10_393_432_0,
    i_10_393_444_0, i_10_393_446_0, i_10_393_514_0, i_10_393_643_0,
    i_10_393_715_0, i_10_393_796_0, i_10_393_829_0, i_10_393_830_0,
    i_10_393_836_0, i_10_393_853_0, i_10_393_896_0, i_10_393_905_0,
    i_10_393_965_0, i_10_393_990_0, i_10_393_991_0, i_10_393_1051_0,
    i_10_393_1233_0, i_10_393_1289_0, i_10_393_1305_0, i_10_393_1306_0,
    i_10_393_1342_0, i_10_393_1366_0, i_10_393_1434_0, i_10_393_1478_0,
    i_10_393_1558_0, i_10_393_1640_0, i_10_393_1913_0, i_10_393_1949_0,
    i_10_393_1991_0, i_10_393_2020_0, i_10_393_2349_0, i_10_393_2351_0,
    i_10_393_2352_0, i_10_393_2353_0, i_10_393_2354_0, i_10_393_2363_0,
    i_10_393_2365_0, i_10_393_2366_0, i_10_393_2470_0, i_10_393_2515_0,
    i_10_393_2527_0, i_10_393_2539_0, i_10_393_2629_0, i_10_393_2675_0,
    i_10_393_2744_0, i_10_393_2817_0, i_10_393_2818_0, i_10_393_2855_0,
    i_10_393_2881_0, i_10_393_2917_0, i_10_393_2918_0, i_10_393_2921_0,
    i_10_393_2980_0, i_10_393_3083_0, i_10_393_3107_0, i_10_393_3114_0,
    i_10_393_3197_0, i_10_393_3269_0, i_10_393_3298_0, i_10_393_3352_0,
    i_10_393_3391_0, i_10_393_3392_0, i_10_393_3403_0, i_10_393_3443_0,
    i_10_393_3460_0, i_10_393_3471_0, i_10_393_3497_0, i_10_393_3502_0,
    i_10_393_3503_0, i_10_393_3539_0, i_10_393_3609_0, i_10_393_3612_0,
    i_10_393_3615_0, i_10_393_3617_0, i_10_393_3625_0, i_10_393_3626_0,
    i_10_393_3683_0, i_10_393_3729_0, i_10_393_3730_0, i_10_393_3731_0,
    i_10_393_3776_0, i_10_393_3833_0, i_10_393_3858_0, i_10_393_3899_0,
    i_10_393_4118_0, i_10_393_4185_0, i_10_393_4276_0, i_10_393_4277_0,
    i_10_393_4403_0, i_10_393_4457_0, i_10_393_4573_0, i_10_393_4583_0;
  output o_10_393_0_0;
  assign o_10_393_0_0 = 0;
endmodule



// Benchmark "kernel_10_394" written by ABC on Sun Jul 19 10:27:53 2020

module kernel_10_394 ( 
    i_10_394_82_0, i_10_394_119_0, i_10_394_122_0, i_10_394_223_0,
    i_10_394_282_0, i_10_394_327_0, i_10_394_328_0, i_10_394_360_0,
    i_10_394_387_0, i_10_394_388_0, i_10_394_390_0, i_10_394_434_0,
    i_10_394_436_0, i_10_394_437_0, i_10_394_446_0, i_10_394_447_0,
    i_10_394_459_0, i_10_394_463_0, i_10_394_464_0, i_10_394_903_0,
    i_10_394_962_0, i_10_394_990_0, i_10_394_1000_0, i_10_394_1027_0,
    i_10_394_1035_0, i_10_394_1036_0, i_10_394_1083_0, i_10_394_1241_0,
    i_10_394_1261_0, i_10_394_1380_0, i_10_394_1449_0, i_10_394_1450_0,
    i_10_394_1452_0, i_10_394_1530_0, i_10_394_1551_0, i_10_394_1654_0,
    i_10_394_1684_0, i_10_394_1685_0, i_10_394_1872_0, i_10_394_1873_0,
    i_10_394_1875_0, i_10_394_1911_0, i_10_394_2000_0, i_10_394_2181_0,
    i_10_394_2182_0, i_10_394_2224_0, i_10_394_2352_0, i_10_394_2377_0,
    i_10_394_2378_0, i_10_394_2403_0, i_10_394_2449_0, i_10_394_2453_0,
    i_10_394_2455_0, i_10_394_2602_0, i_10_394_2603_0, i_10_394_2628_0,
    i_10_394_2658_0, i_10_394_2673_0, i_10_394_2700_0, i_10_394_2718_0,
    i_10_394_2721_0, i_10_394_2731_0, i_10_394_2826_0, i_10_394_2827_0,
    i_10_394_2828_0, i_10_394_2829_0, i_10_394_2920_0, i_10_394_2923_0,
    i_10_394_3036_0, i_10_394_3037_0, i_10_394_3041_0, i_10_394_3042_0,
    i_10_394_3087_0, i_10_394_3159_0, i_10_394_3283_0, i_10_394_3384_0,
    i_10_394_3389_0, i_10_394_3432_0, i_10_394_3470_0, i_10_394_3522_0,
    i_10_394_3537_0, i_10_394_3560_0, i_10_394_3563_0, i_10_394_3685_0,
    i_10_394_3782_0, i_10_394_3784_0, i_10_394_3786_0, i_10_394_3787_0,
    i_10_394_3834_0, i_10_394_3855_0, i_10_394_3856_0, i_10_394_3892_0,
    i_10_394_3981_0, i_10_394_4025_0, i_10_394_4113_0, i_10_394_4213_0,
    i_10_394_4270_0, i_10_394_4279_0, i_10_394_4285_0, i_10_394_4288_0,
    o_10_394_0_0  );
  input  i_10_394_82_0, i_10_394_119_0, i_10_394_122_0, i_10_394_223_0,
    i_10_394_282_0, i_10_394_327_0, i_10_394_328_0, i_10_394_360_0,
    i_10_394_387_0, i_10_394_388_0, i_10_394_390_0, i_10_394_434_0,
    i_10_394_436_0, i_10_394_437_0, i_10_394_446_0, i_10_394_447_0,
    i_10_394_459_0, i_10_394_463_0, i_10_394_464_0, i_10_394_903_0,
    i_10_394_962_0, i_10_394_990_0, i_10_394_1000_0, i_10_394_1027_0,
    i_10_394_1035_0, i_10_394_1036_0, i_10_394_1083_0, i_10_394_1241_0,
    i_10_394_1261_0, i_10_394_1380_0, i_10_394_1449_0, i_10_394_1450_0,
    i_10_394_1452_0, i_10_394_1530_0, i_10_394_1551_0, i_10_394_1654_0,
    i_10_394_1684_0, i_10_394_1685_0, i_10_394_1872_0, i_10_394_1873_0,
    i_10_394_1875_0, i_10_394_1911_0, i_10_394_2000_0, i_10_394_2181_0,
    i_10_394_2182_0, i_10_394_2224_0, i_10_394_2352_0, i_10_394_2377_0,
    i_10_394_2378_0, i_10_394_2403_0, i_10_394_2449_0, i_10_394_2453_0,
    i_10_394_2455_0, i_10_394_2602_0, i_10_394_2603_0, i_10_394_2628_0,
    i_10_394_2658_0, i_10_394_2673_0, i_10_394_2700_0, i_10_394_2718_0,
    i_10_394_2721_0, i_10_394_2731_0, i_10_394_2826_0, i_10_394_2827_0,
    i_10_394_2828_0, i_10_394_2829_0, i_10_394_2920_0, i_10_394_2923_0,
    i_10_394_3036_0, i_10_394_3037_0, i_10_394_3041_0, i_10_394_3042_0,
    i_10_394_3087_0, i_10_394_3159_0, i_10_394_3283_0, i_10_394_3384_0,
    i_10_394_3389_0, i_10_394_3432_0, i_10_394_3470_0, i_10_394_3522_0,
    i_10_394_3537_0, i_10_394_3560_0, i_10_394_3563_0, i_10_394_3685_0,
    i_10_394_3782_0, i_10_394_3784_0, i_10_394_3786_0, i_10_394_3787_0,
    i_10_394_3834_0, i_10_394_3855_0, i_10_394_3856_0, i_10_394_3892_0,
    i_10_394_3981_0, i_10_394_4025_0, i_10_394_4113_0, i_10_394_4213_0,
    i_10_394_4270_0, i_10_394_4279_0, i_10_394_4285_0, i_10_394_4288_0;
  output o_10_394_0_0;
  assign o_10_394_0_0 = 0;
endmodule



// Benchmark "kernel_10_395" written by ABC on Sun Jul 19 10:27:54 2020

module kernel_10_395 ( 
    i_10_395_41_0, i_10_395_42_0, i_10_395_147_0, i_10_395_175_0,
    i_10_395_179_0, i_10_395_224_0, i_10_395_251_0, i_10_395_255_0,
    i_10_395_272_0, i_10_395_282_0, i_10_395_318_0, i_10_395_327_0,
    i_10_395_328_0, i_10_395_439_0, i_10_395_444_0, i_10_395_445_0,
    i_10_395_447_0, i_10_395_516_0, i_10_395_517_0, i_10_395_717_0,
    i_10_395_755_0, i_10_395_798_0, i_10_395_956_0, i_10_395_958_0,
    i_10_395_959_0, i_10_395_961_0, i_10_395_968_0, i_10_395_984_0,
    i_10_395_1028_0, i_10_395_1033_0, i_10_395_1034_0, i_10_395_1206_0,
    i_10_395_1207_0, i_10_395_1306_0, i_10_395_1381_0, i_10_395_1438_0,
    i_10_395_1443_0, i_10_395_1575_0, i_10_395_1581_0, i_10_395_1582_0,
    i_10_395_1645_0, i_10_395_1650_0, i_10_395_1653_0, i_10_395_1654_0,
    i_10_395_1686_0, i_10_395_1713_0, i_10_395_1723_0, i_10_395_1727_0,
    i_10_395_1890_0, i_10_395_2006_0, i_10_395_2017_0, i_10_395_2018_0,
    i_10_395_2179_0, i_10_395_2196_0, i_10_395_2197_0, i_10_395_2204_0,
    i_10_395_2254_0, i_10_395_2327_0, i_10_395_2386_0, i_10_395_2450_0,
    i_10_395_2452_0, i_10_395_2459_0, i_10_395_2471_0, i_10_395_2542_0,
    i_10_395_2564_0, i_10_395_2636_0, i_10_395_2700_0, i_10_395_2702_0,
    i_10_395_2715_0, i_10_395_2721_0, i_10_395_2722_0, i_10_395_2724_0,
    i_10_395_2743_0, i_10_395_2744_0, i_10_395_2922_0, i_10_395_2980_0,
    i_10_395_3038_0, i_10_395_3071_0, i_10_395_3072_0, i_10_395_3079_0,
    i_10_395_3195_0, i_10_395_3196_0, i_10_395_3197_0, i_10_395_3313_0,
    i_10_395_3388_0, i_10_395_3391_0, i_10_395_3392_0, i_10_395_3402_0,
    i_10_395_3473_0, i_10_395_3493_0, i_10_395_3614_0, i_10_395_3646_0,
    i_10_395_3782_0, i_10_395_3798_0, i_10_395_3799_0, i_10_395_3838_0,
    i_10_395_3982_0, i_10_395_4125_0, i_10_395_4170_0, i_10_395_4531_0,
    o_10_395_0_0  );
  input  i_10_395_41_0, i_10_395_42_0, i_10_395_147_0, i_10_395_175_0,
    i_10_395_179_0, i_10_395_224_0, i_10_395_251_0, i_10_395_255_0,
    i_10_395_272_0, i_10_395_282_0, i_10_395_318_0, i_10_395_327_0,
    i_10_395_328_0, i_10_395_439_0, i_10_395_444_0, i_10_395_445_0,
    i_10_395_447_0, i_10_395_516_0, i_10_395_517_0, i_10_395_717_0,
    i_10_395_755_0, i_10_395_798_0, i_10_395_956_0, i_10_395_958_0,
    i_10_395_959_0, i_10_395_961_0, i_10_395_968_0, i_10_395_984_0,
    i_10_395_1028_0, i_10_395_1033_0, i_10_395_1034_0, i_10_395_1206_0,
    i_10_395_1207_0, i_10_395_1306_0, i_10_395_1381_0, i_10_395_1438_0,
    i_10_395_1443_0, i_10_395_1575_0, i_10_395_1581_0, i_10_395_1582_0,
    i_10_395_1645_0, i_10_395_1650_0, i_10_395_1653_0, i_10_395_1654_0,
    i_10_395_1686_0, i_10_395_1713_0, i_10_395_1723_0, i_10_395_1727_0,
    i_10_395_1890_0, i_10_395_2006_0, i_10_395_2017_0, i_10_395_2018_0,
    i_10_395_2179_0, i_10_395_2196_0, i_10_395_2197_0, i_10_395_2204_0,
    i_10_395_2254_0, i_10_395_2327_0, i_10_395_2386_0, i_10_395_2450_0,
    i_10_395_2452_0, i_10_395_2459_0, i_10_395_2471_0, i_10_395_2542_0,
    i_10_395_2564_0, i_10_395_2636_0, i_10_395_2700_0, i_10_395_2702_0,
    i_10_395_2715_0, i_10_395_2721_0, i_10_395_2722_0, i_10_395_2724_0,
    i_10_395_2743_0, i_10_395_2744_0, i_10_395_2922_0, i_10_395_2980_0,
    i_10_395_3038_0, i_10_395_3071_0, i_10_395_3072_0, i_10_395_3079_0,
    i_10_395_3195_0, i_10_395_3196_0, i_10_395_3197_0, i_10_395_3313_0,
    i_10_395_3388_0, i_10_395_3391_0, i_10_395_3392_0, i_10_395_3402_0,
    i_10_395_3473_0, i_10_395_3493_0, i_10_395_3614_0, i_10_395_3646_0,
    i_10_395_3782_0, i_10_395_3798_0, i_10_395_3799_0, i_10_395_3838_0,
    i_10_395_3982_0, i_10_395_4125_0, i_10_395_4170_0, i_10_395_4531_0;
  output o_10_395_0_0;
  assign o_10_395_0_0 = 0;
endmodule



// Benchmark "kernel_10_396" written by ABC on Sun Jul 19 10:27:55 2020

module kernel_10_396 ( 
    i_10_396_160_0, i_10_396_246_0, i_10_396_442_0, i_10_396_461_0,
    i_10_396_464_0, i_10_396_716_0, i_10_396_728_0, i_10_396_749_0,
    i_10_396_899_0, i_10_396_905_0, i_10_396_913_0, i_10_396_962_0,
    i_10_396_995_0, i_10_396_1058_0, i_10_396_1087_0, i_10_396_1129_0,
    i_10_396_1130_0, i_10_396_1220_0, i_10_396_1307_0, i_10_396_1309_0,
    i_10_396_1310_0, i_10_396_1311_0, i_10_396_1312_0, i_10_396_1391_0,
    i_10_396_1442_0, i_10_396_1454_0, i_10_396_1567_0, i_10_396_1577_0,
    i_10_396_1579_0, i_10_396_1814_0, i_10_396_1822_0, i_10_396_1823_0,
    i_10_396_1930_0, i_10_396_2182_0, i_10_396_2204_0, i_10_396_2305_0,
    i_10_396_2306_0, i_10_396_2307_0, i_10_396_2433_0, i_10_396_2449_0,
    i_10_396_2450_0, i_10_396_2451_0, i_10_396_2452_0, i_10_396_2474_0,
    i_10_396_2475_0, i_10_396_2516_0, i_10_396_2609_0, i_10_396_2705_0,
    i_10_396_2722_0, i_10_396_2787_0, i_10_396_2822_0, i_10_396_2828_0,
    i_10_396_2876_0, i_10_396_2886_0, i_10_396_2986_0, i_10_396_2987_0,
    i_10_396_3071_0, i_10_396_3094_0, i_10_396_3227_0, i_10_396_3361_0,
    i_10_396_3389_0, i_10_396_3430_0, i_10_396_3451_0, i_10_396_3452_0,
    i_10_396_3455_0, i_10_396_3589_0, i_10_396_3610_0, i_10_396_3640_0,
    i_10_396_3650_0, i_10_396_3652_0, i_10_396_3686_0, i_10_396_3703_0,
    i_10_396_3721_0, i_10_396_3725_0, i_10_396_3837_0, i_10_396_3840_0,
    i_10_396_3896_0, i_10_396_3920_0, i_10_396_3978_0, i_10_396_4057_0,
    i_10_396_4113_0, i_10_396_4117_0, i_10_396_4118_0, i_10_396_4130_0,
    i_10_396_4145_0, i_10_396_4148_0, i_10_396_4173_0, i_10_396_4174_0,
    i_10_396_4231_0, i_10_396_4238_0, i_10_396_4275_0, i_10_396_4278_0,
    i_10_396_4279_0, i_10_396_4281_0, i_10_396_4379_0, i_10_396_4397_0,
    i_10_396_4517_0, i_10_396_4531_0, i_10_396_4535_0, i_10_396_4560_0,
    o_10_396_0_0  );
  input  i_10_396_160_0, i_10_396_246_0, i_10_396_442_0, i_10_396_461_0,
    i_10_396_464_0, i_10_396_716_0, i_10_396_728_0, i_10_396_749_0,
    i_10_396_899_0, i_10_396_905_0, i_10_396_913_0, i_10_396_962_0,
    i_10_396_995_0, i_10_396_1058_0, i_10_396_1087_0, i_10_396_1129_0,
    i_10_396_1130_0, i_10_396_1220_0, i_10_396_1307_0, i_10_396_1309_0,
    i_10_396_1310_0, i_10_396_1311_0, i_10_396_1312_0, i_10_396_1391_0,
    i_10_396_1442_0, i_10_396_1454_0, i_10_396_1567_0, i_10_396_1577_0,
    i_10_396_1579_0, i_10_396_1814_0, i_10_396_1822_0, i_10_396_1823_0,
    i_10_396_1930_0, i_10_396_2182_0, i_10_396_2204_0, i_10_396_2305_0,
    i_10_396_2306_0, i_10_396_2307_0, i_10_396_2433_0, i_10_396_2449_0,
    i_10_396_2450_0, i_10_396_2451_0, i_10_396_2452_0, i_10_396_2474_0,
    i_10_396_2475_0, i_10_396_2516_0, i_10_396_2609_0, i_10_396_2705_0,
    i_10_396_2722_0, i_10_396_2787_0, i_10_396_2822_0, i_10_396_2828_0,
    i_10_396_2876_0, i_10_396_2886_0, i_10_396_2986_0, i_10_396_2987_0,
    i_10_396_3071_0, i_10_396_3094_0, i_10_396_3227_0, i_10_396_3361_0,
    i_10_396_3389_0, i_10_396_3430_0, i_10_396_3451_0, i_10_396_3452_0,
    i_10_396_3455_0, i_10_396_3589_0, i_10_396_3610_0, i_10_396_3640_0,
    i_10_396_3650_0, i_10_396_3652_0, i_10_396_3686_0, i_10_396_3703_0,
    i_10_396_3721_0, i_10_396_3725_0, i_10_396_3837_0, i_10_396_3840_0,
    i_10_396_3896_0, i_10_396_3920_0, i_10_396_3978_0, i_10_396_4057_0,
    i_10_396_4113_0, i_10_396_4117_0, i_10_396_4118_0, i_10_396_4130_0,
    i_10_396_4145_0, i_10_396_4148_0, i_10_396_4173_0, i_10_396_4174_0,
    i_10_396_4231_0, i_10_396_4238_0, i_10_396_4275_0, i_10_396_4278_0,
    i_10_396_4279_0, i_10_396_4281_0, i_10_396_4379_0, i_10_396_4397_0,
    i_10_396_4517_0, i_10_396_4531_0, i_10_396_4535_0, i_10_396_4560_0;
  output o_10_396_0_0;
  assign o_10_396_0_0 = 0;
endmodule



// Benchmark "kernel_10_397" written by ABC on Sun Jul 19 10:27:56 2020

module kernel_10_397 ( 
    i_10_397_146_0, i_10_397_224_0, i_10_397_263_0, i_10_397_273_0,
    i_10_397_274_0, i_10_397_276_0, i_10_397_279_0, i_10_397_282_0,
    i_10_397_283_0, i_10_397_320_0, i_10_397_392_0, i_10_397_428_0,
    i_10_397_431_0, i_10_397_458_0, i_10_397_460_0, i_10_397_463_0,
    i_10_397_518_0, i_10_397_689_0, i_10_397_1235_0, i_10_397_1237_0,
    i_10_397_1238_0, i_10_397_1241_0, i_10_397_1306_0, i_10_397_1311_0,
    i_10_397_1312_0, i_10_397_1432_0, i_10_397_1435_0, i_10_397_1439_0,
    i_10_397_1541_0, i_10_397_1628_0, i_10_397_1634_0, i_10_397_1643_0,
    i_10_397_1651_0, i_10_397_1652_0, i_10_397_1653_0, i_10_397_1654_0,
    i_10_397_1733_0, i_10_397_1820_0, i_10_397_1826_0, i_10_397_2000_0,
    i_10_397_2006_0, i_10_397_2027_0, i_10_397_2031_0, i_10_397_2033_0,
    i_10_397_2358_0, i_10_397_2361_0, i_10_397_2383_0, i_10_397_2384_0,
    i_10_397_2468_0, i_10_397_2471_0, i_10_397_2474_0, i_10_397_2628_0,
    i_10_397_2702_0, i_10_397_2719_0, i_10_397_2721_0, i_10_397_2723_0,
    i_10_397_2731_0, i_10_397_2782_0, i_10_397_2783_0, i_10_397_2827_0,
    i_10_397_2828_0, i_10_397_2920_0, i_10_397_3037_0, i_10_397_3043_0,
    i_10_397_3050_0, i_10_397_3069_0, i_10_397_3116_0, i_10_397_3276_0,
    i_10_397_3281_0, i_10_397_3314_0, i_10_397_3385_0, i_10_397_3387_0,
    i_10_397_3402_0, i_10_397_3467_0, i_10_397_3470_0, i_10_397_3473_0,
    i_10_397_3506_0, i_10_397_3509_0, i_10_397_3545_0, i_10_397_3583_0,
    i_10_397_3584_0, i_10_397_3587_0, i_10_397_3589_0, i_10_397_3590_0,
    i_10_397_3650_0, i_10_397_3682_0, i_10_397_3787_0, i_10_397_3788_0,
    i_10_397_3800_0, i_10_397_3808_0, i_10_397_3809_0, i_10_397_3838_0,
    i_10_397_3839_0, i_10_397_3842_0, i_10_397_3983_0, i_10_397_3988_0,
    i_10_397_4271_0, i_10_397_4286_0, i_10_397_4289_0, i_10_397_4571_0,
    o_10_397_0_0  );
  input  i_10_397_146_0, i_10_397_224_0, i_10_397_263_0, i_10_397_273_0,
    i_10_397_274_0, i_10_397_276_0, i_10_397_279_0, i_10_397_282_0,
    i_10_397_283_0, i_10_397_320_0, i_10_397_392_0, i_10_397_428_0,
    i_10_397_431_0, i_10_397_458_0, i_10_397_460_0, i_10_397_463_0,
    i_10_397_518_0, i_10_397_689_0, i_10_397_1235_0, i_10_397_1237_0,
    i_10_397_1238_0, i_10_397_1241_0, i_10_397_1306_0, i_10_397_1311_0,
    i_10_397_1312_0, i_10_397_1432_0, i_10_397_1435_0, i_10_397_1439_0,
    i_10_397_1541_0, i_10_397_1628_0, i_10_397_1634_0, i_10_397_1643_0,
    i_10_397_1651_0, i_10_397_1652_0, i_10_397_1653_0, i_10_397_1654_0,
    i_10_397_1733_0, i_10_397_1820_0, i_10_397_1826_0, i_10_397_2000_0,
    i_10_397_2006_0, i_10_397_2027_0, i_10_397_2031_0, i_10_397_2033_0,
    i_10_397_2358_0, i_10_397_2361_0, i_10_397_2383_0, i_10_397_2384_0,
    i_10_397_2468_0, i_10_397_2471_0, i_10_397_2474_0, i_10_397_2628_0,
    i_10_397_2702_0, i_10_397_2719_0, i_10_397_2721_0, i_10_397_2723_0,
    i_10_397_2731_0, i_10_397_2782_0, i_10_397_2783_0, i_10_397_2827_0,
    i_10_397_2828_0, i_10_397_2920_0, i_10_397_3037_0, i_10_397_3043_0,
    i_10_397_3050_0, i_10_397_3069_0, i_10_397_3116_0, i_10_397_3276_0,
    i_10_397_3281_0, i_10_397_3314_0, i_10_397_3385_0, i_10_397_3387_0,
    i_10_397_3402_0, i_10_397_3467_0, i_10_397_3470_0, i_10_397_3473_0,
    i_10_397_3506_0, i_10_397_3509_0, i_10_397_3545_0, i_10_397_3583_0,
    i_10_397_3584_0, i_10_397_3587_0, i_10_397_3589_0, i_10_397_3590_0,
    i_10_397_3650_0, i_10_397_3682_0, i_10_397_3787_0, i_10_397_3788_0,
    i_10_397_3800_0, i_10_397_3808_0, i_10_397_3809_0, i_10_397_3838_0,
    i_10_397_3839_0, i_10_397_3842_0, i_10_397_3983_0, i_10_397_3988_0,
    i_10_397_4271_0, i_10_397_4286_0, i_10_397_4289_0, i_10_397_4571_0;
  output o_10_397_0_0;
  assign o_10_397_0_0 = ~((~i_10_397_3314_0 & ((~i_10_397_146_0 & ~i_10_397_3276_0 & ~i_10_397_3470_0 & ((~i_10_397_1820_0 & ~i_10_397_1826_0 & i_10_397_2719_0) | (~i_10_397_392_0 & ~i_10_397_1235_0 & ~i_10_397_2006_0 & ~i_10_397_3050_0))) | (~i_10_397_392_0 & ~i_10_397_458_0 & ~i_10_397_1306_0 & ~i_10_397_1435_0 & ~i_10_397_1653_0 & ~i_10_397_1820_0 & ~i_10_397_3281_0 & ~i_10_397_3473_0 & ~i_10_397_3509_0 & i_10_397_4271_0))) | (~i_10_397_2471_0 & ((~i_10_397_1435_0 & ~i_10_397_2027_0 & ((~i_10_397_263_0 & ~i_10_397_431_0 & ~i_10_397_1628_0 & ~i_10_397_2000_0 & ~i_10_397_3470_0 & ~i_10_397_3509_0 & ~i_10_397_3545_0) | (i_10_397_2628_0 & ~i_10_397_3402_0 & ~i_10_397_3467_0 & ~i_10_397_3590_0))) | (~i_10_397_458_0 & ~i_10_397_2000_0 & ~i_10_397_2006_0 & ~i_10_397_3509_0 & ~i_10_397_3545_0 & ~i_10_397_3584_0))) | (~i_10_397_431_0 & ((~i_10_397_460_0 & ~i_10_397_2000_0 & ~i_10_397_2031_0 & ~i_10_397_2474_0 & ~i_10_397_3470_0 & ~i_10_397_3545_0 & ~i_10_397_4271_0) | (~i_10_397_282_0 & ~i_10_397_2033_0 & ~i_10_397_2383_0 & i_10_397_2471_0 & ~i_10_397_2723_0 & ~i_10_397_3050_0 & ~i_10_397_3467_0 & ~i_10_397_3842_0 & ~i_10_397_4571_0))) | (~i_10_397_458_0 & ~i_10_397_3983_0 & ((~i_10_397_2000_0 & ~i_10_397_2006_0 & ~i_10_397_2702_0 & ~i_10_397_2719_0 & ~i_10_397_3387_0 & ~i_10_397_3467_0 & ~i_10_397_3839_0 & ~i_10_397_3842_0) | (i_10_397_431_0 & ~i_10_397_3506_0 & ~i_10_397_4271_0))) | (~i_10_397_2006_0 & ((i_10_397_1312_0 & ~i_10_397_3587_0 & i_10_397_3589_0) | (~i_10_397_1235_0 & ~i_10_397_2723_0 & ~i_10_397_3043_0 & ~i_10_397_3276_0 & ~i_10_397_3281_0 & ~i_10_397_3506_0 & ~i_10_397_3839_0 & ~i_10_397_4289_0))) | (~i_10_397_3473_0 & ((~i_10_397_146_0 & ~i_10_397_2000_0 & ~i_10_397_2731_0 & ~i_10_397_3281_0 & ~i_10_397_3387_0 & ~i_10_397_3470_0 & ~i_10_397_3842_0 & ~i_10_397_4271_0) | (i_10_397_2721_0 & i_10_397_4571_0))) | (~i_10_397_3583_0 & ((~i_10_397_2468_0 & ~i_10_397_2474_0 & ~i_10_397_3587_0) | (i_10_397_2828_0 & i_10_397_4289_0))));
endmodule



// Benchmark "kernel_10_398" written by ABC on Sun Jul 19 10:27:57 2020

module kernel_10_398 ( 
    i_10_398_145_0, i_10_398_262_0, i_10_398_284_0, i_10_398_325_0,
    i_10_398_408_0, i_10_398_433_0, i_10_398_436_0, i_10_398_447_0,
    i_10_398_711_0, i_10_398_892_0, i_10_398_893_0, i_10_398_927_0,
    i_10_398_990_0, i_10_398_1036_0, i_10_398_1039_0, i_10_398_1120_0,
    i_10_398_1165_0, i_10_398_1166_0, i_10_398_1236_0, i_10_398_1238_0,
    i_10_398_1247_0, i_10_398_1307_0, i_10_398_1381_0, i_10_398_1440_0,
    i_10_398_1485_0, i_10_398_1554_0, i_10_398_1603_0, i_10_398_1800_0,
    i_10_398_1801_0, i_10_398_1824_0, i_10_398_1825_0, i_10_398_1826_0,
    i_10_398_1908_0, i_10_398_1909_0, i_10_398_1911_0, i_10_398_1981_0,
    i_10_398_1990_0, i_10_398_2206_0, i_10_398_2223_0, i_10_398_2224_0,
    i_10_398_2332_0, i_10_398_2449_0, i_10_398_2450_0, i_10_398_2458_0,
    i_10_398_2481_0, i_10_398_2515_0, i_10_398_2565_0, i_10_398_2567_0,
    i_10_398_2571_0, i_10_398_2635_0, i_10_398_2686_0, i_10_398_2700_0,
    i_10_398_2701_0, i_10_398_2728_0, i_10_398_2827_0, i_10_398_2829_0,
    i_10_398_2831_0, i_10_398_2862_0, i_10_398_2865_0, i_10_398_2866_0,
    i_10_398_2916_0, i_10_398_2917_0, i_10_398_2919_0, i_10_398_2920_0,
    i_10_398_2921_0, i_10_398_2922_0, i_10_398_2923_0, i_10_398_3072_0,
    i_10_398_3199_0, i_10_398_3201_0, i_10_398_3267_0, i_10_398_3278_0,
    i_10_398_3298_0, i_10_398_3299_0, i_10_398_3384_0, i_10_398_3385_0,
    i_10_398_3386_0, i_10_398_3388_0, i_10_398_3406_0, i_10_398_3457_0,
    i_10_398_3523_0, i_10_398_3600_0, i_10_398_3610_0, i_10_398_3611_0,
    i_10_398_3648_0, i_10_398_3851_0, i_10_398_3855_0, i_10_398_3889_0,
    i_10_398_3897_0, i_10_398_3942_0, i_10_398_3943_0, i_10_398_3961_0,
    i_10_398_4120_0, i_10_398_4129_0, i_10_398_4269_0, i_10_398_4270_0,
    i_10_398_4285_0, i_10_398_4306_0, i_10_398_4500_0, i_10_398_4597_0,
    o_10_398_0_0  );
  input  i_10_398_145_0, i_10_398_262_0, i_10_398_284_0, i_10_398_325_0,
    i_10_398_408_0, i_10_398_433_0, i_10_398_436_0, i_10_398_447_0,
    i_10_398_711_0, i_10_398_892_0, i_10_398_893_0, i_10_398_927_0,
    i_10_398_990_0, i_10_398_1036_0, i_10_398_1039_0, i_10_398_1120_0,
    i_10_398_1165_0, i_10_398_1166_0, i_10_398_1236_0, i_10_398_1238_0,
    i_10_398_1247_0, i_10_398_1307_0, i_10_398_1381_0, i_10_398_1440_0,
    i_10_398_1485_0, i_10_398_1554_0, i_10_398_1603_0, i_10_398_1800_0,
    i_10_398_1801_0, i_10_398_1824_0, i_10_398_1825_0, i_10_398_1826_0,
    i_10_398_1908_0, i_10_398_1909_0, i_10_398_1911_0, i_10_398_1981_0,
    i_10_398_1990_0, i_10_398_2206_0, i_10_398_2223_0, i_10_398_2224_0,
    i_10_398_2332_0, i_10_398_2449_0, i_10_398_2450_0, i_10_398_2458_0,
    i_10_398_2481_0, i_10_398_2515_0, i_10_398_2565_0, i_10_398_2567_0,
    i_10_398_2571_0, i_10_398_2635_0, i_10_398_2686_0, i_10_398_2700_0,
    i_10_398_2701_0, i_10_398_2728_0, i_10_398_2827_0, i_10_398_2829_0,
    i_10_398_2831_0, i_10_398_2862_0, i_10_398_2865_0, i_10_398_2866_0,
    i_10_398_2916_0, i_10_398_2917_0, i_10_398_2919_0, i_10_398_2920_0,
    i_10_398_2921_0, i_10_398_2922_0, i_10_398_2923_0, i_10_398_3072_0,
    i_10_398_3199_0, i_10_398_3201_0, i_10_398_3267_0, i_10_398_3278_0,
    i_10_398_3298_0, i_10_398_3299_0, i_10_398_3384_0, i_10_398_3385_0,
    i_10_398_3386_0, i_10_398_3388_0, i_10_398_3406_0, i_10_398_3457_0,
    i_10_398_3523_0, i_10_398_3600_0, i_10_398_3610_0, i_10_398_3611_0,
    i_10_398_3648_0, i_10_398_3851_0, i_10_398_3855_0, i_10_398_3889_0,
    i_10_398_3897_0, i_10_398_3942_0, i_10_398_3943_0, i_10_398_3961_0,
    i_10_398_4120_0, i_10_398_4129_0, i_10_398_4269_0, i_10_398_4270_0,
    i_10_398_4285_0, i_10_398_4306_0, i_10_398_4500_0, i_10_398_4597_0;
  output o_10_398_0_0;
  assign o_10_398_0_0 = 0;
endmodule



// Benchmark "kernel_10_399" written by ABC on Sun Jul 19 10:27:58 2020

module kernel_10_399 ( 
    i_10_399_29_0, i_10_399_41_0, i_10_399_50_0, i_10_399_146_0,
    i_10_399_173_0, i_10_399_174_0, i_10_399_224_0, i_10_399_250_0,
    i_10_399_316_0, i_10_399_319_0, i_10_399_406_0, i_10_399_430_0,
    i_10_399_431_0, i_10_399_508_0, i_10_399_509_0, i_10_399_518_0,
    i_10_399_589_0, i_10_399_590_0, i_10_399_751_0, i_10_399_792_0,
    i_10_399_796_0, i_10_399_800_0, i_10_399_908_0, i_10_399_964_0,
    i_10_399_1032_0, i_10_399_1138_0, i_10_399_1306_0, i_10_399_1448_0,
    i_10_399_1545_0, i_10_399_1643_0, i_10_399_1690_0, i_10_399_1769_0,
    i_10_399_1811_0, i_10_399_1913_0, i_10_399_1937_0, i_10_399_1949_0,
    i_10_399_1999_0, i_10_399_2003_0, i_10_399_2312_0, i_10_399_2350_0,
    i_10_399_2354_0, i_10_399_2365_0, i_10_399_2389_0, i_10_399_2450_0,
    i_10_399_2451_0, i_10_399_2452_0, i_10_399_2453_0, i_10_399_2455_0,
    i_10_399_2469_0, i_10_399_2471_0, i_10_399_2546_0, i_10_399_2628_0,
    i_10_399_2629_0, i_10_399_2661_0, i_10_399_2663_0, i_10_399_2705_0,
    i_10_399_2717_0, i_10_399_2722_0, i_10_399_2723_0, i_10_399_2731_0,
    i_10_399_2732_0, i_10_399_2781_0, i_10_399_2785_0, i_10_399_2821_0,
    i_10_399_2822_0, i_10_399_2824_0, i_10_399_2827_0, i_10_399_2828_0,
    i_10_399_3035_0, i_10_399_3157_0, i_10_399_3236_0, i_10_399_3271_0,
    i_10_399_3280_0, i_10_399_3281_0, i_10_399_3284_0, i_10_399_3322_0,
    i_10_399_3410_0, i_10_399_3466_0, i_10_399_3494_0, i_10_399_3497_0,
    i_10_399_3520_0, i_10_399_3526_0, i_10_399_3584_0, i_10_399_3587_0,
    i_10_399_3613_0, i_10_399_3617_0, i_10_399_3649_0, i_10_399_3788_0,
    i_10_399_3800_0, i_10_399_3838_0, i_10_399_3846_0, i_10_399_3875_0,
    i_10_399_3911_0, i_10_399_3914_0, i_10_399_4123_0, i_10_399_4172_0,
    i_10_399_4268_0, i_10_399_4277_0, i_10_399_4291_0, i_10_399_4292_0,
    o_10_399_0_0  );
  input  i_10_399_29_0, i_10_399_41_0, i_10_399_50_0, i_10_399_146_0,
    i_10_399_173_0, i_10_399_174_0, i_10_399_224_0, i_10_399_250_0,
    i_10_399_316_0, i_10_399_319_0, i_10_399_406_0, i_10_399_430_0,
    i_10_399_431_0, i_10_399_508_0, i_10_399_509_0, i_10_399_518_0,
    i_10_399_589_0, i_10_399_590_0, i_10_399_751_0, i_10_399_792_0,
    i_10_399_796_0, i_10_399_800_0, i_10_399_908_0, i_10_399_964_0,
    i_10_399_1032_0, i_10_399_1138_0, i_10_399_1306_0, i_10_399_1448_0,
    i_10_399_1545_0, i_10_399_1643_0, i_10_399_1690_0, i_10_399_1769_0,
    i_10_399_1811_0, i_10_399_1913_0, i_10_399_1937_0, i_10_399_1949_0,
    i_10_399_1999_0, i_10_399_2003_0, i_10_399_2312_0, i_10_399_2350_0,
    i_10_399_2354_0, i_10_399_2365_0, i_10_399_2389_0, i_10_399_2450_0,
    i_10_399_2451_0, i_10_399_2452_0, i_10_399_2453_0, i_10_399_2455_0,
    i_10_399_2469_0, i_10_399_2471_0, i_10_399_2546_0, i_10_399_2628_0,
    i_10_399_2629_0, i_10_399_2661_0, i_10_399_2663_0, i_10_399_2705_0,
    i_10_399_2717_0, i_10_399_2722_0, i_10_399_2723_0, i_10_399_2731_0,
    i_10_399_2732_0, i_10_399_2781_0, i_10_399_2785_0, i_10_399_2821_0,
    i_10_399_2822_0, i_10_399_2824_0, i_10_399_2827_0, i_10_399_2828_0,
    i_10_399_3035_0, i_10_399_3157_0, i_10_399_3236_0, i_10_399_3271_0,
    i_10_399_3280_0, i_10_399_3281_0, i_10_399_3284_0, i_10_399_3322_0,
    i_10_399_3410_0, i_10_399_3466_0, i_10_399_3494_0, i_10_399_3497_0,
    i_10_399_3520_0, i_10_399_3526_0, i_10_399_3584_0, i_10_399_3587_0,
    i_10_399_3613_0, i_10_399_3617_0, i_10_399_3649_0, i_10_399_3788_0,
    i_10_399_3800_0, i_10_399_3838_0, i_10_399_3846_0, i_10_399_3875_0,
    i_10_399_3911_0, i_10_399_3914_0, i_10_399_4123_0, i_10_399_4172_0,
    i_10_399_4268_0, i_10_399_4277_0, i_10_399_4291_0, i_10_399_4292_0;
  output o_10_399_0_0;
  assign o_10_399_0_0 = ~((i_10_399_174_0 & ((~i_10_399_250_0 & ~i_10_399_1545_0 & ~i_10_399_2781_0 & ~i_10_399_3526_0 & ~i_10_399_3587_0 & ~i_10_399_3649_0) | (~i_10_399_1769_0 & ~i_10_399_2471_0 & ~i_10_399_2785_0 & ~i_10_399_2821_0 & ~i_10_399_3410_0 & ~i_10_399_3617_0 & ~i_10_399_3846_0))) | (~i_10_399_431_0 & ((~i_10_399_224_0 & ((~i_10_399_146_0 & ~i_10_399_319_0 & ~i_10_399_908_0 & ~i_10_399_3271_0 & ~i_10_399_3284_0 & ~i_10_399_3466_0 & ~i_10_399_3526_0 & ~i_10_399_3838_0) | (~i_10_399_518_0 & ~i_10_399_2453_0 & ~i_10_399_2785_0 & ~i_10_399_3911_0 & ~i_10_399_3914_0))) | (~i_10_399_2312_0 & ((~i_10_399_2003_0 & ~i_10_399_2350_0 & ~i_10_399_2451_0 & ~i_10_399_2452_0 & ~i_10_399_2453_0 & ~i_10_399_3280_0 & ~i_10_399_3526_0) | (~i_10_399_316_0 & i_10_399_2781_0 & ~i_10_399_2822_0 & ~i_10_399_4172_0))))) | (~i_10_399_316_0 & ((~i_10_399_796_0 & i_10_399_2450_0 & ~i_10_399_2717_0 & ~i_10_399_2723_0 & i_10_399_2827_0) | (~i_10_399_908_0 & ~i_10_399_1032_0 & i_10_399_2661_0 & ~i_10_399_2722_0 & ~i_10_399_2822_0 & ~i_10_399_3497_0 & ~i_10_399_4172_0 & ~i_10_399_4268_0))) | (~i_10_399_3914_0 & ((~i_10_399_173_0 & ((~i_10_399_319_0 & ~i_10_399_792_0 & ~i_10_399_1032_0 & ~i_10_399_2723_0 & ~i_10_399_2732_0 & ~i_10_399_3584_0 & i_10_399_3838_0) | (~i_10_399_908_0 & ~i_10_399_964_0 & ~i_10_399_2312_0 & ~i_10_399_2471_0 & ~i_10_399_2717_0 & ~i_10_399_3410_0 & ~i_10_399_4172_0))) | (~i_10_399_908_0 & ((i_10_399_319_0 & ~i_10_399_796_0 & ~i_10_399_1690_0 & ~i_10_399_1913_0 & ~i_10_399_1949_0 & ~i_10_399_1999_0 & ~i_10_399_2312_0 & ~i_10_399_2450_0 & ~i_10_399_2451_0 & ~i_10_399_2781_0) | (~i_10_399_146_0 & ~i_10_399_2452_0 & ~i_10_399_2471_0 & ~i_10_399_2663_0 & ~i_10_399_2732_0 & ~i_10_399_2822_0))) | (~i_10_399_146_0 & ((i_10_399_751_0 & ~i_10_399_1448_0 & ~i_10_399_2003_0 & ~i_10_399_2785_0 & ~i_10_399_2827_0) | (~i_10_399_800_0 & ~i_10_399_1545_0 & ~i_10_399_2312_0 & ~i_10_399_2453_0 & i_10_399_2661_0 & ~i_10_399_4268_0))) | (~i_10_399_1769_0 & ~i_10_399_2471_0 & ((~i_10_399_319_0 & ~i_10_399_2450_0 & ~i_10_399_2663_0 & ~i_10_399_3281_0 & ~i_10_399_3587_0 & ~i_10_399_3649_0) | (~i_10_399_1545_0 & ~i_10_399_2821_0 & ~i_10_399_3410_0 & ~i_10_399_3584_0 & ~i_10_399_4291_0 & ~i_10_399_4292_0))))) | (~i_10_399_1690_0 & ((~i_10_399_146_0 & ~i_10_399_406_0 & ~i_10_399_908_0 & ~i_10_399_2312_0 & ~i_10_399_2452_0 & ~i_10_399_2731_0 & ~i_10_399_3284_0) | (~i_10_399_173_0 & i_10_399_1306_0 & ~i_10_399_2003_0 & ~i_10_399_3281_0 & ~i_10_399_3410_0 & ~i_10_399_3466_0 & ~i_10_399_3526_0))) | (~i_10_399_146_0 & ((i_10_399_796_0 & ~i_10_399_2312_0 & ~i_10_399_2354_0 & i_10_399_2451_0 & ~i_10_399_2705_0 & ~i_10_399_2731_0 & ~i_10_399_2824_0 & ~i_10_399_3466_0 & ~i_10_399_3526_0) | (~i_10_399_518_0 & ~i_10_399_3281_0 & i_10_399_3520_0 & i_10_399_3838_0))) | (~i_10_399_2452_0 & ((~i_10_399_406_0 & ~i_10_399_3281_0 & ((~i_10_399_908_0 & ~i_10_399_2717_0 & ~i_10_399_2822_0 & ~i_10_399_3584_0) | (~i_10_399_1769_0 & ~i_10_399_2003_0 & ~i_10_399_2471_0 & ~i_10_399_3497_0 & ~i_10_399_3613_0))) | (i_10_399_29_0 & i_10_399_1949_0 & ~i_10_399_2663_0))) | (~i_10_399_518_0 & ~i_10_399_3911_0 & ((~i_10_399_800_0 & ~i_10_399_1913_0 & ~i_10_399_2450_0 & ~i_10_399_2705_0 & ~i_10_399_2785_0 & ~i_10_399_3284_0) | (i_10_399_1690_0 & ~i_10_399_1999_0 & ~i_10_399_2453_0 & ~i_10_399_2661_0 & ~i_10_399_2723_0 & ~i_10_399_4268_0))) | (~i_10_399_3587_0 & ((~i_10_399_751_0 & ~i_10_399_908_0 & i_10_399_2661_0 & ~i_10_399_3284_0) | i_10_399_3788_0 | (~i_10_399_2663_0 & ~i_10_399_2717_0 & ~i_10_399_2824_0 & ~i_10_399_4292_0))) | (i_10_399_792_0 & ~i_10_399_2453_0 & ~i_10_399_2455_0 & ~i_10_399_3584_0));
endmodule



// Benchmark "kernel_10_400" written by ABC on Sun Jul 19 10:27:59 2020

module kernel_10_400 ( 
    i_10_400_150_0, i_10_400_174_0, i_10_400_175_0, i_10_400_176_0,
    i_10_400_177_0, i_10_400_178_0, i_10_400_179_0, i_10_400_250_0,
    i_10_400_251_0, i_10_400_281_0, i_10_400_282_0, i_10_400_285_0,
    i_10_400_287_0, i_10_400_289_0, i_10_400_318_0, i_10_400_321_0,
    i_10_400_322_0, i_10_400_407_0, i_10_400_408_0, i_10_400_412_0,
    i_10_400_428_0, i_10_400_437_0, i_10_400_439_0, i_10_400_455_0,
    i_10_400_717_0, i_10_400_1002_0, i_10_400_1003_0, i_10_400_1138_0,
    i_10_400_1142_0, i_10_400_1236_0, i_10_400_1237_0, i_10_400_1312_0,
    i_10_400_1344_0, i_10_400_1365_0, i_10_400_1384_0, i_10_400_1441_0,
    i_10_400_1651_0, i_10_400_1684_0, i_10_400_1688_0, i_10_400_1689_0,
    i_10_400_1690_0, i_10_400_1821_0, i_10_400_1823_0, i_10_400_1990_0,
    i_10_400_2022_0, i_10_400_2028_0, i_10_400_2311_0, i_10_400_2349_0,
    i_10_400_2353_0, i_10_400_2410_0, i_10_400_2411_0, i_10_400_2453_0,
    i_10_400_2454_0, i_10_400_2629_0, i_10_400_2632_0, i_10_400_2633_0,
    i_10_400_2635_0, i_10_400_2636_0, i_10_400_2655_0, i_10_400_2660_0,
    i_10_400_2661_0, i_10_400_2704_0, i_10_400_2714_0, i_10_400_2727_0,
    i_10_400_2733_0, i_10_400_2734_0, i_10_400_2735_0, i_10_400_2781_0,
    i_10_400_2785_0, i_10_400_2826_0, i_10_400_2834_0, i_10_400_3039_0,
    i_10_400_3042_0, i_10_400_3075_0, i_10_400_3157_0, i_10_400_3202_0,
    i_10_400_3390_0, i_10_400_3405_0, i_10_400_3468_0, i_10_400_3469_0,
    i_10_400_3496_0, i_10_400_3615_0, i_10_400_3648_0, i_10_400_3651_0,
    i_10_400_3839_0, i_10_400_3846_0, i_10_400_3857_0, i_10_400_3858_0,
    i_10_400_3860_0, i_10_400_3912_0, i_10_400_3984_0, i_10_400_4116_0,
    i_10_400_4117_0, i_10_400_4119_0, i_10_400_4120_0, i_10_400_4122_0,
    i_10_400_4123_0, i_10_400_4125_0, i_10_400_4126_0, i_10_400_4270_0,
    o_10_400_0_0  );
  input  i_10_400_150_0, i_10_400_174_0, i_10_400_175_0, i_10_400_176_0,
    i_10_400_177_0, i_10_400_178_0, i_10_400_179_0, i_10_400_250_0,
    i_10_400_251_0, i_10_400_281_0, i_10_400_282_0, i_10_400_285_0,
    i_10_400_287_0, i_10_400_289_0, i_10_400_318_0, i_10_400_321_0,
    i_10_400_322_0, i_10_400_407_0, i_10_400_408_0, i_10_400_412_0,
    i_10_400_428_0, i_10_400_437_0, i_10_400_439_0, i_10_400_455_0,
    i_10_400_717_0, i_10_400_1002_0, i_10_400_1003_0, i_10_400_1138_0,
    i_10_400_1142_0, i_10_400_1236_0, i_10_400_1237_0, i_10_400_1312_0,
    i_10_400_1344_0, i_10_400_1365_0, i_10_400_1384_0, i_10_400_1441_0,
    i_10_400_1651_0, i_10_400_1684_0, i_10_400_1688_0, i_10_400_1689_0,
    i_10_400_1690_0, i_10_400_1821_0, i_10_400_1823_0, i_10_400_1990_0,
    i_10_400_2022_0, i_10_400_2028_0, i_10_400_2311_0, i_10_400_2349_0,
    i_10_400_2353_0, i_10_400_2410_0, i_10_400_2411_0, i_10_400_2453_0,
    i_10_400_2454_0, i_10_400_2629_0, i_10_400_2632_0, i_10_400_2633_0,
    i_10_400_2635_0, i_10_400_2636_0, i_10_400_2655_0, i_10_400_2660_0,
    i_10_400_2661_0, i_10_400_2704_0, i_10_400_2714_0, i_10_400_2727_0,
    i_10_400_2733_0, i_10_400_2734_0, i_10_400_2735_0, i_10_400_2781_0,
    i_10_400_2785_0, i_10_400_2826_0, i_10_400_2834_0, i_10_400_3039_0,
    i_10_400_3042_0, i_10_400_3075_0, i_10_400_3157_0, i_10_400_3202_0,
    i_10_400_3390_0, i_10_400_3405_0, i_10_400_3468_0, i_10_400_3469_0,
    i_10_400_3496_0, i_10_400_3615_0, i_10_400_3648_0, i_10_400_3651_0,
    i_10_400_3839_0, i_10_400_3846_0, i_10_400_3857_0, i_10_400_3858_0,
    i_10_400_3860_0, i_10_400_3912_0, i_10_400_3984_0, i_10_400_4116_0,
    i_10_400_4117_0, i_10_400_4119_0, i_10_400_4120_0, i_10_400_4122_0,
    i_10_400_4123_0, i_10_400_4125_0, i_10_400_4126_0, i_10_400_4270_0;
  output o_10_400_0_0;
  assign o_10_400_0_0 = ~((~i_10_400_408_0 & ((~i_10_400_178_0 & ((~i_10_400_179_0 & ~i_10_400_3075_0 & ((~i_10_400_174_0 & ~i_10_400_289_0 & ~i_10_400_1237_0 & ~i_10_400_2349_0 & ~i_10_400_2826_0 & ~i_10_400_3468_0 & ~i_10_400_3648_0 & ~i_10_400_3984_0) | (~i_10_400_251_0 & ~i_10_400_2453_0 & i_10_400_3039_0 & ~i_10_400_3846_0 & ~i_10_400_4123_0))) | (~i_10_400_318_0 & ~i_10_400_1236_0 & ~i_10_400_2735_0 & i_10_400_3202_0 & i_10_400_3651_0))) | (~i_10_400_3912_0 & ~i_10_400_4123_0 & ((~i_10_400_250_0 & ((~i_10_400_318_0 & ~i_10_400_322_0 & ~i_10_400_1990_0 & ~i_10_400_2028_0 & ~i_10_400_2636_0 & ~i_10_400_3042_0 & ~i_10_400_3390_0 & ~i_10_400_3496_0) | (~i_10_400_177_0 & ~i_10_400_407_0 & ~i_10_400_1651_0 & ~i_10_400_1689_0 & ~i_10_400_3468_0 & ~i_10_400_4122_0 & ~i_10_400_4126_0))) | (~i_10_400_282_0 & ~i_10_400_407_0 & ~i_10_400_1441_0 & ~i_10_400_2022_0 & ~i_10_400_2734_0 & ~i_10_400_3468_0 & ~i_10_400_3857_0 & ~i_10_400_4122_0))))) | (~i_10_400_321_0 & ((~i_10_400_178_0 & ((~i_10_400_455_0 & i_10_400_1651_0 & ~i_10_400_1684_0 & ~i_10_400_4116_0 & ~i_10_400_4119_0) | (~i_10_400_150_0 & ~i_10_400_2022_0 & ~i_10_400_2633_0 & ~i_10_400_2704_0 & ~i_10_400_3042_0 & ~i_10_400_3468_0 & ~i_10_400_4123_0 & ~i_10_400_4270_0))) | (~i_10_400_1365_0 & ((~i_10_400_281_0 & ~i_10_400_322_0 & ~i_10_400_717_0 & ~i_10_400_1689_0 & ~i_10_400_2704_0 & ~i_10_400_3042_0 & ~i_10_400_3496_0 & ~i_10_400_4122_0) | (~i_10_400_289_0 & ~i_10_400_437_0 & i_10_400_1237_0 & ~i_10_400_1688_0 & ~i_10_400_1690_0 & ~i_10_400_2454_0 & ~i_10_400_2714_0 & ~i_10_400_3075_0 & ~i_10_400_3468_0 & ~i_10_400_4125_0))) | (~i_10_400_2349_0 & ~i_10_400_3468_0 & ((~i_10_400_177_0 & ~i_10_400_251_0 & ~i_10_400_2733_0 & ~i_10_400_3469_0 & ~i_10_400_3846_0 & ~i_10_400_4116_0) | (~i_10_400_175_0 & ~i_10_400_2661_0 & ~i_10_400_3075_0 & ~i_10_400_3648_0 & ~i_10_400_4122_0))) | (~i_10_400_174_0 & ~i_10_400_287_0 & ~i_10_400_1821_0 & ~i_10_400_2660_0 & ~i_10_400_3042_0 & ~i_10_400_3075_0 & ~i_10_400_3469_0 & ~i_10_400_3839_0 & ~i_10_400_4123_0 & ~i_10_400_4126_0))) | (~i_10_400_281_0 & ((~i_10_400_1441_0 & ~i_10_400_1684_0 & ~i_10_400_1821_0 & ~i_10_400_2022_0 & ~i_10_400_2453_0 & i_10_400_2834_0) | (~i_10_400_177_0 & ~i_10_400_285_0 & ~i_10_400_289_0 & i_10_400_2660_0 & ~i_10_400_2714_0 & ~i_10_400_3648_0 & ~i_10_400_4116_0))) | (~i_10_400_177_0 & ((~i_10_400_174_0 & ~i_10_400_175_0 & i_10_400_2636_0 & ~i_10_400_2733_0 & ~i_10_400_2781_0 & ~i_10_400_3468_0) | (~i_10_400_250_0 & ~i_10_400_3042_0 & i_10_400_3860_0))) | (~i_10_400_174_0 & ~i_10_400_3846_0 & ((i_10_400_176_0 & i_10_400_281_0 & ~i_10_400_2785_0 & ~i_10_400_3390_0) | (~i_10_400_250_0 & ~i_10_400_2022_0 & ~i_10_400_2453_0 & ~i_10_400_2704_0 & ~i_10_400_2727_0 & ~i_10_400_2733_0 & ~i_10_400_3912_0))) | (~i_10_400_175_0 & ((i_10_400_2453_0 & ~i_10_400_3839_0) | (~i_10_400_2311_0 & ~i_10_400_2353_0 & ~i_10_400_2785_0 & i_10_400_3858_0 & ~i_10_400_4122_0 & ~i_10_400_4270_0))) | (i_10_400_281_0 & ((~i_10_400_250_0 & ~i_10_400_289_0 & ~i_10_400_1441_0 & ~i_10_400_1823_0 & ~i_10_400_2349_0 & ~i_10_400_2353_0 & ~i_10_400_3469_0) | (~i_10_400_322_0 & ~i_10_400_407_0 & ~i_10_400_1237_0 & ~i_10_400_2781_0 & ~i_10_400_4116_0 & ~i_10_400_4119_0))) | (~i_10_400_1823_0 & ((~i_10_400_318_0 & i_10_400_3468_0 & ~i_10_400_3469_0 & i_10_400_3648_0 & ~i_10_400_3651_0) | (i_10_400_2635_0 & i_10_400_3615_0 & ~i_10_400_4116_0))) | (~i_10_400_318_0 & ((i_10_400_1003_0 & ~i_10_400_2735_0 & ~i_10_400_3039_0) | (~i_10_400_176_0 & ~i_10_400_717_0 & ~i_10_400_1236_0 & ~i_10_400_2714_0 & ~i_10_400_3042_0 & ~i_10_400_4120_0 & ~i_10_400_4125_0))) | (i_10_400_2629_0 & ((~i_10_400_1237_0 & ~i_10_400_1990_0 & ~i_10_400_4116_0 & ~i_10_400_4120_0 & i_10_400_4123_0) | (i_10_400_2353_0 & ~i_10_400_2661_0 & i_10_400_4117_0 & i_10_400_4125_0))) | (~i_10_400_4119_0 & ((~i_10_400_2781_0 & i_10_400_3615_0 & ~i_10_400_3912_0 & i_10_400_4125_0) | (i_10_400_455_0 & i_10_400_4120_0 & ~i_10_400_4126_0))) | (i_10_400_2633_0 & ~i_10_400_2734_0) | (~i_10_400_2349_0 & i_10_400_2727_0 & ~i_10_400_3839_0 & i_10_400_3858_0 & ~i_10_400_4120_0 & i_10_400_4122_0));
endmodule



// Benchmark "kernel_10_401" written by ABC on Sun Jul 19 10:28:01 2020

module kernel_10_401 ( 
    i_10_401_34_0, i_10_401_124_0, i_10_401_177_0, i_10_401_246_0,
    i_10_401_249_0, i_10_401_269_0, i_10_401_282_0, i_10_401_283_0,
    i_10_401_318_0, i_10_401_328_0, i_10_401_329_0, i_10_401_437_0,
    i_10_401_445_0, i_10_401_512_0, i_10_401_962_0, i_10_401_1006_0,
    i_10_401_1135_0, i_10_401_1137_0, i_10_401_1138_0, i_10_401_1241_0,
    i_10_401_1266_0, i_10_401_1348_0, i_10_401_1366_0, i_10_401_1583_0,
    i_10_401_1617_0, i_10_401_1680_0, i_10_401_1687_0, i_10_401_1819_0,
    i_10_401_1821_0, i_10_401_1825_0, i_10_401_1876_0, i_10_401_1912_0,
    i_10_401_1913_0, i_10_401_1951_0, i_10_401_1952_0, i_10_401_2084_0,
    i_10_401_2184_0, i_10_401_2185_0, i_10_401_2186_0, i_10_401_2203_0,
    i_10_401_2312_0, i_10_401_2327_0, i_10_401_2329_0, i_10_401_2338_0,
    i_10_401_2353_0, i_10_401_2354_0, i_10_401_2384_0, i_10_401_2407_0,
    i_10_401_2408_0, i_10_401_2410_0, i_10_401_2411_0, i_10_401_2452_0,
    i_10_401_2453_0, i_10_401_2470_0, i_10_401_2632_0, i_10_401_2655_0,
    i_10_401_2659_0, i_10_401_2660_0, i_10_401_2708_0, i_10_401_2726_0,
    i_10_401_2731_0, i_10_401_2829_0, i_10_401_2884_0, i_10_401_2885_0,
    i_10_401_2921_0, i_10_401_2980_0, i_10_401_2981_0, i_10_401_2986_0,
    i_10_401_3069_0, i_10_401_3274_0, i_10_401_3327_0, i_10_401_3328_0,
    i_10_401_3384_0, i_10_401_3497_0, i_10_401_3590_0, i_10_401_3616_0,
    i_10_401_3787_0, i_10_401_3847_0, i_10_401_3848_0, i_10_401_3853_0,
    i_10_401_3855_0, i_10_401_3859_0, i_10_401_3895_0, i_10_401_3920_0,
    i_10_401_3993_0, i_10_401_4056_0, i_10_401_4057_0, i_10_401_4058_0,
    i_10_401_4116_0, i_10_401_4117_0, i_10_401_4118_0, i_10_401_4124_0,
    i_10_401_4126_0, i_10_401_4127_0, i_10_401_4237_0, i_10_401_4238_0,
    i_10_401_4289_0, i_10_401_4290_0, i_10_401_4568_0, i_10_401_4570_0,
    o_10_401_0_0  );
  input  i_10_401_34_0, i_10_401_124_0, i_10_401_177_0, i_10_401_246_0,
    i_10_401_249_0, i_10_401_269_0, i_10_401_282_0, i_10_401_283_0,
    i_10_401_318_0, i_10_401_328_0, i_10_401_329_0, i_10_401_437_0,
    i_10_401_445_0, i_10_401_512_0, i_10_401_962_0, i_10_401_1006_0,
    i_10_401_1135_0, i_10_401_1137_0, i_10_401_1138_0, i_10_401_1241_0,
    i_10_401_1266_0, i_10_401_1348_0, i_10_401_1366_0, i_10_401_1583_0,
    i_10_401_1617_0, i_10_401_1680_0, i_10_401_1687_0, i_10_401_1819_0,
    i_10_401_1821_0, i_10_401_1825_0, i_10_401_1876_0, i_10_401_1912_0,
    i_10_401_1913_0, i_10_401_1951_0, i_10_401_1952_0, i_10_401_2084_0,
    i_10_401_2184_0, i_10_401_2185_0, i_10_401_2186_0, i_10_401_2203_0,
    i_10_401_2312_0, i_10_401_2327_0, i_10_401_2329_0, i_10_401_2338_0,
    i_10_401_2353_0, i_10_401_2354_0, i_10_401_2384_0, i_10_401_2407_0,
    i_10_401_2408_0, i_10_401_2410_0, i_10_401_2411_0, i_10_401_2452_0,
    i_10_401_2453_0, i_10_401_2470_0, i_10_401_2632_0, i_10_401_2655_0,
    i_10_401_2659_0, i_10_401_2660_0, i_10_401_2708_0, i_10_401_2726_0,
    i_10_401_2731_0, i_10_401_2829_0, i_10_401_2884_0, i_10_401_2885_0,
    i_10_401_2921_0, i_10_401_2980_0, i_10_401_2981_0, i_10_401_2986_0,
    i_10_401_3069_0, i_10_401_3274_0, i_10_401_3327_0, i_10_401_3328_0,
    i_10_401_3384_0, i_10_401_3497_0, i_10_401_3590_0, i_10_401_3616_0,
    i_10_401_3787_0, i_10_401_3847_0, i_10_401_3848_0, i_10_401_3853_0,
    i_10_401_3855_0, i_10_401_3859_0, i_10_401_3895_0, i_10_401_3920_0,
    i_10_401_3993_0, i_10_401_4056_0, i_10_401_4057_0, i_10_401_4058_0,
    i_10_401_4116_0, i_10_401_4117_0, i_10_401_4118_0, i_10_401_4124_0,
    i_10_401_4126_0, i_10_401_4127_0, i_10_401_4237_0, i_10_401_4238_0,
    i_10_401_4289_0, i_10_401_4290_0, i_10_401_4568_0, i_10_401_4570_0;
  output o_10_401_0_0;
  assign o_10_401_0_0 = ~((~i_10_401_2408_0 & ((~i_10_401_4237_0 & ((~i_10_401_34_0 & ((~i_10_401_177_0 & ~i_10_401_445_0 & ~i_10_401_1825_0 & ~i_10_401_2354_0 & ~i_10_401_2981_0) | (~i_10_401_328_0 & ~i_10_401_1952_0 & ~i_10_401_2410_0 & ~i_10_401_2980_0 & ~i_10_401_4056_0 & ~i_10_401_4058_0 & ~i_10_401_4116_0))) | (~i_10_401_1366_0 & ~i_10_401_1951_0 & ~i_10_401_2185_0 & ~i_10_401_2312_0 & ~i_10_401_2327_0 & ~i_10_401_2384_0 & ~i_10_401_2407_0 & ~i_10_401_2655_0 & ~i_10_401_4057_0 & ~i_10_401_4238_0))) | (~i_10_401_2407_0 & ((~i_10_401_2184_0 & ~i_10_401_2329_0 & ((~i_10_401_124_0 & ~i_10_401_2327_0 & ~i_10_401_2354_0 & ~i_10_401_2655_0 & ~i_10_401_2981_0 & ~i_10_401_3274_0 & ~i_10_401_4057_0) | (~i_10_401_962_0 & ~i_10_401_1913_0 & ~i_10_401_2312_0 & ~i_10_401_2980_0 & i_10_401_4568_0))) | (~i_10_401_2185_0 & ~i_10_401_2410_0 & ~i_10_401_2708_0 & ~i_10_401_2980_0 & ~i_10_401_4057_0 & ~i_10_401_4568_0))) | (~i_10_401_177_0 & ~i_10_401_283_0 & i_10_401_1821_0 & ~i_10_401_1951_0 & ~i_10_401_2980_0 & ~i_10_401_4056_0 & ~i_10_401_2327_0 & ~i_10_401_2384_0))) | (~i_10_401_283_0 & ((~i_10_401_269_0 & ~i_10_401_1348_0 & i_10_401_2453_0 & ~i_10_401_4124_0) | (i_10_401_2203_0 & ~i_10_401_2829_0 & i_10_401_4117_0 & ~i_10_401_4568_0))) | (~i_10_401_4058_0 & ((~i_10_401_328_0 & ((~i_10_401_249_0 & ~i_10_401_2407_0 & ~i_10_401_2632_0 & ~i_10_401_2884_0 & ~i_10_401_2981_0 & ~i_10_401_3274_0 & ~i_10_401_4056_0 & ~i_10_401_4238_0) | (~i_10_401_34_0 & ~i_10_401_445_0 & ~i_10_401_1913_0 & ~i_10_401_2327_0 & ~i_10_401_2655_0 & ~i_10_401_2921_0 & ~i_10_401_4289_0))) | (~i_10_401_2353_0 & ~i_10_401_2411_0 & ~i_10_401_2981_0 & i_10_401_3859_0 & ~i_10_401_4056_0) | (~i_10_401_1876_0 & ~i_10_401_2186_0 & ~i_10_401_2327_0 & ~i_10_401_2407_0 & i_10_401_4117_0 & i_10_401_4118_0))) | (~i_10_401_445_0 & ((~i_10_401_1821_0 & ~i_10_401_1913_0 & ((~i_10_401_1266_0 & ~i_10_401_1951_0 & ~i_10_401_2312_0 & i_10_401_3855_0 & ~i_10_401_4056_0) | (~i_10_401_1366_0 & ~i_10_401_2184_0 & ~i_10_401_3590_0 & ~i_10_401_3855_0 & ~i_10_401_3859_0 & i_10_401_4118_0 & ~i_10_401_4238_0))) | (~i_10_401_1876_0 & ((~i_10_401_962_0 & ~i_10_401_1951_0 & ~i_10_401_2354_0 & i_10_401_3853_0 & i_10_401_3855_0) | (~i_10_401_124_0 & i_10_401_283_0 & ~i_10_401_2184_0 & ~i_10_401_2327_0 & ~i_10_401_2452_0 & i_10_401_3859_0))) | (~i_10_401_329_0 & ~i_10_401_1912_0 & ~i_10_401_2186_0 & ~i_10_401_2411_0 & ~i_10_401_2632_0 & ~i_10_401_3274_0 & ~i_10_401_4056_0))) | (~i_10_401_124_0 & ((i_10_401_2203_0 & ~i_10_401_2327_0 & i_10_401_2731_0 & i_10_401_2829_0 & i_10_401_4124_0) | (i_10_401_1825_0 & ~i_10_401_2186_0 & ~i_10_401_2407_0 & ~i_10_401_2410_0 & ~i_10_401_4237_0))) | (i_10_401_3859_0 & ((~i_10_401_2410_0 & i_10_401_2411_0 & i_10_401_2981_0) | (i_10_401_1821_0 & ~i_10_401_3274_0 & ~i_10_401_4056_0 & i_10_401_4116_0))) | (~i_10_401_3274_0 & ((~i_10_401_2184_0 & ~i_10_401_2660_0 & i_10_401_2829_0 & i_10_401_3848_0) | (~i_10_401_2329_0 & ~i_10_401_4057_0 & i_10_401_4290_0 & ~i_10_401_4568_0))) | (~i_10_401_2312_0 & ~i_10_401_2327_0 & ~i_10_401_1821_0 & ~i_10_401_1913_0 & i_10_401_2632_0 & ~i_10_401_2981_0 & ~i_10_401_4056_0 & i_10_401_4118_0));
endmodule



// Benchmark "kernel_10_402" written by ABC on Sun Jul 19 10:28:02 2020

module kernel_10_402 ( 
    i_10_402_175_0, i_10_402_178_0, i_10_402_246_0, i_10_402_247_0,
    i_10_402_249_0, i_10_402_251_0, i_10_402_284_0, i_10_402_286_0,
    i_10_402_293_0, i_10_402_322_0, i_10_402_406_0, i_10_402_409_0,
    i_10_402_410_0, i_10_402_412_0, i_10_402_460_0, i_10_402_461_0,
    i_10_402_462_0, i_10_402_463_0, i_10_402_509_0, i_10_402_800_0,
    i_10_402_964_0, i_10_402_996_0, i_10_402_997_0, i_10_402_1000_0,
    i_10_402_1236_0, i_10_402_1239_0, i_10_402_1241_0, i_10_402_1246_0,
    i_10_402_1260_0, i_10_402_1306_0, i_10_402_1313_0, i_10_402_1432_0,
    i_10_402_1434_0, i_10_402_1687_0, i_10_402_1689_0, i_10_402_1691_0,
    i_10_402_1823_0, i_10_402_2019_0, i_10_402_2020_0, i_10_402_2022_0,
    i_10_402_2023_0, i_10_402_2024_0, i_10_402_2032_0, i_10_402_2356_0,
    i_10_402_2361_0, i_10_402_2405_0, i_10_402_2450_0, i_10_402_2607_0,
    i_10_402_2608_0, i_10_402_2629_0, i_10_402_2631_0, i_10_402_2632_0,
    i_10_402_2636_0, i_10_402_2662_0, i_10_402_2677_0, i_10_402_2700_0,
    i_10_402_2704_0, i_10_402_2707_0, i_10_402_2715_0, i_10_402_2722_0,
    i_10_402_2726_0, i_10_402_2727_0, i_10_402_2781_0, i_10_402_2782_0,
    i_10_402_2784_0, i_10_402_2785_0, i_10_402_3203_0, i_10_402_3436_0,
    i_10_402_3525_0, i_10_402_3526_0, i_10_402_3650_0, i_10_402_3684_0,
    i_10_402_3784_0, i_10_402_3836_0, i_10_402_3841_0, i_10_402_3850_0,
    i_10_402_3856_0, i_10_402_3990_0, i_10_402_3991_0, i_10_402_3995_0,
    i_10_402_4053_0, i_10_402_4117_0, i_10_402_4118_0, i_10_402_4119_0,
    i_10_402_4120_0, i_10_402_4125_0, i_10_402_4126_0, i_10_402_4129_0,
    i_10_402_4130_0, i_10_402_4173_0, i_10_402_4174_0, i_10_402_4266_0,
    i_10_402_4270_0, i_10_402_4272_0, i_10_402_4273_0, i_10_402_4289_0,
    i_10_402_4290_0, i_10_402_4291_0, i_10_402_4292_0, i_10_402_4571_0,
    o_10_402_0_0  );
  input  i_10_402_175_0, i_10_402_178_0, i_10_402_246_0, i_10_402_247_0,
    i_10_402_249_0, i_10_402_251_0, i_10_402_284_0, i_10_402_286_0,
    i_10_402_293_0, i_10_402_322_0, i_10_402_406_0, i_10_402_409_0,
    i_10_402_410_0, i_10_402_412_0, i_10_402_460_0, i_10_402_461_0,
    i_10_402_462_0, i_10_402_463_0, i_10_402_509_0, i_10_402_800_0,
    i_10_402_964_0, i_10_402_996_0, i_10_402_997_0, i_10_402_1000_0,
    i_10_402_1236_0, i_10_402_1239_0, i_10_402_1241_0, i_10_402_1246_0,
    i_10_402_1260_0, i_10_402_1306_0, i_10_402_1313_0, i_10_402_1432_0,
    i_10_402_1434_0, i_10_402_1687_0, i_10_402_1689_0, i_10_402_1691_0,
    i_10_402_1823_0, i_10_402_2019_0, i_10_402_2020_0, i_10_402_2022_0,
    i_10_402_2023_0, i_10_402_2024_0, i_10_402_2032_0, i_10_402_2356_0,
    i_10_402_2361_0, i_10_402_2405_0, i_10_402_2450_0, i_10_402_2607_0,
    i_10_402_2608_0, i_10_402_2629_0, i_10_402_2631_0, i_10_402_2632_0,
    i_10_402_2636_0, i_10_402_2662_0, i_10_402_2677_0, i_10_402_2700_0,
    i_10_402_2704_0, i_10_402_2707_0, i_10_402_2715_0, i_10_402_2722_0,
    i_10_402_2726_0, i_10_402_2727_0, i_10_402_2781_0, i_10_402_2782_0,
    i_10_402_2784_0, i_10_402_2785_0, i_10_402_3203_0, i_10_402_3436_0,
    i_10_402_3525_0, i_10_402_3526_0, i_10_402_3650_0, i_10_402_3684_0,
    i_10_402_3784_0, i_10_402_3836_0, i_10_402_3841_0, i_10_402_3850_0,
    i_10_402_3856_0, i_10_402_3990_0, i_10_402_3991_0, i_10_402_3995_0,
    i_10_402_4053_0, i_10_402_4117_0, i_10_402_4118_0, i_10_402_4119_0,
    i_10_402_4120_0, i_10_402_4125_0, i_10_402_4126_0, i_10_402_4129_0,
    i_10_402_4130_0, i_10_402_4173_0, i_10_402_4174_0, i_10_402_4266_0,
    i_10_402_4270_0, i_10_402_4272_0, i_10_402_4273_0, i_10_402_4289_0,
    i_10_402_4290_0, i_10_402_4291_0, i_10_402_4292_0, i_10_402_4571_0;
  output o_10_402_0_0;
  assign o_10_402_0_0 = ~((~i_10_402_406_0 & ((~i_10_402_293_0 & ~i_10_402_997_0 & ~i_10_402_1236_0 & ~i_10_402_2361_0 & ~i_10_402_2608_0 & ~i_10_402_3203_0 & ~i_10_402_3436_0 & ~i_10_402_3684_0 & ~i_10_402_3990_0 & ~i_10_402_4126_0) | (~i_10_402_2022_0 & ~i_10_402_2023_0 & ~i_10_402_2024_0 & ~i_10_402_2607_0 & ~i_10_402_2704_0 & ~i_10_402_4173_0))) | (~i_10_402_293_0 & ((~i_10_402_246_0 & ~i_10_402_2781_0 & ~i_10_402_3436_0 & ~i_10_402_3836_0 & i_10_402_3856_0 & ~i_10_402_4053_0 & ~i_10_402_4119_0) | (~i_10_402_996_0 & ~i_10_402_1313_0 & ~i_10_402_2019_0 & ~i_10_402_2608_0 & ~i_10_402_2704_0 & ~i_10_402_3684_0 & ~i_10_402_4125_0 & ~i_10_402_4126_0 & ~i_10_402_4266_0))) | (~i_10_402_2022_0 & ((~i_10_402_246_0 & ~i_10_402_3995_0 & ((~i_10_402_251_0 & ~i_10_402_2608_0 & ~i_10_402_2781_0 & ~i_10_402_2785_0) | (~i_10_402_412_0 & ~i_10_402_1000_0 & ~i_10_402_1260_0 & ~i_10_402_3436_0 & ~i_10_402_3525_0 & ~i_10_402_3684_0 & ~i_10_402_3991_0 & ~i_10_402_4053_0 & ~i_10_402_4266_0))) | (~i_10_402_284_0 & ~i_10_402_997_0 & ~i_10_402_2019_0 & ~i_10_402_2023_0 & ~i_10_402_3850_0 & ~i_10_402_3991_0 & ~i_10_402_4053_0) | (~i_10_402_1306_0 & ~i_10_402_1691_0 & ~i_10_402_2024_0 & ~i_10_402_2782_0 & ~i_10_402_2785_0 & ~i_10_402_3525_0 & ~i_10_402_3990_0))) | (~i_10_402_2707_0 & ((~i_10_402_1691_0 & ((~i_10_402_322_0 & ~i_10_402_1823_0 & ~i_10_402_2024_0 & ~i_10_402_2607_0 & ~i_10_402_2608_0 & ~i_10_402_2715_0 & ~i_10_402_3684_0 & ~i_10_402_3990_0) | (~i_10_402_1260_0 & ~i_10_402_3526_0 & i_10_402_3650_0 & ~i_10_402_4126_0))) | (i_10_402_1689_0 & ~i_10_402_2023_0 & ~i_10_402_2782_0 & i_10_402_3841_0))) | (~i_10_402_3525_0 & ((~i_10_402_2023_0 & i_10_402_2450_0 & i_10_402_3836_0 & ~i_10_402_4173_0) | (~i_10_402_175_0 & ~i_10_402_247_0 & ~i_10_402_409_0 & ~i_10_402_2700_0 & ~i_10_402_2784_0 & ~i_10_402_3990_0 & ~i_10_402_3995_0 & ~i_10_402_4571_0))) | (i_10_402_460_0 & i_10_402_2361_0) | (~i_10_402_3991_0 & ~i_10_402_4174_0 & i_10_402_4289_0));
endmodule



// Benchmark "kernel_10_403" written by ABC on Sun Jul 19 10:28:03 2020

module kernel_10_403 ( 
    i_10_403_216_0, i_10_403_223_0, i_10_403_279_0, i_10_403_282_0,
    i_10_403_287_0, i_10_403_327_0, i_10_403_328_0, i_10_403_423_0,
    i_10_403_424_0, i_10_403_426_0, i_10_403_462_0, i_10_403_463_0,
    i_10_403_694_0, i_10_403_696_0, i_10_403_697_0, i_10_403_793_0,
    i_10_403_797_0, i_10_403_799_0, i_10_403_895_0, i_10_403_897_0,
    i_10_403_1030_0, i_10_403_1032_0, i_10_403_1033_0, i_10_403_1034_0,
    i_10_403_1035_0, i_10_403_1117_0, i_10_403_1131_0, i_10_403_1234_0,
    i_10_403_1236_0, i_10_403_1237_0, i_10_403_1346_0, i_10_403_1546_0,
    i_10_403_1548_0, i_10_403_1619_0, i_10_403_1767_0, i_10_403_1821_0,
    i_10_403_1908_0, i_10_403_1909_0, i_10_403_1911_0, i_10_403_1995_0,
    i_10_403_2002_0, i_10_403_2152_0, i_10_403_2309_0, i_10_403_2349_0,
    i_10_403_2352_0, i_10_403_2353_0, i_10_403_2406_0, i_10_403_2430_0,
    i_10_403_2456_0, i_10_403_2457_0, i_10_403_2465_0, i_10_403_2470_0,
    i_10_403_2538_0, i_10_403_2631_0, i_10_403_2634_0, i_10_403_2635_0,
    i_10_403_2636_0, i_10_403_2709_0, i_10_403_2718_0, i_10_403_2722_0,
    i_10_403_2826_0, i_10_403_2827_0, i_10_403_2888_0, i_10_403_2916_0,
    i_10_403_2922_0, i_10_403_2983_0, i_10_403_3089_0, i_10_403_3092_0,
    i_10_403_3195_0, i_10_403_3196_0, i_10_403_3199_0, i_10_403_3276_0,
    i_10_403_3277_0, i_10_403_3306_0, i_10_403_3405_0, i_10_403_3406_0,
    i_10_403_3407_0, i_10_403_3408_0, i_10_403_3409_0, i_10_403_3610_0,
    i_10_403_3613_0, i_10_403_3650_0, i_10_403_3702_0, i_10_403_3852_0,
    i_10_403_3853_0, i_10_403_3855_0, i_10_403_3856_0, i_10_403_3889_0,
    i_10_403_3901_0, i_10_403_3904_0, i_10_403_4126_0, i_10_403_4129_0,
    i_10_403_4130_0, i_10_403_4206_0, i_10_403_4219_0, i_10_403_4233_0,
    i_10_403_4290_0, i_10_403_4565_0, i_10_403_4590_0, i_10_403_4591_0,
    o_10_403_0_0  );
  input  i_10_403_216_0, i_10_403_223_0, i_10_403_279_0, i_10_403_282_0,
    i_10_403_287_0, i_10_403_327_0, i_10_403_328_0, i_10_403_423_0,
    i_10_403_424_0, i_10_403_426_0, i_10_403_462_0, i_10_403_463_0,
    i_10_403_694_0, i_10_403_696_0, i_10_403_697_0, i_10_403_793_0,
    i_10_403_797_0, i_10_403_799_0, i_10_403_895_0, i_10_403_897_0,
    i_10_403_1030_0, i_10_403_1032_0, i_10_403_1033_0, i_10_403_1034_0,
    i_10_403_1035_0, i_10_403_1117_0, i_10_403_1131_0, i_10_403_1234_0,
    i_10_403_1236_0, i_10_403_1237_0, i_10_403_1346_0, i_10_403_1546_0,
    i_10_403_1548_0, i_10_403_1619_0, i_10_403_1767_0, i_10_403_1821_0,
    i_10_403_1908_0, i_10_403_1909_0, i_10_403_1911_0, i_10_403_1995_0,
    i_10_403_2002_0, i_10_403_2152_0, i_10_403_2309_0, i_10_403_2349_0,
    i_10_403_2352_0, i_10_403_2353_0, i_10_403_2406_0, i_10_403_2430_0,
    i_10_403_2456_0, i_10_403_2457_0, i_10_403_2465_0, i_10_403_2470_0,
    i_10_403_2538_0, i_10_403_2631_0, i_10_403_2634_0, i_10_403_2635_0,
    i_10_403_2636_0, i_10_403_2709_0, i_10_403_2718_0, i_10_403_2722_0,
    i_10_403_2826_0, i_10_403_2827_0, i_10_403_2888_0, i_10_403_2916_0,
    i_10_403_2922_0, i_10_403_2983_0, i_10_403_3089_0, i_10_403_3092_0,
    i_10_403_3195_0, i_10_403_3196_0, i_10_403_3199_0, i_10_403_3276_0,
    i_10_403_3277_0, i_10_403_3306_0, i_10_403_3405_0, i_10_403_3406_0,
    i_10_403_3407_0, i_10_403_3408_0, i_10_403_3409_0, i_10_403_3610_0,
    i_10_403_3613_0, i_10_403_3650_0, i_10_403_3702_0, i_10_403_3852_0,
    i_10_403_3853_0, i_10_403_3855_0, i_10_403_3856_0, i_10_403_3889_0,
    i_10_403_3901_0, i_10_403_3904_0, i_10_403_4126_0, i_10_403_4129_0,
    i_10_403_4130_0, i_10_403_4206_0, i_10_403_4219_0, i_10_403_4233_0,
    i_10_403_4290_0, i_10_403_4565_0, i_10_403_4590_0, i_10_403_4591_0;
  output o_10_403_0_0;
  assign o_10_403_0_0 = 0;
endmodule



// Benchmark "kernel_10_404" written by ABC on Sun Jul 19 10:28:04 2020

module kernel_10_404 ( 
    i_10_404_29_0, i_10_404_49_0, i_10_404_172_0, i_10_404_176_0,
    i_10_404_194_0, i_10_404_247_0, i_10_404_280_0, i_10_404_319_0,
    i_10_404_409_0, i_10_404_428_0, i_10_404_433_0, i_10_404_434_0,
    i_10_404_464_0, i_10_404_695_0, i_10_404_700_0, i_10_404_731_0,
    i_10_404_904_0, i_10_404_992_0, i_10_404_1046_0, i_10_404_1048_0,
    i_10_404_1052_0, i_10_404_1109_0, i_10_404_1199_0, i_10_404_1233_0,
    i_10_404_1307_0, i_10_404_1309_0, i_10_404_1312_0, i_10_404_1313_0,
    i_10_404_1345_0, i_10_404_1348_0, i_10_404_1448_0, i_10_404_1550_0,
    i_10_404_1630_0, i_10_404_1650_0, i_10_404_1684_0, i_10_404_1685_0,
    i_10_404_1820_0, i_10_404_1821_0, i_10_404_1824_0, i_10_404_1825_0,
    i_10_404_1908_0, i_10_404_1913_0, i_10_404_1914_0, i_10_404_1916_0,
    i_10_404_1993_0, i_10_404_2002_0, i_10_404_2003_0, i_10_404_2091_0,
    i_10_404_2307_0, i_10_404_2309_0, i_10_404_2350_0, i_10_404_2363_0,
    i_10_404_2451_0, i_10_404_2468_0, i_10_404_2473_0, i_10_404_2515_0,
    i_10_404_2516_0, i_10_404_2601_0, i_10_404_2658_0, i_10_404_2662_0,
    i_10_404_2674_0, i_10_404_2710_0, i_10_404_2721_0, i_10_404_2818_0,
    i_10_404_2832_0, i_10_404_2920_0, i_10_404_2983_0, i_10_404_3073_0,
    i_10_404_3277_0, i_10_404_3279_0, i_10_404_3356_0, i_10_404_3387_0,
    i_10_404_3388_0, i_10_404_3389_0, i_10_404_3391_0, i_10_404_3403_0,
    i_10_404_3404_0, i_10_404_3410_0, i_10_404_3523_0, i_10_404_3583_0,
    i_10_404_3616_0, i_10_404_3617_0, i_10_404_3649_0, i_10_404_3722_0,
    i_10_404_3780_0, i_10_404_3781_0, i_10_404_3782_0, i_10_404_3837_0,
    i_10_404_3838_0, i_10_404_3853_0, i_10_404_3858_0, i_10_404_3859_0,
    i_10_404_3860_0, i_10_404_3985_0, i_10_404_4027_0, i_10_404_4031_0,
    i_10_404_4129_0, i_10_404_4285_0, i_10_404_4290_0, i_10_404_4565_0,
    o_10_404_0_0  );
  input  i_10_404_29_0, i_10_404_49_0, i_10_404_172_0, i_10_404_176_0,
    i_10_404_194_0, i_10_404_247_0, i_10_404_280_0, i_10_404_319_0,
    i_10_404_409_0, i_10_404_428_0, i_10_404_433_0, i_10_404_434_0,
    i_10_404_464_0, i_10_404_695_0, i_10_404_700_0, i_10_404_731_0,
    i_10_404_904_0, i_10_404_992_0, i_10_404_1046_0, i_10_404_1048_0,
    i_10_404_1052_0, i_10_404_1109_0, i_10_404_1199_0, i_10_404_1233_0,
    i_10_404_1307_0, i_10_404_1309_0, i_10_404_1312_0, i_10_404_1313_0,
    i_10_404_1345_0, i_10_404_1348_0, i_10_404_1448_0, i_10_404_1550_0,
    i_10_404_1630_0, i_10_404_1650_0, i_10_404_1684_0, i_10_404_1685_0,
    i_10_404_1820_0, i_10_404_1821_0, i_10_404_1824_0, i_10_404_1825_0,
    i_10_404_1908_0, i_10_404_1913_0, i_10_404_1914_0, i_10_404_1916_0,
    i_10_404_1993_0, i_10_404_2002_0, i_10_404_2003_0, i_10_404_2091_0,
    i_10_404_2307_0, i_10_404_2309_0, i_10_404_2350_0, i_10_404_2363_0,
    i_10_404_2451_0, i_10_404_2468_0, i_10_404_2473_0, i_10_404_2515_0,
    i_10_404_2516_0, i_10_404_2601_0, i_10_404_2658_0, i_10_404_2662_0,
    i_10_404_2674_0, i_10_404_2710_0, i_10_404_2721_0, i_10_404_2818_0,
    i_10_404_2832_0, i_10_404_2920_0, i_10_404_2983_0, i_10_404_3073_0,
    i_10_404_3277_0, i_10_404_3279_0, i_10_404_3356_0, i_10_404_3387_0,
    i_10_404_3388_0, i_10_404_3389_0, i_10_404_3391_0, i_10_404_3403_0,
    i_10_404_3404_0, i_10_404_3410_0, i_10_404_3523_0, i_10_404_3583_0,
    i_10_404_3616_0, i_10_404_3617_0, i_10_404_3649_0, i_10_404_3722_0,
    i_10_404_3780_0, i_10_404_3781_0, i_10_404_3782_0, i_10_404_3837_0,
    i_10_404_3838_0, i_10_404_3853_0, i_10_404_3858_0, i_10_404_3859_0,
    i_10_404_3860_0, i_10_404_3985_0, i_10_404_4027_0, i_10_404_4031_0,
    i_10_404_4129_0, i_10_404_4285_0, i_10_404_4290_0, i_10_404_4565_0;
  output o_10_404_0_0;
  assign o_10_404_0_0 = 0;
endmodule



// Benchmark "kernel_10_405" written by ABC on Sun Jul 19 10:28:05 2020

module kernel_10_405 ( 
    i_10_405_174_0, i_10_405_178_0, i_10_405_280_0, i_10_405_281_0,
    i_10_405_283_0, i_10_405_284_0, i_10_405_320_0, i_10_405_390_0,
    i_10_405_408_0, i_10_405_444_0, i_10_405_520_0, i_10_405_714_0,
    i_10_405_736_0, i_10_405_903_0, i_10_405_952_0, i_10_405_996_0,
    i_10_405_1005_0, i_10_405_1006_0, i_10_405_1039_0, i_10_405_1050_0,
    i_10_405_1051_0, i_10_405_1059_0, i_10_405_1237_0, i_10_405_1246_0,
    i_10_405_1249_0, i_10_405_1250_0, i_10_405_1311_0, i_10_405_1312_0,
    i_10_405_1313_0, i_10_405_1446_0, i_10_405_1455_0, i_10_405_1554_0,
    i_10_405_1555_0, i_10_405_1581_0, i_10_405_1735_0, i_10_405_1823_0,
    i_10_405_1909_0, i_10_405_1914_0, i_10_405_2355_0, i_10_405_2356_0,
    i_10_405_2364_0, i_10_405_2382_0, i_10_405_2383_0, i_10_405_2406_0,
    i_10_405_2407_0, i_10_405_2408_0, i_10_405_2448_0, i_10_405_2449_0,
    i_10_405_2451_0, i_10_405_2452_0, i_10_405_2464_0, i_10_405_2466_0,
    i_10_405_2467_0, i_10_405_2472_0, i_10_405_2473_0, i_10_405_2509_0,
    i_10_405_2607_0, i_10_405_2632_0, i_10_405_2636_0, i_10_405_2641_0,
    i_10_405_2662_0, i_10_405_2705_0, i_10_405_2713_0, i_10_405_2730_0,
    i_10_405_2733_0, i_10_405_2830_0, i_10_405_2834_0, i_10_405_2880_0,
    i_10_405_2884_0, i_10_405_2887_0, i_10_405_2921_0, i_10_405_2922_0,
    i_10_405_2986_0, i_10_405_3033_0, i_10_405_3040_0, i_10_405_3202_0,
    i_10_405_3291_0, i_10_405_3318_0, i_10_405_3390_0, i_10_405_3406_0,
    i_10_405_3613_0, i_10_405_3614_0, i_10_405_3646_0, i_10_405_3685_0,
    i_10_405_3725_0, i_10_405_3840_0, i_10_405_3857_0, i_10_405_3859_0,
    i_10_405_3896_0, i_10_405_3913_0, i_10_405_3914_0, i_10_405_3984_0,
    i_10_405_3985_0, i_10_405_3986_0, i_10_405_4113_0, i_10_405_4118_0,
    i_10_405_4276_0, i_10_405_4280_0, i_10_405_4281_0, i_10_405_4289_0,
    o_10_405_0_0  );
  input  i_10_405_174_0, i_10_405_178_0, i_10_405_280_0, i_10_405_281_0,
    i_10_405_283_0, i_10_405_284_0, i_10_405_320_0, i_10_405_390_0,
    i_10_405_408_0, i_10_405_444_0, i_10_405_520_0, i_10_405_714_0,
    i_10_405_736_0, i_10_405_903_0, i_10_405_952_0, i_10_405_996_0,
    i_10_405_1005_0, i_10_405_1006_0, i_10_405_1039_0, i_10_405_1050_0,
    i_10_405_1051_0, i_10_405_1059_0, i_10_405_1237_0, i_10_405_1246_0,
    i_10_405_1249_0, i_10_405_1250_0, i_10_405_1311_0, i_10_405_1312_0,
    i_10_405_1313_0, i_10_405_1446_0, i_10_405_1455_0, i_10_405_1554_0,
    i_10_405_1555_0, i_10_405_1581_0, i_10_405_1735_0, i_10_405_1823_0,
    i_10_405_1909_0, i_10_405_1914_0, i_10_405_2355_0, i_10_405_2356_0,
    i_10_405_2364_0, i_10_405_2382_0, i_10_405_2383_0, i_10_405_2406_0,
    i_10_405_2407_0, i_10_405_2408_0, i_10_405_2448_0, i_10_405_2449_0,
    i_10_405_2451_0, i_10_405_2452_0, i_10_405_2464_0, i_10_405_2466_0,
    i_10_405_2467_0, i_10_405_2472_0, i_10_405_2473_0, i_10_405_2509_0,
    i_10_405_2607_0, i_10_405_2632_0, i_10_405_2636_0, i_10_405_2641_0,
    i_10_405_2662_0, i_10_405_2705_0, i_10_405_2713_0, i_10_405_2730_0,
    i_10_405_2733_0, i_10_405_2830_0, i_10_405_2834_0, i_10_405_2880_0,
    i_10_405_2884_0, i_10_405_2887_0, i_10_405_2921_0, i_10_405_2922_0,
    i_10_405_2986_0, i_10_405_3033_0, i_10_405_3040_0, i_10_405_3202_0,
    i_10_405_3291_0, i_10_405_3318_0, i_10_405_3390_0, i_10_405_3406_0,
    i_10_405_3613_0, i_10_405_3614_0, i_10_405_3646_0, i_10_405_3685_0,
    i_10_405_3725_0, i_10_405_3840_0, i_10_405_3857_0, i_10_405_3859_0,
    i_10_405_3896_0, i_10_405_3913_0, i_10_405_3914_0, i_10_405_3984_0,
    i_10_405_3985_0, i_10_405_3986_0, i_10_405_4113_0, i_10_405_4118_0,
    i_10_405_4276_0, i_10_405_4280_0, i_10_405_4281_0, i_10_405_4289_0;
  output o_10_405_0_0;
  assign o_10_405_0_0 = 0;
endmodule



// Benchmark "kernel_10_406" written by ABC on Sun Jul 19 10:28:06 2020

module kernel_10_406 ( 
    i_10_406_30_0, i_10_406_174_0, i_10_406_220_0, i_10_406_224_0,
    i_10_406_243_0, i_10_406_246_0, i_10_406_249_0, i_10_406_250_0,
    i_10_406_280_0, i_10_406_288_0, i_10_406_325_0, i_10_406_369_0,
    i_10_406_426_0, i_10_406_438_0, i_10_406_462_0, i_10_406_465_0,
    i_10_406_534_0, i_10_406_796_0, i_10_406_900_0, i_10_406_903_0,
    i_10_406_963_0, i_10_406_1235_0, i_10_406_1260_0, i_10_406_1269_0,
    i_10_406_1270_0, i_10_406_1359_0, i_10_406_1360_0, i_10_406_1390_0,
    i_10_406_1435_0, i_10_406_1443_0, i_10_406_1548_0, i_10_406_1551_0,
    i_10_406_1683_0, i_10_406_1809_0, i_10_406_1812_0, i_10_406_1820_0,
    i_10_406_1872_0, i_10_406_1971_0, i_10_406_2023_0, i_10_406_2197_0,
    i_10_406_2250_0, i_10_406_2259_0, i_10_406_2323_0, i_10_406_2406_0,
    i_10_406_2502_0, i_10_406_2505_0, i_10_406_2515_0, i_10_406_2568_0,
    i_10_406_2604_0, i_10_406_2607_0, i_10_406_2629_0, i_10_406_2634_0,
    i_10_406_2655_0, i_10_406_2660_0, i_10_406_2661_0, i_10_406_2673_0,
    i_10_406_2700_0, i_10_406_2704_0, i_10_406_2712_0, i_10_406_2728_0,
    i_10_406_2731_0, i_10_406_2784_0, i_10_406_2787_0, i_10_406_2828_0,
    i_10_406_2829_0, i_10_406_2921_0, i_10_406_2979_0, i_10_406_3069_0,
    i_10_406_3196_0, i_10_406_3235_0, i_10_406_3270_0, i_10_406_3276_0,
    i_10_406_3277_0, i_10_406_3384_0, i_10_406_3386_0, i_10_406_3430_0,
    i_10_406_3433_0, i_10_406_3492_0, i_10_406_3610_0, i_10_406_3615_0,
    i_10_406_3681_0, i_10_406_3849_0, i_10_406_3857_0, i_10_406_3888_0,
    i_10_406_3978_0, i_10_406_3981_0, i_10_406_3993_0, i_10_406_4050_0,
    i_10_406_4053_0, i_10_406_4117_0, i_10_406_4128_0, i_10_406_4129_0,
    i_10_406_4266_0, i_10_406_4287_0, i_10_406_4365_0, i_10_406_4428_0,
    i_10_406_4429_0, i_10_406_4458_0, i_10_406_4566_0, i_10_406_4571_0,
    o_10_406_0_0  );
  input  i_10_406_30_0, i_10_406_174_0, i_10_406_220_0, i_10_406_224_0,
    i_10_406_243_0, i_10_406_246_0, i_10_406_249_0, i_10_406_250_0,
    i_10_406_280_0, i_10_406_288_0, i_10_406_325_0, i_10_406_369_0,
    i_10_406_426_0, i_10_406_438_0, i_10_406_462_0, i_10_406_465_0,
    i_10_406_534_0, i_10_406_796_0, i_10_406_900_0, i_10_406_903_0,
    i_10_406_963_0, i_10_406_1235_0, i_10_406_1260_0, i_10_406_1269_0,
    i_10_406_1270_0, i_10_406_1359_0, i_10_406_1360_0, i_10_406_1390_0,
    i_10_406_1435_0, i_10_406_1443_0, i_10_406_1548_0, i_10_406_1551_0,
    i_10_406_1683_0, i_10_406_1809_0, i_10_406_1812_0, i_10_406_1820_0,
    i_10_406_1872_0, i_10_406_1971_0, i_10_406_2023_0, i_10_406_2197_0,
    i_10_406_2250_0, i_10_406_2259_0, i_10_406_2323_0, i_10_406_2406_0,
    i_10_406_2502_0, i_10_406_2505_0, i_10_406_2515_0, i_10_406_2568_0,
    i_10_406_2604_0, i_10_406_2607_0, i_10_406_2629_0, i_10_406_2634_0,
    i_10_406_2655_0, i_10_406_2660_0, i_10_406_2661_0, i_10_406_2673_0,
    i_10_406_2700_0, i_10_406_2704_0, i_10_406_2712_0, i_10_406_2728_0,
    i_10_406_2731_0, i_10_406_2784_0, i_10_406_2787_0, i_10_406_2828_0,
    i_10_406_2829_0, i_10_406_2921_0, i_10_406_2979_0, i_10_406_3069_0,
    i_10_406_3196_0, i_10_406_3235_0, i_10_406_3270_0, i_10_406_3276_0,
    i_10_406_3277_0, i_10_406_3384_0, i_10_406_3386_0, i_10_406_3430_0,
    i_10_406_3433_0, i_10_406_3492_0, i_10_406_3610_0, i_10_406_3615_0,
    i_10_406_3681_0, i_10_406_3849_0, i_10_406_3857_0, i_10_406_3888_0,
    i_10_406_3978_0, i_10_406_3981_0, i_10_406_3993_0, i_10_406_4050_0,
    i_10_406_4053_0, i_10_406_4117_0, i_10_406_4128_0, i_10_406_4129_0,
    i_10_406_4266_0, i_10_406_4287_0, i_10_406_4365_0, i_10_406_4428_0,
    i_10_406_4429_0, i_10_406_4458_0, i_10_406_4566_0, i_10_406_4571_0;
  output o_10_406_0_0;
  assign o_10_406_0_0 = 0;
endmodule



// Benchmark "kernel_10_407" written by ABC on Sun Jul 19 10:28:07 2020

module kernel_10_407 ( 
    i_10_407_160_0, i_10_407_175_0, i_10_407_270_0, i_10_407_278_0,
    i_10_407_280_0, i_10_407_281_0, i_10_407_283_0, i_10_407_329_0,
    i_10_407_408_0, i_10_407_431_0, i_10_407_432_0, i_10_407_443_0,
    i_10_407_444_0, i_10_407_445_0, i_10_407_508_0, i_10_407_509_0,
    i_10_407_511_0, i_10_407_711_0, i_10_407_749_0, i_10_407_898_0,
    i_10_407_1142_0, i_10_407_1240_0, i_10_407_1243_0, i_10_407_1244_0,
    i_10_407_1247_0, i_10_407_1310_0, i_10_407_1348_0, i_10_407_1541_0,
    i_10_407_1552_0, i_10_407_1651_0, i_10_407_1652_0, i_10_407_1690_0,
    i_10_407_1821_0, i_10_407_1822_0, i_10_407_1823_0, i_10_407_1826_0,
    i_10_407_1996_0, i_10_407_2349_0, i_10_407_2352_0, i_10_407_2353_0,
    i_10_407_2354_0, i_10_407_2404_0, i_10_407_2455_0, i_10_407_2635_0,
    i_10_407_2659_0, i_10_407_2706_0, i_10_407_2707_0, i_10_407_2721_0,
    i_10_407_2733_0, i_10_407_2735_0, i_10_407_2884_0, i_10_407_2888_0,
    i_10_407_2919_0, i_10_407_2920_0, i_10_407_2921_0, i_10_407_2923_0,
    i_10_407_3035_0, i_10_407_3046_0, i_10_407_3150_0, i_10_407_3154_0,
    i_10_407_3155_0, i_10_407_3166_0, i_10_407_3195_0, i_10_407_3199_0,
    i_10_407_3200_0, i_10_407_3387_0, i_10_407_3388_0, i_10_407_3389_0,
    i_10_407_3390_0, i_10_407_3391_0, i_10_407_3392_0, i_10_407_3405_0,
    i_10_407_3585_0, i_10_407_3586_0, i_10_407_3587_0, i_10_407_3610_0,
    i_10_407_3611_0, i_10_407_3614_0, i_10_407_3782_0, i_10_407_3784_0,
    i_10_407_3785_0, i_10_407_3786_0, i_10_407_3837_0, i_10_407_3838_0,
    i_10_407_3839_0, i_10_407_3846_0, i_10_407_3847_0, i_10_407_3851_0,
    i_10_407_3856_0, i_10_407_3857_0, i_10_407_3980_0, i_10_407_4121_0,
    i_10_407_4123_0, i_10_407_4130_0, i_10_407_4174_0, i_10_407_4175_0,
    i_10_407_4192_0, i_10_407_4283_0, i_10_407_4292_0, i_10_407_4564_0,
    o_10_407_0_0  );
  input  i_10_407_160_0, i_10_407_175_0, i_10_407_270_0, i_10_407_278_0,
    i_10_407_280_0, i_10_407_281_0, i_10_407_283_0, i_10_407_329_0,
    i_10_407_408_0, i_10_407_431_0, i_10_407_432_0, i_10_407_443_0,
    i_10_407_444_0, i_10_407_445_0, i_10_407_508_0, i_10_407_509_0,
    i_10_407_511_0, i_10_407_711_0, i_10_407_749_0, i_10_407_898_0,
    i_10_407_1142_0, i_10_407_1240_0, i_10_407_1243_0, i_10_407_1244_0,
    i_10_407_1247_0, i_10_407_1310_0, i_10_407_1348_0, i_10_407_1541_0,
    i_10_407_1552_0, i_10_407_1651_0, i_10_407_1652_0, i_10_407_1690_0,
    i_10_407_1821_0, i_10_407_1822_0, i_10_407_1823_0, i_10_407_1826_0,
    i_10_407_1996_0, i_10_407_2349_0, i_10_407_2352_0, i_10_407_2353_0,
    i_10_407_2354_0, i_10_407_2404_0, i_10_407_2455_0, i_10_407_2635_0,
    i_10_407_2659_0, i_10_407_2706_0, i_10_407_2707_0, i_10_407_2721_0,
    i_10_407_2733_0, i_10_407_2735_0, i_10_407_2884_0, i_10_407_2888_0,
    i_10_407_2919_0, i_10_407_2920_0, i_10_407_2921_0, i_10_407_2923_0,
    i_10_407_3035_0, i_10_407_3046_0, i_10_407_3150_0, i_10_407_3154_0,
    i_10_407_3155_0, i_10_407_3166_0, i_10_407_3195_0, i_10_407_3199_0,
    i_10_407_3200_0, i_10_407_3387_0, i_10_407_3388_0, i_10_407_3389_0,
    i_10_407_3390_0, i_10_407_3391_0, i_10_407_3392_0, i_10_407_3405_0,
    i_10_407_3585_0, i_10_407_3586_0, i_10_407_3587_0, i_10_407_3610_0,
    i_10_407_3611_0, i_10_407_3614_0, i_10_407_3782_0, i_10_407_3784_0,
    i_10_407_3785_0, i_10_407_3786_0, i_10_407_3837_0, i_10_407_3838_0,
    i_10_407_3839_0, i_10_407_3846_0, i_10_407_3847_0, i_10_407_3851_0,
    i_10_407_3856_0, i_10_407_3857_0, i_10_407_3980_0, i_10_407_4121_0,
    i_10_407_4123_0, i_10_407_4130_0, i_10_407_4174_0, i_10_407_4175_0,
    i_10_407_4192_0, i_10_407_4283_0, i_10_407_4292_0, i_10_407_4564_0;
  output o_10_407_0_0;
  assign o_10_407_0_0 = ~((~i_10_407_175_0 & ((~i_10_407_408_0 & ~i_10_407_431_0 & ~i_10_407_1826_0 & ~i_10_407_2923_0 & ~i_10_407_3166_0 & ~i_10_407_3392_0 & ~i_10_407_3405_0 & ~i_10_407_3782_0 & ~i_10_407_3784_0 & ~i_10_407_3857_0 & ~i_10_407_4130_0) | (~i_10_407_1244_0 & ~i_10_407_1247_0 & ~i_10_407_1996_0 & ~i_10_407_3585_0 & ~i_10_407_3785_0 & ~i_10_407_3838_0 & ~i_10_407_4174_0))) | (~i_10_407_3857_0 & ((~i_10_407_280_0 & ((~i_10_407_431_0 & ~i_10_407_1821_0 & i_10_407_1822_0 & ~i_10_407_3046_0 & ~i_10_407_3784_0 & ~i_10_407_4121_0) | (~i_10_407_1310_0 & ~i_10_407_2659_0 & ~i_10_407_2706_0 & ~i_10_407_3166_0 & ~i_10_407_3405_0 & ~i_10_407_3611_0 & ~i_10_407_3782_0 & i_10_407_3839_0 & ~i_10_407_4174_0))) | (i_10_407_283_0 & ~i_10_407_1651_0 & ~i_10_407_1821_0 & ~i_10_407_3611_0 & ~i_10_407_3856_0) | (~i_10_407_283_0 & ~i_10_407_408_0 & ~i_10_407_1243_0 & ~i_10_407_1822_0 & ~i_10_407_1823_0 & ~i_10_407_2349_0 & ~i_10_407_2735_0 & ~i_10_407_2920_0 & ~i_10_407_2921_0 & ~i_10_407_3387_0 & ~i_10_407_3785_0 & ~i_10_407_4292_0))) | (~i_10_407_3195_0 & ((~i_10_407_281_0 & ((~i_10_407_1823_0 & ~i_10_407_2707_0 & ~i_10_407_2733_0 & ~i_10_407_2920_0 & ~i_10_407_3839_0 & i_10_407_3856_0) | (~i_10_407_2404_0 & ~i_10_407_2706_0 & ~i_10_407_2721_0 & ~i_10_407_2884_0 & ~i_10_407_2919_0 & ~i_10_407_2921_0 & ~i_10_407_3199_0 & ~i_10_407_3785_0 & ~i_10_407_4121_0 & ~i_10_407_4174_0))) | (~i_10_407_3200_0 & ((~i_10_407_1243_0 & ~i_10_407_1244_0 & i_10_407_2721_0 & ~i_10_407_2923_0 & ~i_10_407_3166_0 & ~i_10_407_3390_0) | (~i_10_407_408_0 & i_10_407_1240_0 & ~i_10_407_1826_0 & i_10_407_2659_0 & ~i_10_407_2920_0 & ~i_10_407_4175_0))) | (~i_10_407_3839_0 & ((i_10_407_432_0 & ~i_10_407_2354_0 & ~i_10_407_2888_0 & ~i_10_407_3388_0) | (~i_10_407_711_0 & i_10_407_1652_0 & ~i_10_407_1822_0 & ~i_10_407_3785_0 & ~i_10_407_4130_0))) | (~i_10_407_749_0 & ~i_10_407_2707_0 & i_10_407_3389_0 & ~i_10_407_4130_0))) | (~i_10_407_3166_0 & ((~i_10_407_408_0 & ~i_10_407_3199_0 & ((i_10_407_2455_0 & ~i_10_407_3837_0) | (~i_10_407_898_0 & ~i_10_407_1310_0 & ~i_10_407_2919_0 & ~i_10_407_2920_0 & ~i_10_407_3782_0 & ~i_10_407_4130_0))) | (~i_10_407_1243_0 & ~i_10_407_2707_0 & ~i_10_407_2919_0 & i_10_407_3388_0 & ~i_10_407_4175_0) | (~i_10_407_1821_0 & ~i_10_407_1822_0 & ~i_10_407_1823_0 & i_10_407_3035_0 & ~i_10_407_3614_0 & ~i_10_407_4292_0))) | (~i_10_407_1244_0 & ((~i_10_407_1243_0 & ~i_10_407_2733_0 & i_10_407_2920_0 & ~i_10_407_3389_0 & ~i_10_407_3585_0 & ~i_10_407_3784_0 & ~i_10_407_3839_0) | (~i_10_407_445_0 & ~i_10_407_2354_0 & ~i_10_407_2735_0 & ~i_10_407_2921_0 & ~i_10_407_3586_0 & ~i_10_407_3837_0 & ~i_10_407_4121_0))) | (~i_10_407_1552_0 & ((i_10_407_1240_0 & ~i_10_407_1310_0 & ~i_10_407_1823_0 & ~i_10_407_3199_0) | (i_10_407_445_0 & ~i_10_407_749_0 & ~i_10_407_3838_0 & ~i_10_407_4292_0))) | (~i_10_407_4283_0 & ((~i_10_407_749_0 & ((~i_10_407_431_0 & ~i_10_407_444_0 & ~i_10_407_2884_0 & ~i_10_407_3200_0 & ~i_10_407_3405_0 & ~i_10_407_3784_0) | (i_10_407_3387_0 & ~i_10_407_3839_0))) | (i_10_407_283_0 & ~i_10_407_1690_0 & ~i_10_407_2920_0 & ~i_10_407_2923_0 & ~i_10_407_3587_0 & ~i_10_407_3785_0 & i_10_407_3856_0))) | (~i_10_407_1310_0 & ((~i_10_407_3200_0 & i_10_407_3846_0) | (~i_10_407_1652_0 & ~i_10_407_2733_0 & ~i_10_407_3610_0 & i_10_407_3837_0 & ~i_10_407_3856_0 & ~i_10_407_4130_0))) | (~i_10_407_1821_0 & i_10_407_2349_0 & i_10_407_2919_0) | (~i_10_407_1240_0 & ~i_10_407_1823_0 & ~i_10_407_2707_0 & ~i_10_407_3199_0 & ~i_10_407_3614_0 & ~i_10_407_3784_0) | (~i_10_407_432_0 & i_10_407_443_0 & ~i_10_407_2721_0 & i_10_407_3035_0 & ~i_10_407_3839_0 & i_10_407_4121_0));
endmodule



// Benchmark "kernel_10_408" written by ABC on Sun Jul 19 10:28:09 2020

module kernel_10_408 ( 
    i_10_408_216_0, i_10_408_217_0, i_10_408_218_0, i_10_408_275_0,
    i_10_408_278_0, i_10_408_280_0, i_10_408_281_0, i_10_408_282_0,
    i_10_408_283_0, i_10_408_284_0, i_10_408_316_0, i_10_408_317_0,
    i_10_408_319_0, i_10_408_320_0, i_10_408_444_0, i_10_408_461_0,
    i_10_408_464_0, i_10_408_466_0, i_10_408_467_0, i_10_408_799_0,
    i_10_408_851_0, i_10_408_854_0, i_10_408_1006_0, i_10_408_1027_0,
    i_10_408_1030_0, i_10_408_1034_0, i_10_408_1083_0, i_10_408_1237_0,
    i_10_408_1240_0, i_10_408_1242_0, i_10_408_1243_0, i_10_408_1307_0,
    i_10_408_1648_0, i_10_408_1649_0, i_10_408_1684_0, i_10_408_1685_0,
    i_10_408_1688_0, i_10_408_1819_0, i_10_408_2002_0, i_10_408_2305_0,
    i_10_408_2306_0, i_10_408_2351_0, i_10_408_2358_0, i_10_408_2362_0,
    i_10_408_2363_0, i_10_408_2364_0, i_10_408_2449_0, i_10_408_2460_0,
    i_10_408_2470_0, i_10_408_2701_0, i_10_408_2702_0, i_10_408_2703_0,
    i_10_408_2710_0, i_10_408_2718_0, i_10_408_2719_0, i_10_408_2720_0,
    i_10_408_2722_0, i_10_408_2919_0, i_10_408_2920_0, i_10_408_2921_0,
    i_10_408_2923_0, i_10_408_2924_0, i_10_408_3088_0, i_10_408_3089_0,
    i_10_408_3267_0, i_10_408_3270_0, i_10_408_3277_0, i_10_408_3322_0,
    i_10_408_3328_0, i_10_408_3385_0, i_10_408_3386_0, i_10_408_3402_0,
    i_10_408_3403_0, i_10_408_3404_0, i_10_408_3405_0, i_10_408_3406_0,
    i_10_408_3407_0, i_10_408_3466_0, i_10_408_3469_0, i_10_408_3551_0,
    i_10_408_3611_0, i_10_408_3780_0, i_10_408_3781_0, i_10_408_3783_0,
    i_10_408_3784_0, i_10_408_3844_0, i_10_408_3847_0, i_10_408_3851_0,
    i_10_408_3855_0, i_10_408_3856_0, i_10_408_3857_0, i_10_408_3979_0,
    i_10_408_4212_0, i_10_408_4214_0, i_10_408_4273_0, i_10_408_4284_0,
    i_10_408_4285_0, i_10_408_4565_0, i_10_408_4567_0, i_10_408_4569_0,
    o_10_408_0_0  );
  input  i_10_408_216_0, i_10_408_217_0, i_10_408_218_0, i_10_408_275_0,
    i_10_408_278_0, i_10_408_280_0, i_10_408_281_0, i_10_408_282_0,
    i_10_408_283_0, i_10_408_284_0, i_10_408_316_0, i_10_408_317_0,
    i_10_408_319_0, i_10_408_320_0, i_10_408_444_0, i_10_408_461_0,
    i_10_408_464_0, i_10_408_466_0, i_10_408_467_0, i_10_408_799_0,
    i_10_408_851_0, i_10_408_854_0, i_10_408_1006_0, i_10_408_1027_0,
    i_10_408_1030_0, i_10_408_1034_0, i_10_408_1083_0, i_10_408_1237_0,
    i_10_408_1240_0, i_10_408_1242_0, i_10_408_1243_0, i_10_408_1307_0,
    i_10_408_1648_0, i_10_408_1649_0, i_10_408_1684_0, i_10_408_1685_0,
    i_10_408_1688_0, i_10_408_1819_0, i_10_408_2002_0, i_10_408_2305_0,
    i_10_408_2306_0, i_10_408_2351_0, i_10_408_2358_0, i_10_408_2362_0,
    i_10_408_2363_0, i_10_408_2364_0, i_10_408_2449_0, i_10_408_2460_0,
    i_10_408_2470_0, i_10_408_2701_0, i_10_408_2702_0, i_10_408_2703_0,
    i_10_408_2710_0, i_10_408_2718_0, i_10_408_2719_0, i_10_408_2720_0,
    i_10_408_2722_0, i_10_408_2919_0, i_10_408_2920_0, i_10_408_2921_0,
    i_10_408_2923_0, i_10_408_2924_0, i_10_408_3088_0, i_10_408_3089_0,
    i_10_408_3267_0, i_10_408_3270_0, i_10_408_3277_0, i_10_408_3322_0,
    i_10_408_3328_0, i_10_408_3385_0, i_10_408_3386_0, i_10_408_3402_0,
    i_10_408_3403_0, i_10_408_3404_0, i_10_408_3405_0, i_10_408_3406_0,
    i_10_408_3407_0, i_10_408_3466_0, i_10_408_3469_0, i_10_408_3551_0,
    i_10_408_3611_0, i_10_408_3780_0, i_10_408_3781_0, i_10_408_3783_0,
    i_10_408_3784_0, i_10_408_3844_0, i_10_408_3847_0, i_10_408_3851_0,
    i_10_408_3855_0, i_10_408_3856_0, i_10_408_3857_0, i_10_408_3979_0,
    i_10_408_4212_0, i_10_408_4214_0, i_10_408_4273_0, i_10_408_4284_0,
    i_10_408_4285_0, i_10_408_4565_0, i_10_408_4567_0, i_10_408_4569_0;
  output o_10_408_0_0;
  assign o_10_408_0_0 = ~((~i_10_408_281_0 & ((~i_10_408_316_0 & ~i_10_408_1034_0 & i_10_408_2710_0 & ~i_10_408_2920_0 & ~i_10_408_2921_0 & ~i_10_408_3466_0 & ~i_10_408_3784_0) | (~i_10_408_217_0 & ~i_10_408_283_0 & ~i_10_408_320_0 & ~i_10_408_1307_0 & i_10_408_2722_0 & i_10_408_3386_0 & ~i_10_408_3855_0))) | (~i_10_408_4569_0 & ((~i_10_408_283_0 & ((~i_10_408_2363_0 & ~i_10_408_3385_0 & ~i_10_408_3611_0 & ~i_10_408_3784_0) | (i_10_408_280_0 & ~i_10_408_1242_0 & i_10_408_3385_0 & ~i_10_408_3847_0))) | (~i_10_408_1685_0 & ~i_10_408_2719_0 & ~i_10_408_2722_0 & i_10_408_2919_0 & ~i_10_408_3277_0 & ~i_10_408_3784_0))) | (~i_10_408_284_0 & ((i_10_408_466_0 & ~i_10_408_3270_0 & ~i_10_408_3386_0 & ~i_10_408_3402_0 & ~i_10_408_3844_0) | (i_10_408_281_0 & ~i_10_408_1243_0 & ~i_10_408_2364_0 & i_10_408_3611_0 & ~i_10_408_3847_0))) | (~i_10_408_1034_0 & ((~i_10_408_216_0 & ~i_10_408_217_0 & ~i_10_408_218_0 & ~i_10_408_1030_0 & ~i_10_408_1685_0 & ~i_10_408_2460_0 & ~i_10_408_3089_0) | (~i_10_408_1242_0 & ~i_10_408_2919_0 & ~i_10_408_2920_0 & ~i_10_408_2923_0 & ~i_10_408_3402_0))) | (~i_10_408_217_0 & ((~i_10_408_1243_0 & ~i_10_408_2364_0 & ~i_10_408_2710_0 & ~i_10_408_3403_0 & ~i_10_408_4214_0) | (~i_10_408_461_0 & ~i_10_408_2363_0 & ~i_10_408_3270_0 & ~i_10_408_3385_0 & ~i_10_408_4567_0))) | (~i_10_408_218_0 & ((i_10_408_467_0 & ~i_10_408_3385_0) | (i_10_408_1030_0 & ~i_10_408_1684_0 & ~i_10_408_2305_0 & ~i_10_408_2921_0 & ~i_10_408_3403_0))) | (~i_10_408_1243_0 & ((~i_10_408_1027_0 & ~i_10_408_3405_0 & ~i_10_408_3407_0) | (i_10_408_2919_0 & ~i_10_408_3267_0 & ~i_10_408_3277_0 & ~i_10_408_3847_0 & ~i_10_408_3856_0))) | (~i_10_408_1684_0 & ~i_10_408_2919_0 & ((~i_10_408_1685_0 & ~i_10_408_2306_0 & ~i_10_408_2362_0) | (~i_10_408_2363_0 & ~i_10_408_2460_0 & ~i_10_408_2722_0 & i_10_408_3406_0 & ~i_10_408_3847_0))) | (i_10_408_799_0 & i_10_408_2363_0 & i_10_408_2364_0) | (~i_10_408_282_0 & ~i_10_408_2703_0 & ~i_10_408_3402_0 & ~i_10_408_3406_0 & ~i_10_408_3857_0) | (i_10_408_1027_0 & i_10_408_1684_0 & ~i_10_408_2363_0 & ~i_10_408_3404_0 & ~i_10_408_3781_0 & ~i_10_408_4212_0));
endmodule



// Benchmark "kernel_10_409" written by ABC on Sun Jul 19 10:28:10 2020

module kernel_10_409 ( 
    i_10_409_27_0, i_10_409_28_0, i_10_409_30_0, i_10_409_117_0,
    i_10_409_216_0, i_10_409_220_0, i_10_409_221_0, i_10_409_280_0,
    i_10_409_283_0, i_10_409_285_0, i_10_409_286_0, i_10_409_442_0,
    i_10_409_465_0, i_10_409_508_0, i_10_409_514_0, i_10_409_748_0,
    i_10_409_893_0, i_10_409_955_0, i_10_409_961_0, i_10_409_1238_0,
    i_10_409_1242_0, i_10_409_1243_0, i_10_409_1244_0, i_10_409_1250_0,
    i_10_409_1305_0, i_10_409_1306_0, i_10_409_1308_0, i_10_409_1309_0,
    i_10_409_1310_0, i_10_409_1311_0, i_10_409_1359_0, i_10_409_1360_0,
    i_10_409_1444_0, i_10_409_1552_0, i_10_409_1575_0, i_10_409_1578_0,
    i_10_409_1647_0, i_10_409_1650_0, i_10_409_1819_0, i_10_409_1821_0,
    i_10_409_1823_0, i_10_409_1913_0, i_10_409_1947_0, i_10_409_1998_0,
    i_10_409_2349_0, i_10_409_2449_0, i_10_409_2450_0, i_10_409_2452_0,
    i_10_409_2601_0, i_10_409_2628_0, i_10_409_2629_0, i_10_409_2631_0,
    i_10_409_2658_0, i_10_409_2673_0, i_10_409_2710_0, i_10_409_2711_0,
    i_10_409_2713_0, i_10_409_2714_0, i_10_409_2721_0, i_10_409_2725_0,
    i_10_409_2726_0, i_10_409_2735_0, i_10_409_2784_0, i_10_409_2887_0,
    i_10_409_2982_0, i_10_409_3033_0, i_10_409_3034_0, i_10_409_3036_0,
    i_10_409_3037_0, i_10_409_3038_0, i_10_409_3039_0, i_10_409_3040_0,
    i_10_409_3069_0, i_10_409_3089_0, i_10_409_3281_0, i_10_409_3386_0,
    i_10_409_3387_0, i_10_409_3388_0, i_10_409_3390_0, i_10_409_3391_0,
    i_10_409_3405_0, i_10_409_3502_0, i_10_409_3519_0, i_10_409_3583_0,
    i_10_409_3613_0, i_10_409_3645_0, i_10_409_3646_0, i_10_409_3647_0,
    i_10_409_3648_0, i_10_409_3649_0, i_10_409_3652_0, i_10_409_3780_0,
    i_10_409_3782_0, i_10_409_3783_0, i_10_409_3834_0, i_10_409_3849_0,
    i_10_409_3857_0, i_10_409_4213_0, i_10_409_4292_0, i_10_409_4565_0,
    o_10_409_0_0  );
  input  i_10_409_27_0, i_10_409_28_0, i_10_409_30_0, i_10_409_117_0,
    i_10_409_216_0, i_10_409_220_0, i_10_409_221_0, i_10_409_280_0,
    i_10_409_283_0, i_10_409_285_0, i_10_409_286_0, i_10_409_442_0,
    i_10_409_465_0, i_10_409_508_0, i_10_409_514_0, i_10_409_748_0,
    i_10_409_893_0, i_10_409_955_0, i_10_409_961_0, i_10_409_1238_0,
    i_10_409_1242_0, i_10_409_1243_0, i_10_409_1244_0, i_10_409_1250_0,
    i_10_409_1305_0, i_10_409_1306_0, i_10_409_1308_0, i_10_409_1309_0,
    i_10_409_1310_0, i_10_409_1311_0, i_10_409_1359_0, i_10_409_1360_0,
    i_10_409_1444_0, i_10_409_1552_0, i_10_409_1575_0, i_10_409_1578_0,
    i_10_409_1647_0, i_10_409_1650_0, i_10_409_1819_0, i_10_409_1821_0,
    i_10_409_1823_0, i_10_409_1913_0, i_10_409_1947_0, i_10_409_1998_0,
    i_10_409_2349_0, i_10_409_2449_0, i_10_409_2450_0, i_10_409_2452_0,
    i_10_409_2601_0, i_10_409_2628_0, i_10_409_2629_0, i_10_409_2631_0,
    i_10_409_2658_0, i_10_409_2673_0, i_10_409_2710_0, i_10_409_2711_0,
    i_10_409_2713_0, i_10_409_2714_0, i_10_409_2721_0, i_10_409_2725_0,
    i_10_409_2726_0, i_10_409_2735_0, i_10_409_2784_0, i_10_409_2887_0,
    i_10_409_2982_0, i_10_409_3033_0, i_10_409_3034_0, i_10_409_3036_0,
    i_10_409_3037_0, i_10_409_3038_0, i_10_409_3039_0, i_10_409_3040_0,
    i_10_409_3069_0, i_10_409_3089_0, i_10_409_3281_0, i_10_409_3386_0,
    i_10_409_3387_0, i_10_409_3388_0, i_10_409_3390_0, i_10_409_3391_0,
    i_10_409_3405_0, i_10_409_3502_0, i_10_409_3519_0, i_10_409_3583_0,
    i_10_409_3613_0, i_10_409_3645_0, i_10_409_3646_0, i_10_409_3647_0,
    i_10_409_3648_0, i_10_409_3649_0, i_10_409_3652_0, i_10_409_3780_0,
    i_10_409_3782_0, i_10_409_3783_0, i_10_409_3834_0, i_10_409_3849_0,
    i_10_409_3857_0, i_10_409_4213_0, i_10_409_4292_0, i_10_409_4565_0;
  output o_10_409_0_0;
  assign o_10_409_0_0 = ~((~i_10_409_748_0 & ((i_10_409_1310_0 & ~i_10_409_1647_0 & ~i_10_409_2628_0 & ~i_10_409_3036_0 & ~i_10_409_3037_0 & ~i_10_409_3645_0) | (~i_10_409_221_0 & ~i_10_409_1913_0 & ~i_10_409_2673_0 & ~i_10_409_3033_0 & ~i_10_409_3034_0 & ~i_10_409_3038_0 & ~i_10_409_3648_0))) | (~i_10_409_117_0 & ((~i_10_409_1242_0 & ((~i_10_409_28_0 & ~i_10_409_1308_0 & ~i_10_409_1575_0 & ~i_10_409_1647_0 & ~i_10_409_3036_0) | (~i_10_409_1913_0 & ~i_10_409_2601_0 & ~i_10_409_2784_0 & ~i_10_409_3037_0 & ~i_10_409_3646_0 & ~i_10_409_3783_0))) | (~i_10_409_30_0 & ~i_10_409_216_0 & i_10_409_1238_0 & ~i_10_409_1360_0 & ~i_10_409_1647_0 & ~i_10_409_1998_0 & ~i_10_409_2982_0 & ~i_10_409_3039_0))) | (~i_10_409_2601_0 & ((~i_10_409_1309_0 & ((~i_10_409_286_0 & ~i_10_409_955_0 & ~i_10_409_961_0 & ~i_10_409_1308_0 & ~i_10_409_1821_0 & ~i_10_409_1913_0 & ~i_10_409_2725_0 & ~i_10_409_3040_0) | (~i_10_409_3069_0 & ~i_10_409_3281_0 & i_10_409_3391_0))) | (~i_10_409_1578_0 & ~i_10_409_2452_0 & ~i_10_409_2658_0 & ~i_10_409_2721_0 & ~i_10_409_2887_0 & ~i_10_409_3033_0 & ~i_10_409_3405_0 & ~i_10_409_3647_0 & ~i_10_409_3849_0 & ~i_10_409_3857_0))) | (~i_10_409_1578_0 & ((~i_10_409_1238_0 & i_10_409_1823_0 & ~i_10_409_1947_0 & ~i_10_409_2658_0 & ~i_10_409_3647_0) | (i_10_409_2721_0 & ~i_10_409_3645_0 & ~i_10_409_3646_0 & i_10_409_3857_0))) | (~i_10_409_1998_0 & ((i_10_409_283_0 & ~i_10_409_2628_0 & ~i_10_409_3089_0 & ~i_10_409_3390_0 & ~i_10_409_3652_0 & ~i_10_409_3782_0 & ~i_10_409_3783_0) | (i_10_409_286_0 & ~i_10_409_1305_0 & ~i_10_409_2449_0 & ~i_10_409_2735_0 & ~i_10_409_3647_0 & ~i_10_409_3834_0))) | (~i_10_409_3036_0 & ((i_10_409_3038_0 & ~i_10_409_3040_0 & ~i_10_409_3647_0) | (~i_10_409_220_0 & ~i_10_409_1819_0 & ~i_10_409_2982_0 & ~i_10_409_3386_0 & ~i_10_409_3645_0 & ~i_10_409_3783_0 & ~i_10_409_3857_0))) | (~i_10_409_2982_0 & ((~i_10_409_283_0 & i_10_409_1306_0 & ~i_10_409_2658_0 & ~i_10_409_3645_0) | (~i_10_409_2673_0 & ~i_10_409_3033_0 & i_10_409_3388_0 & ~i_10_409_3780_0))) | (~i_10_409_2658_0 & ((~i_10_409_285_0 & i_10_409_2631_0 & ~i_10_409_2721_0 & ~i_10_409_2784_0 & ~i_10_409_3645_0 & ~i_10_409_3646_0) | (i_10_409_285_0 & i_10_409_2735_0 & i_10_409_3038_0 & ~i_10_409_3647_0))) | (~i_10_409_3039_0 & ((~i_10_409_1359_0 & ~i_10_409_3646_0 & ~i_10_409_3649_0) | (~i_10_409_3783_0 & ~i_10_409_3857_0 & ~i_10_409_1650_0 & ~i_10_409_3645_0))) | (i_10_409_442_0 & ~i_10_409_514_0 & ~i_10_409_3040_0 & i_10_409_3089_0 & ~i_10_409_3645_0) | (~i_10_409_2631_0 & ~i_10_409_3038_0 & i_10_409_3281_0 & ~i_10_409_3646_0));
endmodule



// Benchmark "kernel_10_410" written by ABC on Sun Jul 19 10:28:12 2020

module kernel_10_410 ( 
    i_10_410_171_0, i_10_410_279_0, i_10_410_285_0, i_10_410_286_0,
    i_10_410_292_0, i_10_410_390_0, i_10_410_393_0, i_10_410_394_0,
    i_10_410_412_0, i_10_410_435_0, i_10_410_441_0, i_10_410_442_0,
    i_10_410_462_0, i_10_410_463_0, i_10_410_464_0, i_10_410_466_0,
    i_10_410_467_0, i_10_410_509_0, i_10_410_699_0, i_10_410_700_0,
    i_10_410_750_0, i_10_410_996_0, i_10_410_1237_0, i_10_410_1238_0,
    i_10_410_1239_0, i_10_410_1240_0, i_10_410_1241_0, i_10_410_1308_0,
    i_10_410_1362_0, i_10_410_1363_0, i_10_410_1542_0, i_10_410_1546_0,
    i_10_410_1551_0, i_10_410_1552_0, i_10_410_1554_0, i_10_410_1578_0,
    i_10_410_1579_0, i_10_410_1581_0, i_10_410_1690_0, i_10_410_1824_0,
    i_10_410_1914_0, i_10_410_2158_0, i_10_410_2159_0, i_10_410_2202_0,
    i_10_410_2310_0, i_10_410_2311_0, i_10_410_2312_0, i_10_410_2355_0,
    i_10_410_2356_0, i_10_410_2357_0, i_10_410_2360_0, i_10_410_2382_0,
    i_10_410_2408_0, i_10_410_2452_0, i_10_410_2481_0, i_10_410_2656_0,
    i_10_410_2706_0, i_10_410_2721_0, i_10_410_2880_0, i_10_410_2881_0,
    i_10_410_2884_0, i_10_410_2886_0, i_10_410_2958_0, i_10_410_3039_0,
    i_10_410_3041_0, i_10_410_3153_0, i_10_410_3158_0, i_10_410_3195_0,
    i_10_410_3273_0, i_10_410_3275_0, i_10_410_3279_0, i_10_410_3280_0,
    i_10_410_3283_0, i_10_410_3324_0, i_10_410_3325_0, i_10_410_3328_0,
    i_10_410_3329_0, i_10_410_3387_0, i_10_410_3390_0, i_10_410_3391_0,
    i_10_410_3540_0, i_10_410_3588_0, i_10_410_3782_0, i_10_410_3843_0,
    i_10_410_3856_0, i_10_410_3857_0, i_10_410_3859_0, i_10_410_3964_0,
    i_10_410_3965_0, i_10_410_3981_0, i_10_410_3982_0, i_10_410_3984_0,
    i_10_410_3985_0, i_10_410_4057_0, i_10_410_4115_0, i_10_410_4129_0,
    i_10_410_4173_0, i_10_410_4278_0, i_10_410_4279_0, i_10_410_4281_0,
    o_10_410_0_0  );
  input  i_10_410_171_0, i_10_410_279_0, i_10_410_285_0, i_10_410_286_0,
    i_10_410_292_0, i_10_410_390_0, i_10_410_393_0, i_10_410_394_0,
    i_10_410_412_0, i_10_410_435_0, i_10_410_441_0, i_10_410_442_0,
    i_10_410_462_0, i_10_410_463_0, i_10_410_464_0, i_10_410_466_0,
    i_10_410_467_0, i_10_410_509_0, i_10_410_699_0, i_10_410_700_0,
    i_10_410_750_0, i_10_410_996_0, i_10_410_1237_0, i_10_410_1238_0,
    i_10_410_1239_0, i_10_410_1240_0, i_10_410_1241_0, i_10_410_1308_0,
    i_10_410_1362_0, i_10_410_1363_0, i_10_410_1542_0, i_10_410_1546_0,
    i_10_410_1551_0, i_10_410_1552_0, i_10_410_1554_0, i_10_410_1578_0,
    i_10_410_1579_0, i_10_410_1581_0, i_10_410_1690_0, i_10_410_1824_0,
    i_10_410_1914_0, i_10_410_2158_0, i_10_410_2159_0, i_10_410_2202_0,
    i_10_410_2310_0, i_10_410_2311_0, i_10_410_2312_0, i_10_410_2355_0,
    i_10_410_2356_0, i_10_410_2357_0, i_10_410_2360_0, i_10_410_2382_0,
    i_10_410_2408_0, i_10_410_2452_0, i_10_410_2481_0, i_10_410_2656_0,
    i_10_410_2706_0, i_10_410_2721_0, i_10_410_2880_0, i_10_410_2881_0,
    i_10_410_2884_0, i_10_410_2886_0, i_10_410_2958_0, i_10_410_3039_0,
    i_10_410_3041_0, i_10_410_3153_0, i_10_410_3158_0, i_10_410_3195_0,
    i_10_410_3273_0, i_10_410_3275_0, i_10_410_3279_0, i_10_410_3280_0,
    i_10_410_3283_0, i_10_410_3324_0, i_10_410_3325_0, i_10_410_3328_0,
    i_10_410_3329_0, i_10_410_3387_0, i_10_410_3390_0, i_10_410_3391_0,
    i_10_410_3540_0, i_10_410_3588_0, i_10_410_3782_0, i_10_410_3843_0,
    i_10_410_3856_0, i_10_410_3857_0, i_10_410_3859_0, i_10_410_3964_0,
    i_10_410_3965_0, i_10_410_3981_0, i_10_410_3982_0, i_10_410_3984_0,
    i_10_410_3985_0, i_10_410_4057_0, i_10_410_4115_0, i_10_410_4129_0,
    i_10_410_4173_0, i_10_410_4278_0, i_10_410_4279_0, i_10_410_4281_0;
  output o_10_410_0_0;
  assign o_10_410_0_0 = ~((~i_10_410_3273_0 & ((~i_10_410_390_0 & ((~i_10_410_1579_0 & ~i_10_410_2202_0 & ~i_10_410_2382_0 & ~i_10_410_2884_0 & ~i_10_410_3275_0 & ~i_10_410_3279_0 & ~i_10_410_3390_0 & ~i_10_410_3856_0) | (~i_10_410_699_0 & ~i_10_410_750_0 & ~i_10_410_1546_0 & ~i_10_410_1554_0 & ~i_10_410_1690_0 & ~i_10_410_2310_0 & ~i_10_410_2311_0 & ~i_10_410_2312_0 & ~i_10_410_2481_0 & ~i_10_410_2880_0 & ~i_10_410_4173_0 & ~i_10_410_4278_0 & ~i_10_410_4279_0 & ~i_10_410_4281_0))) | (~i_10_410_393_0 & ~i_10_410_2312_0 & ~i_10_410_2481_0 & ~i_10_410_3985_0 & ~i_10_410_4278_0 & ((~i_10_410_286_0 & ~i_10_410_394_0 & ~i_10_410_435_0 & ~i_10_410_700_0 & ~i_10_410_996_0 & ~i_10_410_1542_0 & ~i_10_410_1546_0 & ~i_10_410_2202_0 & ~i_10_410_3856_0 & ~i_10_410_3981_0) | (~i_10_410_463_0 & ~i_10_410_750_0 & ~i_10_410_1552_0 & ~i_10_410_2886_0 & ~i_10_410_3039_0 & ~i_10_410_3041_0 & ~i_10_410_3195_0 & ~i_10_410_3843_0 & ~i_10_410_4279_0))) | (i_10_410_462_0 & ~i_10_410_699_0 & ~i_10_410_1552_0 & ~i_10_410_1581_0 & ~i_10_410_2356_0 & ~i_10_410_4129_0) | (i_10_410_463_0 & i_10_410_464_0 & i_10_410_467_0 & ~i_10_410_2886_0 & ~i_10_410_4173_0))) | (~i_10_410_2311_0 & ((~i_10_410_171_0 & ((i_10_410_466_0 & i_10_410_467_0 & ~i_10_410_1579_0 & ~i_10_410_2452_0) | (~i_10_410_1554_0 & ~i_10_410_1581_0 & ~i_10_410_2312_0 & ~i_10_410_2481_0 & ~i_10_410_2880_0 & ~i_10_410_2886_0 & i_10_410_3982_0 & ~i_10_410_4129_0))) | (~i_10_410_286_0 & ((~i_10_410_394_0 & ~i_10_410_441_0 & ~i_10_410_1554_0 & ~i_10_410_1578_0 & ~i_10_410_1581_0 & ~i_10_410_2312_0 & ~i_10_410_2356_0 & ~i_10_410_2884_0 & ~i_10_410_3280_0) | (i_10_410_1240_0 & i_10_410_1690_0 & ~i_10_410_2310_0 & ~i_10_410_4279_0 & ~i_10_410_4281_0))) | (~i_10_410_279_0 & ~i_10_410_1552_0 & ~i_10_410_1581_0 & ~i_10_410_1824_0 & ~i_10_410_2356_0 & ~i_10_410_2452_0 & ~i_10_410_2881_0 & ~i_10_410_3856_0 & ~i_10_410_3857_0))) | (~i_10_410_171_0 & ((~i_10_410_467_0 & i_10_410_1238_0 & ~i_10_410_1308_0 & ~i_10_410_1542_0 & ~i_10_410_2382_0 & ~i_10_410_3275_0 & ~i_10_410_3540_0) | (~i_10_410_1552_0 & ~i_10_410_2886_0 & i_10_410_466_0 & ~i_10_410_699_0 & ~i_10_410_3390_0 & ~i_10_410_3843_0 & ~i_10_410_3982_0 & ~i_10_410_3985_0))) | (~i_10_410_1690_0 & ((~i_10_410_279_0 & ((~i_10_410_435_0 & ~i_10_410_1581_0 & i_10_410_1824_0 & ~i_10_410_2355_0 & ~i_10_410_3280_0 & ~i_10_410_3985_0) | (~i_10_410_393_0 & ~i_10_410_1542_0 & ~i_10_410_1551_0 & ~i_10_410_2202_0 & ~i_10_410_2884_0 & i_10_410_3856_0 & ~i_10_410_4278_0))) | (i_10_410_463_0 & ~i_10_410_699_0 & ~i_10_410_996_0 & ~i_10_410_1579_0 & ~i_10_410_3982_0 & ~i_10_410_3985_0 & ~i_10_410_2312_0 & ~i_10_410_3280_0))) | (~i_10_410_2355_0 & ((~i_10_410_467_0 & ((i_10_410_466_0 & i_10_410_2408_0) | (~i_10_410_700_0 & ~i_10_410_1238_0 & ~i_10_410_1542_0 & ~i_10_410_1551_0 & ~i_10_410_1581_0 & ~i_10_410_2356_0 & ~i_10_410_2721_0 & ~i_10_410_3195_0 & ~i_10_410_3982_0 & ~i_10_410_4115_0 & ~i_10_410_4173_0))) | (~i_10_410_700_0 & ~i_10_410_1578_0 & ~i_10_410_1579_0 & ~i_10_410_3275_0 & ~i_10_410_3981_0 & i_10_410_3982_0))) | (~i_10_410_2202_0 & ((~i_10_410_1552_0 & ~i_10_410_3856_0 & ~i_10_410_4278_0 & ((~i_10_410_393_0 & ~i_10_410_750_0 & ~i_10_410_2706_0 & ~i_10_410_2884_0 & ~i_10_410_3390_0 & ~i_10_410_3391_0 & ~i_10_410_3843_0) | (~i_10_410_2312_0 & ~i_10_410_2382_0 & ~i_10_410_3195_0 & ~i_10_410_3387_0 & ~i_10_410_3982_0 & ~i_10_410_3985_0 & ~i_10_410_4115_0))) | (~i_10_410_1578_0 & ~i_10_410_2452_0 & ~i_10_410_2721_0 & i_10_410_2880_0))) | (~i_10_410_2881_0 & ((~i_10_410_1581_0 & i_10_410_3195_0 & ~i_10_410_3280_0 & ~i_10_410_3391_0 & ~i_10_410_4115_0 & ~i_10_410_4279_0) | (i_10_410_286_0 & ~i_10_410_700_0 & ~i_10_410_1239_0 & ~i_10_410_1542_0 & ~i_10_410_3275_0 & ~i_10_410_3279_0 & ~i_10_410_3984_0 & ~i_10_410_4281_0))) | (i_10_410_463_0 & ~i_10_410_1578_0 & ~i_10_410_1824_0 & i_10_410_2656_0 & ~i_10_410_3391_0) | (i_10_410_412_0 & ~i_10_410_435_0 & ~i_10_410_2884_0) | (~i_10_410_3982_0 & ~i_10_410_3985_0 & i_10_410_442_0 & i_10_410_2408_0) | (~i_10_410_1554_0 & ~i_10_410_2310_0 & i_10_410_3588_0 & ~i_10_410_3857_0 & ~i_10_410_3984_0 & ~i_10_410_4278_0));
endmodule



// Benchmark "kernel_10_411" written by ABC on Sun Jul 19 10:28:13 2020

module kernel_10_411 ( 
    i_10_411_145_0, i_10_411_220_0, i_10_411_223_0, i_10_411_271_0,
    i_10_411_272_0, i_10_411_273_0, i_10_411_276_0, i_10_411_283_0,
    i_10_411_293_0, i_10_411_316_0, i_10_411_409_0, i_10_411_410_0,
    i_10_411_444_0, i_10_411_800_0, i_10_411_971_0, i_10_411_1036_0,
    i_10_411_1234_0, i_10_411_1237_0, i_10_411_1238_0, i_10_411_1261_0,
    i_10_411_1288_0, i_10_411_1309_0, i_10_411_1359_0, i_10_411_1360_0,
    i_10_411_1361_0, i_10_411_1431_0, i_10_411_1441_0, i_10_411_1442_0,
    i_10_411_1576_0, i_10_411_1578_0, i_10_411_1655_0, i_10_411_1683_0,
    i_10_411_1684_0, i_10_411_1688_0, i_10_411_1690_0, i_10_411_1819_0,
    i_10_411_1949_0, i_10_411_2180_0, i_10_411_2335_0, i_10_411_2351_0,
    i_10_411_2352_0, i_10_411_2363_0, i_10_411_2404_0, i_10_411_2450_0,
    i_10_411_2451_0, i_10_411_2459_0, i_10_411_2462_0, i_10_411_2467_0,
    i_10_411_2504_0, i_10_411_2634_0, i_10_411_2635_0, i_10_411_2656_0,
    i_10_411_2659_0, i_10_411_2663_0, i_10_411_2673_0, i_10_411_2674_0,
    i_10_411_2675_0, i_10_411_2714_0, i_10_411_2785_0, i_10_411_2831_0,
    i_10_411_2918_0, i_10_411_2919_0, i_10_411_2982_0, i_10_411_3151_0,
    i_10_411_3152_0, i_10_411_3153_0, i_10_411_3154_0, i_10_411_3156_0,
    i_10_411_3195_0, i_10_411_3196_0, i_10_411_3198_0, i_10_411_3268_0,
    i_10_411_3269_0, i_10_411_3271_0, i_10_411_3278_0, i_10_411_3292_0,
    i_10_411_3321_0, i_10_411_3522_0, i_10_411_3541_0, i_10_411_3585_0,
    i_10_411_3586_0, i_10_411_3587_0, i_10_411_3612_0, i_10_411_3613_0,
    i_10_411_3615_0, i_10_411_3651_0, i_10_411_3834_0, i_10_411_3848_0,
    i_10_411_3942_0, i_10_411_3944_0, i_10_411_3994_0, i_10_411_4051_0,
    i_10_411_4052_0, i_10_411_4114_0, i_10_411_4116_0, i_10_411_4288_0,
    i_10_411_4289_0, i_10_411_4563_0, i_10_411_4567_0, i_10_411_4594_0,
    o_10_411_0_0  );
  input  i_10_411_145_0, i_10_411_220_0, i_10_411_223_0, i_10_411_271_0,
    i_10_411_272_0, i_10_411_273_0, i_10_411_276_0, i_10_411_283_0,
    i_10_411_293_0, i_10_411_316_0, i_10_411_409_0, i_10_411_410_0,
    i_10_411_444_0, i_10_411_800_0, i_10_411_971_0, i_10_411_1036_0,
    i_10_411_1234_0, i_10_411_1237_0, i_10_411_1238_0, i_10_411_1261_0,
    i_10_411_1288_0, i_10_411_1309_0, i_10_411_1359_0, i_10_411_1360_0,
    i_10_411_1361_0, i_10_411_1431_0, i_10_411_1441_0, i_10_411_1442_0,
    i_10_411_1576_0, i_10_411_1578_0, i_10_411_1655_0, i_10_411_1683_0,
    i_10_411_1684_0, i_10_411_1688_0, i_10_411_1690_0, i_10_411_1819_0,
    i_10_411_1949_0, i_10_411_2180_0, i_10_411_2335_0, i_10_411_2351_0,
    i_10_411_2352_0, i_10_411_2363_0, i_10_411_2404_0, i_10_411_2450_0,
    i_10_411_2451_0, i_10_411_2459_0, i_10_411_2462_0, i_10_411_2467_0,
    i_10_411_2504_0, i_10_411_2634_0, i_10_411_2635_0, i_10_411_2656_0,
    i_10_411_2659_0, i_10_411_2663_0, i_10_411_2673_0, i_10_411_2674_0,
    i_10_411_2675_0, i_10_411_2714_0, i_10_411_2785_0, i_10_411_2831_0,
    i_10_411_2918_0, i_10_411_2919_0, i_10_411_2982_0, i_10_411_3151_0,
    i_10_411_3152_0, i_10_411_3153_0, i_10_411_3154_0, i_10_411_3156_0,
    i_10_411_3195_0, i_10_411_3196_0, i_10_411_3198_0, i_10_411_3268_0,
    i_10_411_3269_0, i_10_411_3271_0, i_10_411_3278_0, i_10_411_3292_0,
    i_10_411_3321_0, i_10_411_3522_0, i_10_411_3541_0, i_10_411_3585_0,
    i_10_411_3586_0, i_10_411_3587_0, i_10_411_3612_0, i_10_411_3613_0,
    i_10_411_3615_0, i_10_411_3651_0, i_10_411_3834_0, i_10_411_3848_0,
    i_10_411_3942_0, i_10_411_3944_0, i_10_411_3994_0, i_10_411_4051_0,
    i_10_411_4052_0, i_10_411_4114_0, i_10_411_4116_0, i_10_411_4288_0,
    i_10_411_4289_0, i_10_411_4563_0, i_10_411_4567_0, i_10_411_4594_0;
  output o_10_411_0_0;
  assign o_10_411_0_0 = ~((~i_10_411_220_0 & ((~i_10_411_316_0 & i_10_411_2635_0 & ~i_10_411_2673_0 & ~i_10_411_3198_0 & ~i_10_411_3834_0 & ~i_10_411_4052_0) | (~i_10_411_283_0 & ~i_10_411_1359_0 & ~i_10_411_2659_0 & ~i_10_411_2675_0 & ~i_10_411_2982_0 & ~i_10_411_3612_0 & ~i_10_411_3615_0 & ~i_10_411_3994_0 & i_10_411_4116_0))) | (~i_10_411_283_0 & ((~i_10_411_145_0 & ~i_10_411_1442_0 & ~i_10_411_2504_0 & ~i_10_411_2656_0 & ~i_10_411_2673_0 & ~i_10_411_2919_0 & ~i_10_411_3271_0 & ~i_10_411_3587_0) | (~i_10_411_1234_0 & ~i_10_411_1683_0 & ~i_10_411_2674_0 & ~i_10_411_3586_0 & ~i_10_411_3615_0 & ~i_10_411_3942_0 & ~i_10_411_4052_0 & ~i_10_411_4114_0))) | (~i_10_411_409_0 & ((i_10_411_2351_0 & ~i_10_411_2404_0 & ~i_10_411_2674_0) | (~i_10_411_1234_0 & ~i_10_411_1309_0 & ~i_10_411_1949_0 & ~i_10_411_2919_0 & ~i_10_411_3587_0 & ~i_10_411_3942_0 & ~i_10_411_4052_0 & ~i_10_411_4116_0))) | (~i_10_411_800_0 & ((~i_10_411_1359_0 & ~i_10_411_1431_0 & ~i_10_411_1442_0 & ~i_10_411_1576_0 & i_10_411_1690_0 & ~i_10_411_1949_0 & ~i_10_411_2656_0 & ~i_10_411_2673_0 & ~i_10_411_3271_0) | (~i_10_411_2504_0 & ~i_10_411_2982_0 & i_10_411_3269_0 & ~i_10_411_4116_0))) | (~i_10_411_1238_0 & ((~i_10_411_1949_0 & ~i_10_411_2656_0 & i_10_411_2785_0 & i_10_411_3651_0 & ~i_10_411_4114_0) | (~i_10_411_1309_0 & ~i_10_411_2673_0 & i_10_411_3848_0 & ~i_10_411_3944_0 & i_10_411_4567_0))) | (~i_10_411_1309_0 & ((~i_10_411_1441_0 & ~i_10_411_3612_0 & i_10_411_3834_0) | (~i_10_411_145_0 & ~i_10_411_316_0 & ~i_10_411_1361_0 & ~i_10_411_2404_0 & ~i_10_411_3585_0 & ~i_10_411_4051_0 & ~i_10_411_4052_0 & ~i_10_411_4567_0))) | (~i_10_411_1576_0 & ((~i_10_411_2180_0 & ~i_10_411_2404_0 & ~i_10_411_2659_0 & ~i_10_411_2673_0 & ~i_10_411_2675_0 & ~i_10_411_3271_0 & ~i_10_411_3612_0) | (~i_10_411_223_0 & i_10_411_2635_0 & ~i_10_411_3587_0 & ~i_10_411_4051_0))) | (i_10_411_2634_0 & ((~i_10_411_2467_0 & ~i_10_411_2674_0 & ~i_10_411_3587_0 & ~i_10_411_4116_0) | (~i_10_411_2675_0 & i_10_411_4289_0))) | (~i_10_411_2674_0 & ((~i_10_411_4052_0 & ((~i_10_411_145_0 & ~i_10_411_2673_0 & ((~i_10_411_1359_0 & ~i_10_411_2675_0 & ~i_10_411_2785_0 & ~i_10_411_3522_0 & ~i_10_411_3586_0 & ~i_10_411_3615_0) | (~i_10_411_1441_0 & ~i_10_411_2467_0 & ~i_10_411_2504_0 & i_10_411_2656_0 & ~i_10_411_3271_0 & ~i_10_411_3278_0 & ~i_10_411_3994_0 & ~i_10_411_4563_0))) | (i_10_411_2635_0 & ~i_10_411_3522_0 & ~i_10_411_3613_0) | (~i_10_411_410_0 & ~i_10_411_2656_0 & ~i_10_411_3585_0 & i_10_411_3586_0 & ~i_10_411_3848_0 & ~i_10_411_3944_0))) | (~i_10_411_2656_0 & ((~i_10_411_2467_0 & ~i_10_411_2982_0 & i_10_411_3271_0 & ~i_10_411_3615_0 & i_10_411_4567_0) | (~i_10_411_2363_0 & ~i_10_411_2451_0 & i_10_411_2659_0 & ~i_10_411_2675_0 & ~i_10_411_3196_0 & ~i_10_411_3198_0 & ~i_10_411_4563_0 & ~i_10_411_4567_0))) | (i_10_411_2635_0 & ~i_10_411_3586_0 & ~i_10_411_4563_0) | (~i_10_411_1361_0 & ~i_10_411_2450_0 & ~i_10_411_2504_0 & ~i_10_411_2663_0 & ~i_10_411_2673_0 & ~i_10_411_2831_0 & i_10_411_3586_0 & ~i_10_411_4051_0 & ~i_10_411_4567_0))) | (~i_10_411_2656_0 & ((i_10_411_1576_0 & ~i_10_411_2504_0 & ~i_10_411_2673_0 & ~i_10_411_2982_0) | (~i_10_411_4116_0 & i_10_411_4288_0 & i_10_411_4567_0))) | (~i_10_411_2659_0 & ((i_10_411_2352_0 & ~i_10_411_3522_0 & ~i_10_411_3613_0) | (~i_10_411_1442_0 & ~i_10_411_2673_0 & ~i_10_411_3615_0 & i_10_411_4563_0))) | (i_10_411_2714_0 & i_10_411_2831_0 & (~i_10_411_3587_0 | (~i_10_411_3994_0 & ~i_10_411_4567_0))) | (~i_10_411_3522_0 & ~i_10_411_4051_0 & ((i_10_411_1238_0 & ~i_10_411_2675_0 & i_10_411_2785_0 & ~i_10_411_3613_0) | (~i_10_411_2673_0 & i_10_411_3195_0 & ~i_10_411_4052_0))) | (~i_10_411_2673_0 & ((i_10_411_1655_0 & ~i_10_411_1684_0 & ~i_10_411_2467_0 & i_10_411_2674_0 & i_10_411_3278_0) | (~i_10_411_145_0 & ~i_10_411_444_0 & ~i_10_411_1261_0 & ~i_10_411_2404_0 & ~i_10_411_2663_0 & ~i_10_411_2675_0 & ~i_10_411_3942_0 & ~i_10_411_3944_0 & ~i_10_411_4052_0 & ~i_10_411_4116_0 & ~i_10_411_4567_0))) | (~i_10_411_3587_0 & ~i_10_411_3942_0 & i_10_411_2450_0 & ~i_10_411_2675_0) | (i_10_411_2462_0 & ~i_10_411_4114_0) | (i_10_411_2351_0 & i_10_411_3848_0 & ~i_10_411_4563_0 & i_10_411_4567_0));
endmodule



// Benchmark "kernel_10_412" written by ABC on Sun Jul 19 10:28:14 2020

module kernel_10_412 ( 
    i_10_412_121_0, i_10_412_125_0, i_10_412_176_0, i_10_412_220_0,
    i_10_412_247_0, i_10_412_285_0, i_10_412_319_0, i_10_412_408_0,
    i_10_412_409_0, i_10_412_410_0, i_10_412_448_0, i_10_412_565_0,
    i_10_412_955_0, i_10_412_958_0, i_10_412_960_0, i_10_412_962_0,
    i_10_412_1006_0, i_10_412_1007_0, i_10_412_1083_0, i_10_412_1136_0,
    i_10_412_1137_0, i_10_412_1138_0, i_10_412_1181_0, i_10_412_1237_0,
    i_10_412_1308_0, i_10_412_1541_0, i_10_412_1544_0, i_10_412_1552_0,
    i_10_412_1553_0, i_10_412_1575_0, i_10_412_1618_0, i_10_412_1652_0,
    i_10_412_1677_0, i_10_412_1684_0, i_10_412_1687_0, i_10_412_1819_0,
    i_10_412_1951_0, i_10_412_1952_0, i_10_412_2182_0, i_10_412_2184_0,
    i_10_412_2185_0, i_10_412_2186_0, i_10_412_2200_0, i_10_412_2312_0,
    i_10_412_2330_0, i_10_412_2349_0, i_10_412_2353_0, i_10_412_2355_0,
    i_10_412_2361_0, i_10_412_2366_0, i_10_412_2405_0, i_10_412_2411_0,
    i_10_412_2461_0, i_10_412_2470_0, i_10_412_2471_0, i_10_412_2473_0,
    i_10_412_2509_0, i_10_412_2510_0, i_10_412_2632_0, i_10_412_2633_0,
    i_10_412_2681_0, i_10_412_2716_0, i_10_412_2729_0, i_10_412_2833_0,
    i_10_412_2880_0, i_10_412_2881_0, i_10_412_2884_0, i_10_412_2885_0,
    i_10_412_2920_0, i_10_412_2921_0, i_10_412_2924_0, i_10_412_3038_0,
    i_10_412_3151_0, i_10_412_3199_0, i_10_412_3200_0, i_10_412_3203_0,
    i_10_412_3271_0, i_10_412_3275_0, i_10_412_3316_0, i_10_412_3323_0,
    i_10_412_3325_0, i_10_412_3326_0, i_10_412_3328_0, i_10_412_3329_0,
    i_10_412_3497_0, i_10_412_3585_0, i_10_412_3586_0, i_10_412_3617_0,
    i_10_412_3649_0, i_10_412_3653_0, i_10_412_3686_0, i_10_412_3782_0,
    i_10_412_3785_0, i_10_412_3787_0, i_10_412_3834_0, i_10_412_3838_0,
    i_10_412_3856_0, i_10_412_3983_0, i_10_412_4058_0, i_10_412_4567_0,
    o_10_412_0_0  );
  input  i_10_412_121_0, i_10_412_125_0, i_10_412_176_0, i_10_412_220_0,
    i_10_412_247_0, i_10_412_285_0, i_10_412_319_0, i_10_412_408_0,
    i_10_412_409_0, i_10_412_410_0, i_10_412_448_0, i_10_412_565_0,
    i_10_412_955_0, i_10_412_958_0, i_10_412_960_0, i_10_412_962_0,
    i_10_412_1006_0, i_10_412_1007_0, i_10_412_1083_0, i_10_412_1136_0,
    i_10_412_1137_0, i_10_412_1138_0, i_10_412_1181_0, i_10_412_1237_0,
    i_10_412_1308_0, i_10_412_1541_0, i_10_412_1544_0, i_10_412_1552_0,
    i_10_412_1553_0, i_10_412_1575_0, i_10_412_1618_0, i_10_412_1652_0,
    i_10_412_1677_0, i_10_412_1684_0, i_10_412_1687_0, i_10_412_1819_0,
    i_10_412_1951_0, i_10_412_1952_0, i_10_412_2182_0, i_10_412_2184_0,
    i_10_412_2185_0, i_10_412_2186_0, i_10_412_2200_0, i_10_412_2312_0,
    i_10_412_2330_0, i_10_412_2349_0, i_10_412_2353_0, i_10_412_2355_0,
    i_10_412_2361_0, i_10_412_2366_0, i_10_412_2405_0, i_10_412_2411_0,
    i_10_412_2461_0, i_10_412_2470_0, i_10_412_2471_0, i_10_412_2473_0,
    i_10_412_2509_0, i_10_412_2510_0, i_10_412_2632_0, i_10_412_2633_0,
    i_10_412_2681_0, i_10_412_2716_0, i_10_412_2729_0, i_10_412_2833_0,
    i_10_412_2880_0, i_10_412_2881_0, i_10_412_2884_0, i_10_412_2885_0,
    i_10_412_2920_0, i_10_412_2921_0, i_10_412_2924_0, i_10_412_3038_0,
    i_10_412_3151_0, i_10_412_3199_0, i_10_412_3200_0, i_10_412_3203_0,
    i_10_412_3271_0, i_10_412_3275_0, i_10_412_3316_0, i_10_412_3323_0,
    i_10_412_3325_0, i_10_412_3326_0, i_10_412_3328_0, i_10_412_3329_0,
    i_10_412_3497_0, i_10_412_3585_0, i_10_412_3586_0, i_10_412_3617_0,
    i_10_412_3649_0, i_10_412_3653_0, i_10_412_3686_0, i_10_412_3782_0,
    i_10_412_3785_0, i_10_412_3787_0, i_10_412_3834_0, i_10_412_3838_0,
    i_10_412_3856_0, i_10_412_3983_0, i_10_412_4058_0, i_10_412_4567_0;
  output o_10_412_0_0;
  assign o_10_412_0_0 = ~((~i_10_412_2186_0 & ((~i_10_412_960_0 & ((~i_10_412_1006_0 & ~i_10_412_1541_0 & ~i_10_412_1553_0 & ~i_10_412_1684_0 & ~i_10_412_2355_0 & ~i_10_412_2471_0 & ~i_10_412_2881_0 & ~i_10_412_3203_0) | (~i_10_412_1544_0 & ~i_10_412_1819_0 & ~i_10_412_2330_0 & ~i_10_412_2349_0 & ~i_10_412_3271_0 & i_10_412_3617_0 & ~i_10_412_3983_0))) | (~i_10_412_3275_0 & ((~i_10_412_1006_0 & ((~i_10_412_176_0 & ~i_10_412_409_0 & ~i_10_412_1007_0 & ~i_10_412_1083_0 & ~i_10_412_2182_0 & ~i_10_412_2185_0 & i_10_412_2632_0 & ~i_10_412_2881_0 & ~i_10_412_2920_0) | (~i_10_412_962_0 & ~i_10_412_1575_0 & ~i_10_412_1951_0 & i_10_412_2349_0 & ~i_10_412_3617_0 & ~i_10_412_3834_0))) | (~i_10_412_1544_0 & ~i_10_412_2461_0 & ((~i_10_412_1553_0 & ~i_10_412_2184_0 & ~i_10_412_2312_0 & ~i_10_412_3200_0) | (~i_10_412_2182_0 & ~i_10_412_2185_0 & ~i_10_412_2355_0 & ~i_10_412_3983_0))) | (i_10_412_1652_0 & i_10_412_1819_0 & ~i_10_412_2353_0 & ~i_10_412_2366_0 & ~i_10_412_2729_0))) | (~i_10_412_2185_0 & ~i_10_412_2355_0 & ((~i_10_412_247_0 & ~i_10_412_2312_0 & ~i_10_412_2330_0 & ~i_10_412_3649_0) | (i_10_412_2924_0 & ~i_10_412_3038_0 & ~i_10_412_3653_0))) | (~i_10_412_3271_0 & ((~i_10_412_1006_0 & i_10_412_1308_0 & ~i_10_412_1552_0 & ~i_10_412_3203_0 & ~i_10_412_3785_0) | (~i_10_412_410_0 & ~i_10_412_958_0 & ~i_10_412_2510_0 & ~i_10_412_2729_0 & ~i_10_412_2885_0 & ~i_10_412_3316_0 & ~i_10_412_3983_0 & ~i_10_412_4058_0))) | (~i_10_412_1308_0 & ~i_10_412_2411_0 & ~i_10_412_2461_0 & i_10_412_2471_0 & ~i_10_412_3782_0))) | (~i_10_412_958_0 & ((~i_10_412_2182_0 & ~i_10_412_2411_0 & ~i_10_412_2632_0 & i_10_412_3271_0 & ~i_10_412_3649_0) | (~i_10_412_1819_0 & i_10_412_3617_0 & ~i_10_412_3838_0 & ~i_10_412_3983_0))) | (~i_10_412_2185_0 & ((~i_10_412_962_0 & ((~i_10_412_565_0 & ~i_10_412_1544_0 & ~i_10_412_1952_0 & ~i_10_412_2405_0 & ~i_10_412_2729_0 & ~i_10_412_2885_0 & ~i_10_412_3038_0 & ~i_10_412_3838_0) | (~i_10_412_2330_0 & ~i_10_412_3275_0 & ~i_10_412_3649_0 & ~i_10_412_4058_0))) | (~i_10_412_1952_0 & ~i_10_412_2312_0 & ~i_10_412_2366_0 & ~i_10_412_2633_0 & ~i_10_412_3686_0 & ~i_10_412_3787_0))) | (~i_10_412_448_0 & ~i_10_412_2312_0 & i_10_412_2470_0 & ~i_10_412_2510_0 & ~i_10_412_2729_0) | (i_10_412_2880_0 & i_10_412_3275_0) | (i_10_412_1575_0 & ~i_10_412_2632_0 & ~i_10_412_3038_0 & i_10_412_3787_0 & i_10_412_3856_0));
endmodule



// Benchmark "kernel_10_413" written by ABC on Sun Jul 19 10:28:15 2020

module kernel_10_413 ( 
    i_10_413_283_0, i_10_413_296_0, i_10_413_321_0, i_10_413_327_0,
    i_10_413_328_0, i_10_413_329_0, i_10_413_330_0, i_10_413_411_0,
    i_10_413_436_0, i_10_413_459_0, i_10_413_461_0, i_10_413_463_0,
    i_10_413_464_0, i_10_413_749_0, i_10_413_793_0, i_10_413_901_0,
    i_10_413_969_0, i_10_413_1080_0, i_10_413_1083_0, i_10_413_1084_0,
    i_10_413_1217_0, i_10_413_1233_0, i_10_413_1261_0, i_10_413_1263_0,
    i_10_413_1264_0, i_10_413_1277_0, i_10_413_1310_0, i_10_413_1359_0,
    i_10_413_1432_0, i_10_413_1433_0, i_10_413_1638_0, i_10_413_1649_0,
    i_10_413_1655_0, i_10_413_1772_0, i_10_413_1818_0, i_10_413_1822_0,
    i_10_413_1909_0, i_10_413_1912_0, i_10_413_1913_0, i_10_413_2198_0,
    i_10_413_2351_0, i_10_413_2353_0, i_10_413_2357_0, i_10_413_2361_0,
    i_10_413_2379_0, i_10_413_2453_0, i_10_413_2466_0, i_10_413_2467_0,
    i_10_413_2504_0, i_10_413_2629_0, i_10_413_2630_0, i_10_413_2656_0,
    i_10_413_2660_0, i_10_413_2702_0, i_10_413_2705_0, i_10_413_2715_0,
    i_10_413_2717_0, i_10_413_2735_0, i_10_413_2826_0, i_10_413_2827_0,
    i_10_413_2828_0, i_10_413_2877_0, i_10_413_2917_0, i_10_413_2921_0,
    i_10_413_2979_0, i_10_413_2980_0, i_10_413_2981_0, i_10_413_3036_0,
    i_10_413_3040_0, i_10_413_3077_0, i_10_413_3278_0, i_10_413_3326_0,
    i_10_413_3329_0, i_10_413_3384_0, i_10_413_3403_0, i_10_413_3433_0,
    i_10_413_3523_0, i_10_413_3526_0, i_10_413_3611_0, i_10_413_3615_0,
    i_10_413_3646_0, i_10_413_3647_0, i_10_413_3648_0, i_10_413_3650_0,
    i_10_413_3682_0, i_10_413_3719_0, i_10_413_3837_0, i_10_413_3853_0,
    i_10_413_3856_0, i_10_413_3888_0, i_10_413_3889_0, i_10_413_3890_0,
    i_10_413_3987_0, i_10_413_3991_0, i_10_413_4027_0, i_10_413_4124_0,
    i_10_413_4208_0, i_10_413_4211_0, i_10_413_4276_0, i_10_413_4291_0,
    o_10_413_0_0  );
  input  i_10_413_283_0, i_10_413_296_0, i_10_413_321_0, i_10_413_327_0,
    i_10_413_328_0, i_10_413_329_0, i_10_413_330_0, i_10_413_411_0,
    i_10_413_436_0, i_10_413_459_0, i_10_413_461_0, i_10_413_463_0,
    i_10_413_464_0, i_10_413_749_0, i_10_413_793_0, i_10_413_901_0,
    i_10_413_969_0, i_10_413_1080_0, i_10_413_1083_0, i_10_413_1084_0,
    i_10_413_1217_0, i_10_413_1233_0, i_10_413_1261_0, i_10_413_1263_0,
    i_10_413_1264_0, i_10_413_1277_0, i_10_413_1310_0, i_10_413_1359_0,
    i_10_413_1432_0, i_10_413_1433_0, i_10_413_1638_0, i_10_413_1649_0,
    i_10_413_1655_0, i_10_413_1772_0, i_10_413_1818_0, i_10_413_1822_0,
    i_10_413_1909_0, i_10_413_1912_0, i_10_413_1913_0, i_10_413_2198_0,
    i_10_413_2351_0, i_10_413_2353_0, i_10_413_2357_0, i_10_413_2361_0,
    i_10_413_2379_0, i_10_413_2453_0, i_10_413_2466_0, i_10_413_2467_0,
    i_10_413_2504_0, i_10_413_2629_0, i_10_413_2630_0, i_10_413_2656_0,
    i_10_413_2660_0, i_10_413_2702_0, i_10_413_2705_0, i_10_413_2715_0,
    i_10_413_2717_0, i_10_413_2735_0, i_10_413_2826_0, i_10_413_2827_0,
    i_10_413_2828_0, i_10_413_2877_0, i_10_413_2917_0, i_10_413_2921_0,
    i_10_413_2979_0, i_10_413_2980_0, i_10_413_2981_0, i_10_413_3036_0,
    i_10_413_3040_0, i_10_413_3077_0, i_10_413_3278_0, i_10_413_3326_0,
    i_10_413_3329_0, i_10_413_3384_0, i_10_413_3403_0, i_10_413_3433_0,
    i_10_413_3523_0, i_10_413_3526_0, i_10_413_3611_0, i_10_413_3615_0,
    i_10_413_3646_0, i_10_413_3647_0, i_10_413_3648_0, i_10_413_3650_0,
    i_10_413_3682_0, i_10_413_3719_0, i_10_413_3837_0, i_10_413_3853_0,
    i_10_413_3856_0, i_10_413_3888_0, i_10_413_3889_0, i_10_413_3890_0,
    i_10_413_3987_0, i_10_413_3991_0, i_10_413_4027_0, i_10_413_4124_0,
    i_10_413_4208_0, i_10_413_4211_0, i_10_413_4276_0, i_10_413_4291_0;
  output o_10_413_0_0;
  assign o_10_413_0_0 = 0;
endmodule



// Benchmark "kernel_10_414" written by ABC on Sun Jul 19 10:28:17 2020

module kernel_10_414 ( 
    i_10_414_172_0, i_10_414_174_0, i_10_414_175_0, i_10_414_216_0,
    i_10_414_220_0, i_10_414_221_0, i_10_414_224_0, i_10_414_279_0,
    i_10_414_315_0, i_10_414_317_0, i_10_414_387_0, i_10_414_411_0,
    i_10_414_446_0, i_10_414_459_0, i_10_414_461_0, i_10_414_712_0,
    i_10_414_797_0, i_10_414_898_0, i_10_414_962_0, i_10_414_1000_0,
    i_10_414_1003_0, i_10_414_1237_0, i_10_414_1238_0, i_10_414_1310_0,
    i_10_414_1312_0, i_10_414_1431_0, i_10_414_1432_0, i_10_414_1433_0,
    i_10_414_1576_0, i_10_414_1577_0, i_10_414_1580_0, i_10_414_1581_0,
    i_10_414_1651_0, i_10_414_1683_0, i_10_414_1686_0, i_10_414_1820_0,
    i_10_414_1822_0, i_10_414_1913_0, i_10_414_2186_0, i_10_414_2197_0,
    i_10_414_2349_0, i_10_414_2350_0, i_10_414_2356_0, i_10_414_2358_0,
    i_10_414_2410_0, i_10_414_2452_0, i_10_414_2453_0, i_10_414_2460_0,
    i_10_414_2468_0, i_10_414_2502_0, i_10_414_2661_0, i_10_414_2700_0,
    i_10_414_2701_0, i_10_414_2713_0, i_10_414_2714_0, i_10_414_2716_0,
    i_10_414_2717_0, i_10_414_2719_0, i_10_414_2721_0, i_10_414_2722_0,
    i_10_414_2723_0, i_10_414_2885_0, i_10_414_2924_0, i_10_414_3036_0,
    i_10_414_3050_0, i_10_414_3069_0, i_10_414_3070_0, i_10_414_3280_0,
    i_10_414_3384_0, i_10_414_3385_0, i_10_414_3390_0, i_10_414_3391_0,
    i_10_414_3403_0, i_10_414_3405_0, i_10_414_3406_0, i_10_414_3409_0,
    i_10_414_3523_0, i_10_414_3613_0, i_10_414_3647_0, i_10_414_3648_0,
    i_10_414_3651_0, i_10_414_3785_0, i_10_414_3855_0, i_10_414_3856_0,
    i_10_414_3857_0, i_10_414_3860_0, i_10_414_3978_0, i_10_414_3980_0,
    i_10_414_3982_0, i_10_414_3983_0, i_10_414_4029_0, i_10_414_4117_0,
    i_10_414_4118_0, i_10_414_4169_0, i_10_414_4284_0, i_10_414_4285_0,
    i_10_414_4288_0, i_10_414_4290_0, i_10_414_4565_0, i_10_414_4567_0,
    o_10_414_0_0  );
  input  i_10_414_172_0, i_10_414_174_0, i_10_414_175_0, i_10_414_216_0,
    i_10_414_220_0, i_10_414_221_0, i_10_414_224_0, i_10_414_279_0,
    i_10_414_315_0, i_10_414_317_0, i_10_414_387_0, i_10_414_411_0,
    i_10_414_446_0, i_10_414_459_0, i_10_414_461_0, i_10_414_712_0,
    i_10_414_797_0, i_10_414_898_0, i_10_414_962_0, i_10_414_1000_0,
    i_10_414_1003_0, i_10_414_1237_0, i_10_414_1238_0, i_10_414_1310_0,
    i_10_414_1312_0, i_10_414_1431_0, i_10_414_1432_0, i_10_414_1433_0,
    i_10_414_1576_0, i_10_414_1577_0, i_10_414_1580_0, i_10_414_1581_0,
    i_10_414_1651_0, i_10_414_1683_0, i_10_414_1686_0, i_10_414_1820_0,
    i_10_414_1822_0, i_10_414_1913_0, i_10_414_2186_0, i_10_414_2197_0,
    i_10_414_2349_0, i_10_414_2350_0, i_10_414_2356_0, i_10_414_2358_0,
    i_10_414_2410_0, i_10_414_2452_0, i_10_414_2453_0, i_10_414_2460_0,
    i_10_414_2468_0, i_10_414_2502_0, i_10_414_2661_0, i_10_414_2700_0,
    i_10_414_2701_0, i_10_414_2713_0, i_10_414_2714_0, i_10_414_2716_0,
    i_10_414_2717_0, i_10_414_2719_0, i_10_414_2721_0, i_10_414_2722_0,
    i_10_414_2723_0, i_10_414_2885_0, i_10_414_2924_0, i_10_414_3036_0,
    i_10_414_3050_0, i_10_414_3069_0, i_10_414_3070_0, i_10_414_3280_0,
    i_10_414_3384_0, i_10_414_3385_0, i_10_414_3390_0, i_10_414_3391_0,
    i_10_414_3403_0, i_10_414_3405_0, i_10_414_3406_0, i_10_414_3409_0,
    i_10_414_3523_0, i_10_414_3613_0, i_10_414_3647_0, i_10_414_3648_0,
    i_10_414_3651_0, i_10_414_3785_0, i_10_414_3855_0, i_10_414_3856_0,
    i_10_414_3857_0, i_10_414_3860_0, i_10_414_3978_0, i_10_414_3980_0,
    i_10_414_3982_0, i_10_414_3983_0, i_10_414_4029_0, i_10_414_4117_0,
    i_10_414_4118_0, i_10_414_4169_0, i_10_414_4284_0, i_10_414_4285_0,
    i_10_414_4288_0, i_10_414_4290_0, i_10_414_4565_0, i_10_414_4567_0;
  output o_10_414_0_0;
  assign o_10_414_0_0 = ~((~i_10_414_2723_0 & ((i_10_414_174_0 & ((~i_10_414_3856_0 & i_10_414_4117_0 & ~i_10_414_4284_0 & ~i_10_414_4288_0) | (~i_10_414_224_0 & i_10_414_1822_0 & ~i_10_414_2661_0 & ~i_10_414_3050_0 & ~i_10_414_3385_0 & ~i_10_414_3613_0 & i_10_414_4290_0))) | (i_10_414_1822_0 & ((~i_10_414_2716_0 & ~i_10_414_2924_0 & ~i_10_414_3280_0 & ~i_10_414_3385_0 & ~i_10_414_3391_0) | (~i_10_414_712_0 & ~i_10_414_898_0 & ~i_10_414_1238_0 & ~i_10_414_1683_0 & ~i_10_414_2460_0 & ~i_10_414_3036_0 & ~i_10_414_3390_0 & ~i_10_414_3978_0))) | (~i_10_414_898_0 & ((~i_10_414_2717_0 & ~i_10_414_2721_0 & ~i_10_414_2722_0 & ~i_10_414_3280_0) | (~i_10_414_446_0 & ~i_10_414_1310_0 & ~i_10_414_1312_0 & ~i_10_414_2661_0 & ~i_10_414_3036_0 & ~i_10_414_3406_0 & ~i_10_414_3613_0 & ~i_10_414_3856_0 & ~i_10_414_4565_0))) | (~i_10_414_2661_0 & ((i_10_414_2358_0 & ~i_10_414_3391_0 & ~i_10_414_3406_0 & ~i_10_414_4290_0) | (~i_10_414_2713_0 & i_10_414_3855_0 & i_10_414_3857_0 & i_10_414_4567_0))) | (i_10_414_317_0 & ~i_10_414_2716_0) | (~i_10_414_174_0 & i_10_414_446_0 & ~i_10_414_2350_0 & ~i_10_414_3280_0 & ~i_10_414_3406_0))) | (~i_10_414_4290_0 & ((~i_10_414_174_0 & ((~i_10_414_797_0 & ~i_10_414_898_0 & ~i_10_414_2349_0 & ~i_10_414_2713_0 & ~i_10_414_4284_0 & ~i_10_414_4288_0 & ~i_10_414_2717_0 & ~i_10_414_3406_0) | (~i_10_414_1310_0 & i_10_414_2356_0 & ~i_10_414_2460_0 & ~i_10_414_3523_0 & ~i_10_414_4117_0 & i_10_414_4567_0))) | (~i_10_414_220_0 & ~i_10_414_898_0 & ~i_10_414_1686_0 & ~i_10_414_1822_0 & ~i_10_414_3280_0 & ~i_10_414_3406_0 & ~i_10_414_3857_0 & ~i_10_414_3983_0) | (~i_10_414_461_0 & ~i_10_414_1683_0 & ~i_10_414_2452_0 & ~i_10_414_2714_0 & ~i_10_414_3391_0 & ~i_10_414_3409_0 & ~i_10_414_4567_0))) | (~i_10_414_216_0 & ((~i_10_414_221_0 & ~i_10_414_797_0 & i_10_414_1820_0) | (~i_10_414_461_0 & i_10_414_2350_0 & ~i_10_414_2716_0 & ~i_10_414_3391_0 & ~i_10_414_4285_0))) | (~i_10_414_459_0 & ((~i_10_414_224_0 & i_10_414_315_0 & ~i_10_414_898_0 & ~i_10_414_3406_0) | (~i_10_414_2453_0 & i_10_414_2713_0 & i_10_414_2719_0 & ~i_10_414_2722_0 & ~i_10_414_3856_0 & ~i_10_414_4567_0))) | (~i_10_414_461_0 & ((~i_10_414_2716_0 & i_10_414_3983_0 & ~i_10_414_4118_0 & ~i_10_414_4285_0) | (~i_10_414_712_0 & ~i_10_414_1310_0 & ~i_10_414_1651_0 & ~i_10_414_1820_0 & ~i_10_414_2349_0 & ~i_10_414_3050_0 & ~i_10_414_3391_0 & ~i_10_414_3785_0 & ~i_10_414_3982_0 & ~i_10_414_3983_0 & ~i_10_414_4567_0))) | (~i_10_414_1312_0 & ~i_10_414_3523_0 & ((~i_10_414_1820_0 & ~i_10_414_2716_0 & ~i_10_414_2719_0 & ~i_10_414_2722_0 & ~i_10_414_2924_0 & ~i_10_414_3050_0) | (~i_10_414_1822_0 & ~i_10_414_2410_0 & ~i_10_414_2717_0 & ~i_10_414_3403_0 & ~i_10_414_3856_0 & ~i_10_414_4284_0))) | (~i_10_414_2468_0 & ~i_10_414_2713_0 & ((~i_10_414_220_0 & ~i_10_414_1913_0 & ~i_10_414_2717_0 & ~i_10_414_3050_0 & ~i_10_414_3280_0 & ~i_10_414_3855_0) | (~i_10_414_898_0 & ~i_10_414_1237_0 & ~i_10_414_1238_0 & ~i_10_414_2714_0 & ~i_10_414_2716_0 & ~i_10_414_4285_0))) | (~i_10_414_1237_0 & ((~i_10_414_1238_0 & ((~i_10_414_2452_0 & ~i_10_414_2716_0 & ~i_10_414_3050_0 & ~i_10_414_3385_0 & i_10_414_3391_0 & ~i_10_414_3405_0) | (i_10_414_224_0 & ~i_10_414_2714_0 & ~i_10_414_4029_0 & i_10_414_4567_0))) | (~i_10_414_712_0 & ~i_10_414_2349_0 & ~i_10_414_2719_0 & ~i_10_414_3280_0 & ~i_10_414_3648_0 & ~i_10_414_3855_0 & i_10_414_4565_0))) | (~i_10_414_1822_0 & ~i_10_414_2721_0 & i_10_414_3978_0));
endmodule



// Benchmark "kernel_10_415" written by ABC on Sun Jul 19 10:28:17 2020

module kernel_10_415 ( 
    i_10_415_148_0, i_10_415_222_0, i_10_415_247_0, i_10_415_258_0,
    i_10_415_259_0, i_10_415_279_0, i_10_415_282_0, i_10_415_436_0,
    i_10_415_442_0, i_10_415_463_0, i_10_415_464_0, i_10_415_566_0,
    i_10_415_589_0, i_10_415_694_0, i_10_415_718_0, i_10_415_735_0,
    i_10_415_736_0, i_10_415_752_0, i_10_415_792_0, i_10_415_797_0,
    i_10_415_957_0, i_10_415_1029_0, i_10_415_1031_0, i_10_415_1033_0,
    i_10_415_1050_0, i_10_415_1051_0, i_10_415_1052_0, i_10_415_1159_0,
    i_10_415_1160_0, i_10_415_1262_0, i_10_415_1310_0, i_10_415_1311_0,
    i_10_415_1439_0, i_10_415_1443_0, i_10_415_1454_0, i_10_415_1546_0,
    i_10_415_1613_0, i_10_415_1633_0, i_10_415_1634_0, i_10_415_1635_0,
    i_10_415_1636_0, i_10_415_1637_0, i_10_415_1651_0, i_10_415_1652_0,
    i_10_415_1684_0, i_10_415_1688_0, i_10_415_1821_0, i_10_415_1912_0,
    i_10_415_1914_0, i_10_415_1939_0, i_10_415_2002_0, i_10_415_2150_0,
    i_10_415_2181_0, i_10_415_2185_0, i_10_415_2186_0, i_10_415_2366_0,
    i_10_415_2433_0, i_10_415_2435_0, i_10_415_2679_0, i_10_415_2680_0,
    i_10_415_2714_0, i_10_415_2717_0, i_10_415_2725_0, i_10_415_2733_0,
    i_10_415_2829_0, i_10_415_2831_0, i_10_415_2884_0, i_10_415_2888_0,
    i_10_415_3093_0, i_10_415_3094_0, i_10_415_3095_0, i_10_415_3199_0,
    i_10_415_3201_0, i_10_415_3236_0, i_10_415_3271_0, i_10_415_3503_0,
    i_10_415_3562_0, i_10_415_3586_0, i_10_415_3587_0, i_10_415_3588_0,
    i_10_415_3617_0, i_10_415_3653_0, i_10_415_3721_0, i_10_415_3781_0,
    i_10_415_3784_0, i_10_415_3787_0, i_10_415_3838_0, i_10_415_3943_0,
    i_10_415_3944_0, i_10_415_3945_0, i_10_415_3981_0, i_10_415_3983_0,
    i_10_415_3985_0, i_10_415_4031_0, i_10_415_4117_0, i_10_415_4121_0,
    i_10_415_4183_0, i_10_415_4226_0, i_10_415_4270_0, i_10_415_4375_0,
    o_10_415_0_0  );
  input  i_10_415_148_0, i_10_415_222_0, i_10_415_247_0, i_10_415_258_0,
    i_10_415_259_0, i_10_415_279_0, i_10_415_282_0, i_10_415_436_0,
    i_10_415_442_0, i_10_415_463_0, i_10_415_464_0, i_10_415_566_0,
    i_10_415_589_0, i_10_415_694_0, i_10_415_718_0, i_10_415_735_0,
    i_10_415_736_0, i_10_415_752_0, i_10_415_792_0, i_10_415_797_0,
    i_10_415_957_0, i_10_415_1029_0, i_10_415_1031_0, i_10_415_1033_0,
    i_10_415_1050_0, i_10_415_1051_0, i_10_415_1052_0, i_10_415_1159_0,
    i_10_415_1160_0, i_10_415_1262_0, i_10_415_1310_0, i_10_415_1311_0,
    i_10_415_1439_0, i_10_415_1443_0, i_10_415_1454_0, i_10_415_1546_0,
    i_10_415_1613_0, i_10_415_1633_0, i_10_415_1634_0, i_10_415_1635_0,
    i_10_415_1636_0, i_10_415_1637_0, i_10_415_1651_0, i_10_415_1652_0,
    i_10_415_1684_0, i_10_415_1688_0, i_10_415_1821_0, i_10_415_1912_0,
    i_10_415_1914_0, i_10_415_1939_0, i_10_415_2002_0, i_10_415_2150_0,
    i_10_415_2181_0, i_10_415_2185_0, i_10_415_2186_0, i_10_415_2366_0,
    i_10_415_2433_0, i_10_415_2435_0, i_10_415_2679_0, i_10_415_2680_0,
    i_10_415_2714_0, i_10_415_2717_0, i_10_415_2725_0, i_10_415_2733_0,
    i_10_415_2829_0, i_10_415_2831_0, i_10_415_2884_0, i_10_415_2888_0,
    i_10_415_3093_0, i_10_415_3094_0, i_10_415_3095_0, i_10_415_3199_0,
    i_10_415_3201_0, i_10_415_3236_0, i_10_415_3271_0, i_10_415_3503_0,
    i_10_415_3562_0, i_10_415_3586_0, i_10_415_3587_0, i_10_415_3588_0,
    i_10_415_3617_0, i_10_415_3653_0, i_10_415_3721_0, i_10_415_3781_0,
    i_10_415_3784_0, i_10_415_3787_0, i_10_415_3838_0, i_10_415_3943_0,
    i_10_415_3944_0, i_10_415_3945_0, i_10_415_3981_0, i_10_415_3983_0,
    i_10_415_3985_0, i_10_415_4031_0, i_10_415_4117_0, i_10_415_4121_0,
    i_10_415_4183_0, i_10_415_4226_0, i_10_415_4270_0, i_10_415_4375_0;
  output o_10_415_0_0;
  assign o_10_415_0_0 = 0;
endmodule



// Benchmark "kernel_10_416" written by ABC on Sun Jul 19 10:28:18 2020

module kernel_10_416 ( 
    i_10_416_144_0, i_10_416_174_0, i_10_416_216_0, i_10_416_236_0,
    i_10_416_279_0, i_10_416_426_0, i_10_416_433_0, i_10_416_435_0,
    i_10_416_441_0, i_10_416_442_0, i_10_416_443_0, i_10_416_444_0,
    i_10_416_446_0, i_10_416_463_0, i_10_416_515_0, i_10_416_518_0,
    i_10_416_792_0, i_10_416_793_0, i_10_416_794_0, i_10_416_820_0,
    i_10_416_892_0, i_10_416_957_0, i_10_416_967_0, i_10_416_1083_0,
    i_10_416_1084_0, i_10_416_1202_0, i_10_416_1360_0, i_10_416_1377_0,
    i_10_416_1485_0, i_10_416_1546_0, i_10_416_1576_0, i_10_416_1581_0,
    i_10_416_1631_0, i_10_416_1691_0, i_10_416_1728_0, i_10_416_1818_0,
    i_10_416_1820_0, i_10_416_1954_0, i_10_416_2045_0, i_10_416_2200_0,
    i_10_416_2202_0, i_10_416_2225_0, i_10_416_2288_0, i_10_416_2331_0,
    i_10_416_2352_0, i_10_416_2357_0, i_10_416_2358_0, i_10_416_2360_0,
    i_10_416_2377_0, i_10_416_2467_0, i_10_416_2514_0, i_10_416_2568_0,
    i_10_416_2629_0, i_10_416_2631_0, i_10_416_2632_0, i_10_416_2642_0,
    i_10_416_2660_0, i_10_416_2702_0, i_10_416_2713_0, i_10_416_2719_0,
    i_10_416_2722_0, i_10_416_2727_0, i_10_416_2729_0, i_10_416_2746_0,
    i_10_416_2917_0, i_10_416_3033_0, i_10_416_3290_0, i_10_416_3384_0,
    i_10_416_3386_0, i_10_416_3387_0, i_10_416_3388_0, i_10_416_3389_0,
    i_10_416_3448_0, i_10_416_3465_0, i_10_416_3556_0, i_10_416_3584_0,
    i_10_416_3601_0, i_10_416_3614_0, i_10_416_3787_0, i_10_416_3788_0,
    i_10_416_3844_0, i_10_416_3845_0, i_10_416_3848_0, i_10_416_3890_0,
    i_10_416_3974_0, i_10_416_3978_0, i_10_416_3990_0, i_10_416_4126_0,
    i_10_416_4167_0, i_10_416_4168_0, i_10_416_4187_0, i_10_416_4268_0,
    i_10_416_4275_0, i_10_416_4288_0, i_10_416_4307_0, i_10_416_4394_0,
    i_10_416_4395_0, i_10_416_4397_0, i_10_416_4447_0, i_10_416_4572_0,
    o_10_416_0_0  );
  input  i_10_416_144_0, i_10_416_174_0, i_10_416_216_0, i_10_416_236_0,
    i_10_416_279_0, i_10_416_426_0, i_10_416_433_0, i_10_416_435_0,
    i_10_416_441_0, i_10_416_442_0, i_10_416_443_0, i_10_416_444_0,
    i_10_416_446_0, i_10_416_463_0, i_10_416_515_0, i_10_416_518_0,
    i_10_416_792_0, i_10_416_793_0, i_10_416_794_0, i_10_416_820_0,
    i_10_416_892_0, i_10_416_957_0, i_10_416_967_0, i_10_416_1083_0,
    i_10_416_1084_0, i_10_416_1202_0, i_10_416_1360_0, i_10_416_1377_0,
    i_10_416_1485_0, i_10_416_1546_0, i_10_416_1576_0, i_10_416_1581_0,
    i_10_416_1631_0, i_10_416_1691_0, i_10_416_1728_0, i_10_416_1818_0,
    i_10_416_1820_0, i_10_416_1954_0, i_10_416_2045_0, i_10_416_2200_0,
    i_10_416_2202_0, i_10_416_2225_0, i_10_416_2288_0, i_10_416_2331_0,
    i_10_416_2352_0, i_10_416_2357_0, i_10_416_2358_0, i_10_416_2360_0,
    i_10_416_2377_0, i_10_416_2467_0, i_10_416_2514_0, i_10_416_2568_0,
    i_10_416_2629_0, i_10_416_2631_0, i_10_416_2632_0, i_10_416_2642_0,
    i_10_416_2660_0, i_10_416_2702_0, i_10_416_2713_0, i_10_416_2719_0,
    i_10_416_2722_0, i_10_416_2727_0, i_10_416_2729_0, i_10_416_2746_0,
    i_10_416_2917_0, i_10_416_3033_0, i_10_416_3290_0, i_10_416_3384_0,
    i_10_416_3386_0, i_10_416_3387_0, i_10_416_3388_0, i_10_416_3389_0,
    i_10_416_3448_0, i_10_416_3465_0, i_10_416_3556_0, i_10_416_3584_0,
    i_10_416_3601_0, i_10_416_3614_0, i_10_416_3787_0, i_10_416_3788_0,
    i_10_416_3844_0, i_10_416_3845_0, i_10_416_3848_0, i_10_416_3890_0,
    i_10_416_3974_0, i_10_416_3978_0, i_10_416_3990_0, i_10_416_4126_0,
    i_10_416_4167_0, i_10_416_4168_0, i_10_416_4187_0, i_10_416_4268_0,
    i_10_416_4275_0, i_10_416_4288_0, i_10_416_4307_0, i_10_416_4394_0,
    i_10_416_4395_0, i_10_416_4397_0, i_10_416_4447_0, i_10_416_4572_0;
  output o_10_416_0_0;
  assign o_10_416_0_0 = 0;
endmodule



// Benchmark "kernel_10_417" written by ABC on Sun Jul 19 10:28:19 2020

module kernel_10_417 ( 
    i_10_417_46_0, i_10_417_175_0, i_10_417_177_0, i_10_417_219_0,
    i_10_417_222_0, i_10_417_284_0, i_10_417_319_0, i_10_417_322_0,
    i_10_417_327_0, i_10_417_330_0, i_10_417_331_0, i_10_417_442_0,
    i_10_417_751_0, i_10_417_955_0, i_10_417_1032_0, i_10_417_1034_0,
    i_10_417_1237_0, i_10_417_1239_0, i_10_417_1240_0, i_10_417_1248_0,
    i_10_417_1308_0, i_10_417_1311_0, i_10_417_1363_0, i_10_417_1431_0,
    i_10_417_1444_0, i_10_417_1541_0, i_10_417_1549_0, i_10_417_1553_0,
    i_10_417_1556_0, i_10_417_1576_0, i_10_417_1577_0, i_10_417_1683_0,
    i_10_417_1803_0, i_10_417_1820_0, i_10_417_1826_0, i_10_417_1948_0,
    i_10_417_1981_0, i_10_417_1996_0, i_10_417_2017_0, i_10_417_2019_0,
    i_10_417_2028_0, i_10_417_2355_0, i_10_417_2357_0, i_10_417_2462_0,
    i_10_417_2466_0, i_10_417_2508_0, i_10_417_2608_0, i_10_417_2629_0,
    i_10_417_2631_0, i_10_417_2658_0, i_10_417_2659_0, i_10_417_2662_0,
    i_10_417_2663_0, i_10_417_2704_0, i_10_417_2723_0, i_10_417_2724_0,
    i_10_417_2725_0, i_10_417_2726_0, i_10_417_2731_0, i_10_417_2739_0,
    i_10_417_2742_0, i_10_417_2782_0, i_10_417_2823_0, i_10_417_2830_0,
    i_10_417_2831_0, i_10_417_2832_0, i_10_417_2833_0, i_10_417_2834_0,
    i_10_417_2880_0, i_10_417_2982_0, i_10_417_3049_0, i_10_417_3090_0,
    i_10_417_3270_0, i_10_417_3278_0, i_10_417_3279_0, i_10_417_3283_0,
    i_10_417_3469_0, i_10_417_3582_0, i_10_417_3612_0, i_10_417_3645_0,
    i_10_417_3648_0, i_10_417_3649_0, i_10_417_3650_0, i_10_417_3651_0,
    i_10_417_3780_0, i_10_417_3835_0, i_10_417_3837_0, i_10_417_3841_0,
    i_10_417_3860_0, i_10_417_3895_0, i_10_417_3896_0, i_10_417_4113_0,
    i_10_417_4116_0, i_10_417_4123_0, i_10_417_4275_0, i_10_417_4276_0,
    i_10_417_4279_0, i_10_417_4290_0, i_10_417_4291_0, i_10_417_4581_0,
    o_10_417_0_0  );
  input  i_10_417_46_0, i_10_417_175_0, i_10_417_177_0, i_10_417_219_0,
    i_10_417_222_0, i_10_417_284_0, i_10_417_319_0, i_10_417_322_0,
    i_10_417_327_0, i_10_417_330_0, i_10_417_331_0, i_10_417_442_0,
    i_10_417_751_0, i_10_417_955_0, i_10_417_1032_0, i_10_417_1034_0,
    i_10_417_1237_0, i_10_417_1239_0, i_10_417_1240_0, i_10_417_1248_0,
    i_10_417_1308_0, i_10_417_1311_0, i_10_417_1363_0, i_10_417_1431_0,
    i_10_417_1444_0, i_10_417_1541_0, i_10_417_1549_0, i_10_417_1553_0,
    i_10_417_1556_0, i_10_417_1576_0, i_10_417_1577_0, i_10_417_1683_0,
    i_10_417_1803_0, i_10_417_1820_0, i_10_417_1826_0, i_10_417_1948_0,
    i_10_417_1981_0, i_10_417_1996_0, i_10_417_2017_0, i_10_417_2019_0,
    i_10_417_2028_0, i_10_417_2355_0, i_10_417_2357_0, i_10_417_2462_0,
    i_10_417_2466_0, i_10_417_2508_0, i_10_417_2608_0, i_10_417_2629_0,
    i_10_417_2631_0, i_10_417_2658_0, i_10_417_2659_0, i_10_417_2662_0,
    i_10_417_2663_0, i_10_417_2704_0, i_10_417_2723_0, i_10_417_2724_0,
    i_10_417_2725_0, i_10_417_2726_0, i_10_417_2731_0, i_10_417_2739_0,
    i_10_417_2742_0, i_10_417_2782_0, i_10_417_2823_0, i_10_417_2830_0,
    i_10_417_2831_0, i_10_417_2832_0, i_10_417_2833_0, i_10_417_2834_0,
    i_10_417_2880_0, i_10_417_2982_0, i_10_417_3049_0, i_10_417_3090_0,
    i_10_417_3270_0, i_10_417_3278_0, i_10_417_3279_0, i_10_417_3283_0,
    i_10_417_3469_0, i_10_417_3582_0, i_10_417_3612_0, i_10_417_3645_0,
    i_10_417_3648_0, i_10_417_3649_0, i_10_417_3650_0, i_10_417_3651_0,
    i_10_417_3780_0, i_10_417_3835_0, i_10_417_3837_0, i_10_417_3841_0,
    i_10_417_3860_0, i_10_417_3895_0, i_10_417_3896_0, i_10_417_4113_0,
    i_10_417_4116_0, i_10_417_4123_0, i_10_417_4275_0, i_10_417_4276_0,
    i_10_417_4279_0, i_10_417_4290_0, i_10_417_4291_0, i_10_417_4581_0;
  output o_10_417_0_0;
  assign o_10_417_0_0 = 0;
endmodule



// Benchmark "kernel_10_418" written by ABC on Sun Jul 19 10:28:20 2020

module kernel_10_418 ( 
    i_10_418_274_0, i_10_418_275_0, i_10_418_282_0, i_10_418_317_0,
    i_10_418_328_0, i_10_418_432_0, i_10_418_433_0, i_10_418_434_0,
    i_10_418_436_0, i_10_418_437_0, i_10_418_446_0, i_10_418_460_0,
    i_10_418_463_0, i_10_418_464_0, i_10_418_518_0, i_10_418_907_0,
    i_10_418_1032_0, i_10_418_1033_0, i_10_418_1043_0, i_10_418_1138_0,
    i_10_418_1265_0, i_10_418_1309_0, i_10_418_1345_0, i_10_418_1346_0,
    i_10_418_1349_0, i_10_418_1445_0, i_10_418_1546_0, i_10_418_1575_0,
    i_10_418_1654_0, i_10_418_1720_0, i_10_418_1767_0, i_10_418_1768_0,
    i_10_418_1769_0, i_10_418_1821_0, i_10_418_1912_0, i_10_418_1913_0,
    i_10_418_1916_0, i_10_418_2352_0, i_10_418_2365_0, i_10_418_2383_0,
    i_10_418_2384_0, i_10_418_2408_0, i_10_418_2471_0, i_10_418_2512_0,
    i_10_418_2629_0, i_10_418_2630_0, i_10_418_2656_0, i_10_418_2657_0,
    i_10_418_2659_0, i_10_418_2660_0, i_10_418_2661_0, i_10_418_2675_0,
    i_10_418_2678_0, i_10_418_2681_0, i_10_418_2705_0, i_10_418_2723_0,
    i_10_418_2728_0, i_10_418_2729_0, i_10_418_2819_0, i_10_418_2822_0,
    i_10_418_2823_0, i_10_418_2824_0, i_10_418_2828_0, i_10_418_2830_0,
    i_10_418_2831_0, i_10_418_2880_0, i_10_418_2919_0, i_10_418_2980_0,
    i_10_418_3033_0, i_10_418_3034_0, i_10_418_3050_0, i_10_418_3070_0,
    i_10_418_3088_0, i_10_418_3093_0, i_10_418_3150_0, i_10_418_3151_0,
    i_10_418_3160_0, i_10_418_3280_0, i_10_418_3281_0, i_10_418_3322_0,
    i_10_418_3323_0, i_10_418_3349_0, i_10_418_3350_0, i_10_418_3387_0,
    i_10_418_3437_0, i_10_418_3523_0, i_10_418_3587_0, i_10_418_3590_0,
    i_10_418_3613_0, i_10_418_3648_0, i_10_418_3685_0, i_10_418_3842_0,
    i_10_418_3856_0, i_10_418_3857_0, i_10_418_3910_0, i_10_418_4115_0,
    i_10_418_4175_0, i_10_418_4236_0, i_10_418_4267_0, i_10_418_4289_0,
    o_10_418_0_0  );
  input  i_10_418_274_0, i_10_418_275_0, i_10_418_282_0, i_10_418_317_0,
    i_10_418_328_0, i_10_418_432_0, i_10_418_433_0, i_10_418_434_0,
    i_10_418_436_0, i_10_418_437_0, i_10_418_446_0, i_10_418_460_0,
    i_10_418_463_0, i_10_418_464_0, i_10_418_518_0, i_10_418_907_0,
    i_10_418_1032_0, i_10_418_1033_0, i_10_418_1043_0, i_10_418_1138_0,
    i_10_418_1265_0, i_10_418_1309_0, i_10_418_1345_0, i_10_418_1346_0,
    i_10_418_1349_0, i_10_418_1445_0, i_10_418_1546_0, i_10_418_1575_0,
    i_10_418_1654_0, i_10_418_1720_0, i_10_418_1767_0, i_10_418_1768_0,
    i_10_418_1769_0, i_10_418_1821_0, i_10_418_1912_0, i_10_418_1913_0,
    i_10_418_1916_0, i_10_418_2352_0, i_10_418_2365_0, i_10_418_2383_0,
    i_10_418_2384_0, i_10_418_2408_0, i_10_418_2471_0, i_10_418_2512_0,
    i_10_418_2629_0, i_10_418_2630_0, i_10_418_2656_0, i_10_418_2657_0,
    i_10_418_2659_0, i_10_418_2660_0, i_10_418_2661_0, i_10_418_2675_0,
    i_10_418_2678_0, i_10_418_2681_0, i_10_418_2705_0, i_10_418_2723_0,
    i_10_418_2728_0, i_10_418_2729_0, i_10_418_2819_0, i_10_418_2822_0,
    i_10_418_2823_0, i_10_418_2824_0, i_10_418_2828_0, i_10_418_2830_0,
    i_10_418_2831_0, i_10_418_2880_0, i_10_418_2919_0, i_10_418_2980_0,
    i_10_418_3033_0, i_10_418_3034_0, i_10_418_3050_0, i_10_418_3070_0,
    i_10_418_3088_0, i_10_418_3093_0, i_10_418_3150_0, i_10_418_3151_0,
    i_10_418_3160_0, i_10_418_3280_0, i_10_418_3281_0, i_10_418_3322_0,
    i_10_418_3323_0, i_10_418_3349_0, i_10_418_3350_0, i_10_418_3387_0,
    i_10_418_3437_0, i_10_418_3523_0, i_10_418_3587_0, i_10_418_3590_0,
    i_10_418_3613_0, i_10_418_3648_0, i_10_418_3685_0, i_10_418_3842_0,
    i_10_418_3856_0, i_10_418_3857_0, i_10_418_3910_0, i_10_418_4115_0,
    i_10_418_4175_0, i_10_418_4236_0, i_10_418_4267_0, i_10_418_4289_0;
  output o_10_418_0_0;
  assign o_10_418_0_0 = ~((~i_10_418_317_0 & ((~i_10_418_436_0 & ~i_10_418_1345_0 & ~i_10_418_1349_0 & ~i_10_418_1767_0 & ~i_10_418_1769_0 & ~i_10_418_1912_0 & ~i_10_418_1916_0 & ~i_10_418_2823_0 & ~i_10_418_3587_0 & ~i_10_418_3648_0) | (~i_10_418_1445_0 & i_10_418_1821_0 & ~i_10_418_2675_0 & ~i_10_418_2830_0 & ~i_10_418_2880_0 & i_10_418_3280_0 & ~i_10_418_3910_0 & ~i_10_418_4236_0))) | (~i_10_418_4236_0 & ((~i_10_418_2729_0 & ((~i_10_418_436_0 & ((~i_10_418_518_0 & ~i_10_418_1769_0 & ~i_10_418_2681_0 & ~i_10_418_2728_0 & ~i_10_418_2823_0) | (~i_10_418_282_0 & ~i_10_418_2629_0 & ~i_10_418_2830_0 & ~i_10_418_3093_0 & ~i_10_418_3437_0 & ~i_10_418_3648_0 & ~i_10_418_4175_0))) | (i_10_418_436_0 & ~i_10_418_1767_0 & ~i_10_418_1768_0 & ~i_10_418_2384_0 & ~i_10_418_2630_0 & ~i_10_418_2656_0 & ~i_10_418_2660_0 & ~i_10_418_3437_0))) | (~i_10_418_437_0 & ((~i_10_418_2657_0 & i_10_418_2661_0 & ~i_10_418_3280_0 & ~i_10_418_3437_0 & ~i_10_418_3587_0) | (~i_10_418_328_0 & ~i_10_418_518_0 & ~i_10_418_907_0 & ~i_10_418_1767_0 & ~i_10_418_1912_0 & ~i_10_418_2408_0 & ~i_10_418_2823_0 & ~i_10_418_3034_0 & ~i_10_418_3088_0 & ~i_10_418_3093_0 & ~i_10_418_3160_0 & ~i_10_418_4115_0))) | (~i_10_418_2675_0 & ~i_10_418_2824_0 & ((~i_10_418_1346_0 & ~i_10_418_1349_0 & ~i_10_418_2656_0 & ~i_10_418_2678_0 & ~i_10_418_3437_0) | (~i_10_418_1767_0 & ~i_10_418_1769_0 & ~i_10_418_1916_0 & ~i_10_418_2657_0 & ~i_10_418_3034_0 & ~i_10_418_3910_0))))) | (~i_10_418_328_0 & ~i_10_418_1767_0 & ((~i_10_418_2723_0 & ~i_10_418_2824_0 & ~i_10_418_2830_0 & ~i_10_418_3033_0 & ~i_10_418_3093_0 & ~i_10_418_3587_0 & ~i_10_418_3842_0) | (~i_10_418_432_0 & ~i_10_418_1349_0 & ~i_10_418_1916_0 & ~i_10_418_2675_0 & ~i_10_418_2681_0 & ~i_10_418_2822_0 & ~i_10_418_2828_0 & ~i_10_418_3088_0 & ~i_10_418_3280_0 & ~i_10_418_4289_0))) | (~i_10_418_907_0 & ((~i_10_418_1349_0 & ~i_10_418_2629_0 & ~i_10_418_2681_0 & ~i_10_418_3034_0 & ~i_10_418_3280_0 & ~i_10_418_3523_0) | (~i_10_418_460_0 & ~i_10_418_1768_0 & ~i_10_418_2630_0 & ~i_10_418_2678_0 & ~i_10_418_2824_0 & ~i_10_418_3050_0 & ~i_10_418_4289_0))) | (~i_10_418_1916_0 & ((~i_10_418_2657_0 & ~i_10_418_2660_0 & ~i_10_418_2723_0 & ~i_10_418_2822_0 & ~i_10_418_2831_0 & ~i_10_418_3280_0 & ~i_10_418_3281_0) | (~i_10_418_1309_0 & ~i_10_418_2728_0 & ~i_10_418_2828_0 & ~i_10_418_3088_0 & i_10_418_3281_0 & ~i_10_418_3910_0 & i_10_418_4289_0))) | (~i_10_418_1768_0 & ((~i_10_418_2660_0 & ((~i_10_418_433_0 & i_10_418_1767_0 & ~i_10_418_2728_0 & ~i_10_418_3523_0) | (~i_10_418_1345_0 & ~i_10_418_1445_0 & ~i_10_418_2678_0 & ~i_10_418_2819_0 & ~i_10_418_3437_0 & ~i_10_418_3590_0))) | (i_10_418_2384_0 & ~i_10_418_2675_0 & ~i_10_418_2823_0))));
endmodule



// Benchmark "kernel_10_419" written by ABC on Sun Jul 19 10:28:21 2020

module kernel_10_419 ( 
    i_10_419_145_0, i_10_419_174_0, i_10_419_217_0, i_10_419_282_0,
    i_10_419_287_0, i_10_419_293_0, i_10_419_296_0, i_10_419_430_0,
    i_10_419_443_0, i_10_419_459_0, i_10_419_462_0, i_10_419_465_0,
    i_10_419_581_0, i_10_419_699_0, i_10_419_751_0, i_10_419_794_0,
    i_10_419_798_0, i_10_419_835_0, i_10_419_894_0, i_10_419_897_0,
    i_10_419_1030_0, i_10_419_1040_0, i_10_419_1043_0, i_10_419_1234_0,
    i_10_419_1235_0, i_10_419_1236_0, i_10_419_1239_0, i_10_419_1240_0,
    i_10_419_1248_0, i_10_419_1249_0, i_10_419_1309_0, i_10_419_1311_0,
    i_10_419_1312_0, i_10_419_1344_0, i_10_419_1575_0, i_10_419_1637_0,
    i_10_419_1648_0, i_10_419_1650_0, i_10_419_1651_0, i_10_419_1655_0,
    i_10_419_1684_0, i_10_419_1685_0, i_10_419_1686_0, i_10_419_1697_0,
    i_10_419_1798_0, i_10_419_1822_0, i_10_419_2166_0, i_10_419_2201_0,
    i_10_419_2266_0, i_10_419_2327_0, i_10_419_2337_0, i_10_419_2338_0,
    i_10_419_2339_0, i_10_419_2449_0, i_10_419_2451_0, i_10_419_2510_0,
    i_10_419_2559_0, i_10_419_2562_0, i_10_419_2571_0, i_10_419_2636_0,
    i_10_419_2643_0, i_10_419_2652_0, i_10_419_2661_0, i_10_419_2662_0,
    i_10_419_2705_0, i_10_419_2708_0, i_10_419_2717_0, i_10_419_2781_0,
    i_10_419_2782_0, i_10_419_2984_0, i_10_419_3076_0, i_10_419_3201_0,
    i_10_419_3268_0, i_10_419_3270_0, i_10_419_3272_0, i_10_419_3273_0,
    i_10_419_3274_0, i_10_419_3280_0, i_10_419_3405_0, i_10_419_3611_0,
    i_10_419_3612_0, i_10_419_3649_0, i_10_419_3652_0, i_10_419_3703_0,
    i_10_419_3704_0, i_10_419_3783_0, i_10_419_3784_0, i_10_419_3785_0,
    i_10_419_3787_0, i_10_419_3838_0, i_10_419_3859_0, i_10_419_3896_0,
    i_10_419_4027_0, i_10_419_4269_0, i_10_419_4276_0, i_10_419_4277_0,
    i_10_419_4281_0, i_10_419_4292_0, i_10_419_4463_0, i_10_419_4508_0,
    o_10_419_0_0  );
  input  i_10_419_145_0, i_10_419_174_0, i_10_419_217_0, i_10_419_282_0,
    i_10_419_287_0, i_10_419_293_0, i_10_419_296_0, i_10_419_430_0,
    i_10_419_443_0, i_10_419_459_0, i_10_419_462_0, i_10_419_465_0,
    i_10_419_581_0, i_10_419_699_0, i_10_419_751_0, i_10_419_794_0,
    i_10_419_798_0, i_10_419_835_0, i_10_419_894_0, i_10_419_897_0,
    i_10_419_1030_0, i_10_419_1040_0, i_10_419_1043_0, i_10_419_1234_0,
    i_10_419_1235_0, i_10_419_1236_0, i_10_419_1239_0, i_10_419_1240_0,
    i_10_419_1248_0, i_10_419_1249_0, i_10_419_1309_0, i_10_419_1311_0,
    i_10_419_1312_0, i_10_419_1344_0, i_10_419_1575_0, i_10_419_1637_0,
    i_10_419_1648_0, i_10_419_1650_0, i_10_419_1651_0, i_10_419_1655_0,
    i_10_419_1684_0, i_10_419_1685_0, i_10_419_1686_0, i_10_419_1697_0,
    i_10_419_1798_0, i_10_419_1822_0, i_10_419_2166_0, i_10_419_2201_0,
    i_10_419_2266_0, i_10_419_2327_0, i_10_419_2337_0, i_10_419_2338_0,
    i_10_419_2339_0, i_10_419_2449_0, i_10_419_2451_0, i_10_419_2510_0,
    i_10_419_2559_0, i_10_419_2562_0, i_10_419_2571_0, i_10_419_2636_0,
    i_10_419_2643_0, i_10_419_2652_0, i_10_419_2661_0, i_10_419_2662_0,
    i_10_419_2705_0, i_10_419_2708_0, i_10_419_2717_0, i_10_419_2781_0,
    i_10_419_2782_0, i_10_419_2984_0, i_10_419_3076_0, i_10_419_3201_0,
    i_10_419_3268_0, i_10_419_3270_0, i_10_419_3272_0, i_10_419_3273_0,
    i_10_419_3274_0, i_10_419_3280_0, i_10_419_3405_0, i_10_419_3611_0,
    i_10_419_3612_0, i_10_419_3649_0, i_10_419_3652_0, i_10_419_3703_0,
    i_10_419_3704_0, i_10_419_3783_0, i_10_419_3784_0, i_10_419_3785_0,
    i_10_419_3787_0, i_10_419_3838_0, i_10_419_3859_0, i_10_419_3896_0,
    i_10_419_4027_0, i_10_419_4269_0, i_10_419_4276_0, i_10_419_4277_0,
    i_10_419_4281_0, i_10_419_4292_0, i_10_419_4463_0, i_10_419_4508_0;
  output o_10_419_0_0;
  assign o_10_419_0_0 = 0;
endmodule



// Benchmark "kernel_10_420" written by ABC on Sun Jul 19 10:28:22 2020

module kernel_10_420 ( 
    i_10_420_151_0, i_10_420_157_0, i_10_420_268_0, i_10_420_273_0,
    i_10_420_278_0, i_10_420_282_0, i_10_420_283_0, i_10_420_322_0,
    i_10_420_391_0, i_10_420_442_0, i_10_420_508_0, i_10_420_691_0,
    i_10_420_716_0, i_10_420_718_0, i_10_420_719_0, i_10_420_739_0,
    i_10_420_754_0, i_10_420_755_0, i_10_420_795_0, i_10_420_931_0,
    i_10_420_959_0, i_10_420_966_0, i_10_420_968_0, i_10_420_970_0,
    i_10_420_991_0, i_10_420_992_0, i_10_420_1165_0, i_10_420_1166_0,
    i_10_420_1197_0, i_10_420_1198_0, i_10_420_1235_0, i_10_420_1249_0,
    i_10_420_1250_0, i_10_420_1262_0, i_10_420_1359_0, i_10_420_1360_0,
    i_10_420_1440_0, i_10_420_1441_0, i_10_420_1442_0, i_10_420_1491_0,
    i_10_420_1492_0, i_10_420_1536_0, i_10_420_1537_0, i_10_420_1555_0,
    i_10_420_1582_0, i_10_420_1629_0, i_10_420_1691_0, i_10_420_1852_0,
    i_10_420_2002_0, i_10_420_2005_0, i_10_420_2006_0, i_10_420_2019_0,
    i_10_420_2186_0, i_10_420_2351_0, i_10_420_2392_0, i_10_420_2533_0,
    i_10_420_2535_0, i_10_420_2573_0, i_10_420_2609_0, i_10_420_2620_0,
    i_10_420_2621_0, i_10_420_2680_0, i_10_420_2708_0, i_10_420_2725_0,
    i_10_420_2727_0, i_10_420_2735_0, i_10_420_2781_0, i_10_420_2786_0,
    i_10_420_2882_0, i_10_420_2885_0, i_10_420_2919_0, i_10_420_2920_0,
    i_10_420_2982_0, i_10_420_3038_0, i_10_420_3238_0, i_10_420_3384_0,
    i_10_420_3385_0, i_10_420_3386_0, i_10_420_3392_0, i_10_420_3561_0,
    i_10_420_3562_0, i_10_420_3719_0, i_10_420_3786_0, i_10_420_3787_0,
    i_10_420_3846_0, i_10_420_3857_0, i_10_420_3877_0, i_10_420_3897_0,
    i_10_420_3898_0, i_10_420_3912_0, i_10_420_3913_0, i_10_420_3914_0,
    i_10_420_4113_0, i_10_420_4116_0, i_10_420_4118_0, i_10_420_4121_0,
    i_10_420_4204_0, i_10_420_4339_0, i_10_420_4460_0, i_10_420_4463_0,
    o_10_420_0_0  );
  input  i_10_420_151_0, i_10_420_157_0, i_10_420_268_0, i_10_420_273_0,
    i_10_420_278_0, i_10_420_282_0, i_10_420_283_0, i_10_420_322_0,
    i_10_420_391_0, i_10_420_442_0, i_10_420_508_0, i_10_420_691_0,
    i_10_420_716_0, i_10_420_718_0, i_10_420_719_0, i_10_420_739_0,
    i_10_420_754_0, i_10_420_755_0, i_10_420_795_0, i_10_420_931_0,
    i_10_420_959_0, i_10_420_966_0, i_10_420_968_0, i_10_420_970_0,
    i_10_420_991_0, i_10_420_992_0, i_10_420_1165_0, i_10_420_1166_0,
    i_10_420_1197_0, i_10_420_1198_0, i_10_420_1235_0, i_10_420_1249_0,
    i_10_420_1250_0, i_10_420_1262_0, i_10_420_1359_0, i_10_420_1360_0,
    i_10_420_1440_0, i_10_420_1441_0, i_10_420_1442_0, i_10_420_1491_0,
    i_10_420_1492_0, i_10_420_1536_0, i_10_420_1537_0, i_10_420_1555_0,
    i_10_420_1582_0, i_10_420_1629_0, i_10_420_1691_0, i_10_420_1852_0,
    i_10_420_2002_0, i_10_420_2005_0, i_10_420_2006_0, i_10_420_2019_0,
    i_10_420_2186_0, i_10_420_2351_0, i_10_420_2392_0, i_10_420_2533_0,
    i_10_420_2535_0, i_10_420_2573_0, i_10_420_2609_0, i_10_420_2620_0,
    i_10_420_2621_0, i_10_420_2680_0, i_10_420_2708_0, i_10_420_2725_0,
    i_10_420_2727_0, i_10_420_2735_0, i_10_420_2781_0, i_10_420_2786_0,
    i_10_420_2882_0, i_10_420_2885_0, i_10_420_2919_0, i_10_420_2920_0,
    i_10_420_2982_0, i_10_420_3038_0, i_10_420_3238_0, i_10_420_3384_0,
    i_10_420_3385_0, i_10_420_3386_0, i_10_420_3392_0, i_10_420_3561_0,
    i_10_420_3562_0, i_10_420_3719_0, i_10_420_3786_0, i_10_420_3787_0,
    i_10_420_3846_0, i_10_420_3857_0, i_10_420_3877_0, i_10_420_3897_0,
    i_10_420_3898_0, i_10_420_3912_0, i_10_420_3913_0, i_10_420_3914_0,
    i_10_420_4113_0, i_10_420_4116_0, i_10_420_4118_0, i_10_420_4121_0,
    i_10_420_4204_0, i_10_420_4339_0, i_10_420_4460_0, i_10_420_4463_0;
  output o_10_420_0_0;
  assign o_10_420_0_0 = 0;
endmodule



// Benchmark "kernel_10_421" written by ABC on Sun Jul 19 10:28:23 2020

module kernel_10_421 ( 
    i_10_421_49_0, i_10_421_151_0, i_10_421_183_0, i_10_421_184_0,
    i_10_421_222_0, i_10_421_410_0, i_10_421_441_0, i_10_421_442_0,
    i_10_421_444_0, i_10_421_445_0, i_10_421_514_0, i_10_421_515_0,
    i_10_421_588_0, i_10_421_628_0, i_10_421_711_0, i_10_421_745_0,
    i_10_421_797_0, i_10_421_832_0, i_10_421_966_0, i_10_421_982_0,
    i_10_421_983_0, i_10_421_1005_0, i_10_421_1026_0, i_10_421_1033_0,
    i_10_421_1034_0, i_10_421_1086_0, i_10_421_1240_0, i_10_421_1250_0,
    i_10_421_1305_0, i_10_421_1308_0, i_10_421_1309_0, i_10_421_1345_0,
    i_10_421_1383_0, i_10_421_1385_0, i_10_421_1432_0, i_10_421_1438_0,
    i_10_421_1532_0, i_10_421_1647_0, i_10_421_1683_0, i_10_421_1743_0,
    i_10_421_1821_0, i_10_421_1822_0, i_10_421_1823_0, i_10_421_1995_0,
    i_10_421_1996_0, i_10_421_2094_0, i_10_421_2095_0, i_10_421_2180_0,
    i_10_421_2197_0, i_10_421_2243_0, i_10_421_2252_0, i_10_421_2355_0,
    i_10_421_2356_0, i_10_421_2451_0, i_10_421_2452_0, i_10_421_2453_0,
    i_10_421_2474_0, i_10_421_2514_0, i_10_421_2515_0, i_10_421_2516_0,
    i_10_421_2644_0, i_10_421_2679_0, i_10_421_2680_0, i_10_421_2722_0,
    i_10_421_2724_0, i_10_421_2734_0, i_10_421_2735_0, i_10_421_2740_0,
    i_10_421_2741_0, i_10_421_2831_0, i_10_421_2916_0, i_10_421_2917_0,
    i_10_421_2921_0, i_10_421_2922_0, i_10_421_2923_0, i_10_421_3039_0,
    i_10_421_3040_0, i_10_421_3195_0, i_10_421_3388_0, i_10_421_3389_0,
    i_10_421_3405_0, i_10_421_3453_0, i_10_421_3525_0, i_10_421_3586_0,
    i_10_421_3726_0, i_10_421_3781_0, i_10_421_3786_0, i_10_421_3855_0,
    i_10_421_3856_0, i_10_421_3982_0, i_10_421_4026_0, i_10_421_4121_0,
    i_10_421_4182_0, i_10_421_4188_0, i_10_421_4219_0, i_10_421_4220_0,
    i_10_421_4272_0, i_10_421_4292_0, i_10_421_4426_0, i_10_421_4570_0,
    o_10_421_0_0  );
  input  i_10_421_49_0, i_10_421_151_0, i_10_421_183_0, i_10_421_184_0,
    i_10_421_222_0, i_10_421_410_0, i_10_421_441_0, i_10_421_442_0,
    i_10_421_444_0, i_10_421_445_0, i_10_421_514_0, i_10_421_515_0,
    i_10_421_588_0, i_10_421_628_0, i_10_421_711_0, i_10_421_745_0,
    i_10_421_797_0, i_10_421_832_0, i_10_421_966_0, i_10_421_982_0,
    i_10_421_983_0, i_10_421_1005_0, i_10_421_1026_0, i_10_421_1033_0,
    i_10_421_1034_0, i_10_421_1086_0, i_10_421_1240_0, i_10_421_1250_0,
    i_10_421_1305_0, i_10_421_1308_0, i_10_421_1309_0, i_10_421_1345_0,
    i_10_421_1383_0, i_10_421_1385_0, i_10_421_1432_0, i_10_421_1438_0,
    i_10_421_1532_0, i_10_421_1647_0, i_10_421_1683_0, i_10_421_1743_0,
    i_10_421_1821_0, i_10_421_1822_0, i_10_421_1823_0, i_10_421_1995_0,
    i_10_421_1996_0, i_10_421_2094_0, i_10_421_2095_0, i_10_421_2180_0,
    i_10_421_2197_0, i_10_421_2243_0, i_10_421_2252_0, i_10_421_2355_0,
    i_10_421_2356_0, i_10_421_2451_0, i_10_421_2452_0, i_10_421_2453_0,
    i_10_421_2474_0, i_10_421_2514_0, i_10_421_2515_0, i_10_421_2516_0,
    i_10_421_2644_0, i_10_421_2679_0, i_10_421_2680_0, i_10_421_2722_0,
    i_10_421_2724_0, i_10_421_2734_0, i_10_421_2735_0, i_10_421_2740_0,
    i_10_421_2741_0, i_10_421_2831_0, i_10_421_2916_0, i_10_421_2917_0,
    i_10_421_2921_0, i_10_421_2922_0, i_10_421_2923_0, i_10_421_3039_0,
    i_10_421_3040_0, i_10_421_3195_0, i_10_421_3388_0, i_10_421_3389_0,
    i_10_421_3405_0, i_10_421_3453_0, i_10_421_3525_0, i_10_421_3586_0,
    i_10_421_3726_0, i_10_421_3781_0, i_10_421_3786_0, i_10_421_3855_0,
    i_10_421_3856_0, i_10_421_3982_0, i_10_421_4026_0, i_10_421_4121_0,
    i_10_421_4182_0, i_10_421_4188_0, i_10_421_4219_0, i_10_421_4220_0,
    i_10_421_4272_0, i_10_421_4292_0, i_10_421_4426_0, i_10_421_4570_0;
  output o_10_421_0_0;
  assign o_10_421_0_0 = 0;
endmodule



// Benchmark "kernel_10_422" written by ABC on Sun Jul 19 10:28:24 2020

module kernel_10_422 ( 
    i_10_422_32_0, i_10_422_33_0, i_10_422_34_0, i_10_422_53_0,
    i_10_422_143_0, i_10_422_172_0, i_10_422_178_0, i_10_422_179_0,
    i_10_422_188_0, i_10_422_265_0, i_10_422_269_0, i_10_422_274_0,
    i_10_422_277_0, i_10_422_278_0, i_10_422_391_0, i_10_422_440_0,
    i_10_422_462_0, i_10_422_464_0, i_10_422_520_0, i_10_422_755_0,
    i_10_422_934_0, i_10_422_962_0, i_10_422_1033_0, i_10_422_1061_0,
    i_10_422_1236_0, i_10_422_1237_0, i_10_422_1239_0, i_10_422_1240_0,
    i_10_422_1241_0, i_10_422_1246_0, i_10_422_1250_0, i_10_422_1308_0,
    i_10_422_1311_0, i_10_422_1382_0, i_10_422_1385_0, i_10_422_1436_0,
    i_10_422_1547_0, i_10_422_1653_0, i_10_422_1689_0, i_10_422_1819_0,
    i_10_422_1822_0, i_10_422_1824_0, i_10_422_1825_0, i_10_422_1956_0,
    i_10_422_1997_0, i_10_422_2201_0, i_10_422_2357_0, i_10_422_2363_0,
    i_10_422_2452_0, i_10_422_2460_0, i_10_422_2462_0, i_10_422_2469_0,
    i_10_422_2471_0, i_10_422_2474_0, i_10_422_2514_0, i_10_422_2517_0,
    i_10_422_2616_0, i_10_422_2630_0, i_10_422_2663_0, i_10_422_2711_0,
    i_10_422_2733_0, i_10_422_2735_0, i_10_422_2788_0, i_10_422_2789_0,
    i_10_422_2828_0, i_10_422_2832_0, i_10_422_2868_0, i_10_422_3035_0,
    i_10_422_3047_0, i_10_422_3196_0, i_10_422_3199_0, i_10_422_3203_0,
    i_10_422_3281_0, i_10_422_3454_0, i_10_422_3455_0, i_10_422_3470_0,
    i_10_422_3544_0, i_10_422_3552_0, i_10_422_3587_0, i_10_422_3611_0,
    i_10_422_3617_0, i_10_422_3650_0, i_10_422_3653_0, i_10_422_3683_0,
    i_10_422_3704_0, i_10_422_3785_0, i_10_422_3786_0, i_10_422_3788_0,
    i_10_422_3834_0, i_10_422_3835_0, i_10_422_3838_0, i_10_422_3847_0,
    i_10_422_3886_0, i_10_422_3887_0, i_10_422_3995_0, i_10_422_4004_0,
    i_10_422_4055_0, i_10_422_4057_0, i_10_422_4058_0, i_10_422_4382_0,
    o_10_422_0_0  );
  input  i_10_422_32_0, i_10_422_33_0, i_10_422_34_0, i_10_422_53_0,
    i_10_422_143_0, i_10_422_172_0, i_10_422_178_0, i_10_422_179_0,
    i_10_422_188_0, i_10_422_265_0, i_10_422_269_0, i_10_422_274_0,
    i_10_422_277_0, i_10_422_278_0, i_10_422_391_0, i_10_422_440_0,
    i_10_422_462_0, i_10_422_464_0, i_10_422_520_0, i_10_422_755_0,
    i_10_422_934_0, i_10_422_962_0, i_10_422_1033_0, i_10_422_1061_0,
    i_10_422_1236_0, i_10_422_1237_0, i_10_422_1239_0, i_10_422_1240_0,
    i_10_422_1241_0, i_10_422_1246_0, i_10_422_1250_0, i_10_422_1308_0,
    i_10_422_1311_0, i_10_422_1382_0, i_10_422_1385_0, i_10_422_1436_0,
    i_10_422_1547_0, i_10_422_1653_0, i_10_422_1689_0, i_10_422_1819_0,
    i_10_422_1822_0, i_10_422_1824_0, i_10_422_1825_0, i_10_422_1956_0,
    i_10_422_1997_0, i_10_422_2201_0, i_10_422_2357_0, i_10_422_2363_0,
    i_10_422_2452_0, i_10_422_2460_0, i_10_422_2462_0, i_10_422_2469_0,
    i_10_422_2471_0, i_10_422_2474_0, i_10_422_2514_0, i_10_422_2517_0,
    i_10_422_2616_0, i_10_422_2630_0, i_10_422_2663_0, i_10_422_2711_0,
    i_10_422_2733_0, i_10_422_2735_0, i_10_422_2788_0, i_10_422_2789_0,
    i_10_422_2828_0, i_10_422_2832_0, i_10_422_2868_0, i_10_422_3035_0,
    i_10_422_3047_0, i_10_422_3196_0, i_10_422_3199_0, i_10_422_3203_0,
    i_10_422_3281_0, i_10_422_3454_0, i_10_422_3455_0, i_10_422_3470_0,
    i_10_422_3544_0, i_10_422_3552_0, i_10_422_3587_0, i_10_422_3611_0,
    i_10_422_3617_0, i_10_422_3650_0, i_10_422_3653_0, i_10_422_3683_0,
    i_10_422_3704_0, i_10_422_3785_0, i_10_422_3786_0, i_10_422_3788_0,
    i_10_422_3834_0, i_10_422_3835_0, i_10_422_3838_0, i_10_422_3847_0,
    i_10_422_3886_0, i_10_422_3887_0, i_10_422_3995_0, i_10_422_4004_0,
    i_10_422_4055_0, i_10_422_4057_0, i_10_422_4058_0, i_10_422_4382_0;
  output o_10_422_0_0;
  assign o_10_422_0_0 = 0;
endmodule



// Benchmark "kernel_10_423" written by ABC on Sun Jul 19 10:28:25 2020

module kernel_10_423 ( 
    i_10_423_36_0, i_10_423_51_0, i_10_423_172_0, i_10_423_224_0,
    i_10_423_244_0, i_10_423_253_0, i_10_423_256_0, i_10_423_263_0,
    i_10_423_286_0, i_10_423_321_0, i_10_423_410_0, i_10_423_412_0,
    i_10_423_445_0, i_10_423_502_0, i_10_423_906_0, i_10_423_958_0,
    i_10_423_961_0, i_10_423_1030_0, i_10_423_1033_0, i_10_423_1034_0,
    i_10_423_1248_0, i_10_423_1249_0, i_10_423_1260_0, i_10_423_1310_0,
    i_10_423_1311_0, i_10_423_1346_0, i_10_423_1359_0, i_10_423_1434_0,
    i_10_423_1436_0, i_10_423_1451_0, i_10_423_1543_0, i_10_423_1576_0,
    i_10_423_1622_0, i_10_423_1651_0, i_10_423_1683_0, i_10_423_1687_0,
    i_10_423_1818_0, i_10_423_1819_0, i_10_423_1820_0, i_10_423_1821_0,
    i_10_423_1825_0, i_10_423_1909_0, i_10_423_1911_0, i_10_423_1912_0,
    i_10_423_1945_0, i_10_423_1950_0, i_10_423_1951_0, i_10_423_2182_0,
    i_10_423_2183_0, i_10_423_2304_0, i_10_423_2306_0, i_10_423_2350_0,
    i_10_423_2351_0, i_10_423_2356_0, i_10_423_2357_0, i_10_423_2362_0,
    i_10_423_2378_0, i_10_423_2384_0, i_10_423_2405_0, i_10_423_2451_0,
    i_10_423_2452_0, i_10_423_2453_0, i_10_423_2471_0, i_10_423_2518_0,
    i_10_423_2676_0, i_10_423_2715_0, i_10_423_2757_0, i_10_423_2850_0,
    i_10_423_2918_0, i_10_423_2921_0, i_10_423_3033_0, i_10_423_3070_0,
    i_10_423_3167_0, i_10_423_3198_0, i_10_423_3199_0, i_10_423_3278_0,
    i_10_423_3279_0, i_10_423_3326_0, i_10_423_3331_0, i_10_423_3432_0,
    i_10_423_3616_0, i_10_423_3645_0, i_10_423_3653_0, i_10_423_3721_0,
    i_10_423_3733_0, i_10_423_3787_0, i_10_423_3835_0, i_10_423_3839_0,
    i_10_423_3842_0, i_10_423_3852_0, i_10_423_3860_0, i_10_423_3983_0,
    i_10_423_4054_0, i_10_423_4116_0, i_10_423_4117_0, i_10_423_4119_0,
    i_10_423_4120_0, i_10_423_4168_0, i_10_423_4169_0, i_10_423_4277_0,
    o_10_423_0_0  );
  input  i_10_423_36_0, i_10_423_51_0, i_10_423_172_0, i_10_423_224_0,
    i_10_423_244_0, i_10_423_253_0, i_10_423_256_0, i_10_423_263_0,
    i_10_423_286_0, i_10_423_321_0, i_10_423_410_0, i_10_423_412_0,
    i_10_423_445_0, i_10_423_502_0, i_10_423_906_0, i_10_423_958_0,
    i_10_423_961_0, i_10_423_1030_0, i_10_423_1033_0, i_10_423_1034_0,
    i_10_423_1248_0, i_10_423_1249_0, i_10_423_1260_0, i_10_423_1310_0,
    i_10_423_1311_0, i_10_423_1346_0, i_10_423_1359_0, i_10_423_1434_0,
    i_10_423_1436_0, i_10_423_1451_0, i_10_423_1543_0, i_10_423_1576_0,
    i_10_423_1622_0, i_10_423_1651_0, i_10_423_1683_0, i_10_423_1687_0,
    i_10_423_1818_0, i_10_423_1819_0, i_10_423_1820_0, i_10_423_1821_0,
    i_10_423_1825_0, i_10_423_1909_0, i_10_423_1911_0, i_10_423_1912_0,
    i_10_423_1945_0, i_10_423_1950_0, i_10_423_1951_0, i_10_423_2182_0,
    i_10_423_2183_0, i_10_423_2304_0, i_10_423_2306_0, i_10_423_2350_0,
    i_10_423_2351_0, i_10_423_2356_0, i_10_423_2357_0, i_10_423_2362_0,
    i_10_423_2378_0, i_10_423_2384_0, i_10_423_2405_0, i_10_423_2451_0,
    i_10_423_2452_0, i_10_423_2453_0, i_10_423_2471_0, i_10_423_2518_0,
    i_10_423_2676_0, i_10_423_2715_0, i_10_423_2757_0, i_10_423_2850_0,
    i_10_423_2918_0, i_10_423_2921_0, i_10_423_3033_0, i_10_423_3070_0,
    i_10_423_3167_0, i_10_423_3198_0, i_10_423_3199_0, i_10_423_3278_0,
    i_10_423_3279_0, i_10_423_3326_0, i_10_423_3331_0, i_10_423_3432_0,
    i_10_423_3616_0, i_10_423_3645_0, i_10_423_3653_0, i_10_423_3721_0,
    i_10_423_3733_0, i_10_423_3787_0, i_10_423_3835_0, i_10_423_3839_0,
    i_10_423_3842_0, i_10_423_3852_0, i_10_423_3860_0, i_10_423_3983_0,
    i_10_423_4054_0, i_10_423_4116_0, i_10_423_4117_0, i_10_423_4119_0,
    i_10_423_4120_0, i_10_423_4168_0, i_10_423_4169_0, i_10_423_4277_0;
  output o_10_423_0_0;
  assign o_10_423_0_0 = 0;
endmodule



// Benchmark "kernel_10_424" written by ABC on Sun Jul 19 10:28:26 2020

module kernel_10_424 ( 
    i_10_424_150_0, i_10_424_172_0, i_10_424_174_0, i_10_424_182_0,
    i_10_424_285_0, i_10_424_327_0, i_10_424_410_0, i_10_424_444_0,
    i_10_424_447_0, i_10_424_513_0, i_10_424_516_0, i_10_424_717_0,
    i_10_424_795_0, i_10_424_797_0, i_10_424_798_0, i_10_424_963_0,
    i_10_424_964_0, i_10_424_966_0, i_10_424_967_0, i_10_424_1139_0,
    i_10_424_1163_0, i_10_424_1305_0, i_10_424_1308_0, i_10_424_1309_0,
    i_10_424_1311_0, i_10_424_1440_0, i_10_424_1444_0, i_10_424_1447_0,
    i_10_424_1491_0, i_10_424_1492_0, i_10_424_1556_0, i_10_424_1581_0,
    i_10_424_1582_0, i_10_424_1618_0, i_10_424_1635_0, i_10_424_1641_0,
    i_10_424_1726_0, i_10_424_1821_0, i_10_424_1824_0, i_10_424_1951_0,
    i_10_424_2184_0, i_10_424_2310_0, i_10_424_2322_0, i_10_424_2328_0,
    i_10_424_2351_0, i_10_424_2352_0, i_10_424_2377_0, i_10_424_2449_0,
    i_10_424_2472_0, i_10_424_2519_0, i_10_424_2660_0, i_10_424_2673_0,
    i_10_424_2679_0, i_10_424_2701_0, i_10_424_2727_0, i_10_424_2830_0,
    i_10_424_2880_0, i_10_424_2883_0, i_10_424_2885_0, i_10_424_2924_0,
    i_10_424_3035_0, i_10_424_3037_0, i_10_424_3038_0, i_10_424_3120_0,
    i_10_424_3152_0, i_10_424_3196_0, i_10_424_3198_0, i_10_424_3273_0,
    i_10_424_3323_0, i_10_424_3387_0, i_10_424_3405_0, i_10_424_3465_0,
    i_10_424_3468_0, i_10_424_3469_0, i_10_424_3495_0, i_10_424_3496_0,
    i_10_424_3585_0, i_10_424_3588_0, i_10_424_3610_0, i_10_424_3612_0,
    i_10_424_3613_0, i_10_424_3780_0, i_10_424_3805_0, i_10_424_3838_0,
    i_10_424_3840_0, i_10_424_3850_0, i_10_424_3853_0, i_10_424_3948_0,
    i_10_424_4120_0, i_10_424_4123_0, i_10_424_4213_0, i_10_424_4266_0,
    i_10_424_4270_0, i_10_424_4285_0, i_10_424_4287_0, i_10_424_4291_0,
    i_10_424_4458_0, i_10_424_4461_0, i_10_424_4564_0, i_10_424_4567_0,
    o_10_424_0_0  );
  input  i_10_424_150_0, i_10_424_172_0, i_10_424_174_0, i_10_424_182_0,
    i_10_424_285_0, i_10_424_327_0, i_10_424_410_0, i_10_424_444_0,
    i_10_424_447_0, i_10_424_513_0, i_10_424_516_0, i_10_424_717_0,
    i_10_424_795_0, i_10_424_797_0, i_10_424_798_0, i_10_424_963_0,
    i_10_424_964_0, i_10_424_966_0, i_10_424_967_0, i_10_424_1139_0,
    i_10_424_1163_0, i_10_424_1305_0, i_10_424_1308_0, i_10_424_1309_0,
    i_10_424_1311_0, i_10_424_1440_0, i_10_424_1444_0, i_10_424_1447_0,
    i_10_424_1491_0, i_10_424_1492_0, i_10_424_1556_0, i_10_424_1581_0,
    i_10_424_1582_0, i_10_424_1618_0, i_10_424_1635_0, i_10_424_1641_0,
    i_10_424_1726_0, i_10_424_1821_0, i_10_424_1824_0, i_10_424_1951_0,
    i_10_424_2184_0, i_10_424_2310_0, i_10_424_2322_0, i_10_424_2328_0,
    i_10_424_2351_0, i_10_424_2352_0, i_10_424_2377_0, i_10_424_2449_0,
    i_10_424_2472_0, i_10_424_2519_0, i_10_424_2660_0, i_10_424_2673_0,
    i_10_424_2679_0, i_10_424_2701_0, i_10_424_2727_0, i_10_424_2830_0,
    i_10_424_2880_0, i_10_424_2883_0, i_10_424_2885_0, i_10_424_2924_0,
    i_10_424_3035_0, i_10_424_3037_0, i_10_424_3038_0, i_10_424_3120_0,
    i_10_424_3152_0, i_10_424_3196_0, i_10_424_3198_0, i_10_424_3273_0,
    i_10_424_3323_0, i_10_424_3387_0, i_10_424_3405_0, i_10_424_3465_0,
    i_10_424_3468_0, i_10_424_3469_0, i_10_424_3495_0, i_10_424_3496_0,
    i_10_424_3585_0, i_10_424_3588_0, i_10_424_3610_0, i_10_424_3612_0,
    i_10_424_3613_0, i_10_424_3780_0, i_10_424_3805_0, i_10_424_3838_0,
    i_10_424_3840_0, i_10_424_3850_0, i_10_424_3853_0, i_10_424_3948_0,
    i_10_424_4120_0, i_10_424_4123_0, i_10_424_4213_0, i_10_424_4266_0,
    i_10_424_4270_0, i_10_424_4285_0, i_10_424_4287_0, i_10_424_4291_0,
    i_10_424_4458_0, i_10_424_4461_0, i_10_424_4564_0, i_10_424_4567_0;
  output o_10_424_0_0;
  assign o_10_424_0_0 = ~((~i_10_424_150_0 & ((~i_10_424_174_0 & ~i_10_424_513_0 & ~i_10_424_964_0 & ~i_10_424_2352_0 & ~i_10_424_2377_0 & ~i_10_424_3037_0 & ~i_10_424_3387_0 & ~i_10_424_4120_0) | (~i_10_424_447_0 & ~i_10_424_717_0 & ~i_10_424_1444_0 & ~i_10_424_3495_0 & ~i_10_424_4266_0 & ~i_10_424_4285_0 & ~i_10_424_4567_0))) | (~i_10_424_4266_0 & ((i_10_424_285_0 & ~i_10_424_3948_0 & ((~i_10_424_444_0 & i_10_424_1305_0 & ~i_10_424_3495_0) | (~i_10_424_717_0 & i_10_424_797_0 & ~i_10_424_3496_0 & ~i_10_424_4270_0))) | (~i_10_424_4213_0 & ((~i_10_424_516_0 & ((~i_10_424_717_0 & ~i_10_424_798_0 & ~i_10_424_967_0 & ~i_10_424_2377_0 & ~i_10_424_2472_0 & ~i_10_424_3198_0 & ~i_10_424_3469_0 & ~i_10_424_3496_0) | (~i_10_424_2328_0 & ~i_10_424_3585_0 & ~i_10_424_3612_0 & ~i_10_424_4270_0 & ~i_10_424_4287_0))) | (i_10_424_797_0 & ~i_10_424_966_0 & ~i_10_424_1440_0 & ~i_10_424_1447_0 & ~i_10_424_2310_0 & ~i_10_424_2351_0 & ~i_10_424_2449_0 & ~i_10_424_3387_0 & ~i_10_424_3469_0 & ~i_10_424_3496_0))) | (~i_10_424_963_0 & ~i_10_424_3495_0 & ((~i_10_424_447_0 & ~i_10_424_2322_0 & ~i_10_424_2727_0 & ~i_10_424_3588_0) | (~i_10_424_964_0 & ~i_10_424_2377_0 & ~i_10_424_2701_0 & ~i_10_424_3273_0 & ~i_10_424_3465_0 & ~i_10_424_3468_0 & ~i_10_424_3496_0 & ~i_10_424_3840_0 & ~i_10_424_4120_0))))) | (~i_10_424_717_0 & ((~i_10_424_516_0 & ~i_10_424_966_0 & ~i_10_424_1440_0 & ~i_10_424_1491_0 & ~i_10_424_1556_0 & i_10_424_1824_0 & ~i_10_424_2830_0) | (~i_10_424_963_0 & ~i_10_424_1447_0 & ~i_10_424_2310_0 & ~i_10_424_2322_0 & ~i_10_424_3495_0 & ~i_10_424_4123_0 & ~i_10_424_4270_0 & ~i_10_424_4564_0))) | (~i_10_424_798_0 & ((i_10_424_1308_0 & i_10_424_2660_0 & ~i_10_424_4120_0) | (~i_10_424_444_0 & ~i_10_424_513_0 & ~i_10_424_3838_0 & i_10_424_4120_0 & i_10_424_4564_0))) | (~i_10_424_444_0 & ((~i_10_424_964_0 & ~i_10_424_967_0 & i_10_424_1581_0 & ~i_10_424_4285_0) | (i_10_424_2660_0 & ~i_10_424_4213_0 & i_10_424_4287_0))) | (~i_10_424_964_0 & ((i_10_424_797_0 & ~i_10_424_966_0 & ~i_10_424_1444_0 & ~i_10_424_1492_0 & ~i_10_424_1951_0 & ~i_10_424_2673_0 & ~i_10_424_3469_0 & ~i_10_424_3496_0 & ~i_10_424_3850_0) | (~i_10_424_1491_0 & ~i_10_424_1821_0 & ~i_10_424_2322_0 & ~i_10_424_3273_0 & ~i_10_424_3838_0 & i_10_424_4291_0))) | (~i_10_424_967_0 & ((~i_10_424_2322_0 & ~i_10_424_2351_0 & ~i_10_424_3465_0 & i_10_424_3610_0) | (~i_10_424_966_0 & ~i_10_424_2472_0 & ~i_10_424_2679_0 & ~i_10_424_2830_0 & i_10_424_2924_0 & ~i_10_424_3196_0 & ~i_10_424_3273_0 & ~i_10_424_3387_0 & i_10_424_3850_0))) | (i_10_424_1308_0 & ((i_10_424_1305_0 & ~i_10_424_1556_0 & ~i_10_424_2322_0 & ~i_10_424_3495_0) | (~i_10_424_963_0 & ~i_10_424_4120_0 & i_10_424_4123_0))) | (i_10_424_3853_0 & ((~i_10_424_2322_0 & (i_10_424_3405_0 | (i_10_424_3850_0 & i_10_424_4285_0))) | (~i_10_424_3585_0 & ~i_10_424_4567_0))) | (i_10_424_2660_0 & (i_10_424_3198_0 | (i_10_424_4213_0 & ~i_10_424_4287_0))) | (~i_10_424_1821_0 & i_10_424_2377_0 & i_10_424_3198_0) | (i_10_424_172_0 & ~i_10_424_795_0 & ~i_10_424_4270_0 & i_10_424_4567_0) | (~i_10_424_1491_0 & ~i_10_424_2352_0 & ~i_10_424_2449_0 & ~i_10_424_2673_0 & ~i_10_424_3465_0 & ~i_10_424_3496_0 & ~i_10_424_4287_0 & ~i_10_424_4567_0));
endmodule



// Benchmark "kernel_10_425" written by ABC on Sun Jul 19 10:28:27 2020

module kernel_10_425 ( 
    i_10_425_86_0, i_10_425_221_0, i_10_425_286_0, i_10_425_287_0,
    i_10_425_293_0, i_10_425_315_0, i_10_425_410_0, i_10_425_428_0,
    i_10_425_437_0, i_10_425_443_0, i_10_425_444_0, i_10_425_448_0,
    i_10_425_455_0, i_10_425_520_0, i_10_425_700_0, i_10_425_794_0,
    i_10_425_798_0, i_10_425_881_0, i_10_425_971_0, i_10_425_1004_0,
    i_10_425_1026_0, i_10_425_1103_0, i_10_425_1235_0, i_10_425_1238_0,
    i_10_425_1240_0, i_10_425_1364_0, i_10_425_1432_0, i_10_425_1436_0,
    i_10_425_1577_0, i_10_425_1654_0, i_10_425_1688_0, i_10_425_1821_0,
    i_10_425_1875_0, i_10_425_1909_0, i_10_425_1913_0, i_10_425_1925_0,
    i_10_425_1952_0, i_10_425_2186_0, i_10_425_2363_0, i_10_425_2365_0,
    i_10_425_2366_0, i_10_425_2408_0, i_10_425_2451_0, i_10_425_2454_0,
    i_10_425_2455_0, i_10_425_2456_0, i_10_425_2470_0, i_10_425_2519_0,
    i_10_425_2617_0, i_10_425_2630_0, i_10_425_2645_0, i_10_425_2660_0,
    i_10_425_2681_0, i_10_425_2710_0, i_10_425_2719_0, i_10_425_2734_0,
    i_10_425_2882_0, i_10_425_2888_0, i_10_425_2923_0, i_10_425_2924_0,
    i_10_425_2986_0, i_10_425_3040_0, i_10_425_3041_0, i_10_425_3047_0,
    i_10_425_3049_0, i_10_425_3086_0, i_10_425_3153_0, i_10_425_3155_0,
    i_10_425_3156_0, i_10_425_3199_0, i_10_425_3202_0, i_10_425_3277_0,
    i_10_425_3283_0, i_10_425_3284_0, i_10_425_3302_0, i_10_425_3387_0,
    i_10_425_3389_0, i_10_425_3410_0, i_10_425_3465_0, i_10_425_3469_0,
    i_10_425_3503_0, i_10_425_3562_0, i_10_425_3613_0, i_10_425_3733_0,
    i_10_425_3785_0, i_10_425_3839_0, i_10_425_3853_0, i_10_425_3856_0,
    i_10_425_3857_0, i_10_425_3859_0, i_10_425_4030_0, i_10_425_4057_0,
    i_10_425_4058_0, i_10_425_4113_0, i_10_425_4117_0, i_10_425_4129_0,
    i_10_425_4130_0, i_10_425_4148_0, i_10_425_4237_0, i_10_425_4292_0,
    o_10_425_0_0  );
  input  i_10_425_86_0, i_10_425_221_0, i_10_425_286_0, i_10_425_287_0,
    i_10_425_293_0, i_10_425_315_0, i_10_425_410_0, i_10_425_428_0,
    i_10_425_437_0, i_10_425_443_0, i_10_425_444_0, i_10_425_448_0,
    i_10_425_455_0, i_10_425_520_0, i_10_425_700_0, i_10_425_794_0,
    i_10_425_798_0, i_10_425_881_0, i_10_425_971_0, i_10_425_1004_0,
    i_10_425_1026_0, i_10_425_1103_0, i_10_425_1235_0, i_10_425_1238_0,
    i_10_425_1240_0, i_10_425_1364_0, i_10_425_1432_0, i_10_425_1436_0,
    i_10_425_1577_0, i_10_425_1654_0, i_10_425_1688_0, i_10_425_1821_0,
    i_10_425_1875_0, i_10_425_1909_0, i_10_425_1913_0, i_10_425_1925_0,
    i_10_425_1952_0, i_10_425_2186_0, i_10_425_2363_0, i_10_425_2365_0,
    i_10_425_2366_0, i_10_425_2408_0, i_10_425_2451_0, i_10_425_2454_0,
    i_10_425_2455_0, i_10_425_2456_0, i_10_425_2470_0, i_10_425_2519_0,
    i_10_425_2617_0, i_10_425_2630_0, i_10_425_2645_0, i_10_425_2660_0,
    i_10_425_2681_0, i_10_425_2710_0, i_10_425_2719_0, i_10_425_2734_0,
    i_10_425_2882_0, i_10_425_2888_0, i_10_425_2923_0, i_10_425_2924_0,
    i_10_425_2986_0, i_10_425_3040_0, i_10_425_3041_0, i_10_425_3047_0,
    i_10_425_3049_0, i_10_425_3086_0, i_10_425_3153_0, i_10_425_3155_0,
    i_10_425_3156_0, i_10_425_3199_0, i_10_425_3202_0, i_10_425_3277_0,
    i_10_425_3283_0, i_10_425_3284_0, i_10_425_3302_0, i_10_425_3387_0,
    i_10_425_3389_0, i_10_425_3410_0, i_10_425_3465_0, i_10_425_3469_0,
    i_10_425_3503_0, i_10_425_3562_0, i_10_425_3613_0, i_10_425_3733_0,
    i_10_425_3785_0, i_10_425_3839_0, i_10_425_3853_0, i_10_425_3856_0,
    i_10_425_3857_0, i_10_425_3859_0, i_10_425_4030_0, i_10_425_4057_0,
    i_10_425_4058_0, i_10_425_4113_0, i_10_425_4117_0, i_10_425_4129_0,
    i_10_425_4130_0, i_10_425_4148_0, i_10_425_4237_0, i_10_425_4292_0;
  output o_10_425_0_0;
  assign o_10_425_0_0 = ~((~i_10_425_287_0 & ((~i_10_425_1240_0 & ~i_10_425_1913_0 & ~i_10_425_2660_0 & ~i_10_425_3410_0 & ~i_10_425_3859_0) | (~i_10_425_410_0 & ~i_10_425_444_0 & ~i_10_425_798_0 & ~i_10_425_1952_0 & ~i_10_425_4030_0))) | (~i_10_425_437_0 & ((~i_10_425_798_0 & ~i_10_425_1909_0 & ~i_10_425_1913_0 & ~i_10_425_2882_0 & ~i_10_425_3503_0 & ~i_10_425_3613_0 & ~i_10_425_3853_0 & ~i_10_425_4030_0) | (~i_10_425_293_0 & ~i_10_425_2719_0 & ~i_10_425_3041_0 & ~i_10_425_4129_0 & ~i_10_425_4130_0 & ~i_10_425_4237_0))) | (~i_10_425_2617_0 & ((~i_10_425_293_0 & ((~i_10_425_286_0 & ~i_10_425_1235_0 & ~i_10_425_1577_0 & ~i_10_425_4129_0 & ~i_10_425_4130_0) | (i_10_425_1240_0 & ~i_10_425_1952_0 & ~i_10_425_2681_0 & ~i_10_425_3613_0 & ~i_10_425_4292_0))) | (~i_10_425_4058_0 & ((i_10_425_455_0 & ~i_10_425_2630_0 & ~i_10_425_2734_0 & ~i_10_425_2923_0) | (~i_10_425_86_0 & ~i_10_425_1238_0 & ~i_10_425_1364_0 & ~i_10_425_2366_0 & ~i_10_425_3733_0 & ~i_10_425_4130_0))))) | (~i_10_425_86_0 & ((~i_10_425_1909_0 & ~i_10_425_2363_0 & ~i_10_425_3047_0 & ~i_10_425_3049_0 & ~i_10_425_4057_0) | (~i_10_425_1913_0 & ~i_10_425_2408_0 & ~i_10_425_2630_0 & ~i_10_425_3785_0 & ~i_10_425_3857_0 & ~i_10_425_4130_0))) | (~i_10_425_1004_0 & ((~i_10_425_448_0 & ~i_10_425_1913_0 & ~i_10_425_2186_0 & ~i_10_425_2365_0 & ~i_10_425_2719_0 & ~i_10_425_2734_0 & ~i_10_425_2882_0) | (~i_10_425_2455_0 & ~i_10_425_4030_0 & ~i_10_425_4057_0 & ~i_10_425_4058_0 & ~i_10_425_4237_0 & ~i_10_425_4292_0))) | (~i_10_425_2719_0 & ~i_10_425_4030_0 & ((~i_10_425_798_0 & ~i_10_425_1909_0 & ~i_10_425_3049_0 & ~i_10_425_3469_0 & ~i_10_425_4058_0 & i_10_425_4130_0) | (~i_10_425_2734_0 & ~i_10_425_2888_0 & ~i_10_425_2924_0 & ~i_10_425_3857_0 & ~i_10_425_4237_0))) | (~i_10_425_2365_0 & ~i_10_425_2366_0 & ~i_10_425_3040_0 & i_10_425_3199_0) | (~i_10_425_455_0 & ~i_10_425_794_0 & i_10_425_1238_0 & ~i_10_425_1821_0 & ~i_10_425_1913_0 & ~i_10_425_2734_0 & ~i_10_425_2882_0 & ~i_10_425_2888_0 & ~i_10_425_3277_0 & ~i_10_425_4237_0) | (~i_10_425_1952_0 & i_10_425_2455_0 & i_10_425_2456_0 & ~i_10_425_3389_0 & ~i_10_425_3465_0) | (~i_10_425_2710_0 & ~i_10_425_3049_0 & ~i_10_425_3202_0 & ~i_10_425_3856_0 & ~i_10_425_4130_0));
endmodule



// Benchmark "kernel_10_426" written by ABC on Sun Jul 19 10:28:28 2020

module kernel_10_426 ( 
    i_10_426_218_0, i_10_426_244_0, i_10_426_282_0, i_10_426_283_0,
    i_10_426_284_0, i_10_426_285_0, i_10_426_286_0, i_10_426_316_0,
    i_10_426_317_0, i_10_426_318_0, i_10_426_319_0, i_10_426_388_0,
    i_10_426_406_0, i_10_426_432_0, i_10_426_436_0, i_10_426_437_0,
    i_10_426_444_0, i_10_426_445_0, i_10_426_459_0, i_10_426_460_0,
    i_10_426_462_0, i_10_426_463_0, i_10_426_514_0, i_10_426_693_0,
    i_10_426_749_0, i_10_426_793_0, i_10_426_900_0, i_10_426_1000_0,
    i_10_426_1026_0, i_10_426_1027_0, i_10_426_1233_0, i_10_426_1242_0,
    i_10_426_1306_0, i_10_426_1441_0, i_10_426_1442_0, i_10_426_1546_0,
    i_10_426_1549_0, i_10_426_1650_0, i_10_426_1654_0, i_10_426_1819_0,
    i_10_426_1821_0, i_10_426_1822_0, i_10_426_1908_0, i_10_426_1946_0,
    i_10_426_1950_0, i_10_426_2304_0, i_10_426_2305_0, i_10_426_2306_0,
    i_10_426_2350_0, i_10_426_2359_0, i_10_426_2365_0, i_10_426_2404_0,
    i_10_426_2452_0, i_10_426_2454_0, i_10_426_2455_0, i_10_426_2459_0,
    i_10_426_2476_0, i_10_426_2477_0, i_10_426_2628_0, i_10_426_2629_0,
    i_10_426_2630_0, i_10_426_2632_0, i_10_426_2637_0, i_10_426_2638_0,
    i_10_426_2656_0, i_10_426_2657_0, i_10_426_2704_0, i_10_426_2817_0,
    i_10_426_2826_0, i_10_426_2827_0, i_10_426_2880_0, i_10_426_2918_0,
    i_10_426_2981_0, i_10_426_3034_0, i_10_426_3035_0, i_10_426_3047_0,
    i_10_426_3160_0, i_10_426_3200_0, i_10_426_3267_0, i_10_426_3271_0,
    i_10_426_3358_0, i_10_426_3384_0, i_10_426_3389_0, i_10_426_3402_0,
    i_10_426_3403_0, i_10_426_3404_0, i_10_426_3611_0, i_10_426_3613_0,
    i_10_426_3648_0, i_10_426_3682_0, i_10_426_3785_0, i_10_426_3808_0,
    i_10_426_3837_0, i_10_426_3843_0, i_10_426_3852_0, i_10_426_3859_0,
    i_10_426_3899_0, i_10_426_4171_0, i_10_426_4212_0, i_10_426_4276_0,
    o_10_426_0_0  );
  input  i_10_426_218_0, i_10_426_244_0, i_10_426_282_0, i_10_426_283_0,
    i_10_426_284_0, i_10_426_285_0, i_10_426_286_0, i_10_426_316_0,
    i_10_426_317_0, i_10_426_318_0, i_10_426_319_0, i_10_426_388_0,
    i_10_426_406_0, i_10_426_432_0, i_10_426_436_0, i_10_426_437_0,
    i_10_426_444_0, i_10_426_445_0, i_10_426_459_0, i_10_426_460_0,
    i_10_426_462_0, i_10_426_463_0, i_10_426_514_0, i_10_426_693_0,
    i_10_426_749_0, i_10_426_793_0, i_10_426_900_0, i_10_426_1000_0,
    i_10_426_1026_0, i_10_426_1027_0, i_10_426_1233_0, i_10_426_1242_0,
    i_10_426_1306_0, i_10_426_1441_0, i_10_426_1442_0, i_10_426_1546_0,
    i_10_426_1549_0, i_10_426_1650_0, i_10_426_1654_0, i_10_426_1819_0,
    i_10_426_1821_0, i_10_426_1822_0, i_10_426_1908_0, i_10_426_1946_0,
    i_10_426_1950_0, i_10_426_2304_0, i_10_426_2305_0, i_10_426_2306_0,
    i_10_426_2350_0, i_10_426_2359_0, i_10_426_2365_0, i_10_426_2404_0,
    i_10_426_2452_0, i_10_426_2454_0, i_10_426_2455_0, i_10_426_2459_0,
    i_10_426_2476_0, i_10_426_2477_0, i_10_426_2628_0, i_10_426_2629_0,
    i_10_426_2630_0, i_10_426_2632_0, i_10_426_2637_0, i_10_426_2638_0,
    i_10_426_2656_0, i_10_426_2657_0, i_10_426_2704_0, i_10_426_2817_0,
    i_10_426_2826_0, i_10_426_2827_0, i_10_426_2880_0, i_10_426_2918_0,
    i_10_426_2981_0, i_10_426_3034_0, i_10_426_3035_0, i_10_426_3047_0,
    i_10_426_3160_0, i_10_426_3200_0, i_10_426_3267_0, i_10_426_3271_0,
    i_10_426_3358_0, i_10_426_3384_0, i_10_426_3389_0, i_10_426_3402_0,
    i_10_426_3403_0, i_10_426_3404_0, i_10_426_3611_0, i_10_426_3613_0,
    i_10_426_3648_0, i_10_426_3682_0, i_10_426_3785_0, i_10_426_3808_0,
    i_10_426_3837_0, i_10_426_3843_0, i_10_426_3852_0, i_10_426_3859_0,
    i_10_426_3899_0, i_10_426_4171_0, i_10_426_4212_0, i_10_426_4276_0;
  output o_10_426_0_0;
  assign o_10_426_0_0 = 0;
endmodule



// Benchmark "kernel_10_427" written by ABC on Sun Jul 19 10:28:29 2020

module kernel_10_427 ( 
    i_10_427_171_0, i_10_427_243_0, i_10_427_282_0, i_10_427_284_0,
    i_10_427_392_0, i_10_427_425_0, i_10_427_434_0, i_10_427_442_0,
    i_10_427_464_0, i_10_427_748_0, i_10_427_957_0, i_10_427_958_0,
    i_10_427_961_0, i_10_427_1000_0, i_10_427_1003_0, i_10_427_1084_0,
    i_10_427_1307_0, i_10_427_1311_0, i_10_427_1362_0, i_10_427_1378_0,
    i_10_427_1450_0, i_10_427_1451_0, i_10_427_1551_0, i_10_427_1583_0,
    i_10_427_1633_0, i_10_427_1652_0, i_10_427_1653_0, i_10_427_1655_0,
    i_10_427_1686_0, i_10_427_1820_0, i_10_427_1945_0, i_10_427_1946_0,
    i_10_427_1948_0, i_10_427_1949_0, i_10_427_1990_0, i_10_427_1991_0,
    i_10_427_1994_0, i_10_427_2092_0, i_10_427_2201_0, i_10_427_2305_0,
    i_10_427_2306_0, i_10_427_2310_0, i_10_427_2311_0, i_10_427_2324_0,
    i_10_427_2350_0, i_10_427_2351_0, i_10_427_2354_0, i_10_427_2376_0,
    i_10_427_2377_0, i_10_427_2407_0, i_10_427_2449_0, i_10_427_2450_0,
    i_10_427_2506_0, i_10_427_2611_0, i_10_427_2612_0, i_10_427_2634_0,
    i_10_427_2635_0, i_10_427_2656_0, i_10_427_2658_0, i_10_427_2659_0,
    i_10_427_2663_0, i_10_427_2673_0, i_10_427_2674_0, i_10_427_2675_0,
    i_10_427_2703_0, i_10_427_2728_0, i_10_427_2729_0, i_10_427_2827_0,
    i_10_427_2833_0, i_10_427_3037_0, i_10_427_3038_0, i_10_427_3072_0,
    i_10_427_3087_0, i_10_427_3088_0, i_10_427_3089_0, i_10_427_3195_0,
    i_10_427_3270_0, i_10_427_3286_0, i_10_427_3350_0, i_10_427_3384_0,
    i_10_427_3448_0, i_10_427_3542_0, i_10_427_3614_0, i_10_427_3616_0,
    i_10_427_3786_0, i_10_427_3788_0, i_10_427_3838_0, i_10_427_3839_0,
    i_10_427_3857_0, i_10_427_3880_0, i_10_427_3944_0, i_10_427_4006_0,
    i_10_427_4024_0, i_10_427_4113_0, i_10_427_4219_0, i_10_427_4268_0,
    i_10_427_4286_0, i_10_427_4289_0, i_10_427_4474_0, i_10_427_4591_0,
    o_10_427_0_0  );
  input  i_10_427_171_0, i_10_427_243_0, i_10_427_282_0, i_10_427_284_0,
    i_10_427_392_0, i_10_427_425_0, i_10_427_434_0, i_10_427_442_0,
    i_10_427_464_0, i_10_427_748_0, i_10_427_957_0, i_10_427_958_0,
    i_10_427_961_0, i_10_427_1000_0, i_10_427_1003_0, i_10_427_1084_0,
    i_10_427_1307_0, i_10_427_1311_0, i_10_427_1362_0, i_10_427_1378_0,
    i_10_427_1450_0, i_10_427_1451_0, i_10_427_1551_0, i_10_427_1583_0,
    i_10_427_1633_0, i_10_427_1652_0, i_10_427_1653_0, i_10_427_1655_0,
    i_10_427_1686_0, i_10_427_1820_0, i_10_427_1945_0, i_10_427_1946_0,
    i_10_427_1948_0, i_10_427_1949_0, i_10_427_1990_0, i_10_427_1991_0,
    i_10_427_1994_0, i_10_427_2092_0, i_10_427_2201_0, i_10_427_2305_0,
    i_10_427_2306_0, i_10_427_2310_0, i_10_427_2311_0, i_10_427_2324_0,
    i_10_427_2350_0, i_10_427_2351_0, i_10_427_2354_0, i_10_427_2376_0,
    i_10_427_2377_0, i_10_427_2407_0, i_10_427_2449_0, i_10_427_2450_0,
    i_10_427_2506_0, i_10_427_2611_0, i_10_427_2612_0, i_10_427_2634_0,
    i_10_427_2635_0, i_10_427_2656_0, i_10_427_2658_0, i_10_427_2659_0,
    i_10_427_2663_0, i_10_427_2673_0, i_10_427_2674_0, i_10_427_2675_0,
    i_10_427_2703_0, i_10_427_2728_0, i_10_427_2729_0, i_10_427_2827_0,
    i_10_427_2833_0, i_10_427_3037_0, i_10_427_3038_0, i_10_427_3072_0,
    i_10_427_3087_0, i_10_427_3088_0, i_10_427_3089_0, i_10_427_3195_0,
    i_10_427_3270_0, i_10_427_3286_0, i_10_427_3350_0, i_10_427_3384_0,
    i_10_427_3448_0, i_10_427_3542_0, i_10_427_3614_0, i_10_427_3616_0,
    i_10_427_3786_0, i_10_427_3788_0, i_10_427_3838_0, i_10_427_3839_0,
    i_10_427_3857_0, i_10_427_3880_0, i_10_427_3944_0, i_10_427_4006_0,
    i_10_427_4024_0, i_10_427_4113_0, i_10_427_4219_0, i_10_427_4268_0,
    i_10_427_4286_0, i_10_427_4289_0, i_10_427_4474_0, i_10_427_4591_0;
  output o_10_427_0_0;
  assign o_10_427_0_0 = 0;
endmodule



// Benchmark "kernel_10_428" written by ABC on Sun Jul 19 10:28:30 2020

module kernel_10_428 ( 
    i_10_428_19_0, i_10_428_33_0, i_10_428_35_0, i_10_428_69_0,
    i_10_428_393_0, i_10_428_426_0, i_10_428_427_0, i_10_428_429_0,
    i_10_428_467_0, i_10_428_534_0, i_10_428_535_0, i_10_428_538_0,
    i_10_428_539_0, i_10_428_642_0, i_10_428_948_0, i_10_428_1007_0,
    i_10_428_1039_0, i_10_428_1187_0, i_10_428_1200_0, i_10_428_1263_0,
    i_10_428_1305_0, i_10_428_1317_0, i_10_428_1320_0, i_10_428_1321_0,
    i_10_428_1342_0, i_10_428_1348_0, i_10_428_1413_0, i_10_428_1425_0,
    i_10_428_1444_0, i_10_428_1446_0, i_10_428_1447_0, i_10_428_1544_0,
    i_10_428_1552_0, i_10_428_1605_0, i_10_428_1617_0, i_10_428_1648_0,
    i_10_428_1713_0, i_10_428_1761_0, i_10_428_1912_0, i_10_428_1993_0,
    i_10_428_2291_0, i_10_428_2355_0, i_10_428_2436_0, i_10_428_2448_0,
    i_10_428_2556_0, i_10_428_2826_0, i_10_428_2834_0, i_10_428_2880_0,
    i_10_428_2881_0, i_10_428_2917_0, i_10_428_2919_0, i_10_428_2920_0,
    i_10_428_2922_0, i_10_428_2923_0, i_10_428_3034_0, i_10_428_3039_0,
    i_10_428_3040_0, i_10_428_3043_0, i_10_428_3087_0, i_10_428_3090_0,
    i_10_428_3091_0, i_10_428_3093_0, i_10_428_3094_0, i_10_428_3130_0,
    i_10_428_3268_0, i_10_428_3270_0, i_10_428_3279_0, i_10_428_3280_0,
    i_10_428_3283_0, i_10_428_3321_0, i_10_428_3384_0, i_10_428_3408_0,
    i_10_428_3409_0, i_10_428_3436_0, i_10_428_3495_0, i_10_428_3520_0,
    i_10_428_3523_0, i_10_428_3544_0, i_10_428_3609_0, i_10_428_3612_0,
    i_10_428_3615_0, i_10_428_3724_0, i_10_428_3734_0, i_10_428_3816_0,
    i_10_428_3832_0, i_10_428_3855_0, i_10_428_3856_0, i_10_428_3895_0,
    i_10_428_3898_0, i_10_428_4120_0, i_10_428_4121_0, i_10_428_4209_0,
    i_10_428_4219_0, i_10_428_4351_0, i_10_428_4411_0, i_10_428_4458_0,
    i_10_428_4557_0, i_10_428_4569_0, i_10_428_4593_0, i_10_428_4597_0,
    o_10_428_0_0  );
  input  i_10_428_19_0, i_10_428_33_0, i_10_428_35_0, i_10_428_69_0,
    i_10_428_393_0, i_10_428_426_0, i_10_428_427_0, i_10_428_429_0,
    i_10_428_467_0, i_10_428_534_0, i_10_428_535_0, i_10_428_538_0,
    i_10_428_539_0, i_10_428_642_0, i_10_428_948_0, i_10_428_1007_0,
    i_10_428_1039_0, i_10_428_1187_0, i_10_428_1200_0, i_10_428_1263_0,
    i_10_428_1305_0, i_10_428_1317_0, i_10_428_1320_0, i_10_428_1321_0,
    i_10_428_1342_0, i_10_428_1348_0, i_10_428_1413_0, i_10_428_1425_0,
    i_10_428_1444_0, i_10_428_1446_0, i_10_428_1447_0, i_10_428_1544_0,
    i_10_428_1552_0, i_10_428_1605_0, i_10_428_1617_0, i_10_428_1648_0,
    i_10_428_1713_0, i_10_428_1761_0, i_10_428_1912_0, i_10_428_1993_0,
    i_10_428_2291_0, i_10_428_2355_0, i_10_428_2436_0, i_10_428_2448_0,
    i_10_428_2556_0, i_10_428_2826_0, i_10_428_2834_0, i_10_428_2880_0,
    i_10_428_2881_0, i_10_428_2917_0, i_10_428_2919_0, i_10_428_2920_0,
    i_10_428_2922_0, i_10_428_2923_0, i_10_428_3034_0, i_10_428_3039_0,
    i_10_428_3040_0, i_10_428_3043_0, i_10_428_3087_0, i_10_428_3090_0,
    i_10_428_3091_0, i_10_428_3093_0, i_10_428_3094_0, i_10_428_3130_0,
    i_10_428_3268_0, i_10_428_3270_0, i_10_428_3279_0, i_10_428_3280_0,
    i_10_428_3283_0, i_10_428_3321_0, i_10_428_3384_0, i_10_428_3408_0,
    i_10_428_3409_0, i_10_428_3436_0, i_10_428_3495_0, i_10_428_3520_0,
    i_10_428_3523_0, i_10_428_3544_0, i_10_428_3609_0, i_10_428_3612_0,
    i_10_428_3615_0, i_10_428_3724_0, i_10_428_3734_0, i_10_428_3816_0,
    i_10_428_3832_0, i_10_428_3855_0, i_10_428_3856_0, i_10_428_3895_0,
    i_10_428_3898_0, i_10_428_4120_0, i_10_428_4121_0, i_10_428_4209_0,
    i_10_428_4219_0, i_10_428_4351_0, i_10_428_4411_0, i_10_428_4458_0,
    i_10_428_4557_0, i_10_428_4569_0, i_10_428_4593_0, i_10_428_4597_0;
  output o_10_428_0_0;
  assign o_10_428_0_0 = 0;
endmodule



// Benchmark "kernel_10_429" written by ABC on Sun Jul 19 10:28:31 2020

module kernel_10_429 ( 
    i_10_429_89_0, i_10_429_121_0, i_10_429_122_0, i_10_429_156_0,
    i_10_429_157_0, i_10_429_174_0, i_10_429_175_0, i_10_429_177_0,
    i_10_429_185_0, i_10_429_248_0, i_10_429_280_0, i_10_429_287_0,
    i_10_429_388_0, i_10_429_391_0, i_10_429_392_0, i_10_429_410_0,
    i_10_429_445_0, i_10_429_446_0, i_10_429_561_0, i_10_429_629_0,
    i_10_429_795_0, i_10_429_1005_0, i_10_429_1084_0, i_10_429_1305_0,
    i_10_429_1308_0, i_10_429_1432_0, i_10_429_1433_0, i_10_429_1439_0,
    i_10_429_1489_0, i_10_429_1552_0, i_10_429_1578_0, i_10_429_1579_0,
    i_10_429_1650_0, i_10_429_1689_0, i_10_429_1726_0, i_10_429_1771_0,
    i_10_429_1795_0, i_10_429_1796_0, i_10_429_1952_0, i_10_429_2001_0,
    i_10_429_2246_0, i_10_429_2356_0, i_10_429_2357_0, i_10_429_2365_0,
    i_10_429_2403_0, i_10_429_2407_0, i_10_429_2410_0, i_10_429_2446_0,
    i_10_429_2447_0, i_10_429_2453_0, i_10_429_2472_0, i_10_429_2519_0,
    i_10_429_2615_0, i_10_429_2634_0, i_10_429_2643_0, i_10_429_2644_0,
    i_10_429_2731_0, i_10_429_2733_0, i_10_429_2734_0, i_10_429_2735_0,
    i_10_429_2744_0, i_10_429_2829_0, i_10_429_2830_0, i_10_429_2869_0,
    i_10_429_2885_0, i_10_429_2916_0, i_10_429_3235_0, i_10_429_3279_0,
    i_10_429_3280_0, i_10_429_3281_0, i_10_429_3283_0, i_10_429_3284_0,
    i_10_429_3298_0, i_10_429_3299_0, i_10_429_3318_0, i_10_429_3390_0,
    i_10_429_3466_0, i_10_429_3583_0, i_10_429_3614_0, i_10_429_3705_0,
    i_10_429_3729_0, i_10_429_3837_0, i_10_429_3841_0, i_10_429_3860_0,
    i_10_429_3923_0, i_10_429_3981_0, i_10_429_3984_0, i_10_429_3985_0,
    i_10_429_3986_0, i_10_429_4026_0, i_10_429_4028_0, i_10_429_4056_0,
    i_10_429_4120_0, i_10_429_4129_0, i_10_429_4172_0, i_10_429_4175_0,
    i_10_429_4266_0, i_10_429_4267_0, i_10_429_4282_0, i_10_429_4302_0,
    o_10_429_0_0  );
  input  i_10_429_89_0, i_10_429_121_0, i_10_429_122_0, i_10_429_156_0,
    i_10_429_157_0, i_10_429_174_0, i_10_429_175_0, i_10_429_177_0,
    i_10_429_185_0, i_10_429_248_0, i_10_429_280_0, i_10_429_287_0,
    i_10_429_388_0, i_10_429_391_0, i_10_429_392_0, i_10_429_410_0,
    i_10_429_445_0, i_10_429_446_0, i_10_429_561_0, i_10_429_629_0,
    i_10_429_795_0, i_10_429_1005_0, i_10_429_1084_0, i_10_429_1305_0,
    i_10_429_1308_0, i_10_429_1432_0, i_10_429_1433_0, i_10_429_1439_0,
    i_10_429_1489_0, i_10_429_1552_0, i_10_429_1578_0, i_10_429_1579_0,
    i_10_429_1650_0, i_10_429_1689_0, i_10_429_1726_0, i_10_429_1771_0,
    i_10_429_1795_0, i_10_429_1796_0, i_10_429_1952_0, i_10_429_2001_0,
    i_10_429_2246_0, i_10_429_2356_0, i_10_429_2357_0, i_10_429_2365_0,
    i_10_429_2403_0, i_10_429_2407_0, i_10_429_2410_0, i_10_429_2446_0,
    i_10_429_2447_0, i_10_429_2453_0, i_10_429_2472_0, i_10_429_2519_0,
    i_10_429_2615_0, i_10_429_2634_0, i_10_429_2643_0, i_10_429_2644_0,
    i_10_429_2731_0, i_10_429_2733_0, i_10_429_2734_0, i_10_429_2735_0,
    i_10_429_2744_0, i_10_429_2829_0, i_10_429_2830_0, i_10_429_2869_0,
    i_10_429_2885_0, i_10_429_2916_0, i_10_429_3235_0, i_10_429_3279_0,
    i_10_429_3280_0, i_10_429_3281_0, i_10_429_3283_0, i_10_429_3284_0,
    i_10_429_3298_0, i_10_429_3299_0, i_10_429_3318_0, i_10_429_3390_0,
    i_10_429_3466_0, i_10_429_3583_0, i_10_429_3614_0, i_10_429_3705_0,
    i_10_429_3729_0, i_10_429_3837_0, i_10_429_3841_0, i_10_429_3860_0,
    i_10_429_3923_0, i_10_429_3981_0, i_10_429_3984_0, i_10_429_3985_0,
    i_10_429_3986_0, i_10_429_4026_0, i_10_429_4028_0, i_10_429_4056_0,
    i_10_429_4120_0, i_10_429_4129_0, i_10_429_4172_0, i_10_429_4175_0,
    i_10_429_4266_0, i_10_429_4267_0, i_10_429_4282_0, i_10_429_4302_0;
  output o_10_429_0_0;
  assign o_10_429_0_0 = 0;
endmodule



// Benchmark "kernel_10_430" written by ABC on Sun Jul 19 10:28:32 2020

module kernel_10_430 ( 
    i_10_430_50_0, i_10_430_172_0, i_10_430_179_0, i_10_430_217_0,
    i_10_430_218_0, i_10_430_220_0, i_10_430_263_0, i_10_430_287_0,
    i_10_430_325_0, i_10_430_327_0, i_10_430_328_0, i_10_430_392_0,
    i_10_430_500_0, i_10_430_509_0, i_10_430_1000_0, i_10_430_1001_0,
    i_10_430_1030_0, i_10_430_1031_0, i_10_430_1040_0, i_10_430_1088_0,
    i_10_430_1102_0, i_10_430_1234_0, i_10_430_1238_0, i_10_430_1239_0,
    i_10_430_1262_0, i_10_430_1431_0, i_10_430_1433_0, i_10_430_1540_0,
    i_10_430_1578_0, i_10_430_1634_0, i_10_430_1643_0, i_10_430_1651_0,
    i_10_430_1652_0, i_10_430_1654_0, i_10_430_1688_0, i_10_430_1691_0,
    i_10_430_1730_0, i_10_430_1769_0, i_10_430_1820_0, i_10_430_1822_0,
    i_10_430_1982_0, i_10_430_2003_0, i_10_430_2006_0, i_10_430_2030_0,
    i_10_430_2198_0, i_10_430_2201_0, i_10_430_2204_0, i_10_430_2246_0,
    i_10_430_2255_0, i_10_430_2354_0, i_10_430_2364_0, i_10_430_2449_0,
    i_10_430_2450_0, i_10_430_2451_0, i_10_430_2452_0, i_10_430_2455_0,
    i_10_430_2468_0, i_10_430_2474_0, i_10_430_2567_0, i_10_430_2632_0,
    i_10_430_2636_0, i_10_430_2702_0, i_10_430_2704_0, i_10_430_2711_0,
    i_10_430_2714_0, i_10_430_2720_0, i_10_430_2732_0, i_10_430_2733_0,
    i_10_430_2741_0, i_10_430_2825_0, i_10_430_2830_0, i_10_430_2916_0,
    i_10_430_2966_0, i_10_430_3044_0, i_10_430_3071_0, i_10_430_3072_0,
    i_10_430_3268_0, i_10_430_3281_0, i_10_430_3314_0, i_10_430_3317_0,
    i_10_430_3389_0, i_10_430_3390_0, i_10_430_3391_0, i_10_430_3467_0,
    i_10_430_3473_0, i_10_430_3503_0, i_10_430_3506_0, i_10_430_3509_0,
    i_10_430_3584_0, i_10_430_3590_0, i_10_430_3841_0, i_10_430_3848_0,
    i_10_430_4028_0, i_10_430_4121_0, i_10_430_4123_0, i_10_430_4268_0,
    i_10_430_4283_0, i_10_430_4292_0, i_10_430_4565_0, i_10_430_4566_0,
    o_10_430_0_0  );
  input  i_10_430_50_0, i_10_430_172_0, i_10_430_179_0, i_10_430_217_0,
    i_10_430_218_0, i_10_430_220_0, i_10_430_263_0, i_10_430_287_0,
    i_10_430_325_0, i_10_430_327_0, i_10_430_328_0, i_10_430_392_0,
    i_10_430_500_0, i_10_430_509_0, i_10_430_1000_0, i_10_430_1001_0,
    i_10_430_1030_0, i_10_430_1031_0, i_10_430_1040_0, i_10_430_1088_0,
    i_10_430_1102_0, i_10_430_1234_0, i_10_430_1238_0, i_10_430_1239_0,
    i_10_430_1262_0, i_10_430_1431_0, i_10_430_1433_0, i_10_430_1540_0,
    i_10_430_1578_0, i_10_430_1634_0, i_10_430_1643_0, i_10_430_1651_0,
    i_10_430_1652_0, i_10_430_1654_0, i_10_430_1688_0, i_10_430_1691_0,
    i_10_430_1730_0, i_10_430_1769_0, i_10_430_1820_0, i_10_430_1822_0,
    i_10_430_1982_0, i_10_430_2003_0, i_10_430_2006_0, i_10_430_2030_0,
    i_10_430_2198_0, i_10_430_2201_0, i_10_430_2204_0, i_10_430_2246_0,
    i_10_430_2255_0, i_10_430_2354_0, i_10_430_2364_0, i_10_430_2449_0,
    i_10_430_2450_0, i_10_430_2451_0, i_10_430_2452_0, i_10_430_2455_0,
    i_10_430_2468_0, i_10_430_2474_0, i_10_430_2567_0, i_10_430_2632_0,
    i_10_430_2636_0, i_10_430_2702_0, i_10_430_2704_0, i_10_430_2711_0,
    i_10_430_2714_0, i_10_430_2720_0, i_10_430_2732_0, i_10_430_2733_0,
    i_10_430_2741_0, i_10_430_2825_0, i_10_430_2830_0, i_10_430_2916_0,
    i_10_430_2966_0, i_10_430_3044_0, i_10_430_3071_0, i_10_430_3072_0,
    i_10_430_3268_0, i_10_430_3281_0, i_10_430_3314_0, i_10_430_3317_0,
    i_10_430_3389_0, i_10_430_3390_0, i_10_430_3391_0, i_10_430_3467_0,
    i_10_430_3473_0, i_10_430_3503_0, i_10_430_3506_0, i_10_430_3509_0,
    i_10_430_3584_0, i_10_430_3590_0, i_10_430_3841_0, i_10_430_3848_0,
    i_10_430_4028_0, i_10_430_4121_0, i_10_430_4123_0, i_10_430_4268_0,
    i_10_430_4283_0, i_10_430_4292_0, i_10_430_4565_0, i_10_430_4566_0;
  output o_10_430_0_0;
  assign o_10_430_0_0 = 0;
endmodule



// Benchmark "kernel_10_431" written by ABC on Sun Jul 19 10:28:33 2020

module kernel_10_431 ( 
    i_10_431_27_0, i_10_431_148_0, i_10_431_180_0, i_10_431_181_0,
    i_10_431_217_0, i_10_431_221_0, i_10_431_244_0, i_10_431_245_0,
    i_10_431_257_0, i_10_431_280_0, i_10_431_284_0, i_10_431_289_0,
    i_10_431_405_0, i_10_431_407_0, i_10_431_408_0, i_10_431_409_0,
    i_10_431_463_0, i_10_431_516_0, i_10_431_517_0, i_10_431_715_0,
    i_10_431_716_0, i_10_431_748_0, i_10_431_796_0, i_10_431_1009_0,
    i_10_431_1027_0, i_10_431_1028_0, i_10_431_1030_0, i_10_431_1085_0,
    i_10_431_1233_0, i_10_431_1234_0, i_10_431_1243_0, i_10_431_1246_0,
    i_10_431_1247_0, i_10_431_1539_0, i_10_431_1540_0, i_10_431_1550_0,
    i_10_431_1684_0, i_10_431_1685_0, i_10_431_1687_0, i_10_431_1729_0,
    i_10_431_1730_0, i_10_431_1801_0, i_10_431_1818_0, i_10_431_1821_0,
    i_10_431_1912_0, i_10_431_1999_0, i_10_431_2179_0, i_10_431_2288_0,
    i_10_431_2349_0, i_10_431_2353_0, i_10_431_2449_0, i_10_431_2450_0,
    i_10_431_2457_0, i_10_431_2470_0, i_10_431_2511_0, i_10_431_2543_0,
    i_10_431_2601_0, i_10_431_2604_0, i_10_431_2631_0, i_10_431_2660_0,
    i_10_431_2675_0, i_10_431_2728_0, i_10_431_3043_0, i_10_431_3069_0,
    i_10_431_3070_0, i_10_431_3198_0, i_10_431_3199_0, i_10_431_3200_0,
    i_10_431_3268_0, i_10_431_3386_0, i_10_431_3555_0, i_10_431_3583_0,
    i_10_431_3584_0, i_10_431_3587_0, i_10_431_3613_0, i_10_431_3618_0,
    i_10_431_3619_0, i_10_431_3650_0, i_10_431_3682_0, i_10_431_3785_0,
    i_10_431_3838_0, i_10_431_3856_0, i_10_431_3871_0, i_10_431_3946_0,
    i_10_431_3995_0, i_10_431_4010_0, i_10_431_4024_0, i_10_431_4025_0,
    i_10_431_4113_0, i_10_431_4114_0, i_10_431_4168_0, i_10_431_4213_0,
    i_10_431_4216_0, i_10_431_4267_0, i_10_431_4275_0, i_10_431_4276_0,
    i_10_431_4279_0, i_10_431_4285_0, i_10_431_4288_0, i_10_431_4568_0,
    o_10_431_0_0  );
  input  i_10_431_27_0, i_10_431_148_0, i_10_431_180_0, i_10_431_181_0,
    i_10_431_217_0, i_10_431_221_0, i_10_431_244_0, i_10_431_245_0,
    i_10_431_257_0, i_10_431_280_0, i_10_431_284_0, i_10_431_289_0,
    i_10_431_405_0, i_10_431_407_0, i_10_431_408_0, i_10_431_409_0,
    i_10_431_463_0, i_10_431_516_0, i_10_431_517_0, i_10_431_715_0,
    i_10_431_716_0, i_10_431_748_0, i_10_431_796_0, i_10_431_1009_0,
    i_10_431_1027_0, i_10_431_1028_0, i_10_431_1030_0, i_10_431_1085_0,
    i_10_431_1233_0, i_10_431_1234_0, i_10_431_1243_0, i_10_431_1246_0,
    i_10_431_1247_0, i_10_431_1539_0, i_10_431_1540_0, i_10_431_1550_0,
    i_10_431_1684_0, i_10_431_1685_0, i_10_431_1687_0, i_10_431_1729_0,
    i_10_431_1730_0, i_10_431_1801_0, i_10_431_1818_0, i_10_431_1821_0,
    i_10_431_1912_0, i_10_431_1999_0, i_10_431_2179_0, i_10_431_2288_0,
    i_10_431_2349_0, i_10_431_2353_0, i_10_431_2449_0, i_10_431_2450_0,
    i_10_431_2457_0, i_10_431_2470_0, i_10_431_2511_0, i_10_431_2543_0,
    i_10_431_2601_0, i_10_431_2604_0, i_10_431_2631_0, i_10_431_2660_0,
    i_10_431_2675_0, i_10_431_2728_0, i_10_431_3043_0, i_10_431_3069_0,
    i_10_431_3070_0, i_10_431_3198_0, i_10_431_3199_0, i_10_431_3200_0,
    i_10_431_3268_0, i_10_431_3386_0, i_10_431_3555_0, i_10_431_3583_0,
    i_10_431_3584_0, i_10_431_3587_0, i_10_431_3613_0, i_10_431_3618_0,
    i_10_431_3619_0, i_10_431_3650_0, i_10_431_3682_0, i_10_431_3785_0,
    i_10_431_3838_0, i_10_431_3856_0, i_10_431_3871_0, i_10_431_3946_0,
    i_10_431_3995_0, i_10_431_4010_0, i_10_431_4024_0, i_10_431_4025_0,
    i_10_431_4113_0, i_10_431_4114_0, i_10_431_4168_0, i_10_431_4213_0,
    i_10_431_4216_0, i_10_431_4267_0, i_10_431_4275_0, i_10_431_4276_0,
    i_10_431_4279_0, i_10_431_4285_0, i_10_431_4288_0, i_10_431_4568_0;
  output o_10_431_0_0;
  assign o_10_431_0_0 = 0;
endmodule



// Benchmark "kernel_10_432" written by ABC on Sun Jul 19 10:28:34 2020

module kernel_10_432 ( 
    i_10_432_30_0, i_10_432_40_0, i_10_432_123_0, i_10_432_124_0,
    i_10_432_180_0, i_10_432_184_0, i_10_432_186_0, i_10_432_286_0,
    i_10_432_316_0, i_10_432_318_0, i_10_432_393_0, i_10_432_440_0,
    i_10_432_449_0, i_10_432_463_0, i_10_432_465_0, i_10_432_466_0,
    i_10_432_799_0, i_10_432_1137_0, i_10_432_1233_0, i_10_432_1234_0,
    i_10_432_1236_0, i_10_432_1237_0, i_10_432_1239_0, i_10_432_1240_0,
    i_10_432_1248_0, i_10_432_1361_0, i_10_432_1362_0, i_10_432_1363_0,
    i_10_432_1364_0, i_10_432_1365_0, i_10_432_1546_0, i_10_432_1552_0,
    i_10_432_1617_0, i_10_432_1680_0, i_10_432_1686_0, i_10_432_1688_0,
    i_10_432_1820_0, i_10_432_1821_0, i_10_432_1822_0, i_10_432_1947_0,
    i_10_432_1950_0, i_10_432_2355_0, i_10_432_2408_0, i_10_432_2450_0,
    i_10_432_2453_0, i_10_432_2565_0, i_10_432_2631_0, i_10_432_2636_0,
    i_10_432_2656_0, i_10_432_2679_0, i_10_432_2713_0, i_10_432_2719_0,
    i_10_432_2723_0, i_10_432_2727_0, i_10_432_2730_0, i_10_432_2828_0,
    i_10_432_2830_0, i_10_432_2832_0, i_10_432_2880_0, i_10_432_2980_0,
    i_10_432_3035_0, i_10_432_3036_0, i_10_432_3037_0, i_10_432_3039_0,
    i_10_432_3040_0, i_10_432_3048_0, i_10_432_3093_0, i_10_432_3195_0,
    i_10_432_3196_0, i_10_432_3198_0, i_10_432_3276_0, i_10_432_3278_0,
    i_10_432_3279_0, i_10_432_3284_0, i_10_432_3322_0, i_10_432_3325_0,
    i_10_432_3385_0, i_10_432_3386_0, i_10_432_3387_0, i_10_432_3388_0,
    i_10_432_3391_0, i_10_432_3406_0, i_10_432_3430_0, i_10_432_3468_0,
    i_10_432_3522_0, i_10_432_3586_0, i_10_432_3648_0, i_10_432_3649_0,
    i_10_432_3651_0, i_10_432_3681_0, i_10_432_3781_0, i_10_432_3839_0,
    i_10_432_3855_0, i_10_432_3882_0, i_10_432_3894_0, i_10_432_4053_0,
    i_10_432_4056_0, i_10_432_4274_0, i_10_432_4569_0, i_10_432_4570_0,
    o_10_432_0_0  );
  input  i_10_432_30_0, i_10_432_40_0, i_10_432_123_0, i_10_432_124_0,
    i_10_432_180_0, i_10_432_184_0, i_10_432_186_0, i_10_432_286_0,
    i_10_432_316_0, i_10_432_318_0, i_10_432_393_0, i_10_432_440_0,
    i_10_432_449_0, i_10_432_463_0, i_10_432_465_0, i_10_432_466_0,
    i_10_432_799_0, i_10_432_1137_0, i_10_432_1233_0, i_10_432_1234_0,
    i_10_432_1236_0, i_10_432_1237_0, i_10_432_1239_0, i_10_432_1240_0,
    i_10_432_1248_0, i_10_432_1361_0, i_10_432_1362_0, i_10_432_1363_0,
    i_10_432_1364_0, i_10_432_1365_0, i_10_432_1546_0, i_10_432_1552_0,
    i_10_432_1617_0, i_10_432_1680_0, i_10_432_1686_0, i_10_432_1688_0,
    i_10_432_1820_0, i_10_432_1821_0, i_10_432_1822_0, i_10_432_1947_0,
    i_10_432_1950_0, i_10_432_2355_0, i_10_432_2408_0, i_10_432_2450_0,
    i_10_432_2453_0, i_10_432_2565_0, i_10_432_2631_0, i_10_432_2636_0,
    i_10_432_2656_0, i_10_432_2679_0, i_10_432_2713_0, i_10_432_2719_0,
    i_10_432_2723_0, i_10_432_2727_0, i_10_432_2730_0, i_10_432_2828_0,
    i_10_432_2830_0, i_10_432_2832_0, i_10_432_2880_0, i_10_432_2980_0,
    i_10_432_3035_0, i_10_432_3036_0, i_10_432_3037_0, i_10_432_3039_0,
    i_10_432_3040_0, i_10_432_3048_0, i_10_432_3093_0, i_10_432_3195_0,
    i_10_432_3196_0, i_10_432_3198_0, i_10_432_3276_0, i_10_432_3278_0,
    i_10_432_3279_0, i_10_432_3284_0, i_10_432_3322_0, i_10_432_3325_0,
    i_10_432_3385_0, i_10_432_3386_0, i_10_432_3387_0, i_10_432_3388_0,
    i_10_432_3391_0, i_10_432_3406_0, i_10_432_3430_0, i_10_432_3468_0,
    i_10_432_3522_0, i_10_432_3586_0, i_10_432_3648_0, i_10_432_3649_0,
    i_10_432_3651_0, i_10_432_3681_0, i_10_432_3781_0, i_10_432_3839_0,
    i_10_432_3855_0, i_10_432_3882_0, i_10_432_3894_0, i_10_432_4053_0,
    i_10_432_4056_0, i_10_432_4274_0, i_10_432_4569_0, i_10_432_4570_0;
  output o_10_432_0_0;
  assign o_10_432_0_0 = ~((~i_10_432_318_0 & ((~i_10_432_123_0 & ~i_10_432_180_0 & ~i_10_432_184_0 & ~i_10_432_1362_0 & ~i_10_432_1364_0 & ~i_10_432_1947_0 & i_10_432_3386_0) | (~i_10_432_186_0 & ~i_10_432_1236_0 & ~i_10_432_1365_0 & ~i_10_432_1617_0 & ~i_10_432_2730_0 & ~i_10_432_2830_0 & ~i_10_432_3195_0 & ~i_10_432_3430_0 & ~i_10_432_4053_0 & ~i_10_432_4274_0))) | (~i_10_432_4053_0 & ((~i_10_432_123_0 & ((~i_10_432_180_0 & i_10_432_2408_0 & ~i_10_432_2636_0 & ~i_10_432_3040_0) | (~i_10_432_184_0 & ~i_10_432_1237_0 & ~i_10_432_1365_0 & ~i_10_432_1552_0 & ~i_10_432_3284_0 & ~i_10_432_3681_0))) | (~i_10_432_4570_0 & ((~i_10_432_1248_0 & ((~i_10_432_1236_0 & ~i_10_432_1240_0 & i_10_432_3035_0) | (~i_10_432_2408_0 & ~i_10_432_3093_0 & i_10_432_3388_0 & ~i_10_432_3430_0))) | (~i_10_432_1361_0 & ~i_10_432_1686_0 & ~i_10_432_2355_0 & ~i_10_432_2727_0 & ~i_10_432_3198_0 & i_10_432_3649_0 & ~i_10_432_4056_0))) | (~i_10_432_2679_0 & ((~i_10_432_124_0 & ~i_10_432_184_0 & ~i_10_432_1364_0 & ~i_10_432_3036_0 & ~i_10_432_3048_0 & ~i_10_432_3681_0) | (i_10_432_2355_0 & ~i_10_432_2880_0 & i_10_432_3651_0 & ~i_10_432_4274_0))))) | (~i_10_432_4056_0 & ((~i_10_432_3468_0 & ((~i_10_432_180_0 & ~i_10_432_3430_0 & ((~i_10_432_1686_0 & ~i_10_432_2355_0 & ~i_10_432_2828_0 & ~i_10_432_3648_0 & ~i_10_432_3649_0 & ~i_10_432_3781_0) | (~i_10_432_123_0 & ~i_10_432_1363_0 & ~i_10_432_1365_0 & ~i_10_432_3195_0 & ~i_10_432_3279_0 & ~i_10_432_3284_0 & ~i_10_432_3385_0 & i_10_432_3648_0 & ~i_10_432_4274_0 & ~i_10_432_4569_0))) | (~i_10_432_1234_0 & ~i_10_432_1363_0 & ~i_10_432_1686_0 & ~i_10_432_3039_0 & ~i_10_432_3651_0 & ~i_10_432_4569_0))) | (~i_10_432_2679_0 & ((~i_10_432_1362_0 & ~i_10_432_2730_0 & i_10_432_2828_0 & ~i_10_432_3839_0) | (~i_10_432_1233_0 & ~i_10_432_1363_0 & ~i_10_432_2830_0 & ~i_10_432_3039_0 & ~i_10_432_3651_0 & ~i_10_432_3894_0))))) | (~i_10_432_1236_0 & ((~i_10_432_1361_0 & ~i_10_432_1617_0 & ~i_10_432_2355_0 & ~i_10_432_2713_0 & ~i_10_432_2719_0 & ~i_10_432_3037_0 & ~i_10_432_3048_0 & ~i_10_432_3468_0) | (i_10_432_2453_0 & ~i_10_432_3648_0 & ~i_10_432_4570_0))) | (~i_10_432_3039_0 & ((~i_10_432_123_0 & ((~i_10_432_1237_0 & ~i_10_432_1821_0 & ~i_10_432_2723_0 & ~i_10_432_2727_0 & ~i_10_432_3040_0) | (i_10_432_1686_0 & ~i_10_432_3855_0))) | (~i_10_432_393_0 & ~i_10_432_799_0 & ~i_10_432_1234_0 & ~i_10_432_1237_0 & ~i_10_432_1947_0))) | (~i_10_432_1234_0 & ~i_10_432_1239_0 & ((~i_10_432_2679_0 & ~i_10_432_2727_0 & ~i_10_432_3649_0 & ~i_10_432_3681_0) | (~i_10_432_123_0 & ~i_10_432_1947_0 & ~i_10_432_3839_0 & ~i_10_432_4569_0))) | (~i_10_432_4570_0 & ((i_10_432_316_0 & ~i_10_432_3037_0) | (i_10_432_318_0 & i_10_432_3385_0))) | i_10_432_2565_0 | (~i_10_432_1363_0 & i_10_432_2980_0 & ~i_10_432_3196_0 & ~i_10_432_3430_0) | (~i_10_432_1233_0 & ~i_10_432_1365_0 & ~i_10_432_2408_0 & ~i_10_432_2730_0 & ~i_10_432_3284_0 & i_10_432_3388_0 & i_10_432_3586_0) | (~i_10_432_1240_0 & i_10_432_1364_0 & i_10_432_2723_0 & ~i_10_432_3894_0));
endmodule



// Benchmark "kernel_10_433" written by ABC on Sun Jul 19 10:28:35 2020

module kernel_10_433 ( 
    i_10_433_135_0, i_10_433_171_0, i_10_433_174_0, i_10_433_177_0,
    i_10_433_258_0, i_10_433_280_0, i_10_433_285_0, i_10_433_286_0,
    i_10_433_316_0, i_10_433_390_0, i_10_433_463_0, i_10_433_467_0,
    i_10_433_687_0, i_10_433_747_0, i_10_433_796_0, i_10_433_1026_0,
    i_10_433_1027_0, i_10_433_1032_0, i_10_433_1236_0, i_10_433_1237_0,
    i_10_433_1238_0, i_10_433_1240_0, i_10_433_1241_0, i_10_433_1245_0,
    i_10_433_1249_0, i_10_433_1250_0, i_10_433_1308_0, i_10_433_1578_0,
    i_10_433_1582_0, i_10_433_1651_0, i_10_433_1684_0, i_10_433_1686_0,
    i_10_433_1691_0, i_10_433_1819_0, i_10_433_1821_0, i_10_433_1822_0,
    i_10_433_2001_0, i_10_433_2199_0, i_10_433_2304_0, i_10_433_2353_0,
    i_10_433_2356_0, i_10_433_2455_0, i_10_433_2460_0, i_10_433_2463_0,
    i_10_433_2467_0, i_10_433_2470_0, i_10_433_2471_0, i_10_433_2473_0,
    i_10_433_2474_0, i_10_433_2514_0, i_10_433_2535_0, i_10_433_2628_0,
    i_10_433_2631_0, i_10_433_2635_0, i_10_433_2655_0, i_10_433_2656_0,
    i_10_433_2658_0, i_10_433_2659_0, i_10_433_2674_0, i_10_433_2710_0,
    i_10_433_2827_0, i_10_433_2829_0, i_10_433_3034_0, i_10_433_3195_0,
    i_10_433_3196_0, i_10_433_3201_0, i_10_433_3202_0, i_10_433_3277_0,
    i_10_433_3387_0, i_10_433_3389_0, i_10_433_3402_0, i_10_433_3438_0,
    i_10_433_3441_0, i_10_433_3585_0, i_10_433_3586_0, i_10_433_3587_0,
    i_10_433_3609_0, i_10_433_3613_0, i_10_433_3614_0, i_10_433_3615_0,
    i_10_433_3783_0, i_10_433_3786_0, i_10_433_3787_0, i_10_433_3838_0,
    i_10_433_3840_0, i_10_433_3852_0, i_10_433_3858_0, i_10_433_3943_0,
    i_10_433_3982_0, i_10_433_4008_0, i_10_433_4113_0, i_10_433_4126_0,
    i_10_433_4169_0, i_10_433_4219_0, i_10_433_4289_0, i_10_433_4291_0,
    i_10_433_4292_0, i_10_433_4567_0, i_10_433_4569_0, i_10_433_4580_0,
    o_10_433_0_0  );
  input  i_10_433_135_0, i_10_433_171_0, i_10_433_174_0, i_10_433_177_0,
    i_10_433_258_0, i_10_433_280_0, i_10_433_285_0, i_10_433_286_0,
    i_10_433_316_0, i_10_433_390_0, i_10_433_463_0, i_10_433_467_0,
    i_10_433_687_0, i_10_433_747_0, i_10_433_796_0, i_10_433_1026_0,
    i_10_433_1027_0, i_10_433_1032_0, i_10_433_1236_0, i_10_433_1237_0,
    i_10_433_1238_0, i_10_433_1240_0, i_10_433_1241_0, i_10_433_1245_0,
    i_10_433_1249_0, i_10_433_1250_0, i_10_433_1308_0, i_10_433_1578_0,
    i_10_433_1582_0, i_10_433_1651_0, i_10_433_1684_0, i_10_433_1686_0,
    i_10_433_1691_0, i_10_433_1819_0, i_10_433_1821_0, i_10_433_1822_0,
    i_10_433_2001_0, i_10_433_2199_0, i_10_433_2304_0, i_10_433_2353_0,
    i_10_433_2356_0, i_10_433_2455_0, i_10_433_2460_0, i_10_433_2463_0,
    i_10_433_2467_0, i_10_433_2470_0, i_10_433_2471_0, i_10_433_2473_0,
    i_10_433_2474_0, i_10_433_2514_0, i_10_433_2535_0, i_10_433_2628_0,
    i_10_433_2631_0, i_10_433_2635_0, i_10_433_2655_0, i_10_433_2656_0,
    i_10_433_2658_0, i_10_433_2659_0, i_10_433_2674_0, i_10_433_2710_0,
    i_10_433_2827_0, i_10_433_2829_0, i_10_433_3034_0, i_10_433_3195_0,
    i_10_433_3196_0, i_10_433_3201_0, i_10_433_3202_0, i_10_433_3277_0,
    i_10_433_3387_0, i_10_433_3389_0, i_10_433_3402_0, i_10_433_3438_0,
    i_10_433_3441_0, i_10_433_3585_0, i_10_433_3586_0, i_10_433_3587_0,
    i_10_433_3609_0, i_10_433_3613_0, i_10_433_3614_0, i_10_433_3615_0,
    i_10_433_3783_0, i_10_433_3786_0, i_10_433_3787_0, i_10_433_3838_0,
    i_10_433_3840_0, i_10_433_3852_0, i_10_433_3858_0, i_10_433_3943_0,
    i_10_433_3982_0, i_10_433_4008_0, i_10_433_4113_0, i_10_433_4126_0,
    i_10_433_4169_0, i_10_433_4219_0, i_10_433_4289_0, i_10_433_4291_0,
    i_10_433_4292_0, i_10_433_4567_0, i_10_433_4569_0, i_10_433_4580_0;
  output o_10_433_0_0;
  assign o_10_433_0_0 = 0;
endmodule



// Benchmark "kernel_10_434" written by ABC on Sun Jul 19 10:28:37 2020

module kernel_10_434 ( 
    i_10_434_171_0, i_10_434_217_0, i_10_434_218_0, i_10_434_219_0,
    i_10_434_220_0, i_10_434_223_0, i_10_434_251_0, i_10_434_278_0,
    i_10_434_296_0, i_10_434_316_0, i_10_434_317_0, i_10_434_328_0,
    i_10_434_329_0, i_10_434_331_0, i_10_434_408_0, i_10_434_411_0,
    i_10_434_412_0, i_10_434_432_0, i_10_434_441_0, i_10_434_445_0,
    i_10_434_449_0, i_10_434_458_0, i_10_434_467_0, i_10_434_507_0,
    i_10_434_793_0, i_10_434_991_0, i_10_434_1046_0, i_10_434_1234_0,
    i_10_434_1243_0, i_10_434_1261_0, i_10_434_1263_0, i_10_434_1264_0,
    i_10_434_1265_0, i_10_434_1267_0, i_10_434_1308_0, i_10_434_1309_0,
    i_10_434_1311_0, i_10_434_1432_0, i_10_434_1577_0, i_10_434_1579_0,
    i_10_434_1721_0, i_10_434_1809_0, i_10_434_1818_0, i_10_434_1824_0,
    i_10_434_1912_0, i_10_434_1915_0, i_10_434_1916_0, i_10_434_1945_0,
    i_10_434_2018_0, i_10_434_2353_0, i_10_434_2355_0, i_10_434_2358_0,
    i_10_434_2632_0, i_10_434_2635_0, i_10_434_2700_0, i_10_434_2702_0,
    i_10_434_2722_0, i_10_434_2788_0, i_10_434_2817_0, i_10_434_2829_0,
    i_10_434_2830_0, i_10_434_2831_0, i_10_434_2833_0, i_10_434_2919_0,
    i_10_434_2920_0, i_10_434_2923_0, i_10_434_3037_0, i_10_434_3043_0,
    i_10_434_3196_0, i_10_434_3203_0, i_10_434_3279_0, i_10_434_3280_0,
    i_10_434_3321_0, i_10_434_3384_0, i_10_434_3385_0, i_10_434_3392_0,
    i_10_434_3470_0, i_10_434_3614_0, i_10_434_3650_0, i_10_434_3720_0,
    i_10_434_3721_0, i_10_434_3781_0, i_10_434_3785_0, i_10_434_3786_0,
    i_10_434_3787_0, i_10_434_3834_0, i_10_434_3839_0, i_10_434_3844_0,
    i_10_434_3849_0, i_10_434_3852_0, i_10_434_3853_0, i_10_434_3855_0,
    i_10_434_3871_0, i_10_434_3895_0, i_10_434_4266_0, i_10_434_4284_0,
    i_10_434_4286_0, i_10_434_4287_0, i_10_434_4288_0, i_10_434_4289_0,
    o_10_434_0_0  );
  input  i_10_434_171_0, i_10_434_217_0, i_10_434_218_0, i_10_434_219_0,
    i_10_434_220_0, i_10_434_223_0, i_10_434_251_0, i_10_434_278_0,
    i_10_434_296_0, i_10_434_316_0, i_10_434_317_0, i_10_434_328_0,
    i_10_434_329_0, i_10_434_331_0, i_10_434_408_0, i_10_434_411_0,
    i_10_434_412_0, i_10_434_432_0, i_10_434_441_0, i_10_434_445_0,
    i_10_434_449_0, i_10_434_458_0, i_10_434_467_0, i_10_434_507_0,
    i_10_434_793_0, i_10_434_991_0, i_10_434_1046_0, i_10_434_1234_0,
    i_10_434_1243_0, i_10_434_1261_0, i_10_434_1263_0, i_10_434_1264_0,
    i_10_434_1265_0, i_10_434_1267_0, i_10_434_1308_0, i_10_434_1309_0,
    i_10_434_1311_0, i_10_434_1432_0, i_10_434_1577_0, i_10_434_1579_0,
    i_10_434_1721_0, i_10_434_1809_0, i_10_434_1818_0, i_10_434_1824_0,
    i_10_434_1912_0, i_10_434_1915_0, i_10_434_1916_0, i_10_434_1945_0,
    i_10_434_2018_0, i_10_434_2353_0, i_10_434_2355_0, i_10_434_2358_0,
    i_10_434_2632_0, i_10_434_2635_0, i_10_434_2700_0, i_10_434_2702_0,
    i_10_434_2722_0, i_10_434_2788_0, i_10_434_2817_0, i_10_434_2829_0,
    i_10_434_2830_0, i_10_434_2831_0, i_10_434_2833_0, i_10_434_2919_0,
    i_10_434_2920_0, i_10_434_2923_0, i_10_434_3037_0, i_10_434_3043_0,
    i_10_434_3196_0, i_10_434_3203_0, i_10_434_3279_0, i_10_434_3280_0,
    i_10_434_3321_0, i_10_434_3384_0, i_10_434_3385_0, i_10_434_3392_0,
    i_10_434_3470_0, i_10_434_3614_0, i_10_434_3650_0, i_10_434_3720_0,
    i_10_434_3721_0, i_10_434_3781_0, i_10_434_3785_0, i_10_434_3786_0,
    i_10_434_3787_0, i_10_434_3834_0, i_10_434_3839_0, i_10_434_3844_0,
    i_10_434_3849_0, i_10_434_3852_0, i_10_434_3853_0, i_10_434_3855_0,
    i_10_434_3871_0, i_10_434_3895_0, i_10_434_4266_0, i_10_434_4284_0,
    i_10_434_4286_0, i_10_434_4287_0, i_10_434_4288_0, i_10_434_4289_0;
  output o_10_434_0_0;
  assign o_10_434_0_0 = ~((~i_10_434_3650_0 & ((~i_10_434_3787_0 & ((~i_10_434_296_0 & ((~i_10_434_328_0 & ~i_10_434_408_0 & ~i_10_434_3203_0 & i_10_434_3280_0 & ~i_10_434_3834_0) | (~i_10_434_1265_0 & ~i_10_434_1267_0 & ~i_10_434_1577_0 & ~i_10_434_2632_0 & ~i_10_434_2635_0 & ~i_10_434_2788_0 & ~i_10_434_2829_0 & ~i_10_434_3839_0))) | (~i_10_434_328_0 & ~i_10_434_408_0 & ~i_10_434_1265_0 & ~i_10_434_1267_0 & ~i_10_434_1311_0 & i_10_434_2635_0 & ~i_10_434_3614_0))) | (~i_10_434_2355_0 & ~i_10_434_2722_0 & ((~i_10_434_329_0 & ~i_10_434_1309_0 & ~i_10_434_2833_0 & ~i_10_434_3785_0) | (~i_10_434_316_0 & ~i_10_434_331_0 & ~i_10_434_411_0 & i_10_434_1309_0 & ~i_10_434_2829_0 & ~i_10_434_3839_0))))) | (~i_10_434_328_0 & ((~i_10_434_316_0 & ((~i_10_434_1915_0 & i_10_434_2700_0 & ~i_10_434_3279_0 & ~i_10_434_3614_0) | (~i_10_434_329_0 & ~i_10_434_411_0 & ~i_10_434_412_0 & ~i_10_434_1311_0 & ~i_10_434_1579_0 & ~i_10_434_2355_0 & ~i_10_434_2788_0 & ~i_10_434_2831_0 & ~i_10_434_3786_0 & ~i_10_434_3895_0 & ~i_10_434_4286_0))) | (~i_10_434_1265_0 & ~i_10_434_1267_0 & ((~i_10_434_991_0 & ~i_10_434_1264_0 & ~i_10_434_1577_0 & ~i_10_434_2722_0 & i_10_434_3196_0) | (~i_10_434_317_0 & ~i_10_434_1263_0 & ~i_10_434_2788_0 & ~i_10_434_2833_0 & ~i_10_434_2920_0 & ~i_10_434_3037_0 & ~i_10_434_3392_0 & ~i_10_434_3614_0 & ~i_10_434_3895_0 & ~i_10_434_4287_0))) | (~i_10_434_251_0 & ~i_10_434_467_0 & ~i_10_434_1308_0 & ~i_10_434_1309_0 & ~i_10_434_1311_0 & ~i_10_434_2702_0 & ~i_10_434_3785_0))) | (~i_10_434_329_0 & ((~i_10_434_251_0 & ~i_10_434_432_0 & ~i_10_434_458_0 & ~i_10_434_1309_0 & ~i_10_434_2018_0 & ~i_10_434_2829_0) | (~i_10_434_412_0 & ~i_10_434_1809_0 & i_10_434_3853_0))) | (~i_10_434_251_0 & ((~i_10_434_458_0 & ((~i_10_434_331_0 & ~i_10_434_1263_0 & ~i_10_434_1915_0 & ~i_10_434_2018_0 & ~i_10_434_2722_0 & ~i_10_434_2830_0 & ~i_10_434_3203_0 & ~i_10_434_3614_0) | (~i_10_434_991_0 & ~i_10_434_1308_0 & ~i_10_434_2831_0 & i_10_434_3614_0 & ~i_10_434_3787_0))) | (~i_10_434_1263_0 & ~i_10_434_2829_0 & ~i_10_434_3785_0 & ((~i_10_434_449_0 & ~i_10_434_991_0 & ~i_10_434_1265_0 & ~i_10_434_1311_0 & ~i_10_434_1809_0 & ~i_10_434_1916_0 & ~i_10_434_2018_0 & ~i_10_434_3385_0 & ~i_10_434_3787_0) | (i_10_434_1308_0 & ~i_10_434_2700_0 & ~i_10_434_2831_0 & ~i_10_434_3203_0 & ~i_10_434_3392_0 & ~i_10_434_3895_0))))) | (~i_10_434_1263_0 & ((i_10_434_449_0 & ~i_10_434_1824_0 & i_10_434_2788_0 & ~i_10_434_2830_0) | (~i_10_434_331_0 & ~i_10_434_3785_0 & i_10_434_4287_0))) | (~i_10_434_331_0 & ((~i_10_434_1809_0 & ~i_10_434_1912_0 & i_10_434_3781_0) | (i_10_434_441_0 & ~i_10_434_1265_0 & ~i_10_434_3280_0 & ~i_10_434_3839_0))) | (~i_10_434_2831_0 & ((~i_10_434_2829_0 & ((~i_10_434_1265_0 & i_10_434_3385_0) | (~i_10_434_1579_0 & ~i_10_434_3280_0 & i_10_434_3839_0 & i_10_434_3855_0))) | (~i_10_434_458_0 & i_10_434_3043_0 & ~i_10_434_3855_0 & ~i_10_434_3895_0))));
endmodule



// Benchmark "kernel_10_435" written by ABC on Sun Jul 19 10:28:38 2020

module kernel_10_435 ( 
    i_10_435_32_0, i_10_435_121_0, i_10_435_254_0, i_10_435_392_0,
    i_10_435_406_0, i_10_435_434_0, i_10_435_440_0, i_10_435_459_0,
    i_10_435_572_0, i_10_435_694_0, i_10_435_739_0, i_10_435_947_0,
    i_10_435_958_0, i_10_435_990_0, i_10_435_991_0, i_10_435_1002_0,
    i_10_435_1003_0, i_10_435_1157_0, i_10_435_1201_0, i_10_435_1207_0,
    i_10_435_1270_0, i_10_435_1312_0, i_10_435_1313_0, i_10_435_1346_0,
    i_10_435_1451_0, i_10_435_1454_0, i_10_435_1544_0, i_10_435_1549_0,
    i_10_435_1550_0, i_10_435_1553_0, i_10_435_1577_0, i_10_435_1580_0,
    i_10_435_1582_0, i_10_435_1622_0, i_10_435_1633_0, i_10_435_1714_0,
    i_10_435_1803_0, i_10_435_1825_0, i_10_435_1876_0, i_10_435_1909_0,
    i_10_435_1985_0, i_10_435_2003_0, i_10_435_2017_0, i_10_435_2024_0,
    i_10_435_2027_0, i_10_435_2153_0, i_10_435_2155_0, i_10_435_2204_0,
    i_10_435_2291_0, i_10_435_2304_0, i_10_435_2309_0, i_10_435_2351_0,
    i_10_435_2384_0, i_10_435_2458_0, i_10_435_2517_0, i_10_435_2567_0,
    i_10_435_2576_0, i_10_435_2585_0, i_10_435_2593_0, i_10_435_2660_0,
    i_10_435_2714_0, i_10_435_2722_0, i_10_435_2724_0, i_10_435_2725_0,
    i_10_435_2729_0, i_10_435_3164_0, i_10_435_3195_0, i_10_435_3196_0,
    i_10_435_3197_0, i_10_435_3232_0, i_10_435_3233_0, i_10_435_3277_0,
    i_10_435_3278_0, i_10_435_3283_0, i_10_435_3385_0, i_10_435_3389_0,
    i_10_435_3403_0, i_10_435_3503_0, i_10_435_3506_0, i_10_435_3524_0,
    i_10_435_3613_0, i_10_435_3614_0, i_10_435_3673_0, i_10_435_3686_0,
    i_10_435_3691_0, i_10_435_3699_0, i_10_435_3700_0, i_10_435_3727_0,
    i_10_435_3812_0, i_10_435_3839_0, i_10_435_3917_0, i_10_435_4010_0,
    i_10_435_4179_0, i_10_435_4268_0, i_10_435_4271_0, i_10_435_4459_0,
    i_10_435_4528_0, i_10_435_4550_0, i_10_435_4586_0, i_10_435_4591_0,
    o_10_435_0_0  );
  input  i_10_435_32_0, i_10_435_121_0, i_10_435_254_0, i_10_435_392_0,
    i_10_435_406_0, i_10_435_434_0, i_10_435_440_0, i_10_435_459_0,
    i_10_435_572_0, i_10_435_694_0, i_10_435_739_0, i_10_435_947_0,
    i_10_435_958_0, i_10_435_990_0, i_10_435_991_0, i_10_435_1002_0,
    i_10_435_1003_0, i_10_435_1157_0, i_10_435_1201_0, i_10_435_1207_0,
    i_10_435_1270_0, i_10_435_1312_0, i_10_435_1313_0, i_10_435_1346_0,
    i_10_435_1451_0, i_10_435_1454_0, i_10_435_1544_0, i_10_435_1549_0,
    i_10_435_1550_0, i_10_435_1553_0, i_10_435_1577_0, i_10_435_1580_0,
    i_10_435_1582_0, i_10_435_1622_0, i_10_435_1633_0, i_10_435_1714_0,
    i_10_435_1803_0, i_10_435_1825_0, i_10_435_1876_0, i_10_435_1909_0,
    i_10_435_1985_0, i_10_435_2003_0, i_10_435_2017_0, i_10_435_2024_0,
    i_10_435_2027_0, i_10_435_2153_0, i_10_435_2155_0, i_10_435_2204_0,
    i_10_435_2291_0, i_10_435_2304_0, i_10_435_2309_0, i_10_435_2351_0,
    i_10_435_2384_0, i_10_435_2458_0, i_10_435_2517_0, i_10_435_2567_0,
    i_10_435_2576_0, i_10_435_2585_0, i_10_435_2593_0, i_10_435_2660_0,
    i_10_435_2714_0, i_10_435_2722_0, i_10_435_2724_0, i_10_435_2725_0,
    i_10_435_2729_0, i_10_435_3164_0, i_10_435_3195_0, i_10_435_3196_0,
    i_10_435_3197_0, i_10_435_3232_0, i_10_435_3233_0, i_10_435_3277_0,
    i_10_435_3278_0, i_10_435_3283_0, i_10_435_3385_0, i_10_435_3389_0,
    i_10_435_3403_0, i_10_435_3503_0, i_10_435_3506_0, i_10_435_3524_0,
    i_10_435_3613_0, i_10_435_3614_0, i_10_435_3673_0, i_10_435_3686_0,
    i_10_435_3691_0, i_10_435_3699_0, i_10_435_3700_0, i_10_435_3727_0,
    i_10_435_3812_0, i_10_435_3839_0, i_10_435_3917_0, i_10_435_4010_0,
    i_10_435_4179_0, i_10_435_4268_0, i_10_435_4271_0, i_10_435_4459_0,
    i_10_435_4528_0, i_10_435_4550_0, i_10_435_4586_0, i_10_435_4591_0;
  output o_10_435_0_0;
  assign o_10_435_0_0 = 0;
endmodule



// Benchmark "kernel_10_436" written by ABC on Sun Jul 19 10:28:38 2020

module kernel_10_436 ( 
    i_10_436_64_0, i_10_436_261_0, i_10_436_286_0, i_10_436_289_0,
    i_10_436_290_0, i_10_436_320_0, i_10_436_323_0, i_10_436_370_0,
    i_10_436_432_0, i_10_436_433_0, i_10_436_442_0, i_10_436_693_0,
    i_10_436_736_0, i_10_436_737_0, i_10_436_756_0, i_10_436_793_0,
    i_10_436_800_0, i_10_436_843_0, i_10_436_844_0, i_10_436_928_0,
    i_10_436_948_0, i_10_436_954_0, i_10_436_1040_0, i_10_436_1045_0,
    i_10_436_1152_0, i_10_436_1192_0, i_10_436_1199_0, i_10_436_1200_0,
    i_10_436_1238_0, i_10_436_1309_0, i_10_436_1350_0, i_10_436_1354_0,
    i_10_436_1355_0, i_10_436_1363_0, i_10_436_1444_0, i_10_436_1555_0,
    i_10_436_1567_0, i_10_436_1630_0, i_10_436_1685_0, i_10_436_1741_0,
    i_10_436_1800_0, i_10_436_1916_0, i_10_436_1989_0, i_10_436_2205_0,
    i_10_436_2206_0, i_10_436_2207_0, i_10_436_2450_0, i_10_436_2467_0,
    i_10_436_2470_0, i_10_436_2479_0, i_10_436_2506_0, i_10_436_2509_0,
    i_10_436_2514_0, i_10_436_2538_0, i_10_436_2566_0, i_10_436_2569_0,
    i_10_436_2647_0, i_10_436_2659_0, i_10_436_2673_0, i_10_436_2674_0,
    i_10_436_2722_0, i_10_436_2882_0, i_10_436_3074_0, i_10_436_3107_0,
    i_10_436_3201_0, i_10_436_3202_0, i_10_436_3267_0, i_10_436_3268_0,
    i_10_436_3297_0, i_10_436_3360_0, i_10_436_3387_0, i_10_436_3389_0,
    i_10_436_3402_0, i_10_436_3403_0, i_10_436_3405_0, i_10_436_3408_0,
    i_10_436_3525_0, i_10_436_3550_0, i_10_436_3551_0, i_10_436_3553_0,
    i_10_436_3582_0, i_10_436_3604_0, i_10_436_3605_0, i_10_436_3611_0,
    i_10_436_3702_0, i_10_436_3854_0, i_10_436_3855_0, i_10_436_3859_0,
    i_10_436_3901_0, i_10_436_3978_0, i_10_436_3982_0, i_10_436_4185_0,
    i_10_436_4213_0, i_10_436_4216_0, i_10_436_4233_0, i_10_436_4278_0,
    i_10_436_4290_0, i_10_436_4375_0, i_10_436_4376_0, i_10_436_4500_0,
    o_10_436_0_0  );
  input  i_10_436_64_0, i_10_436_261_0, i_10_436_286_0, i_10_436_289_0,
    i_10_436_290_0, i_10_436_320_0, i_10_436_323_0, i_10_436_370_0,
    i_10_436_432_0, i_10_436_433_0, i_10_436_442_0, i_10_436_693_0,
    i_10_436_736_0, i_10_436_737_0, i_10_436_756_0, i_10_436_793_0,
    i_10_436_800_0, i_10_436_843_0, i_10_436_844_0, i_10_436_928_0,
    i_10_436_948_0, i_10_436_954_0, i_10_436_1040_0, i_10_436_1045_0,
    i_10_436_1152_0, i_10_436_1192_0, i_10_436_1199_0, i_10_436_1200_0,
    i_10_436_1238_0, i_10_436_1309_0, i_10_436_1350_0, i_10_436_1354_0,
    i_10_436_1355_0, i_10_436_1363_0, i_10_436_1444_0, i_10_436_1555_0,
    i_10_436_1567_0, i_10_436_1630_0, i_10_436_1685_0, i_10_436_1741_0,
    i_10_436_1800_0, i_10_436_1916_0, i_10_436_1989_0, i_10_436_2205_0,
    i_10_436_2206_0, i_10_436_2207_0, i_10_436_2450_0, i_10_436_2467_0,
    i_10_436_2470_0, i_10_436_2479_0, i_10_436_2506_0, i_10_436_2509_0,
    i_10_436_2514_0, i_10_436_2538_0, i_10_436_2566_0, i_10_436_2569_0,
    i_10_436_2647_0, i_10_436_2659_0, i_10_436_2673_0, i_10_436_2674_0,
    i_10_436_2722_0, i_10_436_2882_0, i_10_436_3074_0, i_10_436_3107_0,
    i_10_436_3201_0, i_10_436_3202_0, i_10_436_3267_0, i_10_436_3268_0,
    i_10_436_3297_0, i_10_436_3360_0, i_10_436_3387_0, i_10_436_3389_0,
    i_10_436_3402_0, i_10_436_3403_0, i_10_436_3405_0, i_10_436_3408_0,
    i_10_436_3525_0, i_10_436_3550_0, i_10_436_3551_0, i_10_436_3553_0,
    i_10_436_3582_0, i_10_436_3604_0, i_10_436_3605_0, i_10_436_3611_0,
    i_10_436_3702_0, i_10_436_3854_0, i_10_436_3855_0, i_10_436_3859_0,
    i_10_436_3901_0, i_10_436_3978_0, i_10_436_3982_0, i_10_436_4185_0,
    i_10_436_4213_0, i_10_436_4216_0, i_10_436_4233_0, i_10_436_4278_0,
    i_10_436_4290_0, i_10_436_4375_0, i_10_436_4376_0, i_10_436_4500_0;
  output o_10_436_0_0;
  assign o_10_436_0_0 = 0;
endmodule



// Benchmark "kernel_10_437" written by ABC on Sun Jul 19 10:28:39 2020

module kernel_10_437 ( 
    i_10_437_30_0, i_10_437_173_0, i_10_437_254_0, i_10_437_390_0,
    i_10_437_407_0, i_10_437_462_0, i_10_437_465_0, i_10_437_631_0,
    i_10_437_633_0, i_10_437_686_0, i_10_437_732_0, i_10_437_733_0,
    i_10_437_736_0, i_10_437_751_0, i_10_437_792_0, i_10_437_793_0,
    i_10_437_795_0, i_10_437_1037_0, i_10_437_1039_0, i_10_437_1087_0,
    i_10_437_1234_0, i_10_437_1305_0, i_10_437_1306_0, i_10_437_1308_0,
    i_10_437_1310_0, i_10_437_1363_0, i_10_437_1397_0, i_10_437_1552_0,
    i_10_437_1714_0, i_10_437_1822_0, i_10_437_1823_0, i_10_437_1824_0,
    i_10_437_1881_0, i_10_437_1882_0, i_10_437_1883_0, i_10_437_1911_0,
    i_10_437_1925_0, i_10_437_2001_0, i_10_437_2026_0, i_10_437_2080_0,
    i_10_437_2093_0, i_10_437_2241_0, i_10_437_2242_0, i_10_437_2243_0,
    i_10_437_2263_0, i_10_437_2309_0, i_10_437_2349_0, i_10_437_2385_0,
    i_10_437_2451_0, i_10_437_2541_0, i_10_437_2612_0, i_10_437_2615_0,
    i_10_437_2628_0, i_10_437_2631_0, i_10_437_2712_0, i_10_437_2742_0,
    i_10_437_2979_0, i_10_437_3072_0, i_10_437_3073_0, i_10_437_3089_0,
    i_10_437_3096_0, i_10_437_3117_0, i_10_437_3121_0, i_10_437_3203_0,
    i_10_437_3232_0, i_10_437_3233_0, i_10_437_3271_0, i_10_437_3387_0,
    i_10_437_3465_0, i_10_437_3519_0, i_10_437_3537_0, i_10_437_3538_0,
    i_10_437_3539_0, i_10_437_3578_0, i_10_437_3609_0, i_10_437_3610_0,
    i_10_437_3645_0, i_10_437_3651_0, i_10_437_3686_0, i_10_437_3798_0,
    i_10_437_3823_0, i_10_437_3844_0, i_10_437_3847_0, i_10_437_3853_0,
    i_10_437_3859_0, i_10_437_3893_0, i_10_437_3942_0, i_10_437_3946_0,
    i_10_437_3997_0, i_10_437_4051_0, i_10_437_4113_0, i_10_437_4116_0,
    i_10_437_4122_0, i_10_437_4125_0, i_10_437_4262_0, i_10_437_4275_0,
    i_10_437_4285_0, i_10_437_4286_0, i_10_437_4459_0, i_10_437_4567_0,
    o_10_437_0_0  );
  input  i_10_437_30_0, i_10_437_173_0, i_10_437_254_0, i_10_437_390_0,
    i_10_437_407_0, i_10_437_462_0, i_10_437_465_0, i_10_437_631_0,
    i_10_437_633_0, i_10_437_686_0, i_10_437_732_0, i_10_437_733_0,
    i_10_437_736_0, i_10_437_751_0, i_10_437_792_0, i_10_437_793_0,
    i_10_437_795_0, i_10_437_1037_0, i_10_437_1039_0, i_10_437_1087_0,
    i_10_437_1234_0, i_10_437_1305_0, i_10_437_1306_0, i_10_437_1308_0,
    i_10_437_1310_0, i_10_437_1363_0, i_10_437_1397_0, i_10_437_1552_0,
    i_10_437_1714_0, i_10_437_1822_0, i_10_437_1823_0, i_10_437_1824_0,
    i_10_437_1881_0, i_10_437_1882_0, i_10_437_1883_0, i_10_437_1911_0,
    i_10_437_1925_0, i_10_437_2001_0, i_10_437_2026_0, i_10_437_2080_0,
    i_10_437_2093_0, i_10_437_2241_0, i_10_437_2242_0, i_10_437_2243_0,
    i_10_437_2263_0, i_10_437_2309_0, i_10_437_2349_0, i_10_437_2385_0,
    i_10_437_2451_0, i_10_437_2541_0, i_10_437_2612_0, i_10_437_2615_0,
    i_10_437_2628_0, i_10_437_2631_0, i_10_437_2712_0, i_10_437_2742_0,
    i_10_437_2979_0, i_10_437_3072_0, i_10_437_3073_0, i_10_437_3089_0,
    i_10_437_3096_0, i_10_437_3117_0, i_10_437_3121_0, i_10_437_3203_0,
    i_10_437_3232_0, i_10_437_3233_0, i_10_437_3271_0, i_10_437_3387_0,
    i_10_437_3465_0, i_10_437_3519_0, i_10_437_3537_0, i_10_437_3538_0,
    i_10_437_3539_0, i_10_437_3578_0, i_10_437_3609_0, i_10_437_3610_0,
    i_10_437_3645_0, i_10_437_3651_0, i_10_437_3686_0, i_10_437_3798_0,
    i_10_437_3823_0, i_10_437_3844_0, i_10_437_3847_0, i_10_437_3853_0,
    i_10_437_3859_0, i_10_437_3893_0, i_10_437_3942_0, i_10_437_3946_0,
    i_10_437_3997_0, i_10_437_4051_0, i_10_437_4113_0, i_10_437_4116_0,
    i_10_437_4122_0, i_10_437_4125_0, i_10_437_4262_0, i_10_437_4275_0,
    i_10_437_4285_0, i_10_437_4286_0, i_10_437_4459_0, i_10_437_4567_0;
  output o_10_437_0_0;
  assign o_10_437_0_0 = 0;
endmodule



// Benchmark "kernel_10_438" written by ABC on Sun Jul 19 10:28:40 2020

module kernel_10_438 ( 
    i_10_438_32_0, i_10_438_171_0, i_10_438_172_0, i_10_438_175_0,
    i_10_438_176_0, i_10_438_179_0, i_10_438_282_0, i_10_438_283_0,
    i_10_438_284_0, i_10_438_411_0, i_10_438_432_0, i_10_438_436_0,
    i_10_438_439_0, i_10_438_466_0, i_10_438_508_0, i_10_438_795_0,
    i_10_438_797_0, i_10_438_800_0, i_10_438_1166_0, i_10_438_1235_0,
    i_10_438_1237_0, i_10_438_1238_0, i_10_438_1240_0, i_10_438_1241_0,
    i_10_438_1296_0, i_10_438_1305_0, i_10_438_1306_0, i_10_438_1346_0,
    i_10_438_1445_0, i_10_438_1622_0, i_10_438_1685_0, i_10_438_1686_0,
    i_10_438_1687_0, i_10_438_1819_0, i_10_438_1821_0, i_10_438_1822_0,
    i_10_438_1823_0, i_10_438_1911_0, i_10_438_1913_0, i_10_438_1945_0,
    i_10_438_2033_0, i_10_438_2353_0, i_10_438_2457_0, i_10_438_2461_0,
    i_10_438_2466_0, i_10_438_2468_0, i_10_438_2567_0, i_10_438_2628_0,
    i_10_438_2629_0, i_10_438_2631_0, i_10_438_2632_0, i_10_438_2633_0,
    i_10_438_2635_0, i_10_438_2658_0, i_10_438_2659_0, i_10_438_2661_0,
    i_10_438_2662_0, i_10_438_2663_0, i_10_438_2710_0, i_10_438_2711_0,
    i_10_438_2714_0, i_10_438_2717_0, i_10_438_2723_0, i_10_438_2728_0,
    i_10_438_2830_0, i_10_438_2831_0, i_10_438_3036_0, i_10_438_3071_0,
    i_10_438_3197_0, i_10_438_3199_0, i_10_438_3200_0, i_10_438_3277_0,
    i_10_438_3278_0, i_10_438_3281_0, i_10_438_3385_0, i_10_438_3386_0,
    i_10_438_3389_0, i_10_438_3467_0, i_10_438_3541_0, i_10_438_3584_0,
    i_10_438_3587_0, i_10_438_3613_0, i_10_438_3617_0, i_10_438_3645_0,
    i_10_438_3647_0, i_10_438_3782_0, i_10_438_3784_0, i_10_438_3785_0,
    i_10_438_3837_0, i_10_438_3839_0, i_10_438_3847_0, i_10_438_3854_0,
    i_10_438_3856_0, i_10_438_3857_0, i_10_438_3914_0, i_10_438_4115_0,
    i_10_438_4123_0, i_10_438_4268_0, i_10_438_4285_0, i_10_438_4286_0,
    o_10_438_0_0  );
  input  i_10_438_32_0, i_10_438_171_0, i_10_438_172_0, i_10_438_175_0,
    i_10_438_176_0, i_10_438_179_0, i_10_438_282_0, i_10_438_283_0,
    i_10_438_284_0, i_10_438_411_0, i_10_438_432_0, i_10_438_436_0,
    i_10_438_439_0, i_10_438_466_0, i_10_438_508_0, i_10_438_795_0,
    i_10_438_797_0, i_10_438_800_0, i_10_438_1166_0, i_10_438_1235_0,
    i_10_438_1237_0, i_10_438_1238_0, i_10_438_1240_0, i_10_438_1241_0,
    i_10_438_1296_0, i_10_438_1305_0, i_10_438_1306_0, i_10_438_1346_0,
    i_10_438_1445_0, i_10_438_1622_0, i_10_438_1685_0, i_10_438_1686_0,
    i_10_438_1687_0, i_10_438_1819_0, i_10_438_1821_0, i_10_438_1822_0,
    i_10_438_1823_0, i_10_438_1911_0, i_10_438_1913_0, i_10_438_1945_0,
    i_10_438_2033_0, i_10_438_2353_0, i_10_438_2457_0, i_10_438_2461_0,
    i_10_438_2466_0, i_10_438_2468_0, i_10_438_2567_0, i_10_438_2628_0,
    i_10_438_2629_0, i_10_438_2631_0, i_10_438_2632_0, i_10_438_2633_0,
    i_10_438_2635_0, i_10_438_2658_0, i_10_438_2659_0, i_10_438_2661_0,
    i_10_438_2662_0, i_10_438_2663_0, i_10_438_2710_0, i_10_438_2711_0,
    i_10_438_2714_0, i_10_438_2717_0, i_10_438_2723_0, i_10_438_2728_0,
    i_10_438_2830_0, i_10_438_2831_0, i_10_438_3036_0, i_10_438_3071_0,
    i_10_438_3197_0, i_10_438_3199_0, i_10_438_3200_0, i_10_438_3277_0,
    i_10_438_3278_0, i_10_438_3281_0, i_10_438_3385_0, i_10_438_3386_0,
    i_10_438_3389_0, i_10_438_3467_0, i_10_438_3541_0, i_10_438_3584_0,
    i_10_438_3587_0, i_10_438_3613_0, i_10_438_3617_0, i_10_438_3645_0,
    i_10_438_3647_0, i_10_438_3782_0, i_10_438_3784_0, i_10_438_3785_0,
    i_10_438_3837_0, i_10_438_3839_0, i_10_438_3847_0, i_10_438_3854_0,
    i_10_438_3856_0, i_10_438_3857_0, i_10_438_3914_0, i_10_438_4115_0,
    i_10_438_4123_0, i_10_438_4268_0, i_10_438_4285_0, i_10_438_4286_0;
  output o_10_438_0_0;
  assign o_10_438_0_0 = ~((~i_10_438_172_0 & ((~i_10_438_283_0 & i_10_438_1821_0 & ~i_10_438_2714_0) | (~i_10_438_171_0 & ~i_10_438_1166_0 & ~i_10_438_1346_0 & ~i_10_438_1911_0 & ~i_10_438_2662_0 & ~i_10_438_2717_0 & ~i_10_438_3071_0 & i_10_438_3386_0 & ~i_10_438_3541_0 & ~i_10_438_4115_0 & ~i_10_438_4268_0))) | (~i_10_438_3584_0 & ((~i_10_438_171_0 & ((~i_10_438_1823_0 & ~i_10_438_1913_0 & ~i_10_438_2723_0 & ~i_10_438_3837_0) | (~i_10_438_176_0 & ~i_10_438_466_0 & i_10_438_1687_0 & ~i_10_438_2466_0 & ~i_10_438_2567_0 & ~i_10_438_3857_0))) | (~i_10_438_3467_0 & ((~i_10_438_1240_0 & ~i_10_438_1445_0 & ~i_10_438_2033_0 & ~i_10_438_2466_0 & ~i_10_438_2567_0 & i_10_438_3386_0 & ~i_10_438_3587_0) | (~i_10_438_1166_0 & i_10_438_1685_0 & ~i_10_438_1821_0 & ~i_10_438_2831_0 & ~i_10_438_3613_0 & ~i_10_438_3782_0 & ~i_10_438_3784_0))))) | (~i_10_438_179_0 & ((~i_10_438_284_0 & ~i_10_438_411_0 & ~i_10_438_2468_0 & ~i_10_438_2710_0) | (i_10_438_1305_0 & ~i_10_438_2659_0 & ~i_10_438_3071_0 & ~i_10_438_3541_0))) | (~i_10_438_282_0 & ((~i_10_438_1445_0 & ~i_10_438_1685_0 & i_10_438_1823_0 & ~i_10_438_2633_0 & ~i_10_438_2831_0 & ~i_10_438_3281_0 & ~i_10_438_3386_0) | (~i_10_438_1237_0 & ~i_10_438_1238_0 & ~i_10_438_1240_0 & ~i_10_438_1819_0 & i_10_438_2723_0 & ~i_10_438_4268_0 & ~i_10_438_4285_0))) | (~i_10_438_284_0 & ((~i_10_438_1237_0 & i_10_438_1240_0 & i_10_438_3839_0) | (~i_10_438_1240_0 & i_10_438_2632_0 & ~i_10_438_2714_0 & i_10_438_3914_0))) | (~i_10_438_1235_0 & ((~i_10_438_176_0 & ~i_10_438_1238_0 & ~i_10_438_2723_0) | (~i_10_438_411_0 & ~i_10_438_1346_0 & ~i_10_438_2714_0 & ~i_10_438_3386_0 & ~i_10_438_3784_0 & ~i_10_438_3839_0 & ~i_10_438_3914_0))) | (~i_10_438_176_0 & ((~i_10_438_1237_0 & ~i_10_438_1346_0 & ~i_10_438_1685_0 & i_10_438_2461_0 & ~i_10_438_2661_0 & ~i_10_438_3613_0) | (~i_10_438_283_0 & ~i_10_438_800_0 & ~i_10_438_1445_0 & i_10_438_1819_0 & ~i_10_438_4123_0))) | (~i_10_438_2033_0 & ~i_10_438_2711_0 & ((~i_10_438_1346_0 & ((~i_10_438_797_0 & ~i_10_438_1686_0 & ~i_10_438_1913_0 & ~i_10_438_2461_0 & ~i_10_438_2567_0 & ~i_10_438_2661_0) | (~i_10_438_1445_0 & ~i_10_438_1685_0 & ~i_10_438_2714_0 & ~i_10_438_2830_0 & ~i_10_438_3200_0 & ~i_10_438_3784_0))) | (i_10_438_176_0 & ~i_10_438_1445_0 & ~i_10_438_2466_0 & ~i_10_438_2723_0 & ~i_10_438_3857_0 & ~i_10_438_4286_0))) | (~i_10_438_4285_0 & ((~i_10_438_1240_0 & i_10_438_2631_0) | (~i_10_438_1241_0 & i_10_438_1819_0 & ~i_10_438_3071_0 & ~i_10_438_3467_0))) | (i_10_438_2461_0 & i_10_438_2632_0 & ~i_10_438_2633_0) | (~i_10_438_795_0 & ~i_10_438_1445_0 & ~i_10_438_2468_0 & i_10_438_2658_0 & ~i_10_438_3587_0 & ~i_10_438_3617_0) | (~i_10_438_1238_0 & i_10_438_2633_0 & ~i_10_438_2662_0 & ~i_10_438_4286_0));
endmodule



// Benchmark "kernel_10_439" written by ABC on Sun Jul 19 10:28:41 2020

module kernel_10_439 ( 
    i_10_439_118_0, i_10_439_175_0, i_10_439_217_0, i_10_439_283_0,
    i_10_439_284_0, i_10_439_288_0, i_10_439_441_0, i_10_439_445_0,
    i_10_439_460_0, i_10_439_463_0, i_10_439_506_0, i_10_439_509_0,
    i_10_439_514_0, i_10_439_793_0, i_10_439_1026_0, i_10_439_1045_0,
    i_10_439_1082_0, i_10_439_1120_0, i_10_439_1234_0, i_10_439_1235_0,
    i_10_439_1237_0, i_10_439_1239_0, i_10_439_1244_0, i_10_439_1359_0,
    i_10_439_1361_0, i_10_439_1364_0, i_10_439_1445_0, i_10_439_1542_0,
    i_10_439_1577_0, i_10_439_1621_0, i_10_439_1648_0, i_10_439_1649_0,
    i_10_439_1650_0, i_10_439_1651_0, i_10_439_1652_0, i_10_439_1653_0,
    i_10_439_1691_0, i_10_439_1767_0, i_10_439_1768_0, i_10_439_1769_0,
    i_10_439_1800_0, i_10_439_1824_0, i_10_439_1910_0, i_10_439_2017_0,
    i_10_439_2232_0, i_10_439_2353_0, i_10_439_2357_0, i_10_439_2448_0,
    i_10_439_2449_0, i_10_439_2450_0, i_10_439_2459_0, i_10_439_2465_0,
    i_10_439_2473_0, i_10_439_2516_0, i_10_439_2565_0, i_10_439_2566_0,
    i_10_439_2630_0, i_10_439_2639_0, i_10_439_2727_0, i_10_439_2729_0,
    i_10_439_2782_0, i_10_439_2831_0, i_10_439_3042_0, i_10_439_3047_0,
    i_10_439_3088_0, i_10_439_3331_0, i_10_439_3388_0, i_10_439_3390_0,
    i_10_439_3406_0, i_10_439_3467_0, i_10_439_3522_0, i_10_439_3555_0,
    i_10_439_3556_0, i_10_439_3584_0, i_10_439_3586_0, i_10_439_3587_0,
    i_10_439_3618_0, i_10_439_3774_0, i_10_439_3840_0, i_10_439_3845_0,
    i_10_439_3847_0, i_10_439_3848_0, i_10_439_3852_0, i_10_439_3853_0,
    i_10_439_3980_0, i_10_439_4024_0, i_10_439_4025_0, i_10_439_4027_0,
    i_10_439_4028_0, i_10_439_4114_0, i_10_439_4115_0, i_10_439_4122_0,
    i_10_439_4123_0, i_10_439_4124_0, i_10_439_4126_0, i_10_439_4150_0,
    i_10_439_4175_0, i_10_439_4285_0, i_10_439_4287_0, i_10_439_4563_0,
    o_10_439_0_0  );
  input  i_10_439_118_0, i_10_439_175_0, i_10_439_217_0, i_10_439_283_0,
    i_10_439_284_0, i_10_439_288_0, i_10_439_441_0, i_10_439_445_0,
    i_10_439_460_0, i_10_439_463_0, i_10_439_506_0, i_10_439_509_0,
    i_10_439_514_0, i_10_439_793_0, i_10_439_1026_0, i_10_439_1045_0,
    i_10_439_1082_0, i_10_439_1120_0, i_10_439_1234_0, i_10_439_1235_0,
    i_10_439_1237_0, i_10_439_1239_0, i_10_439_1244_0, i_10_439_1359_0,
    i_10_439_1361_0, i_10_439_1364_0, i_10_439_1445_0, i_10_439_1542_0,
    i_10_439_1577_0, i_10_439_1621_0, i_10_439_1648_0, i_10_439_1649_0,
    i_10_439_1650_0, i_10_439_1651_0, i_10_439_1652_0, i_10_439_1653_0,
    i_10_439_1691_0, i_10_439_1767_0, i_10_439_1768_0, i_10_439_1769_0,
    i_10_439_1800_0, i_10_439_1824_0, i_10_439_1910_0, i_10_439_2017_0,
    i_10_439_2232_0, i_10_439_2353_0, i_10_439_2357_0, i_10_439_2448_0,
    i_10_439_2449_0, i_10_439_2450_0, i_10_439_2459_0, i_10_439_2465_0,
    i_10_439_2473_0, i_10_439_2516_0, i_10_439_2565_0, i_10_439_2566_0,
    i_10_439_2630_0, i_10_439_2639_0, i_10_439_2727_0, i_10_439_2729_0,
    i_10_439_2782_0, i_10_439_2831_0, i_10_439_3042_0, i_10_439_3047_0,
    i_10_439_3088_0, i_10_439_3331_0, i_10_439_3388_0, i_10_439_3390_0,
    i_10_439_3406_0, i_10_439_3467_0, i_10_439_3522_0, i_10_439_3555_0,
    i_10_439_3556_0, i_10_439_3584_0, i_10_439_3586_0, i_10_439_3587_0,
    i_10_439_3618_0, i_10_439_3774_0, i_10_439_3840_0, i_10_439_3845_0,
    i_10_439_3847_0, i_10_439_3848_0, i_10_439_3852_0, i_10_439_3853_0,
    i_10_439_3980_0, i_10_439_4024_0, i_10_439_4025_0, i_10_439_4027_0,
    i_10_439_4028_0, i_10_439_4114_0, i_10_439_4115_0, i_10_439_4122_0,
    i_10_439_4123_0, i_10_439_4124_0, i_10_439_4126_0, i_10_439_4150_0,
    i_10_439_4175_0, i_10_439_4285_0, i_10_439_4287_0, i_10_439_4563_0;
  output o_10_439_0_0;
  assign o_10_439_0_0 = 0;
endmodule



// Benchmark "kernel_10_440" written by ABC on Sun Jul 19 10:28:42 2020

module kernel_10_440 ( 
    i_10_440_48_0, i_10_440_118_0, i_10_440_119_0, i_10_440_121_0,
    i_10_440_153_0, i_10_440_171_0, i_10_440_172_0, i_10_440_185_0,
    i_10_440_390_0, i_10_440_391_0, i_10_440_433_0, i_10_440_446_0,
    i_10_440_447_0, i_10_440_461_0, i_10_440_463_0, i_10_440_520_0,
    i_10_440_559_0, i_10_440_560_0, i_10_440_694_0, i_10_440_733_0,
    i_10_440_793_0, i_10_440_794_0, i_10_440_797_0, i_10_440_1085_0,
    i_10_440_1235_0, i_10_440_1241_0, i_10_440_1242_0, i_10_440_1361_0,
    i_10_440_1381_0, i_10_440_1433_0, i_10_440_1442_0, i_10_440_1444_0,
    i_10_440_1452_0, i_10_440_1454_0, i_10_440_1532_0, i_10_440_1579_0,
    i_10_440_1613_0, i_10_440_1826_0, i_10_440_1946_0, i_10_440_1949_0,
    i_10_440_2000_0, i_10_440_2090_0, i_10_440_2308_0, i_10_440_2309_0,
    i_10_440_2349_0, i_10_440_2351_0, i_10_440_2352_0, i_10_440_2405_0,
    i_10_440_2407_0, i_10_440_2410_0, i_10_440_2431_0, i_10_440_2454_0,
    i_10_440_2455_0, i_10_440_2456_0, i_10_440_2461_0, i_10_440_2471_0,
    i_10_440_2614_0, i_10_440_2615_0, i_10_440_2629_0, i_10_440_2630_0,
    i_10_440_2642_0, i_10_440_2656_0, i_10_440_2660_0, i_10_440_2674_0,
    i_10_440_2677_0, i_10_440_2678_0, i_10_440_2713_0, i_10_440_2723_0,
    i_10_440_2728_0, i_10_440_2729_0, i_10_440_2817_0, i_10_440_2818_0,
    i_10_440_2827_0, i_10_440_2829_0, i_10_440_2881_0, i_10_440_2884_0,
    i_10_440_2968_0, i_10_440_2980_0, i_10_440_3037_0, i_10_440_3313_0,
    i_10_440_3316_0, i_10_440_3384_0, i_10_440_3387_0, i_10_440_3391_0,
    i_10_440_3470_0, i_10_440_3522_0, i_10_440_3539_0, i_10_440_3586_0,
    i_10_440_3587_0, i_10_440_3717_0, i_10_440_3857_0, i_10_440_3947_0,
    i_10_440_3979_0, i_10_440_3981_0, i_10_440_3989_0, i_10_440_4120_0,
    i_10_440_4144_0, i_10_440_4268_0, i_10_440_4275_0, i_10_440_4276_0,
    o_10_440_0_0  );
  input  i_10_440_48_0, i_10_440_118_0, i_10_440_119_0, i_10_440_121_0,
    i_10_440_153_0, i_10_440_171_0, i_10_440_172_0, i_10_440_185_0,
    i_10_440_390_0, i_10_440_391_0, i_10_440_433_0, i_10_440_446_0,
    i_10_440_447_0, i_10_440_461_0, i_10_440_463_0, i_10_440_520_0,
    i_10_440_559_0, i_10_440_560_0, i_10_440_694_0, i_10_440_733_0,
    i_10_440_793_0, i_10_440_794_0, i_10_440_797_0, i_10_440_1085_0,
    i_10_440_1235_0, i_10_440_1241_0, i_10_440_1242_0, i_10_440_1361_0,
    i_10_440_1381_0, i_10_440_1433_0, i_10_440_1442_0, i_10_440_1444_0,
    i_10_440_1452_0, i_10_440_1454_0, i_10_440_1532_0, i_10_440_1579_0,
    i_10_440_1613_0, i_10_440_1826_0, i_10_440_1946_0, i_10_440_1949_0,
    i_10_440_2000_0, i_10_440_2090_0, i_10_440_2308_0, i_10_440_2309_0,
    i_10_440_2349_0, i_10_440_2351_0, i_10_440_2352_0, i_10_440_2405_0,
    i_10_440_2407_0, i_10_440_2410_0, i_10_440_2431_0, i_10_440_2454_0,
    i_10_440_2455_0, i_10_440_2456_0, i_10_440_2461_0, i_10_440_2471_0,
    i_10_440_2614_0, i_10_440_2615_0, i_10_440_2629_0, i_10_440_2630_0,
    i_10_440_2642_0, i_10_440_2656_0, i_10_440_2660_0, i_10_440_2674_0,
    i_10_440_2677_0, i_10_440_2678_0, i_10_440_2713_0, i_10_440_2723_0,
    i_10_440_2728_0, i_10_440_2729_0, i_10_440_2817_0, i_10_440_2818_0,
    i_10_440_2827_0, i_10_440_2829_0, i_10_440_2881_0, i_10_440_2884_0,
    i_10_440_2968_0, i_10_440_2980_0, i_10_440_3037_0, i_10_440_3313_0,
    i_10_440_3316_0, i_10_440_3384_0, i_10_440_3387_0, i_10_440_3391_0,
    i_10_440_3470_0, i_10_440_3522_0, i_10_440_3539_0, i_10_440_3586_0,
    i_10_440_3587_0, i_10_440_3717_0, i_10_440_3857_0, i_10_440_3947_0,
    i_10_440_3979_0, i_10_440_3981_0, i_10_440_3989_0, i_10_440_4120_0,
    i_10_440_4144_0, i_10_440_4268_0, i_10_440_4275_0, i_10_440_4276_0;
  output o_10_440_0_0;
  assign o_10_440_0_0 = 0;
endmodule



// Benchmark "kernel_10_441" written by ABC on Sun Jul 19 10:28:43 2020

module kernel_10_441 ( 
    i_10_441_67_0, i_10_441_223_0, i_10_441_445_0, i_10_441_464_0,
    i_10_441_466_0, i_10_441_561_0, i_10_441_593_0, i_10_441_712_0,
    i_10_441_736_0, i_10_441_737_0, i_10_441_934_0, i_10_441_957_0,
    i_10_441_999_0, i_10_441_1032_0, i_10_441_1033_0, i_10_441_1034_0,
    i_10_441_1039_0, i_10_441_1088_0, i_10_441_1128_0, i_10_441_1138_0,
    i_10_441_1139_0, i_10_441_1164_0, i_10_441_1165_0, i_10_441_1166_0,
    i_10_441_1233_0, i_10_441_1243_0, i_10_441_1247_0, i_10_441_1248_0,
    i_10_441_1250_0, i_10_441_1307_0, i_10_441_1309_0, i_10_441_1313_0,
    i_10_441_1365_0, i_10_441_1652_0, i_10_441_1653_0, i_10_441_1654_0,
    i_10_441_1823_0, i_10_441_1910_0, i_10_441_1915_0, i_10_441_1917_0,
    i_10_441_1920_0, i_10_441_2154_0, i_10_441_2310_0, i_10_441_2311_0,
    i_10_441_2352_0, i_10_441_2353_0, i_10_441_2454_0, i_10_441_2455_0,
    i_10_441_2512_0, i_10_441_2517_0, i_10_441_2520_0, i_10_441_2521_0,
    i_10_441_2619_0, i_10_441_2631_0, i_10_441_2632_0, i_10_441_2655_0,
    i_10_441_2659_0, i_10_441_2673_0, i_10_441_2722_0, i_10_441_2726_0,
    i_10_441_2831_0, i_10_441_2834_0, i_10_441_2882_0, i_10_441_2884_0,
    i_10_441_2953_0, i_10_441_3071_0, i_10_441_3075_0, i_10_441_3267_0,
    i_10_441_3269_0, i_10_441_3270_0, i_10_441_3275_0, i_10_441_3282_0,
    i_10_441_3390_0, i_10_441_3470_0, i_10_441_3547_0, i_10_441_3548_0,
    i_10_441_3583_0, i_10_441_3585_0, i_10_441_3586_0, i_10_441_3609_0,
    i_10_441_3648_0, i_10_441_3781_0, i_10_441_3782_0, i_10_441_3783_0,
    i_10_441_3784_0, i_10_441_3787_0, i_10_441_3788_0, i_10_441_3835_0,
    i_10_441_3838_0, i_10_441_3839_0, i_10_441_3852_0, i_10_441_3909_0,
    i_10_441_3943_0, i_10_441_3986_0, i_10_441_3999_0, i_10_441_4117_0,
    i_10_441_4118_0, i_10_441_4119_0, i_10_441_4125_0, i_10_441_4303_0,
    o_10_441_0_0  );
  input  i_10_441_67_0, i_10_441_223_0, i_10_441_445_0, i_10_441_464_0,
    i_10_441_466_0, i_10_441_561_0, i_10_441_593_0, i_10_441_712_0,
    i_10_441_736_0, i_10_441_737_0, i_10_441_934_0, i_10_441_957_0,
    i_10_441_999_0, i_10_441_1032_0, i_10_441_1033_0, i_10_441_1034_0,
    i_10_441_1039_0, i_10_441_1088_0, i_10_441_1128_0, i_10_441_1138_0,
    i_10_441_1139_0, i_10_441_1164_0, i_10_441_1165_0, i_10_441_1166_0,
    i_10_441_1233_0, i_10_441_1243_0, i_10_441_1247_0, i_10_441_1248_0,
    i_10_441_1250_0, i_10_441_1307_0, i_10_441_1309_0, i_10_441_1313_0,
    i_10_441_1365_0, i_10_441_1652_0, i_10_441_1653_0, i_10_441_1654_0,
    i_10_441_1823_0, i_10_441_1910_0, i_10_441_1915_0, i_10_441_1917_0,
    i_10_441_1920_0, i_10_441_2154_0, i_10_441_2310_0, i_10_441_2311_0,
    i_10_441_2352_0, i_10_441_2353_0, i_10_441_2454_0, i_10_441_2455_0,
    i_10_441_2512_0, i_10_441_2517_0, i_10_441_2520_0, i_10_441_2521_0,
    i_10_441_2619_0, i_10_441_2631_0, i_10_441_2632_0, i_10_441_2655_0,
    i_10_441_2659_0, i_10_441_2673_0, i_10_441_2722_0, i_10_441_2726_0,
    i_10_441_2831_0, i_10_441_2834_0, i_10_441_2882_0, i_10_441_2884_0,
    i_10_441_2953_0, i_10_441_3071_0, i_10_441_3075_0, i_10_441_3267_0,
    i_10_441_3269_0, i_10_441_3270_0, i_10_441_3275_0, i_10_441_3282_0,
    i_10_441_3390_0, i_10_441_3470_0, i_10_441_3547_0, i_10_441_3548_0,
    i_10_441_3583_0, i_10_441_3585_0, i_10_441_3586_0, i_10_441_3609_0,
    i_10_441_3648_0, i_10_441_3781_0, i_10_441_3782_0, i_10_441_3783_0,
    i_10_441_3784_0, i_10_441_3787_0, i_10_441_3788_0, i_10_441_3835_0,
    i_10_441_3838_0, i_10_441_3839_0, i_10_441_3852_0, i_10_441_3909_0,
    i_10_441_3943_0, i_10_441_3986_0, i_10_441_3999_0, i_10_441_4117_0,
    i_10_441_4118_0, i_10_441_4119_0, i_10_441_4125_0, i_10_441_4303_0;
  output o_10_441_0_0;
  assign o_10_441_0_0 = 0;
endmodule



// Benchmark "kernel_10_442" written by ABC on Sun Jul 19 10:28:44 2020

module kernel_10_442 ( 
    i_10_442_98_0, i_10_442_177_0, i_10_442_250_0, i_10_442_258_0,
    i_10_442_267_0, i_10_442_274_0, i_10_442_280_0, i_10_442_292_0,
    i_10_442_295_0, i_10_442_318_0, i_10_442_321_0, i_10_442_322_0,
    i_10_442_406_0, i_10_442_408_0, i_10_442_409_0, i_10_442_412_0,
    i_10_442_413_0, i_10_442_460_0, i_10_442_463_0, i_10_442_464_0,
    i_10_442_628_0, i_10_442_712_0, i_10_442_714_0, i_10_442_717_0,
    i_10_442_831_0, i_10_442_870_0, i_10_442_871_0, i_10_442_898_0,
    i_10_442_930_0, i_10_442_968_0, i_10_442_989_0, i_10_442_1033_0,
    i_10_442_1233_0, i_10_442_1239_0, i_10_442_1347_0, i_10_442_1363_0,
    i_10_442_1438_0, i_10_442_1543_0, i_10_442_1545_0, i_10_442_1546_0,
    i_10_442_1555_0, i_10_442_1581_0, i_10_442_1626_0, i_10_442_1633_0,
    i_10_442_1635_0, i_10_442_1686_0, i_10_442_1689_0, i_10_442_1806_0,
    i_10_442_1824_0, i_10_442_1885_0, i_10_442_1986_0, i_10_442_2031_0,
    i_10_442_2255_0, i_10_442_2339_0, i_10_442_2356_0, i_10_442_2364_0,
    i_10_442_2383_0, i_10_442_2384_0, i_10_442_2472_0, i_10_442_2514_0,
    i_10_442_2515_0, i_10_442_2572_0, i_10_442_2581_0, i_10_442_2608_0,
    i_10_442_2643_0, i_10_442_2659_0, i_10_442_2678_0, i_10_442_2712_0,
    i_10_442_2713_0, i_10_442_2714_0, i_10_442_2715_0, i_10_442_2716_0,
    i_10_442_2829_0, i_10_442_2884_0, i_10_442_2960_0, i_10_442_3072_0,
    i_10_442_3075_0, i_10_442_3232_0, i_10_442_3281_0, i_10_442_3283_0,
    i_10_442_3315_0, i_10_442_3318_0, i_10_442_3328_0, i_10_442_3337_0,
    i_10_442_3389_0, i_10_442_3405_0, i_10_442_3497_0, i_10_442_3507_0,
    i_10_442_3508_0, i_10_442_3526_0, i_10_442_3543_0, i_10_442_3650_0,
    i_10_442_3685_0, i_10_442_3977_0, i_10_442_4119_0, i_10_442_4120_0,
    i_10_442_4128_0, i_10_442_4210_0, i_10_442_4282_0, i_10_442_4585_0,
    o_10_442_0_0  );
  input  i_10_442_98_0, i_10_442_177_0, i_10_442_250_0, i_10_442_258_0,
    i_10_442_267_0, i_10_442_274_0, i_10_442_280_0, i_10_442_292_0,
    i_10_442_295_0, i_10_442_318_0, i_10_442_321_0, i_10_442_322_0,
    i_10_442_406_0, i_10_442_408_0, i_10_442_409_0, i_10_442_412_0,
    i_10_442_413_0, i_10_442_460_0, i_10_442_463_0, i_10_442_464_0,
    i_10_442_628_0, i_10_442_712_0, i_10_442_714_0, i_10_442_717_0,
    i_10_442_831_0, i_10_442_870_0, i_10_442_871_0, i_10_442_898_0,
    i_10_442_930_0, i_10_442_968_0, i_10_442_989_0, i_10_442_1033_0,
    i_10_442_1233_0, i_10_442_1239_0, i_10_442_1347_0, i_10_442_1363_0,
    i_10_442_1438_0, i_10_442_1543_0, i_10_442_1545_0, i_10_442_1546_0,
    i_10_442_1555_0, i_10_442_1581_0, i_10_442_1626_0, i_10_442_1633_0,
    i_10_442_1635_0, i_10_442_1686_0, i_10_442_1689_0, i_10_442_1806_0,
    i_10_442_1824_0, i_10_442_1885_0, i_10_442_1986_0, i_10_442_2031_0,
    i_10_442_2255_0, i_10_442_2339_0, i_10_442_2356_0, i_10_442_2364_0,
    i_10_442_2383_0, i_10_442_2384_0, i_10_442_2472_0, i_10_442_2514_0,
    i_10_442_2515_0, i_10_442_2572_0, i_10_442_2581_0, i_10_442_2608_0,
    i_10_442_2643_0, i_10_442_2659_0, i_10_442_2678_0, i_10_442_2712_0,
    i_10_442_2713_0, i_10_442_2714_0, i_10_442_2715_0, i_10_442_2716_0,
    i_10_442_2829_0, i_10_442_2884_0, i_10_442_2960_0, i_10_442_3072_0,
    i_10_442_3075_0, i_10_442_3232_0, i_10_442_3281_0, i_10_442_3283_0,
    i_10_442_3315_0, i_10_442_3318_0, i_10_442_3328_0, i_10_442_3337_0,
    i_10_442_3389_0, i_10_442_3405_0, i_10_442_3497_0, i_10_442_3507_0,
    i_10_442_3508_0, i_10_442_3526_0, i_10_442_3543_0, i_10_442_3650_0,
    i_10_442_3685_0, i_10_442_3977_0, i_10_442_4119_0, i_10_442_4120_0,
    i_10_442_4128_0, i_10_442_4210_0, i_10_442_4282_0, i_10_442_4585_0;
  output o_10_442_0_0;
  assign o_10_442_0_0 = 0;
endmodule



// Benchmark "kernel_10_443" written by ABC on Sun Jul 19 10:28:45 2020

module kernel_10_443 ( 
    i_10_443_120_0, i_10_443_174_0, i_10_443_180_0, i_10_443_181_0,
    i_10_443_256_0, i_10_443_275_0, i_10_443_319_0, i_10_443_323_0,
    i_10_443_387_0, i_10_443_388_0, i_10_443_390_0, i_10_443_423_0,
    i_10_443_426_0, i_10_443_462_0, i_10_443_495_0, i_10_443_496_0,
    i_10_443_507_0, i_10_443_508_0, i_10_443_1030_0, i_10_443_1035_0,
    i_10_443_1080_0, i_10_443_1162_0, i_10_443_1215_0, i_10_443_1216_0,
    i_10_443_1233_0, i_10_443_1234_0, i_10_443_1241_0, i_10_443_1359_0,
    i_10_443_1377_0, i_10_443_1578_0, i_10_443_1684_0, i_10_443_1689_0,
    i_10_443_1764_0, i_10_443_1770_0, i_10_443_1822_0, i_10_443_1825_0,
    i_10_443_1908_0, i_10_443_1911_0, i_10_443_1915_0, i_10_443_1989_0,
    i_10_443_1998_0, i_10_443_1999_0, i_10_443_2025_0, i_10_443_2179_0,
    i_10_443_2199_0, i_10_443_2242_0, i_10_443_2305_0, i_10_443_2359_0,
    i_10_443_2361_0, i_10_443_2362_0, i_10_443_2376_0, i_10_443_2379_0,
    i_10_443_2380_0, i_10_443_2457_0, i_10_443_2611_0, i_10_443_2636_0,
    i_10_443_2657_0, i_10_443_2673_0, i_10_443_2711_0, i_10_443_2727_0,
    i_10_443_2817_0, i_10_443_2820_0, i_10_443_2821_0, i_10_443_2919_0,
    i_10_443_2983_0, i_10_443_3152_0, i_10_443_3268_0, i_10_443_3270_0,
    i_10_443_3271_0, i_10_443_3276_0, i_10_443_3277_0, i_10_443_3279_0,
    i_10_443_3282_0, i_10_443_3312_0, i_10_443_3322_0, i_10_443_3387_0,
    i_10_443_3403_0, i_10_443_3466_0, i_10_443_3538_0, i_10_443_3540_0,
    i_10_443_3582_0, i_10_443_3783_0, i_10_443_3784_0, i_10_443_3785_0,
    i_10_443_3787_0, i_10_443_3888_0, i_10_443_3889_0, i_10_443_3978_0,
    i_10_443_3979_0, i_10_443_3980_0, i_10_443_4123_0, i_10_443_4167_0,
    i_10_443_4215_0, i_10_443_4287_0, i_10_443_4288_0, i_10_443_4289_0,
    i_10_443_4290_0, i_10_443_4302_0, i_10_443_4568_0, i_10_443_4569_0,
    o_10_443_0_0  );
  input  i_10_443_120_0, i_10_443_174_0, i_10_443_180_0, i_10_443_181_0,
    i_10_443_256_0, i_10_443_275_0, i_10_443_319_0, i_10_443_323_0,
    i_10_443_387_0, i_10_443_388_0, i_10_443_390_0, i_10_443_423_0,
    i_10_443_426_0, i_10_443_462_0, i_10_443_495_0, i_10_443_496_0,
    i_10_443_507_0, i_10_443_508_0, i_10_443_1030_0, i_10_443_1035_0,
    i_10_443_1080_0, i_10_443_1162_0, i_10_443_1215_0, i_10_443_1216_0,
    i_10_443_1233_0, i_10_443_1234_0, i_10_443_1241_0, i_10_443_1359_0,
    i_10_443_1377_0, i_10_443_1578_0, i_10_443_1684_0, i_10_443_1689_0,
    i_10_443_1764_0, i_10_443_1770_0, i_10_443_1822_0, i_10_443_1825_0,
    i_10_443_1908_0, i_10_443_1911_0, i_10_443_1915_0, i_10_443_1989_0,
    i_10_443_1998_0, i_10_443_1999_0, i_10_443_2025_0, i_10_443_2179_0,
    i_10_443_2199_0, i_10_443_2242_0, i_10_443_2305_0, i_10_443_2359_0,
    i_10_443_2361_0, i_10_443_2362_0, i_10_443_2376_0, i_10_443_2379_0,
    i_10_443_2380_0, i_10_443_2457_0, i_10_443_2611_0, i_10_443_2636_0,
    i_10_443_2657_0, i_10_443_2673_0, i_10_443_2711_0, i_10_443_2727_0,
    i_10_443_2817_0, i_10_443_2820_0, i_10_443_2821_0, i_10_443_2919_0,
    i_10_443_2983_0, i_10_443_3152_0, i_10_443_3268_0, i_10_443_3270_0,
    i_10_443_3271_0, i_10_443_3276_0, i_10_443_3277_0, i_10_443_3279_0,
    i_10_443_3282_0, i_10_443_3312_0, i_10_443_3322_0, i_10_443_3387_0,
    i_10_443_3403_0, i_10_443_3466_0, i_10_443_3538_0, i_10_443_3540_0,
    i_10_443_3582_0, i_10_443_3783_0, i_10_443_3784_0, i_10_443_3785_0,
    i_10_443_3787_0, i_10_443_3888_0, i_10_443_3889_0, i_10_443_3978_0,
    i_10_443_3979_0, i_10_443_3980_0, i_10_443_4123_0, i_10_443_4167_0,
    i_10_443_4215_0, i_10_443_4287_0, i_10_443_4288_0, i_10_443_4289_0,
    i_10_443_4290_0, i_10_443_4302_0, i_10_443_4568_0, i_10_443_4569_0;
  output o_10_443_0_0;
  assign o_10_443_0_0 = ~((~i_10_443_3540_0 & ((~i_10_443_181_0 & ~i_10_443_1915_0 & ((~i_10_443_423_0 & ~i_10_443_1162_0 & ~i_10_443_1822_0 & ~i_10_443_2199_0 & ~i_10_443_2611_0 & ~i_10_443_3276_0) | (~i_10_443_388_0 & ~i_10_443_1359_0 & ~i_10_443_1908_0 & ~i_10_443_2305_0 & ~i_10_443_2376_0 & ~i_10_443_2657_0 & ~i_10_443_2820_0 & ~i_10_443_3279_0 & ~i_10_443_3312_0))) | (~i_10_443_3888_0 & ((~i_10_443_426_0 & ~i_10_443_1162_0 & ~i_10_443_1998_0 & ~i_10_443_2025_0 & ~i_10_443_3980_0 & ~i_10_443_4167_0) | (~i_10_443_323_0 & ~i_10_443_1080_0 & i_10_443_1822_0 & ~i_10_443_2820_0 & ~i_10_443_2919_0 & i_10_443_3582_0 & ~i_10_443_3889_0 & ~i_10_443_4290_0))) | (~i_10_443_1233_0 & ~i_10_443_1911_0 & ~i_10_443_2727_0 & ~i_10_443_2817_0 & ~i_10_443_3312_0))) | (~i_10_443_1035_0 & ((~i_10_443_388_0 & ((~i_10_443_1080_0 & ~i_10_443_1998_0 & ~i_10_443_2727_0 & ~i_10_443_3466_0 & ~i_10_443_3538_0) | (~i_10_443_390_0 & ~i_10_443_423_0 & ~i_10_443_2820_0 & ~i_10_443_2919_0 & ~i_10_443_3979_0))) | (~i_10_443_1684_0 & ((~i_10_443_1998_0 & ~i_10_443_2817_0 & ~i_10_443_2821_0 & ~i_10_443_3889_0 & ~i_10_443_4290_0) | (~i_10_443_2457_0 & ~i_10_443_3466_0 & ~i_10_443_3978_0 & i_10_443_4288_0 & ~i_10_443_4568_0))) | (~i_10_443_1999_0 & ((~i_10_443_387_0 & ~i_10_443_1764_0 & ~i_10_443_1915_0 & ~i_10_443_1998_0 & ~i_10_443_2025_0 & ~i_10_443_2673_0 & ~i_10_443_3279_0 & ~i_10_443_3888_0) | (~i_10_443_2820_0 & ~i_10_443_3978_0 & ~i_10_443_4287_0))) | (~i_10_443_1080_0 & ~i_10_443_1359_0 & ~i_10_443_1689_0 & ~i_10_443_1911_0 & ~i_10_443_2821_0 & i_10_443_2919_0 & ~i_10_443_4167_0))) | (~i_10_443_1359_0 & ((~i_10_443_390_0 & ~i_10_443_3282_0 & ((~i_10_443_387_0 & ~i_10_443_1162_0 & ~i_10_443_1825_0 & ~i_10_443_2711_0 & ~i_10_443_3888_0 & ~i_10_443_3889_0) | (~i_10_443_1998_0 & ~i_10_443_2611_0 & ~i_10_443_2821_0 & ~i_10_443_4167_0 & ~i_10_443_4287_0))) | (~i_10_443_1822_0 & ~i_10_443_1911_0 & ~i_10_443_1998_0 & ~i_10_443_2025_0 & ~i_10_443_3277_0 & ~i_10_443_3980_0 & ~i_10_443_4289_0 & ~i_10_443_4290_0))) | (~i_10_443_387_0 & ((~i_10_443_423_0 & ~i_10_443_1911_0 & ~i_10_443_2380_0 & ~i_10_443_3312_0 & i_10_443_3466_0 & ~i_10_443_3888_0) | (~i_10_443_388_0 & ~i_10_443_2817_0 & ~i_10_443_4287_0 & ~i_10_443_4568_0))) | (~i_10_443_423_0 & ~i_10_443_1234_0 & i_10_443_1915_0 & i_10_443_2636_0 & ~i_10_443_3282_0 & ~i_10_443_3538_0 & ~i_10_443_3978_0 & ~i_10_443_4167_0) | (~i_10_443_4288_0 & i_10_443_4289_0 & i_10_443_4568_0));
endmodule



// Benchmark "kernel_10_444" written by ABC on Sun Jul 19 10:28:46 2020

module kernel_10_444 ( 
    i_10_444_176_0, i_10_444_183_0, i_10_444_223_0, i_10_444_224_0,
    i_10_444_249_0, i_10_444_252_0, i_10_444_282_0, i_10_444_283_0,
    i_10_444_391_0, i_10_444_393_0, i_10_444_408_0, i_10_444_409_0,
    i_10_444_446_0, i_10_444_449_0, i_10_444_515_0, i_10_444_544_0,
    i_10_444_597_0, i_10_444_621_0, i_10_444_689_0, i_10_444_713_0,
    i_10_444_715_0, i_10_444_716_0, i_10_444_753_0, i_10_444_957_0,
    i_10_444_958_0, i_10_444_959_0, i_10_444_962_0, i_10_444_965_0,
    i_10_444_983_0, i_10_444_1000_0, i_10_444_1245_0, i_10_444_1246_0,
    i_10_444_1248_0, i_10_444_1249_0, i_10_444_1260_0, i_10_444_1306_0,
    i_10_444_1307_0, i_10_444_1437_0, i_10_444_1487_0, i_10_444_1492_0,
    i_10_444_1493_0, i_10_444_1532_0, i_10_444_1535_0, i_10_444_1545_0,
    i_10_444_1581_0, i_10_444_1582_0, i_10_444_1683_0, i_10_444_1796_0,
    i_10_444_1823_0, i_10_444_1908_0, i_10_444_1909_0, i_10_444_1912_0,
    i_10_444_2031_0, i_10_444_2185_0, i_10_444_2203_0, i_10_444_2252_0,
    i_10_444_2254_0, i_10_444_2255_0, i_10_444_2327_0, i_10_444_2355_0,
    i_10_444_2362_0, i_10_444_2436_0, i_10_444_2437_0, i_10_444_2451_0,
    i_10_444_2465_0, i_10_444_2506_0, i_10_444_2529_0, i_10_444_2531_0,
    i_10_444_2535_0, i_10_444_2542_0, i_10_444_2704_0, i_10_444_2710_0,
    i_10_444_2731_0, i_10_444_2787_0, i_10_444_2823_0, i_10_444_2985_0,
    i_10_444_3036_0, i_10_444_3038_0, i_10_444_3075_0, i_10_444_3198_0,
    i_10_444_3202_0, i_10_444_3203_0, i_10_444_3238_0, i_10_444_3432_0,
    i_10_444_3588_0, i_10_444_3652_0, i_10_444_3783_0, i_10_444_3786_0,
    i_10_444_3847_0, i_10_444_3855_0, i_10_444_3856_0, i_10_444_3858_0,
    i_10_444_3912_0, i_10_444_3947_0, i_10_444_4002_0, i_10_444_4005_0,
    i_10_444_4011_0, i_10_444_4065_0, i_10_444_4463_0, i_10_444_4567_0,
    o_10_444_0_0  );
  input  i_10_444_176_0, i_10_444_183_0, i_10_444_223_0, i_10_444_224_0,
    i_10_444_249_0, i_10_444_252_0, i_10_444_282_0, i_10_444_283_0,
    i_10_444_391_0, i_10_444_393_0, i_10_444_408_0, i_10_444_409_0,
    i_10_444_446_0, i_10_444_449_0, i_10_444_515_0, i_10_444_544_0,
    i_10_444_597_0, i_10_444_621_0, i_10_444_689_0, i_10_444_713_0,
    i_10_444_715_0, i_10_444_716_0, i_10_444_753_0, i_10_444_957_0,
    i_10_444_958_0, i_10_444_959_0, i_10_444_962_0, i_10_444_965_0,
    i_10_444_983_0, i_10_444_1000_0, i_10_444_1245_0, i_10_444_1246_0,
    i_10_444_1248_0, i_10_444_1249_0, i_10_444_1260_0, i_10_444_1306_0,
    i_10_444_1307_0, i_10_444_1437_0, i_10_444_1487_0, i_10_444_1492_0,
    i_10_444_1493_0, i_10_444_1532_0, i_10_444_1535_0, i_10_444_1545_0,
    i_10_444_1581_0, i_10_444_1582_0, i_10_444_1683_0, i_10_444_1796_0,
    i_10_444_1823_0, i_10_444_1908_0, i_10_444_1909_0, i_10_444_1912_0,
    i_10_444_2031_0, i_10_444_2185_0, i_10_444_2203_0, i_10_444_2252_0,
    i_10_444_2254_0, i_10_444_2255_0, i_10_444_2327_0, i_10_444_2355_0,
    i_10_444_2362_0, i_10_444_2436_0, i_10_444_2437_0, i_10_444_2451_0,
    i_10_444_2465_0, i_10_444_2506_0, i_10_444_2529_0, i_10_444_2531_0,
    i_10_444_2535_0, i_10_444_2542_0, i_10_444_2704_0, i_10_444_2710_0,
    i_10_444_2731_0, i_10_444_2787_0, i_10_444_2823_0, i_10_444_2985_0,
    i_10_444_3036_0, i_10_444_3038_0, i_10_444_3075_0, i_10_444_3198_0,
    i_10_444_3202_0, i_10_444_3203_0, i_10_444_3238_0, i_10_444_3432_0,
    i_10_444_3588_0, i_10_444_3652_0, i_10_444_3783_0, i_10_444_3786_0,
    i_10_444_3847_0, i_10_444_3855_0, i_10_444_3856_0, i_10_444_3858_0,
    i_10_444_3912_0, i_10_444_3947_0, i_10_444_4002_0, i_10_444_4005_0,
    i_10_444_4011_0, i_10_444_4065_0, i_10_444_4463_0, i_10_444_4567_0;
  output o_10_444_0_0;
  assign o_10_444_0_0 = 0;
endmodule



// Benchmark "kernel_10_445" written by ABC on Sun Jul 19 10:28:47 2020

module kernel_10_445 ( 
    i_10_445_220_0, i_10_445_222_0, i_10_445_223_0, i_10_445_250_0,
    i_10_445_279_0, i_10_445_280_0, i_10_445_284_0, i_10_445_318_0,
    i_10_445_322_0, i_10_445_326_0, i_10_445_444_0, i_10_445_445_0,
    i_10_445_448_0, i_10_445_449_0, i_10_445_718_0, i_10_445_751_0,
    i_10_445_752_0, i_10_445_792_0, i_10_445_796_0, i_10_445_898_0,
    i_10_445_963_0, i_10_445_964_0, i_10_445_967_0, i_10_445_997_0,
    i_10_445_1002_0, i_10_445_1003_0, i_10_445_1084_0, i_10_445_1305_0,
    i_10_445_1306_0, i_10_445_1308_0, i_10_445_1437_0, i_10_445_1555_0,
    i_10_445_1580_0, i_10_445_1691_0, i_10_445_1768_0, i_10_445_1819_0,
    i_10_445_1821_0, i_10_445_1822_0, i_10_445_1823_0, i_10_445_1824_0,
    i_10_445_1948_0, i_10_445_2354_0, i_10_445_2362_0, i_10_445_2452_0,
    i_10_445_2453_0, i_10_445_2630_0, i_10_445_2632_0, i_10_445_2633_0,
    i_10_445_2704_0, i_10_445_2706_0, i_10_445_2707_0, i_10_445_2708_0,
    i_10_445_2715_0, i_10_445_2716_0, i_10_445_2717_0, i_10_445_2724_0,
    i_10_445_2725_0, i_10_445_2728_0, i_10_445_2734_0, i_10_445_2782_0,
    i_10_445_2829_0, i_10_445_2830_0, i_10_445_2919_0, i_10_445_2920_0,
    i_10_445_3034_0, i_10_445_3046_0, i_10_445_3076_0, i_10_445_3150_0,
    i_10_445_3154_0, i_10_445_3157_0, i_10_445_3389_0, i_10_445_3390_0,
    i_10_445_3405_0, i_10_445_3406_0, i_10_445_3468_0, i_10_445_3616_0,
    i_10_445_3649_0, i_10_445_3784_0, i_10_445_3787_0, i_10_445_3788_0,
    i_10_445_3815_0, i_10_445_3834_0, i_10_445_3842_0, i_10_445_3848_0,
    i_10_445_3853_0, i_10_445_3856_0, i_10_445_3888_0, i_10_445_3895_0,
    i_10_445_3982_0, i_10_445_3983_0, i_10_445_3985_0, i_10_445_3986_0,
    i_10_445_4116_0, i_10_445_4121_0, i_10_445_4266_0, i_10_445_4273_0,
    i_10_445_4284_0, i_10_445_4287_0, i_10_445_4290_0, i_10_445_4563_0,
    o_10_445_0_0  );
  input  i_10_445_220_0, i_10_445_222_0, i_10_445_223_0, i_10_445_250_0,
    i_10_445_279_0, i_10_445_280_0, i_10_445_284_0, i_10_445_318_0,
    i_10_445_322_0, i_10_445_326_0, i_10_445_444_0, i_10_445_445_0,
    i_10_445_448_0, i_10_445_449_0, i_10_445_718_0, i_10_445_751_0,
    i_10_445_752_0, i_10_445_792_0, i_10_445_796_0, i_10_445_898_0,
    i_10_445_963_0, i_10_445_964_0, i_10_445_967_0, i_10_445_997_0,
    i_10_445_1002_0, i_10_445_1003_0, i_10_445_1084_0, i_10_445_1305_0,
    i_10_445_1306_0, i_10_445_1308_0, i_10_445_1437_0, i_10_445_1555_0,
    i_10_445_1580_0, i_10_445_1691_0, i_10_445_1768_0, i_10_445_1819_0,
    i_10_445_1821_0, i_10_445_1822_0, i_10_445_1823_0, i_10_445_1824_0,
    i_10_445_1948_0, i_10_445_2354_0, i_10_445_2362_0, i_10_445_2452_0,
    i_10_445_2453_0, i_10_445_2630_0, i_10_445_2632_0, i_10_445_2633_0,
    i_10_445_2704_0, i_10_445_2706_0, i_10_445_2707_0, i_10_445_2708_0,
    i_10_445_2715_0, i_10_445_2716_0, i_10_445_2717_0, i_10_445_2724_0,
    i_10_445_2725_0, i_10_445_2728_0, i_10_445_2734_0, i_10_445_2782_0,
    i_10_445_2829_0, i_10_445_2830_0, i_10_445_2919_0, i_10_445_2920_0,
    i_10_445_3034_0, i_10_445_3046_0, i_10_445_3076_0, i_10_445_3150_0,
    i_10_445_3154_0, i_10_445_3157_0, i_10_445_3389_0, i_10_445_3390_0,
    i_10_445_3405_0, i_10_445_3406_0, i_10_445_3468_0, i_10_445_3616_0,
    i_10_445_3649_0, i_10_445_3784_0, i_10_445_3787_0, i_10_445_3788_0,
    i_10_445_3815_0, i_10_445_3834_0, i_10_445_3842_0, i_10_445_3848_0,
    i_10_445_3853_0, i_10_445_3856_0, i_10_445_3888_0, i_10_445_3895_0,
    i_10_445_3982_0, i_10_445_3983_0, i_10_445_3985_0, i_10_445_3986_0,
    i_10_445_4116_0, i_10_445_4121_0, i_10_445_4266_0, i_10_445_4273_0,
    i_10_445_4284_0, i_10_445_4287_0, i_10_445_4290_0, i_10_445_4563_0;
  output o_10_445_0_0;
  assign o_10_445_0_0 = ~((~i_10_445_445_0 & ((~i_10_445_222_0 & ((~i_10_445_796_0 & ~i_10_445_997_0 & ~i_10_445_2452_0 & i_10_445_3853_0) | (~i_10_445_964_0 & ~i_10_445_2633_0 & ~i_10_445_3982_0 & i_10_445_4290_0 & ~i_10_445_4563_0))) | (~i_10_445_448_0 & ~i_10_445_964_0 & ~i_10_445_1819_0 & ~i_10_445_3405_0 & ~i_10_445_3468_0 & ~i_10_445_3856_0))) | (i_10_445_279_0 & ((~i_10_445_718_0 & ~i_10_445_964_0 & ~i_10_445_1822_0 & ~i_10_445_3046_0 & ~i_10_445_3468_0) | (i_10_445_1084_0 & ~i_10_445_4563_0))) | (~i_10_445_967_0 & ((~i_10_445_4563_0 & ((~i_10_445_284_0 & ((~i_10_445_898_0 & ~i_10_445_2630_0 & ~i_10_445_2725_0 & ~i_10_445_3034_0 & ~i_10_445_3848_0 & ~i_10_445_3888_0 & ~i_10_445_4284_0) | (i_10_445_2920_0 & ~i_10_445_3406_0 & ~i_10_445_4287_0))) | (~i_10_445_280_0 & i_10_445_1821_0 & ~i_10_445_2716_0 & ~i_10_445_3405_0 & ~i_10_445_3468_0 & ~i_10_445_4284_0))) | (~i_10_445_718_0 & ~i_10_445_4290_0 & ((~i_10_445_444_0 & ~i_10_445_1308_0 & ~i_10_445_2354_0 & ~i_10_445_2452_0 & ~i_10_445_2704_0 & ~i_10_445_2716_0 & ~i_10_445_3888_0) | (~i_10_445_220_0 & ~i_10_445_223_0 & ~i_10_445_964_0 & ~i_10_445_2920_0 & ~i_10_445_3405_0 & ~i_10_445_4287_0))) | (~i_10_445_2717_0 & ((~i_10_445_963_0 & ~i_10_445_1821_0 & i_10_445_3649_0) | (~i_10_445_752_0 & ~i_10_445_3405_0 & ~i_10_445_3406_0 & ~i_10_445_4116_0 & ~i_10_445_4284_0))))) | (~i_10_445_752_0 & ((~i_10_445_2728_0 & ~i_10_445_2734_0 & i_10_445_3787_0) | (i_10_445_1580_0 & ~i_10_445_2632_0 & ~i_10_445_4284_0))) | (~i_10_445_1822_0 & ((~i_10_445_220_0 & ~i_10_445_964_0 & ~i_10_445_1823_0 & ~i_10_445_2734_0 & ~i_10_445_2919_0 & ~i_10_445_3468_0) | (~i_10_445_223_0 & ~i_10_445_963_0 & ~i_10_445_2829_0 & ~i_10_445_3649_0 & ~i_10_445_3848_0 & ~i_10_445_4284_0))) | (~i_10_445_2728_0 & ((~i_10_445_220_0 & ((~i_10_445_223_0 & ~i_10_445_444_0 & ~i_10_445_718_0 & ~i_10_445_2632_0) | (~i_10_445_449_0 & ~i_10_445_963_0 & ~i_10_445_1002_0 & ~i_10_445_2633_0 & ~i_10_445_2920_0 & ~i_10_445_4116_0))) | (~i_10_445_223_0 & ~i_10_445_796_0 & ~i_10_445_964_0 & i_10_445_1819_0 & ~i_10_445_2782_0 & ~i_10_445_3405_0))) | (~i_10_445_796_0 & ((~i_10_445_444_0 & ~i_10_445_964_0 & ~i_10_445_2715_0 & ~i_10_445_2724_0 & ~i_10_445_2725_0 & ~i_10_445_2920_0 & ~i_10_445_3406_0) | (~i_10_445_898_0 & i_10_445_3853_0 & ~i_10_445_4284_0))) | (~i_10_445_963_0 & ((~i_10_445_444_0 & i_10_445_2630_0 & i_10_445_3842_0 & ~i_10_445_3888_0) | (~i_10_445_964_0 & i_10_445_967_0 & i_10_445_2633_0 & i_10_445_2704_0 & i_10_445_2920_0 & ~i_10_445_4116_0 & ~i_10_445_4287_0 & ~i_10_445_4290_0))) | (~i_10_445_444_0 & ((~i_10_445_2717_0 & i_10_445_2830_0 & ~i_10_445_3034_0) | (~i_10_445_1308_0 & ~i_10_445_1824_0 & ~i_10_445_2633_0 & ~i_10_445_2725_0 & i_10_445_3784_0))) | (~i_10_445_1821_0 & ~i_10_445_2453_0 & i_10_445_2704_0 & ~i_10_445_3034_0) | (i_10_445_280_0 & ~i_10_445_2717_0 & ~i_10_445_2724_0 & ~i_10_445_3405_0 & ~i_10_445_3468_0 & ~i_10_445_3788_0) | (i_10_445_2632_0 & i_10_445_2920_0 & i_10_445_3784_0 & i_10_445_3848_0) | (i_10_445_1580_0 & ~i_10_445_3856_0 & ~i_10_445_4116_0) | (i_10_445_318_0 & ~i_10_445_2919_0 & ~i_10_445_3842_0 & i_10_445_4284_0) | (i_10_445_3983_0 & i_10_445_4563_0));
endmodule



// Benchmark "kernel_10_446" written by ABC on Sun Jul 19 10:28:48 2020

module kernel_10_446 ( 
    i_10_446_32_0, i_10_446_34_0, i_10_446_35_0, i_10_446_124_0,
    i_10_446_125_0, i_10_446_156_0, i_10_446_160_0, i_10_446_178_0,
    i_10_446_248_0, i_10_446_258_0, i_10_446_323_0, i_10_446_431_0,
    i_10_446_519_0, i_10_446_520_0, i_10_446_565_0, i_10_446_566_0,
    i_10_446_628_0, i_10_446_958_0, i_10_446_961_0, i_10_446_962_0,
    i_10_446_996_0, i_10_446_1060_0, i_10_446_1061_0, i_10_446_1070_0,
    i_10_446_1124_0, i_10_446_1129_0, i_10_446_1165_0, i_10_446_1268_0,
    i_10_446_1309_0, i_10_446_1312_0, i_10_446_1347_0, i_10_446_1546_0,
    i_10_446_1555_0, i_10_446_1646_0, i_10_446_1650_0, i_10_446_1651_0,
    i_10_446_1654_0, i_10_446_1812_0, i_10_446_1815_0, i_10_446_1816_0,
    i_10_446_1908_0, i_10_446_1912_0, i_10_446_1914_0, i_10_446_1916_0,
    i_10_446_1952_0, i_10_446_1957_0, i_10_446_1958_0, i_10_446_1961_0,
    i_10_446_2037_0, i_10_446_2084_0, i_10_446_2242_0, i_10_446_2276_0,
    i_10_446_2384_0, i_10_446_2474_0, i_10_446_2481_0, i_10_446_2516_0,
    i_10_446_2632_0, i_10_446_2636_0, i_10_446_2713_0, i_10_446_2722_0,
    i_10_446_2725_0, i_10_446_2734_0, i_10_446_2787_0, i_10_446_2806_0,
    i_10_446_2887_0, i_10_446_3095_0, i_10_446_3166_0, i_10_446_3201_0,
    i_10_446_3286_0, i_10_446_3430_0, i_10_446_3433_0, i_10_446_3542_0,
    i_10_446_3616_0, i_10_446_3650_0, i_10_446_3651_0, i_10_446_3653_0,
    i_10_446_3704_0, i_10_446_3705_0, i_10_446_3718_0, i_10_446_3886_0,
    i_10_446_3887_0, i_10_446_3913_0, i_10_446_3984_0, i_10_446_3985_0,
    i_10_446_3991_0, i_10_446_3992_0, i_10_446_3994_0, i_10_446_3995_0,
    i_10_446_4053_0, i_10_446_4054_0, i_10_446_4057_0, i_10_446_4058_0,
    i_10_446_4118_0, i_10_446_4126_0, i_10_446_4129_0, i_10_446_4237_0,
    i_10_446_4271_0, i_10_446_4283_0, i_10_446_4400_0, i_10_446_4569_0,
    o_10_446_0_0  );
  input  i_10_446_32_0, i_10_446_34_0, i_10_446_35_0, i_10_446_124_0,
    i_10_446_125_0, i_10_446_156_0, i_10_446_160_0, i_10_446_178_0,
    i_10_446_248_0, i_10_446_258_0, i_10_446_323_0, i_10_446_431_0,
    i_10_446_519_0, i_10_446_520_0, i_10_446_565_0, i_10_446_566_0,
    i_10_446_628_0, i_10_446_958_0, i_10_446_961_0, i_10_446_962_0,
    i_10_446_996_0, i_10_446_1060_0, i_10_446_1061_0, i_10_446_1070_0,
    i_10_446_1124_0, i_10_446_1129_0, i_10_446_1165_0, i_10_446_1268_0,
    i_10_446_1309_0, i_10_446_1312_0, i_10_446_1347_0, i_10_446_1546_0,
    i_10_446_1555_0, i_10_446_1646_0, i_10_446_1650_0, i_10_446_1651_0,
    i_10_446_1654_0, i_10_446_1812_0, i_10_446_1815_0, i_10_446_1816_0,
    i_10_446_1908_0, i_10_446_1912_0, i_10_446_1914_0, i_10_446_1916_0,
    i_10_446_1952_0, i_10_446_1957_0, i_10_446_1958_0, i_10_446_1961_0,
    i_10_446_2037_0, i_10_446_2084_0, i_10_446_2242_0, i_10_446_2276_0,
    i_10_446_2384_0, i_10_446_2474_0, i_10_446_2481_0, i_10_446_2516_0,
    i_10_446_2632_0, i_10_446_2636_0, i_10_446_2713_0, i_10_446_2722_0,
    i_10_446_2725_0, i_10_446_2734_0, i_10_446_2787_0, i_10_446_2806_0,
    i_10_446_2887_0, i_10_446_3095_0, i_10_446_3166_0, i_10_446_3201_0,
    i_10_446_3286_0, i_10_446_3430_0, i_10_446_3433_0, i_10_446_3542_0,
    i_10_446_3616_0, i_10_446_3650_0, i_10_446_3651_0, i_10_446_3653_0,
    i_10_446_3704_0, i_10_446_3705_0, i_10_446_3718_0, i_10_446_3886_0,
    i_10_446_3887_0, i_10_446_3913_0, i_10_446_3984_0, i_10_446_3985_0,
    i_10_446_3991_0, i_10_446_3992_0, i_10_446_3994_0, i_10_446_3995_0,
    i_10_446_4053_0, i_10_446_4054_0, i_10_446_4057_0, i_10_446_4058_0,
    i_10_446_4118_0, i_10_446_4126_0, i_10_446_4129_0, i_10_446_4237_0,
    i_10_446_4271_0, i_10_446_4283_0, i_10_446_4400_0, i_10_446_4569_0;
  output o_10_446_0_0;
  assign o_10_446_0_0 = 0;
endmodule



// Benchmark "kernel_10_447" written by ABC on Sun Jul 19 10:28:49 2020

module kernel_10_447 ( 
    i_10_447_88_0, i_10_447_89_0, i_10_447_176_0, i_10_447_219_0,
    i_10_447_224_0, i_10_447_295_0, i_10_447_391_0, i_10_447_395_0,
    i_10_447_408_0, i_10_447_431_0, i_10_447_436_0, i_10_447_439_0,
    i_10_447_440_0, i_10_447_463_0, i_10_447_464_0, i_10_447_500_0,
    i_10_447_511_0, i_10_447_695_0, i_10_447_698_0, i_10_447_853_0,
    i_10_447_854_0, i_10_447_948_0, i_10_447_1027_0, i_10_447_1043_0,
    i_10_447_1056_0, i_10_447_1176_0, i_10_447_1238_0, i_10_447_1240_0,
    i_10_447_1245_0, i_10_447_1321_0, i_10_447_1345_0, i_10_447_1346_0,
    i_10_447_1448_0, i_10_447_1527_0, i_10_447_1552_0, i_10_447_1577_0,
    i_10_447_1649_0, i_10_447_1733_0, i_10_447_1735_0, i_10_447_1736_0,
    i_10_447_1804_0, i_10_447_1807_0, i_10_447_1888_0, i_10_447_2310_0,
    i_10_447_2312_0, i_10_447_2365_0, i_10_447_2374_0, i_10_447_2375_0,
    i_10_447_2451_0, i_10_447_2540_0, i_10_447_2543_0, i_10_447_2558_0,
    i_10_447_2561_0, i_10_447_2631_0, i_10_447_2632_0, i_10_447_2636_0,
    i_10_447_2645_0, i_10_447_2696_0, i_10_447_2714_0, i_10_447_2716_0,
    i_10_447_2733_0, i_10_447_2821_0, i_10_447_2852_0, i_10_447_2882_0,
    i_10_447_2885_0, i_10_447_2919_0, i_10_447_3197_0, i_10_447_3271_0,
    i_10_447_3278_0, i_10_447_3318_0, i_10_447_3319_0, i_10_447_3329_0,
    i_10_447_3356_0, i_10_447_3364_0, i_10_447_3390_0, i_10_447_3391_0,
    i_10_447_3406_0, i_10_447_3409_0, i_10_447_3463_0, i_10_447_3473_0,
    i_10_447_3499_0, i_10_447_3526_0, i_10_447_3620_0, i_10_447_3705_0,
    i_10_447_3706_0, i_10_447_3725_0, i_10_447_3839_0, i_10_447_3841_0,
    i_10_447_3854_0, i_10_447_3893_0, i_10_447_4031_0, i_10_447_4090_0,
    i_10_447_4115_0, i_10_447_4118_0, i_10_447_4129_0, i_10_447_4188_0,
    i_10_447_4277_0, i_10_447_4307_0, i_10_447_4564_0, i_10_447_4585_0,
    o_10_447_0_0  );
  input  i_10_447_88_0, i_10_447_89_0, i_10_447_176_0, i_10_447_219_0,
    i_10_447_224_0, i_10_447_295_0, i_10_447_391_0, i_10_447_395_0,
    i_10_447_408_0, i_10_447_431_0, i_10_447_436_0, i_10_447_439_0,
    i_10_447_440_0, i_10_447_463_0, i_10_447_464_0, i_10_447_500_0,
    i_10_447_511_0, i_10_447_695_0, i_10_447_698_0, i_10_447_853_0,
    i_10_447_854_0, i_10_447_948_0, i_10_447_1027_0, i_10_447_1043_0,
    i_10_447_1056_0, i_10_447_1176_0, i_10_447_1238_0, i_10_447_1240_0,
    i_10_447_1245_0, i_10_447_1321_0, i_10_447_1345_0, i_10_447_1346_0,
    i_10_447_1448_0, i_10_447_1527_0, i_10_447_1552_0, i_10_447_1577_0,
    i_10_447_1649_0, i_10_447_1733_0, i_10_447_1735_0, i_10_447_1736_0,
    i_10_447_1804_0, i_10_447_1807_0, i_10_447_1888_0, i_10_447_2310_0,
    i_10_447_2312_0, i_10_447_2365_0, i_10_447_2374_0, i_10_447_2375_0,
    i_10_447_2451_0, i_10_447_2540_0, i_10_447_2543_0, i_10_447_2558_0,
    i_10_447_2561_0, i_10_447_2631_0, i_10_447_2632_0, i_10_447_2636_0,
    i_10_447_2645_0, i_10_447_2696_0, i_10_447_2714_0, i_10_447_2716_0,
    i_10_447_2733_0, i_10_447_2821_0, i_10_447_2852_0, i_10_447_2882_0,
    i_10_447_2885_0, i_10_447_2919_0, i_10_447_3197_0, i_10_447_3271_0,
    i_10_447_3278_0, i_10_447_3318_0, i_10_447_3319_0, i_10_447_3329_0,
    i_10_447_3356_0, i_10_447_3364_0, i_10_447_3390_0, i_10_447_3391_0,
    i_10_447_3406_0, i_10_447_3409_0, i_10_447_3463_0, i_10_447_3473_0,
    i_10_447_3499_0, i_10_447_3526_0, i_10_447_3620_0, i_10_447_3705_0,
    i_10_447_3706_0, i_10_447_3725_0, i_10_447_3839_0, i_10_447_3841_0,
    i_10_447_3854_0, i_10_447_3893_0, i_10_447_4031_0, i_10_447_4090_0,
    i_10_447_4115_0, i_10_447_4118_0, i_10_447_4129_0, i_10_447_4188_0,
    i_10_447_4277_0, i_10_447_4307_0, i_10_447_4564_0, i_10_447_4585_0;
  output o_10_447_0_0;
  assign o_10_447_0_0 = 0;
endmodule



// Benchmark "kernel_10_448" written by ABC on Sun Jul 19 10:28:50 2020

module kernel_10_448 ( 
    i_10_448_83_0, i_10_448_117_0, i_10_448_152_0, i_10_448_176_0,
    i_10_448_182_0, i_10_448_217_0, i_10_448_279_0, i_10_448_406_0,
    i_10_448_408_0, i_10_448_443_0, i_10_448_445_0, i_10_448_446_0,
    i_10_448_460_0, i_10_448_461_0, i_10_448_463_0, i_10_448_464_0,
    i_10_448_509_0, i_10_448_515_0, i_10_448_686_0, i_10_448_747_0,
    i_10_448_754_0, i_10_448_794_0, i_10_448_795_0, i_10_448_967_0,
    i_10_448_1163_0, i_10_448_1212_0, i_10_448_1235_0, i_10_448_1237_0,
    i_10_448_1243_0, i_10_448_1244_0, i_10_448_1312_0, i_10_448_1361_0,
    i_10_448_1378_0, i_10_448_1487_0, i_10_448_1537_0, i_10_448_1562_0,
    i_10_448_1647_0, i_10_448_1651_0, i_10_448_1652_0, i_10_448_1684_0,
    i_10_448_1685_0, i_10_448_1688_0, i_10_448_1690_0, i_10_448_1768_0,
    i_10_448_1784_0, i_10_448_1808_0, i_10_448_1821_0, i_10_448_1822_0,
    i_10_448_1823_0, i_10_448_1824_0, i_10_448_1937_0, i_10_448_2033_0,
    i_10_448_2252_0, i_10_448_2391_0, i_10_448_2468_0, i_10_448_2509_0,
    i_10_448_2512_0, i_10_448_2631_0, i_10_448_2702_0, i_10_448_2716_0,
    i_10_448_2722_0, i_10_448_2723_0, i_10_448_2725_0, i_10_448_2726_0,
    i_10_448_2728_0, i_10_448_2731_0, i_10_448_2734_0, i_10_448_2735_0,
    i_10_448_2833_0, i_10_448_2916_0, i_10_448_2917_0, i_10_448_2920_0,
    i_10_448_2954_0, i_10_448_3034_0, i_10_448_3268_0, i_10_448_3326_0,
    i_10_448_3384_0, i_10_448_3524_0, i_10_448_3541_0, i_10_448_3586_0,
    i_10_448_3587_0, i_10_448_3645_0, i_10_448_3685_0, i_10_448_3797_0,
    i_10_448_3846_0, i_10_448_3847_0, i_10_448_3854_0, i_10_448_3859_0,
    i_10_448_3870_0, i_10_448_3880_0, i_10_448_3916_0, i_10_448_3961_0,
    i_10_448_4117_0, i_10_448_4118_0, i_10_448_4119_0, i_10_448_4140_0,
    i_10_448_4268_0, i_10_448_4285_0, i_10_448_4286_0, i_10_448_4288_0,
    o_10_448_0_0  );
  input  i_10_448_83_0, i_10_448_117_0, i_10_448_152_0, i_10_448_176_0,
    i_10_448_182_0, i_10_448_217_0, i_10_448_279_0, i_10_448_406_0,
    i_10_448_408_0, i_10_448_443_0, i_10_448_445_0, i_10_448_446_0,
    i_10_448_460_0, i_10_448_461_0, i_10_448_463_0, i_10_448_464_0,
    i_10_448_509_0, i_10_448_515_0, i_10_448_686_0, i_10_448_747_0,
    i_10_448_754_0, i_10_448_794_0, i_10_448_795_0, i_10_448_967_0,
    i_10_448_1163_0, i_10_448_1212_0, i_10_448_1235_0, i_10_448_1237_0,
    i_10_448_1243_0, i_10_448_1244_0, i_10_448_1312_0, i_10_448_1361_0,
    i_10_448_1378_0, i_10_448_1487_0, i_10_448_1537_0, i_10_448_1562_0,
    i_10_448_1647_0, i_10_448_1651_0, i_10_448_1652_0, i_10_448_1684_0,
    i_10_448_1685_0, i_10_448_1688_0, i_10_448_1690_0, i_10_448_1768_0,
    i_10_448_1784_0, i_10_448_1808_0, i_10_448_1821_0, i_10_448_1822_0,
    i_10_448_1823_0, i_10_448_1824_0, i_10_448_1937_0, i_10_448_2033_0,
    i_10_448_2252_0, i_10_448_2391_0, i_10_448_2468_0, i_10_448_2509_0,
    i_10_448_2512_0, i_10_448_2631_0, i_10_448_2702_0, i_10_448_2716_0,
    i_10_448_2722_0, i_10_448_2723_0, i_10_448_2725_0, i_10_448_2726_0,
    i_10_448_2728_0, i_10_448_2731_0, i_10_448_2734_0, i_10_448_2735_0,
    i_10_448_2833_0, i_10_448_2916_0, i_10_448_2917_0, i_10_448_2920_0,
    i_10_448_2954_0, i_10_448_3034_0, i_10_448_3268_0, i_10_448_3326_0,
    i_10_448_3384_0, i_10_448_3524_0, i_10_448_3541_0, i_10_448_3586_0,
    i_10_448_3587_0, i_10_448_3645_0, i_10_448_3685_0, i_10_448_3797_0,
    i_10_448_3846_0, i_10_448_3847_0, i_10_448_3854_0, i_10_448_3859_0,
    i_10_448_3870_0, i_10_448_3880_0, i_10_448_3916_0, i_10_448_3961_0,
    i_10_448_4117_0, i_10_448_4118_0, i_10_448_4119_0, i_10_448_4140_0,
    i_10_448_4268_0, i_10_448_4285_0, i_10_448_4286_0, i_10_448_4288_0;
  output o_10_448_0_0;
  assign o_10_448_0_0 = 0;
endmodule



// Benchmark "kernel_10_449" written by ABC on Sun Jul 19 10:28:51 2020

module kernel_10_449 ( 
    i_10_449_124_0, i_10_449_184_0, i_10_449_224_0, i_10_449_247_0,
    i_10_449_286_0, i_10_449_318_0, i_10_449_408_0, i_10_449_410_0,
    i_10_449_429_0, i_10_449_440_0, i_10_449_446_0, i_10_449_462_0,
    i_10_449_463_0, i_10_449_464_0, i_10_449_466_0, i_10_449_467_0,
    i_10_449_508_0, i_10_449_564_0, i_10_449_796_0, i_10_449_1005_0,
    i_10_449_1006_0, i_10_449_1033_0, i_10_449_1042_0, i_10_449_1043_0,
    i_10_449_1137_0, i_10_449_1138_0, i_10_449_1139_0, i_10_449_1236_0,
    i_10_449_1237_0, i_10_449_1239_0, i_10_449_1307_0, i_10_449_1308_0,
    i_10_449_1313_0, i_10_449_1366_0, i_10_449_1383_0, i_10_449_1384_0,
    i_10_449_1437_0, i_10_449_1653_0, i_10_449_1655_0, i_10_449_1821_0,
    i_10_449_1824_0, i_10_449_1909_0, i_10_449_1912_0, i_10_449_1913_0,
    i_10_449_1950_0, i_10_449_2094_0, i_10_449_2095_0, i_10_449_2350_0,
    i_10_449_2352_0, i_10_449_2356_0, i_10_449_2383_0, i_10_449_2384_0,
    i_10_449_2438_0, i_10_449_2471_0, i_10_449_2508_0, i_10_449_2514_0,
    i_10_449_2628_0, i_10_449_2631_0, i_10_449_2632_0, i_10_449_2634_0,
    i_10_449_2636_0, i_10_449_2655_0, i_10_449_2656_0, i_10_449_2660_0,
    i_10_449_2724_0, i_10_449_2829_0, i_10_449_2830_0, i_10_449_2831_0,
    i_10_449_2922_0, i_10_449_3039_0, i_10_449_3040_0, i_10_449_3154_0,
    i_10_449_3195_0, i_10_449_3197_0, i_10_449_3198_0, i_10_449_3199_0,
    i_10_449_3613_0, i_10_449_3614_0, i_10_449_3645_0, i_10_449_3649_0,
    i_10_449_3651_0, i_10_449_3652_0, i_10_449_3784_0, i_10_449_3788_0,
    i_10_449_3838_0, i_10_449_3847_0, i_10_449_3852_0, i_10_449_3853_0,
    i_10_449_3856_0, i_10_449_3895_0, i_10_449_3896_0, i_10_449_3967_0,
    i_10_449_4056_0, i_10_449_4117_0, i_10_449_4118_0, i_10_449_4120_0,
    i_10_449_4129_0, i_10_449_4278_0, i_10_449_4533_0, i_10_449_4567_0,
    o_10_449_0_0  );
  input  i_10_449_124_0, i_10_449_184_0, i_10_449_224_0, i_10_449_247_0,
    i_10_449_286_0, i_10_449_318_0, i_10_449_408_0, i_10_449_410_0,
    i_10_449_429_0, i_10_449_440_0, i_10_449_446_0, i_10_449_462_0,
    i_10_449_463_0, i_10_449_464_0, i_10_449_466_0, i_10_449_467_0,
    i_10_449_508_0, i_10_449_564_0, i_10_449_796_0, i_10_449_1005_0,
    i_10_449_1006_0, i_10_449_1033_0, i_10_449_1042_0, i_10_449_1043_0,
    i_10_449_1137_0, i_10_449_1138_0, i_10_449_1139_0, i_10_449_1236_0,
    i_10_449_1237_0, i_10_449_1239_0, i_10_449_1307_0, i_10_449_1308_0,
    i_10_449_1313_0, i_10_449_1366_0, i_10_449_1383_0, i_10_449_1384_0,
    i_10_449_1437_0, i_10_449_1653_0, i_10_449_1655_0, i_10_449_1821_0,
    i_10_449_1824_0, i_10_449_1909_0, i_10_449_1912_0, i_10_449_1913_0,
    i_10_449_1950_0, i_10_449_2094_0, i_10_449_2095_0, i_10_449_2350_0,
    i_10_449_2352_0, i_10_449_2356_0, i_10_449_2383_0, i_10_449_2384_0,
    i_10_449_2438_0, i_10_449_2471_0, i_10_449_2508_0, i_10_449_2514_0,
    i_10_449_2628_0, i_10_449_2631_0, i_10_449_2632_0, i_10_449_2634_0,
    i_10_449_2636_0, i_10_449_2655_0, i_10_449_2656_0, i_10_449_2660_0,
    i_10_449_2724_0, i_10_449_2829_0, i_10_449_2830_0, i_10_449_2831_0,
    i_10_449_2922_0, i_10_449_3039_0, i_10_449_3040_0, i_10_449_3154_0,
    i_10_449_3195_0, i_10_449_3197_0, i_10_449_3198_0, i_10_449_3199_0,
    i_10_449_3613_0, i_10_449_3614_0, i_10_449_3645_0, i_10_449_3649_0,
    i_10_449_3651_0, i_10_449_3652_0, i_10_449_3784_0, i_10_449_3788_0,
    i_10_449_3838_0, i_10_449_3847_0, i_10_449_3852_0, i_10_449_3853_0,
    i_10_449_3856_0, i_10_449_3895_0, i_10_449_3896_0, i_10_449_3967_0,
    i_10_449_4056_0, i_10_449_4117_0, i_10_449_4118_0, i_10_449_4120_0,
    i_10_449_4129_0, i_10_449_4278_0, i_10_449_4533_0, i_10_449_4567_0;
  output o_10_449_0_0;
  assign o_10_449_0_0 = ~((~i_10_449_408_0 & ((~i_10_449_429_0 & ~i_10_449_1307_0 & ~i_10_449_2632_0 & ~i_10_449_2831_0 & ~i_10_449_3195_0 & ~i_10_449_3198_0) | (~i_10_449_124_0 & ~i_10_449_1042_0 & ~i_10_449_1043_0 & i_10_449_2830_0 & ~i_10_449_3197_0 & ~i_10_449_4056_0))) | (~i_10_449_124_0 & ((~i_10_449_184_0 & ~i_10_449_1437_0 & ~i_10_449_1913_0 & ~i_10_449_2830_0 & ~i_10_449_3197_0) | (~i_10_449_1909_0 & ~i_10_449_3199_0 & ~i_10_449_3784_0 & ~i_10_449_3856_0))) | (~i_10_449_1043_0 & ((~i_10_449_410_0 & ((~i_10_449_1236_0 & i_10_449_2628_0 & ~i_10_449_3199_0 & ~i_10_449_3651_0) | (~i_10_449_1912_0 & ~i_10_449_2656_0 & i_10_449_2922_0 & i_10_449_3197_0 & ~i_10_449_3852_0))) | (~i_10_449_1006_0 & ~i_10_449_3040_0 & ((~i_10_449_1913_0 & i_10_449_2636_0) | (~i_10_449_1821_0 & ~i_10_449_2831_0 & ~i_10_449_3852_0))) | (i_10_449_440_0 & ~i_10_449_1237_0 & i_10_449_3853_0) | (~i_10_449_440_0 & ~i_10_449_462_0 & ~i_10_449_3853_0) | (~i_10_449_184_0 & ~i_10_449_446_0 & ~i_10_449_464_0 & ~i_10_449_1950_0 & ~i_10_449_2829_0 & ~i_10_449_3895_0))) | (~i_10_449_429_0 & ((~i_10_449_466_0 & ~i_10_449_1236_0 & ~i_10_449_2632_0 & i_10_449_3199_0 & ~i_10_449_3852_0 & ~i_10_449_3853_0) | (i_10_449_466_0 & ~i_10_449_1308_0 & ~i_10_449_3197_0 & ~i_10_449_3784_0 & ~i_10_449_3838_0 & ~i_10_449_4567_0))) | (~i_10_449_184_0 & ((~i_10_449_564_0 & ((~i_10_449_1912_0 & ~i_10_449_2830_0 & ~i_10_449_3039_0 & ~i_10_449_3198_0) | (~i_10_449_446_0 & ~i_10_449_1307_0 & ~i_10_449_1437_0 & ~i_10_449_1909_0 & i_10_449_2631_0 & i_10_449_2632_0 & ~i_10_449_3896_0))) | (~i_10_449_1912_0 & ~i_10_449_2656_0 & ~i_10_449_3039_0 & i_10_449_3613_0 & ~i_10_449_3856_0))) | (~i_10_449_1042_0 & ((~i_10_449_463_0 & ~i_10_449_464_0 & ~i_10_449_2829_0 & ~i_10_449_3853_0) | (~i_10_449_1655_0 & ~i_10_449_1912_0 & ~i_10_449_2471_0 & ~i_10_449_2660_0 & ~i_10_449_3198_0 & ~i_10_449_4056_0))) | (~i_10_449_1236_0 & ((~i_10_449_1239_0 & ~i_10_449_1366_0 & ~i_10_449_1821_0 & ~i_10_449_2831_0 & ~i_10_449_3197_0 & i_10_449_3649_0 & ~i_10_449_3896_0) | (~i_10_449_1307_0 & i_10_449_2632_0 & i_10_449_4117_0))) | (~i_10_449_1239_0 & ((i_10_449_440_0 & ~i_10_449_1912_0 & ~i_10_449_1950_0 & i_10_449_3613_0 & i_10_449_3852_0 & i_10_449_3853_0) | (~i_10_449_4117_0 & i_10_449_4118_0))) | (~i_10_449_1308_0 & ((~i_10_449_3040_0 & ~i_10_449_3614_0) | (~i_10_449_2471_0 & ~i_10_449_2831_0 & i_10_449_3856_0 & ~i_10_449_3895_0))) | (~i_10_449_3652_0 & ((~i_10_449_318_0 & ~i_10_449_1437_0 & ~i_10_449_3614_0 & ~i_10_449_3896_0) | i_10_449_4120_0 | (i_10_449_796_0 & i_10_449_2632_0 & ~i_10_449_2660_0 & ~i_10_449_3195_0 & ~i_10_449_3852_0 & ~i_10_449_3856_0 & i_10_449_3895_0 & ~i_10_449_4567_0))) | (~i_10_449_1909_0 & ~i_10_449_1913_0 & i_10_449_2628_0 & ~i_10_449_3838_0 & ~i_10_449_3853_0 & ~i_10_449_4056_0));
endmodule



// Benchmark "kernel_10_450" written by ABC on Sun Jul 19 10:28:52 2020

module kernel_10_450 ( 
    i_10_450_250_0, i_10_450_251_0, i_10_450_282_0, i_10_450_331_0,
    i_10_450_411_0, i_10_450_412_0, i_10_450_447_0, i_10_450_511_0,
    i_10_450_597_0, i_10_450_794_0, i_10_450_795_0, i_10_450_1030_0,
    i_10_450_1080_0, i_10_450_1083_0, i_10_450_1138_0, i_10_450_1139_0,
    i_10_450_1142_0, i_10_450_1236_0, i_10_450_1240_0, i_10_450_1243_0,
    i_10_450_1305_0, i_10_450_1306_0, i_10_450_1308_0, i_10_450_1309_0,
    i_10_450_1310_0, i_10_450_1312_0, i_10_450_1365_0, i_10_450_1367_0,
    i_10_450_1444_0, i_10_450_1653_0, i_10_450_1687_0, i_10_450_1688_0,
    i_10_450_1767_0, i_10_450_1818_0, i_10_450_1913_0, i_10_450_2158_0,
    i_10_450_2403_0, i_10_450_2406_0, i_10_450_2407_0, i_10_450_2408_0,
    i_10_450_2454_0, i_10_450_2455_0, i_10_450_2456_0, i_10_450_2479_0,
    i_10_450_2518_0, i_10_450_2604_0, i_10_450_2632_0, i_10_450_2634_0,
    i_10_450_2636_0, i_10_450_2658_0, i_10_450_2659_0, i_10_450_2660_0,
    i_10_450_2679_0, i_10_450_2680_0, i_10_450_2681_0, i_10_450_2703_0,
    i_10_450_2726_0, i_10_450_2732_0, i_10_450_2783_0, i_10_450_2784_0,
    i_10_450_2785_0, i_10_450_2787_0, i_10_450_2788_0, i_10_450_2831_0,
    i_10_450_2919_0, i_10_450_3049_0, i_10_450_3150_0, i_10_450_3154_0,
    i_10_450_3277_0, i_10_450_3280_0, i_10_450_3283_0, i_10_450_3385_0,
    i_10_450_3387_0, i_10_450_3388_0, i_10_450_3389_0, i_10_450_3391_0,
    i_10_450_3392_0, i_10_450_3406_0, i_10_450_3494_0, i_10_450_3613_0,
    i_10_450_3650_0, i_10_450_3652_0, i_10_450_3785_0, i_10_450_3835_0,
    i_10_450_3839_0, i_10_450_3841_0, i_10_450_3855_0, i_10_450_3856_0,
    i_10_450_3981_0, i_10_450_4029_0, i_10_450_4054_0, i_10_450_4055_0,
    i_10_450_4056_0, i_10_450_4057_0, i_10_450_4270_0, i_10_450_4284_0,
    i_10_450_4285_0, i_10_450_4288_0, i_10_450_4292_0, i_10_450_4565_0,
    o_10_450_0_0  );
  input  i_10_450_250_0, i_10_450_251_0, i_10_450_282_0, i_10_450_331_0,
    i_10_450_411_0, i_10_450_412_0, i_10_450_447_0, i_10_450_511_0,
    i_10_450_597_0, i_10_450_794_0, i_10_450_795_0, i_10_450_1030_0,
    i_10_450_1080_0, i_10_450_1083_0, i_10_450_1138_0, i_10_450_1139_0,
    i_10_450_1142_0, i_10_450_1236_0, i_10_450_1240_0, i_10_450_1243_0,
    i_10_450_1305_0, i_10_450_1306_0, i_10_450_1308_0, i_10_450_1309_0,
    i_10_450_1310_0, i_10_450_1312_0, i_10_450_1365_0, i_10_450_1367_0,
    i_10_450_1444_0, i_10_450_1653_0, i_10_450_1687_0, i_10_450_1688_0,
    i_10_450_1767_0, i_10_450_1818_0, i_10_450_1913_0, i_10_450_2158_0,
    i_10_450_2403_0, i_10_450_2406_0, i_10_450_2407_0, i_10_450_2408_0,
    i_10_450_2454_0, i_10_450_2455_0, i_10_450_2456_0, i_10_450_2479_0,
    i_10_450_2518_0, i_10_450_2604_0, i_10_450_2632_0, i_10_450_2634_0,
    i_10_450_2636_0, i_10_450_2658_0, i_10_450_2659_0, i_10_450_2660_0,
    i_10_450_2679_0, i_10_450_2680_0, i_10_450_2681_0, i_10_450_2703_0,
    i_10_450_2726_0, i_10_450_2732_0, i_10_450_2783_0, i_10_450_2784_0,
    i_10_450_2785_0, i_10_450_2787_0, i_10_450_2788_0, i_10_450_2831_0,
    i_10_450_2919_0, i_10_450_3049_0, i_10_450_3150_0, i_10_450_3154_0,
    i_10_450_3277_0, i_10_450_3280_0, i_10_450_3283_0, i_10_450_3385_0,
    i_10_450_3387_0, i_10_450_3388_0, i_10_450_3389_0, i_10_450_3391_0,
    i_10_450_3392_0, i_10_450_3406_0, i_10_450_3494_0, i_10_450_3613_0,
    i_10_450_3650_0, i_10_450_3652_0, i_10_450_3785_0, i_10_450_3835_0,
    i_10_450_3839_0, i_10_450_3841_0, i_10_450_3855_0, i_10_450_3856_0,
    i_10_450_3981_0, i_10_450_4029_0, i_10_450_4054_0, i_10_450_4055_0,
    i_10_450_4056_0, i_10_450_4057_0, i_10_450_4270_0, i_10_450_4284_0,
    i_10_450_4285_0, i_10_450_4288_0, i_10_450_4292_0, i_10_450_4565_0;
  output o_10_450_0_0;
  assign o_10_450_0_0 = ~((~i_10_450_447_0 & ((~i_10_450_1080_0 & i_10_450_2456_0 & ~i_10_450_2788_0) | (~i_10_450_1913_0 & ~i_10_450_2726_0 & ~i_10_450_2784_0 & ~i_10_450_3389_0 & ~i_10_450_4055_0))) | (~i_10_450_1365_0 & ((~i_10_450_411_0 & ~i_10_450_1083_0 & ~i_10_450_1367_0 & ~i_10_450_1818_0 & ~i_10_450_3841_0 & ~i_10_450_4029_0) | (~i_10_450_2784_0 & ~i_10_450_3856_0 & ~i_10_450_3981_0 & ~i_10_450_4054_0))) | (~i_10_450_1767_0 & ((~i_10_450_331_0 & ~i_10_450_2408_0 & ~i_10_450_3049_0 & ~i_10_450_3981_0 & ~i_10_450_4029_0) | (~i_10_450_250_0 & ~i_10_450_2732_0 & ~i_10_450_3839_0 & ~i_10_450_4054_0 & ~i_10_450_4057_0))) | (~i_10_450_4056_0 & ((~i_10_450_2407_0 & ((~i_10_450_1312_0 & ~i_10_450_3835_0 & ~i_10_450_3981_0) | (~i_10_450_2680_0 & ~i_10_450_4057_0))) | (~i_10_450_1308_0 & ~i_10_450_2604_0 & ~i_10_450_4057_0 & ~i_10_450_4288_0))) | (i_10_450_3835_0 & ((i_10_450_2632_0 & ~i_10_450_2783_0 & ~i_10_450_2785_0 & ~i_10_450_3280_0) | (i_10_450_2783_0 & ~i_10_450_3049_0 & ~i_10_450_3839_0 & ~i_10_450_4057_0))) | (~i_10_450_1236_0 & ~i_10_450_1444_0 & ~i_10_450_2788_0) | (~i_10_450_2660_0 & ~i_10_450_2787_0 & ~i_10_450_2831_0) | (i_10_450_2456_0 & ~i_10_450_3855_0));
endmodule



// Benchmark "kernel_10_451" written by ABC on Sun Jul 19 10:28:53 2020

module kernel_10_451 ( 
    i_10_451_12_0, i_10_451_174_0, i_10_451_177_0, i_10_451_253_0,
    i_10_451_256_0, i_10_451_261_0, i_10_451_264_0, i_10_451_265_0,
    i_10_451_285_0, i_10_451_286_0, i_10_451_318_0, i_10_451_391_0,
    i_10_451_444_0, i_10_451_460_0, i_10_451_504_0, i_10_451_792_0,
    i_10_451_867_0, i_10_451_999_0, i_10_451_1002_0, i_10_451_1029_0,
    i_10_451_1056_0, i_10_451_1101_0, i_10_451_1104_0, i_10_451_1296_0,
    i_10_451_1299_0, i_10_451_1302_0, i_10_451_1344_0, i_10_451_1347_0,
    i_10_451_1431_0, i_10_451_1434_0, i_10_451_1542_0, i_10_451_1543_0,
    i_10_451_1545_0, i_10_451_1546_0, i_10_451_1575_0, i_10_451_1620_0,
    i_10_451_1623_0, i_10_451_1649_0, i_10_451_1683_0, i_10_451_1686_0,
    i_10_451_1729_0, i_10_451_1731_0, i_10_451_1819_0, i_10_451_1824_0,
    i_10_451_1980_0, i_10_451_2016_0, i_10_451_2028_0, i_10_451_2202_0,
    i_10_451_2349_0, i_10_451_2352_0, i_10_451_2529_0, i_10_451_2532_0,
    i_10_451_2565_0, i_10_451_2568_0, i_10_451_2677_0, i_10_451_2678_0,
    i_10_451_2703_0, i_10_451_2743_0, i_10_451_2820_0, i_10_451_2847_0,
    i_10_451_2881_0, i_10_451_2883_0, i_10_451_2967_0, i_10_451_3045_0,
    i_10_451_3072_0, i_10_451_3267_0, i_10_451_3277_0, i_10_451_3280_0,
    i_10_451_3281_0, i_10_451_3312_0, i_10_451_3390_0, i_10_451_3391_0,
    i_10_451_3471_0, i_10_451_3473_0, i_10_451_3537_0, i_10_451_3540_0,
    i_10_451_3541_0, i_10_451_3543_0, i_10_451_3544_0, i_10_451_3582_0,
    i_10_451_3585_0, i_10_451_3621_0, i_10_451_3652_0, i_10_451_3687_0,
    i_10_451_3795_0, i_10_451_3834_0, i_10_451_3837_0, i_10_451_3842_0,
    i_10_451_3847_0, i_10_451_3850_0, i_10_451_4116_0, i_10_451_4117_0,
    i_10_451_4167_0, i_10_451_4170_0, i_10_451_4275_0, i_10_451_4281_0,
    i_10_451_4287_0, i_10_451_4290_0, i_10_451_4563_0, i_10_451_4585_0,
    o_10_451_0_0  );
  input  i_10_451_12_0, i_10_451_174_0, i_10_451_177_0, i_10_451_253_0,
    i_10_451_256_0, i_10_451_261_0, i_10_451_264_0, i_10_451_265_0,
    i_10_451_285_0, i_10_451_286_0, i_10_451_318_0, i_10_451_391_0,
    i_10_451_444_0, i_10_451_460_0, i_10_451_504_0, i_10_451_792_0,
    i_10_451_867_0, i_10_451_999_0, i_10_451_1002_0, i_10_451_1029_0,
    i_10_451_1056_0, i_10_451_1101_0, i_10_451_1104_0, i_10_451_1296_0,
    i_10_451_1299_0, i_10_451_1302_0, i_10_451_1344_0, i_10_451_1347_0,
    i_10_451_1431_0, i_10_451_1434_0, i_10_451_1542_0, i_10_451_1543_0,
    i_10_451_1545_0, i_10_451_1546_0, i_10_451_1575_0, i_10_451_1620_0,
    i_10_451_1623_0, i_10_451_1649_0, i_10_451_1683_0, i_10_451_1686_0,
    i_10_451_1729_0, i_10_451_1731_0, i_10_451_1819_0, i_10_451_1824_0,
    i_10_451_1980_0, i_10_451_2016_0, i_10_451_2028_0, i_10_451_2202_0,
    i_10_451_2349_0, i_10_451_2352_0, i_10_451_2529_0, i_10_451_2532_0,
    i_10_451_2565_0, i_10_451_2568_0, i_10_451_2677_0, i_10_451_2678_0,
    i_10_451_2703_0, i_10_451_2743_0, i_10_451_2820_0, i_10_451_2847_0,
    i_10_451_2881_0, i_10_451_2883_0, i_10_451_2967_0, i_10_451_3045_0,
    i_10_451_3072_0, i_10_451_3267_0, i_10_451_3277_0, i_10_451_3280_0,
    i_10_451_3281_0, i_10_451_3312_0, i_10_451_3390_0, i_10_451_3391_0,
    i_10_451_3471_0, i_10_451_3473_0, i_10_451_3537_0, i_10_451_3540_0,
    i_10_451_3541_0, i_10_451_3543_0, i_10_451_3544_0, i_10_451_3582_0,
    i_10_451_3585_0, i_10_451_3621_0, i_10_451_3652_0, i_10_451_3687_0,
    i_10_451_3795_0, i_10_451_3834_0, i_10_451_3837_0, i_10_451_3842_0,
    i_10_451_3847_0, i_10_451_3850_0, i_10_451_4116_0, i_10_451_4117_0,
    i_10_451_4167_0, i_10_451_4170_0, i_10_451_4275_0, i_10_451_4281_0,
    i_10_451_4287_0, i_10_451_4290_0, i_10_451_4563_0, i_10_451_4585_0;
  output o_10_451_0_0;
  assign o_10_451_0_0 = 0;
endmodule



// Benchmark "kernel_10_452" written by ABC on Sun Jul 19 10:28:54 2020

module kernel_10_452 ( 
    i_10_452_31_0, i_10_452_33_0, i_10_452_67_0, i_10_452_171_0,
    i_10_452_184_0, i_10_452_212_0, i_10_452_283_0, i_10_452_390_0,
    i_10_452_391_0, i_10_452_405_0, i_10_452_406_0, i_10_452_435_0,
    i_10_452_436_0, i_10_452_439_0, i_10_452_514_0, i_10_452_718_0,
    i_10_452_750_0, i_10_452_1002_0, i_10_452_1030_0, i_10_452_1035_0,
    i_10_452_1038_0, i_10_452_1056_0, i_10_452_1164_0, i_10_452_1261_0,
    i_10_452_1262_0, i_10_452_1264_0, i_10_452_1287_0, i_10_452_1305_0,
    i_10_452_1351_0, i_10_452_1362_0, i_10_452_1363_0, i_10_452_1364_0,
    i_10_452_1366_0, i_10_452_1367_0, i_10_452_1435_0, i_10_452_1542_0,
    i_10_452_1554_0, i_10_452_1606_0, i_10_452_1635_0, i_10_452_1768_0,
    i_10_452_1804_0, i_10_452_1825_0, i_10_452_1872_0, i_10_452_1913_0,
    i_10_452_2041_0, i_10_452_2091_0, i_10_452_2143_0, i_10_452_2196_0,
    i_10_452_2356_0, i_10_452_2374_0, i_10_452_2407_0, i_10_452_2448_0,
    i_10_452_2453_0, i_10_452_2470_0, i_10_452_2512_0, i_10_452_2514_0,
    i_10_452_2526_0, i_10_452_2605_0, i_10_452_2700_0, i_10_452_2722_0,
    i_10_452_2734_0, i_10_452_2754_0, i_10_452_2785_0, i_10_452_2820_0,
    i_10_452_2821_0, i_10_452_2957_0, i_10_452_2982_0, i_10_452_2983_0,
    i_10_452_3033_0, i_10_452_3036_0, i_10_452_3046_0, i_10_452_3234_0,
    i_10_452_3237_0, i_10_452_3268_0, i_10_452_3271_0, i_10_452_3319_0,
    i_10_452_3390_0, i_10_452_3393_0, i_10_452_3586_0, i_10_452_3652_0,
    i_10_452_3653_0, i_10_452_3663_0, i_10_452_3702_0, i_10_452_3717_0,
    i_10_452_3718_0, i_10_452_3719_0, i_10_452_3834_0, i_10_452_3835_0,
    i_10_452_3853_0, i_10_452_3856_0, i_10_452_3982_0, i_10_452_4053_0,
    i_10_452_4174_0, i_10_452_4276_0, i_10_452_4278_0, i_10_452_4373_0,
    i_10_452_4485_0, i_10_452_4528_0, i_10_452_4534_0, i_10_452_4569_0,
    o_10_452_0_0  );
  input  i_10_452_31_0, i_10_452_33_0, i_10_452_67_0, i_10_452_171_0,
    i_10_452_184_0, i_10_452_212_0, i_10_452_283_0, i_10_452_390_0,
    i_10_452_391_0, i_10_452_405_0, i_10_452_406_0, i_10_452_435_0,
    i_10_452_436_0, i_10_452_439_0, i_10_452_514_0, i_10_452_718_0,
    i_10_452_750_0, i_10_452_1002_0, i_10_452_1030_0, i_10_452_1035_0,
    i_10_452_1038_0, i_10_452_1056_0, i_10_452_1164_0, i_10_452_1261_0,
    i_10_452_1262_0, i_10_452_1264_0, i_10_452_1287_0, i_10_452_1305_0,
    i_10_452_1351_0, i_10_452_1362_0, i_10_452_1363_0, i_10_452_1364_0,
    i_10_452_1366_0, i_10_452_1367_0, i_10_452_1435_0, i_10_452_1542_0,
    i_10_452_1554_0, i_10_452_1606_0, i_10_452_1635_0, i_10_452_1768_0,
    i_10_452_1804_0, i_10_452_1825_0, i_10_452_1872_0, i_10_452_1913_0,
    i_10_452_2041_0, i_10_452_2091_0, i_10_452_2143_0, i_10_452_2196_0,
    i_10_452_2356_0, i_10_452_2374_0, i_10_452_2407_0, i_10_452_2448_0,
    i_10_452_2453_0, i_10_452_2470_0, i_10_452_2512_0, i_10_452_2514_0,
    i_10_452_2526_0, i_10_452_2605_0, i_10_452_2700_0, i_10_452_2722_0,
    i_10_452_2734_0, i_10_452_2754_0, i_10_452_2785_0, i_10_452_2820_0,
    i_10_452_2821_0, i_10_452_2957_0, i_10_452_2982_0, i_10_452_2983_0,
    i_10_452_3033_0, i_10_452_3036_0, i_10_452_3046_0, i_10_452_3234_0,
    i_10_452_3237_0, i_10_452_3268_0, i_10_452_3271_0, i_10_452_3319_0,
    i_10_452_3390_0, i_10_452_3393_0, i_10_452_3586_0, i_10_452_3652_0,
    i_10_452_3653_0, i_10_452_3663_0, i_10_452_3702_0, i_10_452_3717_0,
    i_10_452_3718_0, i_10_452_3719_0, i_10_452_3834_0, i_10_452_3835_0,
    i_10_452_3853_0, i_10_452_3856_0, i_10_452_3982_0, i_10_452_4053_0,
    i_10_452_4174_0, i_10_452_4276_0, i_10_452_4278_0, i_10_452_4373_0,
    i_10_452_4485_0, i_10_452_4528_0, i_10_452_4534_0, i_10_452_4569_0;
  output o_10_452_0_0;
  assign o_10_452_0_0 = 0;
endmodule



// Benchmark "kernel_10_453" written by ABC on Sun Jul 19 10:28:55 2020

module kernel_10_453 ( 
    i_10_453_70_0, i_10_453_180_0, i_10_453_181_0, i_10_453_281_0,
    i_10_453_282_0, i_10_453_372_0, i_10_453_407_0, i_10_453_429_0,
    i_10_453_430_0, i_10_453_441_0, i_10_453_442_0, i_10_453_443_0,
    i_10_453_444_0, i_10_453_461_0, i_10_453_464_0, i_10_453_520_0,
    i_10_453_536_0, i_10_453_590_0, i_10_453_629_0, i_10_453_735_0,
    i_10_453_797_0, i_10_453_826_0, i_10_453_967_0, i_10_453_1238_0,
    i_10_453_1243_0, i_10_453_1263_0, i_10_453_1309_0, i_10_453_1321_0,
    i_10_453_1359_0, i_10_453_1581_0, i_10_453_1616_0, i_10_453_1691_0,
    i_10_453_1755_0, i_10_453_1757_0, i_10_453_1805_0, i_10_453_1821_0,
    i_10_453_1823_0, i_10_453_1912_0, i_10_453_1913_0, i_10_453_2083_0,
    i_10_453_2087_0, i_10_453_2159_0, i_10_453_2184_0, i_10_453_2229_0,
    i_10_453_2312_0, i_10_453_2326_0, i_10_453_2327_0, i_10_453_2350_0,
    i_10_453_2408_0, i_10_453_2440_0, i_10_453_2449_0, i_10_453_2453_0,
    i_10_453_2455_0, i_10_453_2456_0, i_10_453_2471_0, i_10_453_2635_0,
    i_10_453_2636_0, i_10_453_2662_0, i_10_453_2663_0, i_10_453_2701_0,
    i_10_453_2704_0, i_10_453_2725_0, i_10_453_2728_0, i_10_453_2729_0,
    i_10_453_2731_0, i_10_453_2831_0, i_10_453_2862_0, i_10_453_2886_0,
    i_10_453_3035_0, i_10_453_3093_0, i_10_453_3094_0, i_10_453_3202_0,
    i_10_453_3234_0, i_10_453_3277_0, i_10_453_3405_0, i_10_453_3409_0,
    i_10_453_3526_0, i_10_453_3527_0, i_10_453_3688_0, i_10_453_3782_0,
    i_10_453_3859_0, i_10_453_3949_0, i_10_453_3980_0, i_10_453_3981_0,
    i_10_453_3982_0, i_10_453_4120_0, i_10_453_4182_0, i_10_453_4185_0,
    i_10_453_4189_0, i_10_453_4190_0, i_10_453_4267_0, i_10_453_4269_0,
    i_10_453_4270_0, i_10_453_4271_0, i_10_453_4274_0, i_10_453_4287_0,
    i_10_453_4458_0, i_10_453_4549_0, i_10_453_4550_0, i_10_453_4571_0,
    o_10_453_0_0  );
  input  i_10_453_70_0, i_10_453_180_0, i_10_453_181_0, i_10_453_281_0,
    i_10_453_282_0, i_10_453_372_0, i_10_453_407_0, i_10_453_429_0,
    i_10_453_430_0, i_10_453_441_0, i_10_453_442_0, i_10_453_443_0,
    i_10_453_444_0, i_10_453_461_0, i_10_453_464_0, i_10_453_520_0,
    i_10_453_536_0, i_10_453_590_0, i_10_453_629_0, i_10_453_735_0,
    i_10_453_797_0, i_10_453_826_0, i_10_453_967_0, i_10_453_1238_0,
    i_10_453_1243_0, i_10_453_1263_0, i_10_453_1309_0, i_10_453_1321_0,
    i_10_453_1359_0, i_10_453_1581_0, i_10_453_1616_0, i_10_453_1691_0,
    i_10_453_1755_0, i_10_453_1757_0, i_10_453_1805_0, i_10_453_1821_0,
    i_10_453_1823_0, i_10_453_1912_0, i_10_453_1913_0, i_10_453_2083_0,
    i_10_453_2087_0, i_10_453_2159_0, i_10_453_2184_0, i_10_453_2229_0,
    i_10_453_2312_0, i_10_453_2326_0, i_10_453_2327_0, i_10_453_2350_0,
    i_10_453_2408_0, i_10_453_2440_0, i_10_453_2449_0, i_10_453_2453_0,
    i_10_453_2455_0, i_10_453_2456_0, i_10_453_2471_0, i_10_453_2635_0,
    i_10_453_2636_0, i_10_453_2662_0, i_10_453_2663_0, i_10_453_2701_0,
    i_10_453_2704_0, i_10_453_2725_0, i_10_453_2728_0, i_10_453_2729_0,
    i_10_453_2731_0, i_10_453_2831_0, i_10_453_2862_0, i_10_453_2886_0,
    i_10_453_3035_0, i_10_453_3093_0, i_10_453_3094_0, i_10_453_3202_0,
    i_10_453_3234_0, i_10_453_3277_0, i_10_453_3405_0, i_10_453_3409_0,
    i_10_453_3526_0, i_10_453_3527_0, i_10_453_3688_0, i_10_453_3782_0,
    i_10_453_3859_0, i_10_453_3949_0, i_10_453_3980_0, i_10_453_3981_0,
    i_10_453_3982_0, i_10_453_4120_0, i_10_453_4182_0, i_10_453_4185_0,
    i_10_453_4189_0, i_10_453_4190_0, i_10_453_4267_0, i_10_453_4269_0,
    i_10_453_4270_0, i_10_453_4271_0, i_10_453_4274_0, i_10_453_4287_0,
    i_10_453_4458_0, i_10_453_4549_0, i_10_453_4550_0, i_10_453_4571_0;
  output o_10_453_0_0;
  assign o_10_453_0_0 = 0;
endmodule



// Benchmark "kernel_10_454" written by ABC on Sun Jul 19 10:28:56 2020

module kernel_10_454 ( 
    i_10_454_171_0, i_10_454_172_0, i_10_454_173_0, i_10_454_175_0,
    i_10_454_176_0, i_10_454_283_0, i_10_454_285_0, i_10_454_320_0,
    i_10_454_321_0, i_10_454_405_0, i_10_454_407_0, i_10_454_433_0,
    i_10_454_435_0, i_10_454_443_0, i_10_454_444_0, i_10_454_445_0,
    i_10_454_461_0, i_10_454_466_0, i_10_454_467_0, i_10_454_505_0,
    i_10_454_518_0, i_10_454_718_0, i_10_454_719_0, i_10_454_960_0,
    i_10_454_962_0, i_10_454_967_0, i_10_454_968_0, i_10_454_1233_0,
    i_10_454_1236_0, i_10_454_1237_0, i_10_454_1240_0, i_10_454_1250_0,
    i_10_454_1306_0, i_10_454_1310_0, i_10_454_1311_0, i_10_454_1579_0,
    i_10_454_1581_0, i_10_454_1653_0, i_10_454_1654_0, i_10_454_1688_0,
    i_10_454_1817_0, i_10_454_1818_0, i_10_454_1819_0, i_10_454_1823_0,
    i_10_454_1825_0, i_10_454_2203_0, i_10_454_2332_0, i_10_454_2338_0,
    i_10_454_2350_0, i_10_454_2363_0, i_10_454_2377_0, i_10_454_2380_0,
    i_10_454_2383_0, i_10_454_2461_0, i_10_454_2462_0, i_10_454_2471_0,
    i_10_454_2633_0, i_10_454_2636_0, i_10_454_2658_0, i_10_454_2659_0,
    i_10_454_2660_0, i_10_454_2700_0, i_10_454_2708_0, i_10_454_2724_0,
    i_10_454_2731_0, i_10_454_2735_0, i_10_454_2881_0, i_10_454_2920_0,
    i_10_454_2921_0, i_10_454_3152_0, i_10_454_3154_0, i_10_454_3322_0,
    i_10_454_3325_0, i_10_454_3385_0, i_10_454_3469_0, i_10_454_3472_0,
    i_10_454_3497_0, i_10_454_3586_0, i_10_454_3612_0, i_10_454_3613_0,
    i_10_454_3616_0, i_10_454_3782_0, i_10_454_3783_0, i_10_454_3847_0,
    i_10_454_3848_0, i_10_454_3853_0, i_10_454_3854_0, i_10_454_3986_0,
    i_10_454_4117_0, i_10_454_4174_0, i_10_454_4267_0, i_10_454_4268_0,
    i_10_454_4270_0, i_10_454_4271_0, i_10_454_4285_0, i_10_454_4286_0,
    i_10_454_4564_0, i_10_454_4566_0, i_10_454_4567_0, i_10_454_4568_0,
    o_10_454_0_0  );
  input  i_10_454_171_0, i_10_454_172_0, i_10_454_173_0, i_10_454_175_0,
    i_10_454_176_0, i_10_454_283_0, i_10_454_285_0, i_10_454_320_0,
    i_10_454_321_0, i_10_454_405_0, i_10_454_407_0, i_10_454_433_0,
    i_10_454_435_0, i_10_454_443_0, i_10_454_444_0, i_10_454_445_0,
    i_10_454_461_0, i_10_454_466_0, i_10_454_467_0, i_10_454_505_0,
    i_10_454_518_0, i_10_454_718_0, i_10_454_719_0, i_10_454_960_0,
    i_10_454_962_0, i_10_454_967_0, i_10_454_968_0, i_10_454_1233_0,
    i_10_454_1236_0, i_10_454_1237_0, i_10_454_1240_0, i_10_454_1250_0,
    i_10_454_1306_0, i_10_454_1310_0, i_10_454_1311_0, i_10_454_1579_0,
    i_10_454_1581_0, i_10_454_1653_0, i_10_454_1654_0, i_10_454_1688_0,
    i_10_454_1817_0, i_10_454_1818_0, i_10_454_1819_0, i_10_454_1823_0,
    i_10_454_1825_0, i_10_454_2203_0, i_10_454_2332_0, i_10_454_2338_0,
    i_10_454_2350_0, i_10_454_2363_0, i_10_454_2377_0, i_10_454_2380_0,
    i_10_454_2383_0, i_10_454_2461_0, i_10_454_2462_0, i_10_454_2471_0,
    i_10_454_2633_0, i_10_454_2636_0, i_10_454_2658_0, i_10_454_2659_0,
    i_10_454_2660_0, i_10_454_2700_0, i_10_454_2708_0, i_10_454_2724_0,
    i_10_454_2731_0, i_10_454_2735_0, i_10_454_2881_0, i_10_454_2920_0,
    i_10_454_2921_0, i_10_454_3152_0, i_10_454_3154_0, i_10_454_3322_0,
    i_10_454_3325_0, i_10_454_3385_0, i_10_454_3469_0, i_10_454_3472_0,
    i_10_454_3497_0, i_10_454_3586_0, i_10_454_3612_0, i_10_454_3613_0,
    i_10_454_3616_0, i_10_454_3782_0, i_10_454_3783_0, i_10_454_3847_0,
    i_10_454_3848_0, i_10_454_3853_0, i_10_454_3854_0, i_10_454_3986_0,
    i_10_454_4117_0, i_10_454_4174_0, i_10_454_4267_0, i_10_454_4268_0,
    i_10_454_4270_0, i_10_454_4271_0, i_10_454_4285_0, i_10_454_4286_0,
    i_10_454_4564_0, i_10_454_4566_0, i_10_454_4567_0, i_10_454_4568_0;
  output o_10_454_0_0;
  assign o_10_454_0_0 = ~((~i_10_454_4567_0 & ((~i_10_454_2735_0 & ((~i_10_454_283_0 & ((~i_10_454_172_0 & ~i_10_454_968_0 & i_10_454_1688_0 & ~i_10_454_2350_0 & ~i_10_454_2383_0) | (i_10_454_2921_0 & i_10_454_3854_0 & ~i_10_454_4564_0))) | (~i_10_454_2363_0 & ~i_10_454_2636_0 & i_10_454_3613_0 & ~i_10_454_3782_0 & ~i_10_454_4271_0 & ~i_10_454_4286_0))) | (~i_10_454_445_0 & ((~i_10_454_176_0 & i_10_454_1819_0 & ~i_10_454_1825_0 & ~i_10_454_2380_0 & ~i_10_454_3848_0) | (~i_10_454_407_0 & i_10_454_1310_0 & ~i_10_454_1817_0 & ~i_10_454_2731_0 & ~i_10_454_2921_0 & ~i_10_454_3586_0 & ~i_10_454_3853_0))) | (i_10_454_283_0 & i_10_454_1306_0 & ~i_10_454_3848_0 & ~i_10_454_4267_0) | (~i_10_454_175_0 & ~i_10_454_461_0 & ~i_10_454_718_0 & ~i_10_454_968_0 & ~i_10_454_1310_0 & ~i_10_454_1579_0 & ~i_10_454_1818_0 & ~i_10_454_2363_0 & ~i_10_454_2383_0 & ~i_10_454_2881_0 & ~i_10_454_4268_0 & ~i_10_454_4271_0) | (~i_10_454_444_0 & ~i_10_454_719_0 & ~i_10_454_1250_0 & ~i_10_454_2338_0 & i_10_454_2660_0 & ~i_10_454_4286_0))) | (~i_10_454_4268_0 & ((~i_10_454_719_0 & ~i_10_454_967_0 & ((~i_10_454_176_0 & ~i_10_454_962_0 & ((~i_10_454_444_0 & ~i_10_454_2735_0 & ~i_10_454_2920_0 & ~i_10_454_2921_0 & ~i_10_454_4267_0 & ~i_10_454_4271_0) | (i_10_454_2203_0 & ~i_10_454_2383_0 & ~i_10_454_4568_0))) | (~i_10_454_1823_0 & i_10_454_1825_0 & ~i_10_454_2380_0 & ~i_10_454_4271_0))) | (~i_10_454_445_0 & ((~i_10_454_2363_0 & ~i_10_454_2633_0 & ~i_10_454_2881_0 & i_10_454_3385_0 & ~i_10_454_4270_0 & ~i_10_454_4271_0 & ~i_10_454_4566_0) | (i_10_454_1240_0 & ~i_10_454_1581_0 & ~i_10_454_2380_0 & ~i_10_454_2700_0 & ~i_10_454_4568_0))) | (~i_10_454_3848_0 & ((i_10_454_405_0 & i_10_454_1654_0 & ~i_10_454_2380_0 & ~i_10_454_3497_0) | (~i_10_454_2636_0 & i_10_454_3853_0 & ~i_10_454_4117_0))) | (~i_10_454_320_0 & ~i_10_454_1823_0 & ~i_10_454_1825_0 & ~i_10_454_2338_0 & ~i_10_454_2377_0 & ~i_10_454_2462_0 & i_10_454_3854_0))) | (i_10_454_285_0 & ((~i_10_454_967_0 & ~i_10_454_1310_0 & i_10_454_2731_0 & ~i_10_454_3848_0 & ~i_10_454_4270_0) | (~i_10_454_2636_0 & ~i_10_454_2921_0 & ~i_10_454_3783_0 & ~i_10_454_3847_0 & ~i_10_454_4566_0))) | (~i_10_454_285_0 & ((i_10_454_433_0 & ~i_10_454_461_0 & ~i_10_454_1823_0 & ~i_10_454_2332_0 & ~i_10_454_2636_0 & ~i_10_454_4117_0) | (i_10_454_1581_0 & ~i_10_454_4270_0 & ~i_10_454_4285_0 & ~i_10_454_4566_0))) | (~i_10_454_4267_0 & ((~i_10_454_518_0 & ((~i_10_454_433_0 & ~i_10_454_968_0 & ~i_10_454_1310_0 & ~i_10_454_2380_0 & i_10_454_3848_0 & ~i_10_454_4270_0 & i_10_454_4564_0) | (i_10_454_171_0 & ~i_10_454_1653_0 & ~i_10_454_2377_0 & ~i_10_454_4286_0 & ~i_10_454_4566_0))) | (~i_10_454_968_0 & i_10_454_3385_0 & i_10_454_3616_0 & ~i_10_454_4271_0) | (~i_10_454_719_0 & ~i_10_454_1823_0 & ~i_10_454_2383_0 & ~i_10_454_3385_0 & ~i_10_454_3469_0 & ~i_10_454_4270_0 & ~i_10_454_4285_0 & i_10_454_4566_0))) | (~i_10_454_718_0 & ((i_10_454_1237_0 & ~i_10_454_2380_0 & i_10_454_2658_0) | (~i_10_454_967_0 & ~i_10_454_2383_0 & ~i_10_454_2920_0 & ~i_10_454_3385_0 & ~i_10_454_4271_0 & i_10_454_4566_0))) | (~i_10_454_1250_0 & ((~i_10_454_719_0 & ~i_10_454_2921_0 & ~i_10_454_3469_0 & i_10_454_3616_0) | (i_10_454_176_0 & ~i_10_454_445_0 & ~i_10_454_1579_0 & i_10_454_2708_0 & ~i_10_454_3847_0))) | (~i_10_454_445_0 & ((i_10_454_466_0 & i_10_454_1825_0 & i_10_454_3613_0) | (i_10_454_443_0 & ~i_10_454_2338_0 & i_10_454_3854_0))) | (~i_10_454_719_0 & ((i_10_454_2708_0 & ~i_10_454_3613_0 & i_10_454_4117_0 & ~i_10_454_4271_0) | (i_10_454_1250_0 & ~i_10_454_1823_0 & ~i_10_454_3848_0 & ~i_10_454_4286_0))) | (~i_10_454_968_0 & ((i_10_454_1818_0 & ((i_10_454_1240_0 & i_10_454_1819_0 & ~i_10_454_3472_0) | (~i_10_454_967_0 & i_10_454_1306_0 & ~i_10_454_4568_0))) | (i_10_454_3783_0 & ((~i_10_454_1581_0 & i_10_454_4117_0 & ~i_10_454_4270_0 & ~i_10_454_4271_0) | (~i_10_454_1688_0 & ~i_10_454_2350_0 & ~i_10_454_2363_0 & ~i_10_454_4566_0))))) | (~i_10_454_2471_0 & ((i_10_454_2203_0 & ~i_10_454_2920_0 & ~i_10_454_3847_0) | (~i_10_454_1823_0 & i_10_454_2658_0 & i_10_454_2660_0 & i_10_454_4117_0))) | (~i_10_454_2724_0 & ((i_10_454_435_0 & ~i_10_454_2350_0) | (~i_10_454_1654_0 & ~i_10_454_2881_0 & i_10_454_3612_0 & ~i_10_454_3848_0))) | (i_10_454_3613_0 & ((i_10_454_2920_0 & i_10_454_3782_0 & i_10_454_4117_0) | (~i_10_454_1579_0 & i_10_454_1654_0 & ~i_10_454_2633_0 & ~i_10_454_2735_0 & ~i_10_454_4117_0 & ~i_10_454_4271_0) | (i_10_454_433_0 & i_10_454_3385_0 & ~i_10_454_4568_0))));
endmodule



// Benchmark "kernel_10_455" written by ABC on Sun Jul 19 10:28:58 2020

module kernel_10_455 ( 
    i_10_455_246_0, i_10_455_249_0, i_10_455_273_0, i_10_455_276_0,
    i_10_455_289_0, i_10_455_294_0, i_10_455_295_0, i_10_455_324_0,
    i_10_455_328_0, i_10_455_330_0, i_10_455_438_0, i_10_455_459_0,
    i_10_455_462_0, i_10_455_463_0, i_10_455_464_0, i_10_455_465_0,
    i_10_455_531_0, i_10_455_534_0, i_10_455_993_0, i_10_455_996_0,
    i_10_455_1000_0, i_10_455_1038_0, i_10_455_1039_0, i_10_455_1041_0,
    i_10_455_1238_0, i_10_455_1240_0, i_10_455_1241_0, i_10_455_1267_0,
    i_10_455_1308_0, i_10_455_1312_0, i_10_455_1344_0, i_10_455_1350_0,
    i_10_455_1435_0, i_10_455_1441_0, i_10_455_1443_0, i_10_455_1446_0,
    i_10_455_1488_0, i_10_455_1546_0, i_10_455_1648_0, i_10_455_1683_0,
    i_10_455_1689_0, i_10_455_1713_0, i_10_455_1818_0, i_10_455_1872_0,
    i_10_455_1946_0, i_10_455_2250_0, i_10_455_2322_0, i_10_455_2325_0,
    i_10_455_2349_0, i_10_455_2351_0, i_10_455_2361_0, i_10_455_2364_0,
    i_10_455_2377_0, i_10_455_2460_0, i_10_455_2469_0, i_10_455_2505_0,
    i_10_455_2607_0, i_10_455_2634_0, i_10_455_2636_0, i_10_455_2658_0,
    i_10_455_2661_0, i_10_455_2676_0, i_10_455_2703_0, i_10_455_2706_0,
    i_10_455_2715_0, i_10_455_2721_0, i_10_455_2724_0, i_10_455_2730_0,
    i_10_455_2781_0, i_10_455_2806_0, i_10_455_2829_0, i_10_455_2831_0,
    i_10_455_2832_0, i_10_455_2834_0, i_10_455_2881_0, i_10_455_2918_0,
    i_10_455_3036_0, i_10_455_3037_0, i_10_455_3039_0, i_10_455_3045_0,
    i_10_455_3153_0, i_10_455_3165_0, i_10_455_3274_0, i_10_455_3281_0,
    i_10_455_3291_0, i_10_455_3403_0, i_10_455_3408_0, i_10_455_3492_0,
    i_10_455_3609_0, i_10_455_3610_0, i_10_455_3616_0, i_10_455_3617_0,
    i_10_455_3849_0, i_10_455_3982_0, i_10_455_3994_0, i_10_455_4028_0,
    i_10_455_4128_0, i_10_455_4291_0, i_10_455_4564_0, i_10_455_4568_0,
    o_10_455_0_0  );
  input  i_10_455_246_0, i_10_455_249_0, i_10_455_273_0, i_10_455_276_0,
    i_10_455_289_0, i_10_455_294_0, i_10_455_295_0, i_10_455_324_0,
    i_10_455_328_0, i_10_455_330_0, i_10_455_438_0, i_10_455_459_0,
    i_10_455_462_0, i_10_455_463_0, i_10_455_464_0, i_10_455_465_0,
    i_10_455_531_0, i_10_455_534_0, i_10_455_993_0, i_10_455_996_0,
    i_10_455_1000_0, i_10_455_1038_0, i_10_455_1039_0, i_10_455_1041_0,
    i_10_455_1238_0, i_10_455_1240_0, i_10_455_1241_0, i_10_455_1267_0,
    i_10_455_1308_0, i_10_455_1312_0, i_10_455_1344_0, i_10_455_1350_0,
    i_10_455_1435_0, i_10_455_1441_0, i_10_455_1443_0, i_10_455_1446_0,
    i_10_455_1488_0, i_10_455_1546_0, i_10_455_1648_0, i_10_455_1683_0,
    i_10_455_1689_0, i_10_455_1713_0, i_10_455_1818_0, i_10_455_1872_0,
    i_10_455_1946_0, i_10_455_2250_0, i_10_455_2322_0, i_10_455_2325_0,
    i_10_455_2349_0, i_10_455_2351_0, i_10_455_2361_0, i_10_455_2364_0,
    i_10_455_2377_0, i_10_455_2460_0, i_10_455_2469_0, i_10_455_2505_0,
    i_10_455_2607_0, i_10_455_2634_0, i_10_455_2636_0, i_10_455_2658_0,
    i_10_455_2661_0, i_10_455_2676_0, i_10_455_2703_0, i_10_455_2706_0,
    i_10_455_2715_0, i_10_455_2721_0, i_10_455_2724_0, i_10_455_2730_0,
    i_10_455_2781_0, i_10_455_2806_0, i_10_455_2829_0, i_10_455_2831_0,
    i_10_455_2832_0, i_10_455_2834_0, i_10_455_2881_0, i_10_455_2918_0,
    i_10_455_3036_0, i_10_455_3037_0, i_10_455_3039_0, i_10_455_3045_0,
    i_10_455_3153_0, i_10_455_3165_0, i_10_455_3274_0, i_10_455_3281_0,
    i_10_455_3291_0, i_10_455_3403_0, i_10_455_3408_0, i_10_455_3492_0,
    i_10_455_3609_0, i_10_455_3610_0, i_10_455_3616_0, i_10_455_3617_0,
    i_10_455_3849_0, i_10_455_3982_0, i_10_455_3994_0, i_10_455_4028_0,
    i_10_455_4128_0, i_10_455_4291_0, i_10_455_4564_0, i_10_455_4568_0;
  output o_10_455_0_0;
  assign o_10_455_0_0 = ~((~i_10_455_246_0 & ((i_10_455_462_0 & ~i_10_455_2834_0 & ~i_10_455_3408_0) | (~i_10_455_295_0 & ~i_10_455_324_0 & ~i_10_455_996_0 & ~i_10_455_1041_0 & ~i_10_455_1488_0 & ~i_10_455_2460_0 & ~i_10_455_2881_0 & ~i_10_455_3994_0))) | (~i_10_455_294_0 & ((~i_10_455_1308_0 & i_10_455_1818_0 & ~i_10_455_3609_0 & ~i_10_455_3849_0) | (~i_10_455_438_0 & ~i_10_455_1038_0 & ~i_10_455_1872_0 & ~i_10_455_2322_0 & ~i_10_455_2607_0 & ~i_10_455_2881_0 & ~i_10_455_3408_0 & ~i_10_455_3982_0 & ~i_10_455_4128_0))) | (~i_10_455_2325_0 & ((~i_10_455_289_0 & ((~i_10_455_295_0 & ~i_10_455_2661_0 & ~i_10_455_2676_0 & ~i_10_455_2706_0 & ~i_10_455_2918_0 & ~i_10_455_3403_0 & ~i_10_455_3616_0) | (~i_10_455_324_0 & ~i_10_455_330_0 & ~i_10_455_438_0 & ~i_10_455_1446_0 & ~i_10_455_1488_0 & ~i_10_455_2377_0 & ~i_10_455_3045_0 & ~i_10_455_3408_0 & ~i_10_455_3994_0))) | (~i_10_455_330_0 & ~i_10_455_993_0 & ~i_10_455_1039_0 & ~i_10_455_1344_0 & ~i_10_455_2377_0 & ~i_10_455_2831_0 & ~i_10_455_3045_0 & ~i_10_455_3609_0 & ~i_10_455_4128_0))) | (~i_10_455_996_0 & ((~i_10_455_993_0 & ((~i_10_455_1038_0 & ~i_10_455_1443_0 & ~i_10_455_2364_0 & ~i_10_455_2832_0) | (~i_10_455_289_0 & ~i_10_455_1039_0 & ~i_10_455_1267_0 & i_10_455_2634_0 & ~i_10_455_2703_0 & ~i_10_455_2881_0 & ~i_10_455_4128_0))) | (~i_10_455_249_0 & ~i_10_455_1041_0 & ~i_10_455_2377_0 & ~i_10_455_2781_0 & ~i_10_455_2881_0 & ~i_10_455_3036_0 & ~i_10_455_3039_0 & ~i_10_455_3165_0 & ~i_10_455_3281_0 & ~i_10_455_3403_0 & ~i_10_455_3982_0))) | (~i_10_455_1038_0 & ((~i_10_455_438_0 & ~i_10_455_1312_0 & ~i_10_455_2715_0 & ~i_10_455_2781_0 & i_10_455_2829_0 & ~i_10_455_3610_0 & ~i_10_455_3994_0) | (~i_10_455_2703_0 & ~i_10_455_2721_0 & ~i_10_455_3616_0 & ~i_10_455_4028_0))) | (i_10_455_3982_0 & ~i_10_455_3994_0 & ~i_10_455_4028_0 & ~i_10_455_4564_0 & i_10_455_4568_0));
endmodule



// Benchmark "kernel_10_456" written by ABC on Sun Jul 19 10:28:59 2020

module kernel_10_456 ( 
    i_10_456_221_0, i_10_456_224_0, i_10_456_319_0, i_10_456_320_0,
    i_10_456_322_0, i_10_456_323_0, i_10_456_329_0, i_10_456_436_0,
    i_10_456_447_0, i_10_456_465_0, i_10_456_466_0, i_10_456_508_0,
    i_10_456_898_0, i_10_456_1004_0, i_10_456_1005_0, i_10_456_1083_0,
    i_10_456_1084_0, i_10_456_1085_0, i_10_456_1086_0, i_10_456_1087_0,
    i_10_456_1088_0, i_10_456_1240_0, i_10_456_1241_0, i_10_456_1242_0,
    i_10_456_1246_0, i_10_456_1249_0, i_10_456_1263_0, i_10_456_1309_0,
    i_10_456_1313_0, i_10_456_1651_0, i_10_456_1652_0, i_10_456_2352_0,
    i_10_456_2382_0, i_10_456_2407_0, i_10_456_2470_0, i_10_456_2509_0,
    i_10_456_2510_0, i_10_456_2629_0, i_10_456_2661_0, i_10_456_2700_0,
    i_10_456_2701_0, i_10_456_2703_0, i_10_456_2704_0, i_10_456_2706_0,
    i_10_456_2707_0, i_10_456_2711_0, i_10_456_2726_0, i_10_456_2782_0,
    i_10_456_2783_0, i_10_456_2785_0, i_10_456_2786_0, i_10_456_2789_0,
    i_10_456_2885_0, i_10_456_2919_0, i_10_456_2920_0, i_10_456_2922_0,
    i_10_456_2923_0, i_10_456_2924_0, i_10_456_2959_0, i_10_456_2987_0,
    i_10_456_3153_0, i_10_456_3279_0, i_10_456_3281_0, i_10_456_3385_0,
    i_10_456_3389_0, i_10_456_3391_0, i_10_456_3406_0, i_10_456_3407_0,
    i_10_456_3408_0, i_10_456_3409_0, i_10_456_3472_0, i_10_456_3496_0,
    i_10_456_3497_0, i_10_456_3586_0, i_10_456_3616_0, i_10_456_3646_0,
    i_10_456_3649_0, i_10_456_3650_0, i_10_456_3653_0, i_10_456_3784_0,
    i_10_456_3786_0, i_10_456_3788_0, i_10_456_3847_0, i_10_456_3848_0,
    i_10_456_3854_0, i_10_456_3860_0, i_10_456_3978_0, i_10_456_3979_0,
    i_10_456_3980_0, i_10_456_3983_0, i_10_456_3985_0, i_10_456_3986_0,
    i_10_456_4057_0, i_10_456_4113_0, i_10_456_4128_0, i_10_456_4130_0,
    i_10_456_4236_0, i_10_456_4237_0, i_10_456_4288_0, i_10_456_4289_0,
    o_10_456_0_0  );
  input  i_10_456_221_0, i_10_456_224_0, i_10_456_319_0, i_10_456_320_0,
    i_10_456_322_0, i_10_456_323_0, i_10_456_329_0, i_10_456_436_0,
    i_10_456_447_0, i_10_456_465_0, i_10_456_466_0, i_10_456_508_0,
    i_10_456_898_0, i_10_456_1004_0, i_10_456_1005_0, i_10_456_1083_0,
    i_10_456_1084_0, i_10_456_1085_0, i_10_456_1086_0, i_10_456_1087_0,
    i_10_456_1088_0, i_10_456_1240_0, i_10_456_1241_0, i_10_456_1242_0,
    i_10_456_1246_0, i_10_456_1249_0, i_10_456_1263_0, i_10_456_1309_0,
    i_10_456_1313_0, i_10_456_1651_0, i_10_456_1652_0, i_10_456_2352_0,
    i_10_456_2382_0, i_10_456_2407_0, i_10_456_2470_0, i_10_456_2509_0,
    i_10_456_2510_0, i_10_456_2629_0, i_10_456_2661_0, i_10_456_2700_0,
    i_10_456_2701_0, i_10_456_2703_0, i_10_456_2704_0, i_10_456_2706_0,
    i_10_456_2707_0, i_10_456_2711_0, i_10_456_2726_0, i_10_456_2782_0,
    i_10_456_2783_0, i_10_456_2785_0, i_10_456_2786_0, i_10_456_2789_0,
    i_10_456_2885_0, i_10_456_2919_0, i_10_456_2920_0, i_10_456_2922_0,
    i_10_456_2923_0, i_10_456_2924_0, i_10_456_2959_0, i_10_456_2987_0,
    i_10_456_3153_0, i_10_456_3279_0, i_10_456_3281_0, i_10_456_3385_0,
    i_10_456_3389_0, i_10_456_3391_0, i_10_456_3406_0, i_10_456_3407_0,
    i_10_456_3408_0, i_10_456_3409_0, i_10_456_3472_0, i_10_456_3496_0,
    i_10_456_3497_0, i_10_456_3586_0, i_10_456_3616_0, i_10_456_3646_0,
    i_10_456_3649_0, i_10_456_3650_0, i_10_456_3653_0, i_10_456_3784_0,
    i_10_456_3786_0, i_10_456_3788_0, i_10_456_3847_0, i_10_456_3848_0,
    i_10_456_3854_0, i_10_456_3860_0, i_10_456_3978_0, i_10_456_3979_0,
    i_10_456_3980_0, i_10_456_3983_0, i_10_456_3985_0, i_10_456_3986_0,
    i_10_456_4057_0, i_10_456_4113_0, i_10_456_4128_0, i_10_456_4130_0,
    i_10_456_4236_0, i_10_456_4237_0, i_10_456_4288_0, i_10_456_4289_0;
  output o_10_456_0_0;
  assign o_10_456_0_0 = ~((~i_10_456_4057_0 & ((~i_10_456_322_0 & ((~i_10_456_466_0 & ~i_10_456_1084_0 & ~i_10_456_1263_0 & ~i_10_456_2704_0 & ~i_10_456_3497_0 & ~i_10_456_3646_0 & ~i_10_456_3860_0) | (~i_10_456_1083_0 & ~i_10_456_1313_0 & ~i_10_456_1652_0 & ~i_10_456_3653_0 & ~i_10_456_3854_0 & ~i_10_456_3983_0 & ~i_10_456_3985_0 & ~i_10_456_4236_0 & ~i_10_456_4237_0))) | (~i_10_456_1083_0 & ((~i_10_456_1087_0 & ~i_10_456_2707_0 & ~i_10_456_2782_0 & i_10_456_3385_0 & ~i_10_456_3649_0) | (~i_10_456_320_0 & ~i_10_456_1004_0 & ~i_10_456_1085_0 & ~i_10_456_1088_0 & ~i_10_456_2352_0 & ~i_10_456_2470_0 & ~i_10_456_2509_0 & ~i_10_456_2510_0 & ~i_10_456_2706_0 & ~i_10_456_3854_0 & ~i_10_456_4128_0))) | (~i_10_456_319_0 & ~i_10_456_1309_0 & ~i_10_456_1313_0 & i_10_456_3854_0 & ~i_10_456_3978_0 & ~i_10_456_3986_0 & ~i_10_456_4113_0 & ~i_10_456_4236_0 & ~i_10_456_4237_0))) | (~i_10_456_1086_0 & ~i_10_456_2789_0 & ((~i_10_456_319_0 & ((~i_10_456_323_0 & ~i_10_456_1005_0 & ~i_10_456_1083_0 & ~i_10_456_1084_0 & ~i_10_456_1085_0 & ~i_10_456_2407_0 & ~i_10_456_3985_0 & ~i_10_456_3986_0 & ~i_10_456_4128_0) | (~i_10_456_221_0 & ~i_10_456_447_0 & ~i_10_456_1088_0 & ~i_10_456_1263_0 & ~i_10_456_2510_0 & ~i_10_456_2701_0 & ~i_10_456_2703_0 & ~i_10_456_2785_0 & ~i_10_456_3854_0 & ~i_10_456_3978_0 & ~i_10_456_4130_0))) | (~i_10_456_1084_0 & ~i_10_456_2382_0 & ~i_10_456_2726_0 & ~i_10_456_2783_0 & ~i_10_456_3472_0 & ~i_10_456_3496_0 & ~i_10_456_3616_0 & ~i_10_456_3653_0 & ~i_10_456_3848_0 & ~i_10_456_3978_0 & ~i_10_456_3979_0 & ~i_10_456_3985_0 & ~i_10_456_3986_0 & ~i_10_456_4237_0))) | (~i_10_456_323_0 & ~i_10_456_2700_0 & ((~i_10_456_1083_0 & ~i_10_456_1084_0 & i_10_456_2407_0 & ~i_10_456_2783_0 & i_10_456_3979_0) | (~i_10_456_1004_0 & ~i_10_456_2382_0 & ~i_10_456_2629_0 & ~i_10_456_2707_0 & ~i_10_456_2785_0 & ~i_10_456_3788_0 & ~i_10_456_3854_0 & ~i_10_456_3860_0 & ~i_10_456_3979_0 & ~i_10_456_4236_0))) | (~i_10_456_1083_0 & ((~i_10_456_1241_0 & ((~i_10_456_1084_0 & ~i_10_456_1088_0 & ~i_10_456_1240_0 & ~i_10_456_1263_0 & ~i_10_456_2707_0 & ~i_10_456_2726_0 & ~i_10_456_3650_0 & ~i_10_456_3979_0) | (~i_10_456_1087_0 & i_10_456_2923_0 & ~i_10_456_4237_0))) | (~i_10_456_329_0 & i_10_456_2629_0 & i_10_456_2923_0 & ~i_10_456_3496_0))) | (~i_10_456_1087_0 & ((~i_10_456_329_0 & ((~i_10_456_2885_0 & i_10_456_2920_0 & ~i_10_456_2987_0 & ~i_10_456_3586_0) | (~i_10_456_436_0 & ~i_10_456_1263_0 & ~i_10_456_1309_0 & i_10_456_1651_0 & ~i_10_456_2509_0 & ~i_10_456_2629_0 & ~i_10_456_3496_0 & ~i_10_456_3854_0 & ~i_10_456_3860_0 & ~i_10_456_3986_0))) | (~i_10_456_1088_0 & ~i_10_456_1263_0 & ~i_10_456_2706_0 & ~i_10_456_2786_0 & i_10_456_2924_0 & ~i_10_456_3985_0))) | (~i_10_456_320_0 & ((~i_10_456_436_0 & ~i_10_456_2661_0 & ~i_10_456_3983_0 & ((i_10_456_2629_0 & ~i_10_456_2786_0 & ~i_10_456_3978_0 & ~i_10_456_3985_0) | (~i_10_456_1084_0 & ~i_10_456_1085_0 & ~i_10_456_2352_0 & ~i_10_456_2470_0 & ~i_10_456_2703_0 & ~i_10_456_2785_0 & ~i_10_456_3860_0 & ~i_10_456_3986_0))) | (~i_10_456_2470_0 & ~i_10_456_3649_0 & i_10_456_3847_0))) | (~i_10_456_3653_0 & ((~i_10_456_1005_0 & i_10_456_1263_0 & ~i_10_456_2701_0 & ~i_10_456_4236_0 & ~i_10_456_4237_0) | (~i_10_456_1084_0 & ~i_10_456_1088_0 & ~i_10_456_2707_0 & ~i_10_456_2785_0 & ~i_10_456_4128_0 & i_10_456_4288_0))) | (~i_10_456_2704_0 & i_10_456_2919_0) | (~i_10_456_2470_0 & i_10_456_3279_0 & i_10_456_4057_0));
endmodule



// Benchmark "kernel_10_457" written by ABC on Sun Jul 19 10:29:00 2020

module kernel_10_457 ( 
    i_10_457_174_0, i_10_457_247_0, i_10_457_248_0, i_10_457_265_0,
    i_10_457_269_0, i_10_457_285_0, i_10_457_286_0, i_10_457_394_0,
    i_10_457_395_0, i_10_457_431_0, i_10_457_436_0, i_10_457_449_0,
    i_10_457_565_0, i_10_457_800_0, i_10_457_966_0, i_10_457_1006_0,
    i_10_457_1007_0, i_10_457_1084_0, i_10_457_1138_0, i_10_457_1237_0,
    i_10_457_1248_0, i_10_457_1303_0, i_10_457_1306_0, i_10_457_1308_0,
    i_10_457_1309_0, i_10_457_1310_0, i_10_457_1366_0, i_10_457_1435_0,
    i_10_457_1438_0, i_10_457_1439_0, i_10_457_1556_0, i_10_457_1654_0,
    i_10_457_1655_0, i_10_457_1717_0, i_10_457_1821_0, i_10_457_1822_0,
    i_10_457_1824_0, i_10_457_1825_0, i_10_457_1826_0, i_10_457_1913_0,
    i_10_457_1996_0, i_10_457_2006_0, i_10_457_2351_0, i_10_457_2352_0,
    i_10_457_2452_0, i_10_457_2474_0, i_10_457_2608_0, i_10_457_2614_0,
    i_10_457_2618_0, i_10_457_2631_0, i_10_457_2654_0, i_10_457_2660_0,
    i_10_457_2703_0, i_10_457_2706_0, i_10_457_2707_0, i_10_457_2722_0,
    i_10_457_2725_0, i_10_457_2730_0, i_10_457_2731_0, i_10_457_2732_0,
    i_10_457_2785_0, i_10_457_2824_0, i_10_457_2825_0, i_10_457_2830_0,
    i_10_457_2885_0, i_10_457_2920_0, i_10_457_2923_0, i_10_457_2924_0,
    i_10_457_3093_0, i_10_457_3094_0, i_10_457_3095_0, i_10_457_3156_0,
    i_10_457_3202_0, i_10_457_3277_0, i_10_457_3281_0, i_10_457_3282_0,
    i_10_457_3283_0, i_10_457_3284_0, i_10_457_3322_0, i_10_457_3473_0,
    i_10_457_3543_0, i_10_457_3587_0, i_10_457_3612_0, i_10_457_3614_0,
    i_10_457_3783_0, i_10_457_3837_0, i_10_457_3855_0, i_10_457_3857_0,
    i_10_457_3858_0, i_10_457_3986_0, i_10_457_3991_0, i_10_457_4114_0,
    i_10_457_4117_0, i_10_457_4118_0, i_10_457_4119_0, i_10_457_4120_0,
    i_10_457_4121_0, i_10_457_4566_0, i_10_457_4567_0, i_10_457_4568_0,
    o_10_457_0_0  );
  input  i_10_457_174_0, i_10_457_247_0, i_10_457_248_0, i_10_457_265_0,
    i_10_457_269_0, i_10_457_285_0, i_10_457_286_0, i_10_457_394_0,
    i_10_457_395_0, i_10_457_431_0, i_10_457_436_0, i_10_457_449_0,
    i_10_457_565_0, i_10_457_800_0, i_10_457_966_0, i_10_457_1006_0,
    i_10_457_1007_0, i_10_457_1084_0, i_10_457_1138_0, i_10_457_1237_0,
    i_10_457_1248_0, i_10_457_1303_0, i_10_457_1306_0, i_10_457_1308_0,
    i_10_457_1309_0, i_10_457_1310_0, i_10_457_1366_0, i_10_457_1435_0,
    i_10_457_1438_0, i_10_457_1439_0, i_10_457_1556_0, i_10_457_1654_0,
    i_10_457_1655_0, i_10_457_1717_0, i_10_457_1821_0, i_10_457_1822_0,
    i_10_457_1824_0, i_10_457_1825_0, i_10_457_1826_0, i_10_457_1913_0,
    i_10_457_1996_0, i_10_457_2006_0, i_10_457_2351_0, i_10_457_2352_0,
    i_10_457_2452_0, i_10_457_2474_0, i_10_457_2608_0, i_10_457_2614_0,
    i_10_457_2618_0, i_10_457_2631_0, i_10_457_2654_0, i_10_457_2660_0,
    i_10_457_2703_0, i_10_457_2706_0, i_10_457_2707_0, i_10_457_2722_0,
    i_10_457_2725_0, i_10_457_2730_0, i_10_457_2731_0, i_10_457_2732_0,
    i_10_457_2785_0, i_10_457_2824_0, i_10_457_2825_0, i_10_457_2830_0,
    i_10_457_2885_0, i_10_457_2920_0, i_10_457_2923_0, i_10_457_2924_0,
    i_10_457_3093_0, i_10_457_3094_0, i_10_457_3095_0, i_10_457_3156_0,
    i_10_457_3202_0, i_10_457_3277_0, i_10_457_3281_0, i_10_457_3282_0,
    i_10_457_3283_0, i_10_457_3284_0, i_10_457_3322_0, i_10_457_3473_0,
    i_10_457_3543_0, i_10_457_3587_0, i_10_457_3612_0, i_10_457_3614_0,
    i_10_457_3783_0, i_10_457_3837_0, i_10_457_3855_0, i_10_457_3857_0,
    i_10_457_3858_0, i_10_457_3986_0, i_10_457_3991_0, i_10_457_4114_0,
    i_10_457_4117_0, i_10_457_4118_0, i_10_457_4119_0, i_10_457_4120_0,
    i_10_457_4121_0, i_10_457_4566_0, i_10_457_4567_0, i_10_457_4568_0;
  output o_10_457_0_0;
  assign o_10_457_0_0 = ~((i_10_457_248_0 & ((~i_10_457_1084_0 & ~i_10_457_3473_0 & ~i_10_457_3855_0) | (i_10_457_436_0 & i_10_457_3857_0))) | (~i_10_457_3855_0 & ((~i_10_457_4114_0 & ((~i_10_457_966_0 & ((~i_10_457_394_0 & ~i_10_457_1309_0 & i_10_457_1821_0 & i_10_457_1822_0 & ~i_10_457_3587_0) | (~i_10_457_1306_0 & ~i_10_457_1439_0 & ~i_10_457_2920_0 & ~i_10_457_3202_0 & ~i_10_457_3543_0 & ~i_10_457_3858_0 & ~i_10_457_3986_0))) | (~i_10_457_1306_0 & i_10_457_2725_0 & ~i_10_457_3284_0 & ~i_10_457_3473_0 & ~i_10_457_3837_0))) | (~i_10_457_1306_0 & ((~i_10_457_1310_0 & ~i_10_457_1438_0 & ~i_10_457_1913_0 & ~i_10_457_3837_0) | (i_10_457_2920_0 & i_10_457_4118_0))) | (i_10_457_286_0 & ~i_10_457_1006_0 & i_10_457_1825_0 & i_10_457_3282_0) | (i_10_457_1309_0 & i_10_457_1821_0 & ~i_10_457_3093_0 & ~i_10_457_3281_0 & ~i_10_457_3282_0 & ~i_10_457_3543_0 & ~i_10_457_3587_0 & ~i_10_457_3614_0) | (i_10_457_1310_0 & ~i_10_457_2730_0 & i_10_457_2731_0 & ~i_10_457_3473_0 & i_10_457_3857_0) | (~i_10_457_2474_0 & ~i_10_457_3857_0 & ~i_10_457_3986_0 & i_10_457_4118_0))) | (~i_10_457_1007_0 & ((~i_10_457_1556_0 & ~i_10_457_1913_0 & ~i_10_457_2006_0 & i_10_457_2351_0 & ~i_10_457_2660_0 & ~i_10_457_2885_0 & ~i_10_457_3614_0 & ~i_10_457_3783_0) | (~i_10_457_1006_0 & ~i_10_457_1306_0 & i_10_457_4567_0))) | (~i_10_457_1821_0 & ((~i_10_457_1237_0 & ~i_10_457_3783_0 & ((~i_10_457_1439_0 & ~i_10_457_2722_0 & ~i_10_457_2785_0 & ~i_10_457_3543_0 & ~i_10_457_3857_0 & ~i_10_457_3986_0 & ~i_10_457_4114_0) | (~i_10_457_2351_0 & i_10_457_3855_0 & i_10_457_4117_0))) | (~i_10_457_394_0 & i_10_457_1237_0 & i_10_457_1825_0 & ~i_10_457_2452_0 & ~i_10_457_3284_0 & ~i_10_457_3857_0) | (~i_10_457_1439_0 & ~i_10_457_3986_0 & i_10_457_4121_0))) | (~i_10_457_1306_0 & ((~i_10_457_1439_0 & i_10_457_1825_0 & ~i_10_457_2722_0 & ~i_10_457_3543_0 & ~i_10_457_3783_0 & ~i_10_457_3858_0) | (~i_10_457_394_0 & ~i_10_457_1435_0 & ~i_10_457_1913_0 & ~i_10_457_2703_0 & ~i_10_457_3202_0 & i_10_457_3858_0 & ~i_10_457_3986_0))) | (~i_10_457_3543_0 & ((~i_10_457_394_0 & ~i_10_457_2474_0 & ((~i_10_457_1435_0 & i_10_457_2923_0 & ~i_10_457_3095_0) | (i_10_457_1824_0 & ~i_10_457_2660_0 & i_10_457_3202_0 & ~i_10_457_3282_0))) | (~i_10_457_1006_0 & ((i_10_457_285_0 & ~i_10_457_395_0 & i_10_457_431_0 & ~i_10_457_3093_0) | (~i_10_457_269_0 & ~i_10_457_565_0 & i_10_457_1825_0 & ~i_10_457_2618_0 & ~i_10_457_3282_0 & ~i_10_457_3612_0 & ~i_10_457_3857_0 & ~i_10_457_3986_0))) | (~i_10_457_431_0 & ~i_10_457_1439_0 & ~i_10_457_2722_0 & i_10_457_2731_0 & ~i_10_457_3093_0))) | (~i_10_457_3473_0 & ((~i_10_457_565_0 & ~i_10_457_3837_0 & ((~i_10_457_1913_0 & i_10_457_2732_0) | (i_10_457_449_0 & ~i_10_457_3095_0 & ~i_10_457_3202_0))) | (~i_10_457_174_0 & ~i_10_457_1006_0 & ~i_10_457_2731_0 & i_10_457_4120_0))) | (i_10_457_1654_0 & ((~i_10_457_2618_0 & i_10_457_2703_0) | (i_10_457_2631_0 & ~i_10_457_3283_0 & ~i_10_457_3857_0))) | (i_10_457_4117_0 & ((~i_10_457_1913_0 & ((~i_10_457_1309_0 & ~i_10_457_2618_0) | (~i_10_457_2352_0 & ~i_10_457_2474_0 & ~i_10_457_3277_0 & ~i_10_457_3783_0))) | (i_10_457_1655_0 & ~i_10_457_2614_0 & ~i_10_457_2618_0) | (i_10_457_2631_0 & ~i_10_457_3612_0) | (~i_10_457_2830_0 & ~i_10_457_3281_0 & ~i_10_457_3587_0 & i_10_457_4118_0))) | (i_10_457_2352_0 & ((~i_10_457_3282_0 & ~i_10_457_3612_0 & ~i_10_457_1439_0 & i_10_457_2706_0) | (i_10_457_1822_0 & i_10_457_2631_0 & ~i_10_457_2722_0 & ~i_10_457_3857_0))) | (~i_10_457_1309_0 & ((i_10_457_2920_0 & (i_10_457_4118_0 | (i_10_457_2722_0 & ~i_10_457_3614_0))) | (~i_10_457_1310_0 & ~i_10_457_1438_0 & ~i_10_457_2920_0 & i_10_457_3277_0 & ~i_10_457_3612_0 & ~i_10_457_3986_0))) | (~i_10_457_2722_0 & i_10_457_2830_0 & ~i_10_457_3612_0 & i_10_457_4114_0) | (i_10_457_247_0 & ~i_10_457_4114_0) | (~i_10_457_1556_0 & ~i_10_457_3587_0 & i_10_457_4568_0));
endmodule



// Benchmark "kernel_10_458" written by ABC on Sun Jul 19 10:29:01 2020

module kernel_10_458 ( 
    i_10_458_204_0, i_10_458_273_0, i_10_458_275_0, i_10_458_279_0,
    i_10_458_343_0, i_10_458_366_0, i_10_458_371_0, i_10_458_385_0,
    i_10_458_406_0, i_10_458_459_0, i_10_458_460_0, i_10_458_496_0,
    i_10_458_500_0, i_10_458_696_0, i_10_458_699_0, i_10_458_731_0,
    i_10_458_818_0, i_10_458_903_0, i_10_458_904_0, i_10_458_906_0,
    i_10_458_930_0, i_10_458_1030_0, i_10_458_1113_0, i_10_458_1166_0,
    i_10_458_1193_0, i_10_458_1221_0, i_10_458_1277_0, i_10_458_1282_0,
    i_10_458_1283_0, i_10_458_1305_0, i_10_458_1306_0, i_10_458_1360_0,
    i_10_458_1361_0, i_10_458_1365_0, i_10_458_1366_0, i_10_458_1371_0,
    i_10_458_1488_0, i_10_458_1548_0, i_10_458_1551_0, i_10_458_1641_0,
    i_10_458_1743_0, i_10_458_1909_0, i_10_458_1914_0, i_10_458_1933_0,
    i_10_458_1979_0, i_10_458_2154_0, i_10_458_2271_0, i_10_458_2272_0,
    i_10_458_2354_0, i_10_458_2376_0, i_10_458_2381_0, i_10_458_2448_0,
    i_10_458_2505_0, i_10_458_2625_0, i_10_458_2703_0, i_10_458_2707_0,
    i_10_458_2727_0, i_10_458_2730_0, i_10_458_2854_0, i_10_458_2857_0,
    i_10_458_2917_0, i_10_458_2941_0, i_10_458_2952_0, i_10_458_2955_0,
    i_10_458_3099_0, i_10_458_3100_0, i_10_458_3103_0, i_10_458_3190_0,
    i_10_458_3208_0, i_10_458_3209_0, i_10_458_3233_0, i_10_458_3236_0,
    i_10_458_3334_0, i_10_458_3362_0, i_10_458_3540_0, i_10_458_3541_0,
    i_10_458_3649_0, i_10_458_3666_0, i_10_458_3722_0, i_10_458_3837_0,
    i_10_458_3852_0, i_10_458_3860_0, i_10_458_3885_0, i_10_458_3919_0,
    i_10_458_4182_0, i_10_458_4186_0, i_10_458_4273_0, i_10_458_4359_0,
    i_10_458_4361_0, i_10_458_4369_0, i_10_458_4381_0, i_10_458_4428_0,
    i_10_458_4429_0, i_10_458_4430_0, i_10_458_4462_0, i_10_458_4523_0,
    i_10_458_4574_0, i_10_458_4590_0, i_10_458_4591_0, i_10_458_4592_0,
    o_10_458_0_0  );
  input  i_10_458_204_0, i_10_458_273_0, i_10_458_275_0, i_10_458_279_0,
    i_10_458_343_0, i_10_458_366_0, i_10_458_371_0, i_10_458_385_0,
    i_10_458_406_0, i_10_458_459_0, i_10_458_460_0, i_10_458_496_0,
    i_10_458_500_0, i_10_458_696_0, i_10_458_699_0, i_10_458_731_0,
    i_10_458_818_0, i_10_458_903_0, i_10_458_904_0, i_10_458_906_0,
    i_10_458_930_0, i_10_458_1030_0, i_10_458_1113_0, i_10_458_1166_0,
    i_10_458_1193_0, i_10_458_1221_0, i_10_458_1277_0, i_10_458_1282_0,
    i_10_458_1283_0, i_10_458_1305_0, i_10_458_1306_0, i_10_458_1360_0,
    i_10_458_1361_0, i_10_458_1365_0, i_10_458_1366_0, i_10_458_1371_0,
    i_10_458_1488_0, i_10_458_1548_0, i_10_458_1551_0, i_10_458_1641_0,
    i_10_458_1743_0, i_10_458_1909_0, i_10_458_1914_0, i_10_458_1933_0,
    i_10_458_1979_0, i_10_458_2154_0, i_10_458_2271_0, i_10_458_2272_0,
    i_10_458_2354_0, i_10_458_2376_0, i_10_458_2381_0, i_10_458_2448_0,
    i_10_458_2505_0, i_10_458_2625_0, i_10_458_2703_0, i_10_458_2707_0,
    i_10_458_2727_0, i_10_458_2730_0, i_10_458_2854_0, i_10_458_2857_0,
    i_10_458_2917_0, i_10_458_2941_0, i_10_458_2952_0, i_10_458_2955_0,
    i_10_458_3099_0, i_10_458_3100_0, i_10_458_3103_0, i_10_458_3190_0,
    i_10_458_3208_0, i_10_458_3209_0, i_10_458_3233_0, i_10_458_3236_0,
    i_10_458_3334_0, i_10_458_3362_0, i_10_458_3540_0, i_10_458_3541_0,
    i_10_458_3649_0, i_10_458_3666_0, i_10_458_3722_0, i_10_458_3837_0,
    i_10_458_3852_0, i_10_458_3860_0, i_10_458_3885_0, i_10_458_3919_0,
    i_10_458_4182_0, i_10_458_4186_0, i_10_458_4273_0, i_10_458_4359_0,
    i_10_458_4361_0, i_10_458_4369_0, i_10_458_4381_0, i_10_458_4428_0,
    i_10_458_4429_0, i_10_458_4430_0, i_10_458_4462_0, i_10_458_4523_0,
    i_10_458_4574_0, i_10_458_4590_0, i_10_458_4591_0, i_10_458_4592_0;
  output o_10_458_0_0;
  assign o_10_458_0_0 = 0;
endmodule



// Benchmark "kernel_10_459" written by ABC on Sun Jul 19 10:29:02 2020

module kernel_10_459 ( 
    i_10_459_172_0, i_10_459_173_0, i_10_459_175_0, i_10_459_244_0,
    i_10_459_286_0, i_10_459_287_0, i_10_459_316_0, i_10_459_317_0,
    i_10_459_329_0, i_10_459_406_0, i_10_459_407_0, i_10_459_461_0,
    i_10_459_515_0, i_10_459_694_0, i_10_459_695_0, i_10_459_748_0,
    i_10_459_958_0, i_10_459_1028_0, i_10_459_1081_0, i_10_459_1234_0,
    i_10_459_1235_0, i_10_459_1237_0, i_10_459_1238_0, i_10_459_1244_0,
    i_10_459_1249_0, i_10_459_1265_0, i_10_459_1306_0, i_10_459_1343_0,
    i_10_459_1541_0, i_10_459_1549_0, i_10_459_1550_0, i_10_459_1576_0,
    i_10_459_1819_0, i_10_459_2018_0, i_10_459_2027_0, i_10_459_2080_0,
    i_10_459_2201_0, i_10_459_2305_0, i_10_459_2306_0, i_10_459_2350_0,
    i_10_459_2351_0, i_10_459_2357_0, i_10_459_2361_0, i_10_459_2431_0,
    i_10_459_2432_0, i_10_459_2452_0, i_10_459_2466_0, i_10_459_2471_0,
    i_10_459_2601_0, i_10_459_2629_0, i_10_459_2630_0, i_10_459_2633_0,
    i_10_459_2661_0, i_10_459_2662_0, i_10_459_2710_0, i_10_459_2730_0,
    i_10_459_2731_0, i_10_459_2783_0, i_10_459_2786_0, i_10_459_2818_0,
    i_10_459_2819_0, i_10_459_2829_0, i_10_459_2884_0, i_10_459_2885_0,
    i_10_459_2917_0, i_10_459_2918_0, i_10_459_2953_0, i_10_459_2980_0,
    i_10_459_2981_0, i_10_459_3042_0, i_10_459_3154_0, i_10_459_3323_0,
    i_10_459_3385_0, i_10_459_3388_0, i_10_459_3389_0, i_10_459_3407_0,
    i_10_459_3526_0, i_10_459_3556_0, i_10_459_3583_0, i_10_459_3586_0,
    i_10_459_3613_0, i_10_459_3614_0, i_10_459_3843_0, i_10_459_3847_0,
    i_10_459_3848_0, i_10_459_3852_0, i_10_459_3853_0, i_10_459_3858_0,
    i_10_459_3888_0, i_10_459_3889_0, i_10_459_3890_0, i_10_459_3908_0,
    i_10_459_3980_0, i_10_459_3981_0, i_10_459_4120_0, i_10_459_4127_0,
    i_10_459_4271_0, i_10_459_4277_0, i_10_459_4285_0, i_10_459_4564_0,
    o_10_459_0_0  );
  input  i_10_459_172_0, i_10_459_173_0, i_10_459_175_0, i_10_459_244_0,
    i_10_459_286_0, i_10_459_287_0, i_10_459_316_0, i_10_459_317_0,
    i_10_459_329_0, i_10_459_406_0, i_10_459_407_0, i_10_459_461_0,
    i_10_459_515_0, i_10_459_694_0, i_10_459_695_0, i_10_459_748_0,
    i_10_459_958_0, i_10_459_1028_0, i_10_459_1081_0, i_10_459_1234_0,
    i_10_459_1235_0, i_10_459_1237_0, i_10_459_1238_0, i_10_459_1244_0,
    i_10_459_1249_0, i_10_459_1265_0, i_10_459_1306_0, i_10_459_1343_0,
    i_10_459_1541_0, i_10_459_1549_0, i_10_459_1550_0, i_10_459_1576_0,
    i_10_459_1819_0, i_10_459_2018_0, i_10_459_2027_0, i_10_459_2080_0,
    i_10_459_2201_0, i_10_459_2305_0, i_10_459_2306_0, i_10_459_2350_0,
    i_10_459_2351_0, i_10_459_2357_0, i_10_459_2361_0, i_10_459_2431_0,
    i_10_459_2432_0, i_10_459_2452_0, i_10_459_2466_0, i_10_459_2471_0,
    i_10_459_2601_0, i_10_459_2629_0, i_10_459_2630_0, i_10_459_2633_0,
    i_10_459_2661_0, i_10_459_2662_0, i_10_459_2710_0, i_10_459_2730_0,
    i_10_459_2731_0, i_10_459_2783_0, i_10_459_2786_0, i_10_459_2818_0,
    i_10_459_2819_0, i_10_459_2829_0, i_10_459_2884_0, i_10_459_2885_0,
    i_10_459_2917_0, i_10_459_2918_0, i_10_459_2953_0, i_10_459_2980_0,
    i_10_459_2981_0, i_10_459_3042_0, i_10_459_3154_0, i_10_459_3323_0,
    i_10_459_3385_0, i_10_459_3388_0, i_10_459_3389_0, i_10_459_3407_0,
    i_10_459_3526_0, i_10_459_3556_0, i_10_459_3583_0, i_10_459_3586_0,
    i_10_459_3613_0, i_10_459_3614_0, i_10_459_3843_0, i_10_459_3847_0,
    i_10_459_3848_0, i_10_459_3852_0, i_10_459_3853_0, i_10_459_3858_0,
    i_10_459_3888_0, i_10_459_3889_0, i_10_459_3890_0, i_10_459_3908_0,
    i_10_459_3980_0, i_10_459_3981_0, i_10_459_4120_0, i_10_459_4127_0,
    i_10_459_4271_0, i_10_459_4277_0, i_10_459_4285_0, i_10_459_4564_0;
  output o_10_459_0_0;
  assign o_10_459_0_0 = ~((~i_10_459_4277_0 & ((~i_10_459_329_0 & ((~i_10_459_244_0 & ~i_10_459_695_0 & ~i_10_459_1550_0 & ~i_10_459_2306_0 & ~i_10_459_3889_0) | (~i_10_459_175_0 & ~i_10_459_316_0 & ~i_10_459_2357_0 & ~i_10_459_2662_0 & ~i_10_459_3389_0 & ~i_10_459_3614_0 & ~i_10_459_3853_0 & ~i_10_459_4285_0 & ~i_10_459_4564_0))) | (~i_10_459_317_0 & i_10_459_3583_0) | (~i_10_459_748_0 & ~i_10_459_2884_0 & ~i_10_459_2980_0 & ~i_10_459_3407_0 & ~i_10_459_3847_0 & ~i_10_459_4120_0))) | (~i_10_459_316_0 & ((i_10_459_1819_0 & ~i_10_459_2630_0) | (~i_10_459_2350_0 & i_10_459_3389_0 & ~i_10_459_3980_0 & ~i_10_459_4564_0))) | (~i_10_459_515_0 & ((i_10_459_1819_0 & i_10_459_3389_0) | (~i_10_459_695_0 & ~i_10_459_1028_0 & ~i_10_459_1244_0 & ~i_10_459_2305_0 & ~i_10_459_2601_0 & ~i_10_459_2884_0 & ~i_10_459_3858_0 & ~i_10_459_3908_0))) | (~i_10_459_3981_0 & ((~i_10_459_694_0 & ~i_10_459_3847_0 & ((~i_10_459_1081_0 & ~i_10_459_1265_0 & ~i_10_459_1550_0 & ~i_10_459_2306_0 & ~i_10_459_3890_0) | (~i_10_459_1576_0 & ~i_10_459_2818_0 & ~i_10_459_2819_0 & ~i_10_459_2884_0 & ~i_10_459_3613_0 & ~i_10_459_4271_0))) | (~i_10_459_2305_0 & ~i_10_459_2819_0 & ~i_10_459_2980_0 & ~i_10_459_3852_0 & i_10_459_3853_0 & ~i_10_459_4285_0))) | (~i_10_459_1081_0 & ((i_10_459_1819_0 & ~i_10_459_2201_0 & ~i_10_459_2361_0 & ~i_10_459_2710_0 & ~i_10_459_3980_0) | (~i_10_459_1549_0 & ~i_10_459_2306_0 & ~i_10_459_4285_0 & i_10_459_4564_0))) | (~i_10_459_2818_0 & (i_10_459_286_0 | (~i_10_459_1550_0 & ((i_10_459_1237_0 & ~i_10_459_1244_0 & ~i_10_459_2027_0 & ~i_10_459_2980_0) | (~i_10_459_748_0 & ~i_10_459_1541_0 & ~i_10_459_2350_0 & ~i_10_459_2819_0 & ~i_10_459_3388_0 & ~i_10_459_3908_0))))) | (~i_10_459_2018_0 & ((~i_10_459_1549_0 & ~i_10_459_2306_0 & ~i_10_459_2351_0 & ~i_10_459_2980_0) | (~i_10_459_1234_0 & ~i_10_459_2731_0 & i_10_459_3388_0 & i_10_459_3847_0))) | (~i_10_459_4285_0 & ((~i_10_459_2629_0 & i_10_459_2917_0) | (~i_10_459_1306_0 & ~i_10_459_2201_0 & ~i_10_459_2351_0 & ~i_10_459_2361_0 & ~i_10_459_2601_0 & ~i_10_459_2633_0 & ~i_10_459_3389_0 & ~i_10_459_4564_0))) | (i_10_459_1819_0 & i_10_459_2471_0 & i_10_459_3583_0) | (~i_10_459_2630_0 & i_10_459_3407_0 & i_10_459_3853_0 & ~i_10_459_3980_0) | (~i_10_459_287_0 & ~i_10_459_1028_0 & ~i_10_459_1265_0 & ~i_10_459_1343_0 & ~i_10_459_3583_0 & ~i_10_459_3843_0 & ~i_10_459_3853_0 & ~i_10_459_3888_0 & ~i_10_459_3890_0 & ~i_10_459_4271_0) | (i_10_459_3847_0 & i_10_459_4120_0 & i_10_459_4564_0));
endmodule



// Benchmark "kernel_10_460" written by ABC on Sun Jul 19 10:29:03 2020

module kernel_10_460 ( 
    i_10_460_125_0, i_10_460_268_0, i_10_460_269_0, i_10_460_283_0,
    i_10_460_286_0, i_10_460_319_0, i_10_460_320_0, i_10_460_392_0,
    i_10_460_395_0, i_10_460_441_0, i_10_460_466_0, i_10_460_539_0,
    i_10_460_581_0, i_10_460_754_0, i_10_460_795_0, i_10_460_953_0,
    i_10_460_1004_0, i_10_460_1006_0, i_10_460_1007_0, i_10_460_1205_0,
    i_10_460_1308_0, i_10_460_1312_0, i_10_460_1345_0, i_10_460_1552_0,
    i_10_460_1577_0, i_10_460_1616_0, i_10_460_1618_0, i_10_460_1619_0,
    i_10_460_1648_0, i_10_460_1650_0, i_10_460_1651_0, i_10_460_1686_0,
    i_10_460_1697_0, i_10_460_1824_0, i_10_460_2158_0, i_10_460_2159_0,
    i_10_460_2310_0, i_10_460_2311_0, i_10_460_2312_0, i_10_460_2336_0,
    i_10_460_2339_0, i_10_460_2354_0, i_10_460_2357_0, i_10_460_2405_0,
    i_10_460_2407_0, i_10_460_2408_0, i_10_460_2410_0, i_10_460_2447_0,
    i_10_460_2455_0, i_10_460_2463_0, i_10_460_2519_0, i_10_460_2536_0,
    i_10_460_2618_0, i_10_460_2629_0, i_10_460_2632_0, i_10_460_2633_0,
    i_10_460_2635_0, i_10_460_2636_0, i_10_460_2705_0, i_10_460_2734_0,
    i_10_460_2788_0, i_10_460_2826_0, i_10_460_2884_0, i_10_460_2885_0,
    i_10_460_2987_0, i_10_460_3058_0, i_10_460_3070_0, i_10_460_3199_0,
    i_10_460_3200_0, i_10_460_3329_0, i_10_460_3365_0, i_10_460_3387_0,
    i_10_460_3391_0, i_10_460_3392_0, i_10_460_3437_0, i_10_460_3587_0,
    i_10_460_3623_0, i_10_460_3645_0, i_10_460_3650_0, i_10_460_3653_0,
    i_10_460_3707_0, i_10_460_3733_0, i_10_460_3734_0, i_10_460_3781_0,
    i_10_460_3838_0, i_10_460_3839_0, i_10_460_3884_0, i_10_460_3986_0,
    i_10_460_4058_0, i_10_460_4094_0, i_10_460_4115_0, i_10_460_4120_0,
    i_10_460_4184_0, i_10_460_4266_0, i_10_460_4268_0, i_10_460_4274_0,
    i_10_460_4382_0, i_10_460_4460_0, i_10_460_4534_0, i_10_460_4567_0,
    o_10_460_0_0  );
  input  i_10_460_125_0, i_10_460_268_0, i_10_460_269_0, i_10_460_283_0,
    i_10_460_286_0, i_10_460_319_0, i_10_460_320_0, i_10_460_392_0,
    i_10_460_395_0, i_10_460_441_0, i_10_460_466_0, i_10_460_539_0,
    i_10_460_581_0, i_10_460_754_0, i_10_460_795_0, i_10_460_953_0,
    i_10_460_1004_0, i_10_460_1006_0, i_10_460_1007_0, i_10_460_1205_0,
    i_10_460_1308_0, i_10_460_1312_0, i_10_460_1345_0, i_10_460_1552_0,
    i_10_460_1577_0, i_10_460_1616_0, i_10_460_1618_0, i_10_460_1619_0,
    i_10_460_1648_0, i_10_460_1650_0, i_10_460_1651_0, i_10_460_1686_0,
    i_10_460_1697_0, i_10_460_1824_0, i_10_460_2158_0, i_10_460_2159_0,
    i_10_460_2310_0, i_10_460_2311_0, i_10_460_2312_0, i_10_460_2336_0,
    i_10_460_2339_0, i_10_460_2354_0, i_10_460_2357_0, i_10_460_2405_0,
    i_10_460_2407_0, i_10_460_2408_0, i_10_460_2410_0, i_10_460_2447_0,
    i_10_460_2455_0, i_10_460_2463_0, i_10_460_2519_0, i_10_460_2536_0,
    i_10_460_2618_0, i_10_460_2629_0, i_10_460_2632_0, i_10_460_2633_0,
    i_10_460_2635_0, i_10_460_2636_0, i_10_460_2705_0, i_10_460_2734_0,
    i_10_460_2788_0, i_10_460_2826_0, i_10_460_2884_0, i_10_460_2885_0,
    i_10_460_2987_0, i_10_460_3058_0, i_10_460_3070_0, i_10_460_3199_0,
    i_10_460_3200_0, i_10_460_3329_0, i_10_460_3365_0, i_10_460_3387_0,
    i_10_460_3391_0, i_10_460_3392_0, i_10_460_3437_0, i_10_460_3587_0,
    i_10_460_3623_0, i_10_460_3645_0, i_10_460_3650_0, i_10_460_3653_0,
    i_10_460_3707_0, i_10_460_3733_0, i_10_460_3734_0, i_10_460_3781_0,
    i_10_460_3838_0, i_10_460_3839_0, i_10_460_3884_0, i_10_460_3986_0,
    i_10_460_4058_0, i_10_460_4094_0, i_10_460_4115_0, i_10_460_4120_0,
    i_10_460_4184_0, i_10_460_4266_0, i_10_460_4268_0, i_10_460_4274_0,
    i_10_460_4382_0, i_10_460_4460_0, i_10_460_4534_0, i_10_460_4567_0;
  output o_10_460_0_0;
  assign o_10_460_0_0 = ~((~i_10_460_269_0 & ((~i_10_460_1006_0 & ~i_10_460_1007_0 & ~i_10_460_2310_0 & ~i_10_460_3645_0 & ~i_10_460_3986_0 & ~i_10_460_4058_0) | (~i_10_460_125_0 & ~i_10_460_2357_0 & ~i_10_460_2408_0 & ~i_10_460_4120_0 & ~i_10_460_4268_0 & ~i_10_460_4567_0))) | (i_10_460_286_0 & ((i_10_460_1345_0 & ~i_10_460_1552_0 & ~i_10_460_2310_0 & ~i_10_460_2407_0 & i_10_460_3387_0) | (~i_10_460_392_0 & ~i_10_460_1577_0 & ~i_10_460_1618_0 & ~i_10_460_1824_0 & ~i_10_460_2312_0 & ~i_10_460_3392_0 & ~i_10_460_3645_0 & ~i_10_460_4120_0 & ~i_10_460_4567_0))) | (~i_10_460_395_0 & ((~i_10_460_283_0 & ~i_10_460_1618_0 & ~i_10_460_2339_0 & ~i_10_460_2407_0) | (~i_10_460_2408_0 & ~i_10_460_2705_0 & ~i_10_460_3437_0))) | (~i_10_460_1618_0 & ((~i_10_460_1619_0 & ~i_10_460_2357_0 & ((~i_10_460_320_0 & ~i_10_460_1650_0 & ~i_10_460_3838_0 & ~i_10_460_4058_0 & ~i_10_460_4266_0) | (~i_10_460_2311_0 & ~i_10_460_2629_0 & ~i_10_460_2826_0 & ~i_10_460_2987_0 & ~i_10_460_4120_0 & ~i_10_460_4274_0))) | (~i_10_460_392_0 & ~i_10_460_2310_0 & ~i_10_460_2339_0 & ~i_10_460_3392_0 & ~i_10_460_3838_0 & ~i_10_460_3986_0))) | (~i_10_460_2312_0 & ((~i_10_460_466_0 & ~i_10_460_1616_0 & ~i_10_460_2788_0 & ~i_10_460_2826_0 & i_10_460_4268_0) | (~i_10_460_1824_0 & i_10_460_2633_0 & ~i_10_460_3437_0 & ~i_10_460_3587_0 & ~i_10_460_4268_0))) | (i_10_460_2407_0 & ((i_10_460_441_0 & i_10_460_3392_0) | (i_10_460_2312_0 & ~i_10_460_2336_0 & ~i_10_460_2618_0 & ~i_10_460_2987_0 & ~i_10_460_3986_0))) | (~i_10_460_2705_0 & ((~i_10_460_268_0 & ~i_10_460_1006_0 & ~i_10_460_2357_0 & ~i_10_460_2618_0) | (~i_10_460_3645_0 & ~i_10_460_4058_0 & ~i_10_460_4567_0))) | (~i_10_460_268_0 & ((i_10_460_1824_0 & ~i_10_460_2407_0 & ~i_10_460_2408_0) | (~i_10_460_1686_0 & i_10_460_3391_0 & ~i_10_460_3437_0 & ~i_10_460_4268_0))) | (~i_10_460_2788_0 & ~i_10_460_3587_0 & ~i_10_460_4058_0 & ~i_10_460_4274_0));
endmodule



// Benchmark "kernel_10_461" written by ABC on Sun Jul 19 10:29:04 2020

module kernel_10_461 ( 
    i_10_461_39_0, i_10_461_149_0, i_10_461_154_0, i_10_461_243_0,
    i_10_461_247_0, i_10_461_263_0, i_10_461_290_0, i_10_461_315_0,
    i_10_461_317_0, i_10_461_318_0, i_10_461_319_0, i_10_461_321_0,
    i_10_461_387_0, i_10_461_409_0, i_10_461_423_0, i_10_461_445_0,
    i_10_461_460_0, i_10_461_462_0, i_10_461_500_0, i_10_461_503_0,
    i_10_461_521_0, i_10_461_639_0, i_10_461_671_0, i_10_461_752_0,
    i_10_461_891_0, i_10_461_1080_0, i_10_461_1237_0, i_10_461_1241_0,
    i_10_461_1270_0, i_10_461_1297_0, i_10_461_1345_0, i_10_461_1432_0,
    i_10_461_1433_0, i_10_461_1442_0, i_10_461_1535_0, i_10_461_1541_0,
    i_10_461_1544_0, i_10_461_1546_0, i_10_461_1596_0, i_10_461_1634_0,
    i_10_461_1643_0, i_10_461_1651_0, i_10_461_1654_0, i_10_461_1684_0,
    i_10_461_1690_0, i_10_461_1810_0, i_10_461_1821_0, i_10_461_1918_0,
    i_10_461_1989_0, i_10_461_2000_0, i_10_461_2003_0, i_10_461_2017_0,
    i_10_461_2018_0, i_10_461_2029_0, i_10_461_2030_0, i_10_461_2033_0,
    i_10_461_2107_0, i_10_461_2108_0, i_10_461_2235_0, i_10_461_2262_0,
    i_10_461_2312_0, i_10_461_2345_0, i_10_461_2348_0, i_10_461_2358_0,
    i_10_461_2361_0, i_10_461_2362_0, i_10_461_2384_0, i_10_461_2448_0,
    i_10_461_2449_0, i_10_461_2454_0, i_10_461_2465_0, i_10_461_2566_0,
    i_10_461_2567_0, i_10_461_2601_0, i_10_461_2635_0, i_10_461_2705_0,
    i_10_461_2785_0, i_10_461_2820_0, i_10_461_2822_0, i_10_461_2915_0,
    i_10_461_3044_0, i_10_461_3070_0, i_10_461_3165_0, i_10_461_3279_0,
    i_10_461_3317_0, i_10_461_3320_0, i_10_461_3335_0, i_10_461_3430_0,
    i_10_461_3467_0, i_10_461_3494_0, i_10_461_3557_0, i_10_461_3560_0,
    i_10_461_3794_0, i_10_461_3841_0, i_10_461_3881_0, i_10_461_3914_0,
    i_10_461_4118_0, i_10_461_4271_0, i_10_461_4274_0, i_10_461_4583_0,
    o_10_461_0_0  );
  input  i_10_461_39_0, i_10_461_149_0, i_10_461_154_0, i_10_461_243_0,
    i_10_461_247_0, i_10_461_263_0, i_10_461_290_0, i_10_461_315_0,
    i_10_461_317_0, i_10_461_318_0, i_10_461_319_0, i_10_461_321_0,
    i_10_461_387_0, i_10_461_409_0, i_10_461_423_0, i_10_461_445_0,
    i_10_461_460_0, i_10_461_462_0, i_10_461_500_0, i_10_461_503_0,
    i_10_461_521_0, i_10_461_639_0, i_10_461_671_0, i_10_461_752_0,
    i_10_461_891_0, i_10_461_1080_0, i_10_461_1237_0, i_10_461_1241_0,
    i_10_461_1270_0, i_10_461_1297_0, i_10_461_1345_0, i_10_461_1432_0,
    i_10_461_1433_0, i_10_461_1442_0, i_10_461_1535_0, i_10_461_1541_0,
    i_10_461_1544_0, i_10_461_1546_0, i_10_461_1596_0, i_10_461_1634_0,
    i_10_461_1643_0, i_10_461_1651_0, i_10_461_1654_0, i_10_461_1684_0,
    i_10_461_1690_0, i_10_461_1810_0, i_10_461_1821_0, i_10_461_1918_0,
    i_10_461_1989_0, i_10_461_2000_0, i_10_461_2003_0, i_10_461_2017_0,
    i_10_461_2018_0, i_10_461_2029_0, i_10_461_2030_0, i_10_461_2033_0,
    i_10_461_2107_0, i_10_461_2108_0, i_10_461_2235_0, i_10_461_2262_0,
    i_10_461_2312_0, i_10_461_2345_0, i_10_461_2348_0, i_10_461_2358_0,
    i_10_461_2361_0, i_10_461_2362_0, i_10_461_2384_0, i_10_461_2448_0,
    i_10_461_2449_0, i_10_461_2454_0, i_10_461_2465_0, i_10_461_2566_0,
    i_10_461_2567_0, i_10_461_2601_0, i_10_461_2635_0, i_10_461_2705_0,
    i_10_461_2785_0, i_10_461_2820_0, i_10_461_2822_0, i_10_461_2915_0,
    i_10_461_3044_0, i_10_461_3070_0, i_10_461_3165_0, i_10_461_3279_0,
    i_10_461_3317_0, i_10_461_3320_0, i_10_461_3335_0, i_10_461_3430_0,
    i_10_461_3467_0, i_10_461_3494_0, i_10_461_3557_0, i_10_461_3560_0,
    i_10_461_3794_0, i_10_461_3841_0, i_10_461_3881_0, i_10_461_3914_0,
    i_10_461_4118_0, i_10_461_4271_0, i_10_461_4274_0, i_10_461_4583_0;
  output o_10_461_0_0;
  assign o_10_461_0_0 = 0;
endmodule



// Benchmark "kernel_10_462" written by ABC on Sun Jul 19 10:29:06 2020

module kernel_10_462 ( 
    i_10_462_40_0, i_10_462_83_0, i_10_462_172_0, i_10_462_282_0,
    i_10_462_289_0, i_10_462_445_0, i_10_462_460_0, i_10_462_461_0,
    i_10_462_463_0, i_10_462_464_0, i_10_462_466_0, i_10_462_504_0,
    i_10_462_715_0, i_10_462_799_0, i_10_462_892_0, i_10_462_967_0,
    i_10_462_1000_0, i_10_462_1042_0, i_10_462_1135_0, i_10_462_1233_0,
    i_10_462_1234_0, i_10_462_1235_0, i_10_462_1241_0, i_10_462_1243_0,
    i_10_462_1344_0, i_10_462_1359_0, i_10_462_1360_0, i_10_462_1361_0,
    i_10_462_1363_0, i_10_462_1364_0, i_10_462_1367_0, i_10_462_1441_0,
    i_10_462_1444_0, i_10_462_1540_0, i_10_462_1543_0, i_10_462_1549_0,
    i_10_462_1576_0, i_10_462_1577_0, i_10_462_1578_0, i_10_462_1580_0,
    i_10_462_1650_0, i_10_462_1678_0, i_10_462_1767_0, i_10_462_1818_0,
    i_10_462_1819_0, i_10_462_1823_0, i_10_462_1908_0, i_10_462_1909_0,
    i_10_462_1911_0, i_10_462_2182_0, i_10_462_2352_0, i_10_462_2357_0,
    i_10_462_2382_0, i_10_462_2455_0, i_10_462_2470_0, i_10_462_2648_0,
    i_10_462_2655_0, i_10_462_2657_0, i_10_462_2673_0, i_10_462_2709_0,
    i_10_462_2710_0, i_10_462_2718_0, i_10_462_2727_0, i_10_462_2728_0,
    i_10_462_2729_0, i_10_462_2826_0, i_10_462_2827_0, i_10_462_2829_0,
    i_10_462_2882_0, i_10_462_2917_0, i_10_462_2918_0, i_10_462_2919_0,
    i_10_462_2920_0, i_10_462_3035_0, i_10_462_3042_0, i_10_462_3231_0,
    i_10_462_3271_0, i_10_462_3321_0, i_10_462_3322_0, i_10_462_3324_0,
    i_10_462_3325_0, i_10_462_3384_0, i_10_462_3385_0, i_10_462_3389_0,
    i_10_462_3523_0, i_10_462_3550_0, i_10_462_3585_0, i_10_462_3586_0,
    i_10_462_3645_0, i_10_462_3781_0, i_10_462_3846_0, i_10_462_3848_0,
    i_10_462_3854_0, i_10_462_3979_0, i_10_462_3980_0, i_10_462_4284_0,
    i_10_462_4285_0, i_10_462_4286_0, i_10_462_4290_0, i_10_462_4565_0,
    o_10_462_0_0  );
  input  i_10_462_40_0, i_10_462_83_0, i_10_462_172_0, i_10_462_282_0,
    i_10_462_289_0, i_10_462_445_0, i_10_462_460_0, i_10_462_461_0,
    i_10_462_463_0, i_10_462_464_0, i_10_462_466_0, i_10_462_504_0,
    i_10_462_715_0, i_10_462_799_0, i_10_462_892_0, i_10_462_967_0,
    i_10_462_1000_0, i_10_462_1042_0, i_10_462_1135_0, i_10_462_1233_0,
    i_10_462_1234_0, i_10_462_1235_0, i_10_462_1241_0, i_10_462_1243_0,
    i_10_462_1344_0, i_10_462_1359_0, i_10_462_1360_0, i_10_462_1361_0,
    i_10_462_1363_0, i_10_462_1364_0, i_10_462_1367_0, i_10_462_1441_0,
    i_10_462_1444_0, i_10_462_1540_0, i_10_462_1543_0, i_10_462_1549_0,
    i_10_462_1576_0, i_10_462_1577_0, i_10_462_1578_0, i_10_462_1580_0,
    i_10_462_1650_0, i_10_462_1678_0, i_10_462_1767_0, i_10_462_1818_0,
    i_10_462_1819_0, i_10_462_1823_0, i_10_462_1908_0, i_10_462_1909_0,
    i_10_462_1911_0, i_10_462_2182_0, i_10_462_2352_0, i_10_462_2357_0,
    i_10_462_2382_0, i_10_462_2455_0, i_10_462_2470_0, i_10_462_2648_0,
    i_10_462_2655_0, i_10_462_2657_0, i_10_462_2673_0, i_10_462_2709_0,
    i_10_462_2710_0, i_10_462_2718_0, i_10_462_2727_0, i_10_462_2728_0,
    i_10_462_2729_0, i_10_462_2826_0, i_10_462_2827_0, i_10_462_2829_0,
    i_10_462_2882_0, i_10_462_2917_0, i_10_462_2918_0, i_10_462_2919_0,
    i_10_462_2920_0, i_10_462_3035_0, i_10_462_3042_0, i_10_462_3231_0,
    i_10_462_3271_0, i_10_462_3321_0, i_10_462_3322_0, i_10_462_3324_0,
    i_10_462_3325_0, i_10_462_3384_0, i_10_462_3385_0, i_10_462_3389_0,
    i_10_462_3523_0, i_10_462_3550_0, i_10_462_3585_0, i_10_462_3586_0,
    i_10_462_3645_0, i_10_462_3781_0, i_10_462_3846_0, i_10_462_3848_0,
    i_10_462_3854_0, i_10_462_3979_0, i_10_462_3980_0, i_10_462_4284_0,
    i_10_462_4285_0, i_10_462_4286_0, i_10_462_4290_0, i_10_462_4565_0;
  output o_10_462_0_0;
  assign o_10_462_0_0 = ~((~i_10_462_445_0 & ((~i_10_462_1042_0 & ~i_10_462_1233_0 & ~i_10_462_1359_0 & ~i_10_462_1360_0 & ~i_10_462_1361_0 & ~i_10_462_2455_0 & ~i_10_462_3271_0 & ~i_10_462_3523_0 & ~i_10_462_3846_0 & ~i_10_462_3848_0) | (~i_10_462_282_0 & ~i_10_462_466_0 & ~i_10_462_1241_0 & ~i_10_462_1444_0 & ~i_10_462_3550_0 & i_10_462_3980_0))) | (~i_10_462_1767_0 & ((~i_10_462_282_0 & ((~i_10_462_289_0 & ~i_10_462_461_0 & ~i_10_462_2657_0 & ~i_10_462_2728_0 & ~i_10_462_2729_0) | (~i_10_462_967_0 & ~i_10_462_1360_0 & ~i_10_462_1361_0 & ~i_10_462_1367_0 & ~i_10_462_1441_0 & ~i_10_462_2727_0 & ~i_10_462_2918_0 & ~i_10_462_3231_0))) | (~i_10_462_1359_0 & ((~i_10_462_289_0 & ~i_10_462_1233_0 & ~i_10_462_1361_0 & ~i_10_462_1367_0 & ~i_10_462_2357_0 & ~i_10_462_2470_0 & ~i_10_462_2709_0 & ~i_10_462_2882_0 & ~i_10_462_3035_0 & ~i_10_462_3231_0 & ~i_10_462_4284_0) | (~i_10_462_1042_0 & ~i_10_462_1364_0 & ~i_10_462_1444_0 & ~i_10_462_1911_0 & i_10_462_2826_0 & ~i_10_462_3980_0 & ~i_10_462_4285_0 & ~i_10_462_4286_0))) | (~i_10_462_3848_0 & ((~i_10_462_460_0 & ~i_10_462_464_0 & ~i_10_462_1363_0 & ~i_10_462_1367_0 & ~i_10_462_1444_0 & ~i_10_462_2920_0) | (~i_10_462_1235_0 & ~i_10_462_1364_0 & ~i_10_462_2826_0 & ~i_10_462_2917_0 & ~i_10_462_3384_0 & ~i_10_462_3585_0))) | (~i_10_462_461_0 & ~i_10_462_463_0 & ~i_10_462_1344_0 & ~i_10_462_2718_0 & ~i_10_462_3231_0 & ~i_10_462_3550_0 & ~i_10_462_4565_0))) | (~i_10_462_1360_0 & ((~i_10_462_1364_0 & ((~i_10_462_282_0 & ((~i_10_462_892_0 & ~i_10_462_1363_0 & ~i_10_462_1367_0 & ~i_10_462_1441_0 & ~i_10_462_2455_0 & ~i_10_462_2470_0 & ~i_10_462_2709_0 & ~i_10_462_3035_0) | (~i_10_462_2655_0 & ~i_10_462_2918_0 & i_10_462_3854_0 & ~i_10_462_4285_0 & ~i_10_462_4565_0))) | (i_10_462_445_0 & ~i_10_462_1042_0 & ~i_10_462_1235_0 & ~i_10_462_1241_0 & ~i_10_462_1361_0 & ~i_10_462_2352_0 & ~i_10_462_3042_0 & ~i_10_462_3231_0 & ~i_10_462_3385_0 & ~i_10_462_3523_0) | (~i_10_462_1344_0 & ~i_10_462_1367_0 & ~i_10_462_2673_0 & ~i_10_462_2729_0 & ~i_10_462_2826_0 & ~i_10_462_3846_0 & ~i_10_462_4286_0))) | (~i_10_462_1367_0 & ~i_10_462_3585_0 & ((~i_10_462_967_0 & ~i_10_462_1577_0 & i_10_462_1819_0 & ~i_10_462_2728_0) | (~i_10_462_1359_0 & ~i_10_462_1363_0 & ~i_10_462_1911_0 & ~i_10_462_2657_0 & ~i_10_462_3042_0 & ~i_10_462_4286_0 & ~i_10_462_4565_0))) | (i_10_462_1650_0 & ~i_10_462_2655_0 & i_10_462_3384_0 & ~i_10_462_3385_0 & ~i_10_462_3586_0))) | (~i_10_462_1359_0 & ((~i_10_462_799_0 & ((~i_10_462_1361_0 & ~i_10_462_1364_0 & i_10_462_1819_0 & ~i_10_462_2709_0 & ~i_10_462_2710_0 & ~i_10_462_2727_0 & ~i_10_462_2826_0 & ~i_10_462_3385_0) | (i_10_462_463_0 & ~i_10_462_1363_0 & ~i_10_462_1911_0 & ~i_10_462_2182_0 & ~i_10_462_2455_0 & ~i_10_462_3231_0 & ~i_10_462_3781_0 & ~i_10_462_3854_0 & ~i_10_462_4565_0))) | (~i_10_462_1361_0 & ~i_10_462_1823_0 & ~i_10_462_2718_0 & ~i_10_462_2729_0 & ~i_10_462_2827_0 & ~i_10_462_2920_0 & ~i_10_462_3585_0))) | (~i_10_462_1361_0 & ((~i_10_462_1367_0 & i_10_462_1577_0) | (~i_10_462_1241_0 & ~i_10_462_1909_0 & ~i_10_462_2728_0 & ~i_10_462_3042_0 & ~i_10_462_3231_0))) | (~i_10_462_2728_0 & ((~i_10_462_289_0 & i_10_462_3389_0 & ~i_10_462_3586_0 & i_10_462_4285_0) | (~i_10_462_1234_0 & ~i_10_462_1363_0 & ~i_10_462_3271_0 & ~i_10_462_3523_0 & ~i_10_462_3550_0 & ~i_10_462_4290_0))) | (i_10_462_3979_0 & ((i_10_462_1650_0 & i_10_462_3585_0) | (~i_10_462_1911_0 & ~i_10_462_3586_0 & i_10_462_3645_0))) | (i_10_462_2470_0 & i_10_462_3271_0 & i_10_462_3389_0 & ~i_10_462_3854_0) | (~i_10_462_1364_0 & ~i_10_462_1367_0 & ~i_10_462_1823_0 & ~i_10_462_2470_0 & ~i_10_462_2655_0 & ~i_10_462_3035_0 & ~i_10_462_3384_0 & ~i_10_462_3550_0 & ~i_10_462_3781_0 & ~i_10_462_4284_0));
endmodule



// Benchmark "kernel_10_463" written by ABC on Sun Jul 19 10:29:07 2020

module kernel_10_463 ( 
    i_10_463_243_0, i_10_463_252_0, i_10_463_263_0, i_10_463_286_0,
    i_10_463_317_0, i_10_463_319_0, i_10_463_320_0, i_10_463_395_0,
    i_10_463_512_0, i_10_463_621_0, i_10_463_687_0, i_10_463_688_0,
    i_10_463_865_0, i_10_463_1001_0, i_10_463_1003_0, i_10_463_1004_0,
    i_10_463_1058_0, i_10_463_1081_0, i_10_463_1084_0, i_10_463_1134_0,
    i_10_463_1135_0, i_10_463_1152_0, i_10_463_1153_0, i_10_463_1223_0,
    i_10_463_1237_0, i_10_463_1263_0, i_10_463_1300_0, i_10_463_1435_0,
    i_10_463_1436_0, i_10_463_1530_0, i_10_463_1535_0, i_10_463_1548_0,
    i_10_463_1551_0, i_10_463_1552_0, i_10_463_1580_0, i_10_463_1625_0,
    i_10_463_1628_0, i_10_463_1730_0, i_10_463_1733_0, i_10_463_1808_0,
    i_10_463_1810_0, i_10_463_1821_0, i_10_463_1906_0, i_10_463_1915_0,
    i_10_463_2020_0, i_10_463_2030_0, i_10_463_2033_0, i_10_463_2064_0,
    i_10_463_2111_0, i_10_463_2200_0, i_10_463_2340_0, i_10_463_2345_0,
    i_10_463_2349_0, i_10_463_2352_0, i_10_463_2353_0, i_10_463_2363_0,
    i_10_463_2380_0, i_10_463_2406_0, i_10_463_2453_0, i_10_463_2468_0,
    i_10_463_2567_0, i_10_463_2570_0, i_10_463_2703_0, i_10_463_2731_0,
    i_10_463_2732_0, i_10_463_2741_0, i_10_463_2744_0, i_10_463_2782_0,
    i_10_463_2808_0, i_10_463_2839_0, i_10_463_2840_0, i_10_463_3043_0,
    i_10_463_3047_0, i_10_463_3091_0, i_10_463_3195_0, i_10_463_3202_0,
    i_10_463_3271_0, i_10_463_3317_0, i_10_463_3320_0, i_10_463_3335_0,
    i_10_463_3353_0, i_10_463_3393_0, i_10_463_3473_0, i_10_463_3545_0,
    i_10_463_3560_0, i_10_463_3612_0, i_10_463_3663_0, i_10_463_3789_0,
    i_10_463_3842_0, i_10_463_3911_0, i_10_463_3942_0, i_10_463_3946_0,
    i_10_463_3999_0, i_10_463_4031_0, i_10_463_4117_0, i_10_463_4127_0,
    i_10_463_4274_0, i_10_463_4280_0, i_10_463_4365_0, i_10_463_4585_0,
    o_10_463_0_0  );
  input  i_10_463_243_0, i_10_463_252_0, i_10_463_263_0, i_10_463_286_0,
    i_10_463_317_0, i_10_463_319_0, i_10_463_320_0, i_10_463_395_0,
    i_10_463_512_0, i_10_463_621_0, i_10_463_687_0, i_10_463_688_0,
    i_10_463_865_0, i_10_463_1001_0, i_10_463_1003_0, i_10_463_1004_0,
    i_10_463_1058_0, i_10_463_1081_0, i_10_463_1084_0, i_10_463_1134_0,
    i_10_463_1135_0, i_10_463_1152_0, i_10_463_1153_0, i_10_463_1223_0,
    i_10_463_1237_0, i_10_463_1263_0, i_10_463_1300_0, i_10_463_1435_0,
    i_10_463_1436_0, i_10_463_1530_0, i_10_463_1535_0, i_10_463_1548_0,
    i_10_463_1551_0, i_10_463_1552_0, i_10_463_1580_0, i_10_463_1625_0,
    i_10_463_1628_0, i_10_463_1730_0, i_10_463_1733_0, i_10_463_1808_0,
    i_10_463_1810_0, i_10_463_1821_0, i_10_463_1906_0, i_10_463_1915_0,
    i_10_463_2020_0, i_10_463_2030_0, i_10_463_2033_0, i_10_463_2064_0,
    i_10_463_2111_0, i_10_463_2200_0, i_10_463_2340_0, i_10_463_2345_0,
    i_10_463_2349_0, i_10_463_2352_0, i_10_463_2353_0, i_10_463_2363_0,
    i_10_463_2380_0, i_10_463_2406_0, i_10_463_2453_0, i_10_463_2468_0,
    i_10_463_2567_0, i_10_463_2570_0, i_10_463_2703_0, i_10_463_2731_0,
    i_10_463_2732_0, i_10_463_2741_0, i_10_463_2744_0, i_10_463_2782_0,
    i_10_463_2808_0, i_10_463_2839_0, i_10_463_2840_0, i_10_463_3043_0,
    i_10_463_3047_0, i_10_463_3091_0, i_10_463_3195_0, i_10_463_3202_0,
    i_10_463_3271_0, i_10_463_3317_0, i_10_463_3320_0, i_10_463_3335_0,
    i_10_463_3353_0, i_10_463_3393_0, i_10_463_3473_0, i_10_463_3545_0,
    i_10_463_3560_0, i_10_463_3612_0, i_10_463_3663_0, i_10_463_3789_0,
    i_10_463_3842_0, i_10_463_3911_0, i_10_463_3942_0, i_10_463_3946_0,
    i_10_463_3999_0, i_10_463_4031_0, i_10_463_4117_0, i_10_463_4127_0,
    i_10_463_4274_0, i_10_463_4280_0, i_10_463_4365_0, i_10_463_4585_0;
  output o_10_463_0_0;
  assign o_10_463_0_0 = 0;
endmodule



// Benchmark "kernel_10_464" written by ABC on Sun Jul 19 10:29:08 2020

module kernel_10_464 ( 
    i_10_464_153_0, i_10_464_172_0, i_10_464_285_0, i_10_464_315_0,
    i_10_464_387_0, i_10_464_393_0, i_10_464_410_0, i_10_464_423_0,
    i_10_464_433_0, i_10_464_910_0, i_10_464_946_0, i_10_464_958_0,
    i_10_464_966_0, i_10_464_1038_0, i_10_464_1051_0, i_10_464_1209_0,
    i_10_464_1240_0, i_10_464_1241_0, i_10_464_1262_0, i_10_464_1307_0,
    i_10_464_1580_0, i_10_464_1614_0, i_10_464_1630_0, i_10_464_1683_0,
    i_10_464_1684_0, i_10_464_1685_0, i_10_464_1688_0, i_10_464_1747_0,
    i_10_464_1819_0, i_10_464_1820_0, i_10_464_1822_0, i_10_464_1825_0,
    i_10_464_1826_0, i_10_464_1893_0, i_10_464_1954_0, i_10_464_2018_0,
    i_10_464_2178_0, i_10_464_2182_0, i_10_464_2244_0, i_10_464_2287_0,
    i_10_464_2291_0, i_10_464_2365_0, i_10_464_2380_0, i_10_464_2382_0,
    i_10_464_2385_0, i_10_464_2386_0, i_10_464_2461_0, i_10_464_2513_0,
    i_10_464_2565_0, i_10_464_2566_0, i_10_464_2569_0, i_10_464_2587_0,
    i_10_464_2660_0, i_10_464_2701_0, i_10_464_2712_0, i_10_464_2718_0,
    i_10_464_2719_0, i_10_464_2724_0, i_10_464_2728_0, i_10_464_2731_0,
    i_10_464_2732_0, i_10_464_2743_0, i_10_464_2834_0, i_10_464_2843_0,
    i_10_464_2866_0, i_10_464_2867_0, i_10_464_2882_0, i_10_464_2920_0,
    i_10_464_2979_0, i_10_464_2982_0, i_10_464_3042_0, i_10_464_3047_0,
    i_10_464_3089_0, i_10_464_3100_0, i_10_464_3166_0, i_10_464_3199_0,
    i_10_464_3202_0, i_10_464_3415_0, i_10_464_3465_0, i_10_464_3540_0,
    i_10_464_3610_0, i_10_464_3613_0, i_10_464_3652_0, i_10_464_3686_0,
    i_10_464_3799_0, i_10_464_3800_0, i_10_464_3820_0, i_10_464_3836_0,
    i_10_464_3839_0, i_10_464_3852_0, i_10_464_3988_0, i_10_464_4053_0,
    i_10_464_4144_0, i_10_464_4192_0, i_10_464_4270_0, i_10_464_4271_0,
    i_10_464_4275_0, i_10_464_4283_0, i_10_464_4308_0, i_10_464_4451_0,
    o_10_464_0_0  );
  input  i_10_464_153_0, i_10_464_172_0, i_10_464_285_0, i_10_464_315_0,
    i_10_464_387_0, i_10_464_393_0, i_10_464_410_0, i_10_464_423_0,
    i_10_464_433_0, i_10_464_910_0, i_10_464_946_0, i_10_464_958_0,
    i_10_464_966_0, i_10_464_1038_0, i_10_464_1051_0, i_10_464_1209_0,
    i_10_464_1240_0, i_10_464_1241_0, i_10_464_1262_0, i_10_464_1307_0,
    i_10_464_1580_0, i_10_464_1614_0, i_10_464_1630_0, i_10_464_1683_0,
    i_10_464_1684_0, i_10_464_1685_0, i_10_464_1688_0, i_10_464_1747_0,
    i_10_464_1819_0, i_10_464_1820_0, i_10_464_1822_0, i_10_464_1825_0,
    i_10_464_1826_0, i_10_464_1893_0, i_10_464_1954_0, i_10_464_2018_0,
    i_10_464_2178_0, i_10_464_2182_0, i_10_464_2244_0, i_10_464_2287_0,
    i_10_464_2291_0, i_10_464_2365_0, i_10_464_2380_0, i_10_464_2382_0,
    i_10_464_2385_0, i_10_464_2386_0, i_10_464_2461_0, i_10_464_2513_0,
    i_10_464_2565_0, i_10_464_2566_0, i_10_464_2569_0, i_10_464_2587_0,
    i_10_464_2660_0, i_10_464_2701_0, i_10_464_2712_0, i_10_464_2718_0,
    i_10_464_2719_0, i_10_464_2724_0, i_10_464_2728_0, i_10_464_2731_0,
    i_10_464_2732_0, i_10_464_2743_0, i_10_464_2834_0, i_10_464_2843_0,
    i_10_464_2866_0, i_10_464_2867_0, i_10_464_2882_0, i_10_464_2920_0,
    i_10_464_2979_0, i_10_464_2982_0, i_10_464_3042_0, i_10_464_3047_0,
    i_10_464_3089_0, i_10_464_3100_0, i_10_464_3166_0, i_10_464_3199_0,
    i_10_464_3202_0, i_10_464_3415_0, i_10_464_3465_0, i_10_464_3540_0,
    i_10_464_3610_0, i_10_464_3613_0, i_10_464_3652_0, i_10_464_3686_0,
    i_10_464_3799_0, i_10_464_3800_0, i_10_464_3820_0, i_10_464_3836_0,
    i_10_464_3839_0, i_10_464_3852_0, i_10_464_3988_0, i_10_464_4053_0,
    i_10_464_4144_0, i_10_464_4192_0, i_10_464_4270_0, i_10_464_4271_0,
    i_10_464_4275_0, i_10_464_4283_0, i_10_464_4308_0, i_10_464_4451_0;
  output o_10_464_0_0;
  assign o_10_464_0_0 = 0;
endmodule



// Benchmark "kernel_10_465" written by ABC on Sun Jul 19 10:29:09 2020

module kernel_10_465 ( 
    i_10_465_121_0, i_10_465_152_0, i_10_465_176_0, i_10_465_186_0,
    i_10_465_187_0, i_10_465_222_0, i_10_465_224_0, i_10_465_318_0,
    i_10_465_441_0, i_10_465_446_0, i_10_465_449_0, i_10_465_460_0,
    i_10_465_463_0, i_10_465_464_0, i_10_465_466_0, i_10_465_467_0,
    i_10_465_510_0, i_10_465_717_0, i_10_465_797_0, i_10_465_800_0,
    i_10_465_908_0, i_10_465_968_0, i_10_465_1040_0, i_10_465_1247_0,
    i_10_465_1250_0, i_10_465_1542_0, i_10_465_1543_0, i_10_465_1578_0,
    i_10_465_1579_0, i_10_465_1652_0, i_10_465_1653_0, i_10_465_1685_0,
    i_10_465_1822_0, i_10_465_1823_0, i_10_465_1824_0, i_10_465_1826_0,
    i_10_465_1912_0, i_10_465_1952_0, i_10_465_1995_0, i_10_465_2004_0,
    i_10_465_2005_0, i_10_465_2006_0, i_10_465_2095_0, i_10_465_2182_0,
    i_10_465_2203_0, i_10_465_2364_0, i_10_465_2379_0, i_10_465_2380_0,
    i_10_465_2381_0, i_10_465_2384_0, i_10_465_2453_0, i_10_465_2456_0,
    i_10_465_2471_0, i_10_465_2473_0, i_10_465_2474_0, i_10_465_2628_0,
    i_10_465_2633_0, i_10_465_2700_0, i_10_465_2703_0, i_10_465_2715_0,
    i_10_465_2717_0, i_10_465_2734_0, i_10_465_2782_0, i_10_465_2830_0,
    i_10_465_2833_0, i_10_465_2834_0, i_10_465_2886_0, i_10_465_3034_0,
    i_10_465_3035_0, i_10_465_3037_0, i_10_465_3038_0, i_10_465_3040_0,
    i_10_465_3041_0, i_10_465_3076_0, i_10_465_3155_0, i_10_465_3199_0,
    i_10_465_3200_0, i_10_465_3269_0, i_10_465_3270_0, i_10_465_3271_0,
    i_10_465_3274_0, i_10_465_3387_0, i_10_465_3389_0, i_10_465_3406_0,
    i_10_465_3587_0, i_10_465_3589_0, i_10_465_3590_0, i_10_465_3615_0,
    i_10_465_3650_0, i_10_465_3651_0, i_10_465_3787_0, i_10_465_3788_0,
    i_10_465_3837_0, i_10_465_3860_0, i_10_465_4121_0, i_10_465_4175_0,
    i_10_465_4286_0, i_10_465_4288_0, i_10_465_4291_0, i_10_465_4568_0,
    o_10_465_0_0  );
  input  i_10_465_121_0, i_10_465_152_0, i_10_465_176_0, i_10_465_186_0,
    i_10_465_187_0, i_10_465_222_0, i_10_465_224_0, i_10_465_318_0,
    i_10_465_441_0, i_10_465_446_0, i_10_465_449_0, i_10_465_460_0,
    i_10_465_463_0, i_10_465_464_0, i_10_465_466_0, i_10_465_467_0,
    i_10_465_510_0, i_10_465_717_0, i_10_465_797_0, i_10_465_800_0,
    i_10_465_908_0, i_10_465_968_0, i_10_465_1040_0, i_10_465_1247_0,
    i_10_465_1250_0, i_10_465_1542_0, i_10_465_1543_0, i_10_465_1578_0,
    i_10_465_1579_0, i_10_465_1652_0, i_10_465_1653_0, i_10_465_1685_0,
    i_10_465_1822_0, i_10_465_1823_0, i_10_465_1824_0, i_10_465_1826_0,
    i_10_465_1912_0, i_10_465_1952_0, i_10_465_1995_0, i_10_465_2004_0,
    i_10_465_2005_0, i_10_465_2006_0, i_10_465_2095_0, i_10_465_2182_0,
    i_10_465_2203_0, i_10_465_2364_0, i_10_465_2379_0, i_10_465_2380_0,
    i_10_465_2381_0, i_10_465_2384_0, i_10_465_2453_0, i_10_465_2456_0,
    i_10_465_2471_0, i_10_465_2473_0, i_10_465_2474_0, i_10_465_2628_0,
    i_10_465_2633_0, i_10_465_2700_0, i_10_465_2703_0, i_10_465_2715_0,
    i_10_465_2717_0, i_10_465_2734_0, i_10_465_2782_0, i_10_465_2830_0,
    i_10_465_2833_0, i_10_465_2834_0, i_10_465_2886_0, i_10_465_3034_0,
    i_10_465_3035_0, i_10_465_3037_0, i_10_465_3038_0, i_10_465_3040_0,
    i_10_465_3041_0, i_10_465_3076_0, i_10_465_3155_0, i_10_465_3199_0,
    i_10_465_3200_0, i_10_465_3269_0, i_10_465_3270_0, i_10_465_3271_0,
    i_10_465_3274_0, i_10_465_3387_0, i_10_465_3389_0, i_10_465_3406_0,
    i_10_465_3587_0, i_10_465_3589_0, i_10_465_3590_0, i_10_465_3615_0,
    i_10_465_3650_0, i_10_465_3651_0, i_10_465_3787_0, i_10_465_3788_0,
    i_10_465_3837_0, i_10_465_3860_0, i_10_465_4121_0, i_10_465_4175_0,
    i_10_465_4286_0, i_10_465_4288_0, i_10_465_4291_0, i_10_465_4568_0;
  output o_10_465_0_0;
  assign o_10_465_0_0 = ~((~i_10_465_446_0 & ((~i_10_465_187_0 & ~i_10_465_467_0 & ~i_10_465_1823_0 & ~i_10_465_2473_0 & ~i_10_465_2703_0 & ~i_10_465_3037_0 & i_10_465_3837_0) | (~i_10_465_449_0 & ~i_10_465_460_0 & i_10_465_2203_0 & ~i_10_465_3041_0 & i_10_465_3199_0 & ~i_10_465_3270_0 & ~i_10_465_4175_0 & ~i_10_465_4288_0))) | (~i_10_465_187_0 & ((~i_10_465_449_0 & ~i_10_465_463_0 & ~i_10_465_464_0 & ~i_10_465_2473_0 & ~i_10_465_2700_0 & ~i_10_465_2717_0 & ~i_10_465_3274_0 & ~i_10_465_3590_0 & ~i_10_465_3787_0) | (~i_10_465_2886_0 & i_10_465_3274_0 & i_10_465_3387_0 & ~i_10_465_4291_0))) | (~i_10_465_2384_0 & ((~i_10_465_800_0 & ((~i_10_465_121_0 & ~i_10_465_968_0 & i_10_465_1824_0 & i_10_465_1826_0 & ~i_10_465_2473_0 & ~i_10_465_2474_0 & ~i_10_465_2703_0 & i_10_465_3650_0) | (~i_10_465_460_0 & ~i_10_465_467_0 & ~i_10_465_908_0 & i_10_465_1652_0 & ~i_10_465_2364_0 & ~i_10_465_3406_0 & ~i_10_465_3587_0 & ~i_10_465_3860_0))) | (~i_10_465_2203_0 & ~i_10_465_2456_0 & ~i_10_465_2734_0 & ~i_10_465_2830_0 & ~i_10_465_3041_0 & i_10_465_3787_0 & ~i_10_465_3860_0 & ~i_10_465_4286_0))) | (~i_10_465_4288_0 & ((~i_10_465_449_0 & ((~i_10_465_467_0 & i_10_465_2715_0 & ~i_10_465_2734_0 & ~i_10_465_3037_0) | (~i_10_465_1250_0 & ~i_10_465_1822_0 & ~i_10_465_1912_0 & ~i_10_465_2628_0 & ~i_10_465_2633_0 & ~i_10_465_3589_0 & ~i_10_465_4291_0))) | (~i_10_465_4175_0 & ((~i_10_465_460_0 & ~i_10_465_467_0 & ~i_10_465_908_0 & ~i_10_465_1250_0 & ~i_10_465_1579_0 & ~i_10_465_2471_0 & ~i_10_465_2628_0 & ~i_10_465_2715_0 & ~i_10_465_2830_0 & ~i_10_465_3041_0 & ~i_10_465_3590_0 & ~i_10_465_3837_0) | (~i_10_465_1824_0 & ~i_10_465_1952_0 & i_10_465_3271_0 & ~i_10_465_3860_0))) | (~i_10_465_121_0 & ~i_10_465_466_0 & ~i_10_465_797_0 & ~i_10_465_1247_0 & i_10_465_1822_0 & i_10_465_2628_0 & ~i_10_465_3035_0 & ~i_10_465_4286_0))) | (~i_10_465_460_0 & ((~i_10_465_467_0 & ~i_10_465_717_0 & ~i_10_465_797_0 & i_10_465_1824_0 & ~i_10_465_3040_0 & ~i_10_465_3389_0) | (~i_10_465_1040_0 & ~i_10_465_2453_0 & ~i_10_465_2473_0 & ~i_10_465_2734_0 & ~i_10_465_2830_0 & ~i_10_465_3034_0 & ~i_10_465_3035_0 & ~i_10_465_3038_0 & ~i_10_465_3587_0 & ~i_10_465_3590_0 & ~i_10_465_4286_0))) | (~i_10_465_1247_0 & ((~i_10_465_152_0 & ~i_10_465_2006_0 & ~i_10_465_2381_0 & i_10_465_2833_0 & i_10_465_2834_0 & ~i_10_465_3034_0 & ~i_10_465_3038_0 & ~i_10_465_3787_0 & ~i_10_465_3788_0) | (i_10_465_463_0 & ~i_10_465_908_0 & ~i_10_465_1685_0 & ~i_10_465_1826_0 & ~i_10_465_2633_0 & ~i_10_465_2782_0 & ~i_10_465_2830_0 & ~i_10_465_3035_0 & ~i_10_465_3037_0 & ~i_10_465_3387_0 & ~i_10_465_3587_0 & ~i_10_465_3589_0 & ~i_10_465_4286_0 & ~i_10_465_4568_0))) | (~i_10_465_4286_0 & ((~i_10_465_449_0 & ((~i_10_465_466_0 & ~i_10_465_1912_0 & ~i_10_465_2717_0 & ~i_10_465_3034_0 & ~i_10_465_3041_0 & ~i_10_465_3389_0 & i_10_465_3837_0) | (~i_10_465_467_0 & ~i_10_465_717_0 & ~i_10_465_908_0 & ~i_10_465_1685_0 & ~i_10_465_1822_0 & ~i_10_465_1823_0 & ~i_10_465_2473_0 & ~i_10_465_2474_0 & ~i_10_465_2700_0 & ~i_10_465_3406_0 & ~i_10_465_3651_0 & ~i_10_465_3860_0))) | (~i_10_465_467_0 & ((~i_10_465_466_0 & ~i_10_465_908_0 & ~i_10_465_968_0 & ~i_10_465_1824_0 & ~i_10_465_2628_0 & ~i_10_465_3034_0 & ~i_10_465_3587_0 & ~i_10_465_3650_0 & ~i_10_465_4121_0) | (~i_10_465_1822_0 & ~i_10_465_3038_0 & ~i_10_465_3040_0 & ~i_10_465_3389_0 & ~i_10_465_3589_0 & ~i_10_465_4568_0))) | (~i_10_465_3651_0 & ((i_10_465_2379_0 & i_10_465_2628_0) | (i_10_465_318_0 & ~i_10_465_1824_0 & ~i_10_465_2005_0 & ~i_10_465_2782_0))) | (~i_10_465_441_0 & ~i_10_465_463_0 & ~i_10_465_1823_0 & i_10_465_1824_0 & ~i_10_465_2004_0 & ~i_10_465_2474_0 & ~i_10_465_2734_0))) | (i_10_465_318_0 & ((~i_10_465_449_0 & i_10_465_1578_0 & i_10_465_2203_0 & ~i_10_465_3590_0) | (~i_10_465_186_0 & i_10_465_4286_0 & i_10_465_4291_0))) | (~i_10_465_449_0 & ((~i_10_465_224_0 & i_10_465_1543_0 & ~i_10_465_2633_0 & ~i_10_465_2715_0 & ~i_10_465_3037_0) | (~i_10_465_121_0 & ~i_10_465_152_0 & ~i_10_465_464_0 & ~i_10_465_797_0 & ~i_10_465_2456_0 & ~i_10_465_2471_0 & ~i_10_465_2734_0 & ~i_10_465_3034_0 & ~i_10_465_3041_0 & ~i_10_465_3271_0 & ~i_10_465_3274_0 & ~i_10_465_3615_0 & ~i_10_465_3837_0))) | (~i_10_465_121_0 & ((~i_10_465_1822_0 & ~i_10_465_1826_0 & ~i_10_465_2703_0 & ~i_10_465_3035_0 & ~i_10_465_3200_0 & i_10_465_3651_0) | (~i_10_465_176_0 & ~i_10_465_466_0 & ~i_10_465_1823_0 & i_10_465_1912_0 & ~i_10_465_3650_0 & ~i_10_465_3837_0 & ~i_10_465_4291_0 & ~i_10_465_4568_0))) | (~i_10_465_1040_0 & ((~i_10_465_152_0 & ~i_10_465_717_0 & ((~i_10_465_466_0 & i_10_465_3270_0) | (~i_10_465_463_0 & ~i_10_465_908_0 & ~i_10_465_968_0 & ~i_10_465_2453_0 & ~i_10_465_2473_0 & ~i_10_465_3590_0))) | (~i_10_465_1823_0 & i_10_465_2380_0 & i_10_465_2700_0 & ~i_10_465_3590_0 & ~i_10_465_3837_0))) | (~i_10_465_463_0 & ((i_10_465_2380_0 & i_10_465_2628_0) | (~i_10_465_2364_0 & i_10_465_2830_0 & i_10_465_3274_0 & ~i_10_465_3788_0 & ~i_10_465_3837_0))) | (~i_10_465_464_0 & ((~i_10_465_467_0 & ~i_10_465_908_0 & ~i_10_465_968_0 & ~i_10_465_1822_0 & ~i_10_465_2005_0 & ~i_10_465_2006_0 & i_10_465_2456_0) | (i_10_465_1579_0 & ~i_10_465_3037_0 & ~i_10_465_3590_0 & ~i_10_465_4121_0))) | (i_10_465_1579_0 & ((~i_10_465_3035_0 & i_10_465_3269_0) | (i_10_465_2700_0 & i_10_465_4288_0))) | (i_10_465_2628_0 & ((i_10_465_1653_0 & ~i_10_465_3199_0 & i_10_465_3615_0 & i_10_465_3651_0) | (~i_10_465_797_0 & ~i_10_465_1822_0 & ~i_10_465_3589_0 & i_10_465_4288_0 & ~i_10_465_4291_0))) | (~i_10_465_797_0 & ((~i_10_465_1823_0 & ~i_10_465_2633_0 & i_10_465_3587_0 & i_10_465_4286_0) | (~i_10_465_1653_0 & i_10_465_2703_0 & i_10_465_4288_0))) | (~i_10_465_466_0 & i_10_465_2182_0 & ~i_10_465_3038_0));
endmodule



// Benchmark "kernel_10_466" written by ABC on Sun Jul 19 10:29:11 2020

module kernel_10_466 ( 
    i_10_466_217_0, i_10_466_220_0, i_10_466_221_0, i_10_466_280_0,
    i_10_466_281_0, i_10_466_282_0, i_10_466_283_0, i_10_466_284_0,
    i_10_466_316_0, i_10_466_324_0, i_10_466_390_0, i_10_466_391_0,
    i_10_466_406_0, i_10_466_443_0, i_10_466_445_0, i_10_466_449_0,
    i_10_466_459_0, i_10_466_464_0, i_10_466_505_0, i_10_466_506_0,
    i_10_466_509_0, i_10_466_749_0, i_10_466_797_0, i_10_466_1135_0,
    i_10_466_1233_0, i_10_466_1236_0, i_10_466_1250_0, i_10_466_1305_0,
    i_10_466_1345_0, i_10_466_1346_0, i_10_466_1431_0, i_10_466_1432_0,
    i_10_466_1433_0, i_10_466_1540_0, i_10_466_1552_0, i_10_466_1621_0,
    i_10_466_1651_0, i_10_466_1654_0, i_10_466_1683_0, i_10_466_1689_0,
    i_10_466_1824_0, i_10_466_1825_0, i_10_466_1981_0, i_10_466_1990_0,
    i_10_466_2017_0, i_10_466_2351_0, i_10_466_2359_0, i_10_466_2380_0,
    i_10_466_2407_0, i_10_466_2451_0, i_10_466_2628_0, i_10_466_2629_0,
    i_10_466_2630_0, i_10_466_2631_0, i_10_466_2632_0, i_10_466_2656_0,
    i_10_466_2701_0, i_10_466_2709_0, i_10_466_2710_0, i_10_466_2718_0,
    i_10_466_2723_0, i_10_466_2884_0, i_10_466_2917_0, i_10_466_2979_0,
    i_10_466_3044_0, i_10_466_3070_0, i_10_466_3152_0, i_10_466_3153_0,
    i_10_466_3156_0, i_10_466_3196_0, i_10_466_3277_0, i_10_466_3278_0,
    i_10_466_3281_0, i_10_466_3385_0, i_10_466_3388_0, i_10_466_3389_0,
    i_10_466_3391_0, i_10_466_3392_0, i_10_466_3523_0, i_10_466_3556_0,
    i_10_466_3728_0, i_10_466_3784_0, i_10_466_3834_0, i_10_466_3837_0,
    i_10_466_3846_0, i_10_466_3859_0, i_10_466_3979_0, i_10_466_3985_0,
    i_10_466_3991_0, i_10_466_4114_0, i_10_466_4115_0, i_10_466_4116_0,
    i_10_466_4117_0, i_10_466_4118_0, i_10_466_4122_0, i_10_466_4168_0,
    i_10_466_4276_0, i_10_466_4566_0, i_10_466_4567_0, i_10_466_4568_0,
    o_10_466_0_0  );
  input  i_10_466_217_0, i_10_466_220_0, i_10_466_221_0, i_10_466_280_0,
    i_10_466_281_0, i_10_466_282_0, i_10_466_283_0, i_10_466_284_0,
    i_10_466_316_0, i_10_466_324_0, i_10_466_390_0, i_10_466_391_0,
    i_10_466_406_0, i_10_466_443_0, i_10_466_445_0, i_10_466_449_0,
    i_10_466_459_0, i_10_466_464_0, i_10_466_505_0, i_10_466_506_0,
    i_10_466_509_0, i_10_466_749_0, i_10_466_797_0, i_10_466_1135_0,
    i_10_466_1233_0, i_10_466_1236_0, i_10_466_1250_0, i_10_466_1305_0,
    i_10_466_1345_0, i_10_466_1346_0, i_10_466_1431_0, i_10_466_1432_0,
    i_10_466_1433_0, i_10_466_1540_0, i_10_466_1552_0, i_10_466_1621_0,
    i_10_466_1651_0, i_10_466_1654_0, i_10_466_1683_0, i_10_466_1689_0,
    i_10_466_1824_0, i_10_466_1825_0, i_10_466_1981_0, i_10_466_1990_0,
    i_10_466_2017_0, i_10_466_2351_0, i_10_466_2359_0, i_10_466_2380_0,
    i_10_466_2407_0, i_10_466_2451_0, i_10_466_2628_0, i_10_466_2629_0,
    i_10_466_2630_0, i_10_466_2631_0, i_10_466_2632_0, i_10_466_2656_0,
    i_10_466_2701_0, i_10_466_2709_0, i_10_466_2710_0, i_10_466_2718_0,
    i_10_466_2723_0, i_10_466_2884_0, i_10_466_2917_0, i_10_466_2979_0,
    i_10_466_3044_0, i_10_466_3070_0, i_10_466_3152_0, i_10_466_3153_0,
    i_10_466_3156_0, i_10_466_3196_0, i_10_466_3277_0, i_10_466_3278_0,
    i_10_466_3281_0, i_10_466_3385_0, i_10_466_3388_0, i_10_466_3389_0,
    i_10_466_3391_0, i_10_466_3392_0, i_10_466_3523_0, i_10_466_3556_0,
    i_10_466_3728_0, i_10_466_3784_0, i_10_466_3834_0, i_10_466_3837_0,
    i_10_466_3846_0, i_10_466_3859_0, i_10_466_3979_0, i_10_466_3985_0,
    i_10_466_3991_0, i_10_466_4114_0, i_10_466_4115_0, i_10_466_4116_0,
    i_10_466_4117_0, i_10_466_4118_0, i_10_466_4122_0, i_10_466_4168_0,
    i_10_466_4276_0, i_10_466_4566_0, i_10_466_4567_0, i_10_466_4568_0;
  output o_10_466_0_0;
  assign o_10_466_0_0 = ~((~i_10_466_316_0 & ((~i_10_466_390_0 & ~i_10_466_1689_0 & ~i_10_466_2451_0 & ~i_10_466_3278_0 & ~i_10_466_3388_0 & ~i_10_466_3846_0 & ~i_10_466_4168_0) | (i_10_466_221_0 & ~i_10_466_2351_0 & ~i_10_466_4276_0))) | (~i_10_466_1233_0 & ((~i_10_466_1433_0 & ~i_10_466_2723_0 & ~i_10_466_2884_0 & ~i_10_466_3281_0 & ~i_10_466_3523_0 & ~i_10_466_3784_0) | (~i_10_466_391_0 & ~i_10_466_2407_0 & ~i_10_466_2451_0 & ~i_10_466_2710_0 & ~i_10_466_3278_0 & ~i_10_466_3392_0 & ~i_10_466_3834_0))) | (~i_10_466_1552_0 & ((i_10_466_1824_0 & ~i_10_466_2709_0 & ~i_10_466_2710_0 & ~i_10_466_3388_0 & ~i_10_466_3389_0 & ~i_10_466_3846_0) | (~i_10_466_1683_0 & ~i_10_466_3277_0 & ~i_10_466_3278_0 & i_10_466_4117_0))) | (~i_10_466_391_0 & ((~i_10_466_1346_0 & ((~i_10_466_1683_0 & ~i_10_466_2351_0 & ~i_10_466_3281_0 & ~i_10_466_3837_0 & ~i_10_466_3985_0) | (~i_10_466_2451_0 & ~i_10_466_2718_0 & ~i_10_466_2884_0 & ~i_10_466_3044_0 & ~i_10_466_3070_0 & i_10_466_3388_0 & ~i_10_466_3784_0 & ~i_10_466_4118_0 & ~i_10_466_4122_0 & ~i_10_466_4568_0))) | (~i_10_466_3985_0 & ((~i_10_466_1432_0 & ((~i_10_466_1824_0 & ~i_10_466_2351_0 & ~i_10_466_3281_0 & ~i_10_466_3392_0) | (~i_10_466_282_0 & ~i_10_466_3277_0 & ~i_10_466_3391_0 & ~i_10_466_4276_0 & ~i_10_466_4568_0))) | (~i_10_466_281_0 & ~i_10_466_1305_0 & i_10_466_1824_0 & ~i_10_466_3044_0 & ~i_10_466_4122_0))) | (~i_10_466_1431_0 & ~i_10_466_2710_0 & ~i_10_466_3044_0 & ~i_10_466_3391_0 & ~i_10_466_3392_0))) | (~i_10_466_282_0 & ((~i_10_466_324_0 & ~i_10_466_1346_0 & ~i_10_466_1540_0 & ~i_10_466_1621_0 & i_10_466_2632_0) | (~i_10_466_2407_0 & ~i_10_466_3278_0 & i_10_466_3784_0 & ~i_10_466_3979_0))) | (~i_10_466_1346_0 & ((~i_10_466_390_0 & ~i_10_466_797_0 & ~i_10_466_1689_0 & ~i_10_466_2710_0 & ~i_10_466_3044_0 & ~i_10_466_3281_0 & ~i_10_466_3846_0) | (~i_10_466_2359_0 & ~i_10_466_3392_0 & ~i_10_466_4276_0 & i_10_466_4567_0))) | (~i_10_466_390_0 & ((~i_10_466_283_0 & i_10_466_464_0 & i_10_466_3277_0 & ~i_10_466_3985_0) | (i_10_466_283_0 & ~i_10_466_445_0 & ~i_10_466_459_0 & ~i_10_466_1433_0 & ~i_10_466_2628_0 & ~i_10_466_2884_0 & ~i_10_466_3389_0 & ~i_10_466_3391_0 & ~i_10_466_4168_0 & ~i_10_466_4567_0))) | (~i_10_466_3281_0 & ((~i_10_466_3391_0 & ~i_10_466_3837_0 & i_10_466_3859_0) | (i_10_466_797_0 & ~i_10_466_1345_0 & ~i_10_466_2656_0 & i_10_466_3523_0 & ~i_10_466_4567_0))) | (~i_10_466_464_0 & ~i_10_466_1432_0 & i_10_466_1825_0 & ~i_10_466_3391_0 & ~i_10_466_3392_0 & ~i_10_466_2380_0 & ~i_10_466_3388_0) | (~i_10_466_280_0 & i_10_466_3196_0 & ~i_10_466_3278_0 & ~i_10_466_3834_0 & ~i_10_466_3985_0) | (i_10_466_3392_0 & i_10_466_4566_0));
endmodule



// Benchmark "kernel_10_467" written by ABC on Sun Jul 19 10:29:12 2020

module kernel_10_467 ( 
    i_10_467_176_0, i_10_467_254_0, i_10_467_263_0, i_10_467_266_0,
    i_10_467_272_0, i_10_467_323_0, i_10_467_407_0, i_10_467_412_0,
    i_10_467_445_0, i_10_467_500_0, i_10_467_502_0, i_10_467_506_0,
    i_10_467_509_0, i_10_467_563_0, i_10_467_595_0, i_10_467_877_0,
    i_10_467_1003_0, i_10_467_1028_0, i_10_467_1109_0, i_10_467_1111_0,
    i_10_467_1112_0, i_10_467_1220_0, i_10_467_1235_0, i_10_467_1239_0,
    i_10_467_1246_0, i_10_467_1283_0, i_10_467_1300_0, i_10_467_1303_0,
    i_10_467_1360_0, i_10_467_1436_0, i_10_467_1451_0, i_10_467_1454_0,
    i_10_467_1541_0, i_10_467_1544_0, i_10_467_1546_0, i_10_467_1580_0,
    i_10_467_1583_0, i_10_467_1622_0, i_10_467_1625_0, i_10_467_1688_0,
    i_10_467_1733_0, i_10_467_1808_0, i_10_467_1824_0, i_10_467_1982_0,
    i_10_467_2003_0, i_10_467_2006_0, i_10_467_2027_0, i_10_467_2108_0,
    i_10_467_2204_0, i_10_467_2351_0, i_10_467_2361_0, i_10_467_2364_0,
    i_10_467_2467_0, i_10_467_2533_0, i_10_467_2534_0, i_10_467_2567_0,
    i_10_467_2570_0, i_10_467_2609_0, i_10_467_2658_0, i_10_467_2705_0,
    i_10_467_2722_0, i_10_467_2731_0, i_10_467_2789_0, i_10_467_2830_0,
    i_10_467_2833_0, i_10_467_2837_0, i_10_467_2867_0, i_10_467_2923_0,
    i_10_467_3034_0, i_10_467_3041_0, i_10_467_3314_0, i_10_467_3316_0,
    i_10_467_3317_0, i_10_467_3332_0, i_10_467_3350_0, i_10_467_3391_0,
    i_10_467_3392_0, i_10_467_3402_0, i_10_467_3443_0, i_10_467_3466_0,
    i_10_467_3583_0, i_10_467_3587_0, i_10_467_3797_0, i_10_467_3835_0,
    i_10_467_3836_0, i_10_467_3842_0, i_10_467_3848_0, i_10_467_3983_0,
    i_10_467_4010_0, i_10_467_4126_0, i_10_467_4127_0, i_10_467_4130_0,
    i_10_467_4154_0, i_10_467_4171_0, i_10_467_4268_0, i_10_467_4288_0,
    i_10_467_4379_0, i_10_467_4550_0, i_10_467_4565_0, i_10_467_4568_0,
    o_10_467_0_0  );
  input  i_10_467_176_0, i_10_467_254_0, i_10_467_263_0, i_10_467_266_0,
    i_10_467_272_0, i_10_467_323_0, i_10_467_407_0, i_10_467_412_0,
    i_10_467_445_0, i_10_467_500_0, i_10_467_502_0, i_10_467_506_0,
    i_10_467_509_0, i_10_467_563_0, i_10_467_595_0, i_10_467_877_0,
    i_10_467_1003_0, i_10_467_1028_0, i_10_467_1109_0, i_10_467_1111_0,
    i_10_467_1112_0, i_10_467_1220_0, i_10_467_1235_0, i_10_467_1239_0,
    i_10_467_1246_0, i_10_467_1283_0, i_10_467_1300_0, i_10_467_1303_0,
    i_10_467_1360_0, i_10_467_1436_0, i_10_467_1451_0, i_10_467_1454_0,
    i_10_467_1541_0, i_10_467_1544_0, i_10_467_1546_0, i_10_467_1580_0,
    i_10_467_1583_0, i_10_467_1622_0, i_10_467_1625_0, i_10_467_1688_0,
    i_10_467_1733_0, i_10_467_1808_0, i_10_467_1824_0, i_10_467_1982_0,
    i_10_467_2003_0, i_10_467_2006_0, i_10_467_2027_0, i_10_467_2108_0,
    i_10_467_2204_0, i_10_467_2351_0, i_10_467_2361_0, i_10_467_2364_0,
    i_10_467_2467_0, i_10_467_2533_0, i_10_467_2534_0, i_10_467_2567_0,
    i_10_467_2570_0, i_10_467_2609_0, i_10_467_2658_0, i_10_467_2705_0,
    i_10_467_2722_0, i_10_467_2731_0, i_10_467_2789_0, i_10_467_2830_0,
    i_10_467_2833_0, i_10_467_2837_0, i_10_467_2867_0, i_10_467_2923_0,
    i_10_467_3034_0, i_10_467_3041_0, i_10_467_3314_0, i_10_467_3316_0,
    i_10_467_3317_0, i_10_467_3332_0, i_10_467_3350_0, i_10_467_3391_0,
    i_10_467_3392_0, i_10_467_3402_0, i_10_467_3443_0, i_10_467_3466_0,
    i_10_467_3583_0, i_10_467_3587_0, i_10_467_3797_0, i_10_467_3835_0,
    i_10_467_3836_0, i_10_467_3842_0, i_10_467_3848_0, i_10_467_3983_0,
    i_10_467_4010_0, i_10_467_4126_0, i_10_467_4127_0, i_10_467_4130_0,
    i_10_467_4154_0, i_10_467_4171_0, i_10_467_4268_0, i_10_467_4288_0,
    i_10_467_4379_0, i_10_467_4550_0, i_10_467_4565_0, i_10_467_4568_0;
  output o_10_467_0_0;
  assign o_10_467_0_0 = 0;
endmodule



// Benchmark "kernel_10_468" written by ABC on Sun Jul 19 10:29:13 2020

module kernel_10_468 ( 
    i_10_468_89_0, i_10_468_171_0, i_10_468_176_0, i_10_468_224_0,
    i_10_468_277_0, i_10_468_281_0, i_10_468_409_0, i_10_468_443_0,
    i_10_468_446_0, i_10_468_459_0, i_10_468_507_0, i_10_468_796_0,
    i_10_468_797_0, i_10_468_955_0, i_10_468_1034_0, i_10_468_1236_0,
    i_10_468_1244_0, i_10_468_1247_0, i_10_468_1248_0, i_10_468_1250_0,
    i_10_468_1343_0, i_10_468_1445_0, i_10_468_1540_0, i_10_468_1544_0,
    i_10_468_1554_0, i_10_468_1577_0, i_10_468_1580_0, i_10_468_1650_0,
    i_10_468_1678_0, i_10_468_1686_0, i_10_468_1688_0, i_10_468_1821_0,
    i_10_468_1822_0, i_10_468_1823_0, i_10_468_2197_0, i_10_468_2201_0,
    i_10_468_2407_0, i_10_468_2410_0, i_10_468_2452_0, i_10_468_2453_0,
    i_10_468_2469_0, i_10_468_2470_0, i_10_468_2472_0, i_10_468_2473_0,
    i_10_468_2474_0, i_10_468_2513_0, i_10_468_2530_0, i_10_468_2656_0,
    i_10_468_2657_0, i_10_468_2659_0, i_10_468_2660_0, i_10_468_2718_0,
    i_10_468_2719_0, i_10_468_2732_0, i_10_468_2828_0, i_10_468_2830_0,
    i_10_468_2831_0, i_10_468_2834_0, i_10_468_2863_0, i_10_468_2920_0,
    i_10_468_2921_0, i_10_468_2923_0, i_10_468_2979_0, i_10_468_3034_0,
    i_10_468_3070_0, i_10_468_3071_0, i_10_468_3198_0, i_10_468_3199_0,
    i_10_468_3200_0, i_10_468_3269_0, i_10_468_3284_0, i_10_468_3321_0,
    i_10_468_3324_0, i_10_468_3325_0, i_10_468_3329_0, i_10_468_3387_0,
    i_10_468_3409_0, i_10_468_3496_0, i_10_468_3497_0, i_10_468_3585_0,
    i_10_468_3586_0, i_10_468_3613_0, i_10_468_3614_0, i_10_468_3650_0,
    i_10_468_3780_0, i_10_468_3781_0, i_10_468_3782_0, i_10_468_3847_0,
    i_10_468_3848_0, i_10_468_3852_0, i_10_468_3853_0, i_10_468_3856_0,
    i_10_468_3992_0, i_10_468_4113_0, i_10_468_4121_0, i_10_468_4266_0,
    i_10_468_4267_0, i_10_468_4270_0, i_10_468_4279_0, i_10_468_4280_0,
    o_10_468_0_0  );
  input  i_10_468_89_0, i_10_468_171_0, i_10_468_176_0, i_10_468_224_0,
    i_10_468_277_0, i_10_468_281_0, i_10_468_409_0, i_10_468_443_0,
    i_10_468_446_0, i_10_468_459_0, i_10_468_507_0, i_10_468_796_0,
    i_10_468_797_0, i_10_468_955_0, i_10_468_1034_0, i_10_468_1236_0,
    i_10_468_1244_0, i_10_468_1247_0, i_10_468_1248_0, i_10_468_1250_0,
    i_10_468_1343_0, i_10_468_1445_0, i_10_468_1540_0, i_10_468_1544_0,
    i_10_468_1554_0, i_10_468_1577_0, i_10_468_1580_0, i_10_468_1650_0,
    i_10_468_1678_0, i_10_468_1686_0, i_10_468_1688_0, i_10_468_1821_0,
    i_10_468_1822_0, i_10_468_1823_0, i_10_468_2197_0, i_10_468_2201_0,
    i_10_468_2407_0, i_10_468_2410_0, i_10_468_2452_0, i_10_468_2453_0,
    i_10_468_2469_0, i_10_468_2470_0, i_10_468_2472_0, i_10_468_2473_0,
    i_10_468_2474_0, i_10_468_2513_0, i_10_468_2530_0, i_10_468_2656_0,
    i_10_468_2657_0, i_10_468_2659_0, i_10_468_2660_0, i_10_468_2718_0,
    i_10_468_2719_0, i_10_468_2732_0, i_10_468_2828_0, i_10_468_2830_0,
    i_10_468_2831_0, i_10_468_2834_0, i_10_468_2863_0, i_10_468_2920_0,
    i_10_468_2921_0, i_10_468_2923_0, i_10_468_2979_0, i_10_468_3034_0,
    i_10_468_3070_0, i_10_468_3071_0, i_10_468_3198_0, i_10_468_3199_0,
    i_10_468_3200_0, i_10_468_3269_0, i_10_468_3284_0, i_10_468_3321_0,
    i_10_468_3324_0, i_10_468_3325_0, i_10_468_3329_0, i_10_468_3387_0,
    i_10_468_3409_0, i_10_468_3496_0, i_10_468_3497_0, i_10_468_3585_0,
    i_10_468_3586_0, i_10_468_3613_0, i_10_468_3614_0, i_10_468_3650_0,
    i_10_468_3780_0, i_10_468_3781_0, i_10_468_3782_0, i_10_468_3847_0,
    i_10_468_3848_0, i_10_468_3852_0, i_10_468_3853_0, i_10_468_3856_0,
    i_10_468_3992_0, i_10_468_4113_0, i_10_468_4121_0, i_10_468_4266_0,
    i_10_468_4267_0, i_10_468_4270_0, i_10_468_4279_0, i_10_468_4280_0;
  output o_10_468_0_0;
  assign o_10_468_0_0 = ~((~i_10_468_1544_0 & ((~i_10_468_171_0 & ((i_10_468_796_0 & ~i_10_468_1821_0 & i_10_468_3852_0 & i_10_468_3853_0) | (~i_10_468_281_0 & ~i_10_468_797_0 & ~i_10_468_1034_0 & ~i_10_468_1580_0 & ~i_10_468_3034_0 & ~i_10_468_3198_0 & ~i_10_468_3200_0 & ~i_10_468_4280_0))) | (~i_10_468_1244_0 & ((~i_10_468_459_0 & ~i_10_468_1250_0 & ~i_10_468_1577_0 & ~i_10_468_2921_0 & i_10_468_3852_0) | (~i_10_468_1343_0 & ~i_10_468_1540_0 & ~i_10_468_1580_0 & ~i_10_468_1821_0 & ~i_10_468_1823_0 & ~i_10_468_2201_0 & ~i_10_468_2452_0 & ~i_10_468_2732_0 & ~i_10_468_3586_0 & ~i_10_468_3852_0 & ~i_10_468_3992_0 & ~i_10_468_4270_0))) | (~i_10_468_1248_0 & ((~i_10_468_1250_0 & i_10_468_2830_0 & ~i_10_468_3614_0 & ~i_10_468_3781_0 & ~i_10_468_4266_0) | (~i_10_468_446_0 & ~i_10_468_797_0 & ~i_10_468_1821_0 & ~i_10_468_1822_0 & ~i_10_468_3848_0 & ~i_10_468_4267_0))) | (~i_10_468_3614_0 & ~i_10_468_3853_0 & ((~i_10_468_409_0 & i_10_468_2474_0 & ~i_10_468_3071_0 & i_10_468_3284_0 & ~i_10_468_3387_0) | (~i_10_468_89_0 & ~i_10_468_1577_0 & i_10_468_1686_0 & ~i_10_468_2921_0 & ~i_10_468_3992_0 & ~i_10_468_4270_0 & ~i_10_468_3034_0 & ~i_10_468_3070_0))))) | (~i_10_468_89_0 & ((i_10_468_171_0 & ~i_10_468_443_0 & ~i_10_468_955_0 & ~i_10_468_3071_0 & ~i_10_468_3200_0 & ~i_10_468_3847_0 & ~i_10_468_4270_0) | (i_10_468_796_0 & i_10_468_797_0 & ~i_10_468_1236_0 & ~i_10_468_1247_0 & ~i_10_468_1343_0 & ~i_10_468_2201_0 & i_10_468_2453_0 & i_10_468_3613_0 & ~i_10_468_4113_0 & ~i_10_468_4279_0))) | (~i_10_468_3614_0 & ((~i_10_468_955_0 & ((~i_10_468_459_0 & ~i_10_468_1244_0 & ~i_10_468_1688_0 & ~i_10_468_2452_0 & ~i_10_468_3200_0 & ~i_10_468_3284_0 & ~i_10_468_3847_0 & ~i_10_468_3992_0) | (~i_10_468_796_0 & ~i_10_468_2201_0 & ~i_10_468_2453_0 & ~i_10_468_3070_0 & ~i_10_468_3650_0 & ~i_10_468_3848_0 & ~i_10_468_4266_0))) | (~i_10_468_2453_0 & ~i_10_468_2719_0 & ~i_10_468_2920_0 & i_10_468_3269_0 & ~i_10_468_3782_0) | (~i_10_468_224_0 & ~i_10_468_281_0 & ~i_10_468_1034_0 & ~i_10_468_1686_0 & ~i_10_468_1823_0 & ~i_10_468_3847_0 & ~i_10_468_4279_0))) | (~i_10_468_224_0 & ((~i_10_468_1248_0 & ~i_10_468_1250_0 & ~i_10_468_1540_0 & i_10_468_3852_0 & i_10_468_3853_0 & ~i_10_468_1577_0 & ~i_10_468_3848_0) | (~i_10_468_409_0 & ~i_10_468_1244_0 & ~i_10_468_1822_0 & ~i_10_468_1823_0 & ~i_10_468_2453_0 & ~i_10_468_3070_0 & ~i_10_468_3409_0 & ~i_10_468_3847_0 & ~i_10_468_4280_0))) | (~i_10_468_281_0 & ((i_10_468_1821_0 & i_10_468_1822_0 & ~i_10_468_2197_0 & ~i_10_468_2921_0 & ~i_10_468_3034_0 & ~i_10_468_3387_0 & ~i_10_468_3650_0 & ~i_10_468_4121_0) | (~i_10_468_443_0 & ~i_10_468_1034_0 & ~i_10_468_1250_0 & ~i_10_468_1540_0 & ~i_10_468_1688_0 & ~i_10_468_2452_0 & ~i_10_468_2453_0 & ~i_10_468_2920_0 & ~i_10_468_2923_0 & ~i_10_468_3070_0 & ~i_10_468_3853_0 & ~i_10_468_4270_0))) | (~i_10_468_1577_0 & ((~i_10_468_443_0 & ((~i_10_468_1244_0 & ~i_10_468_1540_0 & ~i_10_468_1580_0 & ~i_10_468_3071_0 & ~i_10_468_3200_0 & ~i_10_468_1650_0 & ~i_10_468_1823_0) | (~i_10_468_1822_0 & ~i_10_468_2197_0 & i_10_468_2732_0 & ~i_10_468_3199_0 & ~i_10_468_3782_0))) | (~i_10_468_2201_0 & ~i_10_468_2452_0 & ~i_10_468_3034_0 & ~i_10_468_3198_0 & ~i_10_468_3200_0 & ~i_10_468_3585_0 & ~i_10_468_3586_0 & i_10_468_3847_0 & ~i_10_468_3992_0 & ~i_10_468_4266_0))) | (~i_10_468_796_0 & ((~i_10_468_1540_0 & ~i_10_468_1688_0 & ~i_10_468_1821_0 & ~i_10_468_2453_0 & ~i_10_468_2719_0 & ~i_10_468_2831_0 & ~i_10_468_2921_0 & ~i_10_468_3071_0 & ~i_10_468_3992_0 & ~i_10_468_4113_0 & ~i_10_468_4121_0) | (~i_10_468_176_0 & i_10_468_1822_0 & ~i_10_468_1823_0 & ~i_10_468_3199_0 & ~i_10_468_3650_0 & ~i_10_468_4267_0 & ~i_10_468_4279_0))) | (~i_10_468_3848_0 & ((~i_10_468_176_0 & ((~i_10_468_1580_0 & i_10_468_2831_0 & ~i_10_468_2921_0 & ~i_10_468_3782_0) | (~i_10_468_1244_0 & ~i_10_468_1250_0 & ~i_10_468_2452_0 & ~i_10_468_2473_0 & ~i_10_468_3199_0 & ~i_10_468_3780_0 & ~i_10_468_3847_0 & ~i_10_468_3852_0 & ~i_10_468_3853_0))) | (~i_10_468_1686_0 & i_10_468_4113_0 & i_10_468_4266_0))) | (~i_10_468_1034_0 & ~i_10_468_1540_0 & ((~i_10_468_1823_0 & i_10_468_2831_0 & ~i_10_468_2923_0) | (i_10_468_2659_0 & ~i_10_468_3071_0 & ~i_10_468_4280_0))) | (~i_10_468_1247_0 & ((i_10_468_2656_0 & ~i_10_468_3269_0) | (~i_10_468_1580_0 & ~i_10_468_2201_0 & ~i_10_468_3070_0 & ~i_10_468_3071_0 & ~i_10_468_3847_0 & i_10_468_3853_0 & ~i_10_468_3992_0))) | (i_10_468_2979_0 & ((~i_10_468_3269_0 & ~i_10_468_3992_0 & ~i_10_468_4121_0) | (~i_10_468_3034_0 & i_10_468_4270_0))) | (~i_10_468_4121_0 & ((i_10_468_2469_0 & ~i_10_468_2921_0 & ~i_10_468_3782_0) | (i_10_468_2921_0 & ~i_10_468_3847_0 & ~i_10_468_3853_0 & i_10_468_4266_0 & i_10_468_4270_0))) | (~i_10_468_797_0 & ~i_10_468_1580_0 & i_10_468_2718_0 & i_10_468_3387_0) | (~i_10_468_3070_0 & i_10_468_3585_0 & i_10_468_3586_0 & ~i_10_468_3992_0) | (i_10_468_2473_0 & ~i_10_468_2828_0 & ~i_10_468_3613_0 & ~i_10_468_4267_0) | (~i_10_468_1823_0 & ~i_10_468_2732_0 & ~i_10_468_2920_0 & i_10_468_4279_0 & ~i_10_468_4280_0));
endmodule



// Benchmark "kernel_10_469" written by ABC on Sun Jul 19 10:29:14 2020

module kernel_10_469 ( 
    i_10_469_32_0, i_10_469_50_0, i_10_469_52_0, i_10_469_53_0,
    i_10_469_121_0, i_10_469_132_0, i_10_469_146_0, i_10_469_148_0,
    i_10_469_149_0, i_10_469_175_0, i_10_469_224_0, i_10_469_259_0,
    i_10_469_260_0, i_10_469_262_0, i_10_469_393_0, i_10_469_426_0,
    i_10_469_427_0, i_10_469_433_0, i_10_469_443_0, i_10_469_463_0,
    i_10_469_464_0, i_10_469_466_0, i_10_469_745_0, i_10_469_751_0,
    i_10_469_752_0, i_10_469_983_0, i_10_469_1050_0, i_10_469_1237_0,
    i_10_469_1238_0, i_10_469_1240_0, i_10_469_1241_0, i_10_469_1247_0,
    i_10_469_1312_0, i_10_469_1313_0, i_10_469_1534_0, i_10_469_1541_0,
    i_10_469_1544_0, i_10_469_1576_0, i_10_469_1624_0, i_10_469_1634_0,
    i_10_469_1640_0, i_10_469_1643_0, i_10_469_1683_0, i_10_469_1684_0,
    i_10_469_1689_0, i_10_469_1764_0, i_10_469_1819_0, i_10_469_1820_0,
    i_10_469_1957_0, i_10_469_1981_0, i_10_469_2029_0, i_10_469_2436_0,
    i_10_469_2471_0, i_10_469_2511_0, i_10_469_2607_0, i_10_469_2663_0,
    i_10_469_2697_0, i_10_469_2703_0, i_10_469_2704_0, i_10_469_2705_0,
    i_10_469_2707_0, i_10_469_2708_0, i_10_469_2731_0, i_10_469_2821_0,
    i_10_469_2829_0, i_10_469_2831_0, i_10_469_2842_0, i_10_469_2887_0,
    i_10_469_2913_0, i_10_469_2980_0, i_10_469_3045_0, i_10_469_3093_0,
    i_10_469_3130_0, i_10_469_3200_0, i_10_469_3281_0, i_10_469_3308_0,
    i_10_469_3385_0, i_10_469_3414_0, i_10_469_3470_0, i_10_469_3471_0,
    i_10_469_3494_0, i_10_469_3505_0, i_10_469_3587_0, i_10_469_3590_0,
    i_10_469_3611_0, i_10_469_3622_0, i_10_469_3836_0, i_10_469_3855_0,
    i_10_469_3858_0, i_10_469_3860_0, i_10_469_3946_0, i_10_469_3947_0,
    i_10_469_3981_0, i_10_469_4171_0, i_10_469_4204_0, i_10_469_4266_0,
    i_10_469_4267_0, i_10_469_4395_0, i_10_469_4396_0, i_10_469_4582_0,
    o_10_469_0_0  );
  input  i_10_469_32_0, i_10_469_50_0, i_10_469_52_0, i_10_469_53_0,
    i_10_469_121_0, i_10_469_132_0, i_10_469_146_0, i_10_469_148_0,
    i_10_469_149_0, i_10_469_175_0, i_10_469_224_0, i_10_469_259_0,
    i_10_469_260_0, i_10_469_262_0, i_10_469_393_0, i_10_469_426_0,
    i_10_469_427_0, i_10_469_433_0, i_10_469_443_0, i_10_469_463_0,
    i_10_469_464_0, i_10_469_466_0, i_10_469_745_0, i_10_469_751_0,
    i_10_469_752_0, i_10_469_983_0, i_10_469_1050_0, i_10_469_1237_0,
    i_10_469_1238_0, i_10_469_1240_0, i_10_469_1241_0, i_10_469_1247_0,
    i_10_469_1312_0, i_10_469_1313_0, i_10_469_1534_0, i_10_469_1541_0,
    i_10_469_1544_0, i_10_469_1576_0, i_10_469_1624_0, i_10_469_1634_0,
    i_10_469_1640_0, i_10_469_1643_0, i_10_469_1683_0, i_10_469_1684_0,
    i_10_469_1689_0, i_10_469_1764_0, i_10_469_1819_0, i_10_469_1820_0,
    i_10_469_1957_0, i_10_469_1981_0, i_10_469_2029_0, i_10_469_2436_0,
    i_10_469_2471_0, i_10_469_2511_0, i_10_469_2607_0, i_10_469_2663_0,
    i_10_469_2697_0, i_10_469_2703_0, i_10_469_2704_0, i_10_469_2705_0,
    i_10_469_2707_0, i_10_469_2708_0, i_10_469_2731_0, i_10_469_2821_0,
    i_10_469_2829_0, i_10_469_2831_0, i_10_469_2842_0, i_10_469_2887_0,
    i_10_469_2913_0, i_10_469_2980_0, i_10_469_3045_0, i_10_469_3093_0,
    i_10_469_3130_0, i_10_469_3200_0, i_10_469_3281_0, i_10_469_3308_0,
    i_10_469_3385_0, i_10_469_3414_0, i_10_469_3470_0, i_10_469_3471_0,
    i_10_469_3494_0, i_10_469_3505_0, i_10_469_3587_0, i_10_469_3590_0,
    i_10_469_3611_0, i_10_469_3622_0, i_10_469_3836_0, i_10_469_3855_0,
    i_10_469_3858_0, i_10_469_3860_0, i_10_469_3946_0, i_10_469_3947_0,
    i_10_469_3981_0, i_10_469_4171_0, i_10_469_4204_0, i_10_469_4266_0,
    i_10_469_4267_0, i_10_469_4395_0, i_10_469_4396_0, i_10_469_4582_0;
  output o_10_469_0_0;
  assign o_10_469_0_0 = 0;
endmodule



// Benchmark "kernel_10_470" written by ABC on Sun Jul 19 10:29:15 2020

module kernel_10_470 ( 
    i_10_470_221_0, i_10_470_245_0, i_10_470_273_0, i_10_470_320_0,
    i_10_470_329_0, i_10_470_388_0, i_10_470_409_0, i_10_470_432_0,
    i_10_470_433_0, i_10_470_434_0, i_10_470_441_0, i_10_470_443_0,
    i_10_470_444_0, i_10_470_445_0, i_10_470_446_0, i_10_470_459_0,
    i_10_470_463_0, i_10_470_464_0, i_10_470_512_0, i_10_470_713_0,
    i_10_470_875_0, i_10_470_959_0, i_10_470_990_0, i_10_470_991_0,
    i_10_470_992_0, i_10_470_1198_0, i_10_470_1238_0, i_10_470_1265_0,
    i_10_470_1309_0, i_10_470_1313_0, i_10_470_1654_0, i_10_470_1683_0,
    i_10_470_1687_0, i_10_470_1688_0, i_10_470_1819_0, i_10_470_1820_0,
    i_10_470_1821_0, i_10_470_1826_0, i_10_470_1874_0, i_10_470_1990_0,
    i_10_470_1991_0, i_10_470_2018_0, i_10_470_2021_0, i_10_470_2198_0,
    i_10_470_2261_0, i_10_470_2264_0, i_10_470_2353_0, i_10_470_2354_0,
    i_10_470_2359_0, i_10_470_2362_0, i_10_470_2366_0, i_10_470_2377_0,
    i_10_470_2378_0, i_10_470_2381_0, i_10_470_2459_0, i_10_470_2467_0,
    i_10_470_2468_0, i_10_470_2628_0, i_10_470_2660_0, i_10_470_2675_0,
    i_10_470_2720_0, i_10_470_2729_0, i_10_470_2789_0, i_10_470_2826_0,
    i_10_470_2829_0, i_10_470_2830_0, i_10_470_2831_0, i_10_470_2918_0,
    i_10_470_2979_0, i_10_470_3070_0, i_10_470_3076_0, i_10_470_3151_0,
    i_10_470_3155_0, i_10_470_3156_0, i_10_470_3280_0, i_10_470_3281_0,
    i_10_470_3388_0, i_10_470_3389_0, i_10_470_3392_0, i_10_470_3466_0,
    i_10_470_3551_0, i_10_470_3611_0, i_10_470_3612_0, i_10_470_3614_0,
    i_10_470_3785_0, i_10_470_3834_0, i_10_470_3835_0, i_10_470_3838_0,
    i_10_470_3856_0, i_10_470_3978_0, i_10_470_3983_0, i_10_470_4027_0,
    i_10_470_4115_0, i_10_470_4116_0, i_10_470_4126_0, i_10_470_4214_0,
    i_10_470_4268_0, i_10_470_4279_0, i_10_470_4285_0, i_10_470_4291_0,
    o_10_470_0_0  );
  input  i_10_470_221_0, i_10_470_245_0, i_10_470_273_0, i_10_470_320_0,
    i_10_470_329_0, i_10_470_388_0, i_10_470_409_0, i_10_470_432_0,
    i_10_470_433_0, i_10_470_434_0, i_10_470_441_0, i_10_470_443_0,
    i_10_470_444_0, i_10_470_445_0, i_10_470_446_0, i_10_470_459_0,
    i_10_470_463_0, i_10_470_464_0, i_10_470_512_0, i_10_470_713_0,
    i_10_470_875_0, i_10_470_959_0, i_10_470_990_0, i_10_470_991_0,
    i_10_470_992_0, i_10_470_1198_0, i_10_470_1238_0, i_10_470_1265_0,
    i_10_470_1309_0, i_10_470_1313_0, i_10_470_1654_0, i_10_470_1683_0,
    i_10_470_1687_0, i_10_470_1688_0, i_10_470_1819_0, i_10_470_1820_0,
    i_10_470_1821_0, i_10_470_1826_0, i_10_470_1874_0, i_10_470_1990_0,
    i_10_470_1991_0, i_10_470_2018_0, i_10_470_2021_0, i_10_470_2198_0,
    i_10_470_2261_0, i_10_470_2264_0, i_10_470_2353_0, i_10_470_2354_0,
    i_10_470_2359_0, i_10_470_2362_0, i_10_470_2366_0, i_10_470_2377_0,
    i_10_470_2378_0, i_10_470_2381_0, i_10_470_2459_0, i_10_470_2467_0,
    i_10_470_2468_0, i_10_470_2628_0, i_10_470_2660_0, i_10_470_2675_0,
    i_10_470_2720_0, i_10_470_2729_0, i_10_470_2789_0, i_10_470_2826_0,
    i_10_470_2829_0, i_10_470_2830_0, i_10_470_2831_0, i_10_470_2918_0,
    i_10_470_2979_0, i_10_470_3070_0, i_10_470_3076_0, i_10_470_3151_0,
    i_10_470_3155_0, i_10_470_3156_0, i_10_470_3280_0, i_10_470_3281_0,
    i_10_470_3388_0, i_10_470_3389_0, i_10_470_3392_0, i_10_470_3466_0,
    i_10_470_3551_0, i_10_470_3611_0, i_10_470_3612_0, i_10_470_3614_0,
    i_10_470_3785_0, i_10_470_3834_0, i_10_470_3835_0, i_10_470_3838_0,
    i_10_470_3856_0, i_10_470_3978_0, i_10_470_3983_0, i_10_470_4027_0,
    i_10_470_4115_0, i_10_470_4116_0, i_10_470_4126_0, i_10_470_4214_0,
    i_10_470_4268_0, i_10_470_4279_0, i_10_470_4285_0, i_10_470_4291_0;
  output o_10_470_0_0;
  assign o_10_470_0_0 = ~((~i_10_470_329_0 & ((~i_10_470_320_0 & ((~i_10_470_433_0 & ~i_10_470_2353_0 & i_10_470_2359_0 & ~i_10_470_2378_0 & ~i_10_470_2789_0 & ~i_10_470_3612_0 & ~i_10_470_3614_0 & ~i_10_470_3785_0 & ~i_10_470_3835_0) | (~i_10_470_1309_0 & ~i_10_470_2359_0 & ~i_10_470_2377_0 & ~i_10_470_4279_0))) | (~i_10_470_991_0 & ~i_10_470_1265_0 & ~i_10_470_2675_0 & ~i_10_470_2720_0 & ~i_10_470_2729_0 & ~i_10_470_2979_0 & ~i_10_470_4027_0) | (~i_10_470_1826_0 & ~i_10_470_3856_0 & ~i_10_470_4126_0 & i_10_470_4291_0))) | (~i_10_470_434_0 & ((~i_10_470_992_0 & ~i_10_470_2353_0 & ~i_10_470_2377_0 & ~i_10_470_2459_0 & ~i_10_470_2660_0 & ~i_10_470_2789_0) | (~i_10_470_1819_0 & ~i_10_470_2021_0 & ~i_10_470_2830_0 & ~i_10_470_2831_0 & ~i_10_470_2918_0 & ~i_10_470_3281_0 & ~i_10_470_4268_0))) | (~i_10_470_4285_0 & ((i_10_470_463_0 & ((~i_10_470_991_0 & ~i_10_470_4115_0) | (i_10_470_1654_0 & ~i_10_470_3076_0 & i_10_470_4116_0))) | (~i_10_470_433_0 & ~i_10_470_446_0 & ~i_10_470_2354_0 & ~i_10_470_2459_0 & ~i_10_470_2675_0 & ~i_10_470_2826_0 & ~i_10_470_3070_0 & ~i_10_470_3838_0))) | (~i_10_470_2018_0 & ((~i_10_470_433_0 & ~i_10_470_3551_0 & ((~i_10_470_409_0 & ~i_10_470_2366_0 & ~i_10_470_2918_0 & ~i_10_470_3611_0 & ~i_10_470_4027_0) | (~i_10_470_1313_0 & ~i_10_470_2354_0 & ~i_10_470_2378_0 & ~i_10_470_2459_0 & ~i_10_470_2789_0 & ~i_10_470_3076_0 & ~i_10_470_4126_0))) | (~i_10_470_2021_0 & ~i_10_470_2353_0 & ~i_10_470_2377_0 & ~i_10_470_2381_0 & ~i_10_470_3388_0) | (~i_10_470_2359_0 & ~i_10_470_2366_0 & ~i_10_470_2675_0 & ~i_10_470_3392_0 & i_10_470_3834_0))) | (~i_10_470_1265_0 & ((~i_10_470_409_0 & ((~i_10_470_2366_0 & ~i_10_470_2826_0 & ~i_10_470_2829_0 & ~i_10_470_2830_0 & ~i_10_470_2831_0) | (~i_10_470_1874_0 & ~i_10_470_2377_0 & ~i_10_470_2378_0 & ~i_10_470_2459_0 & ~i_10_470_2789_0 & i_10_470_3389_0 & ~i_10_470_3785_0))) | (~i_10_470_1238_0 & i_10_470_1821_0 & ~i_10_470_1990_0 & ~i_10_470_2198_0 & ~i_10_470_2459_0) | (~i_10_470_992_0 & i_10_470_1820_0 & ~i_10_470_2826_0 & ~i_10_470_2918_0) | (i_10_470_1313_0 & i_10_470_2362_0 & i_10_470_3392_0 & i_10_470_3856_0))) | (~i_10_470_991_0 & ((~i_10_470_990_0 & ~i_10_470_1991_0 & ~i_10_470_2354_0 & ~i_10_470_2826_0 & ~i_10_470_3076_0 & ~i_10_470_3389_0) | (~i_10_470_432_0 & ~i_10_470_992_0 & ~i_10_470_2918_0 & i_10_470_3835_0 & ~i_10_470_3856_0))) | (~i_10_470_432_0 & ~i_10_470_1991_0 & ((i_10_470_2021_0 & ~i_10_470_2789_0 & ~i_10_470_2826_0 & i_10_470_4116_0) | (~i_10_470_992_0 & ~i_10_470_1309_0 & ~i_10_470_2381_0 & ~i_10_470_2459_0 & ~i_10_470_2660_0 & ~i_10_470_3281_0 & ~i_10_470_3785_0 & ~i_10_470_3978_0 & ~i_10_470_4291_0))) | (i_10_470_4116_0 & ((i_10_470_3280_0 & ~i_10_470_3983_0) | (i_10_470_3856_0 & ~i_10_470_4115_0 & i_10_470_4279_0))) | (~i_10_470_1238_0 & ~i_10_470_2378_0 & i_10_470_2459_0 & ~i_10_470_2660_0 & i_10_470_2720_0 & ~i_10_470_3281_0 & ~i_10_470_4116_0));
endmodule



// Benchmark "kernel_10_471" written by ABC on Sun Jul 19 10:29:17 2020

module kernel_10_471 ( 
    i_10_471_149_0, i_10_471_172_0, i_10_471_173_0, i_10_471_176_0,
    i_10_471_178_0, i_10_471_250_0, i_10_471_323_0, i_10_471_425_0,
    i_10_471_428_0, i_10_471_429_0, i_10_471_430_0, i_10_471_431_0,
    i_10_471_466_0, i_10_471_467_0, i_10_471_504_0, i_10_471_505_0,
    i_10_471_507_0, i_10_471_508_0, i_10_471_715_0, i_10_471_716_0,
    i_10_471_718_0, i_10_471_794_0, i_10_471_896_0, i_10_471_965_0,
    i_10_471_1233_0, i_10_471_1305_0, i_10_471_1308_0, i_10_471_1310_0,
    i_10_471_1312_0, i_10_471_1313_0, i_10_471_1546_0, i_10_471_1631_0,
    i_10_471_1651_0, i_10_471_1652_0, i_10_471_1654_0, i_10_471_1655_0,
    i_10_471_1684_0, i_10_471_1685_0, i_10_471_1687_0, i_10_471_1768_0,
    i_10_471_1991_0, i_10_471_1994_0, i_10_471_2000_0, i_10_471_2255_0,
    i_10_471_2349_0, i_10_471_2354_0, i_10_471_2357_0, i_10_471_2404_0,
    i_10_471_2450_0, i_10_471_2453_0, i_10_471_2567_0, i_10_471_2570_0,
    i_10_471_2572_0, i_10_471_2628_0, i_10_471_2675_0, i_10_471_2703_0,
    i_10_471_2710_0, i_10_471_2711_0, i_10_471_2714_0, i_10_471_2716_0,
    i_10_471_2717_0, i_10_471_2883_0, i_10_471_3036_0, i_10_471_3037_0,
    i_10_471_3038_0, i_10_471_3072_0, i_10_471_3269_0, i_10_471_3322_0,
    i_10_471_3384_0, i_10_471_3385_0, i_10_471_3386_0, i_10_471_3388_0,
    i_10_471_3389_0, i_10_471_3391_0, i_10_471_3392_0, i_10_471_3404_0,
    i_10_471_3406_0, i_10_471_3410_0, i_10_471_3524_0, i_10_471_3527_0,
    i_10_471_3583_0, i_10_471_3589_0, i_10_471_3650_0, i_10_471_3652_0,
    i_10_471_3684_0, i_10_471_3837_0, i_10_471_3846_0, i_10_471_3847_0,
    i_10_471_3848_0, i_10_471_3857_0, i_10_471_3872_0, i_10_471_3947_0,
    i_10_471_4027_0, i_10_471_4028_0, i_10_471_4123_0, i_10_471_4285_0,
    i_10_471_4286_0, i_10_471_4288_0, i_10_471_4289_0, i_10_471_4291_0,
    o_10_471_0_0  );
  input  i_10_471_149_0, i_10_471_172_0, i_10_471_173_0, i_10_471_176_0,
    i_10_471_178_0, i_10_471_250_0, i_10_471_323_0, i_10_471_425_0,
    i_10_471_428_0, i_10_471_429_0, i_10_471_430_0, i_10_471_431_0,
    i_10_471_466_0, i_10_471_467_0, i_10_471_504_0, i_10_471_505_0,
    i_10_471_507_0, i_10_471_508_0, i_10_471_715_0, i_10_471_716_0,
    i_10_471_718_0, i_10_471_794_0, i_10_471_896_0, i_10_471_965_0,
    i_10_471_1233_0, i_10_471_1305_0, i_10_471_1308_0, i_10_471_1310_0,
    i_10_471_1312_0, i_10_471_1313_0, i_10_471_1546_0, i_10_471_1631_0,
    i_10_471_1651_0, i_10_471_1652_0, i_10_471_1654_0, i_10_471_1655_0,
    i_10_471_1684_0, i_10_471_1685_0, i_10_471_1687_0, i_10_471_1768_0,
    i_10_471_1991_0, i_10_471_1994_0, i_10_471_2000_0, i_10_471_2255_0,
    i_10_471_2349_0, i_10_471_2354_0, i_10_471_2357_0, i_10_471_2404_0,
    i_10_471_2450_0, i_10_471_2453_0, i_10_471_2567_0, i_10_471_2570_0,
    i_10_471_2572_0, i_10_471_2628_0, i_10_471_2675_0, i_10_471_2703_0,
    i_10_471_2710_0, i_10_471_2711_0, i_10_471_2714_0, i_10_471_2716_0,
    i_10_471_2717_0, i_10_471_2883_0, i_10_471_3036_0, i_10_471_3037_0,
    i_10_471_3038_0, i_10_471_3072_0, i_10_471_3269_0, i_10_471_3322_0,
    i_10_471_3384_0, i_10_471_3385_0, i_10_471_3386_0, i_10_471_3388_0,
    i_10_471_3389_0, i_10_471_3391_0, i_10_471_3392_0, i_10_471_3404_0,
    i_10_471_3406_0, i_10_471_3410_0, i_10_471_3524_0, i_10_471_3527_0,
    i_10_471_3583_0, i_10_471_3589_0, i_10_471_3650_0, i_10_471_3652_0,
    i_10_471_3684_0, i_10_471_3837_0, i_10_471_3846_0, i_10_471_3847_0,
    i_10_471_3848_0, i_10_471_3857_0, i_10_471_3872_0, i_10_471_3947_0,
    i_10_471_4027_0, i_10_471_4028_0, i_10_471_4123_0, i_10_471_4285_0,
    i_10_471_4286_0, i_10_471_4288_0, i_10_471_4289_0, i_10_471_4291_0;
  output o_10_471_0_0;
  assign o_10_471_0_0 = ~((~i_10_471_2450_0 & ((~i_10_471_425_0 & ((~i_10_471_250_0 & ~i_10_471_1685_0 & ~i_10_471_1994_0 & ~i_10_471_2354_0 & ~i_10_471_2453_0 & ~i_10_471_2567_0 & ~i_10_471_2716_0 & i_10_471_3846_0) | (~i_10_471_176_0 & ~i_10_471_431_0 & ~i_10_471_2570_0 & ~i_10_471_3072_0 & ~i_10_471_3391_0 & i_10_471_3837_0 & ~i_10_471_3847_0))) | (i_10_471_1651_0 & ~i_10_471_2703_0 & ~i_10_471_2716_0 & i_10_471_3847_0))) | (~i_10_471_176_0 & ((~i_10_471_323_0 & i_10_471_1308_0 & ~i_10_471_3386_0 & i_10_471_3589_0 & ~i_10_471_3848_0) | (~i_10_471_149_0 & ~i_10_471_429_0 & ~i_10_471_1233_0 & ~i_10_471_2349_0 & ~i_10_471_2567_0 & ~i_10_471_2570_0 & ~i_10_471_2572_0 & ~i_10_471_3038_0 & ~i_10_471_3404_0 & ~i_10_471_3410_0 & ~i_10_471_3524_0 & ~i_10_471_3652_0 & ~i_10_471_4123_0))) | (~i_10_471_965_0 & ((~i_10_471_323_0 & ~i_10_471_716_0 & i_10_471_1233_0 & ~i_10_471_1685_0 & ~i_10_471_2711_0) | (~i_10_471_428_0 & ~i_10_471_1994_0 & ~i_10_471_2000_0 & ~i_10_471_2357_0 & ~i_10_471_2570_0 & ~i_10_471_3388_0 & ~i_10_471_3389_0 & ~i_10_471_3410_0 & ~i_10_471_3847_0))) | (~i_10_471_3848_0 & ((~i_10_471_323_0 & ((~i_10_471_1994_0 & ~i_10_471_3410_0 & ~i_10_471_3583_0 & ~i_10_471_4027_0 & ~i_10_471_4289_0) | (~i_10_471_2714_0 & ~i_10_471_3857_0 & ~i_10_471_4028_0 & ~i_10_471_4291_0))) | (~i_10_471_431_0 & ~i_10_471_466_0 & ~i_10_471_2714_0 & i_10_471_2883_0))) | (~i_10_471_2711_0 & ((~i_10_471_428_0 & ~i_10_471_3837_0 & ((~i_10_471_467_0 & ~i_10_471_1685_0 & ~i_10_471_1768_0 & ~i_10_471_2716_0 & ~i_10_471_3583_0) | (~i_10_471_794_0 & ~i_10_471_1308_0 & ~i_10_471_1310_0 & ~i_10_471_1546_0 & ~i_10_471_3589_0 & ~i_10_471_4027_0))) | (~i_10_471_431_0 & ~i_10_471_2714_0 & ~i_10_471_3947_0 & ((~i_10_471_173_0 & ~i_10_471_430_0 & ~i_10_471_2567_0 & ~i_10_471_2572_0 & ~i_10_471_3404_0) | (~i_10_471_2710_0 & ~i_10_471_3392_0 & ~i_10_471_4291_0))))) | (~i_10_471_3392_0 & ((~i_10_471_428_0 & ((~i_10_471_429_0 & ~i_10_471_716_0 & i_10_471_1655_0 & ~i_10_471_1768_0 & ~i_10_471_2570_0 & ~i_10_471_2675_0 & ~i_10_471_3384_0) | (~i_10_471_467_0 & i_10_471_1651_0 & ~i_10_471_2710_0 & ~i_10_471_3589_0 & ~i_10_471_4289_0))) | (~i_10_471_716_0 & ~i_10_471_896_0 & i_10_471_1655_0 & ~i_10_471_2453_0 & ~i_10_471_2567_0 & ~i_10_471_2572_0 & ~i_10_471_4028_0) | (~i_10_471_718_0 & ~i_10_471_1652_0 & ~i_10_471_2349_0 & ~i_10_471_2570_0 & ~i_10_471_3386_0 & ~i_10_471_3410_0 & ~i_10_471_3524_0 & ~i_10_471_4286_0 & ~i_10_471_4288_0))) | (~i_10_471_718_0 & ((~i_10_471_2567_0 & ~i_10_471_2570_0 & ~i_10_471_2572_0 & ~i_10_471_3269_0 & ~i_10_471_3385_0 & ~i_10_471_3388_0 & ~i_10_471_3389_0 & ~i_10_471_3410_0 & ~i_10_471_3527_0 & ~i_10_471_3583_0) | (i_10_471_2404_0 & ~i_10_471_2717_0 & ~i_10_471_3947_0))) | (~i_10_471_467_0 & ~i_10_471_1687_0 & i_10_471_3036_0) | (~i_10_471_1991_0 & ~i_10_471_2000_0 & ~i_10_471_2714_0 & ~i_10_471_2716_0 & ~i_10_471_3391_0 & ~i_10_471_4123_0 & ~i_10_471_4289_0));
endmodule



// Benchmark "kernel_10_472" written by ABC on Sun Jul 19 10:29:18 2020

module kernel_10_472 ( 
    i_10_472_64_0, i_10_472_65_0, i_10_472_68_0, i_10_472_175_0,
    i_10_472_176_0, i_10_472_178_0, i_10_472_179_0, i_10_472_272_0,
    i_10_472_279_0, i_10_472_285_0, i_10_472_316_0, i_10_472_317_0,
    i_10_472_319_0, i_10_472_320_0, i_10_472_408_0, i_10_472_413_0,
    i_10_472_433_0, i_10_472_437_0, i_10_472_533_0, i_10_472_635_0,
    i_10_472_638_0, i_10_472_641_0, i_10_472_644_0, i_10_472_896_0,
    i_10_472_1055_0, i_10_472_1081_0, i_10_472_1233_0, i_10_472_1249_0,
    i_10_472_1298_0, i_10_472_1306_0, i_10_472_1307_0, i_10_472_1309_0,
    i_10_472_1364_0, i_10_472_1433_0, i_10_472_1436_0, i_10_472_1487_0,
    i_10_472_1622_0, i_10_472_1648_0, i_10_472_1651_0, i_10_472_1652_0,
    i_10_472_1655_0, i_10_472_1685_0, i_10_472_1690_0, i_10_472_1768_0,
    i_10_472_1796_0, i_10_472_1874_0, i_10_472_2021_0, i_10_472_2024_0,
    i_10_472_2237_0, i_10_472_2264_0, i_10_472_2351_0, i_10_472_2356_0,
    i_10_472_2381_0, i_10_472_2453_0, i_10_472_2468_0, i_10_472_2470_0,
    i_10_472_2513_0, i_10_472_2519_0, i_10_472_2567_0, i_10_472_2629_0,
    i_10_472_2632_0, i_10_472_2633_0, i_10_472_2704_0, i_10_472_2711_0,
    i_10_472_2717_0, i_10_472_2735_0, i_10_472_2744_0, i_10_472_2831_0,
    i_10_472_2846_0, i_10_472_3044_0, i_10_472_3045_0, i_10_472_3071_0,
    i_10_472_3317_0, i_10_472_3384_0, i_10_472_3386_0, i_10_472_3388_0,
    i_10_472_3389_0, i_10_472_3467_0, i_10_472_3469_0, i_10_472_3470_0,
    i_10_472_3494_0, i_10_472_3539_0, i_10_472_3542_0, i_10_472_3557_0,
    i_10_472_3584_0, i_10_472_3586_0, i_10_472_3587_0, i_10_472_3647_0,
    i_10_472_3775_0, i_10_472_3794_0, i_10_472_3847_0, i_10_472_3848_0,
    i_10_472_3944_0, i_10_472_4114_0, i_10_472_4121_0, i_10_472_4167_0,
    i_10_472_4267_0, i_10_472_4276_0, i_10_472_4289_0, i_10_472_4586_0,
    o_10_472_0_0  );
  input  i_10_472_64_0, i_10_472_65_0, i_10_472_68_0, i_10_472_175_0,
    i_10_472_176_0, i_10_472_178_0, i_10_472_179_0, i_10_472_272_0,
    i_10_472_279_0, i_10_472_285_0, i_10_472_316_0, i_10_472_317_0,
    i_10_472_319_0, i_10_472_320_0, i_10_472_408_0, i_10_472_413_0,
    i_10_472_433_0, i_10_472_437_0, i_10_472_533_0, i_10_472_635_0,
    i_10_472_638_0, i_10_472_641_0, i_10_472_644_0, i_10_472_896_0,
    i_10_472_1055_0, i_10_472_1081_0, i_10_472_1233_0, i_10_472_1249_0,
    i_10_472_1298_0, i_10_472_1306_0, i_10_472_1307_0, i_10_472_1309_0,
    i_10_472_1364_0, i_10_472_1433_0, i_10_472_1436_0, i_10_472_1487_0,
    i_10_472_1622_0, i_10_472_1648_0, i_10_472_1651_0, i_10_472_1652_0,
    i_10_472_1655_0, i_10_472_1685_0, i_10_472_1690_0, i_10_472_1768_0,
    i_10_472_1796_0, i_10_472_1874_0, i_10_472_2021_0, i_10_472_2024_0,
    i_10_472_2237_0, i_10_472_2264_0, i_10_472_2351_0, i_10_472_2356_0,
    i_10_472_2381_0, i_10_472_2453_0, i_10_472_2468_0, i_10_472_2470_0,
    i_10_472_2513_0, i_10_472_2519_0, i_10_472_2567_0, i_10_472_2629_0,
    i_10_472_2632_0, i_10_472_2633_0, i_10_472_2704_0, i_10_472_2711_0,
    i_10_472_2717_0, i_10_472_2735_0, i_10_472_2744_0, i_10_472_2831_0,
    i_10_472_2846_0, i_10_472_3044_0, i_10_472_3045_0, i_10_472_3071_0,
    i_10_472_3317_0, i_10_472_3384_0, i_10_472_3386_0, i_10_472_3388_0,
    i_10_472_3389_0, i_10_472_3467_0, i_10_472_3469_0, i_10_472_3470_0,
    i_10_472_3494_0, i_10_472_3539_0, i_10_472_3542_0, i_10_472_3557_0,
    i_10_472_3584_0, i_10_472_3586_0, i_10_472_3587_0, i_10_472_3647_0,
    i_10_472_3775_0, i_10_472_3794_0, i_10_472_3847_0, i_10_472_3848_0,
    i_10_472_3944_0, i_10_472_4114_0, i_10_472_4121_0, i_10_472_4167_0,
    i_10_472_4267_0, i_10_472_4276_0, i_10_472_4289_0, i_10_472_4586_0;
  output o_10_472_0_0;
  assign o_10_472_0_0 = 0;
endmodule



// Benchmark "kernel_10_473" written by ABC on Sun Jul 19 10:29:18 2020

module kernel_10_473 ( 
    i_10_473_174_0, i_10_473_292_0, i_10_473_295_0, i_10_473_296_0,
    i_10_473_394_0, i_10_473_405_0, i_10_473_429_0, i_10_473_431_0,
    i_10_473_438_0, i_10_473_444_0, i_10_473_445_0, i_10_473_447_0,
    i_10_473_449_0, i_10_473_460_0, i_10_473_795_0, i_10_473_798_0,
    i_10_473_800_0, i_10_473_823_0, i_10_473_826_0, i_10_473_850_0,
    i_10_473_852_0, i_10_473_853_0, i_10_473_1033_0, i_10_473_1052_0,
    i_10_473_1202_0, i_10_473_1235_0, i_10_473_1236_0, i_10_473_1237_0,
    i_10_473_1238_0, i_10_473_1266_0, i_10_473_1309_0, i_10_473_1310_0,
    i_10_473_1342_0, i_10_473_1378_0, i_10_473_1435_0, i_10_473_1436_0,
    i_10_473_1553_0, i_10_473_1579_0, i_10_473_1580_0, i_10_473_1651_0,
    i_10_473_1652_0, i_10_473_1653_0, i_10_473_1680_0, i_10_473_1688_0,
    i_10_473_1823_0, i_10_473_1996_0, i_10_473_2084_0, i_10_473_2158_0,
    i_10_473_2184_0, i_10_473_2309_0, i_10_473_2310_0, i_10_473_2311_0,
    i_10_473_2337_0, i_10_473_2338_0, i_10_473_2351_0, i_10_473_2448_0,
    i_10_473_2450_0, i_10_473_2463_0, i_10_473_2470_0, i_10_473_2482_0,
    i_10_473_2532_0, i_10_473_2562_0, i_10_473_2632_0, i_10_473_2660_0,
    i_10_473_2662_0, i_10_473_2679_0, i_10_473_2697_0, i_10_473_2710_0,
    i_10_473_2718_0, i_10_473_2829_0, i_10_473_2830_0, i_10_473_2880_0,
    i_10_473_2918_0, i_10_473_2922_0, i_10_473_2950_0, i_10_473_3091_0,
    i_10_473_3095_0, i_10_473_3199_0, i_10_473_3278_0, i_10_473_3406_0,
    i_10_473_3539_0, i_10_473_3555_0, i_10_473_3562_0, i_10_473_3601_0,
    i_10_473_3602_0, i_10_473_3637_0, i_10_473_3782_0, i_10_473_3785_0,
    i_10_473_3832_0, i_10_473_3834_0, i_10_473_3840_0, i_10_473_3841_0,
    i_10_473_3853_0, i_10_473_3902_0, i_10_473_3979_0, i_10_473_3983_0,
    i_10_473_3995_0, i_10_473_4116_0, i_10_473_4117_0, i_10_473_4180_0,
    o_10_473_0_0  );
  input  i_10_473_174_0, i_10_473_292_0, i_10_473_295_0, i_10_473_296_0,
    i_10_473_394_0, i_10_473_405_0, i_10_473_429_0, i_10_473_431_0,
    i_10_473_438_0, i_10_473_444_0, i_10_473_445_0, i_10_473_447_0,
    i_10_473_449_0, i_10_473_460_0, i_10_473_795_0, i_10_473_798_0,
    i_10_473_800_0, i_10_473_823_0, i_10_473_826_0, i_10_473_850_0,
    i_10_473_852_0, i_10_473_853_0, i_10_473_1033_0, i_10_473_1052_0,
    i_10_473_1202_0, i_10_473_1235_0, i_10_473_1236_0, i_10_473_1237_0,
    i_10_473_1238_0, i_10_473_1266_0, i_10_473_1309_0, i_10_473_1310_0,
    i_10_473_1342_0, i_10_473_1378_0, i_10_473_1435_0, i_10_473_1436_0,
    i_10_473_1553_0, i_10_473_1579_0, i_10_473_1580_0, i_10_473_1651_0,
    i_10_473_1652_0, i_10_473_1653_0, i_10_473_1680_0, i_10_473_1688_0,
    i_10_473_1823_0, i_10_473_1996_0, i_10_473_2084_0, i_10_473_2158_0,
    i_10_473_2184_0, i_10_473_2309_0, i_10_473_2310_0, i_10_473_2311_0,
    i_10_473_2337_0, i_10_473_2338_0, i_10_473_2351_0, i_10_473_2448_0,
    i_10_473_2450_0, i_10_473_2463_0, i_10_473_2470_0, i_10_473_2482_0,
    i_10_473_2532_0, i_10_473_2562_0, i_10_473_2632_0, i_10_473_2660_0,
    i_10_473_2662_0, i_10_473_2679_0, i_10_473_2697_0, i_10_473_2710_0,
    i_10_473_2718_0, i_10_473_2829_0, i_10_473_2830_0, i_10_473_2880_0,
    i_10_473_2918_0, i_10_473_2922_0, i_10_473_2950_0, i_10_473_3091_0,
    i_10_473_3095_0, i_10_473_3199_0, i_10_473_3278_0, i_10_473_3406_0,
    i_10_473_3539_0, i_10_473_3555_0, i_10_473_3562_0, i_10_473_3601_0,
    i_10_473_3602_0, i_10_473_3637_0, i_10_473_3782_0, i_10_473_3785_0,
    i_10_473_3832_0, i_10_473_3834_0, i_10_473_3840_0, i_10_473_3841_0,
    i_10_473_3853_0, i_10_473_3902_0, i_10_473_3979_0, i_10_473_3983_0,
    i_10_473_3995_0, i_10_473_4116_0, i_10_473_4117_0, i_10_473_4180_0;
  output o_10_473_0_0;
  assign o_10_473_0_0 = 0;
endmodule



// Benchmark "kernel_10_474" written by ABC on Sun Jul 19 10:29:20 2020

module kernel_10_474 ( 
    i_10_474_156_0, i_10_474_175_0, i_10_474_176_0, i_10_474_243_0,
    i_10_474_280_0, i_10_474_328_0, i_10_474_390_0, i_10_474_427_0,
    i_10_474_428_0, i_10_474_438_0, i_10_474_444_0, i_10_474_447_0,
    i_10_474_463_0, i_10_474_506_0, i_10_474_516_0, i_10_474_519_0,
    i_10_474_748_0, i_10_474_752_0, i_10_474_796_0, i_10_474_955_0,
    i_10_474_1032_0, i_10_474_1033_0, i_10_474_1233_0, i_10_474_1307_0,
    i_10_474_1308_0, i_10_474_1311_0, i_10_474_1448_0, i_10_474_1550_0,
    i_10_474_1651_0, i_10_474_1681_0, i_10_474_1682_0, i_10_474_1687_0,
    i_10_474_1822_0, i_10_474_1823_0, i_10_474_1824_0, i_10_474_2016_0,
    i_10_474_2353_0, i_10_474_2354_0, i_10_474_2364_0, i_10_474_2407_0,
    i_10_474_2457_0, i_10_474_2629_0, i_10_474_2631_0, i_10_474_2632_0,
    i_10_474_2636_0, i_10_474_2662_0, i_10_474_2700_0, i_10_474_2701_0,
    i_10_474_2713_0, i_10_474_2714_0, i_10_474_2716_0, i_10_474_2723_0,
    i_10_474_2823_0, i_10_474_2885_0, i_10_474_2920_0, i_10_474_2980_0,
    i_10_474_2981_0, i_10_474_2982_0, i_10_474_2983_0, i_10_474_2984_0,
    i_10_474_2985_0, i_10_474_3036_0, i_10_474_3040_0, i_10_474_3043_0,
    i_10_474_3074_0, i_10_474_3199_0, i_10_474_3276_0, i_10_474_3388_0,
    i_10_474_3405_0, i_10_474_3406_0, i_10_474_3522_0, i_10_474_3613_0,
    i_10_474_3615_0, i_10_474_3650_0, i_10_474_3783_0, i_10_474_3841_0,
    i_10_474_3852_0, i_10_474_3853_0, i_10_474_3854_0, i_10_474_3856_0,
    i_10_474_3888_0, i_10_474_3910_0, i_10_474_3912_0, i_10_474_3982_0,
    i_10_474_3983_0, i_10_474_3990_0, i_10_474_4114_0, i_10_474_4116_0,
    i_10_474_4117_0, i_10_474_4119_0, i_10_474_4266_0, i_10_474_4269_0,
    i_10_474_4271_0, i_10_474_4273_0, i_10_474_4276_0, i_10_474_4277_0,
    i_10_474_4289_0, i_10_474_4292_0, i_10_474_4567_0, i_10_474_4570_0,
    o_10_474_0_0  );
  input  i_10_474_156_0, i_10_474_175_0, i_10_474_176_0, i_10_474_243_0,
    i_10_474_280_0, i_10_474_328_0, i_10_474_390_0, i_10_474_427_0,
    i_10_474_428_0, i_10_474_438_0, i_10_474_444_0, i_10_474_447_0,
    i_10_474_463_0, i_10_474_506_0, i_10_474_516_0, i_10_474_519_0,
    i_10_474_748_0, i_10_474_752_0, i_10_474_796_0, i_10_474_955_0,
    i_10_474_1032_0, i_10_474_1033_0, i_10_474_1233_0, i_10_474_1307_0,
    i_10_474_1308_0, i_10_474_1311_0, i_10_474_1448_0, i_10_474_1550_0,
    i_10_474_1651_0, i_10_474_1681_0, i_10_474_1682_0, i_10_474_1687_0,
    i_10_474_1822_0, i_10_474_1823_0, i_10_474_1824_0, i_10_474_2016_0,
    i_10_474_2353_0, i_10_474_2354_0, i_10_474_2364_0, i_10_474_2407_0,
    i_10_474_2457_0, i_10_474_2629_0, i_10_474_2631_0, i_10_474_2632_0,
    i_10_474_2636_0, i_10_474_2662_0, i_10_474_2700_0, i_10_474_2701_0,
    i_10_474_2713_0, i_10_474_2714_0, i_10_474_2716_0, i_10_474_2723_0,
    i_10_474_2823_0, i_10_474_2885_0, i_10_474_2920_0, i_10_474_2980_0,
    i_10_474_2981_0, i_10_474_2982_0, i_10_474_2983_0, i_10_474_2984_0,
    i_10_474_2985_0, i_10_474_3036_0, i_10_474_3040_0, i_10_474_3043_0,
    i_10_474_3074_0, i_10_474_3199_0, i_10_474_3276_0, i_10_474_3388_0,
    i_10_474_3405_0, i_10_474_3406_0, i_10_474_3522_0, i_10_474_3613_0,
    i_10_474_3615_0, i_10_474_3650_0, i_10_474_3783_0, i_10_474_3841_0,
    i_10_474_3852_0, i_10_474_3853_0, i_10_474_3854_0, i_10_474_3856_0,
    i_10_474_3888_0, i_10_474_3910_0, i_10_474_3912_0, i_10_474_3982_0,
    i_10_474_3983_0, i_10_474_3990_0, i_10_474_4114_0, i_10_474_4116_0,
    i_10_474_4117_0, i_10_474_4119_0, i_10_474_4266_0, i_10_474_4269_0,
    i_10_474_4271_0, i_10_474_4273_0, i_10_474_4276_0, i_10_474_4277_0,
    i_10_474_4289_0, i_10_474_4292_0, i_10_474_4567_0, i_10_474_4570_0;
  output o_10_474_0_0;
  assign o_10_474_0_0 = ~((~i_10_474_175_0 & ((i_10_474_1233_0 & i_10_474_3783_0) | (~i_10_474_2629_0 & ~i_10_474_2632_0 & i_10_474_4277_0))) | (i_10_474_280_0 & ((~i_10_474_2407_0 & ~i_10_474_2982_0 & ~i_10_474_2984_0 & i_10_474_3853_0 & ~i_10_474_4116_0) | (~i_10_474_243_0 & ~i_10_474_328_0 & ~i_10_474_463_0 & ~i_10_474_516_0 & ~i_10_474_4266_0))) | (~i_10_474_328_0 & ((~i_10_474_519_0 & ~i_10_474_2981_0 & ~i_10_474_2982_0 & i_10_474_3040_0 & ~i_10_474_4116_0) | (~i_10_474_516_0 & ~i_10_474_1822_0 & ~i_10_474_2354_0 & ~i_10_474_2631_0 & ~i_10_474_3040_0 & ~i_10_474_3613_0 & ~i_10_474_4119_0))) | (~i_10_474_444_0 & ((~i_10_474_1651_0 & ~i_10_474_2629_0 & ~i_10_474_2980_0 & ~i_10_474_2985_0 & ~i_10_474_3990_0) | (~i_10_474_516_0 & ~i_10_474_796_0 & ~i_10_474_2700_0 & ~i_10_474_2981_0 & ~i_10_474_3522_0 & ~i_10_474_3912_0 & ~i_10_474_4276_0))) | (~i_10_474_3888_0 & ((~i_10_474_519_0 & ~i_10_474_3910_0 & ((i_10_474_1824_0 & ~i_10_474_2457_0 & ~i_10_474_2980_0 & ~i_10_474_2985_0 & ~i_10_474_4269_0) | (~i_10_474_748_0 & ~i_10_474_2981_0 & ~i_10_474_4116_0 & ~i_10_474_4119_0 & ~i_10_474_4567_0))) | (~i_10_474_2354_0 & ((~i_10_474_1307_0 & ~i_10_474_2985_0 & ~i_10_474_3982_0 & ~i_10_474_4266_0 & ((~i_10_474_1233_0 & ~i_10_474_2016_0 & ~i_10_474_2407_0 & ~i_10_474_2980_0 & ~i_10_474_2982_0 & ~i_10_474_3276_0 & ~i_10_474_3406_0 & ~i_10_474_3912_0) | (~i_10_474_1308_0 & ~i_10_474_2716_0 & ~i_10_474_3522_0 & ~i_10_474_4567_0))) | (~i_10_474_438_0 & ~i_10_474_796_0 & i_10_474_1651_0 & ~i_10_474_2981_0 & ~i_10_474_2982_0 & ~i_10_474_3036_0 & ~i_10_474_4276_0 & ~i_10_474_4567_0))) | (i_10_474_444_0 & i_10_474_447_0 & ~i_10_474_2636_0 & ~i_10_474_2982_0 & ~i_10_474_3388_0 & ~i_10_474_3912_0 & ~i_10_474_3982_0 & ~i_10_474_4116_0 & ~i_10_474_4117_0) | (i_10_474_1233_0 & ~i_10_474_2700_0 & ~i_10_474_2980_0 & ~i_10_474_4119_0))) | (~i_10_474_1233_0 & ((i_10_474_1823_0 & i_10_474_3783_0 & ~i_10_474_3912_0 & ~i_10_474_4266_0) | (i_10_474_752_0 & i_10_474_2631_0 & ~i_10_474_2823_0 & ~i_10_474_2982_0 & ~i_10_474_4292_0))) | (~i_10_474_1550_0 & ~i_10_474_4266_0 & ((~i_10_474_748_0 & i_10_474_1307_0 & ~i_10_474_2823_0 & ~i_10_474_4114_0) | (~i_10_474_516_0 & ~i_10_474_2983_0 & ~i_10_474_3522_0 & ~i_10_474_3990_0 & ~i_10_474_4117_0 & ~i_10_474_4277_0))) | (~i_10_474_4269_0 & ((~i_10_474_748_0 & ((~i_10_474_1822_0 & ~i_10_474_2631_0 & i_10_474_2713_0) | (~i_10_474_1448_0 & ~i_10_474_2700_0 & ~i_10_474_2701_0 & ~i_10_474_3040_0 & ~i_10_474_3912_0 & ~i_10_474_4114_0 & ~i_10_474_4116_0 & ~i_10_474_4273_0))) | (~i_10_474_516_0 & ~i_10_474_2631_0 & ~i_10_474_2981_0 & ~i_10_474_4114_0 & ~i_10_474_4119_0 & ~i_10_474_4289_0 & ~i_10_474_4570_0))) | (~i_10_474_516_0 & ~i_10_474_2981_0 & ((i_10_474_3983_0 & i_10_474_4273_0) | (~i_10_474_2631_0 & ~i_10_474_2662_0 & ~i_10_474_2723_0 & ~i_10_474_2984_0 & ~i_10_474_3613_0 & ~i_10_474_4114_0 & ~i_10_474_4289_0))) | (~i_10_474_2985_0 & ((~i_10_474_428_0 & ~i_10_474_752_0 & i_10_474_3406_0 & ~i_10_474_3841_0 & ~i_10_474_3854_0) | (~i_10_474_2353_0 & ~i_10_474_2701_0 & i_10_474_3853_0 & ~i_10_474_3912_0) | (~i_10_474_463_0 & i_10_474_1823_0 & ~i_10_474_2354_0 & ~i_10_474_3650_0 & ~i_10_474_4567_0))) | (i_10_474_2016_0 & i_10_474_2713_0 & i_10_474_2920_0) | (i_10_474_463_0 & ~i_10_474_796_0 & i_10_474_1550_0 & ~i_10_474_4289_0) | (~i_10_474_2700_0 & i_10_474_2981_0 & ~i_10_474_2983_0 & i_10_474_4570_0));
endmodule



// Benchmark "kernel_10_475" written by ABC on Sun Jul 19 10:29:21 2020

module kernel_10_475 ( 
    i_10_475_171_0, i_10_475_216_0, i_10_475_280_0, i_10_475_316_0,
    i_10_475_408_0, i_10_475_425_0, i_10_475_431_0, i_10_475_434_0,
    i_10_475_437_0, i_10_475_439_0, i_10_475_441_0, i_10_475_442_0,
    i_10_475_443_0, i_10_475_445_0, i_10_475_457_0, i_10_475_515_0,
    i_10_475_518_0, i_10_475_749_0, i_10_475_892_0, i_10_475_901_0,
    i_10_475_957_0, i_10_475_958_0, i_10_475_968_0, i_10_475_1036_0,
    i_10_475_1037_0, i_10_475_1038_0, i_10_475_1141_0, i_10_475_1246_0,
    i_10_475_1247_0, i_10_475_1549_0, i_10_475_1579_0, i_10_475_1581_0,
    i_10_475_1648_0, i_10_475_1653_0, i_10_475_1654_0, i_10_475_1686_0,
    i_10_475_1818_0, i_10_475_1823_0, i_10_475_2006_0, i_10_475_2022_0,
    i_10_475_2332_0, i_10_475_2364_0, i_10_475_2383_0, i_10_475_2449_0,
    i_10_475_2510_0, i_10_475_2629_0, i_10_475_2630_0, i_10_475_2632_0,
    i_10_475_2633_0, i_10_475_2634_0, i_10_475_2635_0, i_10_475_2636_0,
    i_10_475_2655_0, i_10_475_2675_0, i_10_475_2678_0, i_10_475_2721_0,
    i_10_475_2818_0, i_10_475_2822_0, i_10_475_2824_0, i_10_475_2880_0,
    i_10_475_2884_0, i_10_475_2885_0, i_10_475_2919_0, i_10_475_2923_0,
    i_10_475_2924_0, i_10_475_2984_0, i_10_475_2987_0, i_10_475_3043_0,
    i_10_475_3074_0, i_10_475_3152_0, i_10_475_3155_0, i_10_475_3196_0,
    i_10_475_3312_0, i_10_475_3391_0, i_10_475_3392_0, i_10_475_3497_0,
    i_10_475_3610_0, i_10_475_3611_0, i_10_475_3645_0, i_10_475_3784_0,
    i_10_475_3785_0, i_10_475_3787_0, i_10_475_3788_0, i_10_475_3834_0,
    i_10_475_3841_0, i_10_475_3849_0, i_10_475_3853_0, i_10_475_3888_0,
    i_10_475_3889_0, i_10_475_3890_0, i_10_475_3906_0, i_10_475_3911_0,
    i_10_475_3980_0, i_10_475_4087_0, i_10_475_4122_0, i_10_475_4127_0,
    i_10_475_4288_0, i_10_475_4289_0, i_10_475_4291_0, i_10_475_4568_0,
    o_10_475_0_0  );
  input  i_10_475_171_0, i_10_475_216_0, i_10_475_280_0, i_10_475_316_0,
    i_10_475_408_0, i_10_475_425_0, i_10_475_431_0, i_10_475_434_0,
    i_10_475_437_0, i_10_475_439_0, i_10_475_441_0, i_10_475_442_0,
    i_10_475_443_0, i_10_475_445_0, i_10_475_457_0, i_10_475_515_0,
    i_10_475_518_0, i_10_475_749_0, i_10_475_892_0, i_10_475_901_0,
    i_10_475_957_0, i_10_475_958_0, i_10_475_968_0, i_10_475_1036_0,
    i_10_475_1037_0, i_10_475_1038_0, i_10_475_1141_0, i_10_475_1246_0,
    i_10_475_1247_0, i_10_475_1549_0, i_10_475_1579_0, i_10_475_1581_0,
    i_10_475_1648_0, i_10_475_1653_0, i_10_475_1654_0, i_10_475_1686_0,
    i_10_475_1818_0, i_10_475_1823_0, i_10_475_2006_0, i_10_475_2022_0,
    i_10_475_2332_0, i_10_475_2364_0, i_10_475_2383_0, i_10_475_2449_0,
    i_10_475_2510_0, i_10_475_2629_0, i_10_475_2630_0, i_10_475_2632_0,
    i_10_475_2633_0, i_10_475_2634_0, i_10_475_2635_0, i_10_475_2636_0,
    i_10_475_2655_0, i_10_475_2675_0, i_10_475_2678_0, i_10_475_2721_0,
    i_10_475_2818_0, i_10_475_2822_0, i_10_475_2824_0, i_10_475_2880_0,
    i_10_475_2884_0, i_10_475_2885_0, i_10_475_2919_0, i_10_475_2923_0,
    i_10_475_2924_0, i_10_475_2984_0, i_10_475_2987_0, i_10_475_3043_0,
    i_10_475_3074_0, i_10_475_3152_0, i_10_475_3155_0, i_10_475_3196_0,
    i_10_475_3312_0, i_10_475_3391_0, i_10_475_3392_0, i_10_475_3497_0,
    i_10_475_3610_0, i_10_475_3611_0, i_10_475_3645_0, i_10_475_3784_0,
    i_10_475_3785_0, i_10_475_3787_0, i_10_475_3788_0, i_10_475_3834_0,
    i_10_475_3841_0, i_10_475_3849_0, i_10_475_3853_0, i_10_475_3888_0,
    i_10_475_3889_0, i_10_475_3890_0, i_10_475_3906_0, i_10_475_3911_0,
    i_10_475_3980_0, i_10_475_4087_0, i_10_475_4122_0, i_10_475_4127_0,
    i_10_475_4288_0, i_10_475_4289_0, i_10_475_4291_0, i_10_475_4568_0;
  output o_10_475_0_0;
  assign o_10_475_0_0 = ~((~i_10_475_2655_0 & ((~i_10_475_2824_0 & ((i_10_475_408_0 & ((~i_10_475_892_0 & ~i_10_475_957_0 & ~i_10_475_958_0 & ~i_10_475_1648_0) | (i_10_475_2678_0 & ~i_10_475_2919_0 & ~i_10_475_2984_0))) | (~i_10_475_425_0 & ~i_10_475_434_0 & ~i_10_475_2510_0 & ~i_10_475_2678_0 & ~i_10_475_2885_0 & i_10_475_3785_0 & ~i_10_475_3889_0 & ~i_10_475_3890_0))) | (i_10_475_280_0 & i_10_475_1818_0 & ~i_10_475_2636_0 & i_10_475_2675_0) | (~i_10_475_445_0 & i_10_475_1247_0 & ~i_10_475_1579_0 & ~i_10_475_2332_0 & i_10_475_3853_0) | (~i_10_475_316_0 & i_10_475_1654_0 & ~i_10_475_2022_0 & ~i_10_475_2510_0 & ~i_10_475_2633_0 & ~i_10_475_2984_0 & ~i_10_475_3611_0 & ~i_10_475_3785_0 & ~i_10_475_3889_0 & ~i_10_475_3890_0 & ~i_10_475_4568_0))) | (~i_10_475_441_0 & ~i_10_475_2885_0 & ((~i_10_475_445_0 & ~i_10_475_892_0 & ~i_10_475_1036_0 & ~i_10_475_1037_0 & ~i_10_475_2510_0 & ~i_10_475_2630_0 & ~i_10_475_2635_0 & ~i_10_475_2822_0 & ~i_10_475_2984_0 & ~i_10_475_3889_0 & ~i_10_475_3906_0 & ~i_10_475_3980_0) | (~i_10_475_316_0 & ~i_10_475_958_0 & ~i_10_475_1549_0 & i_10_475_1654_0 & i_10_475_2924_0 & ~i_10_475_3890_0 & ~i_10_475_3911_0 & ~i_10_475_4288_0))) | (~i_10_475_2630_0 & ((i_10_475_280_0 & ((~i_10_475_515_0 & ~i_10_475_2632_0 & ~i_10_475_2675_0 & ~i_10_475_2822_0 & i_10_475_3043_0) | (~i_10_475_518_0 & i_10_475_1686_0 & ~i_10_475_3312_0))) | (~i_10_475_316_0 & ~i_10_475_518_0 & ~i_10_475_957_0 & ~i_10_475_1818_0 & ~i_10_475_2633_0 & ~i_10_475_2824_0 & ((~i_10_475_443_0 & ~i_10_475_901_0 & ~i_10_475_1653_0 & ~i_10_475_2510_0 & ~i_10_475_2636_0 & ~i_10_475_3888_0) | (~i_10_475_216_0 & ~i_10_475_431_0 & ~i_10_475_2006_0 & ~i_10_475_2675_0 & ~i_10_475_2678_0 & ~i_10_475_2818_0 & ~i_10_475_3889_0))) | (~i_10_475_431_0 & ~i_10_475_3980_0 & ((i_10_475_2632_0 & ~i_10_475_2818_0 & i_10_475_3645_0 & ~i_10_475_3788_0 & i_10_475_3853_0) | (~i_10_475_515_0 & ~i_10_475_1036_0 & ~i_10_475_1037_0 & ~i_10_475_1549_0 & ~i_10_475_2006_0 & ~i_10_475_2636_0 & ~i_10_475_2678_0 & ~i_10_475_2987_0 & ~i_10_475_3888_0 & ~i_10_475_3889_0 & ~i_10_475_4568_0))) | (~i_10_475_1686_0 & ~i_10_475_2006_0 & ~i_10_475_2678_0 & ~i_10_475_2884_0 & ~i_10_475_2924_0 & ~i_10_475_2984_0 & i_10_475_3834_0 & ~i_10_475_3906_0 & ~i_10_475_4127_0))) | (~i_10_475_4289_0 & ((~i_10_475_437_0 & ((i_10_475_518_0 & ~i_10_475_2022_0 & i_10_475_2634_0 & i_10_475_2636_0 & ~i_10_475_2678_0 & ~i_10_475_2984_0 & ~i_10_475_3497_0 & ~i_10_475_3849_0 & ~i_10_475_4288_0) | (~i_10_475_445_0 & ~i_10_475_2632_0 & i_10_475_3392_0 & i_10_475_4291_0))) | (~i_10_475_3890_0 & ((~i_10_475_445_0 & ~i_10_475_2510_0 & ~i_10_475_2675_0 & ~i_10_475_3196_0 & i_10_475_3785_0 & ~i_10_475_3889_0 & ~i_10_475_3980_0) | (i_10_475_443_0 & ~i_10_475_2678_0 & i_10_475_2923_0 & ~i_10_475_2987_0 & ~i_10_475_4291_0))) | (~i_10_475_2383_0 & ~i_10_475_2884_0 & i_10_475_3392_0 & ~i_10_475_3497_0 & ~i_10_475_3610_0 & ~i_10_475_3784_0 & ~i_10_475_4288_0))) | (~i_10_475_2818_0 & ((~i_10_475_437_0 & ((~i_10_475_968_0 & i_10_475_2383_0 & ~i_10_475_2984_0 & ~i_10_475_3611_0 & ~i_10_475_3889_0 & i_10_475_4291_0) | (i_10_475_280_0 & ~i_10_475_425_0 & ~i_10_475_957_0 & ~i_10_475_2633_0 & ~i_10_475_2987_0 & ~i_10_475_3888_0 & ~i_10_475_3980_0 & ~i_10_475_4568_0))) | (~i_10_475_2822_0 & ((~i_10_475_968_0 & ((i_10_475_171_0 & ~i_10_475_515_0 & ~i_10_475_749_0 & ~i_10_475_901_0 & ~i_10_475_3834_0) | (i_10_475_441_0 & ~i_10_475_1037_0 & ~i_10_475_1579_0 & ~i_10_475_2006_0 & i_10_475_2449_0 & ~i_10_475_3890_0))) | (~i_10_475_958_0 & ~i_10_475_2678_0 & i_10_475_3043_0 & i_10_475_3391_0))))) | (~i_10_475_3889_0 & ((~i_10_475_434_0 & ((~i_10_475_1036_0 & ~i_10_475_1579_0 & i_10_475_1648_0 & ~i_10_475_2678_0 & i_10_475_2721_0 & i_10_475_3610_0) | (~i_10_475_431_0 & ~i_10_475_901_0 & ~i_10_475_968_0 & ~i_10_475_2675_0 & ~i_10_475_2884_0 & i_10_475_2923_0 & ~i_10_475_2984_0 & ~i_10_475_3890_0))) | (~i_10_475_2510_0 & ((~i_10_475_518_0 & i_10_475_2022_0 & ~i_10_475_2987_0) | (~i_10_475_457_0 & i_10_475_1654_0 & ~i_10_475_2633_0 & i_10_475_2634_0 & ~i_10_475_3610_0))) | (~i_10_475_892_0 & ~i_10_475_901_0 & ~i_10_475_1549_0 & i_10_475_1648_0 & ~i_10_475_2633_0 & ~i_10_475_2675_0 & ~i_10_475_2822_0 & ~i_10_475_3497_0) | (~i_10_475_1823_0 & ~i_10_475_2635_0 & i_10_475_2721_0 & ~i_10_475_2984_0 & ~i_10_475_3645_0 & ~i_10_475_3906_0 & ~i_10_475_4288_0))) | (~i_10_475_968_0 & ((~i_10_475_434_0 & ~i_10_475_439_0 & ~i_10_475_749_0 & ~i_10_475_1037_0 & ~i_10_475_2629_0 & ~i_10_475_2822_0 & i_10_475_2924_0 & ~i_10_475_2984_0 & ~i_10_475_3787_0 & ~i_10_475_3890_0) | (~i_10_475_2635_0 & ~i_10_475_2987_0 & i_10_475_3391_0 & i_10_475_4291_0))) | (i_10_475_2449_0 & i_10_475_3392_0 & i_10_475_3853_0 & i_10_475_4568_0));
endmodule



// Benchmark "kernel_10_476" written by ABC on Sun Jul 19 10:29:22 2020

module kernel_10_476 ( 
    i_10_476_140_0, i_10_476_223_0, i_10_476_248_0, i_10_476_251_0,
    i_10_476_275_0, i_10_476_276_0, i_10_476_281_0, i_10_476_318_0,
    i_10_476_438_0, i_10_476_442_0, i_10_476_448_0, i_10_476_449_0,
    i_10_476_464_0, i_10_476_467_0, i_10_476_480_0, i_10_476_514_0,
    i_10_476_515_0, i_10_476_518_0, i_10_476_534_0, i_10_476_716_0,
    i_10_476_719_0, i_10_476_732_0, i_10_476_754_0, i_10_476_791_0,
    i_10_476_796_0, i_10_476_799_0, i_10_476_800_0, i_10_476_835_0,
    i_10_476_836_0, i_10_476_967_0, i_10_476_969_0, i_10_476_988_0,
    i_10_476_1115_0, i_10_476_1163_0, i_10_476_1166_0, i_10_476_1214_0,
    i_10_476_1309_0, i_10_476_1446_0, i_10_476_1492_0, i_10_476_1493_0,
    i_10_476_1546_0, i_10_476_1572_0, i_10_476_1653_0, i_10_476_1799_0,
    i_10_476_1808_0, i_10_476_1820_0, i_10_476_1825_0, i_10_476_1943_0,
    i_10_476_1952_0, i_10_476_2030_0, i_10_476_2255_0, i_10_476_2310_0,
    i_10_476_2356_0, i_10_476_2357_0, i_10_476_2363_0, i_10_476_2456_0,
    i_10_476_2534_0, i_10_476_2545_0, i_10_476_2546_0, i_10_476_2562_0,
    i_10_476_2607_0, i_10_476_2609_0, i_10_476_2678_0, i_10_476_2717_0,
    i_10_476_2725_0, i_10_476_2741_0, i_10_476_2876_0, i_10_476_2915_0,
    i_10_476_2919_0, i_10_476_2920_0, i_10_476_2968_0, i_10_476_2982_0,
    i_10_476_2986_0, i_10_476_3030_0, i_10_476_3038_0, i_10_476_3122_0,
    i_10_476_3284_0, i_10_476_3314_0, i_10_476_3315_0, i_10_476_3316_0,
    i_10_476_3320_0, i_10_476_3496_0, i_10_476_3526_0, i_10_476_3590_0,
    i_10_476_3617_0, i_10_476_3803_0, i_10_476_3806_0, i_10_476_3848_0,
    i_10_476_3860_0, i_10_476_3878_0, i_10_476_3946_0, i_10_476_3948_0,
    i_10_476_4182_0, i_10_476_4183_0, i_10_476_4268_0, i_10_476_4292_0,
    i_10_476_4306_0, i_10_476_4371_0, i_10_476_4459_0, i_10_476_4463_0,
    o_10_476_0_0  );
  input  i_10_476_140_0, i_10_476_223_0, i_10_476_248_0, i_10_476_251_0,
    i_10_476_275_0, i_10_476_276_0, i_10_476_281_0, i_10_476_318_0,
    i_10_476_438_0, i_10_476_442_0, i_10_476_448_0, i_10_476_449_0,
    i_10_476_464_0, i_10_476_467_0, i_10_476_480_0, i_10_476_514_0,
    i_10_476_515_0, i_10_476_518_0, i_10_476_534_0, i_10_476_716_0,
    i_10_476_719_0, i_10_476_732_0, i_10_476_754_0, i_10_476_791_0,
    i_10_476_796_0, i_10_476_799_0, i_10_476_800_0, i_10_476_835_0,
    i_10_476_836_0, i_10_476_967_0, i_10_476_969_0, i_10_476_988_0,
    i_10_476_1115_0, i_10_476_1163_0, i_10_476_1166_0, i_10_476_1214_0,
    i_10_476_1309_0, i_10_476_1446_0, i_10_476_1492_0, i_10_476_1493_0,
    i_10_476_1546_0, i_10_476_1572_0, i_10_476_1653_0, i_10_476_1799_0,
    i_10_476_1808_0, i_10_476_1820_0, i_10_476_1825_0, i_10_476_1943_0,
    i_10_476_1952_0, i_10_476_2030_0, i_10_476_2255_0, i_10_476_2310_0,
    i_10_476_2356_0, i_10_476_2357_0, i_10_476_2363_0, i_10_476_2456_0,
    i_10_476_2534_0, i_10_476_2545_0, i_10_476_2546_0, i_10_476_2562_0,
    i_10_476_2607_0, i_10_476_2609_0, i_10_476_2678_0, i_10_476_2717_0,
    i_10_476_2725_0, i_10_476_2741_0, i_10_476_2876_0, i_10_476_2915_0,
    i_10_476_2919_0, i_10_476_2920_0, i_10_476_2968_0, i_10_476_2982_0,
    i_10_476_2986_0, i_10_476_3030_0, i_10_476_3038_0, i_10_476_3122_0,
    i_10_476_3284_0, i_10_476_3314_0, i_10_476_3315_0, i_10_476_3316_0,
    i_10_476_3320_0, i_10_476_3496_0, i_10_476_3526_0, i_10_476_3590_0,
    i_10_476_3617_0, i_10_476_3803_0, i_10_476_3806_0, i_10_476_3848_0,
    i_10_476_3860_0, i_10_476_3878_0, i_10_476_3946_0, i_10_476_3948_0,
    i_10_476_4182_0, i_10_476_4183_0, i_10_476_4268_0, i_10_476_4292_0,
    i_10_476_4306_0, i_10_476_4371_0, i_10_476_4459_0, i_10_476_4463_0;
  output o_10_476_0_0;
  assign o_10_476_0_0 = 0;
endmodule



// Benchmark "kernel_10_477" written by ABC on Sun Jul 19 10:29:23 2020

module kernel_10_477 ( 
    i_10_477_29_0, i_10_477_244_0, i_10_477_254_0, i_10_477_272_0,
    i_10_477_283_0, i_10_477_286_0, i_10_477_391_0, i_10_477_427_0,
    i_10_477_428_0, i_10_477_434_0, i_10_477_435_0, i_10_477_436_0,
    i_10_477_443_0, i_10_477_445_0, i_10_477_463_0, i_10_477_505_0,
    i_10_477_792_0, i_10_477_958_0, i_10_477_1026_0, i_10_477_1027_0,
    i_10_477_1028_0, i_10_477_1080_0, i_10_477_1081_0, i_10_477_1085_0,
    i_10_477_1135_0, i_10_477_1235_0, i_10_477_1305_0, i_10_477_1306_0,
    i_10_477_1307_0, i_10_477_1308_0, i_10_477_1309_0, i_10_477_1364_0,
    i_10_477_1433_0, i_10_477_1436_0, i_10_477_1621_0, i_10_477_1823_0,
    i_10_477_1910_0, i_10_477_1911_0, i_10_477_1913_0, i_10_477_1989_0,
    i_10_477_2030_0, i_10_477_2198_0, i_10_477_2358_0, i_10_477_2408_0,
    i_10_477_2449_0, i_10_477_2470_0, i_10_477_2539_0, i_10_477_2541_0,
    i_10_477_2565_0, i_10_477_2628_0, i_10_477_2629_0, i_10_477_2630_0,
    i_10_477_2631_0, i_10_477_2632_0, i_10_477_2674_0, i_10_477_2675_0,
    i_10_477_2709_0, i_10_477_2710_0, i_10_477_2714_0, i_10_477_2720_0,
    i_10_477_2724_0, i_10_477_2730_0, i_10_477_2827_0, i_10_477_2828_0,
    i_10_477_2830_0, i_10_477_2845_0, i_10_477_2883_0, i_10_477_2919_0,
    i_10_477_3033_0, i_10_477_3069_0, i_10_477_3070_0, i_10_477_3071_0,
    i_10_477_3267_0, i_10_477_3321_0, i_10_477_3322_0, i_10_477_3323_0,
    i_10_477_3328_0, i_10_477_3467_0, i_10_477_3556_0, i_10_477_3584_0,
    i_10_477_3587_0, i_10_477_3609_0, i_10_477_3645_0, i_10_477_3837_0,
    i_10_477_3838_0, i_10_477_3839_0, i_10_477_3843_0, i_10_477_3846_0,
    i_10_477_3847_0, i_10_477_3848_0, i_10_477_3980_0, i_10_477_4030_0,
    i_10_477_4122_0, i_10_477_4123_0, i_10_477_4125_0, i_10_477_4127_0,
    i_10_477_4167_0, i_10_477_4172_0, i_10_477_4266_0, i_10_477_4278_0,
    o_10_477_0_0  );
  input  i_10_477_29_0, i_10_477_244_0, i_10_477_254_0, i_10_477_272_0,
    i_10_477_283_0, i_10_477_286_0, i_10_477_391_0, i_10_477_427_0,
    i_10_477_428_0, i_10_477_434_0, i_10_477_435_0, i_10_477_436_0,
    i_10_477_443_0, i_10_477_445_0, i_10_477_463_0, i_10_477_505_0,
    i_10_477_792_0, i_10_477_958_0, i_10_477_1026_0, i_10_477_1027_0,
    i_10_477_1028_0, i_10_477_1080_0, i_10_477_1081_0, i_10_477_1085_0,
    i_10_477_1135_0, i_10_477_1235_0, i_10_477_1305_0, i_10_477_1306_0,
    i_10_477_1307_0, i_10_477_1308_0, i_10_477_1309_0, i_10_477_1364_0,
    i_10_477_1433_0, i_10_477_1436_0, i_10_477_1621_0, i_10_477_1823_0,
    i_10_477_1910_0, i_10_477_1911_0, i_10_477_1913_0, i_10_477_1989_0,
    i_10_477_2030_0, i_10_477_2198_0, i_10_477_2358_0, i_10_477_2408_0,
    i_10_477_2449_0, i_10_477_2470_0, i_10_477_2539_0, i_10_477_2541_0,
    i_10_477_2565_0, i_10_477_2628_0, i_10_477_2629_0, i_10_477_2630_0,
    i_10_477_2631_0, i_10_477_2632_0, i_10_477_2674_0, i_10_477_2675_0,
    i_10_477_2709_0, i_10_477_2710_0, i_10_477_2714_0, i_10_477_2720_0,
    i_10_477_2724_0, i_10_477_2730_0, i_10_477_2827_0, i_10_477_2828_0,
    i_10_477_2830_0, i_10_477_2845_0, i_10_477_2883_0, i_10_477_2919_0,
    i_10_477_3033_0, i_10_477_3069_0, i_10_477_3070_0, i_10_477_3071_0,
    i_10_477_3267_0, i_10_477_3321_0, i_10_477_3322_0, i_10_477_3323_0,
    i_10_477_3328_0, i_10_477_3467_0, i_10_477_3556_0, i_10_477_3584_0,
    i_10_477_3587_0, i_10_477_3609_0, i_10_477_3645_0, i_10_477_3837_0,
    i_10_477_3838_0, i_10_477_3839_0, i_10_477_3843_0, i_10_477_3846_0,
    i_10_477_3847_0, i_10_477_3848_0, i_10_477_3980_0, i_10_477_4030_0,
    i_10_477_4122_0, i_10_477_4123_0, i_10_477_4125_0, i_10_477_4127_0,
    i_10_477_4167_0, i_10_477_4172_0, i_10_477_4266_0, i_10_477_4278_0;
  output o_10_477_0_0;
  assign o_10_477_0_0 = ~((~i_10_477_2710_0 & ((~i_10_477_29_0 & ((~i_10_477_391_0 & i_10_477_1823_0 & i_10_477_2449_0 & ~i_10_477_3846_0 & ~i_10_477_3848_0) | (~i_10_477_283_0 & ~i_10_477_1085_0 & ~i_10_477_1989_0 & ~i_10_477_3070_0 & ~i_10_477_3847_0 & ~i_10_477_4122_0))) | (~i_10_477_1621_0 & ~i_10_477_2030_0 & ~i_10_477_2709_0 & ~i_10_477_3071_0 & ~i_10_477_3587_0 & ~i_10_477_3848_0 & ~i_10_477_4266_0))) | (~i_10_477_3069_0 & ((~i_10_477_254_0 & ~i_10_477_2030_0 & ((~i_10_477_391_0 & ~i_10_477_1027_0 & ~i_10_477_1028_0 & ~i_10_477_1080_0 & ~i_10_477_1621_0 & ~i_10_477_3070_0) | (~i_10_477_792_0 & i_10_477_2714_0 & ~i_10_477_3071_0 & ~i_10_477_4123_0))) | (~i_10_477_283_0 & ~i_10_477_1433_0 & ((~i_10_477_3071_0 & ~i_10_477_4123_0) | (~i_10_477_1989_0 & ~i_10_477_3839_0))) | (i_10_477_283_0 & ~i_10_477_463_0 & ~i_10_477_792_0 & ~i_10_477_1026_0 & ~i_10_477_1085_0 & ~i_10_477_3467_0 & ~i_10_477_3847_0))) | (~i_10_477_1989_0 & ((~i_10_477_254_0 & ~i_10_477_2565_0 & ((~i_10_477_244_0 & ~i_10_477_1081_0 & ~i_10_477_3071_0 & ~i_10_477_3467_0 & ~i_10_477_3584_0 & ~i_10_477_3837_0) | (~i_10_477_3843_0 & ~i_10_477_3848_0 & ~i_10_477_4172_0 & ~i_10_477_4278_0))) | (~i_10_477_3071_0 & ~i_10_477_3609_0 & ~i_10_477_3838_0 & ~i_10_477_4127_0))) | (~i_10_477_1028_0 & ~i_10_477_3467_0 & ((~i_10_477_1027_0 & ~i_10_477_1433_0 & ~i_10_477_2709_0 & ~i_10_477_3071_0) | (~i_10_477_2629_0 & ~i_10_477_2828_0 & ~i_10_477_3070_0 & ~i_10_477_3267_0 & ~i_10_477_4123_0 & ~i_10_477_4127_0 & ~i_10_477_4167_0 & ~i_10_477_4266_0))) | (i_10_477_1305_0 & ((~i_10_477_1436_0 & i_10_477_3033_0 & ~i_10_477_3846_0) | (i_10_477_1433_0 & ~i_10_477_3267_0 & ~i_10_477_3843_0 & ~i_10_477_3847_0 & ~i_10_477_4278_0))) | (i_10_477_2632_0 & ((i_10_477_436_0 & i_10_477_2628_0) | (~i_10_477_2830_0 & ~i_10_477_3838_0))) | (i_10_477_2630_0 & ((i_10_477_3267_0 & (~i_10_477_2358_0 | (~i_10_477_958_0 & i_10_477_2631_0 & ~i_10_477_4125_0))) | (i_10_477_958_0 & i_10_477_1307_0) | (i_10_477_434_0 & i_10_477_4122_0 & ~i_10_477_4125_0 & ~i_10_477_4127_0))) | (i_10_477_2674_0 & i_10_477_3609_0 & ~i_10_477_3848_0) | (i_10_477_2720_0 & i_10_477_3848_0 & i_10_477_3980_0) | (i_10_477_1306_0 & ~i_10_477_1433_0 & i_10_477_2449_0 & ~i_10_477_3267_0 & ~i_10_477_3846_0 & ~i_10_477_4167_0));
endmodule



// Benchmark "kernel_10_478" written by ABC on Sun Jul 19 10:29:24 2020

module kernel_10_478 ( 
    i_10_478_13_0, i_10_478_31_0, i_10_478_174_0, i_10_478_221_0,
    i_10_478_223_0, i_10_478_224_0, i_10_478_285_0, i_10_478_286_0,
    i_10_478_315_0, i_10_478_316_0, i_10_478_435_0, i_10_478_725_0,
    i_10_478_748_0, i_10_478_820_0, i_10_478_967_0, i_10_478_983_0,
    i_10_478_999_0, i_10_478_1010_0, i_10_478_1107_0, i_10_478_1218_0,
    i_10_478_1233_0, i_10_478_1234_0, i_10_478_1240_0, i_10_478_1279_0,
    i_10_478_1296_0, i_10_478_1302_0, i_10_478_1344_0, i_10_478_1432_0,
    i_10_478_1535_0, i_10_478_1539_0, i_10_478_1540_0, i_10_478_1562_0,
    i_10_478_1683_0, i_10_478_1684_0, i_10_478_1686_0, i_10_478_1689_0,
    i_10_478_1691_0, i_10_478_1795_0, i_10_478_1800_0, i_10_478_1803_0,
    i_10_478_1821_0, i_10_478_1980_0, i_10_478_1982_0, i_10_478_2038_0,
    i_10_478_2089_0, i_10_478_2090_0, i_10_478_2199_0, i_10_478_2235_0,
    i_10_478_2252_0, i_10_478_2255_0, i_10_478_2290_0, i_10_478_2352_0,
    i_10_478_2355_0, i_10_478_2452_0, i_10_478_2466_0, i_10_478_2467_0,
    i_10_478_2471_0, i_10_478_2503_0, i_10_478_2565_0, i_10_478_2567_0,
    i_10_478_2574_0, i_10_478_2631_0, i_10_478_2721_0, i_10_478_2726_0,
    i_10_478_2727_0, i_10_478_2728_0, i_10_478_2730_0, i_10_478_2832_0,
    i_10_478_2847_0, i_10_478_2914_0, i_10_478_2964_0, i_10_478_3045_0,
    i_10_478_3384_0, i_10_478_3432_0, i_10_478_3468_0, i_10_478_3469_0,
    i_10_478_3537_0, i_10_478_3582_0, i_10_478_3612_0, i_10_478_3614_0,
    i_10_478_3793_0, i_10_478_3834_0, i_10_478_3854_0, i_10_478_3855_0,
    i_10_478_3860_0, i_10_478_3873_0, i_10_478_3874_0, i_10_478_3911_0,
    i_10_478_3988_0, i_10_478_4122_0, i_10_478_4125_0, i_10_478_4154_0,
    i_10_478_4168_0, i_10_478_4218_0, i_10_478_4283_0, i_10_478_4287_0,
    i_10_478_4460_0, i_10_478_4502_0, i_10_478_4545_0, i_10_478_4546_0,
    o_10_478_0_0  );
  input  i_10_478_13_0, i_10_478_31_0, i_10_478_174_0, i_10_478_221_0,
    i_10_478_223_0, i_10_478_224_0, i_10_478_285_0, i_10_478_286_0,
    i_10_478_315_0, i_10_478_316_0, i_10_478_435_0, i_10_478_725_0,
    i_10_478_748_0, i_10_478_820_0, i_10_478_967_0, i_10_478_983_0,
    i_10_478_999_0, i_10_478_1010_0, i_10_478_1107_0, i_10_478_1218_0,
    i_10_478_1233_0, i_10_478_1234_0, i_10_478_1240_0, i_10_478_1279_0,
    i_10_478_1296_0, i_10_478_1302_0, i_10_478_1344_0, i_10_478_1432_0,
    i_10_478_1535_0, i_10_478_1539_0, i_10_478_1540_0, i_10_478_1562_0,
    i_10_478_1683_0, i_10_478_1684_0, i_10_478_1686_0, i_10_478_1689_0,
    i_10_478_1691_0, i_10_478_1795_0, i_10_478_1800_0, i_10_478_1803_0,
    i_10_478_1821_0, i_10_478_1980_0, i_10_478_1982_0, i_10_478_2038_0,
    i_10_478_2089_0, i_10_478_2090_0, i_10_478_2199_0, i_10_478_2235_0,
    i_10_478_2252_0, i_10_478_2255_0, i_10_478_2290_0, i_10_478_2352_0,
    i_10_478_2355_0, i_10_478_2452_0, i_10_478_2466_0, i_10_478_2467_0,
    i_10_478_2471_0, i_10_478_2503_0, i_10_478_2565_0, i_10_478_2567_0,
    i_10_478_2574_0, i_10_478_2631_0, i_10_478_2721_0, i_10_478_2726_0,
    i_10_478_2727_0, i_10_478_2728_0, i_10_478_2730_0, i_10_478_2832_0,
    i_10_478_2847_0, i_10_478_2914_0, i_10_478_2964_0, i_10_478_3045_0,
    i_10_478_3384_0, i_10_478_3432_0, i_10_478_3468_0, i_10_478_3469_0,
    i_10_478_3537_0, i_10_478_3582_0, i_10_478_3612_0, i_10_478_3614_0,
    i_10_478_3793_0, i_10_478_3834_0, i_10_478_3854_0, i_10_478_3855_0,
    i_10_478_3860_0, i_10_478_3873_0, i_10_478_3874_0, i_10_478_3911_0,
    i_10_478_3988_0, i_10_478_4122_0, i_10_478_4125_0, i_10_478_4154_0,
    i_10_478_4168_0, i_10_478_4218_0, i_10_478_4283_0, i_10_478_4287_0,
    i_10_478_4460_0, i_10_478_4502_0, i_10_478_4545_0, i_10_478_4546_0;
  output o_10_478_0_0;
  assign o_10_478_0_0 = 0;
endmodule



// Benchmark "kernel_10_479" written by ABC on Sun Jul 19 10:29:25 2020

module kernel_10_479 ( 
    i_10_479_118_0, i_10_479_121_0, i_10_479_248_0, i_10_479_285_0,
    i_10_479_286_0, i_10_479_287_0, i_10_479_315_0, i_10_479_316_0,
    i_10_479_318_0, i_10_479_365_0, i_10_479_406_0, i_10_479_408_0,
    i_10_479_424_0, i_10_479_434_0, i_10_479_443_0, i_10_479_447_0,
    i_10_479_448_0, i_10_479_793_0, i_10_479_794_0, i_10_479_797_0,
    i_10_479_893_0, i_10_479_959_0, i_10_479_1028_0, i_10_479_1031_0,
    i_10_479_1242_0, i_10_479_1243_0, i_10_479_1244_0, i_10_479_1305_0,
    i_10_479_1309_0, i_10_479_1444_0, i_10_479_1445_0, i_10_479_1546_0,
    i_10_479_1547_0, i_10_479_1576_0, i_10_479_1577_0, i_10_479_1580_0,
    i_10_479_1613_0, i_10_479_1650_0, i_10_479_1683_0, i_10_479_1687_0,
    i_10_479_1689_0, i_10_479_1801_0, i_10_479_1821_0, i_10_479_1990_0,
    i_10_479_2197_0, i_10_479_2304_0, i_10_479_2332_0, i_10_479_2361_0,
    i_10_479_2362_0, i_10_479_2363_0, i_10_479_2376_0, i_10_479_2407_0,
    i_10_479_2458_0, i_10_479_2467_0, i_10_479_2475_0, i_10_479_2648_0,
    i_10_479_2663_0, i_10_479_2713_0, i_10_479_2785_0, i_10_479_2828_0,
    i_10_479_2830_0, i_10_479_2831_0, i_10_479_2881_0, i_10_479_2917_0,
    i_10_479_2919_0, i_10_479_2920_0, i_10_479_3201_0, i_10_479_3269_0,
    i_10_479_3276_0, i_10_479_3277_0, i_10_479_3281_0, i_10_479_3294_0,
    i_10_479_3384_0, i_10_479_3386_0, i_10_479_3388_0, i_10_479_3550_0,
    i_10_479_3647_0, i_10_479_3686_0, i_10_479_3717_0, i_10_479_3781_0,
    i_10_479_3783_0, i_10_479_3784_0, i_10_479_3785_0, i_10_479_3786_0,
    i_10_479_3788_0, i_10_479_3842_0, i_10_479_3845_0, i_10_479_3846_0,
    i_10_479_3847_0, i_10_479_3851_0, i_10_479_3852_0, i_10_479_3854_0,
    i_10_479_3855_0, i_10_479_3888_0, i_10_479_3889_0, i_10_479_4061_0,
    i_10_479_4218_0, i_10_479_4219_0, i_10_479_4289_0, i_10_479_4564_0,
    o_10_479_0_0  );
  input  i_10_479_118_0, i_10_479_121_0, i_10_479_248_0, i_10_479_285_0,
    i_10_479_286_0, i_10_479_287_0, i_10_479_315_0, i_10_479_316_0,
    i_10_479_318_0, i_10_479_365_0, i_10_479_406_0, i_10_479_408_0,
    i_10_479_424_0, i_10_479_434_0, i_10_479_443_0, i_10_479_447_0,
    i_10_479_448_0, i_10_479_793_0, i_10_479_794_0, i_10_479_797_0,
    i_10_479_893_0, i_10_479_959_0, i_10_479_1028_0, i_10_479_1031_0,
    i_10_479_1242_0, i_10_479_1243_0, i_10_479_1244_0, i_10_479_1305_0,
    i_10_479_1309_0, i_10_479_1444_0, i_10_479_1445_0, i_10_479_1546_0,
    i_10_479_1547_0, i_10_479_1576_0, i_10_479_1577_0, i_10_479_1580_0,
    i_10_479_1613_0, i_10_479_1650_0, i_10_479_1683_0, i_10_479_1687_0,
    i_10_479_1689_0, i_10_479_1801_0, i_10_479_1821_0, i_10_479_1990_0,
    i_10_479_2197_0, i_10_479_2304_0, i_10_479_2332_0, i_10_479_2361_0,
    i_10_479_2362_0, i_10_479_2363_0, i_10_479_2376_0, i_10_479_2407_0,
    i_10_479_2458_0, i_10_479_2467_0, i_10_479_2475_0, i_10_479_2648_0,
    i_10_479_2663_0, i_10_479_2713_0, i_10_479_2785_0, i_10_479_2828_0,
    i_10_479_2830_0, i_10_479_2831_0, i_10_479_2881_0, i_10_479_2917_0,
    i_10_479_2919_0, i_10_479_2920_0, i_10_479_3201_0, i_10_479_3269_0,
    i_10_479_3276_0, i_10_479_3277_0, i_10_479_3281_0, i_10_479_3294_0,
    i_10_479_3384_0, i_10_479_3386_0, i_10_479_3388_0, i_10_479_3550_0,
    i_10_479_3647_0, i_10_479_3686_0, i_10_479_3717_0, i_10_479_3781_0,
    i_10_479_3783_0, i_10_479_3784_0, i_10_479_3785_0, i_10_479_3786_0,
    i_10_479_3788_0, i_10_479_3842_0, i_10_479_3845_0, i_10_479_3846_0,
    i_10_479_3847_0, i_10_479_3851_0, i_10_479_3852_0, i_10_479_3854_0,
    i_10_479_3855_0, i_10_479_3888_0, i_10_479_3889_0, i_10_479_4061_0,
    i_10_479_4218_0, i_10_479_4219_0, i_10_479_4289_0, i_10_479_4564_0;
  output o_10_479_0_0;
  assign o_10_479_0_0 = 0;
endmodule



// Benchmark "kernel_10_480" written by ABC on Sun Jul 19 10:29:26 2020

module kernel_10_480 ( 
    i_10_480_172_0, i_10_480_186_0, i_10_480_187_0, i_10_480_244_0,
    i_10_480_246_0, i_10_480_247_0, i_10_480_280_0, i_10_480_286_0,
    i_10_480_293_0, i_10_480_423_0, i_10_480_424_0, i_10_480_446_0,
    i_10_480_449_0, i_10_480_460_0, i_10_480_463_0, i_10_480_464_0,
    i_10_480_467_0, i_10_480_712_0, i_10_480_713_0, i_10_480_748_0,
    i_10_480_901_0, i_10_480_902_0, i_10_480_905_0, i_10_480_997_0,
    i_10_480_998_0, i_10_480_1034_0, i_10_480_1168_0, i_10_480_1222_0,
    i_10_480_1234_0, i_10_480_1237_0, i_10_480_1306_0, i_10_480_1309_0,
    i_10_480_1345_0, i_10_480_1361_0, i_10_480_1486_0, i_10_480_1556_0,
    i_10_480_1649_0, i_10_480_1683_0, i_10_480_1684_0, i_10_480_1686_0,
    i_10_480_1765_0, i_10_480_1766_0, i_10_480_1818_0, i_10_480_1825_0,
    i_10_480_1909_0, i_10_480_1914_0, i_10_480_1999_0, i_10_480_2183_0,
    i_10_480_2349_0, i_10_480_2365_0, i_10_480_2366_0, i_10_480_2380_0,
    i_10_480_2449_0, i_10_480_2450_0, i_10_480_2452_0, i_10_480_2470_0,
    i_10_480_2659_0, i_10_480_2725_0, i_10_480_2727_0, i_10_480_2782_0,
    i_10_480_2830_0, i_10_480_2883_0, i_10_480_2886_0, i_10_480_2918_0,
    i_10_480_3044_0, i_10_480_3070_0, i_10_480_3071_0, i_10_480_3115_0,
    i_10_480_3233_0, i_10_480_3276_0, i_10_480_3280_0, i_10_480_3281_0,
    i_10_480_3325_0, i_10_480_3389_0, i_10_480_3392_0, i_10_480_3407_0,
    i_10_480_3408_0, i_10_480_3409_0, i_10_480_3538_0, i_10_480_3583_0,
    i_10_480_3585_0, i_10_480_3586_0, i_10_480_3614_0, i_10_480_3653_0,
    i_10_480_3783_0, i_10_480_3787_0, i_10_480_3788_0, i_10_480_3808_0,
    i_10_480_3811_0, i_10_480_3812_0, i_10_480_3839_0, i_10_480_3855_0,
    i_10_480_3859_0, i_10_480_3966_0, i_10_480_3978_0, i_10_480_3980_0,
    i_10_480_3982_0, i_10_480_4115_0, i_10_480_4289_0, i_10_480_4291_0,
    o_10_480_0_0  );
  input  i_10_480_172_0, i_10_480_186_0, i_10_480_187_0, i_10_480_244_0,
    i_10_480_246_0, i_10_480_247_0, i_10_480_280_0, i_10_480_286_0,
    i_10_480_293_0, i_10_480_423_0, i_10_480_424_0, i_10_480_446_0,
    i_10_480_449_0, i_10_480_460_0, i_10_480_463_0, i_10_480_464_0,
    i_10_480_467_0, i_10_480_712_0, i_10_480_713_0, i_10_480_748_0,
    i_10_480_901_0, i_10_480_902_0, i_10_480_905_0, i_10_480_997_0,
    i_10_480_998_0, i_10_480_1034_0, i_10_480_1168_0, i_10_480_1222_0,
    i_10_480_1234_0, i_10_480_1237_0, i_10_480_1306_0, i_10_480_1309_0,
    i_10_480_1345_0, i_10_480_1361_0, i_10_480_1486_0, i_10_480_1556_0,
    i_10_480_1649_0, i_10_480_1683_0, i_10_480_1684_0, i_10_480_1686_0,
    i_10_480_1765_0, i_10_480_1766_0, i_10_480_1818_0, i_10_480_1825_0,
    i_10_480_1909_0, i_10_480_1914_0, i_10_480_1999_0, i_10_480_2183_0,
    i_10_480_2349_0, i_10_480_2365_0, i_10_480_2366_0, i_10_480_2380_0,
    i_10_480_2449_0, i_10_480_2450_0, i_10_480_2452_0, i_10_480_2470_0,
    i_10_480_2659_0, i_10_480_2725_0, i_10_480_2727_0, i_10_480_2782_0,
    i_10_480_2830_0, i_10_480_2883_0, i_10_480_2886_0, i_10_480_2918_0,
    i_10_480_3044_0, i_10_480_3070_0, i_10_480_3071_0, i_10_480_3115_0,
    i_10_480_3233_0, i_10_480_3276_0, i_10_480_3280_0, i_10_480_3281_0,
    i_10_480_3325_0, i_10_480_3389_0, i_10_480_3392_0, i_10_480_3407_0,
    i_10_480_3408_0, i_10_480_3409_0, i_10_480_3538_0, i_10_480_3583_0,
    i_10_480_3585_0, i_10_480_3586_0, i_10_480_3614_0, i_10_480_3653_0,
    i_10_480_3783_0, i_10_480_3787_0, i_10_480_3788_0, i_10_480_3808_0,
    i_10_480_3811_0, i_10_480_3812_0, i_10_480_3839_0, i_10_480_3855_0,
    i_10_480_3859_0, i_10_480_3966_0, i_10_480_3978_0, i_10_480_3980_0,
    i_10_480_3982_0, i_10_480_4115_0, i_10_480_4289_0, i_10_480_4291_0;
  output o_10_480_0_0;
  assign o_10_480_0_0 = 0;
endmodule



// Benchmark "kernel_10_481" written by ABC on Sun Jul 19 10:29:27 2020

module kernel_10_481 ( 
    i_10_481_44_0, i_10_481_58_0, i_10_481_153_0, i_10_481_208_0,
    i_10_481_257_0, i_10_481_263_0, i_10_481_281_0, i_10_481_283_0,
    i_10_481_317_0, i_10_481_355_0, i_10_481_389_0, i_10_481_392_0,
    i_10_481_499_0, i_10_481_657_0, i_10_481_658_0, i_10_481_893_0,
    i_10_481_1009_0, i_10_481_1010_0, i_10_481_1027_0, i_10_481_1084_0,
    i_10_481_1085_0, i_10_481_1206_0, i_10_481_1234_0, i_10_481_1238_0,
    i_10_481_1271_0, i_10_481_1297_0, i_10_481_1377_0, i_10_481_1396_0,
    i_10_481_1485_0, i_10_481_1550_0, i_10_481_1576_0, i_10_481_1593_0,
    i_10_481_1638_0, i_10_481_1651_0, i_10_481_1697_0, i_10_481_1712_0,
    i_10_481_1716_0, i_10_481_1730_0, i_10_481_1807_0, i_10_481_1809_0,
    i_10_481_1822_0, i_10_481_2000_0, i_10_481_2002_0, i_10_481_2027_0,
    i_10_481_2145_0, i_10_481_2231_0, i_10_481_2269_0, i_10_481_2307_0,
    i_10_481_2341_0, i_10_481_2343_0, i_10_481_2362_0, i_10_481_2467_0,
    i_10_481_2489_0, i_10_481_2504_0, i_10_481_2542_0, i_10_481_2556_0,
    i_10_481_2557_0, i_10_481_2575_0, i_10_481_2885_0, i_10_481_2954_0,
    i_10_481_2961_0, i_10_481_2971_0, i_10_481_2983_0, i_10_481_2984_0,
    i_10_481_3070_0, i_10_481_3071_0, i_10_481_3160_0, i_10_481_3197_0,
    i_10_481_3200_0, i_10_481_3266_0, i_10_481_3332_0, i_10_481_3358_0,
    i_10_481_3404_0, i_10_481_3467_0, i_10_481_3484_0, i_10_481_3539_0,
    i_10_481_3580_0, i_10_481_3584_0, i_10_481_3587_0, i_10_481_3613_0,
    i_10_481_3645_0, i_10_481_3729_0, i_10_481_3792_0, i_10_481_3808_0,
    i_10_481_3842_0, i_10_481_3898_0, i_10_481_3945_0, i_10_481_4069_0,
    i_10_481_4118_0, i_10_481_4144_0, i_10_481_4151_0, i_10_481_4204_0,
    i_10_481_4226_0, i_10_481_4270_0, i_10_481_4273_0, i_10_481_4394_0,
    i_10_481_4421_0, i_10_481_4522_0, i_10_481_4545_0, i_10_481_4546_0,
    o_10_481_0_0  );
  input  i_10_481_44_0, i_10_481_58_0, i_10_481_153_0, i_10_481_208_0,
    i_10_481_257_0, i_10_481_263_0, i_10_481_281_0, i_10_481_283_0,
    i_10_481_317_0, i_10_481_355_0, i_10_481_389_0, i_10_481_392_0,
    i_10_481_499_0, i_10_481_657_0, i_10_481_658_0, i_10_481_893_0,
    i_10_481_1009_0, i_10_481_1010_0, i_10_481_1027_0, i_10_481_1084_0,
    i_10_481_1085_0, i_10_481_1206_0, i_10_481_1234_0, i_10_481_1238_0,
    i_10_481_1271_0, i_10_481_1297_0, i_10_481_1377_0, i_10_481_1396_0,
    i_10_481_1485_0, i_10_481_1550_0, i_10_481_1576_0, i_10_481_1593_0,
    i_10_481_1638_0, i_10_481_1651_0, i_10_481_1697_0, i_10_481_1712_0,
    i_10_481_1716_0, i_10_481_1730_0, i_10_481_1807_0, i_10_481_1809_0,
    i_10_481_1822_0, i_10_481_2000_0, i_10_481_2002_0, i_10_481_2027_0,
    i_10_481_2145_0, i_10_481_2231_0, i_10_481_2269_0, i_10_481_2307_0,
    i_10_481_2341_0, i_10_481_2343_0, i_10_481_2362_0, i_10_481_2467_0,
    i_10_481_2489_0, i_10_481_2504_0, i_10_481_2542_0, i_10_481_2556_0,
    i_10_481_2557_0, i_10_481_2575_0, i_10_481_2885_0, i_10_481_2954_0,
    i_10_481_2961_0, i_10_481_2971_0, i_10_481_2983_0, i_10_481_2984_0,
    i_10_481_3070_0, i_10_481_3071_0, i_10_481_3160_0, i_10_481_3197_0,
    i_10_481_3200_0, i_10_481_3266_0, i_10_481_3332_0, i_10_481_3358_0,
    i_10_481_3404_0, i_10_481_3467_0, i_10_481_3484_0, i_10_481_3539_0,
    i_10_481_3580_0, i_10_481_3584_0, i_10_481_3587_0, i_10_481_3613_0,
    i_10_481_3645_0, i_10_481_3729_0, i_10_481_3792_0, i_10_481_3808_0,
    i_10_481_3842_0, i_10_481_3898_0, i_10_481_3945_0, i_10_481_4069_0,
    i_10_481_4118_0, i_10_481_4144_0, i_10_481_4151_0, i_10_481_4204_0,
    i_10_481_4226_0, i_10_481_4270_0, i_10_481_4273_0, i_10_481_4394_0,
    i_10_481_4421_0, i_10_481_4522_0, i_10_481_4545_0, i_10_481_4546_0;
  output o_10_481_0_0;
  assign o_10_481_0_0 = 0;
endmodule



// Benchmark "kernel_10_482" written by ABC on Sun Jul 19 10:29:28 2020

module kernel_10_482 ( 
    i_10_482_155_0, i_10_482_171_0, i_10_482_172_0, i_10_482_219_0,
    i_10_482_220_0, i_10_482_280_0, i_10_482_320_0, i_10_482_437_0,
    i_10_482_445_0, i_10_482_446_0, i_10_482_448_0, i_10_482_518_0,
    i_10_482_590_0, i_10_482_689_0, i_10_482_992_0, i_10_482_995_0,
    i_10_482_997_0, i_10_482_1026_0, i_10_482_1037_0, i_10_482_1040_0,
    i_10_482_1236_0, i_10_482_1241_0, i_10_482_1289_0, i_10_482_1305_0,
    i_10_482_1342_0, i_10_482_1346_0, i_10_482_1486_0, i_10_482_1487_0,
    i_10_482_1556_0, i_10_482_1595_0, i_10_482_1630_0, i_10_482_1647_0,
    i_10_482_1683_0, i_10_482_1686_0, i_10_482_1687_0, i_10_482_1771_0,
    i_10_482_1819_0, i_10_482_1821_0, i_10_482_1912_0, i_10_482_1913_0,
    i_10_482_1998_0, i_10_482_2002_0, i_10_482_2243_0, i_10_482_2252_0,
    i_10_482_2351_0, i_10_482_2408_0, i_10_482_2454_0, i_10_482_2456_0,
    i_10_482_2512_0, i_10_482_2543_0, i_10_482_2606_0, i_10_482_2609_0,
    i_10_482_2657_0, i_10_482_2660_0, i_10_482_2675_0, i_10_482_2720_0,
    i_10_482_2723_0, i_10_482_2724_0, i_10_482_2728_0, i_10_482_2729_0,
    i_10_482_2819_0, i_10_482_2821_0, i_10_482_2822_0, i_10_482_2885_0,
    i_10_482_2981_0, i_10_482_2984_0, i_10_482_3037_0, i_10_482_3089_0,
    i_10_482_3091_0, i_10_482_3095_0, i_10_482_3160_0, i_10_482_3161_0,
    i_10_482_3235_0, i_10_482_3236_0, i_10_482_3278_0, i_10_482_3281_0,
    i_10_482_3284_0, i_10_482_3388_0, i_10_482_3389_0, i_10_482_3391_0,
    i_10_482_3392_0, i_10_482_3469_0, i_10_482_3470_0, i_10_482_3523_0,
    i_10_482_3524_0, i_10_482_3525_0, i_10_482_3527_0, i_10_482_3554_0,
    i_10_482_3781_0, i_10_482_3785_0, i_10_482_3836_0, i_10_482_3980_0,
    i_10_482_3992_0, i_10_482_4055_0, i_10_482_4114_0, i_10_482_4126_0,
    i_10_482_4268_0, i_10_482_4285_0, i_10_482_4460_0, i_10_482_4565_0,
    o_10_482_0_0  );
  input  i_10_482_155_0, i_10_482_171_0, i_10_482_172_0, i_10_482_219_0,
    i_10_482_220_0, i_10_482_280_0, i_10_482_320_0, i_10_482_437_0,
    i_10_482_445_0, i_10_482_446_0, i_10_482_448_0, i_10_482_518_0,
    i_10_482_590_0, i_10_482_689_0, i_10_482_992_0, i_10_482_995_0,
    i_10_482_997_0, i_10_482_1026_0, i_10_482_1037_0, i_10_482_1040_0,
    i_10_482_1236_0, i_10_482_1241_0, i_10_482_1289_0, i_10_482_1305_0,
    i_10_482_1342_0, i_10_482_1346_0, i_10_482_1486_0, i_10_482_1487_0,
    i_10_482_1556_0, i_10_482_1595_0, i_10_482_1630_0, i_10_482_1647_0,
    i_10_482_1683_0, i_10_482_1686_0, i_10_482_1687_0, i_10_482_1771_0,
    i_10_482_1819_0, i_10_482_1821_0, i_10_482_1912_0, i_10_482_1913_0,
    i_10_482_1998_0, i_10_482_2002_0, i_10_482_2243_0, i_10_482_2252_0,
    i_10_482_2351_0, i_10_482_2408_0, i_10_482_2454_0, i_10_482_2456_0,
    i_10_482_2512_0, i_10_482_2543_0, i_10_482_2606_0, i_10_482_2609_0,
    i_10_482_2657_0, i_10_482_2660_0, i_10_482_2675_0, i_10_482_2720_0,
    i_10_482_2723_0, i_10_482_2724_0, i_10_482_2728_0, i_10_482_2729_0,
    i_10_482_2819_0, i_10_482_2821_0, i_10_482_2822_0, i_10_482_2885_0,
    i_10_482_2981_0, i_10_482_2984_0, i_10_482_3037_0, i_10_482_3089_0,
    i_10_482_3091_0, i_10_482_3095_0, i_10_482_3160_0, i_10_482_3161_0,
    i_10_482_3235_0, i_10_482_3236_0, i_10_482_3278_0, i_10_482_3281_0,
    i_10_482_3284_0, i_10_482_3388_0, i_10_482_3389_0, i_10_482_3391_0,
    i_10_482_3392_0, i_10_482_3469_0, i_10_482_3470_0, i_10_482_3523_0,
    i_10_482_3524_0, i_10_482_3525_0, i_10_482_3527_0, i_10_482_3554_0,
    i_10_482_3781_0, i_10_482_3785_0, i_10_482_3836_0, i_10_482_3980_0,
    i_10_482_3992_0, i_10_482_4055_0, i_10_482_4114_0, i_10_482_4126_0,
    i_10_482_4268_0, i_10_482_4285_0, i_10_482_4460_0, i_10_482_4565_0;
  output o_10_482_0_0;
  assign o_10_482_0_0 = 0;
endmodule



// Benchmark "kernel_10_483" written by ABC on Sun Jul 19 10:29:28 2020

module kernel_10_483 ( 
    i_10_483_284_0, i_10_483_287_0, i_10_483_318_0, i_10_483_323_0,
    i_10_483_388_0, i_10_483_412_0, i_10_483_431_0, i_10_483_443_0,
    i_10_483_465_0, i_10_483_719_0, i_10_483_800_0, i_10_483_1030_0,
    i_10_483_1038_0, i_10_483_1041_0, i_10_483_1043_0, i_10_483_1052_0,
    i_10_483_1053_0, i_10_483_1060_0, i_10_483_1061_0, i_10_483_1084_0,
    i_10_483_1269_0, i_10_483_1308_0, i_10_483_1311_0, i_10_483_1312_0,
    i_10_483_1394_0, i_10_483_1435_0, i_10_483_1439_0, i_10_483_1444_0,
    i_10_483_1539_0, i_10_483_1540_0, i_10_483_1577_0, i_10_483_1624_0,
    i_10_483_1652_0, i_10_483_1654_0, i_10_483_1686_0, i_10_483_1687_0,
    i_10_483_1689_0, i_10_483_1765_0, i_10_483_1769_0, i_10_483_1819_0,
    i_10_483_1824_0, i_10_483_1915_0, i_10_483_1999_0, i_10_483_2001_0,
    i_10_483_2159_0, i_10_483_2349_0, i_10_483_2352_0, i_10_483_2355_0,
    i_10_483_2357_0, i_10_483_2365_0, i_10_483_2376_0, i_10_483_2378_0,
    i_10_483_2405_0, i_10_483_2406_0, i_10_483_2454_0, i_10_483_2456_0,
    i_10_483_2470_0, i_10_483_2516_0, i_10_483_2564_0, i_10_483_2604_0,
    i_10_483_2632_0, i_10_483_2644_0, i_10_483_2677_0, i_10_483_2699_0,
    i_10_483_2714_0, i_10_483_2956_0, i_10_483_2959_0, i_10_483_2980_0,
    i_10_483_2982_0, i_10_483_2983_0, i_10_483_2984_0, i_10_483_2985_0,
    i_10_483_3036_0, i_10_483_3268_0, i_10_483_3272_0, i_10_483_3278_0,
    i_10_483_3297_0, i_10_483_3384_0, i_10_483_3385_0, i_10_483_3388_0,
    i_10_483_3389_0, i_10_483_3472_0, i_10_483_3617_0, i_10_483_3645_0,
    i_10_483_3649_0, i_10_483_3784_0, i_10_483_3785_0, i_10_483_3834_0,
    i_10_483_3852_0, i_10_483_4009_0, i_10_483_4114_0, i_10_483_4125_0,
    i_10_483_4130_0, i_10_483_4170_0, i_10_483_4173_0, i_10_483_4174_0,
    i_10_483_4267_0, i_10_483_4271_0, i_10_483_4278_0, i_10_483_4279_0,
    o_10_483_0_0  );
  input  i_10_483_284_0, i_10_483_287_0, i_10_483_318_0, i_10_483_323_0,
    i_10_483_388_0, i_10_483_412_0, i_10_483_431_0, i_10_483_443_0,
    i_10_483_465_0, i_10_483_719_0, i_10_483_800_0, i_10_483_1030_0,
    i_10_483_1038_0, i_10_483_1041_0, i_10_483_1043_0, i_10_483_1052_0,
    i_10_483_1053_0, i_10_483_1060_0, i_10_483_1061_0, i_10_483_1084_0,
    i_10_483_1269_0, i_10_483_1308_0, i_10_483_1311_0, i_10_483_1312_0,
    i_10_483_1394_0, i_10_483_1435_0, i_10_483_1439_0, i_10_483_1444_0,
    i_10_483_1539_0, i_10_483_1540_0, i_10_483_1577_0, i_10_483_1624_0,
    i_10_483_1652_0, i_10_483_1654_0, i_10_483_1686_0, i_10_483_1687_0,
    i_10_483_1689_0, i_10_483_1765_0, i_10_483_1769_0, i_10_483_1819_0,
    i_10_483_1824_0, i_10_483_1915_0, i_10_483_1999_0, i_10_483_2001_0,
    i_10_483_2159_0, i_10_483_2349_0, i_10_483_2352_0, i_10_483_2355_0,
    i_10_483_2357_0, i_10_483_2365_0, i_10_483_2376_0, i_10_483_2378_0,
    i_10_483_2405_0, i_10_483_2406_0, i_10_483_2454_0, i_10_483_2456_0,
    i_10_483_2470_0, i_10_483_2516_0, i_10_483_2564_0, i_10_483_2604_0,
    i_10_483_2632_0, i_10_483_2644_0, i_10_483_2677_0, i_10_483_2699_0,
    i_10_483_2714_0, i_10_483_2956_0, i_10_483_2959_0, i_10_483_2980_0,
    i_10_483_2982_0, i_10_483_2983_0, i_10_483_2984_0, i_10_483_2985_0,
    i_10_483_3036_0, i_10_483_3268_0, i_10_483_3272_0, i_10_483_3278_0,
    i_10_483_3297_0, i_10_483_3384_0, i_10_483_3385_0, i_10_483_3388_0,
    i_10_483_3389_0, i_10_483_3472_0, i_10_483_3617_0, i_10_483_3645_0,
    i_10_483_3649_0, i_10_483_3784_0, i_10_483_3785_0, i_10_483_3834_0,
    i_10_483_3852_0, i_10_483_4009_0, i_10_483_4114_0, i_10_483_4125_0,
    i_10_483_4130_0, i_10_483_4170_0, i_10_483_4173_0, i_10_483_4174_0,
    i_10_483_4267_0, i_10_483_4271_0, i_10_483_4278_0, i_10_483_4279_0;
  output o_10_483_0_0;
  assign o_10_483_0_0 = 0;
endmodule



// Benchmark "kernel_10_484" written by ABC on Sun Jul 19 10:29:30 2020

module kernel_10_484 ( 
    i_10_484_176_0, i_10_484_284_0, i_10_484_405_0, i_10_484_406_0,
    i_10_484_409_0, i_10_484_459_0, i_10_484_747_0, i_10_484_999_0,
    i_10_484_1000_0, i_10_484_1027_0, i_10_484_1139_0, i_10_484_1141_0,
    i_10_484_1234_0, i_10_484_1238_0, i_10_484_1432_0, i_10_484_1489_0,
    i_10_484_1539_0, i_10_484_1575_0, i_10_484_1576_0, i_10_484_1578_0,
    i_10_484_1647_0, i_10_484_1650_0, i_10_484_1651_0, i_10_484_1691_0,
    i_10_484_1909_0, i_10_484_1945_0, i_10_484_1951_0, i_10_484_2017_0,
    i_10_484_2151_0, i_10_484_2178_0, i_10_484_2179_0, i_10_484_2181_0,
    i_10_484_2185_0, i_10_484_2196_0, i_10_484_2197_0, i_10_484_2199_0,
    i_10_484_2305_0, i_10_484_2306_0, i_10_484_2349_0, i_10_484_2350_0,
    i_10_484_2351_0, i_10_484_2352_0, i_10_484_2353_0, i_10_484_2355_0,
    i_10_484_2377_0, i_10_484_2406_0, i_10_484_2469_0, i_10_484_2662_0,
    i_10_484_2700_0, i_10_484_2711_0, i_10_484_2712_0, i_10_484_2714_0,
    i_10_484_2724_0, i_10_484_2833_0, i_10_484_2887_0, i_10_484_2916_0,
    i_10_484_2917_0, i_10_484_2919_0, i_10_484_2923_0, i_10_484_2954_0,
    i_10_484_2979_0, i_10_484_3069_0, i_10_484_3150_0, i_10_484_3267_0,
    i_10_484_3268_0, i_10_484_3270_0, i_10_484_3271_0, i_10_484_3280_0,
    i_10_484_3330_0, i_10_484_3385_0, i_10_484_3387_0, i_10_484_3522_0,
    i_10_484_3525_0, i_10_484_3526_0, i_10_484_3584_0, i_10_484_3585_0,
    i_10_484_3587_0, i_10_484_3614_0, i_10_484_3615_0, i_10_484_3616_0,
    i_10_484_3617_0, i_10_484_3645_0, i_10_484_3649_0, i_10_484_3685_0,
    i_10_484_3807_0, i_10_484_3837_0, i_10_484_3838_0, i_10_484_3852_0,
    i_10_484_3889_0, i_10_484_3907_0, i_10_484_3980_0, i_10_484_3984_0,
    i_10_484_4266_0, i_10_484_4268_0, i_10_484_4271_0, i_10_484_4275_0,
    i_10_484_4276_0, i_10_484_4287_0, i_10_484_4567_0, i_10_484_4568_0,
    o_10_484_0_0  );
  input  i_10_484_176_0, i_10_484_284_0, i_10_484_405_0, i_10_484_406_0,
    i_10_484_409_0, i_10_484_459_0, i_10_484_747_0, i_10_484_999_0,
    i_10_484_1000_0, i_10_484_1027_0, i_10_484_1139_0, i_10_484_1141_0,
    i_10_484_1234_0, i_10_484_1238_0, i_10_484_1432_0, i_10_484_1489_0,
    i_10_484_1539_0, i_10_484_1575_0, i_10_484_1576_0, i_10_484_1578_0,
    i_10_484_1647_0, i_10_484_1650_0, i_10_484_1651_0, i_10_484_1691_0,
    i_10_484_1909_0, i_10_484_1945_0, i_10_484_1951_0, i_10_484_2017_0,
    i_10_484_2151_0, i_10_484_2178_0, i_10_484_2179_0, i_10_484_2181_0,
    i_10_484_2185_0, i_10_484_2196_0, i_10_484_2197_0, i_10_484_2199_0,
    i_10_484_2305_0, i_10_484_2306_0, i_10_484_2349_0, i_10_484_2350_0,
    i_10_484_2351_0, i_10_484_2352_0, i_10_484_2353_0, i_10_484_2355_0,
    i_10_484_2377_0, i_10_484_2406_0, i_10_484_2469_0, i_10_484_2662_0,
    i_10_484_2700_0, i_10_484_2711_0, i_10_484_2712_0, i_10_484_2714_0,
    i_10_484_2724_0, i_10_484_2833_0, i_10_484_2887_0, i_10_484_2916_0,
    i_10_484_2917_0, i_10_484_2919_0, i_10_484_2923_0, i_10_484_2954_0,
    i_10_484_2979_0, i_10_484_3069_0, i_10_484_3150_0, i_10_484_3267_0,
    i_10_484_3268_0, i_10_484_3270_0, i_10_484_3271_0, i_10_484_3280_0,
    i_10_484_3330_0, i_10_484_3385_0, i_10_484_3387_0, i_10_484_3522_0,
    i_10_484_3525_0, i_10_484_3526_0, i_10_484_3584_0, i_10_484_3585_0,
    i_10_484_3587_0, i_10_484_3614_0, i_10_484_3615_0, i_10_484_3616_0,
    i_10_484_3617_0, i_10_484_3645_0, i_10_484_3649_0, i_10_484_3685_0,
    i_10_484_3807_0, i_10_484_3837_0, i_10_484_3838_0, i_10_484_3852_0,
    i_10_484_3889_0, i_10_484_3907_0, i_10_484_3980_0, i_10_484_3984_0,
    i_10_484_4266_0, i_10_484_4268_0, i_10_484_4271_0, i_10_484_4275_0,
    i_10_484_4276_0, i_10_484_4287_0, i_10_484_4567_0, i_10_484_4568_0;
  output o_10_484_0_0;
  assign o_10_484_0_0 = ~((~i_10_484_2196_0 & ((~i_10_484_2179_0 & ((~i_10_484_2185_0 & ((~i_10_484_405_0 & ((~i_10_484_999_0 & ~i_10_484_1575_0 & ~i_10_484_1945_0 & ~i_10_484_2305_0 & ~i_10_484_2469_0 & ~i_10_484_3889_0 & ~i_10_484_3907_0 & ~i_10_484_3984_0) | (~i_10_484_1576_0 & ~i_10_484_3069_0 & ~i_10_484_3649_0 & ~i_10_484_3685_0 & ~i_10_484_4266_0))) | (~i_10_484_2181_0 & ~i_10_484_2350_0 & ~i_10_484_2352_0 & ~i_10_484_3069_0 & ~i_10_484_4275_0))) | (~i_10_484_1945_0 & ~i_10_484_2181_0 & ~i_10_484_2352_0 & ~i_10_484_2377_0 & ~i_10_484_3271_0 & ~i_10_484_3837_0))) | (~i_10_484_459_0 & ~i_10_484_1027_0 & ~i_10_484_1539_0 & ~i_10_484_1945_0 & ~i_10_484_2349_0 & ~i_10_484_2406_0 & ~i_10_484_3271_0 & ~i_10_484_3526_0) | (i_10_484_1234_0 & ~i_10_484_2178_0 & ~i_10_484_2923_0 & ~i_10_484_2979_0 & ~i_10_484_3069_0 & ~i_10_484_3385_0 & ~i_10_484_4276_0) | (~i_10_484_176_0 & i_10_484_1238_0 & ~i_10_484_1575_0 & ~i_10_484_2185_0 & ~i_10_484_3268_0 & ~i_10_484_4287_0))) | (~i_10_484_999_0 & ((~i_10_484_1000_0 & ((~i_10_484_1539_0 & ~i_10_484_2181_0 & ~i_10_484_2306_0 & ~i_10_484_2350_0 & ~i_10_484_2351_0 & ~i_10_484_2353_0 & ~i_10_484_2355_0 & ~i_10_484_2979_0 & ~i_10_484_3069_0 & ~i_10_484_3615_0) | (~i_10_484_1575_0 & ~i_10_484_1576_0 & ~i_10_484_1578_0 & ~i_10_484_2349_0 & ~i_10_484_3271_0 & ~i_10_484_4568_0))) | (~i_10_484_1539_0 & ~i_10_484_3645_0 & ((~i_10_484_1027_0 & ~i_10_484_1578_0 & ~i_10_484_1945_0 & ~i_10_484_1951_0 & ~i_10_484_2377_0 & ~i_10_484_3280_0 & ~i_10_484_4275_0 & ~i_10_484_4276_0) | (~i_10_484_459_0 & ~i_10_484_2017_0 & ~i_10_484_2179_0 & ~i_10_484_2700_0 & i_10_484_2923_0 & ~i_10_484_3614_0 & ~i_10_484_4568_0))) | (~i_10_484_2349_0 & ((~i_10_484_1575_0 & ((i_10_484_1238_0 & ~i_10_484_2662_0) | (~i_10_484_747_0 & ~i_10_484_2351_0 & ~i_10_484_3837_0 & ~i_10_484_3984_0))) | (~i_10_484_1238_0 & ~i_10_484_1945_0 & ~i_10_484_2178_0 & ~i_10_484_2199_0 & ~i_10_484_3069_0 & ~i_10_484_3271_0 & ~i_10_484_3280_0 & ~i_10_484_4271_0 & ~i_10_484_4275_0))))) | (~i_10_484_1647_0 & ((~i_10_484_1575_0 & ~i_10_484_2185_0 & ~i_10_484_2923_0 & ~i_10_484_3270_0 & ~i_10_484_3280_0 & ~i_10_484_3838_0 & ~i_10_484_3980_0) | (~i_10_484_1539_0 & i_10_484_2724_0 & ~i_10_484_3587_0 & ~i_10_484_4268_0))) | (~i_10_484_1539_0 & ((~i_10_484_1238_0 & ~i_10_484_1576_0 & ~i_10_484_2179_0 & ~i_10_484_2350_0 & i_10_484_3616_0 & i_10_484_3852_0) | (~i_10_484_1951_0 & ~i_10_484_2197_0 & ~i_10_484_2199_0 & ~i_10_484_2919_0 & ~i_10_484_4275_0 & ~i_10_484_4567_0))) | (~i_10_484_2178_0 & ~i_10_484_2181_0 & ~i_10_484_2197_0 & ~i_10_484_2305_0 & ~i_10_484_3271_0 & i_10_484_3980_0 & ~i_10_484_4287_0));
endmodule



// Benchmark "kernel_10_485" written by ABC on Sun Jul 19 10:29:30 2020

module kernel_10_485 ( 
    i_10_485_28_0, i_10_485_45_0, i_10_485_223_0, i_10_485_254_0,
    i_10_485_290_0, i_10_485_299_0, i_10_485_389_0, i_10_485_424_0,
    i_10_485_425_0, i_10_485_434_0, i_10_485_462_0, i_10_485_740_0,
    i_10_485_1003_0, i_10_485_1027_0, i_10_485_1028_0, i_10_485_1034_0,
    i_10_485_1055_0, i_10_485_1082_0, i_10_485_1118_0, i_10_485_1233_0,
    i_10_485_1235_0, i_10_485_1236_0, i_10_485_1238_0, i_10_485_1243_0,
    i_10_485_1244_0, i_10_485_1342_0, i_10_485_1379_0, i_10_485_1541_0,
    i_10_485_1552_0, i_10_485_1577_0, i_10_485_1625_0, i_10_485_1651_0,
    i_10_485_1683_0, i_10_485_1687_0, i_10_485_1710_0, i_10_485_1711_0,
    i_10_485_1914_0, i_10_485_2036_0, i_10_485_2090_0, i_10_485_2179_0,
    i_10_485_2180_0, i_10_485_2200_0, i_10_485_2306_0, i_10_485_2332_0,
    i_10_485_2353_0, i_10_485_2354_0, i_10_485_2359_0, i_10_485_2360_0,
    i_10_485_2362_0, i_10_485_2379_0, i_10_485_2448_0, i_10_485_2451_0,
    i_10_485_2452_0, i_10_485_2456_0, i_10_485_2468_0, i_10_485_2470_0,
    i_10_485_2471_0, i_10_485_2542_0, i_10_485_2653_0, i_10_485_2673_0,
    i_10_485_2713_0, i_10_485_2731_0, i_10_485_2838_0, i_10_485_2920_0,
    i_10_485_2958_0, i_10_485_3070_0, i_10_485_3200_0, i_10_485_3278_0,
    i_10_485_3280_0, i_10_485_3281_0, i_10_485_3403_0, i_10_485_3467_0,
    i_10_485_3548_0, i_10_485_3590_0, i_10_485_3612_0, i_10_485_3649_0,
    i_10_485_3650_0, i_10_485_3683_0, i_10_485_3772_0, i_10_485_3781_0,
    i_10_485_3784_0, i_10_485_3785_0, i_10_485_3835_0, i_10_485_3858_0,
    i_10_485_3859_0, i_10_485_3860_0, i_10_485_3881_0, i_10_485_3907_0,
    i_10_485_3982_0, i_10_485_4114_0, i_10_485_4115_0, i_10_485_4205_0,
    i_10_485_4213_0, i_10_485_4214_0, i_10_485_4217_0, i_10_485_4220_0,
    i_10_485_4270_0, i_10_485_4287_0, i_10_485_4430_0, i_10_485_4529_0,
    o_10_485_0_0  );
  input  i_10_485_28_0, i_10_485_45_0, i_10_485_223_0, i_10_485_254_0,
    i_10_485_290_0, i_10_485_299_0, i_10_485_389_0, i_10_485_424_0,
    i_10_485_425_0, i_10_485_434_0, i_10_485_462_0, i_10_485_740_0,
    i_10_485_1003_0, i_10_485_1027_0, i_10_485_1028_0, i_10_485_1034_0,
    i_10_485_1055_0, i_10_485_1082_0, i_10_485_1118_0, i_10_485_1233_0,
    i_10_485_1235_0, i_10_485_1236_0, i_10_485_1238_0, i_10_485_1243_0,
    i_10_485_1244_0, i_10_485_1342_0, i_10_485_1379_0, i_10_485_1541_0,
    i_10_485_1552_0, i_10_485_1577_0, i_10_485_1625_0, i_10_485_1651_0,
    i_10_485_1683_0, i_10_485_1687_0, i_10_485_1710_0, i_10_485_1711_0,
    i_10_485_1914_0, i_10_485_2036_0, i_10_485_2090_0, i_10_485_2179_0,
    i_10_485_2180_0, i_10_485_2200_0, i_10_485_2306_0, i_10_485_2332_0,
    i_10_485_2353_0, i_10_485_2354_0, i_10_485_2359_0, i_10_485_2360_0,
    i_10_485_2362_0, i_10_485_2379_0, i_10_485_2448_0, i_10_485_2451_0,
    i_10_485_2452_0, i_10_485_2456_0, i_10_485_2468_0, i_10_485_2470_0,
    i_10_485_2471_0, i_10_485_2542_0, i_10_485_2653_0, i_10_485_2673_0,
    i_10_485_2713_0, i_10_485_2731_0, i_10_485_2838_0, i_10_485_2920_0,
    i_10_485_2958_0, i_10_485_3070_0, i_10_485_3200_0, i_10_485_3278_0,
    i_10_485_3280_0, i_10_485_3281_0, i_10_485_3403_0, i_10_485_3467_0,
    i_10_485_3548_0, i_10_485_3590_0, i_10_485_3612_0, i_10_485_3649_0,
    i_10_485_3650_0, i_10_485_3683_0, i_10_485_3772_0, i_10_485_3781_0,
    i_10_485_3784_0, i_10_485_3785_0, i_10_485_3835_0, i_10_485_3858_0,
    i_10_485_3859_0, i_10_485_3860_0, i_10_485_3881_0, i_10_485_3907_0,
    i_10_485_3982_0, i_10_485_4114_0, i_10_485_4115_0, i_10_485_4205_0,
    i_10_485_4213_0, i_10_485_4214_0, i_10_485_4217_0, i_10_485_4220_0,
    i_10_485_4270_0, i_10_485_4287_0, i_10_485_4430_0, i_10_485_4529_0;
  output o_10_485_0_0;
  assign o_10_485_0_0 = 0;
endmodule



// Benchmark "kernel_10_486" written by ABC on Sun Jul 19 10:29:31 2020

module kernel_10_486 ( 
    i_10_486_48_0, i_10_486_144_0, i_10_486_145_0, i_10_486_172_0,
    i_10_486_220_0, i_10_486_261_0, i_10_486_263_0, i_10_486_280_0,
    i_10_486_281_0, i_10_486_285_0, i_10_486_287_0, i_10_486_327_0,
    i_10_486_390_0, i_10_486_406_0, i_10_486_409_0, i_10_486_442_0,
    i_10_486_445_0, i_10_486_461_0, i_10_486_467_0, i_10_486_586_0,
    i_10_486_711_0, i_10_486_712_0, i_10_486_793_0, i_10_486_795_0,
    i_10_486_798_0, i_10_486_799_0, i_10_486_955_0, i_10_486_1237_0,
    i_10_486_1240_0, i_10_486_1266_0, i_10_486_1312_0, i_10_486_1313_0,
    i_10_486_1365_0, i_10_486_1539_0, i_10_486_1553_0, i_10_486_1651_0,
    i_10_486_1685_0, i_10_486_1686_0, i_10_486_1801_0, i_10_486_1802_0,
    i_10_486_1818_0, i_10_486_1825_0, i_10_486_1913_0, i_10_486_1998_0,
    i_10_486_2025_0, i_10_486_2206_0, i_10_486_2223_0, i_10_486_2224_0,
    i_10_486_2356_0, i_10_486_2361_0, i_10_486_2469_0, i_10_486_2471_0,
    i_10_486_2473_0, i_10_486_2601_0, i_10_486_2634_0, i_10_486_2635_0,
    i_10_486_2677_0, i_10_486_2703_0, i_10_486_2704_0, i_10_486_2722_0,
    i_10_486_2723_0, i_10_486_2727_0, i_10_486_2729_0, i_10_486_2731_0,
    i_10_486_2829_0, i_10_486_3034_0, i_10_486_3231_0, i_10_486_3234_0,
    i_10_486_3267_0, i_10_486_3268_0, i_10_486_3277_0, i_10_486_3384_0,
    i_10_486_3391_0, i_10_486_3496_0, i_10_486_3501_0, i_10_486_3507_0,
    i_10_486_3519_0, i_10_486_3522_0, i_10_486_3523_0, i_10_486_3524_0,
    i_10_486_3583_0, i_10_486_3587_0, i_10_486_3588_0, i_10_486_3590_0,
    i_10_486_3783_0, i_10_486_3785_0, i_10_486_3788_0, i_10_486_3834_0,
    i_10_486_3837_0, i_10_486_3838_0, i_10_486_3839_0, i_10_486_3846_0,
    i_10_486_3848_0, i_10_486_3855_0, i_10_486_4114_0, i_10_486_4213_0,
    i_10_486_4269_0, i_10_486_4275_0, i_10_486_4276_0, i_10_486_4289_0,
    o_10_486_0_0  );
  input  i_10_486_48_0, i_10_486_144_0, i_10_486_145_0, i_10_486_172_0,
    i_10_486_220_0, i_10_486_261_0, i_10_486_263_0, i_10_486_280_0,
    i_10_486_281_0, i_10_486_285_0, i_10_486_287_0, i_10_486_327_0,
    i_10_486_390_0, i_10_486_406_0, i_10_486_409_0, i_10_486_442_0,
    i_10_486_445_0, i_10_486_461_0, i_10_486_467_0, i_10_486_586_0,
    i_10_486_711_0, i_10_486_712_0, i_10_486_793_0, i_10_486_795_0,
    i_10_486_798_0, i_10_486_799_0, i_10_486_955_0, i_10_486_1237_0,
    i_10_486_1240_0, i_10_486_1266_0, i_10_486_1312_0, i_10_486_1313_0,
    i_10_486_1365_0, i_10_486_1539_0, i_10_486_1553_0, i_10_486_1651_0,
    i_10_486_1685_0, i_10_486_1686_0, i_10_486_1801_0, i_10_486_1802_0,
    i_10_486_1818_0, i_10_486_1825_0, i_10_486_1913_0, i_10_486_1998_0,
    i_10_486_2025_0, i_10_486_2206_0, i_10_486_2223_0, i_10_486_2224_0,
    i_10_486_2356_0, i_10_486_2361_0, i_10_486_2469_0, i_10_486_2471_0,
    i_10_486_2473_0, i_10_486_2601_0, i_10_486_2634_0, i_10_486_2635_0,
    i_10_486_2677_0, i_10_486_2703_0, i_10_486_2704_0, i_10_486_2722_0,
    i_10_486_2723_0, i_10_486_2727_0, i_10_486_2729_0, i_10_486_2731_0,
    i_10_486_2829_0, i_10_486_3034_0, i_10_486_3231_0, i_10_486_3234_0,
    i_10_486_3267_0, i_10_486_3268_0, i_10_486_3277_0, i_10_486_3384_0,
    i_10_486_3391_0, i_10_486_3496_0, i_10_486_3501_0, i_10_486_3507_0,
    i_10_486_3519_0, i_10_486_3522_0, i_10_486_3523_0, i_10_486_3524_0,
    i_10_486_3583_0, i_10_486_3587_0, i_10_486_3588_0, i_10_486_3590_0,
    i_10_486_3783_0, i_10_486_3785_0, i_10_486_3788_0, i_10_486_3834_0,
    i_10_486_3837_0, i_10_486_3838_0, i_10_486_3839_0, i_10_486_3846_0,
    i_10_486_3848_0, i_10_486_3855_0, i_10_486_4114_0, i_10_486_4213_0,
    i_10_486_4269_0, i_10_486_4275_0, i_10_486_4276_0, i_10_486_4289_0;
  output o_10_486_0_0;
  assign o_10_486_0_0 = 0;
endmodule



// Benchmark "kernel_10_487" written by ABC on Sun Jul 19 10:29:32 2020

module kernel_10_487 ( 
    i_10_487_28_0, i_10_487_70_0, i_10_487_118_0, i_10_487_175_0,
    i_10_487_176_0, i_10_487_260_0, i_10_487_315_0, i_10_487_327_0,
    i_10_487_387_0, i_10_487_391_0, i_10_487_443_0, i_10_487_461_0,
    i_10_487_514_0, i_10_487_797_0, i_10_487_799_0, i_10_487_800_0,
    i_10_487_897_0, i_10_487_899_0, i_10_487_971_0, i_10_487_1240_0,
    i_10_487_1241_0, i_10_487_1243_0, i_10_487_1246_0, i_10_487_1311_0,
    i_10_487_1348_0, i_10_487_1434_0, i_10_487_1539_0, i_10_487_1543_0,
    i_10_487_1549_0, i_10_487_1552_0, i_10_487_1630_0, i_10_487_1650_0,
    i_10_487_1651_0, i_10_487_1686_0, i_10_487_1690_0, i_10_487_1821_0,
    i_10_487_1822_0, i_10_487_1823_0, i_10_487_1913_0, i_10_487_1945_0,
    i_10_487_1949_0, i_10_487_1996_0, i_10_487_2365_0, i_10_487_2404_0,
    i_10_487_2448_0, i_10_487_2449_0, i_10_487_2453_0, i_10_487_2456_0,
    i_10_487_2471_0, i_10_487_2518_0, i_10_487_2660_0, i_10_487_2663_0,
    i_10_487_2708_0, i_10_487_2716_0, i_10_487_2717_0, i_10_487_2723_0,
    i_10_487_2732_0, i_10_487_2733_0, i_10_487_2787_0, i_10_487_2788_0,
    i_10_487_2831_0, i_10_487_2833_0, i_10_487_3033_0, i_10_487_3034_0,
    i_10_487_3036_0, i_10_487_3041_0, i_10_487_3045_0, i_10_487_3199_0,
    i_10_487_3238_0, i_10_487_3269_0, i_10_487_3390_0, i_10_487_3409_0,
    i_10_487_3437_0, i_10_487_3526_0, i_10_487_3613_0, i_10_487_3616_0,
    i_10_487_3617_0, i_10_487_3640_0, i_10_487_3649_0, i_10_487_3650_0,
    i_10_487_3653_0, i_10_487_3781_0, i_10_487_3782_0, i_10_487_3787_0,
    i_10_487_3811_0, i_10_487_3839_0, i_10_487_3840_0, i_10_487_3856_0,
    i_10_487_3857_0, i_10_487_3860_0, i_10_487_3882_0, i_10_487_3949_0,
    i_10_487_3991_0, i_10_487_4025_0, i_10_487_4056_0, i_10_487_4267_0,
    i_10_487_4270_0, i_10_487_4276_0, i_10_487_4283_0, i_10_487_4291_0,
    o_10_487_0_0  );
  input  i_10_487_28_0, i_10_487_70_0, i_10_487_118_0, i_10_487_175_0,
    i_10_487_176_0, i_10_487_260_0, i_10_487_315_0, i_10_487_327_0,
    i_10_487_387_0, i_10_487_391_0, i_10_487_443_0, i_10_487_461_0,
    i_10_487_514_0, i_10_487_797_0, i_10_487_799_0, i_10_487_800_0,
    i_10_487_897_0, i_10_487_899_0, i_10_487_971_0, i_10_487_1240_0,
    i_10_487_1241_0, i_10_487_1243_0, i_10_487_1246_0, i_10_487_1311_0,
    i_10_487_1348_0, i_10_487_1434_0, i_10_487_1539_0, i_10_487_1543_0,
    i_10_487_1549_0, i_10_487_1552_0, i_10_487_1630_0, i_10_487_1650_0,
    i_10_487_1651_0, i_10_487_1686_0, i_10_487_1690_0, i_10_487_1821_0,
    i_10_487_1822_0, i_10_487_1823_0, i_10_487_1913_0, i_10_487_1945_0,
    i_10_487_1949_0, i_10_487_1996_0, i_10_487_2365_0, i_10_487_2404_0,
    i_10_487_2448_0, i_10_487_2449_0, i_10_487_2453_0, i_10_487_2456_0,
    i_10_487_2471_0, i_10_487_2518_0, i_10_487_2660_0, i_10_487_2663_0,
    i_10_487_2708_0, i_10_487_2716_0, i_10_487_2717_0, i_10_487_2723_0,
    i_10_487_2732_0, i_10_487_2733_0, i_10_487_2787_0, i_10_487_2788_0,
    i_10_487_2831_0, i_10_487_2833_0, i_10_487_3033_0, i_10_487_3034_0,
    i_10_487_3036_0, i_10_487_3041_0, i_10_487_3045_0, i_10_487_3199_0,
    i_10_487_3238_0, i_10_487_3269_0, i_10_487_3390_0, i_10_487_3409_0,
    i_10_487_3437_0, i_10_487_3526_0, i_10_487_3613_0, i_10_487_3616_0,
    i_10_487_3617_0, i_10_487_3640_0, i_10_487_3649_0, i_10_487_3650_0,
    i_10_487_3653_0, i_10_487_3781_0, i_10_487_3782_0, i_10_487_3787_0,
    i_10_487_3811_0, i_10_487_3839_0, i_10_487_3840_0, i_10_487_3856_0,
    i_10_487_3857_0, i_10_487_3860_0, i_10_487_3882_0, i_10_487_3949_0,
    i_10_487_3991_0, i_10_487_4025_0, i_10_487_4056_0, i_10_487_4267_0,
    i_10_487_4270_0, i_10_487_4276_0, i_10_487_4283_0, i_10_487_4291_0;
  output o_10_487_0_0;
  assign o_10_487_0_0 = 0;
endmodule



// Benchmark "kernel_10_488" written by ABC on Sun Jul 19 10:29:33 2020

module kernel_10_488 ( 
    i_10_488_139_0, i_10_488_279_0, i_10_488_280_0, i_10_488_361_0,
    i_10_488_441_0, i_10_488_442_0, i_10_488_461_0, i_10_488_496_0,
    i_10_488_585_0, i_10_488_748_0, i_10_488_749_0, i_10_488_754_0,
    i_10_488_792_0, i_10_488_795_0, i_10_488_796_0, i_10_488_828_0,
    i_10_488_830_0, i_10_488_924_0, i_10_488_955_0, i_10_488_983_0,
    i_10_488_1163_0, i_10_488_1239_0, i_10_488_1243_0, i_10_488_1264_0,
    i_10_488_1492_0, i_10_488_1540_0, i_10_488_1629_0, i_10_488_1630_0,
    i_10_488_1631_0, i_10_488_1635_0, i_10_488_1636_0, i_10_488_1644_0,
    i_10_488_1645_0, i_10_488_1654_0, i_10_488_1655_0, i_10_488_1683_0,
    i_10_488_1684_0, i_10_488_1720_0, i_10_488_1801_0, i_10_488_1802_0,
    i_10_488_1818_0, i_10_488_1819_0, i_10_488_2004_0, i_10_488_2005_0,
    i_10_488_2006_0, i_10_488_2031_0, i_10_488_2032_0, i_10_488_2206_0,
    i_10_488_2241_0, i_10_488_2248_0, i_10_488_2386_0, i_10_488_2387_0,
    i_10_488_2472_0, i_10_488_2473_0, i_10_488_2474_0, i_10_488_2539_0,
    i_10_488_2660_0, i_10_488_2661_0, i_10_488_2663_0, i_10_488_2674_0,
    i_10_488_2681_0, i_10_488_2717_0, i_10_488_2733_0, i_10_488_2743_0,
    i_10_488_2817_0, i_10_488_2824_0, i_10_488_2922_0, i_10_488_2979_0,
    i_10_488_2980_0, i_10_488_2982_0, i_10_488_2983_0, i_10_488_2985_0,
    i_10_488_2986_0, i_10_488_3237_0, i_10_488_3238_0, i_10_488_3282_0,
    i_10_488_3283_0, i_10_488_3313_0, i_10_488_3465_0, i_10_488_3493_0,
    i_10_488_3508_0, i_10_488_3520_0, i_10_488_3525_0, i_10_488_3724_0,
    i_10_488_3798_0, i_10_488_3854_0, i_10_488_3912_0, i_10_488_3948_0,
    i_10_488_3949_0, i_10_488_4061_0, i_10_488_4115_0, i_10_488_4269_0,
    i_10_488_4272_0, i_10_488_4284_0, i_10_488_4302_0, i_10_488_4303_0,
    i_10_488_4457_0, i_10_488_4459_0, i_10_488_4582_0, i_10_488_4583_0,
    o_10_488_0_0  );
  input  i_10_488_139_0, i_10_488_279_0, i_10_488_280_0, i_10_488_361_0,
    i_10_488_441_0, i_10_488_442_0, i_10_488_461_0, i_10_488_496_0,
    i_10_488_585_0, i_10_488_748_0, i_10_488_749_0, i_10_488_754_0,
    i_10_488_792_0, i_10_488_795_0, i_10_488_796_0, i_10_488_828_0,
    i_10_488_830_0, i_10_488_924_0, i_10_488_955_0, i_10_488_983_0,
    i_10_488_1163_0, i_10_488_1239_0, i_10_488_1243_0, i_10_488_1264_0,
    i_10_488_1492_0, i_10_488_1540_0, i_10_488_1629_0, i_10_488_1630_0,
    i_10_488_1631_0, i_10_488_1635_0, i_10_488_1636_0, i_10_488_1644_0,
    i_10_488_1645_0, i_10_488_1654_0, i_10_488_1655_0, i_10_488_1683_0,
    i_10_488_1684_0, i_10_488_1720_0, i_10_488_1801_0, i_10_488_1802_0,
    i_10_488_1818_0, i_10_488_1819_0, i_10_488_2004_0, i_10_488_2005_0,
    i_10_488_2006_0, i_10_488_2031_0, i_10_488_2032_0, i_10_488_2206_0,
    i_10_488_2241_0, i_10_488_2248_0, i_10_488_2386_0, i_10_488_2387_0,
    i_10_488_2472_0, i_10_488_2473_0, i_10_488_2474_0, i_10_488_2539_0,
    i_10_488_2660_0, i_10_488_2661_0, i_10_488_2663_0, i_10_488_2674_0,
    i_10_488_2681_0, i_10_488_2717_0, i_10_488_2733_0, i_10_488_2743_0,
    i_10_488_2817_0, i_10_488_2824_0, i_10_488_2922_0, i_10_488_2979_0,
    i_10_488_2980_0, i_10_488_2982_0, i_10_488_2983_0, i_10_488_2985_0,
    i_10_488_2986_0, i_10_488_3237_0, i_10_488_3238_0, i_10_488_3282_0,
    i_10_488_3283_0, i_10_488_3313_0, i_10_488_3465_0, i_10_488_3493_0,
    i_10_488_3508_0, i_10_488_3520_0, i_10_488_3525_0, i_10_488_3724_0,
    i_10_488_3798_0, i_10_488_3854_0, i_10_488_3912_0, i_10_488_3948_0,
    i_10_488_3949_0, i_10_488_4061_0, i_10_488_4115_0, i_10_488_4269_0,
    i_10_488_4272_0, i_10_488_4284_0, i_10_488_4302_0, i_10_488_4303_0,
    i_10_488_4457_0, i_10_488_4459_0, i_10_488_4582_0, i_10_488_4583_0;
  output o_10_488_0_0;
  assign o_10_488_0_0 = 0;
endmodule



// Benchmark "kernel_10_489" written by ABC on Sun Jul 19 10:29:34 2020

module kernel_10_489 ( 
    i_10_489_23_0, i_10_489_137_0, i_10_489_271_0, i_10_489_272_0,
    i_10_489_274_0, i_10_489_275_0, i_10_489_286_0, i_10_489_287_0,
    i_10_489_317_0, i_10_489_388_0, i_10_489_461_0, i_10_489_506_0,
    i_10_489_641_0, i_10_489_692_0, i_10_489_715_0, i_10_489_752_0,
    i_10_489_799_0, i_10_489_821_0, i_10_489_831_0, i_10_489_1157_0,
    i_10_489_1171_0, i_10_489_1209_0, i_10_489_1210_0, i_10_489_1240_0,
    i_10_489_1243_0, i_10_489_1245_0, i_10_489_1308_0, i_10_489_1312_0,
    i_10_489_1328_0, i_10_489_1432_0, i_10_489_1450_0, i_10_489_1522_0,
    i_10_489_1531_0, i_10_489_1534_0, i_10_489_1535_0, i_10_489_1544_0,
    i_10_489_1580_0, i_10_489_1603_0, i_10_489_1622_0, i_10_489_1633_0,
    i_10_489_1688_0, i_10_489_1693_0, i_10_489_1711_0, i_10_489_1717_0,
    i_10_489_1718_0, i_10_489_1805_0, i_10_489_1822_0, i_10_489_1826_0,
    i_10_489_1981_0, i_10_489_2028_0, i_10_489_2029_0, i_10_489_2110_0,
    i_10_489_2113_0, i_10_489_2181_0, i_10_489_2209_0, i_10_489_2228_0,
    i_10_489_2354_0, i_10_489_2376_0, i_10_489_2455_0, i_10_489_2513_0,
    i_10_489_2557_0, i_10_489_2629_0, i_10_489_2632_0, i_10_489_2633_0,
    i_10_489_2665_0, i_10_489_2667_0, i_10_489_2702_0, i_10_489_2704_0,
    i_10_489_2705_0, i_10_489_2714_0, i_10_489_2786_0, i_10_489_2966_0,
    i_10_489_2983_0, i_10_489_3119_0, i_10_489_3166_0, i_10_489_3203_0,
    i_10_489_3296_0, i_10_489_3404_0, i_10_489_3497_0, i_10_489_3500_0,
    i_10_489_3502_0, i_10_489_3538_0, i_10_489_3547_0, i_10_489_3610_0,
    i_10_489_3614_0, i_10_489_3615_0, i_10_489_3688_0, i_10_489_3779_0,
    i_10_489_3808_0, i_10_489_3830_0, i_10_489_3853_0, i_10_489_3854_0,
    i_10_489_3857_0, i_10_489_3859_0, i_10_489_3875_0, i_10_489_4001_0,
    i_10_489_4276_0, i_10_489_4340_0, i_10_489_4456_0, i_10_489_4532_0,
    o_10_489_0_0  );
  input  i_10_489_23_0, i_10_489_137_0, i_10_489_271_0, i_10_489_272_0,
    i_10_489_274_0, i_10_489_275_0, i_10_489_286_0, i_10_489_287_0,
    i_10_489_317_0, i_10_489_388_0, i_10_489_461_0, i_10_489_506_0,
    i_10_489_641_0, i_10_489_692_0, i_10_489_715_0, i_10_489_752_0,
    i_10_489_799_0, i_10_489_821_0, i_10_489_831_0, i_10_489_1157_0,
    i_10_489_1171_0, i_10_489_1209_0, i_10_489_1210_0, i_10_489_1240_0,
    i_10_489_1243_0, i_10_489_1245_0, i_10_489_1308_0, i_10_489_1312_0,
    i_10_489_1328_0, i_10_489_1432_0, i_10_489_1450_0, i_10_489_1522_0,
    i_10_489_1531_0, i_10_489_1534_0, i_10_489_1535_0, i_10_489_1544_0,
    i_10_489_1580_0, i_10_489_1603_0, i_10_489_1622_0, i_10_489_1633_0,
    i_10_489_1688_0, i_10_489_1693_0, i_10_489_1711_0, i_10_489_1717_0,
    i_10_489_1718_0, i_10_489_1805_0, i_10_489_1822_0, i_10_489_1826_0,
    i_10_489_1981_0, i_10_489_2028_0, i_10_489_2029_0, i_10_489_2110_0,
    i_10_489_2113_0, i_10_489_2181_0, i_10_489_2209_0, i_10_489_2228_0,
    i_10_489_2354_0, i_10_489_2376_0, i_10_489_2455_0, i_10_489_2513_0,
    i_10_489_2557_0, i_10_489_2629_0, i_10_489_2632_0, i_10_489_2633_0,
    i_10_489_2665_0, i_10_489_2667_0, i_10_489_2702_0, i_10_489_2704_0,
    i_10_489_2705_0, i_10_489_2714_0, i_10_489_2786_0, i_10_489_2966_0,
    i_10_489_2983_0, i_10_489_3119_0, i_10_489_3166_0, i_10_489_3203_0,
    i_10_489_3296_0, i_10_489_3404_0, i_10_489_3497_0, i_10_489_3500_0,
    i_10_489_3502_0, i_10_489_3538_0, i_10_489_3547_0, i_10_489_3610_0,
    i_10_489_3614_0, i_10_489_3615_0, i_10_489_3688_0, i_10_489_3779_0,
    i_10_489_3808_0, i_10_489_3830_0, i_10_489_3853_0, i_10_489_3854_0,
    i_10_489_3857_0, i_10_489_3859_0, i_10_489_3875_0, i_10_489_4001_0,
    i_10_489_4276_0, i_10_489_4340_0, i_10_489_4456_0, i_10_489_4532_0;
  output o_10_489_0_0;
  assign o_10_489_0_0 = 0;
endmodule



// Benchmark "kernel_10_490" written by ABC on Sun Jul 19 10:29:35 2020

module kernel_10_490 ( 
    i_10_490_34_0, i_10_490_35_0, i_10_490_286_0, i_10_490_315_0,
    i_10_490_319_0, i_10_490_324_0, i_10_490_328_0, i_10_490_330_0,
    i_10_490_393_0, i_10_490_430_0, i_10_490_435_0, i_10_490_438_0,
    i_10_490_439_0, i_10_490_440_0, i_10_490_442_0, i_10_490_457_0,
    i_10_490_516_0, i_10_490_520_0, i_10_490_700_0, i_10_490_951_0,
    i_10_490_996_0, i_10_490_997_0, i_10_490_1006_0, i_10_490_1052_0,
    i_10_490_1138_0, i_10_490_1140_0, i_10_490_1236_0, i_10_490_1237_0,
    i_10_490_1238_0, i_10_490_1250_0, i_10_490_1307_0, i_10_490_1309_0,
    i_10_490_1312_0, i_10_490_1384_0, i_10_490_1385_0, i_10_490_1457_0,
    i_10_490_1554_0, i_10_490_1555_0, i_10_490_1578_0, i_10_490_1600_0,
    i_10_490_1687_0, i_10_490_1688_0, i_10_490_1690_0, i_10_490_1691_0,
    i_10_490_1768_0, i_10_490_1769_0, i_10_490_1815_0, i_10_490_1816_0,
    i_10_490_1825_0, i_10_490_1826_0, i_10_490_2004_0, i_10_490_2310_0,
    i_10_490_2312_0, i_10_490_2350_0, i_10_490_2351_0, i_10_490_2364_0,
    i_10_490_2408_0, i_10_490_2411_0, i_10_490_2464_0, i_10_490_2509_0,
    i_10_490_2510_0, i_10_490_2515_0, i_10_490_2728_0, i_10_490_2831_0,
    i_10_490_2883_0, i_10_490_2887_0, i_10_490_2919_0, i_10_490_2922_0,
    i_10_490_2923_0, i_10_490_2924_0, i_10_490_2959_0, i_10_490_2982_0,
    i_10_490_2983_0, i_10_490_2985_0, i_10_490_2986_0, i_10_490_3093_0,
    i_10_490_3094_0, i_10_490_3156_0, i_10_490_3199_0, i_10_490_3203_0,
    i_10_490_3284_0, i_10_490_3319_0, i_10_490_3389_0, i_10_490_3545_0,
    i_10_490_3613_0, i_10_490_3733_0, i_10_490_3855_0, i_10_490_3857_0,
    i_10_490_3895_0, i_10_490_3981_0, i_10_490_3982_0, i_10_490_3984_0,
    i_10_490_3985_0, i_10_490_3986_0, i_10_490_3992_0, i_10_490_4003_0,
    i_10_490_4217_0, i_10_490_4288_0, i_10_490_4291_0, i_10_490_4292_0,
    o_10_490_0_0  );
  input  i_10_490_34_0, i_10_490_35_0, i_10_490_286_0, i_10_490_315_0,
    i_10_490_319_0, i_10_490_324_0, i_10_490_328_0, i_10_490_330_0,
    i_10_490_393_0, i_10_490_430_0, i_10_490_435_0, i_10_490_438_0,
    i_10_490_439_0, i_10_490_440_0, i_10_490_442_0, i_10_490_457_0,
    i_10_490_516_0, i_10_490_520_0, i_10_490_700_0, i_10_490_951_0,
    i_10_490_996_0, i_10_490_997_0, i_10_490_1006_0, i_10_490_1052_0,
    i_10_490_1138_0, i_10_490_1140_0, i_10_490_1236_0, i_10_490_1237_0,
    i_10_490_1238_0, i_10_490_1250_0, i_10_490_1307_0, i_10_490_1309_0,
    i_10_490_1312_0, i_10_490_1384_0, i_10_490_1385_0, i_10_490_1457_0,
    i_10_490_1554_0, i_10_490_1555_0, i_10_490_1578_0, i_10_490_1600_0,
    i_10_490_1687_0, i_10_490_1688_0, i_10_490_1690_0, i_10_490_1691_0,
    i_10_490_1768_0, i_10_490_1769_0, i_10_490_1815_0, i_10_490_1816_0,
    i_10_490_1825_0, i_10_490_1826_0, i_10_490_2004_0, i_10_490_2310_0,
    i_10_490_2312_0, i_10_490_2350_0, i_10_490_2351_0, i_10_490_2364_0,
    i_10_490_2408_0, i_10_490_2411_0, i_10_490_2464_0, i_10_490_2509_0,
    i_10_490_2510_0, i_10_490_2515_0, i_10_490_2728_0, i_10_490_2831_0,
    i_10_490_2883_0, i_10_490_2887_0, i_10_490_2919_0, i_10_490_2922_0,
    i_10_490_2923_0, i_10_490_2924_0, i_10_490_2959_0, i_10_490_2982_0,
    i_10_490_2983_0, i_10_490_2985_0, i_10_490_2986_0, i_10_490_3093_0,
    i_10_490_3094_0, i_10_490_3156_0, i_10_490_3199_0, i_10_490_3203_0,
    i_10_490_3284_0, i_10_490_3319_0, i_10_490_3389_0, i_10_490_3545_0,
    i_10_490_3613_0, i_10_490_3733_0, i_10_490_3855_0, i_10_490_3857_0,
    i_10_490_3895_0, i_10_490_3981_0, i_10_490_3982_0, i_10_490_3984_0,
    i_10_490_3985_0, i_10_490_3986_0, i_10_490_3992_0, i_10_490_4003_0,
    i_10_490_4217_0, i_10_490_4288_0, i_10_490_4291_0, i_10_490_4292_0;
  output o_10_490_0_0;
  assign o_10_490_0_0 = ~((~i_10_490_328_0 & ((~i_10_490_319_0 & ~i_10_490_1312_0 & ~i_10_490_1555_0 & ~i_10_490_1578_0 & ~i_10_490_1768_0 & ~i_10_490_2411_0 & ~i_10_490_2983_0) | (~i_10_490_439_0 & ~i_10_490_1815_0 & ~i_10_490_1816_0 & ~i_10_490_2510_0 & ~i_10_490_3982_0 & ~i_10_490_3984_0 & ~i_10_490_3986_0))) | (~i_10_490_319_0 & ((~i_10_490_440_0 & ~i_10_490_1554_0 & ~i_10_490_2310_0 & ~i_10_490_2312_0 & ~i_10_490_2728_0 & ~i_10_490_3613_0) | (~i_10_490_996_0 & ~i_10_490_1769_0 & i_10_490_2350_0 & ~i_10_490_2509_0 & ~i_10_490_3895_0))) | (~i_10_490_1816_0 & ((~i_10_490_34_0 & ~i_10_490_2411_0 & ((~i_10_490_435_0 & ~i_10_490_2510_0 & ~i_10_490_2728_0 & ~i_10_490_2883_0 & ~i_10_490_2887_0 & ~i_10_490_2983_0) | (~i_10_490_393_0 & ~i_10_490_440_0 & ~i_10_490_700_0 & ~i_10_490_1578_0 & ~i_10_490_1769_0 & ~i_10_490_2982_0 & ~i_10_490_3857_0))) | (~i_10_490_393_0 & ~i_10_490_997_0 & ~i_10_490_2310_0 & ~i_10_490_2510_0 & ~i_10_490_2831_0 & ~i_10_490_2982_0 & ~i_10_490_3094_0 & ~i_10_490_3199_0 & ~i_10_490_3895_0) | (~i_10_490_435_0 & ~i_10_490_439_0 & ~i_10_490_442_0 & ~i_10_490_516_0 & ~i_10_490_520_0 & ~i_10_490_700_0 & ~i_10_490_1769_0 & ~i_10_490_2986_0 & ~i_10_490_3981_0))) | (~i_10_490_2509_0 & ((~i_10_490_435_0 & ((~i_10_490_996_0 & ~i_10_490_1769_0 & ~i_10_490_330_0 & ~i_10_490_439_0 & ~i_10_490_2887_0 & ~i_10_490_2983_0 & ~i_10_490_1826_0 & ~i_10_490_2408_0) | (i_10_490_286_0 & ~i_10_490_440_0 & ~i_10_490_1307_0 & ~i_10_490_2510_0 & ~i_10_490_3984_0))) | (~i_10_490_996_0 & ((~i_10_490_2728_0 & i_10_490_2923_0 & ~i_10_490_3389_0) | (~i_10_490_315_0 & ~i_10_490_1250_0 & ~i_10_490_2004_0 & ~i_10_490_2312_0 & ~i_10_490_2411_0 & ~i_10_490_2985_0 & ~i_10_490_3093_0 & ~i_10_490_3094_0 & ~i_10_490_3992_0))))) | (~i_10_490_440_0 & ((~i_10_490_996_0 & ~i_10_490_2351_0 & ~i_10_490_2411_0 & ~i_10_490_2983_0 & i_10_490_3855_0 & ~i_10_490_3984_0) | (~i_10_490_1307_0 & ~i_10_490_1578_0 & ~i_10_490_2728_0 & ~i_10_490_2982_0 & ~i_10_490_3389_0 & ~i_10_490_3985_0 & ~i_10_490_3986_0))) | (~i_10_490_3985_0 & ((~i_10_490_35_0 & ~i_10_490_324_0 & ~i_10_490_520_0 & ~i_10_490_2510_0 & ~i_10_490_2982_0 & ~i_10_490_2983_0 & ~i_10_490_2985_0 & ~i_10_490_3093_0 & ~i_10_490_3545_0) | (~i_10_490_516_0 & ~i_10_490_997_0 & i_10_490_2350_0 & ~i_10_490_3613_0 & ~i_10_490_3895_0) | (~i_10_490_1312_0 & ~i_10_490_2728_0 & ~i_10_490_2831_0 & ~i_10_490_3984_0 & ~i_10_490_3986_0))) | (~i_10_490_34_0 & ~i_10_490_996_0 & i_10_490_1687_0 & ~i_10_490_1768_0 & ~i_10_490_1769_0 & ~i_10_490_2986_0));
endmodule



// Benchmark "kernel_10_491" written by ABC on Sun Jul 19 10:29:36 2020

module kernel_10_491 ( 
    i_10_491_30_0, i_10_491_123_0, i_10_491_171_0, i_10_491_243_0,
    i_10_491_281_0, i_10_491_283_0, i_10_491_286_0, i_10_491_287_0,
    i_10_491_432_0, i_10_491_464_0, i_10_491_465_0, i_10_491_711_0,
    i_10_491_747_0, i_10_491_892_0, i_10_491_955_0, i_10_491_956_0,
    i_10_491_1026_0, i_10_491_1233_0, i_10_491_1242_0, i_10_491_1263_0,
    i_10_491_1308_0, i_10_491_1310_0, i_10_491_1381_0, i_10_491_1396_0,
    i_10_491_1434_0, i_10_491_1450_0, i_10_491_1612_0, i_10_491_1652_0,
    i_10_491_1688_0, i_10_491_1766_0, i_10_491_1818_0, i_10_491_1989_0,
    i_10_491_1990_0, i_10_491_2181_0, i_10_491_2182_0, i_10_491_2185_0,
    i_10_491_2196_0, i_10_491_2358_0, i_10_491_2452_0, i_10_491_2453_0,
    i_10_491_2458_0, i_10_491_2566_0, i_10_491_2637_0, i_10_491_2683_0,
    i_10_491_2713_0, i_10_491_2714_0, i_10_491_2728_0, i_10_491_2729_0,
    i_10_491_2826_0, i_10_491_2827_0, i_10_491_2831_0, i_10_491_2869_0,
    i_10_491_2916_0, i_10_491_2917_0, i_10_491_2919_0, i_10_491_3040_0,
    i_10_491_3075_0, i_10_491_3076_0, i_10_491_3199_0, i_10_491_3200_0,
    i_10_491_3276_0, i_10_491_3283_0, i_10_491_3384_0, i_10_491_3385_0,
    i_10_491_3388_0, i_10_491_3408_0, i_10_491_3440_0, i_10_491_3466_0,
    i_10_491_3550_0, i_10_491_3551_0, i_10_491_3585_0, i_10_491_3586_0,
    i_10_491_3645_0, i_10_491_3646_0, i_10_491_3651_0, i_10_491_3726_0,
    i_10_491_3781_0, i_10_491_3782_0, i_10_491_3784_0, i_10_491_3785_0,
    i_10_491_3829_0, i_10_491_3843_0, i_10_491_3844_0, i_10_491_3847_0,
    i_10_491_3852_0, i_10_491_3854_0, i_10_491_3856_0, i_10_491_3857_0,
    i_10_491_3858_0, i_10_491_3860_0, i_10_491_3980_0, i_10_491_3987_0,
    i_10_491_3991_0, i_10_491_4024_0, i_10_491_4115_0, i_10_491_4149_0,
    i_10_491_4172_0, i_10_491_4288_0, i_10_491_4289_0, i_10_491_4291_0,
    o_10_491_0_0  );
  input  i_10_491_30_0, i_10_491_123_0, i_10_491_171_0, i_10_491_243_0,
    i_10_491_281_0, i_10_491_283_0, i_10_491_286_0, i_10_491_287_0,
    i_10_491_432_0, i_10_491_464_0, i_10_491_465_0, i_10_491_711_0,
    i_10_491_747_0, i_10_491_892_0, i_10_491_955_0, i_10_491_956_0,
    i_10_491_1026_0, i_10_491_1233_0, i_10_491_1242_0, i_10_491_1263_0,
    i_10_491_1308_0, i_10_491_1310_0, i_10_491_1381_0, i_10_491_1396_0,
    i_10_491_1434_0, i_10_491_1450_0, i_10_491_1612_0, i_10_491_1652_0,
    i_10_491_1688_0, i_10_491_1766_0, i_10_491_1818_0, i_10_491_1989_0,
    i_10_491_1990_0, i_10_491_2181_0, i_10_491_2182_0, i_10_491_2185_0,
    i_10_491_2196_0, i_10_491_2358_0, i_10_491_2452_0, i_10_491_2453_0,
    i_10_491_2458_0, i_10_491_2566_0, i_10_491_2637_0, i_10_491_2683_0,
    i_10_491_2713_0, i_10_491_2714_0, i_10_491_2728_0, i_10_491_2729_0,
    i_10_491_2826_0, i_10_491_2827_0, i_10_491_2831_0, i_10_491_2869_0,
    i_10_491_2916_0, i_10_491_2917_0, i_10_491_2919_0, i_10_491_3040_0,
    i_10_491_3075_0, i_10_491_3076_0, i_10_491_3199_0, i_10_491_3200_0,
    i_10_491_3276_0, i_10_491_3283_0, i_10_491_3384_0, i_10_491_3385_0,
    i_10_491_3388_0, i_10_491_3408_0, i_10_491_3440_0, i_10_491_3466_0,
    i_10_491_3550_0, i_10_491_3551_0, i_10_491_3585_0, i_10_491_3586_0,
    i_10_491_3645_0, i_10_491_3646_0, i_10_491_3651_0, i_10_491_3726_0,
    i_10_491_3781_0, i_10_491_3782_0, i_10_491_3784_0, i_10_491_3785_0,
    i_10_491_3829_0, i_10_491_3843_0, i_10_491_3844_0, i_10_491_3847_0,
    i_10_491_3852_0, i_10_491_3854_0, i_10_491_3856_0, i_10_491_3857_0,
    i_10_491_3858_0, i_10_491_3860_0, i_10_491_3980_0, i_10_491_3987_0,
    i_10_491_3991_0, i_10_491_4024_0, i_10_491_4115_0, i_10_491_4149_0,
    i_10_491_4172_0, i_10_491_4288_0, i_10_491_4289_0, i_10_491_4291_0;
  output o_10_491_0_0;
  assign o_10_491_0_0 = 0;
endmodule



// Benchmark "kernel_10_492" written by ABC on Sun Jul 19 10:29:37 2020

module kernel_10_492 ( 
    i_10_492_174_0, i_10_492_175_0, i_10_492_184_0, i_10_492_186_0,
    i_10_492_187_0, i_10_492_220_0, i_10_492_223_0, i_10_492_282_0,
    i_10_492_283_0, i_10_492_296_0, i_10_492_321_0, i_10_492_322_0,
    i_10_492_323_0, i_10_492_388_0, i_10_492_449_0, i_10_492_507_0,
    i_10_492_718_0, i_10_492_795_0, i_10_492_796_0, i_10_492_962_0,
    i_10_492_993_0, i_10_492_1041_0, i_10_492_1042_0, i_10_492_1141_0,
    i_10_492_1142_0, i_10_492_1308_0, i_10_492_1309_0, i_10_492_1546_0,
    i_10_492_1582_0, i_10_492_1683_0, i_10_492_1687_0, i_10_492_1688_0,
    i_10_492_1690_0, i_10_492_1821_0, i_10_492_1822_0, i_10_492_1824_0,
    i_10_492_1951_0, i_10_492_2179_0, i_10_492_2180_0, i_10_492_2352_0,
    i_10_492_2353_0, i_10_492_2354_0, i_10_492_2355_0, i_10_492_2364_0,
    i_10_492_2365_0, i_10_492_2407_0, i_10_492_2409_0, i_10_492_2451_0,
    i_10_492_2452_0, i_10_492_2453_0, i_10_492_2662_0, i_10_492_2681_0,
    i_10_492_2700_0, i_10_492_2702_0, i_10_492_2722_0, i_10_492_2725_0,
    i_10_492_2827_0, i_10_492_2883_0, i_10_492_2884_0, i_10_492_2887_0,
    i_10_492_2917_0, i_10_492_2919_0, i_10_492_2979_0, i_10_492_2986_0,
    i_10_492_3043_0, i_10_492_3201_0, i_10_492_3280_0, i_10_492_3283_0,
    i_10_492_3387_0, i_10_492_3405_0, i_10_492_3544_0, i_10_492_3549_0,
    i_10_492_3612_0, i_10_492_3613_0, i_10_492_3614_0, i_10_492_3647_0,
    i_10_492_3652_0, i_10_492_3780_0, i_10_492_3782_0, i_10_492_3783_0,
    i_10_492_3851_0, i_10_492_3855_0, i_10_492_3857_0, i_10_492_3859_0,
    i_10_492_3894_0, i_10_492_3915_0, i_10_492_3985_0, i_10_492_4114_0,
    i_10_492_4119_0, i_10_492_4123_0, i_10_492_4126_0, i_10_492_4127_0,
    i_10_492_4175_0, i_10_492_4282_0, i_10_492_4292_0, i_10_492_4564_0,
    i_10_492_4565_0, i_10_492_4566_0, i_10_492_4567_0, i_10_492_4568_0,
    o_10_492_0_0  );
  input  i_10_492_174_0, i_10_492_175_0, i_10_492_184_0, i_10_492_186_0,
    i_10_492_187_0, i_10_492_220_0, i_10_492_223_0, i_10_492_282_0,
    i_10_492_283_0, i_10_492_296_0, i_10_492_321_0, i_10_492_322_0,
    i_10_492_323_0, i_10_492_388_0, i_10_492_449_0, i_10_492_507_0,
    i_10_492_718_0, i_10_492_795_0, i_10_492_796_0, i_10_492_962_0,
    i_10_492_993_0, i_10_492_1041_0, i_10_492_1042_0, i_10_492_1141_0,
    i_10_492_1142_0, i_10_492_1308_0, i_10_492_1309_0, i_10_492_1546_0,
    i_10_492_1582_0, i_10_492_1683_0, i_10_492_1687_0, i_10_492_1688_0,
    i_10_492_1690_0, i_10_492_1821_0, i_10_492_1822_0, i_10_492_1824_0,
    i_10_492_1951_0, i_10_492_2179_0, i_10_492_2180_0, i_10_492_2352_0,
    i_10_492_2353_0, i_10_492_2354_0, i_10_492_2355_0, i_10_492_2364_0,
    i_10_492_2365_0, i_10_492_2407_0, i_10_492_2409_0, i_10_492_2451_0,
    i_10_492_2452_0, i_10_492_2453_0, i_10_492_2662_0, i_10_492_2681_0,
    i_10_492_2700_0, i_10_492_2702_0, i_10_492_2722_0, i_10_492_2725_0,
    i_10_492_2827_0, i_10_492_2883_0, i_10_492_2884_0, i_10_492_2887_0,
    i_10_492_2917_0, i_10_492_2919_0, i_10_492_2979_0, i_10_492_2986_0,
    i_10_492_3043_0, i_10_492_3201_0, i_10_492_3280_0, i_10_492_3283_0,
    i_10_492_3387_0, i_10_492_3405_0, i_10_492_3544_0, i_10_492_3549_0,
    i_10_492_3612_0, i_10_492_3613_0, i_10_492_3614_0, i_10_492_3647_0,
    i_10_492_3652_0, i_10_492_3780_0, i_10_492_3782_0, i_10_492_3783_0,
    i_10_492_3851_0, i_10_492_3855_0, i_10_492_3857_0, i_10_492_3859_0,
    i_10_492_3894_0, i_10_492_3915_0, i_10_492_3985_0, i_10_492_4114_0,
    i_10_492_4119_0, i_10_492_4123_0, i_10_492_4126_0, i_10_492_4127_0,
    i_10_492_4175_0, i_10_492_4282_0, i_10_492_4292_0, i_10_492_4564_0,
    i_10_492_4565_0, i_10_492_4566_0, i_10_492_4567_0, i_10_492_4568_0;
  output o_10_492_0_0;
  assign o_10_492_0_0 = ~((~i_10_492_3283_0 & ((~i_10_492_186_0 & ((~i_10_492_388_0 & ~i_10_492_1308_0 & ~i_10_492_2451_0 & ~i_10_492_2883_0 & ~i_10_492_3857_0 & ~i_10_492_4114_0 & ~i_10_492_4175_0) | (~i_10_492_187_0 & ~i_10_492_1041_0 & ~i_10_492_1821_0 & ~i_10_492_2180_0 & ~i_10_492_2986_0 & ~i_10_492_3280_0 & ~i_10_492_3544_0 & ~i_10_492_3783_0 & ~i_10_492_3855_0 & ~i_10_492_4282_0))) | (~i_10_492_1042_0 & ~i_10_492_2180_0 & ~i_10_492_2452_0 & ~i_10_492_3405_0 & ~i_10_492_3544_0 & ~i_10_492_3612_0 & ~i_10_492_4175_0) | (~i_10_492_1041_0 & i_10_492_1824_0 & ~i_10_492_2179_0 & ~i_10_492_2453_0 & ~i_10_492_2887_0 & ~i_10_492_3855_0 & ~i_10_492_3985_0))) | (~i_10_492_220_0 & ((~i_10_492_282_0 & ((~i_10_492_1546_0 & ~i_10_492_2451_0 & ~i_10_492_2452_0 & i_10_492_3859_0) | (~i_10_492_1308_0 & ~i_10_492_1821_0 & ~i_10_492_2354_0 & ~i_10_492_2827_0 & ~i_10_492_2917_0 & ~i_10_492_3782_0 & ~i_10_492_3859_0 & ~i_10_492_4175_0 & ~i_10_492_4292_0))) | (~i_10_492_1546_0 & ~i_10_492_3405_0 & ((i_10_492_283_0 & ~i_10_492_322_0 & ~i_10_492_1041_0 & ~i_10_492_1042_0 & ~i_10_492_1687_0 & ~i_10_492_2179_0) | (~i_10_492_388_0 & ~i_10_492_3549_0 & ~i_10_492_3780_0 & ~i_10_492_3782_0 & ~i_10_492_3894_0 & i_10_492_4114_0))) | (i_10_492_3652_0 & ~i_10_492_3780_0 & i_10_492_3782_0 & ~i_10_492_4282_0 & ~i_10_492_4292_0))) | (~i_10_492_4282_0 & ((~i_10_492_283_0 & ((~i_10_492_174_0 & ~i_10_492_2451_0 & ~i_10_492_2452_0 & ~i_10_492_3544_0 & ~i_10_492_3783_0) | (i_10_492_175_0 & ~i_10_492_2883_0 & ~i_10_492_2919_0 & ~i_10_492_3405_0 & ~i_10_492_4175_0))) | (~i_10_492_1309_0 & ~i_10_492_2884_0 & ~i_10_492_3280_0 & ~i_10_492_3780_0 & ~i_10_492_3855_0))) | (~i_10_492_322_0 & ((~i_10_492_187_0 & i_10_492_1309_0 & ~i_10_492_1546_0 & ~i_10_492_1688_0 & i_10_492_2662_0 & ~i_10_492_3405_0 & ~i_10_492_3549_0 & ~i_10_492_4123_0 & ~i_10_492_4564_0) | (~i_10_492_1309_0 & ~i_10_492_2453_0 & i_10_492_2917_0 & ~i_10_492_3387_0 & ~i_10_492_3783_0 & ~i_10_492_4567_0))) | (~i_10_492_1683_0 & ((~i_10_492_187_0 & ~i_10_492_1309_0 & ~i_10_492_2887_0 & i_10_492_3387_0) | (~i_10_492_795_0 & ~i_10_492_1042_0 & i_10_492_1309_0 & ~i_10_492_1688_0 & ~i_10_492_1951_0 & i_10_492_2354_0 & ~i_10_492_2451_0 & ~i_10_492_3387_0))) | (~i_10_492_187_0 & ((i_10_492_449_0 & ~i_10_492_3783_0 & i_10_492_3859_0 & ~i_10_492_4292_0) | (~i_10_492_795_0 & ~i_10_492_1582_0 & ~i_10_492_2681_0 & i_10_492_3387_0 & ~i_10_492_3544_0 & ~i_10_492_3652_0 & ~i_10_492_4568_0))) | (~i_10_492_1821_0 & ((~i_10_492_2451_0 & ~i_10_492_3613_0 & i_10_492_3783_0) | (i_10_492_2702_0 & i_10_492_3857_0))) | (~i_10_492_2179_0 & ~i_10_492_3985_0 & ((~i_10_492_323_0 & ~i_10_492_795_0 & ~i_10_492_1688_0 & ~i_10_492_2352_0 & ~i_10_492_3612_0 & ~i_10_492_3780_0 & ~i_10_492_3782_0) | (i_10_492_2725_0 & ~i_10_492_3544_0 & ~i_10_492_3783_0 & ~i_10_492_4114_0 & ~i_10_492_4175_0))) | (~i_10_492_2452_0 & ((~i_10_492_1309_0 & i_10_492_2883_0 & ~i_10_492_3280_0) | (~i_10_492_2451_0 & ~i_10_492_3612_0 & i_10_492_3647_0 & ~i_10_492_3783_0 & ~i_10_492_4126_0))) | (~i_10_492_1309_0 & ((~i_10_492_1041_0 & ~i_10_492_1042_0 & ~i_10_492_1546_0 & i_10_492_1824_0 & ~i_10_492_2883_0) | (~i_10_492_321_0 & ~i_10_492_3201_0 & ~i_10_492_3544_0 & ~i_10_492_3612_0 & ~i_10_492_3613_0 & ~i_10_492_3855_0))) | (~i_10_492_1042_0 & ((i_10_492_2725_0 & i_10_492_2917_0) | (i_10_492_2352_0 & ~i_10_492_3280_0 & ~i_10_492_3544_0 & ~i_10_492_3614_0 & ~i_10_492_3851_0 & ~i_10_492_4126_0 & ~i_10_492_4566_0))));
endmodule



// Benchmark "kernel_10_493" written by ABC on Sun Jul 19 10:29:38 2020

module kernel_10_493 ( 
    i_10_493_120_0, i_10_493_245_0, i_10_493_257_0, i_10_493_317_0,
    i_10_493_320_0, i_10_493_329_0, i_10_493_390_0, i_10_493_393_0,
    i_10_493_435_0, i_10_493_436_0, i_10_493_437_0, i_10_493_438_0,
    i_10_493_589_0, i_10_493_641_0, i_10_493_688_0, i_10_493_712_0,
    i_10_493_869_0, i_10_493_921_0, i_10_493_992_0, i_10_493_993_0,
    i_10_493_1002_0, i_10_493_1006_0, i_10_493_1135_0, i_10_493_1215_0,
    i_10_493_1216_0, i_10_493_1217_0, i_10_493_1218_0, i_10_493_1219_0,
    i_10_493_1238_0, i_10_493_1267_0, i_10_493_1305_0, i_10_493_1309_0,
    i_10_493_1311_0, i_10_493_1615_0, i_10_493_1618_0, i_10_493_1653_0,
    i_10_493_1804_0, i_10_493_1819_0, i_10_493_1921_0, i_10_493_1947_0,
    i_10_493_1948_0, i_10_493_1950_0, i_10_493_2021_0, i_10_493_2155_0,
    i_10_493_2202_0, i_10_493_2203_0, i_10_493_2355_0, i_10_493_2377_0,
    i_10_493_2513_0, i_10_493_2514_0, i_10_493_2515_0, i_10_493_2540_0,
    i_10_493_2543_0, i_10_493_2582_0, i_10_493_2613_0, i_10_493_2655_0,
    i_10_493_2662_0, i_10_493_2677_0, i_10_493_2744_0, i_10_493_2811_0,
    i_10_493_2812_0, i_10_493_2824_0, i_10_493_2831_0, i_10_493_2834_0,
    i_10_493_2848_0, i_10_493_2880_0, i_10_493_2881_0, i_10_493_2882_0,
    i_10_493_3059_0, i_10_493_3090_0, i_10_493_3332_0, i_10_493_3353_0,
    i_10_493_3397_0, i_10_493_3404_0, i_10_493_3443_0, i_10_493_3445_0,
    i_10_493_3473_0, i_10_493_3525_0, i_10_493_3539_0, i_10_493_3651_0,
    i_10_493_3687_0, i_10_493_3717_0, i_10_493_3718_0, i_10_493_3721_0,
    i_10_493_3815_0, i_10_493_3837_0, i_10_493_3853_0, i_10_493_3893_0,
    i_10_493_3910_0, i_10_493_3912_0, i_10_493_3928_0, i_10_493_3993_0,
    i_10_493_4054_0, i_10_493_4168_0, i_10_493_4185_0, i_10_493_4233_0,
    i_10_493_4276_0, i_10_493_4280_0, i_10_493_4283_0, i_10_493_4519_0,
    o_10_493_0_0  );
  input  i_10_493_120_0, i_10_493_245_0, i_10_493_257_0, i_10_493_317_0,
    i_10_493_320_0, i_10_493_329_0, i_10_493_390_0, i_10_493_393_0,
    i_10_493_435_0, i_10_493_436_0, i_10_493_437_0, i_10_493_438_0,
    i_10_493_589_0, i_10_493_641_0, i_10_493_688_0, i_10_493_712_0,
    i_10_493_869_0, i_10_493_921_0, i_10_493_992_0, i_10_493_993_0,
    i_10_493_1002_0, i_10_493_1006_0, i_10_493_1135_0, i_10_493_1215_0,
    i_10_493_1216_0, i_10_493_1217_0, i_10_493_1218_0, i_10_493_1219_0,
    i_10_493_1238_0, i_10_493_1267_0, i_10_493_1305_0, i_10_493_1309_0,
    i_10_493_1311_0, i_10_493_1615_0, i_10_493_1618_0, i_10_493_1653_0,
    i_10_493_1804_0, i_10_493_1819_0, i_10_493_1921_0, i_10_493_1947_0,
    i_10_493_1948_0, i_10_493_1950_0, i_10_493_2021_0, i_10_493_2155_0,
    i_10_493_2202_0, i_10_493_2203_0, i_10_493_2355_0, i_10_493_2377_0,
    i_10_493_2513_0, i_10_493_2514_0, i_10_493_2515_0, i_10_493_2540_0,
    i_10_493_2543_0, i_10_493_2582_0, i_10_493_2613_0, i_10_493_2655_0,
    i_10_493_2662_0, i_10_493_2677_0, i_10_493_2744_0, i_10_493_2811_0,
    i_10_493_2812_0, i_10_493_2824_0, i_10_493_2831_0, i_10_493_2834_0,
    i_10_493_2848_0, i_10_493_2880_0, i_10_493_2881_0, i_10_493_2882_0,
    i_10_493_3059_0, i_10_493_3090_0, i_10_493_3332_0, i_10_493_3353_0,
    i_10_493_3397_0, i_10_493_3404_0, i_10_493_3443_0, i_10_493_3445_0,
    i_10_493_3473_0, i_10_493_3525_0, i_10_493_3539_0, i_10_493_3651_0,
    i_10_493_3687_0, i_10_493_3717_0, i_10_493_3718_0, i_10_493_3721_0,
    i_10_493_3815_0, i_10_493_3837_0, i_10_493_3853_0, i_10_493_3893_0,
    i_10_493_3910_0, i_10_493_3912_0, i_10_493_3928_0, i_10_493_3993_0,
    i_10_493_4054_0, i_10_493_4168_0, i_10_493_4185_0, i_10_493_4233_0,
    i_10_493_4276_0, i_10_493_4280_0, i_10_493_4283_0, i_10_493_4519_0;
  output o_10_493_0_0;
  assign o_10_493_0_0 = 0;
endmodule



// Benchmark "kernel_10_494" written by ABC on Sun Jul 19 10:29:39 2020

module kernel_10_494 ( 
    i_10_494_171_0, i_10_494_174_0, i_10_494_181_0, i_10_494_283_0,
    i_10_494_285_0, i_10_494_287_0, i_10_494_328_0, i_10_494_388_0,
    i_10_494_424_0, i_10_494_425_0, i_10_494_434_0, i_10_494_438_0,
    i_10_494_451_0, i_10_494_459_0, i_10_494_749_0, i_10_494_753_0,
    i_10_494_754_0, i_10_494_755_0, i_10_494_797_0, i_10_494_968_0,
    i_10_494_1037_0, i_10_494_1234_0, i_10_494_1235_0, i_10_494_1240_0,
    i_10_494_1242_0, i_10_494_1306_0, i_10_494_1309_0, i_10_494_1359_0,
    i_10_494_1650_0, i_10_494_1687_0, i_10_494_1688_0, i_10_494_1819_0,
    i_10_494_1821_0, i_10_494_1822_0, i_10_494_1823_0, i_10_494_1996_0,
    i_10_494_2362_0, i_10_494_2383_0, i_10_494_2448_0, i_10_494_2451_0,
    i_10_494_2628_0, i_10_494_2629_0, i_10_494_2630_0, i_10_494_2634_0,
    i_10_494_2655_0, i_10_494_2656_0, i_10_494_2657_0, i_10_494_2659_0,
    i_10_494_2713_0, i_10_494_2715_0, i_10_494_2716_0, i_10_494_2717_0,
    i_10_494_2919_0, i_10_494_2921_0, i_10_494_2923_0, i_10_494_3036_0,
    i_10_494_3046_0, i_10_494_3050_0, i_10_494_3085_0, i_10_494_3094_0,
    i_10_494_3155_0, i_10_494_3271_0, i_10_494_3280_0, i_10_494_3284_0,
    i_10_494_3402_0, i_10_494_3405_0, i_10_494_3408_0, i_10_494_3586_0,
    i_10_494_3609_0, i_10_494_3613_0, i_10_494_3614_0, i_10_494_3615_0,
    i_10_494_3616_0, i_10_494_3785_0, i_10_494_3834_0, i_10_494_3840_0,
    i_10_494_3841_0, i_10_494_3846_0, i_10_494_3847_0, i_10_494_3848_0,
    i_10_494_3852_0, i_10_494_3856_0, i_10_494_3857_0, i_10_494_3858_0,
    i_10_494_3859_0, i_10_494_3860_0, i_10_494_3990_0, i_10_494_3991_0,
    i_10_494_4116_0, i_10_494_4117_0, i_10_494_4119_0, i_10_494_4120_0,
    i_10_494_4123_0, i_10_494_4269_0, i_10_494_4270_0, i_10_494_4287_0,
    i_10_494_4288_0, i_10_494_4563_0, i_10_494_4567_0, i_10_494_4568_0,
    o_10_494_0_0  );
  input  i_10_494_171_0, i_10_494_174_0, i_10_494_181_0, i_10_494_283_0,
    i_10_494_285_0, i_10_494_287_0, i_10_494_328_0, i_10_494_388_0,
    i_10_494_424_0, i_10_494_425_0, i_10_494_434_0, i_10_494_438_0,
    i_10_494_451_0, i_10_494_459_0, i_10_494_749_0, i_10_494_753_0,
    i_10_494_754_0, i_10_494_755_0, i_10_494_797_0, i_10_494_968_0,
    i_10_494_1037_0, i_10_494_1234_0, i_10_494_1235_0, i_10_494_1240_0,
    i_10_494_1242_0, i_10_494_1306_0, i_10_494_1309_0, i_10_494_1359_0,
    i_10_494_1650_0, i_10_494_1687_0, i_10_494_1688_0, i_10_494_1819_0,
    i_10_494_1821_0, i_10_494_1822_0, i_10_494_1823_0, i_10_494_1996_0,
    i_10_494_2362_0, i_10_494_2383_0, i_10_494_2448_0, i_10_494_2451_0,
    i_10_494_2628_0, i_10_494_2629_0, i_10_494_2630_0, i_10_494_2634_0,
    i_10_494_2655_0, i_10_494_2656_0, i_10_494_2657_0, i_10_494_2659_0,
    i_10_494_2713_0, i_10_494_2715_0, i_10_494_2716_0, i_10_494_2717_0,
    i_10_494_2919_0, i_10_494_2921_0, i_10_494_2923_0, i_10_494_3036_0,
    i_10_494_3046_0, i_10_494_3050_0, i_10_494_3085_0, i_10_494_3094_0,
    i_10_494_3155_0, i_10_494_3271_0, i_10_494_3280_0, i_10_494_3284_0,
    i_10_494_3402_0, i_10_494_3405_0, i_10_494_3408_0, i_10_494_3586_0,
    i_10_494_3609_0, i_10_494_3613_0, i_10_494_3614_0, i_10_494_3615_0,
    i_10_494_3616_0, i_10_494_3785_0, i_10_494_3834_0, i_10_494_3840_0,
    i_10_494_3841_0, i_10_494_3846_0, i_10_494_3847_0, i_10_494_3848_0,
    i_10_494_3852_0, i_10_494_3856_0, i_10_494_3857_0, i_10_494_3858_0,
    i_10_494_3859_0, i_10_494_3860_0, i_10_494_3990_0, i_10_494_3991_0,
    i_10_494_4116_0, i_10_494_4117_0, i_10_494_4119_0, i_10_494_4120_0,
    i_10_494_4123_0, i_10_494_4269_0, i_10_494_4270_0, i_10_494_4287_0,
    i_10_494_4288_0, i_10_494_4563_0, i_10_494_4567_0, i_10_494_4568_0;
  output o_10_494_0_0;
  assign o_10_494_0_0 = ~((~i_10_494_174_0 & ((~i_10_494_2921_0 & ~i_10_494_3405_0 & i_10_494_3841_0 & ~i_10_494_4120_0) | (~i_10_494_181_0 & ~i_10_494_754_0 & ~i_10_494_968_0 & ~i_10_494_1235_0 & ~i_10_494_3036_0 & ~i_10_494_3785_0 & ~i_10_494_3841_0 & ~i_10_494_3856_0 & ~i_10_494_4119_0 & ~i_10_494_4287_0))) | (i_10_494_1240_0 & ((~i_10_494_754_0 & ~i_10_494_968_0 & i_10_494_2713_0 & ~i_10_494_3991_0) | (~i_10_494_434_0 & ~i_10_494_753_0 & ~i_10_494_755_0 & ~i_10_494_1996_0 & i_10_494_3046_0 & ~i_10_494_3785_0 & ~i_10_494_4269_0))) | (~i_10_494_283_0 & ((~i_10_494_1240_0 & ((~i_10_494_388_0 & i_10_494_1819_0 & ~i_10_494_1823_0 & ~i_10_494_3036_0 & ~i_10_494_3990_0) | (~i_10_494_451_0 & ~i_10_494_1037_0 & ~i_10_494_1234_0 & ~i_10_494_1650_0 & ~i_10_494_1687_0 & ~i_10_494_3785_0 & ~i_10_494_4120_0))) | (i_10_494_3841_0 & ~i_10_494_3848_0 & ~i_10_494_3991_0 & ~i_10_494_4287_0 & ~i_10_494_4567_0))) | (~i_10_494_2383_0 & ((~i_10_494_3846_0 & ((~i_10_494_451_0 & ~i_10_494_1688_0 & ((~i_10_494_755_0 & ~i_10_494_1037_0 & i_10_494_1819_0 & ~i_10_494_2362_0 & ~i_10_494_2451_0 & ~i_10_494_3284_0 & ~i_10_494_3615_0 & ~i_10_494_3785_0) | (~i_10_494_968_0 & ~i_10_494_1359_0 & ~i_10_494_2630_0 & ~i_10_494_3614_0 & ~i_10_494_3857_0 & ~i_10_494_4117_0))) | (~i_10_494_753_0 & ~i_10_494_1687_0 & ~i_10_494_1821_0 & ~i_10_494_2921_0 & ~i_10_494_3857_0 & ~i_10_494_4568_0))) | (i_10_494_2628_0 & ~i_10_494_2717_0 & i_10_494_3616_0) | (~i_10_494_753_0 & ~i_10_494_1823_0 & i_10_494_2448_0 & ~i_10_494_2923_0 & ~i_10_494_4567_0))) | (~i_10_494_451_0 & ((~i_10_494_388_0 & ~i_10_494_755_0 & ~i_10_494_968_0 & ~i_10_494_1821_0 & ~i_10_494_1822_0 & ~i_10_494_2716_0 & ~i_10_494_2717_0 & ~i_10_494_4119_0) | (~i_10_494_1037_0 & i_10_494_2628_0 & ~i_10_494_3036_0 & ~i_10_494_3990_0 & ~i_10_494_4269_0 & ~i_10_494_4567_0))) | (~i_10_494_388_0 & ((i_10_494_434_0 & ~i_10_494_754_0) | (~i_10_494_1037_0 & i_10_494_1687_0 & i_10_494_1688_0 & ~i_10_494_3036_0 & ~i_10_494_4123_0 & ~i_10_494_4270_0))) | (~i_10_494_2919_0 & ((~i_10_494_968_0 & ((~i_10_494_754_0 & i_10_494_1823_0 & ~i_10_494_2451_0 & ~i_10_494_3834_0 & ~i_10_494_3847_0 & ~i_10_494_4116_0) | (i_10_494_3615_0 & i_10_494_3858_0 & ~i_10_494_4269_0))) | (~i_10_494_753_0 & ~i_10_494_755_0 & ~i_10_494_1823_0 & ~i_10_494_3847_0 & ~i_10_494_3848_0) | (~i_10_494_4120_0 & i_10_494_4269_0 & i_10_494_4563_0))) | (~i_10_494_3848_0 & ((~i_10_494_754_0 & ((i_10_494_3405_0 & ~i_10_494_4269_0) | (~i_10_494_3847_0 & ~i_10_494_3857_0 & ~i_10_494_4119_0 & ~i_10_494_4123_0 & ~i_10_494_4270_0))) | i_10_494_3860_0 | (~i_10_494_1821_0 & ~i_10_494_4120_0 & ~i_10_494_4123_0))) | (~i_10_494_755_0 & ((i_10_494_797_0 & ~i_10_494_1037_0 & i_10_494_1822_0 & ~i_10_494_2716_0 & ~i_10_494_3857_0 & ~i_10_494_3991_0 & ~i_10_494_4116_0 & ~i_10_494_4270_0) | (~i_10_494_1235_0 & ~i_10_494_1821_0 & ~i_10_494_3036_0 & ~i_10_494_3840_0 & ~i_10_494_4287_0 & ~i_10_494_4567_0 & ~i_10_494_4568_0))) | (~i_10_494_1037_0 & ~i_10_494_3852_0 & ((i_10_494_451_0 & ~i_10_494_2451_0 & ~i_10_494_3847_0 & ~i_10_494_4117_0) | (i_10_494_1819_0 & i_10_494_1822_0 & i_10_494_1823_0 & ~i_10_494_3586_0 & ~i_10_494_3856_0 & ~i_10_494_3990_0 & ~i_10_494_4123_0))) | (~i_10_494_4117_0 & ((i_10_494_424_0 & ~i_10_494_3405_0) | (~i_10_494_3036_0 & i_10_494_3785_0 & i_10_494_3857_0 & ~i_10_494_4568_0))) | (i_10_494_2630_0 & i_10_494_2659_0 & ~i_10_494_3402_0) | (~i_10_494_1650_0 & ~i_10_494_2634_0 & ~i_10_494_3609_0 & i_10_494_3613_0 & i_10_494_3856_0 & ~i_10_494_3991_0 & ~i_10_494_4123_0 & ~i_10_494_4568_0) | (~i_10_494_3785_0 & ~i_10_494_3847_0 & ~i_10_494_4120_0 & ~i_10_494_4270_0 & i_10_494_4567_0));
endmodule



// Benchmark "kernel_10_495" written by ABC on Sun Jul 19 10:29:40 2020

module kernel_10_495 ( 
    i_10_495_32_0, i_10_495_129_0, i_10_495_158_0, i_10_495_161_0,
    i_10_495_264_0, i_10_495_274_0, i_10_495_441_0, i_10_495_446_0,
    i_10_495_518_0, i_10_495_561_0, i_10_495_674_0, i_10_495_718_0,
    i_10_495_755_0, i_10_495_834_0, i_10_495_835_0, i_10_495_922_0,
    i_10_495_986_0, i_10_495_989_0, i_10_495_997_0, i_10_495_998_0,
    i_10_495_1002_0, i_10_495_1005_0, i_10_495_1061_0, i_10_495_1103_0,
    i_10_495_1234_0, i_10_495_1235_0, i_10_495_1248_0, i_10_495_1249_0,
    i_10_495_1340_0, i_10_495_1345_0, i_10_495_1452_0, i_10_495_1488_0,
    i_10_495_1493_0, i_10_495_1538_0, i_10_495_1555_0, i_10_495_1582_0,
    i_10_495_1637_0, i_10_495_1641_0, i_10_495_1646_0, i_10_495_1799_0,
    i_10_495_1818_0, i_10_495_1820_0, i_10_495_1821_0, i_10_495_1822_0,
    i_10_495_1824_0, i_10_495_1940_0, i_10_495_1942_0, i_10_495_1945_0,
    i_10_495_2003_0, i_10_495_2033_0, i_10_495_2069_0, i_10_495_2258_0,
    i_10_495_2408_0, i_10_495_2452_0, i_10_495_2472_0, i_10_495_2605_0,
    i_10_495_2636_0, i_10_495_2681_0, i_10_495_2712_0, i_10_495_2714_0,
    i_10_495_2717_0, i_10_495_2723_0, i_10_495_2734_0, i_10_495_2735_0,
    i_10_495_2804_0, i_10_495_2870_0, i_10_495_2956_0, i_10_495_2986_0,
    i_10_495_2987_0, i_10_495_3011_0, i_10_495_3039_0, i_10_495_3047_0,
    i_10_495_3074_0, i_10_495_3158_0, i_10_495_3238_0, i_10_495_3239_0,
    i_10_495_3282_0, i_10_495_3360_0, i_10_495_3387_0, i_10_495_3406_0,
    i_10_495_3468_0, i_10_495_3470_0, i_10_495_3496_0, i_10_495_3506_0,
    i_10_495_3509_0, i_10_495_3561_0, i_10_495_3617_0, i_10_495_3624_0,
    i_10_495_3806_0, i_10_495_3815_0, i_10_495_3846_0, i_10_495_3884_0,
    i_10_495_3913_0, i_10_495_3946_0, i_10_495_3947_0, i_10_495_3950_0,
    i_10_495_4271_0, i_10_495_4278_0, i_10_495_4290_0, i_10_495_4292_0,
    o_10_495_0_0  );
  input  i_10_495_32_0, i_10_495_129_0, i_10_495_158_0, i_10_495_161_0,
    i_10_495_264_0, i_10_495_274_0, i_10_495_441_0, i_10_495_446_0,
    i_10_495_518_0, i_10_495_561_0, i_10_495_674_0, i_10_495_718_0,
    i_10_495_755_0, i_10_495_834_0, i_10_495_835_0, i_10_495_922_0,
    i_10_495_986_0, i_10_495_989_0, i_10_495_997_0, i_10_495_998_0,
    i_10_495_1002_0, i_10_495_1005_0, i_10_495_1061_0, i_10_495_1103_0,
    i_10_495_1234_0, i_10_495_1235_0, i_10_495_1248_0, i_10_495_1249_0,
    i_10_495_1340_0, i_10_495_1345_0, i_10_495_1452_0, i_10_495_1488_0,
    i_10_495_1493_0, i_10_495_1538_0, i_10_495_1555_0, i_10_495_1582_0,
    i_10_495_1637_0, i_10_495_1641_0, i_10_495_1646_0, i_10_495_1799_0,
    i_10_495_1818_0, i_10_495_1820_0, i_10_495_1821_0, i_10_495_1822_0,
    i_10_495_1824_0, i_10_495_1940_0, i_10_495_1942_0, i_10_495_1945_0,
    i_10_495_2003_0, i_10_495_2033_0, i_10_495_2069_0, i_10_495_2258_0,
    i_10_495_2408_0, i_10_495_2452_0, i_10_495_2472_0, i_10_495_2605_0,
    i_10_495_2636_0, i_10_495_2681_0, i_10_495_2712_0, i_10_495_2714_0,
    i_10_495_2717_0, i_10_495_2723_0, i_10_495_2734_0, i_10_495_2735_0,
    i_10_495_2804_0, i_10_495_2870_0, i_10_495_2956_0, i_10_495_2986_0,
    i_10_495_2987_0, i_10_495_3011_0, i_10_495_3039_0, i_10_495_3047_0,
    i_10_495_3074_0, i_10_495_3158_0, i_10_495_3238_0, i_10_495_3239_0,
    i_10_495_3282_0, i_10_495_3360_0, i_10_495_3387_0, i_10_495_3406_0,
    i_10_495_3468_0, i_10_495_3470_0, i_10_495_3496_0, i_10_495_3506_0,
    i_10_495_3509_0, i_10_495_3561_0, i_10_495_3617_0, i_10_495_3624_0,
    i_10_495_3806_0, i_10_495_3815_0, i_10_495_3846_0, i_10_495_3884_0,
    i_10_495_3913_0, i_10_495_3946_0, i_10_495_3947_0, i_10_495_3950_0,
    i_10_495_4271_0, i_10_495_4278_0, i_10_495_4290_0, i_10_495_4292_0;
  output o_10_495_0_0;
  assign o_10_495_0_0 = 0;
endmodule



// Benchmark "kernel_10_496" written by ABC on Sun Jul 19 10:29:41 2020

module kernel_10_496 ( 
    i_10_496_71_0, i_10_496_119_0, i_10_496_254_0, i_10_496_257_0,
    i_10_496_265_0, i_10_496_266_0, i_10_496_279_0, i_10_496_392_0,
    i_10_496_395_0, i_10_496_448_0, i_10_496_466_0, i_10_496_517_0,
    i_10_496_535_0, i_10_496_560_0, i_10_496_895_0, i_10_496_1000_0,
    i_10_496_1003_0, i_10_496_1004_0, i_10_496_1028_0, i_10_496_1109_0,
    i_10_496_1112_0, i_10_496_1236_0, i_10_496_1239_0, i_10_496_1273_0,
    i_10_496_1298_0, i_10_496_1300_0, i_10_496_1309_0, i_10_496_1311_0,
    i_10_496_1312_0, i_10_496_1360_0, i_10_496_1364_0, i_10_496_1400_0,
    i_10_496_1436_0, i_10_496_1625_0, i_10_496_1648_0, i_10_496_1652_0,
    i_10_496_1712_0, i_10_496_1799_0, i_10_496_1804_0, i_10_496_1805_0,
    i_10_496_1808_0, i_10_496_1909_0, i_10_496_1914_0, i_10_496_1919_0,
    i_10_496_1985_0, i_10_496_2080_0, i_10_496_2178_0, i_10_496_2186_0,
    i_10_496_2188_0, i_10_496_2350_0, i_10_496_2356_0, i_10_496_2379_0,
    i_10_496_2382_0, i_10_496_2430_0, i_10_496_2450_0, i_10_496_2506_0,
    i_10_496_2547_0, i_10_496_2557_0, i_10_496_2558_0, i_10_496_2560_0,
    i_10_496_2561_0, i_10_496_2566_0, i_10_496_2567_0, i_10_496_2569_0,
    i_10_496_2597_0, i_10_496_2641_0, i_10_496_2701_0, i_10_496_2705_0,
    i_10_496_2708_0, i_10_496_2848_0, i_10_496_2849_0, i_10_496_3033_0,
    i_10_496_3034_0, i_10_496_3200_0, i_10_496_3232_0, i_10_496_3235_0,
    i_10_496_3270_0, i_10_496_3274_0, i_10_496_3278_0, i_10_496_3283_0,
    i_10_496_3289_0, i_10_496_3292_0, i_10_496_3429_0, i_10_496_3430_0,
    i_10_496_3466_0, i_10_496_3470_0, i_10_496_3540_0, i_10_496_3542_0,
    i_10_496_3568_0, i_10_496_3652_0, i_10_496_3794_0, i_10_496_3797_0,
    i_10_496_3838_0, i_10_496_3841_0, i_10_496_4148_0, i_10_496_4171_0,
    i_10_496_4277_0, i_10_496_4282_0, i_10_496_4567_0, i_10_496_4589_0,
    o_10_496_0_0  );
  input  i_10_496_71_0, i_10_496_119_0, i_10_496_254_0, i_10_496_257_0,
    i_10_496_265_0, i_10_496_266_0, i_10_496_279_0, i_10_496_392_0,
    i_10_496_395_0, i_10_496_448_0, i_10_496_466_0, i_10_496_517_0,
    i_10_496_535_0, i_10_496_560_0, i_10_496_895_0, i_10_496_1000_0,
    i_10_496_1003_0, i_10_496_1004_0, i_10_496_1028_0, i_10_496_1109_0,
    i_10_496_1112_0, i_10_496_1236_0, i_10_496_1239_0, i_10_496_1273_0,
    i_10_496_1298_0, i_10_496_1300_0, i_10_496_1309_0, i_10_496_1311_0,
    i_10_496_1312_0, i_10_496_1360_0, i_10_496_1364_0, i_10_496_1400_0,
    i_10_496_1436_0, i_10_496_1625_0, i_10_496_1648_0, i_10_496_1652_0,
    i_10_496_1712_0, i_10_496_1799_0, i_10_496_1804_0, i_10_496_1805_0,
    i_10_496_1808_0, i_10_496_1909_0, i_10_496_1914_0, i_10_496_1919_0,
    i_10_496_1985_0, i_10_496_2080_0, i_10_496_2178_0, i_10_496_2186_0,
    i_10_496_2188_0, i_10_496_2350_0, i_10_496_2356_0, i_10_496_2379_0,
    i_10_496_2382_0, i_10_496_2430_0, i_10_496_2450_0, i_10_496_2506_0,
    i_10_496_2547_0, i_10_496_2557_0, i_10_496_2558_0, i_10_496_2560_0,
    i_10_496_2561_0, i_10_496_2566_0, i_10_496_2567_0, i_10_496_2569_0,
    i_10_496_2597_0, i_10_496_2641_0, i_10_496_2701_0, i_10_496_2705_0,
    i_10_496_2708_0, i_10_496_2848_0, i_10_496_2849_0, i_10_496_3033_0,
    i_10_496_3034_0, i_10_496_3200_0, i_10_496_3232_0, i_10_496_3235_0,
    i_10_496_3270_0, i_10_496_3274_0, i_10_496_3278_0, i_10_496_3283_0,
    i_10_496_3289_0, i_10_496_3292_0, i_10_496_3429_0, i_10_496_3430_0,
    i_10_496_3466_0, i_10_496_3470_0, i_10_496_3540_0, i_10_496_3542_0,
    i_10_496_3568_0, i_10_496_3652_0, i_10_496_3794_0, i_10_496_3797_0,
    i_10_496_3838_0, i_10_496_3841_0, i_10_496_4148_0, i_10_496_4171_0,
    i_10_496_4277_0, i_10_496_4282_0, i_10_496_4567_0, i_10_496_4589_0;
  output o_10_496_0_0;
  assign o_10_496_0_0 = 0;
endmodule



// Benchmark "kernel_10_497" written by ABC on Sun Jul 19 10:29:43 2020

module kernel_10_497 ( 
    i_10_497_123_0, i_10_497_216_0, i_10_497_261_0, i_10_497_279_0,
    i_10_497_280_0, i_10_497_281_0, i_10_497_282_0, i_10_497_320_0,
    i_10_497_405_0, i_10_497_443_0, i_10_497_444_0, i_10_497_460_0,
    i_10_497_462_0, i_10_497_904_0, i_10_497_956_0, i_10_497_1053_0,
    i_10_497_1239_0, i_10_497_1263_0, i_10_497_1311_0, i_10_497_1431_0,
    i_10_497_1432_0, i_10_497_1449_0, i_10_497_1539_0, i_10_497_1540_0,
    i_10_497_1542_0, i_10_497_1581_0, i_10_497_1620_0, i_10_497_1629_0,
    i_10_497_1630_0, i_10_497_1651_0, i_10_497_1652_0, i_10_497_1685_0,
    i_10_497_1800_0, i_10_497_1823_0, i_10_497_1944_0, i_10_497_2025_0,
    i_10_497_2026_0, i_10_497_2199_0, i_10_497_2331_0, i_10_497_2351_0,
    i_10_497_2355_0, i_10_497_2403_0, i_10_497_2404_0, i_10_497_2448_0,
    i_10_497_2449_0, i_10_497_2452_0, i_10_497_2470_0, i_10_497_2545_0,
    i_10_497_2565_0, i_10_497_2604_0, i_10_497_2647_0, i_10_497_2662_0,
    i_10_497_2709_0, i_10_497_2718_0, i_10_497_2720_0, i_10_497_2727_0,
    i_10_497_2821_0, i_10_497_2826_0, i_10_497_2844_0, i_10_497_2865_0,
    i_10_497_2961_0, i_10_497_3042_0, i_10_497_3089_0, i_10_497_3278_0,
    i_10_497_3333_0, i_10_497_3386_0, i_10_497_3387_0, i_10_497_3388_0,
    i_10_497_3390_0, i_10_497_3408_0, i_10_497_3468_0, i_10_497_3471_0,
    i_10_497_3537_0, i_10_497_3555_0, i_10_497_3582_0, i_10_497_3610_0,
    i_10_497_3613_0, i_10_497_3618_0, i_10_497_3621_0, i_10_497_3645_0,
    i_10_497_3648_0, i_10_497_3785_0, i_10_497_3840_0, i_10_497_3846_0,
    i_10_497_3847_0, i_10_497_3855_0, i_10_497_3856_0, i_10_497_3858_0,
    i_10_497_3915_0, i_10_497_3978_0, i_10_497_3980_0, i_10_497_4023_0,
    i_10_497_4024_0, i_10_497_4028_0, i_10_497_4113_0, i_10_497_4122_0,
    i_10_497_4169_0, i_10_497_4564_0, i_10_497_4566_0, i_10_497_4581_0,
    o_10_497_0_0  );
  input  i_10_497_123_0, i_10_497_216_0, i_10_497_261_0, i_10_497_279_0,
    i_10_497_280_0, i_10_497_281_0, i_10_497_282_0, i_10_497_320_0,
    i_10_497_405_0, i_10_497_443_0, i_10_497_444_0, i_10_497_460_0,
    i_10_497_462_0, i_10_497_904_0, i_10_497_956_0, i_10_497_1053_0,
    i_10_497_1239_0, i_10_497_1263_0, i_10_497_1311_0, i_10_497_1431_0,
    i_10_497_1432_0, i_10_497_1449_0, i_10_497_1539_0, i_10_497_1540_0,
    i_10_497_1542_0, i_10_497_1581_0, i_10_497_1620_0, i_10_497_1629_0,
    i_10_497_1630_0, i_10_497_1651_0, i_10_497_1652_0, i_10_497_1685_0,
    i_10_497_1800_0, i_10_497_1823_0, i_10_497_1944_0, i_10_497_2025_0,
    i_10_497_2026_0, i_10_497_2199_0, i_10_497_2331_0, i_10_497_2351_0,
    i_10_497_2355_0, i_10_497_2403_0, i_10_497_2404_0, i_10_497_2448_0,
    i_10_497_2449_0, i_10_497_2452_0, i_10_497_2470_0, i_10_497_2545_0,
    i_10_497_2565_0, i_10_497_2604_0, i_10_497_2647_0, i_10_497_2662_0,
    i_10_497_2709_0, i_10_497_2718_0, i_10_497_2720_0, i_10_497_2727_0,
    i_10_497_2821_0, i_10_497_2826_0, i_10_497_2844_0, i_10_497_2865_0,
    i_10_497_2961_0, i_10_497_3042_0, i_10_497_3089_0, i_10_497_3278_0,
    i_10_497_3333_0, i_10_497_3386_0, i_10_497_3387_0, i_10_497_3388_0,
    i_10_497_3390_0, i_10_497_3408_0, i_10_497_3468_0, i_10_497_3471_0,
    i_10_497_3537_0, i_10_497_3555_0, i_10_497_3582_0, i_10_497_3610_0,
    i_10_497_3613_0, i_10_497_3618_0, i_10_497_3621_0, i_10_497_3645_0,
    i_10_497_3648_0, i_10_497_3785_0, i_10_497_3840_0, i_10_497_3846_0,
    i_10_497_3847_0, i_10_497_3855_0, i_10_497_3856_0, i_10_497_3858_0,
    i_10_497_3915_0, i_10_497_3978_0, i_10_497_3980_0, i_10_497_4023_0,
    i_10_497_4024_0, i_10_497_4028_0, i_10_497_4113_0, i_10_497_4122_0,
    i_10_497_4169_0, i_10_497_4564_0, i_10_497_4566_0, i_10_497_4581_0;
  output o_10_497_0_0;
  assign o_10_497_0_0 = ~((~i_10_497_3089_0 & ((~i_10_497_123_0 & ((~i_10_497_405_0 & ~i_10_497_1263_0 & ~i_10_497_1539_0 & ~i_10_497_1542_0 & ~i_10_497_1944_0 & ~i_10_497_2025_0 & ~i_10_497_2565_0 & ~i_10_497_3846_0) | (~i_10_497_282_0 & i_10_497_443_0 & ~i_10_497_3613_0 & ~i_10_497_4122_0))) | (~i_10_497_1944_0 & ~i_10_497_2025_0 & ~i_10_497_1542_0 & ~i_10_497_1581_0 & ~i_10_497_2709_0 & ~i_10_497_3613_0 & ~i_10_497_3840_0 & i_10_497_4028_0 & ~i_10_497_4564_0))) | (i_10_497_1542_0 & ((~i_10_497_443_0 & ~i_10_497_1540_0 & i_10_497_1823_0 & i_10_497_2199_0 & ~i_10_497_3978_0) | (~i_10_497_261_0 & ~i_10_497_1651_0 & ~i_10_497_2025_0 & i_10_497_2709_0 & ~i_10_497_2718_0 & i_10_497_3468_0 & ~i_10_497_3856_0 & ~i_10_497_4113_0))) | (~i_10_497_3978_0 & ((~i_10_497_1581_0 & ~i_10_497_4028_0 & ((~i_10_497_216_0 & ~i_10_497_2025_0 & ~i_10_497_2331_0 & ~i_10_497_2718_0 & ~i_10_497_3648_0) | (i_10_497_3648_0 & ~i_10_497_4024_0 & ~i_10_497_4566_0))) | (~i_10_497_2025_0 & ~i_10_497_2351_0 & ~i_10_497_2826_0 & ~i_10_497_3390_0 & ~i_10_497_3846_0 & ~i_10_497_3858_0 & ~i_10_497_3980_0))) | (~i_10_497_2565_0 & ((~i_10_497_216_0 & ((~i_10_497_1263_0 & i_10_497_2826_0 & i_10_497_3388_0 & ~i_10_497_3471_0) | (~i_10_497_261_0 & i_10_497_280_0 & ~i_10_497_2025_0 & ~i_10_497_3390_0 & ~i_10_497_3537_0 & ~i_10_497_3613_0))) | (~i_10_497_261_0 & ((~i_10_497_444_0 & ~i_10_497_2199_0 & ~i_10_497_2355_0 & ~i_10_497_2662_0 & ~i_10_497_3610_0 & ~i_10_497_4023_0) | (~i_10_497_2727_0 & ~i_10_497_3390_0 & ~i_10_497_3855_0 & ~i_10_497_4566_0))) | (~i_10_497_2709_0 & ~i_10_497_2826_0 & ~i_10_497_3855_0 & ~i_10_497_4023_0 & ~i_10_497_4113_0 & ~i_10_497_4564_0 & ~i_10_497_4566_0))) | (i_10_497_1311_0 & ((~i_10_497_444_0 & ((~i_10_497_1944_0 & ~i_10_497_2449_0 & i_10_497_3855_0 & i_10_497_3858_0) | (~i_10_497_3613_0 & ~i_10_497_4024_0 & i_10_497_4028_0))) | (i_10_497_1823_0 & ~i_10_497_2404_0) | (~i_10_497_1542_0 & i_10_497_2604_0))) | (i_10_497_2604_0 & (i_10_497_1823_0 | (~i_10_497_1542_0 & (i_10_497_3858_0 | (~i_10_497_3408_0 & ~i_10_497_3785_0))))) | (i_10_497_1651_0 & ((~i_10_497_1944_0 & ~i_10_497_3388_0 & ~i_10_497_3537_0) | (~i_10_497_3582_0 & ~i_10_497_4023_0))) | (~i_10_497_261_0 & ((~i_10_497_3042_0 & ((i_10_497_462_0 & ~i_10_497_4023_0) | (~i_10_497_1944_0 & ~i_10_497_3785_0 & ~i_10_497_4566_0))) | (i_10_497_1239_0 & ~i_10_497_2355_0 & ~i_10_497_2826_0 & ~i_10_497_4122_0))) | (~i_10_497_1944_0 & ((~i_10_497_1431_0 & i_10_497_3610_0) | (~i_10_497_2403_0 & ~i_10_497_2727_0 & ~i_10_497_3468_0 & ~i_10_497_3840_0 & ~i_10_497_3847_0 & ~i_10_497_4028_0))) | (~i_10_497_4024_0 & ((~i_10_497_279_0 & i_10_497_3089_0 & i_10_497_3610_0) | (~i_10_497_3390_0 & i_10_497_4023_0))) | (i_10_497_2448_0 & ~i_10_497_2709_0 & ~i_10_497_3537_0 & i_10_497_3582_0));
endmodule



// Benchmark "kernel_10_498" written by ABC on Sun Jul 19 10:29:44 2020

module kernel_10_498 ( 
    i_10_498_30_0, i_10_498_34_0, i_10_498_295_0, i_10_498_296_0,
    i_10_498_320_0, i_10_498_322_0, i_10_498_323_0, i_10_498_437_0,
    i_10_498_460_0, i_10_498_629_0, i_10_498_736_0, i_10_498_796_0,
    i_10_498_893_0, i_10_498_895_0, i_10_498_899_0, i_10_498_1033_0,
    i_10_498_1034_0, i_10_498_1154_0, i_10_498_1174_0, i_10_498_1204_0,
    i_10_498_1205_0, i_10_498_1235_0, i_10_498_1238_0, i_10_498_1248_0,
    i_10_498_1249_0, i_10_498_1250_0, i_10_498_1272_0, i_10_498_1349_0,
    i_10_498_1450_0, i_10_498_1545_0, i_10_498_1549_0, i_10_498_1576_0,
    i_10_498_1627_0, i_10_498_1684_0, i_10_498_1685_0, i_10_498_1873_0,
    i_10_498_1874_0, i_10_498_1916_0, i_10_498_1954_0, i_10_498_1994_0,
    i_10_498_2057_0, i_10_498_2165_0, i_10_498_2202_0, i_10_498_2261_0,
    i_10_498_2336_0, i_10_498_2349_0, i_10_498_2350_0, i_10_498_2351_0,
    i_10_498_2363_0, i_10_498_2365_0, i_10_498_2380_0, i_10_498_2381_0,
    i_10_498_2383_0, i_10_498_2384_0, i_10_498_2454_0, i_10_498_2455_0,
    i_10_498_2465_0, i_10_498_2473_0, i_10_498_2571_0, i_10_498_2572_0,
    i_10_498_2633_0, i_10_498_2710_0, i_10_498_2716_0, i_10_498_2717_0,
    i_10_498_2722_0, i_10_498_2726_0, i_10_498_2730_0, i_10_498_2832_0,
    i_10_498_2869_0, i_10_498_2880_0, i_10_498_2881_0, i_10_498_2882_0,
    i_10_498_2920_0, i_10_498_2957_0, i_10_498_2991_0, i_10_498_3049_0,
    i_10_498_3072_0, i_10_498_3355_0, i_10_498_3403_0, i_10_498_3470_0,
    i_10_498_3571_0, i_10_498_3572_0, i_10_498_3612_0, i_10_498_3723_0,
    i_10_498_3724_0, i_10_498_3732_0, i_10_498_3784_0, i_10_498_3860_0,
    i_10_498_3981_0, i_10_498_4029_0, i_10_498_4030_0, i_10_498_4119_0,
    i_10_498_4129_0, i_10_498_4130_0, i_10_498_4220_0, i_10_498_4272_0,
    i_10_498_4289_0, i_10_498_4426_0, i_10_498_4427_0, i_10_498_4583_0,
    o_10_498_0_0  );
  input  i_10_498_30_0, i_10_498_34_0, i_10_498_295_0, i_10_498_296_0,
    i_10_498_320_0, i_10_498_322_0, i_10_498_323_0, i_10_498_437_0,
    i_10_498_460_0, i_10_498_629_0, i_10_498_736_0, i_10_498_796_0,
    i_10_498_893_0, i_10_498_895_0, i_10_498_899_0, i_10_498_1033_0,
    i_10_498_1034_0, i_10_498_1154_0, i_10_498_1174_0, i_10_498_1204_0,
    i_10_498_1205_0, i_10_498_1235_0, i_10_498_1238_0, i_10_498_1248_0,
    i_10_498_1249_0, i_10_498_1250_0, i_10_498_1272_0, i_10_498_1349_0,
    i_10_498_1450_0, i_10_498_1545_0, i_10_498_1549_0, i_10_498_1576_0,
    i_10_498_1627_0, i_10_498_1684_0, i_10_498_1685_0, i_10_498_1873_0,
    i_10_498_1874_0, i_10_498_1916_0, i_10_498_1954_0, i_10_498_1994_0,
    i_10_498_2057_0, i_10_498_2165_0, i_10_498_2202_0, i_10_498_2261_0,
    i_10_498_2336_0, i_10_498_2349_0, i_10_498_2350_0, i_10_498_2351_0,
    i_10_498_2363_0, i_10_498_2365_0, i_10_498_2380_0, i_10_498_2381_0,
    i_10_498_2383_0, i_10_498_2384_0, i_10_498_2454_0, i_10_498_2455_0,
    i_10_498_2465_0, i_10_498_2473_0, i_10_498_2571_0, i_10_498_2572_0,
    i_10_498_2633_0, i_10_498_2710_0, i_10_498_2716_0, i_10_498_2717_0,
    i_10_498_2722_0, i_10_498_2726_0, i_10_498_2730_0, i_10_498_2832_0,
    i_10_498_2869_0, i_10_498_2880_0, i_10_498_2881_0, i_10_498_2882_0,
    i_10_498_2920_0, i_10_498_2957_0, i_10_498_2991_0, i_10_498_3049_0,
    i_10_498_3072_0, i_10_498_3355_0, i_10_498_3403_0, i_10_498_3470_0,
    i_10_498_3571_0, i_10_498_3572_0, i_10_498_3612_0, i_10_498_3723_0,
    i_10_498_3724_0, i_10_498_3732_0, i_10_498_3784_0, i_10_498_3860_0,
    i_10_498_3981_0, i_10_498_4029_0, i_10_498_4030_0, i_10_498_4119_0,
    i_10_498_4129_0, i_10_498_4130_0, i_10_498_4220_0, i_10_498_4272_0,
    i_10_498_4289_0, i_10_498_4426_0, i_10_498_4427_0, i_10_498_4583_0;
  output o_10_498_0_0;
  assign o_10_498_0_0 = 0;
endmodule



// Benchmark "kernel_10_499" written by ABC on Sun Jul 19 10:29:44 2020

module kernel_10_499 ( 
    i_10_499_36_0, i_10_499_156_0, i_10_499_181_0, i_10_499_216_0,
    i_10_499_245_0, i_10_499_246_0, i_10_499_247_0, i_10_499_284_0,
    i_10_499_316_0, i_10_499_319_0, i_10_499_330_0, i_10_499_393_0,
    i_10_499_409_0, i_10_499_436_0, i_10_499_446_0, i_10_499_459_0,
    i_10_499_460_0, i_10_499_559_0, i_10_499_754_0, i_10_499_792_0,
    i_10_499_892_0, i_10_499_993_0, i_10_499_1000_0, i_10_499_1035_0,
    i_10_499_1039_0, i_10_499_1047_0, i_10_499_1048_0, i_10_499_1059_0,
    i_10_499_1152_0, i_10_499_1164_0, i_10_499_1215_0, i_10_499_1235_0,
    i_10_499_1237_0, i_10_499_1306_0, i_10_499_1307_0, i_10_499_1311_0,
    i_10_499_1312_0, i_10_499_1313_0, i_10_499_1362_0, i_10_499_1539_0,
    i_10_499_1575_0, i_10_499_1594_0, i_10_499_1648_0, i_10_499_1650_0,
    i_10_499_1655_0, i_10_499_1688_0, i_10_499_1690_0, i_10_499_1914_0,
    i_10_499_2016_0, i_10_499_2019_0, i_10_499_2199_0, i_10_499_2349_0,
    i_10_499_2356_0, i_10_499_2601_0, i_10_499_2603_0, i_10_499_2606_0,
    i_10_499_2634_0, i_10_499_2635_0, i_10_499_2705_0, i_10_499_2724_0,
    i_10_499_2728_0, i_10_499_2730_0, i_10_499_2784_0, i_10_499_2785_0,
    i_10_499_2831_0, i_10_499_2881_0, i_10_499_2983_0, i_10_499_2985_0,
    i_10_499_3073_0, i_10_499_3159_0, i_10_499_3162_0, i_10_499_3231_0,
    i_10_499_3270_0, i_10_499_3328_0, i_10_499_3406_0, i_10_499_3429_0,
    i_10_499_3430_0, i_10_499_3501_0, i_10_499_3519_0, i_10_499_3609_0,
    i_10_499_3610_0, i_10_499_3717_0, i_10_499_3721_0, i_10_499_3785_0,
    i_10_499_3787_0, i_10_499_3788_0, i_10_499_3810_0, i_10_499_3850_0,
    i_10_499_3856_0, i_10_499_3859_0, i_10_499_3860_0, i_10_499_3883_0,
    i_10_499_3889_0, i_10_499_3987_0, i_10_499_4062_0, i_10_499_4168_0,
    i_10_499_4173_0, i_10_499_4278_0, i_10_499_4570_0, i_10_499_4586_0,
    o_10_499_0_0  );
  input  i_10_499_36_0, i_10_499_156_0, i_10_499_181_0, i_10_499_216_0,
    i_10_499_245_0, i_10_499_246_0, i_10_499_247_0, i_10_499_284_0,
    i_10_499_316_0, i_10_499_319_0, i_10_499_330_0, i_10_499_393_0,
    i_10_499_409_0, i_10_499_436_0, i_10_499_446_0, i_10_499_459_0,
    i_10_499_460_0, i_10_499_559_0, i_10_499_754_0, i_10_499_792_0,
    i_10_499_892_0, i_10_499_993_0, i_10_499_1000_0, i_10_499_1035_0,
    i_10_499_1039_0, i_10_499_1047_0, i_10_499_1048_0, i_10_499_1059_0,
    i_10_499_1152_0, i_10_499_1164_0, i_10_499_1215_0, i_10_499_1235_0,
    i_10_499_1237_0, i_10_499_1306_0, i_10_499_1307_0, i_10_499_1311_0,
    i_10_499_1312_0, i_10_499_1313_0, i_10_499_1362_0, i_10_499_1539_0,
    i_10_499_1575_0, i_10_499_1594_0, i_10_499_1648_0, i_10_499_1650_0,
    i_10_499_1655_0, i_10_499_1688_0, i_10_499_1690_0, i_10_499_1914_0,
    i_10_499_2016_0, i_10_499_2019_0, i_10_499_2199_0, i_10_499_2349_0,
    i_10_499_2356_0, i_10_499_2601_0, i_10_499_2603_0, i_10_499_2606_0,
    i_10_499_2634_0, i_10_499_2635_0, i_10_499_2705_0, i_10_499_2724_0,
    i_10_499_2728_0, i_10_499_2730_0, i_10_499_2784_0, i_10_499_2785_0,
    i_10_499_2831_0, i_10_499_2881_0, i_10_499_2983_0, i_10_499_2985_0,
    i_10_499_3073_0, i_10_499_3159_0, i_10_499_3162_0, i_10_499_3231_0,
    i_10_499_3270_0, i_10_499_3328_0, i_10_499_3406_0, i_10_499_3429_0,
    i_10_499_3430_0, i_10_499_3501_0, i_10_499_3519_0, i_10_499_3609_0,
    i_10_499_3610_0, i_10_499_3717_0, i_10_499_3721_0, i_10_499_3785_0,
    i_10_499_3787_0, i_10_499_3788_0, i_10_499_3810_0, i_10_499_3850_0,
    i_10_499_3856_0, i_10_499_3859_0, i_10_499_3860_0, i_10_499_3883_0,
    i_10_499_3889_0, i_10_499_3987_0, i_10_499_4062_0, i_10_499_4168_0,
    i_10_499_4173_0, i_10_499_4278_0, i_10_499_4570_0, i_10_499_4586_0;
  output o_10_499_0_0;
  assign o_10_499_0_0 = 0;
endmodule



// Benchmark "kernel_10_500" written by ABC on Sun Jul 19 10:29:45 2020

module kernel_10_500 ( 
    i_10_500_121_0, i_10_500_146_0, i_10_500_175_0, i_10_500_254_0,
    i_10_500_256_0, i_10_500_257_0, i_10_500_283_0, i_10_500_288_0,
    i_10_500_325_0, i_10_500_394_0, i_10_500_441_0, i_10_500_445_0,
    i_10_500_562_0, i_10_500_632_0, i_10_500_796_0, i_10_500_797_0,
    i_10_500_800_0, i_10_500_920_0, i_10_500_955_0, i_10_500_963_0,
    i_10_500_1118_0, i_10_500_1235_0, i_10_500_1236_0, i_10_500_1237_0,
    i_10_500_1238_0, i_10_500_1245_0, i_10_500_1249_0, i_10_500_1250_0,
    i_10_500_1268_0, i_10_500_1313_0, i_10_500_1361_0, i_10_500_1650_0,
    i_10_500_1683_0, i_10_500_1685_0, i_10_500_1687_0, i_10_500_1721_0,
    i_10_500_1724_0, i_10_500_1821_0, i_10_500_1824_0, i_10_500_1825_0,
    i_10_500_1826_0, i_10_500_1883_0, i_10_500_1915_0, i_10_500_1919_0,
    i_10_500_1984_0, i_10_500_2107_0, i_10_500_2243_0, i_10_500_2350_0,
    i_10_500_2352_0, i_10_500_2387_0, i_10_500_2390_0, i_10_500_2453_0,
    i_10_500_2471_0, i_10_500_2659_0, i_10_500_2663_0, i_10_500_2711_0,
    i_10_500_2719_0, i_10_500_2723_0, i_10_500_2737_0, i_10_500_2786_0,
    i_10_500_2827_0, i_10_500_2834_0, i_10_500_2846_0, i_10_500_2981_0,
    i_10_500_3236_0, i_10_500_3280_0, i_10_500_3283_0, i_10_500_3386_0,
    i_10_500_3388_0, i_10_500_3389_0, i_10_500_3431_0, i_10_500_3467_0,
    i_10_500_3494_0, i_10_500_3523_0, i_10_500_3524_0, i_10_500_3539_0,
    i_10_500_3545_0, i_10_500_3584_0, i_10_500_3586_0, i_10_500_3587_0,
    i_10_500_3720_0, i_10_500_3847_0, i_10_500_3872_0, i_10_500_3943_0,
    i_10_500_3944_0, i_10_500_3982_0, i_10_500_3998_0, i_10_500_4054_0,
    i_10_500_4130_0, i_10_500_4151_0, i_10_500_4231_0, i_10_500_4268_0,
    i_10_500_4271_0, i_10_500_4274_0, i_10_500_4275_0, i_10_500_4279_0,
    i_10_500_4460_0, i_10_500_4569_0, i_10_500_4571_0, i_10_500_4583_0,
    o_10_500_0_0  );
  input  i_10_500_121_0, i_10_500_146_0, i_10_500_175_0, i_10_500_254_0,
    i_10_500_256_0, i_10_500_257_0, i_10_500_283_0, i_10_500_288_0,
    i_10_500_325_0, i_10_500_394_0, i_10_500_441_0, i_10_500_445_0,
    i_10_500_562_0, i_10_500_632_0, i_10_500_796_0, i_10_500_797_0,
    i_10_500_800_0, i_10_500_920_0, i_10_500_955_0, i_10_500_963_0,
    i_10_500_1118_0, i_10_500_1235_0, i_10_500_1236_0, i_10_500_1237_0,
    i_10_500_1238_0, i_10_500_1245_0, i_10_500_1249_0, i_10_500_1250_0,
    i_10_500_1268_0, i_10_500_1313_0, i_10_500_1361_0, i_10_500_1650_0,
    i_10_500_1683_0, i_10_500_1685_0, i_10_500_1687_0, i_10_500_1721_0,
    i_10_500_1724_0, i_10_500_1821_0, i_10_500_1824_0, i_10_500_1825_0,
    i_10_500_1826_0, i_10_500_1883_0, i_10_500_1915_0, i_10_500_1919_0,
    i_10_500_1984_0, i_10_500_2107_0, i_10_500_2243_0, i_10_500_2350_0,
    i_10_500_2352_0, i_10_500_2387_0, i_10_500_2390_0, i_10_500_2453_0,
    i_10_500_2471_0, i_10_500_2659_0, i_10_500_2663_0, i_10_500_2711_0,
    i_10_500_2719_0, i_10_500_2723_0, i_10_500_2737_0, i_10_500_2786_0,
    i_10_500_2827_0, i_10_500_2834_0, i_10_500_2846_0, i_10_500_2981_0,
    i_10_500_3236_0, i_10_500_3280_0, i_10_500_3283_0, i_10_500_3386_0,
    i_10_500_3388_0, i_10_500_3389_0, i_10_500_3431_0, i_10_500_3467_0,
    i_10_500_3494_0, i_10_500_3523_0, i_10_500_3524_0, i_10_500_3539_0,
    i_10_500_3545_0, i_10_500_3584_0, i_10_500_3586_0, i_10_500_3587_0,
    i_10_500_3720_0, i_10_500_3847_0, i_10_500_3872_0, i_10_500_3943_0,
    i_10_500_3944_0, i_10_500_3982_0, i_10_500_3998_0, i_10_500_4054_0,
    i_10_500_4130_0, i_10_500_4151_0, i_10_500_4231_0, i_10_500_4268_0,
    i_10_500_4271_0, i_10_500_4274_0, i_10_500_4275_0, i_10_500_4279_0,
    i_10_500_4460_0, i_10_500_4569_0, i_10_500_4571_0, i_10_500_4583_0;
  output o_10_500_0_0;
  assign o_10_500_0_0 = 0;
endmodule



// Benchmark "kernel_10_501" written by ABC on Sun Jul 19 10:29:46 2020

module kernel_10_501 ( 
    i_10_501_27_0, i_10_501_146_0, i_10_501_154_0, i_10_501_173_0,
    i_10_501_289_0, i_10_501_290_0, i_10_501_406_0, i_10_501_423_0,
    i_10_501_428_0, i_10_501_626_0, i_10_501_640_0, i_10_501_821_0,
    i_10_501_848_0, i_10_501_901_0, i_10_501_992_0, i_10_501_1028_0,
    i_10_501_1046_0, i_10_501_1118_0, i_10_501_1238_0, i_10_501_1253_0,
    i_10_501_1289_0, i_10_501_1442_0, i_10_501_1612_0, i_10_501_1613_0,
    i_10_501_1631_0, i_10_501_1648_0, i_10_501_1652_0, i_10_501_1689_0,
    i_10_501_1738_0, i_10_501_1757_0, i_10_501_1759_0, i_10_501_1873_0,
    i_10_501_1874_0, i_10_501_1954_0, i_10_501_1991_0, i_10_501_2216_0,
    i_10_501_2225_0, i_10_501_2288_0, i_10_501_2327_0, i_10_501_2359_0,
    i_10_501_2362_0, i_10_501_2441_0, i_10_501_2469_0, i_10_501_2476_0,
    i_10_501_2477_0, i_10_501_2511_0, i_10_501_2525_0, i_10_501_2566_0,
    i_10_501_2567_0, i_10_501_2603_0, i_10_501_2631_0, i_10_501_2636_0,
    i_10_501_2642_0, i_10_501_2648_0, i_10_501_2651_0, i_10_501_2657_0,
    i_10_501_2675_0, i_10_501_2719_0, i_10_501_2729_0, i_10_501_2738_0,
    i_10_501_2829_0, i_10_501_2833_0, i_10_501_2882_0, i_10_501_2917_0,
    i_10_501_2918_0, i_10_501_2923_0, i_10_501_3161_0, i_10_501_3195_0,
    i_10_501_3233_0, i_10_501_3286_0, i_10_501_3290_0, i_10_501_3405_0,
    i_10_501_3410_0, i_10_501_3440_0, i_10_501_3449_0, i_10_501_3557_0,
    i_10_501_3620_0, i_10_501_3686_0, i_10_501_3728_0, i_10_501_3827_0,
    i_10_501_3830_0, i_10_501_3852_0, i_10_501_3855_0, i_10_501_3899_0,
    i_10_501_4025_0, i_10_501_4028_0, i_10_501_4114_0, i_10_501_4115_0,
    i_10_501_4144_0, i_10_501_4145_0, i_10_501_4151_0, i_10_501_4189_0,
    i_10_501_4214_0, i_10_501_4291_0, i_10_501_4292_0, i_10_501_4307_0,
    i_10_501_4456_0, i_10_501_4501_0, i_10_501_4502_0, i_10_501_4563_0,
    o_10_501_0_0  );
  input  i_10_501_27_0, i_10_501_146_0, i_10_501_154_0, i_10_501_173_0,
    i_10_501_289_0, i_10_501_290_0, i_10_501_406_0, i_10_501_423_0,
    i_10_501_428_0, i_10_501_626_0, i_10_501_640_0, i_10_501_821_0,
    i_10_501_848_0, i_10_501_901_0, i_10_501_992_0, i_10_501_1028_0,
    i_10_501_1046_0, i_10_501_1118_0, i_10_501_1238_0, i_10_501_1253_0,
    i_10_501_1289_0, i_10_501_1442_0, i_10_501_1612_0, i_10_501_1613_0,
    i_10_501_1631_0, i_10_501_1648_0, i_10_501_1652_0, i_10_501_1689_0,
    i_10_501_1738_0, i_10_501_1757_0, i_10_501_1759_0, i_10_501_1873_0,
    i_10_501_1874_0, i_10_501_1954_0, i_10_501_1991_0, i_10_501_2216_0,
    i_10_501_2225_0, i_10_501_2288_0, i_10_501_2327_0, i_10_501_2359_0,
    i_10_501_2362_0, i_10_501_2441_0, i_10_501_2469_0, i_10_501_2476_0,
    i_10_501_2477_0, i_10_501_2511_0, i_10_501_2525_0, i_10_501_2566_0,
    i_10_501_2567_0, i_10_501_2603_0, i_10_501_2631_0, i_10_501_2636_0,
    i_10_501_2642_0, i_10_501_2648_0, i_10_501_2651_0, i_10_501_2657_0,
    i_10_501_2675_0, i_10_501_2719_0, i_10_501_2729_0, i_10_501_2738_0,
    i_10_501_2829_0, i_10_501_2833_0, i_10_501_2882_0, i_10_501_2917_0,
    i_10_501_2918_0, i_10_501_2923_0, i_10_501_3161_0, i_10_501_3195_0,
    i_10_501_3233_0, i_10_501_3286_0, i_10_501_3290_0, i_10_501_3405_0,
    i_10_501_3410_0, i_10_501_3440_0, i_10_501_3449_0, i_10_501_3557_0,
    i_10_501_3620_0, i_10_501_3686_0, i_10_501_3728_0, i_10_501_3827_0,
    i_10_501_3830_0, i_10_501_3852_0, i_10_501_3855_0, i_10_501_3899_0,
    i_10_501_4025_0, i_10_501_4028_0, i_10_501_4114_0, i_10_501_4115_0,
    i_10_501_4144_0, i_10_501_4145_0, i_10_501_4151_0, i_10_501_4189_0,
    i_10_501_4214_0, i_10_501_4291_0, i_10_501_4292_0, i_10_501_4307_0,
    i_10_501_4456_0, i_10_501_4501_0, i_10_501_4502_0, i_10_501_4563_0;
  output o_10_501_0_0;
  assign o_10_501_0_0 = 0;
endmodule



// Benchmark "kernel_10_502" written by ABC on Sun Jul 19 10:29:47 2020

module kernel_10_502 ( 
    i_10_502_33_0, i_10_502_34_0, i_10_502_70_0, i_10_502_179_0,
    i_10_502_208_0, i_10_502_248_0, i_10_502_430_0, i_10_502_431_0,
    i_10_502_444_0, i_10_502_448_0, i_10_502_562_0, i_10_502_563_0,
    i_10_502_719_0, i_10_502_796_0, i_10_502_799_0, i_10_502_820_0,
    i_10_502_823_0, i_10_502_953_0, i_10_502_996_0, i_10_502_1004_0,
    i_10_502_1006_0, i_10_502_1007_0, i_10_502_1052_0, i_10_502_1213_0,
    i_10_502_1247_0, i_10_502_1322_0, i_10_502_1348_0, i_10_502_1349_0,
    i_10_502_1366_0, i_10_502_1367_0, i_10_502_1383_0, i_10_502_1384_0,
    i_10_502_1492_0, i_10_502_1493_0, i_10_502_1565_0, i_10_502_1627_0,
    i_10_502_1628_0, i_10_502_1631_0, i_10_502_1634_0, i_10_502_1655_0,
    i_10_502_1697_0, i_10_502_1736_0, i_10_502_1768_0, i_10_502_1912_0,
    i_10_502_1937_0, i_10_502_2038_0, i_10_502_2041_0, i_10_502_2042_0,
    i_10_502_2159_0, i_10_502_2264_0, i_10_502_2410_0, i_10_502_2437_0,
    i_10_502_2474_0, i_10_502_2508_0, i_10_502_2509_0, i_10_502_2514_0,
    i_10_502_2517_0, i_10_502_2636_0, i_10_502_2661_0, i_10_502_2679_0,
    i_10_502_2698_0, i_10_502_2699_0, i_10_502_2707_0, i_10_502_2708_0,
    i_10_502_2714_0, i_10_502_2744_0, i_10_502_2757_0, i_10_502_2758_0,
    i_10_502_2824_0, i_10_502_2830_0, i_10_502_2852_0, i_10_502_2870_0,
    i_10_502_2885_0, i_10_502_3048_0, i_10_502_3050_0, i_10_502_3094_0,
    i_10_502_3095_0, i_10_502_3284_0, i_10_502_3319_0, i_10_502_3320_0,
    i_10_502_3415_0, i_10_502_3436_0, i_10_502_3472_0, i_10_502_3494_0,
    i_10_502_3588_0, i_10_502_3611_0, i_10_502_3612_0, i_10_502_3625_0,
    i_10_502_3640_0, i_10_502_3704_0, i_10_502_3706_0, i_10_502_3707_0,
    i_10_502_3853_0, i_10_502_3986_0, i_10_502_4237_0, i_10_502_4267_0,
    i_10_502_4268_0, i_10_502_4271_0, i_10_502_4289_0, i_10_502_4454_0,
    o_10_502_0_0  );
  input  i_10_502_33_0, i_10_502_34_0, i_10_502_70_0, i_10_502_179_0,
    i_10_502_208_0, i_10_502_248_0, i_10_502_430_0, i_10_502_431_0,
    i_10_502_444_0, i_10_502_448_0, i_10_502_562_0, i_10_502_563_0,
    i_10_502_719_0, i_10_502_796_0, i_10_502_799_0, i_10_502_820_0,
    i_10_502_823_0, i_10_502_953_0, i_10_502_996_0, i_10_502_1004_0,
    i_10_502_1006_0, i_10_502_1007_0, i_10_502_1052_0, i_10_502_1213_0,
    i_10_502_1247_0, i_10_502_1322_0, i_10_502_1348_0, i_10_502_1349_0,
    i_10_502_1366_0, i_10_502_1367_0, i_10_502_1383_0, i_10_502_1384_0,
    i_10_502_1492_0, i_10_502_1493_0, i_10_502_1565_0, i_10_502_1627_0,
    i_10_502_1628_0, i_10_502_1631_0, i_10_502_1634_0, i_10_502_1655_0,
    i_10_502_1697_0, i_10_502_1736_0, i_10_502_1768_0, i_10_502_1912_0,
    i_10_502_1937_0, i_10_502_2038_0, i_10_502_2041_0, i_10_502_2042_0,
    i_10_502_2159_0, i_10_502_2264_0, i_10_502_2410_0, i_10_502_2437_0,
    i_10_502_2474_0, i_10_502_2508_0, i_10_502_2509_0, i_10_502_2514_0,
    i_10_502_2517_0, i_10_502_2636_0, i_10_502_2661_0, i_10_502_2679_0,
    i_10_502_2698_0, i_10_502_2699_0, i_10_502_2707_0, i_10_502_2708_0,
    i_10_502_2714_0, i_10_502_2744_0, i_10_502_2757_0, i_10_502_2758_0,
    i_10_502_2824_0, i_10_502_2830_0, i_10_502_2852_0, i_10_502_2870_0,
    i_10_502_2885_0, i_10_502_3048_0, i_10_502_3050_0, i_10_502_3094_0,
    i_10_502_3095_0, i_10_502_3284_0, i_10_502_3319_0, i_10_502_3320_0,
    i_10_502_3415_0, i_10_502_3436_0, i_10_502_3472_0, i_10_502_3494_0,
    i_10_502_3588_0, i_10_502_3611_0, i_10_502_3612_0, i_10_502_3625_0,
    i_10_502_3640_0, i_10_502_3704_0, i_10_502_3706_0, i_10_502_3707_0,
    i_10_502_3853_0, i_10_502_3986_0, i_10_502_4237_0, i_10_502_4267_0,
    i_10_502_4268_0, i_10_502_4271_0, i_10_502_4289_0, i_10_502_4454_0;
  output o_10_502_0_0;
  assign o_10_502_0_0 = 0;
endmodule



// Benchmark "kernel_10_503" written by ABC on Sun Jul 19 10:29:48 2020

module kernel_10_503 ( 
    i_10_503_31_0, i_10_503_280_0, i_10_503_282_0, i_10_503_283_0,
    i_10_503_284_0, i_10_503_285_0, i_10_503_290_0, i_10_503_316_0,
    i_10_503_438_0, i_10_503_439_0, i_10_503_463_0, i_10_503_519_0,
    i_10_503_717_0, i_10_503_955_0, i_10_503_1005_0, i_10_503_1234_0,
    i_10_503_1235_0, i_10_503_1236_0, i_10_503_1435_0, i_10_503_1445_0,
    i_10_503_1648_0, i_10_503_1678_0, i_10_503_1679_0, i_10_503_1689_0,
    i_10_503_1819_0, i_10_503_1820_0, i_10_503_1821_0, i_10_503_1915_0,
    i_10_503_2027_0, i_10_503_2029_0, i_10_503_2031_0, i_10_503_2352_0,
    i_10_503_2353_0, i_10_503_2354_0, i_10_503_2357_0, i_10_503_2408_0,
    i_10_503_2449_0, i_10_503_2460_0, i_10_503_2467_0, i_10_503_2628_0,
    i_10_503_2630_0, i_10_503_2660_0, i_10_503_2662_0, i_10_503_2675_0,
    i_10_503_2711_0, i_10_503_2716_0, i_10_503_2722_0, i_10_503_2728_0,
    i_10_503_2729_0, i_10_503_2832_0, i_10_503_2833_0, i_10_503_2881_0,
    i_10_503_2885_0, i_10_503_2888_0, i_10_503_2917_0, i_10_503_2922_0,
    i_10_503_2923_0, i_10_503_2985_0, i_10_503_2987_0, i_10_503_3038_0,
    i_10_503_3040_0, i_10_503_3043_0, i_10_503_3044_0, i_10_503_3196_0,
    i_10_503_3198_0, i_10_503_3199_0, i_10_503_3384_0, i_10_503_3387_0,
    i_10_503_3388_0, i_10_503_3391_0, i_10_503_3405_0, i_10_503_3409_0,
    i_10_503_3497_0, i_10_503_3589_0, i_10_503_3610_0, i_10_503_3611_0,
    i_10_503_3614_0, i_10_503_3650_0, i_10_503_3782_0, i_10_503_3784_0,
    i_10_503_3785_0, i_10_503_3837_0, i_10_503_3840_0, i_10_503_3848_0,
    i_10_503_3858_0, i_10_503_3859_0, i_10_503_3907_0, i_10_503_4025_0,
    i_10_503_4123_0, i_10_503_4124_0, i_10_503_4127_0, i_10_503_4269_0,
    i_10_503_4270_0, i_10_503_4271_0, i_10_503_4278_0, i_10_503_4286_0,
    i_10_503_4292_0, i_10_503_4567_0, i_10_503_4568_0, i_10_503_4569_0,
    o_10_503_0_0  );
  input  i_10_503_31_0, i_10_503_280_0, i_10_503_282_0, i_10_503_283_0,
    i_10_503_284_0, i_10_503_285_0, i_10_503_290_0, i_10_503_316_0,
    i_10_503_438_0, i_10_503_439_0, i_10_503_463_0, i_10_503_519_0,
    i_10_503_717_0, i_10_503_955_0, i_10_503_1005_0, i_10_503_1234_0,
    i_10_503_1235_0, i_10_503_1236_0, i_10_503_1435_0, i_10_503_1445_0,
    i_10_503_1648_0, i_10_503_1678_0, i_10_503_1679_0, i_10_503_1689_0,
    i_10_503_1819_0, i_10_503_1820_0, i_10_503_1821_0, i_10_503_1915_0,
    i_10_503_2027_0, i_10_503_2029_0, i_10_503_2031_0, i_10_503_2352_0,
    i_10_503_2353_0, i_10_503_2354_0, i_10_503_2357_0, i_10_503_2408_0,
    i_10_503_2449_0, i_10_503_2460_0, i_10_503_2467_0, i_10_503_2628_0,
    i_10_503_2630_0, i_10_503_2660_0, i_10_503_2662_0, i_10_503_2675_0,
    i_10_503_2711_0, i_10_503_2716_0, i_10_503_2722_0, i_10_503_2728_0,
    i_10_503_2729_0, i_10_503_2832_0, i_10_503_2833_0, i_10_503_2881_0,
    i_10_503_2885_0, i_10_503_2888_0, i_10_503_2917_0, i_10_503_2922_0,
    i_10_503_2923_0, i_10_503_2985_0, i_10_503_2987_0, i_10_503_3038_0,
    i_10_503_3040_0, i_10_503_3043_0, i_10_503_3044_0, i_10_503_3196_0,
    i_10_503_3198_0, i_10_503_3199_0, i_10_503_3384_0, i_10_503_3387_0,
    i_10_503_3388_0, i_10_503_3391_0, i_10_503_3405_0, i_10_503_3409_0,
    i_10_503_3497_0, i_10_503_3589_0, i_10_503_3610_0, i_10_503_3611_0,
    i_10_503_3614_0, i_10_503_3650_0, i_10_503_3782_0, i_10_503_3784_0,
    i_10_503_3785_0, i_10_503_3837_0, i_10_503_3840_0, i_10_503_3848_0,
    i_10_503_3858_0, i_10_503_3859_0, i_10_503_3907_0, i_10_503_4025_0,
    i_10_503_4123_0, i_10_503_4124_0, i_10_503_4127_0, i_10_503_4269_0,
    i_10_503_4270_0, i_10_503_4271_0, i_10_503_4278_0, i_10_503_4286_0,
    i_10_503_4292_0, i_10_503_4567_0, i_10_503_4568_0, i_10_503_4569_0;
  output o_10_503_0_0;
  assign o_10_503_0_0 = ~((~i_10_503_1689_0 & ((~i_10_503_284_0 & ~i_10_503_3043_0 & i_10_503_3859_0 & ~i_10_503_4127_0 & ~i_10_503_4286_0) | (~i_10_503_1234_0 & ~i_10_503_1235_0 & ~i_10_503_1445_0 & ~i_10_503_2354_0 & ~i_10_503_2467_0 & ~i_10_503_3044_0 & ~i_10_503_4123_0 & ~i_10_503_4567_0))) | (~i_10_503_1821_0 & ((~i_10_503_285_0 & i_10_503_1689_0 & ~i_10_503_3405_0 & ~i_10_503_3614_0 & ~i_10_503_4269_0 & ~i_10_503_4270_0 & ~i_10_503_4568_0) | (~i_10_503_1235_0 & ~i_10_503_2716_0 & ~i_10_503_2722_0 & ~i_10_503_2833_0 & ~i_10_503_3043_0 & ~i_10_503_3388_0 & ~i_10_503_3497_0 & ~i_10_503_3650_0 & ~i_10_503_4569_0))) | (~i_10_503_3391_0 & ((~i_10_503_285_0 & ((i_10_503_1005_0 & ~i_10_503_2354_0 & ~i_10_503_2728_0 & i_10_503_3837_0) | (~i_10_503_283_0 & ~i_10_503_284_0 & ~i_10_503_1445_0 & ~i_10_503_2031_0 & ~i_10_503_2408_0 & ~i_10_503_3497_0 & ~i_10_503_4124_0 & ~i_10_503_4278_0))) | (~i_10_503_316_0 & ~i_10_503_3043_0 & ~i_10_503_4568_0 & ((~i_10_503_280_0 & ~i_10_503_1005_0 & ~i_10_503_1445_0 & ~i_10_503_2408_0 & ~i_10_503_3409_0 & ~i_10_503_3859_0 & ~i_10_503_4025_0 & ~i_10_503_4127_0 & ~i_10_503_4269_0 & ~i_10_503_4270_0) | (~i_10_503_717_0 & ~i_10_503_2031_0 & i_10_503_2352_0 & ~i_10_503_3038_0 & ~i_10_503_4271_0 & ~i_10_503_4569_0))) | (i_10_503_463_0 & ~i_10_503_1235_0 & ~i_10_503_2357_0 & ~i_10_503_3044_0 & ~i_10_503_3384_0 & ~i_10_503_3388_0 & ~i_10_503_3782_0 & ~i_10_503_4123_0 & ~i_10_503_4124_0))) | (~i_10_503_280_0 & ((~i_10_503_284_0 & ~i_10_503_2352_0 & i_10_503_3610_0) | (~i_10_503_439_0 & ~i_10_503_717_0 & ~i_10_503_1234_0 & ~i_10_503_1235_0 & ~i_10_503_1445_0 & ~i_10_503_2031_0 & ~i_10_503_2354_0 & ~i_10_503_2357_0 & ~i_10_503_2467_0 & ~i_10_503_3907_0 & ~i_10_503_4269_0 & ~i_10_503_4286_0))) | (~i_10_503_4127_0 & ((~i_10_503_1234_0 & ((~i_10_503_284_0 & ~i_10_503_2352_0 & ~i_10_503_2711_0 & ~i_10_503_2985_0 & ~i_10_503_2987_0 & ~i_10_503_3043_0 & ~i_10_503_3907_0 & ~i_10_503_4123_0) | (~i_10_503_2353_0 & ~i_10_503_2660_0 & ~i_10_503_2728_0 & ~i_10_503_3497_0 & ~i_10_503_3859_0 & ~i_10_503_4278_0 & ~i_10_503_4286_0))) | (~i_10_503_2027_0 & ~i_10_503_2354_0 & ~i_10_503_2660_0 & i_10_503_3405_0) | (i_10_503_2449_0 & ~i_10_503_3405_0 & i_10_503_3610_0 & ~i_10_503_4124_0) | (~i_10_503_717_0 & ~i_10_503_2729_0 & ~i_10_503_3044_0 & ~i_10_503_3384_0 & ~i_10_503_3388_0 & ~i_10_503_3589_0 & ~i_10_503_3840_0 & ~i_10_503_3907_0 & ~i_10_503_4270_0 & ~i_10_503_4271_0 & ~i_10_503_4567_0))) | (~i_10_503_284_0 & ((~i_10_503_717_0 & ~i_10_503_2027_0 & i_10_503_2922_0 & ~i_10_503_3043_0) | (~i_10_503_283_0 & ~i_10_503_519_0 & ~i_10_503_1819_0 & i_10_503_2353_0 & ~i_10_503_2675_0 & ~i_10_503_3840_0 & ~i_10_503_4124_0 & ~i_10_503_4286_0 & ~i_10_503_4569_0))) | (~i_10_503_2675_0 & ((~i_10_503_283_0 & ((~i_10_503_1005_0 & ~i_10_503_2357_0 & ~i_10_503_2467_0 & ~i_10_503_2728_0 & ~i_10_503_2987_0 & ~i_10_503_3044_0 & ~i_10_503_3589_0 & ~i_10_503_4123_0) | (~i_10_503_2031_0 & ~i_10_503_3388_0 & ~i_10_503_3497_0 & ~i_10_503_3650_0 & ~i_10_503_4025_0 & i_10_503_4270_0 & i_10_503_4567_0))) | (~i_10_503_3497_0 & ((~i_10_503_316_0 & ~i_10_503_1445_0 & ~i_10_503_2353_0 & ~i_10_503_2711_0 & ~i_10_503_2881_0 & ~i_10_503_2985_0 & ~i_10_503_3848_0 & ~i_10_503_4124_0) | (~i_10_503_1005_0 & i_10_503_1648_0 & ~i_10_503_2357_0 & ~i_10_503_4123_0 & ~i_10_503_4278_0))))) | (~i_10_503_1445_0 & ((~i_10_503_290_0 & ((~i_10_503_283_0 & ((i_10_503_1819_0 & ~i_10_503_2029_0 & ~i_10_503_2729_0 & ~i_10_503_2922_0 & ~i_10_503_3384_0 & ~i_10_503_3610_0 & ~i_10_503_3848_0) | (~i_10_503_2408_0 & i_10_503_3610_0 & ~i_10_503_4270_0 & ~i_10_503_4271_0))) | (~i_10_503_316_0 & ~i_10_503_717_0 & ~i_10_503_1005_0 & ~i_10_503_1648_0 & ~i_10_503_2354_0 & ~i_10_503_2660_0 & ~i_10_503_2716_0 & ~i_10_503_3589_0 & ~i_10_503_3784_0 & ~i_10_503_3907_0 & ~i_10_503_4123_0 & ~i_10_503_3785_0 & ~i_10_503_3859_0))) | (~i_10_503_4025_0 & ~i_10_503_4292_0 & ((i_10_503_283_0 & ~i_10_503_1235_0 & ~i_10_503_2352_0 & ~i_10_503_2408_0 & ~i_10_503_2716_0 & ~i_10_503_2833_0 & ~i_10_503_4123_0) | (i_10_503_280_0 & ~i_10_503_316_0 & ~i_10_503_2354_0 & ~i_10_503_2711_0 & ~i_10_503_3387_0 & ~i_10_503_3388_0 & ~i_10_503_3907_0 & ~i_10_503_4269_0 & ~i_10_503_4270_0 & ~i_10_503_4278_0))))) | (i_10_503_1819_0 & ((i_10_503_439_0 & i_10_503_3858_0) | (~i_10_503_2027_0 & i_10_503_2628_0 & ~i_10_503_3044_0 & ~i_10_503_3409_0 & ~i_10_503_4292_0))) | (~i_10_503_4271_0 & ((i_10_503_3859_0 & ((~i_10_503_1915_0 & i_10_503_2354_0 & i_10_503_3388_0 & ~i_10_503_3840_0 & ~i_10_503_4270_0) | (i_10_503_3610_0 & ~i_10_503_4124_0 & ~i_10_503_4286_0))) | (~i_10_503_3044_0 & i_10_503_3199_0 & ~i_10_503_3589_0 & ~i_10_503_4278_0))) | (~i_10_503_2354_0 & i_10_503_3040_0 & ~i_10_503_3650_0));
endmodule



// Benchmark "kernel_10_504" written by ABC on Sun Jul 19 10:29:49 2020

module kernel_10_504 ( 
    i_10_504_175_0, i_10_504_176_0, i_10_504_186_0, i_10_504_187_0,
    i_10_504_188_0, i_10_504_282_0, i_10_504_409_0, i_10_504_464_0,
    i_10_504_467_0, i_10_504_516_0, i_10_504_1165_0, i_10_504_1169_0,
    i_10_504_1236_0, i_10_504_1249_0, i_10_504_1348_0, i_10_504_1435_0,
    i_10_504_1552_0, i_10_504_1556_0, i_10_504_1823_0, i_10_504_1824_0,
    i_10_504_1826_0, i_10_504_1947_0, i_10_504_1993_0, i_10_504_2021_0,
    i_10_504_2309_0, i_10_504_2350_0, i_10_504_2353_0, i_10_504_2450_0,
    i_10_504_2453_0, i_10_504_2467_0, i_10_504_2470_0, i_10_504_2514_0,
    i_10_504_2517_0, i_10_504_2571_0, i_10_504_2572_0, i_10_504_2633_0,
    i_10_504_2704_0, i_10_504_2708_0, i_10_504_2713_0, i_10_504_2714_0,
    i_10_504_2716_0, i_10_504_2717_0, i_10_504_2722_0, i_10_504_2727_0,
    i_10_504_2728_0, i_10_504_2823_0, i_10_504_2831_0, i_10_504_2870_0,
    i_10_504_2883_0, i_10_504_2884_0, i_10_504_2885_0, i_10_504_2886_0,
    i_10_504_2887_0, i_10_504_2921_0, i_10_504_2953_0, i_10_504_2981_0,
    i_10_504_3037_0, i_10_504_3038_0, i_10_504_3047_0, i_10_504_3074_0,
    i_10_504_3198_0, i_10_504_3271_0, i_10_504_3272_0, i_10_504_3274_0,
    i_10_504_3281_0, i_10_504_3386_0, i_10_504_3407_0, i_10_504_3434_0,
    i_10_504_3611_0, i_10_504_3614_0, i_10_504_3653_0, i_10_504_3720_0,
    i_10_504_3771_0, i_10_504_3783_0, i_10_504_3784_0, i_10_504_3785_0,
    i_10_504_3839_0, i_10_504_3853_0, i_10_504_3855_0, i_10_504_3856_0,
    i_10_504_3857_0, i_10_504_3880_0, i_10_504_3885_0, i_10_504_3886_0,
    i_10_504_3890_0, i_10_504_3895_0, i_10_504_3896_0, i_10_504_3984_0,
    i_10_504_3985_0, i_10_504_4051_0, i_10_504_4119_0, i_10_504_4120_0,
    i_10_504_4172_0, i_10_504_4175_0, i_10_504_4189_0, i_10_504_4190_0,
    i_10_504_4191_0, i_10_504_4291_0, i_10_504_4462_0, i_10_504_4571_0,
    o_10_504_0_0  );
  input  i_10_504_175_0, i_10_504_176_0, i_10_504_186_0, i_10_504_187_0,
    i_10_504_188_0, i_10_504_282_0, i_10_504_409_0, i_10_504_464_0,
    i_10_504_467_0, i_10_504_516_0, i_10_504_1165_0, i_10_504_1169_0,
    i_10_504_1236_0, i_10_504_1249_0, i_10_504_1348_0, i_10_504_1435_0,
    i_10_504_1552_0, i_10_504_1556_0, i_10_504_1823_0, i_10_504_1824_0,
    i_10_504_1826_0, i_10_504_1947_0, i_10_504_1993_0, i_10_504_2021_0,
    i_10_504_2309_0, i_10_504_2350_0, i_10_504_2353_0, i_10_504_2450_0,
    i_10_504_2453_0, i_10_504_2467_0, i_10_504_2470_0, i_10_504_2514_0,
    i_10_504_2517_0, i_10_504_2571_0, i_10_504_2572_0, i_10_504_2633_0,
    i_10_504_2704_0, i_10_504_2708_0, i_10_504_2713_0, i_10_504_2714_0,
    i_10_504_2716_0, i_10_504_2717_0, i_10_504_2722_0, i_10_504_2727_0,
    i_10_504_2728_0, i_10_504_2823_0, i_10_504_2831_0, i_10_504_2870_0,
    i_10_504_2883_0, i_10_504_2884_0, i_10_504_2885_0, i_10_504_2886_0,
    i_10_504_2887_0, i_10_504_2921_0, i_10_504_2953_0, i_10_504_2981_0,
    i_10_504_3037_0, i_10_504_3038_0, i_10_504_3047_0, i_10_504_3074_0,
    i_10_504_3198_0, i_10_504_3271_0, i_10_504_3272_0, i_10_504_3274_0,
    i_10_504_3281_0, i_10_504_3386_0, i_10_504_3407_0, i_10_504_3434_0,
    i_10_504_3611_0, i_10_504_3614_0, i_10_504_3653_0, i_10_504_3720_0,
    i_10_504_3771_0, i_10_504_3783_0, i_10_504_3784_0, i_10_504_3785_0,
    i_10_504_3839_0, i_10_504_3853_0, i_10_504_3855_0, i_10_504_3856_0,
    i_10_504_3857_0, i_10_504_3880_0, i_10_504_3885_0, i_10_504_3886_0,
    i_10_504_3890_0, i_10_504_3895_0, i_10_504_3896_0, i_10_504_3984_0,
    i_10_504_3985_0, i_10_504_4051_0, i_10_504_4119_0, i_10_504_4120_0,
    i_10_504_4172_0, i_10_504_4175_0, i_10_504_4189_0, i_10_504_4190_0,
    i_10_504_4191_0, i_10_504_4291_0, i_10_504_4462_0, i_10_504_4571_0;
  output o_10_504_0_0;
  assign o_10_504_0_0 = 0;
endmodule



// Benchmark "kernel_10_505" written by ABC on Sun Jul 19 10:29:50 2020

module kernel_10_505 ( 
    i_10_505_178_0, i_10_505_254_0, i_10_505_260_0, i_10_505_266_0,
    i_10_505_277_0, i_10_505_280_0, i_10_505_283_0, i_10_505_287_0,
    i_10_505_319_0, i_10_505_407_0, i_10_505_442_0, i_10_505_497_0,
    i_10_505_503_0, i_10_505_506_0, i_10_505_509_0, i_10_505_512_0,
    i_10_505_866_0, i_10_505_869_0, i_10_505_1007_0, i_10_505_1083_0,
    i_10_505_1085_0, i_10_505_1086_0, i_10_505_1102_0, i_10_505_1237_0,
    i_10_505_1238_0, i_10_505_1250_0, i_10_505_1297_0, i_10_505_1301_0,
    i_10_505_1303_0, i_10_505_1307_0, i_10_505_1540_0, i_10_505_1541_0,
    i_10_505_1621_0, i_10_505_1622_0, i_10_505_1626_0, i_10_505_1686_0,
    i_10_505_1687_0, i_10_505_1688_0, i_10_505_1764_0, i_10_505_1798_0,
    i_10_505_1807_0, i_10_505_1984_0, i_10_505_2027_0, i_10_505_2030_0,
    i_10_505_2032_0, i_10_505_2033_0, i_10_505_2091_0, i_10_505_2110_0,
    i_10_505_2182_0, i_10_505_2203_0, i_10_505_2354_0, i_10_505_2456_0,
    i_10_505_2471_0, i_10_505_2516_0, i_10_505_2656_0, i_10_505_2701_0,
    i_10_505_2702_0, i_10_505_2703_0, i_10_505_2722_0, i_10_505_2728_0,
    i_10_505_2729_0, i_10_505_2731_0, i_10_505_2734_0, i_10_505_2735_0,
    i_10_505_2965_0, i_10_505_2968_0, i_10_505_2969_0, i_10_505_2984_0,
    i_10_505_3046_0, i_10_505_3314_0, i_10_505_3317_0, i_10_505_3391_0,
    i_10_505_3392_0, i_10_505_3409_0, i_10_505_3410_0, i_10_505_3467_0,
    i_10_505_3470_0, i_10_505_3494_0, i_10_505_3506_0, i_10_505_3525_0,
    i_10_505_3538_0, i_10_505_3587_0, i_10_505_3682_0, i_10_505_3837_0,
    i_10_505_3840_0, i_10_505_3844_0, i_10_505_3850_0, i_10_505_3895_0,
    i_10_505_3982_0, i_10_505_4114_0, i_10_505_4188_0, i_10_505_4208_0,
    i_10_505_4268_0, i_10_505_4271_0, i_10_505_4274_0, i_10_505_4283_0,
    i_10_505_4285_0, i_10_505_4288_0, i_10_505_4292_0, i_10_505_4569_0,
    o_10_505_0_0  );
  input  i_10_505_178_0, i_10_505_254_0, i_10_505_260_0, i_10_505_266_0,
    i_10_505_277_0, i_10_505_280_0, i_10_505_283_0, i_10_505_287_0,
    i_10_505_319_0, i_10_505_407_0, i_10_505_442_0, i_10_505_497_0,
    i_10_505_503_0, i_10_505_506_0, i_10_505_509_0, i_10_505_512_0,
    i_10_505_866_0, i_10_505_869_0, i_10_505_1007_0, i_10_505_1083_0,
    i_10_505_1085_0, i_10_505_1086_0, i_10_505_1102_0, i_10_505_1237_0,
    i_10_505_1238_0, i_10_505_1250_0, i_10_505_1297_0, i_10_505_1301_0,
    i_10_505_1303_0, i_10_505_1307_0, i_10_505_1540_0, i_10_505_1541_0,
    i_10_505_1621_0, i_10_505_1622_0, i_10_505_1626_0, i_10_505_1686_0,
    i_10_505_1687_0, i_10_505_1688_0, i_10_505_1764_0, i_10_505_1798_0,
    i_10_505_1807_0, i_10_505_1984_0, i_10_505_2027_0, i_10_505_2030_0,
    i_10_505_2032_0, i_10_505_2033_0, i_10_505_2091_0, i_10_505_2110_0,
    i_10_505_2182_0, i_10_505_2203_0, i_10_505_2354_0, i_10_505_2456_0,
    i_10_505_2471_0, i_10_505_2516_0, i_10_505_2656_0, i_10_505_2701_0,
    i_10_505_2702_0, i_10_505_2703_0, i_10_505_2722_0, i_10_505_2728_0,
    i_10_505_2729_0, i_10_505_2731_0, i_10_505_2734_0, i_10_505_2735_0,
    i_10_505_2965_0, i_10_505_2968_0, i_10_505_2969_0, i_10_505_2984_0,
    i_10_505_3046_0, i_10_505_3314_0, i_10_505_3317_0, i_10_505_3391_0,
    i_10_505_3392_0, i_10_505_3409_0, i_10_505_3410_0, i_10_505_3467_0,
    i_10_505_3470_0, i_10_505_3494_0, i_10_505_3506_0, i_10_505_3525_0,
    i_10_505_3538_0, i_10_505_3587_0, i_10_505_3682_0, i_10_505_3837_0,
    i_10_505_3840_0, i_10_505_3844_0, i_10_505_3850_0, i_10_505_3895_0,
    i_10_505_3982_0, i_10_505_4114_0, i_10_505_4188_0, i_10_505_4208_0,
    i_10_505_4268_0, i_10_505_4271_0, i_10_505_4274_0, i_10_505_4283_0,
    i_10_505_4285_0, i_10_505_4288_0, i_10_505_4292_0, i_10_505_4569_0;
  output o_10_505_0_0;
  assign o_10_505_0_0 = ~((~i_10_505_3844_0 & ((~i_10_505_266_0 & ((~i_10_505_1007_0 & ~i_10_505_2027_0 & ~i_10_505_2703_0 & ~i_10_505_2731_0 & ~i_10_505_2735_0 & ~i_10_505_3467_0) | (~i_10_505_319_0 & ~i_10_505_1540_0 & ~i_10_505_2032_0 & ~i_10_505_2456_0 & ~i_10_505_2701_0 & ~i_10_505_3506_0 & ~i_10_505_3538_0 & ~i_10_505_4283_0 & ~i_10_505_4569_0))) | (~i_10_505_2729_0 & ~i_10_505_3470_0 & ~i_10_505_4292_0))) | (~i_10_505_1085_0 & ((~i_10_505_1250_0 & i_10_505_2729_0 & ~i_10_505_3317_0 & ~i_10_505_3392_0 & ~i_10_505_3410_0 & ~i_10_505_3467_0) | (~i_10_505_283_0 & ~i_10_505_1621_0 & ~i_10_505_2027_0 & ~i_10_505_2033_0 & ~i_10_505_3494_0 & ~i_10_505_3506_0 & ~i_10_505_3525_0 & ~i_10_505_4283_0))) | (~i_10_505_283_0 & ((~i_10_505_1237_0 & ~i_10_505_1238_0 & ~i_10_505_1250_0 & i_10_505_2456_0 & ~i_10_505_2728_0) | (~i_10_505_407_0 & ~i_10_505_1622_0 & ~i_10_505_2033_0 & ~i_10_505_2354_0 & ~i_10_505_3467_0 & ~i_10_505_4268_0))) | (~i_10_505_3392_0 & ((~i_10_505_1250_0 & ((~i_10_505_1687_0 & ~i_10_505_2728_0) | (~i_10_505_2656_0 & i_10_505_2731_0 & ~i_10_505_3317_0 & ~i_10_505_3506_0 & ~i_10_505_4271_0 & ~i_10_505_4292_0))) | (i_10_505_1307_0 & ~i_10_505_2722_0 & ~i_10_505_3467_0 & ~i_10_505_3506_0 & ~i_10_505_3895_0 & ~i_10_505_4288_0))) | (~i_10_505_2027_0 & ((~i_10_505_319_0 & ~i_10_505_2471_0 & ~i_10_505_2702_0 & ~i_10_505_4271_0) | (~i_10_505_178_0 & ~i_10_505_1688_0 & ~i_10_505_4292_0))) | (~i_10_505_2033_0 & ((~i_10_505_1622_0 & ~i_10_505_2729_0 & ~i_10_505_3314_0 & ~i_10_505_3494_0 & ~i_10_505_4274_0) | (~i_10_505_280_0 & ~i_10_505_1083_0 & ~i_10_505_2030_0 & ~i_10_505_2702_0 & ~i_10_505_4114_0 & i_10_505_4288_0))) | (~i_10_505_1237_0 & ~i_10_505_1238_0 & i_10_505_2735_0 & ~i_10_505_3467_0 & ~i_10_505_4274_0));
endmodule



// Benchmark "kernel_10_506" written by ABC on Sun Jul 19 10:29:51 2020

module kernel_10_506 ( 
    i_10_506_67_0, i_10_506_147_0, i_10_506_151_0, i_10_506_175_0,
    i_10_506_190_0, i_10_506_220_0, i_10_506_318_0, i_10_506_319_0,
    i_10_506_364_0, i_10_506_372_0, i_10_506_410_0, i_10_506_475_0,
    i_10_506_595_0, i_10_506_690_0, i_10_506_733_0, i_10_506_876_0,
    i_10_506_1000_0, i_10_506_1011_0, i_10_506_1069_0, i_10_506_1083_0,
    i_10_506_1099_0, i_10_506_1110_0, i_10_506_1278_0, i_10_506_1293_0,
    i_10_506_1308_0, i_10_506_1309_0, i_10_506_1443_0, i_10_506_1596_0,
    i_10_506_1619_0, i_10_506_1621_0, i_10_506_1623_0, i_10_506_1624_0,
    i_10_506_1635_0, i_10_506_1636_0, i_10_506_1647_0, i_10_506_1651_0,
    i_10_506_1818_0, i_10_506_1821_0, i_10_506_1822_0, i_10_506_1849_0,
    i_10_506_1918_0, i_10_506_1956_0, i_10_506_1959_0, i_10_506_1965_0,
    i_10_506_1987_0, i_10_506_2109_0, i_10_506_2112_0, i_10_506_2226_0,
    i_10_506_2305_0, i_10_506_2353_0, i_10_506_2481_0, i_10_506_2482_0,
    i_10_506_2516_0, i_10_506_2540_0, i_10_506_2561_0, i_10_506_2569_0,
    i_10_506_2588_0, i_10_506_2659_0, i_10_506_2677_0, i_10_506_2680_0,
    i_10_506_2686_0, i_10_506_2713_0, i_10_506_2778_0, i_10_506_2785_0,
    i_10_506_2884_0, i_10_506_2952_0, i_10_506_2953_0, i_10_506_2956_0,
    i_10_506_2980_0, i_10_506_2990_0, i_10_506_3040_0, i_10_506_3276_0,
    i_10_506_3283_0, i_10_506_3297_0, i_10_506_3324_0, i_10_506_3325_0,
    i_10_506_3450_0, i_10_506_3454_0, i_10_506_3550_0, i_10_506_3585_0,
    i_10_506_3649_0, i_10_506_3704_0, i_10_506_3779_0, i_10_506_3838_0,
    i_10_506_3853_0, i_10_506_3854_0, i_10_506_3896_0, i_10_506_4028_0,
    i_10_506_4057_0, i_10_506_4118_0, i_10_506_4120_0, i_10_506_4168_0,
    i_10_506_4279_0, i_10_506_4317_0, i_10_506_4380_0, i_10_506_4459_0,
    i_10_506_4546_0, i_10_506_4570_0, i_10_506_4582_0, i_10_506_4585_0,
    o_10_506_0_0  );
  input  i_10_506_67_0, i_10_506_147_0, i_10_506_151_0, i_10_506_175_0,
    i_10_506_190_0, i_10_506_220_0, i_10_506_318_0, i_10_506_319_0,
    i_10_506_364_0, i_10_506_372_0, i_10_506_410_0, i_10_506_475_0,
    i_10_506_595_0, i_10_506_690_0, i_10_506_733_0, i_10_506_876_0,
    i_10_506_1000_0, i_10_506_1011_0, i_10_506_1069_0, i_10_506_1083_0,
    i_10_506_1099_0, i_10_506_1110_0, i_10_506_1278_0, i_10_506_1293_0,
    i_10_506_1308_0, i_10_506_1309_0, i_10_506_1443_0, i_10_506_1596_0,
    i_10_506_1619_0, i_10_506_1621_0, i_10_506_1623_0, i_10_506_1624_0,
    i_10_506_1635_0, i_10_506_1636_0, i_10_506_1647_0, i_10_506_1651_0,
    i_10_506_1818_0, i_10_506_1821_0, i_10_506_1822_0, i_10_506_1849_0,
    i_10_506_1918_0, i_10_506_1956_0, i_10_506_1959_0, i_10_506_1965_0,
    i_10_506_1987_0, i_10_506_2109_0, i_10_506_2112_0, i_10_506_2226_0,
    i_10_506_2305_0, i_10_506_2353_0, i_10_506_2481_0, i_10_506_2482_0,
    i_10_506_2516_0, i_10_506_2540_0, i_10_506_2561_0, i_10_506_2569_0,
    i_10_506_2588_0, i_10_506_2659_0, i_10_506_2677_0, i_10_506_2680_0,
    i_10_506_2686_0, i_10_506_2713_0, i_10_506_2778_0, i_10_506_2785_0,
    i_10_506_2884_0, i_10_506_2952_0, i_10_506_2953_0, i_10_506_2956_0,
    i_10_506_2980_0, i_10_506_2990_0, i_10_506_3040_0, i_10_506_3276_0,
    i_10_506_3283_0, i_10_506_3297_0, i_10_506_3324_0, i_10_506_3325_0,
    i_10_506_3450_0, i_10_506_3454_0, i_10_506_3550_0, i_10_506_3585_0,
    i_10_506_3649_0, i_10_506_3704_0, i_10_506_3779_0, i_10_506_3838_0,
    i_10_506_3853_0, i_10_506_3854_0, i_10_506_3896_0, i_10_506_4028_0,
    i_10_506_4057_0, i_10_506_4118_0, i_10_506_4120_0, i_10_506_4168_0,
    i_10_506_4279_0, i_10_506_4317_0, i_10_506_4380_0, i_10_506_4459_0,
    i_10_506_4546_0, i_10_506_4570_0, i_10_506_4582_0, i_10_506_4585_0;
  output o_10_506_0_0;
  assign o_10_506_0_0 = 0;
endmodule



// Benchmark "kernel_10_507" written by ABC on Sun Jul 19 10:29:52 2020

module kernel_10_507 ( 
    i_10_507_35_0, i_10_507_118_0, i_10_507_119_0, i_10_507_124_0,
    i_10_507_125_0, i_10_507_175_0, i_10_507_268_0, i_10_507_284_0,
    i_10_507_368_0, i_10_507_391_0, i_10_507_440_0, i_10_507_461_0,
    i_10_507_464_0, i_10_507_521_0, i_10_507_566_0, i_10_507_588_0,
    i_10_507_589_0, i_10_507_590_0, i_10_507_831_0, i_10_507_832_0,
    i_10_507_833_0, i_10_507_899_0, i_10_507_962_0, i_10_507_963_0,
    i_10_507_997_0, i_10_507_1007_0, i_10_507_1055_0, i_10_507_1166_0,
    i_10_507_1310_0, i_10_507_1348_0, i_10_507_1367_0, i_10_507_1382_0,
    i_10_507_1435_0, i_10_507_1436_0, i_10_507_1438_0, i_10_507_1439_0,
    i_10_507_1456_0, i_10_507_1457_0, i_10_507_1616_0, i_10_507_1618_0,
    i_10_507_1619_0, i_10_507_1636_0, i_10_507_1689_0, i_10_507_1822_0,
    i_10_507_1823_0, i_10_507_1922_0, i_10_507_1948_0, i_10_507_1952_0,
    i_10_507_1986_0, i_10_507_2006_0, i_10_507_2213_0, i_10_507_2244_0,
    i_10_507_2356_0, i_10_507_2408_0, i_10_507_2409_0, i_10_507_2430_0,
    i_10_507_2454_0, i_10_507_2515_0, i_10_507_2516_0, i_10_507_2617_0,
    i_10_507_2618_0, i_10_507_2628_0, i_10_507_2629_0, i_10_507_2633_0,
    i_10_507_2660_0, i_10_507_2681_0, i_10_507_2713_0, i_10_507_2731_0,
    i_10_507_2732_0, i_10_507_2882_0, i_10_507_2920_0, i_10_507_2924_0,
    i_10_507_3040_0, i_10_507_3041_0, i_10_507_3043_0, i_10_507_3094_0,
    i_10_507_3117_0, i_10_507_3122_0, i_10_507_3200_0, i_10_507_3351_0,
    i_10_507_3391_0, i_10_507_3526_0, i_10_507_3542_0, i_10_507_3580_0,
    i_10_507_3587_0, i_10_507_3610_0, i_10_507_3613_0, i_10_507_3625_0,
    i_10_507_3647_0, i_10_507_3649_0, i_10_507_3652_0, i_10_507_3653_0,
    i_10_507_3783_0, i_10_507_3837_0, i_10_507_3838_0, i_10_507_3895_0,
    i_10_507_3985_0, i_10_507_4001_0, i_10_507_4172_0, i_10_507_4373_0,
    o_10_507_0_0  );
  input  i_10_507_35_0, i_10_507_118_0, i_10_507_119_0, i_10_507_124_0,
    i_10_507_125_0, i_10_507_175_0, i_10_507_268_0, i_10_507_284_0,
    i_10_507_368_0, i_10_507_391_0, i_10_507_440_0, i_10_507_461_0,
    i_10_507_464_0, i_10_507_521_0, i_10_507_566_0, i_10_507_588_0,
    i_10_507_589_0, i_10_507_590_0, i_10_507_831_0, i_10_507_832_0,
    i_10_507_833_0, i_10_507_899_0, i_10_507_962_0, i_10_507_963_0,
    i_10_507_997_0, i_10_507_1007_0, i_10_507_1055_0, i_10_507_1166_0,
    i_10_507_1310_0, i_10_507_1348_0, i_10_507_1367_0, i_10_507_1382_0,
    i_10_507_1435_0, i_10_507_1436_0, i_10_507_1438_0, i_10_507_1439_0,
    i_10_507_1456_0, i_10_507_1457_0, i_10_507_1616_0, i_10_507_1618_0,
    i_10_507_1619_0, i_10_507_1636_0, i_10_507_1689_0, i_10_507_1822_0,
    i_10_507_1823_0, i_10_507_1922_0, i_10_507_1948_0, i_10_507_1952_0,
    i_10_507_1986_0, i_10_507_2006_0, i_10_507_2213_0, i_10_507_2244_0,
    i_10_507_2356_0, i_10_507_2408_0, i_10_507_2409_0, i_10_507_2430_0,
    i_10_507_2454_0, i_10_507_2515_0, i_10_507_2516_0, i_10_507_2617_0,
    i_10_507_2618_0, i_10_507_2628_0, i_10_507_2629_0, i_10_507_2633_0,
    i_10_507_2660_0, i_10_507_2681_0, i_10_507_2713_0, i_10_507_2731_0,
    i_10_507_2732_0, i_10_507_2882_0, i_10_507_2920_0, i_10_507_2924_0,
    i_10_507_3040_0, i_10_507_3041_0, i_10_507_3043_0, i_10_507_3094_0,
    i_10_507_3117_0, i_10_507_3122_0, i_10_507_3200_0, i_10_507_3351_0,
    i_10_507_3391_0, i_10_507_3526_0, i_10_507_3542_0, i_10_507_3580_0,
    i_10_507_3587_0, i_10_507_3610_0, i_10_507_3613_0, i_10_507_3625_0,
    i_10_507_3647_0, i_10_507_3649_0, i_10_507_3652_0, i_10_507_3653_0,
    i_10_507_3783_0, i_10_507_3837_0, i_10_507_3838_0, i_10_507_3895_0,
    i_10_507_3985_0, i_10_507_4001_0, i_10_507_4172_0, i_10_507_4373_0;
  output o_10_507_0_0;
  assign o_10_507_0_0 = 0;
endmodule



// Benchmark "kernel_10_508" written by ABC on Sun Jul 19 10:29:54 2020

module kernel_10_508 ( 
    i_10_508_171_0, i_10_508_174_0, i_10_508_179_0, i_10_508_221_0,
    i_10_508_245_0, i_10_508_280_0, i_10_508_433_0, i_10_508_435_0,
    i_10_508_436_0, i_10_508_437_0, i_10_508_439_0, i_10_508_440_0,
    i_10_508_444_0, i_10_508_749_0, i_10_508_797_0, i_10_508_1001_0,
    i_10_508_1005_0, i_10_508_1166_0, i_10_508_1234_0, i_10_508_1235_0,
    i_10_508_1246_0, i_10_508_1249_0, i_10_508_1250_0, i_10_508_1309_0,
    i_10_508_1310_0, i_10_508_1550_0, i_10_508_1649_0, i_10_508_1652_0,
    i_10_508_1684_0, i_10_508_1686_0, i_10_508_1687_0, i_10_508_1819_0,
    i_10_508_1822_0, i_10_508_1823_0, i_10_508_1825_0, i_10_508_1946_0,
    i_10_508_2179_0, i_10_508_2180_0, i_10_508_2306_0, i_10_508_2357_0,
    i_10_508_2365_0, i_10_508_2384_0, i_10_508_2470_0, i_10_508_2471_0,
    i_10_508_2516_0, i_10_508_2629_0, i_10_508_2631_0, i_10_508_2633_0,
    i_10_508_2659_0, i_10_508_2675_0, i_10_508_2708_0, i_10_508_2723_0,
    i_10_508_2727_0, i_10_508_2731_0, i_10_508_2830_0, i_10_508_2884_0,
    i_10_508_2885_0, i_10_508_2887_0, i_10_508_2917_0, i_10_508_2918_0,
    i_10_508_3150_0, i_10_508_3151_0, i_10_508_3152_0, i_10_508_3200_0,
    i_10_508_3238_0, i_10_508_3268_0, i_10_508_3269_0, i_10_508_3274_0,
    i_10_508_3322_0, i_10_508_3390_0, i_10_508_3391_0, i_10_508_3406_0,
    i_10_508_3407_0, i_10_508_3410_0, i_10_508_3470_0, i_10_508_3590_0,
    i_10_508_3610_0, i_10_508_3613_0, i_10_508_3614_0, i_10_508_3784_0,
    i_10_508_3835_0, i_10_508_3837_0, i_10_508_3838_0, i_10_508_3839_0,
    i_10_508_3841_0, i_10_508_3846_0, i_10_508_3847_0, i_10_508_3848_0,
    i_10_508_3849_0, i_10_508_3850_0, i_10_508_3853_0, i_10_508_3855_0,
    i_10_508_3859_0, i_10_508_3979_0, i_10_508_3986_0, i_10_508_4117_0,
    i_10_508_4123_0, i_10_508_4285_0, i_10_508_4287_0, i_10_508_4567_0,
    o_10_508_0_0  );
  input  i_10_508_171_0, i_10_508_174_0, i_10_508_179_0, i_10_508_221_0,
    i_10_508_245_0, i_10_508_280_0, i_10_508_433_0, i_10_508_435_0,
    i_10_508_436_0, i_10_508_437_0, i_10_508_439_0, i_10_508_440_0,
    i_10_508_444_0, i_10_508_749_0, i_10_508_797_0, i_10_508_1001_0,
    i_10_508_1005_0, i_10_508_1166_0, i_10_508_1234_0, i_10_508_1235_0,
    i_10_508_1246_0, i_10_508_1249_0, i_10_508_1250_0, i_10_508_1309_0,
    i_10_508_1310_0, i_10_508_1550_0, i_10_508_1649_0, i_10_508_1652_0,
    i_10_508_1684_0, i_10_508_1686_0, i_10_508_1687_0, i_10_508_1819_0,
    i_10_508_1822_0, i_10_508_1823_0, i_10_508_1825_0, i_10_508_1946_0,
    i_10_508_2179_0, i_10_508_2180_0, i_10_508_2306_0, i_10_508_2357_0,
    i_10_508_2365_0, i_10_508_2384_0, i_10_508_2470_0, i_10_508_2471_0,
    i_10_508_2516_0, i_10_508_2629_0, i_10_508_2631_0, i_10_508_2633_0,
    i_10_508_2659_0, i_10_508_2675_0, i_10_508_2708_0, i_10_508_2723_0,
    i_10_508_2727_0, i_10_508_2731_0, i_10_508_2830_0, i_10_508_2884_0,
    i_10_508_2885_0, i_10_508_2887_0, i_10_508_2917_0, i_10_508_2918_0,
    i_10_508_3150_0, i_10_508_3151_0, i_10_508_3152_0, i_10_508_3200_0,
    i_10_508_3238_0, i_10_508_3268_0, i_10_508_3269_0, i_10_508_3274_0,
    i_10_508_3322_0, i_10_508_3390_0, i_10_508_3391_0, i_10_508_3406_0,
    i_10_508_3407_0, i_10_508_3410_0, i_10_508_3470_0, i_10_508_3590_0,
    i_10_508_3610_0, i_10_508_3613_0, i_10_508_3614_0, i_10_508_3784_0,
    i_10_508_3835_0, i_10_508_3837_0, i_10_508_3838_0, i_10_508_3839_0,
    i_10_508_3841_0, i_10_508_3846_0, i_10_508_3847_0, i_10_508_3848_0,
    i_10_508_3849_0, i_10_508_3850_0, i_10_508_3853_0, i_10_508_3855_0,
    i_10_508_3859_0, i_10_508_3979_0, i_10_508_3986_0, i_10_508_4117_0,
    i_10_508_4123_0, i_10_508_4285_0, i_10_508_4287_0, i_10_508_4567_0;
  output o_10_508_0_0;
  assign o_10_508_0_0 = ~((~i_10_508_171_0 & i_10_508_1819_0 & ((~i_10_508_2306_0 & ~i_10_508_2659_0 & ~i_10_508_2675_0 & ~i_10_508_3390_0 & ~i_10_508_3406_0 & ~i_10_508_3410_0 & ~i_10_508_3614_0 & ~i_10_508_3979_0) | (~i_10_508_444_0 & ~i_10_508_749_0 & ~i_10_508_1823_0 & ~i_10_508_2180_0 & i_10_508_3853_0 & ~i_10_508_3986_0))) | (~i_10_508_174_0 & ((~i_10_508_221_0 & ~i_10_508_436_0 & ~i_10_508_1310_0 & ~i_10_508_1550_0 & ~i_10_508_1825_0 & ~i_10_508_2723_0 & ~i_10_508_3784_0 & i_10_508_4117_0) | (~i_10_508_1005_0 & ~i_10_508_1246_0 & i_10_508_1822_0 & i_10_508_1825_0 & ~i_10_508_1946_0 & ~i_10_508_2885_0 & ~i_10_508_3406_0 & ~i_10_508_3590_0 & ~i_10_508_3610_0 & ~i_10_508_3839_0 & ~i_10_508_4285_0))) | (~i_10_508_3406_0 & ((~i_10_508_221_0 & ((~i_10_508_245_0 & ~i_10_508_1005_0 & ~i_10_508_1309_0 & ~i_10_508_1310_0 & ~i_10_508_2179_0 & ~i_10_508_2659_0 & ~i_10_508_2884_0 & ~i_10_508_3274_0 & i_10_508_3838_0) | (~i_10_508_1649_0 & ~i_10_508_2306_0 & ~i_10_508_2723_0 & ~i_10_508_3839_0 & i_10_508_3847_0))) | (~i_10_508_1684_0 & ~i_10_508_3986_0 & ((~i_10_508_437_0 & ~i_10_508_439_0 & ~i_10_508_440_0 & ~i_10_508_1822_0 & i_10_508_1825_0 & ~i_10_508_2884_0 & ~i_10_508_3269_0) | (~i_10_508_1235_0 & ~i_10_508_1825_0 & ~i_10_508_2629_0 & ~i_10_508_2659_0 & ~i_10_508_2885_0 & ~i_10_508_2887_0 & ~i_10_508_3837_0))))) | (~i_10_508_433_0 & ((i_10_508_1825_0 & i_10_508_2731_0 & ~i_10_508_3614_0 & ~i_10_508_3837_0) | (~i_10_508_1234_0 & ~i_10_508_1309_0 & ~i_10_508_1310_0 & ~i_10_508_1946_0 & ~i_10_508_3269_0 & ~i_10_508_3410_0 & ~i_10_508_3838_0 & ~i_10_508_3979_0 & ~i_10_508_4123_0))) | (~i_10_508_3841_0 & ((~i_10_508_436_0 & ~i_10_508_2629_0 & ((i_10_508_1822_0 & ~i_10_508_3200_0 & ~i_10_508_3614_0 & i_10_508_3835_0) | (~i_10_508_439_0 & ~i_10_508_440_0 & ~i_10_508_1005_0 & ~i_10_508_1823_0 & ~i_10_508_1825_0 & ~i_10_508_2384_0 & ~i_10_508_2675_0 & ~i_10_508_3784_0 & ~i_10_508_4287_0))) | (~i_10_508_440_0 & ~i_10_508_1005_0 & ~i_10_508_1649_0 & ~i_10_508_1686_0 & ~i_10_508_2179_0 & ~i_10_508_2180_0 & ~i_10_508_2306_0 & ~i_10_508_2384_0 & ~i_10_508_2884_0 & ~i_10_508_2885_0 & ~i_10_508_3269_0 & ~i_10_508_3391_0 & ~i_10_508_3407_0 & ~i_10_508_3590_0 & ~i_10_508_3979_0 & ~i_10_508_4117_0))) | (~i_10_508_439_0 & ((i_10_508_3835_0 & ~i_10_508_3838_0 & i_10_508_4285_0) | (~i_10_508_1310_0 & ~i_10_508_1822_0 & i_10_508_2629_0 & ~i_10_508_3614_0 & ~i_10_508_3853_0 & ~i_10_508_3859_0 & ~i_10_508_4567_0))) | (~i_10_508_2884_0 & ((~i_10_508_2179_0 & ((~i_10_508_245_0 & ((~i_10_508_1001_0 & ~i_10_508_1823_0 & ~i_10_508_3200_0 & i_10_508_3590_0 & ~i_10_508_3784_0) | (~i_10_508_2180_0 & i_10_508_2918_0 & ~i_10_508_3979_0 & ~i_10_508_3986_0))) | (~i_10_508_1005_0 & ~i_10_508_1310_0 & ~i_10_508_2306_0 & ((i_10_508_1652_0 & ~i_10_508_1822_0 & ~i_10_508_2180_0 & ~i_10_508_2830_0 & ~i_10_508_3407_0) | (~i_10_508_444_0 & ~i_10_508_1550_0 & ~i_10_508_1686_0 & ~i_10_508_3614_0))) | (i_10_508_1249_0 & ~i_10_508_1649_0 & ~i_10_508_3274_0 & i_10_508_3855_0 & ~i_10_508_4287_0))) | (~i_10_508_1309_0 & ~i_10_508_1686_0 & ~i_10_508_1946_0 & ~i_10_508_2180_0 & ~i_10_508_2306_0 & ~i_10_508_2675_0 & ~i_10_508_3407_0 & ~i_10_508_3784_0 & ~i_10_508_3979_0 & ~i_10_508_3986_0) | (~i_10_508_797_0 & ~i_10_508_1001_0 & ~i_10_508_1652_0 & ~i_10_508_1825_0 & ~i_10_508_2365_0 & ~i_10_508_2631_0 & ~i_10_508_2727_0 & ~i_10_508_2885_0 & ~i_10_508_2887_0 & ~i_10_508_3590_0 & ~i_10_508_3610_0 & ~i_10_508_3855_0))) | (~i_10_508_1822_0 & ((~i_10_508_797_0 & ((i_10_508_433_0 & ~i_10_508_1652_0 & ~i_10_508_1946_0 & ~i_10_508_3838_0 & i_10_508_3853_0) | (~i_10_508_437_0 & ~i_10_508_2306_0 & ~i_10_508_2727_0 & ~i_10_508_3269_0 & i_10_508_3610_0 & ~i_10_508_3784_0 & ~i_10_508_3979_0))) | (~i_10_508_749_0 & ~i_10_508_1686_0 & ~i_10_508_2384_0 & ~i_10_508_2675_0 & i_10_508_2731_0 & ~i_10_508_3200_0 & ~i_10_508_3986_0))) | (~i_10_508_437_0 & ((~i_10_508_1310_0 & i_10_508_2917_0 & ~i_10_508_2918_0) | (i_10_508_280_0 & i_10_508_435_0 & ~i_10_508_2675_0 & i_10_508_3853_0))) | (~i_10_508_3613_0 & ((~i_10_508_245_0 & ~i_10_508_1946_0 & ((~i_10_508_1825_0 & i_10_508_2731_0 & ~i_10_508_3839_0 & ~i_10_508_3979_0) | (~i_10_508_1005_0 & ~i_10_508_1309_0 & ~i_10_508_2179_0 & ~i_10_508_2885_0 & ~i_10_508_2918_0 & ~i_10_508_3614_0 & ~i_10_508_3850_0 & ~i_10_508_3986_0))) | (~i_10_508_440_0 & ~i_10_508_1005_0 & ~i_10_508_1649_0 & ~i_10_508_1823_0 & ~i_10_508_2179_0 & ~i_10_508_2180_0 & ~i_10_508_2357_0 & ~i_10_508_2887_0) | (~i_10_508_1309_0 & i_10_508_1825_0 & ~i_10_508_3268_0 & i_10_508_3850_0))) | (~i_10_508_3979_0 & ((~i_10_508_2306_0 & ((~i_10_508_245_0 & ~i_10_508_1235_0 & ~i_10_508_1310_0 & i_10_508_1687_0 & ~i_10_508_2384_0 & i_10_508_2731_0) | (~i_10_508_1005_0 & ~i_10_508_1649_0 & ~i_10_508_2180_0 & ~i_10_508_2887_0 & ~i_10_508_3614_0 & ~i_10_508_3837_0 & ~i_10_508_3838_0))) | (i_10_508_2633_0 & ~i_10_508_2675_0 & ~i_10_508_3839_0 & i_10_508_3859_0 & ~i_10_508_4117_0))) | (i_10_508_1250_0 & ~i_10_508_1686_0 & ~i_10_508_2885_0 & i_10_508_3274_0 & ~i_10_508_3855_0) | (i_10_508_3859_0 & ~i_10_508_4117_0 & i_10_508_2365_0 & ~i_10_508_3839_0));
endmodule



// Benchmark "kernel_10_509" written by ABC on Sun Jul 19 10:29:55 2020

module kernel_10_509 ( 
    i_10_509_34_0, i_10_509_150_0, i_10_509_172_0, i_10_509_174_0,
    i_10_509_175_0, i_10_509_435_0, i_10_509_438_0, i_10_509_444_0,
    i_10_509_447_0, i_10_509_448_0, i_10_509_462_0, i_10_509_467_0,
    i_10_509_508_0, i_10_509_516_0, i_10_509_519_0, i_10_509_717_0,
    i_10_509_799_0, i_10_509_966_0, i_10_509_967_0, i_10_509_996_0,
    i_10_509_1029_0, i_10_509_1141_0, i_10_509_1164_0, i_10_509_1240_0,
    i_10_509_1245_0, i_10_509_1248_0, i_10_509_1309_0, i_10_509_1311_0,
    i_10_509_1366_0, i_10_509_1626_0, i_10_509_1652_0, i_10_509_1653_0,
    i_10_509_1655_0, i_10_509_1689_0, i_10_509_1690_0, i_10_509_1797_0,
    i_10_509_1821_0, i_10_509_1822_0, i_10_509_1912_0, i_10_509_1995_0,
    i_10_509_2005_0, i_10_509_2352_0, i_10_509_2353_0, i_10_509_2455_0,
    i_10_509_2469_0, i_10_509_2472_0, i_10_509_2473_0, i_10_509_2571_0,
    i_10_509_2628_0, i_10_509_2629_0, i_10_509_2659_0, i_10_509_2661_0,
    i_10_509_2706_0, i_10_509_2715_0, i_10_509_2716_0, i_10_509_2722_0,
    i_10_509_2731_0, i_10_509_2734_0, i_10_509_2742_0, i_10_509_2782_0,
    i_10_509_2830_0, i_10_509_2832_0, i_10_509_2883_0, i_10_509_2987_0,
    i_10_509_3037_0, i_10_509_3039_0, i_10_509_3046_0, i_10_509_3048_0,
    i_10_509_3075_0, i_10_509_3093_0, i_10_509_3157_0, i_10_509_3197_0,
    i_10_509_3284_0, i_10_509_3321_0, i_10_509_3322_0, i_10_509_3327_0,
    i_10_509_3391_0, i_10_509_3392_0, i_10_509_3468_0, i_10_509_3495_0,
    i_10_509_3525_0, i_10_509_3583_0, i_10_509_3585_0, i_10_509_3612_0,
    i_10_509_3613_0, i_10_509_3732_0, i_10_509_3780_0, i_10_509_3837_0,
    i_10_509_3876_0, i_10_509_3912_0, i_10_509_3982_0, i_10_509_4113_0,
    i_10_509_4173_0, i_10_509_4269_0, i_10_509_4272_0, i_10_509_4273_0,
    i_10_509_4282_0, i_10_509_4290_0, i_10_509_4317_0, i_10_509_4566_0,
    o_10_509_0_0  );
  input  i_10_509_34_0, i_10_509_150_0, i_10_509_172_0, i_10_509_174_0,
    i_10_509_175_0, i_10_509_435_0, i_10_509_438_0, i_10_509_444_0,
    i_10_509_447_0, i_10_509_448_0, i_10_509_462_0, i_10_509_467_0,
    i_10_509_508_0, i_10_509_516_0, i_10_509_519_0, i_10_509_717_0,
    i_10_509_799_0, i_10_509_966_0, i_10_509_967_0, i_10_509_996_0,
    i_10_509_1029_0, i_10_509_1141_0, i_10_509_1164_0, i_10_509_1240_0,
    i_10_509_1245_0, i_10_509_1248_0, i_10_509_1309_0, i_10_509_1311_0,
    i_10_509_1366_0, i_10_509_1626_0, i_10_509_1652_0, i_10_509_1653_0,
    i_10_509_1655_0, i_10_509_1689_0, i_10_509_1690_0, i_10_509_1797_0,
    i_10_509_1821_0, i_10_509_1822_0, i_10_509_1912_0, i_10_509_1995_0,
    i_10_509_2005_0, i_10_509_2352_0, i_10_509_2353_0, i_10_509_2455_0,
    i_10_509_2469_0, i_10_509_2472_0, i_10_509_2473_0, i_10_509_2571_0,
    i_10_509_2628_0, i_10_509_2629_0, i_10_509_2659_0, i_10_509_2661_0,
    i_10_509_2706_0, i_10_509_2715_0, i_10_509_2716_0, i_10_509_2722_0,
    i_10_509_2731_0, i_10_509_2734_0, i_10_509_2742_0, i_10_509_2782_0,
    i_10_509_2830_0, i_10_509_2832_0, i_10_509_2883_0, i_10_509_2987_0,
    i_10_509_3037_0, i_10_509_3039_0, i_10_509_3046_0, i_10_509_3048_0,
    i_10_509_3075_0, i_10_509_3093_0, i_10_509_3157_0, i_10_509_3197_0,
    i_10_509_3284_0, i_10_509_3321_0, i_10_509_3322_0, i_10_509_3327_0,
    i_10_509_3391_0, i_10_509_3392_0, i_10_509_3468_0, i_10_509_3495_0,
    i_10_509_3525_0, i_10_509_3583_0, i_10_509_3585_0, i_10_509_3612_0,
    i_10_509_3613_0, i_10_509_3732_0, i_10_509_3780_0, i_10_509_3837_0,
    i_10_509_3876_0, i_10_509_3912_0, i_10_509_3982_0, i_10_509_4113_0,
    i_10_509_4173_0, i_10_509_4269_0, i_10_509_4272_0, i_10_509_4273_0,
    i_10_509_4282_0, i_10_509_4290_0, i_10_509_4317_0, i_10_509_4566_0;
  output o_10_509_0_0;
  assign o_10_509_0_0 = ~((~i_10_509_2472_0 & ((~i_10_509_150_0 & ((~i_10_509_966_0 & ~i_10_509_1248_0 & ~i_10_509_2706_0 & ~i_10_509_3046_0) | (~i_10_509_1690_0 & ~i_10_509_4272_0))) | (~i_10_509_3468_0 & ((~i_10_509_444_0 & ~i_10_509_3075_0) | (i_10_509_175_0 & ~i_10_509_1655_0 & ~i_10_509_3837_0))))) | (~i_10_509_516_0 & ((~i_10_509_799_0 & ~i_10_509_1626_0 & ~i_10_509_2571_0 & ~i_10_509_3048_0 & i_10_509_3391_0) | (~i_10_509_172_0 & ~i_10_509_519_0 & ~i_10_509_2715_0 & i_10_509_2734_0 & i_10_509_3048_0 & i_10_509_4282_0))) | (~i_10_509_519_0 & ((~i_10_509_174_0 & ~i_10_509_717_0 & ~i_10_509_966_0 & ~i_10_509_1626_0 & ~i_10_509_2571_0 & ~i_10_509_2706_0) | (i_10_509_2472_0 & ~i_10_509_3391_0 & ~i_10_509_4173_0 & ~i_10_509_4566_0))) | (~i_10_509_1164_0 & ((i_10_509_175_0 & ~i_10_509_1626_0 & ~i_10_509_2473_0 & ~i_10_509_2830_0) | (~i_10_509_1655_0 & ~i_10_509_2352_0 & ~i_10_509_2706_0 & ~i_10_509_3912_0 & i_10_509_4290_0))) | (~i_10_509_1626_0 & ((~i_10_509_966_0 & ~i_10_509_1689_0 & ~i_10_509_3495_0 & ~i_10_509_4269_0) | (~i_10_509_448_0 & ~i_10_509_2706_0 & ~i_10_509_2715_0 & ~i_10_509_3982_0 & ~i_10_509_4566_0))) | (~i_10_509_966_0 & ((~i_10_509_2353_0 & i_10_509_2629_0) | (~i_10_509_1652_0 & ~i_10_509_1821_0 & i_10_509_3039_0 & ~i_10_509_3495_0 & i_10_509_4269_0))) | (i_10_509_1655_0 & ((i_10_509_3039_0 & ~i_10_509_3495_0 & ~i_10_509_4173_0) | (i_10_509_2731_0 & i_10_509_2734_0 & ~i_10_509_4269_0))) | (~i_10_509_3391_0 & ((i_10_509_1822_0 & (i_10_509_3039_0 | (~i_10_509_1652_0 & ~i_10_509_2715_0 & ~i_10_509_4272_0))) | (~i_10_509_1029_0 & i_10_509_1309_0 & ~i_10_509_2473_0 & ~i_10_509_3837_0))) | (i_10_509_4273_0 & ((~i_10_509_799_0 & ~i_10_509_2706_0 & ~i_10_509_2715_0 & ~i_10_509_3048_0) | (~i_10_509_1821_0 & ~i_10_509_3495_0 & i_10_509_3837_0 & i_10_509_3982_0 & ~i_10_509_4282_0))) | (~i_10_509_3495_0 & ((i_10_509_172_0 & i_10_509_467_0 & ~i_10_509_2005_0 & ~i_10_509_2782_0 & ~i_10_509_2987_0) | (~i_10_509_3468_0 & i_10_509_3837_0 & ~i_10_509_3912_0 & ~i_10_509_4173_0 & ~i_10_509_4566_0))) | (i_10_509_2830_0 & i_10_509_3039_0 & i_10_509_3837_0) | (~i_10_509_1689_0 & i_10_509_2731_0 & ~i_10_509_4273_0 & ~i_10_509_4290_0));
endmodule



// Benchmark "kernel_10_510" written by ABC on Sun Jul 19 10:29:56 2020

module kernel_10_510 ( 
    i_10_510_35_0, i_10_510_71_0, i_10_510_124_0, i_10_510_125_0,
    i_10_510_154_0, i_10_510_178_0, i_10_510_215_0, i_10_510_265_0,
    i_10_510_279_0, i_10_510_317_0, i_10_510_390_0, i_10_510_410_0,
    i_10_510_440_0, i_10_510_445_0, i_10_510_465_0, i_10_510_533_0,
    i_10_510_562_0, i_10_510_565_0, i_10_510_566_0, i_10_510_869_0,
    i_10_510_1000_0, i_10_510_1006_0, i_10_510_1163_0, i_10_510_1265_0,
    i_10_510_1277_0, i_10_510_1319_0, i_10_510_1361_0, i_10_510_1363_0,
    i_10_510_1438_0, i_10_510_1439_0, i_10_510_1525_0, i_10_510_1652_0,
    i_10_510_1654_0, i_10_510_1714_0, i_10_510_1769_0, i_10_510_1823_0,
    i_10_510_1913_0, i_10_510_1922_0, i_10_510_1951_0, i_10_510_1952_0,
    i_10_510_2023_0, i_10_510_2033_0, i_10_510_2083_0, i_10_510_2096_0,
    i_10_510_2186_0, i_10_510_2200_0, i_10_510_2201_0, i_10_510_2203_0,
    i_10_510_2237_0, i_10_510_2240_0, i_10_510_2257_0, i_10_510_2312_0,
    i_10_510_2363_0, i_10_510_2378_0, i_10_510_2453_0, i_10_510_2470_0,
    i_10_510_2514_0, i_10_510_2614_0, i_10_510_2615_0, i_10_510_2633_0,
    i_10_510_2636_0, i_10_510_2786_0, i_10_510_2831_0, i_10_510_2881_0,
    i_10_510_2924_0, i_10_510_2960_0, i_10_510_2980_0, i_10_510_2986_0,
    i_10_510_3039_0, i_10_510_3040_0, i_10_510_3041_0, i_10_510_3046_0,
    i_10_510_3070_0, i_10_510_3071_0, i_10_510_3073_0, i_10_510_3159_0,
    i_10_510_3160_0, i_10_510_3434_0, i_10_510_3448_0, i_10_510_3469_0,
    i_10_510_3470_0, i_10_510_3520_0, i_10_510_3544_0, i_10_510_3545_0,
    i_10_510_3562_0, i_10_510_3563_0, i_10_510_3586_0, i_10_510_3590_0,
    i_10_510_3647_0, i_10_510_3652_0, i_10_510_3653_0, i_10_510_3682_0,
    i_10_510_3685_0, i_10_510_3788_0, i_10_510_4167_0, i_10_510_4168_0,
    i_10_510_4169_0, i_10_510_4234_0, i_10_510_4278_0, i_10_510_4531_0,
    o_10_510_0_0  );
  input  i_10_510_35_0, i_10_510_71_0, i_10_510_124_0, i_10_510_125_0,
    i_10_510_154_0, i_10_510_178_0, i_10_510_215_0, i_10_510_265_0,
    i_10_510_279_0, i_10_510_317_0, i_10_510_390_0, i_10_510_410_0,
    i_10_510_440_0, i_10_510_445_0, i_10_510_465_0, i_10_510_533_0,
    i_10_510_562_0, i_10_510_565_0, i_10_510_566_0, i_10_510_869_0,
    i_10_510_1000_0, i_10_510_1006_0, i_10_510_1163_0, i_10_510_1265_0,
    i_10_510_1277_0, i_10_510_1319_0, i_10_510_1361_0, i_10_510_1363_0,
    i_10_510_1438_0, i_10_510_1439_0, i_10_510_1525_0, i_10_510_1652_0,
    i_10_510_1654_0, i_10_510_1714_0, i_10_510_1769_0, i_10_510_1823_0,
    i_10_510_1913_0, i_10_510_1922_0, i_10_510_1951_0, i_10_510_1952_0,
    i_10_510_2023_0, i_10_510_2033_0, i_10_510_2083_0, i_10_510_2096_0,
    i_10_510_2186_0, i_10_510_2200_0, i_10_510_2201_0, i_10_510_2203_0,
    i_10_510_2237_0, i_10_510_2240_0, i_10_510_2257_0, i_10_510_2312_0,
    i_10_510_2363_0, i_10_510_2378_0, i_10_510_2453_0, i_10_510_2470_0,
    i_10_510_2514_0, i_10_510_2614_0, i_10_510_2615_0, i_10_510_2633_0,
    i_10_510_2636_0, i_10_510_2786_0, i_10_510_2831_0, i_10_510_2881_0,
    i_10_510_2924_0, i_10_510_2960_0, i_10_510_2980_0, i_10_510_2986_0,
    i_10_510_3039_0, i_10_510_3040_0, i_10_510_3041_0, i_10_510_3046_0,
    i_10_510_3070_0, i_10_510_3071_0, i_10_510_3073_0, i_10_510_3159_0,
    i_10_510_3160_0, i_10_510_3434_0, i_10_510_3448_0, i_10_510_3469_0,
    i_10_510_3470_0, i_10_510_3520_0, i_10_510_3544_0, i_10_510_3545_0,
    i_10_510_3562_0, i_10_510_3563_0, i_10_510_3586_0, i_10_510_3590_0,
    i_10_510_3647_0, i_10_510_3652_0, i_10_510_3653_0, i_10_510_3682_0,
    i_10_510_3685_0, i_10_510_3788_0, i_10_510_4167_0, i_10_510_4168_0,
    i_10_510_4169_0, i_10_510_4234_0, i_10_510_4278_0, i_10_510_4531_0;
  output o_10_510_0_0;
  assign o_10_510_0_0 = 0;
endmodule



// Benchmark "kernel_10_511" written by ABC on Sun Jul 19 10:29:57 2020

module kernel_10_511 ( 
    i_10_511_174_0, i_10_511_248_0, i_10_511_266_0, i_10_511_270_0,
    i_10_511_273_0, i_10_511_274_0, i_10_511_284_0, i_10_511_285_0,
    i_10_511_293_0, i_10_511_395_0, i_10_511_500_0, i_10_511_503_0,
    i_10_511_629_0, i_10_511_797_0, i_10_511_1003_0, i_10_511_1004_0,
    i_10_511_1086_0, i_10_511_1105_0, i_10_511_1115_0, i_10_511_1120_0,
    i_10_511_1138_0, i_10_511_1223_0, i_10_511_1238_0, i_10_511_1240_0,
    i_10_511_1241_0, i_10_511_1301_0, i_10_511_1303_0, i_10_511_1384_0,
    i_10_511_1436_0, i_10_511_1544_0, i_10_511_1545_0, i_10_511_1547_0,
    i_10_511_1578_0, i_10_511_1581_0, i_10_511_1582_0, i_10_511_1625_0,
    i_10_511_1628_0, i_10_511_1651_0, i_10_511_1690_0, i_10_511_1691_0,
    i_10_511_1733_0, i_10_511_1736_0, i_10_511_1824_0, i_10_511_2003_0,
    i_10_511_2006_0, i_10_511_2030_0, i_10_511_2033_0, i_10_511_2200_0,
    i_10_511_2354_0, i_10_511_2363_0, i_10_511_2453_0, i_10_511_2462_0,
    i_10_511_2471_0, i_10_511_2473_0, i_10_511_2474_0, i_10_511_2510_0,
    i_10_511_2570_0, i_10_511_2573_0, i_10_511_2631_0, i_10_511_2632_0,
    i_10_511_2633_0, i_10_511_2634_0, i_10_511_2635_0, i_10_511_2636_0,
    i_10_511_2641_0, i_10_511_2644_0, i_10_511_2701_0, i_10_511_2705_0,
    i_10_511_2717_0, i_10_511_2785_0, i_10_511_2830_0, i_10_511_2834_0,
    i_10_511_2849_0, i_10_511_2882_0, i_10_511_2883_0, i_10_511_3071_0,
    i_10_511_3278_0, i_10_511_3281_0, i_10_511_3384_0, i_10_511_3388_0,
    i_10_511_3392_0, i_10_511_3408_0, i_10_511_3470_0, i_10_511_3473_0,
    i_10_511_3542_0, i_10_511_3545_0, i_10_511_3584_0, i_10_511_3587_0,
    i_10_511_3613_0, i_10_511_3784_0, i_10_511_3838_0, i_10_511_3839_0,
    i_10_511_3843_0, i_10_511_3853_0, i_10_511_3854_0, i_10_511_4113_0,
    i_10_511_4126_0, i_10_511_4127_0, i_10_511_4283_0, i_10_511_4589_0,
    o_10_511_0_0  );
  input  i_10_511_174_0, i_10_511_248_0, i_10_511_266_0, i_10_511_270_0,
    i_10_511_273_0, i_10_511_274_0, i_10_511_284_0, i_10_511_285_0,
    i_10_511_293_0, i_10_511_395_0, i_10_511_500_0, i_10_511_503_0,
    i_10_511_629_0, i_10_511_797_0, i_10_511_1003_0, i_10_511_1004_0,
    i_10_511_1086_0, i_10_511_1105_0, i_10_511_1115_0, i_10_511_1120_0,
    i_10_511_1138_0, i_10_511_1223_0, i_10_511_1238_0, i_10_511_1240_0,
    i_10_511_1241_0, i_10_511_1301_0, i_10_511_1303_0, i_10_511_1384_0,
    i_10_511_1436_0, i_10_511_1544_0, i_10_511_1545_0, i_10_511_1547_0,
    i_10_511_1578_0, i_10_511_1581_0, i_10_511_1582_0, i_10_511_1625_0,
    i_10_511_1628_0, i_10_511_1651_0, i_10_511_1690_0, i_10_511_1691_0,
    i_10_511_1733_0, i_10_511_1736_0, i_10_511_1824_0, i_10_511_2003_0,
    i_10_511_2006_0, i_10_511_2030_0, i_10_511_2033_0, i_10_511_2200_0,
    i_10_511_2354_0, i_10_511_2363_0, i_10_511_2453_0, i_10_511_2462_0,
    i_10_511_2471_0, i_10_511_2473_0, i_10_511_2474_0, i_10_511_2510_0,
    i_10_511_2570_0, i_10_511_2573_0, i_10_511_2631_0, i_10_511_2632_0,
    i_10_511_2633_0, i_10_511_2634_0, i_10_511_2635_0, i_10_511_2636_0,
    i_10_511_2641_0, i_10_511_2644_0, i_10_511_2701_0, i_10_511_2705_0,
    i_10_511_2717_0, i_10_511_2785_0, i_10_511_2830_0, i_10_511_2834_0,
    i_10_511_2849_0, i_10_511_2882_0, i_10_511_2883_0, i_10_511_3071_0,
    i_10_511_3278_0, i_10_511_3281_0, i_10_511_3384_0, i_10_511_3388_0,
    i_10_511_3392_0, i_10_511_3408_0, i_10_511_3470_0, i_10_511_3473_0,
    i_10_511_3542_0, i_10_511_3545_0, i_10_511_3584_0, i_10_511_3587_0,
    i_10_511_3613_0, i_10_511_3784_0, i_10_511_3838_0, i_10_511_3839_0,
    i_10_511_3843_0, i_10_511_3853_0, i_10_511_3854_0, i_10_511_4113_0,
    i_10_511_4126_0, i_10_511_4127_0, i_10_511_4283_0, i_10_511_4589_0;
  output o_10_511_0_0;
  assign o_10_511_0_0 = ~((~i_10_511_1625_0 & ((~i_10_511_266_0 & ((i_10_511_174_0 & ~i_10_511_1004_0 & ~i_10_511_1628_0) | (~i_10_511_1733_0 & ~i_10_511_2573_0 & ~i_10_511_3584_0))) | (~i_10_511_395_0 & ~i_10_511_1004_0 & ~i_10_511_2030_0 & ~i_10_511_2453_0 & ~i_10_511_2717_0 & ~i_10_511_3388_0 & ~i_10_511_3408_0))) | (~i_10_511_395_0 & i_10_511_1436_0 & ((~i_10_511_797_0 & i_10_511_2200_0 & ~i_10_511_2573_0 & ~i_10_511_3470_0) | (i_10_511_1240_0 & ~i_10_511_1733_0 & ~i_10_511_2717_0 & ~i_10_511_3854_0))) | (~i_10_511_1733_0 & ((i_10_511_2633_0 & i_10_511_3613_0 & ~i_10_511_3853_0) | (~i_10_511_1544_0 & ~i_10_511_2003_0 & ~i_10_511_3545_0 & ~i_10_511_3784_0 & i_10_511_3839_0 & ~i_10_511_4127_0))) | (~i_10_511_1544_0 & ((~i_10_511_3470_0 & ~i_10_511_3587_0) | (i_10_511_1241_0 & ~i_10_511_2003_0 & ~i_10_511_2573_0 & i_10_511_3613_0 & ~i_10_511_4283_0))) | (~i_10_511_3613_0 & ((~i_10_511_1691_0 & i_10_511_2633_0 & i_10_511_3854_0) | (~i_10_511_1628_0 & ~i_10_511_2033_0 & ~i_10_511_3278_0 & ~i_10_511_4283_0))) | (~i_10_511_3278_0 & i_10_511_3854_0 & ((i_10_511_1003_0 & ~i_10_511_1004_0) | (i_10_511_1240_0 & ~i_10_511_2006_0 & ~i_10_511_2453_0))) | (~i_10_511_174_0 & ~i_10_511_1581_0 & i_10_511_2631_0) | (~i_10_511_2471_0 & ~i_10_511_2705_0 & ~i_10_511_3071_0 & ~i_10_511_3384_0 & ~i_10_511_3542_0 & ~i_10_511_3545_0) | (~i_10_511_3470_0 & i_10_511_3587_0 & ~i_10_511_3838_0));
endmodule



module kernel_10 (i_10_0, i_10_1, i_10_2, i_10_3, i_10_4, i_10_5, i_10_6, i_10_7, i_10_8, i_10_9, i_10_10, i_10_11, i_10_12, i_10_13, i_10_14, i_10_15, i_10_16, i_10_17, i_10_18, i_10_19, i_10_20, i_10_21, i_10_22, i_10_23, i_10_24, i_10_25, i_10_26, i_10_27, i_10_28, i_10_29, i_10_30, i_10_31, i_10_32, i_10_33, i_10_34, i_10_35, i_10_36, i_10_37, i_10_38, i_10_39, i_10_40, i_10_41, i_10_42, i_10_43, i_10_44, i_10_45, i_10_46, i_10_47, i_10_48, i_10_49, i_10_50, i_10_51, i_10_52, i_10_53, i_10_54, i_10_55, i_10_56, i_10_57, i_10_58, i_10_59, i_10_60, i_10_61, i_10_62, i_10_63, i_10_64, i_10_65, i_10_66, i_10_67, i_10_68, i_10_69, i_10_70, i_10_71, i_10_72, i_10_73, i_10_74, i_10_75, i_10_76, i_10_77, i_10_78, i_10_79, i_10_80, i_10_81, i_10_82, i_10_83, i_10_84, i_10_85, i_10_86, i_10_87, i_10_88, i_10_89, i_10_90, i_10_91, i_10_92, i_10_93, i_10_94, i_10_95, i_10_96, i_10_97, i_10_98, i_10_99, i_10_100, i_10_101, i_10_102, i_10_103, i_10_104, i_10_105, i_10_106, i_10_107, i_10_108, i_10_109, i_10_110, i_10_111, i_10_112, i_10_113, i_10_114, i_10_115, i_10_116, i_10_117, i_10_118, i_10_119, i_10_120, i_10_121, i_10_122, i_10_123, i_10_124, i_10_125, i_10_126, i_10_127, i_10_128, i_10_129, i_10_130, i_10_131, i_10_132, i_10_133, i_10_134, i_10_135, i_10_136, i_10_137, i_10_138, i_10_139, i_10_140, i_10_141, i_10_142, i_10_143, i_10_144, i_10_145, i_10_146, i_10_147, i_10_148, i_10_149, i_10_150, i_10_151, i_10_152, i_10_153, i_10_154, i_10_155, i_10_156, i_10_157, i_10_158, i_10_159, i_10_160, i_10_161, i_10_162, i_10_163, i_10_164, i_10_165, i_10_166, i_10_167, i_10_168, i_10_169, i_10_170, i_10_171, i_10_172, i_10_173, i_10_174, i_10_175, i_10_176, i_10_177, i_10_178, i_10_179, i_10_180, i_10_181, i_10_182, i_10_183, i_10_184, i_10_185, i_10_186, i_10_187, i_10_188, i_10_189, i_10_190, i_10_191, i_10_192, i_10_193, i_10_194, i_10_195, i_10_196, i_10_197, i_10_198, i_10_199, i_10_200, i_10_201, i_10_202, i_10_203, i_10_204, i_10_205, i_10_206, i_10_207, i_10_208, i_10_209, i_10_210, i_10_211, i_10_212, i_10_213, i_10_214, i_10_215, i_10_216, i_10_217, i_10_218, i_10_219, i_10_220, i_10_221, i_10_222, i_10_223, i_10_224, i_10_225, i_10_226, i_10_227, i_10_228, i_10_229, i_10_230, i_10_231, i_10_232, i_10_233, i_10_234, i_10_235, i_10_236, i_10_237, i_10_238, i_10_239, i_10_240, i_10_241, i_10_242, i_10_243, i_10_244, i_10_245, i_10_246, i_10_247, i_10_248, i_10_249, i_10_250, i_10_251, i_10_252, i_10_253, i_10_254, i_10_255, i_10_256, i_10_257, i_10_258, i_10_259, i_10_260, i_10_261, i_10_262, i_10_263, i_10_264, i_10_265, i_10_266, i_10_267, i_10_268, i_10_269, i_10_270, i_10_271, i_10_272, i_10_273, i_10_274, i_10_275, i_10_276, i_10_277, i_10_278, i_10_279, i_10_280, i_10_281, i_10_282, i_10_283, i_10_284, i_10_285, i_10_286, i_10_287, i_10_288, i_10_289, i_10_290, i_10_291, i_10_292, i_10_293, i_10_294, i_10_295, i_10_296, i_10_297, i_10_298, i_10_299, i_10_300, i_10_301, i_10_302, i_10_303, i_10_304, i_10_305, i_10_306, i_10_307, i_10_308, i_10_309, i_10_310, i_10_311, i_10_312, i_10_313, i_10_314, i_10_315, i_10_316, i_10_317, i_10_318, i_10_319, i_10_320, i_10_321, i_10_322, i_10_323, i_10_324, i_10_325, i_10_326, i_10_327, i_10_328, i_10_329, i_10_330, i_10_331, i_10_332, i_10_333, i_10_334, i_10_335, i_10_336, i_10_337, i_10_338, i_10_339, i_10_340, i_10_341, i_10_342, i_10_343, i_10_344, i_10_345, i_10_346, i_10_347, i_10_348, i_10_349, i_10_350, i_10_351, i_10_352, i_10_353, i_10_354, i_10_355, i_10_356, i_10_357, i_10_358, i_10_359, i_10_360, i_10_361, i_10_362, i_10_363, i_10_364, i_10_365, i_10_366, i_10_367, i_10_368, i_10_369, i_10_370, i_10_371, i_10_372, i_10_373, i_10_374, i_10_375, i_10_376, i_10_377, i_10_378, i_10_379, i_10_380, i_10_381, i_10_382, i_10_383, i_10_384, i_10_385, i_10_386, i_10_387, i_10_388, i_10_389, i_10_390, i_10_391, i_10_392, i_10_393, i_10_394, i_10_395, i_10_396, i_10_397, i_10_398, i_10_399, i_10_400, i_10_401, i_10_402, i_10_403, i_10_404, i_10_405, i_10_406, i_10_407, i_10_408, i_10_409, i_10_410, i_10_411, i_10_412, i_10_413, i_10_414, i_10_415, i_10_416, i_10_417, i_10_418, i_10_419, i_10_420, i_10_421, i_10_422, i_10_423, i_10_424, i_10_425, i_10_426, i_10_427, i_10_428, i_10_429, i_10_430, i_10_431, i_10_432, i_10_433, i_10_434, i_10_435, i_10_436, i_10_437, i_10_438, i_10_439, i_10_440, i_10_441, i_10_442, i_10_443, i_10_444, i_10_445, i_10_446, i_10_447, i_10_448, i_10_449, i_10_450, i_10_451, i_10_452, i_10_453, i_10_454, i_10_455, i_10_456, i_10_457, i_10_458, i_10_459, i_10_460, i_10_461, i_10_462, i_10_463, i_10_464, i_10_465, i_10_466, i_10_467, i_10_468, i_10_469, i_10_470, i_10_471, i_10_472, i_10_473, i_10_474, i_10_475, i_10_476, i_10_477, i_10_478, i_10_479, i_10_480, i_10_481, i_10_482, i_10_483, i_10_484, i_10_485, i_10_486, i_10_487, i_10_488, i_10_489, i_10_490, i_10_491, i_10_492, i_10_493, i_10_494, i_10_495, i_10_496, i_10_497, i_10_498, i_10_499, i_10_500, i_10_501, i_10_502, i_10_503, i_10_504, i_10_505, i_10_506, i_10_507, i_10_508, i_10_509, i_10_510, i_10_511, i_10_512, i_10_513, i_10_514, i_10_515, i_10_516, i_10_517, i_10_518, i_10_519, i_10_520, i_10_521, i_10_522, i_10_523, i_10_524, i_10_525, i_10_526, i_10_527, i_10_528, i_10_529, i_10_530, i_10_531, i_10_532, i_10_533, i_10_534, i_10_535, i_10_536, i_10_537, i_10_538, i_10_539, i_10_540, i_10_541, i_10_542, i_10_543, i_10_544, i_10_545, i_10_546, i_10_547, i_10_548, i_10_549, i_10_550, i_10_551, i_10_552, i_10_553, i_10_554, i_10_555, i_10_556, i_10_557, i_10_558, i_10_559, i_10_560, i_10_561, i_10_562, i_10_563, i_10_564, i_10_565, i_10_566, i_10_567, i_10_568, i_10_569, i_10_570, i_10_571, i_10_572, i_10_573, i_10_574, i_10_575, i_10_576, i_10_577, i_10_578, i_10_579, i_10_580, i_10_581, i_10_582, i_10_583, i_10_584, i_10_585, i_10_586, i_10_587, i_10_588, i_10_589, i_10_590, i_10_591, i_10_592, i_10_593, i_10_594, i_10_595, i_10_596, i_10_597, i_10_598, i_10_599, i_10_600, i_10_601, i_10_602, i_10_603, i_10_604, i_10_605, i_10_606, i_10_607, i_10_608, i_10_609, i_10_610, i_10_611, i_10_612, i_10_613, i_10_614, i_10_615, i_10_616, i_10_617, i_10_618, i_10_619, i_10_620, i_10_621, i_10_622, i_10_623, i_10_624, i_10_625, i_10_626, i_10_627, i_10_628, i_10_629, i_10_630, i_10_631, i_10_632, i_10_633, i_10_634, i_10_635, i_10_636, i_10_637, i_10_638, i_10_639, i_10_640, i_10_641, i_10_642, i_10_643, i_10_644, i_10_645, i_10_646, i_10_647, i_10_648, i_10_649, i_10_650, i_10_651, i_10_652, i_10_653, i_10_654, i_10_655, i_10_656, i_10_657, i_10_658, i_10_659, i_10_660, i_10_661, i_10_662, i_10_663, i_10_664, i_10_665, i_10_666, i_10_667, i_10_668, i_10_669, i_10_670, i_10_671, i_10_672, i_10_673, i_10_674, i_10_675, i_10_676, i_10_677, i_10_678, i_10_679, i_10_680, i_10_681, i_10_682, i_10_683, i_10_684, i_10_685, i_10_686, i_10_687, i_10_688, i_10_689, i_10_690, i_10_691, i_10_692, i_10_693, i_10_694, i_10_695, i_10_696, i_10_697, i_10_698, i_10_699, i_10_700, i_10_701, i_10_702, i_10_703, i_10_704, i_10_705, i_10_706, i_10_707, i_10_708, i_10_709, i_10_710, i_10_711, i_10_712, i_10_713, i_10_714, i_10_715, i_10_716, i_10_717, i_10_718, i_10_719, i_10_720, i_10_721, i_10_722, i_10_723, i_10_724, i_10_725, i_10_726, i_10_727, i_10_728, i_10_729, i_10_730, i_10_731, i_10_732, i_10_733, i_10_734, i_10_735, i_10_736, i_10_737, i_10_738, i_10_739, i_10_740, i_10_741, i_10_742, i_10_743, i_10_744, i_10_745, i_10_746, i_10_747, i_10_748, i_10_749, i_10_750, i_10_751, i_10_752, i_10_753, i_10_754, i_10_755, i_10_756, i_10_757, i_10_758, i_10_759, i_10_760, i_10_761, i_10_762, i_10_763, i_10_764, i_10_765, i_10_766, i_10_767, i_10_768, i_10_769, i_10_770, i_10_771, i_10_772, i_10_773, i_10_774, i_10_775, i_10_776, i_10_777, i_10_778, i_10_779, i_10_780, i_10_781, i_10_782, i_10_783, i_10_784, i_10_785, i_10_786, i_10_787, i_10_788, i_10_789, i_10_790, i_10_791, i_10_792, i_10_793, i_10_794, i_10_795, i_10_796, i_10_797, i_10_798, i_10_799, i_10_800, i_10_801, i_10_802, i_10_803, i_10_804, i_10_805, i_10_806, i_10_807, i_10_808, i_10_809, i_10_810, i_10_811, i_10_812, i_10_813, i_10_814, i_10_815, i_10_816, i_10_817, i_10_818, i_10_819, i_10_820, i_10_821, i_10_822, i_10_823, i_10_824, i_10_825, i_10_826, i_10_827, i_10_828, i_10_829, i_10_830, i_10_831, i_10_832, i_10_833, i_10_834, i_10_835, i_10_836, i_10_837, i_10_838, i_10_839, i_10_840, i_10_841, i_10_842, i_10_843, i_10_844, i_10_845, i_10_846, i_10_847, i_10_848, i_10_849, i_10_850, i_10_851, i_10_852, i_10_853, i_10_854, i_10_855, i_10_856, i_10_857, i_10_858, i_10_859, i_10_860, i_10_861, i_10_862, i_10_863, i_10_864, i_10_865, i_10_866, i_10_867, i_10_868, i_10_869, i_10_870, i_10_871, i_10_872, i_10_873, i_10_874, i_10_875, i_10_876, i_10_877, i_10_878, i_10_879, i_10_880, i_10_881, i_10_882, i_10_883, i_10_884, i_10_885, i_10_886, i_10_887, i_10_888, i_10_889, i_10_890, i_10_891, i_10_892, i_10_893, i_10_894, i_10_895, i_10_896, i_10_897, i_10_898, i_10_899, i_10_900, i_10_901, i_10_902, i_10_903, i_10_904, i_10_905, i_10_906, i_10_907, i_10_908, i_10_909, i_10_910, i_10_911, i_10_912, i_10_913, i_10_914, i_10_915, i_10_916, i_10_917, i_10_918, i_10_919, i_10_920, i_10_921, i_10_922, i_10_923, i_10_924, i_10_925, i_10_926, i_10_927, i_10_928, i_10_929, i_10_930, i_10_931, i_10_932, i_10_933, i_10_934, i_10_935, i_10_936, i_10_937, i_10_938, i_10_939, i_10_940, i_10_941, i_10_942, i_10_943, i_10_944, i_10_945, i_10_946, i_10_947, i_10_948, i_10_949, i_10_950, i_10_951, i_10_952, i_10_953, i_10_954, i_10_955, i_10_956, i_10_957, i_10_958, i_10_959, i_10_960, i_10_961, i_10_962, i_10_963, i_10_964, i_10_965, i_10_966, i_10_967, i_10_968, i_10_969, i_10_970, i_10_971, i_10_972, i_10_973, i_10_974, i_10_975, i_10_976, i_10_977, i_10_978, i_10_979, i_10_980, i_10_981, i_10_982, i_10_983, i_10_984, i_10_985, i_10_986, i_10_987, i_10_988, i_10_989, i_10_990, i_10_991, i_10_992, i_10_993, i_10_994, i_10_995, i_10_996, i_10_997, i_10_998, i_10_999, i_10_1000, i_10_1001, i_10_1002, i_10_1003, i_10_1004, i_10_1005, i_10_1006, i_10_1007, i_10_1008, i_10_1009, i_10_1010, i_10_1011, i_10_1012, i_10_1013, i_10_1014, i_10_1015, i_10_1016, i_10_1017, i_10_1018, i_10_1019, i_10_1020, i_10_1021, i_10_1022, i_10_1023, i_10_1024, i_10_1025, i_10_1026, i_10_1027, i_10_1028, i_10_1029, i_10_1030, i_10_1031, i_10_1032, i_10_1033, i_10_1034, i_10_1035, i_10_1036, i_10_1037, i_10_1038, i_10_1039, i_10_1040, i_10_1041, i_10_1042, i_10_1043, i_10_1044, i_10_1045, i_10_1046, i_10_1047, i_10_1048, i_10_1049, i_10_1050, i_10_1051, i_10_1052, i_10_1053, i_10_1054, i_10_1055, i_10_1056, i_10_1057, i_10_1058, i_10_1059, i_10_1060, i_10_1061, i_10_1062, i_10_1063, i_10_1064, i_10_1065, i_10_1066, i_10_1067, i_10_1068, i_10_1069, i_10_1070, i_10_1071, i_10_1072, i_10_1073, i_10_1074, i_10_1075, i_10_1076, i_10_1077, i_10_1078, i_10_1079, i_10_1080, i_10_1081, i_10_1082, i_10_1083, i_10_1084, i_10_1085, i_10_1086, i_10_1087, i_10_1088, i_10_1089, i_10_1090, i_10_1091, i_10_1092, i_10_1093, i_10_1094, i_10_1095, i_10_1096, i_10_1097, i_10_1098, i_10_1099, i_10_1100, i_10_1101, i_10_1102, i_10_1103, i_10_1104, i_10_1105, i_10_1106, i_10_1107, i_10_1108, i_10_1109, i_10_1110, i_10_1111, i_10_1112, i_10_1113, i_10_1114, i_10_1115, i_10_1116, i_10_1117, i_10_1118, i_10_1119, i_10_1120, i_10_1121, i_10_1122, i_10_1123, i_10_1124, i_10_1125, i_10_1126, i_10_1127, i_10_1128, i_10_1129, i_10_1130, i_10_1131, i_10_1132, i_10_1133, i_10_1134, i_10_1135, i_10_1136, i_10_1137, i_10_1138, i_10_1139, i_10_1140, i_10_1141, i_10_1142, i_10_1143, i_10_1144, i_10_1145, i_10_1146, i_10_1147, i_10_1148, i_10_1149, i_10_1150, i_10_1151, i_10_1152, i_10_1153, i_10_1154, i_10_1155, i_10_1156, i_10_1157, i_10_1158, i_10_1159, i_10_1160, i_10_1161, i_10_1162, i_10_1163, i_10_1164, i_10_1165, i_10_1166, i_10_1167, i_10_1168, i_10_1169, i_10_1170, i_10_1171, i_10_1172, i_10_1173, i_10_1174, i_10_1175, i_10_1176, i_10_1177, i_10_1178, i_10_1179, i_10_1180, i_10_1181, i_10_1182, i_10_1183, i_10_1184, i_10_1185, i_10_1186, i_10_1187, i_10_1188, i_10_1189, i_10_1190, i_10_1191, i_10_1192, i_10_1193, i_10_1194, i_10_1195, i_10_1196, i_10_1197, i_10_1198, i_10_1199, i_10_1200, i_10_1201, i_10_1202, i_10_1203, i_10_1204, i_10_1205, i_10_1206, i_10_1207, i_10_1208, i_10_1209, i_10_1210, i_10_1211, i_10_1212, i_10_1213, i_10_1214, i_10_1215, i_10_1216, i_10_1217, i_10_1218, i_10_1219, i_10_1220, i_10_1221, i_10_1222, i_10_1223, i_10_1224, i_10_1225, i_10_1226, i_10_1227, i_10_1228, i_10_1229, i_10_1230, i_10_1231, i_10_1232, i_10_1233, i_10_1234, i_10_1235, i_10_1236, i_10_1237, i_10_1238, i_10_1239, i_10_1240, i_10_1241, i_10_1242, i_10_1243, i_10_1244, i_10_1245, i_10_1246, i_10_1247, i_10_1248, i_10_1249, i_10_1250, i_10_1251, i_10_1252, i_10_1253, i_10_1254, i_10_1255, i_10_1256, i_10_1257, i_10_1258, i_10_1259, i_10_1260, i_10_1261, i_10_1262, i_10_1263, i_10_1264, i_10_1265, i_10_1266, i_10_1267, i_10_1268, i_10_1269, i_10_1270, i_10_1271, i_10_1272, i_10_1273, i_10_1274, i_10_1275, i_10_1276, i_10_1277, i_10_1278, i_10_1279, i_10_1280, i_10_1281, i_10_1282, i_10_1283, i_10_1284, i_10_1285, i_10_1286, i_10_1287, i_10_1288, i_10_1289, i_10_1290, i_10_1291, i_10_1292, i_10_1293, i_10_1294, i_10_1295, i_10_1296, i_10_1297, i_10_1298, i_10_1299, i_10_1300, i_10_1301, i_10_1302, i_10_1303, i_10_1304, i_10_1305, i_10_1306, i_10_1307, i_10_1308, i_10_1309, i_10_1310, i_10_1311, i_10_1312, i_10_1313, i_10_1314, i_10_1315, i_10_1316, i_10_1317, i_10_1318, i_10_1319, i_10_1320, i_10_1321, i_10_1322, i_10_1323, i_10_1324, i_10_1325, i_10_1326, i_10_1327, i_10_1328, i_10_1329, i_10_1330, i_10_1331, i_10_1332, i_10_1333, i_10_1334, i_10_1335, i_10_1336, i_10_1337, i_10_1338, i_10_1339, i_10_1340, i_10_1341, i_10_1342, i_10_1343, i_10_1344, i_10_1345, i_10_1346, i_10_1347, i_10_1348, i_10_1349, i_10_1350, i_10_1351, i_10_1352, i_10_1353, i_10_1354, i_10_1355, i_10_1356, i_10_1357, i_10_1358, i_10_1359, i_10_1360, i_10_1361, i_10_1362, i_10_1363, i_10_1364, i_10_1365, i_10_1366, i_10_1367, i_10_1368, i_10_1369, i_10_1370, i_10_1371, i_10_1372, i_10_1373, i_10_1374, i_10_1375, i_10_1376, i_10_1377, i_10_1378, i_10_1379, i_10_1380, i_10_1381, i_10_1382, i_10_1383, i_10_1384, i_10_1385, i_10_1386, i_10_1387, i_10_1388, i_10_1389, i_10_1390, i_10_1391, i_10_1392, i_10_1393, i_10_1394, i_10_1395, i_10_1396, i_10_1397, i_10_1398, i_10_1399, i_10_1400, i_10_1401, i_10_1402, i_10_1403, i_10_1404, i_10_1405, i_10_1406, i_10_1407, i_10_1408, i_10_1409, i_10_1410, i_10_1411, i_10_1412, i_10_1413, i_10_1414, i_10_1415, i_10_1416, i_10_1417, i_10_1418, i_10_1419, i_10_1420, i_10_1421, i_10_1422, i_10_1423, i_10_1424, i_10_1425, i_10_1426, i_10_1427, i_10_1428, i_10_1429, i_10_1430, i_10_1431, i_10_1432, i_10_1433, i_10_1434, i_10_1435, i_10_1436, i_10_1437, i_10_1438, i_10_1439, i_10_1440, i_10_1441, i_10_1442, i_10_1443, i_10_1444, i_10_1445, i_10_1446, i_10_1447, i_10_1448, i_10_1449, i_10_1450, i_10_1451, i_10_1452, i_10_1453, i_10_1454, i_10_1455, i_10_1456, i_10_1457, i_10_1458, i_10_1459, i_10_1460, i_10_1461, i_10_1462, i_10_1463, i_10_1464, i_10_1465, i_10_1466, i_10_1467, i_10_1468, i_10_1469, i_10_1470, i_10_1471, i_10_1472, i_10_1473, i_10_1474, i_10_1475, i_10_1476, i_10_1477, i_10_1478, i_10_1479, i_10_1480, i_10_1481, i_10_1482, i_10_1483, i_10_1484, i_10_1485, i_10_1486, i_10_1487, i_10_1488, i_10_1489, i_10_1490, i_10_1491, i_10_1492, i_10_1493, i_10_1494, i_10_1495, i_10_1496, i_10_1497, i_10_1498, i_10_1499, i_10_1500, i_10_1501, i_10_1502, i_10_1503, i_10_1504, i_10_1505, i_10_1506, i_10_1507, i_10_1508, i_10_1509, i_10_1510, i_10_1511, i_10_1512, i_10_1513, i_10_1514, i_10_1515, i_10_1516, i_10_1517, i_10_1518, i_10_1519, i_10_1520, i_10_1521, i_10_1522, i_10_1523, i_10_1524, i_10_1525, i_10_1526, i_10_1527, i_10_1528, i_10_1529, i_10_1530, i_10_1531, i_10_1532, i_10_1533, i_10_1534, i_10_1535, i_10_1536, i_10_1537, i_10_1538, i_10_1539, i_10_1540, i_10_1541, i_10_1542, i_10_1543, i_10_1544, i_10_1545, i_10_1546, i_10_1547, i_10_1548, i_10_1549, i_10_1550, i_10_1551, i_10_1552, i_10_1553, i_10_1554, i_10_1555, i_10_1556, i_10_1557, i_10_1558, i_10_1559, i_10_1560, i_10_1561, i_10_1562, i_10_1563, i_10_1564, i_10_1565, i_10_1566, i_10_1567, i_10_1568, i_10_1569, i_10_1570, i_10_1571, i_10_1572, i_10_1573, i_10_1574, i_10_1575, i_10_1576, i_10_1577, i_10_1578, i_10_1579, i_10_1580, i_10_1581, i_10_1582, i_10_1583, i_10_1584, i_10_1585, i_10_1586, i_10_1587, i_10_1588, i_10_1589, i_10_1590, i_10_1591, i_10_1592, i_10_1593, i_10_1594, i_10_1595, i_10_1596, i_10_1597, i_10_1598, i_10_1599, i_10_1600, i_10_1601, i_10_1602, i_10_1603, i_10_1604, i_10_1605, i_10_1606, i_10_1607, i_10_1608, i_10_1609, i_10_1610, i_10_1611, i_10_1612, i_10_1613, i_10_1614, i_10_1615, i_10_1616, i_10_1617, i_10_1618, i_10_1619, i_10_1620, i_10_1621, i_10_1622, i_10_1623, i_10_1624, i_10_1625, i_10_1626, i_10_1627, i_10_1628, i_10_1629, i_10_1630, i_10_1631, i_10_1632, i_10_1633, i_10_1634, i_10_1635, i_10_1636, i_10_1637, i_10_1638, i_10_1639, i_10_1640, i_10_1641, i_10_1642, i_10_1643, i_10_1644, i_10_1645, i_10_1646, i_10_1647, i_10_1648, i_10_1649, i_10_1650, i_10_1651, i_10_1652, i_10_1653, i_10_1654, i_10_1655, i_10_1656, i_10_1657, i_10_1658, i_10_1659, i_10_1660, i_10_1661, i_10_1662, i_10_1663, i_10_1664, i_10_1665, i_10_1666, i_10_1667, i_10_1668, i_10_1669, i_10_1670, i_10_1671, i_10_1672, i_10_1673, i_10_1674, i_10_1675, i_10_1676, i_10_1677, i_10_1678, i_10_1679, i_10_1680, i_10_1681, i_10_1682, i_10_1683, i_10_1684, i_10_1685, i_10_1686, i_10_1687, i_10_1688, i_10_1689, i_10_1690, i_10_1691, i_10_1692, i_10_1693, i_10_1694, i_10_1695, i_10_1696, i_10_1697, i_10_1698, i_10_1699, i_10_1700, i_10_1701, i_10_1702, i_10_1703, i_10_1704, i_10_1705, i_10_1706, i_10_1707, i_10_1708, i_10_1709, i_10_1710, i_10_1711, i_10_1712, i_10_1713, i_10_1714, i_10_1715, i_10_1716, i_10_1717, i_10_1718, i_10_1719, i_10_1720, i_10_1721, i_10_1722, i_10_1723, i_10_1724, i_10_1725, i_10_1726, i_10_1727, i_10_1728, i_10_1729, i_10_1730, i_10_1731, i_10_1732, i_10_1733, i_10_1734, i_10_1735, i_10_1736, i_10_1737, i_10_1738, i_10_1739, i_10_1740, i_10_1741, i_10_1742, i_10_1743, i_10_1744, i_10_1745, i_10_1746, i_10_1747, i_10_1748, i_10_1749, i_10_1750, i_10_1751, i_10_1752, i_10_1753, i_10_1754, i_10_1755, i_10_1756, i_10_1757, i_10_1758, i_10_1759, i_10_1760, i_10_1761, i_10_1762, i_10_1763, i_10_1764, i_10_1765, i_10_1766, i_10_1767, i_10_1768, i_10_1769, i_10_1770, i_10_1771, i_10_1772, i_10_1773, i_10_1774, i_10_1775, i_10_1776, i_10_1777, i_10_1778, i_10_1779, i_10_1780, i_10_1781, i_10_1782, i_10_1783, i_10_1784, i_10_1785, i_10_1786, i_10_1787, i_10_1788, i_10_1789, i_10_1790, i_10_1791, i_10_1792, i_10_1793, i_10_1794, i_10_1795, i_10_1796, i_10_1797, i_10_1798, i_10_1799, i_10_1800, i_10_1801, i_10_1802, i_10_1803, i_10_1804, i_10_1805, i_10_1806, i_10_1807, i_10_1808, i_10_1809, i_10_1810, i_10_1811, i_10_1812, i_10_1813, i_10_1814, i_10_1815, i_10_1816, i_10_1817, i_10_1818, i_10_1819, i_10_1820, i_10_1821, i_10_1822, i_10_1823, i_10_1824, i_10_1825, i_10_1826, i_10_1827, i_10_1828, i_10_1829, i_10_1830, i_10_1831, i_10_1832, i_10_1833, i_10_1834, i_10_1835, i_10_1836, i_10_1837, i_10_1838, i_10_1839, i_10_1840, i_10_1841, i_10_1842, i_10_1843, i_10_1844, i_10_1845, i_10_1846, i_10_1847, i_10_1848, i_10_1849, i_10_1850, i_10_1851, i_10_1852, i_10_1853, i_10_1854, i_10_1855, i_10_1856, i_10_1857, i_10_1858, i_10_1859, i_10_1860, i_10_1861, i_10_1862, i_10_1863, i_10_1864, i_10_1865, i_10_1866, i_10_1867, i_10_1868, i_10_1869, i_10_1870, i_10_1871, i_10_1872, i_10_1873, i_10_1874, i_10_1875, i_10_1876, i_10_1877, i_10_1878, i_10_1879, i_10_1880, i_10_1881, i_10_1882, i_10_1883, i_10_1884, i_10_1885, i_10_1886, i_10_1887, i_10_1888, i_10_1889, i_10_1890, i_10_1891, i_10_1892, i_10_1893, i_10_1894, i_10_1895, i_10_1896, i_10_1897, i_10_1898, i_10_1899, i_10_1900, i_10_1901, i_10_1902, i_10_1903, i_10_1904, i_10_1905, i_10_1906, i_10_1907, i_10_1908, i_10_1909, i_10_1910, i_10_1911, i_10_1912, i_10_1913, i_10_1914, i_10_1915, i_10_1916, i_10_1917, i_10_1918, i_10_1919, i_10_1920, i_10_1921, i_10_1922, i_10_1923, i_10_1924, i_10_1925, i_10_1926, i_10_1927, i_10_1928, i_10_1929, i_10_1930, i_10_1931, i_10_1932, i_10_1933, i_10_1934, i_10_1935, i_10_1936, i_10_1937, i_10_1938, i_10_1939, i_10_1940, i_10_1941, i_10_1942, i_10_1943, i_10_1944, i_10_1945, i_10_1946, i_10_1947, i_10_1948, i_10_1949, i_10_1950, i_10_1951, i_10_1952, i_10_1953, i_10_1954, i_10_1955, i_10_1956, i_10_1957, i_10_1958, i_10_1959, i_10_1960, i_10_1961, i_10_1962, i_10_1963, i_10_1964, i_10_1965, i_10_1966, i_10_1967, i_10_1968, i_10_1969, i_10_1970, i_10_1971, i_10_1972, i_10_1973, i_10_1974, i_10_1975, i_10_1976, i_10_1977, i_10_1978, i_10_1979, i_10_1980, i_10_1981, i_10_1982, i_10_1983, i_10_1984, i_10_1985, i_10_1986, i_10_1987, i_10_1988, i_10_1989, i_10_1990, i_10_1991, i_10_1992, i_10_1993, i_10_1994, i_10_1995, i_10_1996, i_10_1997, i_10_1998, i_10_1999, i_10_2000, i_10_2001, i_10_2002, i_10_2003, i_10_2004, i_10_2005, i_10_2006, i_10_2007, i_10_2008, i_10_2009, i_10_2010, i_10_2011, i_10_2012, i_10_2013, i_10_2014, i_10_2015, i_10_2016, i_10_2017, i_10_2018, i_10_2019, i_10_2020, i_10_2021, i_10_2022, i_10_2023, i_10_2024, i_10_2025, i_10_2026, i_10_2027, i_10_2028, i_10_2029, i_10_2030, i_10_2031, i_10_2032, i_10_2033, i_10_2034, i_10_2035, i_10_2036, i_10_2037, i_10_2038, i_10_2039, i_10_2040, i_10_2041, i_10_2042, i_10_2043, i_10_2044, i_10_2045, i_10_2046, i_10_2047, i_10_2048, i_10_2049, i_10_2050, i_10_2051, i_10_2052, i_10_2053, i_10_2054, i_10_2055, i_10_2056, i_10_2057, i_10_2058, i_10_2059, i_10_2060, i_10_2061, i_10_2062, i_10_2063, i_10_2064, i_10_2065, i_10_2066, i_10_2067, i_10_2068, i_10_2069, i_10_2070, i_10_2071, i_10_2072, i_10_2073, i_10_2074, i_10_2075, i_10_2076, i_10_2077, i_10_2078, i_10_2079, i_10_2080, i_10_2081, i_10_2082, i_10_2083, i_10_2084, i_10_2085, i_10_2086, i_10_2087, i_10_2088, i_10_2089, i_10_2090, i_10_2091, i_10_2092, i_10_2093, i_10_2094, i_10_2095, i_10_2096, i_10_2097, i_10_2098, i_10_2099, i_10_2100, i_10_2101, i_10_2102, i_10_2103, i_10_2104, i_10_2105, i_10_2106, i_10_2107, i_10_2108, i_10_2109, i_10_2110, i_10_2111, i_10_2112, i_10_2113, i_10_2114, i_10_2115, i_10_2116, i_10_2117, i_10_2118, i_10_2119, i_10_2120, i_10_2121, i_10_2122, i_10_2123, i_10_2124, i_10_2125, i_10_2126, i_10_2127, i_10_2128, i_10_2129, i_10_2130, i_10_2131, i_10_2132, i_10_2133, i_10_2134, i_10_2135, i_10_2136, i_10_2137, i_10_2138, i_10_2139, i_10_2140, i_10_2141, i_10_2142, i_10_2143, i_10_2144, i_10_2145, i_10_2146, i_10_2147, i_10_2148, i_10_2149, i_10_2150, i_10_2151, i_10_2152, i_10_2153, i_10_2154, i_10_2155, i_10_2156, i_10_2157, i_10_2158, i_10_2159, i_10_2160, i_10_2161, i_10_2162, i_10_2163, i_10_2164, i_10_2165, i_10_2166, i_10_2167, i_10_2168, i_10_2169, i_10_2170, i_10_2171, i_10_2172, i_10_2173, i_10_2174, i_10_2175, i_10_2176, i_10_2177, i_10_2178, i_10_2179, i_10_2180, i_10_2181, i_10_2182, i_10_2183, i_10_2184, i_10_2185, i_10_2186, i_10_2187, i_10_2188, i_10_2189, i_10_2190, i_10_2191, i_10_2192, i_10_2193, i_10_2194, i_10_2195, i_10_2196, i_10_2197, i_10_2198, i_10_2199, i_10_2200, i_10_2201, i_10_2202, i_10_2203, i_10_2204, i_10_2205, i_10_2206, i_10_2207, i_10_2208, i_10_2209, i_10_2210, i_10_2211, i_10_2212, i_10_2213, i_10_2214, i_10_2215, i_10_2216, i_10_2217, i_10_2218, i_10_2219, i_10_2220, i_10_2221, i_10_2222, i_10_2223, i_10_2224, i_10_2225, i_10_2226, i_10_2227, i_10_2228, i_10_2229, i_10_2230, i_10_2231, i_10_2232, i_10_2233, i_10_2234, i_10_2235, i_10_2236, i_10_2237, i_10_2238, i_10_2239, i_10_2240, i_10_2241, i_10_2242, i_10_2243, i_10_2244, i_10_2245, i_10_2246, i_10_2247, i_10_2248, i_10_2249, i_10_2250, i_10_2251, i_10_2252, i_10_2253, i_10_2254, i_10_2255, i_10_2256, i_10_2257, i_10_2258, i_10_2259, i_10_2260, i_10_2261, i_10_2262, i_10_2263, i_10_2264, i_10_2265, i_10_2266, i_10_2267, i_10_2268, i_10_2269, i_10_2270, i_10_2271, i_10_2272, i_10_2273, i_10_2274, i_10_2275, i_10_2276, i_10_2277, i_10_2278, i_10_2279, i_10_2280, i_10_2281, i_10_2282, i_10_2283, i_10_2284, i_10_2285, i_10_2286, i_10_2287, i_10_2288, i_10_2289, i_10_2290, i_10_2291, i_10_2292, i_10_2293, i_10_2294, i_10_2295, i_10_2296, i_10_2297, i_10_2298, i_10_2299, i_10_2300, i_10_2301, i_10_2302, i_10_2303, i_10_2304, i_10_2305, i_10_2306, i_10_2307, i_10_2308, i_10_2309, i_10_2310, i_10_2311, i_10_2312, i_10_2313, i_10_2314, i_10_2315, i_10_2316, i_10_2317, i_10_2318, i_10_2319, i_10_2320, i_10_2321, i_10_2322, i_10_2323, i_10_2324, i_10_2325, i_10_2326, i_10_2327, i_10_2328, i_10_2329, i_10_2330, i_10_2331, i_10_2332, i_10_2333, i_10_2334, i_10_2335, i_10_2336, i_10_2337, i_10_2338, i_10_2339, i_10_2340, i_10_2341, i_10_2342, i_10_2343, i_10_2344, i_10_2345, i_10_2346, i_10_2347, i_10_2348, i_10_2349, i_10_2350, i_10_2351, i_10_2352, i_10_2353, i_10_2354, i_10_2355, i_10_2356, i_10_2357, i_10_2358, i_10_2359, i_10_2360, i_10_2361, i_10_2362, i_10_2363, i_10_2364, i_10_2365, i_10_2366, i_10_2367, i_10_2368, i_10_2369, i_10_2370, i_10_2371, i_10_2372, i_10_2373, i_10_2374, i_10_2375, i_10_2376, i_10_2377, i_10_2378, i_10_2379, i_10_2380, i_10_2381, i_10_2382, i_10_2383, i_10_2384, i_10_2385, i_10_2386, i_10_2387, i_10_2388, i_10_2389, i_10_2390, i_10_2391, i_10_2392, i_10_2393, i_10_2394, i_10_2395, i_10_2396, i_10_2397, i_10_2398, i_10_2399, i_10_2400, i_10_2401, i_10_2402, i_10_2403, i_10_2404, i_10_2405, i_10_2406, i_10_2407, i_10_2408, i_10_2409, i_10_2410, i_10_2411, i_10_2412, i_10_2413, i_10_2414, i_10_2415, i_10_2416, i_10_2417, i_10_2418, i_10_2419, i_10_2420, i_10_2421, i_10_2422, i_10_2423, i_10_2424, i_10_2425, i_10_2426, i_10_2427, i_10_2428, i_10_2429, i_10_2430, i_10_2431, i_10_2432, i_10_2433, i_10_2434, i_10_2435, i_10_2436, i_10_2437, i_10_2438, i_10_2439, i_10_2440, i_10_2441, i_10_2442, i_10_2443, i_10_2444, i_10_2445, i_10_2446, i_10_2447, i_10_2448, i_10_2449, i_10_2450, i_10_2451, i_10_2452, i_10_2453, i_10_2454, i_10_2455, i_10_2456, i_10_2457, i_10_2458, i_10_2459, i_10_2460, i_10_2461, i_10_2462, i_10_2463, i_10_2464, i_10_2465, i_10_2466, i_10_2467, i_10_2468, i_10_2469, i_10_2470, i_10_2471, i_10_2472, i_10_2473, i_10_2474, i_10_2475, i_10_2476, i_10_2477, i_10_2478, i_10_2479, i_10_2480, i_10_2481, i_10_2482, i_10_2483, i_10_2484, i_10_2485, i_10_2486, i_10_2487, i_10_2488, i_10_2489, i_10_2490, i_10_2491, i_10_2492, i_10_2493, i_10_2494, i_10_2495, i_10_2496, i_10_2497, i_10_2498, i_10_2499, i_10_2500, i_10_2501, i_10_2502, i_10_2503, i_10_2504, i_10_2505, i_10_2506, i_10_2507, i_10_2508, i_10_2509, i_10_2510, i_10_2511, i_10_2512, i_10_2513, i_10_2514, i_10_2515, i_10_2516, i_10_2517, i_10_2518, i_10_2519, i_10_2520, i_10_2521, i_10_2522, i_10_2523, i_10_2524, i_10_2525, i_10_2526, i_10_2527, i_10_2528, i_10_2529, i_10_2530, i_10_2531, i_10_2532, i_10_2533, i_10_2534, i_10_2535, i_10_2536, i_10_2537, i_10_2538, i_10_2539, i_10_2540, i_10_2541, i_10_2542, i_10_2543, i_10_2544, i_10_2545, i_10_2546, i_10_2547, i_10_2548, i_10_2549, i_10_2550, i_10_2551, i_10_2552, i_10_2553, i_10_2554, i_10_2555, i_10_2556, i_10_2557, i_10_2558, i_10_2559, i_10_2560, i_10_2561, i_10_2562, i_10_2563, i_10_2564, i_10_2565, i_10_2566, i_10_2567, i_10_2568, i_10_2569, i_10_2570, i_10_2571, i_10_2572, i_10_2573, i_10_2574, i_10_2575, i_10_2576, i_10_2577, i_10_2578, i_10_2579, i_10_2580, i_10_2581, i_10_2582, i_10_2583, i_10_2584, i_10_2585, i_10_2586, i_10_2587, i_10_2588, i_10_2589, i_10_2590, i_10_2591, i_10_2592, i_10_2593, i_10_2594, i_10_2595, i_10_2596, i_10_2597, i_10_2598, i_10_2599, i_10_2600, i_10_2601, i_10_2602, i_10_2603, i_10_2604, i_10_2605, i_10_2606, i_10_2607, i_10_2608, i_10_2609, i_10_2610, i_10_2611, i_10_2612, i_10_2613, i_10_2614, i_10_2615, i_10_2616, i_10_2617, i_10_2618, i_10_2619, i_10_2620, i_10_2621, i_10_2622, i_10_2623, i_10_2624, i_10_2625, i_10_2626, i_10_2627, i_10_2628, i_10_2629, i_10_2630, i_10_2631, i_10_2632, i_10_2633, i_10_2634, i_10_2635, i_10_2636, i_10_2637, i_10_2638, i_10_2639, i_10_2640, i_10_2641, i_10_2642, i_10_2643, i_10_2644, i_10_2645, i_10_2646, i_10_2647, i_10_2648, i_10_2649, i_10_2650, i_10_2651, i_10_2652, i_10_2653, i_10_2654, i_10_2655, i_10_2656, i_10_2657, i_10_2658, i_10_2659, i_10_2660, i_10_2661, i_10_2662, i_10_2663, i_10_2664, i_10_2665, i_10_2666, i_10_2667, i_10_2668, i_10_2669, i_10_2670, i_10_2671, i_10_2672, i_10_2673, i_10_2674, i_10_2675, i_10_2676, i_10_2677, i_10_2678, i_10_2679, i_10_2680, i_10_2681, i_10_2682, i_10_2683, i_10_2684, i_10_2685, i_10_2686, i_10_2687, i_10_2688, i_10_2689, i_10_2690, i_10_2691, i_10_2692, i_10_2693, i_10_2694, i_10_2695, i_10_2696, i_10_2697, i_10_2698, i_10_2699, i_10_2700, i_10_2701, i_10_2702, i_10_2703, i_10_2704, i_10_2705, i_10_2706, i_10_2707, i_10_2708, i_10_2709, i_10_2710, i_10_2711, i_10_2712, i_10_2713, i_10_2714, i_10_2715, i_10_2716, i_10_2717, i_10_2718, i_10_2719, i_10_2720, i_10_2721, i_10_2722, i_10_2723, i_10_2724, i_10_2725, i_10_2726, i_10_2727, i_10_2728, i_10_2729, i_10_2730, i_10_2731, i_10_2732, i_10_2733, i_10_2734, i_10_2735, i_10_2736, i_10_2737, i_10_2738, i_10_2739, i_10_2740, i_10_2741, i_10_2742, i_10_2743, i_10_2744, i_10_2745, i_10_2746, i_10_2747, i_10_2748, i_10_2749, i_10_2750, i_10_2751, i_10_2752, i_10_2753, i_10_2754, i_10_2755, i_10_2756, i_10_2757, i_10_2758, i_10_2759, i_10_2760, i_10_2761, i_10_2762, i_10_2763, i_10_2764, i_10_2765, i_10_2766, i_10_2767, i_10_2768, i_10_2769, i_10_2770, i_10_2771, i_10_2772, i_10_2773, i_10_2774, i_10_2775, i_10_2776, i_10_2777, i_10_2778, i_10_2779, i_10_2780, i_10_2781, i_10_2782, i_10_2783, i_10_2784, i_10_2785, i_10_2786, i_10_2787, i_10_2788, i_10_2789, i_10_2790, i_10_2791, i_10_2792, i_10_2793, i_10_2794, i_10_2795, i_10_2796, i_10_2797, i_10_2798, i_10_2799, i_10_2800, i_10_2801, i_10_2802, i_10_2803, i_10_2804, i_10_2805, i_10_2806, i_10_2807, i_10_2808, i_10_2809, i_10_2810, i_10_2811, i_10_2812, i_10_2813, i_10_2814, i_10_2815, i_10_2816, i_10_2817, i_10_2818, i_10_2819, i_10_2820, i_10_2821, i_10_2822, i_10_2823, i_10_2824, i_10_2825, i_10_2826, i_10_2827, i_10_2828, i_10_2829, i_10_2830, i_10_2831, i_10_2832, i_10_2833, i_10_2834, i_10_2835, i_10_2836, i_10_2837, i_10_2838, i_10_2839, i_10_2840, i_10_2841, i_10_2842, i_10_2843, i_10_2844, i_10_2845, i_10_2846, i_10_2847, i_10_2848, i_10_2849, i_10_2850, i_10_2851, i_10_2852, i_10_2853, i_10_2854, i_10_2855, i_10_2856, i_10_2857, i_10_2858, i_10_2859, i_10_2860, i_10_2861, i_10_2862, i_10_2863, i_10_2864, i_10_2865, i_10_2866, i_10_2867, i_10_2868, i_10_2869, i_10_2870, i_10_2871, i_10_2872, i_10_2873, i_10_2874, i_10_2875, i_10_2876, i_10_2877, i_10_2878, i_10_2879, i_10_2880, i_10_2881, i_10_2882, i_10_2883, i_10_2884, i_10_2885, i_10_2886, i_10_2887, i_10_2888, i_10_2889, i_10_2890, i_10_2891, i_10_2892, i_10_2893, i_10_2894, i_10_2895, i_10_2896, i_10_2897, i_10_2898, i_10_2899, i_10_2900, i_10_2901, i_10_2902, i_10_2903, i_10_2904, i_10_2905, i_10_2906, i_10_2907, i_10_2908, i_10_2909, i_10_2910, i_10_2911, i_10_2912, i_10_2913, i_10_2914, i_10_2915, i_10_2916, i_10_2917, i_10_2918, i_10_2919, i_10_2920, i_10_2921, i_10_2922, i_10_2923, i_10_2924, i_10_2925, i_10_2926, i_10_2927, i_10_2928, i_10_2929, i_10_2930, i_10_2931, i_10_2932, i_10_2933, i_10_2934, i_10_2935, i_10_2936, i_10_2937, i_10_2938, i_10_2939, i_10_2940, i_10_2941, i_10_2942, i_10_2943, i_10_2944, i_10_2945, i_10_2946, i_10_2947, i_10_2948, i_10_2949, i_10_2950, i_10_2951, i_10_2952, i_10_2953, i_10_2954, i_10_2955, i_10_2956, i_10_2957, i_10_2958, i_10_2959, i_10_2960, i_10_2961, i_10_2962, i_10_2963, i_10_2964, i_10_2965, i_10_2966, i_10_2967, i_10_2968, i_10_2969, i_10_2970, i_10_2971, i_10_2972, i_10_2973, i_10_2974, i_10_2975, i_10_2976, i_10_2977, i_10_2978, i_10_2979, i_10_2980, i_10_2981, i_10_2982, i_10_2983, i_10_2984, i_10_2985, i_10_2986, i_10_2987, i_10_2988, i_10_2989, i_10_2990, i_10_2991, i_10_2992, i_10_2993, i_10_2994, i_10_2995, i_10_2996, i_10_2997, i_10_2998, i_10_2999, i_10_3000, i_10_3001, i_10_3002, i_10_3003, i_10_3004, i_10_3005, i_10_3006, i_10_3007, i_10_3008, i_10_3009, i_10_3010, i_10_3011, i_10_3012, i_10_3013, i_10_3014, i_10_3015, i_10_3016, i_10_3017, i_10_3018, i_10_3019, i_10_3020, i_10_3021, i_10_3022, i_10_3023, i_10_3024, i_10_3025, i_10_3026, i_10_3027, i_10_3028, i_10_3029, i_10_3030, i_10_3031, i_10_3032, i_10_3033, i_10_3034, i_10_3035, i_10_3036, i_10_3037, i_10_3038, i_10_3039, i_10_3040, i_10_3041, i_10_3042, i_10_3043, i_10_3044, i_10_3045, i_10_3046, i_10_3047, i_10_3048, i_10_3049, i_10_3050, i_10_3051, i_10_3052, i_10_3053, i_10_3054, i_10_3055, i_10_3056, i_10_3057, i_10_3058, i_10_3059, i_10_3060, i_10_3061, i_10_3062, i_10_3063, i_10_3064, i_10_3065, i_10_3066, i_10_3067, i_10_3068, i_10_3069, i_10_3070, i_10_3071, i_10_3072, i_10_3073, i_10_3074, i_10_3075, i_10_3076, i_10_3077, i_10_3078, i_10_3079, i_10_3080, i_10_3081, i_10_3082, i_10_3083, i_10_3084, i_10_3085, i_10_3086, i_10_3087, i_10_3088, i_10_3089, i_10_3090, i_10_3091, i_10_3092, i_10_3093, i_10_3094, i_10_3095, i_10_3096, i_10_3097, i_10_3098, i_10_3099, i_10_3100, i_10_3101, i_10_3102, i_10_3103, i_10_3104, i_10_3105, i_10_3106, i_10_3107, i_10_3108, i_10_3109, i_10_3110, i_10_3111, i_10_3112, i_10_3113, i_10_3114, i_10_3115, i_10_3116, i_10_3117, i_10_3118, i_10_3119, i_10_3120, i_10_3121, i_10_3122, i_10_3123, i_10_3124, i_10_3125, i_10_3126, i_10_3127, i_10_3128, i_10_3129, i_10_3130, i_10_3131, i_10_3132, i_10_3133, i_10_3134, i_10_3135, i_10_3136, i_10_3137, i_10_3138, i_10_3139, i_10_3140, i_10_3141, i_10_3142, i_10_3143, i_10_3144, i_10_3145, i_10_3146, i_10_3147, i_10_3148, i_10_3149, i_10_3150, i_10_3151, i_10_3152, i_10_3153, i_10_3154, i_10_3155, i_10_3156, i_10_3157, i_10_3158, i_10_3159, i_10_3160, i_10_3161, i_10_3162, i_10_3163, i_10_3164, i_10_3165, i_10_3166, i_10_3167, i_10_3168, i_10_3169, i_10_3170, i_10_3171, i_10_3172, i_10_3173, i_10_3174, i_10_3175, i_10_3176, i_10_3177, i_10_3178, i_10_3179, i_10_3180, i_10_3181, i_10_3182, i_10_3183, i_10_3184, i_10_3185, i_10_3186, i_10_3187, i_10_3188, i_10_3189, i_10_3190, i_10_3191, i_10_3192, i_10_3193, i_10_3194, i_10_3195, i_10_3196, i_10_3197, i_10_3198, i_10_3199, i_10_3200, i_10_3201, i_10_3202, i_10_3203, i_10_3204, i_10_3205, i_10_3206, i_10_3207, i_10_3208, i_10_3209, i_10_3210, i_10_3211, i_10_3212, i_10_3213, i_10_3214, i_10_3215, i_10_3216, i_10_3217, i_10_3218, i_10_3219, i_10_3220, i_10_3221, i_10_3222, i_10_3223, i_10_3224, i_10_3225, i_10_3226, i_10_3227, i_10_3228, i_10_3229, i_10_3230, i_10_3231, i_10_3232, i_10_3233, i_10_3234, i_10_3235, i_10_3236, i_10_3237, i_10_3238, i_10_3239, i_10_3240, i_10_3241, i_10_3242, i_10_3243, i_10_3244, i_10_3245, i_10_3246, i_10_3247, i_10_3248, i_10_3249, i_10_3250, i_10_3251, i_10_3252, i_10_3253, i_10_3254, i_10_3255, i_10_3256, i_10_3257, i_10_3258, i_10_3259, i_10_3260, i_10_3261, i_10_3262, i_10_3263, i_10_3264, i_10_3265, i_10_3266, i_10_3267, i_10_3268, i_10_3269, i_10_3270, i_10_3271, i_10_3272, i_10_3273, i_10_3274, i_10_3275, i_10_3276, i_10_3277, i_10_3278, i_10_3279, i_10_3280, i_10_3281, i_10_3282, i_10_3283, i_10_3284, i_10_3285, i_10_3286, i_10_3287, i_10_3288, i_10_3289, i_10_3290, i_10_3291, i_10_3292, i_10_3293, i_10_3294, i_10_3295, i_10_3296, i_10_3297, i_10_3298, i_10_3299, i_10_3300, i_10_3301, i_10_3302, i_10_3303, i_10_3304, i_10_3305, i_10_3306, i_10_3307, i_10_3308, i_10_3309, i_10_3310, i_10_3311, i_10_3312, i_10_3313, i_10_3314, i_10_3315, i_10_3316, i_10_3317, i_10_3318, i_10_3319, i_10_3320, i_10_3321, i_10_3322, i_10_3323, i_10_3324, i_10_3325, i_10_3326, i_10_3327, i_10_3328, i_10_3329, i_10_3330, i_10_3331, i_10_3332, i_10_3333, i_10_3334, i_10_3335, i_10_3336, i_10_3337, i_10_3338, i_10_3339, i_10_3340, i_10_3341, i_10_3342, i_10_3343, i_10_3344, i_10_3345, i_10_3346, i_10_3347, i_10_3348, i_10_3349, i_10_3350, i_10_3351, i_10_3352, i_10_3353, i_10_3354, i_10_3355, i_10_3356, i_10_3357, i_10_3358, i_10_3359, i_10_3360, i_10_3361, i_10_3362, i_10_3363, i_10_3364, i_10_3365, i_10_3366, i_10_3367, i_10_3368, i_10_3369, i_10_3370, i_10_3371, i_10_3372, i_10_3373, i_10_3374, i_10_3375, i_10_3376, i_10_3377, i_10_3378, i_10_3379, i_10_3380, i_10_3381, i_10_3382, i_10_3383, i_10_3384, i_10_3385, i_10_3386, i_10_3387, i_10_3388, i_10_3389, i_10_3390, i_10_3391, i_10_3392, i_10_3393, i_10_3394, i_10_3395, i_10_3396, i_10_3397, i_10_3398, i_10_3399, i_10_3400, i_10_3401, i_10_3402, i_10_3403, i_10_3404, i_10_3405, i_10_3406, i_10_3407, i_10_3408, i_10_3409, i_10_3410, i_10_3411, i_10_3412, i_10_3413, i_10_3414, i_10_3415, i_10_3416, i_10_3417, i_10_3418, i_10_3419, i_10_3420, i_10_3421, i_10_3422, i_10_3423, i_10_3424, i_10_3425, i_10_3426, i_10_3427, i_10_3428, i_10_3429, i_10_3430, i_10_3431, i_10_3432, i_10_3433, i_10_3434, i_10_3435, i_10_3436, i_10_3437, i_10_3438, i_10_3439, i_10_3440, i_10_3441, i_10_3442, i_10_3443, i_10_3444, i_10_3445, i_10_3446, i_10_3447, i_10_3448, i_10_3449, i_10_3450, i_10_3451, i_10_3452, i_10_3453, i_10_3454, i_10_3455, i_10_3456, i_10_3457, i_10_3458, i_10_3459, i_10_3460, i_10_3461, i_10_3462, i_10_3463, i_10_3464, i_10_3465, i_10_3466, i_10_3467, i_10_3468, i_10_3469, i_10_3470, i_10_3471, i_10_3472, i_10_3473, i_10_3474, i_10_3475, i_10_3476, i_10_3477, i_10_3478, i_10_3479, i_10_3480, i_10_3481, i_10_3482, i_10_3483, i_10_3484, i_10_3485, i_10_3486, i_10_3487, i_10_3488, i_10_3489, i_10_3490, i_10_3491, i_10_3492, i_10_3493, i_10_3494, i_10_3495, i_10_3496, i_10_3497, i_10_3498, i_10_3499, i_10_3500, i_10_3501, i_10_3502, i_10_3503, i_10_3504, i_10_3505, i_10_3506, i_10_3507, i_10_3508, i_10_3509, i_10_3510, i_10_3511, i_10_3512, i_10_3513, i_10_3514, i_10_3515, i_10_3516, i_10_3517, i_10_3518, i_10_3519, i_10_3520, i_10_3521, i_10_3522, i_10_3523, i_10_3524, i_10_3525, i_10_3526, i_10_3527, i_10_3528, i_10_3529, i_10_3530, i_10_3531, i_10_3532, i_10_3533, i_10_3534, i_10_3535, i_10_3536, i_10_3537, i_10_3538, i_10_3539, i_10_3540, i_10_3541, i_10_3542, i_10_3543, i_10_3544, i_10_3545, i_10_3546, i_10_3547, i_10_3548, i_10_3549, i_10_3550, i_10_3551, i_10_3552, i_10_3553, i_10_3554, i_10_3555, i_10_3556, i_10_3557, i_10_3558, i_10_3559, i_10_3560, i_10_3561, i_10_3562, i_10_3563, i_10_3564, i_10_3565, i_10_3566, i_10_3567, i_10_3568, i_10_3569, i_10_3570, i_10_3571, i_10_3572, i_10_3573, i_10_3574, i_10_3575, i_10_3576, i_10_3577, i_10_3578, i_10_3579, i_10_3580, i_10_3581, i_10_3582, i_10_3583, i_10_3584, i_10_3585, i_10_3586, i_10_3587, i_10_3588, i_10_3589, i_10_3590, i_10_3591, i_10_3592, i_10_3593, i_10_3594, i_10_3595, i_10_3596, i_10_3597, i_10_3598, i_10_3599, i_10_3600, i_10_3601, i_10_3602, i_10_3603, i_10_3604, i_10_3605, i_10_3606, i_10_3607, i_10_3608, i_10_3609, i_10_3610, i_10_3611, i_10_3612, i_10_3613, i_10_3614, i_10_3615, i_10_3616, i_10_3617, i_10_3618, i_10_3619, i_10_3620, i_10_3621, i_10_3622, i_10_3623, i_10_3624, i_10_3625, i_10_3626, i_10_3627, i_10_3628, i_10_3629, i_10_3630, i_10_3631, i_10_3632, i_10_3633, i_10_3634, i_10_3635, i_10_3636, i_10_3637, i_10_3638, i_10_3639, i_10_3640, i_10_3641, i_10_3642, i_10_3643, i_10_3644, i_10_3645, i_10_3646, i_10_3647, i_10_3648, i_10_3649, i_10_3650, i_10_3651, i_10_3652, i_10_3653, i_10_3654, i_10_3655, i_10_3656, i_10_3657, i_10_3658, i_10_3659, i_10_3660, i_10_3661, i_10_3662, i_10_3663, i_10_3664, i_10_3665, i_10_3666, i_10_3667, i_10_3668, i_10_3669, i_10_3670, i_10_3671, i_10_3672, i_10_3673, i_10_3674, i_10_3675, i_10_3676, i_10_3677, i_10_3678, i_10_3679, i_10_3680, i_10_3681, i_10_3682, i_10_3683, i_10_3684, i_10_3685, i_10_3686, i_10_3687, i_10_3688, i_10_3689, i_10_3690, i_10_3691, i_10_3692, i_10_3693, i_10_3694, i_10_3695, i_10_3696, i_10_3697, i_10_3698, i_10_3699, i_10_3700, i_10_3701, i_10_3702, i_10_3703, i_10_3704, i_10_3705, i_10_3706, i_10_3707, i_10_3708, i_10_3709, i_10_3710, i_10_3711, i_10_3712, i_10_3713, i_10_3714, i_10_3715, i_10_3716, i_10_3717, i_10_3718, i_10_3719, i_10_3720, i_10_3721, i_10_3722, i_10_3723, i_10_3724, i_10_3725, i_10_3726, i_10_3727, i_10_3728, i_10_3729, i_10_3730, i_10_3731, i_10_3732, i_10_3733, i_10_3734, i_10_3735, i_10_3736, i_10_3737, i_10_3738, i_10_3739, i_10_3740, i_10_3741, i_10_3742, i_10_3743, i_10_3744, i_10_3745, i_10_3746, i_10_3747, i_10_3748, i_10_3749, i_10_3750, i_10_3751, i_10_3752, i_10_3753, i_10_3754, i_10_3755, i_10_3756, i_10_3757, i_10_3758, i_10_3759, i_10_3760, i_10_3761, i_10_3762, i_10_3763, i_10_3764, i_10_3765, i_10_3766, i_10_3767, i_10_3768, i_10_3769, i_10_3770, i_10_3771, i_10_3772, i_10_3773, i_10_3774, i_10_3775, i_10_3776, i_10_3777, i_10_3778, i_10_3779, i_10_3780, i_10_3781, i_10_3782, i_10_3783, i_10_3784, i_10_3785, i_10_3786, i_10_3787, i_10_3788, i_10_3789, i_10_3790, i_10_3791, i_10_3792, i_10_3793, i_10_3794, i_10_3795, i_10_3796, i_10_3797, i_10_3798, i_10_3799, i_10_3800, i_10_3801, i_10_3802, i_10_3803, i_10_3804, i_10_3805, i_10_3806, i_10_3807, i_10_3808, i_10_3809, i_10_3810, i_10_3811, i_10_3812, i_10_3813, i_10_3814, i_10_3815, i_10_3816, i_10_3817, i_10_3818, i_10_3819, i_10_3820, i_10_3821, i_10_3822, i_10_3823, i_10_3824, i_10_3825, i_10_3826, i_10_3827, i_10_3828, i_10_3829, i_10_3830, i_10_3831, i_10_3832, i_10_3833, i_10_3834, i_10_3835, i_10_3836, i_10_3837, i_10_3838, i_10_3839, i_10_3840, i_10_3841, i_10_3842, i_10_3843, i_10_3844, i_10_3845, i_10_3846, i_10_3847, i_10_3848, i_10_3849, i_10_3850, i_10_3851, i_10_3852, i_10_3853, i_10_3854, i_10_3855, i_10_3856, i_10_3857, i_10_3858, i_10_3859, i_10_3860, i_10_3861, i_10_3862, i_10_3863, i_10_3864, i_10_3865, i_10_3866, i_10_3867, i_10_3868, i_10_3869, i_10_3870, i_10_3871, i_10_3872, i_10_3873, i_10_3874, i_10_3875, i_10_3876, i_10_3877, i_10_3878, i_10_3879, i_10_3880, i_10_3881, i_10_3882, i_10_3883, i_10_3884, i_10_3885, i_10_3886, i_10_3887, i_10_3888, i_10_3889, i_10_3890, i_10_3891, i_10_3892, i_10_3893, i_10_3894, i_10_3895, i_10_3896, i_10_3897, i_10_3898, i_10_3899, i_10_3900, i_10_3901, i_10_3902, i_10_3903, i_10_3904, i_10_3905, i_10_3906, i_10_3907, i_10_3908, i_10_3909, i_10_3910, i_10_3911, i_10_3912, i_10_3913, i_10_3914, i_10_3915, i_10_3916, i_10_3917, i_10_3918, i_10_3919, i_10_3920, i_10_3921, i_10_3922, i_10_3923, i_10_3924, i_10_3925, i_10_3926, i_10_3927, i_10_3928, i_10_3929, i_10_3930, i_10_3931, i_10_3932, i_10_3933, i_10_3934, i_10_3935, i_10_3936, i_10_3937, i_10_3938, i_10_3939, i_10_3940, i_10_3941, i_10_3942, i_10_3943, i_10_3944, i_10_3945, i_10_3946, i_10_3947, i_10_3948, i_10_3949, i_10_3950, i_10_3951, i_10_3952, i_10_3953, i_10_3954, i_10_3955, i_10_3956, i_10_3957, i_10_3958, i_10_3959, i_10_3960, i_10_3961, i_10_3962, i_10_3963, i_10_3964, i_10_3965, i_10_3966, i_10_3967, i_10_3968, i_10_3969, i_10_3970, i_10_3971, i_10_3972, i_10_3973, i_10_3974, i_10_3975, i_10_3976, i_10_3977, i_10_3978, i_10_3979, i_10_3980, i_10_3981, i_10_3982, i_10_3983, i_10_3984, i_10_3985, i_10_3986, i_10_3987, i_10_3988, i_10_3989, i_10_3990, i_10_3991, i_10_3992, i_10_3993, i_10_3994, i_10_3995, i_10_3996, i_10_3997, i_10_3998, i_10_3999, i_10_4000, i_10_4001, i_10_4002, i_10_4003, i_10_4004, i_10_4005, i_10_4006, i_10_4007, i_10_4008, i_10_4009, i_10_4010, i_10_4011, i_10_4012, i_10_4013, i_10_4014, i_10_4015, i_10_4016, i_10_4017, i_10_4018, i_10_4019, i_10_4020, i_10_4021, i_10_4022, i_10_4023, i_10_4024, i_10_4025, i_10_4026, i_10_4027, i_10_4028, i_10_4029, i_10_4030, i_10_4031, i_10_4032, i_10_4033, i_10_4034, i_10_4035, i_10_4036, i_10_4037, i_10_4038, i_10_4039, i_10_4040, i_10_4041, i_10_4042, i_10_4043, i_10_4044, i_10_4045, i_10_4046, i_10_4047, i_10_4048, i_10_4049, i_10_4050, i_10_4051, i_10_4052, i_10_4053, i_10_4054, i_10_4055, i_10_4056, i_10_4057, i_10_4058, i_10_4059, i_10_4060, i_10_4061, i_10_4062, i_10_4063, i_10_4064, i_10_4065, i_10_4066, i_10_4067, i_10_4068, i_10_4069, i_10_4070, i_10_4071, i_10_4072, i_10_4073, i_10_4074, i_10_4075, i_10_4076, i_10_4077, i_10_4078, i_10_4079, i_10_4080, i_10_4081, i_10_4082, i_10_4083, i_10_4084, i_10_4085, i_10_4086, i_10_4087, i_10_4088, i_10_4089, i_10_4090, i_10_4091, i_10_4092, i_10_4093, i_10_4094, i_10_4095, i_10_4096, i_10_4097, i_10_4098, i_10_4099, i_10_4100, i_10_4101, i_10_4102, i_10_4103, i_10_4104, i_10_4105, i_10_4106, i_10_4107, i_10_4108, i_10_4109, i_10_4110, i_10_4111, i_10_4112, i_10_4113, i_10_4114, i_10_4115, i_10_4116, i_10_4117, i_10_4118, i_10_4119, i_10_4120, i_10_4121, i_10_4122, i_10_4123, i_10_4124, i_10_4125, i_10_4126, i_10_4127, i_10_4128, i_10_4129, i_10_4130, i_10_4131, i_10_4132, i_10_4133, i_10_4134, i_10_4135, i_10_4136, i_10_4137, i_10_4138, i_10_4139, i_10_4140, i_10_4141, i_10_4142, i_10_4143, i_10_4144, i_10_4145, i_10_4146, i_10_4147, i_10_4148, i_10_4149, i_10_4150, i_10_4151, i_10_4152, i_10_4153, i_10_4154, i_10_4155, i_10_4156, i_10_4157, i_10_4158, i_10_4159, i_10_4160, i_10_4161, i_10_4162, i_10_4163, i_10_4164, i_10_4165, i_10_4166, i_10_4167, i_10_4168, i_10_4169, i_10_4170, i_10_4171, i_10_4172, i_10_4173, i_10_4174, i_10_4175, i_10_4176, i_10_4177, i_10_4178, i_10_4179, i_10_4180, i_10_4181, i_10_4182, i_10_4183, i_10_4184, i_10_4185, i_10_4186, i_10_4187, i_10_4188, i_10_4189, i_10_4190, i_10_4191, i_10_4192, i_10_4193, i_10_4194, i_10_4195, i_10_4196, i_10_4197, i_10_4198, i_10_4199, i_10_4200, i_10_4201, i_10_4202, i_10_4203, i_10_4204, i_10_4205, i_10_4206, i_10_4207, i_10_4208, i_10_4209, i_10_4210, i_10_4211, i_10_4212, i_10_4213, i_10_4214, i_10_4215, i_10_4216, i_10_4217, i_10_4218, i_10_4219, i_10_4220, i_10_4221, i_10_4222, i_10_4223, i_10_4224, i_10_4225, i_10_4226, i_10_4227, i_10_4228, i_10_4229, i_10_4230, i_10_4231, i_10_4232, i_10_4233, i_10_4234, i_10_4235, i_10_4236, i_10_4237, i_10_4238, i_10_4239, i_10_4240, i_10_4241, i_10_4242, i_10_4243, i_10_4244, i_10_4245, i_10_4246, i_10_4247, i_10_4248, i_10_4249, i_10_4250, i_10_4251, i_10_4252, i_10_4253, i_10_4254, i_10_4255, i_10_4256, i_10_4257, i_10_4258, i_10_4259, i_10_4260, i_10_4261, i_10_4262, i_10_4263, i_10_4264, i_10_4265, i_10_4266, i_10_4267, i_10_4268, i_10_4269, i_10_4270, i_10_4271, i_10_4272, i_10_4273, i_10_4274, i_10_4275, i_10_4276, i_10_4277, i_10_4278, i_10_4279, i_10_4280, i_10_4281, i_10_4282, i_10_4283, i_10_4284, i_10_4285, i_10_4286, i_10_4287, i_10_4288, i_10_4289, i_10_4290, i_10_4291, i_10_4292, i_10_4293, i_10_4294, i_10_4295, i_10_4296, i_10_4297, i_10_4298, i_10_4299, i_10_4300, i_10_4301, i_10_4302, i_10_4303, i_10_4304, i_10_4305, i_10_4306, i_10_4307, i_10_4308, i_10_4309, i_10_4310, i_10_4311, i_10_4312, i_10_4313, i_10_4314, i_10_4315, i_10_4316, i_10_4317, i_10_4318, i_10_4319, i_10_4320, i_10_4321, i_10_4322, i_10_4323, i_10_4324, i_10_4325, i_10_4326, i_10_4327, i_10_4328, i_10_4329, i_10_4330, i_10_4331, i_10_4332, i_10_4333, i_10_4334, i_10_4335, i_10_4336, i_10_4337, i_10_4338, i_10_4339, i_10_4340, i_10_4341, i_10_4342, i_10_4343, i_10_4344, i_10_4345, i_10_4346, i_10_4347, i_10_4348, i_10_4349, i_10_4350, i_10_4351, i_10_4352, i_10_4353, i_10_4354, i_10_4355, i_10_4356, i_10_4357, i_10_4358, i_10_4359, i_10_4360, i_10_4361, i_10_4362, i_10_4363, i_10_4364, i_10_4365, i_10_4366, i_10_4367, i_10_4368, i_10_4369, i_10_4370, i_10_4371, i_10_4372, i_10_4373, i_10_4374, i_10_4375, i_10_4376, i_10_4377, i_10_4378, i_10_4379, i_10_4380, i_10_4381, i_10_4382, i_10_4383, i_10_4384, i_10_4385, i_10_4386, i_10_4387, i_10_4388, i_10_4389, i_10_4390, i_10_4391, i_10_4392, i_10_4393, i_10_4394, i_10_4395, i_10_4396, i_10_4397, i_10_4398, i_10_4399, i_10_4400, i_10_4401, i_10_4402, i_10_4403, i_10_4404, i_10_4405, i_10_4406, i_10_4407, i_10_4408, i_10_4409, i_10_4410, i_10_4411, i_10_4412, i_10_4413, i_10_4414, i_10_4415, i_10_4416, i_10_4417, i_10_4418, i_10_4419, i_10_4420, i_10_4421, i_10_4422, i_10_4423, i_10_4424, i_10_4425, i_10_4426, i_10_4427, i_10_4428, i_10_4429, i_10_4430, i_10_4431, i_10_4432, i_10_4433, i_10_4434, i_10_4435, i_10_4436, i_10_4437, i_10_4438, i_10_4439, i_10_4440, i_10_4441, i_10_4442, i_10_4443, i_10_4444, i_10_4445, i_10_4446, i_10_4447, i_10_4448, i_10_4449, i_10_4450, i_10_4451, i_10_4452, i_10_4453, i_10_4454, i_10_4455, i_10_4456, i_10_4457, i_10_4458, i_10_4459, i_10_4460, i_10_4461, i_10_4462, i_10_4463, i_10_4464, i_10_4465, i_10_4466, i_10_4467, i_10_4468, i_10_4469, i_10_4470, i_10_4471, i_10_4472, i_10_4473, i_10_4474, i_10_4475, i_10_4476, i_10_4477, i_10_4478, i_10_4479, i_10_4480, i_10_4481, i_10_4482, i_10_4483, i_10_4484, i_10_4485, i_10_4486, i_10_4487, i_10_4488, i_10_4489, i_10_4490, i_10_4491, i_10_4492, i_10_4493, i_10_4494, i_10_4495, i_10_4496, i_10_4497, i_10_4498, i_10_4499, i_10_4500, i_10_4501, i_10_4502, i_10_4503, i_10_4504, i_10_4505, i_10_4506, i_10_4507, i_10_4508, i_10_4509, i_10_4510, i_10_4511, i_10_4512, i_10_4513, i_10_4514, i_10_4515, i_10_4516, i_10_4517, i_10_4518, i_10_4519, i_10_4520, i_10_4521, i_10_4522, i_10_4523, i_10_4524, i_10_4525, i_10_4526, i_10_4527, i_10_4528, i_10_4529, i_10_4530, i_10_4531, i_10_4532, i_10_4533, i_10_4534, i_10_4535, i_10_4536, i_10_4537, i_10_4538, i_10_4539, i_10_4540, i_10_4541, i_10_4542, i_10_4543, i_10_4544, i_10_4545, i_10_4546, i_10_4547, i_10_4548, i_10_4549, i_10_4550, i_10_4551, i_10_4552, i_10_4553, i_10_4554, i_10_4555, i_10_4556, i_10_4557, i_10_4558, i_10_4559, i_10_4560, i_10_4561, i_10_4562, i_10_4563, i_10_4564, i_10_4565, i_10_4566, i_10_4567, i_10_4568, i_10_4569, i_10_4570, i_10_4571, i_10_4572, i_10_4573, i_10_4574, i_10_4575, i_10_4576, i_10_4577, i_10_4578, i_10_4579, i_10_4580, i_10_4581, i_10_4582, i_10_4583, i_10_4584, i_10_4585, i_10_4586, i_10_4587, i_10_4588, i_10_4589, i_10_4590, i_10_4591, i_10_4592, i_10_4593, i_10_4594, i_10_4595, i_10_4596, i_10_4597, i_10_4598, i_10_4599, i_10_4600, i_10_4601, i_10_4602, i_10_4603, i_10_4604, i_10_4605, i_10_4606, i_10_4607, o_10_0, o_10_1, o_10_2, o_10_3, o_10_4, o_10_5, o_10_6, o_10_7, o_10_8, o_10_9, o_10_10, o_10_11, o_10_12, o_10_13, o_10_14, o_10_15, o_10_16, o_10_17, o_10_18, o_10_19, o_10_20, o_10_21, o_10_22, o_10_23, o_10_24, o_10_25, o_10_26, o_10_27, o_10_28, o_10_29, o_10_30, o_10_31, o_10_32, o_10_33, o_10_34, o_10_35, o_10_36, o_10_37, o_10_38, o_10_39, o_10_40, o_10_41, o_10_42, o_10_43, o_10_44, o_10_45, o_10_46, o_10_47, o_10_48, o_10_49, o_10_50, o_10_51, o_10_52, o_10_53, o_10_54, o_10_55, o_10_56, o_10_57, o_10_58, o_10_59, o_10_60, o_10_61, o_10_62, o_10_63, o_10_64, o_10_65, o_10_66, o_10_67, o_10_68, o_10_69, o_10_70, o_10_71, o_10_72, o_10_73, o_10_74, o_10_75, o_10_76, o_10_77, o_10_78, o_10_79, o_10_80, o_10_81, o_10_82, o_10_83, o_10_84, o_10_85, o_10_86, o_10_87, o_10_88, o_10_89, o_10_90, o_10_91, o_10_92, o_10_93, o_10_94, o_10_95, o_10_96, o_10_97, o_10_98, o_10_99, o_10_100, o_10_101, o_10_102, o_10_103, o_10_104, o_10_105, o_10_106, o_10_107, o_10_108, o_10_109, o_10_110, o_10_111, o_10_112, o_10_113, o_10_114, o_10_115, o_10_116, o_10_117, o_10_118, o_10_119, o_10_120, o_10_121, o_10_122, o_10_123, o_10_124, o_10_125, o_10_126, o_10_127, o_10_128, o_10_129, o_10_130, o_10_131, o_10_132, o_10_133, o_10_134, o_10_135, o_10_136, o_10_137, o_10_138, o_10_139, o_10_140, o_10_141, o_10_142, o_10_143, o_10_144, o_10_145, o_10_146, o_10_147, o_10_148, o_10_149, o_10_150, o_10_151, o_10_152, o_10_153, o_10_154, o_10_155, o_10_156, o_10_157, o_10_158, o_10_159, o_10_160, o_10_161, o_10_162, o_10_163, o_10_164, o_10_165, o_10_166, o_10_167, o_10_168, o_10_169, o_10_170, o_10_171, o_10_172, o_10_173, o_10_174, o_10_175, o_10_176, o_10_177, o_10_178, o_10_179, o_10_180, o_10_181, o_10_182, o_10_183, o_10_184, o_10_185, o_10_186, o_10_187, o_10_188, o_10_189, o_10_190, o_10_191, o_10_192, o_10_193, o_10_194, o_10_195, o_10_196, o_10_197, o_10_198, o_10_199, o_10_200, o_10_201, o_10_202, o_10_203, o_10_204, o_10_205, o_10_206, o_10_207, o_10_208, o_10_209, o_10_210, o_10_211, o_10_212, o_10_213, o_10_214, o_10_215, o_10_216, o_10_217, o_10_218, o_10_219, o_10_220, o_10_221, o_10_222, o_10_223, o_10_224, o_10_225, o_10_226, o_10_227, o_10_228, o_10_229, o_10_230, o_10_231, o_10_232, o_10_233, o_10_234, o_10_235, o_10_236, o_10_237, o_10_238, o_10_239, o_10_240, o_10_241, o_10_242, o_10_243, o_10_244, o_10_245, o_10_246, o_10_247, o_10_248, o_10_249, o_10_250, o_10_251, o_10_252, o_10_253, o_10_254, o_10_255, o_10_256, o_10_257, o_10_258, o_10_259, o_10_260, o_10_261, o_10_262, o_10_263, o_10_264, o_10_265, o_10_266, o_10_267, o_10_268, o_10_269, o_10_270, o_10_271, o_10_272, o_10_273, o_10_274, o_10_275, o_10_276, o_10_277, o_10_278, o_10_279, o_10_280, o_10_281, o_10_282, o_10_283, o_10_284, o_10_285, o_10_286, o_10_287, o_10_288, o_10_289, o_10_290, o_10_291, o_10_292, o_10_293, o_10_294, o_10_295, o_10_296, o_10_297, o_10_298, o_10_299, o_10_300, o_10_301, o_10_302, o_10_303, o_10_304, o_10_305, o_10_306, o_10_307, o_10_308, o_10_309, o_10_310, o_10_311, o_10_312, o_10_313, o_10_314, o_10_315, o_10_316, o_10_317, o_10_318, o_10_319, o_10_320, o_10_321, o_10_322, o_10_323, o_10_324, o_10_325, o_10_326, o_10_327, o_10_328, o_10_329, o_10_330, o_10_331, o_10_332, o_10_333, o_10_334, o_10_335, o_10_336, o_10_337, o_10_338, o_10_339, o_10_340, o_10_341, o_10_342, o_10_343, o_10_344, o_10_345, o_10_346, o_10_347, o_10_348, o_10_349, o_10_350, o_10_351, o_10_352, o_10_353, o_10_354, o_10_355, o_10_356, o_10_357, o_10_358, o_10_359, o_10_360, o_10_361, o_10_362, o_10_363, o_10_364, o_10_365, o_10_366, o_10_367, o_10_368, o_10_369, o_10_370, o_10_371, o_10_372, o_10_373, o_10_374, o_10_375, o_10_376, o_10_377, o_10_378, o_10_379, o_10_380, o_10_381, o_10_382, o_10_383, o_10_384, o_10_385, o_10_386, o_10_387, o_10_388, o_10_389, o_10_390, o_10_391, o_10_392, o_10_393, o_10_394, o_10_395, o_10_396, o_10_397, o_10_398, o_10_399, o_10_400, o_10_401, o_10_402, o_10_403, o_10_404, o_10_405, o_10_406, o_10_407, o_10_408, o_10_409, o_10_410, o_10_411, o_10_412, o_10_413, o_10_414, o_10_415, o_10_416, o_10_417, o_10_418, o_10_419, o_10_420, o_10_421, o_10_422, o_10_423, o_10_424, o_10_425, o_10_426, o_10_427, o_10_428, o_10_429, o_10_430, o_10_431, o_10_432, o_10_433, o_10_434, o_10_435, o_10_436, o_10_437, o_10_438, o_10_439, o_10_440, o_10_441, o_10_442, o_10_443, o_10_444, o_10_445, o_10_446, o_10_447, o_10_448, o_10_449, o_10_450, o_10_451, o_10_452, o_10_453, o_10_454, o_10_455, o_10_456, o_10_457, o_10_458, o_10_459, o_10_460, o_10_461, o_10_462, o_10_463, o_10_464, o_10_465, o_10_466, o_10_467, o_10_468, o_10_469, o_10_470, o_10_471, o_10_472, o_10_473, o_10_474, o_10_475, o_10_476, o_10_477, o_10_478, o_10_479, o_10_480, o_10_481, o_10_482, o_10_483, o_10_484, o_10_485, o_10_486, o_10_487, o_10_488, o_10_489, o_10_490, o_10_491, o_10_492, o_10_493, o_10_494, o_10_495, o_10_496, o_10_497, o_10_498, o_10_499, o_10_500, o_10_501, o_10_502, o_10_503, o_10_504, o_10_505, o_10_506, o_10_507, o_10_508, o_10_509, o_10_510, o_10_511);
input i_10_0, i_10_1, i_10_2, i_10_3, i_10_4, i_10_5, i_10_6, i_10_7, i_10_8, i_10_9, i_10_10, i_10_11, i_10_12, i_10_13, i_10_14, i_10_15, i_10_16, i_10_17, i_10_18, i_10_19, i_10_20, i_10_21, i_10_22, i_10_23, i_10_24, i_10_25, i_10_26, i_10_27, i_10_28, i_10_29, i_10_30, i_10_31, i_10_32, i_10_33, i_10_34, i_10_35, i_10_36, i_10_37, i_10_38, i_10_39, i_10_40, i_10_41, i_10_42, i_10_43, i_10_44, i_10_45, i_10_46, i_10_47, i_10_48, i_10_49, i_10_50, i_10_51, i_10_52, i_10_53, i_10_54, i_10_55, i_10_56, i_10_57, i_10_58, i_10_59, i_10_60, i_10_61, i_10_62, i_10_63, i_10_64, i_10_65, i_10_66, i_10_67, i_10_68, i_10_69, i_10_70, i_10_71, i_10_72, i_10_73, i_10_74, i_10_75, i_10_76, i_10_77, i_10_78, i_10_79, i_10_80, i_10_81, i_10_82, i_10_83, i_10_84, i_10_85, i_10_86, i_10_87, i_10_88, i_10_89, i_10_90, i_10_91, i_10_92, i_10_93, i_10_94, i_10_95, i_10_96, i_10_97, i_10_98, i_10_99, i_10_100, i_10_101, i_10_102, i_10_103, i_10_104, i_10_105, i_10_106, i_10_107, i_10_108, i_10_109, i_10_110, i_10_111, i_10_112, i_10_113, i_10_114, i_10_115, i_10_116, i_10_117, i_10_118, i_10_119, i_10_120, i_10_121, i_10_122, i_10_123, i_10_124, i_10_125, i_10_126, i_10_127, i_10_128, i_10_129, i_10_130, i_10_131, i_10_132, i_10_133, i_10_134, i_10_135, i_10_136, i_10_137, i_10_138, i_10_139, i_10_140, i_10_141, i_10_142, i_10_143, i_10_144, i_10_145, i_10_146, i_10_147, i_10_148, i_10_149, i_10_150, i_10_151, i_10_152, i_10_153, i_10_154, i_10_155, i_10_156, i_10_157, i_10_158, i_10_159, i_10_160, i_10_161, i_10_162, i_10_163, i_10_164, i_10_165, i_10_166, i_10_167, i_10_168, i_10_169, i_10_170, i_10_171, i_10_172, i_10_173, i_10_174, i_10_175, i_10_176, i_10_177, i_10_178, i_10_179, i_10_180, i_10_181, i_10_182, i_10_183, i_10_184, i_10_185, i_10_186, i_10_187, i_10_188, i_10_189, i_10_190, i_10_191, i_10_192, i_10_193, i_10_194, i_10_195, i_10_196, i_10_197, i_10_198, i_10_199, i_10_200, i_10_201, i_10_202, i_10_203, i_10_204, i_10_205, i_10_206, i_10_207, i_10_208, i_10_209, i_10_210, i_10_211, i_10_212, i_10_213, i_10_214, i_10_215, i_10_216, i_10_217, i_10_218, i_10_219, i_10_220, i_10_221, i_10_222, i_10_223, i_10_224, i_10_225, i_10_226, i_10_227, i_10_228, i_10_229, i_10_230, i_10_231, i_10_232, i_10_233, i_10_234, i_10_235, i_10_236, i_10_237, i_10_238, i_10_239, i_10_240, i_10_241, i_10_242, i_10_243, i_10_244, i_10_245, i_10_246, i_10_247, i_10_248, i_10_249, i_10_250, i_10_251, i_10_252, i_10_253, i_10_254, i_10_255, i_10_256, i_10_257, i_10_258, i_10_259, i_10_260, i_10_261, i_10_262, i_10_263, i_10_264, i_10_265, i_10_266, i_10_267, i_10_268, i_10_269, i_10_270, i_10_271, i_10_272, i_10_273, i_10_274, i_10_275, i_10_276, i_10_277, i_10_278, i_10_279, i_10_280, i_10_281, i_10_282, i_10_283, i_10_284, i_10_285, i_10_286, i_10_287, i_10_288, i_10_289, i_10_290, i_10_291, i_10_292, i_10_293, i_10_294, i_10_295, i_10_296, i_10_297, i_10_298, i_10_299, i_10_300, i_10_301, i_10_302, i_10_303, i_10_304, i_10_305, i_10_306, i_10_307, i_10_308, i_10_309, i_10_310, i_10_311, i_10_312, i_10_313, i_10_314, i_10_315, i_10_316, i_10_317, i_10_318, i_10_319, i_10_320, i_10_321, i_10_322, i_10_323, i_10_324, i_10_325, i_10_326, i_10_327, i_10_328, i_10_329, i_10_330, i_10_331, i_10_332, i_10_333, i_10_334, i_10_335, i_10_336, i_10_337, i_10_338, i_10_339, i_10_340, i_10_341, i_10_342, i_10_343, i_10_344, i_10_345, i_10_346, i_10_347, i_10_348, i_10_349, i_10_350, i_10_351, i_10_352, i_10_353, i_10_354, i_10_355, i_10_356, i_10_357, i_10_358, i_10_359, i_10_360, i_10_361, i_10_362, i_10_363, i_10_364, i_10_365, i_10_366, i_10_367, i_10_368, i_10_369, i_10_370, i_10_371, i_10_372, i_10_373, i_10_374, i_10_375, i_10_376, i_10_377, i_10_378, i_10_379, i_10_380, i_10_381, i_10_382, i_10_383, i_10_384, i_10_385, i_10_386, i_10_387, i_10_388, i_10_389, i_10_390, i_10_391, i_10_392, i_10_393, i_10_394, i_10_395, i_10_396, i_10_397, i_10_398, i_10_399, i_10_400, i_10_401, i_10_402, i_10_403, i_10_404, i_10_405, i_10_406, i_10_407, i_10_408, i_10_409, i_10_410, i_10_411, i_10_412, i_10_413, i_10_414, i_10_415, i_10_416, i_10_417, i_10_418, i_10_419, i_10_420, i_10_421, i_10_422, i_10_423, i_10_424, i_10_425, i_10_426, i_10_427, i_10_428, i_10_429, i_10_430, i_10_431, i_10_432, i_10_433, i_10_434, i_10_435, i_10_436, i_10_437, i_10_438, i_10_439, i_10_440, i_10_441, i_10_442, i_10_443, i_10_444, i_10_445, i_10_446, i_10_447, i_10_448, i_10_449, i_10_450, i_10_451, i_10_452, i_10_453, i_10_454, i_10_455, i_10_456, i_10_457, i_10_458, i_10_459, i_10_460, i_10_461, i_10_462, i_10_463, i_10_464, i_10_465, i_10_466, i_10_467, i_10_468, i_10_469, i_10_470, i_10_471, i_10_472, i_10_473, i_10_474, i_10_475, i_10_476, i_10_477, i_10_478, i_10_479, i_10_480, i_10_481, i_10_482, i_10_483, i_10_484, i_10_485, i_10_486, i_10_487, i_10_488, i_10_489, i_10_490, i_10_491, i_10_492, i_10_493, i_10_494, i_10_495, i_10_496, i_10_497, i_10_498, i_10_499, i_10_500, i_10_501, i_10_502, i_10_503, i_10_504, i_10_505, i_10_506, i_10_507, i_10_508, i_10_509, i_10_510, i_10_511, i_10_512, i_10_513, i_10_514, i_10_515, i_10_516, i_10_517, i_10_518, i_10_519, i_10_520, i_10_521, i_10_522, i_10_523, i_10_524, i_10_525, i_10_526, i_10_527, i_10_528, i_10_529, i_10_530, i_10_531, i_10_532, i_10_533, i_10_534, i_10_535, i_10_536, i_10_537, i_10_538, i_10_539, i_10_540, i_10_541, i_10_542, i_10_543, i_10_544, i_10_545, i_10_546, i_10_547, i_10_548, i_10_549, i_10_550, i_10_551, i_10_552, i_10_553, i_10_554, i_10_555, i_10_556, i_10_557, i_10_558, i_10_559, i_10_560, i_10_561, i_10_562, i_10_563, i_10_564, i_10_565, i_10_566, i_10_567, i_10_568, i_10_569, i_10_570, i_10_571, i_10_572, i_10_573, i_10_574, i_10_575, i_10_576, i_10_577, i_10_578, i_10_579, i_10_580, i_10_581, i_10_582, i_10_583, i_10_584, i_10_585, i_10_586, i_10_587, i_10_588, i_10_589, i_10_590, i_10_591, i_10_592, i_10_593, i_10_594, i_10_595, i_10_596, i_10_597, i_10_598, i_10_599, i_10_600, i_10_601, i_10_602, i_10_603, i_10_604, i_10_605, i_10_606, i_10_607, i_10_608, i_10_609, i_10_610, i_10_611, i_10_612, i_10_613, i_10_614, i_10_615, i_10_616, i_10_617, i_10_618, i_10_619, i_10_620, i_10_621, i_10_622, i_10_623, i_10_624, i_10_625, i_10_626, i_10_627, i_10_628, i_10_629, i_10_630, i_10_631, i_10_632, i_10_633, i_10_634, i_10_635, i_10_636, i_10_637, i_10_638, i_10_639, i_10_640, i_10_641, i_10_642, i_10_643, i_10_644, i_10_645, i_10_646, i_10_647, i_10_648, i_10_649, i_10_650, i_10_651, i_10_652, i_10_653, i_10_654, i_10_655, i_10_656, i_10_657, i_10_658, i_10_659, i_10_660, i_10_661, i_10_662, i_10_663, i_10_664, i_10_665, i_10_666, i_10_667, i_10_668, i_10_669, i_10_670, i_10_671, i_10_672, i_10_673, i_10_674, i_10_675, i_10_676, i_10_677, i_10_678, i_10_679, i_10_680, i_10_681, i_10_682, i_10_683, i_10_684, i_10_685, i_10_686, i_10_687, i_10_688, i_10_689, i_10_690, i_10_691, i_10_692, i_10_693, i_10_694, i_10_695, i_10_696, i_10_697, i_10_698, i_10_699, i_10_700, i_10_701, i_10_702, i_10_703, i_10_704, i_10_705, i_10_706, i_10_707, i_10_708, i_10_709, i_10_710, i_10_711, i_10_712, i_10_713, i_10_714, i_10_715, i_10_716, i_10_717, i_10_718, i_10_719, i_10_720, i_10_721, i_10_722, i_10_723, i_10_724, i_10_725, i_10_726, i_10_727, i_10_728, i_10_729, i_10_730, i_10_731, i_10_732, i_10_733, i_10_734, i_10_735, i_10_736, i_10_737, i_10_738, i_10_739, i_10_740, i_10_741, i_10_742, i_10_743, i_10_744, i_10_745, i_10_746, i_10_747, i_10_748, i_10_749, i_10_750, i_10_751, i_10_752, i_10_753, i_10_754, i_10_755, i_10_756, i_10_757, i_10_758, i_10_759, i_10_760, i_10_761, i_10_762, i_10_763, i_10_764, i_10_765, i_10_766, i_10_767, i_10_768, i_10_769, i_10_770, i_10_771, i_10_772, i_10_773, i_10_774, i_10_775, i_10_776, i_10_777, i_10_778, i_10_779, i_10_780, i_10_781, i_10_782, i_10_783, i_10_784, i_10_785, i_10_786, i_10_787, i_10_788, i_10_789, i_10_790, i_10_791, i_10_792, i_10_793, i_10_794, i_10_795, i_10_796, i_10_797, i_10_798, i_10_799, i_10_800, i_10_801, i_10_802, i_10_803, i_10_804, i_10_805, i_10_806, i_10_807, i_10_808, i_10_809, i_10_810, i_10_811, i_10_812, i_10_813, i_10_814, i_10_815, i_10_816, i_10_817, i_10_818, i_10_819, i_10_820, i_10_821, i_10_822, i_10_823, i_10_824, i_10_825, i_10_826, i_10_827, i_10_828, i_10_829, i_10_830, i_10_831, i_10_832, i_10_833, i_10_834, i_10_835, i_10_836, i_10_837, i_10_838, i_10_839, i_10_840, i_10_841, i_10_842, i_10_843, i_10_844, i_10_845, i_10_846, i_10_847, i_10_848, i_10_849, i_10_850, i_10_851, i_10_852, i_10_853, i_10_854, i_10_855, i_10_856, i_10_857, i_10_858, i_10_859, i_10_860, i_10_861, i_10_862, i_10_863, i_10_864, i_10_865, i_10_866, i_10_867, i_10_868, i_10_869, i_10_870, i_10_871, i_10_872, i_10_873, i_10_874, i_10_875, i_10_876, i_10_877, i_10_878, i_10_879, i_10_880, i_10_881, i_10_882, i_10_883, i_10_884, i_10_885, i_10_886, i_10_887, i_10_888, i_10_889, i_10_890, i_10_891, i_10_892, i_10_893, i_10_894, i_10_895, i_10_896, i_10_897, i_10_898, i_10_899, i_10_900, i_10_901, i_10_902, i_10_903, i_10_904, i_10_905, i_10_906, i_10_907, i_10_908, i_10_909, i_10_910, i_10_911, i_10_912, i_10_913, i_10_914, i_10_915, i_10_916, i_10_917, i_10_918, i_10_919, i_10_920, i_10_921, i_10_922, i_10_923, i_10_924, i_10_925, i_10_926, i_10_927, i_10_928, i_10_929, i_10_930, i_10_931, i_10_932, i_10_933, i_10_934, i_10_935, i_10_936, i_10_937, i_10_938, i_10_939, i_10_940, i_10_941, i_10_942, i_10_943, i_10_944, i_10_945, i_10_946, i_10_947, i_10_948, i_10_949, i_10_950, i_10_951, i_10_952, i_10_953, i_10_954, i_10_955, i_10_956, i_10_957, i_10_958, i_10_959, i_10_960, i_10_961, i_10_962, i_10_963, i_10_964, i_10_965, i_10_966, i_10_967, i_10_968, i_10_969, i_10_970, i_10_971, i_10_972, i_10_973, i_10_974, i_10_975, i_10_976, i_10_977, i_10_978, i_10_979, i_10_980, i_10_981, i_10_982, i_10_983, i_10_984, i_10_985, i_10_986, i_10_987, i_10_988, i_10_989, i_10_990, i_10_991, i_10_992, i_10_993, i_10_994, i_10_995, i_10_996, i_10_997, i_10_998, i_10_999, i_10_1000, i_10_1001, i_10_1002, i_10_1003, i_10_1004, i_10_1005, i_10_1006, i_10_1007, i_10_1008, i_10_1009, i_10_1010, i_10_1011, i_10_1012, i_10_1013, i_10_1014, i_10_1015, i_10_1016, i_10_1017, i_10_1018, i_10_1019, i_10_1020, i_10_1021, i_10_1022, i_10_1023, i_10_1024, i_10_1025, i_10_1026, i_10_1027, i_10_1028, i_10_1029, i_10_1030, i_10_1031, i_10_1032, i_10_1033, i_10_1034, i_10_1035, i_10_1036, i_10_1037, i_10_1038, i_10_1039, i_10_1040, i_10_1041, i_10_1042, i_10_1043, i_10_1044, i_10_1045, i_10_1046, i_10_1047, i_10_1048, i_10_1049, i_10_1050, i_10_1051, i_10_1052, i_10_1053, i_10_1054, i_10_1055, i_10_1056, i_10_1057, i_10_1058, i_10_1059, i_10_1060, i_10_1061, i_10_1062, i_10_1063, i_10_1064, i_10_1065, i_10_1066, i_10_1067, i_10_1068, i_10_1069, i_10_1070, i_10_1071, i_10_1072, i_10_1073, i_10_1074, i_10_1075, i_10_1076, i_10_1077, i_10_1078, i_10_1079, i_10_1080, i_10_1081, i_10_1082, i_10_1083, i_10_1084, i_10_1085, i_10_1086, i_10_1087, i_10_1088, i_10_1089, i_10_1090, i_10_1091, i_10_1092, i_10_1093, i_10_1094, i_10_1095, i_10_1096, i_10_1097, i_10_1098, i_10_1099, i_10_1100, i_10_1101, i_10_1102, i_10_1103, i_10_1104, i_10_1105, i_10_1106, i_10_1107, i_10_1108, i_10_1109, i_10_1110, i_10_1111, i_10_1112, i_10_1113, i_10_1114, i_10_1115, i_10_1116, i_10_1117, i_10_1118, i_10_1119, i_10_1120, i_10_1121, i_10_1122, i_10_1123, i_10_1124, i_10_1125, i_10_1126, i_10_1127, i_10_1128, i_10_1129, i_10_1130, i_10_1131, i_10_1132, i_10_1133, i_10_1134, i_10_1135, i_10_1136, i_10_1137, i_10_1138, i_10_1139, i_10_1140, i_10_1141, i_10_1142, i_10_1143, i_10_1144, i_10_1145, i_10_1146, i_10_1147, i_10_1148, i_10_1149, i_10_1150, i_10_1151, i_10_1152, i_10_1153, i_10_1154, i_10_1155, i_10_1156, i_10_1157, i_10_1158, i_10_1159, i_10_1160, i_10_1161, i_10_1162, i_10_1163, i_10_1164, i_10_1165, i_10_1166, i_10_1167, i_10_1168, i_10_1169, i_10_1170, i_10_1171, i_10_1172, i_10_1173, i_10_1174, i_10_1175, i_10_1176, i_10_1177, i_10_1178, i_10_1179, i_10_1180, i_10_1181, i_10_1182, i_10_1183, i_10_1184, i_10_1185, i_10_1186, i_10_1187, i_10_1188, i_10_1189, i_10_1190, i_10_1191, i_10_1192, i_10_1193, i_10_1194, i_10_1195, i_10_1196, i_10_1197, i_10_1198, i_10_1199, i_10_1200, i_10_1201, i_10_1202, i_10_1203, i_10_1204, i_10_1205, i_10_1206, i_10_1207, i_10_1208, i_10_1209, i_10_1210, i_10_1211, i_10_1212, i_10_1213, i_10_1214, i_10_1215, i_10_1216, i_10_1217, i_10_1218, i_10_1219, i_10_1220, i_10_1221, i_10_1222, i_10_1223, i_10_1224, i_10_1225, i_10_1226, i_10_1227, i_10_1228, i_10_1229, i_10_1230, i_10_1231, i_10_1232, i_10_1233, i_10_1234, i_10_1235, i_10_1236, i_10_1237, i_10_1238, i_10_1239, i_10_1240, i_10_1241, i_10_1242, i_10_1243, i_10_1244, i_10_1245, i_10_1246, i_10_1247, i_10_1248, i_10_1249, i_10_1250, i_10_1251, i_10_1252, i_10_1253, i_10_1254, i_10_1255, i_10_1256, i_10_1257, i_10_1258, i_10_1259, i_10_1260, i_10_1261, i_10_1262, i_10_1263, i_10_1264, i_10_1265, i_10_1266, i_10_1267, i_10_1268, i_10_1269, i_10_1270, i_10_1271, i_10_1272, i_10_1273, i_10_1274, i_10_1275, i_10_1276, i_10_1277, i_10_1278, i_10_1279, i_10_1280, i_10_1281, i_10_1282, i_10_1283, i_10_1284, i_10_1285, i_10_1286, i_10_1287, i_10_1288, i_10_1289, i_10_1290, i_10_1291, i_10_1292, i_10_1293, i_10_1294, i_10_1295, i_10_1296, i_10_1297, i_10_1298, i_10_1299, i_10_1300, i_10_1301, i_10_1302, i_10_1303, i_10_1304, i_10_1305, i_10_1306, i_10_1307, i_10_1308, i_10_1309, i_10_1310, i_10_1311, i_10_1312, i_10_1313, i_10_1314, i_10_1315, i_10_1316, i_10_1317, i_10_1318, i_10_1319, i_10_1320, i_10_1321, i_10_1322, i_10_1323, i_10_1324, i_10_1325, i_10_1326, i_10_1327, i_10_1328, i_10_1329, i_10_1330, i_10_1331, i_10_1332, i_10_1333, i_10_1334, i_10_1335, i_10_1336, i_10_1337, i_10_1338, i_10_1339, i_10_1340, i_10_1341, i_10_1342, i_10_1343, i_10_1344, i_10_1345, i_10_1346, i_10_1347, i_10_1348, i_10_1349, i_10_1350, i_10_1351, i_10_1352, i_10_1353, i_10_1354, i_10_1355, i_10_1356, i_10_1357, i_10_1358, i_10_1359, i_10_1360, i_10_1361, i_10_1362, i_10_1363, i_10_1364, i_10_1365, i_10_1366, i_10_1367, i_10_1368, i_10_1369, i_10_1370, i_10_1371, i_10_1372, i_10_1373, i_10_1374, i_10_1375, i_10_1376, i_10_1377, i_10_1378, i_10_1379, i_10_1380, i_10_1381, i_10_1382, i_10_1383, i_10_1384, i_10_1385, i_10_1386, i_10_1387, i_10_1388, i_10_1389, i_10_1390, i_10_1391, i_10_1392, i_10_1393, i_10_1394, i_10_1395, i_10_1396, i_10_1397, i_10_1398, i_10_1399, i_10_1400, i_10_1401, i_10_1402, i_10_1403, i_10_1404, i_10_1405, i_10_1406, i_10_1407, i_10_1408, i_10_1409, i_10_1410, i_10_1411, i_10_1412, i_10_1413, i_10_1414, i_10_1415, i_10_1416, i_10_1417, i_10_1418, i_10_1419, i_10_1420, i_10_1421, i_10_1422, i_10_1423, i_10_1424, i_10_1425, i_10_1426, i_10_1427, i_10_1428, i_10_1429, i_10_1430, i_10_1431, i_10_1432, i_10_1433, i_10_1434, i_10_1435, i_10_1436, i_10_1437, i_10_1438, i_10_1439, i_10_1440, i_10_1441, i_10_1442, i_10_1443, i_10_1444, i_10_1445, i_10_1446, i_10_1447, i_10_1448, i_10_1449, i_10_1450, i_10_1451, i_10_1452, i_10_1453, i_10_1454, i_10_1455, i_10_1456, i_10_1457, i_10_1458, i_10_1459, i_10_1460, i_10_1461, i_10_1462, i_10_1463, i_10_1464, i_10_1465, i_10_1466, i_10_1467, i_10_1468, i_10_1469, i_10_1470, i_10_1471, i_10_1472, i_10_1473, i_10_1474, i_10_1475, i_10_1476, i_10_1477, i_10_1478, i_10_1479, i_10_1480, i_10_1481, i_10_1482, i_10_1483, i_10_1484, i_10_1485, i_10_1486, i_10_1487, i_10_1488, i_10_1489, i_10_1490, i_10_1491, i_10_1492, i_10_1493, i_10_1494, i_10_1495, i_10_1496, i_10_1497, i_10_1498, i_10_1499, i_10_1500, i_10_1501, i_10_1502, i_10_1503, i_10_1504, i_10_1505, i_10_1506, i_10_1507, i_10_1508, i_10_1509, i_10_1510, i_10_1511, i_10_1512, i_10_1513, i_10_1514, i_10_1515, i_10_1516, i_10_1517, i_10_1518, i_10_1519, i_10_1520, i_10_1521, i_10_1522, i_10_1523, i_10_1524, i_10_1525, i_10_1526, i_10_1527, i_10_1528, i_10_1529, i_10_1530, i_10_1531, i_10_1532, i_10_1533, i_10_1534, i_10_1535, i_10_1536, i_10_1537, i_10_1538, i_10_1539, i_10_1540, i_10_1541, i_10_1542, i_10_1543, i_10_1544, i_10_1545, i_10_1546, i_10_1547, i_10_1548, i_10_1549, i_10_1550, i_10_1551, i_10_1552, i_10_1553, i_10_1554, i_10_1555, i_10_1556, i_10_1557, i_10_1558, i_10_1559, i_10_1560, i_10_1561, i_10_1562, i_10_1563, i_10_1564, i_10_1565, i_10_1566, i_10_1567, i_10_1568, i_10_1569, i_10_1570, i_10_1571, i_10_1572, i_10_1573, i_10_1574, i_10_1575, i_10_1576, i_10_1577, i_10_1578, i_10_1579, i_10_1580, i_10_1581, i_10_1582, i_10_1583, i_10_1584, i_10_1585, i_10_1586, i_10_1587, i_10_1588, i_10_1589, i_10_1590, i_10_1591, i_10_1592, i_10_1593, i_10_1594, i_10_1595, i_10_1596, i_10_1597, i_10_1598, i_10_1599, i_10_1600, i_10_1601, i_10_1602, i_10_1603, i_10_1604, i_10_1605, i_10_1606, i_10_1607, i_10_1608, i_10_1609, i_10_1610, i_10_1611, i_10_1612, i_10_1613, i_10_1614, i_10_1615, i_10_1616, i_10_1617, i_10_1618, i_10_1619, i_10_1620, i_10_1621, i_10_1622, i_10_1623, i_10_1624, i_10_1625, i_10_1626, i_10_1627, i_10_1628, i_10_1629, i_10_1630, i_10_1631, i_10_1632, i_10_1633, i_10_1634, i_10_1635, i_10_1636, i_10_1637, i_10_1638, i_10_1639, i_10_1640, i_10_1641, i_10_1642, i_10_1643, i_10_1644, i_10_1645, i_10_1646, i_10_1647, i_10_1648, i_10_1649, i_10_1650, i_10_1651, i_10_1652, i_10_1653, i_10_1654, i_10_1655, i_10_1656, i_10_1657, i_10_1658, i_10_1659, i_10_1660, i_10_1661, i_10_1662, i_10_1663, i_10_1664, i_10_1665, i_10_1666, i_10_1667, i_10_1668, i_10_1669, i_10_1670, i_10_1671, i_10_1672, i_10_1673, i_10_1674, i_10_1675, i_10_1676, i_10_1677, i_10_1678, i_10_1679, i_10_1680, i_10_1681, i_10_1682, i_10_1683, i_10_1684, i_10_1685, i_10_1686, i_10_1687, i_10_1688, i_10_1689, i_10_1690, i_10_1691, i_10_1692, i_10_1693, i_10_1694, i_10_1695, i_10_1696, i_10_1697, i_10_1698, i_10_1699, i_10_1700, i_10_1701, i_10_1702, i_10_1703, i_10_1704, i_10_1705, i_10_1706, i_10_1707, i_10_1708, i_10_1709, i_10_1710, i_10_1711, i_10_1712, i_10_1713, i_10_1714, i_10_1715, i_10_1716, i_10_1717, i_10_1718, i_10_1719, i_10_1720, i_10_1721, i_10_1722, i_10_1723, i_10_1724, i_10_1725, i_10_1726, i_10_1727, i_10_1728, i_10_1729, i_10_1730, i_10_1731, i_10_1732, i_10_1733, i_10_1734, i_10_1735, i_10_1736, i_10_1737, i_10_1738, i_10_1739, i_10_1740, i_10_1741, i_10_1742, i_10_1743, i_10_1744, i_10_1745, i_10_1746, i_10_1747, i_10_1748, i_10_1749, i_10_1750, i_10_1751, i_10_1752, i_10_1753, i_10_1754, i_10_1755, i_10_1756, i_10_1757, i_10_1758, i_10_1759, i_10_1760, i_10_1761, i_10_1762, i_10_1763, i_10_1764, i_10_1765, i_10_1766, i_10_1767, i_10_1768, i_10_1769, i_10_1770, i_10_1771, i_10_1772, i_10_1773, i_10_1774, i_10_1775, i_10_1776, i_10_1777, i_10_1778, i_10_1779, i_10_1780, i_10_1781, i_10_1782, i_10_1783, i_10_1784, i_10_1785, i_10_1786, i_10_1787, i_10_1788, i_10_1789, i_10_1790, i_10_1791, i_10_1792, i_10_1793, i_10_1794, i_10_1795, i_10_1796, i_10_1797, i_10_1798, i_10_1799, i_10_1800, i_10_1801, i_10_1802, i_10_1803, i_10_1804, i_10_1805, i_10_1806, i_10_1807, i_10_1808, i_10_1809, i_10_1810, i_10_1811, i_10_1812, i_10_1813, i_10_1814, i_10_1815, i_10_1816, i_10_1817, i_10_1818, i_10_1819, i_10_1820, i_10_1821, i_10_1822, i_10_1823, i_10_1824, i_10_1825, i_10_1826, i_10_1827, i_10_1828, i_10_1829, i_10_1830, i_10_1831, i_10_1832, i_10_1833, i_10_1834, i_10_1835, i_10_1836, i_10_1837, i_10_1838, i_10_1839, i_10_1840, i_10_1841, i_10_1842, i_10_1843, i_10_1844, i_10_1845, i_10_1846, i_10_1847, i_10_1848, i_10_1849, i_10_1850, i_10_1851, i_10_1852, i_10_1853, i_10_1854, i_10_1855, i_10_1856, i_10_1857, i_10_1858, i_10_1859, i_10_1860, i_10_1861, i_10_1862, i_10_1863, i_10_1864, i_10_1865, i_10_1866, i_10_1867, i_10_1868, i_10_1869, i_10_1870, i_10_1871, i_10_1872, i_10_1873, i_10_1874, i_10_1875, i_10_1876, i_10_1877, i_10_1878, i_10_1879, i_10_1880, i_10_1881, i_10_1882, i_10_1883, i_10_1884, i_10_1885, i_10_1886, i_10_1887, i_10_1888, i_10_1889, i_10_1890, i_10_1891, i_10_1892, i_10_1893, i_10_1894, i_10_1895, i_10_1896, i_10_1897, i_10_1898, i_10_1899, i_10_1900, i_10_1901, i_10_1902, i_10_1903, i_10_1904, i_10_1905, i_10_1906, i_10_1907, i_10_1908, i_10_1909, i_10_1910, i_10_1911, i_10_1912, i_10_1913, i_10_1914, i_10_1915, i_10_1916, i_10_1917, i_10_1918, i_10_1919, i_10_1920, i_10_1921, i_10_1922, i_10_1923, i_10_1924, i_10_1925, i_10_1926, i_10_1927, i_10_1928, i_10_1929, i_10_1930, i_10_1931, i_10_1932, i_10_1933, i_10_1934, i_10_1935, i_10_1936, i_10_1937, i_10_1938, i_10_1939, i_10_1940, i_10_1941, i_10_1942, i_10_1943, i_10_1944, i_10_1945, i_10_1946, i_10_1947, i_10_1948, i_10_1949, i_10_1950, i_10_1951, i_10_1952, i_10_1953, i_10_1954, i_10_1955, i_10_1956, i_10_1957, i_10_1958, i_10_1959, i_10_1960, i_10_1961, i_10_1962, i_10_1963, i_10_1964, i_10_1965, i_10_1966, i_10_1967, i_10_1968, i_10_1969, i_10_1970, i_10_1971, i_10_1972, i_10_1973, i_10_1974, i_10_1975, i_10_1976, i_10_1977, i_10_1978, i_10_1979, i_10_1980, i_10_1981, i_10_1982, i_10_1983, i_10_1984, i_10_1985, i_10_1986, i_10_1987, i_10_1988, i_10_1989, i_10_1990, i_10_1991, i_10_1992, i_10_1993, i_10_1994, i_10_1995, i_10_1996, i_10_1997, i_10_1998, i_10_1999, i_10_2000, i_10_2001, i_10_2002, i_10_2003, i_10_2004, i_10_2005, i_10_2006, i_10_2007, i_10_2008, i_10_2009, i_10_2010, i_10_2011, i_10_2012, i_10_2013, i_10_2014, i_10_2015, i_10_2016, i_10_2017, i_10_2018, i_10_2019, i_10_2020, i_10_2021, i_10_2022, i_10_2023, i_10_2024, i_10_2025, i_10_2026, i_10_2027, i_10_2028, i_10_2029, i_10_2030, i_10_2031, i_10_2032, i_10_2033, i_10_2034, i_10_2035, i_10_2036, i_10_2037, i_10_2038, i_10_2039, i_10_2040, i_10_2041, i_10_2042, i_10_2043, i_10_2044, i_10_2045, i_10_2046, i_10_2047, i_10_2048, i_10_2049, i_10_2050, i_10_2051, i_10_2052, i_10_2053, i_10_2054, i_10_2055, i_10_2056, i_10_2057, i_10_2058, i_10_2059, i_10_2060, i_10_2061, i_10_2062, i_10_2063, i_10_2064, i_10_2065, i_10_2066, i_10_2067, i_10_2068, i_10_2069, i_10_2070, i_10_2071, i_10_2072, i_10_2073, i_10_2074, i_10_2075, i_10_2076, i_10_2077, i_10_2078, i_10_2079, i_10_2080, i_10_2081, i_10_2082, i_10_2083, i_10_2084, i_10_2085, i_10_2086, i_10_2087, i_10_2088, i_10_2089, i_10_2090, i_10_2091, i_10_2092, i_10_2093, i_10_2094, i_10_2095, i_10_2096, i_10_2097, i_10_2098, i_10_2099, i_10_2100, i_10_2101, i_10_2102, i_10_2103, i_10_2104, i_10_2105, i_10_2106, i_10_2107, i_10_2108, i_10_2109, i_10_2110, i_10_2111, i_10_2112, i_10_2113, i_10_2114, i_10_2115, i_10_2116, i_10_2117, i_10_2118, i_10_2119, i_10_2120, i_10_2121, i_10_2122, i_10_2123, i_10_2124, i_10_2125, i_10_2126, i_10_2127, i_10_2128, i_10_2129, i_10_2130, i_10_2131, i_10_2132, i_10_2133, i_10_2134, i_10_2135, i_10_2136, i_10_2137, i_10_2138, i_10_2139, i_10_2140, i_10_2141, i_10_2142, i_10_2143, i_10_2144, i_10_2145, i_10_2146, i_10_2147, i_10_2148, i_10_2149, i_10_2150, i_10_2151, i_10_2152, i_10_2153, i_10_2154, i_10_2155, i_10_2156, i_10_2157, i_10_2158, i_10_2159, i_10_2160, i_10_2161, i_10_2162, i_10_2163, i_10_2164, i_10_2165, i_10_2166, i_10_2167, i_10_2168, i_10_2169, i_10_2170, i_10_2171, i_10_2172, i_10_2173, i_10_2174, i_10_2175, i_10_2176, i_10_2177, i_10_2178, i_10_2179, i_10_2180, i_10_2181, i_10_2182, i_10_2183, i_10_2184, i_10_2185, i_10_2186, i_10_2187, i_10_2188, i_10_2189, i_10_2190, i_10_2191, i_10_2192, i_10_2193, i_10_2194, i_10_2195, i_10_2196, i_10_2197, i_10_2198, i_10_2199, i_10_2200, i_10_2201, i_10_2202, i_10_2203, i_10_2204, i_10_2205, i_10_2206, i_10_2207, i_10_2208, i_10_2209, i_10_2210, i_10_2211, i_10_2212, i_10_2213, i_10_2214, i_10_2215, i_10_2216, i_10_2217, i_10_2218, i_10_2219, i_10_2220, i_10_2221, i_10_2222, i_10_2223, i_10_2224, i_10_2225, i_10_2226, i_10_2227, i_10_2228, i_10_2229, i_10_2230, i_10_2231, i_10_2232, i_10_2233, i_10_2234, i_10_2235, i_10_2236, i_10_2237, i_10_2238, i_10_2239, i_10_2240, i_10_2241, i_10_2242, i_10_2243, i_10_2244, i_10_2245, i_10_2246, i_10_2247, i_10_2248, i_10_2249, i_10_2250, i_10_2251, i_10_2252, i_10_2253, i_10_2254, i_10_2255, i_10_2256, i_10_2257, i_10_2258, i_10_2259, i_10_2260, i_10_2261, i_10_2262, i_10_2263, i_10_2264, i_10_2265, i_10_2266, i_10_2267, i_10_2268, i_10_2269, i_10_2270, i_10_2271, i_10_2272, i_10_2273, i_10_2274, i_10_2275, i_10_2276, i_10_2277, i_10_2278, i_10_2279, i_10_2280, i_10_2281, i_10_2282, i_10_2283, i_10_2284, i_10_2285, i_10_2286, i_10_2287, i_10_2288, i_10_2289, i_10_2290, i_10_2291, i_10_2292, i_10_2293, i_10_2294, i_10_2295, i_10_2296, i_10_2297, i_10_2298, i_10_2299, i_10_2300, i_10_2301, i_10_2302, i_10_2303, i_10_2304, i_10_2305, i_10_2306, i_10_2307, i_10_2308, i_10_2309, i_10_2310, i_10_2311, i_10_2312, i_10_2313, i_10_2314, i_10_2315, i_10_2316, i_10_2317, i_10_2318, i_10_2319, i_10_2320, i_10_2321, i_10_2322, i_10_2323, i_10_2324, i_10_2325, i_10_2326, i_10_2327, i_10_2328, i_10_2329, i_10_2330, i_10_2331, i_10_2332, i_10_2333, i_10_2334, i_10_2335, i_10_2336, i_10_2337, i_10_2338, i_10_2339, i_10_2340, i_10_2341, i_10_2342, i_10_2343, i_10_2344, i_10_2345, i_10_2346, i_10_2347, i_10_2348, i_10_2349, i_10_2350, i_10_2351, i_10_2352, i_10_2353, i_10_2354, i_10_2355, i_10_2356, i_10_2357, i_10_2358, i_10_2359, i_10_2360, i_10_2361, i_10_2362, i_10_2363, i_10_2364, i_10_2365, i_10_2366, i_10_2367, i_10_2368, i_10_2369, i_10_2370, i_10_2371, i_10_2372, i_10_2373, i_10_2374, i_10_2375, i_10_2376, i_10_2377, i_10_2378, i_10_2379, i_10_2380, i_10_2381, i_10_2382, i_10_2383, i_10_2384, i_10_2385, i_10_2386, i_10_2387, i_10_2388, i_10_2389, i_10_2390, i_10_2391, i_10_2392, i_10_2393, i_10_2394, i_10_2395, i_10_2396, i_10_2397, i_10_2398, i_10_2399, i_10_2400, i_10_2401, i_10_2402, i_10_2403, i_10_2404, i_10_2405, i_10_2406, i_10_2407, i_10_2408, i_10_2409, i_10_2410, i_10_2411, i_10_2412, i_10_2413, i_10_2414, i_10_2415, i_10_2416, i_10_2417, i_10_2418, i_10_2419, i_10_2420, i_10_2421, i_10_2422, i_10_2423, i_10_2424, i_10_2425, i_10_2426, i_10_2427, i_10_2428, i_10_2429, i_10_2430, i_10_2431, i_10_2432, i_10_2433, i_10_2434, i_10_2435, i_10_2436, i_10_2437, i_10_2438, i_10_2439, i_10_2440, i_10_2441, i_10_2442, i_10_2443, i_10_2444, i_10_2445, i_10_2446, i_10_2447, i_10_2448, i_10_2449, i_10_2450, i_10_2451, i_10_2452, i_10_2453, i_10_2454, i_10_2455, i_10_2456, i_10_2457, i_10_2458, i_10_2459, i_10_2460, i_10_2461, i_10_2462, i_10_2463, i_10_2464, i_10_2465, i_10_2466, i_10_2467, i_10_2468, i_10_2469, i_10_2470, i_10_2471, i_10_2472, i_10_2473, i_10_2474, i_10_2475, i_10_2476, i_10_2477, i_10_2478, i_10_2479, i_10_2480, i_10_2481, i_10_2482, i_10_2483, i_10_2484, i_10_2485, i_10_2486, i_10_2487, i_10_2488, i_10_2489, i_10_2490, i_10_2491, i_10_2492, i_10_2493, i_10_2494, i_10_2495, i_10_2496, i_10_2497, i_10_2498, i_10_2499, i_10_2500, i_10_2501, i_10_2502, i_10_2503, i_10_2504, i_10_2505, i_10_2506, i_10_2507, i_10_2508, i_10_2509, i_10_2510, i_10_2511, i_10_2512, i_10_2513, i_10_2514, i_10_2515, i_10_2516, i_10_2517, i_10_2518, i_10_2519, i_10_2520, i_10_2521, i_10_2522, i_10_2523, i_10_2524, i_10_2525, i_10_2526, i_10_2527, i_10_2528, i_10_2529, i_10_2530, i_10_2531, i_10_2532, i_10_2533, i_10_2534, i_10_2535, i_10_2536, i_10_2537, i_10_2538, i_10_2539, i_10_2540, i_10_2541, i_10_2542, i_10_2543, i_10_2544, i_10_2545, i_10_2546, i_10_2547, i_10_2548, i_10_2549, i_10_2550, i_10_2551, i_10_2552, i_10_2553, i_10_2554, i_10_2555, i_10_2556, i_10_2557, i_10_2558, i_10_2559, i_10_2560, i_10_2561, i_10_2562, i_10_2563, i_10_2564, i_10_2565, i_10_2566, i_10_2567, i_10_2568, i_10_2569, i_10_2570, i_10_2571, i_10_2572, i_10_2573, i_10_2574, i_10_2575, i_10_2576, i_10_2577, i_10_2578, i_10_2579, i_10_2580, i_10_2581, i_10_2582, i_10_2583, i_10_2584, i_10_2585, i_10_2586, i_10_2587, i_10_2588, i_10_2589, i_10_2590, i_10_2591, i_10_2592, i_10_2593, i_10_2594, i_10_2595, i_10_2596, i_10_2597, i_10_2598, i_10_2599, i_10_2600, i_10_2601, i_10_2602, i_10_2603, i_10_2604, i_10_2605, i_10_2606, i_10_2607, i_10_2608, i_10_2609, i_10_2610, i_10_2611, i_10_2612, i_10_2613, i_10_2614, i_10_2615, i_10_2616, i_10_2617, i_10_2618, i_10_2619, i_10_2620, i_10_2621, i_10_2622, i_10_2623, i_10_2624, i_10_2625, i_10_2626, i_10_2627, i_10_2628, i_10_2629, i_10_2630, i_10_2631, i_10_2632, i_10_2633, i_10_2634, i_10_2635, i_10_2636, i_10_2637, i_10_2638, i_10_2639, i_10_2640, i_10_2641, i_10_2642, i_10_2643, i_10_2644, i_10_2645, i_10_2646, i_10_2647, i_10_2648, i_10_2649, i_10_2650, i_10_2651, i_10_2652, i_10_2653, i_10_2654, i_10_2655, i_10_2656, i_10_2657, i_10_2658, i_10_2659, i_10_2660, i_10_2661, i_10_2662, i_10_2663, i_10_2664, i_10_2665, i_10_2666, i_10_2667, i_10_2668, i_10_2669, i_10_2670, i_10_2671, i_10_2672, i_10_2673, i_10_2674, i_10_2675, i_10_2676, i_10_2677, i_10_2678, i_10_2679, i_10_2680, i_10_2681, i_10_2682, i_10_2683, i_10_2684, i_10_2685, i_10_2686, i_10_2687, i_10_2688, i_10_2689, i_10_2690, i_10_2691, i_10_2692, i_10_2693, i_10_2694, i_10_2695, i_10_2696, i_10_2697, i_10_2698, i_10_2699, i_10_2700, i_10_2701, i_10_2702, i_10_2703, i_10_2704, i_10_2705, i_10_2706, i_10_2707, i_10_2708, i_10_2709, i_10_2710, i_10_2711, i_10_2712, i_10_2713, i_10_2714, i_10_2715, i_10_2716, i_10_2717, i_10_2718, i_10_2719, i_10_2720, i_10_2721, i_10_2722, i_10_2723, i_10_2724, i_10_2725, i_10_2726, i_10_2727, i_10_2728, i_10_2729, i_10_2730, i_10_2731, i_10_2732, i_10_2733, i_10_2734, i_10_2735, i_10_2736, i_10_2737, i_10_2738, i_10_2739, i_10_2740, i_10_2741, i_10_2742, i_10_2743, i_10_2744, i_10_2745, i_10_2746, i_10_2747, i_10_2748, i_10_2749, i_10_2750, i_10_2751, i_10_2752, i_10_2753, i_10_2754, i_10_2755, i_10_2756, i_10_2757, i_10_2758, i_10_2759, i_10_2760, i_10_2761, i_10_2762, i_10_2763, i_10_2764, i_10_2765, i_10_2766, i_10_2767, i_10_2768, i_10_2769, i_10_2770, i_10_2771, i_10_2772, i_10_2773, i_10_2774, i_10_2775, i_10_2776, i_10_2777, i_10_2778, i_10_2779, i_10_2780, i_10_2781, i_10_2782, i_10_2783, i_10_2784, i_10_2785, i_10_2786, i_10_2787, i_10_2788, i_10_2789, i_10_2790, i_10_2791, i_10_2792, i_10_2793, i_10_2794, i_10_2795, i_10_2796, i_10_2797, i_10_2798, i_10_2799, i_10_2800, i_10_2801, i_10_2802, i_10_2803, i_10_2804, i_10_2805, i_10_2806, i_10_2807, i_10_2808, i_10_2809, i_10_2810, i_10_2811, i_10_2812, i_10_2813, i_10_2814, i_10_2815, i_10_2816, i_10_2817, i_10_2818, i_10_2819, i_10_2820, i_10_2821, i_10_2822, i_10_2823, i_10_2824, i_10_2825, i_10_2826, i_10_2827, i_10_2828, i_10_2829, i_10_2830, i_10_2831, i_10_2832, i_10_2833, i_10_2834, i_10_2835, i_10_2836, i_10_2837, i_10_2838, i_10_2839, i_10_2840, i_10_2841, i_10_2842, i_10_2843, i_10_2844, i_10_2845, i_10_2846, i_10_2847, i_10_2848, i_10_2849, i_10_2850, i_10_2851, i_10_2852, i_10_2853, i_10_2854, i_10_2855, i_10_2856, i_10_2857, i_10_2858, i_10_2859, i_10_2860, i_10_2861, i_10_2862, i_10_2863, i_10_2864, i_10_2865, i_10_2866, i_10_2867, i_10_2868, i_10_2869, i_10_2870, i_10_2871, i_10_2872, i_10_2873, i_10_2874, i_10_2875, i_10_2876, i_10_2877, i_10_2878, i_10_2879, i_10_2880, i_10_2881, i_10_2882, i_10_2883, i_10_2884, i_10_2885, i_10_2886, i_10_2887, i_10_2888, i_10_2889, i_10_2890, i_10_2891, i_10_2892, i_10_2893, i_10_2894, i_10_2895, i_10_2896, i_10_2897, i_10_2898, i_10_2899, i_10_2900, i_10_2901, i_10_2902, i_10_2903, i_10_2904, i_10_2905, i_10_2906, i_10_2907, i_10_2908, i_10_2909, i_10_2910, i_10_2911, i_10_2912, i_10_2913, i_10_2914, i_10_2915, i_10_2916, i_10_2917, i_10_2918, i_10_2919, i_10_2920, i_10_2921, i_10_2922, i_10_2923, i_10_2924, i_10_2925, i_10_2926, i_10_2927, i_10_2928, i_10_2929, i_10_2930, i_10_2931, i_10_2932, i_10_2933, i_10_2934, i_10_2935, i_10_2936, i_10_2937, i_10_2938, i_10_2939, i_10_2940, i_10_2941, i_10_2942, i_10_2943, i_10_2944, i_10_2945, i_10_2946, i_10_2947, i_10_2948, i_10_2949, i_10_2950, i_10_2951, i_10_2952, i_10_2953, i_10_2954, i_10_2955, i_10_2956, i_10_2957, i_10_2958, i_10_2959, i_10_2960, i_10_2961, i_10_2962, i_10_2963, i_10_2964, i_10_2965, i_10_2966, i_10_2967, i_10_2968, i_10_2969, i_10_2970, i_10_2971, i_10_2972, i_10_2973, i_10_2974, i_10_2975, i_10_2976, i_10_2977, i_10_2978, i_10_2979, i_10_2980, i_10_2981, i_10_2982, i_10_2983, i_10_2984, i_10_2985, i_10_2986, i_10_2987, i_10_2988, i_10_2989, i_10_2990, i_10_2991, i_10_2992, i_10_2993, i_10_2994, i_10_2995, i_10_2996, i_10_2997, i_10_2998, i_10_2999, i_10_3000, i_10_3001, i_10_3002, i_10_3003, i_10_3004, i_10_3005, i_10_3006, i_10_3007, i_10_3008, i_10_3009, i_10_3010, i_10_3011, i_10_3012, i_10_3013, i_10_3014, i_10_3015, i_10_3016, i_10_3017, i_10_3018, i_10_3019, i_10_3020, i_10_3021, i_10_3022, i_10_3023, i_10_3024, i_10_3025, i_10_3026, i_10_3027, i_10_3028, i_10_3029, i_10_3030, i_10_3031, i_10_3032, i_10_3033, i_10_3034, i_10_3035, i_10_3036, i_10_3037, i_10_3038, i_10_3039, i_10_3040, i_10_3041, i_10_3042, i_10_3043, i_10_3044, i_10_3045, i_10_3046, i_10_3047, i_10_3048, i_10_3049, i_10_3050, i_10_3051, i_10_3052, i_10_3053, i_10_3054, i_10_3055, i_10_3056, i_10_3057, i_10_3058, i_10_3059, i_10_3060, i_10_3061, i_10_3062, i_10_3063, i_10_3064, i_10_3065, i_10_3066, i_10_3067, i_10_3068, i_10_3069, i_10_3070, i_10_3071, i_10_3072, i_10_3073, i_10_3074, i_10_3075, i_10_3076, i_10_3077, i_10_3078, i_10_3079, i_10_3080, i_10_3081, i_10_3082, i_10_3083, i_10_3084, i_10_3085, i_10_3086, i_10_3087, i_10_3088, i_10_3089, i_10_3090, i_10_3091, i_10_3092, i_10_3093, i_10_3094, i_10_3095, i_10_3096, i_10_3097, i_10_3098, i_10_3099, i_10_3100, i_10_3101, i_10_3102, i_10_3103, i_10_3104, i_10_3105, i_10_3106, i_10_3107, i_10_3108, i_10_3109, i_10_3110, i_10_3111, i_10_3112, i_10_3113, i_10_3114, i_10_3115, i_10_3116, i_10_3117, i_10_3118, i_10_3119, i_10_3120, i_10_3121, i_10_3122, i_10_3123, i_10_3124, i_10_3125, i_10_3126, i_10_3127, i_10_3128, i_10_3129, i_10_3130, i_10_3131, i_10_3132, i_10_3133, i_10_3134, i_10_3135, i_10_3136, i_10_3137, i_10_3138, i_10_3139, i_10_3140, i_10_3141, i_10_3142, i_10_3143, i_10_3144, i_10_3145, i_10_3146, i_10_3147, i_10_3148, i_10_3149, i_10_3150, i_10_3151, i_10_3152, i_10_3153, i_10_3154, i_10_3155, i_10_3156, i_10_3157, i_10_3158, i_10_3159, i_10_3160, i_10_3161, i_10_3162, i_10_3163, i_10_3164, i_10_3165, i_10_3166, i_10_3167, i_10_3168, i_10_3169, i_10_3170, i_10_3171, i_10_3172, i_10_3173, i_10_3174, i_10_3175, i_10_3176, i_10_3177, i_10_3178, i_10_3179, i_10_3180, i_10_3181, i_10_3182, i_10_3183, i_10_3184, i_10_3185, i_10_3186, i_10_3187, i_10_3188, i_10_3189, i_10_3190, i_10_3191, i_10_3192, i_10_3193, i_10_3194, i_10_3195, i_10_3196, i_10_3197, i_10_3198, i_10_3199, i_10_3200, i_10_3201, i_10_3202, i_10_3203, i_10_3204, i_10_3205, i_10_3206, i_10_3207, i_10_3208, i_10_3209, i_10_3210, i_10_3211, i_10_3212, i_10_3213, i_10_3214, i_10_3215, i_10_3216, i_10_3217, i_10_3218, i_10_3219, i_10_3220, i_10_3221, i_10_3222, i_10_3223, i_10_3224, i_10_3225, i_10_3226, i_10_3227, i_10_3228, i_10_3229, i_10_3230, i_10_3231, i_10_3232, i_10_3233, i_10_3234, i_10_3235, i_10_3236, i_10_3237, i_10_3238, i_10_3239, i_10_3240, i_10_3241, i_10_3242, i_10_3243, i_10_3244, i_10_3245, i_10_3246, i_10_3247, i_10_3248, i_10_3249, i_10_3250, i_10_3251, i_10_3252, i_10_3253, i_10_3254, i_10_3255, i_10_3256, i_10_3257, i_10_3258, i_10_3259, i_10_3260, i_10_3261, i_10_3262, i_10_3263, i_10_3264, i_10_3265, i_10_3266, i_10_3267, i_10_3268, i_10_3269, i_10_3270, i_10_3271, i_10_3272, i_10_3273, i_10_3274, i_10_3275, i_10_3276, i_10_3277, i_10_3278, i_10_3279, i_10_3280, i_10_3281, i_10_3282, i_10_3283, i_10_3284, i_10_3285, i_10_3286, i_10_3287, i_10_3288, i_10_3289, i_10_3290, i_10_3291, i_10_3292, i_10_3293, i_10_3294, i_10_3295, i_10_3296, i_10_3297, i_10_3298, i_10_3299, i_10_3300, i_10_3301, i_10_3302, i_10_3303, i_10_3304, i_10_3305, i_10_3306, i_10_3307, i_10_3308, i_10_3309, i_10_3310, i_10_3311, i_10_3312, i_10_3313, i_10_3314, i_10_3315, i_10_3316, i_10_3317, i_10_3318, i_10_3319, i_10_3320, i_10_3321, i_10_3322, i_10_3323, i_10_3324, i_10_3325, i_10_3326, i_10_3327, i_10_3328, i_10_3329, i_10_3330, i_10_3331, i_10_3332, i_10_3333, i_10_3334, i_10_3335, i_10_3336, i_10_3337, i_10_3338, i_10_3339, i_10_3340, i_10_3341, i_10_3342, i_10_3343, i_10_3344, i_10_3345, i_10_3346, i_10_3347, i_10_3348, i_10_3349, i_10_3350, i_10_3351, i_10_3352, i_10_3353, i_10_3354, i_10_3355, i_10_3356, i_10_3357, i_10_3358, i_10_3359, i_10_3360, i_10_3361, i_10_3362, i_10_3363, i_10_3364, i_10_3365, i_10_3366, i_10_3367, i_10_3368, i_10_3369, i_10_3370, i_10_3371, i_10_3372, i_10_3373, i_10_3374, i_10_3375, i_10_3376, i_10_3377, i_10_3378, i_10_3379, i_10_3380, i_10_3381, i_10_3382, i_10_3383, i_10_3384, i_10_3385, i_10_3386, i_10_3387, i_10_3388, i_10_3389, i_10_3390, i_10_3391, i_10_3392, i_10_3393, i_10_3394, i_10_3395, i_10_3396, i_10_3397, i_10_3398, i_10_3399, i_10_3400, i_10_3401, i_10_3402, i_10_3403, i_10_3404, i_10_3405, i_10_3406, i_10_3407, i_10_3408, i_10_3409, i_10_3410, i_10_3411, i_10_3412, i_10_3413, i_10_3414, i_10_3415, i_10_3416, i_10_3417, i_10_3418, i_10_3419, i_10_3420, i_10_3421, i_10_3422, i_10_3423, i_10_3424, i_10_3425, i_10_3426, i_10_3427, i_10_3428, i_10_3429, i_10_3430, i_10_3431, i_10_3432, i_10_3433, i_10_3434, i_10_3435, i_10_3436, i_10_3437, i_10_3438, i_10_3439, i_10_3440, i_10_3441, i_10_3442, i_10_3443, i_10_3444, i_10_3445, i_10_3446, i_10_3447, i_10_3448, i_10_3449, i_10_3450, i_10_3451, i_10_3452, i_10_3453, i_10_3454, i_10_3455, i_10_3456, i_10_3457, i_10_3458, i_10_3459, i_10_3460, i_10_3461, i_10_3462, i_10_3463, i_10_3464, i_10_3465, i_10_3466, i_10_3467, i_10_3468, i_10_3469, i_10_3470, i_10_3471, i_10_3472, i_10_3473, i_10_3474, i_10_3475, i_10_3476, i_10_3477, i_10_3478, i_10_3479, i_10_3480, i_10_3481, i_10_3482, i_10_3483, i_10_3484, i_10_3485, i_10_3486, i_10_3487, i_10_3488, i_10_3489, i_10_3490, i_10_3491, i_10_3492, i_10_3493, i_10_3494, i_10_3495, i_10_3496, i_10_3497, i_10_3498, i_10_3499, i_10_3500, i_10_3501, i_10_3502, i_10_3503, i_10_3504, i_10_3505, i_10_3506, i_10_3507, i_10_3508, i_10_3509, i_10_3510, i_10_3511, i_10_3512, i_10_3513, i_10_3514, i_10_3515, i_10_3516, i_10_3517, i_10_3518, i_10_3519, i_10_3520, i_10_3521, i_10_3522, i_10_3523, i_10_3524, i_10_3525, i_10_3526, i_10_3527, i_10_3528, i_10_3529, i_10_3530, i_10_3531, i_10_3532, i_10_3533, i_10_3534, i_10_3535, i_10_3536, i_10_3537, i_10_3538, i_10_3539, i_10_3540, i_10_3541, i_10_3542, i_10_3543, i_10_3544, i_10_3545, i_10_3546, i_10_3547, i_10_3548, i_10_3549, i_10_3550, i_10_3551, i_10_3552, i_10_3553, i_10_3554, i_10_3555, i_10_3556, i_10_3557, i_10_3558, i_10_3559, i_10_3560, i_10_3561, i_10_3562, i_10_3563, i_10_3564, i_10_3565, i_10_3566, i_10_3567, i_10_3568, i_10_3569, i_10_3570, i_10_3571, i_10_3572, i_10_3573, i_10_3574, i_10_3575, i_10_3576, i_10_3577, i_10_3578, i_10_3579, i_10_3580, i_10_3581, i_10_3582, i_10_3583, i_10_3584, i_10_3585, i_10_3586, i_10_3587, i_10_3588, i_10_3589, i_10_3590, i_10_3591, i_10_3592, i_10_3593, i_10_3594, i_10_3595, i_10_3596, i_10_3597, i_10_3598, i_10_3599, i_10_3600, i_10_3601, i_10_3602, i_10_3603, i_10_3604, i_10_3605, i_10_3606, i_10_3607, i_10_3608, i_10_3609, i_10_3610, i_10_3611, i_10_3612, i_10_3613, i_10_3614, i_10_3615, i_10_3616, i_10_3617, i_10_3618, i_10_3619, i_10_3620, i_10_3621, i_10_3622, i_10_3623, i_10_3624, i_10_3625, i_10_3626, i_10_3627, i_10_3628, i_10_3629, i_10_3630, i_10_3631, i_10_3632, i_10_3633, i_10_3634, i_10_3635, i_10_3636, i_10_3637, i_10_3638, i_10_3639, i_10_3640, i_10_3641, i_10_3642, i_10_3643, i_10_3644, i_10_3645, i_10_3646, i_10_3647, i_10_3648, i_10_3649, i_10_3650, i_10_3651, i_10_3652, i_10_3653, i_10_3654, i_10_3655, i_10_3656, i_10_3657, i_10_3658, i_10_3659, i_10_3660, i_10_3661, i_10_3662, i_10_3663, i_10_3664, i_10_3665, i_10_3666, i_10_3667, i_10_3668, i_10_3669, i_10_3670, i_10_3671, i_10_3672, i_10_3673, i_10_3674, i_10_3675, i_10_3676, i_10_3677, i_10_3678, i_10_3679, i_10_3680, i_10_3681, i_10_3682, i_10_3683, i_10_3684, i_10_3685, i_10_3686, i_10_3687, i_10_3688, i_10_3689, i_10_3690, i_10_3691, i_10_3692, i_10_3693, i_10_3694, i_10_3695, i_10_3696, i_10_3697, i_10_3698, i_10_3699, i_10_3700, i_10_3701, i_10_3702, i_10_3703, i_10_3704, i_10_3705, i_10_3706, i_10_3707, i_10_3708, i_10_3709, i_10_3710, i_10_3711, i_10_3712, i_10_3713, i_10_3714, i_10_3715, i_10_3716, i_10_3717, i_10_3718, i_10_3719, i_10_3720, i_10_3721, i_10_3722, i_10_3723, i_10_3724, i_10_3725, i_10_3726, i_10_3727, i_10_3728, i_10_3729, i_10_3730, i_10_3731, i_10_3732, i_10_3733, i_10_3734, i_10_3735, i_10_3736, i_10_3737, i_10_3738, i_10_3739, i_10_3740, i_10_3741, i_10_3742, i_10_3743, i_10_3744, i_10_3745, i_10_3746, i_10_3747, i_10_3748, i_10_3749, i_10_3750, i_10_3751, i_10_3752, i_10_3753, i_10_3754, i_10_3755, i_10_3756, i_10_3757, i_10_3758, i_10_3759, i_10_3760, i_10_3761, i_10_3762, i_10_3763, i_10_3764, i_10_3765, i_10_3766, i_10_3767, i_10_3768, i_10_3769, i_10_3770, i_10_3771, i_10_3772, i_10_3773, i_10_3774, i_10_3775, i_10_3776, i_10_3777, i_10_3778, i_10_3779, i_10_3780, i_10_3781, i_10_3782, i_10_3783, i_10_3784, i_10_3785, i_10_3786, i_10_3787, i_10_3788, i_10_3789, i_10_3790, i_10_3791, i_10_3792, i_10_3793, i_10_3794, i_10_3795, i_10_3796, i_10_3797, i_10_3798, i_10_3799, i_10_3800, i_10_3801, i_10_3802, i_10_3803, i_10_3804, i_10_3805, i_10_3806, i_10_3807, i_10_3808, i_10_3809, i_10_3810, i_10_3811, i_10_3812, i_10_3813, i_10_3814, i_10_3815, i_10_3816, i_10_3817, i_10_3818, i_10_3819, i_10_3820, i_10_3821, i_10_3822, i_10_3823, i_10_3824, i_10_3825, i_10_3826, i_10_3827, i_10_3828, i_10_3829, i_10_3830, i_10_3831, i_10_3832, i_10_3833, i_10_3834, i_10_3835, i_10_3836, i_10_3837, i_10_3838, i_10_3839, i_10_3840, i_10_3841, i_10_3842, i_10_3843, i_10_3844, i_10_3845, i_10_3846, i_10_3847, i_10_3848, i_10_3849, i_10_3850, i_10_3851, i_10_3852, i_10_3853, i_10_3854, i_10_3855, i_10_3856, i_10_3857, i_10_3858, i_10_3859, i_10_3860, i_10_3861, i_10_3862, i_10_3863, i_10_3864, i_10_3865, i_10_3866, i_10_3867, i_10_3868, i_10_3869, i_10_3870, i_10_3871, i_10_3872, i_10_3873, i_10_3874, i_10_3875, i_10_3876, i_10_3877, i_10_3878, i_10_3879, i_10_3880, i_10_3881, i_10_3882, i_10_3883, i_10_3884, i_10_3885, i_10_3886, i_10_3887, i_10_3888, i_10_3889, i_10_3890, i_10_3891, i_10_3892, i_10_3893, i_10_3894, i_10_3895, i_10_3896, i_10_3897, i_10_3898, i_10_3899, i_10_3900, i_10_3901, i_10_3902, i_10_3903, i_10_3904, i_10_3905, i_10_3906, i_10_3907, i_10_3908, i_10_3909, i_10_3910, i_10_3911, i_10_3912, i_10_3913, i_10_3914, i_10_3915, i_10_3916, i_10_3917, i_10_3918, i_10_3919, i_10_3920, i_10_3921, i_10_3922, i_10_3923, i_10_3924, i_10_3925, i_10_3926, i_10_3927, i_10_3928, i_10_3929, i_10_3930, i_10_3931, i_10_3932, i_10_3933, i_10_3934, i_10_3935, i_10_3936, i_10_3937, i_10_3938, i_10_3939, i_10_3940, i_10_3941, i_10_3942, i_10_3943, i_10_3944, i_10_3945, i_10_3946, i_10_3947, i_10_3948, i_10_3949, i_10_3950, i_10_3951, i_10_3952, i_10_3953, i_10_3954, i_10_3955, i_10_3956, i_10_3957, i_10_3958, i_10_3959, i_10_3960, i_10_3961, i_10_3962, i_10_3963, i_10_3964, i_10_3965, i_10_3966, i_10_3967, i_10_3968, i_10_3969, i_10_3970, i_10_3971, i_10_3972, i_10_3973, i_10_3974, i_10_3975, i_10_3976, i_10_3977, i_10_3978, i_10_3979, i_10_3980, i_10_3981, i_10_3982, i_10_3983, i_10_3984, i_10_3985, i_10_3986, i_10_3987, i_10_3988, i_10_3989, i_10_3990, i_10_3991, i_10_3992, i_10_3993, i_10_3994, i_10_3995, i_10_3996, i_10_3997, i_10_3998, i_10_3999, i_10_4000, i_10_4001, i_10_4002, i_10_4003, i_10_4004, i_10_4005, i_10_4006, i_10_4007, i_10_4008, i_10_4009, i_10_4010, i_10_4011, i_10_4012, i_10_4013, i_10_4014, i_10_4015, i_10_4016, i_10_4017, i_10_4018, i_10_4019, i_10_4020, i_10_4021, i_10_4022, i_10_4023, i_10_4024, i_10_4025, i_10_4026, i_10_4027, i_10_4028, i_10_4029, i_10_4030, i_10_4031, i_10_4032, i_10_4033, i_10_4034, i_10_4035, i_10_4036, i_10_4037, i_10_4038, i_10_4039, i_10_4040, i_10_4041, i_10_4042, i_10_4043, i_10_4044, i_10_4045, i_10_4046, i_10_4047, i_10_4048, i_10_4049, i_10_4050, i_10_4051, i_10_4052, i_10_4053, i_10_4054, i_10_4055, i_10_4056, i_10_4057, i_10_4058, i_10_4059, i_10_4060, i_10_4061, i_10_4062, i_10_4063, i_10_4064, i_10_4065, i_10_4066, i_10_4067, i_10_4068, i_10_4069, i_10_4070, i_10_4071, i_10_4072, i_10_4073, i_10_4074, i_10_4075, i_10_4076, i_10_4077, i_10_4078, i_10_4079, i_10_4080, i_10_4081, i_10_4082, i_10_4083, i_10_4084, i_10_4085, i_10_4086, i_10_4087, i_10_4088, i_10_4089, i_10_4090, i_10_4091, i_10_4092, i_10_4093, i_10_4094, i_10_4095, i_10_4096, i_10_4097, i_10_4098, i_10_4099, i_10_4100, i_10_4101, i_10_4102, i_10_4103, i_10_4104, i_10_4105, i_10_4106, i_10_4107, i_10_4108, i_10_4109, i_10_4110, i_10_4111, i_10_4112, i_10_4113, i_10_4114, i_10_4115, i_10_4116, i_10_4117, i_10_4118, i_10_4119, i_10_4120, i_10_4121, i_10_4122, i_10_4123, i_10_4124, i_10_4125, i_10_4126, i_10_4127, i_10_4128, i_10_4129, i_10_4130, i_10_4131, i_10_4132, i_10_4133, i_10_4134, i_10_4135, i_10_4136, i_10_4137, i_10_4138, i_10_4139, i_10_4140, i_10_4141, i_10_4142, i_10_4143, i_10_4144, i_10_4145, i_10_4146, i_10_4147, i_10_4148, i_10_4149, i_10_4150, i_10_4151, i_10_4152, i_10_4153, i_10_4154, i_10_4155, i_10_4156, i_10_4157, i_10_4158, i_10_4159, i_10_4160, i_10_4161, i_10_4162, i_10_4163, i_10_4164, i_10_4165, i_10_4166, i_10_4167, i_10_4168, i_10_4169, i_10_4170, i_10_4171, i_10_4172, i_10_4173, i_10_4174, i_10_4175, i_10_4176, i_10_4177, i_10_4178, i_10_4179, i_10_4180, i_10_4181, i_10_4182, i_10_4183, i_10_4184, i_10_4185, i_10_4186, i_10_4187, i_10_4188, i_10_4189, i_10_4190, i_10_4191, i_10_4192, i_10_4193, i_10_4194, i_10_4195, i_10_4196, i_10_4197, i_10_4198, i_10_4199, i_10_4200, i_10_4201, i_10_4202, i_10_4203, i_10_4204, i_10_4205, i_10_4206, i_10_4207, i_10_4208, i_10_4209, i_10_4210, i_10_4211, i_10_4212, i_10_4213, i_10_4214, i_10_4215, i_10_4216, i_10_4217, i_10_4218, i_10_4219, i_10_4220, i_10_4221, i_10_4222, i_10_4223, i_10_4224, i_10_4225, i_10_4226, i_10_4227, i_10_4228, i_10_4229, i_10_4230, i_10_4231, i_10_4232, i_10_4233, i_10_4234, i_10_4235, i_10_4236, i_10_4237, i_10_4238, i_10_4239, i_10_4240, i_10_4241, i_10_4242, i_10_4243, i_10_4244, i_10_4245, i_10_4246, i_10_4247, i_10_4248, i_10_4249, i_10_4250, i_10_4251, i_10_4252, i_10_4253, i_10_4254, i_10_4255, i_10_4256, i_10_4257, i_10_4258, i_10_4259, i_10_4260, i_10_4261, i_10_4262, i_10_4263, i_10_4264, i_10_4265, i_10_4266, i_10_4267, i_10_4268, i_10_4269, i_10_4270, i_10_4271, i_10_4272, i_10_4273, i_10_4274, i_10_4275, i_10_4276, i_10_4277, i_10_4278, i_10_4279, i_10_4280, i_10_4281, i_10_4282, i_10_4283, i_10_4284, i_10_4285, i_10_4286, i_10_4287, i_10_4288, i_10_4289, i_10_4290, i_10_4291, i_10_4292, i_10_4293, i_10_4294, i_10_4295, i_10_4296, i_10_4297, i_10_4298, i_10_4299, i_10_4300, i_10_4301, i_10_4302, i_10_4303, i_10_4304, i_10_4305, i_10_4306, i_10_4307, i_10_4308, i_10_4309, i_10_4310, i_10_4311, i_10_4312, i_10_4313, i_10_4314, i_10_4315, i_10_4316, i_10_4317, i_10_4318, i_10_4319, i_10_4320, i_10_4321, i_10_4322, i_10_4323, i_10_4324, i_10_4325, i_10_4326, i_10_4327, i_10_4328, i_10_4329, i_10_4330, i_10_4331, i_10_4332, i_10_4333, i_10_4334, i_10_4335, i_10_4336, i_10_4337, i_10_4338, i_10_4339, i_10_4340, i_10_4341, i_10_4342, i_10_4343, i_10_4344, i_10_4345, i_10_4346, i_10_4347, i_10_4348, i_10_4349, i_10_4350, i_10_4351, i_10_4352, i_10_4353, i_10_4354, i_10_4355, i_10_4356, i_10_4357, i_10_4358, i_10_4359, i_10_4360, i_10_4361, i_10_4362, i_10_4363, i_10_4364, i_10_4365, i_10_4366, i_10_4367, i_10_4368, i_10_4369, i_10_4370, i_10_4371, i_10_4372, i_10_4373, i_10_4374, i_10_4375, i_10_4376, i_10_4377, i_10_4378, i_10_4379, i_10_4380, i_10_4381, i_10_4382, i_10_4383, i_10_4384, i_10_4385, i_10_4386, i_10_4387, i_10_4388, i_10_4389, i_10_4390, i_10_4391, i_10_4392, i_10_4393, i_10_4394, i_10_4395, i_10_4396, i_10_4397, i_10_4398, i_10_4399, i_10_4400, i_10_4401, i_10_4402, i_10_4403, i_10_4404, i_10_4405, i_10_4406, i_10_4407, i_10_4408, i_10_4409, i_10_4410, i_10_4411, i_10_4412, i_10_4413, i_10_4414, i_10_4415, i_10_4416, i_10_4417, i_10_4418, i_10_4419, i_10_4420, i_10_4421, i_10_4422, i_10_4423, i_10_4424, i_10_4425, i_10_4426, i_10_4427, i_10_4428, i_10_4429, i_10_4430, i_10_4431, i_10_4432, i_10_4433, i_10_4434, i_10_4435, i_10_4436, i_10_4437, i_10_4438, i_10_4439, i_10_4440, i_10_4441, i_10_4442, i_10_4443, i_10_4444, i_10_4445, i_10_4446, i_10_4447, i_10_4448, i_10_4449, i_10_4450, i_10_4451, i_10_4452, i_10_4453, i_10_4454, i_10_4455, i_10_4456, i_10_4457, i_10_4458, i_10_4459, i_10_4460, i_10_4461, i_10_4462, i_10_4463, i_10_4464, i_10_4465, i_10_4466, i_10_4467, i_10_4468, i_10_4469, i_10_4470, i_10_4471, i_10_4472, i_10_4473, i_10_4474, i_10_4475, i_10_4476, i_10_4477, i_10_4478, i_10_4479, i_10_4480, i_10_4481, i_10_4482, i_10_4483, i_10_4484, i_10_4485, i_10_4486, i_10_4487, i_10_4488, i_10_4489, i_10_4490, i_10_4491, i_10_4492, i_10_4493, i_10_4494, i_10_4495, i_10_4496, i_10_4497, i_10_4498, i_10_4499, i_10_4500, i_10_4501, i_10_4502, i_10_4503, i_10_4504, i_10_4505, i_10_4506, i_10_4507, i_10_4508, i_10_4509, i_10_4510, i_10_4511, i_10_4512, i_10_4513, i_10_4514, i_10_4515, i_10_4516, i_10_4517, i_10_4518, i_10_4519, i_10_4520, i_10_4521, i_10_4522, i_10_4523, i_10_4524, i_10_4525, i_10_4526, i_10_4527, i_10_4528, i_10_4529, i_10_4530, i_10_4531, i_10_4532, i_10_4533, i_10_4534, i_10_4535, i_10_4536, i_10_4537, i_10_4538, i_10_4539, i_10_4540, i_10_4541, i_10_4542, i_10_4543, i_10_4544, i_10_4545, i_10_4546, i_10_4547, i_10_4548, i_10_4549, i_10_4550, i_10_4551, i_10_4552, i_10_4553, i_10_4554, i_10_4555, i_10_4556, i_10_4557, i_10_4558, i_10_4559, i_10_4560, i_10_4561, i_10_4562, i_10_4563, i_10_4564, i_10_4565, i_10_4566, i_10_4567, i_10_4568, i_10_4569, i_10_4570, i_10_4571, i_10_4572, i_10_4573, i_10_4574, i_10_4575, i_10_4576, i_10_4577, i_10_4578, i_10_4579, i_10_4580, i_10_4581, i_10_4582, i_10_4583, i_10_4584, i_10_4585, i_10_4586, i_10_4587, i_10_4588, i_10_4589, i_10_4590, i_10_4591, i_10_4592, i_10_4593, i_10_4594, i_10_4595, i_10_4596, i_10_4597, i_10_4598, i_10_4599, i_10_4600, i_10_4601, i_10_4602, i_10_4603, i_10_4604, i_10_4605, i_10_4606, i_10_4607;
output o_10_0, o_10_1, o_10_2, o_10_3, o_10_4, o_10_5, o_10_6, o_10_7, o_10_8, o_10_9, o_10_10, o_10_11, o_10_12, o_10_13, o_10_14, o_10_15, o_10_16, o_10_17, o_10_18, o_10_19, o_10_20, o_10_21, o_10_22, o_10_23, o_10_24, o_10_25, o_10_26, o_10_27, o_10_28, o_10_29, o_10_30, o_10_31, o_10_32, o_10_33, o_10_34, o_10_35, o_10_36, o_10_37, o_10_38, o_10_39, o_10_40, o_10_41, o_10_42, o_10_43, o_10_44, o_10_45, o_10_46, o_10_47, o_10_48, o_10_49, o_10_50, o_10_51, o_10_52, o_10_53, o_10_54, o_10_55, o_10_56, o_10_57, o_10_58, o_10_59, o_10_60, o_10_61, o_10_62, o_10_63, o_10_64, o_10_65, o_10_66, o_10_67, o_10_68, o_10_69, o_10_70, o_10_71, o_10_72, o_10_73, o_10_74, o_10_75, o_10_76, o_10_77, o_10_78, o_10_79, o_10_80, o_10_81, o_10_82, o_10_83, o_10_84, o_10_85, o_10_86, o_10_87, o_10_88, o_10_89, o_10_90, o_10_91, o_10_92, o_10_93, o_10_94, o_10_95, o_10_96, o_10_97, o_10_98, o_10_99, o_10_100, o_10_101, o_10_102, o_10_103, o_10_104, o_10_105, o_10_106, o_10_107, o_10_108, o_10_109, o_10_110, o_10_111, o_10_112, o_10_113, o_10_114, o_10_115, o_10_116, o_10_117, o_10_118, o_10_119, o_10_120, o_10_121, o_10_122, o_10_123, o_10_124, o_10_125, o_10_126, o_10_127, o_10_128, o_10_129, o_10_130, o_10_131, o_10_132, o_10_133, o_10_134, o_10_135, o_10_136, o_10_137, o_10_138, o_10_139, o_10_140, o_10_141, o_10_142, o_10_143, o_10_144, o_10_145, o_10_146, o_10_147, o_10_148, o_10_149, o_10_150, o_10_151, o_10_152, o_10_153, o_10_154, o_10_155, o_10_156, o_10_157, o_10_158, o_10_159, o_10_160, o_10_161, o_10_162, o_10_163, o_10_164, o_10_165, o_10_166, o_10_167, o_10_168, o_10_169, o_10_170, o_10_171, o_10_172, o_10_173, o_10_174, o_10_175, o_10_176, o_10_177, o_10_178, o_10_179, o_10_180, o_10_181, o_10_182, o_10_183, o_10_184, o_10_185, o_10_186, o_10_187, o_10_188, o_10_189, o_10_190, o_10_191, o_10_192, o_10_193, o_10_194, o_10_195, o_10_196, o_10_197, o_10_198, o_10_199, o_10_200, o_10_201, o_10_202, o_10_203, o_10_204, o_10_205, o_10_206, o_10_207, o_10_208, o_10_209, o_10_210, o_10_211, o_10_212, o_10_213, o_10_214, o_10_215, o_10_216, o_10_217, o_10_218, o_10_219, o_10_220, o_10_221, o_10_222, o_10_223, o_10_224, o_10_225, o_10_226, o_10_227, o_10_228, o_10_229, o_10_230, o_10_231, o_10_232, o_10_233, o_10_234, o_10_235, o_10_236, o_10_237, o_10_238, o_10_239, o_10_240, o_10_241, o_10_242, o_10_243, o_10_244, o_10_245, o_10_246, o_10_247, o_10_248, o_10_249, o_10_250, o_10_251, o_10_252, o_10_253, o_10_254, o_10_255, o_10_256, o_10_257, o_10_258, o_10_259, o_10_260, o_10_261, o_10_262, o_10_263, o_10_264, o_10_265, o_10_266, o_10_267, o_10_268, o_10_269, o_10_270, o_10_271, o_10_272, o_10_273, o_10_274, o_10_275, o_10_276, o_10_277, o_10_278, o_10_279, o_10_280, o_10_281, o_10_282, o_10_283, o_10_284, o_10_285, o_10_286, o_10_287, o_10_288, o_10_289, o_10_290, o_10_291, o_10_292, o_10_293, o_10_294, o_10_295, o_10_296, o_10_297, o_10_298, o_10_299, o_10_300, o_10_301, o_10_302, o_10_303, o_10_304, o_10_305, o_10_306, o_10_307, o_10_308, o_10_309, o_10_310, o_10_311, o_10_312, o_10_313, o_10_314, o_10_315, o_10_316, o_10_317, o_10_318, o_10_319, o_10_320, o_10_321, o_10_322, o_10_323, o_10_324, o_10_325, o_10_326, o_10_327, o_10_328, o_10_329, o_10_330, o_10_331, o_10_332, o_10_333, o_10_334, o_10_335, o_10_336, o_10_337, o_10_338, o_10_339, o_10_340, o_10_341, o_10_342, o_10_343, o_10_344, o_10_345, o_10_346, o_10_347, o_10_348, o_10_349, o_10_350, o_10_351, o_10_352, o_10_353, o_10_354, o_10_355, o_10_356, o_10_357, o_10_358, o_10_359, o_10_360, o_10_361, o_10_362, o_10_363, o_10_364, o_10_365, o_10_366, o_10_367, o_10_368, o_10_369, o_10_370, o_10_371, o_10_372, o_10_373, o_10_374, o_10_375, o_10_376, o_10_377, o_10_378, o_10_379, o_10_380, o_10_381, o_10_382, o_10_383, o_10_384, o_10_385, o_10_386, o_10_387, o_10_388, o_10_389, o_10_390, o_10_391, o_10_392, o_10_393, o_10_394, o_10_395, o_10_396, o_10_397, o_10_398, o_10_399, o_10_400, o_10_401, o_10_402, o_10_403, o_10_404, o_10_405, o_10_406, o_10_407, o_10_408, o_10_409, o_10_410, o_10_411, o_10_412, o_10_413, o_10_414, o_10_415, o_10_416, o_10_417, o_10_418, o_10_419, o_10_420, o_10_421, o_10_422, o_10_423, o_10_424, o_10_425, o_10_426, o_10_427, o_10_428, o_10_429, o_10_430, o_10_431, o_10_432, o_10_433, o_10_434, o_10_435, o_10_436, o_10_437, o_10_438, o_10_439, o_10_440, o_10_441, o_10_442, o_10_443, o_10_444, o_10_445, o_10_446, o_10_447, o_10_448, o_10_449, o_10_450, o_10_451, o_10_452, o_10_453, o_10_454, o_10_455, o_10_456, o_10_457, o_10_458, o_10_459, o_10_460, o_10_461, o_10_462, o_10_463, o_10_464, o_10_465, o_10_466, o_10_467, o_10_468, o_10_469, o_10_470, o_10_471, o_10_472, o_10_473, o_10_474, o_10_475, o_10_476, o_10_477, o_10_478, o_10_479, o_10_480, o_10_481, o_10_482, o_10_483, o_10_484, o_10_485, o_10_486, o_10_487, o_10_488, o_10_489, o_10_490, o_10_491, o_10_492, o_10_493, o_10_494, o_10_495, o_10_496, o_10_497, o_10_498, o_10_499, o_10_500, o_10_501, o_10_502, o_10_503, o_10_504, o_10_505, o_10_506, o_10_507, o_10_508, o_10_509, o_10_510, o_10_511;
	kernel_10_0 k_10_0(i_10_31, i_10_180, i_10_185, i_10_216, i_10_277, i_10_278, i_10_286, i_10_324, i_10_408, i_10_424, i_10_427, i_10_432, i_10_433, i_10_444, i_10_465, i_10_514, i_10_697, i_10_954, i_10_955, i_10_956, i_10_957, i_10_970, i_10_994, i_10_1116, i_10_1119, i_10_1167, i_10_1239, i_10_1243, i_10_1244, i_10_1307, i_10_1540, i_10_1541, i_10_1547, i_10_1549, i_10_1550, i_10_1690, i_10_1758, i_10_1760, i_10_1818, i_10_1909, i_10_1911, i_10_1984, i_10_2023, i_10_2029, i_10_2434, i_10_2442, i_10_2443, i_10_2455, i_10_2456, i_10_2534, i_10_2659, i_10_2719, i_10_2821, i_10_2830, i_10_2880, i_10_2881, i_10_2883, i_10_2886, i_10_2887, i_10_2919, i_10_2920, i_10_3034, i_10_3075, i_10_3198, i_10_3384, i_10_3385, i_10_3386, i_10_3387, i_10_3388, i_10_3389, i_10_3437, i_10_3537, i_10_3540, i_10_3647, i_10_3650, i_10_3652, i_10_3685, i_10_3686, i_10_3720, i_10_3783, i_10_3784, i_10_3785, i_10_3787, i_10_3811, i_10_3812, i_10_3842, i_10_3847, i_10_3848, i_10_3908, i_10_3963, i_10_3982, i_10_3994, i_10_3995, i_10_4115, i_10_4172, i_10_4215, i_10_4216, i_10_4218, i_10_4283, i_10_4530, o_10_0);
	kernel_10_1 k_10_1(i_10_53, i_10_86, i_10_118, i_10_280, i_10_424, i_10_427, i_10_436, i_10_437, i_10_442, i_10_444, i_10_459, i_10_463, i_10_467, i_10_514, i_10_518, i_10_587, i_10_706, i_10_746, i_10_764, i_10_793, i_10_794, i_10_832, i_10_833, i_10_964, i_10_989, i_10_991, i_10_1054, i_10_1055, i_10_1361, i_10_1466, i_10_1541, i_10_1619, i_10_1684, i_10_1685, i_10_1768, i_10_1819, i_10_1821, i_10_1862, i_10_2182, i_10_2306, i_10_2330, i_10_2333, i_10_2336, i_10_2357, i_10_2360, i_10_2449, i_10_2453, i_10_2468, i_10_2478, i_10_2482, i_10_2515, i_10_2528, i_10_2539, i_10_2628, i_10_2630, i_10_2676, i_10_2681, i_10_2717, i_10_2728, i_10_2827, i_10_2828, i_10_2830, i_10_2873, i_10_2917, i_10_2918, i_10_2920, i_10_2921, i_10_3195, i_10_3197, i_10_3206, i_10_3208, i_10_3209, i_10_3353, i_10_3384, i_10_3403, i_10_3404, i_10_3434, i_10_3451, i_10_3583, i_10_3584, i_10_3587, i_10_3589, i_10_3610, i_10_3614, i_10_3620, i_10_3688, i_10_3734, i_10_3835, i_10_3836, i_10_3857, i_10_3920, i_10_3988, i_10_4031, i_10_4144, i_10_4147, i_10_4171, i_10_4192, i_10_4279, i_10_4577, i_10_4586, o_10_1);
	kernel_10_2 k_10_2(i_10_171, i_10_174, i_10_175, i_10_176, i_10_216, i_10_217, i_10_316, i_10_317, i_10_318, i_10_321, i_10_322, i_10_412, i_10_429, i_10_442, i_10_467, i_10_797, i_10_800, i_10_892, i_10_958, i_10_959, i_10_1006, i_10_1026, i_10_1027, i_10_1029, i_10_1134, i_10_1233, i_10_1234, i_10_1235, i_10_1236, i_10_1237, i_10_1238, i_10_1242, i_10_1245, i_10_1306, i_10_1307, i_10_1579, i_10_1580, i_10_1651, i_10_1652, i_10_1685, i_10_1819, i_10_1820, i_10_1821, i_10_1951, i_10_1991, i_10_2184, i_10_2185, i_10_2311, i_10_2352, i_10_2359, i_10_2361, i_10_2364, i_10_2376, i_10_2410, i_10_2448, i_10_2450, i_10_2457, i_10_2458, i_10_2461, i_10_2462, i_10_2629, i_10_2631, i_10_2635, i_10_2662, i_10_2719, i_10_2819, i_10_2827, i_10_2829, i_10_2830, i_10_2918, i_10_2920, i_10_3093, i_10_3094, i_10_3151, i_10_3276, i_10_3388, i_10_3391, i_10_3402, i_10_3404, i_10_3551, i_10_3586, i_10_3609, i_10_3616, i_10_3647, i_10_3783, i_10_3784, i_10_3787, i_10_3836, i_10_3838, i_10_3847, i_10_3853, i_10_3855, i_10_3856, i_10_4127, i_10_4212, i_10_4269, i_10_4285, i_10_4564, i_10_4566, i_10_4567, o_10_2);
	kernel_10_3 k_10_3(i_10_176, i_10_289, i_10_316, i_10_325, i_10_391, i_10_406, i_10_409, i_10_433, i_10_442, i_10_444, i_10_466, i_10_622, i_10_725, i_10_792, i_10_955, i_10_1000, i_10_1027, i_10_1028, i_10_1084, i_10_1233, i_10_1235, i_10_1244, i_10_1431, i_10_1432, i_10_1433, i_10_1544, i_10_1577, i_10_1604, i_10_1683, i_10_1684, i_10_1686, i_10_1687, i_10_1914, i_10_1921, i_10_1955, i_10_1981, i_10_2017, i_10_2179, i_10_2349, i_10_2350, i_10_2351, i_10_2360, i_10_2451, i_10_2452, i_10_2453, i_10_2530, i_10_2531, i_10_2567, i_10_2605, i_10_2639, i_10_2655, i_10_2656, i_10_2657, i_10_2728, i_10_2729, i_10_2736, i_10_2737, i_10_2754, i_10_2836, i_10_2844, i_10_2883, i_10_2920, i_10_2921, i_10_3069, i_10_3072, i_10_3073, i_10_3198, i_10_3269, i_10_3315, i_10_3330, i_10_3331, i_10_3332, i_10_3350, i_10_3385, i_10_3386, i_10_3387, i_10_3406, i_10_3458, i_10_3522, i_10_3555, i_10_3556, i_10_3587, i_10_3612, i_10_3837, i_10_3838, i_10_3839, i_10_3848, i_10_3853, i_10_3855, i_10_3945, i_10_4115, i_10_4117, i_10_4122, i_10_4150, i_10_4164, i_10_4172, i_10_4178, i_10_4392, i_10_4428, i_10_4582, o_10_3);
	kernel_10_4 k_10_4(i_10_63, i_10_89, i_10_144, i_10_148, i_10_263, i_10_283, i_10_287, i_10_329, i_10_408, i_10_424, i_10_427, i_10_464, i_10_532, i_10_556, i_10_796, i_10_933, i_10_963, i_10_1003, i_10_1058, i_10_1198, i_10_1267, i_10_1306, i_10_1307, i_10_1308, i_10_1485, i_10_1488, i_10_1489, i_10_1619, i_10_1653, i_10_1654, i_10_1795, i_10_1804, i_10_1818, i_10_1917, i_10_1929, i_10_1937, i_10_1948, i_10_1949, i_10_2028, i_10_2182, i_10_2244, i_10_2247, i_10_2336, i_10_2361, i_10_2364, i_10_2430, i_10_2448, i_10_2449, i_10_2451, i_10_2454, i_10_2469, i_10_2479, i_10_2513, i_10_2515, i_10_2516, i_10_2542, i_10_2544, i_10_2662, i_10_2663, i_10_2710, i_10_2713, i_10_2724, i_10_2789, i_10_2821, i_10_2834, i_10_3043, i_10_3070, i_10_3073, i_10_3235, i_10_3280, i_10_3282, i_10_3283, i_10_3312, i_10_3315, i_10_3384, i_10_3385, i_10_3401, i_10_3454, i_10_3611, i_10_3616, i_10_3645, i_10_3685, i_10_3725, i_10_3856, i_10_3888, i_10_3891, i_10_3909, i_10_3942, i_10_4116, i_10_4156, i_10_4237, i_10_4279, i_10_4287, i_10_4288, i_10_4289, i_10_4396, i_10_4397, i_10_4531, i_10_4582, i_10_4583, o_10_4);
	kernel_10_5 k_10_5(i_10_27, i_10_45, i_10_146, i_10_203, i_10_222, i_10_243, i_10_252, i_10_279, i_10_286, i_10_287, i_10_288, i_10_465, i_10_466, i_10_467, i_10_503, i_10_517, i_10_558, i_10_747, i_10_748, i_10_798, i_10_845, i_10_954, i_10_955, i_10_1026, i_10_1031, i_10_1197, i_10_1233, i_10_1234, i_10_1236, i_10_1237, i_10_1239, i_10_1240, i_10_1241, i_10_1242, i_10_1243, i_10_1274, i_10_1311, i_10_1373, i_10_1378, i_10_1616, i_10_1648, i_10_1649, i_10_1757, i_10_1824, i_10_1912, i_10_1953, i_10_1957, i_10_1961, i_10_2161, i_10_2178, i_10_2196, i_10_2197, i_10_2254, i_10_2303, i_10_2307, i_10_2354, i_10_2357, i_10_2449, i_10_2450, i_10_2451, i_10_2454, i_10_2458, i_10_2469, i_10_2470, i_10_2489, i_10_2605, i_10_2608, i_10_2628, i_10_2629, i_10_2630, i_10_2646, i_10_2680, i_10_2696, i_10_2701, i_10_2732, i_10_2833, i_10_2886, i_10_2948, i_10_2960, i_10_3267, i_10_3268, i_10_3279, i_10_3289, i_10_3292, i_10_3301, i_10_3384, i_10_3387, i_10_3473, i_10_3588, i_10_3589, i_10_3625, i_10_3649, i_10_3724, i_10_3780, i_10_3783, i_10_3853, i_10_4165, i_10_4319, i_10_4586, i_10_4588, o_10_5);
	kernel_10_6 k_10_6(i_10_30, i_10_51, i_10_52, i_10_53, i_10_142, i_10_143, i_10_151, i_10_243, i_10_252, i_10_271, i_10_272, i_10_350, i_10_358, i_10_430, i_10_464, i_10_495, i_10_514, i_10_517, i_10_518, i_10_591, i_10_714, i_10_754, i_10_755, i_10_799, i_10_831, i_10_832, i_10_970, i_10_988, i_10_997, i_10_1082, i_10_1166, i_10_1209, i_10_1240, i_10_1357, i_10_1367, i_10_1384, i_10_1446, i_10_1635, i_10_1636, i_10_1645, i_10_1690, i_10_1764, i_10_1768, i_10_1805, i_10_1808, i_10_1824, i_10_1825, i_10_1918, i_10_1952, i_10_1959, i_10_2004, i_10_2031, i_10_2182, i_10_2185, i_10_2247, i_10_2312, i_10_2329, i_10_2360, i_10_2390, i_10_2452, i_10_2510, i_10_2573, i_10_2602, i_10_2614, i_10_2741, i_10_2882, i_10_2913, i_10_2984, i_10_3122, i_10_3202, i_10_3315, i_10_3410, i_10_3473, i_10_3497, i_10_3547, i_10_3586, i_10_3587, i_10_3684, i_10_3688, i_10_3721, i_10_3822, i_10_3849, i_10_3850, i_10_3851, i_10_3854, i_10_3856, i_10_3878, i_10_3912, i_10_3985, i_10_4028, i_10_4116, i_10_4117, i_10_4119, i_10_4120, i_10_4121, i_10_4266, i_10_4269, i_10_4289, i_10_4459, i_10_4463, o_10_6);
	kernel_10_7 k_10_7(i_10_40, i_10_173, i_10_184, i_10_185, i_10_188, i_10_271, i_10_272, i_10_283, i_10_285, i_10_370, i_10_390, i_10_391, i_10_461, i_10_463, i_10_464, i_10_465, i_10_502, i_10_563, i_10_751, i_10_754, i_10_905, i_10_917, i_10_933, i_10_934, i_10_965, i_10_966, i_10_1056, i_10_1234, i_10_1235, i_10_1241, i_10_1312, i_10_1348, i_10_1366, i_10_1543, i_10_1552, i_10_1645, i_10_1652, i_10_1686, i_10_1714, i_10_1767, i_10_1812, i_10_1813, i_10_1819, i_10_1822, i_10_1907, i_10_1922, i_10_1950, i_10_1957, i_10_1991, i_10_2023, i_10_2184, i_10_2247, i_10_2309, i_10_2388, i_10_2451, i_10_2467, i_10_2511, i_10_2516, i_10_2540, i_10_2602, i_10_2617, i_10_2735, i_10_2743, i_10_2789, i_10_2806, i_10_2807, i_10_2825, i_10_2827, i_10_2980, i_10_3198, i_10_3200, i_10_3328, i_10_3352, i_10_3353, i_10_3454, i_10_3469, i_10_3470, i_10_3525, i_10_3582, i_10_3588, i_10_3590, i_10_3622, i_10_3625, i_10_3685, i_10_3723, i_10_3839, i_10_3855, i_10_3856, i_10_3860, i_10_3881, i_10_3895, i_10_3946, i_10_3950, i_10_4054, i_10_4113, i_10_4118, i_10_4217, i_10_4237, i_10_4267, i_10_4295, o_10_7);
	kernel_10_8 k_10_8(i_10_124, i_10_174, i_10_175, i_10_176, i_10_220, i_10_223, i_10_283, i_10_284, i_10_328, i_10_329, i_10_395, i_10_433, i_10_434, i_10_442, i_10_465, i_10_518, i_10_565, i_10_793, i_10_907, i_10_954, i_10_968, i_10_991, i_10_1006, i_10_1033, i_10_1309, i_10_1310, i_10_1349, i_10_1367, i_10_1379, i_10_1439, i_10_1555, i_10_1556, i_10_1684, i_10_1685, i_10_1687, i_10_1768, i_10_1769, i_10_1810, i_10_1819, i_10_1824, i_10_1951, i_10_1952, i_10_2029, i_10_2185, i_10_2186, i_10_2201, i_10_2311, i_10_2312, i_10_2351, i_10_2353, i_10_2362, i_10_2410, i_10_2411, i_10_2449, i_10_2450, i_10_2451, i_10_2455, i_10_2504, i_10_2572, i_10_2603, i_10_2629, i_10_2632, i_10_2657, i_10_2659, i_10_2660, i_10_2680, i_10_2681, i_10_2705, i_10_2722, i_10_2723, i_10_2725, i_10_2729, i_10_2730, i_10_2731, i_10_2789, i_10_2829, i_10_2830, i_10_2923, i_10_2924, i_10_3047, i_10_3076, i_10_3158, i_10_3497, i_10_3609, i_10_3624, i_10_3650, i_10_3836, i_10_3844, i_10_3846, i_10_3855, i_10_3857, i_10_3912, i_10_3914, i_10_3986, i_10_4058, i_10_4118, i_10_4237, i_10_4285, i_10_4288, i_10_4289, o_10_8);
	kernel_10_9 k_10_9(i_10_47, i_10_146, i_10_171, i_10_176, i_10_191, i_10_224, i_10_247, i_10_279, i_10_281, i_10_287, i_10_315, i_10_317, i_10_443, i_10_459, i_10_462, i_10_463, i_10_464, i_10_509, i_10_635, i_10_821, i_10_891, i_10_894, i_10_1029, i_10_1030, i_10_1031, i_10_1085, i_10_1235, i_10_1238, i_10_1250, i_10_1297, i_10_1298, i_10_1306, i_10_1631, i_10_1634, i_10_1685, i_10_1691, i_10_1822, i_10_1912, i_10_1981, i_10_1992, i_10_2027, i_10_2107, i_10_2197, i_10_2198, i_10_2201, i_10_2288, i_10_2334, i_10_2338, i_10_2352, i_10_2358, i_10_2379, i_10_2380, i_10_2452, i_10_2468, i_10_2470, i_10_2530, i_10_2567, i_10_2650, i_10_2656, i_10_2658, i_10_2711, i_10_2714, i_10_2728, i_10_2729, i_10_2740, i_10_2741, i_10_2783, i_10_2846, i_10_2918, i_10_2990, i_10_3046, i_10_3087, i_10_3313, i_10_3389, i_10_3390, i_10_3391, i_10_3395, i_10_3467, i_10_3502, i_10_3539, i_10_3557, i_10_3587, i_10_3612, i_10_3650, i_10_3652, i_10_3787, i_10_3838, i_10_3841, i_10_3847, i_10_3848, i_10_3910, i_10_3982, i_10_4027, i_10_4028, i_10_4113, i_10_4124, i_10_4172, i_10_4215, i_10_4277, i_10_4280, o_10_9);
	kernel_10_10 k_10_10(i_10_283, i_10_285, i_10_319, i_10_426, i_10_435, i_10_507, i_10_622, i_10_636, i_10_891, i_10_897, i_10_949, i_10_950, i_10_1027, i_10_1029, i_10_1057, i_10_1117, i_10_1118, i_10_1122, i_10_1236, i_10_1243, i_10_1246, i_10_1247, i_10_1354, i_10_1396, i_10_1542, i_10_1575, i_10_1618, i_10_1648, i_10_1649, i_10_1691, i_10_1910, i_10_1945, i_10_1946, i_10_1959, i_10_1989, i_10_1992, i_10_2380, i_10_2454, i_10_2460, i_10_2511, i_10_2556, i_10_2557, i_10_2568, i_10_2608, i_10_2630, i_10_2631, i_10_2646, i_10_2657, i_10_2658, i_10_2659, i_10_2660, i_10_2710, i_10_2720, i_10_2727, i_10_2729, i_10_2829, i_10_2867, i_10_2881, i_10_2921, i_10_2923, i_10_3042, i_10_3045, i_10_3046, i_10_3072, i_10_3161, i_10_3229, i_10_3267, i_10_3269, i_10_3300, i_10_3336, i_10_3386, i_10_3440, i_10_3540, i_10_3549, i_10_3550, i_10_3551, i_10_3557, i_10_3620, i_10_3782, i_10_3848, i_10_3852, i_10_3981, i_10_4025, i_10_4026, i_10_4027, i_10_4118, i_10_4119, i_10_4125, i_10_4149, i_10_4151, i_10_4167, i_10_4191, i_10_4212, i_10_4213, i_10_4214, i_10_4290, i_10_4317, i_10_4565, i_10_4583, i_10_4584, o_10_10);
	kernel_10_11 k_10_11(i_10_89, i_10_172, i_10_174, i_10_319, i_10_322, i_10_391, i_10_443, i_10_460, i_10_562, i_10_753, i_10_960, i_10_1048, i_10_1049, i_10_1088, i_10_1168, i_10_1240, i_10_1432, i_10_1435, i_10_1439, i_10_1545, i_10_1582, i_10_1583, i_10_1627, i_10_1650, i_10_1651, i_10_1686, i_10_1687, i_10_1689, i_10_1690, i_10_1691, i_10_1816, i_10_2023, i_10_2029, i_10_2201, i_10_2203, i_10_2353, i_10_2355, i_10_2356, i_10_2357, i_10_2359, i_10_2453, i_10_2463, i_10_2468, i_10_2471, i_10_2506, i_10_2542, i_10_2661, i_10_2662, i_10_2679, i_10_2707, i_10_2720, i_10_2733, i_10_2735, i_10_2784, i_10_2785, i_10_2789, i_10_2824, i_10_2966, i_10_3046, i_10_3070, i_10_3075, i_10_3238, i_10_3279, i_10_3281, i_10_3316, i_10_3389, i_10_3392, i_10_3431, i_10_3469, i_10_3525, i_10_3541, i_10_3556, i_10_3609, i_10_3683, i_10_3723, i_10_3724, i_10_3725, i_10_3727, i_10_3728, i_10_3780, i_10_3838, i_10_3844, i_10_3846, i_10_3847, i_10_3848, i_10_3946, i_10_4119, i_10_4121, i_10_4126, i_10_4128, i_10_4129, i_10_4207, i_10_4281, i_10_4282, i_10_4283, i_10_4291, i_10_4563, i_10_4566, i_10_4567, i_10_4583, o_10_11);
	kernel_10_12 k_10_12(i_10_44, i_10_147, i_10_151, i_10_177, i_10_430, i_10_448, i_10_518, i_10_521, i_10_637, i_10_714, i_10_717, i_10_735, i_10_798, i_10_832, i_10_903, i_10_931, i_10_967, i_10_970, i_10_1087, i_10_1127, i_10_1165, i_10_1233, i_10_1273, i_10_1306, i_10_1307, i_10_1310, i_10_1535, i_10_1537, i_10_1580, i_10_1637, i_10_1641, i_10_1709, i_10_1768, i_10_1795, i_10_1820, i_10_1874, i_10_1922, i_10_2001, i_10_2004, i_10_2028, i_10_2032, i_10_2186, i_10_2212, i_10_2309, i_10_2310, i_10_2311, i_10_2353, i_10_2354, i_10_2356, i_10_2389, i_10_2390, i_10_2451, i_10_2461, i_10_2472, i_10_2518, i_10_2631, i_10_2678, i_10_2680, i_10_2705, i_10_2914, i_10_2919, i_10_2983, i_10_2987, i_10_3014, i_10_3200, i_10_3234, i_10_3235, i_10_3279, i_10_3280, i_10_3319, i_10_3391, i_10_3470, i_10_3472, i_10_3473, i_10_3495, i_10_3496, i_10_3522, i_10_3525, i_10_3540, i_10_3541, i_10_3584, i_10_3588, i_10_3650, i_10_3776, i_10_3788, i_10_3823, i_10_3854, i_10_4013, i_10_4028, i_10_4051, i_10_4054, i_10_4117, i_10_4118, i_10_4229, i_10_4269, i_10_4282, i_10_4287, i_10_4291, i_10_4435, i_10_4588, o_10_12);
	kernel_10_13 k_10_13(i_10_223, i_10_276, i_10_287, i_10_318, i_10_319, i_10_322, i_10_324, i_10_411, i_10_412, i_10_424, i_10_430, i_10_431, i_10_432, i_10_435, i_10_447, i_10_465, i_10_798, i_10_800, i_10_1249, i_10_1363, i_10_1365, i_10_1431, i_10_1437, i_10_1439, i_10_1546, i_10_1579, i_10_1581, i_10_1582, i_10_1626, i_10_1627, i_10_1653, i_10_1686, i_10_1687, i_10_1688, i_10_1724, i_10_1821, i_10_1822, i_10_1823, i_10_1911, i_10_1912, i_10_1995, i_10_1996, i_10_2005, i_10_2199, i_10_2452, i_10_2454, i_10_2466, i_10_2572, i_10_2604, i_10_2631, i_10_2632, i_10_2634, i_10_2635, i_10_2636, i_10_2705, i_10_2713, i_10_2722, i_10_2723, i_10_2730, i_10_2733, i_10_2734, i_10_2781, i_10_2826, i_10_2827, i_10_2828, i_10_2829, i_10_2830, i_10_2880, i_10_2883, i_10_2884, i_10_2885, i_10_3045, i_10_3070, i_10_3087, i_10_3151, i_10_3202, i_10_3268, i_10_3321, i_10_3387, i_10_3388, i_10_3543, i_10_3582, i_10_3613, i_10_3614, i_10_3616, i_10_3836, i_10_3837, i_10_3859, i_10_3912, i_10_3913, i_10_3978, i_10_3991, i_10_4057, i_10_4128, i_10_4129, i_10_4175, i_10_4281, i_10_4282, i_10_4283, i_10_4569, o_10_13);
	kernel_10_14 k_10_14(i_10_183, i_10_195, i_10_324, i_10_394, i_10_409, i_10_430, i_10_445, i_10_460, i_10_463, i_10_511, i_10_516, i_10_520, i_10_577, i_10_697, i_10_732, i_10_733, i_10_798, i_10_864, i_10_867, i_10_969, i_10_1098, i_10_1119, i_10_1120, i_10_1168, i_10_1239, i_10_1246, i_10_1551, i_10_1581, i_10_1620, i_10_1693, i_10_1696, i_10_1715, i_10_1756, i_10_1767, i_10_1789, i_10_1885, i_10_1908, i_10_1912, i_10_1948, i_10_1950, i_10_2085, i_10_2155, i_10_2334, i_10_2352, i_10_2442, i_10_2452, i_10_2453, i_10_2463, i_10_2481, i_10_2574, i_10_2577, i_10_2631, i_10_2634, i_10_2676, i_10_2680, i_10_2711, i_10_2830, i_10_2866, i_10_2868, i_10_2919, i_10_2922, i_10_2983, i_10_2984, i_10_3036, i_10_3047, i_10_3049, i_10_3198, i_10_3199, i_10_3277, i_10_3298, i_10_3312, i_10_3407, i_10_3540, i_10_3541, i_10_3609, i_10_3686, i_10_3688, i_10_3720, i_10_3724, i_10_3795, i_10_3921, i_10_3931, i_10_3964, i_10_3968, i_10_3981, i_10_3982, i_10_3984, i_10_3985, i_10_4155, i_10_4191, i_10_4192, i_10_4207, i_10_4269, i_10_4271, i_10_4273, i_10_4278, i_10_4279, i_10_4290, i_10_4291, i_10_4515, o_10_14);
	kernel_10_15 k_10_15(i_10_51, i_10_148, i_10_283, i_10_295, i_10_322, i_10_436, i_10_445, i_10_448, i_10_449, i_10_463, i_10_467, i_10_562, i_10_896, i_10_899, i_10_907, i_10_997, i_10_1033, i_10_1034, i_10_1051, i_10_1234, i_10_1249, i_10_1250, i_10_1446, i_10_1447, i_10_1619, i_10_1636, i_10_1637, i_10_1652, i_10_1684, i_10_1686, i_10_1687, i_10_1688, i_10_1690, i_10_1691, i_10_1808, i_10_1819, i_10_1823, i_10_1826, i_10_1910, i_10_1913, i_10_1960, i_10_2015, i_10_2158, i_10_2231, i_10_2353, i_10_2354, i_10_2355, i_10_2357, i_10_2365, i_10_2448, i_10_2456, i_10_2481, i_10_2482, i_10_2528, i_10_2535, i_10_2540, i_10_2546, i_10_2571, i_10_2572, i_10_2608, i_10_2632, i_10_2636, i_10_2654, i_10_2659, i_10_2662, i_10_2689, i_10_2708, i_10_2788, i_10_2832, i_10_2833, i_10_3038, i_10_3076, i_10_3196, i_10_3199, i_10_3200, i_10_3272, i_10_3274, i_10_3275, i_10_3278, i_10_3356, i_10_3384, i_10_3391, i_10_3392, i_10_3463, i_10_3527, i_10_3544, i_10_3721, i_10_3733, i_10_3859, i_10_3894, i_10_3905, i_10_3985, i_10_3986, i_10_3992, i_10_4030, i_10_4031, i_10_4118, i_10_4121, i_10_4154, i_10_4570, o_10_15);
	kernel_10_16 k_10_16(i_10_40, i_10_149, i_10_153, i_10_175, i_10_183, i_10_229, i_10_265, i_10_363, i_10_366, i_10_406, i_10_408, i_10_437, i_10_448, i_10_513, i_10_670, i_10_691, i_10_751, i_10_906, i_10_933, i_10_1029, i_10_1033, i_10_1038, i_10_1135, i_10_1137, i_10_1138, i_10_1139, i_10_1153, i_10_1157, i_10_1158, i_10_1164, i_10_1165, i_10_1218, i_10_1219, i_10_1238, i_10_1239, i_10_1264, i_10_1266, i_10_1267, i_10_1305, i_10_1308, i_10_1310, i_10_1311, i_10_1378, i_10_1399, i_10_1455, i_10_1552, i_10_1554, i_10_1632, i_10_1647, i_10_1815, i_10_1858, i_10_1872, i_10_1914, i_10_1948, i_10_1956, i_10_1998, i_10_2019, i_10_2020, i_10_2068, i_10_2391, i_10_2409, i_10_2505, i_10_2508, i_10_2568, i_10_2589, i_10_2605, i_10_2613, i_10_2634, i_10_2703, i_10_2704, i_10_2705, i_10_2706, i_10_2707, i_10_2713, i_10_2724, i_10_2725, i_10_2733, i_10_2985, i_10_2986, i_10_3234, i_10_3293, i_10_3397, i_10_3435, i_10_3455, i_10_3470, i_10_3498, i_10_3541, i_10_3667, i_10_3717, i_10_3720, i_10_3779, i_10_3789, i_10_3879, i_10_4116, i_10_4117, i_10_4120, i_10_4140, i_10_4278, i_10_4555, i_10_4570, o_10_16);
	kernel_10_17 k_10_17(i_10_37, i_10_49, i_10_68, i_10_128, i_10_155, i_10_244, i_10_282, i_10_286, i_10_406, i_10_407, i_10_438, i_10_441, i_10_443, i_10_463, i_10_464, i_10_824, i_10_959, i_10_994, i_10_1001, i_10_1109, i_10_1241, i_10_1248, i_10_1305, i_10_1306, i_10_1310, i_10_1313, i_10_1432, i_10_1579, i_10_1647, i_10_1648, i_10_1651, i_10_1684, i_10_1688, i_10_1795, i_10_1800, i_10_1913, i_10_1948, i_10_2196, i_10_2197, i_10_2234, i_10_2246, i_10_2352, i_10_2354, i_10_2407, i_10_2449, i_10_2455, i_10_2518, i_10_2534, i_10_2606, i_10_2628, i_10_2677, i_10_2706, i_10_2727, i_10_2730, i_10_2734, i_10_2832, i_10_2880, i_10_3040, i_10_3199, i_10_3232, i_10_3238, i_10_3271, i_10_3281, i_10_3384, i_10_3386, i_10_3387, i_10_3388, i_10_3389, i_10_3523, i_10_3611, i_10_3613, i_10_3614, i_10_3649, i_10_3650, i_10_3652, i_10_3684, i_10_3685, i_10_3781, i_10_3782, i_10_3784, i_10_3787, i_10_3788, i_10_3800, i_10_3834, i_10_3835, i_10_3844, i_10_3847, i_10_3856, i_10_3860, i_10_4027, i_10_4120, i_10_4123, i_10_4143, i_10_4170, i_10_4276, i_10_4285, i_10_4286, i_10_4288, i_10_4289, i_10_4372, o_10_17);
	kernel_10_18 k_10_18(i_10_28, i_10_171, i_10_174, i_10_175, i_10_176, i_10_261, i_10_267, i_10_390, i_10_393, i_10_409, i_10_410, i_10_411, i_10_412, i_10_441, i_10_442, i_10_446, i_10_718, i_10_793, i_10_796, i_10_960, i_10_1003, i_10_1005, i_10_1006, i_10_1026, i_10_1028, i_10_1036, i_10_1238, i_10_1242, i_10_1312, i_10_1431, i_10_1432, i_10_1434, i_10_1440, i_10_1539, i_10_1554, i_10_1575, i_10_1651, i_10_1652, i_10_1655, i_10_1688, i_10_1691, i_10_1819, i_10_1822, i_10_1824, i_10_1825, i_10_1947, i_10_1950, i_10_2001, i_10_2178, i_10_2179, i_10_2184, i_10_2185, i_10_2186, i_10_2355, i_10_2358, i_10_2410, i_10_2460, i_10_2466, i_10_2469, i_10_2565, i_10_2567, i_10_2605, i_10_2656, i_10_2724, i_10_2725, i_10_2731, i_10_2732, i_10_2735, i_10_2832, i_10_2883, i_10_2923, i_10_2987, i_10_3036, i_10_3042, i_10_3045, i_10_3069, i_10_3070, i_10_3095, i_10_3198, i_10_3202, i_10_3276, i_10_3388, i_10_3391, i_10_3467, i_10_3471, i_10_3522, i_10_3523, i_10_3525, i_10_3610, i_10_3780, i_10_3783, i_10_3788, i_10_3834, i_10_3838, i_10_3841, i_10_3855, i_10_3856, i_10_3913, i_10_4291, i_10_4292, o_10_18);
	kernel_10_19 k_10_19(i_10_219, i_10_220, i_10_221, i_10_269, i_10_282, i_10_316, i_10_320, i_10_329, i_10_431, i_10_436, i_10_445, i_10_446, i_10_464, i_10_467, i_10_518, i_10_752, i_10_799, i_10_853, i_10_854, i_10_899, i_10_956, i_10_1030, i_10_1032, i_10_1082, i_10_1123, i_10_1220, i_10_1249, i_10_1308, i_10_1309, i_10_1610, i_10_1618, i_10_1619, i_10_1822, i_10_1916, i_10_1997, i_10_2004, i_10_2021, i_10_2023, i_10_2203, i_10_2228, i_10_2231, i_10_2349, i_10_2350, i_10_2354, i_10_2365, i_10_2382, i_10_2460, i_10_2463, i_10_2464, i_10_2470, i_10_2472, i_10_2473, i_10_2634, i_10_2645, i_10_2678, i_10_2704, i_10_2723, i_10_2832, i_10_2833, i_10_2834, i_10_2886, i_10_2984, i_10_3050, i_10_3072, i_10_3196, i_10_3197, i_10_3278, i_10_3280, i_10_3283, i_10_3384, i_10_3387, i_10_3388, i_10_3469, i_10_3495, i_10_3496, i_10_3523, i_10_3544, i_10_3549, i_10_3651, i_10_3682, i_10_3684, i_10_3729, i_10_3732, i_10_3839, i_10_3842, i_10_3856, i_10_3859, i_10_3860, i_10_3895, i_10_3910, i_10_3913, i_10_3983, i_10_3988, i_10_4027, i_10_4029, i_10_4030, i_10_4216, i_10_4277, i_10_4283, i_10_4568, o_10_19);
	kernel_10_20 k_10_20(i_10_49, i_10_180, i_10_315, i_10_405, i_10_431, i_10_435, i_10_436, i_10_439, i_10_444, i_10_445, i_10_447, i_10_449, i_10_467, i_10_591, i_10_636, i_10_700, i_10_735, i_10_753, i_10_754, i_10_799, i_10_1038, i_10_1039, i_10_1040, i_10_1201, i_10_1236, i_10_1237, i_10_1238, i_10_1240, i_10_1552, i_10_1782, i_10_1821, i_10_1822, i_10_1824, i_10_2147, i_10_2155, i_10_2241, i_10_2244, i_10_2245, i_10_2307, i_10_2309, i_10_2310, i_10_2333, i_10_2334, i_10_2352, i_10_2388, i_10_2460, i_10_2470, i_10_2517, i_10_2542, i_10_2607, i_10_2633, i_10_2634, i_10_2635, i_10_2650, i_10_2651, i_10_2677, i_10_2703, i_10_2704, i_10_2718, i_10_2721, i_10_2730, i_10_2731, i_10_2732, i_10_2820, i_10_2830, i_10_2832, i_10_2919, i_10_3271, i_10_3273, i_10_3387, i_10_3388, i_10_3389, i_10_3500, i_10_3610, i_10_3614, i_10_3646, i_10_3649, i_10_3652, i_10_3684, i_10_3685, i_10_3783, i_10_3786, i_10_3838, i_10_3854, i_10_3856, i_10_3859, i_10_3881, i_10_3882, i_10_3982, i_10_4116, i_10_4117, i_10_4118, i_10_4119, i_10_4120, i_10_4188, i_10_4462, i_10_4485, i_10_4513, i_10_4516, i_10_4602, o_10_20);
	kernel_10_21 k_10_21(i_10_45, i_10_185, i_10_217, i_10_281, i_10_282, i_10_283, i_10_284, i_10_289, i_10_315, i_10_405, i_10_408, i_10_435, i_10_436, i_10_462, i_10_463, i_10_464, i_10_466, i_10_892, i_10_1028, i_10_1233, i_10_1240, i_10_1306, i_10_1307, i_10_1311, i_10_1363, i_10_1432, i_10_1444, i_10_1540, i_10_1543, i_10_1576, i_10_1577, i_10_1648, i_10_1651, i_10_1655, i_10_1675, i_10_1686, i_10_1687, i_10_1689, i_10_1690, i_10_1819, i_10_1989, i_10_1990, i_10_2334, i_10_2358, i_10_2359, i_10_2361, i_10_2362, i_10_2380, i_10_2457, i_10_2467, i_10_2631, i_10_2709, i_10_2710, i_10_2719, i_10_2826, i_10_2829, i_10_2830, i_10_2831, i_10_2834, i_10_2880, i_10_2881, i_10_2918, i_10_2920, i_10_2921, i_10_3034, i_10_3037, i_10_3043, i_10_3072, i_10_3075, i_10_3269, i_10_3277, i_10_3280, i_10_3324, i_10_3327, i_10_3392, i_10_3408, i_10_3409, i_10_3466, i_10_3469, i_10_3611, i_10_3785, i_10_3835, i_10_3838, i_10_3847, i_10_3848, i_10_3849, i_10_3856, i_10_3857, i_10_3892, i_10_4116, i_10_4120, i_10_4122, i_10_4125, i_10_4126, i_10_4212, i_10_4213, i_10_4267, i_10_4276, i_10_4566, i_10_4567, o_10_21);
	kernel_10_22 k_10_22(i_10_21, i_10_22, i_10_48, i_10_134, i_10_180, i_10_181, i_10_184, i_10_185, i_10_428, i_10_433, i_10_515, i_10_599, i_10_639, i_10_640, i_10_716, i_10_759, i_10_793, i_10_798, i_10_799, i_10_950, i_10_1000, i_10_1028, i_10_1131, i_10_1164, i_10_1171, i_10_1238, i_10_1246, i_10_1247, i_10_1312, i_10_1447, i_10_1453, i_10_1541, i_10_1607, i_10_1616, i_10_1632, i_10_1633, i_10_1786, i_10_1823, i_10_1826, i_10_1882, i_10_1909, i_10_1912, i_10_1992, i_10_2011, i_10_2012, i_10_2091, i_10_2162, i_10_2335, i_10_2349, i_10_2365, i_10_2383, i_10_2439, i_10_2441, i_10_2461, i_10_2578, i_10_2604, i_10_2608, i_10_2640, i_10_2649, i_10_2686, i_10_2711, i_10_2747, i_10_2828, i_10_2866, i_10_2885, i_10_2918, i_10_2922, i_10_2923, i_10_3083, i_10_3088, i_10_3107, i_10_3202, i_10_3226, i_10_3234, i_10_3439, i_10_3537, i_10_3538, i_10_3623, i_10_3650, i_10_3721, i_10_3786, i_10_3787, i_10_3788, i_10_3835, i_10_3836, i_10_3889, i_10_3892, i_10_3963, i_10_3964, i_10_4152, i_10_4157, i_10_4185, i_10_4186, i_10_4188, i_10_4190, i_10_4217, i_10_4287, i_10_4435, i_10_4457, i_10_4462, o_10_22);
	kernel_10_23 k_10_23(i_10_224, i_10_293, i_10_409, i_10_410, i_10_444, i_10_445, i_10_447, i_10_643, i_10_646, i_10_797, i_10_1000, i_10_1123, i_10_1172, i_10_1216, i_10_1264, i_10_1313, i_10_1348, i_10_1543, i_10_1578, i_10_1579, i_10_1580, i_10_1582, i_10_1583, i_10_1648, i_10_1724, i_10_1810, i_10_1821, i_10_1826, i_10_1991, i_10_1994, i_10_2023, i_10_2352, i_10_2354, i_10_2360, i_10_2363, i_10_2365, i_10_2366, i_10_2380, i_10_2381, i_10_2384, i_10_2453, i_10_2466, i_10_2656, i_10_2657, i_10_2700, i_10_2708, i_10_2711, i_10_2714, i_10_2717, i_10_2718, i_10_2719, i_10_2720, i_10_2723, i_10_2729, i_10_2730, i_10_2732, i_10_2734, i_10_2735, i_10_2828, i_10_2831, i_10_3038, i_10_3230, i_10_3287, i_10_3290, i_10_3301, i_10_3302, i_10_3384, i_10_3388, i_10_3389, i_10_3403, i_10_3406, i_10_3430, i_10_3461, i_10_3467, i_10_3520, i_10_3523, i_10_3524, i_10_3587, i_10_3611, i_10_3614, i_10_3650, i_10_3689, i_10_3728, i_10_3785, i_10_3852, i_10_3855, i_10_3857, i_10_3893, i_10_3923, i_10_3994, i_10_4118, i_10_4120, i_10_4121, i_10_4169, i_10_4271, i_10_4273, i_10_4275, i_10_4289, i_10_4461, i_10_4571, o_10_23);
	kernel_10_24 k_10_24(i_10_82, i_10_181, i_10_210, i_10_216, i_10_217, i_10_221, i_10_271, i_10_274, i_10_275, i_10_281, i_10_406, i_10_409, i_10_437, i_10_449, i_10_482, i_10_508, i_10_826, i_10_892, i_10_944, i_10_963, i_10_1060, i_10_1080, i_10_1117, i_10_1242, i_10_1243, i_10_1248, i_10_1249, i_10_1310, i_10_1354, i_10_1355, i_10_1359, i_10_1360, i_10_1575, i_10_1576, i_10_1603, i_10_1617, i_10_1688, i_10_1765, i_10_1786, i_10_1881, i_10_1903, i_10_1922, i_10_2020, i_10_2197, i_10_2331, i_10_2332, i_10_2367, i_10_2450, i_10_2502, i_10_2540, i_10_2631, i_10_2638, i_10_2646, i_10_2647, i_10_2704, i_10_2728, i_10_2862, i_10_2869, i_10_2872, i_10_2916, i_10_2919, i_10_2920, i_10_2953, i_10_3054, i_10_3195, i_10_3262, i_10_3384, i_10_3550, i_10_3610, i_10_3611, i_10_3720, i_10_3721, i_10_3846, i_10_3847, i_10_3848, i_10_3851, i_10_3856, i_10_3884, i_10_3888, i_10_3889, i_10_3915, i_10_3960, i_10_3961, i_10_3963, i_10_3964, i_10_4023, i_10_4024, i_10_4025, i_10_4118, i_10_4177, i_10_4185, i_10_4186, i_10_4188, i_10_4287, i_10_4325, i_10_4420, i_10_4428, i_10_4510, i_10_4527, i_10_4600, o_10_24);
	kernel_10_25 k_10_25(i_10_35, i_10_172, i_10_174, i_10_175, i_10_176, i_10_178, i_10_183, i_10_220, i_10_221, i_10_272, i_10_285, i_10_286, i_10_328, i_10_410, i_10_429, i_10_460, i_10_711, i_10_795, i_10_796, i_10_907, i_10_961, i_10_999, i_10_1006, i_10_1168, i_10_1169, i_10_1236, i_10_1244, i_10_1263, i_10_1580, i_10_1583, i_10_1654, i_10_1686, i_10_1689, i_10_1691, i_10_1821, i_10_1822, i_10_1823, i_10_1910, i_10_1913, i_10_2022, i_10_2349, i_10_2350, i_10_2351, i_10_2352, i_10_2353, i_10_2354, i_10_2379, i_10_2407, i_10_2409, i_10_2410, i_10_2451, i_10_2452, i_10_2453, i_10_2681, i_10_2703, i_10_2708, i_10_2711, i_10_2714, i_10_2722, i_10_2725, i_10_2733, i_10_2734, i_10_2735, i_10_2828, i_10_3036, i_10_3153, i_10_3165, i_10_3195, i_10_3196, i_10_3202, i_10_3231, i_10_3237, i_10_3279, i_10_3281, i_10_3325, i_10_3388, i_10_3613, i_10_3614, i_10_3616, i_10_3646, i_10_3649, i_10_3723, i_10_3724, i_10_3781, i_10_3838, i_10_3839, i_10_3846, i_10_3856, i_10_3857, i_10_3859, i_10_3883, i_10_3895, i_10_3913, i_10_3991, i_10_4120, i_10_4121, i_10_4129, i_10_4174, i_10_4269, i_10_4283, o_10_25);
	kernel_10_26 k_10_26(i_10_174, i_10_176, i_10_286, i_10_293, i_10_296, i_10_326, i_10_328, i_10_394, i_10_429, i_10_444, i_10_445, i_10_447, i_10_448, i_10_465, i_10_792, i_10_798, i_10_799, i_10_955, i_10_1002, i_10_1032, i_10_1034, i_10_1240, i_10_1241, i_10_1265, i_10_1305, i_10_1306, i_10_1309, i_10_1651, i_10_1819, i_10_1821, i_10_1826, i_10_1911, i_10_1989, i_10_1995, i_10_1996, i_10_2311, i_10_2349, i_10_2351, i_10_2357, i_10_2364, i_10_2452, i_10_2571, i_10_2655, i_10_2656, i_10_2657, i_10_2658, i_10_2659, i_10_2703, i_10_2704, i_10_2714, i_10_2727, i_10_2728, i_10_2730, i_10_2731, i_10_2732, i_10_2787, i_10_2788, i_10_2819, i_10_2884, i_10_2985, i_10_2987, i_10_3039, i_10_3045, i_10_3046, i_10_3048, i_10_3049, i_10_3075, i_10_3076, i_10_3091, i_10_3094, i_10_3195, i_10_3198, i_10_3271, i_10_3272, i_10_3298, i_10_3326, i_10_3405, i_10_3407, i_10_3408, i_10_3409, i_10_3472, i_10_3613, i_10_3646, i_10_3855, i_10_3857, i_10_3860, i_10_3983, i_10_3985, i_10_3986, i_10_4115, i_10_4116, i_10_4117, i_10_4128, i_10_4216, i_10_4269, i_10_4270, i_10_4271, i_10_4278, i_10_4288, i_10_4568, o_10_26);
	kernel_10_27 k_10_27(i_10_40, i_10_229, i_10_230, i_10_271, i_10_272, i_10_319, i_10_423, i_10_427, i_10_430, i_10_433, i_10_449, i_10_464, i_10_543, i_10_741, i_10_751, i_10_877, i_10_1027, i_10_1054, i_10_1111, i_10_1252, i_10_1265, i_10_1311, i_10_1348, i_10_1354, i_10_1361, i_10_1364, i_10_1416, i_10_1492, i_10_1545, i_10_1552, i_10_1554, i_10_1579, i_10_1642, i_10_1650, i_10_1651, i_10_1652, i_10_1888, i_10_1909, i_10_1948, i_10_2161, i_10_2167, i_10_2168, i_10_2185, i_10_2186, i_10_2453, i_10_2458, i_10_2516, i_10_2641, i_10_2658, i_10_2663, i_10_2731, i_10_2732, i_10_2821, i_10_2865, i_10_2869, i_10_2885, i_10_2912, i_10_2917, i_10_2919, i_10_2924, i_10_2957, i_10_2983, i_10_3040, i_10_3201, i_10_3203, i_10_3270, i_10_3307, i_10_3325, i_10_3469, i_10_3472, i_10_3521, i_10_3523, i_10_3526, i_10_3540, i_10_3541, i_10_3544, i_10_3614, i_10_3718, i_10_3781, i_10_3786, i_10_3828, i_10_3852, i_10_3890, i_10_3910, i_10_3947, i_10_3988, i_10_3990, i_10_4008, i_10_4013, i_10_4054, i_10_4116, i_10_4117, i_10_4149, i_10_4152, i_10_4154, i_10_4190, i_10_4272, i_10_4285, i_10_4570, i_10_4595, o_10_27);
	kernel_10_28 k_10_28(i_10_89, i_10_171, i_10_221, i_10_222, i_10_223, i_10_224, i_10_285, i_10_287, i_10_318, i_10_319, i_10_323, i_10_432, i_10_433, i_10_444, i_10_445, i_10_446, i_10_449, i_10_506, i_10_719, i_10_752, i_10_795, i_10_1037, i_10_1236, i_10_1238, i_10_1242, i_10_1243, i_10_1244, i_10_1246, i_10_1647, i_10_1650, i_10_1651, i_10_1652, i_10_1653, i_10_1819, i_10_1821, i_10_1824, i_10_1825, i_10_1989, i_10_2338, i_10_2359, i_10_2362, i_10_2467, i_10_2468, i_10_2629, i_10_2631, i_10_2633, i_10_2635, i_10_2645, i_10_2657, i_10_2658, i_10_2659, i_10_2660, i_10_2678, i_10_2720, i_10_2785, i_10_2788, i_10_2821, i_10_2888, i_10_2919, i_10_2920, i_10_2922, i_10_2924, i_10_2981, i_10_3033, i_10_3034, i_10_3150, i_10_3151, i_10_3152, i_10_3154, i_10_3155, i_10_3156, i_10_3157, i_10_3195, i_10_3274, i_10_3278, i_10_3385, i_10_3408, i_10_3587, i_10_3685, i_10_3780, i_10_3782, i_10_3788, i_10_3834, i_10_3835, i_10_3836, i_10_3839, i_10_3847, i_10_3848, i_10_3853, i_10_3854, i_10_3856, i_10_3857, i_10_3860, i_10_4116, i_10_4129, i_10_4565, i_10_4567, i_10_4568, i_10_4570, i_10_4571, o_10_28);
	kernel_10_29 k_10_29(i_10_174, i_10_179, i_10_223, i_10_243, i_10_256, i_10_257, i_10_286, i_10_318, i_10_319, i_10_321, i_10_323, i_10_387, i_10_435, i_10_436, i_10_443, i_10_447, i_10_561, i_10_907, i_10_997, i_10_1003, i_10_1004, i_10_1040, i_10_1042, i_10_1043, i_10_1263, i_10_1308, i_10_1344, i_10_1347, i_10_1435, i_10_1444, i_10_1542, i_10_1543, i_10_1544, i_10_1576, i_10_1578, i_10_1579, i_10_1580, i_10_1582, i_10_1611, i_10_1636, i_10_1654, i_10_1689, i_10_1691, i_10_1768, i_10_1816, i_10_1821, i_10_1822, i_10_1913, i_10_1956, i_10_1984, i_10_2003, i_10_2019, i_10_2083, i_10_2291, i_10_2436, i_10_2451, i_10_2453, i_10_2514, i_10_2515, i_10_2631, i_10_2656, i_10_2703, i_10_2704, i_10_2716, i_10_2826, i_10_2882, i_10_2920, i_10_2960, i_10_3036, i_10_3277, i_10_3289, i_10_3298, i_10_3431, i_10_3473, i_10_3541, i_10_3544, i_10_3614, i_10_3649, i_10_3729, i_10_3784, i_10_3786, i_10_3787, i_10_3837, i_10_3848, i_10_3856, i_10_3912, i_10_3946, i_10_3982, i_10_4114, i_10_4115, i_10_4171, i_10_4172, i_10_4175, i_10_4233, i_10_4234, i_10_4279, i_10_4459, i_10_4462, i_10_4568, i_10_4571, o_10_29);
	kernel_10_30 k_10_30(i_10_86, i_10_88, i_10_89, i_10_280, i_10_284, i_10_330, i_10_393, i_10_394, i_10_395, i_10_413, i_10_431, i_10_437, i_10_459, i_10_462, i_10_463, i_10_464, i_10_700, i_10_996, i_10_1033, i_10_1039, i_10_1041, i_10_1168, i_10_1237, i_10_1245, i_10_1246, i_10_1247, i_10_1248, i_10_1249, i_10_1250, i_10_1313, i_10_1367, i_10_1384, i_10_1385, i_10_1582, i_10_1649, i_10_1716, i_10_1717, i_10_1735, i_10_1768, i_10_1769, i_10_1823, i_10_1912, i_10_1913, i_10_2005, i_10_2006, i_10_2201, i_10_2350, i_10_2354, i_10_2355, i_10_2356, i_10_2357, i_10_2361, i_10_2383, i_10_2438, i_10_2449, i_10_2451, i_10_2452, i_10_2455, i_10_2456, i_10_2516, i_10_2653, i_10_2681, i_10_2728, i_10_2918, i_10_2920, i_10_3041, i_10_3043, i_10_3076, i_10_3094, i_10_3200, i_10_3270, i_10_3280, i_10_3386, i_10_3387, i_10_3544, i_10_3611, i_10_3612, i_10_3613, i_10_3614, i_10_3615, i_10_3617, i_10_3781, i_10_3783, i_10_3787, i_10_3788, i_10_3836, i_10_3837, i_10_3838, i_10_3839, i_10_3846, i_10_3855, i_10_3856, i_10_3857, i_10_3886, i_10_3887, i_10_4120, i_10_4130, i_10_4219, i_10_4291, i_10_4292, o_10_30);
	kernel_10_31 k_10_31(i_10_32, i_10_88, i_10_133, i_10_151, i_10_266, i_10_349, i_10_364, i_10_393, i_10_394, i_10_431, i_10_464, i_10_465, i_10_466, i_10_566, i_10_591, i_10_592, i_10_673, i_10_674, i_10_750, i_10_754, i_10_770, i_10_798, i_10_952, i_10_953, i_10_976, i_10_996, i_10_1033, i_10_1052, i_10_1059, i_10_1235, i_10_1236, i_10_1238, i_10_1241, i_10_1312, i_10_1358, i_10_1382, i_10_1457, i_10_1491, i_10_1619, i_10_1822, i_10_1867, i_10_1906, i_10_1912, i_10_1913, i_10_1914, i_10_1952, i_10_1957, i_10_1958, i_10_1960, i_10_1987, i_10_2095, i_10_2275, i_10_2276, i_10_2362, i_10_2465, i_10_2481, i_10_2508, i_10_2516, i_10_2572, i_10_2644, i_10_2661, i_10_2662, i_10_2678, i_10_2712, i_10_2744, i_10_2782, i_10_2786, i_10_2914, i_10_2916, i_10_2948, i_10_2956, i_10_2960, i_10_3093, i_10_3175, i_10_3176, i_10_3198, i_10_3199, i_10_3362, i_10_3446, i_10_3451, i_10_3470, i_10_3472, i_10_3473, i_10_3495, i_10_3508, i_10_3614, i_10_3622, i_10_3642, i_10_3643, i_10_3649, i_10_3652, i_10_3858, i_10_3860, i_10_3885, i_10_4056, i_10_4057, i_10_4058, i_10_4129, i_10_4287, i_10_4526, o_10_31);
	kernel_10_32 k_10_32(i_10_82, i_10_217, i_10_263, i_10_283, i_10_285, i_10_288, i_10_289, i_10_318, i_10_319, i_10_320, i_10_322, i_10_323, i_10_390, i_10_464, i_10_497, i_10_558, i_10_559, i_10_640, i_10_755, i_10_798, i_10_896, i_10_1000, i_10_1007, i_10_1027, i_10_1030, i_10_1234, i_10_1236, i_10_1308, i_10_1454, i_10_1575, i_10_1578, i_10_1579, i_10_1655, i_10_1691, i_10_1767, i_10_1819, i_10_1823, i_10_1909, i_10_1989, i_10_1993, i_10_2153, i_10_2196, i_10_2200, i_10_2297, i_10_2361, i_10_2364, i_10_2448, i_10_2514, i_10_2558, i_10_2566, i_10_2603, i_10_2631, i_10_2632, i_10_2647, i_10_2702, i_10_2711, i_10_2719, i_10_2723, i_10_2728, i_10_2730, i_10_2827, i_10_2831, i_10_2888, i_10_2917, i_10_2921, i_10_3073, i_10_3160, i_10_3234, i_10_3276, i_10_3385, i_10_3388, i_10_3523, i_10_3541, i_10_3543, i_10_3558, i_10_3565, i_10_3613, i_10_3720, i_10_3721, i_10_3785, i_10_3852, i_10_3889, i_10_3986, i_10_4023, i_10_4024, i_10_4096, i_10_4117, i_10_4119, i_10_4122, i_10_4123, i_10_4126, i_10_4153, i_10_4167, i_10_4168, i_10_4170, i_10_4171, i_10_4174, i_10_4275, i_10_4285, i_10_4571, o_10_32);
	kernel_10_33 k_10_33(i_10_279, i_10_441, i_10_442, i_10_445, i_10_446, i_10_469, i_10_590, i_10_733, i_10_736, i_10_737, i_10_784, i_10_901, i_10_932, i_10_1031, i_10_1043, i_10_1120, i_10_1240, i_10_1249, i_10_1343, i_10_1391, i_10_1552, i_10_1683, i_10_1685, i_10_1690, i_10_1765, i_10_1766, i_10_1822, i_10_1888, i_10_1909, i_10_1912, i_10_1913, i_10_2243, i_10_2380, i_10_2462, i_10_2464, i_10_2476, i_10_2514, i_10_2542, i_10_2543, i_10_2571, i_10_2635, i_10_2644, i_10_2645, i_10_2653, i_10_2654, i_10_2663, i_10_2701, i_10_2710, i_10_2719, i_10_2727, i_10_2728, i_10_2729, i_10_2731, i_10_2732, i_10_2734, i_10_2737, i_10_2820, i_10_2831, i_10_2920, i_10_2923, i_10_2983, i_10_3033, i_10_3048, i_10_3076, i_10_3114, i_10_3201, i_10_3202, i_10_3279, i_10_3352, i_10_3353, i_10_3356, i_10_3390, i_10_3391, i_10_3392, i_10_3522, i_10_3538, i_10_3551, i_10_3612, i_10_3614, i_10_3616, i_10_3800, i_10_3839, i_10_3841, i_10_3859, i_10_3860, i_10_3887, i_10_3923, i_10_3981, i_10_4124, i_10_4154, i_10_4156, i_10_4183, i_10_4238, i_10_4270, i_10_4273, i_10_4288, i_10_4459, i_10_4568, i_10_4570, i_10_4594, o_10_33);
	kernel_10_34 k_10_34(i_10_14, i_10_41, i_10_175, i_10_176, i_10_260, i_10_266, i_10_320, i_10_388, i_10_429, i_10_500, i_10_508, i_10_509, i_10_559, i_10_714, i_10_718, i_10_866, i_10_956, i_10_993, i_10_1055, i_10_1112, i_10_1115, i_10_1207, i_10_1211, i_10_1220, i_10_1236, i_10_1301, i_10_1360, i_10_1366, i_10_1379, i_10_1380, i_10_1541, i_10_1544, i_10_1621, i_10_1634, i_10_1650, i_10_1685, i_10_1687, i_10_1691, i_10_1733, i_10_1802, i_10_1877, i_10_1920, i_10_1921, i_10_1981, i_10_1985, i_10_2003, i_10_2027, i_10_2030, i_10_2036, i_10_2089, i_10_2204, i_10_2341, i_10_2359, i_10_2372, i_10_2383, i_10_2467, i_10_2471, i_10_2558, i_10_2576, i_10_2596, i_10_2734, i_10_2836, i_10_2839, i_10_2849, i_10_2851, i_10_2864, i_10_2867, i_10_2963, i_10_2966, i_10_2972, i_10_2975, i_10_3223, i_10_3313, i_10_3352, i_10_3353, i_10_3388, i_10_3466, i_10_3485, i_10_3506, i_10_3519, i_10_3541, i_10_3542, i_10_3545, i_10_3611, i_10_3794, i_10_3841, i_10_3842, i_10_3856, i_10_3908, i_10_3943, i_10_4027, i_10_4028, i_10_4118, i_10_4127, i_10_4148, i_10_4153, i_10_4169, i_10_4205, i_10_4287, i_10_4395, o_10_34);
	kernel_10_35 k_10_35(i_10_174, i_10_176, i_10_407, i_10_409, i_10_443, i_10_520, i_10_697, i_10_798, i_10_799, i_10_956, i_10_958, i_10_998, i_10_1032, i_10_1246, i_10_1248, i_10_1249, i_10_1250, i_10_1308, i_10_1309, i_10_1310, i_10_1311, i_10_1432, i_10_1439, i_10_1552, i_10_1619, i_10_1650, i_10_1651, i_10_1687, i_10_1690, i_10_1691, i_10_1821, i_10_1822, i_10_1825, i_10_1996, i_10_2021, i_10_2023, i_10_2201, i_10_2365, i_10_2366, i_10_2451, i_10_2452, i_10_2463, i_10_2464, i_10_2470, i_10_2473, i_10_2514, i_10_2571, i_10_2702, i_10_2705, i_10_2711, i_10_2722, i_10_2725, i_10_2829, i_10_2832, i_10_2833, i_10_2920, i_10_2923, i_10_2924, i_10_3072, i_10_3074, i_10_3075, i_10_3112, i_10_3199, i_10_3270, i_10_3273, i_10_3277, i_10_3284, i_10_3386, i_10_3407, i_10_3408, i_10_3586, i_10_3609, i_10_3612, i_10_3613, i_10_3614, i_10_3615, i_10_3732, i_10_3733, i_10_3734, i_10_3780, i_10_3781, i_10_3782, i_10_3786, i_10_3787, i_10_3788, i_10_3841, i_10_3856, i_10_4029, i_10_4114, i_10_4116, i_10_4125, i_10_4130, i_10_4216, i_10_4217, i_10_4218, i_10_4269, i_10_4275, i_10_4290, i_10_4564, i_10_4565, o_10_35);
	kernel_10_36 k_10_36(i_10_32, i_10_34, i_10_173, i_10_224, i_10_245, i_10_247, i_10_248, i_10_253, i_10_254, i_10_260, i_10_266, i_10_434, i_10_496, i_10_542, i_10_716, i_10_717, i_10_793, i_10_795, i_10_799, i_10_901, i_10_956, i_10_1030, i_10_1234, i_10_1236, i_10_1237, i_10_1238, i_10_1246, i_10_1247, i_10_1310, i_10_1325, i_10_1349, i_10_1435, i_10_1436, i_10_1437, i_10_1439, i_10_1543, i_10_1579, i_10_1580, i_10_1583, i_10_1653, i_10_1654, i_10_1655, i_10_1685, i_10_1686, i_10_1688, i_10_1689, i_10_1690, i_10_1909, i_10_1937, i_10_1948, i_10_1949, i_10_1954, i_10_2365, i_10_2387, i_10_2449, i_10_2454, i_10_2474, i_10_2477, i_10_2511, i_10_2531, i_10_2532, i_10_2540, i_10_2601, i_10_2660, i_10_2661, i_10_2730, i_10_2735, i_10_2881, i_10_2885, i_10_2918, i_10_3072, i_10_3197, i_10_3199, i_10_3201, i_10_3233, i_10_3281, i_10_3295, i_10_3332, i_10_3341, i_10_3493, i_10_3522, i_10_3523, i_10_3545, i_10_3586, i_10_3611, i_10_3646, i_10_3733, i_10_3784, i_10_3809, i_10_3841, i_10_3842, i_10_3883, i_10_3983, i_10_3997, i_10_4007, i_10_4116, i_10_4126, i_10_4367, i_10_4385, i_10_4585, o_10_36);
	kernel_10_37 k_10_37(i_10_176, i_10_251, i_10_282, i_10_283, i_10_284, i_10_289, i_10_320, i_10_329, i_10_425, i_10_434, i_10_442, i_10_458, i_10_460, i_10_461, i_10_464, i_10_749, i_10_755, i_10_792, i_10_796, i_10_965, i_10_1238, i_10_1239, i_10_1242, i_10_1243, i_10_1250, i_10_1310, i_10_1575, i_10_1576, i_10_1655, i_10_1681, i_10_1686, i_10_1687, i_10_1688, i_10_1768, i_10_1819, i_10_1823, i_10_1824, i_10_1990, i_10_1991, i_10_2197, i_10_2351, i_10_2353, i_10_2354, i_10_2359, i_10_2361, i_10_2362, i_10_2363, i_10_2449, i_10_2452, i_10_2453, i_10_2467, i_10_2468, i_10_2474, i_10_2632, i_10_2633, i_10_2657, i_10_2674, i_10_2710, i_10_2782, i_10_2783, i_10_2830, i_10_2919, i_10_3043, i_10_3044, i_10_3088, i_10_3151, i_10_3199, i_10_3271, i_10_3273, i_10_3277, i_10_3388, i_10_3406, i_10_3409, i_10_3467, i_10_3496, i_10_3550, i_10_3587, i_10_3610, i_10_3617, i_10_3648, i_10_3785, i_10_3786, i_10_3838, i_10_3850, i_10_3853, i_10_3856, i_10_3857, i_10_3858, i_10_3888, i_10_3889, i_10_3949, i_10_3991, i_10_4050, i_10_4115, i_10_4117, i_10_4121, i_10_4267, i_10_4288, i_10_4289, i_10_4568, o_10_37);
	kernel_10_38 k_10_38(i_10_125, i_10_172, i_10_173, i_10_174, i_10_175, i_10_222, i_10_224, i_10_269, i_10_393, i_10_394, i_10_405, i_10_409, i_10_410, i_10_413, i_10_429, i_10_430, i_10_431, i_10_433, i_10_439, i_10_440, i_10_445, i_10_447, i_10_460, i_10_462, i_10_566, i_10_957, i_10_1006, i_10_1241, i_10_1309, i_10_1448, i_10_1550, i_10_1556, i_10_1637, i_10_1649, i_10_1651, i_10_1652, i_10_1653, i_10_1654, i_10_1655, i_10_1823, i_10_1825, i_10_1826, i_10_2006, i_10_2351, i_10_2354, i_10_2355, i_10_2356, i_10_2357, i_10_2358, i_10_2366, i_10_2448, i_10_2458, i_10_2572, i_10_2629, i_10_2632, i_10_2681, i_10_2700, i_10_2705, i_10_2706, i_10_2707, i_10_2708, i_10_2716, i_10_2718, i_10_2721, i_10_2723, i_10_2725, i_10_2728, i_10_2730, i_10_2731, i_10_2732, i_10_2735, i_10_2832, i_10_2833, i_10_2834, i_10_2881, i_10_2884, i_10_2985, i_10_3076, i_10_3087, i_10_3091, i_10_3093, i_10_3094, i_10_3095, i_10_3155, i_10_3198, i_10_3281, i_10_3391, i_10_3408, i_10_3611, i_10_3612, i_10_3615, i_10_3811, i_10_3835, i_10_3838, i_10_3839, i_10_3853, i_10_4120, i_10_4126, i_10_4127, i_10_4128, o_10_38);
	kernel_10_39 k_10_39(i_10_172, i_10_174, i_10_176, i_10_260, i_10_268, i_10_269, i_10_284, i_10_328, i_10_329, i_10_394, i_10_408, i_10_409, i_10_410, i_10_425, i_10_436, i_10_510, i_10_514, i_10_794, i_10_796, i_10_797, i_10_798, i_10_799, i_10_800, i_10_1006, i_10_1029, i_10_1261, i_10_1264, i_10_1308, i_10_1309, i_10_1438, i_10_1439, i_10_1546, i_10_1628, i_10_1651, i_10_1655, i_10_1691, i_10_1727, i_10_1821, i_10_1822, i_10_1823, i_10_1825, i_10_1912, i_10_1996, i_10_2254, i_10_2364, i_10_2451, i_10_2461, i_10_2463, i_10_2470, i_10_2473, i_10_2573, i_10_2634, i_10_2635, i_10_2636, i_10_2659, i_10_2704, i_10_2717, i_10_2720, i_10_2722, i_10_2723, i_10_2725, i_10_2730, i_10_2731, i_10_2826, i_10_2830, i_10_2832, i_10_2884, i_10_2885, i_10_3077, i_10_3087, i_10_3088, i_10_3153, i_10_3195, i_10_3196, i_10_3197, i_10_3200, i_10_3280, i_10_3329, i_10_3388, i_10_3389, i_10_3409, i_10_3473, i_10_3586, i_10_3610, i_10_3611, i_10_3614, i_10_3616, i_10_3648, i_10_3651, i_10_3652, i_10_3860, i_10_4126, i_10_4271, i_10_4289, i_10_4564, i_10_4565, i_10_4567, i_10_4568, i_10_4570, i_10_4571, o_10_39);
	kernel_10_40 k_10_40(i_10_118, i_10_171, i_10_172, i_10_175, i_10_216, i_10_217, i_10_218, i_10_220, i_10_221, i_10_224, i_10_243, i_10_244, i_10_245, i_10_280, i_10_329, i_10_390, i_10_405, i_10_406, i_10_409, i_10_447, i_10_711, i_10_712, i_10_799, i_10_898, i_10_967, i_10_991, i_10_1029, i_10_1030, i_10_1233, i_10_1241, i_10_1306, i_10_1434, i_10_1441, i_10_1648, i_10_1649, i_10_1651, i_10_1683, i_10_1821, i_10_1824, i_10_1990, i_10_2351, i_10_2353, i_10_2354, i_10_2363, i_10_2451, i_10_2473, i_10_2628, i_10_2632, i_10_2635, i_10_2654, i_10_2656, i_10_2709, i_10_2717, i_10_2718, i_10_2735, i_10_2826, i_10_2827, i_10_2831, i_10_2832, i_10_2833, i_10_2834, i_10_2920, i_10_2921, i_10_2924, i_10_2986, i_10_3034, i_10_3151, i_10_3152, i_10_3153, i_10_3162, i_10_3163, i_10_3198, i_10_3322, i_10_3329, i_10_3389, i_10_3406, i_10_3466, i_10_3472, i_10_3547, i_10_3610, i_10_3611, i_10_3613, i_10_3647, i_10_3733, i_10_3782, i_10_3837, i_10_3839, i_10_3856, i_10_3912, i_10_3983, i_10_4113, i_10_4114, i_10_4115, i_10_4116, i_10_4117, i_10_4129, i_10_4271, i_10_4287, i_10_4288, i_10_4289, o_10_40);
	kernel_10_41 k_10_41(i_10_27, i_10_68, i_10_86, i_10_103, i_10_176, i_10_178, i_10_215, i_10_224, i_10_248, i_10_425, i_10_562, i_10_565, i_10_566, i_10_586, i_10_824, i_10_960, i_10_989, i_10_1000, i_10_1001, i_10_1004, i_10_1101, i_10_1223, i_10_1238, i_10_1240, i_10_1349, i_10_1367, i_10_1439, i_10_1544, i_10_1547, i_10_1583, i_10_1651, i_10_1652, i_10_1687, i_10_1715, i_10_1766, i_10_1772, i_10_1778, i_10_1988, i_10_1991, i_10_1997, i_10_2000, i_10_2006, i_10_2023, i_10_2033, i_10_2348, i_10_2449, i_10_2453, i_10_2509, i_10_2510, i_10_2539, i_10_2567, i_10_2570, i_10_2571, i_10_2609, i_10_2636, i_10_2641, i_10_2644, i_10_2645, i_10_2720, i_10_2744, i_10_2834, i_10_2848, i_10_2849, i_10_2851, i_10_2966, i_10_2968, i_10_2999, i_10_3002, i_10_3041, i_10_3071, i_10_3074, i_10_3230, i_10_3238, i_10_3299, i_10_3307, i_10_3308, i_10_3409, i_10_3470, i_10_3506, i_10_3544, i_10_3545, i_10_3611, i_10_3797, i_10_3852, i_10_3853, i_10_3856, i_10_3923, i_10_3944, i_10_3989, i_10_4027, i_10_4129, i_10_4130, i_10_4148, i_10_4175, i_10_4217, i_10_4237, i_10_4238, i_10_4436, i_10_4461, i_10_4463, o_10_41);
	kernel_10_42 k_10_42(i_10_30, i_10_34, i_10_117, i_10_256, i_10_260, i_10_390, i_10_391, i_10_395, i_10_565, i_10_714, i_10_717, i_10_800, i_10_954, i_10_955, i_10_956, i_10_957, i_10_958, i_10_959, i_10_1030, i_10_1235, i_10_1245, i_10_1366, i_10_1439, i_10_1445, i_10_1450, i_10_1576, i_10_1579, i_10_1582, i_10_1619, i_10_1653, i_10_1691, i_10_1823, i_10_1826, i_10_2029, i_10_2030, i_10_2086, i_10_2197, i_10_2200, i_10_2201, i_10_2352, i_10_2353, i_10_2357, i_10_2383, i_10_2470, i_10_2536, i_10_2608, i_10_2614, i_10_2615, i_10_2632, i_10_2705, i_10_2707, i_10_2725, i_10_2869, i_10_3037, i_10_3039, i_10_3072, i_10_3196, i_10_3201, i_10_3202, i_10_3270, i_10_3391, i_10_3408, i_10_3469, i_10_3590, i_10_3612, i_10_3616, i_10_3617, i_10_3645, i_10_3646, i_10_3647, i_10_3649, i_10_3650, i_10_3651, i_10_3652, i_10_3653, i_10_3726, i_10_3729, i_10_3783, i_10_3784, i_10_3785, i_10_3786, i_10_3787, i_10_3788, i_10_3811, i_10_3837, i_10_3843, i_10_3844, i_10_3847, i_10_3856, i_10_3857, i_10_3914, i_10_4012, i_10_4116, i_10_4117, i_10_4118, i_10_4119, i_10_4120, i_10_4267, i_10_4564, i_10_4565, o_10_42);
	kernel_10_43 k_10_43(i_10_27, i_10_28, i_10_48, i_10_117, i_10_118, i_10_121, i_10_218, i_10_315, i_10_317, i_10_388, i_10_390, i_10_391, i_10_445, i_10_463, i_10_748, i_10_892, i_10_946, i_10_956, i_10_958, i_10_1162, i_10_1234, i_10_1237, i_10_1261, i_10_1305, i_10_1309, i_10_1354, i_10_1362, i_10_1377, i_10_1445, i_10_1451, i_10_1576, i_10_1611, i_10_1613, i_10_1640, i_10_1732, i_10_1804, i_10_1820, i_10_1821, i_10_1873, i_10_1882, i_10_1899, i_10_1915, i_10_1917, i_10_1918, i_10_1944, i_10_1946, i_10_1991, i_10_2081, i_10_2155, i_10_2179, i_10_2180, i_10_2241, i_10_2358, i_10_2380, i_10_2468, i_10_2504, i_10_2629, i_10_2630, i_10_2631, i_10_2781, i_10_2782, i_10_2818, i_10_2819, i_10_2881, i_10_2882, i_10_3036, i_10_3038, i_10_3073, i_10_3281, i_10_3430, i_10_3465, i_10_3537, i_10_3582, i_10_3614, i_10_3645, i_10_3646, i_10_3647, i_10_3649, i_10_3650, i_10_3782, i_10_3784, i_10_3785, i_10_3842, i_10_3979, i_10_4050, i_10_4115, i_10_4123, i_10_4126, i_10_4217, i_10_4220, i_10_4261, i_10_4268, i_10_4277, i_10_4279, i_10_4292, i_10_4302, i_10_4527, i_10_4528, i_10_4529, i_10_4583, o_10_43);
	kernel_10_44 k_10_44(i_10_41, i_10_45, i_10_73, i_10_148, i_10_149, i_10_188, i_10_286, i_10_296, i_10_316, i_10_319, i_10_372, i_10_438, i_10_448, i_10_463, i_10_501, i_10_502, i_10_724, i_10_752, i_10_826, i_10_844, i_10_934, i_10_1036, i_10_1083, i_10_1085, i_10_1088, i_10_1166, i_10_1268, i_10_1307, i_10_1327, i_10_1338, i_10_1354, i_10_1534, i_10_1545, i_10_1555, i_10_1616, i_10_1655, i_10_1686, i_10_1689, i_10_1821, i_10_1872, i_10_1909, i_10_1910, i_10_1911, i_10_1914, i_10_1918, i_10_1958, i_10_1986, i_10_2093, i_10_2157, i_10_2166, i_10_2245, i_10_2246, i_10_2284, i_10_2352, i_10_2357, i_10_2380, i_10_2491, i_10_2560, i_10_2563, i_10_2569, i_10_2613, i_10_2629, i_10_2678, i_10_2697, i_10_2731, i_10_2734, i_10_2782, i_10_2865, i_10_2960, i_10_2993, i_10_3011, i_10_3012, i_10_3034, i_10_3036, i_10_3040, i_10_3070, i_10_3084, i_10_3091, i_10_3235, i_10_3264, i_10_3308, i_10_3317, i_10_3433, i_10_3436, i_10_3471, i_10_3540, i_10_3541, i_10_3617, i_10_3624, i_10_3641, i_10_3668, i_10_3853, i_10_3882, i_10_3892, i_10_4073, i_10_4157, i_10_4267, i_10_4534, i_10_4535, i_10_4565, o_10_44);
	kernel_10_45 k_10_45(i_10_30, i_10_33, i_10_34, i_10_121, i_10_123, i_10_124, i_10_132, i_10_146, i_10_157, i_10_183, i_10_184, i_10_185, i_10_248, i_10_269, i_10_317, i_10_320, i_10_431, i_10_444, i_10_449, i_10_462, i_10_466, i_10_758, i_10_921, i_10_958, i_10_1003, i_10_1005, i_10_1013, i_10_1015, i_10_1029, i_10_1048, i_10_1050, i_10_1308, i_10_1365, i_10_1370, i_10_1383, i_10_1500, i_10_1546, i_10_1579, i_10_1612, i_10_1613, i_10_1617, i_10_1651, i_10_1733, i_10_1767, i_10_1768, i_10_1906, i_10_1911, i_10_1912, i_10_1913, i_10_1942, i_10_1950, i_10_1951, i_10_1956, i_10_1957, i_10_1959, i_10_1981, i_10_2000, i_10_2038, i_10_2041, i_10_2094, i_10_2201, i_10_2562, i_10_2570, i_10_2659, i_10_2660, i_10_2721, i_10_2725, i_10_2787, i_10_2833, i_10_2834, i_10_2883, i_10_2921, i_10_2990, i_10_3012, i_10_3013, i_10_3202, i_10_3298, i_10_3299, i_10_3326, i_10_3392, i_10_3473, i_10_3558, i_10_3589, i_10_3617, i_10_3624, i_10_3840, i_10_3841, i_10_3855, i_10_3858, i_10_3945, i_10_3980, i_10_3995, i_10_4053, i_10_4116, i_10_4183, i_10_4288, i_10_4299, i_10_4547, i_10_4569, i_10_4593, o_10_45);
	kernel_10_46 k_10_46(i_10_38, i_10_149, i_10_155, i_10_171, i_10_172, i_10_178, i_10_218, i_10_244, i_10_245, i_10_248, i_10_280, i_10_286, i_10_287, i_10_317, i_10_328, i_10_329, i_10_332, i_10_440, i_10_443, i_10_465, i_10_749, i_10_796, i_10_797, i_10_901, i_10_991, i_10_1028, i_10_1234, i_10_1244, i_10_1247, i_10_1265, i_10_1307, i_10_1309, i_10_1577, i_10_1579, i_10_1580, i_10_1595, i_10_1648, i_10_1649, i_10_1652, i_10_1690, i_10_1691, i_10_1811, i_10_1819, i_10_1824, i_10_1946, i_10_2018, i_10_2024, i_10_2197, i_10_2201, i_10_2312, i_10_2350, i_10_2351, i_10_2353, i_10_2354, i_10_2406, i_10_2467, i_10_2470, i_10_2503, i_10_2602, i_10_2603, i_10_2606, i_10_2634, i_10_2660, i_10_2710, i_10_2711, i_10_2729, i_10_2731, i_10_2827, i_10_2830, i_10_2831, i_10_2834, i_10_3161, i_10_3196, i_10_3197, i_10_3278, i_10_3583, i_10_3585, i_10_3586, i_10_3613, i_10_3650, i_10_3686, i_10_3781, i_10_3786, i_10_3809, i_10_3835, i_10_3841, i_10_3848, i_10_3889, i_10_3908, i_10_4114, i_10_4115, i_10_4172, i_10_4277, i_10_4285, i_10_4286, i_10_4288, i_10_4289, i_10_4291, i_10_4565, i_10_4570, o_10_46);
	kernel_10_47 k_10_47(i_10_174, i_10_175, i_10_177, i_10_244, i_10_245, i_10_247, i_10_276, i_10_289, i_10_290, i_10_292, i_10_293, i_10_361, i_10_364, i_10_405, i_10_406, i_10_409, i_10_410, i_10_411, i_10_412, i_10_435, i_10_445, i_10_456, i_10_460, i_10_461, i_10_463, i_10_467, i_10_510, i_10_749, i_10_792, i_10_796, i_10_797, i_10_799, i_10_800, i_10_1269, i_10_1306, i_10_1359, i_10_1441, i_10_1442, i_10_1649, i_10_1655, i_10_1819, i_10_1822, i_10_1910, i_10_1992, i_10_2178, i_10_2359, i_10_2360, i_10_2361, i_10_2448, i_10_2467, i_10_2468, i_10_2628, i_10_2630, i_10_2631, i_10_2632, i_10_2658, i_10_2659, i_10_2661, i_10_2673, i_10_2680, i_10_2702, i_10_2731, i_10_2781, i_10_2783, i_10_2784, i_10_2882, i_10_2980, i_10_3044, i_10_3069, i_10_3070, i_10_3071, i_10_3073, i_10_3074, i_10_3277, i_10_3278, i_10_3321, i_10_3323, i_10_3328, i_10_3384, i_10_3392, i_10_3523, i_10_3610, i_10_3613, i_10_3787, i_10_3788, i_10_3807, i_10_3808, i_10_3849, i_10_3855, i_10_3858, i_10_3983, i_10_3994, i_10_4119, i_10_4270, i_10_4285, i_10_4288, i_10_4289, i_10_4291, i_10_4292, i_10_4564, o_10_47);
	kernel_10_48 k_10_48(i_10_174, i_10_180, i_10_248, i_10_287, i_10_327, i_10_369, i_10_448, i_10_586, i_10_588, i_10_633, i_10_781, i_10_782, i_10_795, i_10_798, i_10_799, i_10_904, i_10_1087, i_10_1235, i_10_1241, i_10_1249, i_10_1362, i_10_1363, i_10_1450, i_10_1453, i_10_1454, i_10_1490, i_10_1551, i_10_1555, i_10_1577, i_10_1646, i_10_1789, i_10_1882, i_10_1911, i_10_1914, i_10_1979, i_10_2028, i_10_2082, i_10_2085, i_10_2155, i_10_2158, i_10_2159, i_10_2241, i_10_2261, i_10_2264, i_10_2310, i_10_2322, i_10_2337, i_10_2353, i_10_2383, i_10_2385, i_10_2407, i_10_2411, i_10_2442, i_10_2443, i_10_2449, i_10_2451, i_10_2452, i_10_2517, i_10_2518, i_10_2539, i_10_2572, i_10_2573, i_10_2648, i_10_2703, i_10_2707, i_10_2921, i_10_2924, i_10_2954, i_10_2957, i_10_3101, i_10_3228, i_10_3360, i_10_3390, i_10_3492, i_10_3499, i_10_3525, i_10_3577, i_10_3613, i_10_3618, i_10_3649, i_10_3784, i_10_3837, i_10_3838, i_10_3850, i_10_3856, i_10_3895, i_10_3963, i_10_3964, i_10_3983, i_10_4120, i_10_4188, i_10_4273, i_10_4289, i_10_4423, i_10_4458, i_10_4461, i_10_4513, i_10_4525, i_10_4566, i_10_4569, o_10_48);
	kernel_10_49 k_10_49(i_10_30, i_10_117, i_10_171, i_10_172, i_10_173, i_10_174, i_10_175, i_10_285, i_10_315, i_10_318, i_10_325, i_10_424, i_10_427, i_10_432, i_10_448, i_10_796, i_10_797, i_10_800, i_10_955, i_10_957, i_10_958, i_10_959, i_10_968, i_10_1002, i_10_1028, i_10_1029, i_10_1308, i_10_1311, i_10_1361, i_10_1614, i_10_1617, i_10_1652, i_10_1821, i_10_1944, i_10_1945, i_10_1956, i_10_2016, i_10_2178, i_10_2179, i_10_2181, i_10_2184, i_10_2308, i_10_2354, i_10_2358, i_10_2359, i_10_2361, i_10_2362, i_10_2448, i_10_2457, i_10_2613, i_10_2628, i_10_2629, i_10_2631, i_10_2635, i_10_2700, i_10_2701, i_10_2702, i_10_2718, i_10_2782, i_10_2823, i_10_2826, i_10_2885, i_10_3033, i_10_3034, i_10_3036, i_10_3037, i_10_3041, i_10_3045, i_10_3046, i_10_3087, i_10_3151, i_10_3195, i_10_3196, i_10_3197, i_10_3271, i_10_3278, i_10_3403, i_10_3616, i_10_3645, i_10_3648, i_10_3649, i_10_3650, i_10_3651, i_10_3652, i_10_3780, i_10_3786, i_10_3838, i_10_3852, i_10_3853, i_10_3855, i_10_3856, i_10_3858, i_10_4050, i_10_4122, i_10_4123, i_10_4266, i_10_4288, i_10_4458, i_10_4459, i_10_4571, o_10_49);
	kernel_10_50 k_10_50(i_10_171, i_10_172, i_10_178, i_10_223, i_10_254, i_10_270, i_10_279, i_10_282, i_10_289, i_10_317, i_10_391, i_10_392, i_10_395, i_10_409, i_10_410, i_10_447, i_10_461, i_10_464, i_10_715, i_10_793, i_10_799, i_10_956, i_10_992, i_10_1027, i_10_1028, i_10_1030, i_10_1243, i_10_1244, i_10_1305, i_10_1360, i_10_1433, i_10_1435, i_10_1436, i_10_1489, i_10_1540, i_10_1541, i_10_1543, i_10_1544, i_10_1576, i_10_1577, i_10_1580, i_10_1647, i_10_1655, i_10_1684, i_10_1685, i_10_1688, i_10_1690, i_10_1820, i_10_1822, i_10_1823, i_10_2027, i_10_2030, i_10_2352, i_10_2381, i_10_2470, i_10_2530, i_10_2628, i_10_2630, i_10_2631, i_10_2632, i_10_2633, i_10_2634, i_10_2658, i_10_2659, i_10_2732, i_10_2782, i_10_2834, i_10_2846, i_10_2963, i_10_3035, i_10_3044, i_10_3071, i_10_3073, i_10_3155, i_10_3160, i_10_3199, i_10_3203, i_10_3269, i_10_3332, i_10_3386, i_10_3391, i_10_3473, i_10_3494, i_10_3522, i_10_3583, i_10_3586, i_10_3780, i_10_3781, i_10_3787, i_10_3788, i_10_3838, i_10_3839, i_10_3841, i_10_3848, i_10_3853, i_10_3982, i_10_4172, i_10_4277, i_10_4280, i_10_4287, o_10_50);
	kernel_10_51 k_10_51(i_10_174, i_10_279, i_10_280, i_10_316, i_10_318, i_10_319, i_10_330, i_10_331, i_10_393, i_10_409, i_10_425, i_10_432, i_10_625, i_10_712, i_10_749, i_10_864, i_10_901, i_10_902, i_10_958, i_10_1030, i_10_1036, i_10_1037, i_10_1045, i_10_1046, i_10_1080, i_10_1081, i_10_1084, i_10_1152, i_10_1153, i_10_1299, i_10_1306, i_10_1347, i_10_1378, i_10_1433, i_10_1434, i_10_1435, i_10_1450, i_10_1451, i_10_1541, i_10_1542, i_10_1543, i_10_1545, i_10_1611, i_10_1623, i_10_1626, i_10_1629, i_10_1630, i_10_1631, i_10_1683, i_10_1686, i_10_1714, i_10_1818, i_10_1914, i_10_1915, i_10_1956, i_10_2199, i_10_2200, i_10_2201, i_10_2349, i_10_2350, i_10_2355, i_10_2356, i_10_2471, i_10_2565, i_10_2635, i_10_2677, i_10_2706, i_10_2716, i_10_2719, i_10_2721, i_10_2833, i_10_2866, i_10_2881, i_10_3073, i_10_3223, i_10_3276, i_10_3333, i_10_3384, i_10_3388, i_10_3504, i_10_3609, i_10_3615, i_10_3649, i_10_3807, i_10_3841, i_10_3854, i_10_3859, i_10_3860, i_10_3908, i_10_3925, i_10_3946, i_10_3979, i_10_3980, i_10_4025, i_10_4173, i_10_4275, i_10_4276, i_10_4277, i_10_4278, i_10_4281, o_10_51);
	kernel_10_52 k_10_52(i_10_70, i_10_175, i_10_178, i_10_179, i_10_250, i_10_267, i_10_269, i_10_279, i_10_280, i_10_319, i_10_323, i_10_500, i_10_503, i_10_513, i_10_514, i_10_591, i_10_629, i_10_799, i_10_907, i_10_931, i_10_932, i_10_969, i_10_1011, i_10_1029, i_10_1116, i_10_1223, i_10_1238, i_10_1240, i_10_1241, i_10_1304, i_10_1309, i_10_1311, i_10_1313, i_10_1348, i_10_1349, i_10_1436, i_10_1437, i_10_1438, i_10_1547, i_10_1563, i_10_1628, i_10_1687, i_10_1689, i_10_1705, i_10_1808, i_10_1822, i_10_1885, i_10_1908, i_10_1909, i_10_1960, i_10_2006, i_10_2023, i_10_2030, i_10_2113, i_10_2322, i_10_2345, i_10_2348, i_10_2370, i_10_2436, i_10_2451, i_10_2455, i_10_2456, i_10_2471, i_10_2633, i_10_2641, i_10_2649, i_10_2663, i_10_2714, i_10_2725, i_10_2834, i_10_2851, i_10_2883, i_10_2884, i_10_2887, i_10_2896, i_10_2919, i_10_2923, i_10_3058, i_10_3077, i_10_3266, i_10_3270, i_10_3326, i_10_3338, i_10_3469, i_10_3473, i_10_3590, i_10_3611, i_10_3615, i_10_3787, i_10_3963, i_10_3991, i_10_4000, i_10_4011, i_10_4129, i_10_4156, i_10_4175, i_10_4219, i_10_4273, i_10_4422, i_10_4597, o_10_52);
	kernel_10_53 k_10_53(i_10_48, i_10_135, i_10_146, i_10_175, i_10_187, i_10_216, i_10_218, i_10_444, i_10_544, i_10_792, i_10_793, i_10_796, i_10_820, i_10_981, i_10_1138, i_10_1153, i_10_1233, i_10_1242, i_10_1245, i_10_1306, i_10_1307, i_10_1434, i_10_1443, i_10_1444, i_10_1445, i_10_1485, i_10_1539, i_10_1540, i_10_1542, i_10_1557, i_10_1575, i_10_1582, i_10_1632, i_10_1649, i_10_1651, i_10_1791, i_10_1911, i_10_1912, i_10_1913, i_10_1921, i_10_2088, i_10_2200, i_10_2214, i_10_2349, i_10_2352, i_10_2448, i_10_2449, i_10_2469, i_10_2538, i_10_2604, i_10_2608, i_10_2629, i_10_2630, i_10_2631, i_10_2632, i_10_2635, i_10_2658, i_10_2677, i_10_2700, i_10_2703, i_10_2718, i_10_2721, i_10_2727, i_10_2729, i_10_2737, i_10_2817, i_10_2828, i_10_2829, i_10_2910, i_10_3045, i_10_3199, i_10_3231, i_10_3276, i_10_3280, i_10_3297, i_10_3298, i_10_3388, i_10_3431, i_10_3505, i_10_3609, i_10_3612, i_10_3645, i_10_3702, i_10_3729, i_10_3781, i_10_3783, i_10_3838, i_10_3840, i_10_3847, i_10_3848, i_10_3852, i_10_3854, i_10_3874, i_10_4128, i_10_4219, i_10_4266, i_10_4269, i_10_4276, i_10_4277, i_10_4288, o_10_53);
	kernel_10_54 k_10_54(i_10_184, i_10_185, i_10_188, i_10_210, i_10_211, i_10_213, i_10_220, i_10_251, i_10_405, i_10_432, i_10_441, i_10_466, i_10_498, i_10_516, i_10_577, i_10_578, i_10_586, i_10_594, i_10_694, i_10_699, i_10_800, i_10_928, i_10_960, i_10_969, i_10_987, i_10_1065, i_10_1138, i_10_1167, i_10_1204, i_10_1255, i_10_1256, i_10_1435, i_10_1545, i_10_1605, i_10_1650, i_10_1758, i_10_1759, i_10_1826, i_10_1884, i_10_1911, i_10_1978, i_10_1986, i_10_2158, i_10_2254, i_10_2323, i_10_2349, i_10_2352, i_10_2360, i_10_2403, i_10_2455, i_10_2502, i_10_2506, i_10_2507, i_10_2589, i_10_2598, i_10_2604, i_10_2632, i_10_2640, i_10_2649, i_10_2663, i_10_2676, i_10_2701, i_10_2708, i_10_2716, i_10_2875, i_10_2924, i_10_2983, i_10_3033, i_10_3051, i_10_3052, i_10_3054, i_10_3268, i_10_3270, i_10_3271, i_10_3273, i_10_3299, i_10_3300, i_10_3492, i_10_3493, i_10_3540, i_10_3541, i_10_3683, i_10_3850, i_10_3888, i_10_3963, i_10_4090, i_10_4130, i_10_4188, i_10_4219, i_10_4220, i_10_4230, i_10_4233, i_10_4234, i_10_4279, i_10_4459, i_10_4461, i_10_4513, i_10_4564, i_10_4565, i_10_4571, o_10_54);
	kernel_10_55 k_10_55(i_10_29, i_10_89, i_10_120, i_10_387, i_10_388, i_10_390, i_10_391, i_10_426, i_10_459, i_10_460, i_10_461, i_10_558, i_10_559, i_10_689, i_10_747, i_10_748, i_10_750, i_10_752, i_10_919, i_10_985, i_10_999, i_10_1048, i_10_1053, i_10_1054, i_10_1236, i_10_1237, i_10_1305, i_10_1309, i_10_1362, i_10_1381, i_10_1455, i_10_1578, i_10_1611, i_10_1612, i_10_1613, i_10_1643, i_10_1764, i_10_1765, i_10_1822, i_10_1826, i_10_1945, i_10_1947, i_10_1953, i_10_1954, i_10_1996, i_10_2062, i_10_2108, i_10_2179, i_10_2406, i_10_2413, i_10_2455, i_10_2456, i_10_2478, i_10_2613, i_10_2655, i_10_2659, i_10_2661, i_10_2688, i_10_2689, i_10_2710, i_10_2730, i_10_2817, i_10_2911, i_10_3036, i_10_3037, i_10_3043, i_10_3076, i_10_3090, i_10_3195, i_10_3196, i_10_3348, i_10_3349, i_10_3352, i_10_3469, i_10_3470, i_10_3585, i_10_3618, i_10_3619, i_10_3620, i_10_3637, i_10_3645, i_10_3646, i_10_3647, i_10_3732, i_10_3853, i_10_3854, i_10_3879, i_10_3880, i_10_3942, i_10_3988, i_10_4025, i_10_4028, i_10_4029, i_10_4030, i_10_4051, i_10_4053, i_10_4275, i_10_4341, i_10_4530, i_10_4586, o_10_55);
	kernel_10_56 k_10_56(i_10_27, i_10_33, i_10_34, i_10_52, i_10_172, i_10_178, i_10_224, i_10_258, i_10_282, i_10_366, i_10_390, i_10_408, i_10_409, i_10_442, i_10_445, i_10_498, i_10_502, i_10_541, i_10_602, i_10_798, i_10_954, i_10_958, i_10_960, i_10_990, i_10_991, i_10_992, i_10_1033, i_10_1083, i_10_1088, i_10_1164, i_10_1250, i_10_1305, i_10_1306, i_10_1308, i_10_1309, i_10_1381, i_10_1443, i_10_1545, i_10_1686, i_10_1715, i_10_1770, i_10_1813, i_10_1854, i_10_1908, i_10_2005, i_10_2006, i_10_2254, i_10_2353, i_10_2380, i_10_2460, i_10_2536, i_10_2606, i_10_2632, i_10_2634, i_10_2704, i_10_2714, i_10_2722, i_10_2731, i_10_2742, i_10_2826, i_10_2829, i_10_2884, i_10_2920, i_10_2923, i_10_2986, i_10_3033, i_10_3072, i_10_3076, i_10_3165, i_10_3200, i_10_3201, i_10_3282, i_10_3298, i_10_3330, i_10_3333, i_10_3336, i_10_3405, i_10_3406, i_10_3408, i_10_3441, i_10_3466, i_10_3609, i_10_3612, i_10_3616, i_10_3618, i_10_3624, i_10_3625, i_10_3649, i_10_3652, i_10_3653, i_10_3780, i_10_3783, i_10_3784, i_10_3844, i_10_3847, i_10_3853, i_10_3947, i_10_4126, i_10_4288, i_10_4567, o_10_56);
	kernel_10_57 k_10_57(i_10_52, i_10_178, i_10_224, i_10_275, i_10_277, i_10_281, i_10_283, i_10_287, i_10_408, i_10_446, i_10_730, i_10_797, i_10_898, i_10_958, i_10_996, i_10_997, i_10_1033, i_10_1034, i_10_1247, i_10_1306, i_10_1311, i_10_1363, i_10_1543, i_10_1553, i_10_1579, i_10_1626, i_10_1654, i_10_1689, i_10_1690, i_10_1736, i_10_1819, i_10_1820, i_10_1821, i_10_1822, i_10_1826, i_10_1909, i_10_1912, i_10_1996, i_10_1997, i_10_2019, i_10_2028, i_10_2031, i_10_2352, i_10_2353, i_10_2355, i_10_2449, i_10_2452, i_10_2454, i_10_2455, i_10_2474, i_10_2565, i_10_2568, i_10_2572, i_10_2662, i_10_2705, i_10_2716, i_10_2717, i_10_2721, i_10_2725, i_10_2732, i_10_2734, i_10_2880, i_10_2884, i_10_2917, i_10_2918, i_10_2920, i_10_2964, i_10_3038, i_10_3049, i_10_3054, i_10_3197, i_10_3277, i_10_3384, i_10_3385, i_10_3388, i_10_3391, i_10_3405, i_10_3406, i_10_3501, i_10_3525, i_10_3589, i_10_3610, i_10_3613, i_10_3614, i_10_3617, i_10_3653, i_10_3720, i_10_3780, i_10_3781, i_10_3784, i_10_3834, i_10_3837, i_10_3839, i_10_3857, i_10_3896, i_10_3982, i_10_4030, i_10_4266, i_10_4291, i_10_4567, o_10_57);
	kernel_10_58 k_10_58(i_10_174, i_10_179, i_10_279, i_10_280, i_10_290, i_10_317, i_10_328, i_10_406, i_10_407, i_10_443, i_10_712, i_10_713, i_10_748, i_10_749, i_10_797, i_10_893, i_10_955, i_10_1000, i_10_1001, i_10_1033, i_10_1308, i_10_1309, i_10_1310, i_10_1360, i_10_1540, i_10_1541, i_10_1647, i_10_1649, i_10_1651, i_10_1652, i_10_1683, i_10_1684, i_10_1685, i_10_1687, i_10_1688, i_10_1721, i_10_1729, i_10_1819, i_10_1820, i_10_1826, i_10_1946, i_10_1949, i_10_1989, i_10_1999, i_10_2180, i_10_2198, i_10_2351, i_10_2354, i_10_2358, i_10_2377, i_10_2449, i_10_2450, i_10_2452, i_10_2632, i_10_2674, i_10_2716, i_10_2720, i_10_2723, i_10_2738, i_10_2782, i_10_2785, i_10_2828, i_10_2829, i_10_2917, i_10_2918, i_10_3034, i_10_3035, i_10_3036, i_10_3037, i_10_3038, i_10_3042, i_10_3043, i_10_3087, i_10_3153, i_10_3406, i_10_3407, i_10_3550, i_10_3613, i_10_3614, i_10_3648, i_10_3650, i_10_3834, i_10_3838, i_10_3847, i_10_3848, i_10_3852, i_10_3854, i_10_3856, i_10_3857, i_10_3907, i_10_3910, i_10_3992, i_10_4113, i_10_4122, i_10_4125, i_10_4564, i_10_4565, i_10_4566, i_10_4567, i_10_4568, o_10_58);
	kernel_10_59 k_10_59(i_10_150, i_10_180, i_10_286, i_10_319, i_10_461, i_10_588, i_10_592, i_10_633, i_10_692, i_10_735, i_10_798, i_10_799, i_10_828, i_10_831, i_10_929, i_10_961, i_10_962, i_10_1040, i_10_1041, i_10_1120, i_10_1167, i_10_1180, i_10_1306, i_10_1344, i_10_1346, i_10_1365, i_10_1366, i_10_1554, i_10_1570, i_10_1648, i_10_1744, i_10_1769, i_10_1771, i_10_1785, i_10_1788, i_10_1791, i_10_2011, i_10_2012, i_10_2025, i_10_2142, i_10_2380, i_10_2389, i_10_2437, i_10_2438, i_10_2452, i_10_2478, i_10_2479, i_10_2480, i_10_2542, i_10_2636, i_10_2652, i_10_2713, i_10_2818, i_10_2828, i_10_2831, i_10_2844, i_10_2848, i_10_2883, i_10_2910, i_10_2911, i_10_2922, i_10_2923, i_10_2938, i_10_2958, i_10_2959, i_10_2978, i_10_2986, i_10_3046, i_10_3118, i_10_3211, i_10_3228, i_10_3387, i_10_3390, i_10_3404, i_10_3408, i_10_3468, i_10_3525, i_10_3539, i_10_3585, i_10_3598, i_10_3605, i_10_3772, i_10_3808, i_10_3809, i_10_3894, i_10_3905, i_10_3918, i_10_3964, i_10_3967, i_10_3969, i_10_3991, i_10_3994, i_10_4012, i_10_4013, i_10_4294, i_10_4387, i_10_4440, i_10_4455, i_10_4535, i_10_4598, o_10_59);
	kernel_10_60 k_10_60(i_10_51, i_10_246, i_10_247, i_10_254, i_10_287, i_10_290, i_10_315, i_10_316, i_10_319, i_10_320, i_10_327, i_10_392, i_10_393, i_10_467, i_10_908, i_10_1055, i_10_1083, i_10_1160, i_10_1234, i_10_1235, i_10_1238, i_10_1242, i_10_1245, i_10_1308, i_10_1362, i_10_1432, i_10_1441, i_10_1444, i_10_1540, i_10_1551, i_10_1575, i_10_1576, i_10_1577, i_10_1622, i_10_1655, i_10_1730, i_10_1800, i_10_1911, i_10_1981, i_10_1982, i_10_2196, i_10_2197, i_10_2338, i_10_2349, i_10_2352, i_10_2353, i_10_2354, i_10_2448, i_10_2457, i_10_2515, i_10_2516, i_10_2563, i_10_2567, i_10_2608, i_10_2629, i_10_2701, i_10_2712, i_10_2713, i_10_2731, i_10_2820, i_10_2827, i_10_2845, i_10_2955, i_10_2961, i_10_2962, i_10_3042, i_10_3070, i_10_3071, i_10_3277, i_10_3278, i_10_3353, i_10_3384, i_10_3470, i_10_3538, i_10_3557, i_10_3584, i_10_3610, i_10_3611, i_10_3723, i_10_3835, i_10_3836, i_10_3838, i_10_3857, i_10_3906, i_10_4030, i_10_4062, i_10_4113, i_10_4114, i_10_4122, i_10_4123, i_10_4127, i_10_4151, i_10_4168, i_10_4169, i_10_4191, i_10_4275, i_10_4278, i_10_4289, i_10_4581, i_10_4582, o_10_60);
	kernel_10_61 k_10_61(i_10_122, i_10_148, i_10_277, i_10_289, i_10_326, i_10_370, i_10_412, i_10_413, i_10_463, i_10_505, i_10_640, i_10_733, i_10_959, i_10_1009, i_10_1019, i_10_1054, i_10_1055, i_10_1156, i_10_1202, i_10_1243, i_10_1265, i_10_1287, i_10_1382, i_10_1456, i_10_1499, i_10_1540, i_10_1547, i_10_1611, i_10_1615, i_10_1622, i_10_1625, i_10_1648, i_10_1730, i_10_1747, i_10_1783, i_10_1819, i_10_1936, i_10_2018, i_10_2027, i_10_2156, i_10_2197, i_10_2200, i_10_2332, i_10_2336, i_10_2351, i_10_2359, i_10_2360, i_10_2372, i_10_2432, i_10_2435, i_10_2455, i_10_2513, i_10_2525, i_10_2605, i_10_2606, i_10_2630, i_10_2632, i_10_2824, i_10_2827, i_10_2837, i_10_2847, i_10_2864, i_10_2920, i_10_2975, i_10_2993, i_10_3280, i_10_3281, i_10_3298, i_10_3314, i_10_3317, i_10_3402, i_10_3403, i_10_3440, i_10_3469, i_10_3540, i_10_3565, i_10_3613, i_10_3616, i_10_3721, i_10_3800, i_10_3835, i_10_3836, i_10_3839, i_10_3842, i_10_3858, i_10_3898, i_10_3944, i_10_3982, i_10_3998, i_10_4087, i_10_4088, i_10_4130, i_10_4151, i_10_4156, i_10_4243, i_10_4267, i_10_4276, i_10_4277, i_10_4367, i_10_4595, o_10_61);
	kernel_10_62 k_10_62(i_10_221, i_10_243, i_10_244, i_10_250, i_10_281, i_10_283, i_10_286, i_10_322, i_10_323, i_10_439, i_10_467, i_10_755, i_10_796, i_10_799, i_10_800, i_10_904, i_10_991, i_10_992, i_10_1033, i_10_1034, i_10_1233, i_10_1237, i_10_1238, i_10_1240, i_10_1241, i_10_1300, i_10_1309, i_10_1432, i_10_1437, i_10_1438, i_10_1578, i_10_1579, i_10_1583, i_10_1651, i_10_1653, i_10_1655, i_10_1686, i_10_1816, i_10_1817, i_10_1823, i_10_1912, i_10_1913, i_10_2185, i_10_2306, i_10_2351, i_10_2362, i_10_2363, i_10_2448, i_10_2473, i_10_2608, i_10_2631, i_10_2662, i_10_2705, i_10_2719, i_10_2728, i_10_2734, i_10_2735, i_10_2785, i_10_2786, i_10_2828, i_10_2833, i_10_2834, i_10_2888, i_10_2924, i_10_2986, i_10_3154, i_10_3163, i_10_3196, i_10_3197, i_10_3322, i_10_3388, i_10_3406, i_10_3407, i_10_3588, i_10_3589, i_10_3590, i_10_3613, i_10_3616, i_10_3617, i_10_3646, i_10_3652, i_10_3682, i_10_3838, i_10_3839, i_10_3840, i_10_3841, i_10_3856, i_10_3983, i_10_3984, i_10_3991, i_10_3992, i_10_4028, i_10_4117, i_10_4118, i_10_4120, i_10_4130, i_10_4270, i_10_4271, i_10_4290, i_10_4567, o_10_62);
	kernel_10_63 k_10_63(i_10_174, i_10_216, i_10_220, i_10_246, i_10_292, i_10_293, i_10_328, i_10_329, i_10_410, i_10_443, i_10_445, i_10_465, i_10_645, i_10_897, i_10_898, i_10_899, i_10_1168, i_10_1239, i_10_1240, i_10_1308, i_10_1362, i_10_1366, i_10_1444, i_10_1579, i_10_1648, i_10_1650, i_10_1654, i_10_1675, i_10_1684, i_10_1685, i_10_1825, i_10_1915, i_10_1952, i_10_1995, i_10_1996, i_10_2337, i_10_2350, i_10_2352, i_10_2364, i_10_2365, i_10_2382, i_10_2383, i_10_2408, i_10_2411, i_10_2451, i_10_2470, i_10_2481, i_10_2572, i_10_2631, i_10_2632, i_10_2656, i_10_2658, i_10_2661, i_10_2706, i_10_2707, i_10_2716, i_10_2721, i_10_2731, i_10_2734, i_10_2821, i_10_2824, i_10_2831, i_10_2884, i_10_2919, i_10_2920, i_10_2923, i_10_3034, i_10_3035, i_10_3036, i_10_3153, i_10_3196, i_10_3199, i_10_3202, i_10_3270, i_10_3273, i_10_3279, i_10_3282, i_10_3283, i_10_3388, i_10_3404, i_10_3433, i_10_3469, i_10_3472, i_10_3519, i_10_3522, i_10_3647, i_10_3648, i_10_3651, i_10_3653, i_10_3783, i_10_3785, i_10_3835, i_10_3847, i_10_3848, i_10_3985, i_10_4116, i_10_4119, i_10_4120, i_10_4283, i_10_4291, o_10_63);
	kernel_10_64 k_10_64(i_10_34, i_10_65, i_10_172, i_10_224, i_10_281, i_10_284, i_10_330, i_10_331, i_10_442, i_10_448, i_10_541, i_10_542, i_10_544, i_10_545, i_10_596, i_10_712, i_10_713, i_10_715, i_10_736, i_10_794, i_10_797, i_10_955, i_10_956, i_10_990, i_10_1084, i_10_1241, i_10_1247, i_10_1249, i_10_1309, i_10_1514, i_10_1561, i_10_1562, i_10_1578, i_10_1579, i_10_1580, i_10_1615, i_10_1616, i_10_1650, i_10_1687, i_10_1691, i_10_1765, i_10_1819, i_10_1821, i_10_1824, i_10_1825, i_10_1954, i_10_2156, i_10_2164, i_10_2355, i_10_2361, i_10_2362, i_10_2364, i_10_2365, i_10_2432, i_10_2435, i_10_2470, i_10_2603, i_10_2634, i_10_2662, i_10_2728, i_10_2729, i_10_2817, i_10_2820, i_10_2867, i_10_2979, i_10_2982, i_10_3076, i_10_3077, i_10_3116, i_10_3232, i_10_3233, i_10_3235, i_10_3239, i_10_3316, i_10_3385, i_10_3386, i_10_3407, i_10_3410, i_10_3431, i_10_3590, i_10_3611, i_10_3683, i_10_3728, i_10_3808, i_10_3844, i_10_3845, i_10_3906, i_10_3907, i_10_3994, i_10_4008, i_10_4064, i_10_4100, i_10_4117, i_10_4217, i_10_4220, i_10_4267, i_10_4289, i_10_4292, i_10_4475, i_10_4564, o_10_64);
	kernel_10_65 k_10_65(i_10_29, i_10_49, i_10_50, i_10_171, i_10_224, i_10_263, i_10_277, i_10_316, i_10_317, i_10_319, i_10_320, i_10_322, i_10_326, i_10_346, i_10_362, i_10_388, i_10_433, i_10_434, i_10_437, i_10_440, i_10_441, i_10_442, i_10_448, i_10_715, i_10_716, i_10_800, i_10_947, i_10_991, i_10_992, i_10_1001, i_10_1004, i_10_1046, i_10_1084, i_10_1085, i_10_1135, i_10_1136, i_10_1163, i_10_1217, i_10_1220, i_10_1238, i_10_1239, i_10_1306, i_10_1307, i_10_1342, i_10_1346, i_10_1379, i_10_1432, i_10_1544, i_10_1547, i_10_1613, i_10_1652, i_10_1653, i_10_1823, i_10_2000, i_10_2201, i_10_2203, i_10_2204, i_10_2351, i_10_2354, i_10_2357, i_10_2360, i_10_2362, i_10_2380, i_10_2450, i_10_2630, i_10_2675, i_10_2711, i_10_2713, i_10_2720, i_10_2723, i_10_2724, i_10_2783, i_10_2818, i_10_2819, i_10_2822, i_10_2832, i_10_2882, i_10_2884, i_10_2918, i_10_2921, i_10_2980, i_10_2983, i_10_3092, i_10_3152, i_10_3156, i_10_3202, i_10_3203, i_10_3278, i_10_3281, i_10_3584, i_10_3586, i_10_3615, i_10_3835, i_10_3838, i_10_3841, i_10_3893, i_10_3980, i_10_3983, i_10_4280, i_10_4283, o_10_65);
	kernel_10_66 k_10_66(i_10_28, i_10_29, i_10_117, i_10_118, i_10_121, i_10_180, i_10_181, i_10_262, i_10_266, i_10_348, i_10_390, i_10_435, i_10_441, i_10_442, i_10_444, i_10_460, i_10_461, i_10_559, i_10_560, i_10_562, i_10_599, i_10_795, i_10_999, i_10_1027, i_10_1119, i_10_1165, i_10_1305, i_10_1357, i_10_1359, i_10_1360, i_10_1363, i_10_1366, i_10_1401, i_10_1477, i_10_1612, i_10_1652, i_10_1683, i_10_1691, i_10_1821, i_10_1908, i_10_1920, i_10_1947, i_10_1956, i_10_2309, i_10_2408, i_10_2452, i_10_2455, i_10_2482, i_10_2654, i_10_2656, i_10_2657, i_10_2658, i_10_2659, i_10_2703, i_10_2725, i_10_2744, i_10_2754, i_10_2755, i_10_2826, i_10_2828, i_10_3036, i_10_3203, i_10_3235, i_10_3268, i_10_3271, i_10_3284, i_10_3305, i_10_3349, i_10_3392, i_10_3473, i_10_3480, i_10_3494, i_10_3497, i_10_3561, i_10_3585, i_10_3586, i_10_3587, i_10_3589, i_10_3609, i_10_3610, i_10_3614, i_10_3620, i_10_3625, i_10_3646, i_10_3648, i_10_3649, i_10_3702, i_10_3788, i_10_3838, i_10_3853, i_10_3882, i_10_3883, i_10_3983, i_10_3985, i_10_4054, i_10_4055, i_10_4057, i_10_4118, i_10_4144, i_10_4145, o_10_66);
	kernel_10_67 k_10_67(i_10_144, i_10_146, i_10_219, i_10_223, i_10_387, i_10_388, i_10_423, i_10_424, i_10_425, i_10_426, i_10_427, i_10_445, i_10_460, i_10_462, i_10_463, i_10_507, i_10_508, i_10_693, i_10_711, i_10_747, i_10_795, i_10_796, i_10_900, i_10_995, i_10_1234, i_10_1243, i_10_1246, i_10_1248, i_10_1260, i_10_1305, i_10_1341, i_10_1485, i_10_1683, i_10_1819, i_10_1823, i_10_1825, i_10_1911, i_10_1999, i_10_2019, i_10_2241, i_10_2350, i_10_2351, i_10_2352, i_10_2353, i_10_2354, i_10_2356, i_10_2450, i_10_2451, i_10_2452, i_10_2538, i_10_2543, i_10_2678, i_10_2700, i_10_2701, i_10_2702, i_10_2710, i_10_2716, i_10_2820, i_10_2916, i_10_3037, i_10_3087, i_10_3088, i_10_3091, i_10_3114, i_10_3198, i_10_3237, i_10_3276, i_10_3277, i_10_3280, i_10_3312, i_10_3408, i_10_3409, i_10_3465, i_10_3538, i_10_3582, i_10_3583, i_10_3585, i_10_3586, i_10_3612, i_10_3613, i_10_3648, i_10_3682, i_10_3717, i_10_3780, i_10_3781, i_10_3786, i_10_3807, i_10_3808, i_10_3834, i_10_3835, i_10_3838, i_10_3841, i_10_3850, i_10_3857, i_10_3860, i_10_3985, i_10_4117, i_10_4169, i_10_4284, i_10_4290, o_10_67);
	kernel_10_68 k_10_68(i_10_42, i_10_67, i_10_68, i_10_150, i_10_174, i_10_183, i_10_324, i_10_364, i_10_405, i_10_426, i_10_441, i_10_443, i_10_445, i_10_733, i_10_734, i_10_793, i_10_880, i_10_1119, i_10_1237, i_10_1243, i_10_1308, i_10_1309, i_10_1380, i_10_1609, i_10_1617, i_10_1618, i_10_1648, i_10_1649, i_10_1650, i_10_1689, i_10_1910, i_10_1960, i_10_1995, i_10_1996, i_10_2082, i_10_2355, i_10_2380, i_10_2448, i_10_2449, i_10_2450, i_10_2451, i_10_2452, i_10_2460, i_10_2511, i_10_2589, i_10_2590, i_10_2659, i_10_2701, i_10_2705, i_10_2708, i_10_2715, i_10_2716, i_10_2718, i_10_2730, i_10_2734, i_10_2787, i_10_2788, i_10_2828, i_10_2982, i_10_3048, i_10_3049, i_10_3171, i_10_3199, i_10_3271, i_10_3279, i_10_3289, i_10_3292, i_10_3391, i_10_3392, i_10_3471, i_10_3589, i_10_3609, i_10_3610, i_10_3611, i_10_3648, i_10_3649, i_10_3684, i_10_3720, i_10_3814, i_10_3815, i_10_3834, i_10_3837, i_10_3838, i_10_3855, i_10_3882, i_10_3893, i_10_3945, i_10_3987, i_10_4118, i_10_4182, i_10_4216, i_10_4218, i_10_4233, i_10_4234, i_10_4236, i_10_4237, i_10_4425, i_10_4426, i_10_4506, i_10_4507, o_10_68);
	kernel_10_69 k_10_69(i_10_27, i_10_28, i_10_122, i_10_171, i_10_190, i_10_239, i_10_292, i_10_369, i_10_387, i_10_430, i_10_465, i_10_512, i_10_546, i_10_547, i_10_711, i_10_717, i_10_759, i_10_907, i_10_1040, i_10_1120, i_10_1121, i_10_1179, i_10_1251, i_10_1273, i_10_1310, i_10_1345, i_10_1352, i_10_1380, i_10_1441, i_10_1545, i_10_1548, i_10_1578, i_10_1614, i_10_1616, i_10_1620, i_10_1632, i_10_1654, i_10_1803, i_10_2047, i_10_2160, i_10_2178, i_10_2180, i_10_2209, i_10_2290, i_10_2349, i_10_2352, i_10_2372, i_10_2448, i_10_2449, i_10_2452, i_10_2632, i_10_2686, i_10_2725, i_10_2829, i_10_2830, i_10_2834, i_10_2885, i_10_2922, i_10_2935, i_10_2936, i_10_3034, i_10_3035, i_10_3038, i_10_3046, i_10_3067, i_10_3231, i_10_3274, i_10_3291, i_10_3292, i_10_3293, i_10_3523, i_10_3554, i_10_3611, i_10_3612, i_10_3615, i_10_3621, i_10_3637, i_10_3685, i_10_3699, i_10_3703, i_10_3784, i_10_3786, i_10_3787, i_10_3859, i_10_3961, i_10_3965, i_10_4052, i_10_4091, i_10_4126, i_10_4153, i_10_4231, i_10_4233, i_10_4286, i_10_4304, i_10_4309, i_10_4310, i_10_4503, i_10_4529, i_10_4591, i_10_4592, o_10_69);
	kernel_10_70 k_10_70(i_10_37, i_10_40, i_10_52, i_10_247, i_10_286, i_10_315, i_10_316, i_10_320, i_10_321, i_10_322, i_10_323, i_10_408, i_10_409, i_10_410, i_10_430, i_10_439, i_10_691, i_10_832, i_10_833, i_10_994, i_10_1027, i_10_1030, i_10_1031, i_10_1040, i_10_1048, i_10_1082, i_10_1164, i_10_1165, i_10_1166, i_10_1223, i_10_1233, i_10_1243, i_10_1265, i_10_1267, i_10_1268, i_10_1344, i_10_1345, i_10_1543, i_10_1544, i_10_1575, i_10_1578, i_10_1580, i_10_1650, i_10_1651, i_10_1654, i_10_1713, i_10_1825, i_10_1914, i_10_2017, i_10_2024, i_10_2204, i_10_2242, i_10_2251, i_10_2364, i_10_2459, i_10_2607, i_10_2657, i_10_2661, i_10_2662, i_10_2703, i_10_2704, i_10_2705, i_10_2707, i_10_2724, i_10_2833, i_10_2880, i_10_2982, i_10_2983, i_10_3069, i_10_3237, i_10_3279, i_10_3280, i_10_3288, i_10_3496, i_10_3497, i_10_3523, i_10_3525, i_10_3526, i_10_3615, i_10_3787, i_10_3788, i_10_3852, i_10_3856, i_10_3910, i_10_3913, i_10_3987, i_10_4116, i_10_4117, i_10_4118, i_10_4119, i_10_4125, i_10_4129, i_10_4170, i_10_4173, i_10_4215, i_10_4226, i_10_4272, i_10_4275, i_10_4565, i_10_4568, o_10_70);
	kernel_10_71 k_10_71(i_10_29, i_10_118, i_10_259, i_10_260, i_10_280, i_10_317, i_10_331, i_10_332, i_10_373, i_10_387, i_10_388, i_10_391, i_10_439, i_10_462, i_10_517, i_10_518, i_10_959, i_10_967, i_10_1031, i_10_1043, i_10_1057, i_10_1058, i_10_1083, i_10_1084, i_10_1139, i_10_1233, i_10_1234, i_10_1235, i_10_1237, i_10_1238, i_10_1240, i_10_1291, i_10_1312, i_10_1431, i_10_1433, i_10_1539, i_10_1540, i_10_1576, i_10_1577, i_10_1621, i_10_1654, i_10_1717, i_10_1764, i_10_1768, i_10_1769, i_10_1822, i_10_1824, i_10_1825, i_10_1826, i_10_1958, i_10_1980, i_10_1981, i_10_1984, i_10_2017, i_10_2020, i_10_2351, i_10_2356, i_10_2452, i_10_2471, i_10_2546, i_10_2565, i_10_2566, i_10_2581, i_10_2628, i_10_2631, i_10_2632, i_10_2635, i_10_2659, i_10_2704, i_10_2705, i_10_2713, i_10_2734, i_10_2824, i_10_2830, i_10_2921, i_10_3035, i_10_3039, i_10_3050, i_10_3073, i_10_3196, i_10_3323, i_10_3586, i_10_3612, i_10_3619, i_10_3620, i_10_3720, i_10_3786, i_10_3910, i_10_3947, i_10_3983, i_10_4004, i_10_4051, i_10_4054, i_10_4123, i_10_4168, i_10_4169, i_10_4171, i_10_4192, i_10_4282, i_10_4530, o_10_71);
	kernel_10_72 k_10_72(i_10_174, i_10_183, i_10_408, i_10_424, i_10_447, i_10_515, i_10_517, i_10_637, i_10_798, i_10_903, i_10_962, i_10_967, i_10_968, i_10_996, i_10_1032, i_10_1087, i_10_1236, i_10_1237, i_10_1238, i_10_1246, i_10_1247, i_10_1249, i_10_1250, i_10_1491, i_10_1544, i_10_1619, i_10_1647, i_10_1689, i_10_1821, i_10_1823, i_10_1825, i_10_1912, i_10_1945, i_10_2008, i_10_2311, i_10_2382, i_10_2383, i_10_2450, i_10_2452, i_10_2453, i_10_2470, i_10_2471, i_10_2643, i_10_2644, i_10_2681, i_10_2715, i_10_2716, i_10_2721, i_10_2722, i_10_2730, i_10_2732, i_10_2733, i_10_2785, i_10_2827, i_10_2833, i_10_2834, i_10_2880, i_10_2917, i_10_2920, i_10_2921, i_10_3035, i_10_3043, i_10_3044, i_10_3069, i_10_3072, i_10_3164, i_10_3199, i_10_3282, i_10_3387, i_10_3390, i_10_3391, i_10_3406, i_10_3468, i_10_3495, i_10_3496, i_10_3506, i_10_3526, i_10_3583, i_10_3586, i_10_3587, i_10_3589, i_10_3613, i_10_3616, i_10_3617, i_10_3648, i_10_3652, i_10_3653, i_10_3783, i_10_3784, i_10_3785, i_10_3786, i_10_3854, i_10_3878, i_10_4115, i_10_4126, i_10_4213, i_10_4218, i_10_4272, i_10_4273, i_10_4568, o_10_72);
	kernel_10_73 k_10_73(i_10_270, i_10_273, i_10_282, i_10_283, i_10_284, i_10_289, i_10_290, i_10_293, i_10_315, i_10_391, i_10_408, i_10_411, i_10_424, i_10_425, i_10_441, i_10_442, i_10_794, i_10_1163, i_10_1310, i_10_1360, i_10_1361, i_10_1444, i_10_1445, i_10_1540, i_10_1543, i_10_1575, i_10_1577, i_10_1579, i_10_1649, i_10_1650, i_10_1651, i_10_1688, i_10_1721, i_10_1818, i_10_1819, i_10_1821, i_10_1946, i_10_1991, i_10_1993, i_10_2183, i_10_2197, i_10_2350, i_10_2353, i_10_2358, i_10_2359, i_10_2458, i_10_2471, i_10_2629, i_10_2630, i_10_2632, i_10_2634, i_10_2656, i_10_2657, i_10_2659, i_10_2660, i_10_2674, i_10_2675, i_10_2700, i_10_2703, i_10_2710, i_10_2711, i_10_2719, i_10_2721, i_10_2722, i_10_2724, i_10_2828, i_10_2829, i_10_2830, i_10_2885, i_10_2983, i_10_3043, i_10_3088, i_10_3089, i_10_3201, i_10_3232, i_10_3233, i_10_3328, i_10_3349, i_10_3350, i_10_3390, i_10_3431, i_10_3523, i_10_3527, i_10_3549, i_10_3586, i_10_3587, i_10_3609, i_10_3610, i_10_3835, i_10_3845, i_10_3859, i_10_3944, i_10_3983, i_10_4052, i_10_4168, i_10_4169, i_10_4275, i_10_4284, i_10_4567, i_10_4568, o_10_73);
	kernel_10_74 k_10_74(i_10_26, i_10_208, i_10_248, i_10_257, i_10_272, i_10_275, i_10_391, i_10_394, i_10_408, i_10_443, i_10_445, i_10_520, i_10_716, i_10_729, i_10_797, i_10_799, i_10_955, i_10_970, i_10_971, i_10_1037, i_10_1235, i_10_1243, i_10_1244, i_10_1246, i_10_1247, i_10_1310, i_10_1541, i_10_1544, i_10_1550, i_10_1552, i_10_1655, i_10_1688, i_10_1759, i_10_1909, i_10_1910, i_10_1911, i_10_1957, i_10_2008, i_10_2027, i_10_2155, i_10_2180, i_10_2242, i_10_2334, i_10_2336, i_10_2339, i_10_2379, i_10_2405, i_10_2411, i_10_2441, i_10_2442, i_10_2456, i_10_2506, i_10_2531, i_10_2534, i_10_2629, i_10_2637, i_10_2638, i_10_2640, i_10_2647, i_10_2702, i_10_2723, i_10_2729, i_10_2866, i_10_2920, i_10_2954, i_10_3033, i_10_3034, i_10_3036, i_10_3074, i_10_3197, i_10_3205, i_10_3224, i_10_3226, i_10_3286, i_10_3331, i_10_3332, i_10_3585, i_10_3650, i_10_3787, i_10_3817, i_10_3851, i_10_3860, i_10_3944, i_10_3965, i_10_4113, i_10_4117, i_10_4118, i_10_4185, i_10_4186, i_10_4188, i_10_4267, i_10_4268, i_10_4270, i_10_4271, i_10_4286, i_10_4289, i_10_4514, i_10_4528, i_10_4564, i_10_4566, o_10_74);
	kernel_10_75 k_10_75(i_10_38, i_10_49, i_10_66, i_10_69, i_10_155, i_10_191, i_10_194, i_10_218, i_10_237, i_10_246, i_10_425, i_10_442, i_10_460, i_10_595, i_10_621, i_10_794, i_10_958, i_10_995, i_10_1026, i_10_1245, i_10_1246, i_10_1299, i_10_1310, i_10_1314, i_10_1445, i_10_1485, i_10_1549, i_10_1550, i_10_1559, i_10_1798, i_10_1823, i_10_1854, i_10_1876, i_10_2036, i_10_2198, i_10_2324, i_10_2350, i_10_2351, i_10_2353, i_10_2448, i_10_2449, i_10_2450, i_10_2453, i_10_2474, i_10_2475, i_10_2530, i_10_2531, i_10_2532, i_10_2569, i_10_2603, i_10_2674, i_10_2707, i_10_2710, i_10_2713, i_10_2727, i_10_2804, i_10_2818, i_10_2888, i_10_2909, i_10_2980, i_10_2983, i_10_2984, i_10_2989, i_10_2992, i_10_3076, i_10_3077, i_10_3198, i_10_3206, i_10_3277, i_10_3278, i_10_3303, i_10_3333, i_10_3462, i_10_3468, i_10_3469, i_10_3470, i_10_3501, i_10_3503, i_10_3522, i_10_3523, i_10_3524, i_10_3541, i_10_3613, i_10_3649, i_10_3774, i_10_3783, i_10_3853, i_10_3854, i_10_3857, i_10_3859, i_10_3860, i_10_3911, i_10_3926, i_10_4005, i_10_4214, i_10_4249, i_10_4277, i_10_4291, i_10_4457, i_10_4559, o_10_75);
	kernel_10_76 k_10_76(i_10_40, i_10_174, i_10_175, i_10_178, i_10_244, i_10_284, i_10_285, i_10_316, i_10_317, i_10_395, i_10_405, i_10_406, i_10_410, i_10_438, i_10_447, i_10_448, i_10_449, i_10_463, i_10_464, i_10_533, i_10_626, i_10_718, i_10_719, i_10_752, i_10_755, i_10_958, i_10_959, i_10_969, i_10_990, i_10_991, i_10_994, i_10_1051, i_10_1123, i_10_1233, i_10_1238, i_10_1344, i_10_1433, i_10_1445, i_10_1539, i_10_1546, i_10_1621, i_10_1622, i_10_1626, i_10_1635, i_10_1652, i_10_1685, i_10_1766, i_10_1825, i_10_2003, i_10_2019, i_10_2164, i_10_2355, i_10_2356, i_10_2359, i_10_2362, i_10_2514, i_10_2539, i_10_2562, i_10_2563, i_10_2570, i_10_2604, i_10_2632, i_10_2676, i_10_2706, i_10_2733, i_10_2734, i_10_2781, i_10_2866, i_10_2884, i_10_3046, i_10_3069, i_10_3070, i_10_3072, i_10_3073, i_10_3074, i_10_3279, i_10_3283, i_10_3284, i_10_3387, i_10_3540, i_10_3583, i_10_3648, i_10_3651, i_10_3811, i_10_3812, i_10_3840, i_10_3987, i_10_3988, i_10_4114, i_10_4115, i_10_4121, i_10_4129, i_10_4150, i_10_4151, i_10_4172, i_10_4174, i_10_4216, i_10_4276, i_10_4279, i_10_4571, o_10_76);
	kernel_10_77 k_10_77(i_10_71, i_10_83, i_10_217, i_10_254, i_10_277, i_10_320, i_10_322, i_10_388, i_10_409, i_10_423, i_10_424, i_10_425, i_10_427, i_10_428, i_10_434, i_10_532, i_10_693, i_10_904, i_10_991, i_10_1028, i_10_1033, i_10_1040, i_10_1043, i_10_1117, i_10_1171, i_10_1197, i_10_1308, i_10_1399, i_10_1400, i_10_1577, i_10_1733, i_10_1741, i_10_1766, i_10_1768, i_10_1822, i_10_1910, i_10_1944, i_10_1948, i_10_1985, i_10_1991, i_10_1993, i_10_2023, i_10_2377, i_10_2383, i_10_2454, i_10_2455, i_10_2458, i_10_2476, i_10_2557, i_10_2558, i_10_2560, i_10_2569, i_10_2635, i_10_2647, i_10_2648, i_10_2650, i_10_2658, i_10_2659, i_10_2711, i_10_2714, i_10_2720, i_10_2721, i_10_2722, i_10_2881, i_10_2885, i_10_2923, i_10_3071, i_10_3088, i_10_3092, i_10_3195, i_10_3203, i_10_3278, i_10_3353, i_10_3385, i_10_3386, i_10_3387, i_10_3389, i_10_3405, i_10_3440, i_10_3547, i_10_3548, i_10_3550, i_10_3610, i_10_3611, i_10_3834, i_10_3841, i_10_3855, i_10_3856, i_10_3979, i_10_3989, i_10_4024, i_10_4025, i_10_4027, i_10_4029, i_10_4030, i_10_4128, i_10_4171, i_10_4456, i_10_4578, i_10_4590, o_10_77);
	kernel_10_78 k_10_78(i_10_15, i_10_117, i_10_118, i_10_121, i_10_140, i_10_265, i_10_282, i_10_328, i_10_449, i_10_513, i_10_562, i_10_634, i_10_718, i_10_930, i_10_958, i_10_959, i_10_963, i_10_1033, i_10_1162, i_10_1163, i_10_1206, i_10_1239, i_10_1362, i_10_1380, i_10_1451, i_10_1533, i_10_1634, i_10_1642, i_10_1654, i_10_1686, i_10_1687, i_10_1688, i_10_1722, i_10_1723, i_10_1724, i_10_1729, i_10_1730, i_10_1795, i_10_1821, i_10_1914, i_10_1948, i_10_2057, i_10_2065, i_10_2066, i_10_2241, i_10_2244, i_10_2349, i_10_2350, i_10_2365, i_10_2390, i_10_2468, i_10_2469, i_10_2517, i_10_2541, i_10_2542, i_10_2544, i_10_2607, i_10_2608, i_10_2614, i_10_2615, i_10_2666, i_10_2715, i_10_2721, i_10_2722, i_10_2741, i_10_2995, i_10_3035, i_10_3036, i_10_3070, i_10_3390, i_10_3391, i_10_3392, i_10_3449, i_10_3451, i_10_3492, i_10_3493, i_10_3496, i_10_3525, i_10_3541, i_10_3544, i_10_3613, i_10_3648, i_10_3652, i_10_3719, i_10_3777, i_10_3853, i_10_3854, i_10_3878, i_10_3913, i_10_3983, i_10_4114, i_10_4115, i_10_4116, i_10_4129, i_10_4131, i_10_4290, i_10_4450, i_10_4458, i_10_4459, i_10_4531, o_10_78);
	kernel_10_79 k_10_79(i_10_175, i_10_187, i_10_246, i_10_249, i_10_265, i_10_283, i_10_411, i_10_412, i_10_430, i_10_431, i_10_440, i_10_444, i_10_446, i_10_457, i_10_509, i_10_518, i_10_521, i_10_797, i_10_956, i_10_957, i_10_958, i_10_959, i_10_967, i_10_997, i_10_1006, i_10_1007, i_10_1052, i_10_1138, i_10_1140, i_10_1247, i_10_1248, i_10_1493, i_10_1555, i_10_1556, i_10_1653, i_10_1691, i_10_1823, i_10_1913, i_10_1987, i_10_2005, i_10_2006, i_10_2350, i_10_2353, i_10_2364, i_10_2452, i_10_2474, i_10_2509, i_10_2607, i_10_2656, i_10_2662, i_10_2681, i_10_2706, i_10_2716, i_10_2717, i_10_2721, i_10_2732, i_10_2734, i_10_2735, i_10_2852, i_10_2880, i_10_2884, i_10_2885, i_10_2887, i_10_2922, i_10_3039, i_10_3093, i_10_3094, i_10_3095, i_10_3281, i_10_3355, i_10_3387, i_10_3388, i_10_3389, i_10_3406, i_10_3409, i_10_3472, i_10_3473, i_10_3497, i_10_3585, i_10_3587, i_10_3613, i_10_3646, i_10_3648, i_10_3649, i_10_3651, i_10_3784, i_10_3785, i_10_3786, i_10_3787, i_10_3788, i_10_3836, i_10_3847, i_10_3850, i_10_3851, i_10_3913, i_10_3914, i_10_3983, i_10_3986, i_10_4116, i_10_4117, o_10_79);
	kernel_10_80 k_10_80(i_10_52, i_10_224, i_10_293, i_10_319, i_10_425, i_10_427, i_10_464, i_10_694, i_10_793, i_10_845, i_10_849, i_10_927, i_10_1000, i_10_1037, i_10_1045, i_10_1118, i_10_1299, i_10_1341, i_10_1342, i_10_1343, i_10_1352, i_10_1438, i_10_1450, i_10_1549, i_10_1550, i_10_1553, i_10_1616, i_10_1652, i_10_1715, i_10_1728, i_10_1742, i_10_1766, i_10_1822, i_10_1873, i_10_1909, i_10_1910, i_10_1913, i_10_1946, i_10_2091, i_10_2183, i_10_2185, i_10_2186, i_10_2209, i_10_2305, i_10_2309, i_10_2312, i_10_2448, i_10_2450, i_10_2453, i_10_2464, i_10_2479, i_10_2480, i_10_2566, i_10_2640, i_10_2648, i_10_2663, i_10_2674, i_10_2677, i_10_2725, i_10_2740, i_10_2741, i_10_2831, i_10_2880, i_10_2881, i_10_2882, i_10_2918, i_10_2920, i_10_3052, i_10_3091, i_10_3201, i_10_3203, i_10_3268, i_10_3276, i_10_3277, i_10_3278, i_10_3350, i_10_3406, i_10_3410, i_10_3431, i_10_3602, i_10_3604, i_10_3704, i_10_3796, i_10_3828, i_10_3889, i_10_3901, i_10_3902, i_10_3979, i_10_3980, i_10_3983, i_10_4029, i_10_4099, i_10_4115, i_10_4124, i_10_4127, i_10_4175, i_10_4270, i_10_4564, i_10_4591, i_10_4594, o_10_80);
	kernel_10_81 k_10_81(i_10_76, i_10_124, i_10_179, i_10_183, i_10_184, i_10_247, i_10_260, i_10_281, i_10_317, i_10_318, i_10_319, i_10_320, i_10_322, i_10_323, i_10_376, i_10_394, i_10_410, i_10_430, i_10_435, i_10_436, i_10_467, i_10_629, i_10_692, i_10_1032, i_10_1045, i_10_1083, i_10_1138, i_10_1158, i_10_1160, i_10_1166, i_10_1169, i_10_1240, i_10_1241, i_10_1268, i_10_1305, i_10_1312, i_10_1341, i_10_1366, i_10_1385, i_10_1542, i_10_1547, i_10_1713, i_10_1821, i_10_1851, i_10_1852, i_10_1879, i_10_1880, i_10_1912, i_10_1913, i_10_2059, i_10_2202, i_10_2203, i_10_2204, i_10_2355, i_10_2356, i_10_2380, i_10_2456, i_10_2542, i_10_2543, i_10_2580, i_10_2581, i_10_2582, i_10_2605, i_10_2608, i_10_2609, i_10_2636, i_10_2681, i_10_2705, i_10_2717, i_10_2725, i_10_2786, i_10_2834, i_10_2842, i_10_2884, i_10_2919, i_10_2986, i_10_2987, i_10_3072, i_10_3073, i_10_3198, i_10_3237, i_10_3283, i_10_3302, i_10_3391, i_10_3472, i_10_3589, i_10_3610, i_10_3911, i_10_3944, i_10_3948, i_10_3979, i_10_4028, i_10_4116, i_10_4117, i_10_4121, i_10_4126, i_10_4174, i_10_4281, i_10_4282, i_10_4288, o_10_81);
	kernel_10_82 k_10_82(i_10_244, i_10_247, i_10_265, i_10_279, i_10_316, i_10_320, i_10_406, i_10_460, i_10_467, i_10_755, i_10_820, i_10_960, i_10_997, i_10_1084, i_10_1236, i_10_1313, i_10_1345, i_10_1346, i_10_1348, i_10_1360, i_10_1543, i_10_1552, i_10_1580, i_10_1583, i_10_1630, i_10_1648, i_10_1649, i_10_1654, i_10_1655, i_10_1683, i_10_1713, i_10_1768, i_10_1800, i_10_1824, i_10_1825, i_10_1912, i_10_1988, i_10_2025, i_10_2182, i_10_2197, i_10_2198, i_10_2312, i_10_2361, i_10_2384, i_10_2457, i_10_2458, i_10_2468, i_10_2470, i_10_2565, i_10_2659, i_10_2660, i_10_2673, i_10_2701, i_10_2709, i_10_2710, i_10_2719, i_10_2720, i_10_2723, i_10_2729, i_10_2730, i_10_2735, i_10_2757, i_10_2882, i_10_2884, i_10_2887, i_10_2920, i_10_3046, i_10_3049, i_10_3268, i_10_3279, i_10_3280, i_10_3312, i_10_3325, i_10_3406, i_10_3407, i_10_3410, i_10_3541, i_10_3545, i_10_3585, i_10_3586, i_10_3610, i_10_3614, i_10_3650, i_10_3784, i_10_3808, i_10_3838, i_10_3847, i_10_3848, i_10_3854, i_10_3857, i_10_3994, i_10_4113, i_10_4116, i_10_4117, i_10_4118, i_10_4273, i_10_4285, i_10_4291, i_10_4568, i_10_4590, o_10_82);
	kernel_10_83 k_10_83(i_10_82, i_10_117, i_10_118, i_10_120, i_10_172, i_10_173, i_10_174, i_10_175, i_10_247, i_10_280, i_10_281, i_10_315, i_10_322, i_10_444, i_10_447, i_10_499, i_10_515, i_10_564, i_10_740, i_10_758, i_10_932, i_10_1238, i_10_1245, i_10_1306, i_10_1308, i_10_1311, i_10_1312, i_10_1361, i_10_1542, i_10_1611, i_10_1620, i_10_1648, i_10_1683, i_10_1821, i_10_1822, i_10_1918, i_10_1944, i_10_1945, i_10_1946, i_10_1947, i_10_1948, i_10_1951, i_10_1956, i_10_2023, i_10_2179, i_10_2243, i_10_2356, i_10_2380, i_10_2432, i_10_2460, i_10_2466, i_10_2511, i_10_2631, i_10_2635, i_10_2655, i_10_2656, i_10_2673, i_10_2674, i_10_2703, i_10_2711, i_10_2713, i_10_2716, i_10_2722, i_10_2727, i_10_2729, i_10_2819, i_10_2831, i_10_2885, i_10_2987, i_10_3036, i_10_3046, i_10_3089, i_10_3268, i_10_3278, i_10_3281, i_10_3284, i_10_3286, i_10_3296, i_10_3523, i_10_3524, i_10_3561, i_10_3614, i_10_3618, i_10_3649, i_10_3838, i_10_3854, i_10_3860, i_10_4023, i_10_4050, i_10_4117, i_10_4129, i_10_4174, i_10_4283, i_10_4286, i_10_4352, i_10_4460, i_10_4558, i_10_4559, i_10_4568, i_10_4569, o_10_83);
	kernel_10_84 k_10_84(i_10_221, i_10_240, i_10_283, i_10_296, i_10_413, i_10_438, i_10_445, i_10_446, i_10_465, i_10_466, i_10_799, i_10_827, i_10_897, i_10_993, i_10_996, i_10_1033, i_10_1034, i_10_1085, i_10_1153, i_10_1174, i_10_1175, i_10_1205, i_10_1233, i_10_1234, i_10_1238, i_10_1246, i_10_1247, i_10_1248, i_10_1308, i_10_1349, i_10_1363, i_10_1555, i_10_1556, i_10_1610, i_10_1627, i_10_1648, i_10_1687, i_10_1818, i_10_1819, i_10_1825, i_10_1950, i_10_2002, i_10_2003, i_10_2350, i_10_2351, i_10_2357, i_10_2364, i_10_2384, i_10_2411, i_10_2449, i_10_2465, i_10_2519, i_10_2540, i_10_2542, i_10_2543, i_10_2545, i_10_2572, i_10_2573, i_10_2634, i_10_2635, i_10_2708, i_10_2712, i_10_2730, i_10_2818, i_10_2830, i_10_2880, i_10_2887, i_10_2917, i_10_2918, i_10_2921, i_10_2922, i_10_2956, i_10_3039, i_10_3049, i_10_3090, i_10_3091, i_10_3162, i_10_3163, i_10_3277, i_10_3356, i_10_3390, i_10_3392, i_10_3446, i_10_3586, i_10_3613, i_10_3688, i_10_3689, i_10_3717, i_10_3734, i_10_3786, i_10_3850, i_10_3859, i_10_3892, i_10_4168, i_10_4267, i_10_4276, i_10_4277, i_10_4279, i_10_4568, i_10_4571, o_10_84);
	kernel_10_85 k_10_85(i_10_64, i_10_253, i_10_254, i_10_316, i_10_328, i_10_388, i_10_390, i_10_391, i_10_435, i_10_442, i_10_443, i_10_444, i_10_466, i_10_467, i_10_504, i_10_512, i_10_793, i_10_796, i_10_800, i_10_1002, i_10_1027, i_10_1028, i_10_1033, i_10_1034, i_10_1343, i_10_1433, i_10_1436, i_10_1442, i_10_1445, i_10_1539, i_10_1540, i_10_1541, i_10_1576, i_10_1579, i_10_1580, i_10_1620, i_10_1650, i_10_1688, i_10_1689, i_10_1690, i_10_1818, i_10_1819, i_10_1823, i_10_1910, i_10_1984, i_10_1988, i_10_1995, i_10_2198, i_10_2305, i_10_2306, i_10_2349, i_10_2363, i_10_2380, i_10_2530, i_10_2531, i_10_2603, i_10_2655, i_10_2677, i_10_2712, i_10_2721, i_10_2723, i_10_2735, i_10_2829, i_10_2830, i_10_2862, i_10_2863, i_10_2885, i_10_2924, i_10_3036, i_10_3088, i_10_3199, i_10_3201, i_10_3202, i_10_3270, i_10_3277, i_10_3278, i_10_3298, i_10_3321, i_10_3325, i_10_3386, i_10_3392, i_10_3406, i_10_3407, i_10_3614, i_10_3781, i_10_3782, i_10_3783, i_10_3784, i_10_3837, i_10_3853, i_10_3943, i_10_3979, i_10_3980, i_10_4006, i_10_4116, i_10_4286, i_10_4287, i_10_4565, i_10_4591, i_10_4592, o_10_85);
	kernel_10_86 k_10_86(i_10_174, i_10_220, i_10_221, i_10_245, i_10_287, i_10_328, i_10_408, i_10_409, i_10_410, i_10_441, i_10_442, i_10_508, i_10_509, i_10_797, i_10_892, i_10_958, i_10_994, i_10_1026, i_10_1027, i_10_1028, i_10_1242, i_10_1262, i_10_1305, i_10_1432, i_10_1541, i_10_1620, i_10_1621, i_10_1685, i_10_1691, i_10_1819, i_10_1820, i_10_1821, i_10_1909, i_10_1990, i_10_2161, i_10_2353, i_10_2356, i_10_2359, i_10_2362, i_10_2448, i_10_2450, i_10_2566, i_10_2628, i_10_2629, i_10_2630, i_10_2631, i_10_2632, i_10_2633, i_10_2635, i_10_2719, i_10_2722, i_10_2729, i_10_2781, i_10_2785, i_10_2817, i_10_2818, i_10_2826, i_10_2827, i_10_2828, i_10_2834, i_10_2880, i_10_2881, i_10_2882, i_10_2884, i_10_2921, i_10_2923, i_10_2924, i_10_3069, i_10_3070, i_10_3088, i_10_3199, i_10_3272, i_10_3384, i_10_3407, i_10_3523, i_10_3555, i_10_3583, i_10_3584, i_10_3585, i_10_3610, i_10_3612, i_10_3780, i_10_3783, i_10_3785, i_10_3838, i_10_3839, i_10_3844, i_10_3846, i_10_3852, i_10_3889, i_10_4114, i_10_4116, i_10_4122, i_10_4123, i_10_4126, i_10_4168, i_10_4214, i_10_4566, i_10_4590, i_10_4591, o_10_86);
	kernel_10_87 k_10_87(i_10_182, i_10_220, i_10_247, i_10_285, i_10_290, i_10_328, i_10_329, i_10_371, i_10_407, i_10_623, i_10_729, i_10_730, i_10_731, i_10_733, i_10_754, i_10_796, i_10_797, i_10_899, i_10_1030, i_10_1031, i_10_1219, i_10_1264, i_10_1267, i_10_1306, i_10_1307, i_10_1308, i_10_1312, i_10_1345, i_10_1349, i_10_1441, i_10_1442, i_10_1913, i_10_1987, i_10_2017, i_10_2019, i_10_2020, i_10_2197, i_10_2201, i_10_2324, i_10_2358, i_10_2386, i_10_2461, i_10_2463, i_10_2464, i_10_2467, i_10_2471, i_10_2628, i_10_2631, i_10_2632, i_10_2656, i_10_2704, i_10_2722, i_10_2785, i_10_2804, i_10_2827, i_10_2870, i_10_2916, i_10_2917, i_10_2918, i_10_2919, i_10_2920, i_10_2922, i_10_2984, i_10_3035, i_10_3070, i_10_3196, i_10_3203, i_10_3390, i_10_3402, i_10_3430, i_10_3519, i_10_3522, i_10_3588, i_10_3609, i_10_3611, i_10_3614, i_10_3645, i_10_3647, i_10_3648, i_10_3649, i_10_3734, i_10_3783, i_10_3787, i_10_3788, i_10_3842, i_10_3853, i_10_3855, i_10_4028, i_10_4113, i_10_4167, i_10_4170, i_10_4171, i_10_4172, i_10_4212, i_10_4215, i_10_4216, i_10_4217, i_10_4288, i_10_4289, i_10_4462, o_10_87);
	kernel_10_88 k_10_88(i_10_86, i_10_174, i_10_177, i_10_179, i_10_264, i_10_284, i_10_409, i_10_413, i_10_536, i_10_635, i_10_754, i_10_797, i_10_961, i_10_964, i_10_994, i_10_996, i_10_1028, i_10_1160, i_10_1238, i_10_1241, i_10_1274, i_10_1310, i_10_1345, i_10_1346, i_10_1360, i_10_1361, i_10_1364, i_10_1436, i_10_1438, i_10_1439, i_10_1542, i_10_1547, i_10_1549, i_10_1555, i_10_1582, i_10_1625, i_10_1627, i_10_1628, i_10_1650, i_10_1736, i_10_1821, i_10_1823, i_10_1994, i_10_2023, i_10_2024, i_10_2032, i_10_2033, i_10_2201, i_10_2324, i_10_2350, i_10_2364, i_10_2453, i_10_2456, i_10_2507, i_10_2516, i_10_2609, i_10_2628, i_10_2632, i_10_2656, i_10_2674, i_10_2678, i_10_2711, i_10_2717, i_10_2732, i_10_2734, i_10_2783, i_10_2789, i_10_2829, i_10_2831, i_10_2850, i_10_2884, i_10_2885, i_10_2967, i_10_2968, i_10_2969, i_10_3047, i_10_3074, i_10_3077, i_10_3091, i_10_3199, i_10_3277, i_10_3290, i_10_3337, i_10_3431, i_10_3434, i_10_3470, i_10_3494, i_10_3507, i_10_3584, i_10_3652, i_10_3841, i_10_3850, i_10_3860, i_10_4051, i_10_4130, i_10_4175, i_10_4262, i_10_4292, i_10_4460, i_10_4586, o_10_88);
	kernel_10_89 k_10_89(i_10_68, i_10_263, i_10_270, i_10_273, i_10_274, i_10_282, i_10_283, i_10_284, i_10_287, i_10_315, i_10_317, i_10_318, i_10_319, i_10_320, i_10_322, i_10_323, i_10_391, i_10_392, i_10_410, i_10_442, i_10_443, i_10_559, i_10_560, i_10_991, i_10_1001, i_10_1004, i_10_1085, i_10_1111, i_10_1138, i_10_1235, i_10_1238, i_10_1307, i_10_1309, i_10_1310, i_10_1311, i_10_1360, i_10_1379, i_10_1433, i_10_1436, i_10_1442, i_10_1544, i_10_1546, i_10_1547, i_10_1580, i_10_1651, i_10_1652, i_10_1730, i_10_1825, i_10_1826, i_10_2000, i_10_2024, i_10_2312, i_10_2352, i_10_2354, i_10_2356, i_10_2449, i_10_2468, i_10_2538, i_10_2558, i_10_2567, i_10_2605, i_10_2615, i_10_2632, i_10_2703, i_10_2704, i_10_2707, i_10_2713, i_10_2719, i_10_2723, i_10_2727, i_10_2728, i_10_2731, i_10_2833, i_10_2834, i_10_3044, i_10_3072, i_10_3268, i_10_3467, i_10_3542, i_10_3545, i_10_3584, i_10_3647, i_10_3650, i_10_3653, i_10_3775, i_10_3785, i_10_3839, i_10_3840, i_10_3859, i_10_3980, i_10_3983, i_10_3986, i_10_4114, i_10_4115, i_10_4116, i_10_4117, i_10_4121, i_10_4283, i_10_4285, i_10_4288, o_10_89);
	kernel_10_90 k_10_90(i_10_31, i_10_32, i_10_175, i_10_190, i_10_221, i_10_330, i_10_331, i_10_387, i_10_390, i_10_391, i_10_432, i_10_463, i_10_946, i_10_990, i_10_1037, i_10_1056, i_10_1081, i_10_1116, i_10_1233, i_10_1242, i_10_1243, i_10_1366, i_10_1432, i_10_1652, i_10_1654, i_10_1655, i_10_1730, i_10_1913, i_10_1921, i_10_1945, i_10_1949, i_10_1954, i_10_1992, i_10_2182, i_10_2304, i_10_2349, i_10_2350, i_10_2381, i_10_2449, i_10_2450, i_10_2466, i_10_2467, i_10_2469, i_10_2529, i_10_2602, i_10_2606, i_10_2629, i_10_2636, i_10_2701, i_10_2705, i_10_2721, i_10_2722, i_10_2725, i_10_2953, i_10_2979, i_10_3034, i_10_3035, i_10_3044, i_10_3074, i_10_3095, i_10_3231, i_10_3233, i_10_3277, i_10_3281, i_10_3312, i_10_3385, i_10_3402, i_10_3434, i_10_3466, i_10_3586, i_10_3587, i_10_3590, i_10_3610, i_10_3614, i_10_3646, i_10_3648, i_10_3649, i_10_3721, i_10_3839, i_10_3841, i_10_3852, i_10_3856, i_10_3857, i_10_3978, i_10_3979, i_10_3980, i_10_3982, i_10_3987, i_10_3991, i_10_4026, i_10_4027, i_10_4028, i_10_4051, i_10_4053, i_10_4266, i_10_4275, i_10_4276, i_10_4277, i_10_4287, i_10_4554, o_10_90);
	kernel_10_91 k_10_91(i_10_173, i_10_266, i_10_283, i_10_316, i_10_387, i_10_438, i_10_447, i_10_578, i_10_697, i_10_698, i_10_733, i_10_734, i_10_754, i_10_928, i_10_997, i_10_1040, i_10_1043, i_10_1138, i_10_1167, i_10_1205, i_10_1234, i_10_1237, i_10_1309, i_10_1344, i_10_1346, i_10_1384, i_10_1403, i_10_1550, i_10_1552, i_10_1553, i_10_1745, i_10_1766, i_10_1825, i_10_1910, i_10_1958, i_10_2092, i_10_2159, i_10_2209, i_10_2330, i_10_2361, i_10_2377, i_10_2450, i_10_2452, i_10_2527, i_10_2539, i_10_2540, i_10_2543, i_10_2616, i_10_2630, i_10_2632, i_10_2660, i_10_2677, i_10_2714, i_10_2731, i_10_2755, i_10_2817, i_10_2818, i_10_2882, i_10_2920, i_10_3041, i_10_3047, i_10_3074, i_10_3087, i_10_3088, i_10_3089, i_10_3092, i_10_3198, i_10_3199, i_10_3280, i_10_3330, i_10_3331, i_10_3350, i_10_3353, i_10_3359, i_10_3404, i_10_3405, i_10_3503, i_10_3524, i_10_3539, i_10_3551, i_10_3555, i_10_3614, i_10_3859, i_10_3860, i_10_3899, i_10_3983, i_10_3992, i_10_4057, i_10_4167, i_10_4271, i_10_4282, i_10_4292, i_10_4376, i_10_4379, i_10_4382, i_10_4554, i_10_4568, i_10_4574, i_10_4576, i_10_4577, o_10_91);
	kernel_10_92 k_10_92(i_10_27, i_10_156, i_10_180, i_10_258, i_10_267, i_10_268, i_10_280, i_10_292, i_10_331, i_10_348, i_10_363, i_10_425, i_10_444, i_10_446, i_10_449, i_10_562, i_10_564, i_10_565, i_10_669, i_10_910, i_10_918, i_10_933, i_10_958, i_10_988, i_10_999, i_10_1000, i_10_1047, i_10_1052, i_10_1105, i_10_1305, i_10_1306, i_10_1311, i_10_1326, i_10_1457, i_10_1614, i_10_1615, i_10_1684, i_10_1685, i_10_1818, i_10_1899, i_10_1942, i_10_1948, i_10_1992, i_10_2001, i_10_2020, i_10_2079, i_10_2142, i_10_2182, i_10_2186, i_10_2239, i_10_2326, i_10_2350, i_10_2351, i_10_2352, i_10_2409, i_10_2452, i_10_2469, i_10_2582, i_10_2605, i_10_2611, i_10_2614, i_10_2615, i_10_2703, i_10_2754, i_10_2787, i_10_3009, i_10_3039, i_10_3069, i_10_3090, i_10_3195, i_10_3283, i_10_3297, i_10_3301, i_10_3325, i_10_3448, i_10_3495, i_10_3499, i_10_3558, i_10_3561, i_10_3588, i_10_3589, i_10_3609, i_10_3610, i_10_3637, i_10_3695, i_10_3699, i_10_3852, i_10_3882, i_10_3945, i_10_3982, i_10_4027, i_10_4050, i_10_4067, i_10_4186, i_10_4293, i_10_4372, i_10_4373, i_10_4449, i_10_4457, i_10_4530, o_10_92);
	kernel_10_93 k_10_93(i_10_82, i_10_221, i_10_281, i_10_283, i_10_409, i_10_423, i_10_424, i_10_446, i_10_448, i_10_495, i_10_505, i_10_513, i_10_794, i_10_964, i_10_1236, i_10_1240, i_10_1260, i_10_1309, i_10_1342, i_10_1359, i_10_1377, i_10_1444, i_10_1446, i_10_1450, i_10_1540, i_10_1582, i_10_1655, i_10_1683, i_10_1819, i_10_1820, i_10_1821, i_10_1913, i_10_1944, i_10_1945, i_10_1989, i_10_2026, i_10_2331, i_10_2353, i_10_2364, i_10_2377, i_10_2380, i_10_2403, i_10_2404, i_10_2502, i_10_2503, i_10_2504, i_10_2628, i_10_2632, i_10_2637, i_10_2638, i_10_2655, i_10_2658, i_10_2673, i_10_2674, i_10_2675, i_10_2711, i_10_2718, i_10_2722, i_10_2724, i_10_2727, i_10_2728, i_10_2781, i_10_2827, i_10_2830, i_10_2831, i_10_2881, i_10_2920, i_10_2979, i_10_2980, i_10_3042, i_10_3070, i_10_3073, i_10_3076, i_10_3151, i_10_3195, i_10_3198, i_10_3385, i_10_3586, i_10_3609, i_10_3780, i_10_3781, i_10_3835, i_10_3837, i_10_3838, i_10_3841, i_10_3843, i_10_3852, i_10_3889, i_10_3979, i_10_3980, i_10_4054, i_10_4118, i_10_4122, i_10_4123, i_10_4126, i_10_4289, i_10_4564, i_10_4567, i_10_4568, i_10_4570, o_10_93);
	kernel_10_94 k_10_94(i_10_12, i_10_63, i_10_64, i_10_77, i_10_172, i_10_174, i_10_175, i_10_208, i_10_223, i_10_244, i_10_286, i_10_315, i_10_318, i_10_406, i_10_594, i_10_639, i_10_733, i_10_891, i_10_946, i_10_999, i_10_1000, i_10_1041, i_10_1060, i_10_1174, i_10_1239, i_10_1241, i_10_1242, i_10_1244, i_10_1264, i_10_1267, i_10_1268, i_10_1367, i_10_1382, i_10_1545, i_10_1579, i_10_1593, i_10_1611, i_10_1633, i_10_1653, i_10_1654, i_10_1696, i_10_1883, i_10_1912, i_10_1919, i_10_1953, i_10_1989, i_10_1998, i_10_2106, i_10_2203, i_10_2236, i_10_2245, i_10_2246, i_10_2254, i_10_2448, i_10_2459, i_10_2475, i_10_2502, i_10_2514, i_10_2541, i_10_2565, i_10_2611, i_10_2633, i_10_2659, i_10_2662, i_10_2663, i_10_2676, i_10_2730, i_10_2782, i_10_2807, i_10_2882, i_10_3198, i_10_3202, i_10_3454, i_10_3537, i_10_3540, i_10_3618, i_10_3700, i_10_3771, i_10_3847, i_10_3852, i_10_3854, i_10_3857, i_10_3881, i_10_3897, i_10_3901, i_10_3978, i_10_4118, i_10_4150, i_10_4152, i_10_4153, i_10_4155, i_10_4158, i_10_4173, i_10_4174, i_10_4213, i_10_4266, i_10_4410, i_10_4431, i_10_4438, i_10_4528, o_10_94);
	kernel_10_95 k_10_95(i_10_146, i_10_280, i_10_315, i_10_316, i_10_318, i_10_319, i_10_406, i_10_411, i_10_412, i_10_427, i_10_441, i_10_442, i_10_444, i_10_445, i_10_448, i_10_460, i_10_461, i_10_462, i_10_588, i_10_712, i_10_715, i_10_716, i_10_747, i_10_793, i_10_795, i_10_796, i_10_798, i_10_828, i_10_927, i_10_963, i_10_966, i_10_967, i_10_993, i_10_1002, i_10_1003, i_10_1116, i_10_1234, i_10_1235, i_10_1341, i_10_1344, i_10_1444, i_10_1649, i_10_1650, i_10_1651, i_10_1652, i_10_1685, i_10_1686, i_10_1687, i_10_1818, i_10_1821, i_10_1945, i_10_1949, i_10_2154, i_10_2181, i_10_2334, i_10_2335, i_10_2337, i_10_2338, i_10_2350, i_10_2379, i_10_2383, i_10_2407, i_10_2449, i_10_2451, i_10_2452, i_10_2473, i_10_2474, i_10_2629, i_10_2631, i_10_2632, i_10_2634, i_10_2658, i_10_2661, i_10_2662, i_10_2712, i_10_2733, i_10_2734, i_10_2784, i_10_2826, i_10_2880, i_10_2917, i_10_2984, i_10_3039, i_10_3270, i_10_3387, i_10_3402, i_10_3405, i_10_3582, i_10_3583, i_10_3585, i_10_3586, i_10_3589, i_10_3590, i_10_3613, i_10_3727, i_10_3787, i_10_4266, i_10_4284, i_10_4285, i_10_4459, o_10_95);
	kernel_10_96 k_10_96(i_10_174, i_10_175, i_10_176, i_10_177, i_10_221, i_10_224, i_10_283, i_10_328, i_10_329, i_10_331, i_10_391, i_10_408, i_10_410, i_10_428, i_10_797, i_10_898, i_10_1236, i_10_1238, i_10_1544, i_10_1552, i_10_1555, i_10_1579, i_10_1650, i_10_1655, i_10_1690, i_10_1769, i_10_1821, i_10_1822, i_10_1823, i_10_1945, i_10_1997, i_10_2024, i_10_2026, i_10_2311, i_10_2352, i_10_2353, i_10_2354, i_10_2356, i_10_2410, i_10_2453, i_10_2467, i_10_2468, i_10_2473, i_10_2603, i_10_2631, i_10_2632, i_10_2633, i_10_2656, i_10_2680, i_10_2706, i_10_2707, i_10_2783, i_10_2785, i_10_2786, i_10_2827, i_10_2828, i_10_2830, i_10_2920, i_10_2923, i_10_2924, i_10_3038, i_10_3044, i_10_3152, i_10_3153, i_10_3156, i_10_3157, i_10_3201, i_10_3387, i_10_3389, i_10_3583, i_10_3584, i_10_3612, i_10_3613, i_10_3614, i_10_3844, i_10_3846, i_10_3847, i_10_3848, i_10_3851, i_10_3852, i_10_3856, i_10_3991, i_10_3992, i_10_4119, i_10_4122, i_10_4125, i_10_4129, i_10_4130, i_10_4269, i_10_4270, i_10_4271, i_10_4276, i_10_4277, i_10_4286, i_10_4288, i_10_4289, i_10_4563, i_10_4564, i_10_4567, i_10_4568, o_10_96);
	kernel_10_97 k_10_97(i_10_49, i_10_123, i_10_124, i_10_171, i_10_217, i_10_218, i_10_244, i_10_293, i_10_317, i_10_320, i_10_325, i_10_431, i_10_432, i_10_462, i_10_512, i_10_990, i_10_1084, i_10_1306, i_10_1450, i_10_1576, i_10_1577, i_10_1619, i_10_1621, i_10_1649, i_10_1685, i_10_1687, i_10_1767, i_10_1820, i_10_1823, i_10_1990, i_10_1991, i_10_2003, i_10_2312, i_10_2351, i_10_2359, i_10_2360, i_10_2362, i_10_2363, i_10_2377, i_10_2449, i_10_2462, i_10_2468, i_10_2510, i_10_2628, i_10_2636, i_10_2639, i_10_2681, i_10_2711, i_10_2712, i_10_2713, i_10_2723, i_10_2731, i_10_2828, i_10_2831, i_10_2881, i_10_2882, i_10_2916, i_10_2917, i_10_2918, i_10_2919, i_10_2921, i_10_2924, i_10_3069, i_10_3198, i_10_3200, i_10_3269, i_10_3273, i_10_3289, i_10_3290, i_10_3402, i_10_3404, i_10_3406, i_10_3407, i_10_3538, i_10_3610, i_10_3611, i_10_3648, i_10_3649, i_10_3731, i_10_3734, i_10_3787, i_10_3788, i_10_3815, i_10_3835, i_10_3846, i_10_3910, i_10_3981, i_10_3982, i_10_3983, i_10_3986, i_10_3991, i_10_4027, i_10_4028, i_10_4030, i_10_4031, i_10_4121, i_10_4127, i_10_4214, i_10_4274, i_10_4290, o_10_97);
	kernel_10_98 k_10_98(i_10_48, i_10_173, i_10_181, i_10_223, i_10_287, i_10_319, i_10_320, i_10_347, i_10_393, i_10_442, i_10_445, i_10_448, i_10_463, i_10_716, i_10_719, i_10_793, i_10_799, i_10_827, i_10_832, i_10_963, i_10_964, i_10_967, i_10_1081, i_10_1085, i_10_1238, i_10_1248, i_10_1249, i_10_1309, i_10_1313, i_10_1364, i_10_1367, i_10_1438, i_10_1575, i_10_1579, i_10_1616, i_10_1641, i_10_1642, i_10_1648, i_10_1685, i_10_1687, i_10_1689, i_10_1821, i_10_1908, i_10_1916, i_10_1948, i_10_2020, i_10_2455, i_10_2470, i_10_2508, i_10_2520, i_10_2604, i_10_2634, i_10_2704, i_10_2714, i_10_2726, i_10_2729, i_10_2828, i_10_2884, i_10_2885, i_10_2888, i_10_2916, i_10_2923, i_10_2924, i_10_2958, i_10_3037, i_10_3196, i_10_3270, i_10_3284, i_10_3384, i_10_3388, i_10_3429, i_10_3446, i_10_3505, i_10_3522, i_10_3523, i_10_3559, i_10_3561, i_10_3563, i_10_3589, i_10_3614, i_10_3650, i_10_3651, i_10_3652, i_10_3810, i_10_3811, i_10_3859, i_10_3860, i_10_3948, i_10_3949, i_10_3978, i_10_3981, i_10_4050, i_10_4114, i_10_4117, i_10_4204, i_10_4217, i_10_4284, i_10_4288, i_10_4291, i_10_4292, o_10_98);
	kernel_10_99 k_10_99(i_10_39, i_10_121, i_10_148, i_10_149, i_10_157, i_10_188, i_10_244, i_10_256, i_10_257, i_10_271, i_10_394, i_10_395, i_10_445, i_10_544, i_10_585, i_10_598, i_10_601, i_10_602, i_10_688, i_10_734, i_10_800, i_10_880, i_10_1003, i_10_1013, i_10_1154, i_10_1241, i_10_1242, i_10_1249, i_10_1281, i_10_1438, i_10_1441, i_10_1516, i_10_1542, i_10_1544, i_10_1560, i_10_1565, i_10_1580, i_10_1612, i_10_1615, i_10_1616, i_10_1686, i_10_1819, i_10_1822, i_10_1823, i_10_1885, i_10_1920, i_10_1959, i_10_1961, i_10_2020, i_10_2023, i_10_2349, i_10_2350, i_10_2353, i_10_2354, i_10_2408, i_10_2518, i_10_2532, i_10_2535, i_10_2536, i_10_2537, i_10_2629, i_10_2632, i_10_2634, i_10_2696, i_10_2713, i_10_2734, i_10_2735, i_10_2821, i_10_2833, i_10_2870, i_10_2884, i_10_2984, i_10_3199, i_10_3269, i_10_3392, i_10_3431, i_10_3433, i_10_3496, i_10_3524, i_10_3582, i_10_3609, i_10_3784, i_10_3881, i_10_3944, i_10_3982, i_10_4013, i_10_4113, i_10_4114, i_10_4117, i_10_4175, i_10_4178, i_10_4186, i_10_4214, i_10_4267, i_10_4270, i_10_4273, i_10_4522, i_10_4564, i_10_4565, i_10_4566, o_10_99);
	kernel_10_100 k_10_100(i_10_27, i_10_251, i_10_406, i_10_408, i_10_432, i_10_441, i_10_444, i_10_445, i_10_730, i_10_755, i_10_954, i_10_1000, i_10_1001, i_10_1005, i_10_1083, i_10_1234, i_10_1235, i_10_1241, i_10_1274, i_10_1307, i_10_1310, i_10_1313, i_10_1546, i_10_1547, i_10_1549, i_10_1550, i_10_1552, i_10_1612, i_10_1613, i_10_1649, i_10_1655, i_10_1677, i_10_1684, i_10_1690, i_10_1720, i_10_1823, i_10_1944, i_10_1945, i_10_1946, i_10_2083, i_10_2152, i_10_2179, i_10_2180, i_10_2200, i_10_2201, i_10_2306, i_10_2380, i_10_2405, i_10_2407, i_10_2449, i_10_2453, i_10_2459, i_10_2472, i_10_2474, i_10_2632, i_10_2654, i_10_2722, i_10_2723, i_10_2731, i_10_2741, i_10_2826, i_10_2827, i_10_2830, i_10_2831, i_10_2885, i_10_2917, i_10_2952, i_10_2953, i_10_3051, i_10_3054, i_10_3055, i_10_3167, i_10_3277, i_10_3281, i_10_3298, i_10_3387, i_10_3391, i_10_3392, i_10_3467, i_10_3470, i_10_3472, i_10_3584, i_10_3587, i_10_3611, i_10_3612, i_10_3650, i_10_3838, i_10_3854, i_10_3855, i_10_3859, i_10_3990, i_10_3991, i_10_3992, i_10_4052, i_10_4054, i_10_4113, i_10_4117, i_10_4214, i_10_4230, i_10_4266, o_10_100);
	kernel_10_101 k_10_101(i_10_36, i_10_37, i_10_155, i_10_172, i_10_175, i_10_176, i_10_221, i_10_281, i_10_282, i_10_296, i_10_315, i_10_316, i_10_390, i_10_434, i_10_438, i_10_442, i_10_793, i_10_796, i_10_797, i_10_800, i_10_899, i_10_990, i_10_996, i_10_1085, i_10_1153, i_10_1237, i_10_1238, i_10_1239, i_10_1306, i_10_1341, i_10_1345, i_10_1349, i_10_1441, i_10_1551, i_10_1654, i_10_1655, i_10_1676, i_10_1686, i_10_1825, i_10_1910, i_10_1944, i_10_2005, i_10_2019, i_10_2352, i_10_2356, i_10_2365, i_10_2514, i_10_2628, i_10_2629, i_10_2630, i_10_2631, i_10_2632, i_10_2633, i_10_2636, i_10_2657, i_10_2661, i_10_2673, i_10_2703, i_10_2704, i_10_2705, i_10_2711, i_10_2729, i_10_2783, i_10_2829, i_10_2831, i_10_2885, i_10_2916, i_10_2923, i_10_2984, i_10_3034, i_10_3035, i_10_3069, i_10_3070, i_10_3198, i_10_3234, i_10_3270, i_10_3280, i_10_3384, i_10_3522, i_10_3540, i_10_3583, i_10_3609, i_10_3612, i_10_3613, i_10_3647, i_10_3837, i_10_3839, i_10_3853, i_10_3855, i_10_3856, i_10_3860, i_10_3872, i_10_4122, i_10_4123, i_10_4125, i_10_4126, i_10_4167, i_10_4168, i_10_4287, i_10_4566, o_10_101);
	kernel_10_102 k_10_102(i_10_27, i_10_31, i_10_81, i_10_121, i_10_126, i_10_172, i_10_174, i_10_181, i_10_182, i_10_281, i_10_282, i_10_324, i_10_370, i_10_373, i_10_387, i_10_432, i_10_433, i_10_445, i_10_495, i_10_516, i_10_684, i_10_931, i_10_957, i_10_960, i_10_961, i_10_1086, i_10_1233, i_10_1236, i_10_1237, i_10_1324, i_10_1362, i_10_1364, i_10_1432, i_10_1530, i_10_1543, i_10_1548, i_10_1683, i_10_1687, i_10_1822, i_10_1824, i_10_1825, i_10_1917, i_10_1936, i_10_1939, i_10_1944, i_10_1945, i_10_1948, i_10_1949, i_10_1954, i_10_2025, i_10_2179, i_10_2304, i_10_2305, i_10_2329, i_10_2361, i_10_2377, i_10_2403, i_10_2453, i_10_2539, i_10_2556, i_10_2612, i_10_2820, i_10_2827, i_10_2828, i_10_2910, i_10_2911, i_10_3007, i_10_3042, i_10_3087, i_10_3088, i_10_3234, i_10_3313, i_10_3351, i_10_3438, i_10_3439, i_10_3447, i_10_3465, i_10_3466, i_10_3519, i_10_3582, i_10_3585, i_10_3615, i_10_3649, i_10_3786, i_10_3856, i_10_3942, i_10_3943, i_10_3945, i_10_3982, i_10_4023, i_10_4027, i_10_4230, i_10_4232, i_10_4369, i_10_4437, i_10_4446, i_10_4528, i_10_4529, i_10_4566, i_10_4581, o_10_102);
	kernel_10_103 k_10_103(i_10_216, i_10_218, i_10_247, i_10_279, i_10_284, i_10_319, i_10_429, i_10_430, i_10_435, i_10_438, i_10_439, i_10_449, i_10_463, i_10_466, i_10_748, i_10_961, i_10_993, i_10_996, i_10_1059, i_10_1238, i_10_1250, i_10_1354, i_10_1357, i_10_1556, i_10_1684, i_10_1685, i_10_1756, i_10_1818, i_10_1821, i_10_1824, i_10_1825, i_10_1912, i_10_1916, i_10_1947, i_10_1990, i_10_2312, i_10_2353, i_10_2355, i_10_2373, i_10_2451, i_10_2452, i_10_2454, i_10_2469, i_10_2514, i_10_2516, i_10_2546, i_10_2659, i_10_2660, i_10_2701, i_10_2704, i_10_2711, i_10_2720, i_10_2728, i_10_2729, i_10_2820, i_10_2821, i_10_2884, i_10_3039, i_10_3049, i_10_3093, i_10_3094, i_10_3174, i_10_3195, i_10_3235, i_10_3271, i_10_3279, i_10_3280, i_10_3281, i_10_3282, i_10_3283, i_10_3292, i_10_3318, i_10_3384, i_10_3385, i_10_3388, i_10_3389, i_10_3390, i_10_3525, i_10_3526, i_10_3616, i_10_3617, i_10_3685, i_10_3702, i_10_3705, i_10_3850, i_10_3857, i_10_3859, i_10_3885, i_10_3902, i_10_3946, i_10_4027, i_10_4031, i_10_4056, i_10_4116, i_10_4117, i_10_4213, i_10_4271, i_10_4567, i_10_4568, i_10_4589, o_10_103);
	kernel_10_104 k_10_104(i_10_117, i_10_118, i_10_220, i_10_315, i_10_316, i_10_387, i_10_388, i_10_389, i_10_391, i_10_394, i_10_408, i_10_427, i_10_436, i_10_462, i_10_532, i_10_795, i_10_819, i_10_824, i_10_958, i_10_999, i_10_1000, i_10_1026, i_10_1080, i_10_1236, i_10_1296, i_10_1305, i_10_1306, i_10_1308, i_10_1378, i_10_1431, i_10_1448, i_10_1543, i_10_1575, i_10_1576, i_10_1578, i_10_1621, i_10_1651, i_10_1683, i_10_1684, i_10_1685, i_10_1729, i_10_1732, i_10_1733, i_10_1764, i_10_1819, i_10_2022, i_10_2028, i_10_2200, i_10_2203, i_10_2204, i_10_2250, i_10_2352, i_10_2377, i_10_2405, i_10_2410, i_10_2452, i_10_2454, i_10_2455, i_10_2467, i_10_2540, i_10_2556, i_10_2565, i_10_2628, i_10_2629, i_10_2719, i_10_2727, i_10_2729, i_10_2781, i_10_2782, i_10_2785, i_10_2863, i_10_2880, i_10_2980, i_10_3042, i_10_3195, i_10_3313, i_10_3389, i_10_3392, i_10_3466, i_10_3469, i_10_3501, i_10_3522, i_10_3550, i_10_3559, i_10_3582, i_10_3583, i_10_3840, i_10_3841, i_10_3857, i_10_4006, i_10_4023, i_10_4024, i_10_4113, i_10_4115, i_10_4117, i_10_4118, i_10_4204, i_10_4275, i_10_4289, i_10_4581, o_10_104);
	kernel_10_105 k_10_105(i_10_37, i_10_256, i_10_283, i_10_318, i_10_322, i_10_324, i_10_325, i_10_328, i_10_405, i_10_441, i_10_444, i_10_460, i_10_464, i_10_588, i_10_894, i_10_954, i_10_993, i_10_1003, i_10_1031, i_10_1086, i_10_1241, i_10_1377, i_10_1378, i_10_1435, i_10_1542, i_10_1543, i_10_1546, i_10_1579, i_10_1580, i_10_1581, i_10_1582, i_10_1596, i_10_1612, i_10_1647, i_10_1648, i_10_1649, i_10_1654, i_10_1689, i_10_1768, i_10_1822, i_10_1824, i_10_1825, i_10_1947, i_10_1948, i_10_1992, i_10_1995, i_10_2200, i_10_2203, i_10_2242, i_10_2309, i_10_2330, i_10_2352, i_10_2353, i_10_2356, i_10_2364, i_10_2452, i_10_2453, i_10_2454, i_10_2455, i_10_2458, i_10_2471, i_10_2473, i_10_2541, i_10_2604, i_10_2607, i_10_2658, i_10_2714, i_10_2787, i_10_2829, i_10_2831, i_10_2917, i_10_2982, i_10_3270, i_10_3274, i_10_3281, i_10_3282, i_10_3525, i_10_3526, i_10_3614, i_10_3616, i_10_3683, i_10_3780, i_10_3787, i_10_3840, i_10_3841, i_10_3848, i_10_3854, i_10_3857, i_10_3859, i_10_3891, i_10_3893, i_10_3979, i_10_3982, i_10_4233, i_10_4287, i_10_4292, i_10_4456, i_10_4459, i_10_4566, i_10_4570, o_10_105);
	kernel_10_106 k_10_106(i_10_175, i_10_268, i_10_280, i_10_285, i_10_296, i_10_316, i_10_317, i_10_327, i_10_328, i_10_329, i_10_409, i_10_439, i_10_443, i_10_453, i_10_516, i_10_520, i_10_749, i_10_800, i_10_999, i_10_1080, i_10_1081, i_10_1217, i_10_1233, i_10_1234, i_10_1238, i_10_1263, i_10_1264, i_10_1265, i_10_1366, i_10_1438, i_10_1439, i_10_1448, i_10_1546, i_10_1615, i_10_1684, i_10_1687, i_10_1688, i_10_1818, i_10_1819, i_10_1821, i_10_1822, i_10_1826, i_10_2337, i_10_2351, i_10_2352, i_10_2353, i_10_2354, i_10_2408, i_10_2461, i_10_2470, i_10_2606, i_10_2655, i_10_2658, i_10_2659, i_10_2660, i_10_2680, i_10_2707, i_10_2722, i_10_2723, i_10_2729, i_10_2827, i_10_2828, i_10_2831, i_10_2885, i_10_2979, i_10_2980, i_10_2981, i_10_2985, i_10_2986, i_10_2987, i_10_3070, i_10_3074, i_10_3157, i_10_3158, i_10_3198, i_10_3199, i_10_3200, i_10_3201, i_10_3274, i_10_3280, i_10_3281, i_10_3384, i_10_3385, i_10_3388, i_10_3493, i_10_3496, i_10_3497, i_10_3522, i_10_3583, i_10_3837, i_10_3851, i_10_3858, i_10_3872, i_10_3896, i_10_3906, i_10_3979, i_10_4266, i_10_4270, i_10_4277, i_10_4279, o_10_106);
	kernel_10_107 k_10_107(i_10_176, i_10_187, i_10_283, i_10_319, i_10_390, i_10_391, i_10_392, i_10_405, i_10_409, i_10_424, i_10_426, i_10_427, i_10_433, i_10_434, i_10_459, i_10_462, i_10_794, i_10_991, i_10_1026, i_10_1027, i_10_1031, i_10_1043, i_10_1081, i_10_1135, i_10_1306, i_10_1442, i_10_1540, i_10_1541, i_10_1548, i_10_1575, i_10_1577, i_10_1651, i_10_1683, i_10_1684, i_10_1685, i_10_1769, i_10_1825, i_10_1990, i_10_2349, i_10_2353, i_10_2356, i_10_2360, i_10_2404, i_10_2448, i_10_2631, i_10_2632, i_10_2633, i_10_2673, i_10_2674, i_10_2675, i_10_2681, i_10_2701, i_10_2703, i_10_2723, i_10_2727, i_10_2783, i_10_2887, i_10_2918, i_10_2921, i_10_3069, i_10_3071, i_10_3073, i_10_3152, i_10_3153, i_10_3156, i_10_3158, i_10_3268, i_10_3269, i_10_3322, i_10_3328, i_10_3330, i_10_3406, i_10_3585, i_10_3586, i_10_3612, i_10_3614, i_10_3616, i_10_3649, i_10_3780, i_10_3782, i_10_3783, i_10_3784, i_10_3785, i_10_3835, i_10_3837, i_10_3838, i_10_3839, i_10_3855, i_10_3856, i_10_3857, i_10_3980, i_10_4117, i_10_4118, i_10_4119, i_10_4120, i_10_4121, i_10_4266, i_10_4276, i_10_4288, i_10_4567, o_10_107);
	kernel_10_108 k_10_108(i_10_123, i_10_153, i_10_171, i_10_175, i_10_244, i_10_248, i_10_434, i_10_436, i_10_519, i_10_799, i_10_963, i_10_1036, i_10_1120, i_10_1234, i_10_1306, i_10_1308, i_10_1363, i_10_1365, i_10_1431, i_10_1447, i_10_1554, i_10_1612, i_10_1653, i_10_1654, i_10_1655, i_10_1687, i_10_1690, i_10_1820, i_10_1821, i_10_1944, i_10_1945, i_10_1950, i_10_1953, i_10_2199, i_10_2200, i_10_2204, i_10_2307, i_10_2361, i_10_2407, i_10_2470, i_10_2514, i_10_2607, i_10_2630, i_10_2636, i_10_2660, i_10_2679, i_10_2701, i_10_2722, i_10_2724, i_10_2725, i_10_2726, i_10_2727, i_10_2821, i_10_2874, i_10_2885, i_10_2923, i_10_2994, i_10_3036, i_10_3072, i_10_3073, i_10_3090, i_10_3195, i_10_3198, i_10_3203, i_10_3278, i_10_3282, i_10_3298, i_10_3388, i_10_3429, i_10_3430, i_10_3436, i_10_3467, i_10_3468, i_10_3471, i_10_3472, i_10_3498, i_10_3522, i_10_3612, i_10_3621, i_10_3646, i_10_3648, i_10_3649, i_10_3651, i_10_3723, i_10_3726, i_10_3783, i_10_3834, i_10_3853, i_10_3855, i_10_3859, i_10_3860, i_10_3909, i_10_3983, i_10_4171, i_10_4174, i_10_4213, i_10_4216, i_10_4273, i_10_4277, i_10_4291, o_10_108);
	kernel_10_109 k_10_109(i_10_39, i_10_63, i_10_64, i_10_172, i_10_316, i_10_405, i_10_408, i_10_409, i_10_432, i_10_433, i_10_436, i_10_659, i_10_712, i_10_796, i_10_797, i_10_990, i_10_991, i_10_993, i_10_1026, i_10_1154, i_10_1234, i_10_1238, i_10_1306, i_10_1359, i_10_1360, i_10_1362, i_10_1433, i_10_1442, i_10_1539, i_10_1541, i_10_1542, i_10_1544, i_10_1621, i_10_1622, i_10_1683, i_10_1685, i_10_1687, i_10_1688, i_10_1711, i_10_1992, i_10_2016, i_10_2017, i_10_2179, i_10_2197, i_10_2352, i_10_2359, i_10_2362, i_10_2363, i_10_2512, i_10_2566, i_10_2628, i_10_2659, i_10_2718, i_10_2730, i_10_2781, i_10_2829, i_10_2837, i_10_2872, i_10_3042, i_10_3044, i_10_3069, i_10_3070, i_10_3071, i_10_3073, i_10_3074, i_10_3195, i_10_3268, i_10_3331, i_10_3332, i_10_3384, i_10_3538, i_10_3541, i_10_3612, i_10_3785, i_10_3807, i_10_3808, i_10_3838, i_10_3839, i_10_3850, i_10_3853, i_10_3855, i_10_3857, i_10_3880, i_10_3980, i_10_3991, i_10_4113, i_10_4114, i_10_4115, i_10_4116, i_10_4122, i_10_4172, i_10_4175, i_10_4230, i_10_4275, i_10_4285, i_10_4292, i_10_4437, i_10_4567, i_10_4568, i_10_4569, o_10_109);
	kernel_10_110 k_10_110(i_10_31, i_10_37, i_10_178, i_10_218, i_10_220, i_10_224, i_10_319, i_10_406, i_10_407, i_10_448, i_10_514, i_10_602, i_10_711, i_10_713, i_10_714, i_10_732, i_10_794, i_10_797, i_10_800, i_10_828, i_10_830, i_10_963, i_10_1239, i_10_1363, i_10_1454, i_10_1579, i_10_1647, i_10_1649, i_10_1683, i_10_1684, i_10_1685, i_10_1687, i_10_1688, i_10_1691, i_10_1719, i_10_1765, i_10_1766, i_10_1801, i_10_1802, i_10_1805, i_10_1821, i_10_1915, i_10_1939, i_10_2096, i_10_2307, i_10_2308, i_10_2448, i_10_2449, i_10_2450, i_10_2468, i_10_2539, i_10_2542, i_10_2659, i_10_2723, i_10_2725, i_10_2726, i_10_2728, i_10_2734, i_10_2781, i_10_2782, i_10_2784, i_10_2788, i_10_2820, i_10_2832, i_10_2985, i_10_3199, i_10_3270, i_10_3279, i_10_3280, i_10_3281, i_10_3283, i_10_3291, i_10_3325, i_10_3384, i_10_3390, i_10_3406, i_10_3409, i_10_3430, i_10_3494, i_10_3523, i_10_3539, i_10_3616, i_10_3649, i_10_3725, i_10_3727, i_10_3781, i_10_3852, i_10_3854, i_10_3857, i_10_3858, i_10_3906, i_10_3982, i_10_4054, i_10_4121, i_10_4238, i_10_4268, i_10_4285, i_10_4286, i_10_4289, i_10_4477, o_10_110);
	kernel_10_111 k_10_111(i_10_171, i_10_174, i_10_175, i_10_177, i_10_178, i_10_179, i_10_248, i_10_281, i_10_284, i_10_293, i_10_315, i_10_316, i_10_318, i_10_319, i_10_409, i_10_411, i_10_412, i_10_459, i_10_466, i_10_797, i_10_799, i_10_957, i_10_994, i_10_1087, i_10_1156, i_10_1237, i_10_1238, i_10_1240, i_10_1250, i_10_1268, i_10_1313, i_10_1344, i_10_1347, i_10_1348, i_10_1442, i_10_1445, i_10_1577, i_10_1580, i_10_1685, i_10_1686, i_10_1714, i_10_1821, i_10_1825, i_10_1872, i_10_1874, i_10_1995, i_10_2198, i_10_2334, i_10_2358, i_10_2365, i_10_2472, i_10_2517, i_10_2518, i_10_2519, i_10_2605, i_10_2629, i_10_2631, i_10_2632, i_10_2634, i_10_2635, i_10_2636, i_10_2674, i_10_2700, i_10_2704, i_10_2710, i_10_2711, i_10_2723, i_10_2724, i_10_2781, i_10_2782, i_10_2785, i_10_2832, i_10_3072, i_10_3073, i_10_3201, i_10_3279, i_10_3319, i_10_3385, i_10_3431, i_10_3497, i_10_3543, i_10_3562, i_10_3586, i_10_3611, i_10_3617, i_10_3841, i_10_3893, i_10_3942, i_10_3943, i_10_4116, i_10_4117, i_10_4118, i_10_4120, i_10_4121, i_10_4128, i_10_4129, i_10_4130, i_10_4173, i_10_4281, i_10_4291, o_10_111);
	kernel_10_112 k_10_112(i_10_41, i_10_64, i_10_216, i_10_317, i_10_431, i_10_433, i_10_437, i_10_442, i_10_443, i_10_538, i_10_895, i_10_992, i_10_1034, i_10_1119, i_10_1239, i_10_1308, i_10_1309, i_10_1311, i_10_1378, i_10_1456, i_10_1653, i_10_1655, i_10_1676, i_10_1683, i_10_1684, i_10_1690, i_10_1809, i_10_1822, i_10_1824, i_10_1950, i_10_2110, i_10_2202, i_10_2261, i_10_2359, i_10_2361, i_10_2461, i_10_2467, i_10_2572, i_10_2641, i_10_2658, i_10_2659, i_10_2710, i_10_2726, i_10_2727, i_10_2733, i_10_2826, i_10_2827, i_10_2829, i_10_2830, i_10_2831, i_10_2835, i_10_2852, i_10_2920, i_10_2982, i_10_2993, i_10_3042, i_10_3048, i_10_3073, i_10_3093, i_10_3197, i_10_3198, i_10_3199, i_10_3200, i_10_3271, i_10_3454, i_10_3541, i_10_3561, i_10_3609, i_10_3612, i_10_3703, i_10_3775, i_10_3838, i_10_3839, i_10_3854, i_10_3855, i_10_3856, i_10_3859, i_10_3860, i_10_3990, i_10_3991, i_10_4029, i_10_4030, i_10_4031, i_10_4116, i_10_4117, i_10_4119, i_10_4120, i_10_4129, i_10_4159, i_10_4171, i_10_4172, i_10_4173, i_10_4174, i_10_4232, i_10_4279, i_10_4290, i_10_4439, i_10_4529, i_10_4564, i_10_4597, o_10_112);
	kernel_10_113 k_10_113(i_10_35, i_10_124, i_10_178, i_10_249, i_10_282, i_10_283, i_10_284, i_10_286, i_10_319, i_10_322, i_10_324, i_10_408, i_10_409, i_10_430, i_10_437, i_10_444, i_10_445, i_10_446, i_10_460, i_10_967, i_10_993, i_10_1000, i_10_1002, i_10_1005, i_10_1006, i_10_1233, i_10_1237, i_10_1247, i_10_1249, i_10_1310, i_10_1576, i_10_1582, i_10_1617, i_10_1650, i_10_1818, i_10_1819, i_10_1821, i_10_1822, i_10_1823, i_10_1912, i_10_1913, i_10_1950, i_10_1951, i_10_2179, i_10_2180, i_10_2184, i_10_2334, i_10_2338, i_10_2349, i_10_2381, i_10_2382, i_10_2383, i_10_2407, i_10_2409, i_10_2410, i_10_2449, i_10_2454, i_10_2629, i_10_2635, i_10_2636, i_10_2655, i_10_2679, i_10_2706, i_10_2710, i_10_2716, i_10_2728, i_10_2730, i_10_2829, i_10_2917, i_10_3039, i_10_3049, i_10_3094, i_10_3095, i_10_3153, i_10_3154, i_10_3155, i_10_3198, i_10_3200, i_10_3237, i_10_3269, i_10_3270, i_10_3280, i_10_3388, i_10_3389, i_10_3390, i_10_3404, i_10_3405, i_10_3526, i_10_3582, i_10_3613, i_10_3616, i_10_3783, i_10_3837, i_10_3838, i_10_3839, i_10_3847, i_10_3853, i_10_3856, i_10_4120, i_10_4268, o_10_113);
	kernel_10_114 k_10_114(i_10_27, i_10_28, i_10_30, i_10_291, i_10_319, i_10_435, i_10_495, i_10_712, i_10_720, i_10_821, i_10_895, i_10_1026, i_10_1234, i_10_1236, i_10_1237, i_10_1278, i_10_1308, i_10_1362, i_10_1432, i_10_1434, i_10_1435, i_10_1539, i_10_1540, i_10_1547, i_10_1647, i_10_1653, i_10_1683, i_10_1684, i_10_1765, i_10_1805, i_10_1912, i_10_1920, i_10_1985, i_10_2178, i_10_2179, i_10_2224, i_10_2308, i_10_2349, i_10_2352, i_10_2361, i_10_2431, i_10_2451, i_10_2529, i_10_2566, i_10_2610, i_10_2628, i_10_2650, i_10_2659, i_10_2691, i_10_2713, i_10_2718, i_10_2722, i_10_2736, i_10_2743, i_10_2923, i_10_2924, i_10_2926, i_10_2927, i_10_2934, i_10_2943, i_10_2944, i_10_3037, i_10_3078, i_10_3199, i_10_3200, i_10_3279, i_10_3391, i_10_3392, i_10_3406, i_10_3408, i_10_3465, i_10_3466, i_10_3523, i_10_3610, i_10_3612, i_10_3613, i_10_3614, i_10_3645, i_10_3650, i_10_3681, i_10_3682, i_10_3744, i_10_3781, i_10_3782, i_10_3783, i_10_3807, i_10_3817, i_10_3855, i_10_3856, i_10_3857, i_10_3888, i_10_4005, i_10_4006, i_10_4027, i_10_4114, i_10_4117, i_10_4219, i_10_4275, i_10_4276, i_10_4284, o_10_114);
	kernel_10_115 k_10_115(i_10_45, i_10_46, i_10_48, i_10_49, i_10_175, i_10_217, i_10_247, i_10_285, i_10_289, i_10_291, i_10_405, i_10_406, i_10_407, i_10_412, i_10_442, i_10_443, i_10_463, i_10_465, i_10_797, i_10_799, i_10_999, i_10_1002, i_10_1030, i_10_1035, i_10_1234, i_10_1238, i_10_1363, i_10_1436, i_10_1655, i_10_1688, i_10_1821, i_10_1909, i_10_1914, i_10_1915, i_10_1993, i_10_1994, i_10_2186, i_10_2362, i_10_2365, i_10_2449, i_10_2458, i_10_2460, i_10_2468, i_10_2471, i_10_2473, i_10_2474, i_10_2481, i_10_2546, i_10_2572, i_10_2608, i_10_2650, i_10_2661, i_10_2662, i_10_2674, i_10_2710, i_10_2711, i_10_2718, i_10_2720, i_10_2723, i_10_2781, i_10_2820, i_10_2920, i_10_2921, i_10_2924, i_10_3070, i_10_3195, i_10_3267, i_10_3268, i_10_3276, i_10_3388, i_10_3389, i_10_3390, i_10_3402, i_10_3406, i_10_3407, i_10_3467, i_10_3587, i_10_3611, i_10_3619, i_10_3688, i_10_3734, i_10_3842, i_10_3851, i_10_3852, i_10_3858, i_10_3859, i_10_3910, i_10_3929, i_10_3981, i_10_3982, i_10_4117, i_10_4119, i_10_4120, i_10_4121, i_10_4126, i_10_4129, i_10_4290, i_10_4291, i_10_4292, i_10_4459, o_10_115);
	kernel_10_116 k_10_116(i_10_174, i_10_175, i_10_177, i_10_260, i_10_268, i_10_283, i_10_294, i_10_321, i_10_363, i_10_438, i_10_439, i_10_459, i_10_465, i_10_466, i_10_510, i_10_597, i_10_749, i_10_897, i_10_993, i_10_1005, i_10_1033, i_10_1034, i_10_1138, i_10_1236, i_10_1239, i_10_1299, i_10_1306, i_10_1311, i_10_1312, i_10_1347, i_10_1365, i_10_1445, i_10_1446, i_10_1455, i_10_1822, i_10_2022, i_10_2112, i_10_2253, i_10_2265, i_10_2293, i_10_2352, i_10_2353, i_10_2364, i_10_2365, i_10_2452, i_10_2454, i_10_2455, i_10_2474, i_10_2479, i_10_2568, i_10_2571, i_10_2604, i_10_2643, i_10_2663, i_10_2680, i_10_2712, i_10_2715, i_10_2734, i_10_2784, i_10_2882, i_10_2884, i_10_2959, i_10_3045, i_10_3048, i_10_3072, i_10_3075, i_10_3198, i_10_3237, i_10_3273, i_10_3275, i_10_3282, i_10_3318, i_10_3336, i_10_3354, i_10_3388, i_10_3390, i_10_3392, i_10_3407, i_10_3470, i_10_3538, i_10_3543, i_10_3559, i_10_3561, i_10_3585, i_10_3813, i_10_3837, i_10_3845, i_10_3859, i_10_3903, i_10_3984, i_10_3985, i_10_3988, i_10_4056, i_10_4117, i_10_4120, i_10_4128, i_10_4173, i_10_4236, i_10_4292, i_10_4434, o_10_116);
	kernel_10_117 k_10_117(i_10_161, i_10_222, i_10_224, i_10_251, i_10_293, i_10_295, i_10_296, i_10_409, i_10_410, i_10_412, i_10_436, i_10_448, i_10_449, i_10_462, i_10_467, i_10_629, i_10_800, i_10_898, i_10_899, i_10_997, i_10_1033, i_10_1034, i_10_1051, i_10_1239, i_10_1263, i_10_1309, i_10_1365, i_10_1435, i_10_1650, i_10_1652, i_10_1654, i_10_1655, i_10_1687, i_10_1816, i_10_1817, i_10_1818, i_10_1912, i_10_1950, i_10_1997, i_10_2360, i_10_2362, i_10_2383, i_10_2455, i_10_2470, i_10_2471, i_10_2472, i_10_2516, i_10_2654, i_10_2658, i_10_2661, i_10_2662, i_10_2680, i_10_2720, i_10_2724, i_10_2725, i_10_2734, i_10_2735, i_10_2833, i_10_2924, i_10_2986, i_10_3153, i_10_3154, i_10_3155, i_10_3157, i_10_3166, i_10_3281, i_10_3544, i_10_3561, i_10_3586, i_10_3589, i_10_3616, i_10_3617, i_10_3720, i_10_3733, i_10_3734, i_10_3784, i_10_3813, i_10_3814, i_10_3815, i_10_3834, i_10_3835, i_10_3836, i_10_3840, i_10_3841, i_10_3842, i_10_4117, i_10_4121, i_10_4129, i_10_4130, i_10_4173, i_10_4174, i_10_4219, i_10_4220, i_10_4266, i_10_4267, i_10_4270, i_10_4289, i_10_4290, i_10_4292, i_10_4566, o_10_117);
	kernel_10_118 k_10_118(i_10_155, i_10_157, i_10_174, i_10_180, i_10_248, i_10_281, i_10_317, i_10_413, i_10_428, i_10_442, i_10_443, i_10_444, i_10_445, i_10_463, i_10_464, i_10_497, i_10_689, i_10_799, i_10_800, i_10_820, i_10_997, i_10_1235, i_10_1237, i_10_1248, i_10_1306, i_10_1354, i_10_1359, i_10_1489, i_10_1543, i_10_1577, i_10_1580, i_10_1683, i_10_1684, i_10_1685, i_10_1686, i_10_1688, i_10_1689, i_10_1914, i_10_1916, i_10_1946, i_10_2019, i_10_2020, i_10_2026, i_10_2351, i_10_2358, i_10_2365, i_10_2378, i_10_2467, i_10_2470, i_10_2515, i_10_2632, i_10_2662, i_10_2704, i_10_2705, i_10_2710, i_10_2723, i_10_2727, i_10_2728, i_10_2735, i_10_2979, i_10_2986, i_10_2987, i_10_3033, i_10_3036, i_10_3202, i_10_3269, i_10_3274, i_10_3277, i_10_3280, i_10_3281, i_10_3314, i_10_3384, i_10_3387, i_10_3522, i_10_3611, i_10_3614, i_10_3728, i_10_3787, i_10_3800, i_10_3836, i_10_3896, i_10_3946, i_10_4114, i_10_4116, i_10_4118, i_10_4123, i_10_4124, i_10_4126, i_10_4127, i_10_4168, i_10_4169, i_10_4171, i_10_4172, i_10_4173, i_10_4270, i_10_4280, i_10_4283, i_10_4284, i_10_4291, i_10_4415, o_10_118);
	kernel_10_119 k_10_119(i_10_250, i_10_286, i_10_446, i_10_448, i_10_462, i_10_754, i_10_755, i_10_795, i_10_796, i_10_904, i_10_955, i_10_956, i_10_957, i_10_958, i_10_997, i_10_1235, i_10_1240, i_10_1552, i_10_1654, i_10_1684, i_10_1686, i_10_1687, i_10_1911, i_10_1912, i_10_1994, i_10_2312, i_10_2357, i_10_2358, i_10_2359, i_10_2360, i_10_2383, i_10_2407, i_10_2437, i_10_2460, i_10_2464, i_10_2467, i_10_2468, i_10_2470, i_10_2536, i_10_2542, i_10_2604, i_10_2630, i_10_2631, i_10_2635, i_10_2660, i_10_2680, i_10_2701, i_10_2722, i_10_2723, i_10_2728, i_10_2729, i_10_2731, i_10_2781, i_10_2917, i_10_2918, i_10_2921, i_10_2923, i_10_2924, i_10_3041, i_10_3197, i_10_3201, i_10_3277, i_10_3387, i_10_3405, i_10_3406, i_10_3467, i_10_3494, i_10_3523, i_10_3583, i_10_3612, i_10_3614, i_10_3705, i_10_3732, i_10_3783, i_10_3784, i_10_3785, i_10_3786, i_10_3807, i_10_3838, i_10_3847, i_10_3851, i_10_3895, i_10_3980, i_10_4113, i_10_4114, i_10_4116, i_10_4117, i_10_4169, i_10_4267, i_10_4270, i_10_4274, i_10_4282, i_10_4283, i_10_4289, i_10_4292, i_10_4569, i_10_4570, i_10_4571, i_10_4580, i_10_4585, o_10_119);
	kernel_10_120 k_10_120(i_10_28, i_10_119, i_10_122, i_10_172, i_10_174, i_10_175, i_10_280, i_10_281, i_10_424, i_10_425, i_10_432, i_10_433, i_10_434, i_10_436, i_10_437, i_10_449, i_10_459, i_10_992, i_10_1044, i_10_1045, i_10_1197, i_10_1233, i_10_1236, i_10_1239, i_10_1305, i_10_1308, i_10_1309, i_10_1310, i_10_1312, i_10_1540, i_10_1580, i_10_1612, i_10_1651, i_10_1652, i_10_1686, i_10_1687, i_10_1688, i_10_1689, i_10_1824, i_10_1946, i_10_1991, i_10_2030, i_10_2179, i_10_2204, i_10_2349, i_10_2350, i_10_2359, i_10_2360, i_10_2362, i_10_2377, i_10_2448, i_10_2457, i_10_2512, i_10_2513, i_10_2628, i_10_2629, i_10_2630, i_10_2633, i_10_2636, i_10_2659, i_10_2660, i_10_2663, i_10_2675, i_10_2723, i_10_2830, i_10_2831, i_10_2832, i_10_2917, i_10_2919, i_10_2983, i_10_3046, i_10_3050, i_10_3087, i_10_3323, i_10_3326, i_10_3350, i_10_3392, i_10_3402, i_10_3403, i_10_3404, i_10_3406, i_10_3551, i_10_3614, i_10_3650, i_10_3782, i_10_3785, i_10_3834, i_10_3836, i_10_3838, i_10_3848, i_10_3853, i_10_3854, i_10_3855, i_10_3856, i_10_3858, i_10_3980, i_10_3988, i_10_4028, i_10_4216, i_10_4266, o_10_120);
	kernel_10_121 k_10_121(i_10_176, i_10_219, i_10_220, i_10_283, i_10_284, i_10_285, i_10_316, i_10_317, i_10_443, i_10_446, i_10_447, i_10_459, i_10_460, i_10_462, i_10_465, i_10_623, i_10_793, i_10_794, i_10_796, i_10_797, i_10_799, i_10_962, i_10_1026, i_10_1032, i_10_1033, i_10_1081, i_10_1084, i_10_1235, i_10_1313, i_10_1546, i_10_1575, i_10_1577, i_10_1620, i_10_1765, i_10_1819, i_10_1820, i_10_1822, i_10_1825, i_10_1826, i_10_1913, i_10_2025, i_10_2026, i_10_2197, i_10_2199, i_10_2200, i_10_2350, i_10_2351, i_10_2352, i_10_2353, i_10_2354, i_10_2362, i_10_2380, i_10_2448, i_10_2450, i_10_2456, i_10_2631, i_10_2633, i_10_2660, i_10_2712, i_10_2722, i_10_2723, i_10_2727, i_10_2728, i_10_2730, i_10_2732, i_10_2827, i_10_2917, i_10_2920, i_10_2921, i_10_2924, i_10_2980, i_10_3075, i_10_3152, i_10_3203, i_10_3281, i_10_3384, i_10_3389, i_10_3391, i_10_3407, i_10_3616, i_10_3617, i_10_3648, i_10_3787, i_10_3839, i_10_3847, i_10_3857, i_10_3858, i_10_3860, i_10_3906, i_10_3907, i_10_4051, i_10_4118, i_10_4275, i_10_4276, i_10_4277, i_10_4284, i_10_4288, i_10_4564, i_10_4569, i_10_4570, o_10_121);
	kernel_10_122 k_10_122(i_10_31, i_10_153, i_10_171, i_10_223, i_10_279, i_10_282, i_10_285, i_10_327, i_10_329, i_10_413, i_10_444, i_10_445, i_10_463, i_10_513, i_10_594, i_10_633, i_10_750, i_10_795, i_10_797, i_10_799, i_10_800, i_10_900, i_10_955, i_10_1236, i_10_1241, i_10_1245, i_10_1306, i_10_1309, i_10_1313, i_10_1435, i_10_1491, i_10_1580, i_10_1654, i_10_1683, i_10_1686, i_10_1791, i_10_1911, i_10_1936, i_10_1951, i_10_1998, i_10_2028, i_10_2183, i_10_2325, i_10_2349, i_10_2376, i_10_2451, i_10_2452, i_10_2455, i_10_2469, i_10_2506, i_10_2632, i_10_2634, i_10_2635, i_10_2636, i_10_2659, i_10_2661, i_10_2673, i_10_2679, i_10_2709, i_10_2712, i_10_2721, i_10_2722, i_10_2725, i_10_2727, i_10_2733, i_10_2781, i_10_2820, i_10_2910, i_10_3070, i_10_3071, i_10_3088, i_10_3279, i_10_3283, i_10_3297, i_10_3451, i_10_3492, i_10_3495, i_10_3585, i_10_3587, i_10_3612, i_10_3619, i_10_3645, i_10_3649, i_10_3724, i_10_3780, i_10_3781, i_10_3783, i_10_3786, i_10_3853, i_10_3870, i_10_3873, i_10_3912, i_10_3945, i_10_4114, i_10_4150, i_10_4188, i_10_4267, i_10_4269, i_10_4270, i_10_4461, o_10_122);
	kernel_10_123 k_10_123(i_10_395, i_10_405, i_10_725, i_10_728, i_10_799, i_10_820, i_10_928, i_10_929, i_10_957, i_10_958, i_10_959, i_10_961, i_10_989, i_10_1027, i_10_1028, i_10_1116, i_10_1119, i_10_1165, i_10_1239, i_10_1305, i_10_1311, i_10_1352, i_10_1359, i_10_1360, i_10_1363, i_10_1364, i_10_1394, i_10_1605, i_10_1606, i_10_1618, i_10_1621, i_10_1698, i_10_1699, i_10_1768, i_10_1786, i_10_1822, i_10_1823, i_10_1954, i_10_2008, i_10_2196, i_10_2243, i_10_2350, i_10_2353, i_10_2446, i_10_2452, i_10_2641, i_10_2700, i_10_2703, i_10_2828, i_10_2831, i_10_2856, i_10_2857, i_10_2868, i_10_2872, i_10_2916, i_10_2917, i_10_2919, i_10_2920, i_10_2921, i_10_2924, i_10_2935, i_10_3037, i_10_3038, i_10_3070, i_10_3225, i_10_3226, i_10_3234, i_10_3271, i_10_3306, i_10_3316, i_10_3317, i_10_3385, i_10_3404, i_10_3451, i_10_3455, i_10_3542, i_10_3543, i_10_3556, i_10_3596, i_10_3720, i_10_3721, i_10_3726, i_10_3727, i_10_3836, i_10_3848, i_10_3860, i_10_3920, i_10_3960, i_10_3961, i_10_3962, i_10_3964, i_10_3965, i_10_4136, i_10_4143, i_10_4217, i_10_4323, i_10_4529, i_10_4568, i_10_4574, i_10_4591, o_10_123);
	kernel_10_124 k_10_124(i_10_146, i_10_176, i_10_275, i_10_282, i_10_316, i_10_388, i_10_389, i_10_406, i_10_424, i_10_425, i_10_433, i_10_434, i_10_441, i_10_443, i_10_463, i_10_464, i_10_505, i_10_506, i_10_751, i_10_797, i_10_992, i_10_1028, i_10_1030, i_10_1037, i_10_1235, i_10_1238, i_10_1305, i_10_1313, i_10_1342, i_10_1343, i_10_1360, i_10_1361, i_10_1445, i_10_1578, i_10_1579, i_10_1580, i_10_1648, i_10_1650, i_10_1651, i_10_1652, i_10_1653, i_10_1688, i_10_1818, i_10_1821, i_10_2183, i_10_2197, i_10_2324, i_10_2353, i_10_2356, i_10_2379, i_10_2456, i_10_2471, i_10_2629, i_10_2630, i_10_2655, i_10_2656, i_10_2659, i_10_2660, i_10_2675, i_10_2711, i_10_2732, i_10_2919, i_10_3043, i_10_3070, i_10_3071, i_10_3072, i_10_3087, i_10_3088, i_10_3089, i_10_3353, i_10_3385, i_10_3388, i_10_3389, i_10_3403, i_10_3404, i_10_3406, i_10_3467, i_10_3523, i_10_3526, i_10_3584, i_10_3586, i_10_3614, i_10_3782, i_10_3784, i_10_3837, i_10_3838, i_10_3850, i_10_3855, i_10_3859, i_10_3875, i_10_3890, i_10_3944, i_10_3991, i_10_3992, i_10_3994, i_10_4052, i_10_4114, i_10_4115, i_10_4288, i_10_4291, o_10_124);
	kernel_10_125 k_10_125(i_10_31, i_10_32, i_10_53, i_10_86, i_10_178, i_10_179, i_10_329, i_10_409, i_10_463, i_10_465, i_10_466, i_10_467, i_10_507, i_10_518, i_10_628, i_10_729, i_10_799, i_10_955, i_10_956, i_10_1005, i_10_1034, i_10_1235, i_10_1238, i_10_1241, i_10_1247, i_10_1305, i_10_1310, i_10_1348, i_10_1444, i_10_1445, i_10_1653, i_10_1717, i_10_1718, i_10_1765, i_10_1818, i_10_1821, i_10_1929, i_10_1948, i_10_2022, i_10_2023, i_10_2181, i_10_2252, i_10_2254, i_10_2326, i_10_2356, i_10_2357, i_10_2410, i_10_2456, i_10_2467, i_10_2469, i_10_2472, i_10_2514, i_10_2515, i_10_2516, i_10_2519, i_10_2570, i_10_2631, i_10_2632, i_10_2678, i_10_2681, i_10_2704, i_10_2705, i_10_2713, i_10_2714, i_10_2717, i_10_2722, i_10_2760, i_10_2784, i_10_2788, i_10_2830, i_10_2831, i_10_2832, i_10_2884, i_10_3072, i_10_3073, i_10_3201, i_10_3281, i_10_3283, i_10_3386, i_10_3390, i_10_3391, i_10_3392, i_10_3444, i_10_3500, i_10_3507, i_10_3586, i_10_3587, i_10_3589, i_10_3590, i_10_3616, i_10_3617, i_10_3648, i_10_3781, i_10_3782, i_10_3844, i_10_3845, i_10_3858, i_10_4115, i_10_4129, i_10_4568, o_10_125);
	kernel_10_126 k_10_126(i_10_57, i_10_171, i_10_184, i_10_223, i_10_247, i_10_271, i_10_327, i_10_390, i_10_424, i_10_436, i_10_442, i_10_443, i_10_445, i_10_463, i_10_464, i_10_589, i_10_717, i_10_993, i_10_1035, i_10_1041, i_10_1057, i_10_1111, i_10_1207, i_10_1210, i_10_1246, i_10_1264, i_10_1381, i_10_1399, i_10_1400, i_10_1453, i_10_1541, i_10_1614, i_10_1632, i_10_1633, i_10_1650, i_10_1655, i_10_1688, i_10_1692, i_10_1764, i_10_1765, i_10_1766, i_10_1794, i_10_1820, i_10_1893, i_10_1938, i_10_1988, i_10_2031, i_10_2032, i_10_2068, i_10_2208, i_10_2244, i_10_2259, i_10_2308, i_10_2309, i_10_2311, i_10_2353, i_10_2387, i_10_2388, i_10_2452, i_10_2523, i_10_2559, i_10_2658, i_10_2662, i_10_2676, i_10_2704, i_10_2820, i_10_3010, i_10_3046, i_10_3073, i_10_3117, i_10_3209, i_10_3277, i_10_3327, i_10_3451, i_10_3466, i_10_3494, i_10_3497, i_10_3526, i_10_3540, i_10_3570, i_10_3577, i_10_3578, i_10_3616, i_10_3639, i_10_3688, i_10_3725, i_10_3780, i_10_3787, i_10_3838, i_10_3855, i_10_3942, i_10_3946, i_10_3981, i_10_4174, i_10_4192, i_10_4193, i_10_4263, i_10_4282, i_10_4567, i_10_4574, o_10_126);
	kernel_10_127 k_10_127(i_10_145, i_10_146, i_10_172, i_10_173, i_10_176, i_10_217, i_10_222, i_10_224, i_10_262, i_10_284, i_10_432, i_10_442, i_10_443, i_10_444, i_10_445, i_10_446, i_10_455, i_10_461, i_10_514, i_10_515, i_10_793, i_10_794, i_10_796, i_10_797, i_10_965, i_10_967, i_10_968, i_10_1085, i_10_1242, i_10_1305, i_10_1360, i_10_1361, i_10_1364, i_10_1575, i_10_1576, i_10_1577, i_10_1631, i_10_1649, i_10_1651, i_10_1652, i_10_1688, i_10_1819, i_10_1820, i_10_1821, i_10_1822, i_10_1823, i_10_1824, i_10_1945, i_10_1999, i_10_2243, i_10_2350, i_10_2355, i_10_2379, i_10_2380, i_10_2448, i_10_2453, i_10_2458, i_10_2462, i_10_2503, i_10_2504, i_10_2629, i_10_2674, i_10_2675, i_10_2681, i_10_2701, i_10_2718, i_10_2719, i_10_2726, i_10_2734, i_10_2827, i_10_2828, i_10_2830, i_10_2908, i_10_3046, i_10_3232, i_10_3233, i_10_3387, i_10_3389, i_10_3494, i_10_3520, i_10_3524, i_10_3584, i_10_3587, i_10_3610, i_10_3613, i_10_3784, i_10_3809, i_10_3839, i_10_3846, i_10_3853, i_10_3858, i_10_3890, i_10_3913, i_10_3943, i_10_4130, i_10_4268, i_10_4287, i_10_4288, i_10_4291, i_10_4565, o_10_127);
	kernel_10_128 k_10_128(i_10_244, i_10_281, i_10_282, i_10_284, i_10_288, i_10_289, i_10_315, i_10_319, i_10_412, i_10_435, i_10_449, i_10_461, i_10_462, i_10_464, i_10_467, i_10_500, i_10_735, i_10_792, i_10_797, i_10_1118, i_10_1234, i_10_1235, i_10_1238, i_10_1243, i_10_1244, i_10_1245, i_10_1273, i_10_1307, i_10_1361, i_10_1451, i_10_1583, i_10_1651, i_10_1652, i_10_1687, i_10_1688, i_10_1818, i_10_1819, i_10_1820, i_10_1822, i_10_1910, i_10_1945, i_10_1946, i_10_1949, i_10_1951, i_10_1989, i_10_1990, i_10_2178, i_10_2333, i_10_2352, i_10_2353, i_10_2356, i_10_2364, i_10_2376, i_10_2407, i_10_2408, i_10_2441, i_10_2454, i_10_2455, i_10_2459, i_10_2470, i_10_2673, i_10_2679, i_10_2700, i_10_2704, i_10_2709, i_10_2882, i_10_2918, i_10_2921, i_10_2924, i_10_3267, i_10_3268, i_10_3269, i_10_3276, i_10_3277, i_10_3278, i_10_3280, i_10_3281, i_10_3384, i_10_3386, i_10_3406, i_10_3497, i_10_3586, i_10_3615, i_10_3645, i_10_3682, i_10_3728, i_10_3784, i_10_3839, i_10_3846, i_10_3858, i_10_3859, i_10_3894, i_10_3895, i_10_3984, i_10_4054, i_10_4116, i_10_4117, i_10_4119, i_10_4457, i_10_4568, o_10_128);
	kernel_10_129 k_10_129(i_10_51, i_10_52, i_10_153, i_10_156, i_10_181, i_10_237, i_10_251, i_10_283, i_10_293, i_10_327, i_10_354, i_10_355, i_10_357, i_10_589, i_10_633, i_10_636, i_10_687, i_10_688, i_10_732, i_10_828, i_10_930, i_10_993, i_10_1135, i_10_1161, i_10_1209, i_10_1234, i_10_1290, i_10_1306, i_10_1380, i_10_1530, i_10_1531, i_10_1533, i_10_1534, i_10_1543, i_10_1560, i_10_1561, i_10_1632, i_10_1651, i_10_1686, i_10_1791, i_10_1800, i_10_1801, i_10_1848, i_10_1912, i_10_1918, i_10_2163, i_10_2200, i_10_2253, i_10_2256, i_10_2442, i_10_2450, i_10_2529, i_10_2604, i_10_2632, i_10_2674, i_10_2713, i_10_2715, i_10_2716, i_10_2724, i_10_2775, i_10_2832, i_10_2979, i_10_2982, i_10_3096, i_10_3099, i_10_3196, i_10_3198, i_10_3199, i_10_3280, i_10_3282, i_10_3289, i_10_3291, i_10_3315, i_10_3325, i_10_3387, i_10_3388, i_10_3390, i_10_3391, i_10_3465, i_10_3564, i_10_3577, i_10_3609, i_10_3610, i_10_3645, i_10_3646, i_10_3648, i_10_3702, i_10_3703, i_10_3774, i_10_3780, i_10_3783, i_10_3786, i_10_3857, i_10_3870, i_10_3873, i_10_3996, i_10_4131, i_10_4226, i_10_4461, i_10_4582, o_10_129);
	kernel_10_130 k_10_130(i_10_51, i_10_293, i_10_391, i_10_427, i_10_428, i_10_433, i_10_447, i_10_449, i_10_465, i_10_613, i_10_714, i_10_750, i_10_893, i_10_984, i_10_993, i_10_1012, i_10_1029, i_10_1034, i_10_1170, i_10_1171, i_10_1239, i_10_1242, i_10_1244, i_10_1245, i_10_1246, i_10_1247, i_10_1248, i_10_1249, i_10_1445, i_10_1447, i_10_1542, i_10_1632, i_10_1650, i_10_1653, i_10_1654, i_10_1756, i_10_1758, i_10_1759, i_10_1819, i_10_1823, i_10_2012, i_10_2181, i_10_2203, i_10_2207, i_10_2225, i_10_2307, i_10_2362, i_10_2454, i_10_2470, i_10_2471, i_10_2473, i_10_2532, i_10_2628, i_10_2655, i_10_2660, i_10_2686, i_10_2916, i_10_3033, i_10_3034, i_10_3037, i_10_3041, i_10_3166, i_10_3169, i_10_3172, i_10_3307, i_10_3334, i_10_3386, i_10_3429, i_10_3469, i_10_3586, i_10_3590, i_10_3617, i_10_3684, i_10_3685, i_10_3687, i_10_3688, i_10_3717, i_10_3729, i_10_3780, i_10_3784, i_10_3786, i_10_3829, i_10_3844, i_10_4008, i_10_4011, i_10_4066, i_10_4117, i_10_4118, i_10_4174, i_10_4175, i_10_4188, i_10_4219, i_10_4260, i_10_4261, i_10_4269, i_10_4276, i_10_4287, i_10_4477, i_10_4569, i_10_4597, o_10_130);
	kernel_10_131 k_10_131(i_10_48, i_10_118, i_10_136, i_10_171, i_10_182, i_10_246, i_10_282, i_10_283, i_10_285, i_10_286, i_10_291, i_10_292, i_10_293, i_10_315, i_10_330, i_10_390, i_10_391, i_10_407, i_10_409, i_10_410, i_10_448, i_10_625, i_10_634, i_10_689, i_10_792, i_10_826, i_10_957, i_10_963, i_10_967, i_10_993, i_10_1051, i_10_1052, i_10_1163, i_10_1266, i_10_1267, i_10_1302, i_10_1306, i_10_1435, i_10_1444, i_10_1488, i_10_1579, i_10_1581, i_10_1618, i_10_1649, i_10_1653, i_10_1683, i_10_1684, i_10_1800, i_10_2004, i_10_2025, i_10_2082, i_10_2202, i_10_2203, i_10_2353, i_10_2355, i_10_2361, i_10_2377, i_10_2455, i_10_2475, i_10_2541, i_10_2566, i_10_2572, i_10_2605, i_10_2607, i_10_2608, i_10_2611, i_10_2634, i_10_2677, i_10_2679, i_10_2709, i_10_2712, i_10_2718, i_10_2719, i_10_2725, i_10_2734, i_10_2782, i_10_2985, i_10_3198, i_10_3199, i_10_3235, i_10_3282, i_10_3288, i_10_3387, i_10_3388, i_10_3433, i_10_3471, i_10_3585, i_10_3609, i_10_3647, i_10_3721, i_10_3859, i_10_3860, i_10_4030, i_10_4113, i_10_4116, i_10_4275, i_10_4276, i_10_4280, i_10_4459, i_10_4566, o_10_131);
	kernel_10_132 k_10_132(i_10_222, i_10_223, i_10_224, i_10_271, i_10_327, i_10_328, i_10_332, i_10_407, i_10_430, i_10_433, i_10_435, i_10_438, i_10_439, i_10_507, i_10_699, i_10_955, i_10_996, i_10_997, i_10_1001, i_10_1005, i_10_1138, i_10_1237, i_10_1238, i_10_1246, i_10_1247, i_10_1249, i_10_1264, i_10_1307, i_10_1309, i_10_1310, i_10_1312, i_10_1438, i_10_1554, i_10_1654, i_10_1688, i_10_1818, i_10_2020, i_10_2158, i_10_2407, i_10_2508, i_10_2509, i_10_2629, i_10_2630, i_10_2634, i_10_2635, i_10_2657, i_10_2661, i_10_2679, i_10_2680, i_10_2681, i_10_2720, i_10_2724, i_10_2783, i_10_2820, i_10_2823, i_10_2826, i_10_2827, i_10_2828, i_10_2831, i_10_2881, i_10_2882, i_10_2980, i_10_2982, i_10_2985, i_10_3041, i_10_3072, i_10_3199, i_10_3271, i_10_3328, i_10_3387, i_10_3388, i_10_3390, i_10_3391, i_10_3408, i_10_3496, i_10_3614, i_10_3646, i_10_3648, i_10_3652, i_10_3682, i_10_3729, i_10_3780, i_10_3781, i_10_3846, i_10_3848, i_10_3850, i_10_3852, i_10_3853, i_10_3855, i_10_3859, i_10_3981, i_10_3982, i_10_3984, i_10_3985, i_10_3986, i_10_4056, i_10_4129, i_10_4238, i_10_4288, i_10_4289, o_10_132);
	kernel_10_133 k_10_133(i_10_176, i_10_178, i_10_247, i_10_283, i_10_284, i_10_286, i_10_322, i_10_323, i_10_327, i_10_407, i_10_441, i_10_447, i_10_461, i_10_504, i_10_509, i_10_511, i_10_796, i_10_957, i_10_1039, i_10_1043, i_10_1235, i_10_1237, i_10_1246, i_10_1345, i_10_1346, i_10_1442, i_10_1578, i_10_1649, i_10_1655, i_10_1683, i_10_1727, i_10_1768, i_10_1823, i_10_1910, i_10_1912, i_10_1913, i_10_1951, i_10_2000, i_10_2005, i_10_2028, i_10_2186, i_10_2361, i_10_2364, i_10_2365, i_10_2450, i_10_2452, i_10_2453, i_10_2569, i_10_2632, i_10_2710, i_10_2723, i_10_2735, i_10_2884, i_10_2916, i_10_3151, i_10_3195, i_10_3268, i_10_3271, i_10_3274, i_10_3277, i_10_3278, i_10_3279, i_10_3280, i_10_3281, i_10_3283, i_10_3322, i_10_3384, i_10_3392, i_10_3402, i_10_3407, i_10_3520, i_10_3521, i_10_3537, i_10_3542, i_10_3613, i_10_3614, i_10_3647, i_10_3648, i_10_3649, i_10_3784, i_10_3785, i_10_3786, i_10_3787, i_10_3837, i_10_3846, i_10_3858, i_10_3859, i_10_3894, i_10_3895, i_10_3896, i_10_3912, i_10_3913, i_10_3914, i_10_4126, i_10_4281, i_10_4283, i_10_4288, i_10_4290, i_10_4292, i_10_4565, o_10_133);
	kernel_10_134 k_10_134(i_10_31, i_10_37, i_10_67, i_10_117, i_10_125, i_10_259, i_10_264, i_10_266, i_10_284, i_10_317, i_10_394, i_10_405, i_10_406, i_10_688, i_10_715, i_10_756, i_10_865, i_10_866, i_10_952, i_10_991, i_10_993, i_10_1054, i_10_1084, i_10_1135, i_10_1136, i_10_1267, i_10_1269, i_10_1281, i_10_1378, i_10_1438, i_10_1439, i_10_1554, i_10_1577, i_10_1579, i_10_1582, i_10_1583, i_10_1687, i_10_1803, i_10_1810, i_10_1811, i_10_1818, i_10_1846, i_10_1909, i_10_1910, i_10_1912, i_10_1986, i_10_2017, i_10_2018, i_10_2185, i_10_2263, i_10_2351, i_10_2353, i_10_2383, i_10_2404, i_10_2473, i_10_2474, i_10_2487, i_10_2519, i_10_2536, i_10_2563, i_10_2578, i_10_2586, i_10_2596, i_10_2607, i_10_2608, i_10_2702, i_10_2722, i_10_2725, i_10_2726, i_10_2734, i_10_2735, i_10_2787, i_10_2809, i_10_2881, i_10_2884, i_10_2885, i_10_2955, i_10_2983, i_10_2993, i_10_3043, i_10_3048, i_10_3282, i_10_3283, i_10_3284, i_10_3356, i_10_3394, i_10_3395, i_10_3562, i_10_3609, i_10_3841, i_10_3985, i_10_4031, i_10_4063, i_10_4292, i_10_4377, i_10_4378, i_10_4397, i_10_4434, i_10_4588, i_10_4589, o_10_134);
	kernel_10_135 k_10_135(i_10_52, i_10_171, i_10_173, i_10_176, i_10_178, i_10_179, i_10_221, i_10_222, i_10_224, i_10_279, i_10_296, i_10_328, i_10_329, i_10_390, i_10_391, i_10_394, i_10_439, i_10_446, i_10_449, i_10_515, i_10_516, i_10_517, i_10_518, i_10_521, i_10_596, i_10_957, i_10_959, i_10_998, i_10_1138, i_10_1160, i_10_1265, i_10_1268, i_10_1445, i_10_1636, i_10_1651, i_10_1652, i_10_1686, i_10_1687, i_10_1817, i_10_1819, i_10_1821, i_10_1877, i_10_2026, i_10_2179, i_10_2201, i_10_2255, i_10_2330, i_10_2353, i_10_2354, i_10_2364, i_10_2515, i_10_2631, i_10_2636, i_10_2675, i_10_2678, i_10_2681, i_10_2705, i_10_2706, i_10_2725, i_10_2821, i_10_2825, i_10_2829, i_10_2920, i_10_2980, i_10_2984, i_10_3035, i_10_3036, i_10_3038, i_10_3199, i_10_3275, i_10_3281, i_10_3290, i_10_3293, i_10_3494, i_10_3497, i_10_3523, i_10_3524, i_10_3527, i_10_3583, i_10_3616, i_10_3781, i_10_3782, i_10_3784, i_10_3785, i_10_3787, i_10_3788, i_10_3800, i_10_3910, i_10_3911, i_10_3913, i_10_3914, i_10_3950, i_10_4120, i_10_4121, i_10_4127, i_10_4130, i_10_4238, i_10_4268, i_10_4280, i_10_4463, o_10_135);
	kernel_10_136 k_10_136(i_10_174, i_10_219, i_10_286, i_10_318, i_10_328, i_10_424, i_10_444, i_10_446, i_10_793, i_10_799, i_10_896, i_10_955, i_10_1032, i_10_1033, i_10_1308, i_10_1437, i_10_1542, i_10_1583, i_10_1650, i_10_1688, i_10_1765, i_10_1821, i_10_1822, i_10_1912, i_10_1913, i_10_1995, i_10_2178, i_10_2179, i_10_2180, i_10_2305, i_10_2306, i_10_2326, i_10_2350, i_10_2351, i_10_2352, i_10_2353, i_10_2361, i_10_2382, i_10_2404, i_10_2452, i_10_2502, i_10_2571, i_10_2633, i_10_2636, i_10_2673, i_10_2705, i_10_2714, i_10_2727, i_10_2728, i_10_2729, i_10_2733, i_10_2734, i_10_2735, i_10_2826, i_10_2827, i_10_2830, i_10_2832, i_10_2922, i_10_3070, i_10_3153, i_10_3155, i_10_3162, i_10_3196, i_10_3199, i_10_3202, i_10_3268, i_10_3270, i_10_3277, i_10_3326, i_10_3385, i_10_3388, i_10_3389, i_10_3390, i_10_3470, i_10_3612, i_10_3613, i_10_3649, i_10_3652, i_10_3683, i_10_3732, i_10_3780, i_10_3782, i_10_3834, i_10_3857, i_10_3907, i_10_3982, i_10_4050, i_10_4051, i_10_4119, i_10_4128, i_10_4129, i_10_4130, i_10_4168, i_10_4169, i_10_4219, i_10_4270, i_10_4281, i_10_4288, i_10_4566, i_10_4569, o_10_136);
	kernel_10_137 k_10_137(i_10_37, i_10_148, i_10_222, i_10_223, i_10_325, i_10_352, i_10_445, i_10_459, i_10_462, i_10_520, i_10_586, i_10_587, i_10_594, i_10_729, i_10_730, i_10_749, i_10_795, i_10_834, i_10_846, i_10_892, i_10_955, i_10_956, i_10_1026, i_10_1027, i_10_1039, i_10_1042, i_10_1117, i_10_1118, i_10_1161, i_10_1185, i_10_1333, i_10_1342, i_10_1344, i_10_1353, i_10_1362, i_10_1371, i_10_1574, i_10_1579, i_10_1650, i_10_1767, i_10_1801, i_10_1802, i_10_1810, i_10_1818, i_10_1819, i_10_1821, i_10_1875, i_10_1956, i_10_2200, i_10_2338, i_10_2351, i_10_2405, i_10_2451, i_10_2462, i_10_2512, i_10_2538, i_10_2543, i_10_2556, i_10_2568, i_10_2679, i_10_2704, i_10_2730, i_10_2754, i_10_2829, i_10_2830, i_10_2882, i_10_2922, i_10_2955, i_10_2992, i_10_3047, i_10_3049, i_10_3228, i_10_3267, i_10_3272, i_10_3384, i_10_3432, i_10_3433, i_10_3481, i_10_3519, i_10_3520, i_10_3522, i_10_3583, i_10_3584, i_10_3609, i_10_3614, i_10_3684, i_10_3723, i_10_3725, i_10_3857, i_10_4005, i_10_4006, i_10_4007, i_10_4118, i_10_4236, i_10_4285, i_10_4287, i_10_4324, i_10_4425, i_10_4488, i_10_4566, o_10_137);
	kernel_10_138 k_10_138(i_10_34, i_10_171, i_10_178, i_10_250, i_10_283, i_10_318, i_10_392, i_10_409, i_10_410, i_10_441, i_10_448, i_10_449, i_10_514, i_10_751, i_10_963, i_10_1034, i_10_1080, i_10_1242, i_10_1246, i_10_1248, i_10_1249, i_10_1308, i_10_1547, i_10_1575, i_10_1578, i_10_1651, i_10_1760, i_10_1823, i_10_1915, i_10_2006, i_10_2022, i_10_2359, i_10_2411, i_10_2470, i_10_2473, i_10_2474, i_10_2537, i_10_2654, i_10_2659, i_10_2681, i_10_2710, i_10_2728, i_10_2729, i_10_2730, i_10_2833, i_10_2869, i_10_2920, i_10_2921, i_10_3034, i_10_3036, i_10_3037, i_10_3038, i_10_3039, i_10_3162, i_10_3199, i_10_3200, i_10_3202, i_10_3279, i_10_3281, i_10_3284, i_10_3338, i_10_3384, i_10_3386, i_10_3389, i_10_3403, i_10_3408, i_10_3433, i_10_3434, i_10_3466, i_10_3496, i_10_3522, i_10_3526, i_10_3612, i_10_3614, i_10_3648, i_10_3727, i_10_3733, i_10_3782, i_10_3783, i_10_3784, i_10_3785, i_10_3787, i_10_3835, i_10_3836, i_10_3844, i_10_3846, i_10_3848, i_10_3855, i_10_3856, i_10_3857, i_10_3860, i_10_3983, i_10_4120, i_10_4121, i_10_4220, i_10_4286, i_10_4289, i_10_4567, i_10_4568, i_10_4569, o_10_138);
	kernel_10_139 k_10_139(i_10_174, i_10_223, i_10_249, i_10_264, i_10_268, i_10_282, i_10_285, i_10_390, i_10_391, i_10_406, i_10_408, i_10_433, i_10_436, i_10_437, i_10_439, i_10_440, i_10_443, i_10_447, i_10_449, i_10_509, i_10_931, i_10_957, i_10_991, i_10_994, i_10_997, i_10_998, i_10_1002, i_10_1307, i_10_1308, i_10_1309, i_10_1349, i_10_1383, i_10_1435, i_10_1650, i_10_1654, i_10_1713, i_10_1823, i_10_1909, i_10_1910, i_10_1911, i_10_1912, i_10_1913, i_10_1915, i_10_2094, i_10_2184, i_10_2185, i_10_2201, i_10_2350, i_10_2361, i_10_2364, i_10_2451, i_10_2452, i_10_2464, i_10_2469, i_10_2508, i_10_2509, i_10_2604, i_10_2616, i_10_2617, i_10_2635, i_10_2680, i_10_2701, i_10_2705, i_10_2717, i_10_2731, i_10_2734, i_10_2817, i_10_2820, i_10_2821, i_10_2832, i_10_2885, i_10_2886, i_10_2887, i_10_2917, i_10_2919, i_10_3014, i_10_3195, i_10_3275, i_10_3281, i_10_3471, i_10_3472, i_10_3497, i_10_3706, i_10_3787, i_10_3837, i_10_3838, i_10_3850, i_10_3854, i_10_3859, i_10_3982, i_10_3984, i_10_3985, i_10_3986, i_10_4117, i_10_4118, i_10_4119, i_10_4236, i_10_4238, i_10_4533, i_10_4568, o_10_139);
	kernel_10_140 k_10_140(i_10_29, i_10_117, i_10_124, i_10_154, i_10_181, i_10_182, i_10_183, i_10_219, i_10_253, i_10_257, i_10_261, i_10_264, i_10_318, i_10_410, i_10_427, i_10_460, i_10_461, i_10_463, i_10_464, i_10_904, i_10_946, i_10_949, i_10_958, i_10_959, i_10_1219, i_10_1246, i_10_1267, i_10_1297, i_10_1305, i_10_1306, i_10_1311, i_10_1313, i_10_1359, i_10_1361, i_10_1363, i_10_1364, i_10_1539, i_10_1540, i_10_1553, i_10_1683, i_10_1687, i_10_1940, i_10_1942, i_10_1980, i_10_2001, i_10_2202, i_10_2235, i_10_2304, i_10_2349, i_10_2350, i_10_2362, i_10_2376, i_10_2382, i_10_2383, i_10_2411, i_10_2448, i_10_2452, i_10_2453, i_10_2468, i_10_2514, i_10_2529, i_10_2530, i_10_2614, i_10_2615, i_10_2631, i_10_2636, i_10_2657, i_10_2738, i_10_2785, i_10_2832, i_10_2881, i_10_2920, i_10_2921, i_10_3073, i_10_3197, i_10_3278, i_10_3315, i_10_3408, i_10_3469, i_10_3609, i_10_3610, i_10_3611, i_10_3617, i_10_3647, i_10_3834, i_10_3838, i_10_3853, i_10_4050, i_10_4114, i_10_4117, i_10_4125, i_10_4129, i_10_4186, i_10_4217, i_10_4288, i_10_4289, i_10_4291, i_10_4563, i_10_4564, i_10_4567, o_10_140);
	kernel_10_141 k_10_141(i_10_136, i_10_172, i_10_183, i_10_253, i_10_318, i_10_321, i_10_328, i_10_409, i_10_430, i_10_436, i_10_459, i_10_460, i_10_585, i_10_586, i_10_795, i_10_919, i_10_996, i_10_997, i_10_1039, i_10_1041, i_10_1042, i_10_1086, i_10_1087, i_10_1163, i_10_1238, i_10_1240, i_10_1241, i_10_1307, i_10_1308, i_10_1345, i_10_1361, i_10_1439, i_10_1551, i_10_1615, i_10_1630, i_10_1633, i_10_1651, i_10_1690, i_10_1691, i_10_1719, i_10_1729, i_10_1818, i_10_1873, i_10_1881, i_10_1911, i_10_2000, i_10_2233, i_10_2354, i_10_2407, i_10_2468, i_10_2473, i_10_2509, i_10_2566, i_10_2606, i_10_2718, i_10_2720, i_10_2787, i_10_2826, i_10_2827, i_10_2830, i_10_2833, i_10_2834, i_10_2908, i_10_2911, i_10_2920, i_10_3038, i_10_3070, i_10_3071, i_10_3116, i_10_3279, i_10_3406, i_10_3447, i_10_3587, i_10_3588, i_10_3589, i_10_3613, i_10_3615, i_10_3616, i_10_3622, i_10_3650, i_10_3774, i_10_3780, i_10_3782, i_10_3798, i_10_3840, i_10_3860, i_10_3891, i_10_3894, i_10_3895, i_10_4096, i_10_4115, i_10_4131, i_10_4230, i_10_4261, i_10_4312, i_10_4460, i_10_4519, i_10_4529, i_10_4567, i_10_4585, o_10_141);
	kernel_10_142 k_10_142(i_10_171, i_10_175, i_10_279, i_10_280, i_10_281, i_10_282, i_10_283, i_10_284, i_10_286, i_10_429, i_10_445, i_10_460, i_10_506, i_10_517, i_10_518, i_10_519, i_10_794, i_10_799, i_10_967, i_10_968, i_10_1032, i_10_1037, i_10_1238, i_10_1349, i_10_1491, i_10_1550, i_10_1580, i_10_1650, i_10_1681, i_10_1686, i_10_1687, i_10_1688, i_10_1821, i_10_1822, i_10_1823, i_10_2001, i_10_2004, i_10_2152, i_10_2304, i_10_2305, i_10_2306, i_10_2351, i_10_2354, i_10_2364, i_10_2452, i_10_2467, i_10_2571, i_10_2630, i_10_2632, i_10_2655, i_10_2658, i_10_2659, i_10_2701, i_10_2715, i_10_2717, i_10_2721, i_10_2831, i_10_2883, i_10_2884, i_10_2920, i_10_2922, i_10_3043, i_10_3070, i_10_3071, i_10_3151, i_10_3165, i_10_3267, i_10_3270, i_10_3271, i_10_3280, i_10_3388, i_10_3389, i_10_3390, i_10_3404, i_10_3406, i_10_3408, i_10_3582, i_10_3612, i_10_3614, i_10_3784, i_10_3786, i_10_3787, i_10_3839, i_10_3841, i_10_3852, i_10_3853, i_10_3857, i_10_3889, i_10_3890, i_10_3912, i_10_3913, i_10_3914, i_10_4117, i_10_4130, i_10_4287, i_10_4288, i_10_4289, i_10_4290, i_10_4563, i_10_4570, o_10_142);
	kernel_10_143 k_10_143(i_10_173, i_10_176, i_10_245, i_10_272, i_10_275, i_10_283, i_10_316, i_10_317, i_10_319, i_10_320, i_10_391, i_10_413, i_10_434, i_10_445, i_10_461, i_10_464, i_10_716, i_10_749, i_10_752, i_10_794, i_10_797, i_10_892, i_10_893, i_10_992, i_10_995, i_10_1084, i_10_1154, i_10_1305, i_10_1310, i_10_1313, i_10_1342, i_10_1343, i_10_1346, i_10_1360, i_10_1361, i_10_1442, i_10_1622, i_10_1648, i_10_1652, i_10_1684, i_10_1685, i_10_1712, i_10_1823, i_10_1874, i_10_1916, i_10_1990, i_10_2017, i_10_2018, i_10_2198, i_10_2359, i_10_2381, i_10_2432, i_10_2468, i_10_2469, i_10_2470, i_10_2628, i_10_2630, i_10_2631, i_10_2632, i_10_2633, i_10_2636, i_10_2659, i_10_2674, i_10_2702, i_10_2711, i_10_2722, i_10_2782, i_10_2783, i_10_2827, i_10_2828, i_10_3044, i_10_3070, i_10_3071, i_10_3272, i_10_3278, i_10_3326, i_10_3328, i_10_3329, i_10_3392, i_10_3467, i_10_3523, i_10_3647, i_10_3837, i_10_3847, i_10_3848, i_10_3853, i_10_3854, i_10_3991, i_10_4114, i_10_4116, i_10_4117, i_10_4121, i_10_4127, i_10_4169, i_10_4276, i_10_4277, i_10_4286, i_10_4292, i_10_4568, i_10_4571, o_10_143);
	kernel_10_144 k_10_144(i_10_145, i_10_177, i_10_246, i_10_252, i_10_282, i_10_315, i_10_316, i_10_322, i_10_327, i_10_443, i_10_444, i_10_498, i_10_501, i_10_504, i_10_505, i_10_508, i_10_712, i_10_1059, i_10_1084, i_10_1236, i_10_1239, i_10_1241, i_10_1299, i_10_1302, i_10_1312, i_10_1363, i_10_1434, i_10_1444, i_10_1542, i_10_1576, i_10_1578, i_10_1618, i_10_1623, i_10_1686, i_10_1688, i_10_1689, i_10_1731, i_10_1734, i_10_1803, i_10_1820, i_10_1822, i_10_1823, i_10_1978, i_10_2028, i_10_2031, i_10_2202, i_10_2376, i_10_2451, i_10_2455, i_10_2466, i_10_2469, i_10_2470, i_10_2472, i_10_2568, i_10_2700, i_10_2715, i_10_2721, i_10_2725, i_10_2733, i_10_2826, i_10_2832, i_10_2964, i_10_2967, i_10_3196, i_10_3268, i_10_3277, i_10_3279, i_10_3281, i_10_3282, i_10_3283, i_10_3315, i_10_3318, i_10_3325, i_10_3327, i_10_3385, i_10_3501, i_10_3504, i_10_3543, i_10_3544, i_10_3582, i_10_3585, i_10_3588, i_10_3646, i_10_3651, i_10_3781, i_10_3795, i_10_3840, i_10_3909, i_10_4030, i_10_4114, i_10_4119, i_10_4266, i_10_4269, i_10_4272, i_10_4281, i_10_4290, i_10_4548, i_10_4567, i_10_4570, i_10_4585, o_10_144);
	kernel_10_145 k_10_145(i_10_21, i_10_22, i_10_58, i_10_89, i_10_181, i_10_213, i_10_277, i_10_280, i_10_388, i_10_445, i_10_500, i_10_507, i_10_584, i_10_595, i_10_597, i_10_598, i_10_659, i_10_679, i_10_729, i_10_967, i_10_1011, i_10_1187, i_10_1201, i_10_1326, i_10_1327, i_10_1345, i_10_1366, i_10_1444, i_10_1480, i_10_1488, i_10_1526, i_10_1536, i_10_1543, i_10_1548, i_10_1614, i_10_1624, i_10_1651, i_10_1652, i_10_1713, i_10_1750, i_10_1761, i_10_1789, i_10_1826, i_10_1875, i_10_1919, i_10_1930, i_10_2001, i_10_2152, i_10_2226, i_10_2227, i_10_2272, i_10_2507, i_10_2601, i_10_2604, i_10_2653, i_10_2667, i_10_2668, i_10_2732, i_10_2767, i_10_2803, i_10_2877, i_10_2879, i_10_2953, i_10_2963, i_10_3028, i_10_3029, i_10_3040, i_10_3043, i_10_3057, i_10_3135, i_10_3189, i_10_3190, i_10_3191, i_10_3201, i_10_3224, i_10_3297, i_10_3402, i_10_3403, i_10_3544, i_10_3604, i_10_3610, i_10_3616, i_10_3723, i_10_3724, i_10_3729, i_10_3838, i_10_3863, i_10_3922, i_10_3975, i_10_4068, i_10_4069, i_10_4182, i_10_4218, i_10_4407, i_10_4446, i_10_4447, i_10_4455, i_10_4459, i_10_4516, i_10_4517, o_10_145);
	kernel_10_146 k_10_146(i_10_43, i_10_176, i_10_178, i_10_283, i_10_284, i_10_287, i_10_293, i_10_315, i_10_316, i_10_317, i_10_390, i_10_426, i_10_429, i_10_435, i_10_436, i_10_445, i_10_499, i_10_588, i_10_589, i_10_693, i_10_694, i_10_928, i_10_990, i_10_991, i_10_1033, i_10_1233, i_10_1234, i_10_1235, i_10_1238, i_10_1309, i_10_1310, i_10_1445, i_10_1541, i_10_1581, i_10_1685, i_10_1688, i_10_1764, i_10_1821, i_10_1823, i_10_1909, i_10_1910, i_10_2353, i_10_2449, i_10_2451, i_10_2452, i_10_2460, i_10_2463, i_10_2467, i_10_2468, i_10_2514, i_10_2634, i_10_2733, i_10_2817, i_10_2831, i_10_2880, i_10_2881, i_10_2883, i_10_2884, i_10_2919, i_10_2920, i_10_2921, i_10_2979, i_10_2980, i_10_3090, i_10_3091, i_10_3159, i_10_3169, i_10_3199, i_10_3200, i_10_3356, i_10_3388, i_10_3445, i_10_3446, i_10_3519, i_10_3520, i_10_3522, i_10_3613, i_10_3614, i_10_3699, i_10_3703, i_10_3826, i_10_3850, i_10_3853, i_10_3889, i_10_3890, i_10_3898, i_10_3899, i_10_3905, i_10_3906, i_10_3984, i_10_4026, i_10_4028, i_10_4031, i_10_4052, i_10_4097, i_10_4216, i_10_4531, i_10_4591, i_10_4592, i_10_4594, o_10_146);
	kernel_10_147 k_10_147(i_10_176, i_10_218, i_10_221, i_10_270, i_10_275, i_10_285, i_10_319, i_10_435, i_10_442, i_10_464, i_10_506, i_10_507, i_10_955, i_10_956, i_10_959, i_10_961, i_10_1027, i_10_1028, i_10_1030, i_10_1031, i_10_1034, i_10_1086, i_10_1087, i_10_1134, i_10_1141, i_10_1237, i_10_1246, i_10_1307, i_10_1308, i_10_1540, i_10_1541, i_10_1543, i_10_1552, i_10_1553, i_10_1580, i_10_1649, i_10_1691, i_10_1820, i_10_1826, i_10_1994, i_10_2201, i_10_2204, i_10_2358, i_10_2363, i_10_2365, i_10_2461, i_10_2464, i_10_2466, i_10_2470, i_10_2628, i_10_2663, i_10_2674, i_10_2678, i_10_2700, i_10_2701, i_10_2722, i_10_2723, i_10_2833, i_10_2834, i_10_2885, i_10_2924, i_10_3196, i_10_3197, i_10_3199, i_10_3202, i_10_3203, i_10_3268, i_10_3280, i_10_3323, i_10_3392, i_10_3403, i_10_3466, i_10_3469, i_10_3470, i_10_3522, i_10_3583, i_10_3586, i_10_3587, i_10_3589, i_10_3731, i_10_3781, i_10_3782, i_10_3784, i_10_3785, i_10_3786, i_10_3787, i_10_3788, i_10_3844, i_10_3849, i_10_3854, i_10_3856, i_10_3857, i_10_3859, i_10_3860, i_10_3979, i_10_3980, i_10_3982, i_10_4121, i_10_4291, i_10_4567, o_10_147);
	kernel_10_148 k_10_148(i_10_178, i_10_283, i_10_327, i_10_406, i_10_429, i_10_446, i_10_461, i_10_463, i_10_464, i_10_465, i_10_466, i_10_467, i_10_498, i_10_795, i_10_796, i_10_994, i_10_1123, i_10_1236, i_10_1237, i_10_1238, i_10_1240, i_10_1241, i_10_1491, i_10_1575, i_10_1650, i_10_1651, i_10_1683, i_10_1685, i_10_1689, i_10_1690, i_10_1914, i_10_1915, i_10_1948, i_10_2001, i_10_2005, i_10_2028, i_10_2244, i_10_2351, i_10_2353, i_10_2355, i_10_2356, i_10_2357, i_10_2359, i_10_2362, i_10_2363, i_10_2364, i_10_2451, i_10_2452, i_10_2453, i_10_2466, i_10_2478, i_10_2515, i_10_2565, i_10_2571, i_10_2677, i_10_2728, i_10_2781, i_10_2784, i_10_2823, i_10_2826, i_10_2827, i_10_2828, i_10_2869, i_10_3271, i_10_3273, i_10_3278, i_10_3279, i_10_3280, i_10_3281, i_10_3282, i_10_3283, i_10_3328, i_10_3430, i_10_3466, i_10_3471, i_10_3544, i_10_3582, i_10_3585, i_10_3586, i_10_3587, i_10_3590, i_10_3610, i_10_3684, i_10_3685, i_10_3721, i_10_3781, i_10_3788, i_10_3845, i_10_3983, i_10_4114, i_10_4119, i_10_4120, i_10_4128, i_10_4174, i_10_4269, i_10_4272, i_10_4287, i_10_4290, i_10_4291, i_10_4584, o_10_148);
	kernel_10_149 k_10_149(i_10_29, i_10_86, i_10_122, i_10_280, i_10_435, i_10_438, i_10_503, i_10_585, i_10_739, i_10_751, i_10_800, i_10_853, i_10_854, i_10_930, i_10_995, i_10_1006, i_10_1054, i_10_1223, i_10_1234, i_10_1239, i_10_1354, i_10_1579, i_10_1733, i_10_1736, i_10_1807, i_10_1819, i_10_1914, i_10_1916, i_10_1919, i_10_1925, i_10_1981, i_10_1995, i_10_1996, i_10_2002, i_10_2093, i_10_2096, i_10_2306, i_10_2354, i_10_2362, i_10_2452, i_10_2470, i_10_2475, i_10_2542, i_10_2543, i_10_2567, i_10_2573, i_10_2629, i_10_2641, i_10_2704, i_10_2724, i_10_2725, i_10_2801, i_10_2828, i_10_2831, i_10_2882, i_10_2883, i_10_2884, i_10_2917, i_10_2919, i_10_3082, i_10_3088, i_10_3090, i_10_3091, i_10_3124, i_10_3173, i_10_3278, i_10_3281, i_10_3353, i_10_3385, i_10_3406, i_10_3407, i_10_3409, i_10_3465, i_10_3473, i_10_3508, i_10_3586, i_10_3612, i_10_3650, i_10_3685, i_10_3686, i_10_3702, i_10_3748, i_10_3786, i_10_3832, i_10_3834, i_10_3849, i_10_3853, i_10_3901, i_10_3984, i_10_3988, i_10_4029, i_10_4030, i_10_4128, i_10_4130, i_10_4211, i_10_4216, i_10_4236, i_10_4272, i_10_4289, i_10_4566, o_10_149);
	kernel_10_150 k_10_150(i_10_263, i_10_280, i_10_282, i_10_327, i_10_393, i_10_411, i_10_438, i_10_509, i_10_511, i_10_512, i_10_718, i_10_961, i_10_1026, i_10_1035, i_10_1135, i_10_1239, i_10_1431, i_10_1576, i_10_1683, i_10_1684, i_10_1686, i_10_1689, i_10_1690, i_10_1821, i_10_1822, i_10_1825, i_10_1980, i_10_1998, i_10_2001, i_10_2006, i_10_2025, i_10_2028, i_10_2032, i_10_2199, i_10_2361, i_10_2362, i_10_2364, i_10_2365, i_10_2407, i_10_2452, i_10_2461, i_10_2466, i_10_2469, i_10_2506, i_10_2630, i_10_2658, i_10_2659, i_10_2680, i_10_2700, i_10_2701, i_10_2703, i_10_2704, i_10_2716, i_10_2718, i_10_2719, i_10_2727, i_10_2730, i_10_2733, i_10_2734, i_10_2785, i_10_2788, i_10_2827, i_10_2831, i_10_2885, i_10_3037, i_10_3153, i_10_3154, i_10_3195, i_10_3196, i_10_3198, i_10_3277, i_10_3279, i_10_3280, i_10_3283, i_10_3312, i_10_3386, i_10_3388, i_10_3391, i_10_3465, i_10_3468, i_10_3507, i_10_3588, i_10_3646, i_10_3647, i_10_3650, i_10_3684, i_10_3783, i_10_3786, i_10_3840, i_10_3846, i_10_3982, i_10_3983, i_10_4116, i_10_4117, i_10_4120, i_10_4126, i_10_4266, i_10_4281, i_10_4290, i_10_4570, o_10_150);
	kernel_10_151 k_10_151(i_10_48, i_10_82, i_10_216, i_10_219, i_10_245, i_10_270, i_10_280, i_10_281, i_10_282, i_10_283, i_10_322, i_10_405, i_10_424, i_10_435, i_10_436, i_10_459, i_10_460, i_10_467, i_10_891, i_10_902, i_10_1026, i_10_1163, i_10_1236, i_10_1263, i_10_1307, i_10_1432, i_10_1433, i_10_1441, i_10_1444, i_10_1485, i_10_1539, i_10_1540, i_10_1579, i_10_1652, i_10_1687, i_10_1688, i_10_1767, i_10_1768, i_10_1824, i_10_1825, i_10_1826, i_10_1911, i_10_1912, i_10_2200, i_10_2325, i_10_2351, i_10_2449, i_10_2628, i_10_2631, i_10_2637, i_10_2655, i_10_2656, i_10_2658, i_10_2659, i_10_2660, i_10_2673, i_10_2674, i_10_2700, i_10_2702, i_10_2718, i_10_2719, i_10_2720, i_10_2721, i_10_2722, i_10_2723, i_10_2729, i_10_2781, i_10_2826, i_10_2884, i_10_2885, i_10_2921, i_10_2985, i_10_3033, i_10_3045, i_10_3070, i_10_3071, i_10_3154, i_10_3159, i_10_3196, i_10_3326, i_10_3388, i_10_3391, i_10_3405, i_10_3470, i_10_3522, i_10_3523, i_10_3645, i_10_3682, i_10_3782, i_10_3847, i_10_3855, i_10_3856, i_10_3857, i_10_3906, i_10_3907, i_10_3979, i_10_4117, i_10_4118, i_10_4123, i_10_4287, o_10_151);
	kernel_10_152 k_10_152(i_10_153, i_10_175, i_10_220, i_10_257, i_10_315, i_10_316, i_10_392, i_10_432, i_10_437, i_10_464, i_10_561, i_10_588, i_10_799, i_10_1034, i_10_1039, i_10_1087, i_10_1234, i_10_1236, i_10_1239, i_10_1310, i_10_1355, i_10_1385, i_10_1432, i_10_1436, i_10_1448, i_10_1542, i_10_1543, i_10_1549, i_10_1551, i_10_1576, i_10_1655, i_10_1686, i_10_1687, i_10_1729, i_10_1732, i_10_1824, i_10_1826, i_10_1880, i_10_1951, i_10_1982, i_10_1984, i_10_1987, i_10_2107, i_10_2108, i_10_2158, i_10_2204, i_10_2331, i_10_2338, i_10_2352, i_10_2364, i_10_2383, i_10_2468, i_10_2538, i_10_2541, i_10_2632, i_10_2640, i_10_2731, i_10_2734, i_10_2820, i_10_2826, i_10_2827, i_10_2831, i_10_2881, i_10_2884, i_10_3043, i_10_3070, i_10_3071, i_10_3074, i_10_3075, i_10_3271, i_10_3277, i_10_3278, i_10_3282, i_10_3318, i_10_3354, i_10_3384, i_10_3433, i_10_3471, i_10_3540, i_10_3541, i_10_3542, i_10_3645, i_10_3652, i_10_3811, i_10_3851, i_10_3944, i_10_4086, i_10_4127, i_10_4172, i_10_4173, i_10_4174, i_10_4175, i_10_4219, i_10_4279, i_10_4280, i_10_4281, i_10_4282, i_10_4459, i_10_4533, i_10_4568, o_10_152);
	kernel_10_153 k_10_153(i_10_171, i_10_244, i_10_245, i_10_253, i_10_254, i_10_279, i_10_283, i_10_284, i_10_329, i_10_392, i_10_434, i_10_441, i_10_442, i_10_443, i_10_514, i_10_515, i_10_542, i_10_712, i_10_713, i_10_748, i_10_793, i_10_794, i_10_797, i_10_956, i_10_1000, i_10_1027, i_10_1028, i_10_1162, i_10_1234, i_10_1235, i_10_1237, i_10_1243, i_10_1244, i_10_1306, i_10_1310, i_10_1347, i_10_1540, i_10_1541, i_10_1549, i_10_1580, i_10_1650, i_10_1655, i_10_1684, i_10_1687, i_10_1688, i_10_1821, i_10_1823, i_10_2305, i_10_2306, i_10_2333, i_10_2349, i_10_2359, i_10_2361, i_10_2377, i_10_2452, i_10_2467, i_10_2512, i_10_2531, i_10_2603, i_10_2629, i_10_2632, i_10_2657, i_10_2660, i_10_2701, i_10_2711, i_10_2730, i_10_2732, i_10_2783, i_10_2827, i_10_3072, i_10_3073, i_10_3074, i_10_3196, i_10_3199, i_10_3200, i_10_3332, i_10_3384, i_10_3385, i_10_3388, i_10_3391, i_10_3409, i_10_3586, i_10_3587, i_10_3613, i_10_3614, i_10_3650, i_10_3781, i_10_3782, i_10_3784, i_10_3785, i_10_3788, i_10_3835, i_10_3838, i_10_3841, i_10_3842, i_10_4115, i_10_4123, i_10_4125, i_10_4126, i_10_4565, o_10_153);
	kernel_10_154 k_10_154(i_10_27, i_10_187, i_10_188, i_10_223, i_10_284, i_10_315, i_10_316, i_10_317, i_10_323, i_10_329, i_10_409, i_10_445, i_10_446, i_10_458, i_10_515, i_10_793, i_10_797, i_10_798, i_10_800, i_10_954, i_10_966, i_10_1001, i_10_1028, i_10_1234, i_10_1309, i_10_1310, i_10_1345, i_10_1432, i_10_1444, i_10_1547, i_10_1555, i_10_1582, i_10_1583, i_10_1648, i_10_1822, i_10_1823, i_10_1952, i_10_2179, i_10_2353, i_10_2354, i_10_2356, i_10_2357, i_10_2363, i_10_2381, i_10_2450, i_10_2453, i_10_2632, i_10_2659, i_10_2702, i_10_2707, i_10_2718, i_10_2719, i_10_2720, i_10_2722, i_10_2828, i_10_2833, i_10_2884, i_10_2920, i_10_2923, i_10_2924, i_10_3037, i_10_3070, i_10_3071, i_10_3152, i_10_3277, i_10_3278, i_10_3281, i_10_3324, i_10_3390, i_10_3391, i_10_3466, i_10_3467, i_10_3519, i_10_3586, i_10_3612, i_10_3613, i_10_3614, i_10_3617, i_10_3653, i_10_3780, i_10_3781, i_10_3784, i_10_3786, i_10_3788, i_10_3835, i_10_3837, i_10_3838, i_10_3848, i_10_3856, i_10_3857, i_10_3890, i_10_3907, i_10_4114, i_10_4115, i_10_4282, i_10_4283, i_10_4287, i_10_4288, i_10_4289, i_10_4564, o_10_154);
	kernel_10_155 k_10_155(i_10_177, i_10_246, i_10_249, i_10_252, i_10_264, i_10_318, i_10_320, i_10_321, i_10_322, i_10_327, i_10_413, i_10_462, i_10_933, i_10_1002, i_10_1007, i_10_1030, i_10_1032, i_10_1107, i_10_1110, i_10_1299, i_10_1302, i_10_1307, i_10_1431, i_10_1434, i_10_1437, i_10_1545, i_10_1581, i_10_1626, i_10_1654, i_10_1686, i_10_1731, i_10_1734, i_10_1735, i_10_1764, i_10_1806, i_10_1818, i_10_1821, i_10_1823, i_10_1983, i_10_1986, i_10_2031, i_10_2202, i_10_2349, i_10_2350, i_10_2351, i_10_2353, i_10_2358, i_10_2450, i_10_2472, i_10_2565, i_10_2568, i_10_2571, i_10_2604, i_10_2617, i_10_2663, i_10_2676, i_10_2680, i_10_2708, i_10_2712, i_10_2722, i_10_2734, i_10_2760, i_10_2826, i_10_2828, i_10_2847, i_10_2850, i_10_2920, i_10_2924, i_10_3045, i_10_3072, i_10_3073, i_10_3075, i_10_3202, i_10_3280, i_10_3390, i_10_3391, i_10_3434, i_10_3525, i_10_3540, i_10_3543, i_10_3544, i_10_3585, i_10_3617, i_10_3622, i_10_3645, i_10_3650, i_10_3787, i_10_3837, i_10_3854, i_10_3990, i_10_4029, i_10_4113, i_10_4115, i_10_4116, i_10_4117, i_10_4128, i_10_4168, i_10_4273, i_10_4584, i_10_4588, o_10_155);
	kernel_10_156 k_10_156(i_10_182, i_10_248, i_10_249, i_10_271, i_10_280, i_10_286, i_10_317, i_10_327, i_10_328, i_10_408, i_10_428, i_10_434, i_10_443, i_10_448, i_10_796, i_10_825, i_10_1029, i_10_1031, i_10_1033, i_10_1034, i_10_1118, i_10_1245, i_10_1441, i_10_1443, i_10_1492, i_10_1554, i_10_1582, i_10_1650, i_10_1675, i_10_1680, i_10_1682, i_10_1686, i_10_1818, i_10_1820, i_10_1822, i_10_1826, i_10_1909, i_10_1911, i_10_1947, i_10_2311, i_10_2354, i_10_2358, i_10_2407, i_10_2449, i_10_2450, i_10_2470, i_10_2471, i_10_2473, i_10_2633, i_10_2657, i_10_2658, i_10_2662, i_10_2704, i_10_2709, i_10_2710, i_10_2711, i_10_2714, i_10_2717, i_10_2722, i_10_2723, i_10_2731, i_10_2732, i_10_2826, i_10_2828, i_10_2872, i_10_2917, i_10_2918, i_10_2919, i_10_2921, i_10_3034, i_10_3035, i_10_3036, i_10_3163, i_10_3196, i_10_3199, i_10_3283, i_10_3326, i_10_3389, i_10_3392, i_10_3436, i_10_3470, i_10_3471, i_10_3585, i_10_3586, i_10_3588, i_10_3589, i_10_3647, i_10_3783, i_10_3854, i_10_3894, i_10_3947, i_10_3984, i_10_3985, i_10_3991, i_10_4121, i_10_4126, i_10_4216, i_10_4279, i_10_4284, i_10_4566, o_10_156);
	kernel_10_157 k_10_157(i_10_40, i_10_64, i_10_67, i_10_151, i_10_181, i_10_221, i_10_223, i_10_271, i_10_283, i_10_290, i_10_319, i_10_320, i_10_362, i_10_412, i_10_424, i_10_432, i_10_437, i_10_444, i_10_448, i_10_496, i_10_559, i_10_635, i_10_718, i_10_900, i_10_907, i_10_927, i_10_928, i_10_958, i_10_990, i_10_1009, i_10_1200, i_10_1236, i_10_1238, i_10_1241, i_10_1272, i_10_1275, i_10_1278, i_10_1310, i_10_1363, i_10_1364, i_10_1491, i_10_1579, i_10_1705, i_10_1783, i_10_1824, i_10_1849, i_10_1940, i_10_1943, i_10_2003, i_10_2052, i_10_2089, i_10_2264, i_10_2338, i_10_2350, i_10_2385, i_10_2452, i_10_2455, i_10_2476, i_10_2512, i_10_2596, i_10_2711, i_10_2714, i_10_2783, i_10_2830, i_10_2831, i_10_2910, i_10_2953, i_10_3011, i_10_3045, i_10_3050, i_10_3163, i_10_3198, i_10_3273, i_10_3275, i_10_3276, i_10_3281, i_10_3284, i_10_3286, i_10_3317, i_10_3386, i_10_3391, i_10_3469, i_10_3584, i_10_3585, i_10_3612, i_10_3648, i_10_3649, i_10_3682, i_10_3856, i_10_3860, i_10_3947, i_10_4050, i_10_4126, i_10_4157, i_10_4162, i_10_4192, i_10_4217, i_10_4282, i_10_4307, i_10_4519, o_10_157);
	kernel_10_158 k_10_158(i_10_172, i_10_223, i_10_245, i_10_251, i_10_254, i_10_282, i_10_284, i_10_390, i_10_406, i_10_426, i_10_441, i_10_443, i_10_459, i_10_460, i_10_463, i_10_747, i_10_748, i_10_749, i_10_793, i_10_794, i_10_796, i_10_797, i_10_1004, i_10_1026, i_10_1027, i_10_1033, i_10_1240, i_10_1306, i_10_1310, i_10_1365, i_10_1432, i_10_1433, i_10_1539, i_10_1540, i_10_1541, i_10_1543, i_10_1544, i_10_1576, i_10_1649, i_10_1683, i_10_1687, i_10_1821, i_10_1822, i_10_1954, i_10_2180, i_10_2351, i_10_2361, i_10_2450, i_10_2453, i_10_2461, i_10_2572, i_10_2628, i_10_2657, i_10_2674, i_10_2675, i_10_2701, i_10_2720, i_10_2733, i_10_2734, i_10_2817, i_10_2818, i_10_2821, i_10_2884, i_10_2923, i_10_2924, i_10_3035, i_10_3048, i_10_3049, i_10_3069, i_10_3070, i_10_3198, i_10_3199, i_10_3200, i_10_3270, i_10_3331, i_10_3405, i_10_3522, i_10_3525, i_10_3611, i_10_3612, i_10_3685, i_10_3686, i_10_3780, i_10_3782, i_10_3783, i_10_3784, i_10_3785, i_10_3837, i_10_3838, i_10_3842, i_10_3857, i_10_3858, i_10_3859, i_10_4117, i_10_4120, i_10_4121, i_10_4266, i_10_4269, i_10_4276, i_10_4568, o_10_158);
	kernel_10_159 k_10_159(i_10_29, i_10_172, i_10_273, i_10_284, i_10_388, i_10_409, i_10_410, i_10_442, i_10_459, i_10_508, i_10_511, i_10_512, i_10_796, i_10_800, i_10_958, i_10_1001, i_10_1004, i_10_1034, i_10_1081, i_10_1267, i_10_1433, i_10_1439, i_10_1576, i_10_1654, i_10_1655, i_10_1683, i_10_1690, i_10_1691, i_10_1736, i_10_1821, i_10_1822, i_10_1823, i_10_1824, i_10_1825, i_10_1913, i_10_1916, i_10_1946, i_10_2006, i_10_2030, i_10_2033, i_10_2381, i_10_2408, i_10_2449, i_10_2455, i_10_2472, i_10_2474, i_10_2608, i_10_2634, i_10_2635, i_10_2675, i_10_2722, i_10_2723, i_10_2730, i_10_2734, i_10_2735, i_10_2830, i_10_2831, i_10_2833, i_10_2885, i_10_2887, i_10_2922, i_10_2923, i_10_2986, i_10_3035, i_10_3049, i_10_3088, i_10_3320, i_10_3323, i_10_3384, i_10_3385, i_10_3386, i_10_3388, i_10_3389, i_10_3437, i_10_3470, i_10_3473, i_10_3509, i_10_3539, i_10_3584, i_10_3587, i_10_3590, i_10_3617, i_10_3784, i_10_3837, i_10_3839, i_10_3841, i_10_3842, i_10_3843, i_10_3853, i_10_3860, i_10_3890, i_10_3980, i_10_4114, i_10_4115, i_10_4174, i_10_4268, i_10_4271, i_10_4274, i_10_4287, i_10_4568, o_10_159);
	kernel_10_160 k_10_160(i_10_34, i_10_153, i_10_220, i_10_248, i_10_256, i_10_272, i_10_286, i_10_327, i_10_330, i_10_358, i_10_466, i_10_495, i_10_504, i_10_513, i_10_637, i_10_711, i_10_954, i_10_963, i_10_1026, i_10_1031, i_10_1032, i_10_1162, i_10_1165, i_10_1241, i_10_1242, i_10_1309, i_10_1545, i_10_1546, i_10_1561, i_10_1635, i_10_1651, i_10_1690, i_10_1691, i_10_1794, i_10_1821, i_10_1823, i_10_1909, i_10_1947, i_10_1984, i_10_2182, i_10_2256, i_10_2257, i_10_2323, i_10_2353, i_10_2385, i_10_2386, i_10_2455, i_10_2629, i_10_2633, i_10_2824, i_10_2833, i_10_2871, i_10_2893, i_10_2923, i_10_2924, i_10_2953, i_10_2986, i_10_3036, i_10_3037, i_10_3069, i_10_3073, i_10_3202, i_10_3203, i_10_3234, i_10_3291, i_10_3385, i_10_3387, i_10_3390, i_10_3409, i_10_3465, i_10_3492, i_10_3537, i_10_3580, i_10_3612, i_10_3682, i_10_3683, i_10_3730, i_10_3732, i_10_3774, i_10_3786, i_10_3787, i_10_3801, i_10_3807, i_10_3826, i_10_3844, i_10_3858, i_10_3860, i_10_3992, i_10_4009, i_10_4117, i_10_4134, i_10_4216, i_10_4219, i_10_4263, i_10_4264, i_10_4305, i_10_4436, i_10_4486, i_10_4567, i_10_4584, o_10_160);
	kernel_10_161 k_10_161(i_10_185, i_10_221, i_10_254, i_10_269, i_10_279, i_10_280, i_10_281, i_10_282, i_10_285, i_10_319, i_10_320, i_10_321, i_10_327, i_10_328, i_10_438, i_10_439, i_10_443, i_10_445, i_10_446, i_10_462, i_10_463, i_10_464, i_10_466, i_10_467, i_10_511, i_10_1030, i_10_1037, i_10_1240, i_10_1244, i_10_1245, i_10_1247, i_10_1248, i_10_1250, i_10_1363, i_10_1365, i_10_1546, i_10_1552, i_10_1554, i_10_1690, i_10_1819, i_10_1821, i_10_1822, i_10_1823, i_10_1945, i_10_1952, i_10_2185, i_10_2306, i_10_2323, i_10_2351, i_10_2353, i_10_2354, i_10_2355, i_10_2356, i_10_2467, i_10_2470, i_10_2515, i_10_2617, i_10_2630, i_10_2632, i_10_2634, i_10_2654, i_10_2662, i_10_2720, i_10_2724, i_10_2734, i_10_2735, i_10_2833, i_10_2887, i_10_2916, i_10_2919, i_10_2920, i_10_2921, i_10_2924, i_10_2986, i_10_3037, i_10_3038, i_10_3093, i_10_3154, i_10_3155, i_10_3163, i_10_3196, i_10_3197, i_10_3198, i_10_3199, i_10_3200, i_10_3281, i_10_3283, i_10_3328, i_10_3390, i_10_3407, i_10_3611, i_10_3650, i_10_3785, i_10_3838, i_10_3839, i_10_3842, i_10_4183, i_10_4569, i_10_4570, i_10_4571, o_10_161);
	kernel_10_162 k_10_162(i_10_30, i_10_123, i_10_174, i_10_178, i_10_183, i_10_221, i_10_429, i_10_430, i_10_464, i_10_500, i_10_535, i_10_564, i_10_898, i_10_951, i_10_996, i_10_1033, i_10_1114, i_10_1119, i_10_1237, i_10_1241, i_10_1309, i_10_1312, i_10_1345, i_10_1349, i_10_1489, i_10_1541, i_10_1542, i_10_1576, i_10_1618, i_10_1623, i_10_1624, i_10_1683, i_10_1684, i_10_1686, i_10_1768, i_10_1770, i_10_1824, i_10_1908, i_10_1912, i_10_1957, i_10_2004, i_10_2348, i_10_2364, i_10_2471, i_10_2515, i_10_2517, i_10_2519, i_10_2562, i_10_2567, i_10_2651, i_10_2652, i_10_2653, i_10_2658, i_10_2662, i_10_2715, i_10_2716, i_10_2722, i_10_2723, i_10_2725, i_10_2829, i_10_2830, i_10_2919, i_10_2966, i_10_2980, i_10_3071, i_10_3090, i_10_3093, i_10_3094, i_10_3166, i_10_3198, i_10_3199, i_10_3407, i_10_3410, i_10_3434, i_10_3472, i_10_3611, i_10_3612, i_10_3615, i_10_3624, i_10_3702, i_10_3705, i_10_3723, i_10_3797, i_10_3837, i_10_3855, i_10_3857, i_10_3883, i_10_3922, i_10_3982, i_10_3985, i_10_4026, i_10_4114, i_10_4117, i_10_4156, i_10_4175, i_10_4219, i_10_4236, i_10_4270, i_10_4425, i_10_4582, o_10_162);
	kernel_10_163 k_10_163(i_10_322, i_10_393, i_10_409, i_10_429, i_10_437, i_10_438, i_10_442, i_10_445, i_10_447, i_10_460, i_10_589, i_10_699, i_10_700, i_10_732, i_10_733, i_10_736, i_10_750, i_10_795, i_10_827, i_10_956, i_10_960, i_10_994, i_10_995, i_10_997, i_10_1060, i_10_1237, i_10_1238, i_10_1240, i_10_1241, i_10_1308, i_10_1343, i_10_1346, i_10_1576, i_10_1651, i_10_1684, i_10_1685, i_10_1688, i_10_1957, i_10_2184, i_10_2185, i_10_2364, i_10_2461, i_10_2463, i_10_2469, i_10_2470, i_10_2473, i_10_2632, i_10_2635, i_10_2659, i_10_2660, i_10_2698, i_10_2701, i_10_2702, i_10_2727, i_10_2728, i_10_2735, i_10_2821, i_10_2883, i_10_2884, i_10_2885, i_10_2886, i_10_2887, i_10_2888, i_10_2920, i_10_2922, i_10_2958, i_10_2959, i_10_3036, i_10_3037, i_10_3038, i_10_3198, i_10_3201, i_10_3202, i_10_3271, i_10_3279, i_10_3282, i_10_3283, i_10_3354, i_10_3406, i_10_3522, i_10_3543, i_10_3544, i_10_3588, i_10_3612, i_10_3702, i_10_3784, i_10_3787, i_10_3814, i_10_3837, i_10_3853, i_10_3854, i_10_3981, i_10_3984, i_10_3985, i_10_3989, i_10_4028, i_10_4119, i_10_4273, i_10_4285, i_10_4519, o_10_163);
	kernel_10_164 k_10_164(i_10_46, i_10_223, i_10_243, i_10_244, i_10_245, i_10_285, i_10_315, i_10_316, i_10_360, i_10_445, i_10_712, i_10_956, i_10_1026, i_10_1028, i_10_1044, i_10_1235, i_10_1243, i_10_1308, i_10_1309, i_10_1539, i_10_1540, i_10_1541, i_10_1576, i_10_1579, i_10_1649, i_10_1650, i_10_1651, i_10_1683, i_10_1685, i_10_1686, i_10_1955, i_10_2016, i_10_2178, i_10_2179, i_10_2180, i_10_2199, i_10_2304, i_10_2305, i_10_2307, i_10_2351, i_10_2353, i_10_2354, i_10_2451, i_10_2452, i_10_2455, i_10_2470, i_10_2471, i_10_2545, i_10_2569, i_10_2601, i_10_2602, i_10_2605, i_10_2662, i_10_2678, i_10_2703, i_10_2704, i_10_2719, i_10_2726, i_10_2728, i_10_2730, i_10_2738, i_10_2826, i_10_2827, i_10_3071, i_10_3196, i_10_3199, i_10_3200, i_10_3270, i_10_3331, i_10_3403, i_10_3405, i_10_3406, i_10_3493, i_10_3583, i_10_3585, i_10_3586, i_10_3588, i_10_3612, i_10_3613, i_10_3614, i_10_3615, i_10_3616, i_10_3646, i_10_3647, i_10_3720, i_10_3780, i_10_3781, i_10_3782, i_10_3783, i_10_3784, i_10_3785, i_10_3834, i_10_3844, i_10_3857, i_10_3909, i_10_4114, i_10_4115, i_10_4169, i_10_4171, i_10_4212, o_10_164);
	kernel_10_165 k_10_165(i_10_31, i_10_42, i_10_223, i_10_255, i_10_263, i_10_284, i_10_390, i_10_409, i_10_428, i_10_446, i_10_448, i_10_459, i_10_460, i_10_501, i_10_504, i_10_733, i_10_993, i_10_999, i_10_1001, i_10_1002, i_10_1180, i_10_1235, i_10_1238, i_10_1246, i_10_1542, i_10_1551, i_10_1552, i_10_1578, i_10_1582, i_10_1583, i_10_1623, i_10_1649, i_10_1651, i_10_1684, i_10_1731, i_10_1732, i_10_1734, i_10_1764, i_10_1806, i_10_1813, i_10_1823, i_10_1981, i_10_1983, i_10_1991, i_10_2154, i_10_2304, i_10_2352, i_10_2353, i_10_2377, i_10_2378, i_10_2379, i_10_2455, i_10_2456, i_10_2565, i_10_2567, i_10_2568, i_10_2658, i_10_2661, i_10_2701, i_10_2727, i_10_2829, i_10_2881, i_10_2884, i_10_2952, i_10_2953, i_10_2982, i_10_3033, i_10_3054, i_10_3232, i_10_3277, i_10_3316, i_10_3318, i_10_3384, i_10_3472, i_10_3538, i_10_3610, i_10_3614, i_10_3616, i_10_3782, i_10_3835, i_10_3851, i_10_3906, i_10_3978, i_10_3979, i_10_3988, i_10_4114, i_10_4116, i_10_4117, i_10_4124, i_10_4266, i_10_4267, i_10_4269, i_10_4272, i_10_4275, i_10_4278, i_10_4281, i_10_4287, i_10_4288, i_10_4290, i_10_4566, o_10_165);
	kernel_10_166 k_10_166(i_10_174, i_10_175, i_10_179, i_10_220, i_10_262, i_10_282, i_10_283, i_10_321, i_10_322, i_10_450, i_10_711, i_10_797, i_10_799, i_10_957, i_10_958, i_10_960, i_10_967, i_10_999, i_10_1000, i_10_1083, i_10_1135, i_10_1169, i_10_1237, i_10_1240, i_10_1308, i_10_1310, i_10_1438, i_10_1679, i_10_1684, i_10_1687, i_10_1688, i_10_1819, i_10_1821, i_10_1822, i_10_1909, i_10_1911, i_10_1944, i_10_1945, i_10_1946, i_10_2184, i_10_2185, i_10_2203, i_10_2331, i_10_2350, i_10_2352, i_10_2353, i_10_2356, i_10_2376, i_10_2377, i_10_2404, i_10_2449, i_10_2452, i_10_2470, i_10_2502, i_10_2504, i_10_2711, i_10_2713, i_10_2716, i_10_2729, i_10_2734, i_10_2788, i_10_2880, i_10_2881, i_10_2885, i_10_2923, i_10_3034, i_10_3036, i_10_3042, i_10_3044, i_10_3150, i_10_3279, i_10_3280, i_10_3493, i_10_3610, i_10_3614, i_10_3687, i_10_3783, i_10_3786, i_10_3838, i_10_3840, i_10_3841, i_10_3843, i_10_3847, i_10_3851, i_10_3860, i_10_3877, i_10_3889, i_10_3978, i_10_3979, i_10_4050, i_10_4117, i_10_4122, i_10_4123, i_10_4129, i_10_4290, i_10_4291, i_10_4292, i_10_4564, i_10_4566, i_10_4567, o_10_166);
	kernel_10_167 k_10_167(i_10_33, i_10_174, i_10_175, i_10_178, i_10_285, i_10_286, i_10_332, i_10_390, i_10_442, i_10_447, i_10_448, i_10_459, i_10_460, i_10_467, i_10_800, i_10_1029, i_10_1034, i_10_1237, i_10_1238, i_10_1239, i_10_1308, i_10_1309, i_10_1545, i_10_1619, i_10_1648, i_10_1651, i_10_1687, i_10_1767, i_10_1769, i_10_1824, i_10_1825, i_10_1912, i_10_1950, i_10_1951, i_10_1952, i_10_1961, i_10_2004, i_10_2019, i_10_2185, i_10_2186, i_10_2436, i_10_2455, i_10_2515, i_10_2516, i_10_2631, i_10_2634, i_10_2635, i_10_2656, i_10_2707, i_10_2708, i_10_2710, i_10_2718, i_10_2723, i_10_2731, i_10_2757, i_10_2782, i_10_2788, i_10_2827, i_10_3036, i_10_3037, i_10_3040, i_10_3093, i_10_3094, i_10_3095, i_10_3198, i_10_3199, i_10_3202, i_10_3277, i_10_3278, i_10_3279, i_10_3280, i_10_3328, i_10_3407, i_10_3433, i_10_3466, i_10_3468, i_10_3469, i_10_3494, i_10_3496, i_10_3610, i_10_3613, i_10_3614, i_10_3650, i_10_3652, i_10_3702, i_10_3783, i_10_3784, i_10_3786, i_10_3838, i_10_3842, i_10_3855, i_10_3856, i_10_3857, i_10_3985, i_10_3991, i_10_4126, i_10_4129, i_10_4130, i_10_4273, i_10_4565, o_10_167);
	kernel_10_168 k_10_168(i_10_30, i_10_69, i_10_193, i_10_279, i_10_285, i_10_387, i_10_390, i_10_393, i_10_426, i_10_445, i_10_462, i_10_463, i_10_465, i_10_480, i_10_759, i_10_826, i_10_950, i_10_1029, i_10_1030, i_10_1031, i_10_1034, i_10_1260, i_10_1261, i_10_1262, i_10_1308, i_10_1353, i_10_1435, i_10_1498, i_10_1548, i_10_1579, i_10_1581, i_10_1617, i_10_1623, i_10_1650, i_10_1687, i_10_1691, i_10_1743, i_10_1756, i_10_1759, i_10_1803, i_10_1918, i_10_2164, i_10_2196, i_10_2198, i_10_2307, i_10_2311, i_10_2312, i_10_2338, i_10_2351, i_10_2352, i_10_2362, i_10_2433, i_10_2457, i_10_2460, i_10_2472, i_10_2559, i_10_2565, i_10_2568, i_10_2631, i_10_2634, i_10_2661, i_10_2830, i_10_2845, i_10_2865, i_10_3072, i_10_3201, i_10_3202, i_10_3267, i_10_3268, i_10_3333, i_10_3334, i_10_3392, i_10_3406, i_10_3465, i_10_3468, i_10_3609, i_10_3612, i_10_3615, i_10_3681, i_10_3685, i_10_3686, i_10_3688, i_10_3706, i_10_3727, i_10_3777, i_10_3781, i_10_3843, i_10_3844, i_10_3993, i_10_4098, i_10_4113, i_10_4121, i_10_4175, i_10_4218, i_10_4236, i_10_4290, i_10_4458, i_10_4477, i_10_4478, i_10_4561, o_10_168);
	kernel_10_169 k_10_169(i_10_172, i_10_178, i_10_279, i_10_280, i_10_282, i_10_423, i_10_428, i_10_429, i_10_430, i_10_433, i_10_435, i_10_436, i_10_438, i_10_439, i_10_440, i_10_441, i_10_447, i_10_465, i_10_507, i_10_717, i_10_748, i_10_751, i_10_793, i_10_800, i_10_1137, i_10_1138, i_10_1237, i_10_1238, i_10_1249, i_10_1305, i_10_1306, i_10_1308, i_10_1309, i_10_1579, i_10_1647, i_10_1683, i_10_1687, i_10_1819, i_10_1820, i_10_1823, i_10_2350, i_10_2351, i_10_2352, i_10_2353, i_10_2354, i_10_2453, i_10_2514, i_10_2516, i_10_2629, i_10_2634, i_10_2636, i_10_2703, i_10_2704, i_10_2706, i_10_2715, i_10_2718, i_10_2884, i_10_2885, i_10_2980, i_10_2986, i_10_3034, i_10_3036, i_10_3087, i_10_3093, i_10_3094, i_10_3154, i_10_3155, i_10_3165, i_10_3196, i_10_3198, i_10_3199, i_10_3200, i_10_3321, i_10_3322, i_10_3384, i_10_3405, i_10_3406, i_10_3407, i_10_3408, i_10_3409, i_10_3610, i_10_3613, i_10_3614, i_10_3615, i_10_3650, i_10_3702, i_10_3780, i_10_3782, i_10_3788, i_10_3837, i_10_3846, i_10_3856, i_10_3859, i_10_3982, i_10_4115, i_10_4273, i_10_4288, i_10_4564, i_10_4565, i_10_4568, o_10_169);
	kernel_10_170 k_10_170(i_10_51, i_10_83, i_10_223, i_10_280, i_10_281, i_10_282, i_10_286, i_10_289, i_10_394, i_10_430, i_10_512, i_10_516, i_10_743, i_10_751, i_10_823, i_10_824, i_10_852, i_10_896, i_10_1003, i_10_1030, i_10_1031, i_10_1112, i_10_1219, i_10_1300, i_10_1306, i_10_1309, i_10_1345, i_10_1346, i_10_1349, i_10_1357, i_10_1435, i_10_1439, i_10_1445, i_10_1493, i_10_1544, i_10_1556, i_10_1607, i_10_1652, i_10_1654, i_10_1803, i_10_1804, i_10_1820, i_10_1915, i_10_1996, i_10_1997, i_10_2184, i_10_2185, i_10_2291, i_10_2380, i_10_2444, i_10_2566, i_10_2567, i_10_2570, i_10_2604, i_10_2644, i_10_2674, i_10_2712, i_10_2713, i_10_2714, i_10_2730, i_10_2734, i_10_2742, i_10_2827, i_10_2867, i_10_2882, i_10_2965, i_10_2990, i_10_3046, i_10_3091, i_10_3162, i_10_3197, i_10_3391, i_10_3505, i_10_3558, i_10_3609, i_10_3653, i_10_3797, i_10_3841, i_10_3842, i_10_3859, i_10_3892, i_10_3893, i_10_3979, i_10_4026, i_10_4027, i_10_4028, i_10_4030, i_10_4129, i_10_4153, i_10_4154, i_10_4175, i_10_4193, i_10_4208, i_10_4237, i_10_4271, i_10_4278, i_10_4400, i_10_4455, i_10_4535, i_10_4553, o_10_170);
	kernel_10_171 k_10_171(i_10_177, i_10_184, i_10_220, i_10_223, i_10_291, i_10_321, i_10_329, i_10_394, i_10_411, i_10_426, i_10_427, i_10_430, i_10_444, i_10_448, i_10_467, i_10_511, i_10_693, i_10_694, i_10_730, i_10_733, i_10_796, i_10_797, i_10_800, i_10_961, i_10_970, i_10_999, i_10_1233, i_10_1234, i_10_1235, i_10_1238, i_10_1243, i_10_1363, i_10_1548, i_10_1549, i_10_1552, i_10_1578, i_10_1617, i_10_1734, i_10_1821, i_10_1823, i_10_1909, i_10_1912, i_10_1990, i_10_2358, i_10_2361, i_10_2362, i_10_2364, i_10_2365, i_10_2376, i_10_2383, i_10_2448, i_10_2716, i_10_2719, i_10_2823, i_10_2827, i_10_2829, i_10_2883, i_10_2884, i_10_2917, i_10_2953, i_10_2980, i_10_2982, i_10_2985, i_10_3034, i_10_3036, i_10_3038, i_10_3153, i_10_3154, i_10_3200, i_10_3273, i_10_3276, i_10_3279, i_10_3281, i_10_3282, i_10_3283, i_10_3324, i_10_3326, i_10_3784, i_10_3850, i_10_3852, i_10_3853, i_10_3855, i_10_3858, i_10_3859, i_10_3860, i_10_3888, i_10_3895, i_10_3912, i_10_3978, i_10_3979, i_10_3981, i_10_3982, i_10_3984, i_10_3985, i_10_3990, i_10_4113, i_10_4121, i_10_4281, i_10_4292, i_10_4570, o_10_171);
	kernel_10_172 k_10_172(i_10_70, i_10_71, i_10_157, i_10_185, i_10_283, i_10_285, i_10_286, i_10_316, i_10_434, i_10_445, i_10_447, i_10_562, i_10_563, i_10_953, i_10_1045, i_10_1080, i_10_1081, i_10_1160, i_10_1236, i_10_1237, i_10_1238, i_10_1267, i_10_1363, i_10_1544, i_10_1555, i_10_1577, i_10_1614, i_10_1627, i_10_1642, i_10_1654, i_10_1772, i_10_1922, i_10_2017, i_10_2159, i_10_2203, i_10_2240, i_10_2354, i_10_2356, i_10_2357, i_10_2361, i_10_2364, i_10_2365, i_10_2407, i_10_2436, i_10_2451, i_10_2452, i_10_2458, i_10_2461, i_10_2463, i_10_2464, i_10_2516, i_10_2518, i_10_2564, i_10_2570, i_10_2573, i_10_2602, i_10_2607, i_10_2633, i_10_2656, i_10_2658, i_10_2717, i_10_2826, i_10_2829, i_10_2830, i_10_2831, i_10_2834, i_10_2885, i_10_3036, i_10_3046, i_10_3074, i_10_3160, i_10_3199, i_10_3392, i_10_3519, i_10_3545, i_10_3563, i_10_3585, i_10_3586, i_10_3613, i_10_3721, i_10_3722, i_10_3788, i_10_3842, i_10_3850, i_10_3856, i_10_3857, i_10_3907, i_10_3923, i_10_3988, i_10_4120, i_10_4122, i_10_4123, i_10_4168, i_10_4169, i_10_4282, i_10_4283, i_10_4310, i_10_4435, i_10_4521, i_10_4565, o_10_172);
	kernel_10_173 k_10_173(i_10_133, i_10_221, i_10_257, i_10_263, i_10_269, i_10_282, i_10_405, i_10_409, i_10_442, i_10_566, i_10_626, i_10_793, i_10_1003, i_10_1004, i_10_1007, i_10_1016, i_10_1052, i_10_1106, i_10_1213, i_10_1234, i_10_1235, i_10_1237, i_10_1238, i_10_1267, i_10_1300, i_10_1303, i_10_1304, i_10_1305, i_10_1345, i_10_1540, i_10_1628, i_10_1683, i_10_1685, i_10_1686, i_10_1728, i_10_1729, i_10_1769, i_10_1771, i_10_1804, i_10_1823, i_10_1922, i_10_2006, i_10_2200, i_10_2362, i_10_2365, i_10_2436, i_10_2449, i_10_2453, i_10_2461, i_10_2563, i_10_2564, i_10_2607, i_10_2608, i_10_2631, i_10_2636, i_10_2658, i_10_2660, i_10_2711, i_10_2716, i_10_2734, i_10_2759, i_10_2762, i_10_2824, i_10_2831, i_10_2845, i_10_2870, i_10_2962, i_10_2963, i_10_3033, i_10_3036, i_10_3185, i_10_3200, i_10_3317, i_10_3389, i_10_3473, i_10_3526, i_10_3538, i_10_3540, i_10_3541, i_10_3542, i_10_3614, i_10_3702, i_10_3838, i_10_3839, i_10_3840, i_10_3843, i_10_3844, i_10_3858, i_10_3913, i_10_3986, i_10_4118, i_10_4151, i_10_4168, i_10_4169, i_10_4266, i_10_4274, i_10_4287, i_10_4428, i_10_4553, i_10_4565, o_10_173);
	kernel_10_174 k_10_174(i_10_89, i_10_177, i_10_179, i_10_267, i_10_283, i_10_317, i_10_389, i_10_390, i_10_407, i_10_441, i_10_460, i_10_713, i_10_795, i_10_993, i_10_1003, i_10_1121, i_10_1260, i_10_1360, i_10_1431, i_10_1540, i_10_1552, i_10_1683, i_10_1684, i_10_1685, i_10_1687, i_10_1688, i_10_1740, i_10_1771, i_10_1800, i_10_1801, i_10_1803, i_10_1804, i_10_1819, i_10_1821, i_10_1981, i_10_2000, i_10_2365, i_10_2449, i_10_2452, i_10_2539, i_10_2543, i_10_2565, i_10_2566, i_10_2608, i_10_2629, i_10_2631, i_10_2657, i_10_2673, i_10_2700, i_10_2702, i_10_2703, i_10_2704, i_10_2705, i_10_2709, i_10_2710, i_10_2713, i_10_2728, i_10_2729, i_10_2737, i_10_2782, i_10_2785, i_10_2786, i_10_2821, i_10_2828, i_10_2829, i_10_3040, i_10_3043, i_10_3073, i_10_3091, i_10_3114, i_10_3166, i_10_3233, i_10_3281, i_10_3385, i_10_3386, i_10_3388, i_10_3406, i_10_3407, i_10_3410, i_10_3542, i_10_3584, i_10_3645, i_10_3647, i_10_3648, i_10_3649, i_10_3650, i_10_3652, i_10_3811, i_10_3834, i_10_3837, i_10_3855, i_10_3902, i_10_3904, i_10_3906, i_10_4025, i_10_4115, i_10_4214, i_10_4290, i_10_4291, i_10_4568, o_10_174);
	kernel_10_175 k_10_175(i_10_221, i_10_248, i_10_280, i_10_281, i_10_284, i_10_328, i_10_388, i_10_391, i_10_536, i_10_621, i_10_635, i_10_639, i_10_659, i_10_716, i_10_722, i_10_946, i_10_967, i_10_998, i_10_1237, i_10_1296, i_10_1305, i_10_1378, i_10_1453, i_10_1540, i_10_1544, i_10_1546, i_10_1562, i_10_1565, i_10_1617, i_10_1705, i_10_1809, i_10_1877, i_10_1917, i_10_1999, i_10_2000, i_10_2008, i_10_2020, i_10_2021, i_10_2039, i_10_2054, i_10_2057, i_10_2109, i_10_2183, i_10_2305, i_10_2306, i_10_2326, i_10_2452, i_10_2454, i_10_2455, i_10_2456, i_10_2507, i_10_2515, i_10_2557, i_10_2602, i_10_2605, i_10_2663, i_10_2674, i_10_2675, i_10_2848, i_10_2909, i_10_2911, i_10_2953, i_10_2961, i_10_3073, i_10_3106, i_10_3203, i_10_3278, i_10_3284, i_10_3285, i_10_3376, i_10_3386, i_10_3410, i_10_3431, i_10_3604, i_10_3609, i_10_3699, i_10_3777, i_10_3785, i_10_3788, i_10_3857, i_10_3902, i_10_3919, i_10_3947, i_10_3979, i_10_4023, i_10_4024, i_10_4025, i_10_4114, i_10_4117, i_10_4122, i_10_4123, i_10_4149, i_10_4150, i_10_4216, i_10_4220, i_10_4267, i_10_4275, i_10_4411, i_10_4522, i_10_4523, o_10_175);
	kernel_10_176 k_10_176(i_10_34, i_10_121, i_10_122, i_10_124, i_10_132, i_10_133, i_10_177, i_10_178, i_10_183, i_10_331, i_10_367, i_10_374, i_10_386, i_10_429, i_10_437, i_10_439, i_10_440, i_10_462, i_10_599, i_10_600, i_10_602, i_10_634, i_10_754, i_10_755, i_10_906, i_10_967, i_10_971, i_10_1160, i_10_1240, i_10_1483, i_10_1499, i_10_1543, i_10_1627, i_10_1644, i_10_1645, i_10_1700, i_10_1727, i_10_1765, i_10_1781, i_10_1795, i_10_1796, i_10_1826, i_10_1913, i_10_2004, i_10_2060, i_10_2095, i_10_2245, i_10_2246, i_10_2248, i_10_2470, i_10_2473, i_10_2474, i_10_2512, i_10_2516, i_10_2534, i_10_2571, i_10_2572, i_10_2633, i_10_2708, i_10_2715, i_10_2789, i_10_2913, i_10_2914, i_10_2915, i_10_2958, i_10_2983, i_10_2984, i_10_3069, i_10_3095, i_10_3229, i_10_3356, i_10_3431, i_10_3451, i_10_3452, i_10_3471, i_10_3472, i_10_3473, i_10_3496, i_10_3545, i_10_3586, i_10_3589, i_10_3590, i_10_3603, i_10_3624, i_10_3625, i_10_3856, i_10_3857, i_10_3885, i_10_3949, i_10_3950, i_10_3979, i_10_4004, i_10_4058, i_10_4117, i_10_4120, i_10_4171, i_10_4265, i_10_4291, i_10_4426, i_10_4481, o_10_176);
	kernel_10_177 k_10_177(i_10_317, i_10_325, i_10_372, i_10_373, i_10_376, i_10_388, i_10_405, i_10_434, i_10_444, i_10_446, i_10_447, i_10_448, i_10_459, i_10_462, i_10_466, i_10_467, i_10_578, i_10_736, i_10_737, i_10_792, i_10_793, i_10_794, i_10_799, i_10_800, i_10_970, i_10_1002, i_10_1003, i_10_1006, i_10_1116, i_10_1163, i_10_1183, i_10_1242, i_10_1305, i_10_1306, i_10_1315, i_10_1344, i_10_1363, i_10_1441, i_10_1442, i_10_1543, i_10_1549, i_10_1642, i_10_1729, i_10_1730, i_10_1823, i_10_1826, i_10_1910, i_10_1948, i_10_2083, i_10_2154, i_10_2157, i_10_2158, i_10_2305, i_10_2309, i_10_2353, i_10_2404, i_10_2407, i_10_2408, i_10_2539, i_10_2633, i_10_2635, i_10_2705, i_10_2782, i_10_2880, i_10_2881, i_10_2887, i_10_2953, i_10_2956, i_10_2983, i_10_3058, i_10_3236, i_10_3316, i_10_3390, i_10_3494, i_10_3508, i_10_3688, i_10_3835, i_10_3859, i_10_3860, i_10_3889, i_10_3890, i_10_3919, i_10_3920, i_10_3928, i_10_3983, i_10_4087, i_10_4088, i_10_4266, i_10_4268, i_10_4270, i_10_4271, i_10_4273, i_10_4274, i_10_4288, i_10_4379, i_10_4460, i_10_4477, i_10_4569, i_10_4570, i_10_4571, o_10_177);
	kernel_10_178 k_10_178(i_10_28, i_10_82, i_10_174, i_10_176, i_10_246, i_10_289, i_10_793, i_10_954, i_10_955, i_10_961, i_10_993, i_10_1272, i_10_1359, i_10_1378, i_10_1575, i_10_1647, i_10_1648, i_10_1650, i_10_1683, i_10_1684, i_10_1686, i_10_1687, i_10_1691, i_10_1818, i_10_1819, i_10_1820, i_10_1916, i_10_1944, i_10_1945, i_10_1947, i_10_2178, i_10_2325, i_10_2361, i_10_2376, i_10_2379, i_10_2404, i_10_2448, i_10_2449, i_10_2450, i_10_2452, i_10_2453, i_10_2470, i_10_2502, i_10_2503, i_10_2505, i_10_2514, i_10_2601, i_10_2602, i_10_2610, i_10_2628, i_10_2631, i_10_2634, i_10_2637, i_10_2655, i_10_2663, i_10_2673, i_10_2674, i_10_2676, i_10_2700, i_10_2701, i_10_2703, i_10_2712, i_10_2727, i_10_2781, i_10_2882, i_10_2887, i_10_3033, i_10_3036, i_10_3042, i_10_3051, i_10_3267, i_10_3277, i_10_3280, i_10_3385, i_10_3386, i_10_3387, i_10_3388, i_10_3389, i_10_3447, i_10_3448, i_10_3611, i_10_3645, i_10_3646, i_10_3648, i_10_3649, i_10_3681, i_10_3783, i_10_3845, i_10_3852, i_10_3853, i_10_3854, i_10_3860, i_10_3894, i_10_3979, i_10_3981, i_10_4050, i_10_4113, i_10_4287, i_10_4564, i_10_4566, o_10_178);
	kernel_10_179 k_10_179(i_10_248, i_10_250, i_10_268, i_10_321, i_10_408, i_10_409, i_10_410, i_10_425, i_10_441, i_10_444, i_10_447, i_10_463, i_10_466, i_10_566, i_10_799, i_10_958, i_10_969, i_10_990, i_10_996, i_10_1031, i_10_1239, i_10_1250, i_10_1263, i_10_1307, i_10_1344, i_10_1345, i_10_1348, i_10_1439, i_10_1546, i_10_1576, i_10_1577, i_10_1686, i_10_1687, i_10_1818, i_10_1819, i_10_1909, i_10_1912, i_10_2022, i_10_2023, i_10_2032, i_10_2200, i_10_2201, i_10_2358, i_10_2359, i_10_2384, i_10_2456, i_10_2474, i_10_2633, i_10_2700, i_10_2709, i_10_2710, i_10_2713, i_10_2727, i_10_2731, i_10_2784, i_10_2785, i_10_2817, i_10_2818, i_10_2883, i_10_2884, i_10_2887, i_10_3034, i_10_3037, i_10_3038, i_10_3040, i_10_3069, i_10_3150, i_10_3151, i_10_3152, i_10_3155, i_10_3157, i_10_3284, i_10_3384, i_10_3385, i_10_3403, i_10_3472, i_10_3520, i_10_3522, i_10_3523, i_10_3525, i_10_3612, i_10_3613, i_10_3781, i_10_3784, i_10_3847, i_10_3856, i_10_3859, i_10_3983, i_10_3990, i_10_4114, i_10_4116, i_10_4119, i_10_4120, i_10_4121, i_10_4266, i_10_4267, i_10_4271, i_10_4273, i_10_4288, i_10_4290, o_10_179);
	kernel_10_180 k_10_180(i_10_22, i_10_23, i_10_86, i_10_245, i_10_248, i_10_262, i_10_283, i_10_284, i_10_317, i_10_319, i_10_320, i_10_391, i_10_439, i_10_460, i_10_464, i_10_479, i_10_496, i_10_497, i_10_832, i_10_932, i_10_947, i_10_1001, i_10_1085, i_10_1223, i_10_1240, i_10_1243, i_10_1267, i_10_1301, i_10_1328, i_10_1346, i_10_1433, i_10_1445, i_10_1487, i_10_1541, i_10_1544, i_10_1577, i_10_1607, i_10_1622, i_10_1624, i_10_1625, i_10_1687, i_10_1714, i_10_1741, i_10_1805, i_10_1821, i_10_1826, i_10_1931, i_10_2017, i_10_2018, i_10_2026, i_10_2027, i_10_2110, i_10_2111, i_10_2162, i_10_2198, i_10_2204, i_10_2359, i_10_2366, i_10_2453, i_10_2567, i_10_2602, i_10_2605, i_10_2606, i_10_2663, i_10_2702, i_10_2705, i_10_2719, i_10_2725, i_10_2732, i_10_2846, i_10_2924, i_10_3025, i_10_3044, i_10_3070, i_10_3077, i_10_3167, i_10_3317, i_10_3332, i_10_3377, i_10_3389, i_10_3523, i_10_3557, i_10_3602, i_10_3613, i_10_3722, i_10_3725, i_10_3772, i_10_3835, i_10_3841, i_10_3851, i_10_3856, i_10_3916, i_10_3989, i_10_4096, i_10_4097, i_10_4114, i_10_4117, i_10_4123, i_10_4124, i_10_4276, o_10_180);
	kernel_10_181 k_10_181(i_10_85, i_10_86, i_10_155, i_10_158, i_10_243, i_10_245, i_10_246, i_10_287, i_10_319, i_10_374, i_10_405, i_10_423, i_10_436, i_10_460, i_10_462, i_10_463, i_10_466, i_10_948, i_10_990, i_10_991, i_10_992, i_10_1031, i_10_1053, i_10_1173, i_10_1201, i_10_1202, i_10_1217, i_10_1260, i_10_1307, i_10_1358, i_10_1443, i_10_1444, i_10_1543, i_10_1596, i_10_1608, i_10_1622, i_10_1647, i_10_1648, i_10_1649, i_10_1651, i_10_1713, i_10_1994, i_10_2000, i_10_2016, i_10_2018, i_10_2201, i_10_2204, i_10_2324, i_10_2357, i_10_2459, i_10_2460, i_10_2512, i_10_2513, i_10_2606, i_10_2641, i_10_2659, i_10_2660, i_10_2720, i_10_2721, i_10_2725, i_10_2726, i_10_2782, i_10_2828, i_10_2834, i_10_2884, i_10_2964, i_10_2965, i_10_2981, i_10_2984, i_10_3044, i_10_3083, i_10_3201, i_10_3259, i_10_3272, i_10_3442, i_10_3443, i_10_3611, i_10_3721, i_10_3722, i_10_3788, i_10_3807, i_10_3830, i_10_3857, i_10_3860, i_10_3893, i_10_3910, i_10_3926, i_10_3980, i_10_3988, i_10_4030, i_10_4031, i_10_4114, i_10_4115, i_10_4169, i_10_4214, i_10_4277, i_10_4286, i_10_4317, i_10_4456, i_10_4521, o_10_181);
	kernel_10_182 k_10_182(i_10_172, i_10_244, i_10_246, i_10_247, i_10_253, i_10_276, i_10_286, i_10_405, i_10_426, i_10_427, i_10_460, i_10_467, i_10_747, i_10_748, i_10_954, i_10_955, i_10_956, i_10_962, i_10_1026, i_10_1029, i_10_1234, i_10_1236, i_10_1237, i_10_1241, i_10_1243, i_10_1308, i_10_1309, i_10_1311, i_10_1312, i_10_1540, i_10_1542, i_10_1545, i_10_1650, i_10_1686, i_10_1688, i_10_1818, i_10_1819, i_10_1820, i_10_1826, i_10_1953, i_10_2196, i_10_2351, i_10_2354, i_10_2450, i_10_2452, i_10_2469, i_10_2474, i_10_2601, i_10_2674, i_10_2677, i_10_2710, i_10_2711, i_10_2719, i_10_2731, i_10_2917, i_10_2924, i_10_2980, i_10_3036, i_10_3072, i_10_3075, i_10_3198, i_10_3199, i_10_3200, i_10_3202, i_10_3385, i_10_3408, i_10_3522, i_10_3523, i_10_3582, i_10_3585, i_10_3586, i_10_3612, i_10_3613, i_10_3615, i_10_3646, i_10_3648, i_10_3649, i_10_3780, i_10_3781, i_10_3782, i_10_3783, i_10_3784, i_10_3786, i_10_3787, i_10_3788, i_10_3835, i_10_3840, i_10_3856, i_10_4113, i_10_4114, i_10_4116, i_10_4117, i_10_4216, i_10_4267, i_10_4284, i_10_4288, i_10_4563, i_10_4564, i_10_4567, i_10_4568, o_10_182);
	kernel_10_183 k_10_183(i_10_117, i_10_118, i_10_136, i_10_146, i_10_175, i_10_216, i_10_220, i_10_263, i_10_284, i_10_308, i_10_347, i_10_390, i_10_391, i_10_435, i_10_508, i_10_509, i_10_689, i_10_748, i_10_892, i_10_901, i_10_902, i_10_963, i_10_1045, i_10_1046, i_10_1083, i_10_1234, i_10_1238, i_10_1246, i_10_1247, i_10_1432, i_10_1433, i_10_1451, i_10_1534, i_10_1621, i_10_1622, i_10_1683, i_10_1686, i_10_1689, i_10_1691, i_10_1821, i_10_1901, i_10_1908, i_10_1909, i_10_1944, i_10_2035, i_10_2161, i_10_2243, i_10_2246, i_10_2252, i_10_2326, i_10_2448, i_10_2449, i_10_2453, i_10_2467, i_10_2468, i_10_2469, i_10_2512, i_10_2513, i_10_2544, i_10_2565, i_10_2629, i_10_2630, i_10_2632, i_10_2638, i_10_2655, i_10_2656, i_10_2663, i_10_2700, i_10_2718, i_10_2723, i_10_2728, i_10_2911, i_10_3043, i_10_3069, i_10_3071, i_10_3170, i_10_3392, i_10_3408, i_10_3409, i_10_3449, i_10_3465, i_10_3469, i_10_3527, i_10_3538, i_10_3555, i_10_3562, i_10_3583, i_10_3609, i_10_3837, i_10_3856, i_10_4121, i_10_4122, i_10_4278, i_10_4285, i_10_4286, i_10_4288, i_10_4289, i_10_4428, i_10_4570, i_10_4582, o_10_183);
	kernel_10_184 k_10_184(i_10_64, i_10_180, i_10_243, i_10_262, i_10_408, i_10_424, i_10_429, i_10_430, i_10_444, i_10_445, i_10_462, i_10_467, i_10_831, i_10_921, i_10_954, i_10_955, i_10_956, i_10_957, i_10_959, i_10_962, i_10_1002, i_10_1026, i_10_1034, i_10_1080, i_10_1161, i_10_1162, i_10_1233, i_10_1287, i_10_1488, i_10_1494, i_10_1533, i_10_1579, i_10_1614, i_10_1638, i_10_1854, i_10_1872, i_10_1910, i_10_1914, i_10_1944, i_10_1945, i_10_2088, i_10_2202, i_10_2304, i_10_2323, i_10_2349, i_10_2350, i_10_2365, i_10_2376, i_10_2406, i_10_2409, i_10_2472, i_10_2473, i_10_2563, i_10_2604, i_10_2629, i_10_2632, i_10_2657, i_10_2658, i_10_2662, i_10_2676, i_10_2700, i_10_2705, i_10_2734, i_10_2740, i_10_2754, i_10_2982, i_10_3034, i_10_3037, i_10_3070, i_10_3195, i_10_3196, i_10_3283, i_10_3294, i_10_3312, i_10_3384, i_10_3385, i_10_3387, i_10_3391, i_10_3432, i_10_3465, i_10_3469, i_10_3499, i_10_3585, i_10_3609, i_10_3616, i_10_3645, i_10_3651, i_10_3877, i_10_3996, i_10_4000, i_10_4113, i_10_4114, i_10_4115, i_10_4188, i_10_4275, i_10_4287, i_10_4297, i_10_4369, i_10_4554, i_10_4581, o_10_184);
	kernel_10_185 k_10_185(i_10_32, i_10_174, i_10_223, i_10_224, i_10_245, i_10_319, i_10_320, i_10_361, i_10_393, i_10_443, i_10_460, i_10_461, i_10_463, i_10_467, i_10_499, i_10_514, i_10_931, i_10_996, i_10_999, i_10_1237, i_10_1245, i_10_1246, i_10_1249, i_10_1297, i_10_1399, i_10_1432, i_10_1434, i_10_1435, i_10_1502, i_10_1543, i_10_1580, i_10_1624, i_10_1625, i_10_1689, i_10_1690, i_10_1807, i_10_1818, i_10_1819, i_10_1912, i_10_1983, i_10_1994, i_10_1996, i_10_2003, i_10_2006, i_10_2337, i_10_2353, i_10_2450, i_10_2474, i_10_2556, i_10_2629, i_10_2631, i_10_2634, i_10_2642, i_10_2705, i_10_2731, i_10_2733, i_10_2734, i_10_2735, i_10_2786, i_10_3041, i_10_3157, i_10_3284, i_10_3313, i_10_3316, i_10_3333, i_10_3387, i_10_3434, i_10_3451, i_10_3470, i_10_3473, i_10_3500, i_10_3525, i_10_3526, i_10_3543, i_10_3544, i_10_3725, i_10_3834, i_10_3835, i_10_3838, i_10_3839, i_10_3841, i_10_3852, i_10_3855, i_10_3883, i_10_3884, i_10_3895, i_10_3896, i_10_3988, i_10_4054, i_10_4055, i_10_4115, i_10_4121, i_10_4207, i_10_4208, i_10_4211, i_10_4282, i_10_4292, i_10_4588, i_10_4589, i_10_4592, o_10_185);
	kernel_10_186 k_10_186(i_10_46, i_10_47, i_10_49, i_10_50, i_10_154, i_10_179, i_10_220, i_10_221, i_10_222, i_10_280, i_10_291, i_10_318, i_10_327, i_10_328, i_10_406, i_10_410, i_10_440, i_10_445, i_10_795, i_10_798, i_10_893, i_10_1028, i_10_1037, i_10_1118, i_10_1121, i_10_1202, i_10_1239, i_10_1242, i_10_1264, i_10_1266, i_10_1276, i_10_1306, i_10_1445, i_10_1539, i_10_1653, i_10_1683, i_10_1685, i_10_1691, i_10_1765, i_10_1767, i_10_1768, i_10_1769, i_10_1771, i_10_1772, i_10_1819, i_10_1822, i_10_2201, i_10_2327, i_10_2361, i_10_2362, i_10_2378, i_10_2381, i_10_2449, i_10_2460, i_10_2603, i_10_2607, i_10_2629, i_10_2631, i_10_2635, i_10_2718, i_10_2723, i_10_2826, i_10_2829, i_10_2831, i_10_2834, i_10_2917, i_10_2918, i_10_2919, i_10_2921, i_10_2923, i_10_2924, i_10_2980, i_10_3048, i_10_3070, i_10_3072, i_10_3091, i_10_3092, i_10_3283, i_10_3388, i_10_3403, i_10_3407, i_10_3523, i_10_3551, i_10_3614, i_10_3809, i_10_3837, i_10_3846, i_10_3850, i_10_3852, i_10_3853, i_10_3855, i_10_3856, i_10_3857, i_10_4123, i_10_4284, i_10_4286, i_10_4288, i_10_4564, i_10_4570, i_10_4571, o_10_186);
	kernel_10_187 k_10_187(i_10_144, i_10_147, i_10_148, i_10_172, i_10_177, i_10_222, i_10_223, i_10_250, i_10_260, i_10_266, i_10_293, i_10_330, i_10_405, i_10_408, i_10_411, i_10_447, i_10_628, i_10_629, i_10_687, i_10_741, i_10_742, i_10_745, i_10_747, i_10_798, i_10_967, i_10_970, i_10_1002, i_10_1218, i_10_1221, i_10_1222, i_10_1236, i_10_1239, i_10_1240, i_10_1275, i_10_1365, i_10_1434, i_10_1438, i_10_1444, i_10_1446, i_10_1447, i_10_1488, i_10_1502, i_10_1821, i_10_1920, i_10_2001, i_10_2031, i_10_2032, i_10_2037, i_10_2040, i_10_2110, i_10_2290, i_10_2349, i_10_2353, i_10_2354, i_10_2383, i_10_2384, i_10_2406, i_10_2470, i_10_2559, i_10_2608, i_10_2711, i_10_2715, i_10_2734, i_10_2742, i_10_2787, i_10_2841, i_10_2847, i_10_2885, i_10_2960, i_10_2967, i_10_3076, i_10_3077, i_10_3273, i_10_3283, i_10_3319, i_10_3384, i_10_3387, i_10_3492, i_10_3504, i_10_3507, i_10_3508, i_10_3544, i_10_3718, i_10_3721, i_10_3836, i_10_3840, i_10_4012, i_10_4119, i_10_4129, i_10_4211, i_10_4220, i_10_4266, i_10_4269, i_10_4272, i_10_4281, i_10_4292, i_10_4435, i_10_4564, i_10_4567, i_10_4585, o_10_187);
	kernel_10_188 k_10_188(i_10_172, i_10_177, i_10_183, i_10_249, i_10_267, i_10_285, i_10_286, i_10_319, i_10_324, i_10_328, i_10_408, i_10_410, i_10_460, i_10_507, i_10_753, i_10_754, i_10_797, i_10_996, i_10_1006, i_10_1041, i_10_1042, i_10_1309, i_10_1437, i_10_1442, i_10_1578, i_10_1579, i_10_1654, i_10_1655, i_10_1684, i_10_1687, i_10_1690, i_10_1815, i_10_1821, i_10_1823, i_10_1825, i_10_1947, i_10_1951, i_10_1996, i_10_2019, i_10_2022, i_10_2349, i_10_2350, i_10_2352, i_10_2353, i_10_2355, i_10_2451, i_10_2453, i_10_2469, i_10_2607, i_10_2632, i_10_2633, i_10_2673, i_10_2703, i_10_2704, i_10_2713, i_10_2715, i_10_2729, i_10_2734, i_10_2735, i_10_2823, i_10_2829, i_10_2985, i_10_2986, i_10_3076, i_10_3270, i_10_3271, i_10_3272, i_10_3274, i_10_3388, i_10_3391, i_10_3409, i_10_3469, i_10_3472, i_10_3525, i_10_3582, i_10_3588, i_10_3589, i_10_3612, i_10_3613, i_10_3780, i_10_3837, i_10_3841, i_10_3852, i_10_3855, i_10_3857, i_10_3858, i_10_3894, i_10_3895, i_10_3990, i_10_3991, i_10_4116, i_10_4127, i_10_4129, i_10_4267, i_10_4281, i_10_4282, i_10_4283, i_10_4288, i_10_4290, i_10_4567, o_10_188);
	kernel_10_189 k_10_189(i_10_172, i_10_173, i_10_219, i_10_222, i_10_224, i_10_271, i_10_279, i_10_286, i_10_315, i_10_316, i_10_318, i_10_319, i_10_320, i_10_408, i_10_442, i_10_463, i_10_464, i_10_467, i_10_716, i_10_900, i_10_967, i_10_1084, i_10_1245, i_10_1246, i_10_1247, i_10_1248, i_10_1249, i_10_1250, i_10_1305, i_10_1307, i_10_1308, i_10_1311, i_10_1365, i_10_1651, i_10_1652, i_10_1653, i_10_1678, i_10_1685, i_10_1687, i_10_1802, i_10_1822, i_10_1825, i_10_1911, i_10_1912, i_10_1913, i_10_2198, i_10_2355, i_10_2403, i_10_2452, i_10_2460, i_10_2506, i_10_2628, i_10_2629, i_10_2632, i_10_2636, i_10_2701, i_10_2721, i_10_2722, i_10_2724, i_10_2725, i_10_2726, i_10_2731, i_10_2782, i_10_2828, i_10_2829, i_10_2833, i_10_2916, i_10_2919, i_10_2920, i_10_2922, i_10_2923, i_10_3034, i_10_3163, i_10_3195, i_10_3284, i_10_3323, i_10_3325, i_10_3390, i_10_3391, i_10_3402, i_10_3403, i_10_3586, i_10_3855, i_10_3856, i_10_3858, i_10_3860, i_10_3979, i_10_3980, i_10_3982, i_10_3983, i_10_3986, i_10_4117, i_10_4279, i_10_4285, i_10_4286, i_10_4287, i_10_4288, i_10_4290, i_10_4291, i_10_4566, o_10_189);
	kernel_10_190 k_10_190(i_10_14, i_10_49, i_10_86, i_10_176, i_10_179, i_10_221, i_10_254, i_10_283, i_10_287, i_10_317, i_10_391, i_10_464, i_10_509, i_10_689, i_10_869, i_10_1084, i_10_1085, i_10_1088, i_10_1103, i_10_1235, i_10_1237, i_10_1238, i_10_1271, i_10_1298, i_10_1301, i_10_1439, i_10_1454, i_10_1541, i_10_1544, i_10_1583, i_10_1622, i_10_1648, i_10_1651, i_10_1684, i_10_1685, i_10_1687, i_10_1688, i_10_1981, i_10_1982, i_10_1990, i_10_1994, i_10_2003, i_10_2020, i_10_2021, i_10_2030, i_10_2189, i_10_2201, i_10_2204, i_10_2351, i_10_2356, i_10_2465, i_10_2468, i_10_2471, i_10_2473, i_10_2479, i_10_2567, i_10_2629, i_10_2636, i_10_2650, i_10_2651, i_10_2654, i_10_2660, i_10_2711, i_10_2714, i_10_2821, i_10_2830, i_10_2831, i_10_2846, i_10_2917, i_10_2919, i_10_2924, i_10_2966, i_10_2969, i_10_3043, i_10_3070, i_10_3073, i_10_3088, i_10_3197, i_10_3323, i_10_3391, i_10_3503, i_10_3526, i_10_3584, i_10_3733, i_10_3734, i_10_3786, i_10_3794, i_10_3835, i_10_3847, i_10_3979, i_10_4028, i_10_4126, i_10_4127, i_10_4130, i_10_4154, i_10_4172, i_10_4175, i_10_4279, i_10_4291, i_10_4565, o_10_190);
	kernel_10_191 k_10_191(i_10_87, i_10_152, i_10_172, i_10_176, i_10_221, i_10_224, i_10_259, i_10_260, i_10_325, i_10_433, i_10_443, i_10_445, i_10_446, i_10_448, i_10_449, i_10_454, i_10_461, i_10_463, i_10_467, i_10_716, i_10_794, i_10_797, i_10_800, i_10_899, i_10_904, i_10_905, i_10_908, i_10_965, i_10_971, i_10_999, i_10_1000, i_10_1135, i_10_1165, i_10_1166, i_10_1237, i_10_1240, i_10_1244, i_10_1245, i_10_1246, i_10_1247, i_10_1248, i_10_1308, i_10_1311, i_10_1553, i_10_1818, i_10_1822, i_10_1823, i_10_2181, i_10_2249, i_10_2309, i_10_2335, i_10_2355, i_10_2410, i_10_2450, i_10_2453, i_10_2470, i_10_2630, i_10_2635, i_10_2662, i_10_2663, i_10_2700, i_10_2713, i_10_2720, i_10_2728, i_10_2729, i_10_2731, i_10_2735, i_10_2785, i_10_2824, i_10_2881, i_10_2884, i_10_2917, i_10_2919, i_10_2920, i_10_3038, i_10_3073, i_10_3274, i_10_3334, i_10_3387, i_10_3391, i_10_3493, i_10_3494, i_10_3541, i_10_3649, i_10_3788, i_10_3836, i_10_3858, i_10_3859, i_10_3986, i_10_4120, i_10_4121, i_10_4220, i_10_4270, i_10_4271, i_10_4274, i_10_4291, i_10_4292, i_10_4564, i_10_4565, i_10_4571, o_10_191);
	kernel_10_192 k_10_192(i_10_217, i_10_223, i_10_224, i_10_245, i_10_280, i_10_281, i_10_283, i_10_284, i_10_316, i_10_318, i_10_319, i_10_413, i_10_435, i_10_443, i_10_460, i_10_748, i_10_749, i_10_792, i_10_793, i_10_795, i_10_898, i_10_956, i_10_1026, i_10_1027, i_10_1028, i_10_1033, i_10_1137, i_10_1139, i_10_1233, i_10_1234, i_10_1243, i_10_1539, i_10_1541, i_10_1549, i_10_1651, i_10_1654, i_10_1683, i_10_1684, i_10_1685, i_10_1686, i_10_1687, i_10_1688, i_10_1689, i_10_1691, i_10_1818, i_10_1819, i_10_1820, i_10_1821, i_10_1826, i_10_1913, i_10_2180, i_10_2243, i_10_2352, i_10_2358, i_10_2452, i_10_2470, i_10_2628, i_10_2631, i_10_2674, i_10_2675, i_10_2677, i_10_2701, i_10_2702, i_10_2710, i_10_2718, i_10_2728, i_10_2983, i_10_3073, i_10_3195, i_10_3198, i_10_3199, i_10_3203, i_10_3322, i_10_3407, i_10_3408, i_10_3409, i_10_3519, i_10_3585, i_10_3588, i_10_3589, i_10_3609, i_10_3610, i_10_3612, i_10_3614, i_10_3781, i_10_3784, i_10_3785, i_10_3786, i_10_3787, i_10_3837, i_10_3855, i_10_3856, i_10_3857, i_10_3979, i_10_3980, i_10_3987, i_10_4113, i_10_4287, i_10_4567, i_10_4568, o_10_192);
	kernel_10_193 k_10_193(i_10_89, i_10_219, i_10_220, i_10_224, i_10_286, i_10_388, i_10_405, i_10_410, i_10_445, i_10_511, i_10_519, i_10_628, i_10_696, i_10_697, i_10_698, i_10_797, i_10_799, i_10_846, i_10_850, i_10_853, i_10_949, i_10_963, i_10_976, i_10_1060, i_10_1124, i_10_1237, i_10_1247, i_10_1249, i_10_1250, i_10_1308, i_10_1478, i_10_1651, i_10_1652, i_10_1688, i_10_1691, i_10_1711, i_10_1755, i_10_1776, i_10_1819, i_10_1820, i_10_1821, i_10_1823, i_10_1826, i_10_1913, i_10_1952, i_10_2020, i_10_2083, i_10_2272, i_10_2381, i_10_2382, i_10_2514, i_10_2517, i_10_2518, i_10_2533, i_10_2543, i_10_2563, i_10_2635, i_10_2653, i_10_2654, i_10_2722, i_10_2724, i_10_2732, i_10_2758, i_10_2820, i_10_2830, i_10_2833, i_10_2918, i_10_3049, i_10_3118, i_10_3165, i_10_3166, i_10_3198, i_10_3200, i_10_3273, i_10_3275, i_10_3358, i_10_3388, i_10_3392, i_10_3407, i_10_3409, i_10_3410, i_10_3544, i_10_3640, i_10_3705, i_10_3706, i_10_3732, i_10_3832, i_10_3838, i_10_3840, i_10_3851, i_10_3860, i_10_3905, i_10_3978, i_10_3979, i_10_4129, i_10_4184, i_10_4288, i_10_4460, i_10_4480, i_10_4570, o_10_193);
	kernel_10_194 k_10_194(i_10_28, i_10_118, i_10_119, i_10_122, i_10_220, i_10_221, i_10_250, i_10_281, i_10_284, i_10_316, i_10_329, i_10_388, i_10_431, i_10_433, i_10_437, i_10_460, i_10_520, i_10_749, i_10_754, i_10_793, i_10_794, i_10_797, i_10_968, i_10_990, i_10_1000, i_10_1236, i_10_1240, i_10_1241, i_10_1261, i_10_1308, i_10_1309, i_10_1578, i_10_1647, i_10_1650, i_10_1651, i_10_1652, i_10_1686, i_10_1687, i_10_1732, i_10_1821, i_10_1822, i_10_1912, i_10_1944, i_10_2186, i_10_2242, i_10_2350, i_10_2352, i_10_2354, i_10_2355, i_10_2357, i_10_2467, i_10_2473, i_10_2632, i_10_2633, i_10_2658, i_10_2660, i_10_2701, i_10_2732, i_10_2788, i_10_2827, i_10_2832, i_10_2886, i_10_2888, i_10_2922, i_10_3036, i_10_3037, i_10_3038, i_10_3046, i_10_3049, i_10_3075, i_10_3076, i_10_3088, i_10_3198, i_10_3199, i_10_3276, i_10_3390, i_10_3391, i_10_3406, i_10_3466, i_10_3587, i_10_3609, i_10_3649, i_10_3650, i_10_3653, i_10_3782, i_10_3785, i_10_3788, i_10_3855, i_10_3856, i_10_3893, i_10_3979, i_10_3980, i_10_4114, i_10_4115, i_10_4117, i_10_4127, i_10_4270, i_10_4288, i_10_4289, i_10_4567, o_10_194);
	kernel_10_195 k_10_195(i_10_45, i_10_144, i_10_219, i_10_280, i_10_283, i_10_287, i_10_316, i_10_320, i_10_328, i_10_390, i_10_392, i_10_437, i_10_440, i_10_442, i_10_463, i_10_464, i_10_711, i_10_712, i_10_821, i_10_1234, i_10_1240, i_10_1241, i_10_1245, i_10_1246, i_10_1298, i_10_1363, i_10_1433, i_10_1441, i_10_1445, i_10_1551, i_10_1552, i_10_1553, i_10_1580, i_10_1622, i_10_1649, i_10_1655, i_10_1683, i_10_1684, i_10_1686, i_10_1687, i_10_1769, i_10_1943, i_10_1952, i_10_1982, i_10_2003, i_10_2185, i_10_2312, i_10_2349, i_10_2358, i_10_2361, i_10_2362, i_10_2448, i_10_2449, i_10_2450, i_10_2456, i_10_2468, i_10_2473, i_10_2516, i_10_2593, i_10_2629, i_10_2630, i_10_2631, i_10_2632, i_10_2638, i_10_2655, i_10_2658, i_10_2660, i_10_2661, i_10_2718, i_10_2720, i_10_2723, i_10_2728, i_10_2781, i_10_2818, i_10_2887, i_10_2963, i_10_3071, i_10_3231, i_10_3388, i_10_3389, i_10_3469, i_10_3540, i_10_3583, i_10_3586, i_10_3587, i_10_3650, i_10_3784, i_10_3835, i_10_3838, i_10_3839, i_10_3884, i_10_3910, i_10_4028, i_10_4119, i_10_4124, i_10_4127, i_10_4142, i_10_4145, i_10_4266, i_10_4289, o_10_195);
	kernel_10_196 k_10_196(i_10_83, i_10_283, i_10_284, i_10_289, i_10_325, i_10_442, i_10_446, i_10_461, i_10_464, i_10_504, i_10_508, i_10_514, i_10_545, i_10_892, i_10_893, i_10_1027, i_10_1028, i_10_1135, i_10_1139, i_10_1233, i_10_1234, i_10_1236, i_10_1238, i_10_1243, i_10_1244, i_10_1264, i_10_1306, i_10_1313, i_10_1650, i_10_1652, i_10_1690, i_10_1818, i_10_1819, i_10_1823, i_10_1909, i_10_1910, i_10_1912, i_10_1913, i_10_1989, i_10_1990, i_10_1991, i_10_2017, i_10_2198, i_10_2353, i_10_2358, i_10_2359, i_10_2360, i_10_2361, i_10_2362, i_10_2408, i_10_2449, i_10_2457, i_10_2458, i_10_2459, i_10_2462, i_10_2470, i_10_2601, i_10_2700, i_10_2709, i_10_2728, i_10_2818, i_10_2828, i_10_2830, i_10_2882, i_10_2918, i_10_2920, i_10_2921, i_10_3150, i_10_3269, i_10_3272, i_10_3277, i_10_3386, i_10_3388, i_10_3389, i_10_3402, i_10_3406, i_10_3523, i_10_3587, i_10_3722, i_10_3783, i_10_3784, i_10_3785, i_10_3787, i_10_3830, i_10_3834, i_10_3848, i_10_3849, i_10_3850, i_10_3854, i_10_3855, i_10_3856, i_10_3857, i_10_3890, i_10_3892, i_10_3982, i_10_3986, i_10_4024, i_10_4233, i_10_4565, i_10_4567, o_10_196);
	kernel_10_197 k_10_197(i_10_89, i_10_177, i_10_214, i_10_259, i_10_325, i_10_329, i_10_370, i_10_446, i_10_518, i_10_543, i_10_738, i_10_793, i_10_797, i_10_799, i_10_827, i_10_963, i_10_967, i_10_999, i_10_1083, i_10_1087, i_10_1120, i_10_1205, i_10_1237, i_10_1245, i_10_1248, i_10_1306, i_10_1312, i_10_1313, i_10_1344, i_10_1542, i_10_1553, i_10_1647, i_10_1650, i_10_1685, i_10_1689, i_10_1690, i_10_1818, i_10_2019, i_10_2182, i_10_2338, i_10_2350, i_10_2378, i_10_2404, i_10_2407, i_10_2451, i_10_2472, i_10_2629, i_10_2631, i_10_2632, i_10_2636, i_10_2707, i_10_2713, i_10_2714, i_10_2718, i_10_2727, i_10_2731, i_10_2781, i_10_2823, i_10_2824, i_10_2828, i_10_2832, i_10_2850, i_10_2868, i_10_2887, i_10_2922, i_10_2954, i_10_2957, i_10_2983, i_10_3037, i_10_3038, i_10_3092, i_10_3268, i_10_3274, i_10_3280, i_10_3328, i_10_3388, i_10_3405, i_10_3432, i_10_3444, i_10_3447, i_10_3526, i_10_3583, i_10_3589, i_10_3612, i_10_3613, i_10_3616, i_10_3672, i_10_3687, i_10_3813, i_10_3841, i_10_3843, i_10_3844, i_10_3946, i_10_4156, i_10_4157, i_10_4175, i_10_4215, i_10_4272, i_10_4273, i_10_4565, o_10_197);
	kernel_10_198 k_10_198(i_10_24, i_10_64, i_10_67, i_10_70, i_10_175, i_10_183, i_10_272, i_10_283, i_10_319, i_10_408, i_10_410, i_10_434, i_10_458, i_10_536, i_10_817, i_10_905, i_10_906, i_10_947, i_10_951, i_10_956, i_10_1064, i_10_1119, i_10_1172, i_10_1286, i_10_1375, i_10_1445, i_10_1482, i_10_1484, i_10_1551, i_10_1554, i_10_1632, i_10_1641, i_10_1647, i_10_1684, i_10_1790, i_10_1819, i_10_1822, i_10_1887, i_10_1911, i_10_1912, i_10_1915, i_10_1916, i_10_1918, i_10_1919, i_10_1932, i_10_1933, i_10_2027, i_10_2059, i_10_2063, i_10_2094, i_10_2095, i_10_2154, i_10_2157, i_10_2158, i_10_2274, i_10_2275, i_10_2311, i_10_2312, i_10_2337, i_10_2351, i_10_2352, i_10_2353, i_10_2354, i_10_2357, i_10_2452, i_10_2453, i_10_2508, i_10_2509, i_10_2541, i_10_2557, i_10_2605, i_10_2635, i_10_2640, i_10_2663, i_10_2698, i_10_2770, i_10_2820, i_10_2848, i_10_2856, i_10_2857, i_10_2919, i_10_2922, i_10_3031, i_10_3032, i_10_3074, i_10_3102, i_10_3103, i_10_3104, i_10_3229, i_10_3545, i_10_3610, i_10_3647, i_10_3775, i_10_3805, i_10_3806, i_10_3859, i_10_3982, i_10_4126, i_10_4364, i_10_4534, o_10_198);
	kernel_10_199 k_10_199(i_10_27, i_10_124, i_10_175, i_10_285, i_10_369, i_10_433, i_10_443, i_10_444, i_10_467, i_10_501, i_10_532, i_10_729, i_10_730, i_10_732, i_10_733, i_10_901, i_10_961, i_10_999, i_10_1052, i_10_1201, i_10_1263, i_10_1265, i_10_1270, i_10_1271, i_10_1308, i_10_1309, i_10_1353, i_10_1361, i_10_1363, i_10_1638, i_10_1741, i_10_1765, i_10_1823, i_10_1912, i_10_1947, i_10_1948, i_10_1957, i_10_2079, i_10_2151, i_10_2166, i_10_2167, i_10_2304, i_10_2306, i_10_2307, i_10_2310, i_10_2333, i_10_2335, i_10_2357, i_10_2436, i_10_2475, i_10_2478, i_10_2511, i_10_2608, i_10_2614, i_10_2615, i_10_2628, i_10_2630, i_10_2638, i_10_2655, i_10_2658, i_10_2659, i_10_2700, i_10_2832, i_10_2871, i_10_2881, i_10_2916, i_10_2920, i_10_2923, i_10_2952, i_10_2953, i_10_3037, i_10_3038, i_10_3040, i_10_3055, i_10_3087, i_10_3204, i_10_3229, i_10_3356, i_10_3358, i_10_3560, i_10_3651, i_10_3682, i_10_3683, i_10_3684, i_10_3685, i_10_3774, i_10_3853, i_10_3889, i_10_3892, i_10_3894, i_10_3924, i_10_3984, i_10_4124, i_10_4192, i_10_4230, i_10_4231, i_10_4374, i_10_4375, i_10_4376, i_10_4580, o_10_199);
	kernel_10_200 k_10_200(i_10_33, i_10_123, i_10_174, i_10_177, i_10_260, i_10_286, i_10_319, i_10_328, i_10_408, i_10_412, i_10_438, i_10_439, i_10_440, i_10_511, i_10_512, i_10_796, i_10_967, i_10_1003, i_10_1236, i_10_1239, i_10_1311, i_10_1439, i_10_1546, i_10_1619, i_10_1626, i_10_1627, i_10_1686, i_10_1689, i_10_1690, i_10_1691, i_10_1821, i_10_1822, i_10_1823, i_10_1986, i_10_1996, i_10_2031, i_10_2032, i_10_2361, i_10_2364, i_10_2407, i_10_2410, i_10_2451, i_10_2452, i_10_2455, i_10_2472, i_10_2473, i_10_2605, i_10_2634, i_10_2635, i_10_2636, i_10_2663, i_10_2704, i_10_2706, i_10_2713, i_10_2716, i_10_2717, i_10_2722, i_10_2733, i_10_2734, i_10_2788, i_10_2826, i_10_2827, i_10_2829, i_10_2830, i_10_2831, i_10_2833, i_10_2883, i_10_2884, i_10_2885, i_10_2985, i_10_2986, i_10_3049, i_10_3151, i_10_3202, i_10_3280, i_10_3283, i_10_3318, i_10_3325, i_10_3328, i_10_3391, i_10_3403, i_10_3525, i_10_3585, i_10_3615, i_10_3616, i_10_3617, i_10_3649, i_10_3653, i_10_3783, i_10_3786, i_10_3834, i_10_3835, i_10_3856, i_10_3858, i_10_3859, i_10_3912, i_10_3913, i_10_4281, i_10_4289, i_10_4571, o_10_200);
	kernel_10_201 k_10_201(i_10_24, i_10_33, i_10_184, i_10_283, i_10_320, i_10_323, i_10_330, i_10_332, i_10_393, i_10_394, i_10_436, i_10_440, i_10_444, i_10_461, i_10_500, i_10_503, i_10_696, i_10_732, i_10_733, i_10_734, i_10_931, i_10_952, i_10_1002, i_10_1043, i_10_1047, i_10_1348, i_10_1349, i_10_1482, i_10_1488, i_10_1528, i_10_1548, i_10_1551, i_10_1555, i_10_1556, i_10_1655, i_10_1686, i_10_1767, i_10_1768, i_10_1823, i_10_1869, i_10_1957, i_10_2003, i_10_2004, i_10_2029, i_10_2083, i_10_2088, i_10_2156, i_10_2186, i_10_2204, i_10_2212, i_10_2312, i_10_2382, i_10_2409, i_10_2453, i_10_2571, i_10_2631, i_10_2632, i_10_2636, i_10_2659, i_10_2721, i_10_2722, i_10_2761, i_10_2806, i_10_2917, i_10_2923, i_10_2956, i_10_2983, i_10_2987, i_10_3030, i_10_3041, i_10_3131, i_10_3275, i_10_3361, i_10_3362, i_10_3388, i_10_3537, i_10_3538, i_10_3554, i_10_3588, i_10_3605, i_10_3608, i_10_3612, i_10_3615, i_10_3616, i_10_3837, i_10_3856, i_10_3865, i_10_3981, i_10_3982, i_10_3984, i_10_3990, i_10_3991, i_10_3993, i_10_4287, i_10_4288, i_10_4289, i_10_4292, i_10_4372, i_10_4570, i_10_4571, o_10_201);
	kernel_10_202 k_10_202(i_10_42, i_10_177, i_10_220, i_10_222, i_10_246, i_10_247, i_10_249, i_10_250, i_10_283, i_10_292, i_10_442, i_10_463, i_10_466, i_10_467, i_10_566, i_10_597, i_10_894, i_10_996, i_10_1032, i_10_1033, i_10_1141, i_10_1239, i_10_1241, i_10_1266, i_10_1444, i_10_1545, i_10_1578, i_10_1648, i_10_1653, i_10_1654, i_10_1825, i_10_2004, i_10_2019, i_10_2022, i_10_2351, i_10_2353, i_10_2359, i_10_2361, i_10_2364, i_10_2469, i_10_2470, i_10_2471, i_10_2472, i_10_2473, i_10_2604, i_10_2607, i_10_2632, i_10_2657, i_10_2658, i_10_2703, i_10_2704, i_10_2706, i_10_2721, i_10_2727, i_10_2731, i_10_2781, i_10_2826, i_10_2833, i_10_2917, i_10_3033, i_10_3043, i_10_3045, i_10_3072, i_10_3075, i_10_3158, i_10_3162, i_10_3267, i_10_3270, i_10_3278, i_10_3279, i_10_3280, i_10_3388, i_10_3406, i_10_3430, i_10_3493, i_10_3652, i_10_3684, i_10_3687, i_10_3782, i_10_3787, i_10_3810, i_10_3811, i_10_3813, i_10_3839, i_10_3846, i_10_3855, i_10_3858, i_10_4116, i_10_4117, i_10_4119, i_10_4125, i_10_4128, i_10_4129, i_10_4215, i_10_4218, i_10_4289, i_10_4291, i_10_4292, i_10_4564, i_10_4567, o_10_202);
	kernel_10_203 k_10_203(i_10_34, i_10_176, i_10_221, i_10_254, i_10_280, i_10_328, i_10_374, i_10_394, i_10_445, i_10_446, i_10_715, i_10_718, i_10_754, i_10_792, i_10_797, i_10_798, i_10_829, i_10_830, i_10_832, i_10_957, i_10_959, i_10_1012, i_10_1031, i_10_1119, i_10_1234, i_10_1235, i_10_1313, i_10_1544, i_10_1578, i_10_1579, i_10_1683, i_10_1687, i_10_1814, i_10_1819, i_10_1820, i_10_1823, i_10_1919, i_10_1939, i_10_2026, i_10_2178, i_10_2179, i_10_2309, i_10_2311, i_10_2350, i_10_2353, i_10_2354, i_10_2365, i_10_2380, i_10_2404, i_10_2569, i_10_2708, i_10_2721, i_10_2722, i_10_2731, i_10_2783, i_10_2785, i_10_2834, i_10_3011, i_10_3099, i_10_3200, i_10_3202, i_10_3236, i_10_3239, i_10_3275, i_10_3298, i_10_3352, i_10_3386, i_10_3389, i_10_3493, i_10_3494, i_10_3542, i_10_3581, i_10_3583, i_10_3584, i_10_3615, i_10_3616, i_10_3617, i_10_3636, i_10_3650, i_10_3653, i_10_3711, i_10_3724, i_10_3781, i_10_3782, i_10_3783, i_10_3784, i_10_3785, i_10_3786, i_10_3787, i_10_3788, i_10_3809, i_10_3860, i_10_3947, i_10_4024, i_10_4118, i_10_4120, i_10_4121, i_10_4130, i_10_4175, i_10_4214, o_10_203);
	kernel_10_204 k_10_204(i_10_17, i_10_68, i_10_134, i_10_152, i_10_170, i_10_223, i_10_239, i_10_275, i_10_331, i_10_373, i_10_376, i_10_392, i_10_440, i_10_445, i_10_446, i_10_447, i_10_462, i_10_518, i_10_548, i_10_637, i_10_718, i_10_719, i_10_737, i_10_799, i_10_950, i_10_989, i_10_1166, i_10_1245, i_10_1246, i_10_1267, i_10_1312, i_10_1313, i_10_1438, i_10_1491, i_10_1493, i_10_1538, i_10_1539, i_10_1583, i_10_1616, i_10_1637, i_10_1643, i_10_1646, i_10_1651, i_10_1653, i_10_1691, i_10_1824, i_10_1873, i_10_1940, i_10_1942, i_10_1951, i_10_1961, i_10_2032, i_10_2069, i_10_2183, i_10_2231, i_10_2326, i_10_2330, i_10_2359, i_10_2452, i_10_2474, i_10_2521, i_10_2535, i_10_2636, i_10_2663, i_10_2672, i_10_2705, i_10_2865, i_10_2883, i_10_2884, i_10_2986, i_10_2987, i_10_3072, i_10_3075, i_10_3122, i_10_3195, i_10_3199, i_10_3356, i_10_3455, i_10_3469, i_10_3495, i_10_3509, i_10_3590, i_10_3617, i_10_3650, i_10_3788, i_10_3801, i_10_3804, i_10_3860, i_10_3877, i_10_3878, i_10_3910, i_10_3950, i_10_3991, i_10_3994, i_10_3995, i_10_4138, i_10_4154, i_10_4183, i_10_4288, i_10_4291, o_10_204);
	kernel_10_205 k_10_205(i_10_39, i_10_159, i_10_251, i_10_282, i_10_284, i_10_292, i_10_296, i_10_320, i_10_328, i_10_329, i_10_368, i_10_394, i_10_411, i_10_412, i_10_413, i_10_439, i_10_440, i_10_444, i_10_447, i_10_448, i_10_449, i_10_512, i_10_800, i_10_962, i_10_1015, i_10_1016, i_10_1034, i_10_1221, i_10_1222, i_10_1237, i_10_1346, i_10_1348, i_10_1687, i_10_1688, i_10_1690, i_10_1691, i_10_1729, i_10_1730, i_10_1733, i_10_1984, i_10_2003, i_10_2006, i_10_2030, i_10_2357, i_10_2383, i_10_2384, i_10_2450, i_10_2454, i_10_2455, i_10_2456, i_10_2464, i_10_2471, i_10_2512, i_10_2516, i_10_2536, i_10_2537, i_10_2571, i_10_2601, i_10_2604, i_10_2673, i_10_2676, i_10_2704, i_10_2714, i_10_2716, i_10_2717, i_10_2728, i_10_2734, i_10_2743, i_10_2788, i_10_2831, i_10_2833, i_10_2834, i_10_2885, i_10_2969, i_10_2980, i_10_3199, i_10_3278, i_10_3281, i_10_3301, i_10_3506, i_10_3551, i_10_3561, i_10_3562, i_10_3586, i_10_3587, i_10_3590, i_10_3613, i_10_3614, i_10_3616, i_10_3784, i_10_3787, i_10_3840, i_10_3913, i_10_3983, i_10_4120, i_10_4155, i_10_4277, i_10_4291, i_10_4292, i_10_4567, o_10_205);
	kernel_10_206 k_10_206(i_10_152, i_10_172, i_10_222, i_10_268, i_10_280, i_10_284, i_10_285, i_10_392, i_10_409, i_10_413, i_10_431, i_10_439, i_10_565, i_10_751, i_10_754, i_10_755, i_10_799, i_10_899, i_10_954, i_10_957, i_10_958, i_10_967, i_10_1032, i_10_1033, i_10_1236, i_10_1238, i_10_1242, i_10_1243, i_10_1244, i_10_1245, i_10_1249, i_10_1306, i_10_1345, i_10_1360, i_10_1366, i_10_1549, i_10_1683, i_10_1823, i_10_1825, i_10_1913, i_10_1916, i_10_1949, i_10_1952, i_10_1997, i_10_2311, i_10_2353, i_10_2364, i_10_2410, i_10_2450, i_10_2457, i_10_2470, i_10_2472, i_10_2474, i_10_2513, i_10_2705, i_10_2725, i_10_2735, i_10_2830, i_10_2834, i_10_2917, i_10_2919, i_10_2923, i_10_2924, i_10_2992, i_10_3037, i_10_3038, i_10_3039, i_10_3091, i_10_3199, i_10_3200, i_10_3270, i_10_3283, i_10_3388, i_10_3525, i_10_3563, i_10_3615, i_10_3617, i_10_3651, i_10_3780, i_10_3783, i_10_3784, i_10_3786, i_10_3787, i_10_3788, i_10_3844, i_10_3847, i_10_3854, i_10_3859, i_10_3982, i_10_3983, i_10_3986, i_10_3994, i_10_4116, i_10_4117, i_10_4118, i_10_4267, i_10_4273, i_10_4564, i_10_4571, i_10_4597, o_10_206);
	kernel_10_207 k_10_207(i_10_171, i_10_178, i_10_179, i_10_253, i_10_328, i_10_329, i_10_364, i_10_409, i_10_410, i_10_443, i_10_444, i_10_462, i_10_463, i_10_466, i_10_960, i_10_962, i_10_1032, i_10_1033, i_10_1034, i_10_1165, i_10_1233, i_10_1242, i_10_1296, i_10_1307, i_10_1431, i_10_1432, i_10_1443, i_10_1444, i_10_1539, i_10_1576, i_10_1683, i_10_1686, i_10_1728, i_10_1818, i_10_1819, i_10_2021, i_10_2223, i_10_2352, i_10_2359, i_10_2361, i_10_2364, i_10_2431, i_10_2442, i_10_2449, i_10_2450, i_10_2451, i_10_2454, i_10_2628, i_10_2629, i_10_2655, i_10_2658, i_10_2659, i_10_2661, i_10_2681, i_10_2701, i_10_2714, i_10_2727, i_10_2784, i_10_2862, i_10_2916, i_10_3038, i_10_3074, i_10_3267, i_10_3271, i_10_3277, i_10_3279, i_10_3280, i_10_3282, i_10_3316, i_10_3331, i_10_3349, i_10_3450, i_10_3497, i_10_3537, i_10_3538, i_10_3614, i_10_3617, i_10_3650, i_10_3786, i_10_3787, i_10_3834, i_10_3846, i_10_3854, i_10_4116, i_10_4119, i_10_4171, i_10_4172, i_10_4204, i_10_4219, i_10_4267, i_10_4269, i_10_4270, i_10_4279, i_10_4284, i_10_4285, i_10_4288, i_10_4428, i_10_4459, i_10_4582, i_10_4591, o_10_207);
	kernel_10_208 k_10_208(i_10_28, i_10_89, i_10_224, i_10_247, i_10_283, i_10_315, i_10_324, i_10_325, i_10_408, i_10_446, i_10_447, i_10_463, i_10_464, i_10_467, i_10_508, i_10_510, i_10_737, i_10_755, i_10_798, i_10_800, i_10_966, i_10_1027, i_10_1030, i_10_1034, i_10_1039, i_10_1140, i_10_1233, i_10_1234, i_10_1235, i_10_1238, i_10_1241, i_10_1307, i_10_1313, i_10_1363, i_10_1579, i_10_1650, i_10_1652, i_10_1820, i_10_1825, i_10_1910, i_10_1995, i_10_1996, i_10_2179, i_10_2186, i_10_2338, i_10_2382, i_10_2383, i_10_2384, i_10_2463, i_10_2464, i_10_2470, i_10_2474, i_10_2629, i_10_2661, i_10_2680, i_10_2706, i_10_2707, i_10_2714, i_10_2721, i_10_2730, i_10_2832, i_10_2833, i_10_2985, i_10_3039, i_10_3040, i_10_3049, i_10_3162, i_10_3165, i_10_3196, i_10_3197, i_10_3268, i_10_3270, i_10_3271, i_10_3321, i_10_3388, i_10_3389, i_10_3391, i_10_3402, i_10_3406, i_10_3468, i_10_3582, i_10_3609, i_10_3615, i_10_3785, i_10_3787, i_10_3834, i_10_3837, i_10_3846, i_10_3847, i_10_3889, i_10_3984, i_10_3985, i_10_4030, i_10_4031, i_10_4116, i_10_4128, i_10_4155, i_10_4217, i_10_4292, i_10_4567, o_10_208);
	kernel_10_209 k_10_209(i_10_197, i_10_202, i_10_273, i_10_274, i_10_276, i_10_277, i_10_279, i_10_293, i_10_392, i_10_408, i_10_447, i_10_509, i_10_515, i_10_792, i_10_959, i_10_985, i_10_1256, i_10_1322, i_10_1363, i_10_1394, i_10_1444, i_10_1462, i_10_1463, i_10_1484, i_10_1526, i_10_1552, i_10_1570, i_10_1573, i_10_1610, i_10_1643, i_10_1713, i_10_1716, i_10_1744, i_10_1764, i_10_1772, i_10_1820, i_10_1915, i_10_2005, i_10_2011, i_10_2019, i_10_2020, i_10_2022, i_10_2028, i_10_2182, i_10_2185, i_10_2186, i_10_2303, i_10_2327, i_10_2329, i_10_2330, i_10_2359, i_10_2434, i_10_2482, i_10_2483, i_10_2505, i_10_2506, i_10_2510, i_10_2634, i_10_2642, i_10_2675, i_10_2824, i_10_2874, i_10_2884, i_10_2965, i_10_2986, i_10_2987, i_10_3032, i_10_3039, i_10_3076, i_10_3320, i_10_3362, i_10_3364, i_10_3365, i_10_3431, i_10_3437, i_10_3496, i_10_3521, i_10_3717, i_10_3720, i_10_3806, i_10_3838, i_10_3841, i_10_3889, i_10_3890, i_10_3896, i_10_3920, i_10_3965, i_10_3982, i_10_3989, i_10_3992, i_10_4143, i_10_4144, i_10_4283, i_10_4360, i_10_4445, i_10_4526, i_10_4568, i_10_4574, i_10_4577, i_10_4596, o_10_209);
	kernel_10_210 k_10_210(i_10_175, i_10_283, i_10_284, i_10_285, i_10_286, i_10_289, i_10_318, i_10_325, i_10_390, i_10_425, i_10_460, i_10_463, i_10_464, i_10_514, i_10_639, i_10_752, i_10_892, i_10_893, i_10_965, i_10_967, i_10_990, i_10_1003, i_10_1026, i_10_1235, i_10_1241, i_10_1296, i_10_1305, i_10_1306, i_10_1307, i_10_1342, i_10_1542, i_10_1603, i_10_1629, i_10_1651, i_10_1652, i_10_1653, i_10_1655, i_10_1720, i_10_1721, i_10_1821, i_10_1822, i_10_1823, i_10_1909, i_10_1910, i_10_1916, i_10_1989, i_10_1990, i_10_2026, i_10_2288, i_10_2359, i_10_2361, i_10_2362, i_10_2377, i_10_2378, i_10_2566, i_10_2631, i_10_2656, i_10_2657, i_10_2675, i_10_2702, i_10_2710, i_10_2725, i_10_2726, i_10_2828, i_10_2918, i_10_2919, i_10_2980, i_10_3035, i_10_3069, i_10_3269, i_10_3384, i_10_3389, i_10_3403, i_10_3405, i_10_3555, i_10_3556, i_10_3582, i_10_3613, i_10_3615, i_10_3616, i_10_3617, i_10_3647, i_10_3683, i_10_3846, i_10_3848, i_10_3856, i_10_3888, i_10_3889, i_10_3980, i_10_4023, i_10_4096, i_10_4123, i_10_4125, i_10_4127, i_10_4214, i_10_4287, i_10_4288, i_10_4565, i_10_4567, i_10_4568, o_10_210);
	kernel_10_211 k_10_211(i_10_9, i_10_153, i_10_174, i_10_175, i_10_223, i_10_280, i_10_284, i_10_315, i_10_316, i_10_327, i_10_390, i_10_437, i_10_445, i_10_448, i_10_459, i_10_460, i_10_621, i_10_687, i_10_688, i_10_820, i_10_903, i_10_990, i_10_1030, i_10_1080, i_10_1083, i_10_1107, i_10_1215, i_10_1218, i_10_1236, i_10_1237, i_10_1239, i_10_1241, i_10_1264, i_10_1582, i_10_1800, i_10_1818, i_10_1826, i_10_1945, i_10_2016, i_10_2017, i_10_2026, i_10_2181, i_10_2199, i_10_2336, i_10_2352, i_10_2353, i_10_2355, i_10_2377, i_10_2378, i_10_2379, i_10_2406, i_10_2460, i_10_2466, i_10_2468, i_10_2471, i_10_2511, i_10_2514, i_10_2605, i_10_2611, i_10_2657, i_10_2700, i_10_2709, i_10_2718, i_10_2734, i_10_2783, i_10_2831, i_10_2881, i_10_3042, i_10_3069, i_10_3094, i_10_3392, i_10_3409, i_10_3468, i_10_3493, i_10_3610, i_10_3614, i_10_3616, i_10_3717, i_10_3720, i_10_3846, i_10_3855, i_10_3857, i_10_3894, i_10_3905, i_10_3906, i_10_3907, i_10_3909, i_10_4030, i_10_4122, i_10_4123, i_10_4168, i_10_4170, i_10_4176, i_10_4276, i_10_4291, i_10_4410, i_10_4566, i_10_4567, i_10_4568, i_10_4581, o_10_211);
	kernel_10_212 k_10_212(i_10_28, i_10_175, i_10_178, i_10_286, i_10_327, i_10_444, i_10_461, i_10_463, i_10_464, i_10_514, i_10_794, i_10_797, i_10_901, i_10_956, i_10_958, i_10_959, i_10_999, i_10_1000, i_10_1009, i_10_1162, i_10_1241, i_10_1306, i_10_1378, i_10_1379, i_10_1486, i_10_1576, i_10_1654, i_10_1655, i_10_1685, i_10_1687, i_10_1688, i_10_1813, i_10_1821, i_10_1944, i_10_1945, i_10_1946, i_10_2090, i_10_2183, i_10_2203, i_10_2305, i_10_2378, i_10_2448, i_10_2449, i_10_2450, i_10_2455, i_10_2456, i_10_2470, i_10_2471, i_10_2635, i_10_2636, i_10_2638, i_10_2639, i_10_2674, i_10_2711, i_10_2717, i_10_2720, i_10_2727, i_10_2728, i_10_3034, i_10_3035, i_10_3037, i_10_3042, i_10_3043, i_10_3046, i_10_3074, i_10_3087, i_10_3203, i_10_3267, i_10_3271, i_10_3278, i_10_3281, i_10_3384, i_10_3390, i_10_3392, i_10_3409, i_10_3431, i_10_3495, i_10_3539, i_10_3725, i_10_3781, i_10_3786, i_10_3837, i_10_3838, i_10_3857, i_10_3888, i_10_3890, i_10_3911, i_10_3979, i_10_3992, i_10_4055, i_10_4117, i_10_4118, i_10_4119, i_10_4121, i_10_4126, i_10_4280, i_10_4284, i_10_4370, i_10_4429, i_10_4583, o_10_212);
	kernel_10_213 k_10_213(i_10_64, i_10_176, i_10_177, i_10_178, i_10_183, i_10_214, i_10_262, i_10_284, i_10_316, i_10_521, i_10_757, i_10_758, i_10_794, i_10_798, i_10_799, i_10_907, i_10_994, i_10_1000, i_10_1012, i_10_1039, i_10_1058, i_10_1114, i_10_1300, i_10_1354, i_10_1355, i_10_1367, i_10_1434, i_10_1577, i_10_1579, i_10_1622, i_10_1625, i_10_1649, i_10_1651, i_10_1652, i_10_1684, i_10_1685, i_10_1689, i_10_1691, i_10_1730, i_10_1822, i_10_1919, i_10_1982, i_10_2027, i_10_2030, i_10_2153, i_10_2180, i_10_2201, i_10_2288, i_10_2360, i_10_2449, i_10_2506, i_10_2533, i_10_2566, i_10_2567, i_10_2570, i_10_2641, i_10_2663, i_10_2714, i_10_2719, i_10_2720, i_10_2728, i_10_2731, i_10_2826, i_10_2829, i_10_2849, i_10_2924, i_10_2963, i_10_3041, i_10_3044, i_10_3269, i_10_3280, i_10_3314, i_10_3316, i_10_3317, i_10_3387, i_10_3406, i_10_3461, i_10_3539, i_10_3560, i_10_3584, i_10_3689, i_10_3797, i_10_3834, i_10_3835, i_10_3839, i_10_3842, i_10_3849, i_10_3852, i_10_3894, i_10_3895, i_10_3982, i_10_4025, i_10_4028, i_10_4127, i_10_4172, i_10_4267, i_10_4283, i_10_4289, i_10_4583, i_10_4596, o_10_213);
	kernel_10_214 k_10_214(i_10_42, i_10_43, i_10_144, i_10_145, i_10_159, i_10_175, i_10_250, i_10_287, i_10_293, i_10_296, i_10_327, i_10_328, i_10_391, i_10_409, i_10_411, i_10_430, i_10_539, i_10_898, i_10_1084, i_10_1131, i_10_1132, i_10_1234, i_10_1237, i_10_1239, i_10_1241, i_10_1269, i_10_1270, i_10_1306, i_10_1307, i_10_1357, i_10_1362, i_10_1365, i_10_1444, i_10_1445, i_10_1447, i_10_1448, i_10_1651, i_10_1654, i_10_1680, i_10_1726, i_10_1816, i_10_1875, i_10_2019, i_10_2020, i_10_2022, i_10_2050, i_10_2253, i_10_2256, i_10_2257, i_10_2258, i_10_2259, i_10_2325, i_10_2354, i_10_2364, i_10_2454, i_10_2467, i_10_2514, i_10_2527, i_10_2546, i_10_2571, i_10_2660, i_10_2675, i_10_2787, i_10_2839, i_10_2913, i_10_2914, i_10_2979, i_10_3047, i_10_3237, i_10_3284, i_10_3291, i_10_3389, i_10_3399, i_10_3433, i_10_3495, i_10_3499, i_10_3583, i_10_3585, i_10_3586, i_10_3590, i_10_3687, i_10_3814, i_10_3837, i_10_3846, i_10_3855, i_10_3856, i_10_3873, i_10_3887, i_10_3945, i_10_3948, i_10_3973, i_10_4028, i_10_4055, i_10_4119, i_10_4123, i_10_4128, i_10_4220, i_10_4236, i_10_4267, i_10_4269, o_10_214);
	kernel_10_215 k_10_215(i_10_144, i_10_282, i_10_283, i_10_284, i_10_288, i_10_289, i_10_290, i_10_316, i_10_423, i_10_424, i_10_425, i_10_446, i_10_449, i_10_639, i_10_718, i_10_793, i_10_794, i_10_891, i_10_1003, i_10_1080, i_10_1083, i_10_1247, i_10_1262, i_10_1360, i_10_1440, i_10_1441, i_10_1442, i_10_1443, i_10_1444, i_10_1539, i_10_1543, i_10_1575, i_10_1576, i_10_1577, i_10_1579, i_10_1581, i_10_1653, i_10_1654, i_10_1679, i_10_1821, i_10_1822, i_10_1913, i_10_1945, i_10_1989, i_10_1990, i_10_2197, i_10_2200, i_10_2349, i_10_2351, i_10_2355, i_10_2362, i_10_2461, i_10_2659, i_10_2673, i_10_2674, i_10_2701, i_10_2709, i_10_2710, i_10_2711, i_10_2826, i_10_2881, i_10_2918, i_10_2920, i_10_3034, i_10_3038, i_10_3088, i_10_3196, i_10_3232, i_10_3267, i_10_3278, i_10_3294, i_10_3384, i_10_3405, i_10_3430, i_10_3431, i_10_3440, i_10_3522, i_10_3550, i_10_3584, i_10_3612, i_10_3614, i_10_3649, i_10_3781, i_10_3788, i_10_3835, i_10_3839, i_10_3859, i_10_3897, i_10_3910, i_10_3942, i_10_3990, i_10_3991, i_10_4051, i_10_4057, i_10_4119, i_10_4168, i_10_4276, i_10_4279, i_10_4565, i_10_4568, o_10_215);
	kernel_10_216 k_10_216(i_10_64, i_10_171, i_10_175, i_10_223, i_10_224, i_10_286, i_10_290, i_10_461, i_10_517, i_10_532, i_10_533, i_10_748, i_10_797, i_10_1026, i_10_1027, i_10_1029, i_10_1035, i_10_1236, i_10_1242, i_10_1243, i_10_1315, i_10_1547, i_10_1578, i_10_1579, i_10_1614, i_10_1687, i_10_1691, i_10_1822, i_10_1854, i_10_1915, i_10_1916, i_10_1954, i_10_1989, i_10_1991, i_10_1998, i_10_2151, i_10_2154, i_10_2179, i_10_2224, i_10_2304, i_10_2305, i_10_2307, i_10_2358, i_10_2361, i_10_2362, i_10_2364, i_10_2368, i_10_2448, i_10_2456, i_10_2457, i_10_2460, i_10_2461, i_10_2466, i_10_2467, i_10_2629, i_10_2631, i_10_2632, i_10_2677, i_10_2726, i_10_2730, i_10_2862, i_10_2983, i_10_3088, i_10_3196, i_10_3199, i_10_3231, i_10_3283, i_10_3303, i_10_3330, i_10_3333, i_10_3385, i_10_3442, i_10_3468, i_10_3520, i_10_3522, i_10_3609, i_10_3612, i_10_3613, i_10_3614, i_10_3681, i_10_3682, i_10_3684, i_10_3686, i_10_3840, i_10_3844, i_10_3856, i_10_3889, i_10_3930, i_10_3980, i_10_4024, i_10_4113, i_10_4124, i_10_4143, i_10_4212, i_10_4213, i_10_4216, i_10_4284, i_10_4350, i_10_4351, i_10_4590, o_10_216);
	kernel_10_217 k_10_217(i_10_172, i_10_177, i_10_223, i_10_283, i_10_316, i_10_318, i_10_330, i_10_409, i_10_410, i_10_411, i_10_412, i_10_413, i_10_512, i_10_993, i_10_1236, i_10_1238, i_10_1239, i_10_1240, i_10_1241, i_10_1243, i_10_1310, i_10_1365, i_10_1549, i_10_1552, i_10_1577, i_10_1581, i_10_1647, i_10_1683, i_10_1687, i_10_1820, i_10_1821, i_10_1945, i_10_2244, i_10_2339, i_10_2353, i_10_2381, i_10_2451, i_10_2453, i_10_2455, i_10_2466, i_10_2467, i_10_2468, i_10_2469, i_10_2473, i_10_2629, i_10_2630, i_10_2631, i_10_2632, i_10_2633, i_10_2635, i_10_2636, i_10_2659, i_10_2674, i_10_2703, i_10_2706, i_10_2728, i_10_2731, i_10_2732, i_10_2733, i_10_2781, i_10_2782, i_10_2785, i_10_2787, i_10_2788, i_10_2827, i_10_2834, i_10_2886, i_10_3042, i_10_3043, i_10_3044, i_10_3047, i_10_3151, i_10_3157, i_10_3158, i_10_3198, i_10_3237, i_10_3405, i_10_3408, i_10_3468, i_10_3472, i_10_3582, i_10_3585, i_10_3586, i_10_3588, i_10_3589, i_10_3617, i_10_3651, i_10_3652, i_10_3781, i_10_3785, i_10_3847, i_10_3853, i_10_3907, i_10_4054, i_10_4118, i_10_4119, i_10_4289, i_10_4292, i_10_4567, i_10_4584, o_10_217);
	kernel_10_218 k_10_218(i_10_42, i_10_89, i_10_180, i_10_181, i_10_183, i_10_184, i_10_250, i_10_280, i_10_287, i_10_292, i_10_293, i_10_408, i_10_409, i_10_412, i_10_426, i_10_436, i_10_444, i_10_795, i_10_796, i_10_798, i_10_957, i_10_958, i_10_997, i_10_1119, i_10_1167, i_10_1168, i_10_1237, i_10_1238, i_10_1239, i_10_1240, i_10_1247, i_10_1249, i_10_1250, i_10_1354, i_10_1363, i_10_1543, i_10_1758, i_10_1763, i_10_1824, i_10_1826, i_10_1909, i_10_1915, i_10_1995, i_10_1996, i_10_2005, i_10_2022, i_10_2023, i_10_2334, i_10_2353, i_10_2474, i_10_2608, i_10_2629, i_10_2633, i_10_2636, i_10_2677, i_10_2707, i_10_2719, i_10_2721, i_10_2722, i_10_2723, i_10_2729, i_10_2785, i_10_2788, i_10_2827, i_10_2829, i_10_2830, i_10_2923, i_10_2924, i_10_2983, i_10_3038, i_10_3048, i_10_3076, i_10_3270, i_10_3271, i_10_3283, i_10_3385, i_10_3387, i_10_3433, i_10_3612, i_10_3647, i_10_3649, i_10_3688, i_10_3689, i_10_3720, i_10_3835, i_10_3836, i_10_3841, i_10_3886, i_10_3982, i_10_3986, i_10_4027, i_10_4095, i_10_4120, i_10_4153, i_10_4180, i_10_4188, i_10_4189, i_10_4191, i_10_4272, i_10_4565, o_10_218);
	kernel_10_219 k_10_219(i_10_34, i_10_66, i_10_174, i_10_175, i_10_197, i_10_260, i_10_268, i_10_269, i_10_499, i_10_538, i_10_718, i_10_797, i_10_966, i_10_967, i_10_971, i_10_1030, i_10_1195, i_10_1196, i_10_1223, i_10_1241, i_10_1276, i_10_1277, i_10_1285, i_10_1302, i_10_1545, i_10_1556, i_10_1618, i_10_1641, i_10_1696, i_10_1697, i_10_1766, i_10_1767, i_10_1769, i_10_1822, i_10_1908, i_10_1943, i_10_1949, i_10_1957, i_10_2022, i_10_2023, i_10_2032, i_10_2033, i_10_2192, i_10_2203, i_10_2204, i_10_2348, i_10_2355, i_10_2356, i_10_2357, i_10_2456, i_10_2572, i_10_2580, i_10_2591, i_10_2599, i_10_2636, i_10_2705, i_10_2734, i_10_2761, i_10_2784, i_10_2785, i_10_2869, i_10_2883, i_10_2923, i_10_2959, i_10_2986, i_10_3026, i_10_3058, i_10_3059, i_10_3273, i_10_3281, i_10_3329, i_10_3473, i_10_3506, i_10_3571, i_10_3586, i_10_3605, i_10_3608, i_10_3616, i_10_3688, i_10_3839, i_10_3977, i_10_3984, i_10_3985, i_10_4013, i_10_4094, i_10_4126, i_10_4173, i_10_4183, i_10_4271, i_10_4272, i_10_4280, i_10_4281, i_10_4282, i_10_4283, i_10_4360, i_10_4379, i_10_4381, i_10_4461, i_10_4568, i_10_4569, o_10_219);
	kernel_10_220 k_10_220(i_10_51, i_10_88, i_10_150, i_10_186, i_10_187, i_10_258, i_10_269, i_10_372, i_10_408, i_10_464, i_10_565, i_10_642, i_10_762, i_10_793, i_10_794, i_10_826, i_10_853, i_10_854, i_10_898, i_10_996, i_10_1083, i_10_1086, i_10_1223, i_10_1305, i_10_1309, i_10_1396, i_10_1443, i_10_1551, i_10_1555, i_10_1556, i_10_1635, i_10_1636, i_10_1650, i_10_1651, i_10_1652, i_10_1653, i_10_1691, i_10_1713, i_10_1714, i_10_1732, i_10_1822, i_10_1883, i_10_1984, i_10_1986, i_10_2014, i_10_2026, i_10_2062, i_10_2157, i_10_2159, i_10_2227, i_10_2266, i_10_2290, i_10_2339, i_10_2365, i_10_2446, i_10_2451, i_10_2465, i_10_2568, i_10_2572, i_10_2634, i_10_2652, i_10_2661, i_10_2680, i_10_2711, i_10_2717, i_10_2730, i_10_2731, i_10_2734, i_10_2806, i_10_2850, i_10_3040, i_10_3091, i_10_3165, i_10_3166, i_10_3174, i_10_3273, i_10_3391, i_10_3408, i_10_3409, i_10_3410, i_10_3561, i_10_3611, i_10_3612, i_10_3613, i_10_3642, i_10_3803, i_10_3813, i_10_3854, i_10_3855, i_10_3856, i_10_3905, i_10_3923, i_10_4102, i_10_4120, i_10_4157, i_10_4174, i_10_4191, i_10_4269, i_10_4287, i_10_4552, o_10_220);
	kernel_10_221 k_10_221(i_10_34, i_10_172, i_10_224, i_10_247, i_10_259, i_10_280, i_10_283, i_10_319, i_10_409, i_10_410, i_10_447, i_10_448, i_10_466, i_10_749, i_10_752, i_10_792, i_10_795, i_10_799, i_10_955, i_10_956, i_10_1032, i_10_1033, i_10_1034, i_10_1234, i_10_1235, i_10_1240, i_10_1248, i_10_1305, i_10_1312, i_10_1432, i_10_1438, i_10_1442, i_10_1577, i_10_1579, i_10_1647, i_10_1648, i_10_1650, i_10_1651, i_10_1652, i_10_1687, i_10_1688, i_10_1689, i_10_1822, i_10_1996, i_10_2001, i_10_2022, i_10_2025, i_10_2230, i_10_2324, i_10_2358, i_10_2359, i_10_2361, i_10_2365, i_10_2455, i_10_2471, i_10_2473, i_10_2474, i_10_2631, i_10_2655, i_10_2657, i_10_2661, i_10_2701, i_10_2703, i_10_2713, i_10_2724, i_10_2923, i_10_3033, i_10_3070, i_10_3196, i_10_3202, i_10_3203, i_10_3277, i_10_3279, i_10_3384, i_10_3386, i_10_3391, i_10_3405, i_10_3406, i_10_3609, i_10_3616, i_10_3717, i_10_3780, i_10_3782, i_10_3783, i_10_3785, i_10_3786, i_10_3787, i_10_3808, i_10_3811, i_10_3839, i_10_3844, i_10_3845, i_10_3847, i_10_3860, i_10_4114, i_10_4273, i_10_4278, i_10_4285, i_10_4289, i_10_4291, o_10_221);
	kernel_10_222 k_10_222(i_10_218, i_10_219, i_10_220, i_10_221, i_10_279, i_10_280, i_10_391, i_10_424, i_10_425, i_10_431, i_10_460, i_10_461, i_10_462, i_10_463, i_10_464, i_10_712, i_10_713, i_10_794, i_10_899, i_10_990, i_10_999, i_10_1236, i_10_1237, i_10_1243, i_10_1244, i_10_1247, i_10_1250, i_10_1310, i_10_1365, i_10_1650, i_10_1652, i_10_1686, i_10_1688, i_10_1821, i_10_1824, i_10_1825, i_10_1915, i_10_2022, i_10_2180, i_10_2306, i_10_2350, i_10_2352, i_10_2353, i_10_2354, i_10_2359, i_10_2452, i_10_2454, i_10_2455, i_10_2464, i_10_2468, i_10_2471, i_10_2571, i_10_2628, i_10_2654, i_10_2660, i_10_2700, i_10_2701, i_10_2702, i_10_2723, i_10_2726, i_10_2734, i_10_2880, i_10_2887, i_10_2923, i_10_3037, i_10_3049, i_10_3050, i_10_3073, i_10_3165, i_10_3196, i_10_3200, i_10_3271, i_10_3387, i_10_3406, i_10_3408, i_10_3409, i_10_3613, i_10_3614, i_10_3645, i_10_3653, i_10_3732, i_10_3783, i_10_3784, i_10_3785, i_10_3837, i_10_3848, i_10_3854, i_10_3855, i_10_3856, i_10_3857, i_10_3991, i_10_4119, i_10_4120, i_10_4121, i_10_4270, i_10_4288, i_10_4289, i_10_4564, i_10_4565, i_10_4568, o_10_222);
	kernel_10_223 k_10_223(i_10_174, i_10_175, i_10_216, i_10_268, i_10_279, i_10_287, i_10_443, i_10_466, i_10_508, i_10_511, i_10_697, i_10_797, i_10_798, i_10_1005, i_10_1006, i_10_1234, i_10_1237, i_10_1240, i_10_1249, i_10_1310, i_10_1311, i_10_1647, i_10_1648, i_10_1650, i_10_1651, i_10_1652, i_10_1654, i_10_1684, i_10_1686, i_10_1820, i_10_1821, i_10_1823, i_10_1824, i_10_1825, i_10_1910, i_10_1913, i_10_1952, i_10_1994, i_10_1996, i_10_2179, i_10_2185, i_10_2203, i_10_2332, i_10_2337, i_10_2338, i_10_2339, i_10_2353, i_10_2366, i_10_2377, i_10_2380, i_10_2383, i_10_2384, i_10_2407, i_10_2408, i_10_2410, i_10_2451, i_10_2456, i_10_2569, i_10_2571, i_10_2572, i_10_2711, i_10_2730, i_10_2735, i_10_2883, i_10_3034, i_10_3037, i_10_3046, i_10_3047, i_10_3048, i_10_3049, i_10_3050, i_10_3069, i_10_3072, i_10_3074, i_10_3151, i_10_3153, i_10_3155, i_10_3158, i_10_3199, i_10_3267, i_10_3268, i_10_3271, i_10_3327, i_10_3405, i_10_3469, i_10_3497, i_10_3617, i_10_3650, i_10_3837, i_10_3838, i_10_3839, i_10_3846, i_10_3847, i_10_4056, i_10_4117, i_10_4118, i_10_4119, i_10_4120, i_10_4121, i_10_4285, o_10_223);
	kernel_10_224 k_10_224(i_10_29, i_10_216, i_10_283, i_10_284, i_10_308, i_10_374, i_10_433, i_10_444, i_10_505, i_10_558, i_10_623, i_10_794, i_10_821, i_10_847, i_10_893, i_10_895, i_10_901, i_10_1030, i_10_1031, i_10_1084, i_10_1085, i_10_1233, i_10_1235, i_10_1243, i_10_1548, i_10_1575, i_10_1606, i_10_1612, i_10_1616, i_10_1684, i_10_1825, i_10_1911, i_10_1956, i_10_1990, i_10_1991, i_10_2090, i_10_2225, i_10_2242, i_10_2304, i_10_2332, i_10_2335, i_10_2336, i_10_2361, i_10_2462, i_10_2556, i_10_2567, i_10_2632, i_10_2638, i_10_2639, i_10_2660, i_10_2675, i_10_2701, i_10_2702, i_10_2709, i_10_2728, i_10_2729, i_10_2783, i_10_2827, i_10_2829, i_10_2830, i_10_2867, i_10_2880, i_10_2917, i_10_2920, i_10_3160, i_10_3161, i_10_3315, i_10_3353, i_10_3385, i_10_3389, i_10_3440, i_10_3448, i_10_3457, i_10_3458, i_10_3551, i_10_3553, i_10_3557, i_10_3611, i_10_3614, i_10_3646, i_10_3784, i_10_3834, i_10_3837, i_10_3848, i_10_3856, i_10_3857, i_10_3880, i_10_3920, i_10_3978, i_10_4009, i_10_4010, i_10_4028, i_10_4051, i_10_4052, i_10_4213, i_10_4214, i_10_4291, i_10_4302, i_10_4564, i_10_4565, o_10_224);
	kernel_10_225 k_10_225(i_10_171, i_10_174, i_10_185, i_10_217, i_10_218, i_10_221, i_10_223, i_10_255, i_10_271, i_10_276, i_10_315, i_10_370, i_10_395, i_10_427, i_10_433, i_10_436, i_10_460, i_10_461, i_10_712, i_10_904, i_10_1027, i_10_1084, i_10_1120, i_10_1162, i_10_1237, i_10_1240, i_10_1242, i_10_1243, i_10_1246, i_10_1264, i_10_1308, i_10_1542, i_10_1544, i_10_1583, i_10_1650, i_10_1688, i_10_1908, i_10_1910, i_10_2304, i_10_2310, i_10_2312, i_10_2356, i_10_2359, i_10_2363, i_10_2367, i_10_2452, i_10_2458, i_10_2470, i_10_2471, i_10_2513, i_10_2713, i_10_2714, i_10_2721, i_10_2727, i_10_2730, i_10_2831, i_10_2884, i_10_2923, i_10_2982, i_10_3034, i_10_3036, i_10_3198, i_10_3199, i_10_3280, i_10_3297, i_10_3335, i_10_3390, i_10_3402, i_10_3405, i_10_3406, i_10_3410, i_10_3430, i_10_3586, i_10_3609, i_10_3612, i_10_3616, i_10_3652, i_10_3689, i_10_3730, i_10_3731, i_10_3780, i_10_3783, i_10_3784, i_10_3821, i_10_3840, i_10_3855, i_10_3858, i_10_3892, i_10_3943, i_10_3991, i_10_3992, i_10_3998, i_10_4173, i_10_4174, i_10_4213, i_10_4214, i_10_4274, i_10_4288, i_10_4289, i_10_4567, o_10_225);
	kernel_10_226 k_10_226(i_10_223, i_10_269, i_10_292, i_10_320, i_10_323, i_10_432, i_10_437, i_10_446, i_10_448, i_10_462, i_10_466, i_10_503, i_10_509, i_10_628, i_10_629, i_10_711, i_10_716, i_10_799, i_10_896, i_10_968, i_10_1011, i_10_1034, i_10_1106, i_10_1124, i_10_1156, i_10_1223, i_10_1270, i_10_1354, i_10_1439, i_10_1441, i_10_1442, i_10_1448, i_10_1492, i_10_1545, i_10_1581, i_10_1582, i_10_1637, i_10_1689, i_10_1690, i_10_1691, i_10_1736, i_10_1808, i_10_1822, i_10_1984, i_10_1994, i_10_2005, i_10_2006, i_10_2033, i_10_2202, i_10_2223, i_10_2347, i_10_2352, i_10_2365, i_10_2366, i_10_2451, i_10_2474, i_10_2635, i_10_2659, i_10_2679, i_10_2680, i_10_2704, i_10_2715, i_10_2722, i_10_2732, i_10_2762, i_10_2782, i_10_2833, i_10_2919, i_10_2924, i_10_2969, i_10_2978, i_10_3077, i_10_3199, i_10_3281, i_10_3389, i_10_3409, i_10_3465, i_10_3467, i_10_3473, i_10_3494, i_10_3497, i_10_3538, i_10_3545, i_10_3587, i_10_3590, i_10_3649, i_10_3853, i_10_3914, i_10_3923, i_10_4122, i_10_4210, i_10_4211, i_10_4269, i_10_4271, i_10_4273, i_10_4281, i_10_4291, i_10_4395, i_10_4584, i_10_4589, o_10_226);
	kernel_10_227 k_10_227(i_10_122, i_10_171, i_10_174, i_10_175, i_10_176, i_10_282, i_10_283, i_10_319, i_10_387, i_10_409, i_10_434, i_10_445, i_10_460, i_10_461, i_10_462, i_10_464, i_10_497, i_10_713, i_10_752, i_10_900, i_10_1048, i_10_1084, i_10_1237, i_10_1238, i_10_1279, i_10_1310, i_10_1342, i_10_1354, i_10_1435, i_10_1539, i_10_1540, i_10_1580, i_10_1651, i_10_1687, i_10_1688, i_10_1690, i_10_1691, i_10_1909, i_10_2033, i_10_2201, i_10_2359, i_10_2379, i_10_2452, i_10_2455, i_10_2468, i_10_2629, i_10_2630, i_10_2644, i_10_2656, i_10_2657, i_10_2658, i_10_2659, i_10_2679, i_10_2711, i_10_2720, i_10_2722, i_10_2789, i_10_2817, i_10_3070, i_10_3071, i_10_3200, i_10_3276, i_10_3277, i_10_3278, i_10_3279, i_10_3280, i_10_3281, i_10_3283, i_10_3316, i_10_3385, i_10_3387, i_10_3392, i_10_3496, i_10_3538, i_10_3541, i_10_3587, i_10_3686, i_10_3837, i_10_3838, i_10_3839, i_10_3849, i_10_3856, i_10_3857, i_10_3859, i_10_3860, i_10_3888, i_10_3889, i_10_3981, i_10_3982, i_10_4114, i_10_4118, i_10_4167, i_10_4170, i_10_4171, i_10_4269, i_10_4270, i_10_4287, i_10_4288, i_10_4289, i_10_4290, o_10_227);
	kernel_10_228 k_10_228(i_10_38, i_10_148, i_10_286, i_10_287, i_10_356, i_10_358, i_10_359, i_10_365, i_10_374, i_10_410, i_10_428, i_10_446, i_10_464, i_10_635, i_10_719, i_10_734, i_10_736, i_10_737, i_10_755, i_10_793, i_10_800, i_10_832, i_10_905, i_10_955, i_10_959, i_10_994, i_10_1054, i_10_1088, i_10_1136, i_10_1162, i_10_1163, i_10_1166, i_10_1219, i_10_1235, i_10_1238, i_10_1262, i_10_1289, i_10_1292, i_10_1349, i_10_1355, i_10_1493, i_10_1535, i_10_1651, i_10_1652, i_10_1694, i_10_1823, i_10_1847, i_10_1850, i_10_1913, i_10_1958, i_10_2003, i_10_2207, i_10_2213, i_10_2249, i_10_2386, i_10_2387, i_10_2390, i_10_2408, i_10_2452, i_10_2454, i_10_2455, i_10_2495, i_10_2519, i_10_2543, i_10_2609, i_10_2611, i_10_2632, i_10_2633, i_10_2659, i_10_2678, i_10_2833, i_10_2980, i_10_2984, i_10_3119, i_10_3278, i_10_3283, i_10_3292, i_10_3293, i_10_3317, i_10_3326, i_10_3362, i_10_3385, i_10_3386, i_10_3388, i_10_3526, i_10_3539, i_10_3581, i_10_3584, i_10_3616, i_10_3638, i_10_3777, i_10_3824, i_10_4001, i_10_4061, i_10_4064, i_10_4115, i_10_4306, i_10_4382, i_10_4484, i_10_4571, o_10_228);
	kernel_10_229 k_10_229(i_10_174, i_10_175, i_10_176, i_10_184, i_10_270, i_10_286, i_10_287, i_10_319, i_10_409, i_10_410, i_10_436, i_10_438, i_10_440, i_10_446, i_10_447, i_10_448, i_10_449, i_10_466, i_10_467, i_10_518, i_10_717, i_10_718, i_10_719, i_10_755, i_10_793, i_10_797, i_10_798, i_10_799, i_10_958, i_10_968, i_10_971, i_10_1003, i_10_1006, i_10_1164, i_10_1165, i_10_1166, i_10_1169, i_10_1237, i_10_1245, i_10_1247, i_10_1249, i_10_1250, i_10_1309, i_10_1311, i_10_1435, i_10_1624, i_10_1654, i_10_1655, i_10_1765, i_10_1822, i_10_1823, i_10_1909, i_10_2095, i_10_2179, i_10_2308, i_10_2350, i_10_2351, i_10_2407, i_10_2634, i_10_2635, i_10_2636, i_10_2724, i_10_2727, i_10_2728, i_10_2734, i_10_2783, i_10_2784, i_10_2830, i_10_2834, i_10_2883, i_10_2920, i_10_2986, i_10_3038, i_10_3039, i_10_3041, i_10_3048, i_10_3271, i_10_3273, i_10_3617, i_10_3652, i_10_3653, i_10_3783, i_10_3839, i_10_3840, i_10_3846, i_10_3851, i_10_3895, i_10_3982, i_10_3983, i_10_3985, i_10_4116, i_10_4120, i_10_4121, i_10_4125, i_10_4188, i_10_4192, i_10_4270, i_10_4272, i_10_4290, i_10_4291, o_10_229);
	kernel_10_230 k_10_230(i_10_268, i_10_269, i_10_282, i_10_283, i_10_315, i_10_316, i_10_321, i_10_327, i_10_390, i_10_408, i_10_412, i_10_439, i_10_440, i_10_501, i_10_516, i_10_664, i_10_685, i_10_826, i_10_960, i_10_969, i_10_1030, i_10_1105, i_10_1113, i_10_1242, i_10_1248, i_10_1264, i_10_1302, i_10_1303, i_10_1357, i_10_1447, i_10_1547, i_10_1556, i_10_1578, i_10_1579, i_10_1580, i_10_1618, i_10_1627, i_10_1683, i_10_1689, i_10_1734, i_10_1735, i_10_1806, i_10_1819, i_10_1821, i_10_1945, i_10_1984, i_10_1986, i_10_2005, i_10_2035, i_10_2243, i_10_2353, i_10_2355, i_10_2356, i_10_2383, i_10_2384, i_10_2449, i_10_2451, i_10_2452, i_10_2472, i_10_2569, i_10_2572, i_10_2631, i_10_2635, i_10_2662, i_10_2733, i_10_2734, i_10_2832, i_10_2919, i_10_2920, i_10_3037, i_10_3069, i_10_3280, i_10_3281, i_10_3283, i_10_3329, i_10_3390, i_10_3391, i_10_3472, i_10_3501, i_10_3504, i_10_3508, i_10_3540, i_10_3541, i_10_3612, i_10_3613, i_10_3785, i_10_3837, i_10_3839, i_10_3841, i_10_3850, i_10_3852, i_10_3859, i_10_3860, i_10_3871, i_10_4030, i_10_4116, i_10_4117, i_10_4120, i_10_4171, i_10_4173, o_10_230);
	kernel_10_231 k_10_231(i_10_28, i_10_29, i_10_146, i_10_172, i_10_220, i_10_243, i_10_252, i_10_387, i_10_433, i_10_519, i_10_570, i_10_687, i_10_711, i_10_712, i_10_747, i_10_748, i_10_752, i_10_846, i_10_954, i_10_1029, i_10_1237, i_10_1305, i_10_1309, i_10_1313, i_10_1377, i_10_1539, i_10_1575, i_10_1614, i_10_1617, i_10_1683, i_10_1686, i_10_1688, i_10_1823, i_10_1826, i_10_2178, i_10_2179, i_10_2308, i_10_2451, i_10_2462, i_10_2463, i_10_2470, i_10_2471, i_10_2529, i_10_2530, i_10_2535, i_10_2601, i_10_2602, i_10_2604, i_10_2628, i_10_2640, i_10_2662, i_10_2728, i_10_2830, i_10_2831, i_10_2924, i_10_2995, i_10_3070, i_10_3072, i_10_3156, i_10_3195, i_10_3196, i_10_3234, i_10_3278, i_10_3385, i_10_3386, i_10_3389, i_10_3405, i_10_3406, i_10_3408, i_10_3441, i_10_3444, i_10_3523, i_10_3525, i_10_3552, i_10_3586, i_10_3609, i_10_3612, i_10_3616, i_10_3646, i_10_3649, i_10_3726, i_10_3780, i_10_3781, i_10_3807, i_10_3808, i_10_3839, i_10_3845, i_10_3849, i_10_3879, i_10_3880, i_10_4113, i_10_4114, i_10_4116, i_10_4117, i_10_4118, i_10_4212, i_10_4216, i_10_4284, i_10_4456, i_10_4582, o_10_231);
	kernel_10_232 k_10_232(i_10_177, i_10_183, i_10_184, i_10_186, i_10_187, i_10_188, i_10_220, i_10_244, i_10_282, i_10_283, i_10_284, i_10_316, i_10_406, i_10_410, i_10_429, i_10_436, i_10_437, i_10_438, i_10_439, i_10_442, i_10_459, i_10_794, i_10_996, i_10_1026, i_10_1027, i_10_1033, i_10_1042, i_10_1043, i_10_1236, i_10_1247, i_10_1250, i_10_1435, i_10_1444, i_10_1445, i_10_1447, i_10_1540, i_10_1543, i_10_1544, i_10_1547, i_10_1575, i_10_1576, i_10_1579, i_10_1582, i_10_1583, i_10_1650, i_10_1652, i_10_1653, i_10_1683, i_10_1684, i_10_1686, i_10_1820, i_10_1821, i_10_1915, i_10_2183, i_10_2407, i_10_2473, i_10_2478, i_10_2566, i_10_2628, i_10_2630, i_10_2633, i_10_2657, i_10_2658, i_10_2659, i_10_2660, i_10_2662, i_10_2663, i_10_2680, i_10_2708, i_10_2716, i_10_2728, i_10_2732, i_10_2883, i_10_2922, i_10_3040, i_10_3069, i_10_3070, i_10_3152, i_10_3278, i_10_3329, i_10_3386, i_10_3408, i_10_3465, i_10_3544, i_10_3783, i_10_3837, i_10_3838, i_10_3839, i_10_3842, i_10_3846, i_10_3847, i_10_3895, i_10_4114, i_10_4273, i_10_4278, i_10_4282, i_10_4286, i_10_4291, i_10_4292, i_10_4563, o_10_232);
	kernel_10_233 k_10_233(i_10_153, i_10_243, i_10_318, i_10_442, i_10_460, i_10_463, i_10_498, i_10_513, i_10_516, i_10_565, i_10_622, i_10_864, i_10_865, i_10_903, i_10_993, i_10_1026, i_10_1045, i_10_1080, i_10_1235, i_10_1263, i_10_1264, i_10_1449, i_10_1450, i_10_1551, i_10_1623, i_10_1683, i_10_1690, i_10_1809, i_10_1812, i_10_1819, i_10_1825, i_10_1826, i_10_1878, i_10_1909, i_10_1910, i_10_1913, i_10_1989, i_10_2002, i_10_2199, i_10_2200, i_10_2308, i_10_2349, i_10_2353, i_10_2357, i_10_2376, i_10_2377, i_10_2450, i_10_2451, i_10_2452, i_10_2453, i_10_2469, i_10_2505, i_10_2565, i_10_2574, i_10_2657, i_10_2673, i_10_2700, i_10_2701, i_10_2703, i_10_2723, i_10_2732, i_10_2735, i_10_2827, i_10_2880, i_10_2952, i_10_2961, i_10_2983, i_10_3042, i_10_3159, i_10_3196, i_10_3283, i_10_3284, i_10_3315, i_10_3388, i_10_3389, i_10_3555, i_10_3613, i_10_3614, i_10_3649, i_10_3685, i_10_3780, i_10_3784, i_10_3810, i_10_3839, i_10_3843, i_10_3858, i_10_3876, i_10_3979, i_10_4118, i_10_4121, i_10_4122, i_10_4123, i_10_4126, i_10_4128, i_10_4186, i_10_4266, i_10_4286, i_10_4289, i_10_4564, i_10_4566, o_10_233);
	kernel_10_234 k_10_234(i_10_31, i_10_318, i_10_393, i_10_444, i_10_447, i_10_459, i_10_460, i_10_463, i_10_467, i_10_792, i_10_849, i_10_970, i_10_1036, i_10_1039, i_10_1040, i_10_1242, i_10_1308, i_10_1360, i_10_1382, i_10_1409, i_10_1444, i_10_1447, i_10_1465, i_10_1552, i_10_1650, i_10_1757, i_10_1912, i_10_1918, i_10_2012, i_10_2029, i_10_2096, i_10_2157, i_10_2332, i_10_2338, i_10_2339, i_10_2434, i_10_2445, i_10_2461, i_10_2470, i_10_2526, i_10_2579, i_10_2632, i_10_2659, i_10_2702, i_10_2705, i_10_2709, i_10_2710, i_10_2711, i_10_2714, i_10_2887, i_10_2916, i_10_2917, i_10_2919, i_10_2924, i_10_2954, i_10_3033, i_10_3057, i_10_3208, i_10_3277, i_10_3279, i_10_3284, i_10_3297, i_10_3386, i_10_3387, i_10_3388, i_10_3391, i_10_3403, i_10_3408, i_10_3409, i_10_3451, i_10_3496, i_10_3497, i_10_3500, i_10_3550, i_10_3577, i_10_3611, i_10_3615, i_10_3684, i_10_3717, i_10_3719, i_10_3720, i_10_3722, i_10_3854, i_10_3860, i_10_3889, i_10_3965, i_10_4030, i_10_4119, i_10_4186, i_10_4188, i_10_4189, i_10_4204, i_10_4270, i_10_4271, i_10_4272, i_10_4273, i_10_4274, i_10_4290, i_10_4291, i_10_4531, o_10_234);
	kernel_10_235 k_10_235(i_10_49, i_10_173, i_10_174, i_10_175, i_10_176, i_10_244, i_10_257, i_10_315, i_10_371, i_10_389, i_10_394, i_10_395, i_10_407, i_10_411, i_10_412, i_10_427, i_10_435, i_10_439, i_10_500, i_10_503, i_10_520, i_10_521, i_10_590, i_10_716, i_10_792, i_10_989, i_10_1031, i_10_1235, i_10_1244, i_10_1306, i_10_1313, i_10_1362, i_10_1436, i_10_1583, i_10_1634, i_10_1654, i_10_1655, i_10_1685, i_10_1686, i_10_1687, i_10_1688, i_10_1719, i_10_1720, i_10_1824, i_10_1826, i_10_1909, i_10_2003, i_10_2198, i_10_2351, i_10_2352, i_10_2380, i_10_2456, i_10_2468, i_10_2471, i_10_2531, i_10_2634, i_10_2690, i_10_2719, i_10_2722, i_10_2732, i_10_2833, i_10_2834, i_10_2923, i_10_3074, i_10_3200, i_10_3271, i_10_3278, i_10_3332, i_10_3466, i_10_3506, i_10_3509, i_10_3610, i_10_3613, i_10_3616, i_10_3646, i_10_3648, i_10_3649, i_10_3651, i_10_3652, i_10_3653, i_10_3721, i_10_3780, i_10_3781, i_10_3782, i_10_3840, i_10_3841, i_10_3842, i_10_3855, i_10_3856, i_10_3910, i_10_3911, i_10_4029, i_10_4126, i_10_4171, i_10_4189, i_10_4268, i_10_4270, i_10_4271, i_10_4288, i_10_4289, o_10_235);
	kernel_10_236 k_10_236(i_10_71, i_10_89, i_10_145, i_10_146, i_10_172, i_10_174, i_10_175, i_10_224, i_10_248, i_10_286, i_10_287, i_10_393, i_10_408, i_10_439, i_10_446, i_10_462, i_10_464, i_10_466, i_10_691, i_10_794, i_10_796, i_10_800, i_10_1042, i_10_1043, i_10_1165, i_10_1168, i_10_1237, i_10_1240, i_10_1241, i_10_1306, i_10_1308, i_10_1364, i_10_1450, i_10_1540, i_10_1555, i_10_1613, i_10_1653, i_10_1654, i_10_1735, i_10_1760, i_10_1821, i_10_1823, i_10_1824, i_10_1915, i_10_2159, i_10_2246, i_10_2248, i_10_2249, i_10_2309, i_10_2329, i_10_2350, i_10_2352, i_10_2361, i_10_2380, i_10_2451, i_10_2456, i_10_2473, i_10_2581, i_10_2658, i_10_2730, i_10_2734, i_10_2841, i_10_2881, i_10_2922, i_10_2923, i_10_2941, i_10_2942, i_10_3036, i_10_3037, i_10_3073, i_10_3198, i_10_3202, i_10_3388, i_10_3405, i_10_3470, i_10_3610, i_10_3613, i_10_3614, i_10_3615, i_10_3649, i_10_3674, i_10_3686, i_10_3703, i_10_3788, i_10_3810, i_10_3838, i_10_3853, i_10_3855, i_10_3856, i_10_3858, i_10_3859, i_10_3860, i_10_3883, i_10_3967, i_10_4267, i_10_4270, i_10_4271, i_10_4292, i_10_4463, i_10_4606, o_10_236);
	kernel_10_237 k_10_237(i_10_66, i_10_121, i_10_177, i_10_193, i_10_252, i_10_253, i_10_256, i_10_262, i_10_393, i_10_499, i_10_558, i_10_561, i_10_562, i_10_606, i_10_693, i_10_694, i_10_696, i_10_759, i_10_946, i_10_1002, i_10_1107, i_10_1110, i_10_1129, i_10_1233, i_10_1236, i_10_1281, i_10_1282, i_10_1296, i_10_1299, i_10_1432, i_10_1434, i_10_1435, i_10_1438, i_10_1539, i_10_1540, i_10_1542, i_10_1549, i_10_1550, i_10_1552, i_10_1553, i_10_1624, i_10_1625, i_10_1651, i_10_1654, i_10_1820, i_10_2092, i_10_2155, i_10_2156, i_10_2235, i_10_2238, i_10_2244, i_10_2289, i_10_2290, i_10_2350, i_10_2352, i_10_2353, i_10_2529, i_10_2531, i_10_2556, i_10_2565, i_10_2566, i_10_2570, i_10_2584, i_10_2587, i_10_2595, i_10_2694, i_10_2757, i_10_2782, i_10_2881, i_10_2944, i_10_2957, i_10_2989, i_10_3055, i_10_3070, i_10_3171, i_10_3198, i_10_3277, i_10_3279, i_10_3462, i_10_3567, i_10_3793, i_10_3858, i_10_3979, i_10_4027, i_10_4053, i_10_4153, i_10_4156, i_10_4167, i_10_4170, i_10_4171, i_10_4180, i_10_4189, i_10_4266, i_10_4275, i_10_4279, i_10_4378, i_10_4545, i_10_4549, i_10_4563, i_10_4564, o_10_237);
	kernel_10_238 k_10_238(i_10_171, i_10_247, i_10_282, i_10_286, i_10_287, i_10_390, i_10_406, i_10_408, i_10_429, i_10_435, i_10_444, i_10_445, i_10_448, i_10_449, i_10_521, i_10_793, i_10_966, i_10_967, i_10_992, i_10_1001, i_10_1007, i_10_1233, i_10_1238, i_10_1241, i_10_1246, i_10_1311, i_10_1360, i_10_1541, i_10_1552, i_10_1553, i_10_1555, i_10_1622, i_10_1655, i_10_1721, i_10_1730, i_10_1820, i_10_1824, i_10_1825, i_10_1826, i_10_1913, i_10_2030, i_10_2332, i_10_2333, i_10_2337, i_10_2338, i_10_2351, i_10_2352, i_10_2353, i_10_2377, i_10_2379, i_10_2380, i_10_2381, i_10_2383, i_10_2384, i_10_2405, i_10_2410, i_10_2570, i_10_2638, i_10_2656, i_10_2658, i_10_2659, i_10_2660, i_10_2701, i_10_2716, i_10_2721, i_10_2734, i_10_2917, i_10_2953, i_10_2963, i_10_2979, i_10_2980, i_10_2985, i_10_3038, i_10_3045, i_10_3151, i_10_3152, i_10_3153, i_10_3154, i_10_3155, i_10_3199, i_10_3268, i_10_3317, i_10_3388, i_10_3389, i_10_3437, i_10_3495, i_10_3497, i_10_3582, i_10_3650, i_10_3837, i_10_3842, i_10_3856, i_10_3857, i_10_3982, i_10_4114, i_10_4267, i_10_4270, i_10_4271, i_10_4274, i_10_4565, o_10_238);
	kernel_10_239 k_10_239(i_10_30, i_10_61, i_10_64, i_10_249, i_10_250, i_10_258, i_10_282, i_10_292, i_10_318, i_10_319, i_10_324, i_10_327, i_10_361, i_10_405, i_10_436, i_10_438, i_10_444, i_10_445, i_10_448, i_10_627, i_10_663, i_10_870, i_10_877, i_10_954, i_10_959, i_10_1156, i_10_1159, i_10_1234, i_10_1260, i_10_1308, i_10_1309, i_10_1347, i_10_1437, i_10_1441, i_10_1542, i_10_1545, i_10_1546, i_10_1581, i_10_1626, i_10_1641, i_10_1689, i_10_1690, i_10_1765, i_10_1766, i_10_1992, i_10_2022, i_10_2031, i_10_2094, i_10_2199, i_10_2292, i_10_2323, i_10_2346, i_10_2352, i_10_2355, i_10_2452, i_10_2470, i_10_2506, i_10_2535, i_10_2634, i_10_2635, i_10_2712, i_10_2731, i_10_2742, i_10_2850, i_10_2868, i_10_2888, i_10_2919, i_10_2967, i_10_2989, i_10_3075, i_10_3076, i_10_3166, i_10_3279, i_10_3281, i_10_3328, i_10_3336, i_10_3391, i_10_3431, i_10_3468, i_10_3469, i_10_3498, i_10_3586, i_10_3588, i_10_3609, i_10_3616, i_10_3846, i_10_3913, i_10_3984, i_10_4011, i_10_4113, i_10_4114, i_10_4116, i_10_4119, i_10_4209, i_10_4216, i_10_4231, i_10_4272, i_10_4502, i_10_4505, i_10_4568, o_10_239);
	kernel_10_240 k_10_240(i_10_159, i_10_264, i_10_265, i_10_273, i_10_274, i_10_284, i_10_286, i_10_439, i_10_444, i_10_446, i_10_447, i_10_465, i_10_467, i_10_754, i_10_755, i_10_797, i_10_799, i_10_800, i_10_898, i_10_899, i_10_964, i_10_996, i_10_1002, i_10_1027, i_10_1031, i_10_1032, i_10_1033, i_10_1034, i_10_1236, i_10_1241, i_10_1245, i_10_1246, i_10_1306, i_10_1308, i_10_1309, i_10_1312, i_10_1431, i_10_1576, i_10_1579, i_10_1597, i_10_1650, i_10_1651, i_10_1652, i_10_1689, i_10_1813, i_10_1913, i_10_1920, i_10_2202, i_10_2363, i_10_2383, i_10_2469, i_10_2473, i_10_2571, i_10_2609, i_10_2635, i_10_2702, i_10_2717, i_10_2719, i_10_2734, i_10_2829, i_10_2833, i_10_2880, i_10_2883, i_10_2918, i_10_2919, i_10_2921, i_10_3074, i_10_3151, i_10_3163, i_10_3165, i_10_3166, i_10_3196, i_10_3200, i_10_3274, i_10_3403, i_10_3409, i_10_3410, i_10_3589, i_10_3610, i_10_3612, i_10_3616, i_10_3649, i_10_3653, i_10_3781, i_10_3782, i_10_3855, i_10_3856, i_10_3880, i_10_3913, i_10_4116, i_10_4117, i_10_4120, i_10_4126, i_10_4128, i_10_4129, i_10_4130, i_10_4219, i_10_4273, i_10_4287, i_10_4288, o_10_240);
	kernel_10_241 k_10_241(i_10_171, i_10_172, i_10_175, i_10_176, i_10_220, i_10_221, i_10_223, i_10_250, i_10_282, i_10_283, i_10_284, i_10_432, i_10_433, i_10_434, i_10_441, i_10_463, i_10_794, i_10_797, i_10_892, i_10_968, i_10_1082, i_10_1236, i_10_1243, i_10_1244, i_10_1248, i_10_1347, i_10_1348, i_10_1360, i_10_1365, i_10_1441, i_10_1575, i_10_1652, i_10_1683, i_10_1687, i_10_1688, i_10_1768, i_10_1818, i_10_1819, i_10_1824, i_10_1825, i_10_2186, i_10_2354, i_10_2361, i_10_2382, i_10_2384, i_10_2448, i_10_2449, i_10_2450, i_10_2461, i_10_2469, i_10_2629, i_10_2632, i_10_2633, i_10_2656, i_10_2657, i_10_2658, i_10_2659, i_10_2721, i_10_2725, i_10_2727, i_10_2728, i_10_2729, i_10_2787, i_10_2827, i_10_2829, i_10_2830, i_10_2831, i_10_2883, i_10_2916, i_10_2983, i_10_3037, i_10_3039, i_10_3040, i_10_3075, i_10_3151, i_10_3153, i_10_3156, i_10_3195, i_10_3198, i_10_3238, i_10_3384, i_10_3387, i_10_3434, i_10_3610, i_10_3647, i_10_3648, i_10_3649, i_10_3652, i_10_3653, i_10_3784, i_10_3786, i_10_3835, i_10_3840, i_10_3855, i_10_3856, i_10_3857, i_10_3988, i_10_4056, i_10_4266, i_10_4269, o_10_241);
	kernel_10_242 k_10_242(i_10_22, i_10_172, i_10_217, i_10_273, i_10_274, i_10_282, i_10_508, i_10_531, i_10_586, i_10_729, i_10_730, i_10_733, i_10_792, i_10_828, i_10_1120, i_10_1243, i_10_1245, i_10_1377, i_10_1378, i_10_1386, i_10_1440, i_10_1521, i_10_1522, i_10_1559, i_10_1602, i_10_1649, i_10_1651, i_10_1652, i_10_1684, i_10_1685, i_10_1693, i_10_1767, i_10_1768, i_10_1824, i_10_1882, i_10_1913, i_10_1926, i_10_1929, i_10_1944, i_10_1945, i_10_1947, i_10_1981, i_10_2181, i_10_2331, i_10_2334, i_10_2376, i_10_2377, i_10_2380, i_10_2443, i_10_2475, i_10_2542, i_10_2630, i_10_2640, i_10_2673, i_10_2674, i_10_2689, i_10_2728, i_10_2729, i_10_2865, i_10_2872, i_10_2935, i_10_2965, i_10_2990, i_10_3096, i_10_3224, i_10_3231, i_10_3404, i_10_3519, i_10_3520, i_10_3521, i_10_3592, i_10_3614, i_10_3646, i_10_3726, i_10_3846, i_10_3847, i_10_3849, i_10_3850, i_10_3861, i_10_3889, i_10_3906, i_10_3961, i_10_4120, i_10_4176, i_10_4177, i_10_4266, i_10_4267, i_10_4269, i_10_4275, i_10_4302, i_10_4305, i_10_4306, i_10_4432, i_10_4437, i_10_4458, i_10_4459, i_10_4509, i_10_4510, i_10_4519, i_10_4567, o_10_242);
	kernel_10_243 k_10_243(i_10_48, i_10_49, i_10_50, i_10_145, i_10_244, i_10_253, i_10_274, i_10_281, i_10_283, i_10_284, i_10_320, i_10_425, i_10_433, i_10_450, i_10_515, i_10_711, i_10_712, i_10_796, i_10_800, i_10_956, i_10_963, i_10_1000, i_10_1237, i_10_1239, i_10_1241, i_10_1311, i_10_1360, i_10_1433, i_10_1532, i_10_1539, i_10_1577, i_10_1653, i_10_1718, i_10_1768, i_10_1769, i_10_1818, i_10_1819, i_10_1821, i_10_1911, i_10_1912, i_10_1913, i_10_1916, i_10_1917, i_10_2366, i_10_2383, i_10_2450, i_10_2452, i_10_2453, i_10_2459, i_10_2468, i_10_2470, i_10_2543, i_10_2629, i_10_2630, i_10_2659, i_10_2710, i_10_2711, i_10_2715, i_10_2717, i_10_2719, i_10_2721, i_10_2722, i_10_2723, i_10_2728, i_10_2729, i_10_2781, i_10_2782, i_10_2783, i_10_2827, i_10_2829, i_10_2830, i_10_2833, i_10_2916, i_10_2953, i_10_3069, i_10_3155, i_10_3196, i_10_3278, i_10_3281, i_10_3384, i_10_3385, i_10_3386, i_10_3405, i_10_3406, i_10_3466, i_10_3467, i_10_3522, i_10_3523, i_10_3615, i_10_3616, i_10_3647, i_10_3648, i_10_3685, i_10_3834, i_10_3848, i_10_3856, i_10_3857, i_10_4171, i_10_4231, i_10_4279, o_10_243);
	kernel_10_244 k_10_244(i_10_277, i_10_279, i_10_282, i_10_286, i_10_287, i_10_328, i_10_329, i_10_405, i_10_408, i_10_410, i_10_413, i_10_424, i_10_425, i_10_430, i_10_436, i_10_439, i_10_440, i_10_464, i_10_518, i_10_713, i_10_796, i_10_958, i_10_959, i_10_996, i_10_997, i_10_1138, i_10_1234, i_10_1238, i_10_1265, i_10_1346, i_10_1546, i_10_1552, i_10_1555, i_10_1556, i_10_1768, i_10_1818, i_10_1819, i_10_1823, i_10_1825, i_10_1826, i_10_1912, i_10_1915, i_10_2021, i_10_2407, i_10_2408, i_10_2471, i_10_2474, i_10_2508, i_10_2515, i_10_2542, i_10_2633, i_10_2656, i_10_2658, i_10_2679, i_10_2680, i_10_2681, i_10_2705, i_10_2707, i_10_2723, i_10_2726, i_10_2730, i_10_2732, i_10_2785, i_10_2823, i_10_2829, i_10_2830, i_10_2831, i_10_2959, i_10_2979, i_10_2983, i_10_2984, i_10_2986, i_10_3034, i_10_3039, i_10_3070, i_10_3072, i_10_3157, i_10_3158, i_10_3387, i_10_3391, i_10_3496, i_10_3497, i_10_3499, i_10_3519, i_10_3522, i_10_3523, i_10_3525, i_10_3586, i_10_3612, i_10_3613, i_10_3614, i_10_3648, i_10_3784, i_10_3786, i_10_3839, i_10_3847, i_10_3849, i_10_3855, i_10_3985, i_10_3986, o_10_244);
	kernel_10_245 k_10_245(i_10_17, i_10_149, i_10_187, i_10_242, i_10_263, i_10_431, i_10_448, i_10_463, i_10_563, i_10_586, i_10_587, i_10_659, i_10_694, i_10_712, i_10_824, i_10_892, i_10_893, i_10_896, i_10_899, i_10_950, i_10_997, i_10_1000, i_10_1109, i_10_1111, i_10_1112, i_10_1237, i_10_1270, i_10_1283, i_10_1300, i_10_1301, i_10_1304, i_10_1345, i_10_1346, i_10_1388, i_10_1439, i_10_1577, i_10_1579, i_10_1606, i_10_1732, i_10_1765, i_10_1799, i_10_1807, i_10_1883, i_10_1913, i_10_1940, i_10_1985, i_10_2011, i_10_2030, i_10_2152, i_10_2200, i_10_2210, i_10_2291, i_10_2350, i_10_2351, i_10_2450, i_10_2453, i_10_2515, i_10_2533, i_10_2556, i_10_2558, i_10_2560, i_10_2567, i_10_2570, i_10_2573, i_10_2660, i_10_2711, i_10_2713, i_10_2833, i_10_2846, i_10_2876, i_10_2885, i_10_2888, i_10_2957, i_10_3173, i_10_3277, i_10_3359, i_10_3395, i_10_3406, i_10_3464, i_10_3470, i_10_3520, i_10_3521, i_10_3560, i_10_3614, i_10_3649, i_10_3652, i_10_3841, i_10_3842, i_10_3920, i_10_3974, i_10_3983, i_10_4031, i_10_4117, i_10_4145, i_10_4151, i_10_4169, i_10_4172, i_10_4181, i_10_4268, i_10_4286, o_10_245);
	kernel_10_246 k_10_246(i_10_35, i_10_122, i_10_161, i_10_251, i_10_323, i_10_349, i_10_390, i_10_391, i_10_436, i_10_446, i_10_448, i_10_449, i_10_462, i_10_465, i_10_601, i_10_754, i_10_957, i_10_998, i_10_1004, i_10_1033, i_10_1034, i_10_1052, i_10_1058, i_10_1083, i_10_1084, i_10_1223, i_10_1291, i_10_1308, i_10_1382, i_10_1385, i_10_1579, i_10_1580, i_10_1651, i_10_1655, i_10_1736, i_10_1816, i_10_1818, i_10_1822, i_10_1823, i_10_1913, i_10_1961, i_10_2024, i_10_2086, i_10_2264, i_10_2384, i_10_2452, i_10_2453, i_10_2474, i_10_2609, i_10_2617, i_10_2657, i_10_2658, i_10_2700, i_10_2707, i_10_2715, i_10_2786, i_10_2788, i_10_2789, i_10_2824, i_10_2825, i_10_2959, i_10_2995, i_10_3094, i_10_3167, i_10_3238, i_10_3239, i_10_3269, i_10_3280, i_10_3281, i_10_3419, i_10_3434, i_10_3473, i_10_3505, i_10_3508, i_10_3526, i_10_3527, i_10_3587, i_10_3647, i_10_3848, i_10_3883, i_10_3913, i_10_3914, i_10_3950, i_10_3985, i_10_3991, i_10_3992, i_10_4004, i_10_4057, i_10_4113, i_10_4118, i_10_4120, i_10_4130, i_10_4168, i_10_4172, i_10_4174, i_10_4276, i_10_4279, i_10_4281, i_10_4454, i_10_4568, o_10_246);
	kernel_10_247 k_10_247(i_10_123, i_10_181, i_10_183, i_10_319, i_10_320, i_10_323, i_10_328, i_10_330, i_10_390, i_10_391, i_10_408, i_10_437, i_10_442, i_10_449, i_10_755, i_10_850, i_10_965, i_10_998, i_10_1031, i_10_1048, i_10_1240, i_10_1241, i_10_1264, i_10_1265, i_10_1268, i_10_1310, i_10_1345, i_10_1362, i_10_1363, i_10_1464, i_10_1555, i_10_1651, i_10_1653, i_10_1684, i_10_1687, i_10_1878, i_10_1915, i_10_1983, i_10_2056, i_10_2183, i_10_2200, i_10_2361, i_10_2464, i_10_2466, i_10_2471, i_10_2474, i_10_2505, i_10_2508, i_10_2509, i_10_2515, i_10_2632, i_10_2634, i_10_2635, i_10_2636, i_10_2655, i_10_2661, i_10_2679, i_10_2681, i_10_2705, i_10_2706, i_10_2711, i_10_2716, i_10_2718, i_10_2719, i_10_2728, i_10_2734, i_10_2787, i_10_2826, i_10_2833, i_10_2886, i_10_2923, i_10_3036, i_10_3074, i_10_3075, i_10_3076, i_10_3077, i_10_3165, i_10_3280, i_10_3283, i_10_3315, i_10_3385, i_10_3388, i_10_3617, i_10_3808, i_10_3848, i_10_3860, i_10_3892, i_10_3894, i_10_3982, i_10_4118, i_10_4119, i_10_4130, i_10_4219, i_10_4261, i_10_4279, i_10_4289, i_10_4566, i_10_4585, i_10_4586, i_10_4598, o_10_247);
	kernel_10_248 k_10_248(i_10_123, i_10_124, i_10_149, i_10_220, i_10_245, i_10_265, i_10_282, i_10_286, i_10_326, i_10_329, i_10_447, i_10_448, i_10_449, i_10_459, i_10_467, i_10_515, i_10_518, i_10_599, i_10_713, i_10_715, i_10_716, i_10_751, i_10_755, i_10_796, i_10_964, i_10_965, i_10_1004, i_10_1239, i_10_1266, i_10_1384, i_10_1583, i_10_1634, i_10_1726, i_10_1764, i_10_1822, i_10_1916, i_10_1945, i_10_1991, i_10_2255, i_10_2349, i_10_2353, i_10_2354, i_10_2377, i_10_2378, i_10_2453, i_10_2455, i_10_2469, i_10_2471, i_10_2504, i_10_2512, i_10_2605, i_10_2606, i_10_2633, i_10_2657, i_10_2663, i_10_2710, i_10_2714, i_10_2728, i_10_2729, i_10_2818, i_10_2918, i_10_2920, i_10_2980, i_10_2982, i_10_3043, i_10_3044, i_10_3047, i_10_3070, i_10_3275, i_10_3279, i_10_3391, i_10_3467, i_10_3473, i_10_3589, i_10_3590, i_10_3609, i_10_3649, i_10_3650, i_10_3652, i_10_3653, i_10_3781, i_10_3786, i_10_3809, i_10_3835, i_10_3842, i_10_3845, i_10_3854, i_10_3875, i_10_3947, i_10_4115, i_10_4117, i_10_4119, i_10_4121, i_10_4124, i_10_4214, i_10_4269, i_10_4285, i_10_4287, i_10_4460, i_10_4569, o_10_248);
	kernel_10_249 k_10_249(i_10_221, i_10_280, i_10_282, i_10_283, i_10_284, i_10_286, i_10_287, i_10_433, i_10_435, i_10_436, i_10_441, i_10_442, i_10_445, i_10_446, i_10_448, i_10_466, i_10_507, i_10_510, i_10_755, i_10_793, i_10_794, i_10_798, i_10_902, i_10_957, i_10_958, i_10_961, i_10_1032, i_10_1033, i_10_1237, i_10_1240, i_10_1241, i_10_1365, i_10_1366, i_10_1545, i_10_1578, i_10_1648, i_10_1649, i_10_1650, i_10_1651, i_10_1654, i_10_1686, i_10_1687, i_10_1689, i_10_1819, i_10_1824, i_10_1825, i_10_1909, i_10_1915, i_10_1990, i_10_2312, i_10_2338, i_10_2354, i_10_2366, i_10_2380, i_10_2382, i_10_2454, i_10_2457, i_10_2460, i_10_2461, i_10_2662, i_10_2679, i_10_2703, i_10_2704, i_10_2706, i_10_2707, i_10_2708, i_10_2719, i_10_2731, i_10_2783, i_10_2827, i_10_2830, i_10_2831, i_10_2832, i_10_2833, i_10_2919, i_10_2923, i_10_3038, i_10_3158, i_10_3271, i_10_3387, i_10_3388, i_10_3389, i_10_3391, i_10_3392, i_10_3406, i_10_3472, i_10_3588, i_10_3616, i_10_3783, i_10_3786, i_10_3787, i_10_3838, i_10_3840, i_10_3841, i_10_3847, i_10_3855, i_10_3860, i_10_4118, i_10_4121, i_10_4274, o_10_249);
	kernel_10_250 k_10_250(i_10_157, i_10_174, i_10_248, i_10_273, i_10_274, i_10_277, i_10_285, i_10_286, i_10_324, i_10_428, i_10_436, i_10_439, i_10_467, i_10_793, i_10_796, i_10_959, i_10_967, i_10_968, i_10_995, i_10_999, i_10_1027, i_10_1033, i_10_1217, i_10_1241, i_10_1245, i_10_1250, i_10_1306, i_10_1309, i_10_1310, i_10_1313, i_10_1432, i_10_1444, i_10_1647, i_10_1649, i_10_1945, i_10_1949, i_10_1950, i_10_2019, i_10_2308, i_10_2327, i_10_2350, i_10_2452, i_10_2471, i_10_2508, i_10_2509, i_10_2541, i_10_2542, i_10_2628, i_10_2629, i_10_2630, i_10_2633, i_10_2635, i_10_2657, i_10_2663, i_10_2713, i_10_2734, i_10_2735, i_10_2785, i_10_2828, i_10_2830, i_10_2920, i_10_3033, i_10_3037, i_10_3038, i_10_3092, i_10_3268, i_10_3271, i_10_3281, i_10_3384, i_10_3385, i_10_3388, i_10_3433, i_10_3465, i_10_3472, i_10_3586, i_10_3587, i_10_3613, i_10_3614, i_10_3616, i_10_3626, i_10_3646, i_10_3647, i_10_3649, i_10_3650, i_10_3836, i_10_3838, i_10_3839, i_10_3846, i_10_3847, i_10_3848, i_10_3857, i_10_3890, i_10_3980, i_10_3988, i_10_3994, i_10_4055, i_10_4114, i_10_4116, i_10_4118, i_10_4284, o_10_250);
	kernel_10_251 k_10_251(i_10_124, i_10_222, i_10_246, i_10_247, i_10_249, i_10_250, i_10_280, i_10_315, i_10_317, i_10_327, i_10_329, i_10_331, i_10_395, i_10_406, i_10_409, i_10_751, i_10_797, i_10_955, i_10_956, i_10_993, i_10_1040, i_10_1129, i_10_1234, i_10_1235, i_10_1238, i_10_1241, i_10_1244, i_10_1246, i_10_1264, i_10_1309, i_10_1341, i_10_1363, i_10_1579, i_10_1600, i_10_1651, i_10_1686, i_10_1689, i_10_1819, i_10_1824, i_10_1950, i_10_2182, i_10_2203, i_10_2350, i_10_2353, i_10_2354, i_10_2356, i_10_2357, i_10_2361, i_10_2364, i_10_2365, i_10_2366, i_10_2454, i_10_2455, i_10_2456, i_10_2461, i_10_2721, i_10_2722, i_10_2723, i_10_2725, i_10_2728, i_10_2885, i_10_2888, i_10_2916, i_10_2922, i_10_2923, i_10_3034, i_10_3038, i_10_3043, i_10_3202, i_10_3203, i_10_3275, i_10_3281, i_10_3284, i_10_3386, i_10_3389, i_10_3392, i_10_3542, i_10_3586, i_10_3589, i_10_3616, i_10_3617, i_10_3653, i_10_3780, i_10_3781, i_10_3785, i_10_3788, i_10_3808, i_10_3814, i_10_3844, i_10_3845, i_10_3848, i_10_3858, i_10_3914, i_10_3983, i_10_4117, i_10_4120, i_10_4286, i_10_4288, i_10_4289, i_10_4563, o_10_251);
	kernel_10_252 k_10_252(i_10_150, i_10_175, i_10_183, i_10_219, i_10_220, i_10_224, i_10_260, i_10_281, i_10_286, i_10_319, i_10_320, i_10_409, i_10_432, i_10_435, i_10_436, i_10_441, i_10_444, i_10_445, i_10_448, i_10_461, i_10_462, i_10_519, i_10_697, i_10_795, i_10_796, i_10_898, i_10_966, i_10_967, i_10_1033, i_10_1237, i_10_1238, i_10_1241, i_10_1243, i_10_1305, i_10_1308, i_10_1309, i_10_1437, i_10_1650, i_10_1651, i_10_1681, i_10_1682, i_10_1819, i_10_1821, i_10_1822, i_10_1825, i_10_2182, i_10_2331, i_10_2334, i_10_2382, i_10_2384, i_10_2405, i_10_2452, i_10_2453, i_10_2455, i_10_2631, i_10_2635, i_10_2658, i_10_2659, i_10_2660, i_10_2710, i_10_2733, i_10_2831, i_10_2919, i_10_2920, i_10_3036, i_10_3037, i_10_3045, i_10_3046, i_10_3150, i_10_3153, i_10_3165, i_10_3166, i_10_3270, i_10_3274, i_10_3278, i_10_3280, i_10_3281, i_10_3326, i_10_3469, i_10_3583, i_10_3649, i_10_3781, i_10_3846, i_10_3847, i_10_3853, i_10_3858, i_10_3912, i_10_3915, i_10_3980, i_10_3985, i_10_4116, i_10_4118, i_10_4120, i_10_4219, i_10_4269, i_10_4271, i_10_4283, i_10_4564, i_10_4566, i_10_4567, o_10_252);
	kernel_10_253 k_10_253(i_10_88, i_10_148, i_10_217, i_10_269, i_10_408, i_10_424, i_10_434, i_10_435, i_10_441, i_10_442, i_10_459, i_10_533, i_10_559, i_10_733, i_10_794, i_10_990, i_10_1036, i_10_1085, i_10_1164, i_10_1222, i_10_1234, i_10_1241, i_10_1309, i_10_1310, i_10_1341, i_10_1384, i_10_1552, i_10_1579, i_10_1580, i_10_1582, i_10_1687, i_10_1688, i_10_1737, i_10_1806, i_10_1818, i_10_1819, i_10_2016, i_10_2206, i_10_2250, i_10_2355, i_10_2356, i_10_2364, i_10_2389, i_10_2451, i_10_2469, i_10_2470, i_10_2515, i_10_2563, i_10_2602, i_10_2604, i_10_2606, i_10_2628, i_10_2629, i_10_2701, i_10_2711, i_10_2725, i_10_2782, i_10_2789, i_10_2817, i_10_2820, i_10_2841, i_10_2862, i_10_2863, i_10_2883, i_10_2884, i_10_2921, i_10_3048, i_10_3124, i_10_3200, i_10_3268, i_10_3269, i_10_3277, i_10_3295, i_10_3297, i_10_3357, i_10_3384, i_10_3387, i_10_3388, i_10_3389, i_10_3408, i_10_3430, i_10_3520, i_10_3544, i_10_3610, i_10_3612, i_10_3640, i_10_3649, i_10_3808, i_10_3835, i_10_3855, i_10_3889, i_10_3920, i_10_3981, i_10_3991, i_10_4129, i_10_4272, i_10_4273, i_10_4281, i_10_4290, i_10_4292, o_10_253);
	kernel_10_254 k_10_254(i_10_40, i_10_41, i_10_175, i_10_185, i_10_197, i_10_251, i_10_268, i_10_269, i_10_280, i_10_286, i_10_319, i_10_320, i_10_410, i_10_447, i_10_462, i_10_463, i_10_533, i_10_697, i_10_700, i_10_701, i_10_737, i_10_794, i_10_995, i_10_997, i_10_998, i_10_1003, i_10_1043, i_10_1088, i_10_1236, i_10_1237, i_10_1240, i_10_1349, i_10_1445, i_10_1582, i_10_1601, i_10_1653, i_10_1654, i_10_1655, i_10_1685, i_10_1817, i_10_1823, i_10_1946, i_10_1949, i_10_2006, i_10_2158, i_10_2311, i_10_2334, i_10_2339, i_10_2355, i_10_2383, i_10_2384, i_10_2453, i_10_2470, i_10_2471, i_10_2510, i_10_2635, i_10_2636, i_10_2680, i_10_2681, i_10_2707, i_10_2729, i_10_2786, i_10_2825, i_10_2828, i_10_2830, i_10_2883, i_10_2887, i_10_2983, i_10_2985, i_10_3038, i_10_3073, i_10_3076, i_10_3196, i_10_3274, i_10_3284, i_10_3290, i_10_3302, i_10_3409, i_10_3410, i_10_3472, i_10_3611, i_10_3616, i_10_3649, i_10_3650, i_10_3688, i_10_3784, i_10_3837, i_10_3853, i_10_3854, i_10_3857, i_10_3859, i_10_3896, i_10_3919, i_10_3985, i_10_3986, i_10_3991, i_10_3994, i_10_4220, i_10_4283, i_10_4289, o_10_254);
	kernel_10_255 k_10_255(i_10_35, i_10_175, i_10_176, i_10_218, i_10_223, i_10_282, i_10_410, i_10_444, i_10_460, i_10_462, i_10_463, i_10_464, i_10_798, i_10_799, i_10_969, i_10_970, i_10_994, i_10_1005, i_10_1030, i_10_1138, i_10_1236, i_10_1237, i_10_1238, i_10_1260, i_10_1305, i_10_1309, i_10_1310, i_10_1362, i_10_1654, i_10_1686, i_10_1687, i_10_1819, i_10_1820, i_10_1823, i_10_1909, i_10_1911, i_10_1944, i_10_1989, i_10_1990, i_10_2180, i_10_2183, i_10_2305, i_10_2310, i_10_2409, i_10_2450, i_10_2472, i_10_2632, i_10_2657, i_10_2659, i_10_2701, i_10_2711, i_10_2713, i_10_2727, i_10_2785, i_10_2830, i_10_2833, i_10_2881, i_10_2883, i_10_2885, i_10_2920, i_10_3034, i_10_3036, i_10_3037, i_10_3038, i_10_3039, i_10_3040, i_10_3069, i_10_3199, i_10_3200, i_10_3323, i_10_3386, i_10_3389, i_10_3403, i_10_3405, i_10_3406, i_10_3585, i_10_3588, i_10_3590, i_10_3649, i_10_3652, i_10_3653, i_10_3835, i_10_3842, i_10_3846, i_10_3848, i_10_3857, i_10_3882, i_10_3981, i_10_3982, i_10_3985, i_10_4116, i_10_4118, i_10_4125, i_10_4126, i_10_4127, i_10_4218, i_10_4269, i_10_4273, i_10_4289, i_10_4566, o_10_255);
	kernel_10_256 k_10_256(i_10_41, i_10_255, i_10_282, i_10_409, i_10_423, i_10_430, i_10_431, i_10_436, i_10_444, i_10_445, i_10_446, i_10_447, i_10_448, i_10_466, i_10_716, i_10_794, i_10_796, i_10_800, i_10_967, i_10_968, i_10_969, i_10_970, i_10_1240, i_10_1241, i_10_1243, i_10_1266, i_10_1365, i_10_1452, i_10_1453, i_10_1548, i_10_1580, i_10_1582, i_10_1583, i_10_1629, i_10_1650, i_10_1651, i_10_1655, i_10_1683, i_10_1690, i_10_1691, i_10_2203, i_10_2352, i_10_2362, i_10_2363, i_10_2364, i_10_2365, i_10_2366, i_10_2376, i_10_2410, i_10_2411, i_10_2469, i_10_2470, i_10_2472, i_10_2473, i_10_2474, i_10_2631, i_10_2632, i_10_2659, i_10_2660, i_10_2661, i_10_2662, i_10_2663, i_10_2702, i_10_2716, i_10_2734, i_10_2735, i_10_2831, i_10_2832, i_10_2982, i_10_3049, i_10_3087, i_10_3165, i_10_3385, i_10_3386, i_10_3388, i_10_3389, i_10_3390, i_10_3391, i_10_3392, i_10_3468, i_10_3469, i_10_3470, i_10_3586, i_10_3587, i_10_3588, i_10_3589, i_10_3590, i_10_3783, i_10_3784, i_10_3787, i_10_3834, i_10_3843, i_10_4058, i_10_4116, i_10_4117, i_10_4119, i_10_4165, i_10_4270, i_10_4365, i_10_4585, o_10_256);
	kernel_10_257 k_10_257(i_10_149, i_10_174, i_10_175, i_10_177, i_10_178, i_10_183, i_10_184, i_10_185, i_10_187, i_10_286, i_10_319, i_10_328, i_10_329, i_10_408, i_10_409, i_10_410, i_10_442, i_10_463, i_10_510, i_10_753, i_10_754, i_10_796, i_10_967, i_10_1032, i_10_1042, i_10_1043, i_10_1169, i_10_1250, i_10_1263, i_10_1582, i_10_1651, i_10_1652, i_10_1653, i_10_1654, i_10_1655, i_10_1684, i_10_1821, i_10_1822, i_10_1824, i_10_1825, i_10_1826, i_10_1910, i_10_1952, i_10_2185, i_10_2307, i_10_2352, i_10_2353, i_10_2354, i_10_2355, i_10_2410, i_10_2452, i_10_2454, i_10_2470, i_10_2473, i_10_2474, i_10_2608, i_10_2701, i_10_2704, i_10_2713, i_10_2716, i_10_2735, i_10_2833, i_10_2916, i_10_2919, i_10_2920, i_10_2921, i_10_2980, i_10_2985, i_10_3035, i_10_3050, i_10_3152, i_10_3162, i_10_3271, i_10_3279, i_10_3280, i_10_3387, i_10_3388, i_10_3390, i_10_3391, i_10_3405, i_10_3472, i_10_3611, i_10_3613, i_10_3614, i_10_3615, i_10_3646, i_10_3647, i_10_3653, i_10_3725, i_10_3834, i_10_3837, i_10_3840, i_10_3857, i_10_3895, i_10_3990, i_10_3991, i_10_4115, i_10_4182, i_10_4189, i_10_4282, o_10_257);
	kernel_10_258 k_10_258(i_10_177, i_10_252, i_10_282, i_10_284, i_10_290, i_10_324, i_10_370, i_10_430, i_10_438, i_10_442, i_10_464, i_10_504, i_10_595, i_10_717, i_10_793, i_10_891, i_10_999, i_10_1000, i_10_1053, i_10_1245, i_10_1313, i_10_1443, i_10_1445, i_10_1654, i_10_1655, i_10_1719, i_10_1809, i_10_1819, i_10_1824, i_10_1825, i_10_1948, i_10_1990, i_10_1991, i_10_2181, i_10_2184, i_10_2245, i_10_2322, i_10_2331, i_10_2353, i_10_2356, i_10_2361, i_10_2379, i_10_2380, i_10_2453, i_10_2461, i_10_2566, i_10_2638, i_10_2680, i_10_2700, i_10_2704, i_10_2709, i_10_2881, i_10_2882, i_10_2885, i_10_2953, i_10_3033, i_10_3042, i_10_3043, i_10_3044, i_10_3045, i_10_3156, i_10_3196, i_10_3200, i_10_3267, i_10_3268, i_10_3277, i_10_3280, i_10_3288, i_10_3385, i_10_3386, i_10_3406, i_10_3465, i_10_3468, i_10_3495, i_10_3496, i_10_3525, i_10_3609, i_10_3610, i_10_3617, i_10_3647, i_10_3651, i_10_3780, i_10_3785, i_10_3836, i_10_3837, i_10_3851, i_10_3856, i_10_3859, i_10_4113, i_10_4122, i_10_4123, i_10_4126, i_10_4213, i_10_4231, i_10_4269, i_10_4290, i_10_4564, i_10_4566, i_10_4567, i_10_4568, o_10_258);
	kernel_10_259 k_10_259(i_10_119, i_10_174, i_10_331, i_10_332, i_10_361, i_10_409, i_10_446, i_10_519, i_10_895, i_10_906, i_10_951, i_10_1039, i_10_1041, i_10_1042, i_10_1122, i_10_1204, i_10_1241, i_10_1266, i_10_1267, i_10_1271, i_10_1308, i_10_1309, i_10_1311, i_10_1312, i_10_1353, i_10_1354, i_10_1546, i_10_1647, i_10_1651, i_10_1654, i_10_1824, i_10_1911, i_10_1912, i_10_1950, i_10_2002, i_10_2326, i_10_2355, i_10_2356, i_10_2357, i_10_2454, i_10_2467, i_10_2515, i_10_2607, i_10_2630, i_10_2632, i_10_2655, i_10_2656, i_10_2676, i_10_2679, i_10_2703, i_10_2704, i_10_2722, i_10_2733, i_10_2784, i_10_2788, i_10_2820, i_10_2823, i_10_2833, i_10_2834, i_10_2883, i_10_2919, i_10_2955, i_10_2985, i_10_2986, i_10_3088, i_10_3163, i_10_3272, i_10_3297, i_10_3388, i_10_3406, i_10_3407, i_10_3433, i_10_3434, i_10_3450, i_10_3496, i_10_3614, i_10_3700, i_10_3723, i_10_3834, i_10_3852, i_10_3859, i_10_3860, i_10_3894, i_10_3895, i_10_3896, i_10_3964, i_10_3980, i_10_3981, i_10_3982, i_10_3987, i_10_4116, i_10_4129, i_10_4130, i_10_4281, i_10_4282, i_10_4285, i_10_4288, i_10_4291, i_10_4292, i_10_4579, o_10_259);
	kernel_10_260 k_10_260(i_10_28, i_10_55, i_10_56, i_10_250, i_10_251, i_10_282, i_10_294, i_10_321, i_10_322, i_10_430, i_10_431, i_10_463, i_10_517, i_10_593, i_10_706, i_10_797, i_10_799, i_10_876, i_10_898, i_10_906, i_10_921, i_10_930, i_10_945, i_10_969, i_10_1029, i_10_1165, i_10_1237, i_10_1238, i_10_1239, i_10_1347, i_10_1364, i_10_1369, i_10_1385, i_10_1489, i_10_1543, i_10_1546, i_10_1547, i_10_1628, i_10_1630, i_10_1695, i_10_1718, i_10_1908, i_10_1996, i_10_2023, i_10_2326, i_10_2353, i_10_2356, i_10_2357, i_10_2568, i_10_2571, i_10_2608, i_10_2609, i_10_2632, i_10_2679, i_10_2691, i_10_2694, i_10_2695, i_10_2710, i_10_2716, i_10_2782, i_10_2788, i_10_2789, i_10_2828, i_10_2830, i_10_2850, i_10_2851, i_10_2921, i_10_2982, i_10_3072, i_10_3073, i_10_3076, i_10_3093, i_10_3271, i_10_3293, i_10_3301, i_10_3359, i_10_3390, i_10_3391, i_10_3434, i_10_3561, i_10_3582, i_10_3583, i_10_3590, i_10_3784, i_10_3813, i_10_3815, i_10_3855, i_10_3856, i_10_3877, i_10_3889, i_10_3945, i_10_4031, i_10_4119, i_10_4173, i_10_4236, i_10_4266, i_10_4278, i_10_4281, i_10_4461, i_10_4566, o_10_260);
	kernel_10_261 k_10_261(i_10_123, i_10_148, i_10_178, i_10_267, i_10_277, i_10_282, i_10_283, i_10_292, i_10_408, i_10_510, i_10_520, i_10_663, i_10_1005, i_10_1006, i_10_1236, i_10_1266, i_10_1309, i_10_1312, i_10_1437, i_10_1438, i_10_1546, i_10_1552, i_10_1555, i_10_1579, i_10_1626, i_10_1689, i_10_1716, i_10_1734, i_10_1735, i_10_1806, i_10_1951, i_10_1992, i_10_2031, i_10_2311, i_10_2353, i_10_2355, i_10_2356, i_10_2408, i_10_2453, i_10_2469, i_10_2472, i_10_2571, i_10_2632, i_10_2662, i_10_2663, i_10_2715, i_10_2716, i_10_2730, i_10_2731, i_10_2734, i_10_2785, i_10_2827, i_10_2850, i_10_2884, i_10_2887, i_10_2922, i_10_2967, i_10_2985, i_10_3045, i_10_3072, i_10_3075, i_10_3196, i_10_3199, i_10_3201, i_10_3278, i_10_3279, i_10_3283, i_10_3318, i_10_3386, i_10_3391, i_10_3471, i_10_3507, i_10_3525, i_10_3540, i_10_3585, i_10_3613, i_10_3616, i_10_3688, i_10_3782, i_10_3783, i_10_3784, i_10_3787, i_10_3811, i_10_3837, i_10_3838, i_10_3846, i_10_3859, i_10_3909, i_10_3985, i_10_4056, i_10_4116, i_10_4117, i_10_4120, i_10_4121, i_10_4173, i_10_4272, i_10_4273, i_10_4281, i_10_4282, i_10_4290, o_10_261);
	kernel_10_262 k_10_262(i_10_319, i_10_390, i_10_408, i_10_409, i_10_410, i_10_411, i_10_413, i_10_441, i_10_444, i_10_499, i_10_586, i_10_736, i_10_737, i_10_797, i_10_853, i_10_931, i_10_1034, i_10_1119, i_10_1181, i_10_1239, i_10_1240, i_10_1241, i_10_1276, i_10_1308, i_10_1347, i_10_1438, i_10_1439, i_10_1545, i_10_1552, i_10_1579, i_10_1583, i_10_1650, i_10_1651, i_10_1766, i_10_1804, i_10_1807, i_10_1819, i_10_1821, i_10_1822, i_10_2200, i_10_2223, i_10_2355, i_10_2356, i_10_2380, i_10_2389, i_10_2391, i_10_2392, i_10_2410, i_10_2435, i_10_2441, i_10_2443, i_10_2444, i_10_2450, i_10_2452, i_10_2459, i_10_2635, i_10_2650, i_10_2658, i_10_2660, i_10_2679, i_10_2695, i_10_2704, i_10_2716, i_10_2733, i_10_2734, i_10_2784, i_10_2821, i_10_2884, i_10_2888, i_10_2983, i_10_3072, i_10_3075, i_10_3076, i_10_3117, i_10_3166, i_10_3202, i_10_3468, i_10_3471, i_10_3539, i_10_3541, i_10_3544, i_10_3609, i_10_3684, i_10_3775, i_10_3805, i_10_3840, i_10_3846, i_10_3857, i_10_3893, i_10_4013, i_10_4173, i_10_4175, i_10_4182, i_10_4475, i_10_4524, i_10_4563, i_10_4564, i_10_4568, i_10_4588, i_10_4598, o_10_262);
	kernel_10_263 k_10_263(i_10_243, i_10_283, i_10_444, i_10_459, i_10_460, i_10_464, i_10_751, i_10_793, i_10_795, i_10_966, i_10_968, i_10_999, i_10_1000, i_10_1041, i_10_1235, i_10_1236, i_10_1243, i_10_1246, i_10_1247, i_10_1249, i_10_1445, i_10_1539, i_10_1541, i_10_1819, i_10_1821, i_10_1823, i_10_1911, i_10_1912, i_10_1913, i_10_2004, i_10_2179, i_10_2180, i_10_2354, i_10_2377, i_10_2467, i_10_2473, i_10_2628, i_10_2630, i_10_2631, i_10_2634, i_10_2655, i_10_2657, i_10_2658, i_10_2660, i_10_2680, i_10_2681, i_10_2700, i_10_2701, i_10_2720, i_10_2721, i_10_2722, i_10_2727, i_10_2728, i_10_2732, i_10_2733, i_10_2735, i_10_2818, i_10_2827, i_10_2829, i_10_2830, i_10_2833, i_10_2883, i_10_2884, i_10_2919, i_10_2920, i_10_3034, i_10_3038, i_10_3069, i_10_3070, i_10_3071, i_10_3087, i_10_3198, i_10_3268, i_10_3270, i_10_3385, i_10_3388, i_10_3389, i_10_3469, i_10_3537, i_10_3589, i_10_3612, i_10_3681, i_10_3687, i_10_3781, i_10_3787, i_10_3852, i_10_3853, i_10_3854, i_10_3860, i_10_3888, i_10_3889, i_10_3912, i_10_3978, i_10_3990, i_10_3991, i_10_4266, i_10_4267, i_10_4290, i_10_4429, i_10_4571, o_10_263);
	kernel_10_264 k_10_264(i_10_155, i_10_177, i_10_220, i_10_223, i_10_224, i_10_247, i_10_249, i_10_272, i_10_281, i_10_290, i_10_291, i_10_292, i_10_318, i_10_326, i_10_329, i_10_406, i_10_407, i_10_408, i_10_497, i_10_593, i_10_797, i_10_830, i_10_832, i_10_833, i_10_896, i_10_899, i_10_931, i_10_954, i_10_955, i_10_957, i_10_1057, i_10_1121, i_10_1264, i_10_1273, i_10_1305, i_10_1308, i_10_1345, i_10_1363, i_10_1364, i_10_1367, i_10_1444, i_10_1648, i_10_1651, i_10_1688, i_10_1724, i_10_1765, i_10_1913, i_10_1921, i_10_1996, i_10_1997, i_10_2023, i_10_2255, i_10_2310, i_10_2351, i_10_2362, i_10_2365, i_10_2452, i_10_2516, i_10_2518, i_10_2655, i_10_2656, i_10_2657, i_10_2714, i_10_2718, i_10_2719, i_10_2720, i_10_2731, i_10_2782, i_10_2784, i_10_2787, i_10_2884, i_10_2984, i_10_3047, i_10_3050, i_10_3077, i_10_3092, i_10_3281, i_10_3290, i_10_3302, i_10_3356, i_10_3406, i_10_3407, i_10_3494, i_10_3497, i_10_3526, i_10_3527, i_10_3542, i_10_3641, i_10_3688, i_10_3780, i_10_3852, i_10_3854, i_10_3984, i_10_3995, i_10_4054, i_10_4055, i_10_4121, i_10_4171, i_10_4237, i_10_4268, o_10_264);
	kernel_10_265 k_10_265(i_10_210, i_10_277, i_10_279, i_10_280, i_10_287, i_10_444, i_10_447, i_10_499, i_10_517, i_10_586, i_10_587, i_10_607, i_10_792, i_10_793, i_10_796, i_10_798, i_10_799, i_10_904, i_10_1049, i_10_1123, i_10_1164, i_10_1171, i_10_1200, i_10_1201, i_10_1234, i_10_1305, i_10_1362, i_10_1444, i_10_1447, i_10_1448, i_10_1602, i_10_1651, i_10_1652, i_10_1732, i_10_1818, i_10_1822, i_10_1881, i_10_1882, i_10_2155, i_10_2329, i_10_2338, i_10_2362, i_10_2382, i_10_2448, i_10_2449, i_10_2451, i_10_2475, i_10_2543, i_10_2659, i_10_2660, i_10_2662, i_10_2663, i_10_2728, i_10_2731, i_10_2814, i_10_2888, i_10_2916, i_10_2917, i_10_2919, i_10_2922, i_10_2979, i_10_3039, i_10_3047, i_10_3049, i_10_3050, i_10_3092, i_10_3109, i_10_3169, i_10_3172, i_10_3282, i_10_3294, i_10_3388, i_10_3496, i_10_3615, i_10_3684, i_10_3720, i_10_3721, i_10_3729, i_10_3787, i_10_3851, i_10_3854, i_10_3859, i_10_3892, i_10_3919, i_10_3950, i_10_4024, i_10_4117, i_10_4170, i_10_4189, i_10_4277, i_10_4290, i_10_4326, i_10_4354, i_10_4371, i_10_4449, i_10_4476, i_10_4477, i_10_4539, i_10_4575, i_10_4593, o_10_265);
	kernel_10_266 k_10_266(i_10_33, i_10_39, i_10_69, i_10_144, i_10_146, i_10_178, i_10_248, i_10_257, i_10_271, i_10_282, i_10_406, i_10_429, i_10_445, i_10_502, i_10_520, i_10_561, i_10_585, i_10_598, i_10_642, i_10_730, i_10_731, i_10_733, i_10_734, i_10_737, i_10_832, i_10_847, i_10_848, i_10_1003, i_10_1039, i_10_1233, i_10_1234, i_10_1239, i_10_1268, i_10_1307, i_10_1347, i_10_1353, i_10_1365, i_10_1441, i_10_1442, i_10_1611, i_10_1650, i_10_1697, i_10_1717, i_10_1824, i_10_1825, i_10_1872, i_10_1942, i_10_2079, i_10_2179, i_10_2206, i_10_2376, i_10_2379, i_10_2434, i_10_2452, i_10_2457, i_10_2463, i_10_2471, i_10_2504, i_10_2602, i_10_2617, i_10_2632, i_10_2658, i_10_2724, i_10_2730, i_10_2789, i_10_2829, i_10_2869, i_10_2920, i_10_2922, i_10_3038, i_10_3076, i_10_3097, i_10_3098, i_10_3101, i_10_3198, i_10_3201, i_10_3203, i_10_3282, i_10_3351, i_10_3469, i_10_3472, i_10_3473, i_10_3496, i_10_3525, i_10_3612, i_10_3650, i_10_3685, i_10_3717, i_10_3783, i_10_3786, i_10_3787, i_10_3788, i_10_3810, i_10_3834, i_10_3835, i_10_3857, i_10_4054, i_10_4101, i_10_4279, i_10_4563, o_10_266);
	kernel_10_267 k_10_267(i_10_34, i_10_85, i_10_86, i_10_89, i_10_121, i_10_151, i_10_172, i_10_249, i_10_283, i_10_330, i_10_427, i_10_431, i_10_438, i_10_445, i_10_465, i_10_520, i_10_565, i_10_898, i_10_996, i_10_1003, i_10_1032, i_10_1033, i_10_1165, i_10_1166, i_10_1168, i_10_1173, i_10_1174, i_10_1233, i_10_1237, i_10_1239, i_10_1293, i_10_1365, i_10_1381, i_10_1488, i_10_1491, i_10_1536, i_10_1537, i_10_1583, i_10_1691, i_10_1821, i_10_1824, i_10_1997, i_10_2004, i_10_2352, i_10_2382, i_10_2391, i_10_2392, i_10_2463, i_10_2508, i_10_2542, i_10_2607, i_10_2634, i_10_2635, i_10_2653, i_10_2654, i_10_2660, i_10_2680, i_10_2703, i_10_2705, i_10_2724, i_10_2725, i_10_2729, i_10_2730, i_10_2731, i_10_2733, i_10_2734, i_10_2787, i_10_2828, i_10_2834, i_10_2920, i_10_2986, i_10_3120, i_10_3150, i_10_3151, i_10_3152, i_10_3162, i_10_3163, i_10_3165, i_10_3195, i_10_3202, i_10_3300, i_10_3496, i_10_3522, i_10_3616, i_10_3617, i_10_3688, i_10_3689, i_10_3733, i_10_3839, i_10_3846, i_10_3847, i_10_3856, i_10_4116, i_10_4117, i_10_4120, i_10_4128, i_10_4288, i_10_4290, i_10_4566, i_10_4567, o_10_267);
	kernel_10_268 k_10_268(i_10_34, i_10_42, i_10_51, i_10_52, i_10_53, i_10_142, i_10_151, i_10_177, i_10_184, i_10_287, i_10_294, i_10_321, i_10_430, i_10_431, i_10_445, i_10_447, i_10_464, i_10_465, i_10_637, i_10_699, i_10_834, i_10_897, i_10_934, i_10_957, i_10_961, i_10_966, i_10_971, i_10_1087, i_10_1236, i_10_1239, i_10_1241, i_10_1311, i_10_1543, i_10_1582, i_10_1583, i_10_1636, i_10_1645, i_10_1687, i_10_1688, i_10_1696, i_10_1725, i_10_1816, i_10_1823, i_10_1957, i_10_2040, i_10_2391, i_10_2471, i_10_2472, i_10_2535, i_10_2545, i_10_2632, i_10_2633, i_10_2679, i_10_2706, i_10_2707, i_10_2708, i_10_2716, i_10_2717, i_10_2730, i_10_2830, i_10_2913, i_10_3198, i_10_3238, i_10_3390, i_10_3468, i_10_3469, i_10_3495, i_10_3496, i_10_3497, i_10_3498, i_10_3500, i_10_3509, i_10_3541, i_10_3588, i_10_3648, i_10_3651, i_10_3783, i_10_3784, i_10_3785, i_10_3787, i_10_3846, i_10_3849, i_10_3851, i_10_3859, i_10_3886, i_10_3949, i_10_3999, i_10_4119, i_10_4121, i_10_4165, i_10_4242, i_10_4269, i_10_4270, i_10_4287, i_10_4462, i_10_4463, i_10_4566, i_10_4567, i_10_4570, i_10_4588, o_10_268);
	kernel_10_269 k_10_269(i_10_25, i_10_187, i_10_249, i_10_258, i_10_259, i_10_260, i_10_276, i_10_277, i_10_282, i_10_283, i_10_321, i_10_426, i_10_517, i_10_600, i_10_717, i_10_728, i_10_754, i_10_800, i_10_850, i_10_853, i_10_997, i_10_998, i_10_1033, i_10_1034, i_10_1124, i_10_1194, i_10_1195, i_10_1239, i_10_1240, i_10_1249, i_10_1250, i_10_1356, i_10_1515, i_10_1579, i_10_1583, i_10_1618, i_10_1619, i_10_1653, i_10_1654, i_10_1687, i_10_1688, i_10_1819, i_10_1820, i_10_1821, i_10_1823, i_10_1826, i_10_1833, i_10_1960, i_10_2352, i_10_2355, i_10_2356, i_10_2357, i_10_2436, i_10_2457, i_10_2458, i_10_2460, i_10_2509, i_10_2563, i_10_2634, i_10_2716, i_10_2823, i_10_2868, i_10_2887, i_10_2895, i_10_3192, i_10_3195, i_10_3273, i_10_3319, i_10_3391, i_10_3401, i_10_3434, i_10_3508, i_10_3562, i_10_3610, i_10_3651, i_10_3687, i_10_3775, i_10_3783, i_10_3787, i_10_3813, i_10_3814, i_10_3815, i_10_3846, i_10_3910, i_10_3946, i_10_3947, i_10_3948, i_10_4012, i_10_4013, i_10_4055, i_10_4117, i_10_4118, i_10_4171, i_10_4279, i_10_4280, i_10_4290, i_10_4291, i_10_4369, i_10_4461, i_10_4462, o_10_269);
	kernel_10_270 k_10_270(i_10_29, i_10_145, i_10_146, i_10_176, i_10_221, i_10_247, i_10_254, i_10_281, i_10_318, i_10_319, i_10_391, i_10_434, i_10_461, i_10_462, i_10_463, i_10_464, i_10_513, i_10_711, i_10_713, i_10_749, i_10_800, i_10_954, i_10_992, i_10_1027, i_10_1046, i_10_1049, i_10_1083, i_10_1220, i_10_1349, i_10_1361, i_10_1396, i_10_1397, i_10_1451, i_10_1539, i_10_1616, i_10_1622, i_10_1685, i_10_1821, i_10_1822, i_10_1954, i_10_1981, i_10_2066, i_10_2201, i_10_2349, i_10_2351, i_10_2353, i_10_2453, i_10_2471, i_10_2601, i_10_2612, i_10_2660, i_10_2701, i_10_2702, i_10_2704, i_10_2711, i_10_2722, i_10_2723, i_10_2783, i_10_2920, i_10_3038, i_10_3044, i_10_3196, i_10_3198, i_10_3199, i_10_3232, i_10_3278, i_10_3314, i_10_3388, i_10_3407, i_10_3503, i_10_3519, i_10_3520, i_10_3584, i_10_3586, i_10_3620, i_10_3645, i_10_3646, i_10_3683, i_10_3728, i_10_3783, i_10_3785, i_10_3837, i_10_3838, i_10_3839, i_10_3852, i_10_3859, i_10_3980, i_10_4115, i_10_4117, i_10_4126, i_10_4153, i_10_4171, i_10_4172, i_10_4275, i_10_4279, i_10_4280, i_10_4288, i_10_4289, i_10_4566, i_10_4568, o_10_270);
	kernel_10_271 k_10_271(i_10_161, i_10_175, i_10_183, i_10_187, i_10_220, i_10_246, i_10_248, i_10_251, i_10_268, i_10_279, i_10_285, i_10_410, i_10_431, i_10_446, i_10_462, i_10_463, i_10_464, i_10_465, i_10_466, i_10_467, i_10_754, i_10_755, i_10_799, i_10_995, i_10_997, i_10_1237, i_10_1238, i_10_1239, i_10_1240, i_10_1241, i_10_1312, i_10_1362, i_10_1363, i_10_1434, i_10_1436, i_10_1438, i_10_1439, i_10_1545, i_10_1654, i_10_1655, i_10_1685, i_10_1821, i_10_1825, i_10_1911, i_10_1912, i_10_2338, i_10_2339, i_10_2349, i_10_2350, i_10_2351, i_10_2356, i_10_2357, i_10_2361, i_10_2364, i_10_2383, i_10_2384, i_10_2455, i_10_2463, i_10_2464, i_10_2470, i_10_2609, i_10_2635, i_10_2636, i_10_2658, i_10_2662, i_10_2713, i_10_2732, i_10_2735, i_10_2916, i_10_2921, i_10_2985, i_10_2986, i_10_2987, i_10_3070, i_10_3151, i_10_3163, i_10_3195, i_10_3237, i_10_3238, i_10_3271, i_10_3275, i_10_3278, i_10_3390, i_10_3686, i_10_3837, i_10_3839, i_10_3840, i_10_3841, i_10_3852, i_10_3860, i_10_3892, i_10_4116, i_10_4117, i_10_4118, i_10_4121, i_10_4130, i_10_4269, i_10_4270, i_10_4288, i_10_4289, o_10_271);
	kernel_10_272 k_10_272(i_10_22, i_10_135, i_10_144, i_10_193, i_10_218, i_10_274, i_10_284, i_10_289, i_10_371, i_10_460, i_10_461, i_10_694, i_10_792, i_10_846, i_10_900, i_10_901, i_10_949, i_10_1280, i_10_1315, i_10_1360, i_10_1369, i_10_1370, i_10_1391, i_10_1441, i_10_1442, i_10_1479, i_10_1566, i_10_1567, i_10_1568, i_10_1651, i_10_1714, i_10_1818, i_10_1911, i_10_1924, i_10_1927, i_10_1930, i_10_1979, i_10_1984, i_10_2080, i_10_2089, i_10_2125, i_10_2151, i_10_2155, i_10_2269, i_10_2305, i_10_2306, i_10_2324, i_10_2350, i_10_2460, i_10_2475, i_10_2502, i_10_2503, i_10_2504, i_10_2506, i_10_2550, i_10_2629, i_10_2630, i_10_2677, i_10_2692, i_10_2729, i_10_2767, i_10_2803, i_10_2804, i_10_2953, i_10_2957, i_10_2959, i_10_3025, i_10_3026, i_10_3029, i_10_3096, i_10_3097, i_10_3214, i_10_3258, i_10_3298, i_10_3321, i_10_3357, i_10_3358, i_10_3540, i_10_3602, i_10_3651, i_10_3802, i_10_3838, i_10_3848, i_10_3979, i_10_3980, i_10_3994, i_10_4068, i_10_4089, i_10_4090, i_10_4114, i_10_4230, i_10_4266, i_10_4270, i_10_4279, i_10_4280, i_10_4357, i_10_4358, i_10_4403, i_10_4433, i_10_4440, o_10_272);
	kernel_10_273 k_10_273(i_10_281, i_10_282, i_10_283, i_10_296, i_10_327, i_10_328, i_10_408, i_10_411, i_10_413, i_10_425, i_10_443, i_10_712, i_10_748, i_10_800, i_10_1134, i_10_1235, i_10_1240, i_10_1248, i_10_1263, i_10_1264, i_10_1309, i_10_1366, i_10_1445, i_10_1580, i_10_1649, i_10_1819, i_10_1821, i_10_1823, i_10_1824, i_10_1876, i_10_1910, i_10_1911, i_10_1912, i_10_1913, i_10_1948, i_10_1989, i_10_2180, i_10_2186, i_10_2353, i_10_2354, i_10_2362, i_10_2380, i_10_2453, i_10_2468, i_10_2632, i_10_2634, i_10_2635, i_10_2636, i_10_2659, i_10_2660, i_10_2677, i_10_2711, i_10_2718, i_10_2719, i_10_2721, i_10_2722, i_10_2731, i_10_2781, i_10_2916, i_10_2921, i_10_2979, i_10_2980, i_10_2981, i_10_3033, i_10_3034, i_10_3035, i_10_3039, i_10_3040, i_10_3069, i_10_3196, i_10_3281, i_10_3283, i_10_3284, i_10_3324, i_10_3384, i_10_3388, i_10_3389, i_10_3392, i_10_3406, i_10_3437, i_10_3519, i_10_3520, i_10_3523, i_10_3613, i_10_3649, i_10_3650, i_10_3835, i_10_3849, i_10_3850, i_10_3855, i_10_3856, i_10_3857, i_10_3859, i_10_3906, i_10_3991, i_10_4114, i_10_4121, i_10_4563, i_10_4566, i_10_4568, o_10_273);
	kernel_10_274 k_10_274(i_10_27, i_10_28, i_10_29, i_10_117, i_10_118, i_10_119, i_10_122, i_10_153, i_10_174, i_10_279, i_10_280, i_10_286, i_10_316, i_10_462, i_10_464, i_10_514, i_10_559, i_10_793, i_10_958, i_10_1235, i_10_1240, i_10_1242, i_10_1309, i_10_1310, i_10_1549, i_10_1652, i_10_1686, i_10_1687, i_10_1820, i_10_1822, i_10_2018, i_10_2026, i_10_2029, i_10_2179, i_10_2180, i_10_2200, i_10_2350, i_10_2352, i_10_2380, i_10_2449, i_10_2452, i_10_2453, i_10_2466, i_10_2467, i_10_2470, i_10_2471, i_10_2502, i_10_2610, i_10_2628, i_10_2631, i_10_2659, i_10_2663, i_10_2700, i_10_2701, i_10_2719, i_10_2782, i_10_2827, i_10_2919, i_10_3036, i_10_3037, i_10_3088, i_10_3089, i_10_3155, i_10_3200, i_10_3385, i_10_3390, i_10_3519, i_10_3520, i_10_3525, i_10_3583, i_10_3586, i_10_3587, i_10_3613, i_10_3646, i_10_3649, i_10_3785, i_10_3837, i_10_3842, i_10_3847, i_10_3851, i_10_3854, i_10_3855, i_10_3856, i_10_3857, i_10_3860, i_10_3907, i_10_3978, i_10_4051, i_10_4052, i_10_4113, i_10_4114, i_10_4120, i_10_4168, i_10_4276, i_10_4288, i_10_4289, i_10_4564, i_10_4565, i_10_4568, i_10_4570, o_10_274);
	kernel_10_275 k_10_275(i_10_69, i_10_176, i_10_178, i_10_283, i_10_284, i_10_328, i_10_329, i_10_406, i_10_409, i_10_410, i_10_412, i_10_458, i_10_462, i_10_463, i_10_464, i_10_466, i_10_467, i_10_511, i_10_799, i_10_800, i_10_959, i_10_962, i_10_1002, i_10_1233, i_10_1307, i_10_1312, i_10_1547, i_10_1552, i_10_1553, i_10_1555, i_10_1556, i_10_1626, i_10_1652, i_10_1691, i_10_1716, i_10_1717, i_10_1726, i_10_1821, i_10_1822, i_10_1825, i_10_1949, i_10_2005, i_10_2159, i_10_2199, i_10_2311, i_10_2312, i_10_2352, i_10_2353, i_10_2354, i_10_2355, i_10_2407, i_10_2473, i_10_2631, i_10_2632, i_10_2635, i_10_2656, i_10_2661, i_10_2663, i_10_2725, i_10_2730, i_10_2731, i_10_2827, i_10_2832, i_10_2834, i_10_2880, i_10_2881, i_10_2921, i_10_2923, i_10_2924, i_10_3075, i_10_3076, i_10_3094, i_10_3155, i_10_3385, i_10_3388, i_10_3389, i_10_3391, i_10_3392, i_10_3497, i_10_3541, i_10_3545, i_10_3551, i_10_3614, i_10_3783, i_10_3788, i_10_3835, i_10_3854, i_10_3856, i_10_3859, i_10_3860, i_10_3894, i_10_3982, i_10_3994, i_10_4050, i_10_4124, i_10_4220, i_10_4237, i_10_4270, i_10_4273, i_10_4564, o_10_275);
	kernel_10_276 k_10_276(i_10_160, i_10_259, i_10_282, i_10_283, i_10_315, i_10_320, i_10_328, i_10_367, i_10_393, i_10_425, i_10_436, i_10_445, i_10_446, i_10_447, i_10_463, i_10_464, i_10_715, i_10_750, i_10_864, i_10_1005, i_10_1104, i_10_1237, i_10_1296, i_10_1308, i_10_1309, i_10_1341, i_10_1365, i_10_1432, i_10_1575, i_10_1576, i_10_1626, i_10_1648, i_10_1651, i_10_1653, i_10_1683, i_10_1684, i_10_1687, i_10_1688, i_10_1689, i_10_1690, i_10_1710, i_10_1711, i_10_1821, i_10_1824, i_10_1826, i_10_1995, i_10_2349, i_10_2362, i_10_2364, i_10_2365, i_10_2453, i_10_2456, i_10_2460, i_10_2463, i_10_2468, i_10_2479, i_10_2511, i_10_2513, i_10_2565, i_10_2628, i_10_2631, i_10_2633, i_10_2657, i_10_2658, i_10_2660, i_10_2728, i_10_2731, i_10_2742, i_10_2754, i_10_2830, i_10_2831, i_10_2834, i_10_2869, i_10_2924, i_10_2953, i_10_2976, i_10_3036, i_10_3038, i_10_3075, i_10_3268, i_10_3280, i_10_3281, i_10_3501, i_10_3537, i_10_3582, i_10_3610, i_10_3611, i_10_3855, i_10_3856, i_10_3858, i_10_3860, i_10_3893, i_10_3919, i_10_4114, i_10_4116, i_10_4123, i_10_4156, i_10_4167, i_10_4275, i_10_4582, o_10_276);
	kernel_10_277 k_10_277(i_10_47, i_10_179, i_10_254, i_10_281, i_10_285, i_10_388, i_10_391, i_10_406, i_10_506, i_10_542, i_10_560, i_10_623, i_10_712, i_10_983, i_10_1000, i_10_1001, i_10_1003, i_10_1028, i_10_1100, i_10_1190, i_10_1207, i_10_1243, i_10_1280, i_10_1362, i_10_1363, i_10_1366, i_10_1397, i_10_1436, i_10_1541, i_10_1568, i_10_1577, i_10_1582, i_10_1613, i_10_1654, i_10_1655, i_10_1687, i_10_1688, i_10_1693, i_10_1730, i_10_1819, i_10_1820, i_10_1826, i_10_1828, i_10_1955, i_10_2020, i_10_2027, i_10_2350, i_10_2362, i_10_2365, i_10_2377, i_10_2435, i_10_2467, i_10_2470, i_10_2476, i_10_2531, i_10_2533, i_10_2534, i_10_2567, i_10_2661, i_10_2702, i_10_2705, i_10_2711, i_10_2713, i_10_2719, i_10_2755, i_10_2836, i_10_2846, i_10_2863, i_10_2867, i_10_3041, i_10_3042, i_10_3045, i_10_3074, i_10_3196, i_10_3232, i_10_3332, i_10_3350, i_10_3387, i_10_3388, i_10_3407, i_10_3439, i_10_3440, i_10_3449, i_10_3484, i_10_3503, i_10_3519, i_10_3609, i_10_3808, i_10_3837, i_10_3842, i_10_3908, i_10_3911, i_10_3982, i_10_4113, i_10_4114, i_10_4124, i_10_4145, i_10_4151, i_10_4268, i_10_4286, o_10_277);
	kernel_10_278 k_10_278(i_10_21, i_10_22, i_10_23, i_10_27, i_10_55, i_10_82, i_10_171, i_10_270, i_10_373, i_10_460, i_10_461, i_10_468, i_10_469, i_10_477, i_10_478, i_10_495, i_10_498, i_10_567, i_10_568, i_10_569, i_10_675, i_10_676, i_10_730, i_10_901, i_10_945, i_10_999, i_10_1171, i_10_1235, i_10_1280, i_10_1368, i_10_1521, i_10_1522, i_10_1566, i_10_1569, i_10_1570, i_10_1690, i_10_1691, i_10_1728, i_10_1729, i_10_1737, i_10_1768, i_10_1845, i_10_1927, i_10_1944, i_10_1945, i_10_2025, i_10_2180, i_10_2244, i_10_2322, i_10_2325, i_10_2333, i_10_2334, i_10_2358, i_10_2538, i_10_2569, i_10_2602, i_10_2610, i_10_2709, i_10_2764, i_10_2817, i_10_2839, i_10_2919, i_10_2981, i_10_3025, i_10_3096, i_10_3186, i_10_3258, i_10_3268, i_10_3288, i_10_3357, i_10_3358, i_10_3359, i_10_3474, i_10_3583, i_10_3600, i_10_3601, i_10_3615, i_10_3651, i_10_3727, i_10_3799, i_10_3802, i_10_3850, i_10_3860, i_10_3861, i_10_3870, i_10_3892, i_10_3927, i_10_3942, i_10_4068, i_10_4069, i_10_4086, i_10_4095, i_10_4116, i_10_4185, i_10_4231, i_10_4430, i_10_4432, i_10_4433, i_10_4437, i_10_4446, o_10_278);
	kernel_10_279 k_10_279(i_10_33, i_10_34, i_10_40, i_10_82, i_10_124, i_10_185, i_10_187, i_10_196, i_10_272, i_10_275, i_10_282, i_10_321, i_10_374, i_10_390, i_10_393, i_10_394, i_10_465, i_10_499, i_10_564, i_10_629, i_10_700, i_10_906, i_10_988, i_10_1048, i_10_1201, i_10_1234, i_10_1241, i_10_1249, i_10_1312, i_10_1365, i_10_1366, i_10_1543, i_10_1547, i_10_1641, i_10_1646, i_10_1651, i_10_1756, i_10_1905, i_10_1906, i_10_1930, i_10_1931, i_10_1933, i_10_1934, i_10_1941, i_10_1942, i_10_1951, i_10_1952, i_10_2094, i_10_2095, i_10_2245, i_10_2275, i_10_2276, i_10_2330, i_10_2380, i_10_2464, i_10_2515, i_10_2518, i_10_2632, i_10_2678, i_10_2726, i_10_2823, i_10_2851, i_10_2947, i_10_2982, i_10_2986, i_10_3050, i_10_3076, i_10_3093, i_10_3100, i_10_3208, i_10_3315, i_10_3316, i_10_3356, i_10_3392, i_10_3466, i_10_3471, i_10_3472, i_10_3495, i_10_3544, i_10_3585, i_10_3588, i_10_3589, i_10_3613, i_10_3624, i_10_3625, i_10_3649, i_10_3653, i_10_3751, i_10_3805, i_10_3931, i_10_3985, i_10_4189, i_10_4237, i_10_4287, i_10_4292, i_10_4524, i_10_4525, i_10_4526, i_10_4533, i_10_4534, o_10_279);
	kernel_10_280 k_10_280(i_10_27, i_10_117, i_10_207, i_10_262, i_10_282, i_10_283, i_10_284, i_10_287, i_10_325, i_10_369, i_10_390, i_10_423, i_10_426, i_10_433, i_10_434, i_10_558, i_10_730, i_10_793, i_10_797, i_10_945, i_10_958, i_10_969, i_10_996, i_10_1044, i_10_1163, i_10_1236, i_10_1341, i_10_1359, i_10_1377, i_10_1449, i_10_1450, i_10_1494, i_10_1611, i_10_1620, i_10_1630, i_10_1651, i_10_1684, i_10_1686, i_10_1689, i_10_1768, i_10_1818, i_10_1820, i_10_1822, i_10_1823, i_10_1825, i_10_1899, i_10_1944, i_10_2019, i_10_2089, i_10_2091, i_10_2178, i_10_2350, i_10_2403, i_10_2502, i_10_2505, i_10_2514, i_10_2601, i_10_2610, i_10_2611, i_10_2655, i_10_2661, i_10_2673, i_10_2700, i_10_2721, i_10_2729, i_10_2784, i_10_2817, i_10_2880, i_10_2907, i_10_2919, i_10_3036, i_10_3198, i_10_3231, i_10_3384, i_10_3385, i_10_3387, i_10_3402, i_10_3409, i_10_3468, i_10_3496, i_10_3555, i_10_3590, i_10_3618, i_10_3646, i_10_3786, i_10_3787, i_10_3837, i_10_3851, i_10_3895, i_10_3942, i_10_3978, i_10_3979, i_10_4053, i_10_4125, i_10_4176, i_10_4230, i_10_4419, i_10_4527, i_10_4567, i_10_4581, o_10_280);
	kernel_10_281 k_10_281(i_10_40, i_10_171, i_10_174, i_10_253, i_10_280, i_10_282, i_10_283, i_10_424, i_10_444, i_10_463, i_10_464, i_10_713, i_10_749, i_10_820, i_10_967, i_10_1027, i_10_1028, i_10_1040, i_10_1235, i_10_1236, i_10_1237, i_10_1243, i_10_1296, i_10_1305, i_10_1359, i_10_1444, i_10_1540, i_10_1541, i_10_1650, i_10_1683, i_10_1684, i_10_1686, i_10_1687, i_10_1691, i_10_1730, i_10_1765, i_10_1801, i_10_1821, i_10_1824, i_10_1954, i_10_2027, i_10_2199, i_10_2350, i_10_2467, i_10_2470, i_10_2557, i_10_2566, i_10_2602, i_10_2628, i_10_2631, i_10_2632, i_10_2633, i_10_2659, i_10_2728, i_10_2731, i_10_2818, i_10_2828, i_10_2920, i_10_2921, i_10_3037, i_10_3070, i_10_3198, i_10_3199, i_10_3200, i_10_3277, i_10_3278, i_10_3281, i_10_3386, i_10_3389, i_10_3406, i_10_3407, i_10_3522, i_10_3523, i_10_3538, i_10_3541, i_10_3584, i_10_3613, i_10_3615, i_10_3646, i_10_3650, i_10_3781, i_10_3782, i_10_3784, i_10_3837, i_10_3846, i_10_3853, i_10_3854, i_10_3856, i_10_3857, i_10_4115, i_10_4121, i_10_4171, i_10_4204, i_10_4267, i_10_4275, i_10_4276, i_10_4285, i_10_4286, i_10_4567, i_10_4582, o_10_281);
	kernel_10_282 k_10_282(i_10_64, i_10_144, i_10_177, i_10_189, i_10_190, i_10_275, i_10_315, i_10_369, i_10_388, i_10_391, i_10_443, i_10_447, i_10_459, i_10_460, i_10_463, i_10_465, i_10_535, i_10_536, i_10_585, i_10_588, i_10_698, i_10_700, i_10_800, i_10_967, i_10_994, i_10_1233, i_10_1290, i_10_1307, i_10_1312, i_10_1343, i_10_1417, i_10_1444, i_10_1447, i_10_1476, i_10_1551, i_10_1552, i_10_1556, i_10_1618, i_10_1648, i_10_1651, i_10_1801, i_10_1820, i_10_1826, i_10_1980, i_10_1982, i_10_2304, i_10_2305, i_10_2352, i_10_2430, i_10_2451, i_10_2514, i_10_2607, i_10_2608, i_10_2609, i_10_2629, i_10_2630, i_10_2641, i_10_2655, i_10_2660, i_10_2679, i_10_2722, i_10_2726, i_10_2734, i_10_2829, i_10_2830, i_10_2832, i_10_2923, i_10_3034, i_10_3036, i_10_3199, i_10_3271, i_10_3317, i_10_3402, i_10_3403, i_10_3405, i_10_3408, i_10_3469, i_10_3492, i_10_3493, i_10_3495, i_10_3523, i_10_3540, i_10_3639, i_10_3649, i_10_3682, i_10_3706, i_10_3846, i_10_3855, i_10_3857, i_10_3978, i_10_3979, i_10_3986, i_10_4030, i_10_4171, i_10_4266, i_10_4352, i_10_4354, i_10_4567, i_10_4582, i_10_4595, o_10_282);
	kernel_10_283 k_10_283(i_10_222, i_10_324, i_10_433, i_10_442, i_10_444, i_10_463, i_10_513, i_10_516, i_10_793, i_10_794, i_10_796, i_10_900, i_10_954, i_10_959, i_10_966, i_10_967, i_10_968, i_10_990, i_10_1027, i_10_1028, i_10_1031, i_10_1036, i_10_1235, i_10_1263, i_10_1359, i_10_1444, i_10_1651, i_10_1654, i_10_1683, i_10_1684, i_10_1689, i_10_1812, i_10_1818, i_10_1819, i_10_1823, i_10_1825, i_10_1872, i_10_2322, i_10_2325, i_10_2351, i_10_2356, i_10_2461, i_10_2502, i_10_2604, i_10_2635, i_10_2673, i_10_2674, i_10_2700, i_10_2701, i_10_2723, i_10_2781, i_10_2782, i_10_2817, i_10_2828, i_10_2919, i_10_2921, i_10_2979, i_10_2980, i_10_3043, i_10_3071, i_10_3073, i_10_3200, i_10_3201, i_10_3387, i_10_3389, i_10_3391, i_10_3405, i_10_3406, i_10_3519, i_10_3522, i_10_3582, i_10_3585, i_10_3684, i_10_3780, i_10_3781, i_10_3783, i_10_3784, i_10_3788, i_10_3838, i_10_3839, i_10_3841, i_10_3854, i_10_3855, i_10_3889, i_10_3979, i_10_3980, i_10_3991, i_10_4027, i_10_4030, i_10_4116, i_10_4117, i_10_4230, i_10_4266, i_10_4267, i_10_4285, i_10_4292, i_10_4458, i_10_4461, i_10_4564, i_10_4566, o_10_283);
	kernel_10_284 k_10_284(i_10_65, i_10_178, i_10_181, i_10_220, i_10_280, i_10_425, i_10_434, i_10_448, i_10_460, i_10_796, i_10_1036, i_10_1200, i_10_1233, i_10_1234, i_10_1240, i_10_1242, i_10_1342, i_10_1359, i_10_1550, i_10_1576, i_10_1651, i_10_1819, i_10_1913, i_10_1945, i_10_1946, i_10_1949, i_10_1991, i_10_2178, i_10_2179, i_10_2305, i_10_2306, i_10_2324, i_10_2333, i_10_2354, i_10_2358, i_10_2359, i_10_2362, i_10_2363, i_10_2378, i_10_2381, i_10_2404, i_10_2451, i_10_2453, i_10_2463, i_10_2467, i_10_2475, i_10_2476, i_10_2503, i_10_2628, i_10_2634, i_10_2635, i_10_2659, i_10_2660, i_10_2674, i_10_2704, i_10_2709, i_10_2710, i_10_2711, i_10_2721, i_10_2727, i_10_2730, i_10_2731, i_10_2732, i_10_2828, i_10_2886, i_10_2916, i_10_2924, i_10_3034, i_10_3035, i_10_3040, i_10_3087, i_10_3088, i_10_3203, i_10_3268, i_10_3269, i_10_3384, i_10_3403, i_10_3404, i_10_3405, i_10_3406, i_10_3407, i_10_3648, i_10_3682, i_10_3838, i_10_3848, i_10_3858, i_10_3893, i_10_3908, i_10_3978, i_10_3991, i_10_4051, i_10_4052, i_10_4116, i_10_4121, i_10_4129, i_10_4214, i_10_4231, i_10_4232, i_10_4270, i_10_4528, o_10_284);
	kernel_10_285 k_10_285(i_10_121, i_10_148, i_10_171, i_10_174, i_10_175, i_10_219, i_10_220, i_10_244, i_10_271, i_10_279, i_10_280, i_10_281, i_10_328, i_10_390, i_10_435, i_10_439, i_10_447, i_10_507, i_10_747, i_10_748, i_10_750, i_10_793, i_10_891, i_10_1000, i_10_1026, i_10_1027, i_10_1028, i_10_1029, i_10_1233, i_10_1242, i_10_1306, i_10_1307, i_10_1308, i_10_1309, i_10_1311, i_10_1312, i_10_1539, i_10_1540, i_10_1575, i_10_1576, i_10_1647, i_10_1648, i_10_1651, i_10_1655, i_10_1711, i_10_1818, i_10_1822, i_10_2196, i_10_2199, i_10_2202, i_10_2349, i_10_2350, i_10_2364, i_10_2406, i_10_2463, i_10_2466, i_10_2467, i_10_2468, i_10_2470, i_10_2512, i_10_2530, i_10_2604, i_10_2628, i_10_2629, i_10_2674, i_10_2710, i_10_2711, i_10_2720, i_10_2722, i_10_2727, i_10_2732, i_10_2829, i_10_2830, i_10_2981, i_10_3038, i_10_3154, i_10_3159, i_10_3198, i_10_3270, i_10_3271, i_10_3322, i_10_3408, i_10_3409, i_10_3465, i_10_3466, i_10_3582, i_10_3586, i_10_3785, i_10_3807, i_10_3808, i_10_3841, i_10_3842, i_10_3853, i_10_3855, i_10_3857, i_10_4113, i_10_4114, i_10_4119, i_10_4269, i_10_4288, o_10_285);
	kernel_10_286 k_10_286(i_10_208, i_10_209, i_10_218, i_10_270, i_10_271, i_10_272, i_10_281, i_10_283, i_10_407, i_10_424, i_10_425, i_10_433, i_10_437, i_10_445, i_10_465, i_10_508, i_10_902, i_10_986, i_10_1036, i_10_1117, i_10_1118, i_10_1217, i_10_1235, i_10_1243, i_10_1244, i_10_1361, i_10_1444, i_10_1445, i_10_1822, i_10_1823, i_10_1882, i_10_1883, i_10_1990, i_10_2089, i_10_2323, i_10_2327, i_10_2333, i_10_2351, i_10_2368, i_10_2369, i_10_2432, i_10_2441, i_10_2462, i_10_2606, i_10_2630, i_10_2634, i_10_2639, i_10_2674, i_10_2675, i_10_2701, i_10_2702, i_10_2705, i_10_2728, i_10_2819, i_10_2831, i_10_2863, i_10_2864, i_10_2917, i_10_2920, i_10_2921, i_10_3034, i_10_3224, i_10_3281, i_10_3298, i_10_3349, i_10_3406, i_10_3466, i_10_3647, i_10_3682, i_10_3782, i_10_3785, i_10_3847, i_10_3848, i_10_3849, i_10_3857, i_10_3889, i_10_3890, i_10_3893, i_10_3980, i_10_4028, i_10_4118, i_10_4142, i_10_4185, i_10_4186, i_10_4187, i_10_4276, i_10_4277, i_10_4285, i_10_4286, i_10_4288, i_10_4289, i_10_4290, i_10_4291, i_10_4510, i_10_4511, i_10_4563, i_10_4564, i_10_4571, i_10_4583, i_10_4601, o_10_286);
	kernel_10_287 k_10_287(i_10_34, i_10_89, i_10_174, i_10_175, i_10_176, i_10_177, i_10_178, i_10_249, i_10_267, i_10_277, i_10_283, i_10_284, i_10_412, i_10_440, i_10_509, i_10_796, i_10_898, i_10_963, i_10_1033, i_10_1034, i_10_1165, i_10_1237, i_10_1311, i_10_1362, i_10_1440, i_10_1491, i_10_1549, i_10_1550, i_10_1651, i_10_1654, i_10_1655, i_10_1821, i_10_1822, i_10_1823, i_10_2026, i_10_2334, i_10_2350, i_10_2351, i_10_2353, i_10_2354, i_10_2407, i_10_2408, i_10_2449, i_10_2452, i_10_2453, i_10_2465, i_10_2608, i_10_2609, i_10_2631, i_10_2635, i_10_2636, i_10_2644, i_10_2678, i_10_2725, i_10_2733, i_10_2735, i_10_2829, i_10_2919, i_10_3076, i_10_3154, i_10_3155, i_10_3156, i_10_3162, i_10_3165, i_10_3166, i_10_3167, i_10_3201, i_10_3237, i_10_3279, i_10_3280, i_10_3282, i_10_3385, i_10_3386, i_10_3388, i_10_3389, i_10_3390, i_10_3525, i_10_3586, i_10_3587, i_10_3613, i_10_3614, i_10_3853, i_10_3855, i_10_3891, i_10_3912, i_10_3991, i_10_4113, i_10_4117, i_10_4118, i_10_4119, i_10_4121, i_10_4125, i_10_4126, i_10_4128, i_10_4129, i_10_4130, i_10_4174, i_10_4219, i_10_4272, i_10_4292, o_10_287);
	kernel_10_288 k_10_288(i_10_48, i_10_63, i_10_81, i_10_117, i_10_174, i_10_178, i_10_219, i_10_220, i_10_222, i_10_223, i_10_224, i_10_261, i_10_285, i_10_286, i_10_367, i_10_406, i_10_427, i_10_439, i_10_531, i_10_534, i_10_736, i_10_901, i_10_957, i_10_999, i_10_1041, i_10_1156, i_10_1233, i_10_1236, i_10_1296, i_10_1310, i_10_1341, i_10_1359, i_10_1440, i_10_1441, i_10_1476, i_10_1540, i_10_1614, i_10_1653, i_10_1655, i_10_1711, i_10_1719, i_10_1764, i_10_1765, i_10_1821, i_10_1890, i_10_1909, i_10_1912, i_10_1916, i_10_1945, i_10_2019, i_10_2109, i_10_2160, i_10_2178, i_10_2236, i_10_2254, i_10_2350, i_10_2361, i_10_2377, i_10_2466, i_10_2469, i_10_2515, i_10_2541, i_10_2655, i_10_2676, i_10_2704, i_10_2709, i_10_2742, i_10_2844, i_10_2923, i_10_3033, i_10_3040, i_10_3095, i_10_3114, i_10_3231, i_10_3270, i_10_3277, i_10_3289, i_10_3331, i_10_3434, i_10_3465, i_10_3492, i_10_3523, i_10_3526, i_10_3538, i_10_3561, i_10_3582, i_10_3837, i_10_3852, i_10_3853, i_10_3859, i_10_3901, i_10_4114, i_10_4161, i_10_4218, i_10_4219, i_10_4222, i_10_4234, i_10_4311, i_10_4554, i_10_4580, o_10_288);
	kernel_10_289 k_10_289(i_10_124, i_10_125, i_10_174, i_10_177, i_10_183, i_10_184, i_10_280, i_10_285, i_10_286, i_10_287, i_10_317, i_10_318, i_10_319, i_10_446, i_10_449, i_10_460, i_10_462, i_10_463, i_10_464, i_10_510, i_10_511, i_10_514, i_10_749, i_10_955, i_10_993, i_10_1006, i_10_1034, i_10_1037, i_10_1244, i_10_1247, i_10_1308, i_10_1310, i_10_1363, i_10_1380, i_10_1552, i_10_1653, i_10_1685, i_10_1819, i_10_1820, i_10_1822, i_10_1823, i_10_1825, i_10_1826, i_10_1950, i_10_1995, i_10_2095, i_10_2351, i_10_2354, i_10_2356, i_10_2361, i_10_2362, i_10_2455, i_10_2469, i_10_2632, i_10_2702, i_10_2713, i_10_2715, i_10_2722, i_10_2724, i_10_2725, i_10_2731, i_10_2734, i_10_2829, i_10_2830, i_10_2834, i_10_2920, i_10_3040, i_10_3041, i_10_3151, i_10_3195, i_10_3196, i_10_3197, i_10_3198, i_10_3199, i_10_3270, i_10_3271, i_10_3328, i_10_3387, i_10_3388, i_10_3389, i_10_3391, i_10_3392, i_10_3610, i_10_3613, i_10_3647, i_10_3649, i_10_3653, i_10_3780, i_10_3781, i_10_3782, i_10_3837, i_10_3838, i_10_3839, i_10_3842, i_10_3856, i_10_3967, i_10_3985, i_10_4114, i_10_4291, i_10_4427, o_10_289);
	kernel_10_290 k_10_290(i_10_36, i_10_64, i_10_68, i_10_119, i_10_191, i_10_254, i_10_262, i_10_316, i_10_319, i_10_411, i_10_433, i_10_443, i_10_448, i_10_497, i_10_514, i_10_515, i_10_695, i_10_712, i_10_829, i_10_830, i_10_1036, i_10_1037, i_10_1082, i_10_1099, i_10_1108, i_10_1109, i_10_1235, i_10_1265, i_10_1273, i_10_1301, i_10_1360, i_10_1361, i_10_1433, i_10_1451, i_10_1540, i_10_1541, i_10_1544, i_10_1621, i_10_1622, i_10_1739, i_10_1801, i_10_1802, i_10_1804, i_10_1874, i_10_1981, i_10_1996, i_10_1997, i_10_2018, i_10_2111, i_10_2153, i_10_2198, i_10_2201, i_10_2305, i_10_2306, i_10_2350, i_10_2351, i_10_2365, i_10_2376, i_10_2377, i_10_2467, i_10_2531, i_10_2558, i_10_2567, i_10_2585, i_10_2594, i_10_2609, i_10_2612, i_10_2615, i_10_2629, i_10_2653, i_10_2654, i_10_2675, i_10_2714, i_10_2830, i_10_2935, i_10_3092, i_10_3199, i_10_3280, i_10_3404, i_10_3410, i_10_3467, i_10_3494, i_10_3538, i_10_3584, i_10_3686, i_10_3692, i_10_3699, i_10_3794, i_10_3836, i_10_3839, i_10_3851, i_10_4115, i_10_4151, i_10_4154, i_10_4275, i_10_4278, i_10_4291, i_10_4547, i_10_4569, i_10_4571, o_10_290);
	kernel_10_291 k_10_291(i_10_41, i_10_43, i_10_46, i_10_63, i_10_65, i_10_155, i_10_246, i_10_248, i_10_249, i_10_289, i_10_409, i_10_595, i_10_608, i_10_712, i_10_713, i_10_756, i_10_875, i_10_901, i_10_947, i_10_993, i_10_1010, i_10_1120, i_10_1157, i_10_1433, i_10_1488, i_10_1540, i_10_1614, i_10_1649, i_10_1703, i_10_1710, i_10_1802, i_10_1873, i_10_1915, i_10_1916, i_10_1947, i_10_2021, i_10_2030, i_10_2054, i_10_2109, i_10_2162, i_10_2180, i_10_2218, i_10_2304, i_10_2333, i_10_2336, i_10_2351, i_10_2359, i_10_2366, i_10_2431, i_10_2450, i_10_2451, i_10_2529, i_10_2602, i_10_2702, i_10_2705, i_10_2709, i_10_2713, i_10_2720, i_10_2863, i_10_2864, i_10_2923, i_10_3024, i_10_3071, i_10_3073, i_10_3074, i_10_3223, i_10_3227, i_10_3269, i_10_3278, i_10_3280, i_10_3287, i_10_3304, i_10_3330, i_10_3331, i_10_3385, i_10_3387, i_10_3403, i_10_3431, i_10_3523, i_10_3619, i_10_3647, i_10_3651, i_10_3730, i_10_3771, i_10_3774, i_10_3807, i_10_3834, i_10_3838, i_10_3839, i_10_3840, i_10_3849, i_10_3893, i_10_3902, i_10_3989, i_10_3993, i_10_4118, i_10_4188, i_10_4217, i_10_4302, i_10_4430, o_10_291);
	kernel_10_292 k_10_292(i_10_68, i_10_175, i_10_247, i_10_273, i_10_319, i_10_328, i_10_355, i_10_363, i_10_390, i_10_425, i_10_435, i_10_442, i_10_443, i_10_465, i_10_518, i_10_608, i_10_631, i_10_734, i_10_736, i_10_793, i_10_794, i_10_796, i_10_799, i_10_908, i_10_956, i_10_977, i_10_993, i_10_1041, i_10_1163, i_10_1184, i_10_1194, i_10_1195, i_10_1220, i_10_1276, i_10_1360, i_10_1583, i_10_1683, i_10_1790, i_10_1894, i_10_1900, i_10_1911, i_10_1912, i_10_2003, i_10_2027, i_10_2030, i_10_2083, i_10_2158, i_10_2308, i_10_2309, i_10_2336, i_10_2359, i_10_2379, i_10_2381, i_10_2389, i_10_2480, i_10_2498, i_10_2542, i_10_2543, i_10_2603, i_10_2606, i_10_2629, i_10_2662, i_10_2727, i_10_2859, i_10_2923, i_10_2952, i_10_2983, i_10_2984, i_10_3044, i_10_3047, i_10_3056, i_10_3195, i_10_3196, i_10_3231, i_10_3273, i_10_3275, i_10_3300, i_10_3302, i_10_3325, i_10_3362, i_10_3363, i_10_3541, i_10_3647, i_10_3653, i_10_3684, i_10_3857, i_10_3875, i_10_3893, i_10_3945, i_10_3995, i_10_4113, i_10_4122, i_10_4220, i_10_4237, i_10_4275, i_10_4278, i_10_4295, i_10_4378, i_10_4381, i_10_4478, o_10_292);
	kernel_10_293 k_10_293(i_10_28, i_10_29, i_10_31, i_10_32, i_10_45, i_10_46, i_10_124, i_10_224, i_10_408, i_10_437, i_10_443, i_10_444, i_10_461, i_10_465, i_10_466, i_10_516, i_10_517, i_10_732, i_10_733, i_10_753, i_10_754, i_10_755, i_10_928, i_10_961, i_10_1032, i_10_1305, i_10_1306, i_10_1310, i_10_1312, i_10_1313, i_10_1546, i_10_1559, i_10_1616, i_10_1648, i_10_1800, i_10_1818, i_10_1948, i_10_1949, i_10_1951, i_10_1952, i_10_2006, i_10_2366, i_10_2407, i_10_2473, i_10_2603, i_10_2632, i_10_2633, i_10_2635, i_10_2655, i_10_2656, i_10_2657, i_10_2660, i_10_2718, i_10_2719, i_10_2722, i_10_2723, i_10_2724, i_10_2726, i_10_2735, i_10_2826, i_10_2827, i_10_2828, i_10_2887, i_10_2924, i_10_2986, i_10_3036, i_10_3039, i_10_3040, i_10_3041, i_10_3045, i_10_3046, i_10_3196, i_10_3276, i_10_3278, i_10_3279, i_10_3349, i_10_3390, i_10_3391, i_10_3392, i_10_3494, i_10_3522, i_10_3587, i_10_3610, i_10_3611, i_10_3646, i_10_3649, i_10_3651, i_10_3653, i_10_3688, i_10_3689, i_10_3727, i_10_3728, i_10_3780, i_10_3781, i_10_3852, i_10_3853, i_10_3856, i_10_3859, i_10_4025, i_10_4127, o_10_293);
	kernel_10_294 k_10_294(i_10_118, i_10_175, i_10_186, i_10_243, i_10_282, i_10_283, i_10_284, i_10_285, i_10_318, i_10_319, i_10_408, i_10_409, i_10_410, i_10_412, i_10_430, i_10_431, i_10_460, i_10_461, i_10_508, i_10_511, i_10_737, i_10_1002, i_10_1135, i_10_1168, i_10_1234, i_10_1235, i_10_1237, i_10_1238, i_10_1307, i_10_1309, i_10_1310, i_10_1552, i_10_1555, i_10_1575, i_10_1582, i_10_1615, i_10_1647, i_10_1652, i_10_1653, i_10_1681, i_10_1687, i_10_1821, i_10_1822, i_10_1823, i_10_1825, i_10_1826, i_10_1914, i_10_1915, i_10_1916, i_10_2022, i_10_2311, i_10_2355, i_10_2362, i_10_2383, i_10_2453, i_10_2456, i_10_2473, i_10_2631, i_10_2634, i_10_2655, i_10_2656, i_10_2658, i_10_2659, i_10_2679, i_10_2704, i_10_2706, i_10_2707, i_10_2715, i_10_2716, i_10_2719, i_10_2735, i_10_2788, i_10_2831, i_10_2888, i_10_2983, i_10_3034, i_10_3040, i_10_3044, i_10_3046, i_10_3196, i_10_3197, i_10_3279, i_10_3319, i_10_3387, i_10_3392, i_10_3405, i_10_3409, i_10_3613, i_10_3783, i_10_3835, i_10_3840, i_10_3842, i_10_3847, i_10_3854, i_10_3981, i_10_4050, i_10_4119, i_10_4130, i_10_4191, i_10_4289, o_10_294);
	kernel_10_295 k_10_295(i_10_28, i_10_171, i_10_174, i_10_178, i_10_183, i_10_185, i_10_317, i_10_390, i_10_410, i_10_427, i_10_442, i_10_443, i_10_459, i_10_566, i_10_748, i_10_792, i_10_798, i_10_1027, i_10_1033, i_10_1034, i_10_1042, i_10_1043, i_10_1236, i_10_1245, i_10_1246, i_10_1247, i_10_1539, i_10_1542, i_10_1543, i_10_1575, i_10_1576, i_10_1650, i_10_1655, i_10_1683, i_10_1684, i_10_1686, i_10_1688, i_10_1769, i_10_1911, i_10_1912, i_10_1913, i_10_1915, i_10_1948, i_10_1949, i_10_1997, i_10_2201, i_10_2353, i_10_2380, i_10_2448, i_10_2470, i_10_2632, i_10_2636, i_10_2659, i_10_2661, i_10_2662, i_10_2701, i_10_2706, i_10_2709, i_10_2721, i_10_2723, i_10_2728, i_10_2729, i_10_2827, i_10_2828, i_10_2831, i_10_3035, i_10_3040, i_10_3041, i_10_3043, i_10_3152, i_10_3198, i_10_3199, i_10_3277, i_10_3329, i_10_3388, i_10_3497, i_10_3525, i_10_3583, i_10_3586, i_10_3614, i_10_3649, i_10_3653, i_10_3780, i_10_3783, i_10_3837, i_10_3839, i_10_3855, i_10_3858, i_10_3894, i_10_3895, i_10_3896, i_10_3985, i_10_4116, i_10_4128, i_10_4129, i_10_4169, i_10_4276, i_10_4290, i_10_4291, i_10_4535, o_10_295);
	kernel_10_296 k_10_296(i_10_9, i_10_223, i_10_270, i_10_272, i_10_279, i_10_285, i_10_447, i_10_462, i_10_464, i_10_505, i_10_506, i_10_507, i_10_508, i_10_513, i_10_516, i_10_711, i_10_712, i_10_749, i_10_957, i_10_967, i_10_999, i_10_1080, i_10_1083, i_10_1098, i_10_1215, i_10_1239, i_10_1263, i_10_1306, i_10_1539, i_10_1549, i_10_1578, i_10_1653, i_10_1686, i_10_1782, i_10_1821, i_10_1822, i_10_1990, i_10_2016, i_10_2088, i_10_2179, i_10_2196, i_10_2197, i_10_2199, i_10_2352, i_10_2376, i_10_2448, i_10_2502, i_10_2574, i_10_2604, i_10_2610, i_10_2629, i_10_2630, i_10_2631, i_10_2655, i_10_2659, i_10_2662, i_10_2673, i_10_2700, i_10_2701, i_10_2703, i_10_2713, i_10_2882, i_10_2917, i_10_2979, i_10_3046, i_10_3054, i_10_3055, i_10_3088, i_10_3158, i_10_3328, i_10_3329, i_10_3385, i_10_3387, i_10_3538, i_10_3616, i_10_3681, i_10_3781, i_10_3785, i_10_3844, i_10_3852, i_10_3853, i_10_3854, i_10_3855, i_10_3858, i_10_3859, i_10_3860, i_10_3978, i_10_3979, i_10_4122, i_10_4123, i_10_4126, i_10_4167, i_10_4168, i_10_4170, i_10_4266, i_10_4267, i_10_4269, i_10_4275, i_10_4278, i_10_4567, o_10_296);
	kernel_10_297 k_10_297(i_10_175, i_10_283, i_10_287, i_10_390, i_10_426, i_10_429, i_10_430, i_10_467, i_10_506, i_10_516, i_10_518, i_10_519, i_10_714, i_10_735, i_10_799, i_10_958, i_10_967, i_10_1000, i_10_1002, i_10_1263, i_10_1264, i_10_1309, i_10_1492, i_10_1552, i_10_1554, i_10_1578, i_10_1635, i_10_1651, i_10_1690, i_10_1695, i_10_1820, i_10_1823, i_10_1824, i_10_1875, i_10_1913, i_10_1938, i_10_1995, i_10_2184, i_10_2253, i_10_2310, i_10_2311, i_10_2329, i_10_2352, i_10_2452, i_10_2453, i_10_2467, i_10_2481, i_10_2508, i_10_2541, i_10_2628, i_10_2629, i_10_2630, i_10_2676, i_10_2679, i_10_2680, i_10_2708, i_10_2710, i_10_2715, i_10_2716, i_10_2824, i_10_2833, i_10_2919, i_10_3038, i_10_3041, i_10_3237, i_10_3315, i_10_3318, i_10_3321, i_10_3322, i_10_3325, i_10_3326, i_10_3388, i_10_3471, i_10_3495, i_10_3496, i_10_3504, i_10_3525, i_10_3541, i_10_3586, i_10_3588, i_10_3611, i_10_3648, i_10_3652, i_10_3782, i_10_3783, i_10_3784, i_10_3786, i_10_3836, i_10_3840, i_10_3848, i_10_3853, i_10_3859, i_10_3948, i_10_3949, i_10_3985, i_10_4057, i_10_4270, i_10_4272, i_10_4287, i_10_4291, o_10_297);
	kernel_10_298 k_10_298(i_10_118, i_10_217, i_10_221, i_10_279, i_10_280, i_10_281, i_10_284, i_10_329, i_10_389, i_10_410, i_10_463, i_10_711, i_10_712, i_10_748, i_10_749, i_10_794, i_10_796, i_10_990, i_10_999, i_10_1000, i_10_1086, i_10_1234, i_10_1237, i_10_1246, i_10_1308, i_10_1309, i_10_1310, i_10_1359, i_10_1541, i_10_1577, i_10_1613, i_10_1647, i_10_1648, i_10_1649, i_10_1651, i_10_1654, i_10_1655, i_10_1684, i_10_1687, i_10_1820, i_10_1911, i_10_1912, i_10_1913, i_10_1916, i_10_1949, i_10_2352, i_10_2353, i_10_2354, i_10_2358, i_10_2359, i_10_2361, i_10_2449, i_10_2455, i_10_2630, i_10_2633, i_10_2635, i_10_2659, i_10_2660, i_10_2718, i_10_2721, i_10_2722, i_10_2723, i_10_2727, i_10_2729, i_10_2817, i_10_2818, i_10_2919, i_10_2920, i_10_2921, i_10_2980, i_10_3034, i_10_3035, i_10_3038, i_10_3042, i_10_3043, i_10_3157, i_10_3277, i_10_3278, i_10_3279, i_10_3388, i_10_3466, i_10_3523, i_10_3556, i_10_3613, i_10_3645, i_10_3834, i_10_3840, i_10_3846, i_10_3857, i_10_3906, i_10_3907, i_10_3908, i_10_3979, i_10_4051, i_10_4113, i_10_4114, i_10_4118, i_10_4271, i_10_4288, i_10_4289, o_10_298);
	kernel_10_299 k_10_299(i_10_175, i_10_221, i_10_280, i_10_285, i_10_286, i_10_390, i_10_465, i_10_466, i_10_753, i_10_796, i_10_957, i_10_967, i_10_1032, i_10_1035, i_10_1236, i_10_1237, i_10_1239, i_10_1240, i_10_1242, i_10_1243, i_10_1248, i_10_1249, i_10_1263, i_10_1341, i_10_1359, i_10_1444, i_10_1545, i_10_1555, i_10_1576, i_10_1647, i_10_1650, i_10_1651, i_10_1683, i_10_1812, i_10_1819, i_10_1913, i_10_1915, i_10_1945, i_10_2185, i_10_2197, i_10_2199, i_10_2352, i_10_2353, i_10_2361, i_10_2449, i_10_2456, i_10_2467, i_10_2471, i_10_2601, i_10_2602, i_10_2604, i_10_2607, i_10_2628, i_10_2629, i_10_2634, i_10_2636, i_10_2659, i_10_2662, i_10_2700, i_10_2709, i_10_2731, i_10_2827, i_10_2830, i_10_2833, i_10_2981, i_10_3033, i_10_3034, i_10_3036, i_10_3037, i_10_3329, i_10_3389, i_10_3466, i_10_3549, i_10_3583, i_10_3586, i_10_3624, i_10_3645, i_10_3646, i_10_3647, i_10_3648, i_10_3649, i_10_3717, i_10_3718, i_10_3840, i_10_3843, i_10_3847, i_10_3848, i_10_3850, i_10_3852, i_10_3860, i_10_3870, i_10_3888, i_10_3982, i_10_4116, i_10_4117, i_10_4217, i_10_4275, i_10_4276, i_10_4564, i_10_4566, o_10_299);
	kernel_10_300 k_10_300(i_10_171, i_10_172, i_10_175, i_10_222, i_10_244, i_10_279, i_10_283, i_10_328, i_10_409, i_10_436, i_10_441, i_10_442, i_10_443, i_10_462, i_10_696, i_10_748, i_10_990, i_10_991, i_10_1026, i_10_1029, i_10_1233, i_10_1234, i_10_1238, i_10_1262, i_10_1265, i_10_1308, i_10_1309, i_10_1310, i_10_1445, i_10_1539, i_10_1540, i_10_1541, i_10_1575, i_10_1576, i_10_1651, i_10_1819, i_10_1822, i_10_1911, i_10_1912, i_10_1944, i_10_2179, i_10_2180, i_10_2197, i_10_2198, i_10_2201, i_10_2351, i_10_2450, i_10_2453, i_10_2468, i_10_2469, i_10_2470, i_10_2471, i_10_2629, i_10_2630, i_10_2633, i_10_2636, i_10_2661, i_10_2702, i_10_2817, i_10_2820, i_10_2827, i_10_2830, i_10_2881, i_10_2882, i_10_2884, i_10_2885, i_10_2888, i_10_3071, i_10_3078, i_10_3196, i_10_3198, i_10_3199, i_10_3200, i_10_3202, i_10_3203, i_10_3391, i_10_3403, i_10_3583, i_10_3586, i_10_3611, i_10_3613, i_10_3614, i_10_3645, i_10_3788, i_10_3834, i_10_3839, i_10_3846, i_10_3851, i_10_3853, i_10_3854, i_10_3888, i_10_3994, i_10_4113, i_10_4114, i_10_4116, i_10_4129, i_10_4278, i_10_4291, i_10_4292, i_10_4457, o_10_300);
	kernel_10_301 k_10_301(i_10_44, i_10_152, i_10_171, i_10_179, i_10_187, i_10_188, i_10_251, i_10_327, i_10_329, i_10_332, i_10_394, i_10_463, i_10_465, i_10_518, i_10_520, i_10_521, i_10_565, i_10_566, i_10_638, i_10_796, i_10_799, i_10_800, i_10_899, i_10_908, i_10_959, i_10_995, i_10_998, i_10_1166, i_10_1204, i_10_1235, i_10_1241, i_10_1264, i_10_1276, i_10_1313, i_10_1653, i_10_1817, i_10_1826, i_10_1889, i_10_1913, i_10_1997, i_10_2006, i_10_2024, i_10_2032, i_10_2033, i_10_2041, i_10_2353, i_10_2365, i_10_2450, i_10_2452, i_10_2464, i_10_2468, i_10_2510, i_10_2515, i_10_2568, i_10_2609, i_10_2681, i_10_2717, i_10_2734, i_10_2830, i_10_2882, i_10_2885, i_10_2888, i_10_2986, i_10_3033, i_10_3059, i_10_3200, i_10_3239, i_10_3270, i_10_3280, i_10_3283, i_10_3302, i_10_3409, i_10_3473, i_10_3497, i_10_3509, i_10_3526, i_10_3552, i_10_3613, i_10_3689, i_10_3783, i_10_3851, i_10_3852, i_10_3859, i_10_3878, i_10_3913, i_10_3914, i_10_3923, i_10_3983, i_10_3995, i_10_4023, i_10_4168, i_10_4237, i_10_4271, i_10_4272, i_10_4274, i_10_4287, i_10_4463, i_10_4568, i_10_4569, i_10_4571, o_10_301);
	kernel_10_302 k_10_302(i_10_118, i_10_171, i_10_172, i_10_244, i_10_249, i_10_282, i_10_285, i_10_410, i_10_431, i_10_462, i_10_467, i_10_800, i_10_957, i_10_958, i_10_959, i_10_1236, i_10_1237, i_10_1238, i_10_1240, i_10_1241, i_10_1246, i_10_1308, i_10_1309, i_10_1581, i_10_1582, i_10_1648, i_10_1649, i_10_1687, i_10_1819, i_10_1820, i_10_1821, i_10_1911, i_10_1916, i_10_1944, i_10_1945, i_10_1946, i_10_2027, i_10_2178, i_10_2179, i_10_2181, i_10_2184, i_10_2185, i_10_2186, i_10_2333, i_10_2364, i_10_2404, i_10_2407, i_10_2448, i_10_2503, i_10_2629, i_10_2630, i_10_2632, i_10_2658, i_10_2673, i_10_2700, i_10_2710, i_10_2712, i_10_2713, i_10_2722, i_10_2724, i_10_2731, i_10_2733, i_10_2882, i_10_2920, i_10_2923, i_10_2986, i_10_3034, i_10_3036, i_10_3037, i_10_3150, i_10_3156, i_10_3160, i_10_3195, i_10_3231, i_10_3276, i_10_3277, i_10_3278, i_10_3282, i_10_3409, i_10_3586, i_10_3611, i_10_3612, i_10_3613, i_10_3646, i_10_3648, i_10_3649, i_10_3784, i_10_3786, i_10_3787, i_10_3834, i_10_3835, i_10_3838, i_10_3849, i_10_4052, i_10_4267, i_10_4563, i_10_4566, i_10_4567, i_10_4568, i_10_4593, o_10_302);
	kernel_10_303 k_10_303(i_10_175, i_10_217, i_10_221, i_10_262, i_10_282, i_10_283, i_10_315, i_10_320, i_10_426, i_10_432, i_10_466, i_10_510, i_10_626, i_10_631, i_10_830, i_10_954, i_10_990, i_10_991, i_10_1026, i_10_1027, i_10_1030, i_10_1117, i_10_1236, i_10_1264, i_10_1300, i_10_1307, i_10_1341, i_10_1431, i_10_1432, i_10_1539, i_10_1578, i_10_1579, i_10_1620, i_10_1683, i_10_1684, i_10_1818, i_10_2197, i_10_2359, i_10_2361, i_10_2362, i_10_2376, i_10_2377, i_10_2408, i_10_2565, i_10_2566, i_10_2638, i_10_2659, i_10_2704, i_10_2729, i_10_2740, i_10_2743, i_10_2844, i_10_2845, i_10_2885, i_10_2918, i_10_2919, i_10_2921, i_10_3042, i_10_3196, i_10_3223, i_10_3268, i_10_3384, i_10_3386, i_10_3387, i_10_3402, i_10_3403, i_10_3431, i_10_3452, i_10_3469, i_10_3485, i_10_3538, i_10_3649, i_10_3650, i_10_3652, i_10_3682, i_10_3781, i_10_3782, i_10_3783, i_10_3784, i_10_3785, i_10_3838, i_10_3844, i_10_3852, i_10_3853, i_10_3854, i_10_3961, i_10_3980, i_10_4023, i_10_4052, i_10_4143, i_10_4168, i_10_4173, i_10_4175, i_10_4213, i_10_4214, i_10_4270, i_10_4420, i_10_4511, i_10_4581, i_10_4600, o_10_303);
	kernel_10_304 k_10_304(i_10_29, i_10_154, i_10_181, i_10_282, i_10_315, i_10_316, i_10_319, i_10_390, i_10_436, i_10_464, i_10_465, i_10_467, i_10_505, i_10_820, i_10_829, i_10_999, i_10_1053, i_10_1081, i_10_1083, i_10_1084, i_10_1154, i_10_1239, i_10_1240, i_10_1241, i_10_1265, i_10_1360, i_10_1539, i_10_1540, i_10_1542, i_10_1575, i_10_1579, i_10_1620, i_10_1621, i_10_1622, i_10_1650, i_10_1686, i_10_1687, i_10_1688, i_10_1909, i_10_1999, i_10_2008, i_10_2025, i_10_2183, i_10_2196, i_10_2197, i_10_2198, i_10_2199, i_10_2236, i_10_2350, i_10_2352, i_10_2353, i_10_2364, i_10_2406, i_10_2407, i_10_2572, i_10_2636, i_10_2659, i_10_2674, i_10_2675, i_10_2700, i_10_2701, i_10_2831, i_10_2882, i_10_2884, i_10_2922, i_10_2923, i_10_3276, i_10_3277, i_10_3278, i_10_3279, i_10_3280, i_10_3281, i_10_3316, i_10_3429, i_10_3448, i_10_3468, i_10_3469, i_10_3538, i_10_3541, i_10_3542, i_10_3555, i_10_3558, i_10_3559, i_10_3586, i_10_3836, i_10_3979, i_10_3980, i_10_4050, i_10_4113, i_10_4119, i_10_4125, i_10_4126, i_10_4127, i_10_4167, i_10_4170, i_10_4172, i_10_4276, i_10_4282, i_10_4546, i_10_4565, o_10_304);
	kernel_10_305 k_10_305(i_10_32, i_10_152, i_10_157, i_10_174, i_10_179, i_10_256, i_10_257, i_10_262, i_10_266, i_10_281, i_10_394, i_10_410, i_10_430, i_10_440, i_10_441, i_10_464, i_10_548, i_10_796, i_10_800, i_10_962, i_10_1003, i_10_1004, i_10_1031, i_10_1039, i_10_1084, i_10_1234, i_10_1236, i_10_1250, i_10_1344, i_10_1432, i_10_1433, i_10_1546, i_10_1555, i_10_1556, i_10_1655, i_10_1687, i_10_1689, i_10_1690, i_10_1813, i_10_1826, i_10_1915, i_10_1945, i_10_1946, i_10_1948, i_10_2332, i_10_2356, i_10_2382, i_10_2448, i_10_2452, i_10_2456, i_10_2468, i_10_2516, i_10_2519, i_10_2628, i_10_2632, i_10_2633, i_10_2636, i_10_2657, i_10_2660, i_10_2707, i_10_2719, i_10_2721, i_10_2727, i_10_2730, i_10_2731, i_10_2781, i_10_2785, i_10_2829, i_10_2830, i_10_2832, i_10_2833, i_10_3013, i_10_3033, i_10_3034, i_10_3076, i_10_3199, i_10_3200, i_10_3201, i_10_3316, i_10_3386, i_10_3469, i_10_3473, i_10_3493, i_10_3541, i_10_3587, i_10_3615, i_10_3626, i_10_3646, i_10_3841, i_10_3849, i_10_3850, i_10_3853, i_10_3859, i_10_3990, i_10_4052, i_10_4114, i_10_4115, i_10_4117, i_10_4121, i_10_4288, o_10_305);
	kernel_10_306 k_10_306(i_10_118, i_10_153, i_10_243, i_10_244, i_10_253, i_10_284, i_10_388, i_10_390, i_10_460, i_10_462, i_10_513, i_10_687, i_10_711, i_10_747, i_10_748, i_10_794, i_10_1000, i_10_1035, i_10_1242, i_10_1246, i_10_1261, i_10_1263, i_10_1307, i_10_1308, i_10_1359, i_10_1360, i_10_1530, i_10_1612, i_10_1647, i_10_1648, i_10_1650, i_10_1651, i_10_1652, i_10_1654, i_10_1674, i_10_1683, i_10_1711, i_10_1809, i_10_1810, i_10_1819, i_10_1822, i_10_1911, i_10_1913, i_10_2178, i_10_2179, i_10_2199, i_10_2202, i_10_2308, i_10_2349, i_10_2350, i_10_2355, i_10_2380, i_10_2406, i_10_2451, i_10_2452, i_10_2467, i_10_2513, i_10_2601, i_10_2628, i_10_2631, i_10_2658, i_10_2659, i_10_2660, i_10_2718, i_10_2721, i_10_2722, i_10_2727, i_10_2740, i_10_2817, i_10_2818, i_10_2820, i_10_2829, i_10_2834, i_10_2881, i_10_3088, i_10_3231, i_10_3386, i_10_3466, i_10_3519, i_10_3522, i_10_3583, i_10_3646, i_10_3647, i_10_3788, i_10_3834, i_10_3847, i_10_3848, i_10_3856, i_10_3889, i_10_3906, i_10_3980, i_10_4023, i_10_4113, i_10_4122, i_10_4267, i_10_4269, i_10_4273, i_10_4284, i_10_4287, i_10_4571, o_10_306);
	kernel_10_307 k_10_307(i_10_177, i_10_266, i_10_268, i_10_269, i_10_276, i_10_282, i_10_319, i_10_323, i_10_388, i_10_391, i_10_393, i_10_431, i_10_439, i_10_464, i_10_560, i_10_798, i_10_799, i_10_800, i_10_1026, i_10_1136, i_10_1233, i_10_1241, i_10_1246, i_10_1267, i_10_1308, i_10_1309, i_10_1310, i_10_1312, i_10_1582, i_10_1583, i_10_1655, i_10_1821, i_10_1822, i_10_1823, i_10_1912, i_10_1915, i_10_2006, i_10_2179, i_10_2354, i_10_2356, i_10_2357, i_10_2365, i_10_2452, i_10_2453, i_10_2471, i_10_2472, i_10_2473, i_10_2516, i_10_2611, i_10_2631, i_10_2632, i_10_2635, i_10_2663, i_10_2721, i_10_2722, i_10_2723, i_10_2731, i_10_2732, i_10_2733, i_10_2734, i_10_2735, i_10_2834, i_10_2883, i_10_2884, i_10_2923, i_10_3035, i_10_3037, i_10_3045, i_10_3048, i_10_3049, i_10_3151, i_10_3154, i_10_3155, i_10_3201, i_10_3388, i_10_3389, i_10_3472, i_10_3523, i_10_3613, i_10_3688, i_10_3780, i_10_3783, i_10_3785, i_10_3837, i_10_3847, i_10_3850, i_10_3851, i_10_3855, i_10_3984, i_10_3985, i_10_3986, i_10_4128, i_10_4129, i_10_4130, i_10_4271, i_10_4282, i_10_4290, i_10_4291, i_10_4568, i_10_4571, o_10_307);
	kernel_10_308 k_10_308(i_10_89, i_10_146, i_10_221, i_10_284, i_10_286, i_10_320, i_10_327, i_10_329, i_10_330, i_10_331, i_10_437, i_10_443, i_10_462, i_10_463, i_10_464, i_10_467, i_10_514, i_10_711, i_10_719, i_10_748, i_10_749, i_10_797, i_10_800, i_10_990, i_10_991, i_10_1036, i_10_1174, i_10_1235, i_10_1239, i_10_1240, i_10_1241, i_10_1263, i_10_1265, i_10_1310, i_10_1342, i_10_1397, i_10_1610, i_10_1685, i_10_1826, i_10_1908, i_10_1911, i_10_1916, i_10_1990, i_10_1998, i_10_2200, i_10_2201, i_10_2335, i_10_2354, i_10_2407, i_10_2454, i_10_2456, i_10_2470, i_10_2503, i_10_2516, i_10_2567, i_10_2602, i_10_2605, i_10_2606, i_10_2629, i_10_2630, i_10_2661, i_10_2716, i_10_2720, i_10_2722, i_10_2724, i_10_2729, i_10_2782, i_10_2817, i_10_2829, i_10_2883, i_10_2953, i_10_3087, i_10_3088, i_10_3128, i_10_3199, i_10_3201, i_10_3202, i_10_3267, i_10_3385, i_10_3404, i_10_3523, i_10_3544, i_10_3557, i_10_3613, i_10_3614, i_10_3720, i_10_3733, i_10_3837, i_10_3847, i_10_3856, i_10_3881, i_10_4115, i_10_4277, i_10_4280, i_10_4284, i_10_4289, i_10_4351, i_10_4432, i_10_4569, i_10_4570, o_10_308);
	kernel_10_309 k_10_309(i_10_175, i_10_218, i_10_244, i_10_245, i_10_409, i_10_410, i_10_436, i_10_439, i_10_445, i_10_459, i_10_467, i_10_507, i_10_796, i_10_896, i_10_990, i_10_991, i_10_992, i_10_997, i_10_1000, i_10_1003, i_10_1006, i_10_1042, i_10_1043, i_10_1234, i_10_1236, i_10_1308, i_10_1309, i_10_1310, i_10_1312, i_10_1487, i_10_1649, i_10_1652, i_10_1654, i_10_1690, i_10_1769, i_10_1819, i_10_1820, i_10_1821, i_10_1824, i_10_1909, i_10_1916, i_10_1951, i_10_1952, i_10_2185, i_10_2452, i_10_2453, i_10_2473, i_10_2566, i_10_2628, i_10_2629, i_10_2704, i_10_2723, i_10_2724, i_10_2782, i_10_2817, i_10_2829, i_10_2831, i_10_2832, i_10_2833, i_10_2884, i_10_2885, i_10_2917, i_10_3034, i_10_3070, i_10_3151, i_10_3197, i_10_3198, i_10_3200, i_10_3272, i_10_3326, i_10_3385, i_10_3407, i_10_3466, i_10_3467, i_10_3499, i_10_3523, i_10_3585, i_10_3589, i_10_3610, i_10_3613, i_10_3614, i_10_3616, i_10_3617, i_10_3689, i_10_3785, i_10_3788, i_10_3835, i_10_3843, i_10_3986, i_10_3991, i_10_3992, i_10_4113, i_10_4114, i_10_4115, i_10_4122, i_10_4123, i_10_4284, i_10_4287, i_10_4563, i_10_4564, o_10_309);
	kernel_10_310 k_10_310(i_10_33, i_10_247, i_10_248, i_10_249, i_10_282, i_10_283, i_10_287, i_10_430, i_10_435, i_10_436, i_10_438, i_10_444, i_10_445, i_10_449, i_10_462, i_10_465, i_10_466, i_10_517, i_10_747, i_10_748, i_10_754, i_10_795, i_10_796, i_10_956, i_10_959, i_10_1233, i_10_1243, i_10_1246, i_10_1267, i_10_1306, i_10_1311, i_10_1360, i_10_1442, i_10_1578, i_10_1651, i_10_1654, i_10_1684, i_10_1689, i_10_1823, i_10_2254, i_10_2304, i_10_2310, i_10_2311, i_10_2312, i_10_2350, i_10_2454, i_10_2473, i_10_2474, i_10_2628, i_10_2631, i_10_2632, i_10_2634, i_10_2705, i_10_2727, i_10_2728, i_10_2821, i_10_2881, i_10_2887, i_10_2888, i_10_2913, i_10_2916, i_10_2923, i_10_3033, i_10_3034, i_10_3036, i_10_3037, i_10_3038, i_10_3040, i_10_3041, i_10_3074, i_10_3196, i_10_3197, i_10_3198, i_10_3202, i_10_3280, i_10_3387, i_10_3390, i_10_3392, i_10_3402, i_10_3403, i_10_3469, i_10_3493, i_10_3497, i_10_3614, i_10_3615, i_10_3649, i_10_3727, i_10_3780, i_10_3781, i_10_3837, i_10_3860, i_10_3906, i_10_3907, i_10_3972, i_10_3994, i_10_4113, i_10_4278, i_10_4279, i_10_4462, i_10_4525, o_10_310);
	kernel_10_311 k_10_311(i_10_86, i_10_387, i_10_388, i_10_409, i_10_423, i_10_433, i_10_461, i_10_496, i_10_514, i_10_693, i_10_694, i_10_714, i_10_733, i_10_734, i_10_735, i_10_796, i_10_799, i_10_800, i_10_901, i_10_993, i_10_999, i_10_1037, i_10_1237, i_10_1238, i_10_1239, i_10_1278, i_10_1307, i_10_1341, i_10_1342, i_10_1343, i_10_1354, i_10_1549, i_10_1576, i_10_1621, i_10_1650, i_10_1651, i_10_1685, i_10_1714, i_10_1818, i_10_1825, i_10_1826, i_10_1908, i_10_1909, i_10_1910, i_10_1944, i_10_2080, i_10_2263, i_10_2312, i_10_2327, i_10_2349, i_10_2350, i_10_2351, i_10_2383, i_10_2448, i_10_2454, i_10_2458, i_10_2566, i_10_2632, i_10_2635, i_10_2636, i_10_2720, i_10_2721, i_10_2820, i_10_2821, i_10_2882, i_10_2884, i_10_2885, i_10_2983, i_10_3197, i_10_3276, i_10_3277, i_10_3385, i_10_3613, i_10_3614, i_10_3615, i_10_3616, i_10_3650, i_10_3837, i_10_3840, i_10_3842, i_10_3853, i_10_3856, i_10_3859, i_10_3888, i_10_3889, i_10_3891, i_10_3979, i_10_3988, i_10_4027, i_10_4113, i_10_4154, i_10_4176, i_10_4177, i_10_4216, i_10_4275, i_10_4288, i_10_4291, i_10_4568, i_10_4587, i_10_4592, o_10_311);
	kernel_10_312 k_10_312(i_10_118, i_10_218, i_10_282, i_10_283, i_10_287, i_10_316, i_10_407, i_10_409, i_10_432, i_10_433, i_10_434, i_10_435, i_10_437, i_10_448, i_10_799, i_10_800, i_10_962, i_10_1029, i_10_1030, i_10_1033, i_10_1241, i_10_1309, i_10_1310, i_10_1365, i_10_1556, i_10_1650, i_10_1651, i_10_1654, i_10_1684, i_10_1685, i_10_1821, i_10_1825, i_10_1996, i_10_2179, i_10_2349, i_10_2350, i_10_2351, i_10_2361, i_10_2364, i_10_2365, i_10_2407, i_10_2453, i_10_2458, i_10_2461, i_10_2463, i_10_2467, i_10_2474, i_10_2571, i_10_2611, i_10_2634, i_10_2657, i_10_2661, i_10_2701, i_10_2704, i_10_2707, i_10_2714, i_10_2721, i_10_2731, i_10_2733, i_10_2788, i_10_2821, i_10_2824, i_10_2825, i_10_2831, i_10_2881, i_10_2882, i_10_2919, i_10_3036, i_10_3037, i_10_3038, i_10_3041, i_10_3050, i_10_3088, i_10_3196, i_10_3199, i_10_3391, i_10_3403, i_10_3404, i_10_3583, i_10_3613, i_10_3614, i_10_3648, i_10_3786, i_10_3839, i_10_3840, i_10_3843, i_10_3855, i_10_3856, i_10_3857, i_10_3858, i_10_3859, i_10_3994, i_10_4128, i_10_4168, i_10_4170, i_10_4172, i_10_4267, i_10_4273, i_10_4565, i_10_4570, o_10_312);
	kernel_10_313 k_10_313(i_10_48, i_10_156, i_10_216, i_10_223, i_10_252, i_10_327, i_10_387, i_10_408, i_10_409, i_10_410, i_10_445, i_10_463, i_10_498, i_10_504, i_10_516, i_10_531, i_10_532, i_10_748, i_10_750, i_10_753, i_10_867, i_10_906, i_10_957, i_10_958, i_10_990, i_10_1084, i_10_1134, i_10_1162, i_10_1218, i_10_1221, i_10_1236, i_10_1238, i_10_1262, i_10_1263, i_10_1266, i_10_1290, i_10_1310, i_10_1312, i_10_1347, i_10_1348, i_10_1398, i_10_1485, i_10_1545, i_10_1655, i_10_1683, i_10_1690, i_10_1822, i_10_1848, i_10_1947, i_10_1999, i_10_2361, i_10_2380, i_10_2452, i_10_2541, i_10_2577, i_10_2632, i_10_2634, i_10_2657, i_10_2660, i_10_2661, i_10_2677, i_10_2723, i_10_2728, i_10_2817, i_10_2881, i_10_2979, i_10_2983, i_10_3038, i_10_3040, i_10_3231, i_10_3232, i_10_3276, i_10_3277, i_10_3279, i_10_3281, i_10_3283, i_10_3388, i_10_3391, i_10_3466, i_10_3467, i_10_3496, i_10_3522, i_10_3613, i_10_3614, i_10_3648, i_10_3684, i_10_3782, i_10_3785, i_10_3786, i_10_3852, i_10_3910, i_10_3979, i_10_4113, i_10_4114, i_10_4266, i_10_4270, i_10_4275, i_10_4290, i_10_4291, i_10_4584, o_10_313);
	kernel_10_314 k_10_314(i_10_174, i_10_179, i_10_220, i_10_221, i_10_224, i_10_283, i_10_321, i_10_371, i_10_501, i_10_734, i_10_799, i_10_957, i_10_958, i_10_1054, i_10_1234, i_10_1236, i_10_1237, i_10_1431, i_10_1432, i_10_1541, i_10_1544, i_10_1578, i_10_1626, i_10_1635, i_10_1651, i_10_1655, i_10_1683, i_10_1684, i_10_1689, i_10_1690, i_10_1714, i_10_1735, i_10_1804, i_10_1805, i_10_1807, i_10_2003, i_10_2019, i_10_2029, i_10_2200, i_10_2201, i_10_2330, i_10_2353, i_10_2365, i_10_2366, i_10_2452, i_10_2481, i_10_2599, i_10_2605, i_10_2628, i_10_2631, i_10_2716, i_10_2718, i_10_2730, i_10_2731, i_10_2732, i_10_2733, i_10_2734, i_10_2757, i_10_2886, i_10_2966, i_10_2968, i_10_3162, i_10_3269, i_10_3278, i_10_3280, i_10_3282, i_10_3283, i_10_3284, i_10_3315, i_10_3387, i_10_3410, i_10_3430, i_10_3468, i_10_3469, i_10_3525, i_10_3545, i_10_3583, i_10_3612, i_10_3646, i_10_3648, i_10_3649, i_10_3811, i_10_3841, i_10_3855, i_10_3913, i_10_3988, i_10_4051, i_10_4099, i_10_4113, i_10_4114, i_10_4121, i_10_4129, i_10_4130, i_10_4215, i_10_4276, i_10_4291, i_10_4306, i_10_4565, i_10_4567, i_10_4568, o_10_314);
	kernel_10_315 k_10_315(i_10_173, i_10_328, i_10_410, i_10_427, i_10_443, i_10_445, i_10_463, i_10_466, i_10_515, i_10_716, i_10_892, i_10_958, i_10_1027, i_10_1028, i_10_1237, i_10_1244, i_10_1246, i_10_1249, i_10_1308, i_10_1310, i_10_1312, i_10_1313, i_10_1541, i_10_1631, i_10_1652, i_10_1675, i_10_1676, i_10_1685, i_10_1687, i_10_1691, i_10_1820, i_10_1825, i_10_1910, i_10_1916, i_10_2026, i_10_2027, i_10_2243, i_10_2378, i_10_2468, i_10_2566, i_10_2567, i_10_2608, i_10_2635, i_10_2701, i_10_2711, i_10_2719, i_10_2720, i_10_2722, i_10_2723, i_10_2727, i_10_2728, i_10_2729, i_10_2731, i_10_2786, i_10_2829, i_10_2917, i_10_2919, i_10_2920, i_10_2924, i_10_2980, i_10_3042, i_10_3044, i_10_3277, i_10_3281, i_10_3385, i_10_3387, i_10_3389, i_10_3392, i_10_3539, i_10_3542, i_10_3586, i_10_3611, i_10_3646, i_10_3727, i_10_3787, i_10_3839, i_10_3843, i_10_3844, i_10_3846, i_10_3848, i_10_3851, i_10_3852, i_10_3855, i_10_3857, i_10_3906, i_10_3908, i_10_3979, i_10_4213, i_10_4216, i_10_4268, i_10_4271, i_10_4284, i_10_4285, i_10_4286, i_10_4288, i_10_4289, i_10_4290, i_10_4563, i_10_4564, i_10_4566, o_10_315);
	kernel_10_316 k_10_316(i_10_81, i_10_224, i_10_280, i_10_284, i_10_286, i_10_316, i_10_317, i_10_328, i_10_390, i_10_464, i_10_796, i_10_799, i_10_800, i_10_957, i_10_1000, i_10_1153, i_10_1236, i_10_1241, i_10_1248, i_10_1263, i_10_1267, i_10_1307, i_10_1308, i_10_1309, i_10_1310, i_10_1544, i_10_1575, i_10_1579, i_10_1655, i_10_1810, i_10_1821, i_10_2017, i_10_2197, i_10_2312, i_10_2349, i_10_2350, i_10_2351, i_10_2352, i_10_2353, i_10_2354, i_10_2355, i_10_2359, i_10_2377, i_10_2378, i_10_2379, i_10_2380, i_10_2381, i_10_2383, i_10_2407, i_10_2409, i_10_2448, i_10_2449, i_10_2452, i_10_2453, i_10_2454, i_10_2471, i_10_2503, i_10_2506, i_10_2507, i_10_2604, i_10_2605, i_10_2657, i_10_2659, i_10_2700, i_10_2701, i_10_2727, i_10_2880, i_10_2882, i_10_2919, i_10_2965, i_10_3280, i_10_3283, i_10_3384, i_10_3385, i_10_3403, i_10_3537, i_10_3586, i_10_3587, i_10_3610, i_10_3613, i_10_3616, i_10_3836, i_10_3841, i_10_3853, i_10_3854, i_10_3856, i_10_3890, i_10_3982, i_10_4113, i_10_4115, i_10_4119, i_10_4127, i_10_4168, i_10_4271, i_10_4276, i_10_4277, i_10_4288, i_10_4566, i_10_4567, i_10_4568, o_10_316);
	kernel_10_317 k_10_317(i_10_88, i_10_89, i_10_117, i_10_149, i_10_178, i_10_182, i_10_276, i_10_277, i_10_282, i_10_375, i_10_409, i_10_410, i_10_436, i_10_449, i_10_459, i_10_460, i_10_461, i_10_467, i_10_473, i_10_515, i_10_578, i_10_581, i_10_800, i_10_906, i_10_1010, i_10_1040, i_10_1041, i_10_1168, i_10_1233, i_10_1240, i_10_1241, i_10_1292, i_10_1310, i_10_1348, i_10_1634, i_10_1650, i_10_1724, i_10_1767, i_10_1773, i_10_1822, i_10_1823, i_10_1912, i_10_1950, i_10_1951, i_10_2038, i_10_2183, i_10_2308, i_10_2337, i_10_2351, i_10_2352, i_10_2353, i_10_2378, i_10_2408, i_10_2451, i_10_2470, i_10_2474, i_10_2509, i_10_2606, i_10_2638, i_10_2711, i_10_2715, i_10_2741, i_10_2788, i_10_2865, i_10_2914, i_10_2915, i_10_2924, i_10_2957, i_10_2983, i_10_3001, i_10_3041, i_10_3046, i_10_3208, i_10_3209, i_10_3272, i_10_3329, i_10_3432, i_10_3494, i_10_3500, i_10_3585, i_10_3588, i_10_3589, i_10_3617, i_10_3733, i_10_3785, i_10_3806, i_10_3855, i_10_3886, i_10_3895, i_10_3946, i_10_3967, i_10_4054, i_10_4182, i_10_4183, i_10_4270, i_10_4273, i_10_4274, i_10_4463, i_10_4477, i_10_4478, o_10_317);
	kernel_10_318 k_10_318(i_10_28, i_10_37, i_10_155, i_10_193, i_10_273, i_10_280, i_10_282, i_10_332, i_10_424, i_10_432, i_10_435, i_10_436, i_10_437, i_10_521, i_10_629, i_10_752, i_10_779, i_10_847, i_10_929, i_10_1095, i_10_1121, i_10_1129, i_10_1239, i_10_1266, i_10_1268, i_10_1315, i_10_1343, i_10_1355, i_10_1441, i_10_1548, i_10_1549, i_10_1552, i_10_1555, i_10_1766, i_10_1797, i_10_1813, i_10_1814, i_10_1817, i_10_1880, i_10_1992, i_10_2007, i_10_2206, i_10_2242, i_10_2243, i_10_2349, i_10_2351, i_10_2353, i_10_2355, i_10_2356, i_10_2432, i_10_2476, i_10_2541, i_10_2556, i_10_2565, i_10_2583, i_10_2606, i_10_2701, i_10_2720, i_10_2727, i_10_2728, i_10_2756, i_10_2803, i_10_2804, i_10_2844, i_10_2864, i_10_2883, i_10_2920, i_10_2954, i_10_3033, i_10_3089, i_10_3238, i_10_3276, i_10_3277, i_10_3312, i_10_3521, i_10_3523, i_10_3602, i_10_3700, i_10_3746, i_10_3748, i_10_3812, i_10_3854, i_10_3855, i_10_3882, i_10_3989, i_10_4007, i_10_4114, i_10_4115, i_10_4125, i_10_4147, i_10_4171, i_10_4304, i_10_4439, i_10_4457, i_10_4522, i_10_4525, i_10_4532, i_10_4573, i_10_4574, i_10_4591, o_10_318);
	kernel_10_319 k_10_319(i_10_28, i_10_30, i_10_147, i_10_259, i_10_292, i_10_387, i_10_390, i_10_391, i_10_462, i_10_501, i_10_633, i_10_642, i_10_961, i_10_999, i_10_1002, i_10_1056, i_10_1236, i_10_1237, i_10_1239, i_10_1365, i_10_1391, i_10_1431, i_10_1434, i_10_1578, i_10_1579, i_10_1614, i_10_1623, i_10_1650, i_10_1696, i_10_1731, i_10_1821, i_10_1915, i_10_1920, i_10_1923, i_10_1938, i_10_1951, i_10_1992, i_10_2204, i_10_2235, i_10_2267, i_10_2291, i_10_2325, i_10_2355, i_10_2365, i_10_2448, i_10_2454, i_10_2466, i_10_2469, i_10_2470, i_10_2478, i_10_2514, i_10_2565, i_10_2571, i_10_2590, i_10_2607, i_10_2679, i_10_2709, i_10_2733, i_10_2742, i_10_2781, i_10_2784, i_10_2833, i_10_2994, i_10_2995, i_10_3040, i_10_3042, i_10_3045, i_10_3235, i_10_3280, i_10_3283, i_10_3318, i_10_3384, i_10_3387, i_10_3450, i_10_3469, i_10_3471, i_10_3472, i_10_3500, i_10_3504, i_10_3562, i_10_3610, i_10_3616, i_10_3625, i_10_3774, i_10_3807, i_10_3876, i_10_3882, i_10_3942, i_10_3981, i_10_3982, i_10_4053, i_10_4098, i_10_4102, i_10_4113, i_10_4189, i_10_4219, i_10_4226, i_10_4289, i_10_4372, i_10_4585, o_10_319);
	kernel_10_320 k_10_320(i_10_223, i_10_224, i_10_269, i_10_281, i_10_316, i_10_319, i_10_323, i_10_328, i_10_410, i_10_433, i_10_435, i_10_444, i_10_445, i_10_447, i_10_464, i_10_465, i_10_518, i_10_749, i_10_993, i_10_1006, i_10_1042, i_10_1043, i_10_1081, i_10_1237, i_10_1238, i_10_1241, i_10_1246, i_10_1296, i_10_1308, i_10_1309, i_10_1310, i_10_1348, i_10_1363, i_10_1543, i_10_1579, i_10_1582, i_10_1628, i_10_1653, i_10_1821, i_10_1824, i_10_1825, i_10_1911, i_10_1912, i_10_1913, i_10_1990, i_10_2186, i_10_2358, i_10_2380, i_10_2383, i_10_2633, i_10_2635, i_10_2657, i_10_2659, i_10_2660, i_10_2707, i_10_2708, i_10_2710, i_10_2718, i_10_2732, i_10_2789, i_10_2817, i_10_2818, i_10_2819, i_10_2828, i_10_2882, i_10_2920, i_10_2921, i_10_2924, i_10_3033, i_10_3076, i_10_3155, i_10_3199, i_10_3276, i_10_3338, i_10_3386, i_10_3389, i_10_3407, i_10_3523, i_10_3544, i_10_3584, i_10_3612, i_10_3613, i_10_3614, i_10_3649, i_10_3785, i_10_3834, i_10_3847, i_10_3848, i_10_3850, i_10_3857, i_10_3907, i_10_3986, i_10_4116, i_10_4117, i_10_4118, i_10_4119, i_10_4120, i_10_4125, i_10_4564, i_10_4565, o_10_320);
	kernel_10_321 k_10_321(i_10_117, i_10_175, i_10_180, i_10_268, i_10_279, i_10_319, i_10_407, i_10_408, i_10_427, i_10_428, i_10_440, i_10_444, i_10_445, i_10_461, i_10_462, i_10_712, i_10_748, i_10_796, i_10_897, i_10_958, i_10_1005, i_10_1166, i_10_1233, i_10_1238, i_10_1242, i_10_1366, i_10_1367, i_10_1385, i_10_1444, i_10_1612, i_10_1654, i_10_1655, i_10_1683, i_10_1821, i_10_1822, i_10_1823, i_10_1824, i_10_1911, i_10_1946, i_10_2001, i_10_2004, i_10_2020, i_10_2199, i_10_2311, i_10_2355, i_10_2451, i_10_2452, i_10_2460, i_10_2629, i_10_2631, i_10_2633, i_10_2643, i_10_2662, i_10_2721, i_10_2730, i_10_2733, i_10_2830, i_10_2882, i_10_2885, i_10_2916, i_10_2917, i_10_2985, i_10_2986, i_10_3035, i_10_3036, i_10_3040, i_10_3087, i_10_3094, i_10_3195, i_10_3196, i_10_3280, i_10_3284, i_10_3403, i_10_3469, i_10_3497, i_10_3541, i_10_3590, i_10_3609, i_10_3614, i_10_3682, i_10_3683, i_10_3721, i_10_3843, i_10_3847, i_10_3855, i_10_3858, i_10_3859, i_10_3918, i_10_3980, i_10_3983, i_10_4113, i_10_4119, i_10_4120, i_10_4122, i_10_4183, i_10_4189, i_10_4275, i_10_4288, i_10_4517, i_10_4566, o_10_321);
	kernel_10_322 k_10_322(i_10_40, i_10_41, i_10_43, i_10_120, i_10_124, i_10_172, i_10_179, i_10_224, i_10_293, i_10_315, i_10_324, i_10_325, i_10_328, i_10_390, i_10_391, i_10_407, i_10_410, i_10_413, i_10_446, i_10_539, i_10_561, i_10_796, i_10_800, i_10_826, i_10_905, i_10_961, i_10_998, i_10_1006, i_10_1087, i_10_1157, i_10_1160, i_10_1239, i_10_1241, i_10_1307, i_10_1309, i_10_1310, i_10_1349, i_10_1364, i_10_1432, i_10_1448, i_10_1451, i_10_1649, i_10_1715, i_10_1874, i_10_1903, i_10_1921, i_10_1947, i_10_2267, i_10_2363, i_10_2365, i_10_2366, i_10_2411, i_10_2471, i_10_2510, i_10_2557, i_10_2561, i_10_2606, i_10_2609, i_10_2611, i_10_2616, i_10_2617, i_10_2629, i_10_2632, i_10_2702, i_10_2704, i_10_2705, i_10_2710, i_10_2735, i_10_2786, i_10_2823, i_10_2882, i_10_2920, i_10_2957, i_10_3047, i_10_3049, i_10_3090, i_10_3093, i_10_3236, i_10_3239, i_10_3292, i_10_3401, i_10_3473, i_10_3527, i_10_3563, i_10_3781, i_10_3793, i_10_3811, i_10_3812, i_10_3835, i_10_3836, i_10_4052, i_10_4055, i_10_4121, i_10_4130, i_10_4171, i_10_4175, i_10_4281, i_10_4372, i_10_4571, i_10_4586, o_10_322);
	kernel_10_323 k_10_323(i_10_175, i_10_178, i_10_287, i_10_315, i_10_405, i_10_496, i_10_506, i_10_638, i_10_766, i_10_796, i_10_797, i_10_821, i_10_874, i_10_899, i_10_1000, i_10_1001, i_10_1103, i_10_1112, i_10_1207, i_10_1211, i_10_1235, i_10_1240, i_10_1274, i_10_1283, i_10_1301, i_10_1306, i_10_1363, i_10_1400, i_10_1541, i_10_1562, i_10_1565, i_10_1634, i_10_1688, i_10_1724, i_10_1729, i_10_1733, i_10_1799, i_10_1802, i_10_1804, i_10_1805, i_10_1916, i_10_1981, i_10_1984, i_10_2006, i_10_2186, i_10_2198, i_10_2201, i_10_2237, i_10_2249, i_10_2258, i_10_2566, i_10_2714, i_10_2717, i_10_2722, i_10_2728, i_10_2729, i_10_2747, i_10_2848, i_10_2890, i_10_2915, i_10_2965, i_10_2966, i_10_2975, i_10_3025, i_10_3053, i_10_3233, i_10_3281, i_10_3293, i_10_3296, i_10_3384, i_10_3433, i_10_3436, i_10_3470, i_10_3503, i_10_3539, i_10_3542, i_10_3566, i_10_3569, i_10_3586, i_10_3587, i_10_3620, i_10_3646, i_10_3682, i_10_3715, i_10_3787, i_10_3793, i_10_3796, i_10_3803, i_10_3839, i_10_3844, i_10_4007, i_10_4028, i_10_4150, i_10_4168, i_10_4169, i_10_4277, i_10_4547, i_10_4570, i_10_4571, i_10_4586, o_10_323);
	kernel_10_324 k_10_324(i_10_220, i_10_223, i_10_247, i_10_248, i_10_446, i_10_462, i_10_520, i_10_733, i_10_736, i_10_797, i_10_927, i_10_928, i_10_929, i_10_971, i_10_1028, i_10_1040, i_10_1083, i_10_1117, i_10_1233, i_10_1236, i_10_1237, i_10_1239, i_10_1243, i_10_1305, i_10_1306, i_10_1342, i_10_1446, i_10_1546, i_10_1547, i_10_1549, i_10_1551, i_10_1552, i_10_1648, i_10_1649, i_10_1683, i_10_1684, i_10_1685, i_10_1688, i_10_1691, i_10_1818, i_10_1819, i_10_1823, i_10_1826, i_10_1910, i_10_1915, i_10_1916, i_10_1991, i_10_2006, i_10_2309, i_10_2353, i_10_2357, i_10_2362, i_10_2379, i_10_2380, i_10_2430, i_10_2450, i_10_2451, i_10_2452, i_10_2569, i_10_2573, i_10_2725, i_10_2727, i_10_2832, i_10_2923, i_10_3072, i_10_3073, i_10_3087, i_10_3195, i_10_3196, i_10_3278, i_10_3385, i_10_3388, i_10_3391, i_10_3407, i_10_3433, i_10_3538, i_10_3550, i_10_3551, i_10_3586, i_10_3612, i_10_3648, i_10_3649, i_10_3650, i_10_3787, i_10_3838, i_10_3839, i_10_3847, i_10_3848, i_10_3855, i_10_3856, i_10_4009, i_10_4027, i_10_4057, i_10_4153, i_10_4175, i_10_4286, i_10_4375, i_10_4376, i_10_4564, i_10_4568, o_10_324);
	kernel_10_325 k_10_325(i_10_31, i_10_33, i_10_40, i_10_43, i_10_151, i_10_222, i_10_248, i_10_251, i_10_285, i_10_286, i_10_287, i_10_318, i_10_319, i_10_409, i_10_410, i_10_412, i_10_413, i_10_428, i_10_434, i_10_436, i_10_437, i_10_439, i_10_520, i_10_964, i_10_996, i_10_997, i_10_1004, i_10_1030, i_10_1041, i_10_1042, i_10_1043, i_10_1169, i_10_1236, i_10_1294, i_10_1311, i_10_1343, i_10_1344, i_10_1346, i_10_1546, i_10_1653, i_10_1655, i_10_1735, i_10_1815, i_10_1880, i_10_1908, i_10_1909, i_10_1913, i_10_2023, i_10_2245, i_10_2352, i_10_2353, i_10_2354, i_10_2355, i_10_2365, i_10_2452, i_10_2453, i_10_2455, i_10_2469, i_10_2471, i_10_2705, i_10_2724, i_10_2731, i_10_2832, i_10_2833, i_10_2869, i_10_2886, i_10_2887, i_10_3036, i_10_3037, i_10_3039, i_10_3045, i_10_3164, i_10_3166, i_10_3272, i_10_3280, i_10_3301, i_10_3433, i_10_3523, i_10_3526, i_10_3527, i_10_3585, i_10_3586, i_10_3611, i_10_3613, i_10_3616, i_10_3650, i_10_3784, i_10_3838, i_10_3893, i_10_3994, i_10_3995, i_10_4030, i_10_4116, i_10_4117, i_10_4172, i_10_4220, i_10_4273, i_10_4274, i_10_4282, i_10_4283, o_10_325);
	kernel_10_326 k_10_326(i_10_171, i_10_174, i_10_221, i_10_244, i_10_263, i_10_280, i_10_282, i_10_283, i_10_320, i_10_390, i_10_393, i_10_406, i_10_409, i_10_445, i_10_446, i_10_448, i_10_451, i_10_460, i_10_466, i_10_560, i_10_589, i_10_699, i_10_748, i_10_797, i_10_906, i_10_954, i_10_1002, i_10_1005, i_10_1027, i_10_1032, i_10_1238, i_10_1305, i_10_1307, i_10_1348, i_10_1447, i_10_1626, i_10_1651, i_10_1652, i_10_1655, i_10_1767, i_10_1768, i_10_1769, i_10_1818, i_10_1819, i_10_1821, i_10_1824, i_10_1910, i_10_1911, i_10_1949, i_10_1995, i_10_2310, i_10_2334, i_10_2376, i_10_2384, i_10_2460, i_10_2461, i_10_2565, i_10_2647, i_10_2658, i_10_2679, i_10_2704, i_10_2718, i_10_2721, i_10_2728, i_10_2826, i_10_2829, i_10_2830, i_10_2831, i_10_2921, i_10_2924, i_10_3157, i_10_3280, i_10_3386, i_10_3387, i_10_3388, i_10_3403, i_10_3436, i_10_3437, i_10_3540, i_10_3541, i_10_3550, i_10_3610, i_10_3835, i_10_3853, i_10_3854, i_10_3855, i_10_3856, i_10_3860, i_10_3984, i_10_4025, i_10_4026, i_10_4027, i_10_4117, i_10_4118, i_10_4120, i_10_4122, i_10_4128, i_10_4174, i_10_4548, i_10_4571, o_10_326);
	kernel_10_327 k_10_327(i_10_32, i_10_158, i_10_185, i_10_284, i_10_390, i_10_391, i_10_392, i_10_436, i_10_437, i_10_443, i_10_464, i_10_718, i_10_854, i_10_955, i_10_961, i_10_964, i_10_992, i_10_1003, i_10_1036, i_10_1043, i_10_1045, i_10_1058, i_10_1082, i_10_1083, i_10_1120, i_10_1240, i_10_1247, i_10_1268, i_10_1365, i_10_1366, i_10_1367, i_10_1380, i_10_1436, i_10_1443, i_10_1448, i_10_1489, i_10_1597, i_10_1651, i_10_1772, i_10_1797, i_10_1806, i_10_1919, i_10_1954, i_10_2018, i_10_2095, i_10_2096, i_10_2349, i_10_2357, i_10_2362, i_10_2366, i_10_2381, i_10_2465, i_10_2492, i_10_2511, i_10_2514, i_10_2560, i_10_2565, i_10_2603, i_10_2659, i_10_2660, i_10_2702, i_10_2743, i_10_2744, i_10_2781, i_10_2782, i_10_2831, i_10_2834, i_10_3159, i_10_3162, i_10_3283, i_10_3284, i_10_3450, i_10_3452, i_10_3470, i_10_3703, i_10_3704, i_10_3747, i_10_3835, i_10_3853, i_10_3879, i_10_3923, i_10_4056, i_10_4057, i_10_4114, i_10_4144, i_10_4220, i_10_4237, i_10_4238, i_10_4268, i_10_4275, i_10_4278, i_10_4280, i_10_4282, i_10_4342, i_10_4436, i_10_4521, i_10_4522, i_10_4523, i_10_4565, i_10_4571, o_10_327);
	kernel_10_328 k_10_328(i_10_48, i_10_174, i_10_175, i_10_220, i_10_279, i_10_282, i_10_283, i_10_329, i_10_445, i_10_446, i_10_459, i_10_460, i_10_462, i_10_463, i_10_685, i_10_686, i_10_748, i_10_828, i_10_963, i_10_990, i_10_997, i_10_1026, i_10_1035, i_10_1036, i_10_1161, i_10_1162, i_10_1266, i_10_1268, i_10_1288, i_10_1306, i_10_1307, i_10_1486, i_10_1532, i_10_1551, i_10_1562, i_10_1647, i_10_1648, i_10_1649, i_10_1683, i_10_1766, i_10_1823, i_10_1825, i_10_1917, i_10_1946, i_10_2353, i_10_2448, i_10_2451, i_10_2452, i_10_2454, i_10_2472, i_10_2473, i_10_2503, i_10_2539, i_10_2603, i_10_2605, i_10_2629, i_10_2630, i_10_2632, i_10_2657, i_10_2658, i_10_2661, i_10_2726, i_10_2727, i_10_2787, i_10_2817, i_10_2820, i_10_2822, i_10_2826, i_10_2827, i_10_2828, i_10_2880, i_10_2881, i_10_3034, i_10_3035, i_10_3282, i_10_3312, i_10_3313, i_10_3384, i_10_3388, i_10_3522, i_10_3523, i_10_3525, i_10_3526, i_10_3646, i_10_3840, i_10_3980, i_10_3987, i_10_3998, i_10_4113, i_10_4115, i_10_4117, i_10_4168, i_10_4275, i_10_4284, i_10_4285, i_10_4287, i_10_4288, i_10_4456, i_10_4563, i_10_4564, o_10_328);
	kernel_10_329 k_10_329(i_10_175, i_10_267, i_10_281, i_10_284, i_10_286, i_10_393, i_10_405, i_10_406, i_10_408, i_10_409, i_10_412, i_10_439, i_10_444, i_10_447, i_10_448, i_10_462, i_10_467, i_10_713, i_10_793, i_10_798, i_10_1002, i_10_1005, i_10_1054, i_10_1061, i_10_1122, i_10_1215, i_10_1239, i_10_1247, i_10_1249, i_10_1296, i_10_1313, i_10_1437, i_10_1542, i_10_1626, i_10_1650, i_10_1684, i_10_1685, i_10_1686, i_10_1728, i_10_1730, i_10_1768, i_10_1821, i_10_1914, i_10_1915, i_10_1952, i_10_2025, i_10_2029, i_10_2324, i_10_2327, i_10_2355, i_10_2453, i_10_2454, i_10_2455, i_10_2469, i_10_2517, i_10_2565, i_10_2628, i_10_2632, i_10_2634, i_10_2636, i_10_2655, i_10_2658, i_10_2659, i_10_2662, i_10_2663, i_10_2678, i_10_2702, i_10_2704, i_10_2706, i_10_2711, i_10_2725, i_10_2730, i_10_2732, i_10_2737, i_10_2784, i_10_2785, i_10_2804, i_10_2954, i_10_2979, i_10_2996, i_10_3033, i_10_3071, i_10_3279, i_10_3284, i_10_3320, i_10_3388, i_10_3389, i_10_3471, i_10_3525, i_10_3545, i_10_3561, i_10_3586, i_10_3613, i_10_3780, i_10_3784, i_10_3837, i_10_3859, i_10_4117, i_10_4124, i_10_4272, o_10_329);
	kernel_10_330 k_10_330(i_10_33, i_10_34, i_10_123, i_10_143, i_10_256, i_10_265, i_10_266, i_10_272, i_10_274, i_10_275, i_10_283, i_10_432, i_10_448, i_10_449, i_10_498, i_10_501, i_10_502, i_10_506, i_10_564, i_10_565, i_10_628, i_10_719, i_10_745, i_10_753, i_10_1005, i_10_1030, i_10_1034, i_10_1111, i_10_1115, i_10_1165, i_10_1213, i_10_1240, i_10_1243, i_10_1261, i_10_1302, i_10_1303, i_10_1326, i_10_1348, i_10_1435, i_10_1439, i_10_1542, i_10_1583, i_10_1732, i_10_1820, i_10_1821, i_10_1950, i_10_1959, i_10_2035, i_10_2204, i_10_2294, i_10_2350, i_10_2351, i_10_2354, i_10_2355, i_10_2408, i_10_2515, i_10_2533, i_10_2560, i_10_2714, i_10_2744, i_10_2760, i_10_2761, i_10_2785, i_10_2839, i_10_2840, i_10_2851, i_10_2869, i_10_2870, i_10_2885, i_10_2968, i_10_2969, i_10_3048, i_10_3049, i_10_3195, i_10_3200, i_10_3337, i_10_3388, i_10_3435, i_10_3504, i_10_3543, i_10_3544, i_10_3649, i_10_3651, i_10_3747, i_10_3797, i_10_3804, i_10_3853, i_10_3857, i_10_3984, i_10_4000, i_10_4117, i_10_4210, i_10_4211, i_10_4269, i_10_4272, i_10_4273, i_10_4291, i_10_4392, i_10_4564, i_10_4589, o_10_330);
	kernel_10_331 k_10_331(i_10_49, i_10_173, i_10_409, i_10_460, i_10_464, i_10_496, i_10_700, i_10_712, i_10_713, i_10_718, i_10_748, i_10_749, i_10_752, i_10_893, i_10_949, i_10_1028, i_10_1163, i_10_1235, i_10_1236, i_10_1237, i_10_1264, i_10_1306, i_10_1307, i_10_1308, i_10_1309, i_10_1310, i_10_1313, i_10_1577, i_10_1612, i_10_1684, i_10_1685, i_10_1688, i_10_1766, i_10_1812, i_10_1813, i_10_1821, i_10_2180, i_10_2359, i_10_2448, i_10_2467, i_10_2526, i_10_2606, i_10_2631, i_10_2641, i_10_2657, i_10_2660, i_10_2701, i_10_2702, i_10_2711, i_10_2719, i_10_2720, i_10_2728, i_10_2733, i_10_2818, i_10_2830, i_10_2831, i_10_2833, i_10_2884, i_10_2885, i_10_2921, i_10_2923, i_10_3070, i_10_3233, i_10_3268, i_10_3269, i_10_3280, i_10_3297, i_10_3385, i_10_3386, i_10_3390, i_10_3391, i_10_3392, i_10_3406, i_10_3462, i_10_3523, i_10_3585, i_10_3613, i_10_3614, i_10_3647, i_10_3649, i_10_3650, i_10_3727, i_10_3732, i_10_3781, i_10_3782, i_10_3783, i_10_3784, i_10_3787, i_10_3835, i_10_3837, i_10_3888, i_10_3909, i_10_4115, i_10_4125, i_10_4169, i_10_4212, i_10_4285, i_10_4286, i_10_4518, i_10_4565, o_10_331);
	kernel_10_332 k_10_332(i_10_11, i_10_254, i_10_320, i_10_344, i_10_392, i_10_394, i_10_433, i_10_464, i_10_497, i_10_821, i_10_824, i_10_931, i_10_1100, i_10_1210, i_10_1220, i_10_1235, i_10_1238, i_10_1297, i_10_1298, i_10_1300, i_10_1307, i_10_1433, i_10_1540, i_10_1541, i_10_1622, i_10_1625, i_10_1684, i_10_1685, i_10_1688, i_10_1730, i_10_1733, i_10_1805, i_10_1822, i_10_1825, i_10_1985, i_10_1990, i_10_2108, i_10_2162, i_10_2201, i_10_2288, i_10_2345, i_10_2351, i_10_2358, i_10_2359, i_10_2360, i_10_2408, i_10_2466, i_10_2467, i_10_2470, i_10_2507, i_10_2530, i_10_2558, i_10_2561, i_10_2566, i_10_2567, i_10_2570, i_10_2606, i_10_2632, i_10_2638, i_10_2641, i_10_2702, i_10_2705, i_10_2710, i_10_2722, i_10_2729, i_10_2755, i_10_2852, i_10_2963, i_10_3043, i_10_3070, i_10_3290, i_10_3317, i_10_3332, i_10_3461, i_10_3503, i_10_3539, i_10_3545, i_10_3548, i_10_3556, i_10_3557, i_10_3584, i_10_3586, i_10_3835, i_10_3836, i_10_3839, i_10_3847, i_10_3848, i_10_3854, i_10_3908, i_10_4007, i_10_4060, i_10_4123, i_10_4154, i_10_4169, i_10_4172, i_10_4267, i_10_4277, i_10_4429, i_10_4433, i_10_4566, o_10_332);
	kernel_10_333 k_10_333(i_10_14, i_10_35, i_10_80, i_10_160, i_10_223, i_10_268, i_10_269, i_10_296, i_10_410, i_10_413, i_10_439, i_10_440, i_10_463, i_10_511, i_10_512, i_10_692, i_10_755, i_10_872, i_10_1033, i_10_1034, i_10_1041, i_10_1042, i_10_1043, i_10_1052, i_10_1059, i_10_1139, i_10_1157, i_10_1160, i_10_1175, i_10_1205, i_10_1241, i_10_1249, i_10_1294, i_10_1303, i_10_1312, i_10_1348, i_10_1356, i_10_1362, i_10_1366, i_10_1367, i_10_1439, i_10_1457, i_10_1545, i_10_1546, i_10_1547, i_10_1582, i_10_1583, i_10_1627, i_10_1651, i_10_1655, i_10_1690, i_10_1733, i_10_1735, i_10_1736, i_10_1772, i_10_1781, i_10_1817, i_10_1850, i_10_1913, i_10_1915, i_10_1984, i_10_1987, i_10_1988, i_10_2356, i_10_2453, i_10_2467, i_10_2560, i_10_2609, i_10_2660, i_10_2702, i_10_2723, i_10_2743, i_10_2816, i_10_2829, i_10_2830, i_10_2839, i_10_2851, i_10_2965, i_10_2968, i_10_2969, i_10_2987, i_10_3049, i_10_3274, i_10_3392, i_10_3409, i_10_3437, i_10_3508, i_10_3544, i_10_3614, i_10_3859, i_10_3984, i_10_3985, i_10_4117, i_10_4118, i_10_4119, i_10_4238, i_10_4288, i_10_4462, i_10_4570, i_10_4571, o_10_333);
	kernel_10_334 k_10_334(i_10_13, i_10_15, i_10_16, i_10_22, i_10_39, i_10_40, i_10_121, i_10_160, i_10_281, i_10_286, i_10_433, i_10_434, i_10_513, i_10_514, i_10_595, i_10_598, i_10_635, i_10_661, i_10_691, i_10_800, i_10_872, i_10_907, i_10_1060, i_10_1159, i_10_1169, i_10_1175, i_10_1399, i_10_1439, i_10_1487, i_10_1542, i_10_1545, i_10_1713, i_10_1850, i_10_1877, i_10_1879, i_10_1880, i_10_2020, i_10_2023, i_10_2024, i_10_2029, i_10_2030, i_10_2037, i_10_2112, i_10_2203, i_10_2204, i_10_2222, i_10_2243, i_10_2245, i_10_2380, i_10_2410, i_10_2411, i_10_2467, i_10_2468, i_10_2472, i_10_2598, i_10_2599, i_10_2608, i_10_2616, i_10_2660, i_10_2663, i_10_2678, i_10_2707, i_10_2708, i_10_2711, i_10_2714, i_10_2722, i_10_2733, i_10_2735, i_10_2789, i_10_2821, i_10_2824, i_10_2884, i_10_2885, i_10_2987, i_10_3046, i_10_3072, i_10_3075, i_10_3076, i_10_3077, i_10_3109, i_10_3163, i_10_3199, i_10_3407, i_10_3469, i_10_3472, i_10_3473, i_10_3522, i_10_3586, i_10_3589, i_10_3590, i_10_3622, i_10_3653, i_10_3683, i_10_3724, i_10_3839, i_10_3909, i_10_3910, i_10_4121, i_10_4124, i_10_4526, o_10_334);
	kernel_10_335 k_10_335(i_10_146, i_10_175, i_10_284, i_10_407, i_10_441, i_10_442, i_10_443, i_10_444, i_10_793, i_10_794, i_10_800, i_10_964, i_10_966, i_10_1117, i_10_1205, i_10_1264, i_10_1307, i_10_1308, i_10_1346, i_10_1575, i_10_1620, i_10_1636, i_10_1647, i_10_1651, i_10_1652, i_10_1683, i_10_1684, i_10_1685, i_10_1820, i_10_1826, i_10_1915, i_10_1947, i_10_2000, i_10_2158, i_10_2159, i_10_2333, i_10_2350, i_10_2352, i_10_2454, i_10_2470, i_10_2514, i_10_2556, i_10_2631, i_10_2632, i_10_2701, i_10_2711, i_10_2719, i_10_2789, i_10_2831, i_10_2850, i_10_2884, i_10_2888, i_10_2920, i_10_2921, i_10_2923, i_10_2924, i_10_2952, i_10_2979, i_10_3090, i_10_3239, i_10_3270, i_10_3387, i_10_3388, i_10_3391, i_10_3406, i_10_3434, i_10_3522, i_10_3523, i_10_3524, i_10_3525, i_10_3526, i_10_3527, i_10_3590, i_10_3610, i_10_3611, i_10_3613, i_10_3614, i_10_3682, i_10_3683, i_10_3704, i_10_3730, i_10_3783, i_10_3835, i_10_3844, i_10_3854, i_10_3860, i_10_3995, i_10_4191, i_10_4192, i_10_4215, i_10_4216, i_10_4218, i_10_4269, i_10_4290, i_10_4291, i_10_4459, i_10_4460, i_10_4462, i_10_4560, i_10_4570, o_10_335);
	kernel_10_336 k_10_336(i_10_70, i_10_71, i_10_174, i_10_175, i_10_278, i_10_286, i_10_328, i_10_329, i_10_442, i_10_445, i_10_446, i_10_448, i_10_449, i_10_466, i_10_505, i_10_623, i_10_700, i_10_794, i_10_958, i_10_960, i_10_961, i_10_1031, i_10_1043, i_10_1233, i_10_1239, i_10_1308, i_10_1312, i_10_1313, i_10_1347, i_10_1348, i_10_1349, i_10_1547, i_10_1556, i_10_1653, i_10_1684, i_10_1717, i_10_1718, i_10_1768, i_10_1822, i_10_1823, i_10_1824, i_10_1825, i_10_1877, i_10_1991, i_10_2021, i_10_2166, i_10_2167, i_10_2198, i_10_2200, i_10_2363, i_10_2382, i_10_2449, i_10_2450, i_10_2452, i_10_2460, i_10_2461, i_10_2631, i_10_2634, i_10_2661, i_10_2663, i_10_2703, i_10_2704, i_10_2716, i_10_2717, i_10_2722, i_10_2723, i_10_2733, i_10_2734, i_10_2825, i_10_2829, i_10_2887, i_10_2923, i_10_2924, i_10_3046, i_10_3047, i_10_3076, i_10_3077, i_10_3151, i_10_3153, i_10_3284, i_10_3388, i_10_3389, i_10_3390, i_10_3391, i_10_3392, i_10_3434, i_10_3472, i_10_3616, i_10_3617, i_10_3650, i_10_3653, i_10_3775, i_10_3786, i_10_3835, i_10_3841, i_10_3851, i_10_3856, i_10_4117, i_10_4287, i_10_4571, o_10_336);
	kernel_10_337 k_10_337(i_10_276, i_10_282, i_10_320, i_10_321, i_10_328, i_10_442, i_10_443, i_10_447, i_10_448, i_10_462, i_10_514, i_10_516, i_10_519, i_10_561, i_10_718, i_10_795, i_10_798, i_10_969, i_10_970, i_10_993, i_10_1164, i_10_1234, i_10_1438, i_10_1445, i_10_1492, i_10_1578, i_10_1581, i_10_1641, i_10_1652, i_10_1653, i_10_1807, i_10_1815, i_10_1822, i_10_1946, i_10_2030, i_10_2182, i_10_2251, i_10_2308, i_10_2310, i_10_2311, i_10_2349, i_10_2350, i_10_2351, i_10_2352, i_10_2353, i_10_2356, i_10_2383, i_10_2410, i_10_2450, i_10_2454, i_10_2544, i_10_2634, i_10_2676, i_10_2717, i_10_2724, i_10_2727, i_10_2730, i_10_2743, i_10_2784, i_10_2785, i_10_2955, i_10_2982, i_10_2985, i_10_2986, i_10_3040, i_10_3091, i_10_3102, i_10_3103, i_10_3120, i_10_3156, i_10_3198, i_10_3232, i_10_3283, i_10_3298, i_10_3468, i_10_3493, i_10_3494, i_10_3496, i_10_3525, i_10_3588, i_10_3611, i_10_3649, i_10_3653, i_10_3786, i_10_3805, i_10_3857, i_10_3874, i_10_3896, i_10_3949, i_10_3979, i_10_4113, i_10_4117, i_10_4119, i_10_4146, i_10_4266, i_10_4270, i_10_4271, i_10_4281, i_10_4285, i_10_4288, o_10_337);
	kernel_10_338 k_10_338(i_10_171, i_10_172, i_10_177, i_10_220, i_10_223, i_10_271, i_10_272, i_10_274, i_10_282, i_10_318, i_10_427, i_10_430, i_10_435, i_10_438, i_10_442, i_10_446, i_10_463, i_10_711, i_10_712, i_10_1030, i_10_1037, i_10_1238, i_10_1305, i_10_1311, i_10_1343, i_10_1346, i_10_1548, i_10_1549, i_10_1551, i_10_1552, i_10_1651, i_10_1652, i_10_1654, i_10_1655, i_10_1683, i_10_1764, i_10_1765, i_10_1819, i_10_1822, i_10_1824, i_10_1910, i_10_2197, i_10_2358, i_10_2381, i_10_2382, i_10_2383, i_10_2410, i_10_2635, i_10_2636, i_10_2662, i_10_2704, i_10_2707, i_10_2710, i_10_2712, i_10_2728, i_10_2731, i_10_2732, i_10_2783, i_10_2821, i_10_2832, i_10_2880, i_10_2883, i_10_2884, i_10_2885, i_10_2886, i_10_2887, i_10_2888, i_10_3040, i_10_3070, i_10_3151, i_10_3198, i_10_3277, i_10_3326, i_10_3384, i_10_3385, i_10_3386, i_10_3387, i_10_3405, i_10_3406, i_10_3409, i_10_3410, i_10_3588, i_10_3614, i_10_3684, i_10_3842, i_10_3856, i_10_3857, i_10_3859, i_10_3860, i_10_3891, i_10_3983, i_10_3994, i_10_3995, i_10_4118, i_10_4126, i_10_4287, i_10_4288, i_10_4290, i_10_4292, i_10_4594, o_10_338);
	kernel_10_339 k_10_339(i_10_255, i_10_277, i_10_280, i_10_281, i_10_315, i_10_318, i_10_322, i_10_387, i_10_393, i_10_406, i_10_408, i_10_441, i_10_442, i_10_462, i_10_465, i_10_519, i_10_747, i_10_795, i_10_798, i_10_963, i_10_1026, i_10_1029, i_10_1241, i_10_1308, i_10_1362, i_10_1431, i_10_1434, i_10_1435, i_10_1444, i_10_1539, i_10_1540, i_10_1542, i_10_1545, i_10_1578, i_10_1626, i_10_1648, i_10_1683, i_10_1684, i_10_1686, i_10_1689, i_10_1719, i_10_1806, i_10_1819, i_10_1821, i_10_1823, i_10_1826, i_10_2028, i_10_2179, i_10_2180, i_10_2349, i_10_2350, i_10_2407, i_10_2451, i_10_2469, i_10_2628, i_10_2631, i_10_2632, i_10_2636, i_10_2656, i_10_2659, i_10_2660, i_10_2661, i_10_2728, i_10_2731, i_10_2733, i_10_2785, i_10_2829, i_10_2880, i_10_2921, i_10_2967, i_10_3034, i_10_3069, i_10_3072, i_10_3151, i_10_3153, i_10_3154, i_10_3270, i_10_3271, i_10_3280, i_10_3318, i_10_3325, i_10_3336, i_10_3468, i_10_3523, i_10_3543, i_10_3615, i_10_3648, i_10_3835, i_10_3837, i_10_3847, i_10_3909, i_10_3910, i_10_3993, i_10_3994, i_10_4118, i_10_4170, i_10_4270, i_10_4272, i_10_4275, i_10_4566, o_10_339);
	kernel_10_340 k_10_340(i_10_34, i_10_61, i_10_259, i_10_273, i_10_282, i_10_283, i_10_284, i_10_301, i_10_444, i_10_637, i_10_642, i_10_717, i_10_718, i_10_755, i_10_958, i_10_962, i_10_1030, i_10_1034, i_10_1243, i_10_1248, i_10_1249, i_10_1250, i_10_1265, i_10_1309, i_10_1385, i_10_1448, i_10_1546, i_10_1547, i_10_1582, i_10_1619, i_10_1689, i_10_1690, i_10_1691, i_10_1760, i_10_1824, i_10_1825, i_10_1961, i_10_2167, i_10_2168, i_10_2185, i_10_2186, i_10_2199, i_10_2203, i_10_2204, i_10_2273, i_10_2338, i_10_2352, i_10_2355, i_10_2356, i_10_2357, i_10_2472, i_10_2536, i_10_2609, i_10_2632, i_10_2662, i_10_2694, i_10_2955, i_10_3038, i_10_3075, i_10_3076, i_10_3177, i_10_3199, i_10_3202, i_10_3239, i_10_3268, i_10_3274, i_10_3275, i_10_3306, i_10_3337, i_10_3389, i_10_3390, i_10_3434, i_10_3468, i_10_3551, i_10_3613, i_10_3626, i_10_3650, i_10_3734, i_10_3786, i_10_3795, i_10_3810, i_10_3814, i_10_3815, i_10_3846, i_10_3847, i_10_3848, i_10_3850, i_10_3851, i_10_3856, i_10_3877, i_10_4000, i_10_4013, i_10_4116, i_10_4119, i_10_4120, i_10_4174, i_10_4220, i_10_4264, i_10_4292, i_10_4585, o_10_340);
	kernel_10_341 k_10_341(i_10_30, i_10_34, i_10_175, i_10_282, i_10_283, i_10_319, i_10_390, i_10_410, i_10_412, i_10_445, i_10_466, i_10_542, i_10_714, i_10_798, i_10_799, i_10_954, i_10_958, i_10_968, i_10_1026, i_10_1027, i_10_1028, i_10_1029, i_10_1233, i_10_1234, i_10_1264, i_10_1265, i_10_1305, i_10_1306, i_10_1313, i_10_1542, i_10_1596, i_10_1653, i_10_1655, i_10_1691, i_10_1824, i_10_1825, i_10_2006, i_10_2016, i_10_2081, i_10_2185, i_10_2198, i_10_2307, i_10_2310, i_10_2350, i_10_2352, i_10_2353, i_10_2361, i_10_2471, i_10_2629, i_10_2635, i_10_2657, i_10_2677, i_10_2713, i_10_2714, i_10_2718, i_10_2726, i_10_2739, i_10_2824, i_10_2829, i_10_2922, i_10_2952, i_10_3033, i_10_3034, i_10_3076, i_10_3231, i_10_3232, i_10_3270, i_10_3331, i_10_3333, i_10_3429, i_10_3546, i_10_3616, i_10_3617, i_10_3626, i_10_3649, i_10_3650, i_10_3689, i_10_3718, i_10_3780, i_10_3783, i_10_3784, i_10_3786, i_10_3787, i_10_3788, i_10_3808, i_10_3810, i_10_3811, i_10_3843, i_10_3844, i_10_3846, i_10_3854, i_10_4115, i_10_4116, i_10_4119, i_10_4121, i_10_4122, i_10_4123, i_10_4126, i_10_4167, i_10_4275, o_10_341);
	kernel_10_342 k_10_342(i_10_48, i_10_51, i_10_52, i_10_219, i_10_221, i_10_223, i_10_267, i_10_284, i_10_286, i_10_295, i_10_461, i_10_462, i_10_463, i_10_699, i_10_796, i_10_852, i_10_897, i_10_898, i_10_1037, i_10_1050, i_10_1113, i_10_1195, i_10_1250, i_10_1346, i_10_1435, i_10_1575, i_10_1616, i_10_1623, i_10_1685, i_10_1688, i_10_1771, i_10_1821, i_10_1824, i_10_2211, i_10_2263, i_10_2357, i_10_2365, i_10_2438, i_10_2454, i_10_2455, i_10_2465, i_10_2474, i_10_2514, i_10_2515, i_10_2568, i_10_2631, i_10_2632, i_10_2641, i_10_2652, i_10_2653, i_10_2705, i_10_2712, i_10_2715, i_10_2723, i_10_2828, i_10_2832, i_10_2885, i_10_2888, i_10_2923, i_10_2924, i_10_2982, i_10_2986, i_10_3093, i_10_3094, i_10_3270, i_10_3273, i_10_3275, i_10_3276, i_10_3277, i_10_3390, i_10_3391, i_10_3392, i_10_3407, i_10_3561, i_10_3612, i_10_3613, i_10_3617, i_10_3732, i_10_3839, i_10_3841, i_10_3847, i_10_3855, i_10_3856, i_10_3858, i_10_3892, i_10_3893, i_10_3894, i_10_3982, i_10_3983, i_10_3985, i_10_3992, i_10_4027, i_10_4029, i_10_4031, i_10_4120, i_10_4154, i_10_4156, i_10_4218, i_10_4219, i_10_4506, o_10_342);
	kernel_10_343 k_10_343(i_10_37, i_10_63, i_10_91, i_10_221, i_10_261, i_10_292, i_10_327, i_10_413, i_10_440, i_10_464, i_10_585, i_10_589, i_10_632, i_10_697, i_10_725, i_10_733, i_10_792, i_10_793, i_10_832, i_10_833, i_10_877, i_10_891, i_10_892, i_10_920, i_10_931, i_10_964, i_10_967, i_10_968, i_10_970, i_10_1008, i_10_1029, i_10_1031, i_10_1117, i_10_1163, i_10_1216, i_10_1270, i_10_1288, i_10_1291, i_10_1310, i_10_1311, i_10_1363, i_10_1687, i_10_1766, i_10_1801, i_10_1810, i_10_1819, i_10_1823, i_10_1980, i_10_1999, i_10_2002, i_10_2224, i_10_2308, i_10_2351, i_10_2407, i_10_2449, i_10_2489, i_10_2517, i_10_2518, i_10_2539, i_10_2565, i_10_2678, i_10_2710, i_10_2721, i_10_2722, i_10_2821, i_10_2822, i_10_2980, i_10_2984, i_10_3010, i_10_3013, i_10_3274, i_10_3298, i_10_3331, i_10_3332, i_10_3349, i_10_3470, i_10_3539, i_10_3587, i_10_3610, i_10_3622, i_10_3623, i_10_3651, i_10_3685, i_10_3820, i_10_3970, i_10_3992, i_10_3997, i_10_4009, i_10_4060, i_10_4061, i_10_4118, i_10_4226, i_10_4387, i_10_4429, i_10_4522, i_10_4525, i_10_4571, i_10_4582, i_10_4583, i_10_4588, o_10_343);
	kernel_10_344 k_10_344(i_10_86, i_10_144, i_10_149, i_10_172, i_10_173, i_10_184, i_10_185, i_10_253, i_10_254, i_10_311, i_10_374, i_10_423, i_10_424, i_10_428, i_10_465, i_10_560, i_10_692, i_10_734, i_10_779, i_10_792, i_10_900, i_10_901, i_10_923, i_10_963, i_10_997, i_10_1003, i_10_1030, i_10_1053, i_10_1123, i_10_1162, i_10_1205, i_10_1328, i_10_1486, i_10_1654, i_10_1683, i_10_1685, i_10_1768, i_10_1792, i_10_1801, i_10_1854, i_10_1864, i_10_1905, i_10_1942, i_10_1949, i_10_2002, i_10_2090, i_10_2255, i_10_2356, i_10_2383, i_10_2450, i_10_2453, i_10_2461, i_10_2479, i_10_2513, i_10_2531, i_10_2578, i_10_2663, i_10_2709, i_10_2713, i_10_2722, i_10_2727, i_10_2740, i_10_2783, i_10_2804, i_10_2823, i_10_2827, i_10_2880, i_10_2887, i_10_2998, i_10_3007, i_10_3119, i_10_3197, i_10_3231, i_10_3290, i_10_3386, i_10_3451, i_10_3452, i_10_3466, i_10_3493, i_10_3501, i_10_3552, i_10_3589, i_10_3590, i_10_3616, i_10_3702, i_10_3788, i_10_3838, i_10_3858, i_10_3880, i_10_3883, i_10_3943, i_10_4055, i_10_4114, i_10_4115, i_10_4213, i_10_4217, i_10_4220, i_10_4281, i_10_4340, i_10_4451, o_10_344);
	kernel_10_345 k_10_345(i_10_269, i_10_283, i_10_284, i_10_286, i_10_327, i_10_408, i_10_409, i_10_410, i_10_413, i_10_441, i_10_444, i_10_520, i_10_521, i_10_718, i_10_793, i_10_797, i_10_1237, i_10_1238, i_10_1299, i_10_1310, i_10_1312, i_10_1313, i_10_1552, i_10_1555, i_10_1652, i_10_1819, i_10_1824, i_10_1826, i_10_1995, i_10_1996, i_10_2022, i_10_2185, i_10_2197, i_10_2200, i_10_2311, i_10_2312, i_10_2332, i_10_2352, i_10_2353, i_10_2354, i_10_2361, i_10_2376, i_10_2377, i_10_2378, i_10_2382, i_10_2383, i_10_2407, i_10_2410, i_10_2411, i_10_2462, i_10_2628, i_10_2632, i_10_2633, i_10_2658, i_10_2661, i_10_2718, i_10_2735, i_10_2782, i_10_2785, i_10_2788, i_10_2827, i_10_2828, i_10_2831, i_10_2922, i_10_2923, i_10_2924, i_10_2983, i_10_2986, i_10_3049, i_10_3050, i_10_3203, i_10_3271, i_10_3272, i_10_3282, i_10_3387, i_10_3389, i_10_3391, i_10_3392, i_10_3405, i_10_3408, i_10_3497, i_10_3652, i_10_3846, i_10_3847, i_10_3848, i_10_3851, i_10_3857, i_10_3858, i_10_3859, i_10_3895, i_10_3986, i_10_4129, i_10_4269, i_10_4270, i_10_4271, i_10_4277, i_10_4292, i_10_4567, i_10_4568, i_10_4569, o_10_345);
	kernel_10_346 k_10_346(i_10_86, i_10_172, i_10_173, i_10_181, i_10_185, i_10_326, i_10_446, i_10_449, i_10_499, i_10_588, i_10_591, i_10_800, i_10_971, i_10_1234, i_10_1238, i_10_1246, i_10_1273, i_10_1363, i_10_1367, i_10_1412, i_10_1543, i_10_1553, i_10_1648, i_10_1651, i_10_1655, i_10_1760, i_10_1765, i_10_1777, i_10_1819, i_10_1820, i_10_1822, i_10_1825, i_10_1886, i_10_1888, i_10_1909, i_10_1949, i_10_2093, i_10_2096, i_10_2311, i_10_2336, i_10_2339, i_10_2448, i_10_2449, i_10_2450, i_10_2456, i_10_2543, i_10_2606, i_10_2638, i_10_2642, i_10_2702, i_10_2703, i_10_2725, i_10_2731, i_10_2788, i_10_2833, i_10_2866, i_10_2867, i_10_2869, i_10_2870, i_10_2917, i_10_2920, i_10_2923, i_10_3033, i_10_3037, i_10_3040, i_10_3092, i_10_3196, i_10_3197, i_10_3199, i_10_3202, i_10_3203, i_10_3386, i_10_3390, i_10_3392, i_10_3471, i_10_3586, i_10_3587, i_10_3588, i_10_3589, i_10_3611, i_10_3683, i_10_3731, i_10_3734, i_10_3884, i_10_3923, i_10_3964, i_10_3965, i_10_4117, i_10_4118, i_10_4120, i_10_4180, i_10_4267, i_10_4274, i_10_4283, i_10_4310, i_10_4561, i_10_4588, i_10_4592, i_10_4603, i_10_4604, o_10_346);
	kernel_10_347 k_10_347(i_10_247, i_10_330, i_10_393, i_10_405, i_10_423, i_10_424, i_10_438, i_10_442, i_10_444, i_10_459, i_10_463, i_10_464, i_10_467, i_10_507, i_10_562, i_10_711, i_10_792, i_10_956, i_10_1026, i_10_1305, i_10_1438, i_10_1548, i_10_1579, i_10_1654, i_10_1655, i_10_1683, i_10_1819, i_10_1821, i_10_1913, i_10_2202, i_10_2337, i_10_2350, i_10_2351, i_10_2352, i_10_2353, i_10_2354, i_10_2355, i_10_2365, i_10_2379, i_10_2451, i_10_2452, i_10_2571, i_10_2633, i_10_2634, i_10_2658, i_10_2701, i_10_2710, i_10_2732, i_10_2733, i_10_2781, i_10_2830, i_10_2883, i_10_2884, i_10_2888, i_10_2922, i_10_2985, i_10_3038, i_10_3048, i_10_3087, i_10_3152, i_10_3154, i_10_3165, i_10_3198, i_10_3199, i_10_3277, i_10_3280, i_10_3283, i_10_3385, i_10_3386, i_10_3405, i_10_3406, i_10_3408, i_10_3471, i_10_3610, i_10_3612, i_10_3613, i_10_3616, i_10_3702, i_10_3834, i_10_3837, i_10_3847, i_10_3850, i_10_3851, i_10_3855, i_10_3894, i_10_3982, i_10_4027, i_10_4116, i_10_4117, i_10_4120, i_10_4125, i_10_4126, i_10_4127, i_10_4285, i_10_4292, i_10_4563, i_10_4564, i_10_4566, i_10_4567, i_10_4568, o_10_347);
	kernel_10_348 k_10_348(i_10_171, i_10_174, i_10_175, i_10_184, i_10_220, i_10_223, i_10_247, i_10_265, i_10_269, i_10_270, i_10_271, i_10_273, i_10_283, i_10_284, i_10_287, i_10_395, i_10_405, i_10_408, i_10_412, i_10_436, i_10_798, i_10_958, i_10_1004, i_10_1006, i_10_1085, i_10_1310, i_10_1434, i_10_1435, i_10_1438, i_10_1451, i_10_1547, i_10_1554, i_10_1555, i_10_1619, i_10_1877, i_10_1945, i_10_1947, i_10_1948, i_10_1949, i_10_1951, i_10_1952, i_10_2185, i_10_2310, i_10_2312, i_10_2350, i_10_2353, i_10_2354, i_10_2356, i_10_2357, i_10_2407, i_10_2408, i_10_2411, i_10_2449, i_10_2470, i_10_2471, i_10_2510, i_10_2663, i_10_2681, i_10_2730, i_10_2781, i_10_2821, i_10_2920, i_10_2921, i_10_2923, i_10_2924, i_10_3034, i_10_3047, i_10_3050, i_10_3077, i_10_3090, i_10_3151, i_10_3157, i_10_3199, i_10_3272, i_10_3275, i_10_3281, i_10_3301, i_10_3384, i_10_3385, i_10_3392, i_10_3472, i_10_3473, i_10_3545, i_10_3560, i_10_3586, i_10_3588, i_10_3590, i_10_3784, i_10_3859, i_10_3895, i_10_3986, i_10_4054, i_10_4115, i_10_4116, i_10_4117, i_10_4118, i_10_4273, i_10_4283, i_10_4285, i_10_4567, o_10_348);
	kernel_10_349 k_10_349(i_10_17, i_10_67, i_10_118, i_10_245, i_10_252, i_10_279, i_10_281, i_10_317, i_10_320, i_10_325, i_10_326, i_10_389, i_10_395, i_10_410, i_10_428, i_10_434, i_10_442, i_10_464, i_10_506, i_10_792, i_10_968, i_10_994, i_10_1098, i_10_1235, i_10_1307, i_10_1311, i_10_1313, i_10_1343, i_10_1379, i_10_1454, i_10_1456, i_10_1544, i_10_1547, i_10_1576, i_10_1625, i_10_1655, i_10_1985, i_10_1993, i_10_1994, i_10_1997, i_10_2201, i_10_2203, i_10_2443, i_10_2444, i_10_2448, i_10_2450, i_10_2455, i_10_2456, i_10_2471, i_10_2529, i_10_2534, i_10_2584, i_10_2592, i_10_2639, i_10_2703, i_10_2705, i_10_2713, i_10_2716, i_10_2717, i_10_2828, i_10_2830, i_10_2834, i_10_2867, i_10_2870, i_10_2881, i_10_2882, i_10_2884, i_10_2885, i_10_2984, i_10_3041, i_10_3277, i_10_3278, i_10_3317, i_10_3384, i_10_3388, i_10_3409, i_10_3452, i_10_3523, i_10_3610, i_10_3611, i_10_3615, i_10_3653, i_10_3700, i_10_3703, i_10_3775, i_10_3836, i_10_3837, i_10_3857, i_10_3860, i_10_3912, i_10_3914, i_10_3983, i_10_4163, i_10_4175, i_10_4214, i_10_4273, i_10_4283, i_10_4288, i_10_4588, i_10_4592, o_10_349);
	kernel_10_350 k_10_350(i_10_27, i_10_220, i_10_249, i_10_282, i_10_284, i_10_293, i_10_327, i_10_412, i_10_428, i_10_517, i_10_518, i_10_520, i_10_798, i_10_800, i_10_955, i_10_957, i_10_961, i_10_1033, i_10_1035, i_10_1152, i_10_1243, i_10_1245, i_10_1246, i_10_1247, i_10_1310, i_10_1311, i_10_1384, i_10_1539, i_10_1617, i_10_1683, i_10_1686, i_10_1690, i_10_1691, i_10_1820, i_10_1822, i_10_1825, i_10_1908, i_10_1911, i_10_1912, i_10_2186, i_10_2349, i_10_2350, i_10_2360, i_10_2361, i_10_2406, i_10_2452, i_10_2467, i_10_2468, i_10_2470, i_10_2473, i_10_2655, i_10_2679, i_10_2719, i_10_2725, i_10_2726, i_10_2740, i_10_2827, i_10_3036, i_10_3048, i_10_3074, i_10_3075, i_10_3201, i_10_3269, i_10_3387, i_10_3391, i_10_3392, i_10_3453, i_10_3520, i_10_3523, i_10_3609, i_10_3612, i_10_3613, i_10_3614, i_10_3617, i_10_3624, i_10_3648, i_10_3651, i_10_3652, i_10_3706, i_10_3723, i_10_3730, i_10_3780, i_10_3834, i_10_3835, i_10_3839, i_10_3840, i_10_3860, i_10_3993, i_10_4114, i_10_4120, i_10_4126, i_10_4215, i_10_4216, i_10_4219, i_10_4236, i_10_4273, i_10_4291, i_10_4563, i_10_4566, i_10_4568, o_10_350);
	kernel_10_351 k_10_351(i_10_131, i_10_182, i_10_220, i_10_307, i_10_350, i_10_361, i_10_374, i_10_388, i_10_433, i_10_560, i_10_563, i_10_566, i_10_716, i_10_751, i_10_819, i_10_907, i_10_931, i_10_955, i_10_1046, i_10_1049, i_10_1084, i_10_1237, i_10_1247, i_10_1305, i_10_1308, i_10_1309, i_10_1310, i_10_1454, i_10_1488, i_10_1489, i_10_1543, i_10_1616, i_10_1648, i_10_1649, i_10_1652, i_10_1654, i_10_1688, i_10_1689, i_10_1864, i_10_2026, i_10_2038, i_10_2061, i_10_2080, i_10_2081, i_10_2201, i_10_2254, i_10_2514, i_10_2515, i_10_2533, i_10_2610, i_10_2657, i_10_2660, i_10_2729, i_10_2731, i_10_2740, i_10_2741, i_10_2830, i_10_2999, i_10_3039, i_10_3070, i_10_3292, i_10_3388, i_10_3389, i_10_3492, i_10_3542, i_10_3583, i_10_3587, i_10_3618, i_10_3646, i_10_3647, i_10_3649, i_10_3650, i_10_3682, i_10_3788, i_10_3807, i_10_3853, i_10_3854, i_10_3856, i_10_3857, i_10_3910, i_10_3911, i_10_3978, i_10_3979, i_10_4051, i_10_4052, i_10_4054, i_10_4055, i_10_4113, i_10_4114, i_10_4117, i_10_4191, i_10_4216, i_10_4311, i_10_4394, i_10_4400, i_10_4451, i_10_4528, i_10_4529, i_10_4531, i_10_4567, o_10_351);
	kernel_10_352 k_10_352(i_10_281, i_10_282, i_10_284, i_10_293, i_10_320, i_10_322, i_10_328, i_10_329, i_10_405, i_10_409, i_10_410, i_10_412, i_10_436, i_10_445, i_10_446, i_10_448, i_10_466, i_10_467, i_10_796, i_10_959, i_10_960, i_10_961, i_10_991, i_10_992, i_10_994, i_10_996, i_10_1233, i_10_1237, i_10_1263, i_10_1264, i_10_1309, i_10_1348, i_10_1653, i_10_1769, i_10_1819, i_10_1820, i_10_1821, i_10_1822, i_10_1876, i_10_1877, i_10_1912, i_10_1913, i_10_1989, i_10_1990, i_10_2351, i_10_2352, i_10_2357, i_10_2362, i_10_2382, i_10_2383, i_10_2456, i_10_2603, i_10_2634, i_10_2655, i_10_2656, i_10_2657, i_10_2659, i_10_2663, i_10_2713, i_10_2714, i_10_2715, i_10_2716, i_10_2717, i_10_2718, i_10_2719, i_10_2722, i_10_2730, i_10_2819, i_10_2826, i_10_2827, i_10_2829, i_10_2830, i_10_2883, i_10_2919, i_10_2923, i_10_2981, i_10_3034, i_10_3035, i_10_3037, i_10_3070, i_10_3076, i_10_3094, i_10_3385, i_10_3388, i_10_3390, i_10_3406, i_10_3407, i_10_3434, i_10_3520, i_10_3521, i_10_3523, i_10_3610, i_10_3834, i_10_3835, i_10_3855, i_10_3859, i_10_4268, i_10_4271, i_10_4277, i_10_4570, o_10_352);
	kernel_10_353 k_10_353(i_10_43, i_10_44, i_10_49, i_10_89, i_10_176, i_10_179, i_10_224, i_10_248, i_10_279, i_10_281, i_10_282, i_10_295, i_10_316, i_10_317, i_10_319, i_10_320, i_10_328, i_10_412, i_10_413, i_10_434, i_10_441, i_10_467, i_10_643, i_10_715, i_10_716, i_10_795, i_10_796, i_10_896, i_10_898, i_10_958, i_10_997, i_10_1004, i_10_1236, i_10_1238, i_10_1241, i_10_1244, i_10_1247, i_10_1261, i_10_1262, i_10_1313, i_10_1365, i_10_1366, i_10_1645, i_10_1654, i_10_1687, i_10_1732, i_10_1824, i_10_1994, i_10_1999, i_10_2002, i_10_2005, i_10_2024, i_10_2057, i_10_2165, i_10_2351, i_10_2362, i_10_2363, i_10_2365, i_10_2366, i_10_2377, i_10_2449, i_10_2467, i_10_2470, i_10_2471, i_10_2603, i_10_2630, i_10_2675, i_10_2678, i_10_2680, i_10_2723, i_10_2725, i_10_2785, i_10_2786, i_10_2884, i_10_2981, i_10_3074, i_10_3077, i_10_3272, i_10_3613, i_10_3616, i_10_3617, i_10_3721, i_10_3722, i_10_3809, i_10_3841, i_10_3853, i_10_3875, i_10_3911, i_10_3949, i_10_3993, i_10_3994, i_10_3995, i_10_4115, i_10_4117, i_10_4120, i_10_4121, i_10_4130, i_10_4175, i_10_4220, i_10_4276, o_10_353);
	kernel_10_354 k_10_354(i_10_83, i_10_89, i_10_172, i_10_177, i_10_187, i_10_188, i_10_214, i_10_224, i_10_283, i_10_284, i_10_318, i_10_371, i_10_406, i_10_410, i_10_413, i_10_446, i_10_799, i_10_800, i_10_906, i_10_907, i_10_908, i_10_919, i_10_920, i_10_1237, i_10_1238, i_10_1239, i_10_1240, i_10_1245, i_10_1249, i_10_1250, i_10_1367, i_10_1618, i_10_1651, i_10_1686, i_10_1687, i_10_1688, i_10_1767, i_10_1768, i_10_1802, i_10_1888, i_10_1907, i_10_1909, i_10_1912, i_10_1914, i_10_1940, i_10_1951, i_10_1952, i_10_1960, i_10_2020, i_10_2312, i_10_2452, i_10_2455, i_10_2462, i_10_2463, i_10_2464, i_10_2509, i_10_2629, i_10_2632, i_10_2634, i_10_2707, i_10_2708, i_10_2730, i_10_2732, i_10_2758, i_10_2783, i_10_2922, i_10_2924, i_10_3011, i_10_3014, i_10_3038, i_10_3185, i_10_3198, i_10_3199, i_10_3320, i_10_3387, i_10_3613, i_10_3614, i_10_3689, i_10_3707, i_10_3839, i_10_3857, i_10_3884, i_10_3887, i_10_3895, i_10_3967, i_10_3982, i_10_4183, i_10_4184, i_10_4193, i_10_4270, i_10_4272, i_10_4273, i_10_4274, i_10_4279, i_10_4298, i_10_4534, i_10_4567, i_10_4568, i_10_4606, i_10_4607, o_10_354);
	kernel_10_355 k_10_355(i_10_27, i_10_48, i_10_49, i_10_130, i_10_144, i_10_145, i_10_172, i_10_176, i_10_283, i_10_324, i_10_495, i_10_513, i_10_586, i_10_587, i_10_623, i_10_711, i_10_733, i_10_792, i_10_795, i_10_821, i_10_918, i_10_963, i_10_981, i_10_999, i_10_1027, i_10_1044, i_10_1081, i_10_1161, i_10_1215, i_10_1216, i_10_1218, i_10_1236, i_10_1237, i_10_1280, i_10_1446, i_10_1476, i_10_1477, i_10_1478, i_10_1548, i_10_1617, i_10_1639, i_10_1764, i_10_1812, i_10_1822, i_10_1911, i_10_1915, i_10_1953, i_10_1956, i_10_1990, i_10_1998, i_10_2089, i_10_2179, i_10_2180, i_10_2199, i_10_2201, i_10_2304, i_10_2410, i_10_2485, i_10_2493, i_10_2631, i_10_2659, i_10_2662, i_10_2688, i_10_2922, i_10_2955, i_10_2981, i_10_3070, i_10_3097, i_10_3114, i_10_3115, i_10_3277, i_10_3278, i_10_3312, i_10_3331, i_10_3348, i_10_3439, i_10_3492, i_10_3493, i_10_3539, i_10_3589, i_10_3645, i_10_3646, i_10_3794, i_10_3871, i_10_3879, i_10_3997, i_10_4007, i_10_4059, i_10_4060, i_10_4063, i_10_4114, i_10_4126, i_10_4267, i_10_4286, i_10_4293, i_10_4294, i_10_4311, i_10_4314, i_10_4581, i_10_4582, o_10_355);
	kernel_10_356 k_10_356(i_10_122, i_10_124, i_10_175, i_10_220, i_10_246, i_10_248, i_10_319, i_10_423, i_10_426, i_10_427, i_10_442, i_10_445, i_10_459, i_10_460, i_10_461, i_10_463, i_10_464, i_10_466, i_10_795, i_10_800, i_10_896, i_10_956, i_10_959, i_10_1030, i_10_1233, i_10_1234, i_10_1241, i_10_1312, i_10_1362, i_10_1379, i_10_1381, i_10_1445, i_10_1541, i_10_1551, i_10_1552, i_10_1579, i_10_1583, i_10_1654, i_10_1690, i_10_1825, i_10_1826, i_10_1909, i_10_1948, i_10_2203, i_10_2350, i_10_2351, i_10_2353, i_10_2360, i_10_2377, i_10_2452, i_10_2459, i_10_2467, i_10_2471, i_10_2629, i_10_2660, i_10_2661, i_10_2710, i_10_2713, i_10_2721, i_10_2725, i_10_2728, i_10_2731, i_10_2830, i_10_2831, i_10_2917, i_10_3037, i_10_3038, i_10_3046, i_10_3075, i_10_3196, i_10_3199, i_10_3202, i_10_3270, i_10_3271, i_10_3272, i_10_3281, i_10_3387, i_10_3388, i_10_3467, i_10_3493, i_10_3611, i_10_3613, i_10_3647, i_10_3650, i_10_3781, i_10_3785, i_10_3835, i_10_3837, i_10_3838, i_10_3844, i_10_3845, i_10_3846, i_10_3853, i_10_3855, i_10_3880, i_10_4121, i_10_4267, i_10_4269, i_10_4279, i_10_4286, o_10_356);
	kernel_10_357 k_10_357(i_10_145, i_10_151, i_10_178, i_10_179, i_10_186, i_10_284, i_10_285, i_10_443, i_10_445, i_10_446, i_10_449, i_10_465, i_10_466, i_10_519, i_10_520, i_10_719, i_10_755, i_10_793, i_10_798, i_10_799, i_10_966, i_10_967, i_10_971, i_10_997, i_10_1026, i_10_1166, i_10_1242, i_10_1246, i_10_1247, i_10_1250, i_10_1308, i_10_1309, i_10_1363, i_10_1537, i_10_1543, i_10_1580, i_10_1582, i_10_1583, i_10_1613, i_10_1616, i_10_1617, i_10_1686, i_10_1819, i_10_2004, i_10_2005, i_10_2248, i_10_2359, i_10_2361, i_10_2456, i_10_2607, i_10_2634, i_10_2635, i_10_2637, i_10_2638, i_10_2660, i_10_2701, i_10_2703, i_10_2704, i_10_2705, i_10_2718, i_10_2719, i_10_2725, i_10_2727, i_10_2729, i_10_2923, i_10_3039, i_10_3041, i_10_3198, i_10_3199, i_10_3200, i_10_3276, i_10_3277, i_10_3278, i_10_3392, i_10_3410, i_10_3493, i_10_3617, i_10_3721, i_10_3783, i_10_3785, i_10_3788, i_10_3848, i_10_3856, i_10_3857, i_10_3899, i_10_3913, i_10_3914, i_10_4027, i_10_4087, i_10_4117, i_10_4118, i_10_4119, i_10_4121, i_10_4150, i_10_4267, i_10_4269, i_10_4273, i_10_4289, i_10_4462, i_10_4527, o_10_357);
	kernel_10_358 k_10_358(i_10_66, i_10_119, i_10_121, i_10_175, i_10_181, i_10_287, i_10_316, i_10_346, i_10_432, i_10_433, i_10_443, i_10_446, i_10_515, i_10_535, i_10_800, i_10_909, i_10_957, i_10_959, i_10_1008, i_10_1048, i_10_1055, i_10_1119, i_10_1187, i_10_1234, i_10_1288, i_10_1305, i_10_1361, i_10_1363, i_10_1364, i_10_1371, i_10_1447, i_10_1495, i_10_1581, i_10_1607, i_10_1746, i_10_1882, i_10_1949, i_10_1955, i_10_1979, i_10_2200, i_10_2308, i_10_2309, i_10_2354, i_10_2365, i_10_2458, i_10_2464, i_10_2476, i_10_2565, i_10_2566, i_10_2610, i_10_2641, i_10_2673, i_10_2677, i_10_2710, i_10_2711, i_10_2729, i_10_2731, i_10_2782, i_10_3008, i_10_3037, i_10_3043, i_10_3088, i_10_3202, i_10_3211, i_10_3222, i_10_3226, i_10_3238, i_10_3239, i_10_3267, i_10_3268, i_10_3291, i_10_3319, i_10_3350, i_10_3384, i_10_3447, i_10_3448, i_10_3549, i_10_3550, i_10_3551, i_10_3681, i_10_3686, i_10_3775, i_10_3835, i_10_3837, i_10_3879, i_10_3919, i_10_3980, i_10_3987, i_10_4052, i_10_4213, i_10_4232, i_10_4286, i_10_4306, i_10_4366, i_10_4369, i_10_4370, i_10_4455, i_10_4460, i_10_4563, i_10_4564, o_10_358);
	kernel_10_359 k_10_359(i_10_173, i_10_196, i_10_280, i_10_315, i_10_388, i_10_394, i_10_395, i_10_437, i_10_513, i_10_722, i_10_854, i_10_948, i_10_949, i_10_964, i_10_965, i_10_1035, i_10_1036, i_10_1112, i_10_1121, i_10_1131, i_10_1237, i_10_1308, i_10_1309, i_10_1353, i_10_1354, i_10_1357, i_10_1363, i_10_1435, i_10_1438, i_10_1579, i_10_1650, i_10_1652, i_10_1653, i_10_1820, i_10_1909, i_10_1912, i_10_1929, i_10_1947, i_10_1950, i_10_1984, i_10_1985, i_10_2016, i_10_2209, i_10_2351, i_10_2512, i_10_2651, i_10_2656, i_10_2657, i_10_2659, i_10_2695, i_10_2709, i_10_2710, i_10_2732, i_10_2754, i_10_2826, i_10_2828, i_10_2831, i_10_2832, i_10_2840, i_10_2880, i_10_2916, i_10_2918, i_10_2919, i_10_2920, i_10_2921, i_10_2922, i_10_3046, i_10_3087, i_10_3090, i_10_3235, i_10_3269, i_10_3272, i_10_3313, i_10_3315, i_10_3321, i_10_3356, i_10_3432, i_10_3538, i_10_3585, i_10_3610, i_10_3651, i_10_3652, i_10_3664, i_10_3699, i_10_3718, i_10_3775, i_10_3786, i_10_3811, i_10_3901, i_10_3981, i_10_3982, i_10_3984, i_10_4091, i_10_4118, i_10_4268, i_10_4285, i_10_4288, i_10_4290, i_10_4291, i_10_4593, o_10_359);
	kernel_10_360 k_10_360(i_10_177, i_10_178, i_10_279, i_10_282, i_10_283, i_10_296, i_10_328, i_10_329, i_10_410, i_10_438, i_10_459, i_10_466, i_10_467, i_10_506, i_10_509, i_10_799, i_10_955, i_10_1005, i_10_1006, i_10_1007, i_10_1236, i_10_1239, i_10_1248, i_10_1249, i_10_1263, i_10_1264, i_10_1305, i_10_1448, i_10_1551, i_10_1552, i_10_1554, i_10_1556, i_10_1582, i_10_1626, i_10_1651, i_10_1678, i_10_1683, i_10_1689, i_10_1691, i_10_1716, i_10_1822, i_10_1823, i_10_1825, i_10_1912, i_10_2204, i_10_2310, i_10_2311, i_10_2312, i_10_2352, i_10_2354, i_10_2357, i_10_2364, i_10_2408, i_10_2469, i_10_2470, i_10_2481, i_10_2633, i_10_2635, i_10_2661, i_10_2663, i_10_2704, i_10_2708, i_10_2715, i_10_2716, i_10_2717, i_10_2727, i_10_2731, i_10_2732, i_10_2735, i_10_2832, i_10_2923, i_10_3072, i_10_3157, i_10_3158, i_10_3279, i_10_3280, i_10_3386, i_10_3497, i_10_3501, i_10_3540, i_10_3543, i_10_3585, i_10_3586, i_10_3649, i_10_3650, i_10_3653, i_10_3784, i_10_3788, i_10_3847, i_10_3859, i_10_3895, i_10_3896, i_10_3906, i_10_3985, i_10_4116, i_10_4117, i_10_4118, i_10_4121, i_10_4236, i_10_4237, o_10_360);
	kernel_10_361 k_10_361(i_10_172, i_10_244, i_10_430, i_10_431, i_10_444, i_10_447, i_10_466, i_10_467, i_10_589, i_10_744, i_10_798, i_10_820, i_10_1007, i_10_1032, i_10_1043, i_10_1060, i_10_1061, i_10_1083, i_10_1132, i_10_1215, i_10_1233, i_10_1237, i_10_1241, i_10_1349, i_10_1580, i_10_1582, i_10_1648, i_10_1649, i_10_1652, i_10_1654, i_10_1684, i_10_1687, i_10_1690, i_10_1736, i_10_1772, i_10_1821, i_10_1822, i_10_2023, i_10_2201, i_10_2349, i_10_2352, i_10_2355, i_10_2374, i_10_2450, i_10_2468, i_10_2516, i_10_2584, i_10_2632, i_10_2634, i_10_2659, i_10_2701, i_10_2707, i_10_2727, i_10_2729, i_10_2741, i_10_2743, i_10_2829, i_10_2831, i_10_2919, i_10_2921, i_10_2923, i_10_3073, i_10_3075, i_10_3199, i_10_3271, i_10_3283, i_10_3326, i_10_3384, i_10_3387, i_10_3388, i_10_3390, i_10_3391, i_10_3468, i_10_3470, i_10_3522, i_10_3523, i_10_3544, i_10_3613, i_10_3615, i_10_3616, i_10_3617, i_10_3649, i_10_3668, i_10_3726, i_10_3784, i_10_3838, i_10_3848, i_10_3853, i_10_3855, i_10_3857, i_10_3990, i_10_4173, i_10_4174, i_10_4208, i_10_4238, i_10_4281, i_10_4287, i_10_4288, i_10_4289, i_10_4571, o_10_361);
	kernel_10_362 k_10_362(i_10_85, i_10_261, i_10_279, i_10_281, i_10_284, i_10_285, i_10_393, i_10_436, i_10_498, i_10_502, i_10_558, i_10_600, i_10_643, i_10_698, i_10_711, i_10_724, i_10_727, i_10_822, i_10_852, i_10_876, i_10_1029, i_10_1086, i_10_1133, i_10_1222, i_10_1239, i_10_1299, i_10_1332, i_10_1348, i_10_1434, i_10_1449, i_10_1542, i_10_1551, i_10_1579, i_10_1605, i_10_1623, i_10_1624, i_10_1711, i_10_1803, i_10_1804, i_10_1954, i_10_1956, i_10_2001, i_10_2002, i_10_2010, i_10_2028, i_10_2091, i_10_2109, i_10_2155, i_10_2162, i_10_2202, i_10_2349, i_10_2356, i_10_2451, i_10_2452, i_10_2515, i_10_2599, i_10_2730, i_10_2731, i_10_2732, i_10_2737, i_10_2742, i_10_2743, i_10_2744, i_10_2832, i_10_2880, i_10_2884, i_10_2955, i_10_2958, i_10_2974, i_10_3048, i_10_3109, i_10_3162, i_10_3272, i_10_3392, i_10_3472, i_10_3492, i_10_3504, i_10_3544, i_10_3546, i_10_3729, i_10_3777, i_10_3840, i_10_3851, i_10_3859, i_10_3860, i_10_3922, i_10_3978, i_10_4126, i_10_4216, i_10_4218, i_10_4269, i_10_4270, i_10_4278, i_10_4287, i_10_4392, i_10_4563, i_10_4571, i_10_4582, i_10_4585, i_10_4588, o_10_362);
	kernel_10_363 k_10_363(i_10_52, i_10_160, i_10_276, i_10_319, i_10_328, i_10_388, i_10_393, i_10_439, i_10_446, i_10_463, i_10_466, i_10_634, i_10_635, i_10_718, i_10_793, i_10_795, i_10_796, i_10_797, i_10_799, i_10_830, i_10_832, i_10_919, i_10_996, i_10_1116, i_10_1209, i_10_1210, i_10_1270, i_10_1295, i_10_1305, i_10_1477, i_10_1492, i_10_1493, i_10_1580, i_10_1655, i_10_1690, i_10_1821, i_10_1822, i_10_1823, i_10_1885, i_10_1889, i_10_1937, i_10_1939, i_10_1940, i_10_1957, i_10_2002, i_10_2004, i_10_2006, i_10_2086, i_10_2245, i_10_2386, i_10_2453, i_10_2455, i_10_2467, i_10_2474, i_10_2516, i_10_2582, i_10_2681, i_10_2701, i_10_2715, i_10_2716, i_10_2740, i_10_2825, i_10_2923, i_10_2983, i_10_2987, i_10_3119, i_10_3122, i_10_3270, i_10_3274, i_10_3387, i_10_3392, i_10_3466, i_10_3467, i_10_3496, i_10_3497, i_10_3538, i_10_3539, i_10_3541, i_10_3586, i_10_3622, i_10_3644, i_10_3645, i_10_3786, i_10_3878, i_10_3879, i_10_3946, i_10_4061, i_10_4116, i_10_4118, i_10_4119, i_10_4120, i_10_4121, i_10_4125, i_10_4155, i_10_4156, i_10_4269, i_10_4270, i_10_4273, i_10_4566, i_10_4569, o_10_363);
	kernel_10_364 k_10_364(i_10_38, i_10_43, i_10_47, i_10_118, i_10_127, i_10_130, i_10_131, i_10_171, i_10_181, i_10_244, i_10_349, i_10_361, i_10_391, i_10_424, i_10_427, i_10_437, i_10_439, i_10_442, i_10_459, i_10_560, i_10_740, i_10_794, i_10_820, i_10_956, i_10_982, i_10_999, i_10_1000, i_10_1084, i_10_1088, i_10_1215, i_10_1234, i_10_1235, i_10_1236, i_10_1237, i_10_1296, i_10_1345, i_10_1378, i_10_1546, i_10_1579, i_10_1693, i_10_1909, i_10_1944, i_10_1947, i_10_2025, i_10_2037, i_10_2089, i_10_2113, i_10_2204, i_10_2270, i_10_2272, i_10_2305, i_10_2341, i_10_2351, i_10_2354, i_10_2361, i_10_2453, i_10_2455, i_10_2459, i_10_2468, i_10_2606, i_10_2631, i_10_2634, i_10_2700, i_10_2703, i_10_2725, i_10_2783, i_10_2863, i_10_2910, i_10_2961, i_10_3036, i_10_3037, i_10_3038, i_10_3042, i_10_3154, i_10_3163, i_10_3232, i_10_3352, i_10_3356, i_10_3466, i_10_3523, i_10_3541, i_10_3553, i_10_3556, i_10_3582, i_10_3584, i_10_3617, i_10_3686, i_10_3838, i_10_3860, i_10_4023, i_10_4053, i_10_4118, i_10_4154, i_10_4169, i_10_4204, i_10_4367, i_10_4394, i_10_4395, i_10_4432, i_10_4593, o_10_364);
	kernel_10_365 k_10_365(i_10_216, i_10_246, i_10_249, i_10_275, i_10_278, i_10_282, i_10_283, i_10_287, i_10_324, i_10_329, i_10_465, i_10_508, i_10_750, i_10_751, i_10_799, i_10_898, i_10_957, i_10_1002, i_10_1029, i_10_1032, i_10_1128, i_10_1138, i_10_1139, i_10_1162, i_10_1239, i_10_1240, i_10_1241, i_10_1242, i_10_1243, i_10_1244, i_10_1245, i_10_1265, i_10_1308, i_10_1345, i_10_1575, i_10_1578, i_10_1579, i_10_1581, i_10_1614, i_10_1647, i_10_1650, i_10_1651, i_10_1655, i_10_1687, i_10_1764, i_10_1819, i_10_1826, i_10_2355, i_10_2449, i_10_2456, i_10_2463, i_10_2604, i_10_2628, i_10_2631, i_10_2632, i_10_2643, i_10_2718, i_10_2724, i_10_2832, i_10_2833, i_10_2916, i_10_2917, i_10_2919, i_10_2922, i_10_2979, i_10_3034, i_10_3037, i_10_3162, i_10_3203, i_10_3277, i_10_3280, i_10_3325, i_10_3386, i_10_3402, i_10_3409, i_10_3588, i_10_3645, i_10_3648, i_10_3653, i_10_3729, i_10_3781, i_10_3783, i_10_3785, i_10_3786, i_10_3841, i_10_3844, i_10_3852, i_10_3855, i_10_4115, i_10_4116, i_10_4117, i_10_4118, i_10_4119, i_10_4120, i_10_4129, i_10_4278, i_10_4290, i_10_4564, i_10_4565, i_10_4566, o_10_365);
	kernel_10_366 k_10_366(i_10_28, i_10_70, i_10_102, i_10_103, i_10_120, i_10_214, i_10_220, i_10_223, i_10_279, i_10_280, i_10_372, i_10_373, i_10_375, i_10_408, i_10_424, i_10_459, i_10_461, i_10_463, i_10_499, i_10_586, i_10_588, i_10_724, i_10_792, i_10_795, i_10_798, i_10_919, i_10_922, i_10_957, i_10_960, i_10_999, i_10_1002, i_10_1039, i_10_1045, i_10_1164, i_10_1201, i_10_1233, i_10_1237, i_10_1240, i_10_1263, i_10_1380, i_10_1429, i_10_1648, i_10_1653, i_10_1785, i_10_1821, i_10_1866, i_10_1940, i_10_2004, i_10_2032, i_10_2094, i_10_2248, i_10_2329, i_10_2337, i_10_2450, i_10_2452, i_10_2470, i_10_2509, i_10_2510, i_10_2673, i_10_2676, i_10_2713, i_10_2782, i_10_2783, i_10_2839, i_10_2865, i_10_2869, i_10_2874, i_10_2881, i_10_2919, i_10_2923, i_10_2992, i_10_3070, i_10_3210, i_10_3238, i_10_3336, i_10_3433, i_10_3450, i_10_3470, i_10_3480, i_10_3496, i_10_3497, i_10_3559, i_10_3562, i_10_3645, i_10_3687, i_10_3837, i_10_3838, i_10_3841, i_10_3874, i_10_4055, i_10_4152, i_10_4234, i_10_4422, i_10_4423, i_10_4426, i_10_4434, i_10_4446, i_10_4447, i_10_4578, i_10_4579, o_10_366);
	kernel_10_367 k_10_367(i_10_150, i_10_181, i_10_201, i_10_291, i_10_427, i_10_434, i_10_463, i_10_465, i_10_496, i_10_507, i_10_558, i_10_589, i_10_604, i_10_607, i_10_792, i_10_819, i_10_839, i_10_903, i_10_928, i_10_945, i_10_981, i_10_1080, i_10_1092, i_10_1120, i_10_1279, i_10_1353, i_10_1397, i_10_1440, i_10_1452, i_10_1548, i_10_1566, i_10_1652, i_10_1796, i_10_1819, i_10_1820, i_10_1825, i_10_1875, i_10_1999, i_10_2016, i_10_2018, i_10_2025, i_10_2107, i_10_2178, i_10_2180, i_10_2334, i_10_2341, i_10_2450, i_10_2502, i_10_2511, i_10_2556, i_10_2595, i_10_2596, i_10_2614, i_10_2629, i_10_2632, i_10_2635, i_10_2638, i_10_2664, i_10_2700, i_10_2707, i_10_2714, i_10_2718, i_10_2821, i_10_2831, i_10_2866, i_10_2881, i_10_2917, i_10_2918, i_10_2944, i_10_2947, i_10_2952, i_10_2953, i_10_3106, i_10_3235, i_10_3238, i_10_3267, i_10_3279, i_10_3465, i_10_3493, i_10_3520, i_10_3540, i_10_3541, i_10_3612, i_10_3619, i_10_3684, i_10_3685, i_10_3838, i_10_3855, i_10_3856, i_10_3883, i_10_3943, i_10_3988, i_10_3993, i_10_4113, i_10_4122, i_10_4194, i_10_4213, i_10_4268, i_10_4393, i_10_4594, o_10_367);
	kernel_10_368 k_10_368(i_10_29, i_10_253, i_10_270, i_10_271, i_10_284, i_10_287, i_10_390, i_10_391, i_10_392, i_10_495, i_10_558, i_10_694, i_10_963, i_10_1002, i_10_1029, i_10_1045, i_10_1107, i_10_1108, i_10_1206, i_10_1235, i_10_1238, i_10_1243, i_10_1244, i_10_1296, i_10_1297, i_10_1310, i_10_1528, i_10_1550, i_10_1575, i_10_1576, i_10_1621, i_10_1630, i_10_1683, i_10_1685, i_10_1686, i_10_1687, i_10_1688, i_10_1735, i_10_1794, i_10_1798, i_10_1800, i_10_1801, i_10_1820, i_10_1911, i_10_1912, i_10_1981, i_10_1999, i_10_2107, i_10_2349, i_10_2351, i_10_2380, i_10_2439, i_10_2440, i_10_2443, i_10_2467, i_10_2542, i_10_2548, i_10_2556, i_10_2566, i_10_2621, i_10_2701, i_10_2702, i_10_2719, i_10_2720, i_10_2730, i_10_2755, i_10_2817, i_10_2882, i_10_2969, i_10_3070, i_10_3171, i_10_3278, i_10_3321, i_10_3323, i_10_3355, i_10_3386, i_10_3407, i_10_3463, i_10_3525, i_10_3555, i_10_3574, i_10_3583, i_10_3647, i_10_3703, i_10_3704, i_10_3707, i_10_3783, i_10_3785, i_10_3817, i_10_3857, i_10_3871, i_10_3909, i_10_3910, i_10_4140, i_10_4177, i_10_4270, i_10_4284, i_10_4307, i_10_4431, i_10_4582, o_10_368);
	kernel_10_369 k_10_369(i_10_263, i_10_271, i_10_286, i_10_326, i_10_412, i_10_424, i_10_425, i_10_427, i_10_464, i_10_640, i_10_712, i_10_1082, i_10_1084, i_10_1136, i_10_1238, i_10_1241, i_10_1305, i_10_1306, i_10_1309, i_10_1310, i_10_1313, i_10_1445, i_10_1543, i_10_1549, i_10_1550, i_10_1603, i_10_1648, i_10_1650, i_10_1651, i_10_1654, i_10_1685, i_10_1687, i_10_1690, i_10_1818, i_10_1819, i_10_1825, i_10_1994, i_10_2306, i_10_2349, i_10_2350, i_10_2362, i_10_2363, i_10_2377, i_10_2407, i_10_2448, i_10_2629, i_10_2630, i_10_2705, i_10_2710, i_10_2711, i_10_2827, i_10_2828, i_10_2832, i_10_2884, i_10_2888, i_10_2919, i_10_2920, i_10_2921, i_10_2922, i_10_2980, i_10_3033, i_10_3092, i_10_3152, i_10_3277, i_10_3386, i_10_3388, i_10_3403, i_10_3404, i_10_3523, i_10_3547, i_10_3613, i_10_3617, i_10_3646, i_10_3649, i_10_3787, i_10_3834, i_10_3841, i_10_3847, i_10_3851, i_10_3852, i_10_3853, i_10_3854, i_10_3857, i_10_3890, i_10_3982, i_10_3990, i_10_4121, i_10_4122, i_10_4123, i_10_4189, i_10_4231, i_10_4270, i_10_4271, i_10_4285, i_10_4286, i_10_4287, i_10_4288, i_10_4567, i_10_4568, i_10_4592, o_10_369);
	kernel_10_370 k_10_370(i_10_39, i_10_48, i_10_171, i_10_174, i_10_175, i_10_193, i_10_247, i_10_249, i_10_289, i_10_318, i_10_327, i_10_330, i_10_364, i_10_405, i_10_406, i_10_412, i_10_435, i_10_520, i_10_594, i_10_633, i_10_793, i_10_832, i_10_877, i_10_1002, i_10_1155, i_10_1266, i_10_1270, i_10_1293, i_10_1306, i_10_1327, i_10_1329, i_10_1341, i_10_1344, i_10_1365, i_10_1366, i_10_1441, i_10_1576, i_10_1714, i_10_1825, i_10_1873, i_10_1878, i_10_1992, i_10_1996, i_10_2016, i_10_2020, i_10_2202, i_10_2241, i_10_2250, i_10_2317, i_10_2326, i_10_2352, i_10_2359, i_10_2364, i_10_2380, i_10_2406, i_10_2449, i_10_2473, i_10_2586, i_10_2604, i_10_2605, i_10_2608, i_10_2643, i_10_2676, i_10_2701, i_10_2704, i_10_2720, i_10_2721, i_10_2724, i_10_2782, i_10_2785, i_10_2786, i_10_2834, i_10_2881, i_10_2882, i_10_2994, i_10_3030, i_10_3075, i_10_3165, i_10_3198, i_10_3199, i_10_3273, i_10_3297, i_10_3300, i_10_3588, i_10_3589, i_10_3703, i_10_3714, i_10_3975, i_10_4126, i_10_4156, i_10_4233, i_10_4260, i_10_4273, i_10_4276, i_10_4378, i_10_4505, i_10_4522, i_10_4524, i_10_4581, i_10_4585, o_10_370);
	kernel_10_371 k_10_371(i_10_156, i_10_220, i_10_249, i_10_279, i_10_390, i_10_391, i_10_423, i_10_441, i_10_447, i_10_459, i_10_513, i_10_516, i_10_519, i_10_600, i_10_636, i_10_637, i_10_718, i_10_795, i_10_796, i_10_898, i_10_1087, i_10_1122, i_10_1248, i_10_1306, i_10_1307, i_10_1308, i_10_1339, i_10_1359, i_10_1377, i_10_1485, i_10_1486, i_10_1541, i_10_1642, i_10_1683, i_10_1684, i_10_1685, i_10_1824, i_10_1915, i_10_1950, i_10_2061, i_10_2185, i_10_2247, i_10_2384, i_10_2391, i_10_2451, i_10_2452, i_10_2468, i_10_2562, i_10_2634, i_10_2679, i_10_2715, i_10_2718, i_10_2719, i_10_2721, i_10_2727, i_10_2742, i_10_2743, i_10_2781, i_10_2785, i_10_2786, i_10_2832, i_10_2833, i_10_2916, i_10_2919, i_10_2982, i_10_3047, i_10_3201, i_10_3234, i_10_3237, i_10_3276, i_10_3279, i_10_3312, i_10_3390, i_10_3468, i_10_3471, i_10_3472, i_10_3495, i_10_3519, i_10_3522, i_10_3525, i_10_3586, i_10_3589, i_10_3590, i_10_3834, i_10_3841, i_10_3844, i_10_3853, i_10_3858, i_10_3877, i_10_3906, i_10_3949, i_10_3985, i_10_4114, i_10_4228, i_10_4229, i_10_4271, i_10_4287, i_10_4317, i_10_4318, i_10_4588, o_10_371);
	kernel_10_372 k_10_372(i_10_40, i_10_43, i_10_176, i_10_257, i_10_266, i_10_269, i_10_323, i_10_374, i_10_394, i_10_395, i_10_410, i_10_413, i_10_439, i_10_440, i_10_449, i_10_640, i_10_743, i_10_797, i_10_1004, i_10_1007, i_10_1034, i_10_1042, i_10_1222, i_10_1223, i_10_1235, i_10_1237, i_10_1238, i_10_1240, i_10_1303, i_10_1308, i_10_1310, i_10_1366, i_10_1385, i_10_1435, i_10_1436, i_10_1439, i_10_1544, i_10_1552, i_10_1612, i_10_1717, i_10_1736, i_10_1823, i_10_1916, i_10_1919, i_10_1956, i_10_1988, i_10_2006, i_10_2023, i_10_2029, i_10_2033, i_10_2204, i_10_2312, i_10_2348, i_10_2354, i_10_2608, i_10_2633, i_10_2635, i_10_2636, i_10_2735, i_10_2761, i_10_2786, i_10_2789, i_10_2830, i_10_2843, i_10_2870, i_10_2966, i_10_3024, i_10_3040, i_10_3049, i_10_3050, i_10_3074, i_10_3077, i_10_3391, i_10_3392, i_10_3473, i_10_3506, i_10_3563, i_10_3584, i_10_3586, i_10_3587, i_10_3589, i_10_3590, i_10_3612, i_10_3721, i_10_3722, i_10_3734, i_10_3854, i_10_3860, i_10_3986, i_10_4004, i_10_4161, i_10_4175, i_10_4210, i_10_4211, i_10_4217, i_10_4268, i_10_4271, i_10_4273, i_10_4489, i_10_4535, o_10_372);
	kernel_10_373 k_10_373(i_10_150, i_10_176, i_10_390, i_10_394, i_10_395, i_10_409, i_10_412, i_10_429, i_10_430, i_10_431, i_10_445, i_10_448, i_10_457, i_10_460, i_10_505, i_10_508, i_10_717, i_10_796, i_10_799, i_10_907, i_10_908, i_10_957, i_10_966, i_10_967, i_10_1005, i_10_1307, i_10_1312, i_10_1313, i_10_1583, i_10_1652, i_10_1653, i_10_1655, i_10_1689, i_10_1690, i_10_1823, i_10_1826, i_10_1995, i_10_2033, i_10_2351, i_10_2365, i_10_2407, i_10_2451, i_10_2452, i_10_2453, i_10_2455, i_10_2469, i_10_2472, i_10_2473, i_10_2636, i_10_2659, i_10_2660, i_10_2703, i_10_2704, i_10_2706, i_10_2707, i_10_2708, i_10_2786, i_10_2788, i_10_2789, i_10_2824, i_10_2830, i_10_2833, i_10_2922, i_10_2923, i_10_3071, i_10_3157, i_10_3158, i_10_3196, i_10_3197, i_10_3272, i_10_3283, i_10_3284, i_10_3315, i_10_3328, i_10_3329, i_10_3388, i_10_3391, i_10_3392, i_10_3468, i_10_3469, i_10_3470, i_10_3542, i_10_3544, i_10_3545, i_10_3589, i_10_3613, i_10_3787, i_10_3837, i_10_3840, i_10_3846, i_10_3847, i_10_3859, i_10_3860, i_10_4057, i_10_4121, i_10_4129, i_10_4270, i_10_4274, i_10_4287, i_10_4292, o_10_373);
	kernel_10_374 k_10_374(i_10_117, i_10_171, i_10_173, i_10_222, i_10_249, i_10_250, i_10_282, i_10_283, i_10_295, i_10_316, i_10_423, i_10_425, i_10_431, i_10_433, i_10_449, i_10_467, i_10_748, i_10_795, i_10_799, i_10_892, i_10_893, i_10_957, i_10_958, i_10_959, i_10_960, i_10_1239, i_10_1309, i_10_1360, i_10_1578, i_10_1619, i_10_1648, i_10_1650, i_10_1652, i_10_1822, i_10_1913, i_10_1944, i_10_2178, i_10_2358, i_10_2361, i_10_2382, i_10_2409, i_10_2452, i_10_2454, i_10_2456, i_10_2632, i_10_2658, i_10_2661, i_10_2663, i_10_2702, i_10_2721, i_10_2725, i_10_2729, i_10_2731, i_10_2732, i_10_2734, i_10_2827, i_10_2884, i_10_3033, i_10_3036, i_10_3037, i_10_3042, i_10_3075, i_10_3085, i_10_3087, i_10_3150, i_10_3152, i_10_3154, i_10_3195, i_10_3196, i_10_3276, i_10_3279, i_10_3388, i_10_3583, i_10_3589, i_10_3612, i_10_3617, i_10_3645, i_10_3646, i_10_3647, i_10_3653, i_10_3783, i_10_3785, i_10_3835, i_10_3837, i_10_3838, i_10_3839, i_10_3848, i_10_3854, i_10_3855, i_10_3856, i_10_3857, i_10_3889, i_10_4024, i_10_4051, i_10_4120, i_10_4168, i_10_4212, i_10_4288, i_10_4291, i_10_4566, o_10_374);
	kernel_10_375 k_10_375(i_10_189, i_10_220, i_10_283, i_10_284, i_10_318, i_10_361, i_10_364, i_10_390, i_10_433, i_10_444, i_10_467, i_10_505, i_10_639, i_10_739, i_10_750, i_10_945, i_10_946, i_10_948, i_10_949, i_10_1000, i_10_1002, i_10_1027, i_10_1028, i_10_1030, i_10_1056, i_10_1152, i_10_1153, i_10_1236, i_10_1237, i_10_1238, i_10_1244, i_10_1270, i_10_1311, i_10_1312, i_10_1315, i_10_1360, i_10_1362, i_10_1395, i_10_1440, i_10_1620, i_10_1650, i_10_1651, i_10_1713, i_10_1737, i_10_1740, i_10_1981, i_10_1990, i_10_2019, i_10_2028, i_10_2152, i_10_2153, i_10_2233, i_10_2359, i_10_2364, i_10_2430, i_10_2456, i_10_2473, i_10_2556, i_10_2567, i_10_2632, i_10_2754, i_10_2784, i_10_2817, i_10_2844, i_10_2863, i_10_2961, i_10_3070, i_10_3071, i_10_3087, i_10_3088, i_10_3127, i_10_3196, i_10_3312, i_10_3313, i_10_3472, i_10_3541, i_10_3583, i_10_3653, i_10_3682, i_10_3683, i_10_3700, i_10_3784, i_10_3838, i_10_3846, i_10_3889, i_10_3979, i_10_3991, i_10_4123, i_10_4126, i_10_4169, i_10_4214, i_10_4230, i_10_4258, i_10_4269, i_10_4292, i_10_4350, i_10_4370, i_10_4375, i_10_4437, i_10_4456, o_10_375);
	kernel_10_376 k_10_376(i_10_178, i_10_184, i_10_220, i_10_221, i_10_282, i_10_283, i_10_284, i_10_287, i_10_317, i_10_319, i_10_393, i_10_430, i_10_441, i_10_445, i_10_463, i_10_466, i_10_504, i_10_511, i_10_512, i_10_520, i_10_755, i_10_797, i_10_964, i_10_1033, i_10_1124, i_10_1136, i_10_1138, i_10_1236, i_10_1237, i_10_1249, i_10_1260, i_10_1365, i_10_1366, i_10_1555, i_10_1556, i_10_1575, i_10_1684, i_10_1689, i_10_1821, i_10_1824, i_10_1825, i_10_1826, i_10_1912, i_10_1914, i_10_1915, i_10_2017, i_10_2357, i_10_2451, i_10_2454, i_10_2455, i_10_2456, i_10_2466, i_10_2467, i_10_2635, i_10_2658, i_10_2659, i_10_2660, i_10_2680, i_10_2701, i_10_2721, i_10_2723, i_10_2731, i_10_2787, i_10_2818, i_10_2824, i_10_2826, i_10_2827, i_10_2830, i_10_2883, i_10_2884, i_10_2885, i_10_2982, i_10_3035, i_10_3039, i_10_3041, i_10_3069, i_10_3150, i_10_3151, i_10_3158, i_10_3267, i_10_3271, i_10_3328, i_10_3391, i_10_3409, i_10_3586, i_10_3587, i_10_3612, i_10_3613, i_10_3615, i_10_3783, i_10_3847, i_10_3850, i_10_3855, i_10_3856, i_10_3858, i_10_3982, i_10_4117, i_10_4118, i_10_4119, i_10_4270, o_10_376);
	kernel_10_377 k_10_377(i_10_180, i_10_222, i_10_276, i_10_283, i_10_284, i_10_324, i_10_325, i_10_388, i_10_426, i_10_435, i_10_436, i_10_442, i_10_443, i_10_459, i_10_465, i_10_466, i_10_514, i_10_958, i_10_959, i_10_960, i_10_961, i_10_962, i_10_1163, i_10_1164, i_10_1233, i_10_1236, i_10_1245, i_10_1248, i_10_1432, i_10_1546, i_10_1582, i_10_1652, i_10_1690, i_10_1720, i_10_1759, i_10_1760, i_10_1820, i_10_1822, i_10_1823, i_10_1824, i_10_1826, i_10_2029, i_10_2352, i_10_2380, i_10_2452, i_10_2453, i_10_2630, i_10_2658, i_10_2659, i_10_2660, i_10_2702, i_10_2708, i_10_2713, i_10_2721, i_10_2722, i_10_2724, i_10_2727, i_10_2728, i_10_2730, i_10_2731, i_10_2735, i_10_2982, i_10_3033, i_10_3034, i_10_3035, i_10_3036, i_10_3037, i_10_3069, i_10_3150, i_10_3231, i_10_3268, i_10_3271, i_10_3316, i_10_3332, i_10_3388, i_10_3389, i_10_3391, i_10_3469, i_10_3494, i_10_3537, i_10_3616, i_10_3649, i_10_3783, i_10_3837, i_10_3847, i_10_3848, i_10_3849, i_10_3850, i_10_3857, i_10_3983, i_10_4113, i_10_4120, i_10_4121, i_10_4185, i_10_4269, i_10_4279, i_10_4285, i_10_4286, i_10_4289, i_10_4563, o_10_377);
	kernel_10_378 k_10_378(i_10_145, i_10_171, i_10_173, i_10_223, i_10_247, i_10_261, i_10_262, i_10_263, i_10_270, i_10_273, i_10_282, i_10_315, i_10_316, i_10_317, i_10_319, i_10_320, i_10_388, i_10_389, i_10_391, i_10_392, i_10_406, i_10_407, i_10_428, i_10_433, i_10_434, i_10_437, i_10_442, i_10_445, i_10_623, i_10_792, i_10_892, i_10_994, i_10_1000, i_10_1001, i_10_1081, i_10_1082, i_10_1100, i_10_1103, i_10_1138, i_10_1217, i_10_1219, i_10_1233, i_10_1296, i_10_1299, i_10_1307, i_10_1343, i_10_1433, i_10_1544, i_10_1553, i_10_1580, i_10_1650, i_10_1652, i_10_1655, i_10_1765, i_10_1823, i_10_1825, i_10_1826, i_10_1910, i_10_2000, i_10_2198, i_10_2200, i_10_2362, i_10_2448, i_10_2518, i_10_2602, i_10_2657, i_10_2660, i_10_2721, i_10_2781, i_10_2830, i_10_2832, i_10_2918, i_10_3038, i_10_3072, i_10_3151, i_10_3196, i_10_3197, i_10_3200, i_10_3202, i_10_3203, i_10_3323, i_10_3405, i_10_3431, i_10_3470, i_10_3538, i_10_3539, i_10_3610, i_10_3647, i_10_3793, i_10_3834, i_10_3836, i_10_3838, i_10_3844, i_10_3880, i_10_3979, i_10_3980, i_10_4117, i_10_4169, i_10_4277, i_10_4283, o_10_378);
	kernel_10_379 k_10_379(i_10_31, i_10_247, i_10_346, i_10_391, i_10_394, i_10_435, i_10_438, i_10_443, i_10_518, i_10_560, i_10_563, i_10_597, i_10_623, i_10_714, i_10_798, i_10_968, i_10_1010, i_10_1051, i_10_1236, i_10_1238, i_10_1240, i_10_1241, i_10_1269, i_10_1310, i_10_1359, i_10_1362, i_10_1364, i_10_1498, i_10_1543, i_10_1550, i_10_1632, i_10_1652, i_10_1684, i_10_1807, i_10_1822, i_10_1874, i_10_2021, i_10_2329, i_10_2354, i_10_2454, i_10_2468, i_10_2507, i_10_2513, i_10_2531, i_10_2566, i_10_2569, i_10_2612, i_10_2621, i_10_2635, i_10_2659, i_10_2660, i_10_2674, i_10_2707, i_10_2718, i_10_2719, i_10_2720, i_10_2722, i_10_2729, i_10_2821, i_10_2827, i_10_2830, i_10_2918, i_10_2919, i_10_2920, i_10_2921, i_10_3034, i_10_3072, i_10_3233, i_10_3285, i_10_3286, i_10_3355, i_10_3402, i_10_3434, i_10_3436, i_10_3437, i_10_3493, i_10_3505, i_10_3544, i_10_3613, i_10_3625, i_10_3653, i_10_3683, i_10_3688, i_10_3728, i_10_3827, i_10_3837, i_10_3846, i_10_3857, i_10_3890, i_10_4025, i_10_4122, i_10_4123, i_10_4124, i_10_4279, i_10_4288, i_10_4289, i_10_4307, i_10_4564, i_10_4582, i_10_4590, o_10_379);
	kernel_10_380 k_10_380(i_10_174, i_10_175, i_10_178, i_10_264, i_10_265, i_10_268, i_10_284, i_10_289, i_10_315, i_10_316, i_10_324, i_10_446, i_10_464, i_10_503, i_10_629, i_10_718, i_10_748, i_10_754, i_10_931, i_10_997, i_10_1121, i_10_1221, i_10_1237, i_10_1239, i_10_1361, i_10_1432, i_10_1435, i_10_1438, i_10_1539, i_10_1581, i_10_1627, i_10_1650, i_10_1651, i_10_1652, i_10_1683, i_10_1686, i_10_1687, i_10_1689, i_10_1713, i_10_1717, i_10_1769, i_10_1819, i_10_1821, i_10_1823, i_10_1948, i_10_2032, i_10_2346, i_10_2347, i_10_2352, i_10_2362, i_10_2363, i_10_2451, i_10_2452, i_10_2471, i_10_2631, i_10_2632, i_10_2659, i_10_2709, i_10_2710, i_10_2727, i_10_2734, i_10_2735, i_10_2823, i_10_2850, i_10_2888, i_10_2919, i_10_2965, i_10_2967, i_10_2968, i_10_2980, i_10_3043, i_10_3049, i_10_3070, i_10_3199, i_10_3281, i_10_3283, i_10_3284, i_10_3380, i_10_3392, i_10_3504, i_10_3612, i_10_3781, i_10_3784, i_10_3840, i_10_3985, i_10_3993, i_10_4026, i_10_4113, i_10_4115, i_10_4119, i_10_4149, i_10_4173, i_10_4174, i_10_4212, i_10_4219, i_10_4269, i_10_4272, i_10_4276, i_10_4288, i_10_4571, o_10_380);
	kernel_10_381 k_10_381(i_10_176, i_10_178, i_10_185, i_10_187, i_10_188, i_10_213, i_10_390, i_10_408, i_10_410, i_10_430, i_10_431, i_10_508, i_10_511, i_10_512, i_10_795, i_10_796, i_10_957, i_10_997, i_10_1028, i_10_1032, i_10_1042, i_10_1043, i_10_1141, i_10_1142, i_10_1237, i_10_1238, i_10_1261, i_10_1305, i_10_1308, i_10_1310, i_10_1365, i_10_1366, i_10_1367, i_10_1487, i_10_1580, i_10_1582, i_10_1583, i_10_1653, i_10_1683, i_10_1823, i_10_1824, i_10_1825, i_10_1913, i_10_2021, i_10_2185, i_10_2186, i_10_2309, i_10_2355, i_10_2453, i_10_2703, i_10_2705, i_10_2706, i_10_2707, i_10_2708, i_10_2716, i_10_2717, i_10_2730, i_10_2732, i_10_2734, i_10_2830, i_10_2831, i_10_2833, i_10_2870, i_10_2919, i_10_3037, i_10_3041, i_10_3151, i_10_3152, i_10_3199, i_10_3200, i_10_3270, i_10_3271, i_10_3284, i_10_3387, i_10_3388, i_10_3389, i_10_3390, i_10_3406, i_10_3523, i_10_3611, i_10_3614, i_10_3617, i_10_3651, i_10_3788, i_10_3895, i_10_3896, i_10_3991, i_10_4031, i_10_4119, i_10_4171, i_10_4172, i_10_4175, i_10_4182, i_10_4183, i_10_4192, i_10_4272, i_10_4273, i_10_4280, i_10_4282, i_10_4283, o_10_381);
	kernel_10_382 k_10_382(i_10_15, i_10_48, i_10_219, i_10_222, i_10_264, i_10_285, i_10_286, i_10_316, i_10_321, i_10_374, i_10_387, i_10_390, i_10_408, i_10_623, i_10_626, i_10_750, i_10_800, i_10_961, i_10_1049, i_10_1233, i_10_1234, i_10_1240, i_10_1296, i_10_1312, i_10_1346, i_10_1544, i_10_1549, i_10_1550, i_10_1686, i_10_1731, i_10_1732, i_10_1764, i_10_1810, i_10_1980, i_10_1990, i_10_2028, i_10_2031, i_10_2198, i_10_2199, i_10_2201, i_10_2349, i_10_2350, i_10_2352, i_10_2353, i_10_2364, i_10_2448, i_10_2458, i_10_2466, i_10_2469, i_10_2470, i_10_2472, i_10_2514, i_10_2565, i_10_2568, i_10_2570, i_10_2571, i_10_2628, i_10_2730, i_10_2781, i_10_2819, i_10_2822, i_10_2839, i_10_2880, i_10_2881, i_10_2982, i_10_3039, i_10_3087, i_10_3277, i_10_3283, i_10_3315, i_10_3318, i_10_3353, i_10_3392, i_10_3465, i_10_3468, i_10_3471, i_10_3507, i_10_3519, i_10_3543, i_10_3555, i_10_3582, i_10_3583, i_10_3585, i_10_3616, i_10_3838, i_10_3840, i_10_3980, i_10_4113, i_10_4115, i_10_4123, i_10_4168, i_10_4170, i_10_4266, i_10_4276, i_10_4285, i_10_4289, i_10_4290, i_10_4374, i_10_4461, i_10_4585, o_10_382);
	kernel_10_383 k_10_383(i_10_9, i_10_16, i_10_66, i_10_67, i_10_69, i_10_148, i_10_159, i_10_160, i_10_224, i_10_237, i_10_245, i_10_251, i_10_253, i_10_256, i_10_261, i_10_270, i_10_290, i_10_293, i_10_318, i_10_321, i_10_331, i_10_368, i_10_373, i_10_393, i_10_519, i_10_541, i_10_627, i_10_688, i_10_721, i_10_823, i_10_1029, i_10_1030, i_10_1042, i_10_1110, i_10_1221, i_10_1239, i_10_1296, i_10_1299, i_10_1306, i_10_1359, i_10_1362, i_10_1431, i_10_1435, i_10_1438, i_10_1445, i_10_1513, i_10_1540, i_10_1553, i_10_1612, i_10_1798, i_10_1876, i_10_1879, i_10_1956, i_10_1966, i_10_2019, i_10_2022, i_10_2023, i_10_2196, i_10_2202, i_10_2203, i_10_2207, i_10_2326, i_10_2533, i_10_2535, i_10_2554, i_10_2565, i_10_2569, i_10_2587, i_10_2676, i_10_2709, i_10_2713, i_10_2724, i_10_2806, i_10_2913, i_10_2914, i_10_2989, i_10_2992, i_10_3072, i_10_3073, i_10_3177, i_10_3201, i_10_3268, i_10_3297, i_10_3469, i_10_3470, i_10_3472, i_10_3473, i_10_3504, i_10_3615, i_10_3777, i_10_3793, i_10_3814, i_10_3815, i_10_3840, i_10_3850, i_10_4120, i_10_4171, i_10_4174, i_10_4400, i_10_4587, o_10_383);
	kernel_10_384 k_10_384(i_10_118, i_10_124, i_10_247, i_10_280, i_10_321, i_10_322, i_10_323, i_10_388, i_10_389, i_10_424, i_10_433, i_10_436, i_10_445, i_10_446, i_10_506, i_10_507, i_10_508, i_10_509, i_10_565, i_10_713, i_10_755, i_10_797, i_10_893, i_10_954, i_10_990, i_10_1027, i_10_1031, i_10_1043, i_10_1237, i_10_1309, i_10_1310, i_10_1575, i_10_1647, i_10_1648, i_10_1650, i_10_1691, i_10_1818, i_10_1819, i_10_1821, i_10_1822, i_10_2002, i_10_2197, i_10_2199, i_10_2357, i_10_2361, i_10_2410, i_10_2451, i_10_2452, i_10_2453, i_10_2467, i_10_2468, i_10_2700, i_10_2701, i_10_2702, i_10_2707, i_10_2709, i_10_2716, i_10_2817, i_10_2818, i_10_2826, i_10_2830, i_10_2883, i_10_2884, i_10_3037, i_10_3069, i_10_3088, i_10_3152, i_10_3278, i_10_3280, i_10_3281, i_10_3385, i_10_3386, i_10_3389, i_10_3390, i_10_3403, i_10_3404, i_10_3409, i_10_3583, i_10_3613, i_10_3614, i_10_3648, i_10_3650, i_10_3682, i_10_3835, i_10_3839, i_10_3847, i_10_3848, i_10_3851, i_10_3856, i_10_3860, i_10_3983, i_10_3992, i_10_4126, i_10_4127, i_10_4277, i_10_4292, i_10_4564, i_10_4565, i_10_4567, i_10_4568, o_10_384);
	kernel_10_385 k_10_385(i_10_125, i_10_132, i_10_174, i_10_178, i_10_250, i_10_251, i_10_268, i_10_282, i_10_318, i_10_391, i_10_393, i_10_394, i_10_395, i_10_409, i_10_436, i_10_441, i_10_442, i_10_448, i_10_561, i_10_564, i_10_733, i_10_734, i_10_736, i_10_795, i_10_798, i_10_800, i_10_825, i_10_967, i_10_970, i_10_1002, i_10_1005, i_10_1006, i_10_1033, i_10_1113, i_10_1164, i_10_1233, i_10_1247, i_10_1306, i_10_1500, i_10_1689, i_10_1767, i_10_1821, i_10_1822, i_10_1920, i_10_2004, i_10_2351, i_10_2354, i_10_2361, i_10_2362, i_10_2381, i_10_2407, i_10_2448, i_10_2449, i_10_2453, i_10_2455, i_10_2518, i_10_2562, i_10_2630, i_10_2636, i_10_2662, i_10_2711, i_10_2725, i_10_2730, i_10_2732, i_10_2734, i_10_2833, i_10_2888, i_10_2955, i_10_2983, i_10_3042, i_10_3043, i_10_3049, i_10_3074, i_10_3283, i_10_3390, i_10_3437, i_10_3471, i_10_3472, i_10_3541, i_10_3542, i_10_3586, i_10_3588, i_10_3589, i_10_3612, i_10_3814, i_10_3850, i_10_3930, i_10_3985, i_10_3990, i_10_4024, i_10_4056, i_10_4057, i_10_4116, i_10_4117, i_10_4272, i_10_4292, i_10_4374, i_10_4570, i_10_4597, i_10_4598, o_10_385);
	kernel_10_386 k_10_386(i_10_172, i_10_183, i_10_265, i_10_275, i_10_327, i_10_328, i_10_390, i_10_393, i_10_394, i_10_408, i_10_427, i_10_429, i_10_437, i_10_440, i_10_538, i_10_539, i_10_701, i_10_735, i_10_755, i_10_996, i_10_997, i_10_1002, i_10_1003, i_10_1087, i_10_1138, i_10_1141, i_10_1168, i_10_1233, i_10_1264, i_10_1348, i_10_1349, i_10_1434, i_10_1435, i_10_1445, i_10_1555, i_10_1652, i_10_1655, i_10_1717, i_10_1769, i_10_1772, i_10_1818, i_10_1822, i_10_1823, i_10_1912, i_10_1913, i_10_1948, i_10_1949, i_10_2181, i_10_2184, i_10_2185, i_10_2199, i_10_2204, i_10_2311, i_10_2312, i_10_2329, i_10_2406, i_10_2407, i_10_2408, i_10_2455, i_10_2469, i_10_2481, i_10_2629, i_10_2631, i_10_2657, i_10_2679, i_10_2713, i_10_2716, i_10_2833, i_10_2919, i_10_2921, i_10_2922, i_10_2923, i_10_2982, i_10_2983, i_10_3041, i_10_3047, i_10_3093, i_10_3094, i_10_3152, i_10_3154, i_10_3155, i_10_3210, i_10_3472, i_10_3473, i_10_3497, i_10_3543, i_10_3544, i_10_3588, i_10_3855, i_10_3856, i_10_3859, i_10_4057, i_10_4114, i_10_4117, i_10_4175, i_10_4236, i_10_4238, i_10_4290, i_10_4291, i_10_4533, o_10_386);
	kernel_10_387 k_10_387(i_10_45, i_10_48, i_10_120, i_10_144, i_10_145, i_10_177, i_10_219, i_10_246, i_10_280, i_10_285, i_10_286, i_10_315, i_10_373, i_10_448, i_10_449, i_10_461, i_10_462, i_10_467, i_10_747, i_10_796, i_10_797, i_10_798, i_10_799, i_10_967, i_10_981, i_10_1030, i_10_1242, i_10_1266, i_10_1305, i_10_1309, i_10_1342, i_10_1446, i_10_1482, i_10_1578, i_10_1629, i_10_1632, i_10_1638, i_10_1686, i_10_1689, i_10_1791, i_10_1916, i_10_1925, i_10_1951, i_10_1952, i_10_2025, i_10_2311, i_10_2312, i_10_2349, i_10_2350, i_10_2469, i_10_2565, i_10_2628, i_10_2638, i_10_2658, i_10_2659, i_10_2673, i_10_2700, i_10_2721, i_10_2727, i_10_2728, i_10_2817, i_10_2969, i_10_3043, i_10_3114, i_10_3277, i_10_3283, i_10_3312, i_10_3348, i_10_3360, i_10_3384, i_10_3387, i_10_3388, i_10_3393, i_10_3468, i_10_3471, i_10_3504, i_10_3585, i_10_3619, i_10_3652, i_10_3784, i_10_3843, i_10_3844, i_10_3845, i_10_3847, i_10_3856, i_10_3870, i_10_3913, i_10_4030, i_10_4116, i_10_4117, i_10_4125, i_10_4129, i_10_4152, i_10_4153, i_10_4170, i_10_4267, i_10_4275, i_10_4284, i_10_4290, i_10_4565, o_10_387);
	kernel_10_388 k_10_388(i_10_150, i_10_256, i_10_294, i_10_409, i_10_410, i_10_429, i_10_430, i_10_438, i_10_439, i_10_447, i_10_627, i_10_645, i_10_796, i_10_798, i_10_799, i_10_897, i_10_1033, i_10_1051, i_10_1203, i_10_1245, i_10_1249, i_10_1364, i_10_1367, i_10_1384, i_10_1444, i_10_1552, i_10_1608, i_10_1618, i_10_1650, i_10_1653, i_10_1808, i_10_1822, i_10_1915, i_10_1951, i_10_1995, i_10_1996, i_10_2265, i_10_2338, i_10_2350, i_10_2351, i_10_2352, i_10_2355, i_10_2356, i_10_2364, i_10_2446, i_10_2447, i_10_2451, i_10_2463, i_10_2481, i_10_2482, i_10_2514, i_10_2515, i_10_2543, i_10_2607, i_10_2634, i_10_2643, i_10_2644, i_10_2716, i_10_2717, i_10_2718, i_10_2720, i_10_2726, i_10_2731, i_10_2735, i_10_2866, i_10_2919, i_10_2920, i_10_2922, i_10_3165, i_10_3166, i_10_3175, i_10_3196, i_10_3228, i_10_3270, i_10_3276, i_10_3280, i_10_3281, i_10_3283, i_10_3544, i_10_3561, i_10_3610, i_10_3612, i_10_3613, i_10_3706, i_10_3785, i_10_3838, i_10_3855, i_10_3904, i_10_3991, i_10_3992, i_10_4026, i_10_4027, i_10_4028, i_10_4029, i_10_4215, i_10_4219, i_10_4236, i_10_4276, i_10_4291, i_10_4480, o_10_388);
	kernel_10_389 k_10_389(i_10_35, i_10_71, i_10_242, i_10_251, i_10_275, i_10_283, i_10_284, i_10_285, i_10_368, i_10_448, i_10_466, i_10_467, i_10_545, i_10_719, i_10_752, i_10_800, i_10_954, i_10_959, i_10_1031, i_10_1032, i_10_1033, i_10_1034, i_10_1244, i_10_1248, i_10_1250, i_10_1345, i_10_1439, i_10_1448, i_10_1619, i_10_1687, i_10_1819, i_10_1822, i_10_1823, i_10_1825, i_10_1958, i_10_1961, i_10_1995, i_10_1996, i_10_2185, i_10_2186, i_10_2311, i_10_2312, i_10_2361, i_10_2363, i_10_2365, i_10_2470, i_10_2573, i_10_2609, i_10_2632, i_10_2658, i_10_2663, i_10_2704, i_10_2705, i_10_2708, i_10_2711, i_10_2714, i_10_2717, i_10_2732, i_10_2735, i_10_2744, i_10_2830, i_10_2831, i_10_3034, i_10_3037, i_10_3038, i_10_3077, i_10_3198, i_10_3199, i_10_3272, i_10_3275, i_10_3384, i_10_3389, i_10_3443, i_10_3446, i_10_3472, i_10_3525, i_10_3584, i_10_3613, i_10_3614, i_10_3784, i_10_3785, i_10_3787, i_10_3788, i_10_3840, i_10_3842, i_10_3848, i_10_3849, i_10_3855, i_10_3949, i_10_3991, i_10_4113, i_10_4114, i_10_4118, i_10_4121, i_10_4127, i_10_4170, i_10_4220, i_10_4280, i_10_4291, i_10_4571, o_10_389);
	kernel_10_390 k_10_390(i_10_47, i_10_49, i_10_50, i_10_137, i_10_171, i_10_172, i_10_178, i_10_216, i_10_221, i_10_245, i_10_248, i_10_287, i_10_515, i_10_544, i_10_545, i_10_662, i_10_689, i_10_716, i_10_748, i_10_749, i_10_796, i_10_954, i_10_964, i_10_965, i_10_983, i_10_1028, i_10_1031, i_10_1181, i_10_1184, i_10_1217, i_10_1242, i_10_1244, i_10_1310, i_10_1355, i_10_1487, i_10_1531, i_10_1532, i_10_1541, i_10_1559, i_10_1580, i_10_1616, i_10_1653, i_10_1685, i_10_2003, i_10_2035, i_10_2081, i_10_2161, i_10_2305, i_10_2306, i_10_2308, i_10_2327, i_10_2330, i_10_2363, i_10_2458, i_10_2459, i_10_2463, i_10_2471, i_10_2473, i_10_2567, i_10_2602, i_10_2603, i_10_2630, i_10_2659, i_10_2660, i_10_2737, i_10_2738, i_10_3074, i_10_3199, i_10_3200, i_10_3233, i_10_3281, i_10_3290, i_10_3388, i_10_3406, i_10_3407, i_10_3445, i_10_3550, i_10_3584, i_10_3587, i_10_3610, i_10_3613, i_10_3614, i_10_3619, i_10_3620, i_10_3647, i_10_3800, i_10_3871, i_10_3908, i_10_3998, i_10_4064, i_10_4115, i_10_4126, i_10_4217, i_10_4220, i_10_4268, i_10_4276, i_10_4285, i_10_4287, i_10_4288, i_10_4289, o_10_390);
	kernel_10_391 k_10_391(i_10_47, i_10_51, i_10_83, i_10_155, i_10_217, i_10_220, i_10_245, i_10_281, i_10_283, i_10_286, i_10_319, i_10_329, i_10_389, i_10_409, i_10_434, i_10_436, i_10_441, i_10_442, i_10_462, i_10_465, i_10_639, i_10_640, i_10_643, i_10_985, i_10_1026, i_10_1029, i_10_1046, i_10_1059, i_10_1207, i_10_1237, i_10_1250, i_10_1264, i_10_1492, i_10_1543, i_10_1683, i_10_1689, i_10_1824, i_10_1825, i_10_1826, i_10_1915, i_10_1992, i_10_1999, i_10_2000, i_10_2016, i_10_2352, i_10_2436, i_10_2448, i_10_2449, i_10_2452, i_10_2464, i_10_2465, i_10_2628, i_10_2631, i_10_2642, i_10_2656, i_10_2659, i_10_2660, i_10_2674, i_10_2727, i_10_2728, i_10_2729, i_10_2819, i_10_2829, i_10_2830, i_10_2833, i_10_2963, i_10_2964, i_10_2982, i_10_2986, i_10_3045, i_10_3087, i_10_3088, i_10_3089, i_10_3094, i_10_3161, i_10_3233, i_10_3289, i_10_3388, i_10_3391, i_10_3434, i_10_3504, i_10_3522, i_10_3523, i_10_3524, i_10_3682, i_10_3700, i_10_3783, i_10_3809, i_10_3838, i_10_3856, i_10_3857, i_10_4029, i_10_4054, i_10_4127, i_10_4153, i_10_4172, i_10_4275, i_10_4280, i_10_4282, i_10_4292, o_10_391);
	kernel_10_392 k_10_392(i_10_281, i_10_282, i_10_295, i_10_296, i_10_327, i_10_328, i_10_329, i_10_407, i_10_433, i_10_434, i_10_441, i_10_442, i_10_443, i_10_444, i_10_445, i_10_749, i_10_796, i_10_960, i_10_1233, i_10_1234, i_10_1235, i_10_1239, i_10_1263, i_10_1311, i_10_1312, i_10_1348, i_10_1431, i_10_1432, i_10_1447, i_10_1654, i_10_1767, i_10_1768, i_10_1819, i_10_1822, i_10_1823, i_10_1824, i_10_1825, i_10_1911, i_10_1912, i_10_1913, i_10_1946, i_10_2180, i_10_2457, i_10_2458, i_10_2470, i_10_2629, i_10_2630, i_10_2656, i_10_2658, i_10_2659, i_10_2663, i_10_2711, i_10_2716, i_10_2718, i_10_2719, i_10_2722, i_10_2723, i_10_2781, i_10_2782, i_10_2783, i_10_2817, i_10_2819, i_10_2826, i_10_2827, i_10_2830, i_10_2831, i_10_2923, i_10_2981, i_10_3033, i_10_3034, i_10_3035, i_10_3047, i_10_3196, i_10_3323, i_10_3392, i_10_3403, i_10_3409, i_10_3523, i_10_3583, i_10_3609, i_10_3612, i_10_3613, i_10_3682, i_10_3783, i_10_3785, i_10_3838, i_10_3839, i_10_3852, i_10_3853, i_10_3857, i_10_3906, i_10_3907, i_10_3991, i_10_4113, i_10_4116, i_10_4118, i_10_4267, i_10_4285, i_10_4288, i_10_4566, o_10_392);
	kernel_10_393 k_10_393(i_10_100, i_10_133, i_10_134, i_10_174, i_10_175, i_10_190, i_10_282, i_10_432, i_10_444, i_10_446, i_10_514, i_10_643, i_10_715, i_10_796, i_10_829, i_10_830, i_10_836, i_10_853, i_10_896, i_10_905, i_10_965, i_10_990, i_10_991, i_10_1051, i_10_1233, i_10_1289, i_10_1305, i_10_1306, i_10_1342, i_10_1366, i_10_1434, i_10_1478, i_10_1558, i_10_1640, i_10_1913, i_10_1949, i_10_1991, i_10_2020, i_10_2349, i_10_2351, i_10_2352, i_10_2353, i_10_2354, i_10_2363, i_10_2365, i_10_2366, i_10_2470, i_10_2515, i_10_2527, i_10_2539, i_10_2629, i_10_2675, i_10_2744, i_10_2817, i_10_2818, i_10_2855, i_10_2881, i_10_2917, i_10_2918, i_10_2921, i_10_2980, i_10_3083, i_10_3107, i_10_3114, i_10_3197, i_10_3269, i_10_3298, i_10_3352, i_10_3391, i_10_3392, i_10_3403, i_10_3443, i_10_3460, i_10_3471, i_10_3497, i_10_3502, i_10_3503, i_10_3539, i_10_3609, i_10_3612, i_10_3615, i_10_3617, i_10_3625, i_10_3626, i_10_3683, i_10_3729, i_10_3730, i_10_3731, i_10_3776, i_10_3833, i_10_3858, i_10_3899, i_10_4118, i_10_4185, i_10_4276, i_10_4277, i_10_4403, i_10_4457, i_10_4573, i_10_4583, o_10_393);
	kernel_10_394 k_10_394(i_10_82, i_10_119, i_10_122, i_10_223, i_10_282, i_10_327, i_10_328, i_10_360, i_10_387, i_10_388, i_10_390, i_10_434, i_10_436, i_10_437, i_10_446, i_10_447, i_10_459, i_10_463, i_10_464, i_10_903, i_10_962, i_10_990, i_10_1000, i_10_1027, i_10_1035, i_10_1036, i_10_1083, i_10_1241, i_10_1261, i_10_1380, i_10_1449, i_10_1450, i_10_1452, i_10_1530, i_10_1551, i_10_1654, i_10_1684, i_10_1685, i_10_1872, i_10_1873, i_10_1875, i_10_1911, i_10_2000, i_10_2181, i_10_2182, i_10_2224, i_10_2352, i_10_2377, i_10_2378, i_10_2403, i_10_2449, i_10_2453, i_10_2455, i_10_2602, i_10_2603, i_10_2628, i_10_2658, i_10_2673, i_10_2700, i_10_2718, i_10_2721, i_10_2731, i_10_2826, i_10_2827, i_10_2828, i_10_2829, i_10_2920, i_10_2923, i_10_3036, i_10_3037, i_10_3041, i_10_3042, i_10_3087, i_10_3159, i_10_3283, i_10_3384, i_10_3389, i_10_3432, i_10_3470, i_10_3522, i_10_3537, i_10_3560, i_10_3563, i_10_3685, i_10_3782, i_10_3784, i_10_3786, i_10_3787, i_10_3834, i_10_3855, i_10_3856, i_10_3892, i_10_3981, i_10_4025, i_10_4113, i_10_4213, i_10_4270, i_10_4279, i_10_4285, i_10_4288, o_10_394);
	kernel_10_395 k_10_395(i_10_41, i_10_42, i_10_147, i_10_175, i_10_179, i_10_224, i_10_251, i_10_255, i_10_272, i_10_282, i_10_318, i_10_327, i_10_328, i_10_439, i_10_444, i_10_445, i_10_447, i_10_516, i_10_517, i_10_717, i_10_755, i_10_798, i_10_956, i_10_958, i_10_959, i_10_961, i_10_968, i_10_984, i_10_1028, i_10_1033, i_10_1034, i_10_1206, i_10_1207, i_10_1306, i_10_1381, i_10_1438, i_10_1443, i_10_1575, i_10_1581, i_10_1582, i_10_1645, i_10_1650, i_10_1653, i_10_1654, i_10_1686, i_10_1713, i_10_1723, i_10_1727, i_10_1890, i_10_2006, i_10_2017, i_10_2018, i_10_2179, i_10_2196, i_10_2197, i_10_2204, i_10_2254, i_10_2327, i_10_2386, i_10_2450, i_10_2452, i_10_2459, i_10_2471, i_10_2542, i_10_2564, i_10_2636, i_10_2700, i_10_2702, i_10_2715, i_10_2721, i_10_2722, i_10_2724, i_10_2743, i_10_2744, i_10_2922, i_10_2980, i_10_3038, i_10_3071, i_10_3072, i_10_3079, i_10_3195, i_10_3196, i_10_3197, i_10_3313, i_10_3388, i_10_3391, i_10_3392, i_10_3402, i_10_3473, i_10_3493, i_10_3614, i_10_3646, i_10_3782, i_10_3798, i_10_3799, i_10_3838, i_10_3982, i_10_4125, i_10_4170, i_10_4531, o_10_395);
	kernel_10_396 k_10_396(i_10_160, i_10_246, i_10_442, i_10_461, i_10_464, i_10_716, i_10_728, i_10_749, i_10_899, i_10_905, i_10_913, i_10_962, i_10_995, i_10_1058, i_10_1087, i_10_1129, i_10_1130, i_10_1220, i_10_1307, i_10_1309, i_10_1310, i_10_1311, i_10_1312, i_10_1391, i_10_1442, i_10_1454, i_10_1567, i_10_1577, i_10_1579, i_10_1814, i_10_1822, i_10_1823, i_10_1930, i_10_2182, i_10_2204, i_10_2305, i_10_2306, i_10_2307, i_10_2433, i_10_2449, i_10_2450, i_10_2451, i_10_2452, i_10_2474, i_10_2475, i_10_2516, i_10_2609, i_10_2705, i_10_2722, i_10_2787, i_10_2822, i_10_2828, i_10_2876, i_10_2886, i_10_2986, i_10_2987, i_10_3071, i_10_3094, i_10_3227, i_10_3361, i_10_3389, i_10_3430, i_10_3451, i_10_3452, i_10_3455, i_10_3589, i_10_3610, i_10_3640, i_10_3650, i_10_3652, i_10_3686, i_10_3703, i_10_3721, i_10_3725, i_10_3837, i_10_3840, i_10_3896, i_10_3920, i_10_3978, i_10_4057, i_10_4113, i_10_4117, i_10_4118, i_10_4130, i_10_4145, i_10_4148, i_10_4173, i_10_4174, i_10_4231, i_10_4238, i_10_4275, i_10_4278, i_10_4279, i_10_4281, i_10_4379, i_10_4397, i_10_4517, i_10_4531, i_10_4535, i_10_4560, o_10_396);
	kernel_10_397 k_10_397(i_10_146, i_10_224, i_10_263, i_10_273, i_10_274, i_10_276, i_10_279, i_10_282, i_10_283, i_10_320, i_10_392, i_10_428, i_10_431, i_10_458, i_10_460, i_10_463, i_10_518, i_10_689, i_10_1235, i_10_1237, i_10_1238, i_10_1241, i_10_1306, i_10_1311, i_10_1312, i_10_1432, i_10_1435, i_10_1439, i_10_1541, i_10_1628, i_10_1634, i_10_1643, i_10_1651, i_10_1652, i_10_1653, i_10_1654, i_10_1733, i_10_1820, i_10_1826, i_10_2000, i_10_2006, i_10_2027, i_10_2031, i_10_2033, i_10_2358, i_10_2361, i_10_2383, i_10_2384, i_10_2468, i_10_2471, i_10_2474, i_10_2628, i_10_2702, i_10_2719, i_10_2721, i_10_2723, i_10_2731, i_10_2782, i_10_2783, i_10_2827, i_10_2828, i_10_2920, i_10_3037, i_10_3043, i_10_3050, i_10_3069, i_10_3116, i_10_3276, i_10_3281, i_10_3314, i_10_3385, i_10_3387, i_10_3402, i_10_3467, i_10_3470, i_10_3473, i_10_3506, i_10_3509, i_10_3545, i_10_3583, i_10_3584, i_10_3587, i_10_3589, i_10_3590, i_10_3650, i_10_3682, i_10_3787, i_10_3788, i_10_3800, i_10_3808, i_10_3809, i_10_3838, i_10_3839, i_10_3842, i_10_3983, i_10_3988, i_10_4271, i_10_4286, i_10_4289, i_10_4571, o_10_397);
	kernel_10_398 k_10_398(i_10_145, i_10_262, i_10_284, i_10_325, i_10_408, i_10_433, i_10_436, i_10_447, i_10_711, i_10_892, i_10_893, i_10_927, i_10_990, i_10_1036, i_10_1039, i_10_1120, i_10_1165, i_10_1166, i_10_1236, i_10_1238, i_10_1247, i_10_1307, i_10_1381, i_10_1440, i_10_1485, i_10_1554, i_10_1603, i_10_1800, i_10_1801, i_10_1824, i_10_1825, i_10_1826, i_10_1908, i_10_1909, i_10_1911, i_10_1981, i_10_1990, i_10_2206, i_10_2223, i_10_2224, i_10_2332, i_10_2449, i_10_2450, i_10_2458, i_10_2481, i_10_2515, i_10_2565, i_10_2567, i_10_2571, i_10_2635, i_10_2686, i_10_2700, i_10_2701, i_10_2728, i_10_2827, i_10_2829, i_10_2831, i_10_2862, i_10_2865, i_10_2866, i_10_2916, i_10_2917, i_10_2919, i_10_2920, i_10_2921, i_10_2922, i_10_2923, i_10_3072, i_10_3199, i_10_3201, i_10_3267, i_10_3278, i_10_3298, i_10_3299, i_10_3384, i_10_3385, i_10_3386, i_10_3388, i_10_3406, i_10_3457, i_10_3523, i_10_3600, i_10_3610, i_10_3611, i_10_3648, i_10_3851, i_10_3855, i_10_3889, i_10_3897, i_10_3942, i_10_3943, i_10_3961, i_10_4120, i_10_4129, i_10_4269, i_10_4270, i_10_4285, i_10_4306, i_10_4500, i_10_4597, o_10_398);
	kernel_10_399 k_10_399(i_10_29, i_10_41, i_10_50, i_10_146, i_10_173, i_10_174, i_10_224, i_10_250, i_10_316, i_10_319, i_10_406, i_10_430, i_10_431, i_10_508, i_10_509, i_10_518, i_10_589, i_10_590, i_10_751, i_10_792, i_10_796, i_10_800, i_10_908, i_10_964, i_10_1032, i_10_1138, i_10_1306, i_10_1448, i_10_1545, i_10_1643, i_10_1690, i_10_1769, i_10_1811, i_10_1913, i_10_1937, i_10_1949, i_10_1999, i_10_2003, i_10_2312, i_10_2350, i_10_2354, i_10_2365, i_10_2389, i_10_2450, i_10_2451, i_10_2452, i_10_2453, i_10_2455, i_10_2469, i_10_2471, i_10_2546, i_10_2628, i_10_2629, i_10_2661, i_10_2663, i_10_2705, i_10_2717, i_10_2722, i_10_2723, i_10_2731, i_10_2732, i_10_2781, i_10_2785, i_10_2821, i_10_2822, i_10_2824, i_10_2827, i_10_2828, i_10_3035, i_10_3157, i_10_3236, i_10_3271, i_10_3280, i_10_3281, i_10_3284, i_10_3322, i_10_3410, i_10_3466, i_10_3494, i_10_3497, i_10_3520, i_10_3526, i_10_3584, i_10_3587, i_10_3613, i_10_3617, i_10_3649, i_10_3788, i_10_3800, i_10_3838, i_10_3846, i_10_3875, i_10_3911, i_10_3914, i_10_4123, i_10_4172, i_10_4268, i_10_4277, i_10_4291, i_10_4292, o_10_399);
	kernel_10_400 k_10_400(i_10_150, i_10_174, i_10_175, i_10_176, i_10_177, i_10_178, i_10_179, i_10_250, i_10_251, i_10_281, i_10_282, i_10_285, i_10_287, i_10_289, i_10_318, i_10_321, i_10_322, i_10_407, i_10_408, i_10_412, i_10_428, i_10_437, i_10_439, i_10_455, i_10_717, i_10_1002, i_10_1003, i_10_1138, i_10_1142, i_10_1236, i_10_1237, i_10_1312, i_10_1344, i_10_1365, i_10_1384, i_10_1441, i_10_1651, i_10_1684, i_10_1688, i_10_1689, i_10_1690, i_10_1821, i_10_1823, i_10_1990, i_10_2022, i_10_2028, i_10_2311, i_10_2349, i_10_2353, i_10_2410, i_10_2411, i_10_2453, i_10_2454, i_10_2629, i_10_2632, i_10_2633, i_10_2635, i_10_2636, i_10_2655, i_10_2660, i_10_2661, i_10_2704, i_10_2714, i_10_2727, i_10_2733, i_10_2734, i_10_2735, i_10_2781, i_10_2785, i_10_2826, i_10_2834, i_10_3039, i_10_3042, i_10_3075, i_10_3157, i_10_3202, i_10_3390, i_10_3405, i_10_3468, i_10_3469, i_10_3496, i_10_3615, i_10_3648, i_10_3651, i_10_3839, i_10_3846, i_10_3857, i_10_3858, i_10_3860, i_10_3912, i_10_3984, i_10_4116, i_10_4117, i_10_4119, i_10_4120, i_10_4122, i_10_4123, i_10_4125, i_10_4126, i_10_4270, o_10_400);
	kernel_10_401 k_10_401(i_10_34, i_10_124, i_10_177, i_10_246, i_10_249, i_10_269, i_10_282, i_10_283, i_10_318, i_10_328, i_10_329, i_10_437, i_10_445, i_10_512, i_10_962, i_10_1006, i_10_1135, i_10_1137, i_10_1138, i_10_1241, i_10_1266, i_10_1348, i_10_1366, i_10_1583, i_10_1617, i_10_1680, i_10_1687, i_10_1819, i_10_1821, i_10_1825, i_10_1876, i_10_1912, i_10_1913, i_10_1951, i_10_1952, i_10_2084, i_10_2184, i_10_2185, i_10_2186, i_10_2203, i_10_2312, i_10_2327, i_10_2329, i_10_2338, i_10_2353, i_10_2354, i_10_2384, i_10_2407, i_10_2408, i_10_2410, i_10_2411, i_10_2452, i_10_2453, i_10_2470, i_10_2632, i_10_2655, i_10_2659, i_10_2660, i_10_2708, i_10_2726, i_10_2731, i_10_2829, i_10_2884, i_10_2885, i_10_2921, i_10_2980, i_10_2981, i_10_2986, i_10_3069, i_10_3274, i_10_3327, i_10_3328, i_10_3384, i_10_3497, i_10_3590, i_10_3616, i_10_3787, i_10_3847, i_10_3848, i_10_3853, i_10_3855, i_10_3859, i_10_3895, i_10_3920, i_10_3993, i_10_4056, i_10_4057, i_10_4058, i_10_4116, i_10_4117, i_10_4118, i_10_4124, i_10_4126, i_10_4127, i_10_4237, i_10_4238, i_10_4289, i_10_4290, i_10_4568, i_10_4570, o_10_401);
	kernel_10_402 k_10_402(i_10_175, i_10_178, i_10_246, i_10_247, i_10_249, i_10_251, i_10_284, i_10_286, i_10_293, i_10_322, i_10_406, i_10_409, i_10_410, i_10_412, i_10_460, i_10_461, i_10_462, i_10_463, i_10_509, i_10_800, i_10_964, i_10_996, i_10_997, i_10_1000, i_10_1236, i_10_1239, i_10_1241, i_10_1246, i_10_1260, i_10_1306, i_10_1313, i_10_1432, i_10_1434, i_10_1687, i_10_1689, i_10_1691, i_10_1823, i_10_2019, i_10_2020, i_10_2022, i_10_2023, i_10_2024, i_10_2032, i_10_2356, i_10_2361, i_10_2405, i_10_2450, i_10_2607, i_10_2608, i_10_2629, i_10_2631, i_10_2632, i_10_2636, i_10_2662, i_10_2677, i_10_2700, i_10_2704, i_10_2707, i_10_2715, i_10_2722, i_10_2726, i_10_2727, i_10_2781, i_10_2782, i_10_2784, i_10_2785, i_10_3203, i_10_3436, i_10_3525, i_10_3526, i_10_3650, i_10_3684, i_10_3784, i_10_3836, i_10_3841, i_10_3850, i_10_3856, i_10_3990, i_10_3991, i_10_3995, i_10_4053, i_10_4117, i_10_4118, i_10_4119, i_10_4120, i_10_4125, i_10_4126, i_10_4129, i_10_4130, i_10_4173, i_10_4174, i_10_4266, i_10_4270, i_10_4272, i_10_4273, i_10_4289, i_10_4290, i_10_4291, i_10_4292, i_10_4571, o_10_402);
	kernel_10_403 k_10_403(i_10_216, i_10_223, i_10_279, i_10_282, i_10_287, i_10_327, i_10_328, i_10_423, i_10_424, i_10_426, i_10_462, i_10_463, i_10_694, i_10_696, i_10_697, i_10_793, i_10_797, i_10_799, i_10_895, i_10_897, i_10_1030, i_10_1032, i_10_1033, i_10_1034, i_10_1035, i_10_1117, i_10_1131, i_10_1234, i_10_1236, i_10_1237, i_10_1346, i_10_1546, i_10_1548, i_10_1619, i_10_1767, i_10_1821, i_10_1908, i_10_1909, i_10_1911, i_10_1995, i_10_2002, i_10_2152, i_10_2309, i_10_2349, i_10_2352, i_10_2353, i_10_2406, i_10_2430, i_10_2456, i_10_2457, i_10_2465, i_10_2470, i_10_2538, i_10_2631, i_10_2634, i_10_2635, i_10_2636, i_10_2709, i_10_2718, i_10_2722, i_10_2826, i_10_2827, i_10_2888, i_10_2916, i_10_2922, i_10_2983, i_10_3089, i_10_3092, i_10_3195, i_10_3196, i_10_3199, i_10_3276, i_10_3277, i_10_3306, i_10_3405, i_10_3406, i_10_3407, i_10_3408, i_10_3409, i_10_3610, i_10_3613, i_10_3650, i_10_3702, i_10_3852, i_10_3853, i_10_3855, i_10_3856, i_10_3889, i_10_3901, i_10_3904, i_10_4126, i_10_4129, i_10_4130, i_10_4206, i_10_4219, i_10_4233, i_10_4290, i_10_4565, i_10_4590, i_10_4591, o_10_403);
	kernel_10_404 k_10_404(i_10_29, i_10_49, i_10_172, i_10_176, i_10_194, i_10_247, i_10_280, i_10_319, i_10_409, i_10_428, i_10_433, i_10_434, i_10_464, i_10_695, i_10_700, i_10_731, i_10_904, i_10_992, i_10_1046, i_10_1048, i_10_1052, i_10_1109, i_10_1199, i_10_1233, i_10_1307, i_10_1309, i_10_1312, i_10_1313, i_10_1345, i_10_1348, i_10_1448, i_10_1550, i_10_1630, i_10_1650, i_10_1684, i_10_1685, i_10_1820, i_10_1821, i_10_1824, i_10_1825, i_10_1908, i_10_1913, i_10_1914, i_10_1916, i_10_1993, i_10_2002, i_10_2003, i_10_2091, i_10_2307, i_10_2309, i_10_2350, i_10_2363, i_10_2451, i_10_2468, i_10_2473, i_10_2515, i_10_2516, i_10_2601, i_10_2658, i_10_2662, i_10_2674, i_10_2710, i_10_2721, i_10_2818, i_10_2832, i_10_2920, i_10_2983, i_10_3073, i_10_3277, i_10_3279, i_10_3356, i_10_3387, i_10_3388, i_10_3389, i_10_3391, i_10_3403, i_10_3404, i_10_3410, i_10_3523, i_10_3583, i_10_3616, i_10_3617, i_10_3649, i_10_3722, i_10_3780, i_10_3781, i_10_3782, i_10_3837, i_10_3838, i_10_3853, i_10_3858, i_10_3859, i_10_3860, i_10_3985, i_10_4027, i_10_4031, i_10_4129, i_10_4285, i_10_4290, i_10_4565, o_10_404);
	kernel_10_405 k_10_405(i_10_174, i_10_178, i_10_280, i_10_281, i_10_283, i_10_284, i_10_320, i_10_390, i_10_408, i_10_444, i_10_520, i_10_714, i_10_736, i_10_903, i_10_952, i_10_996, i_10_1005, i_10_1006, i_10_1039, i_10_1050, i_10_1051, i_10_1059, i_10_1237, i_10_1246, i_10_1249, i_10_1250, i_10_1311, i_10_1312, i_10_1313, i_10_1446, i_10_1455, i_10_1554, i_10_1555, i_10_1581, i_10_1735, i_10_1823, i_10_1909, i_10_1914, i_10_2355, i_10_2356, i_10_2364, i_10_2382, i_10_2383, i_10_2406, i_10_2407, i_10_2408, i_10_2448, i_10_2449, i_10_2451, i_10_2452, i_10_2464, i_10_2466, i_10_2467, i_10_2472, i_10_2473, i_10_2509, i_10_2607, i_10_2632, i_10_2636, i_10_2641, i_10_2662, i_10_2705, i_10_2713, i_10_2730, i_10_2733, i_10_2830, i_10_2834, i_10_2880, i_10_2884, i_10_2887, i_10_2921, i_10_2922, i_10_2986, i_10_3033, i_10_3040, i_10_3202, i_10_3291, i_10_3318, i_10_3390, i_10_3406, i_10_3613, i_10_3614, i_10_3646, i_10_3685, i_10_3725, i_10_3840, i_10_3857, i_10_3859, i_10_3896, i_10_3913, i_10_3914, i_10_3984, i_10_3985, i_10_3986, i_10_4113, i_10_4118, i_10_4276, i_10_4280, i_10_4281, i_10_4289, o_10_405);
	kernel_10_406 k_10_406(i_10_30, i_10_174, i_10_220, i_10_224, i_10_243, i_10_246, i_10_249, i_10_250, i_10_280, i_10_288, i_10_325, i_10_369, i_10_426, i_10_438, i_10_462, i_10_465, i_10_534, i_10_796, i_10_900, i_10_903, i_10_963, i_10_1235, i_10_1260, i_10_1269, i_10_1270, i_10_1359, i_10_1360, i_10_1390, i_10_1435, i_10_1443, i_10_1548, i_10_1551, i_10_1683, i_10_1809, i_10_1812, i_10_1820, i_10_1872, i_10_1971, i_10_2023, i_10_2197, i_10_2250, i_10_2259, i_10_2323, i_10_2406, i_10_2502, i_10_2505, i_10_2515, i_10_2568, i_10_2604, i_10_2607, i_10_2629, i_10_2634, i_10_2655, i_10_2660, i_10_2661, i_10_2673, i_10_2700, i_10_2704, i_10_2712, i_10_2728, i_10_2731, i_10_2784, i_10_2787, i_10_2828, i_10_2829, i_10_2921, i_10_2979, i_10_3069, i_10_3196, i_10_3235, i_10_3270, i_10_3276, i_10_3277, i_10_3384, i_10_3386, i_10_3430, i_10_3433, i_10_3492, i_10_3610, i_10_3615, i_10_3681, i_10_3849, i_10_3857, i_10_3888, i_10_3978, i_10_3981, i_10_3993, i_10_4050, i_10_4053, i_10_4117, i_10_4128, i_10_4129, i_10_4266, i_10_4287, i_10_4365, i_10_4428, i_10_4429, i_10_4458, i_10_4566, i_10_4571, o_10_406);
	kernel_10_407 k_10_407(i_10_160, i_10_175, i_10_270, i_10_278, i_10_280, i_10_281, i_10_283, i_10_329, i_10_408, i_10_431, i_10_432, i_10_443, i_10_444, i_10_445, i_10_508, i_10_509, i_10_511, i_10_711, i_10_749, i_10_898, i_10_1142, i_10_1240, i_10_1243, i_10_1244, i_10_1247, i_10_1310, i_10_1348, i_10_1541, i_10_1552, i_10_1651, i_10_1652, i_10_1690, i_10_1821, i_10_1822, i_10_1823, i_10_1826, i_10_1996, i_10_2349, i_10_2352, i_10_2353, i_10_2354, i_10_2404, i_10_2455, i_10_2635, i_10_2659, i_10_2706, i_10_2707, i_10_2721, i_10_2733, i_10_2735, i_10_2884, i_10_2888, i_10_2919, i_10_2920, i_10_2921, i_10_2923, i_10_3035, i_10_3046, i_10_3150, i_10_3154, i_10_3155, i_10_3166, i_10_3195, i_10_3199, i_10_3200, i_10_3387, i_10_3388, i_10_3389, i_10_3390, i_10_3391, i_10_3392, i_10_3405, i_10_3585, i_10_3586, i_10_3587, i_10_3610, i_10_3611, i_10_3614, i_10_3782, i_10_3784, i_10_3785, i_10_3786, i_10_3837, i_10_3838, i_10_3839, i_10_3846, i_10_3847, i_10_3851, i_10_3856, i_10_3857, i_10_3980, i_10_4121, i_10_4123, i_10_4130, i_10_4174, i_10_4175, i_10_4192, i_10_4283, i_10_4292, i_10_4564, o_10_407);
	kernel_10_408 k_10_408(i_10_216, i_10_217, i_10_218, i_10_275, i_10_278, i_10_280, i_10_281, i_10_282, i_10_283, i_10_284, i_10_316, i_10_317, i_10_319, i_10_320, i_10_444, i_10_461, i_10_464, i_10_466, i_10_467, i_10_799, i_10_851, i_10_854, i_10_1006, i_10_1027, i_10_1030, i_10_1034, i_10_1083, i_10_1237, i_10_1240, i_10_1242, i_10_1243, i_10_1307, i_10_1648, i_10_1649, i_10_1684, i_10_1685, i_10_1688, i_10_1819, i_10_2002, i_10_2305, i_10_2306, i_10_2351, i_10_2358, i_10_2362, i_10_2363, i_10_2364, i_10_2449, i_10_2460, i_10_2470, i_10_2701, i_10_2702, i_10_2703, i_10_2710, i_10_2718, i_10_2719, i_10_2720, i_10_2722, i_10_2919, i_10_2920, i_10_2921, i_10_2923, i_10_2924, i_10_3088, i_10_3089, i_10_3267, i_10_3270, i_10_3277, i_10_3322, i_10_3328, i_10_3385, i_10_3386, i_10_3402, i_10_3403, i_10_3404, i_10_3405, i_10_3406, i_10_3407, i_10_3466, i_10_3469, i_10_3551, i_10_3611, i_10_3780, i_10_3781, i_10_3783, i_10_3784, i_10_3844, i_10_3847, i_10_3851, i_10_3855, i_10_3856, i_10_3857, i_10_3979, i_10_4212, i_10_4214, i_10_4273, i_10_4284, i_10_4285, i_10_4565, i_10_4567, i_10_4569, o_10_408);
	kernel_10_409 k_10_409(i_10_27, i_10_28, i_10_30, i_10_117, i_10_216, i_10_220, i_10_221, i_10_280, i_10_283, i_10_285, i_10_286, i_10_442, i_10_465, i_10_508, i_10_514, i_10_748, i_10_893, i_10_955, i_10_961, i_10_1238, i_10_1242, i_10_1243, i_10_1244, i_10_1250, i_10_1305, i_10_1306, i_10_1308, i_10_1309, i_10_1310, i_10_1311, i_10_1359, i_10_1360, i_10_1444, i_10_1552, i_10_1575, i_10_1578, i_10_1647, i_10_1650, i_10_1819, i_10_1821, i_10_1823, i_10_1913, i_10_1947, i_10_1998, i_10_2349, i_10_2449, i_10_2450, i_10_2452, i_10_2601, i_10_2628, i_10_2629, i_10_2631, i_10_2658, i_10_2673, i_10_2710, i_10_2711, i_10_2713, i_10_2714, i_10_2721, i_10_2725, i_10_2726, i_10_2735, i_10_2784, i_10_2887, i_10_2982, i_10_3033, i_10_3034, i_10_3036, i_10_3037, i_10_3038, i_10_3039, i_10_3040, i_10_3069, i_10_3089, i_10_3281, i_10_3386, i_10_3387, i_10_3388, i_10_3390, i_10_3391, i_10_3405, i_10_3502, i_10_3519, i_10_3583, i_10_3613, i_10_3645, i_10_3646, i_10_3647, i_10_3648, i_10_3649, i_10_3652, i_10_3780, i_10_3782, i_10_3783, i_10_3834, i_10_3849, i_10_3857, i_10_4213, i_10_4292, i_10_4565, o_10_409);
	kernel_10_410 k_10_410(i_10_171, i_10_279, i_10_285, i_10_286, i_10_292, i_10_390, i_10_393, i_10_394, i_10_412, i_10_435, i_10_441, i_10_442, i_10_462, i_10_463, i_10_464, i_10_466, i_10_467, i_10_509, i_10_699, i_10_700, i_10_750, i_10_996, i_10_1237, i_10_1238, i_10_1239, i_10_1240, i_10_1241, i_10_1308, i_10_1362, i_10_1363, i_10_1542, i_10_1546, i_10_1551, i_10_1552, i_10_1554, i_10_1578, i_10_1579, i_10_1581, i_10_1690, i_10_1824, i_10_1914, i_10_2158, i_10_2159, i_10_2202, i_10_2310, i_10_2311, i_10_2312, i_10_2355, i_10_2356, i_10_2357, i_10_2360, i_10_2382, i_10_2408, i_10_2452, i_10_2481, i_10_2656, i_10_2706, i_10_2721, i_10_2880, i_10_2881, i_10_2884, i_10_2886, i_10_2958, i_10_3039, i_10_3041, i_10_3153, i_10_3158, i_10_3195, i_10_3273, i_10_3275, i_10_3279, i_10_3280, i_10_3283, i_10_3324, i_10_3325, i_10_3328, i_10_3329, i_10_3387, i_10_3390, i_10_3391, i_10_3540, i_10_3588, i_10_3782, i_10_3843, i_10_3856, i_10_3857, i_10_3859, i_10_3964, i_10_3965, i_10_3981, i_10_3982, i_10_3984, i_10_3985, i_10_4057, i_10_4115, i_10_4129, i_10_4173, i_10_4278, i_10_4279, i_10_4281, o_10_410);
	kernel_10_411 k_10_411(i_10_145, i_10_220, i_10_223, i_10_271, i_10_272, i_10_273, i_10_276, i_10_283, i_10_293, i_10_316, i_10_409, i_10_410, i_10_444, i_10_800, i_10_971, i_10_1036, i_10_1234, i_10_1237, i_10_1238, i_10_1261, i_10_1288, i_10_1309, i_10_1359, i_10_1360, i_10_1361, i_10_1431, i_10_1441, i_10_1442, i_10_1576, i_10_1578, i_10_1655, i_10_1683, i_10_1684, i_10_1688, i_10_1690, i_10_1819, i_10_1949, i_10_2180, i_10_2335, i_10_2351, i_10_2352, i_10_2363, i_10_2404, i_10_2450, i_10_2451, i_10_2459, i_10_2462, i_10_2467, i_10_2504, i_10_2634, i_10_2635, i_10_2656, i_10_2659, i_10_2663, i_10_2673, i_10_2674, i_10_2675, i_10_2714, i_10_2785, i_10_2831, i_10_2918, i_10_2919, i_10_2982, i_10_3151, i_10_3152, i_10_3153, i_10_3154, i_10_3156, i_10_3195, i_10_3196, i_10_3198, i_10_3268, i_10_3269, i_10_3271, i_10_3278, i_10_3292, i_10_3321, i_10_3522, i_10_3541, i_10_3585, i_10_3586, i_10_3587, i_10_3612, i_10_3613, i_10_3615, i_10_3651, i_10_3834, i_10_3848, i_10_3942, i_10_3944, i_10_3994, i_10_4051, i_10_4052, i_10_4114, i_10_4116, i_10_4288, i_10_4289, i_10_4563, i_10_4567, i_10_4594, o_10_411);
	kernel_10_412 k_10_412(i_10_121, i_10_125, i_10_176, i_10_220, i_10_247, i_10_285, i_10_319, i_10_408, i_10_409, i_10_410, i_10_448, i_10_565, i_10_955, i_10_958, i_10_960, i_10_962, i_10_1006, i_10_1007, i_10_1083, i_10_1136, i_10_1137, i_10_1138, i_10_1181, i_10_1237, i_10_1308, i_10_1541, i_10_1544, i_10_1552, i_10_1553, i_10_1575, i_10_1618, i_10_1652, i_10_1677, i_10_1684, i_10_1687, i_10_1819, i_10_1951, i_10_1952, i_10_2182, i_10_2184, i_10_2185, i_10_2186, i_10_2200, i_10_2312, i_10_2330, i_10_2349, i_10_2353, i_10_2355, i_10_2361, i_10_2366, i_10_2405, i_10_2411, i_10_2461, i_10_2470, i_10_2471, i_10_2473, i_10_2509, i_10_2510, i_10_2632, i_10_2633, i_10_2681, i_10_2716, i_10_2729, i_10_2833, i_10_2880, i_10_2881, i_10_2884, i_10_2885, i_10_2920, i_10_2921, i_10_2924, i_10_3038, i_10_3151, i_10_3199, i_10_3200, i_10_3203, i_10_3271, i_10_3275, i_10_3316, i_10_3323, i_10_3325, i_10_3326, i_10_3328, i_10_3329, i_10_3497, i_10_3585, i_10_3586, i_10_3617, i_10_3649, i_10_3653, i_10_3686, i_10_3782, i_10_3785, i_10_3787, i_10_3834, i_10_3838, i_10_3856, i_10_3983, i_10_4058, i_10_4567, o_10_412);
	kernel_10_413 k_10_413(i_10_283, i_10_296, i_10_321, i_10_327, i_10_328, i_10_329, i_10_330, i_10_411, i_10_436, i_10_459, i_10_461, i_10_463, i_10_464, i_10_749, i_10_793, i_10_901, i_10_969, i_10_1080, i_10_1083, i_10_1084, i_10_1217, i_10_1233, i_10_1261, i_10_1263, i_10_1264, i_10_1277, i_10_1310, i_10_1359, i_10_1432, i_10_1433, i_10_1638, i_10_1649, i_10_1655, i_10_1772, i_10_1818, i_10_1822, i_10_1909, i_10_1912, i_10_1913, i_10_2198, i_10_2351, i_10_2353, i_10_2357, i_10_2361, i_10_2379, i_10_2453, i_10_2466, i_10_2467, i_10_2504, i_10_2629, i_10_2630, i_10_2656, i_10_2660, i_10_2702, i_10_2705, i_10_2715, i_10_2717, i_10_2735, i_10_2826, i_10_2827, i_10_2828, i_10_2877, i_10_2917, i_10_2921, i_10_2979, i_10_2980, i_10_2981, i_10_3036, i_10_3040, i_10_3077, i_10_3278, i_10_3326, i_10_3329, i_10_3384, i_10_3403, i_10_3433, i_10_3523, i_10_3526, i_10_3611, i_10_3615, i_10_3646, i_10_3647, i_10_3648, i_10_3650, i_10_3682, i_10_3719, i_10_3837, i_10_3853, i_10_3856, i_10_3888, i_10_3889, i_10_3890, i_10_3987, i_10_3991, i_10_4027, i_10_4124, i_10_4208, i_10_4211, i_10_4276, i_10_4291, o_10_413);
	kernel_10_414 k_10_414(i_10_172, i_10_174, i_10_175, i_10_216, i_10_220, i_10_221, i_10_224, i_10_279, i_10_315, i_10_317, i_10_387, i_10_411, i_10_446, i_10_459, i_10_461, i_10_712, i_10_797, i_10_898, i_10_962, i_10_1000, i_10_1003, i_10_1237, i_10_1238, i_10_1310, i_10_1312, i_10_1431, i_10_1432, i_10_1433, i_10_1576, i_10_1577, i_10_1580, i_10_1581, i_10_1651, i_10_1683, i_10_1686, i_10_1820, i_10_1822, i_10_1913, i_10_2186, i_10_2197, i_10_2349, i_10_2350, i_10_2356, i_10_2358, i_10_2410, i_10_2452, i_10_2453, i_10_2460, i_10_2468, i_10_2502, i_10_2661, i_10_2700, i_10_2701, i_10_2713, i_10_2714, i_10_2716, i_10_2717, i_10_2719, i_10_2721, i_10_2722, i_10_2723, i_10_2885, i_10_2924, i_10_3036, i_10_3050, i_10_3069, i_10_3070, i_10_3280, i_10_3384, i_10_3385, i_10_3390, i_10_3391, i_10_3403, i_10_3405, i_10_3406, i_10_3409, i_10_3523, i_10_3613, i_10_3647, i_10_3648, i_10_3651, i_10_3785, i_10_3855, i_10_3856, i_10_3857, i_10_3860, i_10_3978, i_10_3980, i_10_3982, i_10_3983, i_10_4029, i_10_4117, i_10_4118, i_10_4169, i_10_4284, i_10_4285, i_10_4288, i_10_4290, i_10_4565, i_10_4567, o_10_414);
	kernel_10_415 k_10_415(i_10_148, i_10_222, i_10_247, i_10_258, i_10_259, i_10_279, i_10_282, i_10_436, i_10_442, i_10_463, i_10_464, i_10_566, i_10_589, i_10_694, i_10_718, i_10_735, i_10_736, i_10_752, i_10_792, i_10_797, i_10_957, i_10_1029, i_10_1031, i_10_1033, i_10_1050, i_10_1051, i_10_1052, i_10_1159, i_10_1160, i_10_1262, i_10_1310, i_10_1311, i_10_1439, i_10_1443, i_10_1454, i_10_1546, i_10_1613, i_10_1633, i_10_1634, i_10_1635, i_10_1636, i_10_1637, i_10_1651, i_10_1652, i_10_1684, i_10_1688, i_10_1821, i_10_1912, i_10_1914, i_10_1939, i_10_2002, i_10_2150, i_10_2181, i_10_2185, i_10_2186, i_10_2366, i_10_2433, i_10_2435, i_10_2679, i_10_2680, i_10_2714, i_10_2717, i_10_2725, i_10_2733, i_10_2829, i_10_2831, i_10_2884, i_10_2888, i_10_3093, i_10_3094, i_10_3095, i_10_3199, i_10_3201, i_10_3236, i_10_3271, i_10_3503, i_10_3562, i_10_3586, i_10_3587, i_10_3588, i_10_3617, i_10_3653, i_10_3721, i_10_3781, i_10_3784, i_10_3787, i_10_3838, i_10_3943, i_10_3944, i_10_3945, i_10_3981, i_10_3983, i_10_3985, i_10_4031, i_10_4117, i_10_4121, i_10_4183, i_10_4226, i_10_4270, i_10_4375, o_10_415);
	kernel_10_416 k_10_416(i_10_144, i_10_174, i_10_216, i_10_236, i_10_279, i_10_426, i_10_433, i_10_435, i_10_441, i_10_442, i_10_443, i_10_444, i_10_446, i_10_463, i_10_515, i_10_518, i_10_792, i_10_793, i_10_794, i_10_820, i_10_892, i_10_957, i_10_967, i_10_1083, i_10_1084, i_10_1202, i_10_1360, i_10_1377, i_10_1485, i_10_1546, i_10_1576, i_10_1581, i_10_1631, i_10_1691, i_10_1728, i_10_1818, i_10_1820, i_10_1954, i_10_2045, i_10_2200, i_10_2202, i_10_2225, i_10_2288, i_10_2331, i_10_2352, i_10_2357, i_10_2358, i_10_2360, i_10_2377, i_10_2467, i_10_2514, i_10_2568, i_10_2629, i_10_2631, i_10_2632, i_10_2642, i_10_2660, i_10_2702, i_10_2713, i_10_2719, i_10_2722, i_10_2727, i_10_2729, i_10_2746, i_10_2917, i_10_3033, i_10_3290, i_10_3384, i_10_3386, i_10_3387, i_10_3388, i_10_3389, i_10_3448, i_10_3465, i_10_3556, i_10_3584, i_10_3601, i_10_3614, i_10_3787, i_10_3788, i_10_3844, i_10_3845, i_10_3848, i_10_3890, i_10_3974, i_10_3978, i_10_3990, i_10_4126, i_10_4167, i_10_4168, i_10_4187, i_10_4268, i_10_4275, i_10_4288, i_10_4307, i_10_4394, i_10_4395, i_10_4397, i_10_4447, i_10_4572, o_10_416);
	kernel_10_417 k_10_417(i_10_46, i_10_175, i_10_177, i_10_219, i_10_222, i_10_284, i_10_319, i_10_322, i_10_327, i_10_330, i_10_331, i_10_442, i_10_751, i_10_955, i_10_1032, i_10_1034, i_10_1237, i_10_1239, i_10_1240, i_10_1248, i_10_1308, i_10_1311, i_10_1363, i_10_1431, i_10_1444, i_10_1541, i_10_1549, i_10_1553, i_10_1556, i_10_1576, i_10_1577, i_10_1683, i_10_1803, i_10_1820, i_10_1826, i_10_1948, i_10_1981, i_10_1996, i_10_2017, i_10_2019, i_10_2028, i_10_2355, i_10_2357, i_10_2462, i_10_2466, i_10_2508, i_10_2608, i_10_2629, i_10_2631, i_10_2658, i_10_2659, i_10_2662, i_10_2663, i_10_2704, i_10_2723, i_10_2724, i_10_2725, i_10_2726, i_10_2731, i_10_2739, i_10_2742, i_10_2782, i_10_2823, i_10_2830, i_10_2831, i_10_2832, i_10_2833, i_10_2834, i_10_2880, i_10_2982, i_10_3049, i_10_3090, i_10_3270, i_10_3278, i_10_3279, i_10_3283, i_10_3469, i_10_3582, i_10_3612, i_10_3645, i_10_3648, i_10_3649, i_10_3650, i_10_3651, i_10_3780, i_10_3835, i_10_3837, i_10_3841, i_10_3860, i_10_3895, i_10_3896, i_10_4113, i_10_4116, i_10_4123, i_10_4275, i_10_4276, i_10_4279, i_10_4290, i_10_4291, i_10_4581, o_10_417);
	kernel_10_418 k_10_418(i_10_274, i_10_275, i_10_282, i_10_317, i_10_328, i_10_432, i_10_433, i_10_434, i_10_436, i_10_437, i_10_446, i_10_460, i_10_463, i_10_464, i_10_518, i_10_907, i_10_1032, i_10_1033, i_10_1043, i_10_1138, i_10_1265, i_10_1309, i_10_1345, i_10_1346, i_10_1349, i_10_1445, i_10_1546, i_10_1575, i_10_1654, i_10_1720, i_10_1767, i_10_1768, i_10_1769, i_10_1821, i_10_1912, i_10_1913, i_10_1916, i_10_2352, i_10_2365, i_10_2383, i_10_2384, i_10_2408, i_10_2471, i_10_2512, i_10_2629, i_10_2630, i_10_2656, i_10_2657, i_10_2659, i_10_2660, i_10_2661, i_10_2675, i_10_2678, i_10_2681, i_10_2705, i_10_2723, i_10_2728, i_10_2729, i_10_2819, i_10_2822, i_10_2823, i_10_2824, i_10_2828, i_10_2830, i_10_2831, i_10_2880, i_10_2919, i_10_2980, i_10_3033, i_10_3034, i_10_3050, i_10_3070, i_10_3088, i_10_3093, i_10_3150, i_10_3151, i_10_3160, i_10_3280, i_10_3281, i_10_3322, i_10_3323, i_10_3349, i_10_3350, i_10_3387, i_10_3437, i_10_3523, i_10_3587, i_10_3590, i_10_3613, i_10_3648, i_10_3685, i_10_3842, i_10_3856, i_10_3857, i_10_3910, i_10_4115, i_10_4175, i_10_4236, i_10_4267, i_10_4289, o_10_418);
	kernel_10_419 k_10_419(i_10_145, i_10_174, i_10_217, i_10_282, i_10_287, i_10_293, i_10_296, i_10_430, i_10_443, i_10_459, i_10_462, i_10_465, i_10_581, i_10_699, i_10_751, i_10_794, i_10_798, i_10_835, i_10_894, i_10_897, i_10_1030, i_10_1040, i_10_1043, i_10_1234, i_10_1235, i_10_1236, i_10_1239, i_10_1240, i_10_1248, i_10_1249, i_10_1309, i_10_1311, i_10_1312, i_10_1344, i_10_1575, i_10_1637, i_10_1648, i_10_1650, i_10_1651, i_10_1655, i_10_1684, i_10_1685, i_10_1686, i_10_1697, i_10_1798, i_10_1822, i_10_2166, i_10_2201, i_10_2266, i_10_2327, i_10_2337, i_10_2338, i_10_2339, i_10_2449, i_10_2451, i_10_2510, i_10_2559, i_10_2562, i_10_2571, i_10_2636, i_10_2643, i_10_2652, i_10_2661, i_10_2662, i_10_2705, i_10_2708, i_10_2717, i_10_2781, i_10_2782, i_10_2984, i_10_3076, i_10_3201, i_10_3268, i_10_3270, i_10_3272, i_10_3273, i_10_3274, i_10_3280, i_10_3405, i_10_3611, i_10_3612, i_10_3649, i_10_3652, i_10_3703, i_10_3704, i_10_3783, i_10_3784, i_10_3785, i_10_3787, i_10_3838, i_10_3859, i_10_3896, i_10_4027, i_10_4269, i_10_4276, i_10_4277, i_10_4281, i_10_4292, i_10_4463, i_10_4508, o_10_419);
	kernel_10_420 k_10_420(i_10_151, i_10_157, i_10_268, i_10_273, i_10_278, i_10_282, i_10_283, i_10_322, i_10_391, i_10_442, i_10_508, i_10_691, i_10_716, i_10_718, i_10_719, i_10_739, i_10_754, i_10_755, i_10_795, i_10_931, i_10_959, i_10_966, i_10_968, i_10_970, i_10_991, i_10_992, i_10_1165, i_10_1166, i_10_1197, i_10_1198, i_10_1235, i_10_1249, i_10_1250, i_10_1262, i_10_1359, i_10_1360, i_10_1440, i_10_1441, i_10_1442, i_10_1491, i_10_1492, i_10_1536, i_10_1537, i_10_1555, i_10_1582, i_10_1629, i_10_1691, i_10_1852, i_10_2002, i_10_2005, i_10_2006, i_10_2019, i_10_2186, i_10_2351, i_10_2392, i_10_2533, i_10_2535, i_10_2573, i_10_2609, i_10_2620, i_10_2621, i_10_2680, i_10_2708, i_10_2725, i_10_2727, i_10_2735, i_10_2781, i_10_2786, i_10_2882, i_10_2885, i_10_2919, i_10_2920, i_10_2982, i_10_3038, i_10_3238, i_10_3384, i_10_3385, i_10_3386, i_10_3392, i_10_3561, i_10_3562, i_10_3719, i_10_3786, i_10_3787, i_10_3846, i_10_3857, i_10_3877, i_10_3897, i_10_3898, i_10_3912, i_10_3913, i_10_3914, i_10_4113, i_10_4116, i_10_4118, i_10_4121, i_10_4204, i_10_4339, i_10_4460, i_10_4463, o_10_420);
	kernel_10_421 k_10_421(i_10_49, i_10_151, i_10_183, i_10_184, i_10_222, i_10_410, i_10_441, i_10_442, i_10_444, i_10_445, i_10_514, i_10_515, i_10_588, i_10_628, i_10_711, i_10_745, i_10_797, i_10_832, i_10_966, i_10_982, i_10_983, i_10_1005, i_10_1026, i_10_1033, i_10_1034, i_10_1086, i_10_1240, i_10_1250, i_10_1305, i_10_1308, i_10_1309, i_10_1345, i_10_1383, i_10_1385, i_10_1432, i_10_1438, i_10_1532, i_10_1647, i_10_1683, i_10_1743, i_10_1821, i_10_1822, i_10_1823, i_10_1995, i_10_1996, i_10_2094, i_10_2095, i_10_2180, i_10_2197, i_10_2243, i_10_2252, i_10_2355, i_10_2356, i_10_2451, i_10_2452, i_10_2453, i_10_2474, i_10_2514, i_10_2515, i_10_2516, i_10_2644, i_10_2679, i_10_2680, i_10_2722, i_10_2724, i_10_2734, i_10_2735, i_10_2740, i_10_2741, i_10_2831, i_10_2916, i_10_2917, i_10_2921, i_10_2922, i_10_2923, i_10_3039, i_10_3040, i_10_3195, i_10_3388, i_10_3389, i_10_3405, i_10_3453, i_10_3525, i_10_3586, i_10_3726, i_10_3781, i_10_3786, i_10_3855, i_10_3856, i_10_3982, i_10_4026, i_10_4121, i_10_4182, i_10_4188, i_10_4219, i_10_4220, i_10_4272, i_10_4292, i_10_4426, i_10_4570, o_10_421);
	kernel_10_422 k_10_422(i_10_32, i_10_33, i_10_34, i_10_53, i_10_143, i_10_172, i_10_178, i_10_179, i_10_188, i_10_265, i_10_269, i_10_274, i_10_277, i_10_278, i_10_391, i_10_440, i_10_462, i_10_464, i_10_520, i_10_755, i_10_934, i_10_962, i_10_1033, i_10_1061, i_10_1236, i_10_1237, i_10_1239, i_10_1240, i_10_1241, i_10_1246, i_10_1250, i_10_1308, i_10_1311, i_10_1382, i_10_1385, i_10_1436, i_10_1547, i_10_1653, i_10_1689, i_10_1819, i_10_1822, i_10_1824, i_10_1825, i_10_1956, i_10_1997, i_10_2201, i_10_2357, i_10_2363, i_10_2452, i_10_2460, i_10_2462, i_10_2469, i_10_2471, i_10_2474, i_10_2514, i_10_2517, i_10_2616, i_10_2630, i_10_2663, i_10_2711, i_10_2733, i_10_2735, i_10_2788, i_10_2789, i_10_2828, i_10_2832, i_10_2868, i_10_3035, i_10_3047, i_10_3196, i_10_3199, i_10_3203, i_10_3281, i_10_3454, i_10_3455, i_10_3470, i_10_3544, i_10_3552, i_10_3587, i_10_3611, i_10_3617, i_10_3650, i_10_3653, i_10_3683, i_10_3704, i_10_3785, i_10_3786, i_10_3788, i_10_3834, i_10_3835, i_10_3838, i_10_3847, i_10_3886, i_10_3887, i_10_3995, i_10_4004, i_10_4055, i_10_4057, i_10_4058, i_10_4382, o_10_422);
	kernel_10_423 k_10_423(i_10_36, i_10_51, i_10_172, i_10_224, i_10_244, i_10_253, i_10_256, i_10_263, i_10_286, i_10_321, i_10_410, i_10_412, i_10_445, i_10_502, i_10_906, i_10_958, i_10_961, i_10_1030, i_10_1033, i_10_1034, i_10_1248, i_10_1249, i_10_1260, i_10_1310, i_10_1311, i_10_1346, i_10_1359, i_10_1434, i_10_1436, i_10_1451, i_10_1543, i_10_1576, i_10_1622, i_10_1651, i_10_1683, i_10_1687, i_10_1818, i_10_1819, i_10_1820, i_10_1821, i_10_1825, i_10_1909, i_10_1911, i_10_1912, i_10_1945, i_10_1950, i_10_1951, i_10_2182, i_10_2183, i_10_2304, i_10_2306, i_10_2350, i_10_2351, i_10_2356, i_10_2357, i_10_2362, i_10_2378, i_10_2384, i_10_2405, i_10_2451, i_10_2452, i_10_2453, i_10_2471, i_10_2518, i_10_2676, i_10_2715, i_10_2757, i_10_2850, i_10_2918, i_10_2921, i_10_3033, i_10_3070, i_10_3167, i_10_3198, i_10_3199, i_10_3278, i_10_3279, i_10_3326, i_10_3331, i_10_3432, i_10_3616, i_10_3645, i_10_3653, i_10_3721, i_10_3733, i_10_3787, i_10_3835, i_10_3839, i_10_3842, i_10_3852, i_10_3860, i_10_3983, i_10_4054, i_10_4116, i_10_4117, i_10_4119, i_10_4120, i_10_4168, i_10_4169, i_10_4277, o_10_423);
	kernel_10_424 k_10_424(i_10_150, i_10_172, i_10_174, i_10_182, i_10_285, i_10_327, i_10_410, i_10_444, i_10_447, i_10_513, i_10_516, i_10_717, i_10_795, i_10_797, i_10_798, i_10_963, i_10_964, i_10_966, i_10_967, i_10_1139, i_10_1163, i_10_1305, i_10_1308, i_10_1309, i_10_1311, i_10_1440, i_10_1444, i_10_1447, i_10_1491, i_10_1492, i_10_1556, i_10_1581, i_10_1582, i_10_1618, i_10_1635, i_10_1641, i_10_1726, i_10_1821, i_10_1824, i_10_1951, i_10_2184, i_10_2310, i_10_2322, i_10_2328, i_10_2351, i_10_2352, i_10_2377, i_10_2449, i_10_2472, i_10_2519, i_10_2660, i_10_2673, i_10_2679, i_10_2701, i_10_2727, i_10_2830, i_10_2880, i_10_2883, i_10_2885, i_10_2924, i_10_3035, i_10_3037, i_10_3038, i_10_3120, i_10_3152, i_10_3196, i_10_3198, i_10_3273, i_10_3323, i_10_3387, i_10_3405, i_10_3465, i_10_3468, i_10_3469, i_10_3495, i_10_3496, i_10_3585, i_10_3588, i_10_3610, i_10_3612, i_10_3613, i_10_3780, i_10_3805, i_10_3838, i_10_3840, i_10_3850, i_10_3853, i_10_3948, i_10_4120, i_10_4123, i_10_4213, i_10_4266, i_10_4270, i_10_4285, i_10_4287, i_10_4291, i_10_4458, i_10_4461, i_10_4564, i_10_4567, o_10_424);
	kernel_10_425 k_10_425(i_10_86, i_10_221, i_10_286, i_10_287, i_10_293, i_10_315, i_10_410, i_10_428, i_10_437, i_10_443, i_10_444, i_10_448, i_10_455, i_10_520, i_10_700, i_10_794, i_10_798, i_10_881, i_10_971, i_10_1004, i_10_1026, i_10_1103, i_10_1235, i_10_1238, i_10_1240, i_10_1364, i_10_1432, i_10_1436, i_10_1577, i_10_1654, i_10_1688, i_10_1821, i_10_1875, i_10_1909, i_10_1913, i_10_1925, i_10_1952, i_10_2186, i_10_2363, i_10_2365, i_10_2366, i_10_2408, i_10_2451, i_10_2454, i_10_2455, i_10_2456, i_10_2470, i_10_2519, i_10_2617, i_10_2630, i_10_2645, i_10_2660, i_10_2681, i_10_2710, i_10_2719, i_10_2734, i_10_2882, i_10_2888, i_10_2923, i_10_2924, i_10_2986, i_10_3040, i_10_3041, i_10_3047, i_10_3049, i_10_3086, i_10_3153, i_10_3155, i_10_3156, i_10_3199, i_10_3202, i_10_3277, i_10_3283, i_10_3284, i_10_3302, i_10_3387, i_10_3389, i_10_3410, i_10_3465, i_10_3469, i_10_3503, i_10_3562, i_10_3613, i_10_3733, i_10_3785, i_10_3839, i_10_3853, i_10_3856, i_10_3857, i_10_3859, i_10_4030, i_10_4057, i_10_4058, i_10_4113, i_10_4117, i_10_4129, i_10_4130, i_10_4148, i_10_4237, i_10_4292, o_10_425);
	kernel_10_426 k_10_426(i_10_218, i_10_244, i_10_282, i_10_283, i_10_284, i_10_285, i_10_286, i_10_316, i_10_317, i_10_318, i_10_319, i_10_388, i_10_406, i_10_432, i_10_436, i_10_437, i_10_444, i_10_445, i_10_459, i_10_460, i_10_462, i_10_463, i_10_514, i_10_693, i_10_749, i_10_793, i_10_900, i_10_1000, i_10_1026, i_10_1027, i_10_1233, i_10_1242, i_10_1306, i_10_1441, i_10_1442, i_10_1546, i_10_1549, i_10_1650, i_10_1654, i_10_1819, i_10_1821, i_10_1822, i_10_1908, i_10_1946, i_10_1950, i_10_2304, i_10_2305, i_10_2306, i_10_2350, i_10_2359, i_10_2365, i_10_2404, i_10_2452, i_10_2454, i_10_2455, i_10_2459, i_10_2476, i_10_2477, i_10_2628, i_10_2629, i_10_2630, i_10_2632, i_10_2637, i_10_2638, i_10_2656, i_10_2657, i_10_2704, i_10_2817, i_10_2826, i_10_2827, i_10_2880, i_10_2918, i_10_2981, i_10_3034, i_10_3035, i_10_3047, i_10_3160, i_10_3200, i_10_3267, i_10_3271, i_10_3358, i_10_3384, i_10_3389, i_10_3402, i_10_3403, i_10_3404, i_10_3611, i_10_3613, i_10_3648, i_10_3682, i_10_3785, i_10_3808, i_10_3837, i_10_3843, i_10_3852, i_10_3859, i_10_3899, i_10_4171, i_10_4212, i_10_4276, o_10_426);
	kernel_10_427 k_10_427(i_10_171, i_10_243, i_10_282, i_10_284, i_10_392, i_10_425, i_10_434, i_10_442, i_10_464, i_10_748, i_10_957, i_10_958, i_10_961, i_10_1000, i_10_1003, i_10_1084, i_10_1307, i_10_1311, i_10_1362, i_10_1378, i_10_1450, i_10_1451, i_10_1551, i_10_1583, i_10_1633, i_10_1652, i_10_1653, i_10_1655, i_10_1686, i_10_1820, i_10_1945, i_10_1946, i_10_1948, i_10_1949, i_10_1990, i_10_1991, i_10_1994, i_10_2092, i_10_2201, i_10_2305, i_10_2306, i_10_2310, i_10_2311, i_10_2324, i_10_2350, i_10_2351, i_10_2354, i_10_2376, i_10_2377, i_10_2407, i_10_2449, i_10_2450, i_10_2506, i_10_2611, i_10_2612, i_10_2634, i_10_2635, i_10_2656, i_10_2658, i_10_2659, i_10_2663, i_10_2673, i_10_2674, i_10_2675, i_10_2703, i_10_2728, i_10_2729, i_10_2827, i_10_2833, i_10_3037, i_10_3038, i_10_3072, i_10_3087, i_10_3088, i_10_3089, i_10_3195, i_10_3270, i_10_3286, i_10_3350, i_10_3384, i_10_3448, i_10_3542, i_10_3614, i_10_3616, i_10_3786, i_10_3788, i_10_3838, i_10_3839, i_10_3857, i_10_3880, i_10_3944, i_10_4006, i_10_4024, i_10_4113, i_10_4219, i_10_4268, i_10_4286, i_10_4289, i_10_4474, i_10_4591, o_10_427);
	kernel_10_428 k_10_428(i_10_19, i_10_33, i_10_35, i_10_69, i_10_393, i_10_426, i_10_427, i_10_429, i_10_467, i_10_534, i_10_535, i_10_538, i_10_539, i_10_642, i_10_948, i_10_1007, i_10_1039, i_10_1187, i_10_1200, i_10_1263, i_10_1305, i_10_1317, i_10_1320, i_10_1321, i_10_1342, i_10_1348, i_10_1413, i_10_1425, i_10_1444, i_10_1446, i_10_1447, i_10_1544, i_10_1552, i_10_1605, i_10_1617, i_10_1648, i_10_1713, i_10_1761, i_10_1912, i_10_1993, i_10_2291, i_10_2355, i_10_2436, i_10_2448, i_10_2556, i_10_2826, i_10_2834, i_10_2880, i_10_2881, i_10_2917, i_10_2919, i_10_2920, i_10_2922, i_10_2923, i_10_3034, i_10_3039, i_10_3040, i_10_3043, i_10_3087, i_10_3090, i_10_3091, i_10_3093, i_10_3094, i_10_3130, i_10_3268, i_10_3270, i_10_3279, i_10_3280, i_10_3283, i_10_3321, i_10_3384, i_10_3408, i_10_3409, i_10_3436, i_10_3495, i_10_3520, i_10_3523, i_10_3544, i_10_3609, i_10_3612, i_10_3615, i_10_3724, i_10_3734, i_10_3816, i_10_3832, i_10_3855, i_10_3856, i_10_3895, i_10_3898, i_10_4120, i_10_4121, i_10_4209, i_10_4219, i_10_4351, i_10_4411, i_10_4458, i_10_4557, i_10_4569, i_10_4593, i_10_4597, o_10_428);
	kernel_10_429 k_10_429(i_10_89, i_10_121, i_10_122, i_10_156, i_10_157, i_10_174, i_10_175, i_10_177, i_10_185, i_10_248, i_10_280, i_10_287, i_10_388, i_10_391, i_10_392, i_10_410, i_10_445, i_10_446, i_10_561, i_10_629, i_10_795, i_10_1005, i_10_1084, i_10_1305, i_10_1308, i_10_1432, i_10_1433, i_10_1439, i_10_1489, i_10_1552, i_10_1578, i_10_1579, i_10_1650, i_10_1689, i_10_1726, i_10_1771, i_10_1795, i_10_1796, i_10_1952, i_10_2001, i_10_2246, i_10_2356, i_10_2357, i_10_2365, i_10_2403, i_10_2407, i_10_2410, i_10_2446, i_10_2447, i_10_2453, i_10_2472, i_10_2519, i_10_2615, i_10_2634, i_10_2643, i_10_2644, i_10_2731, i_10_2733, i_10_2734, i_10_2735, i_10_2744, i_10_2829, i_10_2830, i_10_2869, i_10_2885, i_10_2916, i_10_3235, i_10_3279, i_10_3280, i_10_3281, i_10_3283, i_10_3284, i_10_3298, i_10_3299, i_10_3318, i_10_3390, i_10_3466, i_10_3583, i_10_3614, i_10_3705, i_10_3729, i_10_3837, i_10_3841, i_10_3860, i_10_3923, i_10_3981, i_10_3984, i_10_3985, i_10_3986, i_10_4026, i_10_4028, i_10_4056, i_10_4120, i_10_4129, i_10_4172, i_10_4175, i_10_4266, i_10_4267, i_10_4282, i_10_4302, o_10_429);
	kernel_10_430 k_10_430(i_10_50, i_10_172, i_10_179, i_10_217, i_10_218, i_10_220, i_10_263, i_10_287, i_10_325, i_10_327, i_10_328, i_10_392, i_10_500, i_10_509, i_10_1000, i_10_1001, i_10_1030, i_10_1031, i_10_1040, i_10_1088, i_10_1102, i_10_1234, i_10_1238, i_10_1239, i_10_1262, i_10_1431, i_10_1433, i_10_1540, i_10_1578, i_10_1634, i_10_1643, i_10_1651, i_10_1652, i_10_1654, i_10_1688, i_10_1691, i_10_1730, i_10_1769, i_10_1820, i_10_1822, i_10_1982, i_10_2003, i_10_2006, i_10_2030, i_10_2198, i_10_2201, i_10_2204, i_10_2246, i_10_2255, i_10_2354, i_10_2364, i_10_2449, i_10_2450, i_10_2451, i_10_2452, i_10_2455, i_10_2468, i_10_2474, i_10_2567, i_10_2632, i_10_2636, i_10_2702, i_10_2704, i_10_2711, i_10_2714, i_10_2720, i_10_2732, i_10_2733, i_10_2741, i_10_2825, i_10_2830, i_10_2916, i_10_2966, i_10_3044, i_10_3071, i_10_3072, i_10_3268, i_10_3281, i_10_3314, i_10_3317, i_10_3389, i_10_3390, i_10_3391, i_10_3467, i_10_3473, i_10_3503, i_10_3506, i_10_3509, i_10_3584, i_10_3590, i_10_3841, i_10_3848, i_10_4028, i_10_4121, i_10_4123, i_10_4268, i_10_4283, i_10_4292, i_10_4565, i_10_4566, o_10_430);
	kernel_10_431 k_10_431(i_10_27, i_10_148, i_10_180, i_10_181, i_10_217, i_10_221, i_10_244, i_10_245, i_10_257, i_10_280, i_10_284, i_10_289, i_10_405, i_10_407, i_10_408, i_10_409, i_10_463, i_10_516, i_10_517, i_10_715, i_10_716, i_10_748, i_10_796, i_10_1009, i_10_1027, i_10_1028, i_10_1030, i_10_1085, i_10_1233, i_10_1234, i_10_1243, i_10_1246, i_10_1247, i_10_1539, i_10_1540, i_10_1550, i_10_1684, i_10_1685, i_10_1687, i_10_1729, i_10_1730, i_10_1801, i_10_1818, i_10_1821, i_10_1912, i_10_1999, i_10_2179, i_10_2288, i_10_2349, i_10_2353, i_10_2449, i_10_2450, i_10_2457, i_10_2470, i_10_2511, i_10_2543, i_10_2601, i_10_2604, i_10_2631, i_10_2660, i_10_2675, i_10_2728, i_10_3043, i_10_3069, i_10_3070, i_10_3198, i_10_3199, i_10_3200, i_10_3268, i_10_3386, i_10_3555, i_10_3583, i_10_3584, i_10_3587, i_10_3613, i_10_3618, i_10_3619, i_10_3650, i_10_3682, i_10_3785, i_10_3838, i_10_3856, i_10_3871, i_10_3946, i_10_3995, i_10_4010, i_10_4024, i_10_4025, i_10_4113, i_10_4114, i_10_4168, i_10_4213, i_10_4216, i_10_4267, i_10_4275, i_10_4276, i_10_4279, i_10_4285, i_10_4288, i_10_4568, o_10_431);
	kernel_10_432 k_10_432(i_10_30, i_10_40, i_10_123, i_10_124, i_10_180, i_10_184, i_10_186, i_10_286, i_10_316, i_10_318, i_10_393, i_10_440, i_10_449, i_10_463, i_10_465, i_10_466, i_10_799, i_10_1137, i_10_1233, i_10_1234, i_10_1236, i_10_1237, i_10_1239, i_10_1240, i_10_1248, i_10_1361, i_10_1362, i_10_1363, i_10_1364, i_10_1365, i_10_1546, i_10_1552, i_10_1617, i_10_1680, i_10_1686, i_10_1688, i_10_1820, i_10_1821, i_10_1822, i_10_1947, i_10_1950, i_10_2355, i_10_2408, i_10_2450, i_10_2453, i_10_2565, i_10_2631, i_10_2636, i_10_2656, i_10_2679, i_10_2713, i_10_2719, i_10_2723, i_10_2727, i_10_2730, i_10_2828, i_10_2830, i_10_2832, i_10_2880, i_10_2980, i_10_3035, i_10_3036, i_10_3037, i_10_3039, i_10_3040, i_10_3048, i_10_3093, i_10_3195, i_10_3196, i_10_3198, i_10_3276, i_10_3278, i_10_3279, i_10_3284, i_10_3322, i_10_3325, i_10_3385, i_10_3386, i_10_3387, i_10_3388, i_10_3391, i_10_3406, i_10_3430, i_10_3468, i_10_3522, i_10_3586, i_10_3648, i_10_3649, i_10_3651, i_10_3681, i_10_3781, i_10_3839, i_10_3855, i_10_3882, i_10_3894, i_10_4053, i_10_4056, i_10_4274, i_10_4569, i_10_4570, o_10_432);
	kernel_10_433 k_10_433(i_10_135, i_10_171, i_10_174, i_10_177, i_10_258, i_10_280, i_10_285, i_10_286, i_10_316, i_10_390, i_10_463, i_10_467, i_10_687, i_10_747, i_10_796, i_10_1026, i_10_1027, i_10_1032, i_10_1236, i_10_1237, i_10_1238, i_10_1240, i_10_1241, i_10_1245, i_10_1249, i_10_1250, i_10_1308, i_10_1578, i_10_1582, i_10_1651, i_10_1684, i_10_1686, i_10_1691, i_10_1819, i_10_1821, i_10_1822, i_10_2001, i_10_2199, i_10_2304, i_10_2353, i_10_2356, i_10_2455, i_10_2460, i_10_2463, i_10_2467, i_10_2470, i_10_2471, i_10_2473, i_10_2474, i_10_2514, i_10_2535, i_10_2628, i_10_2631, i_10_2635, i_10_2655, i_10_2656, i_10_2658, i_10_2659, i_10_2674, i_10_2710, i_10_2827, i_10_2829, i_10_3034, i_10_3195, i_10_3196, i_10_3201, i_10_3202, i_10_3277, i_10_3387, i_10_3389, i_10_3402, i_10_3438, i_10_3441, i_10_3585, i_10_3586, i_10_3587, i_10_3609, i_10_3613, i_10_3614, i_10_3615, i_10_3783, i_10_3786, i_10_3787, i_10_3838, i_10_3840, i_10_3852, i_10_3858, i_10_3943, i_10_3982, i_10_4008, i_10_4113, i_10_4126, i_10_4169, i_10_4219, i_10_4289, i_10_4291, i_10_4292, i_10_4567, i_10_4569, i_10_4580, o_10_433);
	kernel_10_434 k_10_434(i_10_171, i_10_217, i_10_218, i_10_219, i_10_220, i_10_223, i_10_251, i_10_278, i_10_296, i_10_316, i_10_317, i_10_328, i_10_329, i_10_331, i_10_408, i_10_411, i_10_412, i_10_432, i_10_441, i_10_445, i_10_449, i_10_458, i_10_467, i_10_507, i_10_793, i_10_991, i_10_1046, i_10_1234, i_10_1243, i_10_1261, i_10_1263, i_10_1264, i_10_1265, i_10_1267, i_10_1308, i_10_1309, i_10_1311, i_10_1432, i_10_1577, i_10_1579, i_10_1721, i_10_1809, i_10_1818, i_10_1824, i_10_1912, i_10_1915, i_10_1916, i_10_1945, i_10_2018, i_10_2353, i_10_2355, i_10_2358, i_10_2632, i_10_2635, i_10_2700, i_10_2702, i_10_2722, i_10_2788, i_10_2817, i_10_2829, i_10_2830, i_10_2831, i_10_2833, i_10_2919, i_10_2920, i_10_2923, i_10_3037, i_10_3043, i_10_3196, i_10_3203, i_10_3279, i_10_3280, i_10_3321, i_10_3384, i_10_3385, i_10_3392, i_10_3470, i_10_3614, i_10_3650, i_10_3720, i_10_3721, i_10_3781, i_10_3785, i_10_3786, i_10_3787, i_10_3834, i_10_3839, i_10_3844, i_10_3849, i_10_3852, i_10_3853, i_10_3855, i_10_3871, i_10_3895, i_10_4266, i_10_4284, i_10_4286, i_10_4287, i_10_4288, i_10_4289, o_10_434);
	kernel_10_435 k_10_435(i_10_32, i_10_121, i_10_254, i_10_392, i_10_406, i_10_434, i_10_440, i_10_459, i_10_572, i_10_694, i_10_739, i_10_947, i_10_958, i_10_990, i_10_991, i_10_1002, i_10_1003, i_10_1157, i_10_1201, i_10_1207, i_10_1270, i_10_1312, i_10_1313, i_10_1346, i_10_1451, i_10_1454, i_10_1544, i_10_1549, i_10_1550, i_10_1553, i_10_1577, i_10_1580, i_10_1582, i_10_1622, i_10_1633, i_10_1714, i_10_1803, i_10_1825, i_10_1876, i_10_1909, i_10_1985, i_10_2003, i_10_2017, i_10_2024, i_10_2027, i_10_2153, i_10_2155, i_10_2204, i_10_2291, i_10_2304, i_10_2309, i_10_2351, i_10_2384, i_10_2458, i_10_2517, i_10_2567, i_10_2576, i_10_2585, i_10_2593, i_10_2660, i_10_2714, i_10_2722, i_10_2724, i_10_2725, i_10_2729, i_10_3164, i_10_3195, i_10_3196, i_10_3197, i_10_3232, i_10_3233, i_10_3277, i_10_3278, i_10_3283, i_10_3385, i_10_3389, i_10_3403, i_10_3503, i_10_3506, i_10_3524, i_10_3613, i_10_3614, i_10_3673, i_10_3686, i_10_3691, i_10_3699, i_10_3700, i_10_3727, i_10_3812, i_10_3839, i_10_3917, i_10_4010, i_10_4179, i_10_4268, i_10_4271, i_10_4459, i_10_4528, i_10_4550, i_10_4586, i_10_4591, o_10_435);
	kernel_10_436 k_10_436(i_10_64, i_10_261, i_10_286, i_10_289, i_10_290, i_10_320, i_10_323, i_10_370, i_10_432, i_10_433, i_10_442, i_10_693, i_10_736, i_10_737, i_10_756, i_10_793, i_10_800, i_10_843, i_10_844, i_10_928, i_10_948, i_10_954, i_10_1040, i_10_1045, i_10_1152, i_10_1192, i_10_1199, i_10_1200, i_10_1238, i_10_1309, i_10_1350, i_10_1354, i_10_1355, i_10_1363, i_10_1444, i_10_1555, i_10_1567, i_10_1630, i_10_1685, i_10_1741, i_10_1800, i_10_1916, i_10_1989, i_10_2205, i_10_2206, i_10_2207, i_10_2450, i_10_2467, i_10_2470, i_10_2479, i_10_2506, i_10_2509, i_10_2514, i_10_2538, i_10_2566, i_10_2569, i_10_2647, i_10_2659, i_10_2673, i_10_2674, i_10_2722, i_10_2882, i_10_3074, i_10_3107, i_10_3201, i_10_3202, i_10_3267, i_10_3268, i_10_3297, i_10_3360, i_10_3387, i_10_3389, i_10_3402, i_10_3403, i_10_3405, i_10_3408, i_10_3525, i_10_3550, i_10_3551, i_10_3553, i_10_3582, i_10_3604, i_10_3605, i_10_3611, i_10_3702, i_10_3854, i_10_3855, i_10_3859, i_10_3901, i_10_3978, i_10_3982, i_10_4185, i_10_4213, i_10_4216, i_10_4233, i_10_4278, i_10_4290, i_10_4375, i_10_4376, i_10_4500, o_10_436);
	kernel_10_437 k_10_437(i_10_30, i_10_173, i_10_254, i_10_390, i_10_407, i_10_462, i_10_465, i_10_631, i_10_633, i_10_686, i_10_732, i_10_733, i_10_736, i_10_751, i_10_792, i_10_793, i_10_795, i_10_1037, i_10_1039, i_10_1087, i_10_1234, i_10_1305, i_10_1306, i_10_1308, i_10_1310, i_10_1363, i_10_1397, i_10_1552, i_10_1714, i_10_1822, i_10_1823, i_10_1824, i_10_1881, i_10_1882, i_10_1883, i_10_1911, i_10_1925, i_10_2001, i_10_2026, i_10_2080, i_10_2093, i_10_2241, i_10_2242, i_10_2243, i_10_2263, i_10_2309, i_10_2349, i_10_2385, i_10_2451, i_10_2541, i_10_2612, i_10_2615, i_10_2628, i_10_2631, i_10_2712, i_10_2742, i_10_2979, i_10_3072, i_10_3073, i_10_3089, i_10_3096, i_10_3117, i_10_3121, i_10_3203, i_10_3232, i_10_3233, i_10_3271, i_10_3387, i_10_3465, i_10_3519, i_10_3537, i_10_3538, i_10_3539, i_10_3578, i_10_3609, i_10_3610, i_10_3645, i_10_3651, i_10_3686, i_10_3798, i_10_3823, i_10_3844, i_10_3847, i_10_3853, i_10_3859, i_10_3893, i_10_3942, i_10_3946, i_10_3997, i_10_4051, i_10_4113, i_10_4116, i_10_4122, i_10_4125, i_10_4262, i_10_4275, i_10_4285, i_10_4286, i_10_4459, i_10_4567, o_10_437);
	kernel_10_438 k_10_438(i_10_32, i_10_171, i_10_172, i_10_175, i_10_176, i_10_179, i_10_282, i_10_283, i_10_284, i_10_411, i_10_432, i_10_436, i_10_439, i_10_466, i_10_508, i_10_795, i_10_797, i_10_800, i_10_1166, i_10_1235, i_10_1237, i_10_1238, i_10_1240, i_10_1241, i_10_1296, i_10_1305, i_10_1306, i_10_1346, i_10_1445, i_10_1622, i_10_1685, i_10_1686, i_10_1687, i_10_1819, i_10_1821, i_10_1822, i_10_1823, i_10_1911, i_10_1913, i_10_1945, i_10_2033, i_10_2353, i_10_2457, i_10_2461, i_10_2466, i_10_2468, i_10_2567, i_10_2628, i_10_2629, i_10_2631, i_10_2632, i_10_2633, i_10_2635, i_10_2658, i_10_2659, i_10_2661, i_10_2662, i_10_2663, i_10_2710, i_10_2711, i_10_2714, i_10_2717, i_10_2723, i_10_2728, i_10_2830, i_10_2831, i_10_3036, i_10_3071, i_10_3197, i_10_3199, i_10_3200, i_10_3277, i_10_3278, i_10_3281, i_10_3385, i_10_3386, i_10_3389, i_10_3467, i_10_3541, i_10_3584, i_10_3587, i_10_3613, i_10_3617, i_10_3645, i_10_3647, i_10_3782, i_10_3784, i_10_3785, i_10_3837, i_10_3839, i_10_3847, i_10_3854, i_10_3856, i_10_3857, i_10_3914, i_10_4115, i_10_4123, i_10_4268, i_10_4285, i_10_4286, o_10_438);
	kernel_10_439 k_10_439(i_10_118, i_10_175, i_10_217, i_10_283, i_10_284, i_10_288, i_10_441, i_10_445, i_10_460, i_10_463, i_10_506, i_10_509, i_10_514, i_10_793, i_10_1026, i_10_1045, i_10_1082, i_10_1120, i_10_1234, i_10_1235, i_10_1237, i_10_1239, i_10_1244, i_10_1359, i_10_1361, i_10_1364, i_10_1445, i_10_1542, i_10_1577, i_10_1621, i_10_1648, i_10_1649, i_10_1650, i_10_1651, i_10_1652, i_10_1653, i_10_1691, i_10_1767, i_10_1768, i_10_1769, i_10_1800, i_10_1824, i_10_1910, i_10_2017, i_10_2232, i_10_2353, i_10_2357, i_10_2448, i_10_2449, i_10_2450, i_10_2459, i_10_2465, i_10_2473, i_10_2516, i_10_2565, i_10_2566, i_10_2630, i_10_2639, i_10_2727, i_10_2729, i_10_2782, i_10_2831, i_10_3042, i_10_3047, i_10_3088, i_10_3331, i_10_3388, i_10_3390, i_10_3406, i_10_3467, i_10_3522, i_10_3555, i_10_3556, i_10_3584, i_10_3586, i_10_3587, i_10_3618, i_10_3774, i_10_3840, i_10_3845, i_10_3847, i_10_3848, i_10_3852, i_10_3853, i_10_3980, i_10_4024, i_10_4025, i_10_4027, i_10_4028, i_10_4114, i_10_4115, i_10_4122, i_10_4123, i_10_4124, i_10_4126, i_10_4150, i_10_4175, i_10_4285, i_10_4287, i_10_4563, o_10_439);
	kernel_10_440 k_10_440(i_10_48, i_10_118, i_10_119, i_10_121, i_10_153, i_10_171, i_10_172, i_10_185, i_10_390, i_10_391, i_10_433, i_10_446, i_10_447, i_10_461, i_10_463, i_10_520, i_10_559, i_10_560, i_10_694, i_10_733, i_10_793, i_10_794, i_10_797, i_10_1085, i_10_1235, i_10_1241, i_10_1242, i_10_1361, i_10_1381, i_10_1433, i_10_1442, i_10_1444, i_10_1452, i_10_1454, i_10_1532, i_10_1579, i_10_1613, i_10_1826, i_10_1946, i_10_1949, i_10_2000, i_10_2090, i_10_2308, i_10_2309, i_10_2349, i_10_2351, i_10_2352, i_10_2405, i_10_2407, i_10_2410, i_10_2431, i_10_2454, i_10_2455, i_10_2456, i_10_2461, i_10_2471, i_10_2614, i_10_2615, i_10_2629, i_10_2630, i_10_2642, i_10_2656, i_10_2660, i_10_2674, i_10_2677, i_10_2678, i_10_2713, i_10_2723, i_10_2728, i_10_2729, i_10_2817, i_10_2818, i_10_2827, i_10_2829, i_10_2881, i_10_2884, i_10_2968, i_10_2980, i_10_3037, i_10_3313, i_10_3316, i_10_3384, i_10_3387, i_10_3391, i_10_3470, i_10_3522, i_10_3539, i_10_3586, i_10_3587, i_10_3717, i_10_3857, i_10_3947, i_10_3979, i_10_3981, i_10_3989, i_10_4120, i_10_4144, i_10_4268, i_10_4275, i_10_4276, o_10_440);
	kernel_10_441 k_10_441(i_10_67, i_10_223, i_10_445, i_10_464, i_10_466, i_10_561, i_10_593, i_10_712, i_10_736, i_10_737, i_10_934, i_10_957, i_10_999, i_10_1032, i_10_1033, i_10_1034, i_10_1039, i_10_1088, i_10_1128, i_10_1138, i_10_1139, i_10_1164, i_10_1165, i_10_1166, i_10_1233, i_10_1243, i_10_1247, i_10_1248, i_10_1250, i_10_1307, i_10_1309, i_10_1313, i_10_1365, i_10_1652, i_10_1653, i_10_1654, i_10_1823, i_10_1910, i_10_1915, i_10_1917, i_10_1920, i_10_2154, i_10_2310, i_10_2311, i_10_2352, i_10_2353, i_10_2454, i_10_2455, i_10_2512, i_10_2517, i_10_2520, i_10_2521, i_10_2619, i_10_2631, i_10_2632, i_10_2655, i_10_2659, i_10_2673, i_10_2722, i_10_2726, i_10_2831, i_10_2834, i_10_2882, i_10_2884, i_10_2953, i_10_3071, i_10_3075, i_10_3267, i_10_3269, i_10_3270, i_10_3275, i_10_3282, i_10_3390, i_10_3470, i_10_3547, i_10_3548, i_10_3583, i_10_3585, i_10_3586, i_10_3609, i_10_3648, i_10_3781, i_10_3782, i_10_3783, i_10_3784, i_10_3787, i_10_3788, i_10_3835, i_10_3838, i_10_3839, i_10_3852, i_10_3909, i_10_3943, i_10_3986, i_10_3999, i_10_4117, i_10_4118, i_10_4119, i_10_4125, i_10_4303, o_10_441);
	kernel_10_442 k_10_442(i_10_98, i_10_177, i_10_250, i_10_258, i_10_267, i_10_274, i_10_280, i_10_292, i_10_295, i_10_318, i_10_321, i_10_322, i_10_406, i_10_408, i_10_409, i_10_412, i_10_413, i_10_460, i_10_463, i_10_464, i_10_628, i_10_712, i_10_714, i_10_717, i_10_831, i_10_870, i_10_871, i_10_898, i_10_930, i_10_968, i_10_989, i_10_1033, i_10_1233, i_10_1239, i_10_1347, i_10_1363, i_10_1438, i_10_1543, i_10_1545, i_10_1546, i_10_1555, i_10_1581, i_10_1626, i_10_1633, i_10_1635, i_10_1686, i_10_1689, i_10_1806, i_10_1824, i_10_1885, i_10_1986, i_10_2031, i_10_2255, i_10_2339, i_10_2356, i_10_2364, i_10_2383, i_10_2384, i_10_2472, i_10_2514, i_10_2515, i_10_2572, i_10_2581, i_10_2608, i_10_2643, i_10_2659, i_10_2678, i_10_2712, i_10_2713, i_10_2714, i_10_2715, i_10_2716, i_10_2829, i_10_2884, i_10_2960, i_10_3072, i_10_3075, i_10_3232, i_10_3281, i_10_3283, i_10_3315, i_10_3318, i_10_3328, i_10_3337, i_10_3389, i_10_3405, i_10_3497, i_10_3507, i_10_3508, i_10_3526, i_10_3543, i_10_3650, i_10_3685, i_10_3977, i_10_4119, i_10_4120, i_10_4128, i_10_4210, i_10_4282, i_10_4585, o_10_442);
	kernel_10_443 k_10_443(i_10_120, i_10_174, i_10_180, i_10_181, i_10_256, i_10_275, i_10_319, i_10_323, i_10_387, i_10_388, i_10_390, i_10_423, i_10_426, i_10_462, i_10_495, i_10_496, i_10_507, i_10_508, i_10_1030, i_10_1035, i_10_1080, i_10_1162, i_10_1215, i_10_1216, i_10_1233, i_10_1234, i_10_1241, i_10_1359, i_10_1377, i_10_1578, i_10_1684, i_10_1689, i_10_1764, i_10_1770, i_10_1822, i_10_1825, i_10_1908, i_10_1911, i_10_1915, i_10_1989, i_10_1998, i_10_1999, i_10_2025, i_10_2179, i_10_2199, i_10_2242, i_10_2305, i_10_2359, i_10_2361, i_10_2362, i_10_2376, i_10_2379, i_10_2380, i_10_2457, i_10_2611, i_10_2636, i_10_2657, i_10_2673, i_10_2711, i_10_2727, i_10_2817, i_10_2820, i_10_2821, i_10_2919, i_10_2983, i_10_3152, i_10_3268, i_10_3270, i_10_3271, i_10_3276, i_10_3277, i_10_3279, i_10_3282, i_10_3312, i_10_3322, i_10_3387, i_10_3403, i_10_3466, i_10_3538, i_10_3540, i_10_3582, i_10_3783, i_10_3784, i_10_3785, i_10_3787, i_10_3888, i_10_3889, i_10_3978, i_10_3979, i_10_3980, i_10_4123, i_10_4167, i_10_4215, i_10_4287, i_10_4288, i_10_4289, i_10_4290, i_10_4302, i_10_4568, i_10_4569, o_10_443);
	kernel_10_444 k_10_444(i_10_176, i_10_183, i_10_223, i_10_224, i_10_249, i_10_252, i_10_282, i_10_283, i_10_391, i_10_393, i_10_408, i_10_409, i_10_446, i_10_449, i_10_515, i_10_544, i_10_597, i_10_621, i_10_689, i_10_713, i_10_715, i_10_716, i_10_753, i_10_957, i_10_958, i_10_959, i_10_962, i_10_965, i_10_983, i_10_1000, i_10_1245, i_10_1246, i_10_1248, i_10_1249, i_10_1260, i_10_1306, i_10_1307, i_10_1437, i_10_1487, i_10_1492, i_10_1493, i_10_1532, i_10_1535, i_10_1545, i_10_1581, i_10_1582, i_10_1683, i_10_1796, i_10_1823, i_10_1908, i_10_1909, i_10_1912, i_10_2031, i_10_2185, i_10_2203, i_10_2252, i_10_2254, i_10_2255, i_10_2327, i_10_2355, i_10_2362, i_10_2436, i_10_2437, i_10_2451, i_10_2465, i_10_2506, i_10_2529, i_10_2531, i_10_2535, i_10_2542, i_10_2704, i_10_2710, i_10_2731, i_10_2787, i_10_2823, i_10_2985, i_10_3036, i_10_3038, i_10_3075, i_10_3198, i_10_3202, i_10_3203, i_10_3238, i_10_3432, i_10_3588, i_10_3652, i_10_3783, i_10_3786, i_10_3847, i_10_3855, i_10_3856, i_10_3858, i_10_3912, i_10_3947, i_10_4002, i_10_4005, i_10_4011, i_10_4065, i_10_4463, i_10_4567, o_10_444);
	kernel_10_445 k_10_445(i_10_220, i_10_222, i_10_223, i_10_250, i_10_279, i_10_280, i_10_284, i_10_318, i_10_322, i_10_326, i_10_444, i_10_445, i_10_448, i_10_449, i_10_718, i_10_751, i_10_752, i_10_792, i_10_796, i_10_898, i_10_963, i_10_964, i_10_967, i_10_997, i_10_1002, i_10_1003, i_10_1084, i_10_1305, i_10_1306, i_10_1308, i_10_1437, i_10_1555, i_10_1580, i_10_1691, i_10_1768, i_10_1819, i_10_1821, i_10_1822, i_10_1823, i_10_1824, i_10_1948, i_10_2354, i_10_2362, i_10_2452, i_10_2453, i_10_2630, i_10_2632, i_10_2633, i_10_2704, i_10_2706, i_10_2707, i_10_2708, i_10_2715, i_10_2716, i_10_2717, i_10_2724, i_10_2725, i_10_2728, i_10_2734, i_10_2782, i_10_2829, i_10_2830, i_10_2919, i_10_2920, i_10_3034, i_10_3046, i_10_3076, i_10_3150, i_10_3154, i_10_3157, i_10_3389, i_10_3390, i_10_3405, i_10_3406, i_10_3468, i_10_3616, i_10_3649, i_10_3784, i_10_3787, i_10_3788, i_10_3815, i_10_3834, i_10_3842, i_10_3848, i_10_3853, i_10_3856, i_10_3888, i_10_3895, i_10_3982, i_10_3983, i_10_3985, i_10_3986, i_10_4116, i_10_4121, i_10_4266, i_10_4273, i_10_4284, i_10_4287, i_10_4290, i_10_4563, o_10_445);
	kernel_10_446 k_10_446(i_10_32, i_10_34, i_10_35, i_10_124, i_10_125, i_10_156, i_10_160, i_10_178, i_10_248, i_10_258, i_10_323, i_10_431, i_10_519, i_10_520, i_10_565, i_10_566, i_10_628, i_10_958, i_10_961, i_10_962, i_10_996, i_10_1060, i_10_1061, i_10_1070, i_10_1124, i_10_1129, i_10_1165, i_10_1268, i_10_1309, i_10_1312, i_10_1347, i_10_1546, i_10_1555, i_10_1646, i_10_1650, i_10_1651, i_10_1654, i_10_1812, i_10_1815, i_10_1816, i_10_1908, i_10_1912, i_10_1914, i_10_1916, i_10_1952, i_10_1957, i_10_1958, i_10_1961, i_10_2037, i_10_2084, i_10_2242, i_10_2276, i_10_2384, i_10_2474, i_10_2481, i_10_2516, i_10_2632, i_10_2636, i_10_2713, i_10_2722, i_10_2725, i_10_2734, i_10_2787, i_10_2806, i_10_2887, i_10_3095, i_10_3166, i_10_3201, i_10_3286, i_10_3430, i_10_3433, i_10_3542, i_10_3616, i_10_3650, i_10_3651, i_10_3653, i_10_3704, i_10_3705, i_10_3718, i_10_3886, i_10_3887, i_10_3913, i_10_3984, i_10_3985, i_10_3991, i_10_3992, i_10_3994, i_10_3995, i_10_4053, i_10_4054, i_10_4057, i_10_4058, i_10_4118, i_10_4126, i_10_4129, i_10_4237, i_10_4271, i_10_4283, i_10_4400, i_10_4569, o_10_446);
	kernel_10_447 k_10_447(i_10_88, i_10_89, i_10_176, i_10_219, i_10_224, i_10_295, i_10_391, i_10_395, i_10_408, i_10_431, i_10_436, i_10_439, i_10_440, i_10_463, i_10_464, i_10_500, i_10_511, i_10_695, i_10_698, i_10_853, i_10_854, i_10_948, i_10_1027, i_10_1043, i_10_1056, i_10_1176, i_10_1238, i_10_1240, i_10_1245, i_10_1321, i_10_1345, i_10_1346, i_10_1448, i_10_1527, i_10_1552, i_10_1577, i_10_1649, i_10_1733, i_10_1735, i_10_1736, i_10_1804, i_10_1807, i_10_1888, i_10_2310, i_10_2312, i_10_2365, i_10_2374, i_10_2375, i_10_2451, i_10_2540, i_10_2543, i_10_2558, i_10_2561, i_10_2631, i_10_2632, i_10_2636, i_10_2645, i_10_2696, i_10_2714, i_10_2716, i_10_2733, i_10_2821, i_10_2852, i_10_2882, i_10_2885, i_10_2919, i_10_3197, i_10_3271, i_10_3278, i_10_3318, i_10_3319, i_10_3329, i_10_3356, i_10_3364, i_10_3390, i_10_3391, i_10_3406, i_10_3409, i_10_3463, i_10_3473, i_10_3499, i_10_3526, i_10_3620, i_10_3705, i_10_3706, i_10_3725, i_10_3839, i_10_3841, i_10_3854, i_10_3893, i_10_4031, i_10_4090, i_10_4115, i_10_4118, i_10_4129, i_10_4188, i_10_4277, i_10_4307, i_10_4564, i_10_4585, o_10_447);
	kernel_10_448 k_10_448(i_10_83, i_10_117, i_10_152, i_10_176, i_10_182, i_10_217, i_10_279, i_10_406, i_10_408, i_10_443, i_10_445, i_10_446, i_10_460, i_10_461, i_10_463, i_10_464, i_10_509, i_10_515, i_10_686, i_10_747, i_10_754, i_10_794, i_10_795, i_10_967, i_10_1163, i_10_1212, i_10_1235, i_10_1237, i_10_1243, i_10_1244, i_10_1312, i_10_1361, i_10_1378, i_10_1487, i_10_1537, i_10_1562, i_10_1647, i_10_1651, i_10_1652, i_10_1684, i_10_1685, i_10_1688, i_10_1690, i_10_1768, i_10_1784, i_10_1808, i_10_1821, i_10_1822, i_10_1823, i_10_1824, i_10_1937, i_10_2033, i_10_2252, i_10_2391, i_10_2468, i_10_2509, i_10_2512, i_10_2631, i_10_2702, i_10_2716, i_10_2722, i_10_2723, i_10_2725, i_10_2726, i_10_2728, i_10_2731, i_10_2734, i_10_2735, i_10_2833, i_10_2916, i_10_2917, i_10_2920, i_10_2954, i_10_3034, i_10_3268, i_10_3326, i_10_3384, i_10_3524, i_10_3541, i_10_3586, i_10_3587, i_10_3645, i_10_3685, i_10_3797, i_10_3846, i_10_3847, i_10_3854, i_10_3859, i_10_3870, i_10_3880, i_10_3916, i_10_3961, i_10_4117, i_10_4118, i_10_4119, i_10_4140, i_10_4268, i_10_4285, i_10_4286, i_10_4288, o_10_448);
	kernel_10_449 k_10_449(i_10_124, i_10_184, i_10_224, i_10_247, i_10_286, i_10_318, i_10_408, i_10_410, i_10_429, i_10_440, i_10_446, i_10_462, i_10_463, i_10_464, i_10_466, i_10_467, i_10_508, i_10_564, i_10_796, i_10_1005, i_10_1006, i_10_1033, i_10_1042, i_10_1043, i_10_1137, i_10_1138, i_10_1139, i_10_1236, i_10_1237, i_10_1239, i_10_1307, i_10_1308, i_10_1313, i_10_1366, i_10_1383, i_10_1384, i_10_1437, i_10_1653, i_10_1655, i_10_1821, i_10_1824, i_10_1909, i_10_1912, i_10_1913, i_10_1950, i_10_2094, i_10_2095, i_10_2350, i_10_2352, i_10_2356, i_10_2383, i_10_2384, i_10_2438, i_10_2471, i_10_2508, i_10_2514, i_10_2628, i_10_2631, i_10_2632, i_10_2634, i_10_2636, i_10_2655, i_10_2656, i_10_2660, i_10_2724, i_10_2829, i_10_2830, i_10_2831, i_10_2922, i_10_3039, i_10_3040, i_10_3154, i_10_3195, i_10_3197, i_10_3198, i_10_3199, i_10_3613, i_10_3614, i_10_3645, i_10_3649, i_10_3651, i_10_3652, i_10_3784, i_10_3788, i_10_3838, i_10_3847, i_10_3852, i_10_3853, i_10_3856, i_10_3895, i_10_3896, i_10_3967, i_10_4056, i_10_4117, i_10_4118, i_10_4120, i_10_4129, i_10_4278, i_10_4533, i_10_4567, o_10_449);
	kernel_10_450 k_10_450(i_10_250, i_10_251, i_10_282, i_10_331, i_10_411, i_10_412, i_10_447, i_10_511, i_10_597, i_10_794, i_10_795, i_10_1030, i_10_1080, i_10_1083, i_10_1138, i_10_1139, i_10_1142, i_10_1236, i_10_1240, i_10_1243, i_10_1305, i_10_1306, i_10_1308, i_10_1309, i_10_1310, i_10_1312, i_10_1365, i_10_1367, i_10_1444, i_10_1653, i_10_1687, i_10_1688, i_10_1767, i_10_1818, i_10_1913, i_10_2158, i_10_2403, i_10_2406, i_10_2407, i_10_2408, i_10_2454, i_10_2455, i_10_2456, i_10_2479, i_10_2518, i_10_2604, i_10_2632, i_10_2634, i_10_2636, i_10_2658, i_10_2659, i_10_2660, i_10_2679, i_10_2680, i_10_2681, i_10_2703, i_10_2726, i_10_2732, i_10_2783, i_10_2784, i_10_2785, i_10_2787, i_10_2788, i_10_2831, i_10_2919, i_10_3049, i_10_3150, i_10_3154, i_10_3277, i_10_3280, i_10_3283, i_10_3385, i_10_3387, i_10_3388, i_10_3389, i_10_3391, i_10_3392, i_10_3406, i_10_3494, i_10_3613, i_10_3650, i_10_3652, i_10_3785, i_10_3835, i_10_3839, i_10_3841, i_10_3855, i_10_3856, i_10_3981, i_10_4029, i_10_4054, i_10_4055, i_10_4056, i_10_4057, i_10_4270, i_10_4284, i_10_4285, i_10_4288, i_10_4292, i_10_4565, o_10_450);
	kernel_10_451 k_10_451(i_10_12, i_10_174, i_10_177, i_10_253, i_10_256, i_10_261, i_10_264, i_10_265, i_10_285, i_10_286, i_10_318, i_10_391, i_10_444, i_10_460, i_10_504, i_10_792, i_10_867, i_10_999, i_10_1002, i_10_1029, i_10_1056, i_10_1101, i_10_1104, i_10_1296, i_10_1299, i_10_1302, i_10_1344, i_10_1347, i_10_1431, i_10_1434, i_10_1542, i_10_1543, i_10_1545, i_10_1546, i_10_1575, i_10_1620, i_10_1623, i_10_1649, i_10_1683, i_10_1686, i_10_1729, i_10_1731, i_10_1819, i_10_1824, i_10_1980, i_10_2016, i_10_2028, i_10_2202, i_10_2349, i_10_2352, i_10_2529, i_10_2532, i_10_2565, i_10_2568, i_10_2677, i_10_2678, i_10_2703, i_10_2743, i_10_2820, i_10_2847, i_10_2881, i_10_2883, i_10_2967, i_10_3045, i_10_3072, i_10_3267, i_10_3277, i_10_3280, i_10_3281, i_10_3312, i_10_3390, i_10_3391, i_10_3471, i_10_3473, i_10_3537, i_10_3540, i_10_3541, i_10_3543, i_10_3544, i_10_3582, i_10_3585, i_10_3621, i_10_3652, i_10_3687, i_10_3795, i_10_3834, i_10_3837, i_10_3842, i_10_3847, i_10_3850, i_10_4116, i_10_4117, i_10_4167, i_10_4170, i_10_4275, i_10_4281, i_10_4287, i_10_4290, i_10_4563, i_10_4585, o_10_451);
	kernel_10_452 k_10_452(i_10_31, i_10_33, i_10_67, i_10_171, i_10_184, i_10_212, i_10_283, i_10_390, i_10_391, i_10_405, i_10_406, i_10_435, i_10_436, i_10_439, i_10_514, i_10_718, i_10_750, i_10_1002, i_10_1030, i_10_1035, i_10_1038, i_10_1056, i_10_1164, i_10_1261, i_10_1262, i_10_1264, i_10_1287, i_10_1305, i_10_1351, i_10_1362, i_10_1363, i_10_1364, i_10_1366, i_10_1367, i_10_1435, i_10_1542, i_10_1554, i_10_1606, i_10_1635, i_10_1768, i_10_1804, i_10_1825, i_10_1872, i_10_1913, i_10_2041, i_10_2091, i_10_2143, i_10_2196, i_10_2356, i_10_2374, i_10_2407, i_10_2448, i_10_2453, i_10_2470, i_10_2512, i_10_2514, i_10_2526, i_10_2605, i_10_2700, i_10_2722, i_10_2734, i_10_2754, i_10_2785, i_10_2820, i_10_2821, i_10_2957, i_10_2982, i_10_2983, i_10_3033, i_10_3036, i_10_3046, i_10_3234, i_10_3237, i_10_3268, i_10_3271, i_10_3319, i_10_3390, i_10_3393, i_10_3586, i_10_3652, i_10_3653, i_10_3663, i_10_3702, i_10_3717, i_10_3718, i_10_3719, i_10_3834, i_10_3835, i_10_3853, i_10_3856, i_10_3982, i_10_4053, i_10_4174, i_10_4276, i_10_4278, i_10_4373, i_10_4485, i_10_4528, i_10_4534, i_10_4569, o_10_452);
	kernel_10_453 k_10_453(i_10_70, i_10_180, i_10_181, i_10_281, i_10_282, i_10_372, i_10_407, i_10_429, i_10_430, i_10_441, i_10_442, i_10_443, i_10_444, i_10_461, i_10_464, i_10_520, i_10_536, i_10_590, i_10_629, i_10_735, i_10_797, i_10_826, i_10_967, i_10_1238, i_10_1243, i_10_1263, i_10_1309, i_10_1321, i_10_1359, i_10_1581, i_10_1616, i_10_1691, i_10_1755, i_10_1757, i_10_1805, i_10_1821, i_10_1823, i_10_1912, i_10_1913, i_10_2083, i_10_2087, i_10_2159, i_10_2184, i_10_2229, i_10_2312, i_10_2326, i_10_2327, i_10_2350, i_10_2408, i_10_2440, i_10_2449, i_10_2453, i_10_2455, i_10_2456, i_10_2471, i_10_2635, i_10_2636, i_10_2662, i_10_2663, i_10_2701, i_10_2704, i_10_2725, i_10_2728, i_10_2729, i_10_2731, i_10_2831, i_10_2862, i_10_2886, i_10_3035, i_10_3093, i_10_3094, i_10_3202, i_10_3234, i_10_3277, i_10_3405, i_10_3409, i_10_3526, i_10_3527, i_10_3688, i_10_3782, i_10_3859, i_10_3949, i_10_3980, i_10_3981, i_10_3982, i_10_4120, i_10_4182, i_10_4185, i_10_4189, i_10_4190, i_10_4267, i_10_4269, i_10_4270, i_10_4271, i_10_4274, i_10_4287, i_10_4458, i_10_4549, i_10_4550, i_10_4571, o_10_453);
	kernel_10_454 k_10_454(i_10_171, i_10_172, i_10_173, i_10_175, i_10_176, i_10_283, i_10_285, i_10_320, i_10_321, i_10_405, i_10_407, i_10_433, i_10_435, i_10_443, i_10_444, i_10_445, i_10_461, i_10_466, i_10_467, i_10_505, i_10_518, i_10_718, i_10_719, i_10_960, i_10_962, i_10_967, i_10_968, i_10_1233, i_10_1236, i_10_1237, i_10_1240, i_10_1250, i_10_1306, i_10_1310, i_10_1311, i_10_1579, i_10_1581, i_10_1653, i_10_1654, i_10_1688, i_10_1817, i_10_1818, i_10_1819, i_10_1823, i_10_1825, i_10_2203, i_10_2332, i_10_2338, i_10_2350, i_10_2363, i_10_2377, i_10_2380, i_10_2383, i_10_2461, i_10_2462, i_10_2471, i_10_2633, i_10_2636, i_10_2658, i_10_2659, i_10_2660, i_10_2700, i_10_2708, i_10_2724, i_10_2731, i_10_2735, i_10_2881, i_10_2920, i_10_2921, i_10_3152, i_10_3154, i_10_3322, i_10_3325, i_10_3385, i_10_3469, i_10_3472, i_10_3497, i_10_3586, i_10_3612, i_10_3613, i_10_3616, i_10_3782, i_10_3783, i_10_3847, i_10_3848, i_10_3853, i_10_3854, i_10_3986, i_10_4117, i_10_4174, i_10_4267, i_10_4268, i_10_4270, i_10_4271, i_10_4285, i_10_4286, i_10_4564, i_10_4566, i_10_4567, i_10_4568, o_10_454);
	kernel_10_455 k_10_455(i_10_246, i_10_249, i_10_273, i_10_276, i_10_289, i_10_294, i_10_295, i_10_324, i_10_328, i_10_330, i_10_438, i_10_459, i_10_462, i_10_463, i_10_464, i_10_465, i_10_531, i_10_534, i_10_993, i_10_996, i_10_1000, i_10_1038, i_10_1039, i_10_1041, i_10_1238, i_10_1240, i_10_1241, i_10_1267, i_10_1308, i_10_1312, i_10_1344, i_10_1350, i_10_1435, i_10_1441, i_10_1443, i_10_1446, i_10_1488, i_10_1546, i_10_1648, i_10_1683, i_10_1689, i_10_1713, i_10_1818, i_10_1872, i_10_1946, i_10_2250, i_10_2322, i_10_2325, i_10_2349, i_10_2351, i_10_2361, i_10_2364, i_10_2377, i_10_2460, i_10_2469, i_10_2505, i_10_2607, i_10_2634, i_10_2636, i_10_2658, i_10_2661, i_10_2676, i_10_2703, i_10_2706, i_10_2715, i_10_2721, i_10_2724, i_10_2730, i_10_2781, i_10_2806, i_10_2829, i_10_2831, i_10_2832, i_10_2834, i_10_2881, i_10_2918, i_10_3036, i_10_3037, i_10_3039, i_10_3045, i_10_3153, i_10_3165, i_10_3274, i_10_3281, i_10_3291, i_10_3403, i_10_3408, i_10_3492, i_10_3609, i_10_3610, i_10_3616, i_10_3617, i_10_3849, i_10_3982, i_10_3994, i_10_4028, i_10_4128, i_10_4291, i_10_4564, i_10_4568, o_10_455);
	kernel_10_456 k_10_456(i_10_221, i_10_224, i_10_319, i_10_320, i_10_322, i_10_323, i_10_329, i_10_436, i_10_447, i_10_465, i_10_466, i_10_508, i_10_898, i_10_1004, i_10_1005, i_10_1083, i_10_1084, i_10_1085, i_10_1086, i_10_1087, i_10_1088, i_10_1240, i_10_1241, i_10_1242, i_10_1246, i_10_1249, i_10_1263, i_10_1309, i_10_1313, i_10_1651, i_10_1652, i_10_2352, i_10_2382, i_10_2407, i_10_2470, i_10_2509, i_10_2510, i_10_2629, i_10_2661, i_10_2700, i_10_2701, i_10_2703, i_10_2704, i_10_2706, i_10_2707, i_10_2711, i_10_2726, i_10_2782, i_10_2783, i_10_2785, i_10_2786, i_10_2789, i_10_2885, i_10_2919, i_10_2920, i_10_2922, i_10_2923, i_10_2924, i_10_2959, i_10_2987, i_10_3153, i_10_3279, i_10_3281, i_10_3385, i_10_3389, i_10_3391, i_10_3406, i_10_3407, i_10_3408, i_10_3409, i_10_3472, i_10_3496, i_10_3497, i_10_3586, i_10_3616, i_10_3646, i_10_3649, i_10_3650, i_10_3653, i_10_3784, i_10_3786, i_10_3788, i_10_3847, i_10_3848, i_10_3854, i_10_3860, i_10_3978, i_10_3979, i_10_3980, i_10_3983, i_10_3985, i_10_3986, i_10_4057, i_10_4113, i_10_4128, i_10_4130, i_10_4236, i_10_4237, i_10_4288, i_10_4289, o_10_456);
	kernel_10_457 k_10_457(i_10_174, i_10_247, i_10_248, i_10_265, i_10_269, i_10_285, i_10_286, i_10_394, i_10_395, i_10_431, i_10_436, i_10_449, i_10_565, i_10_800, i_10_966, i_10_1006, i_10_1007, i_10_1084, i_10_1138, i_10_1237, i_10_1248, i_10_1303, i_10_1306, i_10_1308, i_10_1309, i_10_1310, i_10_1366, i_10_1435, i_10_1438, i_10_1439, i_10_1556, i_10_1654, i_10_1655, i_10_1717, i_10_1821, i_10_1822, i_10_1824, i_10_1825, i_10_1826, i_10_1913, i_10_1996, i_10_2006, i_10_2351, i_10_2352, i_10_2452, i_10_2474, i_10_2608, i_10_2614, i_10_2618, i_10_2631, i_10_2654, i_10_2660, i_10_2703, i_10_2706, i_10_2707, i_10_2722, i_10_2725, i_10_2730, i_10_2731, i_10_2732, i_10_2785, i_10_2824, i_10_2825, i_10_2830, i_10_2885, i_10_2920, i_10_2923, i_10_2924, i_10_3093, i_10_3094, i_10_3095, i_10_3156, i_10_3202, i_10_3277, i_10_3281, i_10_3282, i_10_3283, i_10_3284, i_10_3322, i_10_3473, i_10_3543, i_10_3587, i_10_3612, i_10_3614, i_10_3783, i_10_3837, i_10_3855, i_10_3857, i_10_3858, i_10_3986, i_10_3991, i_10_4114, i_10_4117, i_10_4118, i_10_4119, i_10_4120, i_10_4121, i_10_4566, i_10_4567, i_10_4568, o_10_457);
	kernel_10_458 k_10_458(i_10_204, i_10_273, i_10_275, i_10_279, i_10_343, i_10_366, i_10_371, i_10_385, i_10_406, i_10_459, i_10_460, i_10_496, i_10_500, i_10_696, i_10_699, i_10_731, i_10_818, i_10_903, i_10_904, i_10_906, i_10_930, i_10_1030, i_10_1113, i_10_1166, i_10_1193, i_10_1221, i_10_1277, i_10_1282, i_10_1283, i_10_1305, i_10_1306, i_10_1360, i_10_1361, i_10_1365, i_10_1366, i_10_1371, i_10_1488, i_10_1548, i_10_1551, i_10_1641, i_10_1743, i_10_1909, i_10_1914, i_10_1933, i_10_1979, i_10_2154, i_10_2271, i_10_2272, i_10_2354, i_10_2376, i_10_2381, i_10_2448, i_10_2505, i_10_2625, i_10_2703, i_10_2707, i_10_2727, i_10_2730, i_10_2854, i_10_2857, i_10_2917, i_10_2941, i_10_2952, i_10_2955, i_10_3099, i_10_3100, i_10_3103, i_10_3190, i_10_3208, i_10_3209, i_10_3233, i_10_3236, i_10_3334, i_10_3362, i_10_3540, i_10_3541, i_10_3649, i_10_3666, i_10_3722, i_10_3837, i_10_3852, i_10_3860, i_10_3885, i_10_3919, i_10_4182, i_10_4186, i_10_4273, i_10_4359, i_10_4361, i_10_4369, i_10_4381, i_10_4428, i_10_4429, i_10_4430, i_10_4462, i_10_4523, i_10_4574, i_10_4590, i_10_4591, i_10_4592, o_10_458);
	kernel_10_459 k_10_459(i_10_172, i_10_173, i_10_175, i_10_244, i_10_286, i_10_287, i_10_316, i_10_317, i_10_329, i_10_406, i_10_407, i_10_461, i_10_515, i_10_694, i_10_695, i_10_748, i_10_958, i_10_1028, i_10_1081, i_10_1234, i_10_1235, i_10_1237, i_10_1238, i_10_1244, i_10_1249, i_10_1265, i_10_1306, i_10_1343, i_10_1541, i_10_1549, i_10_1550, i_10_1576, i_10_1819, i_10_2018, i_10_2027, i_10_2080, i_10_2201, i_10_2305, i_10_2306, i_10_2350, i_10_2351, i_10_2357, i_10_2361, i_10_2431, i_10_2432, i_10_2452, i_10_2466, i_10_2471, i_10_2601, i_10_2629, i_10_2630, i_10_2633, i_10_2661, i_10_2662, i_10_2710, i_10_2730, i_10_2731, i_10_2783, i_10_2786, i_10_2818, i_10_2819, i_10_2829, i_10_2884, i_10_2885, i_10_2917, i_10_2918, i_10_2953, i_10_2980, i_10_2981, i_10_3042, i_10_3154, i_10_3323, i_10_3385, i_10_3388, i_10_3389, i_10_3407, i_10_3526, i_10_3556, i_10_3583, i_10_3586, i_10_3613, i_10_3614, i_10_3843, i_10_3847, i_10_3848, i_10_3852, i_10_3853, i_10_3858, i_10_3888, i_10_3889, i_10_3890, i_10_3908, i_10_3980, i_10_3981, i_10_4120, i_10_4127, i_10_4271, i_10_4277, i_10_4285, i_10_4564, o_10_459);
	kernel_10_460 k_10_460(i_10_125, i_10_268, i_10_269, i_10_283, i_10_286, i_10_319, i_10_320, i_10_392, i_10_395, i_10_441, i_10_466, i_10_539, i_10_581, i_10_754, i_10_795, i_10_953, i_10_1004, i_10_1006, i_10_1007, i_10_1205, i_10_1308, i_10_1312, i_10_1345, i_10_1552, i_10_1577, i_10_1616, i_10_1618, i_10_1619, i_10_1648, i_10_1650, i_10_1651, i_10_1686, i_10_1697, i_10_1824, i_10_2158, i_10_2159, i_10_2310, i_10_2311, i_10_2312, i_10_2336, i_10_2339, i_10_2354, i_10_2357, i_10_2405, i_10_2407, i_10_2408, i_10_2410, i_10_2447, i_10_2455, i_10_2463, i_10_2519, i_10_2536, i_10_2618, i_10_2629, i_10_2632, i_10_2633, i_10_2635, i_10_2636, i_10_2705, i_10_2734, i_10_2788, i_10_2826, i_10_2884, i_10_2885, i_10_2987, i_10_3058, i_10_3070, i_10_3199, i_10_3200, i_10_3329, i_10_3365, i_10_3387, i_10_3391, i_10_3392, i_10_3437, i_10_3587, i_10_3623, i_10_3645, i_10_3650, i_10_3653, i_10_3707, i_10_3733, i_10_3734, i_10_3781, i_10_3838, i_10_3839, i_10_3884, i_10_3986, i_10_4058, i_10_4094, i_10_4115, i_10_4120, i_10_4184, i_10_4266, i_10_4268, i_10_4274, i_10_4382, i_10_4460, i_10_4534, i_10_4567, o_10_460);
	kernel_10_461 k_10_461(i_10_39, i_10_149, i_10_154, i_10_243, i_10_247, i_10_263, i_10_290, i_10_315, i_10_317, i_10_318, i_10_319, i_10_321, i_10_387, i_10_409, i_10_423, i_10_445, i_10_460, i_10_462, i_10_500, i_10_503, i_10_521, i_10_639, i_10_671, i_10_752, i_10_891, i_10_1080, i_10_1237, i_10_1241, i_10_1270, i_10_1297, i_10_1345, i_10_1432, i_10_1433, i_10_1442, i_10_1535, i_10_1541, i_10_1544, i_10_1546, i_10_1596, i_10_1634, i_10_1643, i_10_1651, i_10_1654, i_10_1684, i_10_1690, i_10_1810, i_10_1821, i_10_1918, i_10_1989, i_10_2000, i_10_2003, i_10_2017, i_10_2018, i_10_2029, i_10_2030, i_10_2033, i_10_2107, i_10_2108, i_10_2235, i_10_2262, i_10_2312, i_10_2345, i_10_2348, i_10_2358, i_10_2361, i_10_2362, i_10_2384, i_10_2448, i_10_2449, i_10_2454, i_10_2465, i_10_2566, i_10_2567, i_10_2601, i_10_2635, i_10_2705, i_10_2785, i_10_2820, i_10_2822, i_10_2915, i_10_3044, i_10_3070, i_10_3165, i_10_3279, i_10_3317, i_10_3320, i_10_3335, i_10_3430, i_10_3467, i_10_3494, i_10_3557, i_10_3560, i_10_3794, i_10_3841, i_10_3881, i_10_3914, i_10_4118, i_10_4271, i_10_4274, i_10_4583, o_10_461);
	kernel_10_462 k_10_462(i_10_40, i_10_83, i_10_172, i_10_282, i_10_289, i_10_445, i_10_460, i_10_461, i_10_463, i_10_464, i_10_466, i_10_504, i_10_715, i_10_799, i_10_892, i_10_967, i_10_1000, i_10_1042, i_10_1135, i_10_1233, i_10_1234, i_10_1235, i_10_1241, i_10_1243, i_10_1344, i_10_1359, i_10_1360, i_10_1361, i_10_1363, i_10_1364, i_10_1367, i_10_1441, i_10_1444, i_10_1540, i_10_1543, i_10_1549, i_10_1576, i_10_1577, i_10_1578, i_10_1580, i_10_1650, i_10_1678, i_10_1767, i_10_1818, i_10_1819, i_10_1823, i_10_1908, i_10_1909, i_10_1911, i_10_2182, i_10_2352, i_10_2357, i_10_2382, i_10_2455, i_10_2470, i_10_2648, i_10_2655, i_10_2657, i_10_2673, i_10_2709, i_10_2710, i_10_2718, i_10_2727, i_10_2728, i_10_2729, i_10_2826, i_10_2827, i_10_2829, i_10_2882, i_10_2917, i_10_2918, i_10_2919, i_10_2920, i_10_3035, i_10_3042, i_10_3231, i_10_3271, i_10_3321, i_10_3322, i_10_3324, i_10_3325, i_10_3384, i_10_3385, i_10_3389, i_10_3523, i_10_3550, i_10_3585, i_10_3586, i_10_3645, i_10_3781, i_10_3846, i_10_3848, i_10_3854, i_10_3979, i_10_3980, i_10_4284, i_10_4285, i_10_4286, i_10_4290, i_10_4565, o_10_462);
	kernel_10_463 k_10_463(i_10_243, i_10_252, i_10_263, i_10_286, i_10_317, i_10_319, i_10_320, i_10_395, i_10_512, i_10_621, i_10_687, i_10_688, i_10_865, i_10_1001, i_10_1003, i_10_1004, i_10_1058, i_10_1081, i_10_1084, i_10_1134, i_10_1135, i_10_1152, i_10_1153, i_10_1223, i_10_1237, i_10_1263, i_10_1300, i_10_1435, i_10_1436, i_10_1530, i_10_1535, i_10_1548, i_10_1551, i_10_1552, i_10_1580, i_10_1625, i_10_1628, i_10_1730, i_10_1733, i_10_1808, i_10_1810, i_10_1821, i_10_1906, i_10_1915, i_10_2020, i_10_2030, i_10_2033, i_10_2064, i_10_2111, i_10_2200, i_10_2340, i_10_2345, i_10_2349, i_10_2352, i_10_2353, i_10_2363, i_10_2380, i_10_2406, i_10_2453, i_10_2468, i_10_2567, i_10_2570, i_10_2703, i_10_2731, i_10_2732, i_10_2741, i_10_2744, i_10_2782, i_10_2808, i_10_2839, i_10_2840, i_10_3043, i_10_3047, i_10_3091, i_10_3195, i_10_3202, i_10_3271, i_10_3317, i_10_3320, i_10_3335, i_10_3353, i_10_3393, i_10_3473, i_10_3545, i_10_3560, i_10_3612, i_10_3663, i_10_3789, i_10_3842, i_10_3911, i_10_3942, i_10_3946, i_10_3999, i_10_4031, i_10_4117, i_10_4127, i_10_4274, i_10_4280, i_10_4365, i_10_4585, o_10_463);
	kernel_10_464 k_10_464(i_10_153, i_10_172, i_10_285, i_10_315, i_10_387, i_10_393, i_10_410, i_10_423, i_10_433, i_10_910, i_10_946, i_10_958, i_10_966, i_10_1038, i_10_1051, i_10_1209, i_10_1240, i_10_1241, i_10_1262, i_10_1307, i_10_1580, i_10_1614, i_10_1630, i_10_1683, i_10_1684, i_10_1685, i_10_1688, i_10_1747, i_10_1819, i_10_1820, i_10_1822, i_10_1825, i_10_1826, i_10_1893, i_10_1954, i_10_2018, i_10_2178, i_10_2182, i_10_2244, i_10_2287, i_10_2291, i_10_2365, i_10_2380, i_10_2382, i_10_2385, i_10_2386, i_10_2461, i_10_2513, i_10_2565, i_10_2566, i_10_2569, i_10_2587, i_10_2660, i_10_2701, i_10_2712, i_10_2718, i_10_2719, i_10_2724, i_10_2728, i_10_2731, i_10_2732, i_10_2743, i_10_2834, i_10_2843, i_10_2866, i_10_2867, i_10_2882, i_10_2920, i_10_2979, i_10_2982, i_10_3042, i_10_3047, i_10_3089, i_10_3100, i_10_3166, i_10_3199, i_10_3202, i_10_3415, i_10_3465, i_10_3540, i_10_3610, i_10_3613, i_10_3652, i_10_3686, i_10_3799, i_10_3800, i_10_3820, i_10_3836, i_10_3839, i_10_3852, i_10_3988, i_10_4053, i_10_4144, i_10_4192, i_10_4270, i_10_4271, i_10_4275, i_10_4283, i_10_4308, i_10_4451, o_10_464);
	kernel_10_465 k_10_465(i_10_121, i_10_152, i_10_176, i_10_186, i_10_187, i_10_222, i_10_224, i_10_318, i_10_441, i_10_446, i_10_449, i_10_460, i_10_463, i_10_464, i_10_466, i_10_467, i_10_510, i_10_717, i_10_797, i_10_800, i_10_908, i_10_968, i_10_1040, i_10_1247, i_10_1250, i_10_1542, i_10_1543, i_10_1578, i_10_1579, i_10_1652, i_10_1653, i_10_1685, i_10_1822, i_10_1823, i_10_1824, i_10_1826, i_10_1912, i_10_1952, i_10_1995, i_10_2004, i_10_2005, i_10_2006, i_10_2095, i_10_2182, i_10_2203, i_10_2364, i_10_2379, i_10_2380, i_10_2381, i_10_2384, i_10_2453, i_10_2456, i_10_2471, i_10_2473, i_10_2474, i_10_2628, i_10_2633, i_10_2700, i_10_2703, i_10_2715, i_10_2717, i_10_2734, i_10_2782, i_10_2830, i_10_2833, i_10_2834, i_10_2886, i_10_3034, i_10_3035, i_10_3037, i_10_3038, i_10_3040, i_10_3041, i_10_3076, i_10_3155, i_10_3199, i_10_3200, i_10_3269, i_10_3270, i_10_3271, i_10_3274, i_10_3387, i_10_3389, i_10_3406, i_10_3587, i_10_3589, i_10_3590, i_10_3615, i_10_3650, i_10_3651, i_10_3787, i_10_3788, i_10_3837, i_10_3860, i_10_4121, i_10_4175, i_10_4286, i_10_4288, i_10_4291, i_10_4568, o_10_465);
	kernel_10_466 k_10_466(i_10_217, i_10_220, i_10_221, i_10_280, i_10_281, i_10_282, i_10_283, i_10_284, i_10_316, i_10_324, i_10_390, i_10_391, i_10_406, i_10_443, i_10_445, i_10_449, i_10_459, i_10_464, i_10_505, i_10_506, i_10_509, i_10_749, i_10_797, i_10_1135, i_10_1233, i_10_1236, i_10_1250, i_10_1305, i_10_1345, i_10_1346, i_10_1431, i_10_1432, i_10_1433, i_10_1540, i_10_1552, i_10_1621, i_10_1651, i_10_1654, i_10_1683, i_10_1689, i_10_1824, i_10_1825, i_10_1981, i_10_1990, i_10_2017, i_10_2351, i_10_2359, i_10_2380, i_10_2407, i_10_2451, i_10_2628, i_10_2629, i_10_2630, i_10_2631, i_10_2632, i_10_2656, i_10_2701, i_10_2709, i_10_2710, i_10_2718, i_10_2723, i_10_2884, i_10_2917, i_10_2979, i_10_3044, i_10_3070, i_10_3152, i_10_3153, i_10_3156, i_10_3196, i_10_3277, i_10_3278, i_10_3281, i_10_3385, i_10_3388, i_10_3389, i_10_3391, i_10_3392, i_10_3523, i_10_3556, i_10_3728, i_10_3784, i_10_3834, i_10_3837, i_10_3846, i_10_3859, i_10_3979, i_10_3985, i_10_3991, i_10_4114, i_10_4115, i_10_4116, i_10_4117, i_10_4118, i_10_4122, i_10_4168, i_10_4276, i_10_4566, i_10_4567, i_10_4568, o_10_466);
	kernel_10_467 k_10_467(i_10_176, i_10_254, i_10_263, i_10_266, i_10_272, i_10_323, i_10_407, i_10_412, i_10_445, i_10_500, i_10_502, i_10_506, i_10_509, i_10_563, i_10_595, i_10_877, i_10_1003, i_10_1028, i_10_1109, i_10_1111, i_10_1112, i_10_1220, i_10_1235, i_10_1239, i_10_1246, i_10_1283, i_10_1300, i_10_1303, i_10_1360, i_10_1436, i_10_1451, i_10_1454, i_10_1541, i_10_1544, i_10_1546, i_10_1580, i_10_1583, i_10_1622, i_10_1625, i_10_1688, i_10_1733, i_10_1808, i_10_1824, i_10_1982, i_10_2003, i_10_2006, i_10_2027, i_10_2108, i_10_2204, i_10_2351, i_10_2361, i_10_2364, i_10_2467, i_10_2533, i_10_2534, i_10_2567, i_10_2570, i_10_2609, i_10_2658, i_10_2705, i_10_2722, i_10_2731, i_10_2789, i_10_2830, i_10_2833, i_10_2837, i_10_2867, i_10_2923, i_10_3034, i_10_3041, i_10_3314, i_10_3316, i_10_3317, i_10_3332, i_10_3350, i_10_3391, i_10_3392, i_10_3402, i_10_3443, i_10_3466, i_10_3583, i_10_3587, i_10_3797, i_10_3835, i_10_3836, i_10_3842, i_10_3848, i_10_3983, i_10_4010, i_10_4126, i_10_4127, i_10_4130, i_10_4154, i_10_4171, i_10_4268, i_10_4288, i_10_4379, i_10_4550, i_10_4565, i_10_4568, o_10_467);
	kernel_10_468 k_10_468(i_10_89, i_10_171, i_10_176, i_10_224, i_10_277, i_10_281, i_10_409, i_10_443, i_10_446, i_10_459, i_10_507, i_10_796, i_10_797, i_10_955, i_10_1034, i_10_1236, i_10_1244, i_10_1247, i_10_1248, i_10_1250, i_10_1343, i_10_1445, i_10_1540, i_10_1544, i_10_1554, i_10_1577, i_10_1580, i_10_1650, i_10_1678, i_10_1686, i_10_1688, i_10_1821, i_10_1822, i_10_1823, i_10_2197, i_10_2201, i_10_2407, i_10_2410, i_10_2452, i_10_2453, i_10_2469, i_10_2470, i_10_2472, i_10_2473, i_10_2474, i_10_2513, i_10_2530, i_10_2656, i_10_2657, i_10_2659, i_10_2660, i_10_2718, i_10_2719, i_10_2732, i_10_2828, i_10_2830, i_10_2831, i_10_2834, i_10_2863, i_10_2920, i_10_2921, i_10_2923, i_10_2979, i_10_3034, i_10_3070, i_10_3071, i_10_3198, i_10_3199, i_10_3200, i_10_3269, i_10_3284, i_10_3321, i_10_3324, i_10_3325, i_10_3329, i_10_3387, i_10_3409, i_10_3496, i_10_3497, i_10_3585, i_10_3586, i_10_3613, i_10_3614, i_10_3650, i_10_3780, i_10_3781, i_10_3782, i_10_3847, i_10_3848, i_10_3852, i_10_3853, i_10_3856, i_10_3992, i_10_4113, i_10_4121, i_10_4266, i_10_4267, i_10_4270, i_10_4279, i_10_4280, o_10_468);
	kernel_10_469 k_10_469(i_10_32, i_10_50, i_10_52, i_10_53, i_10_121, i_10_132, i_10_146, i_10_148, i_10_149, i_10_175, i_10_224, i_10_259, i_10_260, i_10_262, i_10_393, i_10_426, i_10_427, i_10_433, i_10_443, i_10_463, i_10_464, i_10_466, i_10_745, i_10_751, i_10_752, i_10_983, i_10_1050, i_10_1237, i_10_1238, i_10_1240, i_10_1241, i_10_1247, i_10_1312, i_10_1313, i_10_1534, i_10_1541, i_10_1544, i_10_1576, i_10_1624, i_10_1634, i_10_1640, i_10_1643, i_10_1683, i_10_1684, i_10_1689, i_10_1764, i_10_1819, i_10_1820, i_10_1957, i_10_1981, i_10_2029, i_10_2436, i_10_2471, i_10_2511, i_10_2607, i_10_2663, i_10_2697, i_10_2703, i_10_2704, i_10_2705, i_10_2707, i_10_2708, i_10_2731, i_10_2821, i_10_2829, i_10_2831, i_10_2842, i_10_2887, i_10_2913, i_10_2980, i_10_3045, i_10_3093, i_10_3130, i_10_3200, i_10_3281, i_10_3308, i_10_3385, i_10_3414, i_10_3470, i_10_3471, i_10_3494, i_10_3505, i_10_3587, i_10_3590, i_10_3611, i_10_3622, i_10_3836, i_10_3855, i_10_3858, i_10_3860, i_10_3946, i_10_3947, i_10_3981, i_10_4171, i_10_4204, i_10_4266, i_10_4267, i_10_4395, i_10_4396, i_10_4582, o_10_469);
	kernel_10_470 k_10_470(i_10_221, i_10_245, i_10_273, i_10_320, i_10_329, i_10_388, i_10_409, i_10_432, i_10_433, i_10_434, i_10_441, i_10_443, i_10_444, i_10_445, i_10_446, i_10_459, i_10_463, i_10_464, i_10_512, i_10_713, i_10_875, i_10_959, i_10_990, i_10_991, i_10_992, i_10_1198, i_10_1238, i_10_1265, i_10_1309, i_10_1313, i_10_1654, i_10_1683, i_10_1687, i_10_1688, i_10_1819, i_10_1820, i_10_1821, i_10_1826, i_10_1874, i_10_1990, i_10_1991, i_10_2018, i_10_2021, i_10_2198, i_10_2261, i_10_2264, i_10_2353, i_10_2354, i_10_2359, i_10_2362, i_10_2366, i_10_2377, i_10_2378, i_10_2381, i_10_2459, i_10_2467, i_10_2468, i_10_2628, i_10_2660, i_10_2675, i_10_2720, i_10_2729, i_10_2789, i_10_2826, i_10_2829, i_10_2830, i_10_2831, i_10_2918, i_10_2979, i_10_3070, i_10_3076, i_10_3151, i_10_3155, i_10_3156, i_10_3280, i_10_3281, i_10_3388, i_10_3389, i_10_3392, i_10_3466, i_10_3551, i_10_3611, i_10_3612, i_10_3614, i_10_3785, i_10_3834, i_10_3835, i_10_3838, i_10_3856, i_10_3978, i_10_3983, i_10_4027, i_10_4115, i_10_4116, i_10_4126, i_10_4214, i_10_4268, i_10_4279, i_10_4285, i_10_4291, o_10_470);
	kernel_10_471 k_10_471(i_10_149, i_10_172, i_10_173, i_10_176, i_10_178, i_10_250, i_10_323, i_10_425, i_10_428, i_10_429, i_10_430, i_10_431, i_10_466, i_10_467, i_10_504, i_10_505, i_10_507, i_10_508, i_10_715, i_10_716, i_10_718, i_10_794, i_10_896, i_10_965, i_10_1233, i_10_1305, i_10_1308, i_10_1310, i_10_1312, i_10_1313, i_10_1546, i_10_1631, i_10_1651, i_10_1652, i_10_1654, i_10_1655, i_10_1684, i_10_1685, i_10_1687, i_10_1768, i_10_1991, i_10_1994, i_10_2000, i_10_2255, i_10_2349, i_10_2354, i_10_2357, i_10_2404, i_10_2450, i_10_2453, i_10_2567, i_10_2570, i_10_2572, i_10_2628, i_10_2675, i_10_2703, i_10_2710, i_10_2711, i_10_2714, i_10_2716, i_10_2717, i_10_2883, i_10_3036, i_10_3037, i_10_3038, i_10_3072, i_10_3269, i_10_3322, i_10_3384, i_10_3385, i_10_3386, i_10_3388, i_10_3389, i_10_3391, i_10_3392, i_10_3404, i_10_3406, i_10_3410, i_10_3524, i_10_3527, i_10_3583, i_10_3589, i_10_3650, i_10_3652, i_10_3684, i_10_3837, i_10_3846, i_10_3847, i_10_3848, i_10_3857, i_10_3872, i_10_3947, i_10_4027, i_10_4028, i_10_4123, i_10_4285, i_10_4286, i_10_4288, i_10_4289, i_10_4291, o_10_471);
	kernel_10_472 k_10_472(i_10_64, i_10_65, i_10_68, i_10_175, i_10_176, i_10_178, i_10_179, i_10_272, i_10_279, i_10_285, i_10_316, i_10_317, i_10_319, i_10_320, i_10_408, i_10_413, i_10_433, i_10_437, i_10_533, i_10_635, i_10_638, i_10_641, i_10_644, i_10_896, i_10_1055, i_10_1081, i_10_1233, i_10_1249, i_10_1298, i_10_1306, i_10_1307, i_10_1309, i_10_1364, i_10_1433, i_10_1436, i_10_1487, i_10_1622, i_10_1648, i_10_1651, i_10_1652, i_10_1655, i_10_1685, i_10_1690, i_10_1768, i_10_1796, i_10_1874, i_10_2021, i_10_2024, i_10_2237, i_10_2264, i_10_2351, i_10_2356, i_10_2381, i_10_2453, i_10_2468, i_10_2470, i_10_2513, i_10_2519, i_10_2567, i_10_2629, i_10_2632, i_10_2633, i_10_2704, i_10_2711, i_10_2717, i_10_2735, i_10_2744, i_10_2831, i_10_2846, i_10_3044, i_10_3045, i_10_3071, i_10_3317, i_10_3384, i_10_3386, i_10_3388, i_10_3389, i_10_3467, i_10_3469, i_10_3470, i_10_3494, i_10_3539, i_10_3542, i_10_3557, i_10_3584, i_10_3586, i_10_3587, i_10_3647, i_10_3775, i_10_3794, i_10_3847, i_10_3848, i_10_3944, i_10_4114, i_10_4121, i_10_4167, i_10_4267, i_10_4276, i_10_4289, i_10_4586, o_10_472);
	kernel_10_473 k_10_473(i_10_174, i_10_292, i_10_295, i_10_296, i_10_394, i_10_405, i_10_429, i_10_431, i_10_438, i_10_444, i_10_445, i_10_447, i_10_449, i_10_460, i_10_795, i_10_798, i_10_800, i_10_823, i_10_826, i_10_850, i_10_852, i_10_853, i_10_1033, i_10_1052, i_10_1202, i_10_1235, i_10_1236, i_10_1237, i_10_1238, i_10_1266, i_10_1309, i_10_1310, i_10_1342, i_10_1378, i_10_1435, i_10_1436, i_10_1553, i_10_1579, i_10_1580, i_10_1651, i_10_1652, i_10_1653, i_10_1680, i_10_1688, i_10_1823, i_10_1996, i_10_2084, i_10_2158, i_10_2184, i_10_2309, i_10_2310, i_10_2311, i_10_2337, i_10_2338, i_10_2351, i_10_2448, i_10_2450, i_10_2463, i_10_2470, i_10_2482, i_10_2532, i_10_2562, i_10_2632, i_10_2660, i_10_2662, i_10_2679, i_10_2697, i_10_2710, i_10_2718, i_10_2829, i_10_2830, i_10_2880, i_10_2918, i_10_2922, i_10_2950, i_10_3091, i_10_3095, i_10_3199, i_10_3278, i_10_3406, i_10_3539, i_10_3555, i_10_3562, i_10_3601, i_10_3602, i_10_3637, i_10_3782, i_10_3785, i_10_3832, i_10_3834, i_10_3840, i_10_3841, i_10_3853, i_10_3902, i_10_3979, i_10_3983, i_10_3995, i_10_4116, i_10_4117, i_10_4180, o_10_473);
	kernel_10_474 k_10_474(i_10_156, i_10_175, i_10_176, i_10_243, i_10_280, i_10_328, i_10_390, i_10_427, i_10_428, i_10_438, i_10_444, i_10_447, i_10_463, i_10_506, i_10_516, i_10_519, i_10_748, i_10_752, i_10_796, i_10_955, i_10_1032, i_10_1033, i_10_1233, i_10_1307, i_10_1308, i_10_1311, i_10_1448, i_10_1550, i_10_1651, i_10_1681, i_10_1682, i_10_1687, i_10_1822, i_10_1823, i_10_1824, i_10_2016, i_10_2353, i_10_2354, i_10_2364, i_10_2407, i_10_2457, i_10_2629, i_10_2631, i_10_2632, i_10_2636, i_10_2662, i_10_2700, i_10_2701, i_10_2713, i_10_2714, i_10_2716, i_10_2723, i_10_2823, i_10_2885, i_10_2920, i_10_2980, i_10_2981, i_10_2982, i_10_2983, i_10_2984, i_10_2985, i_10_3036, i_10_3040, i_10_3043, i_10_3074, i_10_3199, i_10_3276, i_10_3388, i_10_3405, i_10_3406, i_10_3522, i_10_3613, i_10_3615, i_10_3650, i_10_3783, i_10_3841, i_10_3852, i_10_3853, i_10_3854, i_10_3856, i_10_3888, i_10_3910, i_10_3912, i_10_3982, i_10_3983, i_10_3990, i_10_4114, i_10_4116, i_10_4117, i_10_4119, i_10_4266, i_10_4269, i_10_4271, i_10_4273, i_10_4276, i_10_4277, i_10_4289, i_10_4292, i_10_4567, i_10_4570, o_10_474);
	kernel_10_475 k_10_475(i_10_171, i_10_216, i_10_280, i_10_316, i_10_408, i_10_425, i_10_431, i_10_434, i_10_437, i_10_439, i_10_441, i_10_442, i_10_443, i_10_445, i_10_457, i_10_515, i_10_518, i_10_749, i_10_892, i_10_901, i_10_957, i_10_958, i_10_968, i_10_1036, i_10_1037, i_10_1038, i_10_1141, i_10_1246, i_10_1247, i_10_1549, i_10_1579, i_10_1581, i_10_1648, i_10_1653, i_10_1654, i_10_1686, i_10_1818, i_10_1823, i_10_2006, i_10_2022, i_10_2332, i_10_2364, i_10_2383, i_10_2449, i_10_2510, i_10_2629, i_10_2630, i_10_2632, i_10_2633, i_10_2634, i_10_2635, i_10_2636, i_10_2655, i_10_2675, i_10_2678, i_10_2721, i_10_2818, i_10_2822, i_10_2824, i_10_2880, i_10_2884, i_10_2885, i_10_2919, i_10_2923, i_10_2924, i_10_2984, i_10_2987, i_10_3043, i_10_3074, i_10_3152, i_10_3155, i_10_3196, i_10_3312, i_10_3391, i_10_3392, i_10_3497, i_10_3610, i_10_3611, i_10_3645, i_10_3784, i_10_3785, i_10_3787, i_10_3788, i_10_3834, i_10_3841, i_10_3849, i_10_3853, i_10_3888, i_10_3889, i_10_3890, i_10_3906, i_10_3911, i_10_3980, i_10_4087, i_10_4122, i_10_4127, i_10_4288, i_10_4289, i_10_4291, i_10_4568, o_10_475);
	kernel_10_476 k_10_476(i_10_140, i_10_223, i_10_248, i_10_251, i_10_275, i_10_276, i_10_281, i_10_318, i_10_438, i_10_442, i_10_448, i_10_449, i_10_464, i_10_467, i_10_480, i_10_514, i_10_515, i_10_518, i_10_534, i_10_716, i_10_719, i_10_732, i_10_754, i_10_791, i_10_796, i_10_799, i_10_800, i_10_835, i_10_836, i_10_967, i_10_969, i_10_988, i_10_1115, i_10_1163, i_10_1166, i_10_1214, i_10_1309, i_10_1446, i_10_1492, i_10_1493, i_10_1546, i_10_1572, i_10_1653, i_10_1799, i_10_1808, i_10_1820, i_10_1825, i_10_1943, i_10_1952, i_10_2030, i_10_2255, i_10_2310, i_10_2356, i_10_2357, i_10_2363, i_10_2456, i_10_2534, i_10_2545, i_10_2546, i_10_2562, i_10_2607, i_10_2609, i_10_2678, i_10_2717, i_10_2725, i_10_2741, i_10_2876, i_10_2915, i_10_2919, i_10_2920, i_10_2968, i_10_2982, i_10_2986, i_10_3030, i_10_3038, i_10_3122, i_10_3284, i_10_3314, i_10_3315, i_10_3316, i_10_3320, i_10_3496, i_10_3526, i_10_3590, i_10_3617, i_10_3803, i_10_3806, i_10_3848, i_10_3860, i_10_3878, i_10_3946, i_10_3948, i_10_4182, i_10_4183, i_10_4268, i_10_4292, i_10_4306, i_10_4371, i_10_4459, i_10_4463, o_10_476);
	kernel_10_477 k_10_477(i_10_29, i_10_244, i_10_254, i_10_272, i_10_283, i_10_286, i_10_391, i_10_427, i_10_428, i_10_434, i_10_435, i_10_436, i_10_443, i_10_445, i_10_463, i_10_505, i_10_792, i_10_958, i_10_1026, i_10_1027, i_10_1028, i_10_1080, i_10_1081, i_10_1085, i_10_1135, i_10_1235, i_10_1305, i_10_1306, i_10_1307, i_10_1308, i_10_1309, i_10_1364, i_10_1433, i_10_1436, i_10_1621, i_10_1823, i_10_1910, i_10_1911, i_10_1913, i_10_1989, i_10_2030, i_10_2198, i_10_2358, i_10_2408, i_10_2449, i_10_2470, i_10_2539, i_10_2541, i_10_2565, i_10_2628, i_10_2629, i_10_2630, i_10_2631, i_10_2632, i_10_2674, i_10_2675, i_10_2709, i_10_2710, i_10_2714, i_10_2720, i_10_2724, i_10_2730, i_10_2827, i_10_2828, i_10_2830, i_10_2845, i_10_2883, i_10_2919, i_10_3033, i_10_3069, i_10_3070, i_10_3071, i_10_3267, i_10_3321, i_10_3322, i_10_3323, i_10_3328, i_10_3467, i_10_3556, i_10_3584, i_10_3587, i_10_3609, i_10_3645, i_10_3837, i_10_3838, i_10_3839, i_10_3843, i_10_3846, i_10_3847, i_10_3848, i_10_3980, i_10_4030, i_10_4122, i_10_4123, i_10_4125, i_10_4127, i_10_4167, i_10_4172, i_10_4266, i_10_4278, o_10_477);
	kernel_10_478 k_10_478(i_10_13, i_10_31, i_10_174, i_10_221, i_10_223, i_10_224, i_10_285, i_10_286, i_10_315, i_10_316, i_10_435, i_10_725, i_10_748, i_10_820, i_10_967, i_10_983, i_10_999, i_10_1010, i_10_1107, i_10_1218, i_10_1233, i_10_1234, i_10_1240, i_10_1279, i_10_1296, i_10_1302, i_10_1344, i_10_1432, i_10_1535, i_10_1539, i_10_1540, i_10_1562, i_10_1683, i_10_1684, i_10_1686, i_10_1689, i_10_1691, i_10_1795, i_10_1800, i_10_1803, i_10_1821, i_10_1980, i_10_1982, i_10_2038, i_10_2089, i_10_2090, i_10_2199, i_10_2235, i_10_2252, i_10_2255, i_10_2290, i_10_2352, i_10_2355, i_10_2452, i_10_2466, i_10_2467, i_10_2471, i_10_2503, i_10_2565, i_10_2567, i_10_2574, i_10_2631, i_10_2721, i_10_2726, i_10_2727, i_10_2728, i_10_2730, i_10_2832, i_10_2847, i_10_2914, i_10_2964, i_10_3045, i_10_3384, i_10_3432, i_10_3468, i_10_3469, i_10_3537, i_10_3582, i_10_3612, i_10_3614, i_10_3793, i_10_3834, i_10_3854, i_10_3855, i_10_3860, i_10_3873, i_10_3874, i_10_3911, i_10_3988, i_10_4122, i_10_4125, i_10_4154, i_10_4168, i_10_4218, i_10_4283, i_10_4287, i_10_4460, i_10_4502, i_10_4545, i_10_4546, o_10_478);
	kernel_10_479 k_10_479(i_10_118, i_10_121, i_10_248, i_10_285, i_10_286, i_10_287, i_10_315, i_10_316, i_10_318, i_10_365, i_10_406, i_10_408, i_10_424, i_10_434, i_10_443, i_10_447, i_10_448, i_10_793, i_10_794, i_10_797, i_10_893, i_10_959, i_10_1028, i_10_1031, i_10_1242, i_10_1243, i_10_1244, i_10_1305, i_10_1309, i_10_1444, i_10_1445, i_10_1546, i_10_1547, i_10_1576, i_10_1577, i_10_1580, i_10_1613, i_10_1650, i_10_1683, i_10_1687, i_10_1689, i_10_1801, i_10_1821, i_10_1990, i_10_2197, i_10_2304, i_10_2332, i_10_2361, i_10_2362, i_10_2363, i_10_2376, i_10_2407, i_10_2458, i_10_2467, i_10_2475, i_10_2648, i_10_2663, i_10_2713, i_10_2785, i_10_2828, i_10_2830, i_10_2831, i_10_2881, i_10_2917, i_10_2919, i_10_2920, i_10_3201, i_10_3269, i_10_3276, i_10_3277, i_10_3281, i_10_3294, i_10_3384, i_10_3386, i_10_3388, i_10_3550, i_10_3647, i_10_3686, i_10_3717, i_10_3781, i_10_3783, i_10_3784, i_10_3785, i_10_3786, i_10_3788, i_10_3842, i_10_3845, i_10_3846, i_10_3847, i_10_3851, i_10_3852, i_10_3854, i_10_3855, i_10_3888, i_10_3889, i_10_4061, i_10_4218, i_10_4219, i_10_4289, i_10_4564, o_10_479);
	kernel_10_480 k_10_480(i_10_172, i_10_186, i_10_187, i_10_244, i_10_246, i_10_247, i_10_280, i_10_286, i_10_293, i_10_423, i_10_424, i_10_446, i_10_449, i_10_460, i_10_463, i_10_464, i_10_467, i_10_712, i_10_713, i_10_748, i_10_901, i_10_902, i_10_905, i_10_997, i_10_998, i_10_1034, i_10_1168, i_10_1222, i_10_1234, i_10_1237, i_10_1306, i_10_1309, i_10_1345, i_10_1361, i_10_1486, i_10_1556, i_10_1649, i_10_1683, i_10_1684, i_10_1686, i_10_1765, i_10_1766, i_10_1818, i_10_1825, i_10_1909, i_10_1914, i_10_1999, i_10_2183, i_10_2349, i_10_2365, i_10_2366, i_10_2380, i_10_2449, i_10_2450, i_10_2452, i_10_2470, i_10_2659, i_10_2725, i_10_2727, i_10_2782, i_10_2830, i_10_2883, i_10_2886, i_10_2918, i_10_3044, i_10_3070, i_10_3071, i_10_3115, i_10_3233, i_10_3276, i_10_3280, i_10_3281, i_10_3325, i_10_3389, i_10_3392, i_10_3407, i_10_3408, i_10_3409, i_10_3538, i_10_3583, i_10_3585, i_10_3586, i_10_3614, i_10_3653, i_10_3783, i_10_3787, i_10_3788, i_10_3808, i_10_3811, i_10_3812, i_10_3839, i_10_3855, i_10_3859, i_10_3966, i_10_3978, i_10_3980, i_10_3982, i_10_4115, i_10_4289, i_10_4291, o_10_480);
	kernel_10_481 k_10_481(i_10_44, i_10_58, i_10_153, i_10_208, i_10_257, i_10_263, i_10_281, i_10_283, i_10_317, i_10_355, i_10_389, i_10_392, i_10_499, i_10_657, i_10_658, i_10_893, i_10_1009, i_10_1010, i_10_1027, i_10_1084, i_10_1085, i_10_1206, i_10_1234, i_10_1238, i_10_1271, i_10_1297, i_10_1377, i_10_1396, i_10_1485, i_10_1550, i_10_1576, i_10_1593, i_10_1638, i_10_1651, i_10_1697, i_10_1712, i_10_1716, i_10_1730, i_10_1807, i_10_1809, i_10_1822, i_10_2000, i_10_2002, i_10_2027, i_10_2145, i_10_2231, i_10_2269, i_10_2307, i_10_2341, i_10_2343, i_10_2362, i_10_2467, i_10_2489, i_10_2504, i_10_2542, i_10_2556, i_10_2557, i_10_2575, i_10_2885, i_10_2954, i_10_2961, i_10_2971, i_10_2983, i_10_2984, i_10_3070, i_10_3071, i_10_3160, i_10_3197, i_10_3200, i_10_3266, i_10_3332, i_10_3358, i_10_3404, i_10_3467, i_10_3484, i_10_3539, i_10_3580, i_10_3584, i_10_3587, i_10_3613, i_10_3645, i_10_3729, i_10_3792, i_10_3808, i_10_3842, i_10_3898, i_10_3945, i_10_4069, i_10_4118, i_10_4144, i_10_4151, i_10_4204, i_10_4226, i_10_4270, i_10_4273, i_10_4394, i_10_4421, i_10_4522, i_10_4545, i_10_4546, o_10_481);
	kernel_10_482 k_10_482(i_10_155, i_10_171, i_10_172, i_10_219, i_10_220, i_10_280, i_10_320, i_10_437, i_10_445, i_10_446, i_10_448, i_10_518, i_10_590, i_10_689, i_10_992, i_10_995, i_10_997, i_10_1026, i_10_1037, i_10_1040, i_10_1236, i_10_1241, i_10_1289, i_10_1305, i_10_1342, i_10_1346, i_10_1486, i_10_1487, i_10_1556, i_10_1595, i_10_1630, i_10_1647, i_10_1683, i_10_1686, i_10_1687, i_10_1771, i_10_1819, i_10_1821, i_10_1912, i_10_1913, i_10_1998, i_10_2002, i_10_2243, i_10_2252, i_10_2351, i_10_2408, i_10_2454, i_10_2456, i_10_2512, i_10_2543, i_10_2606, i_10_2609, i_10_2657, i_10_2660, i_10_2675, i_10_2720, i_10_2723, i_10_2724, i_10_2728, i_10_2729, i_10_2819, i_10_2821, i_10_2822, i_10_2885, i_10_2981, i_10_2984, i_10_3037, i_10_3089, i_10_3091, i_10_3095, i_10_3160, i_10_3161, i_10_3235, i_10_3236, i_10_3278, i_10_3281, i_10_3284, i_10_3388, i_10_3389, i_10_3391, i_10_3392, i_10_3469, i_10_3470, i_10_3523, i_10_3524, i_10_3525, i_10_3527, i_10_3554, i_10_3781, i_10_3785, i_10_3836, i_10_3980, i_10_3992, i_10_4055, i_10_4114, i_10_4126, i_10_4268, i_10_4285, i_10_4460, i_10_4565, o_10_482);
	kernel_10_483 k_10_483(i_10_284, i_10_287, i_10_318, i_10_323, i_10_388, i_10_412, i_10_431, i_10_443, i_10_465, i_10_719, i_10_800, i_10_1030, i_10_1038, i_10_1041, i_10_1043, i_10_1052, i_10_1053, i_10_1060, i_10_1061, i_10_1084, i_10_1269, i_10_1308, i_10_1311, i_10_1312, i_10_1394, i_10_1435, i_10_1439, i_10_1444, i_10_1539, i_10_1540, i_10_1577, i_10_1624, i_10_1652, i_10_1654, i_10_1686, i_10_1687, i_10_1689, i_10_1765, i_10_1769, i_10_1819, i_10_1824, i_10_1915, i_10_1999, i_10_2001, i_10_2159, i_10_2349, i_10_2352, i_10_2355, i_10_2357, i_10_2365, i_10_2376, i_10_2378, i_10_2405, i_10_2406, i_10_2454, i_10_2456, i_10_2470, i_10_2516, i_10_2564, i_10_2604, i_10_2632, i_10_2644, i_10_2677, i_10_2699, i_10_2714, i_10_2956, i_10_2959, i_10_2980, i_10_2982, i_10_2983, i_10_2984, i_10_2985, i_10_3036, i_10_3268, i_10_3272, i_10_3278, i_10_3297, i_10_3384, i_10_3385, i_10_3388, i_10_3389, i_10_3472, i_10_3617, i_10_3645, i_10_3649, i_10_3784, i_10_3785, i_10_3834, i_10_3852, i_10_4009, i_10_4114, i_10_4125, i_10_4130, i_10_4170, i_10_4173, i_10_4174, i_10_4267, i_10_4271, i_10_4278, i_10_4279, o_10_483);
	kernel_10_484 k_10_484(i_10_176, i_10_284, i_10_405, i_10_406, i_10_409, i_10_459, i_10_747, i_10_999, i_10_1000, i_10_1027, i_10_1139, i_10_1141, i_10_1234, i_10_1238, i_10_1432, i_10_1489, i_10_1539, i_10_1575, i_10_1576, i_10_1578, i_10_1647, i_10_1650, i_10_1651, i_10_1691, i_10_1909, i_10_1945, i_10_1951, i_10_2017, i_10_2151, i_10_2178, i_10_2179, i_10_2181, i_10_2185, i_10_2196, i_10_2197, i_10_2199, i_10_2305, i_10_2306, i_10_2349, i_10_2350, i_10_2351, i_10_2352, i_10_2353, i_10_2355, i_10_2377, i_10_2406, i_10_2469, i_10_2662, i_10_2700, i_10_2711, i_10_2712, i_10_2714, i_10_2724, i_10_2833, i_10_2887, i_10_2916, i_10_2917, i_10_2919, i_10_2923, i_10_2954, i_10_2979, i_10_3069, i_10_3150, i_10_3267, i_10_3268, i_10_3270, i_10_3271, i_10_3280, i_10_3330, i_10_3385, i_10_3387, i_10_3522, i_10_3525, i_10_3526, i_10_3584, i_10_3585, i_10_3587, i_10_3614, i_10_3615, i_10_3616, i_10_3617, i_10_3645, i_10_3649, i_10_3685, i_10_3807, i_10_3837, i_10_3838, i_10_3852, i_10_3889, i_10_3907, i_10_3980, i_10_3984, i_10_4266, i_10_4268, i_10_4271, i_10_4275, i_10_4276, i_10_4287, i_10_4567, i_10_4568, o_10_484);
	kernel_10_485 k_10_485(i_10_28, i_10_45, i_10_223, i_10_254, i_10_290, i_10_299, i_10_389, i_10_424, i_10_425, i_10_434, i_10_462, i_10_740, i_10_1003, i_10_1027, i_10_1028, i_10_1034, i_10_1055, i_10_1082, i_10_1118, i_10_1233, i_10_1235, i_10_1236, i_10_1238, i_10_1243, i_10_1244, i_10_1342, i_10_1379, i_10_1541, i_10_1552, i_10_1577, i_10_1625, i_10_1651, i_10_1683, i_10_1687, i_10_1710, i_10_1711, i_10_1914, i_10_2036, i_10_2090, i_10_2179, i_10_2180, i_10_2200, i_10_2306, i_10_2332, i_10_2353, i_10_2354, i_10_2359, i_10_2360, i_10_2362, i_10_2379, i_10_2448, i_10_2451, i_10_2452, i_10_2456, i_10_2468, i_10_2470, i_10_2471, i_10_2542, i_10_2653, i_10_2673, i_10_2713, i_10_2731, i_10_2838, i_10_2920, i_10_2958, i_10_3070, i_10_3200, i_10_3278, i_10_3280, i_10_3281, i_10_3403, i_10_3467, i_10_3548, i_10_3590, i_10_3612, i_10_3649, i_10_3650, i_10_3683, i_10_3772, i_10_3781, i_10_3784, i_10_3785, i_10_3835, i_10_3858, i_10_3859, i_10_3860, i_10_3881, i_10_3907, i_10_3982, i_10_4114, i_10_4115, i_10_4205, i_10_4213, i_10_4214, i_10_4217, i_10_4220, i_10_4270, i_10_4287, i_10_4430, i_10_4529, o_10_485);
	kernel_10_486 k_10_486(i_10_48, i_10_144, i_10_145, i_10_172, i_10_220, i_10_261, i_10_263, i_10_280, i_10_281, i_10_285, i_10_287, i_10_327, i_10_390, i_10_406, i_10_409, i_10_442, i_10_445, i_10_461, i_10_467, i_10_586, i_10_711, i_10_712, i_10_793, i_10_795, i_10_798, i_10_799, i_10_955, i_10_1237, i_10_1240, i_10_1266, i_10_1312, i_10_1313, i_10_1365, i_10_1539, i_10_1553, i_10_1651, i_10_1685, i_10_1686, i_10_1801, i_10_1802, i_10_1818, i_10_1825, i_10_1913, i_10_1998, i_10_2025, i_10_2206, i_10_2223, i_10_2224, i_10_2356, i_10_2361, i_10_2469, i_10_2471, i_10_2473, i_10_2601, i_10_2634, i_10_2635, i_10_2677, i_10_2703, i_10_2704, i_10_2722, i_10_2723, i_10_2727, i_10_2729, i_10_2731, i_10_2829, i_10_3034, i_10_3231, i_10_3234, i_10_3267, i_10_3268, i_10_3277, i_10_3384, i_10_3391, i_10_3496, i_10_3501, i_10_3507, i_10_3519, i_10_3522, i_10_3523, i_10_3524, i_10_3583, i_10_3587, i_10_3588, i_10_3590, i_10_3783, i_10_3785, i_10_3788, i_10_3834, i_10_3837, i_10_3838, i_10_3839, i_10_3846, i_10_3848, i_10_3855, i_10_4114, i_10_4213, i_10_4269, i_10_4275, i_10_4276, i_10_4289, o_10_486);
	kernel_10_487 k_10_487(i_10_28, i_10_70, i_10_118, i_10_175, i_10_176, i_10_260, i_10_315, i_10_327, i_10_387, i_10_391, i_10_443, i_10_461, i_10_514, i_10_797, i_10_799, i_10_800, i_10_897, i_10_899, i_10_971, i_10_1240, i_10_1241, i_10_1243, i_10_1246, i_10_1311, i_10_1348, i_10_1434, i_10_1539, i_10_1543, i_10_1549, i_10_1552, i_10_1630, i_10_1650, i_10_1651, i_10_1686, i_10_1690, i_10_1821, i_10_1822, i_10_1823, i_10_1913, i_10_1945, i_10_1949, i_10_1996, i_10_2365, i_10_2404, i_10_2448, i_10_2449, i_10_2453, i_10_2456, i_10_2471, i_10_2518, i_10_2660, i_10_2663, i_10_2708, i_10_2716, i_10_2717, i_10_2723, i_10_2732, i_10_2733, i_10_2787, i_10_2788, i_10_2831, i_10_2833, i_10_3033, i_10_3034, i_10_3036, i_10_3041, i_10_3045, i_10_3199, i_10_3238, i_10_3269, i_10_3390, i_10_3409, i_10_3437, i_10_3526, i_10_3613, i_10_3616, i_10_3617, i_10_3640, i_10_3649, i_10_3650, i_10_3653, i_10_3781, i_10_3782, i_10_3787, i_10_3811, i_10_3839, i_10_3840, i_10_3856, i_10_3857, i_10_3860, i_10_3882, i_10_3949, i_10_3991, i_10_4025, i_10_4056, i_10_4267, i_10_4270, i_10_4276, i_10_4283, i_10_4291, o_10_487);
	kernel_10_488 k_10_488(i_10_139, i_10_279, i_10_280, i_10_361, i_10_441, i_10_442, i_10_461, i_10_496, i_10_585, i_10_748, i_10_749, i_10_754, i_10_792, i_10_795, i_10_796, i_10_828, i_10_830, i_10_924, i_10_955, i_10_983, i_10_1163, i_10_1239, i_10_1243, i_10_1264, i_10_1492, i_10_1540, i_10_1629, i_10_1630, i_10_1631, i_10_1635, i_10_1636, i_10_1644, i_10_1645, i_10_1654, i_10_1655, i_10_1683, i_10_1684, i_10_1720, i_10_1801, i_10_1802, i_10_1818, i_10_1819, i_10_2004, i_10_2005, i_10_2006, i_10_2031, i_10_2032, i_10_2206, i_10_2241, i_10_2248, i_10_2386, i_10_2387, i_10_2472, i_10_2473, i_10_2474, i_10_2539, i_10_2660, i_10_2661, i_10_2663, i_10_2674, i_10_2681, i_10_2717, i_10_2733, i_10_2743, i_10_2817, i_10_2824, i_10_2922, i_10_2979, i_10_2980, i_10_2982, i_10_2983, i_10_2985, i_10_2986, i_10_3237, i_10_3238, i_10_3282, i_10_3283, i_10_3313, i_10_3465, i_10_3493, i_10_3508, i_10_3520, i_10_3525, i_10_3724, i_10_3798, i_10_3854, i_10_3912, i_10_3948, i_10_3949, i_10_4061, i_10_4115, i_10_4269, i_10_4272, i_10_4284, i_10_4302, i_10_4303, i_10_4457, i_10_4459, i_10_4582, i_10_4583, o_10_488);
	kernel_10_489 k_10_489(i_10_23, i_10_137, i_10_271, i_10_272, i_10_274, i_10_275, i_10_286, i_10_287, i_10_317, i_10_388, i_10_461, i_10_506, i_10_641, i_10_692, i_10_715, i_10_752, i_10_799, i_10_821, i_10_831, i_10_1157, i_10_1171, i_10_1209, i_10_1210, i_10_1240, i_10_1243, i_10_1245, i_10_1308, i_10_1312, i_10_1328, i_10_1432, i_10_1450, i_10_1522, i_10_1531, i_10_1534, i_10_1535, i_10_1544, i_10_1580, i_10_1603, i_10_1622, i_10_1633, i_10_1688, i_10_1693, i_10_1711, i_10_1717, i_10_1718, i_10_1805, i_10_1822, i_10_1826, i_10_1981, i_10_2028, i_10_2029, i_10_2110, i_10_2113, i_10_2181, i_10_2209, i_10_2228, i_10_2354, i_10_2376, i_10_2455, i_10_2513, i_10_2557, i_10_2629, i_10_2632, i_10_2633, i_10_2665, i_10_2667, i_10_2702, i_10_2704, i_10_2705, i_10_2714, i_10_2786, i_10_2966, i_10_2983, i_10_3119, i_10_3166, i_10_3203, i_10_3296, i_10_3404, i_10_3497, i_10_3500, i_10_3502, i_10_3538, i_10_3547, i_10_3610, i_10_3614, i_10_3615, i_10_3688, i_10_3779, i_10_3808, i_10_3830, i_10_3853, i_10_3854, i_10_3857, i_10_3859, i_10_3875, i_10_4001, i_10_4276, i_10_4340, i_10_4456, i_10_4532, o_10_489);
	kernel_10_490 k_10_490(i_10_34, i_10_35, i_10_286, i_10_315, i_10_319, i_10_324, i_10_328, i_10_330, i_10_393, i_10_430, i_10_435, i_10_438, i_10_439, i_10_440, i_10_442, i_10_457, i_10_516, i_10_520, i_10_700, i_10_951, i_10_996, i_10_997, i_10_1006, i_10_1052, i_10_1138, i_10_1140, i_10_1236, i_10_1237, i_10_1238, i_10_1250, i_10_1307, i_10_1309, i_10_1312, i_10_1384, i_10_1385, i_10_1457, i_10_1554, i_10_1555, i_10_1578, i_10_1600, i_10_1687, i_10_1688, i_10_1690, i_10_1691, i_10_1768, i_10_1769, i_10_1815, i_10_1816, i_10_1825, i_10_1826, i_10_2004, i_10_2310, i_10_2312, i_10_2350, i_10_2351, i_10_2364, i_10_2408, i_10_2411, i_10_2464, i_10_2509, i_10_2510, i_10_2515, i_10_2728, i_10_2831, i_10_2883, i_10_2887, i_10_2919, i_10_2922, i_10_2923, i_10_2924, i_10_2959, i_10_2982, i_10_2983, i_10_2985, i_10_2986, i_10_3093, i_10_3094, i_10_3156, i_10_3199, i_10_3203, i_10_3284, i_10_3319, i_10_3389, i_10_3545, i_10_3613, i_10_3733, i_10_3855, i_10_3857, i_10_3895, i_10_3981, i_10_3982, i_10_3984, i_10_3985, i_10_3986, i_10_3992, i_10_4003, i_10_4217, i_10_4288, i_10_4291, i_10_4292, o_10_490);
	kernel_10_491 k_10_491(i_10_30, i_10_123, i_10_171, i_10_243, i_10_281, i_10_283, i_10_286, i_10_287, i_10_432, i_10_464, i_10_465, i_10_711, i_10_747, i_10_892, i_10_955, i_10_956, i_10_1026, i_10_1233, i_10_1242, i_10_1263, i_10_1308, i_10_1310, i_10_1381, i_10_1396, i_10_1434, i_10_1450, i_10_1612, i_10_1652, i_10_1688, i_10_1766, i_10_1818, i_10_1989, i_10_1990, i_10_2181, i_10_2182, i_10_2185, i_10_2196, i_10_2358, i_10_2452, i_10_2453, i_10_2458, i_10_2566, i_10_2637, i_10_2683, i_10_2713, i_10_2714, i_10_2728, i_10_2729, i_10_2826, i_10_2827, i_10_2831, i_10_2869, i_10_2916, i_10_2917, i_10_2919, i_10_3040, i_10_3075, i_10_3076, i_10_3199, i_10_3200, i_10_3276, i_10_3283, i_10_3384, i_10_3385, i_10_3388, i_10_3408, i_10_3440, i_10_3466, i_10_3550, i_10_3551, i_10_3585, i_10_3586, i_10_3645, i_10_3646, i_10_3651, i_10_3726, i_10_3781, i_10_3782, i_10_3784, i_10_3785, i_10_3829, i_10_3843, i_10_3844, i_10_3847, i_10_3852, i_10_3854, i_10_3856, i_10_3857, i_10_3858, i_10_3860, i_10_3980, i_10_3987, i_10_3991, i_10_4024, i_10_4115, i_10_4149, i_10_4172, i_10_4288, i_10_4289, i_10_4291, o_10_491);
	kernel_10_492 k_10_492(i_10_174, i_10_175, i_10_184, i_10_186, i_10_187, i_10_220, i_10_223, i_10_282, i_10_283, i_10_296, i_10_321, i_10_322, i_10_323, i_10_388, i_10_449, i_10_507, i_10_718, i_10_795, i_10_796, i_10_962, i_10_993, i_10_1041, i_10_1042, i_10_1141, i_10_1142, i_10_1308, i_10_1309, i_10_1546, i_10_1582, i_10_1683, i_10_1687, i_10_1688, i_10_1690, i_10_1821, i_10_1822, i_10_1824, i_10_1951, i_10_2179, i_10_2180, i_10_2352, i_10_2353, i_10_2354, i_10_2355, i_10_2364, i_10_2365, i_10_2407, i_10_2409, i_10_2451, i_10_2452, i_10_2453, i_10_2662, i_10_2681, i_10_2700, i_10_2702, i_10_2722, i_10_2725, i_10_2827, i_10_2883, i_10_2884, i_10_2887, i_10_2917, i_10_2919, i_10_2979, i_10_2986, i_10_3043, i_10_3201, i_10_3280, i_10_3283, i_10_3387, i_10_3405, i_10_3544, i_10_3549, i_10_3612, i_10_3613, i_10_3614, i_10_3647, i_10_3652, i_10_3780, i_10_3782, i_10_3783, i_10_3851, i_10_3855, i_10_3857, i_10_3859, i_10_3894, i_10_3915, i_10_3985, i_10_4114, i_10_4119, i_10_4123, i_10_4126, i_10_4127, i_10_4175, i_10_4282, i_10_4292, i_10_4564, i_10_4565, i_10_4566, i_10_4567, i_10_4568, o_10_492);
	kernel_10_493 k_10_493(i_10_120, i_10_245, i_10_257, i_10_317, i_10_320, i_10_329, i_10_390, i_10_393, i_10_435, i_10_436, i_10_437, i_10_438, i_10_589, i_10_641, i_10_688, i_10_712, i_10_869, i_10_921, i_10_992, i_10_993, i_10_1002, i_10_1006, i_10_1135, i_10_1215, i_10_1216, i_10_1217, i_10_1218, i_10_1219, i_10_1238, i_10_1267, i_10_1305, i_10_1309, i_10_1311, i_10_1615, i_10_1618, i_10_1653, i_10_1804, i_10_1819, i_10_1921, i_10_1947, i_10_1948, i_10_1950, i_10_2021, i_10_2155, i_10_2202, i_10_2203, i_10_2355, i_10_2377, i_10_2513, i_10_2514, i_10_2515, i_10_2540, i_10_2543, i_10_2582, i_10_2613, i_10_2655, i_10_2662, i_10_2677, i_10_2744, i_10_2811, i_10_2812, i_10_2824, i_10_2831, i_10_2834, i_10_2848, i_10_2880, i_10_2881, i_10_2882, i_10_3059, i_10_3090, i_10_3332, i_10_3353, i_10_3397, i_10_3404, i_10_3443, i_10_3445, i_10_3473, i_10_3525, i_10_3539, i_10_3651, i_10_3687, i_10_3717, i_10_3718, i_10_3721, i_10_3815, i_10_3837, i_10_3853, i_10_3893, i_10_3910, i_10_3912, i_10_3928, i_10_3993, i_10_4054, i_10_4168, i_10_4185, i_10_4233, i_10_4276, i_10_4280, i_10_4283, i_10_4519, o_10_493);
	kernel_10_494 k_10_494(i_10_171, i_10_174, i_10_181, i_10_283, i_10_285, i_10_287, i_10_328, i_10_388, i_10_424, i_10_425, i_10_434, i_10_438, i_10_451, i_10_459, i_10_749, i_10_753, i_10_754, i_10_755, i_10_797, i_10_968, i_10_1037, i_10_1234, i_10_1235, i_10_1240, i_10_1242, i_10_1306, i_10_1309, i_10_1359, i_10_1650, i_10_1687, i_10_1688, i_10_1819, i_10_1821, i_10_1822, i_10_1823, i_10_1996, i_10_2362, i_10_2383, i_10_2448, i_10_2451, i_10_2628, i_10_2629, i_10_2630, i_10_2634, i_10_2655, i_10_2656, i_10_2657, i_10_2659, i_10_2713, i_10_2715, i_10_2716, i_10_2717, i_10_2919, i_10_2921, i_10_2923, i_10_3036, i_10_3046, i_10_3050, i_10_3085, i_10_3094, i_10_3155, i_10_3271, i_10_3280, i_10_3284, i_10_3402, i_10_3405, i_10_3408, i_10_3586, i_10_3609, i_10_3613, i_10_3614, i_10_3615, i_10_3616, i_10_3785, i_10_3834, i_10_3840, i_10_3841, i_10_3846, i_10_3847, i_10_3848, i_10_3852, i_10_3856, i_10_3857, i_10_3858, i_10_3859, i_10_3860, i_10_3990, i_10_3991, i_10_4116, i_10_4117, i_10_4119, i_10_4120, i_10_4123, i_10_4269, i_10_4270, i_10_4287, i_10_4288, i_10_4563, i_10_4567, i_10_4568, o_10_494);
	kernel_10_495 k_10_495(i_10_32, i_10_129, i_10_158, i_10_161, i_10_264, i_10_274, i_10_441, i_10_446, i_10_518, i_10_561, i_10_674, i_10_718, i_10_755, i_10_834, i_10_835, i_10_922, i_10_986, i_10_989, i_10_997, i_10_998, i_10_1002, i_10_1005, i_10_1061, i_10_1103, i_10_1234, i_10_1235, i_10_1248, i_10_1249, i_10_1340, i_10_1345, i_10_1452, i_10_1488, i_10_1493, i_10_1538, i_10_1555, i_10_1582, i_10_1637, i_10_1641, i_10_1646, i_10_1799, i_10_1818, i_10_1820, i_10_1821, i_10_1822, i_10_1824, i_10_1940, i_10_1942, i_10_1945, i_10_2003, i_10_2033, i_10_2069, i_10_2258, i_10_2408, i_10_2452, i_10_2472, i_10_2605, i_10_2636, i_10_2681, i_10_2712, i_10_2714, i_10_2717, i_10_2723, i_10_2734, i_10_2735, i_10_2804, i_10_2870, i_10_2956, i_10_2986, i_10_2987, i_10_3011, i_10_3039, i_10_3047, i_10_3074, i_10_3158, i_10_3238, i_10_3239, i_10_3282, i_10_3360, i_10_3387, i_10_3406, i_10_3468, i_10_3470, i_10_3496, i_10_3506, i_10_3509, i_10_3561, i_10_3617, i_10_3624, i_10_3806, i_10_3815, i_10_3846, i_10_3884, i_10_3913, i_10_3946, i_10_3947, i_10_3950, i_10_4271, i_10_4278, i_10_4290, i_10_4292, o_10_495);
	kernel_10_496 k_10_496(i_10_71, i_10_119, i_10_254, i_10_257, i_10_265, i_10_266, i_10_279, i_10_392, i_10_395, i_10_448, i_10_466, i_10_517, i_10_535, i_10_560, i_10_895, i_10_1000, i_10_1003, i_10_1004, i_10_1028, i_10_1109, i_10_1112, i_10_1236, i_10_1239, i_10_1273, i_10_1298, i_10_1300, i_10_1309, i_10_1311, i_10_1312, i_10_1360, i_10_1364, i_10_1400, i_10_1436, i_10_1625, i_10_1648, i_10_1652, i_10_1712, i_10_1799, i_10_1804, i_10_1805, i_10_1808, i_10_1909, i_10_1914, i_10_1919, i_10_1985, i_10_2080, i_10_2178, i_10_2186, i_10_2188, i_10_2350, i_10_2356, i_10_2379, i_10_2382, i_10_2430, i_10_2450, i_10_2506, i_10_2547, i_10_2557, i_10_2558, i_10_2560, i_10_2561, i_10_2566, i_10_2567, i_10_2569, i_10_2597, i_10_2641, i_10_2701, i_10_2705, i_10_2708, i_10_2848, i_10_2849, i_10_3033, i_10_3034, i_10_3200, i_10_3232, i_10_3235, i_10_3270, i_10_3274, i_10_3278, i_10_3283, i_10_3289, i_10_3292, i_10_3429, i_10_3430, i_10_3466, i_10_3470, i_10_3540, i_10_3542, i_10_3568, i_10_3652, i_10_3794, i_10_3797, i_10_3838, i_10_3841, i_10_4148, i_10_4171, i_10_4277, i_10_4282, i_10_4567, i_10_4589, o_10_496);
	kernel_10_497 k_10_497(i_10_123, i_10_216, i_10_261, i_10_279, i_10_280, i_10_281, i_10_282, i_10_320, i_10_405, i_10_443, i_10_444, i_10_460, i_10_462, i_10_904, i_10_956, i_10_1053, i_10_1239, i_10_1263, i_10_1311, i_10_1431, i_10_1432, i_10_1449, i_10_1539, i_10_1540, i_10_1542, i_10_1581, i_10_1620, i_10_1629, i_10_1630, i_10_1651, i_10_1652, i_10_1685, i_10_1800, i_10_1823, i_10_1944, i_10_2025, i_10_2026, i_10_2199, i_10_2331, i_10_2351, i_10_2355, i_10_2403, i_10_2404, i_10_2448, i_10_2449, i_10_2452, i_10_2470, i_10_2545, i_10_2565, i_10_2604, i_10_2647, i_10_2662, i_10_2709, i_10_2718, i_10_2720, i_10_2727, i_10_2821, i_10_2826, i_10_2844, i_10_2865, i_10_2961, i_10_3042, i_10_3089, i_10_3278, i_10_3333, i_10_3386, i_10_3387, i_10_3388, i_10_3390, i_10_3408, i_10_3468, i_10_3471, i_10_3537, i_10_3555, i_10_3582, i_10_3610, i_10_3613, i_10_3618, i_10_3621, i_10_3645, i_10_3648, i_10_3785, i_10_3840, i_10_3846, i_10_3847, i_10_3855, i_10_3856, i_10_3858, i_10_3915, i_10_3978, i_10_3980, i_10_4023, i_10_4024, i_10_4028, i_10_4113, i_10_4122, i_10_4169, i_10_4564, i_10_4566, i_10_4581, o_10_497);
	kernel_10_498 k_10_498(i_10_30, i_10_34, i_10_295, i_10_296, i_10_320, i_10_322, i_10_323, i_10_437, i_10_460, i_10_629, i_10_736, i_10_796, i_10_893, i_10_895, i_10_899, i_10_1033, i_10_1034, i_10_1154, i_10_1174, i_10_1204, i_10_1205, i_10_1235, i_10_1238, i_10_1248, i_10_1249, i_10_1250, i_10_1272, i_10_1349, i_10_1450, i_10_1545, i_10_1549, i_10_1576, i_10_1627, i_10_1684, i_10_1685, i_10_1873, i_10_1874, i_10_1916, i_10_1954, i_10_1994, i_10_2057, i_10_2165, i_10_2202, i_10_2261, i_10_2336, i_10_2349, i_10_2350, i_10_2351, i_10_2363, i_10_2365, i_10_2380, i_10_2381, i_10_2383, i_10_2384, i_10_2454, i_10_2455, i_10_2465, i_10_2473, i_10_2571, i_10_2572, i_10_2633, i_10_2710, i_10_2716, i_10_2717, i_10_2722, i_10_2726, i_10_2730, i_10_2832, i_10_2869, i_10_2880, i_10_2881, i_10_2882, i_10_2920, i_10_2957, i_10_2991, i_10_3049, i_10_3072, i_10_3355, i_10_3403, i_10_3470, i_10_3571, i_10_3572, i_10_3612, i_10_3723, i_10_3724, i_10_3732, i_10_3784, i_10_3860, i_10_3981, i_10_4029, i_10_4030, i_10_4119, i_10_4129, i_10_4130, i_10_4220, i_10_4272, i_10_4289, i_10_4426, i_10_4427, i_10_4583, o_10_498);
	kernel_10_499 k_10_499(i_10_36, i_10_156, i_10_181, i_10_216, i_10_245, i_10_246, i_10_247, i_10_284, i_10_316, i_10_319, i_10_330, i_10_393, i_10_409, i_10_436, i_10_446, i_10_459, i_10_460, i_10_559, i_10_754, i_10_792, i_10_892, i_10_993, i_10_1000, i_10_1035, i_10_1039, i_10_1047, i_10_1048, i_10_1059, i_10_1152, i_10_1164, i_10_1215, i_10_1235, i_10_1237, i_10_1306, i_10_1307, i_10_1311, i_10_1312, i_10_1313, i_10_1362, i_10_1539, i_10_1575, i_10_1594, i_10_1648, i_10_1650, i_10_1655, i_10_1688, i_10_1690, i_10_1914, i_10_2016, i_10_2019, i_10_2199, i_10_2349, i_10_2356, i_10_2601, i_10_2603, i_10_2606, i_10_2634, i_10_2635, i_10_2705, i_10_2724, i_10_2728, i_10_2730, i_10_2784, i_10_2785, i_10_2831, i_10_2881, i_10_2983, i_10_2985, i_10_3073, i_10_3159, i_10_3162, i_10_3231, i_10_3270, i_10_3328, i_10_3406, i_10_3429, i_10_3430, i_10_3501, i_10_3519, i_10_3609, i_10_3610, i_10_3717, i_10_3721, i_10_3785, i_10_3787, i_10_3788, i_10_3810, i_10_3850, i_10_3856, i_10_3859, i_10_3860, i_10_3883, i_10_3889, i_10_3987, i_10_4062, i_10_4168, i_10_4173, i_10_4278, i_10_4570, i_10_4586, o_10_499);
	kernel_10_500 k_10_500(i_10_121, i_10_146, i_10_175, i_10_254, i_10_256, i_10_257, i_10_283, i_10_288, i_10_325, i_10_394, i_10_441, i_10_445, i_10_562, i_10_632, i_10_796, i_10_797, i_10_800, i_10_920, i_10_955, i_10_963, i_10_1118, i_10_1235, i_10_1236, i_10_1237, i_10_1238, i_10_1245, i_10_1249, i_10_1250, i_10_1268, i_10_1313, i_10_1361, i_10_1650, i_10_1683, i_10_1685, i_10_1687, i_10_1721, i_10_1724, i_10_1821, i_10_1824, i_10_1825, i_10_1826, i_10_1883, i_10_1915, i_10_1919, i_10_1984, i_10_2107, i_10_2243, i_10_2350, i_10_2352, i_10_2387, i_10_2390, i_10_2453, i_10_2471, i_10_2659, i_10_2663, i_10_2711, i_10_2719, i_10_2723, i_10_2737, i_10_2786, i_10_2827, i_10_2834, i_10_2846, i_10_2981, i_10_3236, i_10_3280, i_10_3283, i_10_3386, i_10_3388, i_10_3389, i_10_3431, i_10_3467, i_10_3494, i_10_3523, i_10_3524, i_10_3539, i_10_3545, i_10_3584, i_10_3586, i_10_3587, i_10_3720, i_10_3847, i_10_3872, i_10_3943, i_10_3944, i_10_3982, i_10_3998, i_10_4054, i_10_4130, i_10_4151, i_10_4231, i_10_4268, i_10_4271, i_10_4274, i_10_4275, i_10_4279, i_10_4460, i_10_4569, i_10_4571, i_10_4583, o_10_500);
	kernel_10_501 k_10_501(i_10_27, i_10_146, i_10_154, i_10_173, i_10_289, i_10_290, i_10_406, i_10_423, i_10_428, i_10_626, i_10_640, i_10_821, i_10_848, i_10_901, i_10_992, i_10_1028, i_10_1046, i_10_1118, i_10_1238, i_10_1253, i_10_1289, i_10_1442, i_10_1612, i_10_1613, i_10_1631, i_10_1648, i_10_1652, i_10_1689, i_10_1738, i_10_1757, i_10_1759, i_10_1873, i_10_1874, i_10_1954, i_10_1991, i_10_2216, i_10_2225, i_10_2288, i_10_2327, i_10_2359, i_10_2362, i_10_2441, i_10_2469, i_10_2476, i_10_2477, i_10_2511, i_10_2525, i_10_2566, i_10_2567, i_10_2603, i_10_2631, i_10_2636, i_10_2642, i_10_2648, i_10_2651, i_10_2657, i_10_2675, i_10_2719, i_10_2729, i_10_2738, i_10_2829, i_10_2833, i_10_2882, i_10_2917, i_10_2918, i_10_2923, i_10_3161, i_10_3195, i_10_3233, i_10_3286, i_10_3290, i_10_3405, i_10_3410, i_10_3440, i_10_3449, i_10_3557, i_10_3620, i_10_3686, i_10_3728, i_10_3827, i_10_3830, i_10_3852, i_10_3855, i_10_3899, i_10_4025, i_10_4028, i_10_4114, i_10_4115, i_10_4144, i_10_4145, i_10_4151, i_10_4189, i_10_4214, i_10_4291, i_10_4292, i_10_4307, i_10_4456, i_10_4501, i_10_4502, i_10_4563, o_10_501);
	kernel_10_502 k_10_502(i_10_33, i_10_34, i_10_70, i_10_179, i_10_208, i_10_248, i_10_430, i_10_431, i_10_444, i_10_448, i_10_562, i_10_563, i_10_719, i_10_796, i_10_799, i_10_820, i_10_823, i_10_953, i_10_996, i_10_1004, i_10_1006, i_10_1007, i_10_1052, i_10_1213, i_10_1247, i_10_1322, i_10_1348, i_10_1349, i_10_1366, i_10_1367, i_10_1383, i_10_1384, i_10_1492, i_10_1493, i_10_1565, i_10_1627, i_10_1628, i_10_1631, i_10_1634, i_10_1655, i_10_1697, i_10_1736, i_10_1768, i_10_1912, i_10_1937, i_10_2038, i_10_2041, i_10_2042, i_10_2159, i_10_2264, i_10_2410, i_10_2437, i_10_2474, i_10_2508, i_10_2509, i_10_2514, i_10_2517, i_10_2636, i_10_2661, i_10_2679, i_10_2698, i_10_2699, i_10_2707, i_10_2708, i_10_2714, i_10_2744, i_10_2757, i_10_2758, i_10_2824, i_10_2830, i_10_2852, i_10_2870, i_10_2885, i_10_3048, i_10_3050, i_10_3094, i_10_3095, i_10_3284, i_10_3319, i_10_3320, i_10_3415, i_10_3436, i_10_3472, i_10_3494, i_10_3588, i_10_3611, i_10_3612, i_10_3625, i_10_3640, i_10_3704, i_10_3706, i_10_3707, i_10_3853, i_10_3986, i_10_4237, i_10_4267, i_10_4268, i_10_4271, i_10_4289, i_10_4454, o_10_502);
	kernel_10_503 k_10_503(i_10_31, i_10_280, i_10_282, i_10_283, i_10_284, i_10_285, i_10_290, i_10_316, i_10_438, i_10_439, i_10_463, i_10_519, i_10_717, i_10_955, i_10_1005, i_10_1234, i_10_1235, i_10_1236, i_10_1435, i_10_1445, i_10_1648, i_10_1678, i_10_1679, i_10_1689, i_10_1819, i_10_1820, i_10_1821, i_10_1915, i_10_2027, i_10_2029, i_10_2031, i_10_2352, i_10_2353, i_10_2354, i_10_2357, i_10_2408, i_10_2449, i_10_2460, i_10_2467, i_10_2628, i_10_2630, i_10_2660, i_10_2662, i_10_2675, i_10_2711, i_10_2716, i_10_2722, i_10_2728, i_10_2729, i_10_2832, i_10_2833, i_10_2881, i_10_2885, i_10_2888, i_10_2917, i_10_2922, i_10_2923, i_10_2985, i_10_2987, i_10_3038, i_10_3040, i_10_3043, i_10_3044, i_10_3196, i_10_3198, i_10_3199, i_10_3384, i_10_3387, i_10_3388, i_10_3391, i_10_3405, i_10_3409, i_10_3497, i_10_3589, i_10_3610, i_10_3611, i_10_3614, i_10_3650, i_10_3782, i_10_3784, i_10_3785, i_10_3837, i_10_3840, i_10_3848, i_10_3858, i_10_3859, i_10_3907, i_10_4025, i_10_4123, i_10_4124, i_10_4127, i_10_4269, i_10_4270, i_10_4271, i_10_4278, i_10_4286, i_10_4292, i_10_4567, i_10_4568, i_10_4569, o_10_503);
	kernel_10_504 k_10_504(i_10_175, i_10_176, i_10_186, i_10_187, i_10_188, i_10_282, i_10_409, i_10_464, i_10_467, i_10_516, i_10_1165, i_10_1169, i_10_1236, i_10_1249, i_10_1348, i_10_1435, i_10_1552, i_10_1556, i_10_1823, i_10_1824, i_10_1826, i_10_1947, i_10_1993, i_10_2021, i_10_2309, i_10_2350, i_10_2353, i_10_2450, i_10_2453, i_10_2467, i_10_2470, i_10_2514, i_10_2517, i_10_2571, i_10_2572, i_10_2633, i_10_2704, i_10_2708, i_10_2713, i_10_2714, i_10_2716, i_10_2717, i_10_2722, i_10_2727, i_10_2728, i_10_2823, i_10_2831, i_10_2870, i_10_2883, i_10_2884, i_10_2885, i_10_2886, i_10_2887, i_10_2921, i_10_2953, i_10_2981, i_10_3037, i_10_3038, i_10_3047, i_10_3074, i_10_3198, i_10_3271, i_10_3272, i_10_3274, i_10_3281, i_10_3386, i_10_3407, i_10_3434, i_10_3611, i_10_3614, i_10_3653, i_10_3720, i_10_3771, i_10_3783, i_10_3784, i_10_3785, i_10_3839, i_10_3853, i_10_3855, i_10_3856, i_10_3857, i_10_3880, i_10_3885, i_10_3886, i_10_3890, i_10_3895, i_10_3896, i_10_3984, i_10_3985, i_10_4051, i_10_4119, i_10_4120, i_10_4172, i_10_4175, i_10_4189, i_10_4190, i_10_4191, i_10_4291, i_10_4462, i_10_4571, o_10_504);
	kernel_10_505 k_10_505(i_10_178, i_10_254, i_10_260, i_10_266, i_10_277, i_10_280, i_10_283, i_10_287, i_10_319, i_10_407, i_10_442, i_10_497, i_10_503, i_10_506, i_10_509, i_10_512, i_10_866, i_10_869, i_10_1007, i_10_1083, i_10_1085, i_10_1086, i_10_1102, i_10_1237, i_10_1238, i_10_1250, i_10_1297, i_10_1301, i_10_1303, i_10_1307, i_10_1540, i_10_1541, i_10_1621, i_10_1622, i_10_1626, i_10_1686, i_10_1687, i_10_1688, i_10_1764, i_10_1798, i_10_1807, i_10_1984, i_10_2027, i_10_2030, i_10_2032, i_10_2033, i_10_2091, i_10_2110, i_10_2182, i_10_2203, i_10_2354, i_10_2456, i_10_2471, i_10_2516, i_10_2656, i_10_2701, i_10_2702, i_10_2703, i_10_2722, i_10_2728, i_10_2729, i_10_2731, i_10_2734, i_10_2735, i_10_2965, i_10_2968, i_10_2969, i_10_2984, i_10_3046, i_10_3314, i_10_3317, i_10_3391, i_10_3392, i_10_3409, i_10_3410, i_10_3467, i_10_3470, i_10_3494, i_10_3506, i_10_3525, i_10_3538, i_10_3587, i_10_3682, i_10_3837, i_10_3840, i_10_3844, i_10_3850, i_10_3895, i_10_3982, i_10_4114, i_10_4188, i_10_4208, i_10_4268, i_10_4271, i_10_4274, i_10_4283, i_10_4285, i_10_4288, i_10_4292, i_10_4569, o_10_505);
	kernel_10_506 k_10_506(i_10_67, i_10_147, i_10_151, i_10_175, i_10_190, i_10_220, i_10_318, i_10_319, i_10_364, i_10_372, i_10_410, i_10_475, i_10_595, i_10_690, i_10_733, i_10_876, i_10_1000, i_10_1011, i_10_1069, i_10_1083, i_10_1099, i_10_1110, i_10_1278, i_10_1293, i_10_1308, i_10_1309, i_10_1443, i_10_1596, i_10_1619, i_10_1621, i_10_1623, i_10_1624, i_10_1635, i_10_1636, i_10_1647, i_10_1651, i_10_1818, i_10_1821, i_10_1822, i_10_1849, i_10_1918, i_10_1956, i_10_1959, i_10_1965, i_10_1987, i_10_2109, i_10_2112, i_10_2226, i_10_2305, i_10_2353, i_10_2481, i_10_2482, i_10_2516, i_10_2540, i_10_2561, i_10_2569, i_10_2588, i_10_2659, i_10_2677, i_10_2680, i_10_2686, i_10_2713, i_10_2778, i_10_2785, i_10_2884, i_10_2952, i_10_2953, i_10_2956, i_10_2980, i_10_2990, i_10_3040, i_10_3276, i_10_3283, i_10_3297, i_10_3324, i_10_3325, i_10_3450, i_10_3454, i_10_3550, i_10_3585, i_10_3649, i_10_3704, i_10_3779, i_10_3838, i_10_3853, i_10_3854, i_10_3896, i_10_4028, i_10_4057, i_10_4118, i_10_4120, i_10_4168, i_10_4279, i_10_4317, i_10_4380, i_10_4459, i_10_4546, i_10_4570, i_10_4582, i_10_4585, o_10_506);
	kernel_10_507 k_10_507(i_10_35, i_10_118, i_10_119, i_10_124, i_10_125, i_10_175, i_10_268, i_10_284, i_10_368, i_10_391, i_10_440, i_10_461, i_10_464, i_10_521, i_10_566, i_10_588, i_10_589, i_10_590, i_10_831, i_10_832, i_10_833, i_10_899, i_10_962, i_10_963, i_10_997, i_10_1007, i_10_1055, i_10_1166, i_10_1310, i_10_1348, i_10_1367, i_10_1382, i_10_1435, i_10_1436, i_10_1438, i_10_1439, i_10_1456, i_10_1457, i_10_1616, i_10_1618, i_10_1619, i_10_1636, i_10_1689, i_10_1822, i_10_1823, i_10_1922, i_10_1948, i_10_1952, i_10_1986, i_10_2006, i_10_2213, i_10_2244, i_10_2356, i_10_2408, i_10_2409, i_10_2430, i_10_2454, i_10_2515, i_10_2516, i_10_2617, i_10_2618, i_10_2628, i_10_2629, i_10_2633, i_10_2660, i_10_2681, i_10_2713, i_10_2731, i_10_2732, i_10_2882, i_10_2920, i_10_2924, i_10_3040, i_10_3041, i_10_3043, i_10_3094, i_10_3117, i_10_3122, i_10_3200, i_10_3351, i_10_3391, i_10_3526, i_10_3542, i_10_3580, i_10_3587, i_10_3610, i_10_3613, i_10_3625, i_10_3647, i_10_3649, i_10_3652, i_10_3653, i_10_3783, i_10_3837, i_10_3838, i_10_3895, i_10_3985, i_10_4001, i_10_4172, i_10_4373, o_10_507);
	kernel_10_508 k_10_508(i_10_171, i_10_174, i_10_179, i_10_221, i_10_245, i_10_280, i_10_433, i_10_435, i_10_436, i_10_437, i_10_439, i_10_440, i_10_444, i_10_749, i_10_797, i_10_1001, i_10_1005, i_10_1166, i_10_1234, i_10_1235, i_10_1246, i_10_1249, i_10_1250, i_10_1309, i_10_1310, i_10_1550, i_10_1649, i_10_1652, i_10_1684, i_10_1686, i_10_1687, i_10_1819, i_10_1822, i_10_1823, i_10_1825, i_10_1946, i_10_2179, i_10_2180, i_10_2306, i_10_2357, i_10_2365, i_10_2384, i_10_2470, i_10_2471, i_10_2516, i_10_2629, i_10_2631, i_10_2633, i_10_2659, i_10_2675, i_10_2708, i_10_2723, i_10_2727, i_10_2731, i_10_2830, i_10_2884, i_10_2885, i_10_2887, i_10_2917, i_10_2918, i_10_3150, i_10_3151, i_10_3152, i_10_3200, i_10_3238, i_10_3268, i_10_3269, i_10_3274, i_10_3322, i_10_3390, i_10_3391, i_10_3406, i_10_3407, i_10_3410, i_10_3470, i_10_3590, i_10_3610, i_10_3613, i_10_3614, i_10_3784, i_10_3835, i_10_3837, i_10_3838, i_10_3839, i_10_3841, i_10_3846, i_10_3847, i_10_3848, i_10_3849, i_10_3850, i_10_3853, i_10_3855, i_10_3859, i_10_3979, i_10_3986, i_10_4117, i_10_4123, i_10_4285, i_10_4287, i_10_4567, o_10_508);
	kernel_10_509 k_10_509(i_10_34, i_10_150, i_10_172, i_10_174, i_10_175, i_10_435, i_10_438, i_10_444, i_10_447, i_10_448, i_10_462, i_10_467, i_10_508, i_10_516, i_10_519, i_10_717, i_10_799, i_10_966, i_10_967, i_10_996, i_10_1029, i_10_1141, i_10_1164, i_10_1240, i_10_1245, i_10_1248, i_10_1309, i_10_1311, i_10_1366, i_10_1626, i_10_1652, i_10_1653, i_10_1655, i_10_1689, i_10_1690, i_10_1797, i_10_1821, i_10_1822, i_10_1912, i_10_1995, i_10_2005, i_10_2352, i_10_2353, i_10_2455, i_10_2469, i_10_2472, i_10_2473, i_10_2571, i_10_2628, i_10_2629, i_10_2659, i_10_2661, i_10_2706, i_10_2715, i_10_2716, i_10_2722, i_10_2731, i_10_2734, i_10_2742, i_10_2782, i_10_2830, i_10_2832, i_10_2883, i_10_2987, i_10_3037, i_10_3039, i_10_3046, i_10_3048, i_10_3075, i_10_3093, i_10_3157, i_10_3197, i_10_3284, i_10_3321, i_10_3322, i_10_3327, i_10_3391, i_10_3392, i_10_3468, i_10_3495, i_10_3525, i_10_3583, i_10_3585, i_10_3612, i_10_3613, i_10_3732, i_10_3780, i_10_3837, i_10_3876, i_10_3912, i_10_3982, i_10_4113, i_10_4173, i_10_4269, i_10_4272, i_10_4273, i_10_4282, i_10_4290, i_10_4317, i_10_4566, o_10_509);
	kernel_10_510 k_10_510(i_10_35, i_10_71, i_10_124, i_10_125, i_10_154, i_10_178, i_10_215, i_10_265, i_10_279, i_10_317, i_10_390, i_10_410, i_10_440, i_10_445, i_10_465, i_10_533, i_10_562, i_10_565, i_10_566, i_10_869, i_10_1000, i_10_1006, i_10_1163, i_10_1265, i_10_1277, i_10_1319, i_10_1361, i_10_1363, i_10_1438, i_10_1439, i_10_1525, i_10_1652, i_10_1654, i_10_1714, i_10_1769, i_10_1823, i_10_1913, i_10_1922, i_10_1951, i_10_1952, i_10_2023, i_10_2033, i_10_2083, i_10_2096, i_10_2186, i_10_2200, i_10_2201, i_10_2203, i_10_2237, i_10_2240, i_10_2257, i_10_2312, i_10_2363, i_10_2378, i_10_2453, i_10_2470, i_10_2514, i_10_2614, i_10_2615, i_10_2633, i_10_2636, i_10_2786, i_10_2831, i_10_2881, i_10_2924, i_10_2960, i_10_2980, i_10_2986, i_10_3039, i_10_3040, i_10_3041, i_10_3046, i_10_3070, i_10_3071, i_10_3073, i_10_3159, i_10_3160, i_10_3434, i_10_3448, i_10_3469, i_10_3470, i_10_3520, i_10_3544, i_10_3545, i_10_3562, i_10_3563, i_10_3586, i_10_3590, i_10_3647, i_10_3652, i_10_3653, i_10_3682, i_10_3685, i_10_3788, i_10_4167, i_10_4168, i_10_4169, i_10_4234, i_10_4278, i_10_4531, o_10_510);
	kernel_10_511 k_10_511(i_10_174, i_10_248, i_10_266, i_10_270, i_10_273, i_10_274, i_10_284, i_10_285, i_10_293, i_10_395, i_10_500, i_10_503, i_10_629, i_10_797, i_10_1003, i_10_1004, i_10_1086, i_10_1105, i_10_1115, i_10_1120, i_10_1138, i_10_1223, i_10_1238, i_10_1240, i_10_1241, i_10_1301, i_10_1303, i_10_1384, i_10_1436, i_10_1544, i_10_1545, i_10_1547, i_10_1578, i_10_1581, i_10_1582, i_10_1625, i_10_1628, i_10_1651, i_10_1690, i_10_1691, i_10_1733, i_10_1736, i_10_1824, i_10_2003, i_10_2006, i_10_2030, i_10_2033, i_10_2200, i_10_2354, i_10_2363, i_10_2453, i_10_2462, i_10_2471, i_10_2473, i_10_2474, i_10_2510, i_10_2570, i_10_2573, i_10_2631, i_10_2632, i_10_2633, i_10_2634, i_10_2635, i_10_2636, i_10_2641, i_10_2644, i_10_2701, i_10_2705, i_10_2717, i_10_2785, i_10_2830, i_10_2834, i_10_2849, i_10_2882, i_10_2883, i_10_3071, i_10_3278, i_10_3281, i_10_3384, i_10_3388, i_10_3392, i_10_3408, i_10_3470, i_10_3473, i_10_3542, i_10_3545, i_10_3584, i_10_3587, i_10_3613, i_10_3784, i_10_3838, i_10_3839, i_10_3843, i_10_3853, i_10_3854, i_10_4113, i_10_4126, i_10_4127, i_10_4283, i_10_4589, o_10_511);
endmodule


module kernel_10_wrapper (input ap_clk, ap_rst, ap_ce, ap_start, ap_continue,
                        input [4607:0] in_reg,
                        output ap_idle, ap_done, ap_ready,
                        output out_reg_ap_vld,
                        output reg [511:0] out_reg);

  wire ce = ap_ce;
  reg i_10_0, i_10_1, i_10_2, i_10_3, i_10_4, i_10_5, i_10_6, i_10_7, i_10_8, i_10_9, i_10_10, i_10_11, i_10_12, i_10_13, i_10_14, i_10_15, i_10_16, i_10_17, i_10_18, i_10_19, i_10_20, i_10_21, i_10_22, i_10_23, i_10_24, i_10_25, i_10_26, i_10_27, i_10_28, i_10_29, i_10_30, i_10_31, i_10_32, i_10_33, i_10_34, i_10_35, i_10_36, i_10_37, i_10_38, i_10_39, i_10_40, i_10_41, i_10_42, i_10_43, i_10_44, i_10_45, i_10_46, i_10_47, i_10_48, i_10_49, i_10_50, i_10_51, i_10_52, i_10_53, i_10_54, i_10_55, i_10_56, i_10_57, i_10_58, i_10_59, i_10_60, i_10_61, i_10_62, i_10_63, i_10_64, i_10_65, i_10_66, i_10_67, i_10_68, i_10_69, i_10_70, i_10_71, i_10_72, i_10_73, i_10_74, i_10_75, i_10_76, i_10_77, i_10_78, i_10_79, i_10_80, i_10_81, i_10_82, i_10_83, i_10_84, i_10_85, i_10_86, i_10_87, i_10_88, i_10_89, i_10_90, i_10_91, i_10_92, i_10_93, i_10_94, i_10_95, i_10_96, i_10_97, i_10_98, i_10_99, i_10_100, i_10_101, i_10_102, i_10_103, i_10_104, i_10_105, i_10_106, i_10_107, i_10_108, i_10_109, i_10_110, i_10_111, i_10_112, i_10_113, i_10_114, i_10_115, i_10_116, i_10_117, i_10_118, i_10_119, i_10_120, i_10_121, i_10_122, i_10_123, i_10_124, i_10_125, i_10_126, i_10_127, i_10_128, i_10_129, i_10_130, i_10_131, i_10_132, i_10_133, i_10_134, i_10_135, i_10_136, i_10_137, i_10_138, i_10_139, i_10_140, i_10_141, i_10_142, i_10_143, i_10_144, i_10_145, i_10_146, i_10_147, i_10_148, i_10_149, i_10_150, i_10_151, i_10_152, i_10_153, i_10_154, i_10_155, i_10_156, i_10_157, i_10_158, i_10_159, i_10_160, i_10_161, i_10_162, i_10_163, i_10_164, i_10_165, i_10_166, i_10_167, i_10_168, i_10_169, i_10_170, i_10_171, i_10_172, i_10_173, i_10_174, i_10_175, i_10_176, i_10_177, i_10_178, i_10_179, i_10_180, i_10_181, i_10_182, i_10_183, i_10_184, i_10_185, i_10_186, i_10_187, i_10_188, i_10_189, i_10_190, i_10_191, i_10_192, i_10_193, i_10_194, i_10_195, i_10_196, i_10_197, i_10_198, i_10_199, i_10_200, i_10_201, i_10_202, i_10_203, i_10_204, i_10_205, i_10_206, i_10_207, i_10_208, i_10_209, i_10_210, i_10_211, i_10_212, i_10_213, i_10_214, i_10_215, i_10_216, i_10_217, i_10_218, i_10_219, i_10_220, i_10_221, i_10_222, i_10_223, i_10_224, i_10_225, i_10_226, i_10_227, i_10_228, i_10_229, i_10_230, i_10_231, i_10_232, i_10_233, i_10_234, i_10_235, i_10_236, i_10_237, i_10_238, i_10_239, i_10_240, i_10_241, i_10_242, i_10_243, i_10_244, i_10_245, i_10_246, i_10_247, i_10_248, i_10_249, i_10_250, i_10_251, i_10_252, i_10_253, i_10_254, i_10_255, i_10_256, i_10_257, i_10_258, i_10_259, i_10_260, i_10_261, i_10_262, i_10_263, i_10_264, i_10_265, i_10_266, i_10_267, i_10_268, i_10_269, i_10_270, i_10_271, i_10_272, i_10_273, i_10_274, i_10_275, i_10_276, i_10_277, i_10_278, i_10_279, i_10_280, i_10_281, i_10_282, i_10_283, i_10_284, i_10_285, i_10_286, i_10_287, i_10_288, i_10_289, i_10_290, i_10_291, i_10_292, i_10_293, i_10_294, i_10_295, i_10_296, i_10_297, i_10_298, i_10_299, i_10_300, i_10_301, i_10_302, i_10_303, i_10_304, i_10_305, i_10_306, i_10_307, i_10_308, i_10_309, i_10_310, i_10_311, i_10_312, i_10_313, i_10_314, i_10_315, i_10_316, i_10_317, i_10_318, i_10_319, i_10_320, i_10_321, i_10_322, i_10_323, i_10_324, i_10_325, i_10_326, i_10_327, i_10_328, i_10_329, i_10_330, i_10_331, i_10_332, i_10_333, i_10_334, i_10_335, i_10_336, i_10_337, i_10_338, i_10_339, i_10_340, i_10_341, i_10_342, i_10_343, i_10_344, i_10_345, i_10_346, i_10_347, i_10_348, i_10_349, i_10_350, i_10_351, i_10_352, i_10_353, i_10_354, i_10_355, i_10_356, i_10_357, i_10_358, i_10_359, i_10_360, i_10_361, i_10_362, i_10_363, i_10_364, i_10_365, i_10_366, i_10_367, i_10_368, i_10_369, i_10_370, i_10_371, i_10_372, i_10_373, i_10_374, i_10_375, i_10_376, i_10_377, i_10_378, i_10_379, i_10_380, i_10_381, i_10_382, i_10_383, i_10_384, i_10_385, i_10_386, i_10_387, i_10_388, i_10_389, i_10_390, i_10_391, i_10_392, i_10_393, i_10_394, i_10_395, i_10_396, i_10_397, i_10_398, i_10_399, i_10_400, i_10_401, i_10_402, i_10_403, i_10_404, i_10_405, i_10_406, i_10_407, i_10_408, i_10_409, i_10_410, i_10_411, i_10_412, i_10_413, i_10_414, i_10_415, i_10_416, i_10_417, i_10_418, i_10_419, i_10_420, i_10_421, i_10_422, i_10_423, i_10_424, i_10_425, i_10_426, i_10_427, i_10_428, i_10_429, i_10_430, i_10_431, i_10_432, i_10_433, i_10_434, i_10_435, i_10_436, i_10_437, i_10_438, i_10_439, i_10_440, i_10_441, i_10_442, i_10_443, i_10_444, i_10_445, i_10_446, i_10_447, i_10_448, i_10_449, i_10_450, i_10_451, i_10_452, i_10_453, i_10_454, i_10_455, i_10_456, i_10_457, i_10_458, i_10_459, i_10_460, i_10_461, i_10_462, i_10_463, i_10_464, i_10_465, i_10_466, i_10_467, i_10_468, i_10_469, i_10_470, i_10_471, i_10_472, i_10_473, i_10_474, i_10_475, i_10_476, i_10_477, i_10_478, i_10_479, i_10_480, i_10_481, i_10_482, i_10_483, i_10_484, i_10_485, i_10_486, i_10_487, i_10_488, i_10_489, i_10_490, i_10_491, i_10_492, i_10_493, i_10_494, i_10_495, i_10_496, i_10_497, i_10_498, i_10_499, i_10_500, i_10_501, i_10_502, i_10_503, i_10_504, i_10_505, i_10_506, i_10_507, i_10_508, i_10_509, i_10_510, i_10_511, i_10_512, i_10_513, i_10_514, i_10_515, i_10_516, i_10_517, i_10_518, i_10_519, i_10_520, i_10_521, i_10_522, i_10_523, i_10_524, i_10_525, i_10_526, i_10_527, i_10_528, i_10_529, i_10_530, i_10_531, i_10_532, i_10_533, i_10_534, i_10_535, i_10_536, i_10_537, i_10_538, i_10_539, i_10_540, i_10_541, i_10_542, i_10_543, i_10_544, i_10_545, i_10_546, i_10_547, i_10_548, i_10_549, i_10_550, i_10_551, i_10_552, i_10_553, i_10_554, i_10_555, i_10_556, i_10_557, i_10_558, i_10_559, i_10_560, i_10_561, i_10_562, i_10_563, i_10_564, i_10_565, i_10_566, i_10_567, i_10_568, i_10_569, i_10_570, i_10_571, i_10_572, i_10_573, i_10_574, i_10_575, i_10_576, i_10_577, i_10_578, i_10_579, i_10_580, i_10_581, i_10_582, i_10_583, i_10_584, i_10_585, i_10_586, i_10_587, i_10_588, i_10_589, i_10_590, i_10_591, i_10_592, i_10_593, i_10_594, i_10_595, i_10_596, i_10_597, i_10_598, i_10_599, i_10_600, i_10_601, i_10_602, i_10_603, i_10_604, i_10_605, i_10_606, i_10_607, i_10_608, i_10_609, i_10_610, i_10_611, i_10_612, i_10_613, i_10_614, i_10_615, i_10_616, i_10_617, i_10_618, i_10_619, i_10_620, i_10_621, i_10_622, i_10_623, i_10_624, i_10_625, i_10_626, i_10_627, i_10_628, i_10_629, i_10_630, i_10_631, i_10_632, i_10_633, i_10_634, i_10_635, i_10_636, i_10_637, i_10_638, i_10_639, i_10_640, i_10_641, i_10_642, i_10_643, i_10_644, i_10_645, i_10_646, i_10_647, i_10_648, i_10_649, i_10_650, i_10_651, i_10_652, i_10_653, i_10_654, i_10_655, i_10_656, i_10_657, i_10_658, i_10_659, i_10_660, i_10_661, i_10_662, i_10_663, i_10_664, i_10_665, i_10_666, i_10_667, i_10_668, i_10_669, i_10_670, i_10_671, i_10_672, i_10_673, i_10_674, i_10_675, i_10_676, i_10_677, i_10_678, i_10_679, i_10_680, i_10_681, i_10_682, i_10_683, i_10_684, i_10_685, i_10_686, i_10_687, i_10_688, i_10_689, i_10_690, i_10_691, i_10_692, i_10_693, i_10_694, i_10_695, i_10_696, i_10_697, i_10_698, i_10_699, i_10_700, i_10_701, i_10_702, i_10_703, i_10_704, i_10_705, i_10_706, i_10_707, i_10_708, i_10_709, i_10_710, i_10_711, i_10_712, i_10_713, i_10_714, i_10_715, i_10_716, i_10_717, i_10_718, i_10_719, i_10_720, i_10_721, i_10_722, i_10_723, i_10_724, i_10_725, i_10_726, i_10_727, i_10_728, i_10_729, i_10_730, i_10_731, i_10_732, i_10_733, i_10_734, i_10_735, i_10_736, i_10_737, i_10_738, i_10_739, i_10_740, i_10_741, i_10_742, i_10_743, i_10_744, i_10_745, i_10_746, i_10_747, i_10_748, i_10_749, i_10_750, i_10_751, i_10_752, i_10_753, i_10_754, i_10_755, i_10_756, i_10_757, i_10_758, i_10_759, i_10_760, i_10_761, i_10_762, i_10_763, i_10_764, i_10_765, i_10_766, i_10_767, i_10_768, i_10_769, i_10_770, i_10_771, i_10_772, i_10_773, i_10_774, i_10_775, i_10_776, i_10_777, i_10_778, i_10_779, i_10_780, i_10_781, i_10_782, i_10_783, i_10_784, i_10_785, i_10_786, i_10_787, i_10_788, i_10_789, i_10_790, i_10_791, i_10_792, i_10_793, i_10_794, i_10_795, i_10_796, i_10_797, i_10_798, i_10_799, i_10_800, i_10_801, i_10_802, i_10_803, i_10_804, i_10_805, i_10_806, i_10_807, i_10_808, i_10_809, i_10_810, i_10_811, i_10_812, i_10_813, i_10_814, i_10_815, i_10_816, i_10_817, i_10_818, i_10_819, i_10_820, i_10_821, i_10_822, i_10_823, i_10_824, i_10_825, i_10_826, i_10_827, i_10_828, i_10_829, i_10_830, i_10_831, i_10_832, i_10_833, i_10_834, i_10_835, i_10_836, i_10_837, i_10_838, i_10_839, i_10_840, i_10_841, i_10_842, i_10_843, i_10_844, i_10_845, i_10_846, i_10_847, i_10_848, i_10_849, i_10_850, i_10_851, i_10_852, i_10_853, i_10_854, i_10_855, i_10_856, i_10_857, i_10_858, i_10_859, i_10_860, i_10_861, i_10_862, i_10_863, i_10_864, i_10_865, i_10_866, i_10_867, i_10_868, i_10_869, i_10_870, i_10_871, i_10_872, i_10_873, i_10_874, i_10_875, i_10_876, i_10_877, i_10_878, i_10_879, i_10_880, i_10_881, i_10_882, i_10_883, i_10_884, i_10_885, i_10_886, i_10_887, i_10_888, i_10_889, i_10_890, i_10_891, i_10_892, i_10_893, i_10_894, i_10_895, i_10_896, i_10_897, i_10_898, i_10_899, i_10_900, i_10_901, i_10_902, i_10_903, i_10_904, i_10_905, i_10_906, i_10_907, i_10_908, i_10_909, i_10_910, i_10_911, i_10_912, i_10_913, i_10_914, i_10_915, i_10_916, i_10_917, i_10_918, i_10_919, i_10_920, i_10_921, i_10_922, i_10_923, i_10_924, i_10_925, i_10_926, i_10_927, i_10_928, i_10_929, i_10_930, i_10_931, i_10_932, i_10_933, i_10_934, i_10_935, i_10_936, i_10_937, i_10_938, i_10_939, i_10_940, i_10_941, i_10_942, i_10_943, i_10_944, i_10_945, i_10_946, i_10_947, i_10_948, i_10_949, i_10_950, i_10_951, i_10_952, i_10_953, i_10_954, i_10_955, i_10_956, i_10_957, i_10_958, i_10_959, i_10_960, i_10_961, i_10_962, i_10_963, i_10_964, i_10_965, i_10_966, i_10_967, i_10_968, i_10_969, i_10_970, i_10_971, i_10_972, i_10_973, i_10_974, i_10_975, i_10_976, i_10_977, i_10_978, i_10_979, i_10_980, i_10_981, i_10_982, i_10_983, i_10_984, i_10_985, i_10_986, i_10_987, i_10_988, i_10_989, i_10_990, i_10_991, i_10_992, i_10_993, i_10_994, i_10_995, i_10_996, i_10_997, i_10_998, i_10_999, i_10_1000, i_10_1001, i_10_1002, i_10_1003, i_10_1004, i_10_1005, i_10_1006, i_10_1007, i_10_1008, i_10_1009, i_10_1010, i_10_1011, i_10_1012, i_10_1013, i_10_1014, i_10_1015, i_10_1016, i_10_1017, i_10_1018, i_10_1019, i_10_1020, i_10_1021, i_10_1022, i_10_1023, i_10_1024, i_10_1025, i_10_1026, i_10_1027, i_10_1028, i_10_1029, i_10_1030, i_10_1031, i_10_1032, i_10_1033, i_10_1034, i_10_1035, i_10_1036, i_10_1037, i_10_1038, i_10_1039, i_10_1040, i_10_1041, i_10_1042, i_10_1043, i_10_1044, i_10_1045, i_10_1046, i_10_1047, i_10_1048, i_10_1049, i_10_1050, i_10_1051, i_10_1052, i_10_1053, i_10_1054, i_10_1055, i_10_1056, i_10_1057, i_10_1058, i_10_1059, i_10_1060, i_10_1061, i_10_1062, i_10_1063, i_10_1064, i_10_1065, i_10_1066, i_10_1067, i_10_1068, i_10_1069, i_10_1070, i_10_1071, i_10_1072, i_10_1073, i_10_1074, i_10_1075, i_10_1076, i_10_1077, i_10_1078, i_10_1079, i_10_1080, i_10_1081, i_10_1082, i_10_1083, i_10_1084, i_10_1085, i_10_1086, i_10_1087, i_10_1088, i_10_1089, i_10_1090, i_10_1091, i_10_1092, i_10_1093, i_10_1094, i_10_1095, i_10_1096, i_10_1097, i_10_1098, i_10_1099, i_10_1100, i_10_1101, i_10_1102, i_10_1103, i_10_1104, i_10_1105, i_10_1106, i_10_1107, i_10_1108, i_10_1109, i_10_1110, i_10_1111, i_10_1112, i_10_1113, i_10_1114, i_10_1115, i_10_1116, i_10_1117, i_10_1118, i_10_1119, i_10_1120, i_10_1121, i_10_1122, i_10_1123, i_10_1124, i_10_1125, i_10_1126, i_10_1127, i_10_1128, i_10_1129, i_10_1130, i_10_1131, i_10_1132, i_10_1133, i_10_1134, i_10_1135, i_10_1136, i_10_1137, i_10_1138, i_10_1139, i_10_1140, i_10_1141, i_10_1142, i_10_1143, i_10_1144, i_10_1145, i_10_1146, i_10_1147, i_10_1148, i_10_1149, i_10_1150, i_10_1151, i_10_1152, i_10_1153, i_10_1154, i_10_1155, i_10_1156, i_10_1157, i_10_1158, i_10_1159, i_10_1160, i_10_1161, i_10_1162, i_10_1163, i_10_1164, i_10_1165, i_10_1166, i_10_1167, i_10_1168, i_10_1169, i_10_1170, i_10_1171, i_10_1172, i_10_1173, i_10_1174, i_10_1175, i_10_1176, i_10_1177, i_10_1178, i_10_1179, i_10_1180, i_10_1181, i_10_1182, i_10_1183, i_10_1184, i_10_1185, i_10_1186, i_10_1187, i_10_1188, i_10_1189, i_10_1190, i_10_1191, i_10_1192, i_10_1193, i_10_1194, i_10_1195, i_10_1196, i_10_1197, i_10_1198, i_10_1199, i_10_1200, i_10_1201, i_10_1202, i_10_1203, i_10_1204, i_10_1205, i_10_1206, i_10_1207, i_10_1208, i_10_1209, i_10_1210, i_10_1211, i_10_1212, i_10_1213, i_10_1214, i_10_1215, i_10_1216, i_10_1217, i_10_1218, i_10_1219, i_10_1220, i_10_1221, i_10_1222, i_10_1223, i_10_1224, i_10_1225, i_10_1226, i_10_1227, i_10_1228, i_10_1229, i_10_1230, i_10_1231, i_10_1232, i_10_1233, i_10_1234, i_10_1235, i_10_1236, i_10_1237, i_10_1238, i_10_1239, i_10_1240, i_10_1241, i_10_1242, i_10_1243, i_10_1244, i_10_1245, i_10_1246, i_10_1247, i_10_1248, i_10_1249, i_10_1250, i_10_1251, i_10_1252, i_10_1253, i_10_1254, i_10_1255, i_10_1256, i_10_1257, i_10_1258, i_10_1259, i_10_1260, i_10_1261, i_10_1262, i_10_1263, i_10_1264, i_10_1265, i_10_1266, i_10_1267, i_10_1268, i_10_1269, i_10_1270, i_10_1271, i_10_1272, i_10_1273, i_10_1274, i_10_1275, i_10_1276, i_10_1277, i_10_1278, i_10_1279, i_10_1280, i_10_1281, i_10_1282, i_10_1283, i_10_1284, i_10_1285, i_10_1286, i_10_1287, i_10_1288, i_10_1289, i_10_1290, i_10_1291, i_10_1292, i_10_1293, i_10_1294, i_10_1295, i_10_1296, i_10_1297, i_10_1298, i_10_1299, i_10_1300, i_10_1301, i_10_1302, i_10_1303, i_10_1304, i_10_1305, i_10_1306, i_10_1307, i_10_1308, i_10_1309, i_10_1310, i_10_1311, i_10_1312, i_10_1313, i_10_1314, i_10_1315, i_10_1316, i_10_1317, i_10_1318, i_10_1319, i_10_1320, i_10_1321, i_10_1322, i_10_1323, i_10_1324, i_10_1325, i_10_1326, i_10_1327, i_10_1328, i_10_1329, i_10_1330, i_10_1331, i_10_1332, i_10_1333, i_10_1334, i_10_1335, i_10_1336, i_10_1337, i_10_1338, i_10_1339, i_10_1340, i_10_1341, i_10_1342, i_10_1343, i_10_1344, i_10_1345, i_10_1346, i_10_1347, i_10_1348, i_10_1349, i_10_1350, i_10_1351, i_10_1352, i_10_1353, i_10_1354, i_10_1355, i_10_1356, i_10_1357, i_10_1358, i_10_1359, i_10_1360, i_10_1361, i_10_1362, i_10_1363, i_10_1364, i_10_1365, i_10_1366, i_10_1367, i_10_1368, i_10_1369, i_10_1370, i_10_1371, i_10_1372, i_10_1373, i_10_1374, i_10_1375, i_10_1376, i_10_1377, i_10_1378, i_10_1379, i_10_1380, i_10_1381, i_10_1382, i_10_1383, i_10_1384, i_10_1385, i_10_1386, i_10_1387, i_10_1388, i_10_1389, i_10_1390, i_10_1391, i_10_1392, i_10_1393, i_10_1394, i_10_1395, i_10_1396, i_10_1397, i_10_1398, i_10_1399, i_10_1400, i_10_1401, i_10_1402, i_10_1403, i_10_1404, i_10_1405, i_10_1406, i_10_1407, i_10_1408, i_10_1409, i_10_1410, i_10_1411, i_10_1412, i_10_1413, i_10_1414, i_10_1415, i_10_1416, i_10_1417, i_10_1418, i_10_1419, i_10_1420, i_10_1421, i_10_1422, i_10_1423, i_10_1424, i_10_1425, i_10_1426, i_10_1427, i_10_1428, i_10_1429, i_10_1430, i_10_1431, i_10_1432, i_10_1433, i_10_1434, i_10_1435, i_10_1436, i_10_1437, i_10_1438, i_10_1439, i_10_1440, i_10_1441, i_10_1442, i_10_1443, i_10_1444, i_10_1445, i_10_1446, i_10_1447, i_10_1448, i_10_1449, i_10_1450, i_10_1451, i_10_1452, i_10_1453, i_10_1454, i_10_1455, i_10_1456, i_10_1457, i_10_1458, i_10_1459, i_10_1460, i_10_1461, i_10_1462, i_10_1463, i_10_1464, i_10_1465, i_10_1466, i_10_1467, i_10_1468, i_10_1469, i_10_1470, i_10_1471, i_10_1472, i_10_1473, i_10_1474, i_10_1475, i_10_1476, i_10_1477, i_10_1478, i_10_1479, i_10_1480, i_10_1481, i_10_1482, i_10_1483, i_10_1484, i_10_1485, i_10_1486, i_10_1487, i_10_1488, i_10_1489, i_10_1490, i_10_1491, i_10_1492, i_10_1493, i_10_1494, i_10_1495, i_10_1496, i_10_1497, i_10_1498, i_10_1499, i_10_1500, i_10_1501, i_10_1502, i_10_1503, i_10_1504, i_10_1505, i_10_1506, i_10_1507, i_10_1508, i_10_1509, i_10_1510, i_10_1511, i_10_1512, i_10_1513, i_10_1514, i_10_1515, i_10_1516, i_10_1517, i_10_1518, i_10_1519, i_10_1520, i_10_1521, i_10_1522, i_10_1523, i_10_1524, i_10_1525, i_10_1526, i_10_1527, i_10_1528, i_10_1529, i_10_1530, i_10_1531, i_10_1532, i_10_1533, i_10_1534, i_10_1535, i_10_1536, i_10_1537, i_10_1538, i_10_1539, i_10_1540, i_10_1541, i_10_1542, i_10_1543, i_10_1544, i_10_1545, i_10_1546, i_10_1547, i_10_1548, i_10_1549, i_10_1550, i_10_1551, i_10_1552, i_10_1553, i_10_1554, i_10_1555, i_10_1556, i_10_1557, i_10_1558, i_10_1559, i_10_1560, i_10_1561, i_10_1562, i_10_1563, i_10_1564, i_10_1565, i_10_1566, i_10_1567, i_10_1568, i_10_1569, i_10_1570, i_10_1571, i_10_1572, i_10_1573, i_10_1574, i_10_1575, i_10_1576, i_10_1577, i_10_1578, i_10_1579, i_10_1580, i_10_1581, i_10_1582, i_10_1583, i_10_1584, i_10_1585, i_10_1586, i_10_1587, i_10_1588, i_10_1589, i_10_1590, i_10_1591, i_10_1592, i_10_1593, i_10_1594, i_10_1595, i_10_1596, i_10_1597, i_10_1598, i_10_1599, i_10_1600, i_10_1601, i_10_1602, i_10_1603, i_10_1604, i_10_1605, i_10_1606, i_10_1607, i_10_1608, i_10_1609, i_10_1610, i_10_1611, i_10_1612, i_10_1613, i_10_1614, i_10_1615, i_10_1616, i_10_1617, i_10_1618, i_10_1619, i_10_1620, i_10_1621, i_10_1622, i_10_1623, i_10_1624, i_10_1625, i_10_1626, i_10_1627, i_10_1628, i_10_1629, i_10_1630, i_10_1631, i_10_1632, i_10_1633, i_10_1634, i_10_1635, i_10_1636, i_10_1637, i_10_1638, i_10_1639, i_10_1640, i_10_1641, i_10_1642, i_10_1643, i_10_1644, i_10_1645, i_10_1646, i_10_1647, i_10_1648, i_10_1649, i_10_1650, i_10_1651, i_10_1652, i_10_1653, i_10_1654, i_10_1655, i_10_1656, i_10_1657, i_10_1658, i_10_1659, i_10_1660, i_10_1661, i_10_1662, i_10_1663, i_10_1664, i_10_1665, i_10_1666, i_10_1667, i_10_1668, i_10_1669, i_10_1670, i_10_1671, i_10_1672, i_10_1673, i_10_1674, i_10_1675, i_10_1676, i_10_1677, i_10_1678, i_10_1679, i_10_1680, i_10_1681, i_10_1682, i_10_1683, i_10_1684, i_10_1685, i_10_1686, i_10_1687, i_10_1688, i_10_1689, i_10_1690, i_10_1691, i_10_1692, i_10_1693, i_10_1694, i_10_1695, i_10_1696, i_10_1697, i_10_1698, i_10_1699, i_10_1700, i_10_1701, i_10_1702, i_10_1703, i_10_1704, i_10_1705, i_10_1706, i_10_1707, i_10_1708, i_10_1709, i_10_1710, i_10_1711, i_10_1712, i_10_1713, i_10_1714, i_10_1715, i_10_1716, i_10_1717, i_10_1718, i_10_1719, i_10_1720, i_10_1721, i_10_1722, i_10_1723, i_10_1724, i_10_1725, i_10_1726, i_10_1727, i_10_1728, i_10_1729, i_10_1730, i_10_1731, i_10_1732, i_10_1733, i_10_1734, i_10_1735, i_10_1736, i_10_1737, i_10_1738, i_10_1739, i_10_1740, i_10_1741, i_10_1742, i_10_1743, i_10_1744, i_10_1745, i_10_1746, i_10_1747, i_10_1748, i_10_1749, i_10_1750, i_10_1751, i_10_1752, i_10_1753, i_10_1754, i_10_1755, i_10_1756, i_10_1757, i_10_1758, i_10_1759, i_10_1760, i_10_1761, i_10_1762, i_10_1763, i_10_1764, i_10_1765, i_10_1766, i_10_1767, i_10_1768, i_10_1769, i_10_1770, i_10_1771, i_10_1772, i_10_1773, i_10_1774, i_10_1775, i_10_1776, i_10_1777, i_10_1778, i_10_1779, i_10_1780, i_10_1781, i_10_1782, i_10_1783, i_10_1784, i_10_1785, i_10_1786, i_10_1787, i_10_1788, i_10_1789, i_10_1790, i_10_1791, i_10_1792, i_10_1793, i_10_1794, i_10_1795, i_10_1796, i_10_1797, i_10_1798, i_10_1799, i_10_1800, i_10_1801, i_10_1802, i_10_1803, i_10_1804, i_10_1805, i_10_1806, i_10_1807, i_10_1808, i_10_1809, i_10_1810, i_10_1811, i_10_1812, i_10_1813, i_10_1814, i_10_1815, i_10_1816, i_10_1817, i_10_1818, i_10_1819, i_10_1820, i_10_1821, i_10_1822, i_10_1823, i_10_1824, i_10_1825, i_10_1826, i_10_1827, i_10_1828, i_10_1829, i_10_1830, i_10_1831, i_10_1832, i_10_1833, i_10_1834, i_10_1835, i_10_1836, i_10_1837, i_10_1838, i_10_1839, i_10_1840, i_10_1841, i_10_1842, i_10_1843, i_10_1844, i_10_1845, i_10_1846, i_10_1847, i_10_1848, i_10_1849, i_10_1850, i_10_1851, i_10_1852, i_10_1853, i_10_1854, i_10_1855, i_10_1856, i_10_1857, i_10_1858, i_10_1859, i_10_1860, i_10_1861, i_10_1862, i_10_1863, i_10_1864, i_10_1865, i_10_1866, i_10_1867, i_10_1868, i_10_1869, i_10_1870, i_10_1871, i_10_1872, i_10_1873, i_10_1874, i_10_1875, i_10_1876, i_10_1877, i_10_1878, i_10_1879, i_10_1880, i_10_1881, i_10_1882, i_10_1883, i_10_1884, i_10_1885, i_10_1886, i_10_1887, i_10_1888, i_10_1889, i_10_1890, i_10_1891, i_10_1892, i_10_1893, i_10_1894, i_10_1895, i_10_1896, i_10_1897, i_10_1898, i_10_1899, i_10_1900, i_10_1901, i_10_1902, i_10_1903, i_10_1904, i_10_1905, i_10_1906, i_10_1907, i_10_1908, i_10_1909, i_10_1910, i_10_1911, i_10_1912, i_10_1913, i_10_1914, i_10_1915, i_10_1916, i_10_1917, i_10_1918, i_10_1919, i_10_1920, i_10_1921, i_10_1922, i_10_1923, i_10_1924, i_10_1925, i_10_1926, i_10_1927, i_10_1928, i_10_1929, i_10_1930, i_10_1931, i_10_1932, i_10_1933, i_10_1934, i_10_1935, i_10_1936, i_10_1937, i_10_1938, i_10_1939, i_10_1940, i_10_1941, i_10_1942, i_10_1943, i_10_1944, i_10_1945, i_10_1946, i_10_1947, i_10_1948, i_10_1949, i_10_1950, i_10_1951, i_10_1952, i_10_1953, i_10_1954, i_10_1955, i_10_1956, i_10_1957, i_10_1958, i_10_1959, i_10_1960, i_10_1961, i_10_1962, i_10_1963, i_10_1964, i_10_1965, i_10_1966, i_10_1967, i_10_1968, i_10_1969, i_10_1970, i_10_1971, i_10_1972, i_10_1973, i_10_1974, i_10_1975, i_10_1976, i_10_1977, i_10_1978, i_10_1979, i_10_1980, i_10_1981, i_10_1982, i_10_1983, i_10_1984, i_10_1985, i_10_1986, i_10_1987, i_10_1988, i_10_1989, i_10_1990, i_10_1991, i_10_1992, i_10_1993, i_10_1994, i_10_1995, i_10_1996, i_10_1997, i_10_1998, i_10_1999, i_10_2000, i_10_2001, i_10_2002, i_10_2003, i_10_2004, i_10_2005, i_10_2006, i_10_2007, i_10_2008, i_10_2009, i_10_2010, i_10_2011, i_10_2012, i_10_2013, i_10_2014, i_10_2015, i_10_2016, i_10_2017, i_10_2018, i_10_2019, i_10_2020, i_10_2021, i_10_2022, i_10_2023, i_10_2024, i_10_2025, i_10_2026, i_10_2027, i_10_2028, i_10_2029, i_10_2030, i_10_2031, i_10_2032, i_10_2033, i_10_2034, i_10_2035, i_10_2036, i_10_2037, i_10_2038, i_10_2039, i_10_2040, i_10_2041, i_10_2042, i_10_2043, i_10_2044, i_10_2045, i_10_2046, i_10_2047, i_10_2048, i_10_2049, i_10_2050, i_10_2051, i_10_2052, i_10_2053, i_10_2054, i_10_2055, i_10_2056, i_10_2057, i_10_2058, i_10_2059, i_10_2060, i_10_2061, i_10_2062, i_10_2063, i_10_2064, i_10_2065, i_10_2066, i_10_2067, i_10_2068, i_10_2069, i_10_2070, i_10_2071, i_10_2072, i_10_2073, i_10_2074, i_10_2075, i_10_2076, i_10_2077, i_10_2078, i_10_2079, i_10_2080, i_10_2081, i_10_2082, i_10_2083, i_10_2084, i_10_2085, i_10_2086, i_10_2087, i_10_2088, i_10_2089, i_10_2090, i_10_2091, i_10_2092, i_10_2093, i_10_2094, i_10_2095, i_10_2096, i_10_2097, i_10_2098, i_10_2099, i_10_2100, i_10_2101, i_10_2102, i_10_2103, i_10_2104, i_10_2105, i_10_2106, i_10_2107, i_10_2108, i_10_2109, i_10_2110, i_10_2111, i_10_2112, i_10_2113, i_10_2114, i_10_2115, i_10_2116, i_10_2117, i_10_2118, i_10_2119, i_10_2120, i_10_2121, i_10_2122, i_10_2123, i_10_2124, i_10_2125, i_10_2126, i_10_2127, i_10_2128, i_10_2129, i_10_2130, i_10_2131, i_10_2132, i_10_2133, i_10_2134, i_10_2135, i_10_2136, i_10_2137, i_10_2138, i_10_2139, i_10_2140, i_10_2141, i_10_2142, i_10_2143, i_10_2144, i_10_2145, i_10_2146, i_10_2147, i_10_2148, i_10_2149, i_10_2150, i_10_2151, i_10_2152, i_10_2153, i_10_2154, i_10_2155, i_10_2156, i_10_2157, i_10_2158, i_10_2159, i_10_2160, i_10_2161, i_10_2162, i_10_2163, i_10_2164, i_10_2165, i_10_2166, i_10_2167, i_10_2168, i_10_2169, i_10_2170, i_10_2171, i_10_2172, i_10_2173, i_10_2174, i_10_2175, i_10_2176, i_10_2177, i_10_2178, i_10_2179, i_10_2180, i_10_2181, i_10_2182, i_10_2183, i_10_2184, i_10_2185, i_10_2186, i_10_2187, i_10_2188, i_10_2189, i_10_2190, i_10_2191, i_10_2192, i_10_2193, i_10_2194, i_10_2195, i_10_2196, i_10_2197, i_10_2198, i_10_2199, i_10_2200, i_10_2201, i_10_2202, i_10_2203, i_10_2204, i_10_2205, i_10_2206, i_10_2207, i_10_2208, i_10_2209, i_10_2210, i_10_2211, i_10_2212, i_10_2213, i_10_2214, i_10_2215, i_10_2216, i_10_2217, i_10_2218, i_10_2219, i_10_2220, i_10_2221, i_10_2222, i_10_2223, i_10_2224, i_10_2225, i_10_2226, i_10_2227, i_10_2228, i_10_2229, i_10_2230, i_10_2231, i_10_2232, i_10_2233, i_10_2234, i_10_2235, i_10_2236, i_10_2237, i_10_2238, i_10_2239, i_10_2240, i_10_2241, i_10_2242, i_10_2243, i_10_2244, i_10_2245, i_10_2246, i_10_2247, i_10_2248, i_10_2249, i_10_2250, i_10_2251, i_10_2252, i_10_2253, i_10_2254, i_10_2255, i_10_2256, i_10_2257, i_10_2258, i_10_2259, i_10_2260, i_10_2261, i_10_2262, i_10_2263, i_10_2264, i_10_2265, i_10_2266, i_10_2267, i_10_2268, i_10_2269, i_10_2270, i_10_2271, i_10_2272, i_10_2273, i_10_2274, i_10_2275, i_10_2276, i_10_2277, i_10_2278, i_10_2279, i_10_2280, i_10_2281, i_10_2282, i_10_2283, i_10_2284, i_10_2285, i_10_2286, i_10_2287, i_10_2288, i_10_2289, i_10_2290, i_10_2291, i_10_2292, i_10_2293, i_10_2294, i_10_2295, i_10_2296, i_10_2297, i_10_2298, i_10_2299, i_10_2300, i_10_2301, i_10_2302, i_10_2303, i_10_2304, i_10_2305, i_10_2306, i_10_2307, i_10_2308, i_10_2309, i_10_2310, i_10_2311, i_10_2312, i_10_2313, i_10_2314, i_10_2315, i_10_2316, i_10_2317, i_10_2318, i_10_2319, i_10_2320, i_10_2321, i_10_2322, i_10_2323, i_10_2324, i_10_2325, i_10_2326, i_10_2327, i_10_2328, i_10_2329, i_10_2330, i_10_2331, i_10_2332, i_10_2333, i_10_2334, i_10_2335, i_10_2336, i_10_2337, i_10_2338, i_10_2339, i_10_2340, i_10_2341, i_10_2342, i_10_2343, i_10_2344, i_10_2345, i_10_2346, i_10_2347, i_10_2348, i_10_2349, i_10_2350, i_10_2351, i_10_2352, i_10_2353, i_10_2354, i_10_2355, i_10_2356, i_10_2357, i_10_2358, i_10_2359, i_10_2360, i_10_2361, i_10_2362, i_10_2363, i_10_2364, i_10_2365, i_10_2366, i_10_2367, i_10_2368, i_10_2369, i_10_2370, i_10_2371, i_10_2372, i_10_2373, i_10_2374, i_10_2375, i_10_2376, i_10_2377, i_10_2378, i_10_2379, i_10_2380, i_10_2381, i_10_2382, i_10_2383, i_10_2384, i_10_2385, i_10_2386, i_10_2387, i_10_2388, i_10_2389, i_10_2390, i_10_2391, i_10_2392, i_10_2393, i_10_2394, i_10_2395, i_10_2396, i_10_2397, i_10_2398, i_10_2399, i_10_2400, i_10_2401, i_10_2402, i_10_2403, i_10_2404, i_10_2405, i_10_2406, i_10_2407, i_10_2408, i_10_2409, i_10_2410, i_10_2411, i_10_2412, i_10_2413, i_10_2414, i_10_2415, i_10_2416, i_10_2417, i_10_2418, i_10_2419, i_10_2420, i_10_2421, i_10_2422, i_10_2423, i_10_2424, i_10_2425, i_10_2426, i_10_2427, i_10_2428, i_10_2429, i_10_2430, i_10_2431, i_10_2432, i_10_2433, i_10_2434, i_10_2435, i_10_2436, i_10_2437, i_10_2438, i_10_2439, i_10_2440, i_10_2441, i_10_2442, i_10_2443, i_10_2444, i_10_2445, i_10_2446, i_10_2447, i_10_2448, i_10_2449, i_10_2450, i_10_2451, i_10_2452, i_10_2453, i_10_2454, i_10_2455, i_10_2456, i_10_2457, i_10_2458, i_10_2459, i_10_2460, i_10_2461, i_10_2462, i_10_2463, i_10_2464, i_10_2465, i_10_2466, i_10_2467, i_10_2468, i_10_2469, i_10_2470, i_10_2471, i_10_2472, i_10_2473, i_10_2474, i_10_2475, i_10_2476, i_10_2477, i_10_2478, i_10_2479, i_10_2480, i_10_2481, i_10_2482, i_10_2483, i_10_2484, i_10_2485, i_10_2486, i_10_2487, i_10_2488, i_10_2489, i_10_2490, i_10_2491, i_10_2492, i_10_2493, i_10_2494, i_10_2495, i_10_2496, i_10_2497, i_10_2498, i_10_2499, i_10_2500, i_10_2501, i_10_2502, i_10_2503, i_10_2504, i_10_2505, i_10_2506, i_10_2507, i_10_2508, i_10_2509, i_10_2510, i_10_2511, i_10_2512, i_10_2513, i_10_2514, i_10_2515, i_10_2516, i_10_2517, i_10_2518, i_10_2519, i_10_2520, i_10_2521, i_10_2522, i_10_2523, i_10_2524, i_10_2525, i_10_2526, i_10_2527, i_10_2528, i_10_2529, i_10_2530, i_10_2531, i_10_2532, i_10_2533, i_10_2534, i_10_2535, i_10_2536, i_10_2537, i_10_2538, i_10_2539, i_10_2540, i_10_2541, i_10_2542, i_10_2543, i_10_2544, i_10_2545, i_10_2546, i_10_2547, i_10_2548, i_10_2549, i_10_2550, i_10_2551, i_10_2552, i_10_2553, i_10_2554, i_10_2555, i_10_2556, i_10_2557, i_10_2558, i_10_2559, i_10_2560, i_10_2561, i_10_2562, i_10_2563, i_10_2564, i_10_2565, i_10_2566, i_10_2567, i_10_2568, i_10_2569, i_10_2570, i_10_2571, i_10_2572, i_10_2573, i_10_2574, i_10_2575, i_10_2576, i_10_2577, i_10_2578, i_10_2579, i_10_2580, i_10_2581, i_10_2582, i_10_2583, i_10_2584, i_10_2585, i_10_2586, i_10_2587, i_10_2588, i_10_2589, i_10_2590, i_10_2591, i_10_2592, i_10_2593, i_10_2594, i_10_2595, i_10_2596, i_10_2597, i_10_2598, i_10_2599, i_10_2600, i_10_2601, i_10_2602, i_10_2603, i_10_2604, i_10_2605, i_10_2606, i_10_2607, i_10_2608, i_10_2609, i_10_2610, i_10_2611, i_10_2612, i_10_2613, i_10_2614, i_10_2615, i_10_2616, i_10_2617, i_10_2618, i_10_2619, i_10_2620, i_10_2621, i_10_2622, i_10_2623, i_10_2624, i_10_2625, i_10_2626, i_10_2627, i_10_2628, i_10_2629, i_10_2630, i_10_2631, i_10_2632, i_10_2633, i_10_2634, i_10_2635, i_10_2636, i_10_2637, i_10_2638, i_10_2639, i_10_2640, i_10_2641, i_10_2642, i_10_2643, i_10_2644, i_10_2645, i_10_2646, i_10_2647, i_10_2648, i_10_2649, i_10_2650, i_10_2651, i_10_2652, i_10_2653, i_10_2654, i_10_2655, i_10_2656, i_10_2657, i_10_2658, i_10_2659, i_10_2660, i_10_2661, i_10_2662, i_10_2663, i_10_2664, i_10_2665, i_10_2666, i_10_2667, i_10_2668, i_10_2669, i_10_2670, i_10_2671, i_10_2672, i_10_2673, i_10_2674, i_10_2675, i_10_2676, i_10_2677, i_10_2678, i_10_2679, i_10_2680, i_10_2681, i_10_2682, i_10_2683, i_10_2684, i_10_2685, i_10_2686, i_10_2687, i_10_2688, i_10_2689, i_10_2690, i_10_2691, i_10_2692, i_10_2693, i_10_2694, i_10_2695, i_10_2696, i_10_2697, i_10_2698, i_10_2699, i_10_2700, i_10_2701, i_10_2702, i_10_2703, i_10_2704, i_10_2705, i_10_2706, i_10_2707, i_10_2708, i_10_2709, i_10_2710, i_10_2711, i_10_2712, i_10_2713, i_10_2714, i_10_2715, i_10_2716, i_10_2717, i_10_2718, i_10_2719, i_10_2720, i_10_2721, i_10_2722, i_10_2723, i_10_2724, i_10_2725, i_10_2726, i_10_2727, i_10_2728, i_10_2729, i_10_2730, i_10_2731, i_10_2732, i_10_2733, i_10_2734, i_10_2735, i_10_2736, i_10_2737, i_10_2738, i_10_2739, i_10_2740, i_10_2741, i_10_2742, i_10_2743, i_10_2744, i_10_2745, i_10_2746, i_10_2747, i_10_2748, i_10_2749, i_10_2750, i_10_2751, i_10_2752, i_10_2753, i_10_2754, i_10_2755, i_10_2756, i_10_2757, i_10_2758, i_10_2759, i_10_2760, i_10_2761, i_10_2762, i_10_2763, i_10_2764, i_10_2765, i_10_2766, i_10_2767, i_10_2768, i_10_2769, i_10_2770, i_10_2771, i_10_2772, i_10_2773, i_10_2774, i_10_2775, i_10_2776, i_10_2777, i_10_2778, i_10_2779, i_10_2780, i_10_2781, i_10_2782, i_10_2783, i_10_2784, i_10_2785, i_10_2786, i_10_2787, i_10_2788, i_10_2789, i_10_2790, i_10_2791, i_10_2792, i_10_2793, i_10_2794, i_10_2795, i_10_2796, i_10_2797, i_10_2798, i_10_2799, i_10_2800, i_10_2801, i_10_2802, i_10_2803, i_10_2804, i_10_2805, i_10_2806, i_10_2807, i_10_2808, i_10_2809, i_10_2810, i_10_2811, i_10_2812, i_10_2813, i_10_2814, i_10_2815, i_10_2816, i_10_2817, i_10_2818, i_10_2819, i_10_2820, i_10_2821, i_10_2822, i_10_2823, i_10_2824, i_10_2825, i_10_2826, i_10_2827, i_10_2828, i_10_2829, i_10_2830, i_10_2831, i_10_2832, i_10_2833, i_10_2834, i_10_2835, i_10_2836, i_10_2837, i_10_2838, i_10_2839, i_10_2840, i_10_2841, i_10_2842, i_10_2843, i_10_2844, i_10_2845, i_10_2846, i_10_2847, i_10_2848, i_10_2849, i_10_2850, i_10_2851, i_10_2852, i_10_2853, i_10_2854, i_10_2855, i_10_2856, i_10_2857, i_10_2858, i_10_2859, i_10_2860, i_10_2861, i_10_2862, i_10_2863, i_10_2864, i_10_2865, i_10_2866, i_10_2867, i_10_2868, i_10_2869, i_10_2870, i_10_2871, i_10_2872, i_10_2873, i_10_2874, i_10_2875, i_10_2876, i_10_2877, i_10_2878, i_10_2879, i_10_2880, i_10_2881, i_10_2882, i_10_2883, i_10_2884, i_10_2885, i_10_2886, i_10_2887, i_10_2888, i_10_2889, i_10_2890, i_10_2891, i_10_2892, i_10_2893, i_10_2894, i_10_2895, i_10_2896, i_10_2897, i_10_2898, i_10_2899, i_10_2900, i_10_2901, i_10_2902, i_10_2903, i_10_2904, i_10_2905, i_10_2906, i_10_2907, i_10_2908, i_10_2909, i_10_2910, i_10_2911, i_10_2912, i_10_2913, i_10_2914, i_10_2915, i_10_2916, i_10_2917, i_10_2918, i_10_2919, i_10_2920, i_10_2921, i_10_2922, i_10_2923, i_10_2924, i_10_2925, i_10_2926, i_10_2927, i_10_2928, i_10_2929, i_10_2930, i_10_2931, i_10_2932, i_10_2933, i_10_2934, i_10_2935, i_10_2936, i_10_2937, i_10_2938, i_10_2939, i_10_2940, i_10_2941, i_10_2942, i_10_2943, i_10_2944, i_10_2945, i_10_2946, i_10_2947, i_10_2948, i_10_2949, i_10_2950, i_10_2951, i_10_2952, i_10_2953, i_10_2954, i_10_2955, i_10_2956, i_10_2957, i_10_2958, i_10_2959, i_10_2960, i_10_2961, i_10_2962, i_10_2963, i_10_2964, i_10_2965, i_10_2966, i_10_2967, i_10_2968, i_10_2969, i_10_2970, i_10_2971, i_10_2972, i_10_2973, i_10_2974, i_10_2975, i_10_2976, i_10_2977, i_10_2978, i_10_2979, i_10_2980, i_10_2981, i_10_2982, i_10_2983, i_10_2984, i_10_2985, i_10_2986, i_10_2987, i_10_2988, i_10_2989, i_10_2990, i_10_2991, i_10_2992, i_10_2993, i_10_2994, i_10_2995, i_10_2996, i_10_2997, i_10_2998, i_10_2999, i_10_3000, i_10_3001, i_10_3002, i_10_3003, i_10_3004, i_10_3005, i_10_3006, i_10_3007, i_10_3008, i_10_3009, i_10_3010, i_10_3011, i_10_3012, i_10_3013, i_10_3014, i_10_3015, i_10_3016, i_10_3017, i_10_3018, i_10_3019, i_10_3020, i_10_3021, i_10_3022, i_10_3023, i_10_3024, i_10_3025, i_10_3026, i_10_3027, i_10_3028, i_10_3029, i_10_3030, i_10_3031, i_10_3032, i_10_3033, i_10_3034, i_10_3035, i_10_3036, i_10_3037, i_10_3038, i_10_3039, i_10_3040, i_10_3041, i_10_3042, i_10_3043, i_10_3044, i_10_3045, i_10_3046, i_10_3047, i_10_3048, i_10_3049, i_10_3050, i_10_3051, i_10_3052, i_10_3053, i_10_3054, i_10_3055, i_10_3056, i_10_3057, i_10_3058, i_10_3059, i_10_3060, i_10_3061, i_10_3062, i_10_3063, i_10_3064, i_10_3065, i_10_3066, i_10_3067, i_10_3068, i_10_3069, i_10_3070, i_10_3071, i_10_3072, i_10_3073, i_10_3074, i_10_3075, i_10_3076, i_10_3077, i_10_3078, i_10_3079, i_10_3080, i_10_3081, i_10_3082, i_10_3083, i_10_3084, i_10_3085, i_10_3086, i_10_3087, i_10_3088, i_10_3089, i_10_3090, i_10_3091, i_10_3092, i_10_3093, i_10_3094, i_10_3095, i_10_3096, i_10_3097, i_10_3098, i_10_3099, i_10_3100, i_10_3101, i_10_3102, i_10_3103, i_10_3104, i_10_3105, i_10_3106, i_10_3107, i_10_3108, i_10_3109, i_10_3110, i_10_3111, i_10_3112, i_10_3113, i_10_3114, i_10_3115, i_10_3116, i_10_3117, i_10_3118, i_10_3119, i_10_3120, i_10_3121, i_10_3122, i_10_3123, i_10_3124, i_10_3125, i_10_3126, i_10_3127, i_10_3128, i_10_3129, i_10_3130, i_10_3131, i_10_3132, i_10_3133, i_10_3134, i_10_3135, i_10_3136, i_10_3137, i_10_3138, i_10_3139, i_10_3140, i_10_3141, i_10_3142, i_10_3143, i_10_3144, i_10_3145, i_10_3146, i_10_3147, i_10_3148, i_10_3149, i_10_3150, i_10_3151, i_10_3152, i_10_3153, i_10_3154, i_10_3155, i_10_3156, i_10_3157, i_10_3158, i_10_3159, i_10_3160, i_10_3161, i_10_3162, i_10_3163, i_10_3164, i_10_3165, i_10_3166, i_10_3167, i_10_3168, i_10_3169, i_10_3170, i_10_3171, i_10_3172, i_10_3173, i_10_3174, i_10_3175, i_10_3176, i_10_3177, i_10_3178, i_10_3179, i_10_3180, i_10_3181, i_10_3182, i_10_3183, i_10_3184, i_10_3185, i_10_3186, i_10_3187, i_10_3188, i_10_3189, i_10_3190, i_10_3191, i_10_3192, i_10_3193, i_10_3194, i_10_3195, i_10_3196, i_10_3197, i_10_3198, i_10_3199, i_10_3200, i_10_3201, i_10_3202, i_10_3203, i_10_3204, i_10_3205, i_10_3206, i_10_3207, i_10_3208, i_10_3209, i_10_3210, i_10_3211, i_10_3212, i_10_3213, i_10_3214, i_10_3215, i_10_3216, i_10_3217, i_10_3218, i_10_3219, i_10_3220, i_10_3221, i_10_3222, i_10_3223, i_10_3224, i_10_3225, i_10_3226, i_10_3227, i_10_3228, i_10_3229, i_10_3230, i_10_3231, i_10_3232, i_10_3233, i_10_3234, i_10_3235, i_10_3236, i_10_3237, i_10_3238, i_10_3239, i_10_3240, i_10_3241, i_10_3242, i_10_3243, i_10_3244, i_10_3245, i_10_3246, i_10_3247, i_10_3248, i_10_3249, i_10_3250, i_10_3251, i_10_3252, i_10_3253, i_10_3254, i_10_3255, i_10_3256, i_10_3257, i_10_3258, i_10_3259, i_10_3260, i_10_3261, i_10_3262, i_10_3263, i_10_3264, i_10_3265, i_10_3266, i_10_3267, i_10_3268, i_10_3269, i_10_3270, i_10_3271, i_10_3272, i_10_3273, i_10_3274, i_10_3275, i_10_3276, i_10_3277, i_10_3278, i_10_3279, i_10_3280, i_10_3281, i_10_3282, i_10_3283, i_10_3284, i_10_3285, i_10_3286, i_10_3287, i_10_3288, i_10_3289, i_10_3290, i_10_3291, i_10_3292, i_10_3293, i_10_3294, i_10_3295, i_10_3296, i_10_3297, i_10_3298, i_10_3299, i_10_3300, i_10_3301, i_10_3302, i_10_3303, i_10_3304, i_10_3305, i_10_3306, i_10_3307, i_10_3308, i_10_3309, i_10_3310, i_10_3311, i_10_3312, i_10_3313, i_10_3314, i_10_3315, i_10_3316, i_10_3317, i_10_3318, i_10_3319, i_10_3320, i_10_3321, i_10_3322, i_10_3323, i_10_3324, i_10_3325, i_10_3326, i_10_3327, i_10_3328, i_10_3329, i_10_3330, i_10_3331, i_10_3332, i_10_3333, i_10_3334, i_10_3335, i_10_3336, i_10_3337, i_10_3338, i_10_3339, i_10_3340, i_10_3341, i_10_3342, i_10_3343, i_10_3344, i_10_3345, i_10_3346, i_10_3347, i_10_3348, i_10_3349, i_10_3350, i_10_3351, i_10_3352, i_10_3353, i_10_3354, i_10_3355, i_10_3356, i_10_3357, i_10_3358, i_10_3359, i_10_3360, i_10_3361, i_10_3362, i_10_3363, i_10_3364, i_10_3365, i_10_3366, i_10_3367, i_10_3368, i_10_3369, i_10_3370, i_10_3371, i_10_3372, i_10_3373, i_10_3374, i_10_3375, i_10_3376, i_10_3377, i_10_3378, i_10_3379, i_10_3380, i_10_3381, i_10_3382, i_10_3383, i_10_3384, i_10_3385, i_10_3386, i_10_3387, i_10_3388, i_10_3389, i_10_3390, i_10_3391, i_10_3392, i_10_3393, i_10_3394, i_10_3395, i_10_3396, i_10_3397, i_10_3398, i_10_3399, i_10_3400, i_10_3401, i_10_3402, i_10_3403, i_10_3404, i_10_3405, i_10_3406, i_10_3407, i_10_3408, i_10_3409, i_10_3410, i_10_3411, i_10_3412, i_10_3413, i_10_3414, i_10_3415, i_10_3416, i_10_3417, i_10_3418, i_10_3419, i_10_3420, i_10_3421, i_10_3422, i_10_3423, i_10_3424, i_10_3425, i_10_3426, i_10_3427, i_10_3428, i_10_3429, i_10_3430, i_10_3431, i_10_3432, i_10_3433, i_10_3434, i_10_3435, i_10_3436, i_10_3437, i_10_3438, i_10_3439, i_10_3440, i_10_3441, i_10_3442, i_10_3443, i_10_3444, i_10_3445, i_10_3446, i_10_3447, i_10_3448, i_10_3449, i_10_3450, i_10_3451, i_10_3452, i_10_3453, i_10_3454, i_10_3455, i_10_3456, i_10_3457, i_10_3458, i_10_3459, i_10_3460, i_10_3461, i_10_3462, i_10_3463, i_10_3464, i_10_3465, i_10_3466, i_10_3467, i_10_3468, i_10_3469, i_10_3470, i_10_3471, i_10_3472, i_10_3473, i_10_3474, i_10_3475, i_10_3476, i_10_3477, i_10_3478, i_10_3479, i_10_3480, i_10_3481, i_10_3482, i_10_3483, i_10_3484, i_10_3485, i_10_3486, i_10_3487, i_10_3488, i_10_3489, i_10_3490, i_10_3491, i_10_3492, i_10_3493, i_10_3494, i_10_3495, i_10_3496, i_10_3497, i_10_3498, i_10_3499, i_10_3500, i_10_3501, i_10_3502, i_10_3503, i_10_3504, i_10_3505, i_10_3506, i_10_3507, i_10_3508, i_10_3509, i_10_3510, i_10_3511, i_10_3512, i_10_3513, i_10_3514, i_10_3515, i_10_3516, i_10_3517, i_10_3518, i_10_3519, i_10_3520, i_10_3521, i_10_3522, i_10_3523, i_10_3524, i_10_3525, i_10_3526, i_10_3527, i_10_3528, i_10_3529, i_10_3530, i_10_3531, i_10_3532, i_10_3533, i_10_3534, i_10_3535, i_10_3536, i_10_3537, i_10_3538, i_10_3539, i_10_3540, i_10_3541, i_10_3542, i_10_3543, i_10_3544, i_10_3545, i_10_3546, i_10_3547, i_10_3548, i_10_3549, i_10_3550, i_10_3551, i_10_3552, i_10_3553, i_10_3554, i_10_3555, i_10_3556, i_10_3557, i_10_3558, i_10_3559, i_10_3560, i_10_3561, i_10_3562, i_10_3563, i_10_3564, i_10_3565, i_10_3566, i_10_3567, i_10_3568, i_10_3569, i_10_3570, i_10_3571, i_10_3572, i_10_3573, i_10_3574, i_10_3575, i_10_3576, i_10_3577, i_10_3578, i_10_3579, i_10_3580, i_10_3581, i_10_3582, i_10_3583, i_10_3584, i_10_3585, i_10_3586, i_10_3587, i_10_3588, i_10_3589, i_10_3590, i_10_3591, i_10_3592, i_10_3593, i_10_3594, i_10_3595, i_10_3596, i_10_3597, i_10_3598, i_10_3599, i_10_3600, i_10_3601, i_10_3602, i_10_3603, i_10_3604, i_10_3605, i_10_3606, i_10_3607, i_10_3608, i_10_3609, i_10_3610, i_10_3611, i_10_3612, i_10_3613, i_10_3614, i_10_3615, i_10_3616, i_10_3617, i_10_3618, i_10_3619, i_10_3620, i_10_3621, i_10_3622, i_10_3623, i_10_3624, i_10_3625, i_10_3626, i_10_3627, i_10_3628, i_10_3629, i_10_3630, i_10_3631, i_10_3632, i_10_3633, i_10_3634, i_10_3635, i_10_3636, i_10_3637, i_10_3638, i_10_3639, i_10_3640, i_10_3641, i_10_3642, i_10_3643, i_10_3644, i_10_3645, i_10_3646, i_10_3647, i_10_3648, i_10_3649, i_10_3650, i_10_3651, i_10_3652, i_10_3653, i_10_3654, i_10_3655, i_10_3656, i_10_3657, i_10_3658, i_10_3659, i_10_3660, i_10_3661, i_10_3662, i_10_3663, i_10_3664, i_10_3665, i_10_3666, i_10_3667, i_10_3668, i_10_3669, i_10_3670, i_10_3671, i_10_3672, i_10_3673, i_10_3674, i_10_3675, i_10_3676, i_10_3677, i_10_3678, i_10_3679, i_10_3680, i_10_3681, i_10_3682, i_10_3683, i_10_3684, i_10_3685, i_10_3686, i_10_3687, i_10_3688, i_10_3689, i_10_3690, i_10_3691, i_10_3692, i_10_3693, i_10_3694, i_10_3695, i_10_3696, i_10_3697, i_10_3698, i_10_3699, i_10_3700, i_10_3701, i_10_3702, i_10_3703, i_10_3704, i_10_3705, i_10_3706, i_10_3707, i_10_3708, i_10_3709, i_10_3710, i_10_3711, i_10_3712, i_10_3713, i_10_3714, i_10_3715, i_10_3716, i_10_3717, i_10_3718, i_10_3719, i_10_3720, i_10_3721, i_10_3722, i_10_3723, i_10_3724, i_10_3725, i_10_3726, i_10_3727, i_10_3728, i_10_3729, i_10_3730, i_10_3731, i_10_3732, i_10_3733, i_10_3734, i_10_3735, i_10_3736, i_10_3737, i_10_3738, i_10_3739, i_10_3740, i_10_3741, i_10_3742, i_10_3743, i_10_3744, i_10_3745, i_10_3746, i_10_3747, i_10_3748, i_10_3749, i_10_3750, i_10_3751, i_10_3752, i_10_3753, i_10_3754, i_10_3755, i_10_3756, i_10_3757, i_10_3758, i_10_3759, i_10_3760, i_10_3761, i_10_3762, i_10_3763, i_10_3764, i_10_3765, i_10_3766, i_10_3767, i_10_3768, i_10_3769, i_10_3770, i_10_3771, i_10_3772, i_10_3773, i_10_3774, i_10_3775, i_10_3776, i_10_3777, i_10_3778, i_10_3779, i_10_3780, i_10_3781, i_10_3782, i_10_3783, i_10_3784, i_10_3785, i_10_3786, i_10_3787, i_10_3788, i_10_3789, i_10_3790, i_10_3791, i_10_3792, i_10_3793, i_10_3794, i_10_3795, i_10_3796, i_10_3797, i_10_3798, i_10_3799, i_10_3800, i_10_3801, i_10_3802, i_10_3803, i_10_3804, i_10_3805, i_10_3806, i_10_3807, i_10_3808, i_10_3809, i_10_3810, i_10_3811, i_10_3812, i_10_3813, i_10_3814, i_10_3815, i_10_3816, i_10_3817, i_10_3818, i_10_3819, i_10_3820, i_10_3821, i_10_3822, i_10_3823, i_10_3824, i_10_3825, i_10_3826, i_10_3827, i_10_3828, i_10_3829, i_10_3830, i_10_3831, i_10_3832, i_10_3833, i_10_3834, i_10_3835, i_10_3836, i_10_3837, i_10_3838, i_10_3839, i_10_3840, i_10_3841, i_10_3842, i_10_3843, i_10_3844, i_10_3845, i_10_3846, i_10_3847, i_10_3848, i_10_3849, i_10_3850, i_10_3851, i_10_3852, i_10_3853, i_10_3854, i_10_3855, i_10_3856, i_10_3857, i_10_3858, i_10_3859, i_10_3860, i_10_3861, i_10_3862, i_10_3863, i_10_3864, i_10_3865, i_10_3866, i_10_3867, i_10_3868, i_10_3869, i_10_3870, i_10_3871, i_10_3872, i_10_3873, i_10_3874, i_10_3875, i_10_3876, i_10_3877, i_10_3878, i_10_3879, i_10_3880, i_10_3881, i_10_3882, i_10_3883, i_10_3884, i_10_3885, i_10_3886, i_10_3887, i_10_3888, i_10_3889, i_10_3890, i_10_3891, i_10_3892, i_10_3893, i_10_3894, i_10_3895, i_10_3896, i_10_3897, i_10_3898, i_10_3899, i_10_3900, i_10_3901, i_10_3902, i_10_3903, i_10_3904, i_10_3905, i_10_3906, i_10_3907, i_10_3908, i_10_3909, i_10_3910, i_10_3911, i_10_3912, i_10_3913, i_10_3914, i_10_3915, i_10_3916, i_10_3917, i_10_3918, i_10_3919, i_10_3920, i_10_3921, i_10_3922, i_10_3923, i_10_3924, i_10_3925, i_10_3926, i_10_3927, i_10_3928, i_10_3929, i_10_3930, i_10_3931, i_10_3932, i_10_3933, i_10_3934, i_10_3935, i_10_3936, i_10_3937, i_10_3938, i_10_3939, i_10_3940, i_10_3941, i_10_3942, i_10_3943, i_10_3944, i_10_3945, i_10_3946, i_10_3947, i_10_3948, i_10_3949, i_10_3950, i_10_3951, i_10_3952, i_10_3953, i_10_3954, i_10_3955, i_10_3956, i_10_3957, i_10_3958, i_10_3959, i_10_3960, i_10_3961, i_10_3962, i_10_3963, i_10_3964, i_10_3965, i_10_3966, i_10_3967, i_10_3968, i_10_3969, i_10_3970, i_10_3971, i_10_3972, i_10_3973, i_10_3974, i_10_3975, i_10_3976, i_10_3977, i_10_3978, i_10_3979, i_10_3980, i_10_3981, i_10_3982, i_10_3983, i_10_3984, i_10_3985, i_10_3986, i_10_3987, i_10_3988, i_10_3989, i_10_3990, i_10_3991, i_10_3992, i_10_3993, i_10_3994, i_10_3995, i_10_3996, i_10_3997, i_10_3998, i_10_3999, i_10_4000, i_10_4001, i_10_4002, i_10_4003, i_10_4004, i_10_4005, i_10_4006, i_10_4007, i_10_4008, i_10_4009, i_10_4010, i_10_4011, i_10_4012, i_10_4013, i_10_4014, i_10_4015, i_10_4016, i_10_4017, i_10_4018, i_10_4019, i_10_4020, i_10_4021, i_10_4022, i_10_4023, i_10_4024, i_10_4025, i_10_4026, i_10_4027, i_10_4028, i_10_4029, i_10_4030, i_10_4031, i_10_4032, i_10_4033, i_10_4034, i_10_4035, i_10_4036, i_10_4037, i_10_4038, i_10_4039, i_10_4040, i_10_4041, i_10_4042, i_10_4043, i_10_4044, i_10_4045, i_10_4046, i_10_4047, i_10_4048, i_10_4049, i_10_4050, i_10_4051, i_10_4052, i_10_4053, i_10_4054, i_10_4055, i_10_4056, i_10_4057, i_10_4058, i_10_4059, i_10_4060, i_10_4061, i_10_4062, i_10_4063, i_10_4064, i_10_4065, i_10_4066, i_10_4067, i_10_4068, i_10_4069, i_10_4070, i_10_4071, i_10_4072, i_10_4073, i_10_4074, i_10_4075, i_10_4076, i_10_4077, i_10_4078, i_10_4079, i_10_4080, i_10_4081, i_10_4082, i_10_4083, i_10_4084, i_10_4085, i_10_4086, i_10_4087, i_10_4088, i_10_4089, i_10_4090, i_10_4091, i_10_4092, i_10_4093, i_10_4094, i_10_4095, i_10_4096, i_10_4097, i_10_4098, i_10_4099, i_10_4100, i_10_4101, i_10_4102, i_10_4103, i_10_4104, i_10_4105, i_10_4106, i_10_4107, i_10_4108, i_10_4109, i_10_4110, i_10_4111, i_10_4112, i_10_4113, i_10_4114, i_10_4115, i_10_4116, i_10_4117, i_10_4118, i_10_4119, i_10_4120, i_10_4121, i_10_4122, i_10_4123, i_10_4124, i_10_4125, i_10_4126, i_10_4127, i_10_4128, i_10_4129, i_10_4130, i_10_4131, i_10_4132, i_10_4133, i_10_4134, i_10_4135, i_10_4136, i_10_4137, i_10_4138, i_10_4139, i_10_4140, i_10_4141, i_10_4142, i_10_4143, i_10_4144, i_10_4145, i_10_4146, i_10_4147, i_10_4148, i_10_4149, i_10_4150, i_10_4151, i_10_4152, i_10_4153, i_10_4154, i_10_4155, i_10_4156, i_10_4157, i_10_4158, i_10_4159, i_10_4160, i_10_4161, i_10_4162, i_10_4163, i_10_4164, i_10_4165, i_10_4166, i_10_4167, i_10_4168, i_10_4169, i_10_4170, i_10_4171, i_10_4172, i_10_4173, i_10_4174, i_10_4175, i_10_4176, i_10_4177, i_10_4178, i_10_4179, i_10_4180, i_10_4181, i_10_4182, i_10_4183, i_10_4184, i_10_4185, i_10_4186, i_10_4187, i_10_4188, i_10_4189, i_10_4190, i_10_4191, i_10_4192, i_10_4193, i_10_4194, i_10_4195, i_10_4196, i_10_4197, i_10_4198, i_10_4199, i_10_4200, i_10_4201, i_10_4202, i_10_4203, i_10_4204, i_10_4205, i_10_4206, i_10_4207, i_10_4208, i_10_4209, i_10_4210, i_10_4211, i_10_4212, i_10_4213, i_10_4214, i_10_4215, i_10_4216, i_10_4217, i_10_4218, i_10_4219, i_10_4220, i_10_4221, i_10_4222, i_10_4223, i_10_4224, i_10_4225, i_10_4226, i_10_4227, i_10_4228, i_10_4229, i_10_4230, i_10_4231, i_10_4232, i_10_4233, i_10_4234, i_10_4235, i_10_4236, i_10_4237, i_10_4238, i_10_4239, i_10_4240, i_10_4241, i_10_4242, i_10_4243, i_10_4244, i_10_4245, i_10_4246, i_10_4247, i_10_4248, i_10_4249, i_10_4250, i_10_4251, i_10_4252, i_10_4253, i_10_4254, i_10_4255, i_10_4256, i_10_4257, i_10_4258, i_10_4259, i_10_4260, i_10_4261, i_10_4262, i_10_4263, i_10_4264, i_10_4265, i_10_4266, i_10_4267, i_10_4268, i_10_4269, i_10_4270, i_10_4271, i_10_4272, i_10_4273, i_10_4274, i_10_4275, i_10_4276, i_10_4277, i_10_4278, i_10_4279, i_10_4280, i_10_4281, i_10_4282, i_10_4283, i_10_4284, i_10_4285, i_10_4286, i_10_4287, i_10_4288, i_10_4289, i_10_4290, i_10_4291, i_10_4292, i_10_4293, i_10_4294, i_10_4295, i_10_4296, i_10_4297, i_10_4298, i_10_4299, i_10_4300, i_10_4301, i_10_4302, i_10_4303, i_10_4304, i_10_4305, i_10_4306, i_10_4307, i_10_4308, i_10_4309, i_10_4310, i_10_4311, i_10_4312, i_10_4313, i_10_4314, i_10_4315, i_10_4316, i_10_4317, i_10_4318, i_10_4319, i_10_4320, i_10_4321, i_10_4322, i_10_4323, i_10_4324, i_10_4325, i_10_4326, i_10_4327, i_10_4328, i_10_4329, i_10_4330, i_10_4331, i_10_4332, i_10_4333, i_10_4334, i_10_4335, i_10_4336, i_10_4337, i_10_4338, i_10_4339, i_10_4340, i_10_4341, i_10_4342, i_10_4343, i_10_4344, i_10_4345, i_10_4346, i_10_4347, i_10_4348, i_10_4349, i_10_4350, i_10_4351, i_10_4352, i_10_4353, i_10_4354, i_10_4355, i_10_4356, i_10_4357, i_10_4358, i_10_4359, i_10_4360, i_10_4361, i_10_4362, i_10_4363, i_10_4364, i_10_4365, i_10_4366, i_10_4367, i_10_4368, i_10_4369, i_10_4370, i_10_4371, i_10_4372, i_10_4373, i_10_4374, i_10_4375, i_10_4376, i_10_4377, i_10_4378, i_10_4379, i_10_4380, i_10_4381, i_10_4382, i_10_4383, i_10_4384, i_10_4385, i_10_4386, i_10_4387, i_10_4388, i_10_4389, i_10_4390, i_10_4391, i_10_4392, i_10_4393, i_10_4394, i_10_4395, i_10_4396, i_10_4397, i_10_4398, i_10_4399, i_10_4400, i_10_4401, i_10_4402, i_10_4403, i_10_4404, i_10_4405, i_10_4406, i_10_4407, i_10_4408, i_10_4409, i_10_4410, i_10_4411, i_10_4412, i_10_4413, i_10_4414, i_10_4415, i_10_4416, i_10_4417, i_10_4418, i_10_4419, i_10_4420, i_10_4421, i_10_4422, i_10_4423, i_10_4424, i_10_4425, i_10_4426, i_10_4427, i_10_4428, i_10_4429, i_10_4430, i_10_4431, i_10_4432, i_10_4433, i_10_4434, i_10_4435, i_10_4436, i_10_4437, i_10_4438, i_10_4439, i_10_4440, i_10_4441, i_10_4442, i_10_4443, i_10_4444, i_10_4445, i_10_4446, i_10_4447, i_10_4448, i_10_4449, i_10_4450, i_10_4451, i_10_4452, i_10_4453, i_10_4454, i_10_4455, i_10_4456, i_10_4457, i_10_4458, i_10_4459, i_10_4460, i_10_4461, i_10_4462, i_10_4463, i_10_4464, i_10_4465, i_10_4466, i_10_4467, i_10_4468, i_10_4469, i_10_4470, i_10_4471, i_10_4472, i_10_4473, i_10_4474, i_10_4475, i_10_4476, i_10_4477, i_10_4478, i_10_4479, i_10_4480, i_10_4481, i_10_4482, i_10_4483, i_10_4484, i_10_4485, i_10_4486, i_10_4487, i_10_4488, i_10_4489, i_10_4490, i_10_4491, i_10_4492, i_10_4493, i_10_4494, i_10_4495, i_10_4496, i_10_4497, i_10_4498, i_10_4499, i_10_4500, i_10_4501, i_10_4502, i_10_4503, i_10_4504, i_10_4505, i_10_4506, i_10_4507, i_10_4508, i_10_4509, i_10_4510, i_10_4511, i_10_4512, i_10_4513, i_10_4514, i_10_4515, i_10_4516, i_10_4517, i_10_4518, i_10_4519, i_10_4520, i_10_4521, i_10_4522, i_10_4523, i_10_4524, i_10_4525, i_10_4526, i_10_4527, i_10_4528, i_10_4529, i_10_4530, i_10_4531, i_10_4532, i_10_4533, i_10_4534, i_10_4535, i_10_4536, i_10_4537, i_10_4538, i_10_4539, i_10_4540, i_10_4541, i_10_4542, i_10_4543, i_10_4544, i_10_4545, i_10_4546, i_10_4547, i_10_4548, i_10_4549, i_10_4550, i_10_4551, i_10_4552, i_10_4553, i_10_4554, i_10_4555, i_10_4556, i_10_4557, i_10_4558, i_10_4559, i_10_4560, i_10_4561, i_10_4562, i_10_4563, i_10_4564, i_10_4565, i_10_4566, i_10_4567, i_10_4568, i_10_4569, i_10_4570, i_10_4571, i_10_4572, i_10_4573, i_10_4574, i_10_4575, i_10_4576, i_10_4577, i_10_4578, i_10_4579, i_10_4580, i_10_4581, i_10_4582, i_10_4583, i_10_4584, i_10_4585, i_10_4586, i_10_4587, i_10_4588, i_10_4589, i_10_4590, i_10_4591, i_10_4592, i_10_4593, i_10_4594, i_10_4595, i_10_4596, i_10_4597, i_10_4598, i_10_4599, i_10_4600, i_10_4601, i_10_4602, i_10_4603, i_10_4604, i_10_4605, i_10_4606, i_10_4607;
  reg dly1, dly2;
  wire o_10_0, o_10_1, o_10_2, o_10_3, o_10_4, o_10_5, o_10_6, o_10_7, o_10_8, o_10_9, o_10_10, o_10_11, o_10_12, o_10_13, o_10_14, o_10_15, o_10_16, o_10_17, o_10_18, o_10_19, o_10_20, o_10_21, o_10_22, o_10_23, o_10_24, o_10_25, o_10_26, o_10_27, o_10_28, o_10_29, o_10_30, o_10_31, o_10_32, o_10_33, o_10_34, o_10_35, o_10_36, o_10_37, o_10_38, o_10_39, o_10_40, o_10_41, o_10_42, o_10_43, o_10_44, o_10_45, o_10_46, o_10_47, o_10_48, o_10_49, o_10_50, o_10_51, o_10_52, o_10_53, o_10_54, o_10_55, o_10_56, o_10_57, o_10_58, o_10_59, o_10_60, o_10_61, o_10_62, o_10_63, o_10_64, o_10_65, o_10_66, o_10_67, o_10_68, o_10_69, o_10_70, o_10_71, o_10_72, o_10_73, o_10_74, o_10_75, o_10_76, o_10_77, o_10_78, o_10_79, o_10_80, o_10_81, o_10_82, o_10_83, o_10_84, o_10_85, o_10_86, o_10_87, o_10_88, o_10_89, o_10_90, o_10_91, o_10_92, o_10_93, o_10_94, o_10_95, o_10_96, o_10_97, o_10_98, o_10_99, o_10_100, o_10_101, o_10_102, o_10_103, o_10_104, o_10_105, o_10_106, o_10_107, o_10_108, o_10_109, o_10_110, o_10_111, o_10_112, o_10_113, o_10_114, o_10_115, o_10_116, o_10_117, o_10_118, o_10_119, o_10_120, o_10_121, o_10_122, o_10_123, o_10_124, o_10_125, o_10_126, o_10_127, o_10_128, o_10_129, o_10_130, o_10_131, o_10_132, o_10_133, o_10_134, o_10_135, o_10_136, o_10_137, o_10_138, o_10_139, o_10_140, o_10_141, o_10_142, o_10_143, o_10_144, o_10_145, o_10_146, o_10_147, o_10_148, o_10_149, o_10_150, o_10_151, o_10_152, o_10_153, o_10_154, o_10_155, o_10_156, o_10_157, o_10_158, o_10_159, o_10_160, o_10_161, o_10_162, o_10_163, o_10_164, o_10_165, o_10_166, o_10_167, o_10_168, o_10_169, o_10_170, o_10_171, o_10_172, o_10_173, o_10_174, o_10_175, o_10_176, o_10_177, o_10_178, o_10_179, o_10_180, o_10_181, o_10_182, o_10_183, o_10_184, o_10_185, o_10_186, o_10_187, o_10_188, o_10_189, o_10_190, o_10_191, o_10_192, o_10_193, o_10_194, o_10_195, o_10_196, o_10_197, o_10_198, o_10_199, o_10_200, o_10_201, o_10_202, o_10_203, o_10_204, o_10_205, o_10_206, o_10_207, o_10_208, o_10_209, o_10_210, o_10_211, o_10_212, o_10_213, o_10_214, o_10_215, o_10_216, o_10_217, o_10_218, o_10_219, o_10_220, o_10_221, o_10_222, o_10_223, o_10_224, o_10_225, o_10_226, o_10_227, o_10_228, o_10_229, o_10_230, o_10_231, o_10_232, o_10_233, o_10_234, o_10_235, o_10_236, o_10_237, o_10_238, o_10_239, o_10_240, o_10_241, o_10_242, o_10_243, o_10_244, o_10_245, o_10_246, o_10_247, o_10_248, o_10_249, o_10_250, o_10_251, o_10_252, o_10_253, o_10_254, o_10_255, o_10_256, o_10_257, o_10_258, o_10_259, o_10_260, o_10_261, o_10_262, o_10_263, o_10_264, o_10_265, o_10_266, o_10_267, o_10_268, o_10_269, o_10_270, o_10_271, o_10_272, o_10_273, o_10_274, o_10_275, o_10_276, o_10_277, o_10_278, o_10_279, o_10_280, o_10_281, o_10_282, o_10_283, o_10_284, o_10_285, o_10_286, o_10_287, o_10_288, o_10_289, o_10_290, o_10_291, o_10_292, o_10_293, o_10_294, o_10_295, o_10_296, o_10_297, o_10_298, o_10_299, o_10_300, o_10_301, o_10_302, o_10_303, o_10_304, o_10_305, o_10_306, o_10_307, o_10_308, o_10_309, o_10_310, o_10_311, o_10_312, o_10_313, o_10_314, o_10_315, o_10_316, o_10_317, o_10_318, o_10_319, o_10_320, o_10_321, o_10_322, o_10_323, o_10_324, o_10_325, o_10_326, o_10_327, o_10_328, o_10_329, o_10_330, o_10_331, o_10_332, o_10_333, o_10_334, o_10_335, o_10_336, o_10_337, o_10_338, o_10_339, o_10_340, o_10_341, o_10_342, o_10_343, o_10_344, o_10_345, o_10_346, o_10_347, o_10_348, o_10_349, o_10_350, o_10_351, o_10_352, o_10_353, o_10_354, o_10_355, o_10_356, o_10_357, o_10_358, o_10_359, o_10_360, o_10_361, o_10_362, o_10_363, o_10_364, o_10_365, o_10_366, o_10_367, o_10_368, o_10_369, o_10_370, o_10_371, o_10_372, o_10_373, o_10_374, o_10_375, o_10_376, o_10_377, o_10_378, o_10_379, o_10_380, o_10_381, o_10_382, o_10_383, o_10_384, o_10_385, o_10_386, o_10_387, o_10_388, o_10_389, o_10_390, o_10_391, o_10_392, o_10_393, o_10_394, o_10_395, o_10_396, o_10_397, o_10_398, o_10_399, o_10_400, o_10_401, o_10_402, o_10_403, o_10_404, o_10_405, o_10_406, o_10_407, o_10_408, o_10_409, o_10_410, o_10_411, o_10_412, o_10_413, o_10_414, o_10_415, o_10_416, o_10_417, o_10_418, o_10_419, o_10_420, o_10_421, o_10_422, o_10_423, o_10_424, o_10_425, o_10_426, o_10_427, o_10_428, o_10_429, o_10_430, o_10_431, o_10_432, o_10_433, o_10_434, o_10_435, o_10_436, o_10_437, o_10_438, o_10_439, o_10_440, o_10_441, o_10_442, o_10_443, o_10_444, o_10_445, o_10_446, o_10_447, o_10_448, o_10_449, o_10_450, o_10_451, o_10_452, o_10_453, o_10_454, o_10_455, o_10_456, o_10_457, o_10_458, o_10_459, o_10_460, o_10_461, o_10_462, o_10_463, o_10_464, o_10_465, o_10_466, o_10_467, o_10_468, o_10_469, o_10_470, o_10_471, o_10_472, o_10_473, o_10_474, o_10_475, o_10_476, o_10_477, o_10_478, o_10_479, o_10_480, o_10_481, o_10_482, o_10_483, o_10_484, o_10_485, o_10_486, o_10_487, o_10_488, o_10_489, o_10_490, o_10_491, o_10_492, o_10_493, o_10_494, o_10_495, o_10_496, o_10_497, o_10_498, o_10_499, o_10_500, o_10_501, o_10_502, o_10_503, o_10_504, o_10_505, o_10_506, o_10_507, o_10_508, o_10_509, o_10_510, o_10_511;

  kernel_10 kernel_nulla( i_10_0, i_10_1, i_10_2, i_10_3, i_10_4, i_10_5, i_10_6, i_10_7, i_10_8, i_10_9, i_10_10, i_10_11, i_10_12, i_10_13, i_10_14, i_10_15, i_10_16, i_10_17, i_10_18, i_10_19, i_10_20, i_10_21, i_10_22, i_10_23, i_10_24, i_10_25, i_10_26, i_10_27, i_10_28, i_10_29, i_10_30, i_10_31, i_10_32, i_10_33, i_10_34, i_10_35, i_10_36, i_10_37, i_10_38, i_10_39, i_10_40, i_10_41, i_10_42, i_10_43, i_10_44, i_10_45, i_10_46, i_10_47, i_10_48, i_10_49, i_10_50, i_10_51, i_10_52, i_10_53, i_10_54, i_10_55, i_10_56, i_10_57, i_10_58, i_10_59, i_10_60, i_10_61, i_10_62, i_10_63, i_10_64, i_10_65, i_10_66, i_10_67, i_10_68, i_10_69, i_10_70, i_10_71, i_10_72, i_10_73, i_10_74, i_10_75, i_10_76, i_10_77, i_10_78, i_10_79, i_10_80, i_10_81, i_10_82, i_10_83, i_10_84, i_10_85, i_10_86, i_10_87, i_10_88, i_10_89, i_10_90, i_10_91, i_10_92, i_10_93, i_10_94, i_10_95, i_10_96, i_10_97, i_10_98, i_10_99, i_10_100, i_10_101, i_10_102, i_10_103, i_10_104, i_10_105, i_10_106, i_10_107, i_10_108, i_10_109, i_10_110, i_10_111, i_10_112, i_10_113, i_10_114, i_10_115, i_10_116, i_10_117, i_10_118, i_10_119, i_10_120, i_10_121, i_10_122, i_10_123, i_10_124, i_10_125, i_10_126, i_10_127, i_10_128, i_10_129, i_10_130, i_10_131, i_10_132, i_10_133, i_10_134, i_10_135, i_10_136, i_10_137, i_10_138, i_10_139, i_10_140, i_10_141, i_10_142, i_10_143, i_10_144, i_10_145, i_10_146, i_10_147, i_10_148, i_10_149, i_10_150, i_10_151, i_10_152, i_10_153, i_10_154, i_10_155, i_10_156, i_10_157, i_10_158, i_10_159, i_10_160, i_10_161, i_10_162, i_10_163, i_10_164, i_10_165, i_10_166, i_10_167, i_10_168, i_10_169, i_10_170, i_10_171, i_10_172, i_10_173, i_10_174, i_10_175, i_10_176, i_10_177, i_10_178, i_10_179, i_10_180, i_10_181, i_10_182, i_10_183, i_10_184, i_10_185, i_10_186, i_10_187, i_10_188, i_10_189, i_10_190, i_10_191, i_10_192, i_10_193, i_10_194, i_10_195, i_10_196, i_10_197, i_10_198, i_10_199, i_10_200, i_10_201, i_10_202, i_10_203, i_10_204, i_10_205, i_10_206, i_10_207, i_10_208, i_10_209, i_10_210, i_10_211, i_10_212, i_10_213, i_10_214, i_10_215, i_10_216, i_10_217, i_10_218, i_10_219, i_10_220, i_10_221, i_10_222, i_10_223, i_10_224, i_10_225, i_10_226, i_10_227, i_10_228, i_10_229, i_10_230, i_10_231, i_10_232, i_10_233, i_10_234, i_10_235, i_10_236, i_10_237, i_10_238, i_10_239, i_10_240, i_10_241, i_10_242, i_10_243, i_10_244, i_10_245, i_10_246, i_10_247, i_10_248, i_10_249, i_10_250, i_10_251, i_10_252, i_10_253, i_10_254, i_10_255, i_10_256, i_10_257, i_10_258, i_10_259, i_10_260, i_10_261, i_10_262, i_10_263, i_10_264, i_10_265, i_10_266, i_10_267, i_10_268, i_10_269, i_10_270, i_10_271, i_10_272, i_10_273, i_10_274, i_10_275, i_10_276, i_10_277, i_10_278, i_10_279, i_10_280, i_10_281, i_10_282, i_10_283, i_10_284, i_10_285, i_10_286, i_10_287, i_10_288, i_10_289, i_10_290, i_10_291, i_10_292, i_10_293, i_10_294, i_10_295, i_10_296, i_10_297, i_10_298, i_10_299, i_10_300, i_10_301, i_10_302, i_10_303, i_10_304, i_10_305, i_10_306, i_10_307, i_10_308, i_10_309, i_10_310, i_10_311, i_10_312, i_10_313, i_10_314, i_10_315, i_10_316, i_10_317, i_10_318, i_10_319, i_10_320, i_10_321, i_10_322, i_10_323, i_10_324, i_10_325, i_10_326, i_10_327, i_10_328, i_10_329, i_10_330, i_10_331, i_10_332, i_10_333, i_10_334, i_10_335, i_10_336, i_10_337, i_10_338, i_10_339, i_10_340, i_10_341, i_10_342, i_10_343, i_10_344, i_10_345, i_10_346, i_10_347, i_10_348, i_10_349, i_10_350, i_10_351, i_10_352, i_10_353, i_10_354, i_10_355, i_10_356, i_10_357, i_10_358, i_10_359, i_10_360, i_10_361, i_10_362, i_10_363, i_10_364, i_10_365, i_10_366, i_10_367, i_10_368, i_10_369, i_10_370, i_10_371, i_10_372, i_10_373, i_10_374, i_10_375, i_10_376, i_10_377, i_10_378, i_10_379, i_10_380, i_10_381, i_10_382, i_10_383, i_10_384, i_10_385, i_10_386, i_10_387, i_10_388, i_10_389, i_10_390, i_10_391, i_10_392, i_10_393, i_10_394, i_10_395, i_10_396, i_10_397, i_10_398, i_10_399, i_10_400, i_10_401, i_10_402, i_10_403, i_10_404, i_10_405, i_10_406, i_10_407, i_10_408, i_10_409, i_10_410, i_10_411, i_10_412, i_10_413, i_10_414, i_10_415, i_10_416, i_10_417, i_10_418, i_10_419, i_10_420, i_10_421, i_10_422, i_10_423, i_10_424, i_10_425, i_10_426, i_10_427, i_10_428, i_10_429, i_10_430, i_10_431, i_10_432, i_10_433, i_10_434, i_10_435, i_10_436, i_10_437, i_10_438, i_10_439, i_10_440, i_10_441, i_10_442, i_10_443, i_10_444, i_10_445, i_10_446, i_10_447, i_10_448, i_10_449, i_10_450, i_10_451, i_10_452, i_10_453, i_10_454, i_10_455, i_10_456, i_10_457, i_10_458, i_10_459, i_10_460, i_10_461, i_10_462, i_10_463, i_10_464, i_10_465, i_10_466, i_10_467, i_10_468, i_10_469, i_10_470, i_10_471, i_10_472, i_10_473, i_10_474, i_10_475, i_10_476, i_10_477, i_10_478, i_10_479, i_10_480, i_10_481, i_10_482, i_10_483, i_10_484, i_10_485, i_10_486, i_10_487, i_10_488, i_10_489, i_10_490, i_10_491, i_10_492, i_10_493, i_10_494, i_10_495, i_10_496, i_10_497, i_10_498, i_10_499, i_10_500, i_10_501, i_10_502, i_10_503, i_10_504, i_10_505, i_10_506, i_10_507, i_10_508, i_10_509, i_10_510, i_10_511, i_10_512, i_10_513, i_10_514, i_10_515, i_10_516, i_10_517, i_10_518, i_10_519, i_10_520, i_10_521, i_10_522, i_10_523, i_10_524, i_10_525, i_10_526, i_10_527, i_10_528, i_10_529, i_10_530, i_10_531, i_10_532, i_10_533, i_10_534, i_10_535, i_10_536, i_10_537, i_10_538, i_10_539, i_10_540, i_10_541, i_10_542, i_10_543, i_10_544, i_10_545, i_10_546, i_10_547, i_10_548, i_10_549, i_10_550, i_10_551, i_10_552, i_10_553, i_10_554, i_10_555, i_10_556, i_10_557, i_10_558, i_10_559, i_10_560, i_10_561, i_10_562, i_10_563, i_10_564, i_10_565, i_10_566, i_10_567, i_10_568, i_10_569, i_10_570, i_10_571, i_10_572, i_10_573, i_10_574, i_10_575, i_10_576, i_10_577, i_10_578, i_10_579, i_10_580, i_10_581, i_10_582, i_10_583, i_10_584, i_10_585, i_10_586, i_10_587, i_10_588, i_10_589, i_10_590, i_10_591, i_10_592, i_10_593, i_10_594, i_10_595, i_10_596, i_10_597, i_10_598, i_10_599, i_10_600, i_10_601, i_10_602, i_10_603, i_10_604, i_10_605, i_10_606, i_10_607, i_10_608, i_10_609, i_10_610, i_10_611, i_10_612, i_10_613, i_10_614, i_10_615, i_10_616, i_10_617, i_10_618, i_10_619, i_10_620, i_10_621, i_10_622, i_10_623, i_10_624, i_10_625, i_10_626, i_10_627, i_10_628, i_10_629, i_10_630, i_10_631, i_10_632, i_10_633, i_10_634, i_10_635, i_10_636, i_10_637, i_10_638, i_10_639, i_10_640, i_10_641, i_10_642, i_10_643, i_10_644, i_10_645, i_10_646, i_10_647, i_10_648, i_10_649, i_10_650, i_10_651, i_10_652, i_10_653, i_10_654, i_10_655, i_10_656, i_10_657, i_10_658, i_10_659, i_10_660, i_10_661, i_10_662, i_10_663, i_10_664, i_10_665, i_10_666, i_10_667, i_10_668, i_10_669, i_10_670, i_10_671, i_10_672, i_10_673, i_10_674, i_10_675, i_10_676, i_10_677, i_10_678, i_10_679, i_10_680, i_10_681, i_10_682, i_10_683, i_10_684, i_10_685, i_10_686, i_10_687, i_10_688, i_10_689, i_10_690, i_10_691, i_10_692, i_10_693, i_10_694, i_10_695, i_10_696, i_10_697, i_10_698, i_10_699, i_10_700, i_10_701, i_10_702, i_10_703, i_10_704, i_10_705, i_10_706, i_10_707, i_10_708, i_10_709, i_10_710, i_10_711, i_10_712, i_10_713, i_10_714, i_10_715, i_10_716, i_10_717, i_10_718, i_10_719, i_10_720, i_10_721, i_10_722, i_10_723, i_10_724, i_10_725, i_10_726, i_10_727, i_10_728, i_10_729, i_10_730, i_10_731, i_10_732, i_10_733, i_10_734, i_10_735, i_10_736, i_10_737, i_10_738, i_10_739, i_10_740, i_10_741, i_10_742, i_10_743, i_10_744, i_10_745, i_10_746, i_10_747, i_10_748, i_10_749, i_10_750, i_10_751, i_10_752, i_10_753, i_10_754, i_10_755, i_10_756, i_10_757, i_10_758, i_10_759, i_10_760, i_10_761, i_10_762, i_10_763, i_10_764, i_10_765, i_10_766, i_10_767, i_10_768, i_10_769, i_10_770, i_10_771, i_10_772, i_10_773, i_10_774, i_10_775, i_10_776, i_10_777, i_10_778, i_10_779, i_10_780, i_10_781, i_10_782, i_10_783, i_10_784, i_10_785, i_10_786, i_10_787, i_10_788, i_10_789, i_10_790, i_10_791, i_10_792, i_10_793, i_10_794, i_10_795, i_10_796, i_10_797, i_10_798, i_10_799, i_10_800, i_10_801, i_10_802, i_10_803, i_10_804, i_10_805, i_10_806, i_10_807, i_10_808, i_10_809, i_10_810, i_10_811, i_10_812, i_10_813, i_10_814, i_10_815, i_10_816, i_10_817, i_10_818, i_10_819, i_10_820, i_10_821, i_10_822, i_10_823, i_10_824, i_10_825, i_10_826, i_10_827, i_10_828, i_10_829, i_10_830, i_10_831, i_10_832, i_10_833, i_10_834, i_10_835, i_10_836, i_10_837, i_10_838, i_10_839, i_10_840, i_10_841, i_10_842, i_10_843, i_10_844, i_10_845, i_10_846, i_10_847, i_10_848, i_10_849, i_10_850, i_10_851, i_10_852, i_10_853, i_10_854, i_10_855, i_10_856, i_10_857, i_10_858, i_10_859, i_10_860, i_10_861, i_10_862, i_10_863, i_10_864, i_10_865, i_10_866, i_10_867, i_10_868, i_10_869, i_10_870, i_10_871, i_10_872, i_10_873, i_10_874, i_10_875, i_10_876, i_10_877, i_10_878, i_10_879, i_10_880, i_10_881, i_10_882, i_10_883, i_10_884, i_10_885, i_10_886, i_10_887, i_10_888, i_10_889, i_10_890, i_10_891, i_10_892, i_10_893, i_10_894, i_10_895, i_10_896, i_10_897, i_10_898, i_10_899, i_10_900, i_10_901, i_10_902, i_10_903, i_10_904, i_10_905, i_10_906, i_10_907, i_10_908, i_10_909, i_10_910, i_10_911, i_10_912, i_10_913, i_10_914, i_10_915, i_10_916, i_10_917, i_10_918, i_10_919, i_10_920, i_10_921, i_10_922, i_10_923, i_10_924, i_10_925, i_10_926, i_10_927, i_10_928, i_10_929, i_10_930, i_10_931, i_10_932, i_10_933, i_10_934, i_10_935, i_10_936, i_10_937, i_10_938, i_10_939, i_10_940, i_10_941, i_10_942, i_10_943, i_10_944, i_10_945, i_10_946, i_10_947, i_10_948, i_10_949, i_10_950, i_10_951, i_10_952, i_10_953, i_10_954, i_10_955, i_10_956, i_10_957, i_10_958, i_10_959, i_10_960, i_10_961, i_10_962, i_10_963, i_10_964, i_10_965, i_10_966, i_10_967, i_10_968, i_10_969, i_10_970, i_10_971, i_10_972, i_10_973, i_10_974, i_10_975, i_10_976, i_10_977, i_10_978, i_10_979, i_10_980, i_10_981, i_10_982, i_10_983, i_10_984, i_10_985, i_10_986, i_10_987, i_10_988, i_10_989, i_10_990, i_10_991, i_10_992, i_10_993, i_10_994, i_10_995, i_10_996, i_10_997, i_10_998, i_10_999, i_10_1000, i_10_1001, i_10_1002, i_10_1003, i_10_1004, i_10_1005, i_10_1006, i_10_1007, i_10_1008, i_10_1009, i_10_1010, i_10_1011, i_10_1012, i_10_1013, i_10_1014, i_10_1015, i_10_1016, i_10_1017, i_10_1018, i_10_1019, i_10_1020, i_10_1021, i_10_1022, i_10_1023, i_10_1024, i_10_1025, i_10_1026, i_10_1027, i_10_1028, i_10_1029, i_10_1030, i_10_1031, i_10_1032, i_10_1033, i_10_1034, i_10_1035, i_10_1036, i_10_1037, i_10_1038, i_10_1039, i_10_1040, i_10_1041, i_10_1042, i_10_1043, i_10_1044, i_10_1045, i_10_1046, i_10_1047, i_10_1048, i_10_1049, i_10_1050, i_10_1051, i_10_1052, i_10_1053, i_10_1054, i_10_1055, i_10_1056, i_10_1057, i_10_1058, i_10_1059, i_10_1060, i_10_1061, i_10_1062, i_10_1063, i_10_1064, i_10_1065, i_10_1066, i_10_1067, i_10_1068, i_10_1069, i_10_1070, i_10_1071, i_10_1072, i_10_1073, i_10_1074, i_10_1075, i_10_1076, i_10_1077, i_10_1078, i_10_1079, i_10_1080, i_10_1081, i_10_1082, i_10_1083, i_10_1084, i_10_1085, i_10_1086, i_10_1087, i_10_1088, i_10_1089, i_10_1090, i_10_1091, i_10_1092, i_10_1093, i_10_1094, i_10_1095, i_10_1096, i_10_1097, i_10_1098, i_10_1099, i_10_1100, i_10_1101, i_10_1102, i_10_1103, i_10_1104, i_10_1105, i_10_1106, i_10_1107, i_10_1108, i_10_1109, i_10_1110, i_10_1111, i_10_1112, i_10_1113, i_10_1114, i_10_1115, i_10_1116, i_10_1117, i_10_1118, i_10_1119, i_10_1120, i_10_1121, i_10_1122, i_10_1123, i_10_1124, i_10_1125, i_10_1126, i_10_1127, i_10_1128, i_10_1129, i_10_1130, i_10_1131, i_10_1132, i_10_1133, i_10_1134, i_10_1135, i_10_1136, i_10_1137, i_10_1138, i_10_1139, i_10_1140, i_10_1141, i_10_1142, i_10_1143, i_10_1144, i_10_1145, i_10_1146, i_10_1147, i_10_1148, i_10_1149, i_10_1150, i_10_1151, i_10_1152, i_10_1153, i_10_1154, i_10_1155, i_10_1156, i_10_1157, i_10_1158, i_10_1159, i_10_1160, i_10_1161, i_10_1162, i_10_1163, i_10_1164, i_10_1165, i_10_1166, i_10_1167, i_10_1168, i_10_1169, i_10_1170, i_10_1171, i_10_1172, i_10_1173, i_10_1174, i_10_1175, i_10_1176, i_10_1177, i_10_1178, i_10_1179, i_10_1180, i_10_1181, i_10_1182, i_10_1183, i_10_1184, i_10_1185, i_10_1186, i_10_1187, i_10_1188, i_10_1189, i_10_1190, i_10_1191, i_10_1192, i_10_1193, i_10_1194, i_10_1195, i_10_1196, i_10_1197, i_10_1198, i_10_1199, i_10_1200, i_10_1201, i_10_1202, i_10_1203, i_10_1204, i_10_1205, i_10_1206, i_10_1207, i_10_1208, i_10_1209, i_10_1210, i_10_1211, i_10_1212, i_10_1213, i_10_1214, i_10_1215, i_10_1216, i_10_1217, i_10_1218, i_10_1219, i_10_1220, i_10_1221, i_10_1222, i_10_1223, i_10_1224, i_10_1225, i_10_1226, i_10_1227, i_10_1228, i_10_1229, i_10_1230, i_10_1231, i_10_1232, i_10_1233, i_10_1234, i_10_1235, i_10_1236, i_10_1237, i_10_1238, i_10_1239, i_10_1240, i_10_1241, i_10_1242, i_10_1243, i_10_1244, i_10_1245, i_10_1246, i_10_1247, i_10_1248, i_10_1249, i_10_1250, i_10_1251, i_10_1252, i_10_1253, i_10_1254, i_10_1255, i_10_1256, i_10_1257, i_10_1258, i_10_1259, i_10_1260, i_10_1261, i_10_1262, i_10_1263, i_10_1264, i_10_1265, i_10_1266, i_10_1267, i_10_1268, i_10_1269, i_10_1270, i_10_1271, i_10_1272, i_10_1273, i_10_1274, i_10_1275, i_10_1276, i_10_1277, i_10_1278, i_10_1279, i_10_1280, i_10_1281, i_10_1282, i_10_1283, i_10_1284, i_10_1285, i_10_1286, i_10_1287, i_10_1288, i_10_1289, i_10_1290, i_10_1291, i_10_1292, i_10_1293, i_10_1294, i_10_1295, i_10_1296, i_10_1297, i_10_1298, i_10_1299, i_10_1300, i_10_1301, i_10_1302, i_10_1303, i_10_1304, i_10_1305, i_10_1306, i_10_1307, i_10_1308, i_10_1309, i_10_1310, i_10_1311, i_10_1312, i_10_1313, i_10_1314, i_10_1315, i_10_1316, i_10_1317, i_10_1318, i_10_1319, i_10_1320, i_10_1321, i_10_1322, i_10_1323, i_10_1324, i_10_1325, i_10_1326, i_10_1327, i_10_1328, i_10_1329, i_10_1330, i_10_1331, i_10_1332, i_10_1333, i_10_1334, i_10_1335, i_10_1336, i_10_1337, i_10_1338, i_10_1339, i_10_1340, i_10_1341, i_10_1342, i_10_1343, i_10_1344, i_10_1345, i_10_1346, i_10_1347, i_10_1348, i_10_1349, i_10_1350, i_10_1351, i_10_1352, i_10_1353, i_10_1354, i_10_1355, i_10_1356, i_10_1357, i_10_1358, i_10_1359, i_10_1360, i_10_1361, i_10_1362, i_10_1363, i_10_1364, i_10_1365, i_10_1366, i_10_1367, i_10_1368, i_10_1369, i_10_1370, i_10_1371, i_10_1372, i_10_1373, i_10_1374, i_10_1375, i_10_1376, i_10_1377, i_10_1378, i_10_1379, i_10_1380, i_10_1381, i_10_1382, i_10_1383, i_10_1384, i_10_1385, i_10_1386, i_10_1387, i_10_1388, i_10_1389, i_10_1390, i_10_1391, i_10_1392, i_10_1393, i_10_1394, i_10_1395, i_10_1396, i_10_1397, i_10_1398, i_10_1399, i_10_1400, i_10_1401, i_10_1402, i_10_1403, i_10_1404, i_10_1405, i_10_1406, i_10_1407, i_10_1408, i_10_1409, i_10_1410, i_10_1411, i_10_1412, i_10_1413, i_10_1414, i_10_1415, i_10_1416, i_10_1417, i_10_1418, i_10_1419, i_10_1420, i_10_1421, i_10_1422, i_10_1423, i_10_1424, i_10_1425, i_10_1426, i_10_1427, i_10_1428, i_10_1429, i_10_1430, i_10_1431, i_10_1432, i_10_1433, i_10_1434, i_10_1435, i_10_1436, i_10_1437, i_10_1438, i_10_1439, i_10_1440, i_10_1441, i_10_1442, i_10_1443, i_10_1444, i_10_1445, i_10_1446, i_10_1447, i_10_1448, i_10_1449, i_10_1450, i_10_1451, i_10_1452, i_10_1453, i_10_1454, i_10_1455, i_10_1456, i_10_1457, i_10_1458, i_10_1459, i_10_1460, i_10_1461, i_10_1462, i_10_1463, i_10_1464, i_10_1465, i_10_1466, i_10_1467, i_10_1468, i_10_1469, i_10_1470, i_10_1471, i_10_1472, i_10_1473, i_10_1474, i_10_1475, i_10_1476, i_10_1477, i_10_1478, i_10_1479, i_10_1480, i_10_1481, i_10_1482, i_10_1483, i_10_1484, i_10_1485, i_10_1486, i_10_1487, i_10_1488, i_10_1489, i_10_1490, i_10_1491, i_10_1492, i_10_1493, i_10_1494, i_10_1495, i_10_1496, i_10_1497, i_10_1498, i_10_1499, i_10_1500, i_10_1501, i_10_1502, i_10_1503, i_10_1504, i_10_1505, i_10_1506, i_10_1507, i_10_1508, i_10_1509, i_10_1510, i_10_1511, i_10_1512, i_10_1513, i_10_1514, i_10_1515, i_10_1516, i_10_1517, i_10_1518, i_10_1519, i_10_1520, i_10_1521, i_10_1522, i_10_1523, i_10_1524, i_10_1525, i_10_1526, i_10_1527, i_10_1528, i_10_1529, i_10_1530, i_10_1531, i_10_1532, i_10_1533, i_10_1534, i_10_1535, i_10_1536, i_10_1537, i_10_1538, i_10_1539, i_10_1540, i_10_1541, i_10_1542, i_10_1543, i_10_1544, i_10_1545, i_10_1546, i_10_1547, i_10_1548, i_10_1549, i_10_1550, i_10_1551, i_10_1552, i_10_1553, i_10_1554, i_10_1555, i_10_1556, i_10_1557, i_10_1558, i_10_1559, i_10_1560, i_10_1561, i_10_1562, i_10_1563, i_10_1564, i_10_1565, i_10_1566, i_10_1567, i_10_1568, i_10_1569, i_10_1570, i_10_1571, i_10_1572, i_10_1573, i_10_1574, i_10_1575, i_10_1576, i_10_1577, i_10_1578, i_10_1579, i_10_1580, i_10_1581, i_10_1582, i_10_1583, i_10_1584, i_10_1585, i_10_1586, i_10_1587, i_10_1588, i_10_1589, i_10_1590, i_10_1591, i_10_1592, i_10_1593, i_10_1594, i_10_1595, i_10_1596, i_10_1597, i_10_1598, i_10_1599, i_10_1600, i_10_1601, i_10_1602, i_10_1603, i_10_1604, i_10_1605, i_10_1606, i_10_1607, i_10_1608, i_10_1609, i_10_1610, i_10_1611, i_10_1612, i_10_1613, i_10_1614, i_10_1615, i_10_1616, i_10_1617, i_10_1618, i_10_1619, i_10_1620, i_10_1621, i_10_1622, i_10_1623, i_10_1624, i_10_1625, i_10_1626, i_10_1627, i_10_1628, i_10_1629, i_10_1630, i_10_1631, i_10_1632, i_10_1633, i_10_1634, i_10_1635, i_10_1636, i_10_1637, i_10_1638, i_10_1639, i_10_1640, i_10_1641, i_10_1642, i_10_1643, i_10_1644, i_10_1645, i_10_1646, i_10_1647, i_10_1648, i_10_1649, i_10_1650, i_10_1651, i_10_1652, i_10_1653, i_10_1654, i_10_1655, i_10_1656, i_10_1657, i_10_1658, i_10_1659, i_10_1660, i_10_1661, i_10_1662, i_10_1663, i_10_1664, i_10_1665, i_10_1666, i_10_1667, i_10_1668, i_10_1669, i_10_1670, i_10_1671, i_10_1672, i_10_1673, i_10_1674, i_10_1675, i_10_1676, i_10_1677, i_10_1678, i_10_1679, i_10_1680, i_10_1681, i_10_1682, i_10_1683, i_10_1684, i_10_1685, i_10_1686, i_10_1687, i_10_1688, i_10_1689, i_10_1690, i_10_1691, i_10_1692, i_10_1693, i_10_1694, i_10_1695, i_10_1696, i_10_1697, i_10_1698, i_10_1699, i_10_1700, i_10_1701, i_10_1702, i_10_1703, i_10_1704, i_10_1705, i_10_1706, i_10_1707, i_10_1708, i_10_1709, i_10_1710, i_10_1711, i_10_1712, i_10_1713, i_10_1714, i_10_1715, i_10_1716, i_10_1717, i_10_1718, i_10_1719, i_10_1720, i_10_1721, i_10_1722, i_10_1723, i_10_1724, i_10_1725, i_10_1726, i_10_1727, i_10_1728, i_10_1729, i_10_1730, i_10_1731, i_10_1732, i_10_1733, i_10_1734, i_10_1735, i_10_1736, i_10_1737, i_10_1738, i_10_1739, i_10_1740, i_10_1741, i_10_1742, i_10_1743, i_10_1744, i_10_1745, i_10_1746, i_10_1747, i_10_1748, i_10_1749, i_10_1750, i_10_1751, i_10_1752, i_10_1753, i_10_1754, i_10_1755, i_10_1756, i_10_1757, i_10_1758, i_10_1759, i_10_1760, i_10_1761, i_10_1762, i_10_1763, i_10_1764, i_10_1765, i_10_1766, i_10_1767, i_10_1768, i_10_1769, i_10_1770, i_10_1771, i_10_1772, i_10_1773, i_10_1774, i_10_1775, i_10_1776, i_10_1777, i_10_1778, i_10_1779, i_10_1780, i_10_1781, i_10_1782, i_10_1783, i_10_1784, i_10_1785, i_10_1786, i_10_1787, i_10_1788, i_10_1789, i_10_1790, i_10_1791, i_10_1792, i_10_1793, i_10_1794, i_10_1795, i_10_1796, i_10_1797, i_10_1798, i_10_1799, i_10_1800, i_10_1801, i_10_1802, i_10_1803, i_10_1804, i_10_1805, i_10_1806, i_10_1807, i_10_1808, i_10_1809, i_10_1810, i_10_1811, i_10_1812, i_10_1813, i_10_1814, i_10_1815, i_10_1816, i_10_1817, i_10_1818, i_10_1819, i_10_1820, i_10_1821, i_10_1822, i_10_1823, i_10_1824, i_10_1825, i_10_1826, i_10_1827, i_10_1828, i_10_1829, i_10_1830, i_10_1831, i_10_1832, i_10_1833, i_10_1834, i_10_1835, i_10_1836, i_10_1837, i_10_1838, i_10_1839, i_10_1840, i_10_1841, i_10_1842, i_10_1843, i_10_1844, i_10_1845, i_10_1846, i_10_1847, i_10_1848, i_10_1849, i_10_1850, i_10_1851, i_10_1852, i_10_1853, i_10_1854, i_10_1855, i_10_1856, i_10_1857, i_10_1858, i_10_1859, i_10_1860, i_10_1861, i_10_1862, i_10_1863, i_10_1864, i_10_1865, i_10_1866, i_10_1867, i_10_1868, i_10_1869, i_10_1870, i_10_1871, i_10_1872, i_10_1873, i_10_1874, i_10_1875, i_10_1876, i_10_1877, i_10_1878, i_10_1879, i_10_1880, i_10_1881, i_10_1882, i_10_1883, i_10_1884, i_10_1885, i_10_1886, i_10_1887, i_10_1888, i_10_1889, i_10_1890, i_10_1891, i_10_1892, i_10_1893, i_10_1894, i_10_1895, i_10_1896, i_10_1897, i_10_1898, i_10_1899, i_10_1900, i_10_1901, i_10_1902, i_10_1903, i_10_1904, i_10_1905, i_10_1906, i_10_1907, i_10_1908, i_10_1909, i_10_1910, i_10_1911, i_10_1912, i_10_1913, i_10_1914, i_10_1915, i_10_1916, i_10_1917, i_10_1918, i_10_1919, i_10_1920, i_10_1921, i_10_1922, i_10_1923, i_10_1924, i_10_1925, i_10_1926, i_10_1927, i_10_1928, i_10_1929, i_10_1930, i_10_1931, i_10_1932, i_10_1933, i_10_1934, i_10_1935, i_10_1936, i_10_1937, i_10_1938, i_10_1939, i_10_1940, i_10_1941, i_10_1942, i_10_1943, i_10_1944, i_10_1945, i_10_1946, i_10_1947, i_10_1948, i_10_1949, i_10_1950, i_10_1951, i_10_1952, i_10_1953, i_10_1954, i_10_1955, i_10_1956, i_10_1957, i_10_1958, i_10_1959, i_10_1960, i_10_1961, i_10_1962, i_10_1963, i_10_1964, i_10_1965, i_10_1966, i_10_1967, i_10_1968, i_10_1969, i_10_1970, i_10_1971, i_10_1972, i_10_1973, i_10_1974, i_10_1975, i_10_1976, i_10_1977, i_10_1978, i_10_1979, i_10_1980, i_10_1981, i_10_1982, i_10_1983, i_10_1984, i_10_1985, i_10_1986, i_10_1987, i_10_1988, i_10_1989, i_10_1990, i_10_1991, i_10_1992, i_10_1993, i_10_1994, i_10_1995, i_10_1996, i_10_1997, i_10_1998, i_10_1999, i_10_2000, i_10_2001, i_10_2002, i_10_2003, i_10_2004, i_10_2005, i_10_2006, i_10_2007, i_10_2008, i_10_2009, i_10_2010, i_10_2011, i_10_2012, i_10_2013, i_10_2014, i_10_2015, i_10_2016, i_10_2017, i_10_2018, i_10_2019, i_10_2020, i_10_2021, i_10_2022, i_10_2023, i_10_2024, i_10_2025, i_10_2026, i_10_2027, i_10_2028, i_10_2029, i_10_2030, i_10_2031, i_10_2032, i_10_2033, i_10_2034, i_10_2035, i_10_2036, i_10_2037, i_10_2038, i_10_2039, i_10_2040, i_10_2041, i_10_2042, i_10_2043, i_10_2044, i_10_2045, i_10_2046, i_10_2047, i_10_2048, i_10_2049, i_10_2050, i_10_2051, i_10_2052, i_10_2053, i_10_2054, i_10_2055, i_10_2056, i_10_2057, i_10_2058, i_10_2059, i_10_2060, i_10_2061, i_10_2062, i_10_2063, i_10_2064, i_10_2065, i_10_2066, i_10_2067, i_10_2068, i_10_2069, i_10_2070, i_10_2071, i_10_2072, i_10_2073, i_10_2074, i_10_2075, i_10_2076, i_10_2077, i_10_2078, i_10_2079, i_10_2080, i_10_2081, i_10_2082, i_10_2083, i_10_2084, i_10_2085, i_10_2086, i_10_2087, i_10_2088, i_10_2089, i_10_2090, i_10_2091, i_10_2092, i_10_2093, i_10_2094, i_10_2095, i_10_2096, i_10_2097, i_10_2098, i_10_2099, i_10_2100, i_10_2101, i_10_2102, i_10_2103, i_10_2104, i_10_2105, i_10_2106, i_10_2107, i_10_2108, i_10_2109, i_10_2110, i_10_2111, i_10_2112, i_10_2113, i_10_2114, i_10_2115, i_10_2116, i_10_2117, i_10_2118, i_10_2119, i_10_2120, i_10_2121, i_10_2122, i_10_2123, i_10_2124, i_10_2125, i_10_2126, i_10_2127, i_10_2128, i_10_2129, i_10_2130, i_10_2131, i_10_2132, i_10_2133, i_10_2134, i_10_2135, i_10_2136, i_10_2137, i_10_2138, i_10_2139, i_10_2140, i_10_2141, i_10_2142, i_10_2143, i_10_2144, i_10_2145, i_10_2146, i_10_2147, i_10_2148, i_10_2149, i_10_2150, i_10_2151, i_10_2152, i_10_2153, i_10_2154, i_10_2155, i_10_2156, i_10_2157, i_10_2158, i_10_2159, i_10_2160, i_10_2161, i_10_2162, i_10_2163, i_10_2164, i_10_2165, i_10_2166, i_10_2167, i_10_2168, i_10_2169, i_10_2170, i_10_2171, i_10_2172, i_10_2173, i_10_2174, i_10_2175, i_10_2176, i_10_2177, i_10_2178, i_10_2179, i_10_2180, i_10_2181, i_10_2182, i_10_2183, i_10_2184, i_10_2185, i_10_2186, i_10_2187, i_10_2188, i_10_2189, i_10_2190, i_10_2191, i_10_2192, i_10_2193, i_10_2194, i_10_2195, i_10_2196, i_10_2197, i_10_2198, i_10_2199, i_10_2200, i_10_2201, i_10_2202, i_10_2203, i_10_2204, i_10_2205, i_10_2206, i_10_2207, i_10_2208, i_10_2209, i_10_2210, i_10_2211, i_10_2212, i_10_2213, i_10_2214, i_10_2215, i_10_2216, i_10_2217, i_10_2218, i_10_2219, i_10_2220, i_10_2221, i_10_2222, i_10_2223, i_10_2224, i_10_2225, i_10_2226, i_10_2227, i_10_2228, i_10_2229, i_10_2230, i_10_2231, i_10_2232, i_10_2233, i_10_2234, i_10_2235, i_10_2236, i_10_2237, i_10_2238, i_10_2239, i_10_2240, i_10_2241, i_10_2242, i_10_2243, i_10_2244, i_10_2245, i_10_2246, i_10_2247, i_10_2248, i_10_2249, i_10_2250, i_10_2251, i_10_2252, i_10_2253, i_10_2254, i_10_2255, i_10_2256, i_10_2257, i_10_2258, i_10_2259, i_10_2260, i_10_2261, i_10_2262, i_10_2263, i_10_2264, i_10_2265, i_10_2266, i_10_2267, i_10_2268, i_10_2269, i_10_2270, i_10_2271, i_10_2272, i_10_2273, i_10_2274, i_10_2275, i_10_2276, i_10_2277, i_10_2278, i_10_2279, i_10_2280, i_10_2281, i_10_2282, i_10_2283, i_10_2284, i_10_2285, i_10_2286, i_10_2287, i_10_2288, i_10_2289, i_10_2290, i_10_2291, i_10_2292, i_10_2293, i_10_2294, i_10_2295, i_10_2296, i_10_2297, i_10_2298, i_10_2299, i_10_2300, i_10_2301, i_10_2302, i_10_2303, i_10_2304, i_10_2305, i_10_2306, i_10_2307, i_10_2308, i_10_2309, i_10_2310, i_10_2311, i_10_2312, i_10_2313, i_10_2314, i_10_2315, i_10_2316, i_10_2317, i_10_2318, i_10_2319, i_10_2320, i_10_2321, i_10_2322, i_10_2323, i_10_2324, i_10_2325, i_10_2326, i_10_2327, i_10_2328, i_10_2329, i_10_2330, i_10_2331, i_10_2332, i_10_2333, i_10_2334, i_10_2335, i_10_2336, i_10_2337, i_10_2338, i_10_2339, i_10_2340, i_10_2341, i_10_2342, i_10_2343, i_10_2344, i_10_2345, i_10_2346, i_10_2347, i_10_2348, i_10_2349, i_10_2350, i_10_2351, i_10_2352, i_10_2353, i_10_2354, i_10_2355, i_10_2356, i_10_2357, i_10_2358, i_10_2359, i_10_2360, i_10_2361, i_10_2362, i_10_2363, i_10_2364, i_10_2365, i_10_2366, i_10_2367, i_10_2368, i_10_2369, i_10_2370, i_10_2371, i_10_2372, i_10_2373, i_10_2374, i_10_2375, i_10_2376, i_10_2377, i_10_2378, i_10_2379, i_10_2380, i_10_2381, i_10_2382, i_10_2383, i_10_2384, i_10_2385, i_10_2386, i_10_2387, i_10_2388, i_10_2389, i_10_2390, i_10_2391, i_10_2392, i_10_2393, i_10_2394, i_10_2395, i_10_2396, i_10_2397, i_10_2398, i_10_2399, i_10_2400, i_10_2401, i_10_2402, i_10_2403, i_10_2404, i_10_2405, i_10_2406, i_10_2407, i_10_2408, i_10_2409, i_10_2410, i_10_2411, i_10_2412, i_10_2413, i_10_2414, i_10_2415, i_10_2416, i_10_2417, i_10_2418, i_10_2419, i_10_2420, i_10_2421, i_10_2422, i_10_2423, i_10_2424, i_10_2425, i_10_2426, i_10_2427, i_10_2428, i_10_2429, i_10_2430, i_10_2431, i_10_2432, i_10_2433, i_10_2434, i_10_2435, i_10_2436, i_10_2437, i_10_2438, i_10_2439, i_10_2440, i_10_2441, i_10_2442, i_10_2443, i_10_2444, i_10_2445, i_10_2446, i_10_2447, i_10_2448, i_10_2449, i_10_2450, i_10_2451, i_10_2452, i_10_2453, i_10_2454, i_10_2455, i_10_2456, i_10_2457, i_10_2458, i_10_2459, i_10_2460, i_10_2461, i_10_2462, i_10_2463, i_10_2464, i_10_2465, i_10_2466, i_10_2467, i_10_2468, i_10_2469, i_10_2470, i_10_2471, i_10_2472, i_10_2473, i_10_2474, i_10_2475, i_10_2476, i_10_2477, i_10_2478, i_10_2479, i_10_2480, i_10_2481, i_10_2482, i_10_2483, i_10_2484, i_10_2485, i_10_2486, i_10_2487, i_10_2488, i_10_2489, i_10_2490, i_10_2491, i_10_2492, i_10_2493, i_10_2494, i_10_2495, i_10_2496, i_10_2497, i_10_2498, i_10_2499, i_10_2500, i_10_2501, i_10_2502, i_10_2503, i_10_2504, i_10_2505, i_10_2506, i_10_2507, i_10_2508, i_10_2509, i_10_2510, i_10_2511, i_10_2512, i_10_2513, i_10_2514, i_10_2515, i_10_2516, i_10_2517, i_10_2518, i_10_2519, i_10_2520, i_10_2521, i_10_2522, i_10_2523, i_10_2524, i_10_2525, i_10_2526, i_10_2527, i_10_2528, i_10_2529, i_10_2530, i_10_2531, i_10_2532, i_10_2533, i_10_2534, i_10_2535, i_10_2536, i_10_2537, i_10_2538, i_10_2539, i_10_2540, i_10_2541, i_10_2542, i_10_2543, i_10_2544, i_10_2545, i_10_2546, i_10_2547, i_10_2548, i_10_2549, i_10_2550, i_10_2551, i_10_2552, i_10_2553, i_10_2554, i_10_2555, i_10_2556, i_10_2557, i_10_2558, i_10_2559, i_10_2560, i_10_2561, i_10_2562, i_10_2563, i_10_2564, i_10_2565, i_10_2566, i_10_2567, i_10_2568, i_10_2569, i_10_2570, i_10_2571, i_10_2572, i_10_2573, i_10_2574, i_10_2575, i_10_2576, i_10_2577, i_10_2578, i_10_2579, i_10_2580, i_10_2581, i_10_2582, i_10_2583, i_10_2584, i_10_2585, i_10_2586, i_10_2587, i_10_2588, i_10_2589, i_10_2590, i_10_2591, i_10_2592, i_10_2593, i_10_2594, i_10_2595, i_10_2596, i_10_2597, i_10_2598, i_10_2599, i_10_2600, i_10_2601, i_10_2602, i_10_2603, i_10_2604, i_10_2605, i_10_2606, i_10_2607, i_10_2608, i_10_2609, i_10_2610, i_10_2611, i_10_2612, i_10_2613, i_10_2614, i_10_2615, i_10_2616, i_10_2617, i_10_2618, i_10_2619, i_10_2620, i_10_2621, i_10_2622, i_10_2623, i_10_2624, i_10_2625, i_10_2626, i_10_2627, i_10_2628, i_10_2629, i_10_2630, i_10_2631, i_10_2632, i_10_2633, i_10_2634, i_10_2635, i_10_2636, i_10_2637, i_10_2638, i_10_2639, i_10_2640, i_10_2641, i_10_2642, i_10_2643, i_10_2644, i_10_2645, i_10_2646, i_10_2647, i_10_2648, i_10_2649, i_10_2650, i_10_2651, i_10_2652, i_10_2653, i_10_2654, i_10_2655, i_10_2656, i_10_2657, i_10_2658, i_10_2659, i_10_2660, i_10_2661, i_10_2662, i_10_2663, i_10_2664, i_10_2665, i_10_2666, i_10_2667, i_10_2668, i_10_2669, i_10_2670, i_10_2671, i_10_2672, i_10_2673, i_10_2674, i_10_2675, i_10_2676, i_10_2677, i_10_2678, i_10_2679, i_10_2680, i_10_2681, i_10_2682, i_10_2683, i_10_2684, i_10_2685, i_10_2686, i_10_2687, i_10_2688, i_10_2689, i_10_2690, i_10_2691, i_10_2692, i_10_2693, i_10_2694, i_10_2695, i_10_2696, i_10_2697, i_10_2698, i_10_2699, i_10_2700, i_10_2701, i_10_2702, i_10_2703, i_10_2704, i_10_2705, i_10_2706, i_10_2707, i_10_2708, i_10_2709, i_10_2710, i_10_2711, i_10_2712, i_10_2713, i_10_2714, i_10_2715, i_10_2716, i_10_2717, i_10_2718, i_10_2719, i_10_2720, i_10_2721, i_10_2722, i_10_2723, i_10_2724, i_10_2725, i_10_2726, i_10_2727, i_10_2728, i_10_2729, i_10_2730, i_10_2731, i_10_2732, i_10_2733, i_10_2734, i_10_2735, i_10_2736, i_10_2737, i_10_2738, i_10_2739, i_10_2740, i_10_2741, i_10_2742, i_10_2743, i_10_2744, i_10_2745, i_10_2746, i_10_2747, i_10_2748, i_10_2749, i_10_2750, i_10_2751, i_10_2752, i_10_2753, i_10_2754, i_10_2755, i_10_2756, i_10_2757, i_10_2758, i_10_2759, i_10_2760, i_10_2761, i_10_2762, i_10_2763, i_10_2764, i_10_2765, i_10_2766, i_10_2767, i_10_2768, i_10_2769, i_10_2770, i_10_2771, i_10_2772, i_10_2773, i_10_2774, i_10_2775, i_10_2776, i_10_2777, i_10_2778, i_10_2779, i_10_2780, i_10_2781, i_10_2782, i_10_2783, i_10_2784, i_10_2785, i_10_2786, i_10_2787, i_10_2788, i_10_2789, i_10_2790, i_10_2791, i_10_2792, i_10_2793, i_10_2794, i_10_2795, i_10_2796, i_10_2797, i_10_2798, i_10_2799, i_10_2800, i_10_2801, i_10_2802, i_10_2803, i_10_2804, i_10_2805, i_10_2806, i_10_2807, i_10_2808, i_10_2809, i_10_2810, i_10_2811, i_10_2812, i_10_2813, i_10_2814, i_10_2815, i_10_2816, i_10_2817, i_10_2818, i_10_2819, i_10_2820, i_10_2821, i_10_2822, i_10_2823, i_10_2824, i_10_2825, i_10_2826, i_10_2827, i_10_2828, i_10_2829, i_10_2830, i_10_2831, i_10_2832, i_10_2833, i_10_2834, i_10_2835, i_10_2836, i_10_2837, i_10_2838, i_10_2839, i_10_2840, i_10_2841, i_10_2842, i_10_2843, i_10_2844, i_10_2845, i_10_2846, i_10_2847, i_10_2848, i_10_2849, i_10_2850, i_10_2851, i_10_2852, i_10_2853, i_10_2854, i_10_2855, i_10_2856, i_10_2857, i_10_2858, i_10_2859, i_10_2860, i_10_2861, i_10_2862, i_10_2863, i_10_2864, i_10_2865, i_10_2866, i_10_2867, i_10_2868, i_10_2869, i_10_2870, i_10_2871, i_10_2872, i_10_2873, i_10_2874, i_10_2875, i_10_2876, i_10_2877, i_10_2878, i_10_2879, i_10_2880, i_10_2881, i_10_2882, i_10_2883, i_10_2884, i_10_2885, i_10_2886, i_10_2887, i_10_2888, i_10_2889, i_10_2890, i_10_2891, i_10_2892, i_10_2893, i_10_2894, i_10_2895, i_10_2896, i_10_2897, i_10_2898, i_10_2899, i_10_2900, i_10_2901, i_10_2902, i_10_2903, i_10_2904, i_10_2905, i_10_2906, i_10_2907, i_10_2908, i_10_2909, i_10_2910, i_10_2911, i_10_2912, i_10_2913, i_10_2914, i_10_2915, i_10_2916, i_10_2917, i_10_2918, i_10_2919, i_10_2920, i_10_2921, i_10_2922, i_10_2923, i_10_2924, i_10_2925, i_10_2926, i_10_2927, i_10_2928, i_10_2929, i_10_2930, i_10_2931, i_10_2932, i_10_2933, i_10_2934, i_10_2935, i_10_2936, i_10_2937, i_10_2938, i_10_2939, i_10_2940, i_10_2941, i_10_2942, i_10_2943, i_10_2944, i_10_2945, i_10_2946, i_10_2947, i_10_2948, i_10_2949, i_10_2950, i_10_2951, i_10_2952, i_10_2953, i_10_2954, i_10_2955, i_10_2956, i_10_2957, i_10_2958, i_10_2959, i_10_2960, i_10_2961, i_10_2962, i_10_2963, i_10_2964, i_10_2965, i_10_2966, i_10_2967, i_10_2968, i_10_2969, i_10_2970, i_10_2971, i_10_2972, i_10_2973, i_10_2974, i_10_2975, i_10_2976, i_10_2977, i_10_2978, i_10_2979, i_10_2980, i_10_2981, i_10_2982, i_10_2983, i_10_2984, i_10_2985, i_10_2986, i_10_2987, i_10_2988, i_10_2989, i_10_2990, i_10_2991, i_10_2992, i_10_2993, i_10_2994, i_10_2995, i_10_2996, i_10_2997, i_10_2998, i_10_2999, i_10_3000, i_10_3001, i_10_3002, i_10_3003, i_10_3004, i_10_3005, i_10_3006, i_10_3007, i_10_3008, i_10_3009, i_10_3010, i_10_3011, i_10_3012, i_10_3013, i_10_3014, i_10_3015, i_10_3016, i_10_3017, i_10_3018, i_10_3019, i_10_3020, i_10_3021, i_10_3022, i_10_3023, i_10_3024, i_10_3025, i_10_3026, i_10_3027, i_10_3028, i_10_3029, i_10_3030, i_10_3031, i_10_3032, i_10_3033, i_10_3034, i_10_3035, i_10_3036, i_10_3037, i_10_3038, i_10_3039, i_10_3040, i_10_3041, i_10_3042, i_10_3043, i_10_3044, i_10_3045, i_10_3046, i_10_3047, i_10_3048, i_10_3049, i_10_3050, i_10_3051, i_10_3052, i_10_3053, i_10_3054, i_10_3055, i_10_3056, i_10_3057, i_10_3058, i_10_3059, i_10_3060, i_10_3061, i_10_3062, i_10_3063, i_10_3064, i_10_3065, i_10_3066, i_10_3067, i_10_3068, i_10_3069, i_10_3070, i_10_3071, i_10_3072, i_10_3073, i_10_3074, i_10_3075, i_10_3076, i_10_3077, i_10_3078, i_10_3079, i_10_3080, i_10_3081, i_10_3082, i_10_3083, i_10_3084, i_10_3085, i_10_3086, i_10_3087, i_10_3088, i_10_3089, i_10_3090, i_10_3091, i_10_3092, i_10_3093, i_10_3094, i_10_3095, i_10_3096, i_10_3097, i_10_3098, i_10_3099, i_10_3100, i_10_3101, i_10_3102, i_10_3103, i_10_3104, i_10_3105, i_10_3106, i_10_3107, i_10_3108, i_10_3109, i_10_3110, i_10_3111, i_10_3112, i_10_3113, i_10_3114, i_10_3115, i_10_3116, i_10_3117, i_10_3118, i_10_3119, i_10_3120, i_10_3121, i_10_3122, i_10_3123, i_10_3124, i_10_3125, i_10_3126, i_10_3127, i_10_3128, i_10_3129, i_10_3130, i_10_3131, i_10_3132, i_10_3133, i_10_3134, i_10_3135, i_10_3136, i_10_3137, i_10_3138, i_10_3139, i_10_3140, i_10_3141, i_10_3142, i_10_3143, i_10_3144, i_10_3145, i_10_3146, i_10_3147, i_10_3148, i_10_3149, i_10_3150, i_10_3151, i_10_3152, i_10_3153, i_10_3154, i_10_3155, i_10_3156, i_10_3157, i_10_3158, i_10_3159, i_10_3160, i_10_3161, i_10_3162, i_10_3163, i_10_3164, i_10_3165, i_10_3166, i_10_3167, i_10_3168, i_10_3169, i_10_3170, i_10_3171, i_10_3172, i_10_3173, i_10_3174, i_10_3175, i_10_3176, i_10_3177, i_10_3178, i_10_3179, i_10_3180, i_10_3181, i_10_3182, i_10_3183, i_10_3184, i_10_3185, i_10_3186, i_10_3187, i_10_3188, i_10_3189, i_10_3190, i_10_3191, i_10_3192, i_10_3193, i_10_3194, i_10_3195, i_10_3196, i_10_3197, i_10_3198, i_10_3199, i_10_3200, i_10_3201, i_10_3202, i_10_3203, i_10_3204, i_10_3205, i_10_3206, i_10_3207, i_10_3208, i_10_3209, i_10_3210, i_10_3211, i_10_3212, i_10_3213, i_10_3214, i_10_3215, i_10_3216, i_10_3217, i_10_3218, i_10_3219, i_10_3220, i_10_3221, i_10_3222, i_10_3223, i_10_3224, i_10_3225, i_10_3226, i_10_3227, i_10_3228, i_10_3229, i_10_3230, i_10_3231, i_10_3232, i_10_3233, i_10_3234, i_10_3235, i_10_3236, i_10_3237, i_10_3238, i_10_3239, i_10_3240, i_10_3241, i_10_3242, i_10_3243, i_10_3244, i_10_3245, i_10_3246, i_10_3247, i_10_3248, i_10_3249, i_10_3250, i_10_3251, i_10_3252, i_10_3253, i_10_3254, i_10_3255, i_10_3256, i_10_3257, i_10_3258, i_10_3259, i_10_3260, i_10_3261, i_10_3262, i_10_3263, i_10_3264, i_10_3265, i_10_3266, i_10_3267, i_10_3268, i_10_3269, i_10_3270, i_10_3271, i_10_3272, i_10_3273, i_10_3274, i_10_3275, i_10_3276, i_10_3277, i_10_3278, i_10_3279, i_10_3280, i_10_3281, i_10_3282, i_10_3283, i_10_3284, i_10_3285, i_10_3286, i_10_3287, i_10_3288, i_10_3289, i_10_3290, i_10_3291, i_10_3292, i_10_3293, i_10_3294, i_10_3295, i_10_3296, i_10_3297, i_10_3298, i_10_3299, i_10_3300, i_10_3301, i_10_3302, i_10_3303, i_10_3304, i_10_3305, i_10_3306, i_10_3307, i_10_3308, i_10_3309, i_10_3310, i_10_3311, i_10_3312, i_10_3313, i_10_3314, i_10_3315, i_10_3316, i_10_3317, i_10_3318, i_10_3319, i_10_3320, i_10_3321, i_10_3322, i_10_3323, i_10_3324, i_10_3325, i_10_3326, i_10_3327, i_10_3328, i_10_3329, i_10_3330, i_10_3331, i_10_3332, i_10_3333, i_10_3334, i_10_3335, i_10_3336, i_10_3337, i_10_3338, i_10_3339, i_10_3340, i_10_3341, i_10_3342, i_10_3343, i_10_3344, i_10_3345, i_10_3346, i_10_3347, i_10_3348, i_10_3349, i_10_3350, i_10_3351, i_10_3352, i_10_3353, i_10_3354, i_10_3355, i_10_3356, i_10_3357, i_10_3358, i_10_3359, i_10_3360, i_10_3361, i_10_3362, i_10_3363, i_10_3364, i_10_3365, i_10_3366, i_10_3367, i_10_3368, i_10_3369, i_10_3370, i_10_3371, i_10_3372, i_10_3373, i_10_3374, i_10_3375, i_10_3376, i_10_3377, i_10_3378, i_10_3379, i_10_3380, i_10_3381, i_10_3382, i_10_3383, i_10_3384, i_10_3385, i_10_3386, i_10_3387, i_10_3388, i_10_3389, i_10_3390, i_10_3391, i_10_3392, i_10_3393, i_10_3394, i_10_3395, i_10_3396, i_10_3397, i_10_3398, i_10_3399, i_10_3400, i_10_3401, i_10_3402, i_10_3403, i_10_3404, i_10_3405, i_10_3406, i_10_3407, i_10_3408, i_10_3409, i_10_3410, i_10_3411, i_10_3412, i_10_3413, i_10_3414, i_10_3415, i_10_3416, i_10_3417, i_10_3418, i_10_3419, i_10_3420, i_10_3421, i_10_3422, i_10_3423, i_10_3424, i_10_3425, i_10_3426, i_10_3427, i_10_3428, i_10_3429, i_10_3430, i_10_3431, i_10_3432, i_10_3433, i_10_3434, i_10_3435, i_10_3436, i_10_3437, i_10_3438, i_10_3439, i_10_3440, i_10_3441, i_10_3442, i_10_3443, i_10_3444, i_10_3445, i_10_3446, i_10_3447, i_10_3448, i_10_3449, i_10_3450, i_10_3451, i_10_3452, i_10_3453, i_10_3454, i_10_3455, i_10_3456, i_10_3457, i_10_3458, i_10_3459, i_10_3460, i_10_3461, i_10_3462, i_10_3463, i_10_3464, i_10_3465, i_10_3466, i_10_3467, i_10_3468, i_10_3469, i_10_3470, i_10_3471, i_10_3472, i_10_3473, i_10_3474, i_10_3475, i_10_3476, i_10_3477, i_10_3478, i_10_3479, i_10_3480, i_10_3481, i_10_3482, i_10_3483, i_10_3484, i_10_3485, i_10_3486, i_10_3487, i_10_3488, i_10_3489, i_10_3490, i_10_3491, i_10_3492, i_10_3493, i_10_3494, i_10_3495, i_10_3496, i_10_3497, i_10_3498, i_10_3499, i_10_3500, i_10_3501, i_10_3502, i_10_3503, i_10_3504, i_10_3505, i_10_3506, i_10_3507, i_10_3508, i_10_3509, i_10_3510, i_10_3511, i_10_3512, i_10_3513, i_10_3514, i_10_3515, i_10_3516, i_10_3517, i_10_3518, i_10_3519, i_10_3520, i_10_3521, i_10_3522, i_10_3523, i_10_3524, i_10_3525, i_10_3526, i_10_3527, i_10_3528, i_10_3529, i_10_3530, i_10_3531, i_10_3532, i_10_3533, i_10_3534, i_10_3535, i_10_3536, i_10_3537, i_10_3538, i_10_3539, i_10_3540, i_10_3541, i_10_3542, i_10_3543, i_10_3544, i_10_3545, i_10_3546, i_10_3547, i_10_3548, i_10_3549, i_10_3550, i_10_3551, i_10_3552, i_10_3553, i_10_3554, i_10_3555, i_10_3556, i_10_3557, i_10_3558, i_10_3559, i_10_3560, i_10_3561, i_10_3562, i_10_3563, i_10_3564, i_10_3565, i_10_3566, i_10_3567, i_10_3568, i_10_3569, i_10_3570, i_10_3571, i_10_3572, i_10_3573, i_10_3574, i_10_3575, i_10_3576, i_10_3577, i_10_3578, i_10_3579, i_10_3580, i_10_3581, i_10_3582, i_10_3583, i_10_3584, i_10_3585, i_10_3586, i_10_3587, i_10_3588, i_10_3589, i_10_3590, i_10_3591, i_10_3592, i_10_3593, i_10_3594, i_10_3595, i_10_3596, i_10_3597, i_10_3598, i_10_3599, i_10_3600, i_10_3601, i_10_3602, i_10_3603, i_10_3604, i_10_3605, i_10_3606, i_10_3607, i_10_3608, i_10_3609, i_10_3610, i_10_3611, i_10_3612, i_10_3613, i_10_3614, i_10_3615, i_10_3616, i_10_3617, i_10_3618, i_10_3619, i_10_3620, i_10_3621, i_10_3622, i_10_3623, i_10_3624, i_10_3625, i_10_3626, i_10_3627, i_10_3628, i_10_3629, i_10_3630, i_10_3631, i_10_3632, i_10_3633, i_10_3634, i_10_3635, i_10_3636, i_10_3637, i_10_3638, i_10_3639, i_10_3640, i_10_3641, i_10_3642, i_10_3643, i_10_3644, i_10_3645, i_10_3646, i_10_3647, i_10_3648, i_10_3649, i_10_3650, i_10_3651, i_10_3652, i_10_3653, i_10_3654, i_10_3655, i_10_3656, i_10_3657, i_10_3658, i_10_3659, i_10_3660, i_10_3661, i_10_3662, i_10_3663, i_10_3664, i_10_3665, i_10_3666, i_10_3667, i_10_3668, i_10_3669, i_10_3670, i_10_3671, i_10_3672, i_10_3673, i_10_3674, i_10_3675, i_10_3676, i_10_3677, i_10_3678, i_10_3679, i_10_3680, i_10_3681, i_10_3682, i_10_3683, i_10_3684, i_10_3685, i_10_3686, i_10_3687, i_10_3688, i_10_3689, i_10_3690, i_10_3691, i_10_3692, i_10_3693, i_10_3694, i_10_3695, i_10_3696, i_10_3697, i_10_3698, i_10_3699, i_10_3700, i_10_3701, i_10_3702, i_10_3703, i_10_3704, i_10_3705, i_10_3706, i_10_3707, i_10_3708, i_10_3709, i_10_3710, i_10_3711, i_10_3712, i_10_3713, i_10_3714, i_10_3715, i_10_3716, i_10_3717, i_10_3718, i_10_3719, i_10_3720, i_10_3721, i_10_3722, i_10_3723, i_10_3724, i_10_3725, i_10_3726, i_10_3727, i_10_3728, i_10_3729, i_10_3730, i_10_3731, i_10_3732, i_10_3733, i_10_3734, i_10_3735, i_10_3736, i_10_3737, i_10_3738, i_10_3739, i_10_3740, i_10_3741, i_10_3742, i_10_3743, i_10_3744, i_10_3745, i_10_3746, i_10_3747, i_10_3748, i_10_3749, i_10_3750, i_10_3751, i_10_3752, i_10_3753, i_10_3754, i_10_3755, i_10_3756, i_10_3757, i_10_3758, i_10_3759, i_10_3760, i_10_3761, i_10_3762, i_10_3763, i_10_3764, i_10_3765, i_10_3766, i_10_3767, i_10_3768, i_10_3769, i_10_3770, i_10_3771, i_10_3772, i_10_3773, i_10_3774, i_10_3775, i_10_3776, i_10_3777, i_10_3778, i_10_3779, i_10_3780, i_10_3781, i_10_3782, i_10_3783, i_10_3784, i_10_3785, i_10_3786, i_10_3787, i_10_3788, i_10_3789, i_10_3790, i_10_3791, i_10_3792, i_10_3793, i_10_3794, i_10_3795, i_10_3796, i_10_3797, i_10_3798, i_10_3799, i_10_3800, i_10_3801, i_10_3802, i_10_3803, i_10_3804, i_10_3805, i_10_3806, i_10_3807, i_10_3808, i_10_3809, i_10_3810, i_10_3811, i_10_3812, i_10_3813, i_10_3814, i_10_3815, i_10_3816, i_10_3817, i_10_3818, i_10_3819, i_10_3820, i_10_3821, i_10_3822, i_10_3823, i_10_3824, i_10_3825, i_10_3826, i_10_3827, i_10_3828, i_10_3829, i_10_3830, i_10_3831, i_10_3832, i_10_3833, i_10_3834, i_10_3835, i_10_3836, i_10_3837, i_10_3838, i_10_3839, i_10_3840, i_10_3841, i_10_3842, i_10_3843, i_10_3844, i_10_3845, i_10_3846, i_10_3847, i_10_3848, i_10_3849, i_10_3850, i_10_3851, i_10_3852, i_10_3853, i_10_3854, i_10_3855, i_10_3856, i_10_3857, i_10_3858, i_10_3859, i_10_3860, i_10_3861, i_10_3862, i_10_3863, i_10_3864, i_10_3865, i_10_3866, i_10_3867, i_10_3868, i_10_3869, i_10_3870, i_10_3871, i_10_3872, i_10_3873, i_10_3874, i_10_3875, i_10_3876, i_10_3877, i_10_3878, i_10_3879, i_10_3880, i_10_3881, i_10_3882, i_10_3883, i_10_3884, i_10_3885, i_10_3886, i_10_3887, i_10_3888, i_10_3889, i_10_3890, i_10_3891, i_10_3892, i_10_3893, i_10_3894, i_10_3895, i_10_3896, i_10_3897, i_10_3898, i_10_3899, i_10_3900, i_10_3901, i_10_3902, i_10_3903, i_10_3904, i_10_3905, i_10_3906, i_10_3907, i_10_3908, i_10_3909, i_10_3910, i_10_3911, i_10_3912, i_10_3913, i_10_3914, i_10_3915, i_10_3916, i_10_3917, i_10_3918, i_10_3919, i_10_3920, i_10_3921, i_10_3922, i_10_3923, i_10_3924, i_10_3925, i_10_3926, i_10_3927, i_10_3928, i_10_3929, i_10_3930, i_10_3931, i_10_3932, i_10_3933, i_10_3934, i_10_3935, i_10_3936, i_10_3937, i_10_3938, i_10_3939, i_10_3940, i_10_3941, i_10_3942, i_10_3943, i_10_3944, i_10_3945, i_10_3946, i_10_3947, i_10_3948, i_10_3949, i_10_3950, i_10_3951, i_10_3952, i_10_3953, i_10_3954, i_10_3955, i_10_3956, i_10_3957, i_10_3958, i_10_3959, i_10_3960, i_10_3961, i_10_3962, i_10_3963, i_10_3964, i_10_3965, i_10_3966, i_10_3967, i_10_3968, i_10_3969, i_10_3970, i_10_3971, i_10_3972, i_10_3973, i_10_3974, i_10_3975, i_10_3976, i_10_3977, i_10_3978, i_10_3979, i_10_3980, i_10_3981, i_10_3982, i_10_3983, i_10_3984, i_10_3985, i_10_3986, i_10_3987, i_10_3988, i_10_3989, i_10_3990, i_10_3991, i_10_3992, i_10_3993, i_10_3994, i_10_3995, i_10_3996, i_10_3997, i_10_3998, i_10_3999, i_10_4000, i_10_4001, i_10_4002, i_10_4003, i_10_4004, i_10_4005, i_10_4006, i_10_4007, i_10_4008, i_10_4009, i_10_4010, i_10_4011, i_10_4012, i_10_4013, i_10_4014, i_10_4015, i_10_4016, i_10_4017, i_10_4018, i_10_4019, i_10_4020, i_10_4021, i_10_4022, i_10_4023, i_10_4024, i_10_4025, i_10_4026, i_10_4027, i_10_4028, i_10_4029, i_10_4030, i_10_4031, i_10_4032, i_10_4033, i_10_4034, i_10_4035, i_10_4036, i_10_4037, i_10_4038, i_10_4039, i_10_4040, i_10_4041, i_10_4042, i_10_4043, i_10_4044, i_10_4045, i_10_4046, i_10_4047, i_10_4048, i_10_4049, i_10_4050, i_10_4051, i_10_4052, i_10_4053, i_10_4054, i_10_4055, i_10_4056, i_10_4057, i_10_4058, i_10_4059, i_10_4060, i_10_4061, i_10_4062, i_10_4063, i_10_4064, i_10_4065, i_10_4066, i_10_4067, i_10_4068, i_10_4069, i_10_4070, i_10_4071, i_10_4072, i_10_4073, i_10_4074, i_10_4075, i_10_4076, i_10_4077, i_10_4078, i_10_4079, i_10_4080, i_10_4081, i_10_4082, i_10_4083, i_10_4084, i_10_4085, i_10_4086, i_10_4087, i_10_4088, i_10_4089, i_10_4090, i_10_4091, i_10_4092, i_10_4093, i_10_4094, i_10_4095, i_10_4096, i_10_4097, i_10_4098, i_10_4099, i_10_4100, i_10_4101, i_10_4102, i_10_4103, i_10_4104, i_10_4105, i_10_4106, i_10_4107, i_10_4108, i_10_4109, i_10_4110, i_10_4111, i_10_4112, i_10_4113, i_10_4114, i_10_4115, i_10_4116, i_10_4117, i_10_4118, i_10_4119, i_10_4120, i_10_4121, i_10_4122, i_10_4123, i_10_4124, i_10_4125, i_10_4126, i_10_4127, i_10_4128, i_10_4129, i_10_4130, i_10_4131, i_10_4132, i_10_4133, i_10_4134, i_10_4135, i_10_4136, i_10_4137, i_10_4138, i_10_4139, i_10_4140, i_10_4141, i_10_4142, i_10_4143, i_10_4144, i_10_4145, i_10_4146, i_10_4147, i_10_4148, i_10_4149, i_10_4150, i_10_4151, i_10_4152, i_10_4153, i_10_4154, i_10_4155, i_10_4156, i_10_4157, i_10_4158, i_10_4159, i_10_4160, i_10_4161, i_10_4162, i_10_4163, i_10_4164, i_10_4165, i_10_4166, i_10_4167, i_10_4168, i_10_4169, i_10_4170, i_10_4171, i_10_4172, i_10_4173, i_10_4174, i_10_4175, i_10_4176, i_10_4177, i_10_4178, i_10_4179, i_10_4180, i_10_4181, i_10_4182, i_10_4183, i_10_4184, i_10_4185, i_10_4186, i_10_4187, i_10_4188, i_10_4189, i_10_4190, i_10_4191, i_10_4192, i_10_4193, i_10_4194, i_10_4195, i_10_4196, i_10_4197, i_10_4198, i_10_4199, i_10_4200, i_10_4201, i_10_4202, i_10_4203, i_10_4204, i_10_4205, i_10_4206, i_10_4207, i_10_4208, i_10_4209, i_10_4210, i_10_4211, i_10_4212, i_10_4213, i_10_4214, i_10_4215, i_10_4216, i_10_4217, i_10_4218, i_10_4219, i_10_4220, i_10_4221, i_10_4222, i_10_4223, i_10_4224, i_10_4225, i_10_4226, i_10_4227, i_10_4228, i_10_4229, i_10_4230, i_10_4231, i_10_4232, i_10_4233, i_10_4234, i_10_4235, i_10_4236, i_10_4237, i_10_4238, i_10_4239, i_10_4240, i_10_4241, i_10_4242, i_10_4243, i_10_4244, i_10_4245, i_10_4246, i_10_4247, i_10_4248, i_10_4249, i_10_4250, i_10_4251, i_10_4252, i_10_4253, i_10_4254, i_10_4255, i_10_4256, i_10_4257, i_10_4258, i_10_4259, i_10_4260, i_10_4261, i_10_4262, i_10_4263, i_10_4264, i_10_4265, i_10_4266, i_10_4267, i_10_4268, i_10_4269, i_10_4270, i_10_4271, i_10_4272, i_10_4273, i_10_4274, i_10_4275, i_10_4276, i_10_4277, i_10_4278, i_10_4279, i_10_4280, i_10_4281, i_10_4282, i_10_4283, i_10_4284, i_10_4285, i_10_4286, i_10_4287, i_10_4288, i_10_4289, i_10_4290, i_10_4291, i_10_4292, i_10_4293, i_10_4294, i_10_4295, i_10_4296, i_10_4297, i_10_4298, i_10_4299, i_10_4300, i_10_4301, i_10_4302, i_10_4303, i_10_4304, i_10_4305, i_10_4306, i_10_4307, i_10_4308, i_10_4309, i_10_4310, i_10_4311, i_10_4312, i_10_4313, i_10_4314, i_10_4315, i_10_4316, i_10_4317, i_10_4318, i_10_4319, i_10_4320, i_10_4321, i_10_4322, i_10_4323, i_10_4324, i_10_4325, i_10_4326, i_10_4327, i_10_4328, i_10_4329, i_10_4330, i_10_4331, i_10_4332, i_10_4333, i_10_4334, i_10_4335, i_10_4336, i_10_4337, i_10_4338, i_10_4339, i_10_4340, i_10_4341, i_10_4342, i_10_4343, i_10_4344, i_10_4345, i_10_4346, i_10_4347, i_10_4348, i_10_4349, i_10_4350, i_10_4351, i_10_4352, i_10_4353, i_10_4354, i_10_4355, i_10_4356, i_10_4357, i_10_4358, i_10_4359, i_10_4360, i_10_4361, i_10_4362, i_10_4363, i_10_4364, i_10_4365, i_10_4366, i_10_4367, i_10_4368, i_10_4369, i_10_4370, i_10_4371, i_10_4372, i_10_4373, i_10_4374, i_10_4375, i_10_4376, i_10_4377, i_10_4378, i_10_4379, i_10_4380, i_10_4381, i_10_4382, i_10_4383, i_10_4384, i_10_4385, i_10_4386, i_10_4387, i_10_4388, i_10_4389, i_10_4390, i_10_4391, i_10_4392, i_10_4393, i_10_4394, i_10_4395, i_10_4396, i_10_4397, i_10_4398, i_10_4399, i_10_4400, i_10_4401, i_10_4402, i_10_4403, i_10_4404, i_10_4405, i_10_4406, i_10_4407, i_10_4408, i_10_4409, i_10_4410, i_10_4411, i_10_4412, i_10_4413, i_10_4414, i_10_4415, i_10_4416, i_10_4417, i_10_4418, i_10_4419, i_10_4420, i_10_4421, i_10_4422, i_10_4423, i_10_4424, i_10_4425, i_10_4426, i_10_4427, i_10_4428, i_10_4429, i_10_4430, i_10_4431, i_10_4432, i_10_4433, i_10_4434, i_10_4435, i_10_4436, i_10_4437, i_10_4438, i_10_4439, i_10_4440, i_10_4441, i_10_4442, i_10_4443, i_10_4444, i_10_4445, i_10_4446, i_10_4447, i_10_4448, i_10_4449, i_10_4450, i_10_4451, i_10_4452, i_10_4453, i_10_4454, i_10_4455, i_10_4456, i_10_4457, i_10_4458, i_10_4459, i_10_4460, i_10_4461, i_10_4462, i_10_4463, i_10_4464, i_10_4465, i_10_4466, i_10_4467, i_10_4468, i_10_4469, i_10_4470, i_10_4471, i_10_4472, i_10_4473, i_10_4474, i_10_4475, i_10_4476, i_10_4477, i_10_4478, i_10_4479, i_10_4480, i_10_4481, i_10_4482, i_10_4483, i_10_4484, i_10_4485, i_10_4486, i_10_4487, i_10_4488, i_10_4489, i_10_4490, i_10_4491, i_10_4492, i_10_4493, i_10_4494, i_10_4495, i_10_4496, i_10_4497, i_10_4498, i_10_4499, i_10_4500, i_10_4501, i_10_4502, i_10_4503, i_10_4504, i_10_4505, i_10_4506, i_10_4507, i_10_4508, i_10_4509, i_10_4510, i_10_4511, i_10_4512, i_10_4513, i_10_4514, i_10_4515, i_10_4516, i_10_4517, i_10_4518, i_10_4519, i_10_4520, i_10_4521, i_10_4522, i_10_4523, i_10_4524, i_10_4525, i_10_4526, i_10_4527, i_10_4528, i_10_4529, i_10_4530, i_10_4531, i_10_4532, i_10_4533, i_10_4534, i_10_4535, i_10_4536, i_10_4537, i_10_4538, i_10_4539, i_10_4540, i_10_4541, i_10_4542, i_10_4543, i_10_4544, i_10_4545, i_10_4546, i_10_4547, i_10_4548, i_10_4549, i_10_4550, i_10_4551, i_10_4552, i_10_4553, i_10_4554, i_10_4555, i_10_4556, i_10_4557, i_10_4558, i_10_4559, i_10_4560, i_10_4561, i_10_4562, i_10_4563, i_10_4564, i_10_4565, i_10_4566, i_10_4567, i_10_4568, i_10_4569, i_10_4570, i_10_4571, i_10_4572, i_10_4573, i_10_4574, i_10_4575, i_10_4576, i_10_4577, i_10_4578, i_10_4579, i_10_4580, i_10_4581, i_10_4582, i_10_4583, i_10_4584, i_10_4585, i_10_4586, i_10_4587, i_10_4588, i_10_4589, i_10_4590, i_10_4591, i_10_4592, i_10_4593, i_10_4594, i_10_4595, i_10_4596, i_10_4597, i_10_4598, i_10_4599, i_10_4600, i_10_4601, i_10_4602, i_10_4603, i_10_4604, i_10_4605, i_10_4606, i_10_4607, o_10_0, o_10_1, o_10_2, o_10_3, o_10_4, o_10_5, o_10_6, o_10_7, o_10_8, o_10_9, o_10_10, o_10_11, o_10_12, o_10_13, o_10_14, o_10_15, o_10_16, o_10_17, o_10_18, o_10_19, o_10_20, o_10_21, o_10_22, o_10_23, o_10_24, o_10_25, o_10_26, o_10_27, o_10_28, o_10_29, o_10_30, o_10_31, o_10_32, o_10_33, o_10_34, o_10_35, o_10_36, o_10_37, o_10_38, o_10_39, o_10_40, o_10_41, o_10_42, o_10_43, o_10_44, o_10_45, o_10_46, o_10_47, o_10_48, o_10_49, o_10_50, o_10_51, o_10_52, o_10_53, o_10_54, o_10_55, o_10_56, o_10_57, o_10_58, o_10_59, o_10_60, o_10_61, o_10_62, o_10_63, o_10_64, o_10_65, o_10_66, o_10_67, o_10_68, o_10_69, o_10_70, o_10_71, o_10_72, o_10_73, o_10_74, o_10_75, o_10_76, o_10_77, o_10_78, o_10_79, o_10_80, o_10_81, o_10_82, o_10_83, o_10_84, o_10_85, o_10_86, o_10_87, o_10_88, o_10_89, o_10_90, o_10_91, o_10_92, o_10_93, o_10_94, o_10_95, o_10_96, o_10_97, o_10_98, o_10_99, o_10_100, o_10_101, o_10_102, o_10_103, o_10_104, o_10_105, o_10_106, o_10_107, o_10_108, o_10_109, o_10_110, o_10_111, o_10_112, o_10_113, o_10_114, o_10_115, o_10_116, o_10_117, o_10_118, o_10_119, o_10_120, o_10_121, o_10_122, o_10_123, o_10_124, o_10_125, o_10_126, o_10_127, o_10_128, o_10_129, o_10_130, o_10_131, o_10_132, o_10_133, o_10_134, o_10_135, o_10_136, o_10_137, o_10_138, o_10_139, o_10_140, o_10_141, o_10_142, o_10_143, o_10_144, o_10_145, o_10_146, o_10_147, o_10_148, o_10_149, o_10_150, o_10_151, o_10_152, o_10_153, o_10_154, o_10_155, o_10_156, o_10_157, o_10_158, o_10_159, o_10_160, o_10_161, o_10_162, o_10_163, o_10_164, o_10_165, o_10_166, o_10_167, o_10_168, o_10_169, o_10_170, o_10_171, o_10_172, o_10_173, o_10_174, o_10_175, o_10_176, o_10_177, o_10_178, o_10_179, o_10_180, o_10_181, o_10_182, o_10_183, o_10_184, o_10_185, o_10_186, o_10_187, o_10_188, o_10_189, o_10_190, o_10_191, o_10_192, o_10_193, o_10_194, o_10_195, o_10_196, o_10_197, o_10_198, o_10_199, o_10_200, o_10_201, o_10_202, o_10_203, o_10_204, o_10_205, o_10_206, o_10_207, o_10_208, o_10_209, o_10_210, o_10_211, o_10_212, o_10_213, o_10_214, o_10_215, o_10_216, o_10_217, o_10_218, o_10_219, o_10_220, o_10_221, o_10_222, o_10_223, o_10_224, o_10_225, o_10_226, o_10_227, o_10_228, o_10_229, o_10_230, o_10_231, o_10_232, o_10_233, o_10_234, o_10_235, o_10_236, o_10_237, o_10_238, o_10_239, o_10_240, o_10_241, o_10_242, o_10_243, o_10_244, o_10_245, o_10_246, o_10_247, o_10_248, o_10_249, o_10_250, o_10_251, o_10_252, o_10_253, o_10_254, o_10_255, o_10_256, o_10_257, o_10_258, o_10_259, o_10_260, o_10_261, o_10_262, o_10_263, o_10_264, o_10_265, o_10_266, o_10_267, o_10_268, o_10_269, o_10_270, o_10_271, o_10_272, o_10_273, o_10_274, o_10_275, o_10_276, o_10_277, o_10_278, o_10_279, o_10_280, o_10_281, o_10_282, o_10_283, o_10_284, o_10_285, o_10_286, o_10_287, o_10_288, o_10_289, o_10_290, o_10_291, o_10_292, o_10_293, o_10_294, o_10_295, o_10_296, o_10_297, o_10_298, o_10_299, o_10_300, o_10_301, o_10_302, o_10_303, o_10_304, o_10_305, o_10_306, o_10_307, o_10_308, o_10_309, o_10_310, o_10_311, o_10_312, o_10_313, o_10_314, o_10_315, o_10_316, o_10_317, o_10_318, o_10_319, o_10_320, o_10_321, o_10_322, o_10_323, o_10_324, o_10_325, o_10_326, o_10_327, o_10_328, o_10_329, o_10_330, o_10_331, o_10_332, o_10_333, o_10_334, o_10_335, o_10_336, o_10_337, o_10_338, o_10_339, o_10_340, o_10_341, o_10_342, o_10_343, o_10_344, o_10_345, o_10_346, o_10_347, o_10_348, o_10_349, o_10_350, o_10_351, o_10_352, o_10_353, o_10_354, o_10_355, o_10_356, o_10_357, o_10_358, o_10_359, o_10_360, o_10_361, o_10_362, o_10_363, o_10_364, o_10_365, o_10_366, o_10_367, o_10_368, o_10_369, o_10_370, o_10_371, o_10_372, o_10_373, o_10_374, o_10_375, o_10_376, o_10_377, o_10_378, o_10_379, o_10_380, o_10_381, o_10_382, o_10_383, o_10_384, o_10_385, o_10_386, o_10_387, o_10_388, o_10_389, o_10_390, o_10_391, o_10_392, o_10_393, o_10_394, o_10_395, o_10_396, o_10_397, o_10_398, o_10_399, o_10_400, o_10_401, o_10_402, o_10_403, o_10_404, o_10_405, o_10_406, o_10_407, o_10_408, o_10_409, o_10_410, o_10_411, o_10_412, o_10_413, o_10_414, o_10_415, o_10_416, o_10_417, o_10_418, o_10_419, o_10_420, o_10_421, o_10_422, o_10_423, o_10_424, o_10_425, o_10_426, o_10_427, o_10_428, o_10_429, o_10_430, o_10_431, o_10_432, o_10_433, o_10_434, o_10_435, o_10_436, o_10_437, o_10_438, o_10_439, o_10_440, o_10_441, o_10_442, o_10_443, o_10_444, o_10_445, o_10_446, o_10_447, o_10_448, o_10_449, o_10_450, o_10_451, o_10_452, o_10_453, o_10_454, o_10_455, o_10_456, o_10_457, o_10_458, o_10_459, o_10_460, o_10_461, o_10_462, o_10_463, o_10_464, o_10_465, o_10_466, o_10_467, o_10_468, o_10_469, o_10_470, o_10_471, o_10_472, o_10_473, o_10_474, o_10_475, o_10_476, o_10_477, o_10_478, o_10_479, o_10_480, o_10_481, o_10_482, o_10_483, o_10_484, o_10_485, o_10_486, o_10_487, o_10_488, o_10_489, o_10_490, o_10_491, o_10_492, o_10_493, o_10_494, o_10_495, o_10_496, o_10_497, o_10_498, o_10_499, o_10_500, o_10_501, o_10_502, o_10_503, o_10_504, o_10_505, o_10_506, o_10_507, o_10_508, o_10_509, o_10_510, o_10_511);

  always @ (posedge ap_clk)
    if (ap_rst)
      begin
        out_reg <= 0;
        i_10_0 <= 0;
        i_10_1 <= 0;
        i_10_2 <= 0;
        i_10_3 <= 0;
        i_10_4 <= 0;
        i_10_5 <= 0;
        i_10_6 <= 0;
        i_10_7 <= 0;
        i_10_8 <= 0;
        i_10_9 <= 0;
        i_10_10 <= 0;
        i_10_11 <= 0;
        i_10_12 <= 0;
        i_10_13 <= 0;
        i_10_14 <= 0;
        i_10_15 <= 0;
        i_10_16 <= 0;
        i_10_17 <= 0;
        i_10_18 <= 0;
        i_10_19 <= 0;
        i_10_20 <= 0;
        i_10_21 <= 0;
        i_10_22 <= 0;
        i_10_23 <= 0;
        i_10_24 <= 0;
        i_10_25 <= 0;
        i_10_26 <= 0;
        i_10_27 <= 0;
        i_10_28 <= 0;
        i_10_29 <= 0;
        i_10_30 <= 0;
        i_10_31 <= 0;
        i_10_32 <= 0;
        i_10_33 <= 0;
        i_10_34 <= 0;
        i_10_35 <= 0;
        i_10_36 <= 0;
        i_10_37 <= 0;
        i_10_38 <= 0;
        i_10_39 <= 0;
        i_10_40 <= 0;
        i_10_41 <= 0;
        i_10_42 <= 0;
        i_10_43 <= 0;
        i_10_44 <= 0;
        i_10_45 <= 0;
        i_10_46 <= 0;
        i_10_47 <= 0;
        i_10_48 <= 0;
        i_10_49 <= 0;
        i_10_50 <= 0;
        i_10_51 <= 0;
        i_10_52 <= 0;
        i_10_53 <= 0;
        i_10_54 <= 0;
        i_10_55 <= 0;
        i_10_56 <= 0;
        i_10_57 <= 0;
        i_10_58 <= 0;
        i_10_59 <= 0;
        i_10_60 <= 0;
        i_10_61 <= 0;
        i_10_62 <= 0;
        i_10_63 <= 0;
        i_10_64 <= 0;
        i_10_65 <= 0;
        i_10_66 <= 0;
        i_10_67 <= 0;
        i_10_68 <= 0;
        i_10_69 <= 0;
        i_10_70 <= 0;
        i_10_71 <= 0;
        i_10_72 <= 0;
        i_10_73 <= 0;
        i_10_74 <= 0;
        i_10_75 <= 0;
        i_10_76 <= 0;
        i_10_77 <= 0;
        i_10_78 <= 0;
        i_10_79 <= 0;
        i_10_80 <= 0;
        i_10_81 <= 0;
        i_10_82 <= 0;
        i_10_83 <= 0;
        i_10_84 <= 0;
        i_10_85 <= 0;
        i_10_86 <= 0;
        i_10_87 <= 0;
        i_10_88 <= 0;
        i_10_89 <= 0;
        i_10_90 <= 0;
        i_10_91 <= 0;
        i_10_92 <= 0;
        i_10_93 <= 0;
        i_10_94 <= 0;
        i_10_95 <= 0;
        i_10_96 <= 0;
        i_10_97 <= 0;
        i_10_98 <= 0;
        i_10_99 <= 0;
        i_10_100 <= 0;
        i_10_101 <= 0;
        i_10_102 <= 0;
        i_10_103 <= 0;
        i_10_104 <= 0;
        i_10_105 <= 0;
        i_10_106 <= 0;
        i_10_107 <= 0;
        i_10_108 <= 0;
        i_10_109 <= 0;
        i_10_110 <= 0;
        i_10_111 <= 0;
        i_10_112 <= 0;
        i_10_113 <= 0;
        i_10_114 <= 0;
        i_10_115 <= 0;
        i_10_116 <= 0;
        i_10_117 <= 0;
        i_10_118 <= 0;
        i_10_119 <= 0;
        i_10_120 <= 0;
        i_10_121 <= 0;
        i_10_122 <= 0;
        i_10_123 <= 0;
        i_10_124 <= 0;
        i_10_125 <= 0;
        i_10_126 <= 0;
        i_10_127 <= 0;
        i_10_128 <= 0;
        i_10_129 <= 0;
        i_10_130 <= 0;
        i_10_131 <= 0;
        i_10_132 <= 0;
        i_10_133 <= 0;
        i_10_134 <= 0;
        i_10_135 <= 0;
        i_10_136 <= 0;
        i_10_137 <= 0;
        i_10_138 <= 0;
        i_10_139 <= 0;
        i_10_140 <= 0;
        i_10_141 <= 0;
        i_10_142 <= 0;
        i_10_143 <= 0;
        i_10_144 <= 0;
        i_10_145 <= 0;
        i_10_146 <= 0;
        i_10_147 <= 0;
        i_10_148 <= 0;
        i_10_149 <= 0;
        i_10_150 <= 0;
        i_10_151 <= 0;
        i_10_152 <= 0;
        i_10_153 <= 0;
        i_10_154 <= 0;
        i_10_155 <= 0;
        i_10_156 <= 0;
        i_10_157 <= 0;
        i_10_158 <= 0;
        i_10_159 <= 0;
        i_10_160 <= 0;
        i_10_161 <= 0;
        i_10_162 <= 0;
        i_10_163 <= 0;
        i_10_164 <= 0;
        i_10_165 <= 0;
        i_10_166 <= 0;
        i_10_167 <= 0;
        i_10_168 <= 0;
        i_10_169 <= 0;
        i_10_170 <= 0;
        i_10_171 <= 0;
        i_10_172 <= 0;
        i_10_173 <= 0;
        i_10_174 <= 0;
        i_10_175 <= 0;
        i_10_176 <= 0;
        i_10_177 <= 0;
        i_10_178 <= 0;
        i_10_179 <= 0;
        i_10_180 <= 0;
        i_10_181 <= 0;
        i_10_182 <= 0;
        i_10_183 <= 0;
        i_10_184 <= 0;
        i_10_185 <= 0;
        i_10_186 <= 0;
        i_10_187 <= 0;
        i_10_188 <= 0;
        i_10_189 <= 0;
        i_10_190 <= 0;
        i_10_191 <= 0;
        i_10_192 <= 0;
        i_10_193 <= 0;
        i_10_194 <= 0;
        i_10_195 <= 0;
        i_10_196 <= 0;
        i_10_197 <= 0;
        i_10_198 <= 0;
        i_10_199 <= 0;
        i_10_200 <= 0;
        i_10_201 <= 0;
        i_10_202 <= 0;
        i_10_203 <= 0;
        i_10_204 <= 0;
        i_10_205 <= 0;
        i_10_206 <= 0;
        i_10_207 <= 0;
        i_10_208 <= 0;
        i_10_209 <= 0;
        i_10_210 <= 0;
        i_10_211 <= 0;
        i_10_212 <= 0;
        i_10_213 <= 0;
        i_10_214 <= 0;
        i_10_215 <= 0;
        i_10_216 <= 0;
        i_10_217 <= 0;
        i_10_218 <= 0;
        i_10_219 <= 0;
        i_10_220 <= 0;
        i_10_221 <= 0;
        i_10_222 <= 0;
        i_10_223 <= 0;
        i_10_224 <= 0;
        i_10_225 <= 0;
        i_10_226 <= 0;
        i_10_227 <= 0;
        i_10_228 <= 0;
        i_10_229 <= 0;
        i_10_230 <= 0;
        i_10_231 <= 0;
        i_10_232 <= 0;
        i_10_233 <= 0;
        i_10_234 <= 0;
        i_10_235 <= 0;
        i_10_236 <= 0;
        i_10_237 <= 0;
        i_10_238 <= 0;
        i_10_239 <= 0;
        i_10_240 <= 0;
        i_10_241 <= 0;
        i_10_242 <= 0;
        i_10_243 <= 0;
        i_10_244 <= 0;
        i_10_245 <= 0;
        i_10_246 <= 0;
        i_10_247 <= 0;
        i_10_248 <= 0;
        i_10_249 <= 0;
        i_10_250 <= 0;
        i_10_251 <= 0;
        i_10_252 <= 0;
        i_10_253 <= 0;
        i_10_254 <= 0;
        i_10_255 <= 0;
        i_10_256 <= 0;
        i_10_257 <= 0;
        i_10_258 <= 0;
        i_10_259 <= 0;
        i_10_260 <= 0;
        i_10_261 <= 0;
        i_10_262 <= 0;
        i_10_263 <= 0;
        i_10_264 <= 0;
        i_10_265 <= 0;
        i_10_266 <= 0;
        i_10_267 <= 0;
        i_10_268 <= 0;
        i_10_269 <= 0;
        i_10_270 <= 0;
        i_10_271 <= 0;
        i_10_272 <= 0;
        i_10_273 <= 0;
        i_10_274 <= 0;
        i_10_275 <= 0;
        i_10_276 <= 0;
        i_10_277 <= 0;
        i_10_278 <= 0;
        i_10_279 <= 0;
        i_10_280 <= 0;
        i_10_281 <= 0;
        i_10_282 <= 0;
        i_10_283 <= 0;
        i_10_284 <= 0;
        i_10_285 <= 0;
        i_10_286 <= 0;
        i_10_287 <= 0;
        i_10_288 <= 0;
        i_10_289 <= 0;
        i_10_290 <= 0;
        i_10_291 <= 0;
        i_10_292 <= 0;
        i_10_293 <= 0;
        i_10_294 <= 0;
        i_10_295 <= 0;
        i_10_296 <= 0;
        i_10_297 <= 0;
        i_10_298 <= 0;
        i_10_299 <= 0;
        i_10_300 <= 0;
        i_10_301 <= 0;
        i_10_302 <= 0;
        i_10_303 <= 0;
        i_10_304 <= 0;
        i_10_305 <= 0;
        i_10_306 <= 0;
        i_10_307 <= 0;
        i_10_308 <= 0;
        i_10_309 <= 0;
        i_10_310 <= 0;
        i_10_311 <= 0;
        i_10_312 <= 0;
        i_10_313 <= 0;
        i_10_314 <= 0;
        i_10_315 <= 0;
        i_10_316 <= 0;
        i_10_317 <= 0;
        i_10_318 <= 0;
        i_10_319 <= 0;
        i_10_320 <= 0;
        i_10_321 <= 0;
        i_10_322 <= 0;
        i_10_323 <= 0;
        i_10_324 <= 0;
        i_10_325 <= 0;
        i_10_326 <= 0;
        i_10_327 <= 0;
        i_10_328 <= 0;
        i_10_329 <= 0;
        i_10_330 <= 0;
        i_10_331 <= 0;
        i_10_332 <= 0;
        i_10_333 <= 0;
        i_10_334 <= 0;
        i_10_335 <= 0;
        i_10_336 <= 0;
        i_10_337 <= 0;
        i_10_338 <= 0;
        i_10_339 <= 0;
        i_10_340 <= 0;
        i_10_341 <= 0;
        i_10_342 <= 0;
        i_10_343 <= 0;
        i_10_344 <= 0;
        i_10_345 <= 0;
        i_10_346 <= 0;
        i_10_347 <= 0;
        i_10_348 <= 0;
        i_10_349 <= 0;
        i_10_350 <= 0;
        i_10_351 <= 0;
        i_10_352 <= 0;
        i_10_353 <= 0;
        i_10_354 <= 0;
        i_10_355 <= 0;
        i_10_356 <= 0;
        i_10_357 <= 0;
        i_10_358 <= 0;
        i_10_359 <= 0;
        i_10_360 <= 0;
        i_10_361 <= 0;
        i_10_362 <= 0;
        i_10_363 <= 0;
        i_10_364 <= 0;
        i_10_365 <= 0;
        i_10_366 <= 0;
        i_10_367 <= 0;
        i_10_368 <= 0;
        i_10_369 <= 0;
        i_10_370 <= 0;
        i_10_371 <= 0;
        i_10_372 <= 0;
        i_10_373 <= 0;
        i_10_374 <= 0;
        i_10_375 <= 0;
        i_10_376 <= 0;
        i_10_377 <= 0;
        i_10_378 <= 0;
        i_10_379 <= 0;
        i_10_380 <= 0;
        i_10_381 <= 0;
        i_10_382 <= 0;
        i_10_383 <= 0;
        i_10_384 <= 0;
        i_10_385 <= 0;
        i_10_386 <= 0;
        i_10_387 <= 0;
        i_10_388 <= 0;
        i_10_389 <= 0;
        i_10_390 <= 0;
        i_10_391 <= 0;
        i_10_392 <= 0;
        i_10_393 <= 0;
        i_10_394 <= 0;
        i_10_395 <= 0;
        i_10_396 <= 0;
        i_10_397 <= 0;
        i_10_398 <= 0;
        i_10_399 <= 0;
        i_10_400 <= 0;
        i_10_401 <= 0;
        i_10_402 <= 0;
        i_10_403 <= 0;
        i_10_404 <= 0;
        i_10_405 <= 0;
        i_10_406 <= 0;
        i_10_407 <= 0;
        i_10_408 <= 0;
        i_10_409 <= 0;
        i_10_410 <= 0;
        i_10_411 <= 0;
        i_10_412 <= 0;
        i_10_413 <= 0;
        i_10_414 <= 0;
        i_10_415 <= 0;
        i_10_416 <= 0;
        i_10_417 <= 0;
        i_10_418 <= 0;
        i_10_419 <= 0;
        i_10_420 <= 0;
        i_10_421 <= 0;
        i_10_422 <= 0;
        i_10_423 <= 0;
        i_10_424 <= 0;
        i_10_425 <= 0;
        i_10_426 <= 0;
        i_10_427 <= 0;
        i_10_428 <= 0;
        i_10_429 <= 0;
        i_10_430 <= 0;
        i_10_431 <= 0;
        i_10_432 <= 0;
        i_10_433 <= 0;
        i_10_434 <= 0;
        i_10_435 <= 0;
        i_10_436 <= 0;
        i_10_437 <= 0;
        i_10_438 <= 0;
        i_10_439 <= 0;
        i_10_440 <= 0;
        i_10_441 <= 0;
        i_10_442 <= 0;
        i_10_443 <= 0;
        i_10_444 <= 0;
        i_10_445 <= 0;
        i_10_446 <= 0;
        i_10_447 <= 0;
        i_10_448 <= 0;
        i_10_449 <= 0;
        i_10_450 <= 0;
        i_10_451 <= 0;
        i_10_452 <= 0;
        i_10_453 <= 0;
        i_10_454 <= 0;
        i_10_455 <= 0;
        i_10_456 <= 0;
        i_10_457 <= 0;
        i_10_458 <= 0;
        i_10_459 <= 0;
        i_10_460 <= 0;
        i_10_461 <= 0;
        i_10_462 <= 0;
        i_10_463 <= 0;
        i_10_464 <= 0;
        i_10_465 <= 0;
        i_10_466 <= 0;
        i_10_467 <= 0;
        i_10_468 <= 0;
        i_10_469 <= 0;
        i_10_470 <= 0;
        i_10_471 <= 0;
        i_10_472 <= 0;
        i_10_473 <= 0;
        i_10_474 <= 0;
        i_10_475 <= 0;
        i_10_476 <= 0;
        i_10_477 <= 0;
        i_10_478 <= 0;
        i_10_479 <= 0;
        i_10_480 <= 0;
        i_10_481 <= 0;
        i_10_482 <= 0;
        i_10_483 <= 0;
        i_10_484 <= 0;
        i_10_485 <= 0;
        i_10_486 <= 0;
        i_10_487 <= 0;
        i_10_488 <= 0;
        i_10_489 <= 0;
        i_10_490 <= 0;
        i_10_491 <= 0;
        i_10_492 <= 0;
        i_10_493 <= 0;
        i_10_494 <= 0;
        i_10_495 <= 0;
        i_10_496 <= 0;
        i_10_497 <= 0;
        i_10_498 <= 0;
        i_10_499 <= 0;
        i_10_500 <= 0;
        i_10_501 <= 0;
        i_10_502 <= 0;
        i_10_503 <= 0;
        i_10_504 <= 0;
        i_10_505 <= 0;
        i_10_506 <= 0;
        i_10_507 <= 0;
        i_10_508 <= 0;
        i_10_509 <= 0;
        i_10_510 <= 0;
        i_10_511 <= 0;
        i_10_512 <= 0;
        i_10_513 <= 0;
        i_10_514 <= 0;
        i_10_515 <= 0;
        i_10_516 <= 0;
        i_10_517 <= 0;
        i_10_518 <= 0;
        i_10_519 <= 0;
        i_10_520 <= 0;
        i_10_521 <= 0;
        i_10_522 <= 0;
        i_10_523 <= 0;
        i_10_524 <= 0;
        i_10_525 <= 0;
        i_10_526 <= 0;
        i_10_527 <= 0;
        i_10_528 <= 0;
        i_10_529 <= 0;
        i_10_530 <= 0;
        i_10_531 <= 0;
        i_10_532 <= 0;
        i_10_533 <= 0;
        i_10_534 <= 0;
        i_10_535 <= 0;
        i_10_536 <= 0;
        i_10_537 <= 0;
        i_10_538 <= 0;
        i_10_539 <= 0;
        i_10_540 <= 0;
        i_10_541 <= 0;
        i_10_542 <= 0;
        i_10_543 <= 0;
        i_10_544 <= 0;
        i_10_545 <= 0;
        i_10_546 <= 0;
        i_10_547 <= 0;
        i_10_548 <= 0;
        i_10_549 <= 0;
        i_10_550 <= 0;
        i_10_551 <= 0;
        i_10_552 <= 0;
        i_10_553 <= 0;
        i_10_554 <= 0;
        i_10_555 <= 0;
        i_10_556 <= 0;
        i_10_557 <= 0;
        i_10_558 <= 0;
        i_10_559 <= 0;
        i_10_560 <= 0;
        i_10_561 <= 0;
        i_10_562 <= 0;
        i_10_563 <= 0;
        i_10_564 <= 0;
        i_10_565 <= 0;
        i_10_566 <= 0;
        i_10_567 <= 0;
        i_10_568 <= 0;
        i_10_569 <= 0;
        i_10_570 <= 0;
        i_10_571 <= 0;
        i_10_572 <= 0;
        i_10_573 <= 0;
        i_10_574 <= 0;
        i_10_575 <= 0;
        i_10_576 <= 0;
        i_10_577 <= 0;
        i_10_578 <= 0;
        i_10_579 <= 0;
        i_10_580 <= 0;
        i_10_581 <= 0;
        i_10_582 <= 0;
        i_10_583 <= 0;
        i_10_584 <= 0;
        i_10_585 <= 0;
        i_10_586 <= 0;
        i_10_587 <= 0;
        i_10_588 <= 0;
        i_10_589 <= 0;
        i_10_590 <= 0;
        i_10_591 <= 0;
        i_10_592 <= 0;
        i_10_593 <= 0;
        i_10_594 <= 0;
        i_10_595 <= 0;
        i_10_596 <= 0;
        i_10_597 <= 0;
        i_10_598 <= 0;
        i_10_599 <= 0;
        i_10_600 <= 0;
        i_10_601 <= 0;
        i_10_602 <= 0;
        i_10_603 <= 0;
        i_10_604 <= 0;
        i_10_605 <= 0;
        i_10_606 <= 0;
        i_10_607 <= 0;
        i_10_608 <= 0;
        i_10_609 <= 0;
        i_10_610 <= 0;
        i_10_611 <= 0;
        i_10_612 <= 0;
        i_10_613 <= 0;
        i_10_614 <= 0;
        i_10_615 <= 0;
        i_10_616 <= 0;
        i_10_617 <= 0;
        i_10_618 <= 0;
        i_10_619 <= 0;
        i_10_620 <= 0;
        i_10_621 <= 0;
        i_10_622 <= 0;
        i_10_623 <= 0;
        i_10_624 <= 0;
        i_10_625 <= 0;
        i_10_626 <= 0;
        i_10_627 <= 0;
        i_10_628 <= 0;
        i_10_629 <= 0;
        i_10_630 <= 0;
        i_10_631 <= 0;
        i_10_632 <= 0;
        i_10_633 <= 0;
        i_10_634 <= 0;
        i_10_635 <= 0;
        i_10_636 <= 0;
        i_10_637 <= 0;
        i_10_638 <= 0;
        i_10_639 <= 0;
        i_10_640 <= 0;
        i_10_641 <= 0;
        i_10_642 <= 0;
        i_10_643 <= 0;
        i_10_644 <= 0;
        i_10_645 <= 0;
        i_10_646 <= 0;
        i_10_647 <= 0;
        i_10_648 <= 0;
        i_10_649 <= 0;
        i_10_650 <= 0;
        i_10_651 <= 0;
        i_10_652 <= 0;
        i_10_653 <= 0;
        i_10_654 <= 0;
        i_10_655 <= 0;
        i_10_656 <= 0;
        i_10_657 <= 0;
        i_10_658 <= 0;
        i_10_659 <= 0;
        i_10_660 <= 0;
        i_10_661 <= 0;
        i_10_662 <= 0;
        i_10_663 <= 0;
        i_10_664 <= 0;
        i_10_665 <= 0;
        i_10_666 <= 0;
        i_10_667 <= 0;
        i_10_668 <= 0;
        i_10_669 <= 0;
        i_10_670 <= 0;
        i_10_671 <= 0;
        i_10_672 <= 0;
        i_10_673 <= 0;
        i_10_674 <= 0;
        i_10_675 <= 0;
        i_10_676 <= 0;
        i_10_677 <= 0;
        i_10_678 <= 0;
        i_10_679 <= 0;
        i_10_680 <= 0;
        i_10_681 <= 0;
        i_10_682 <= 0;
        i_10_683 <= 0;
        i_10_684 <= 0;
        i_10_685 <= 0;
        i_10_686 <= 0;
        i_10_687 <= 0;
        i_10_688 <= 0;
        i_10_689 <= 0;
        i_10_690 <= 0;
        i_10_691 <= 0;
        i_10_692 <= 0;
        i_10_693 <= 0;
        i_10_694 <= 0;
        i_10_695 <= 0;
        i_10_696 <= 0;
        i_10_697 <= 0;
        i_10_698 <= 0;
        i_10_699 <= 0;
        i_10_700 <= 0;
        i_10_701 <= 0;
        i_10_702 <= 0;
        i_10_703 <= 0;
        i_10_704 <= 0;
        i_10_705 <= 0;
        i_10_706 <= 0;
        i_10_707 <= 0;
        i_10_708 <= 0;
        i_10_709 <= 0;
        i_10_710 <= 0;
        i_10_711 <= 0;
        i_10_712 <= 0;
        i_10_713 <= 0;
        i_10_714 <= 0;
        i_10_715 <= 0;
        i_10_716 <= 0;
        i_10_717 <= 0;
        i_10_718 <= 0;
        i_10_719 <= 0;
        i_10_720 <= 0;
        i_10_721 <= 0;
        i_10_722 <= 0;
        i_10_723 <= 0;
        i_10_724 <= 0;
        i_10_725 <= 0;
        i_10_726 <= 0;
        i_10_727 <= 0;
        i_10_728 <= 0;
        i_10_729 <= 0;
        i_10_730 <= 0;
        i_10_731 <= 0;
        i_10_732 <= 0;
        i_10_733 <= 0;
        i_10_734 <= 0;
        i_10_735 <= 0;
        i_10_736 <= 0;
        i_10_737 <= 0;
        i_10_738 <= 0;
        i_10_739 <= 0;
        i_10_740 <= 0;
        i_10_741 <= 0;
        i_10_742 <= 0;
        i_10_743 <= 0;
        i_10_744 <= 0;
        i_10_745 <= 0;
        i_10_746 <= 0;
        i_10_747 <= 0;
        i_10_748 <= 0;
        i_10_749 <= 0;
        i_10_750 <= 0;
        i_10_751 <= 0;
        i_10_752 <= 0;
        i_10_753 <= 0;
        i_10_754 <= 0;
        i_10_755 <= 0;
        i_10_756 <= 0;
        i_10_757 <= 0;
        i_10_758 <= 0;
        i_10_759 <= 0;
        i_10_760 <= 0;
        i_10_761 <= 0;
        i_10_762 <= 0;
        i_10_763 <= 0;
        i_10_764 <= 0;
        i_10_765 <= 0;
        i_10_766 <= 0;
        i_10_767 <= 0;
        i_10_768 <= 0;
        i_10_769 <= 0;
        i_10_770 <= 0;
        i_10_771 <= 0;
        i_10_772 <= 0;
        i_10_773 <= 0;
        i_10_774 <= 0;
        i_10_775 <= 0;
        i_10_776 <= 0;
        i_10_777 <= 0;
        i_10_778 <= 0;
        i_10_779 <= 0;
        i_10_780 <= 0;
        i_10_781 <= 0;
        i_10_782 <= 0;
        i_10_783 <= 0;
        i_10_784 <= 0;
        i_10_785 <= 0;
        i_10_786 <= 0;
        i_10_787 <= 0;
        i_10_788 <= 0;
        i_10_789 <= 0;
        i_10_790 <= 0;
        i_10_791 <= 0;
        i_10_792 <= 0;
        i_10_793 <= 0;
        i_10_794 <= 0;
        i_10_795 <= 0;
        i_10_796 <= 0;
        i_10_797 <= 0;
        i_10_798 <= 0;
        i_10_799 <= 0;
        i_10_800 <= 0;
        i_10_801 <= 0;
        i_10_802 <= 0;
        i_10_803 <= 0;
        i_10_804 <= 0;
        i_10_805 <= 0;
        i_10_806 <= 0;
        i_10_807 <= 0;
        i_10_808 <= 0;
        i_10_809 <= 0;
        i_10_810 <= 0;
        i_10_811 <= 0;
        i_10_812 <= 0;
        i_10_813 <= 0;
        i_10_814 <= 0;
        i_10_815 <= 0;
        i_10_816 <= 0;
        i_10_817 <= 0;
        i_10_818 <= 0;
        i_10_819 <= 0;
        i_10_820 <= 0;
        i_10_821 <= 0;
        i_10_822 <= 0;
        i_10_823 <= 0;
        i_10_824 <= 0;
        i_10_825 <= 0;
        i_10_826 <= 0;
        i_10_827 <= 0;
        i_10_828 <= 0;
        i_10_829 <= 0;
        i_10_830 <= 0;
        i_10_831 <= 0;
        i_10_832 <= 0;
        i_10_833 <= 0;
        i_10_834 <= 0;
        i_10_835 <= 0;
        i_10_836 <= 0;
        i_10_837 <= 0;
        i_10_838 <= 0;
        i_10_839 <= 0;
        i_10_840 <= 0;
        i_10_841 <= 0;
        i_10_842 <= 0;
        i_10_843 <= 0;
        i_10_844 <= 0;
        i_10_845 <= 0;
        i_10_846 <= 0;
        i_10_847 <= 0;
        i_10_848 <= 0;
        i_10_849 <= 0;
        i_10_850 <= 0;
        i_10_851 <= 0;
        i_10_852 <= 0;
        i_10_853 <= 0;
        i_10_854 <= 0;
        i_10_855 <= 0;
        i_10_856 <= 0;
        i_10_857 <= 0;
        i_10_858 <= 0;
        i_10_859 <= 0;
        i_10_860 <= 0;
        i_10_861 <= 0;
        i_10_862 <= 0;
        i_10_863 <= 0;
        i_10_864 <= 0;
        i_10_865 <= 0;
        i_10_866 <= 0;
        i_10_867 <= 0;
        i_10_868 <= 0;
        i_10_869 <= 0;
        i_10_870 <= 0;
        i_10_871 <= 0;
        i_10_872 <= 0;
        i_10_873 <= 0;
        i_10_874 <= 0;
        i_10_875 <= 0;
        i_10_876 <= 0;
        i_10_877 <= 0;
        i_10_878 <= 0;
        i_10_879 <= 0;
        i_10_880 <= 0;
        i_10_881 <= 0;
        i_10_882 <= 0;
        i_10_883 <= 0;
        i_10_884 <= 0;
        i_10_885 <= 0;
        i_10_886 <= 0;
        i_10_887 <= 0;
        i_10_888 <= 0;
        i_10_889 <= 0;
        i_10_890 <= 0;
        i_10_891 <= 0;
        i_10_892 <= 0;
        i_10_893 <= 0;
        i_10_894 <= 0;
        i_10_895 <= 0;
        i_10_896 <= 0;
        i_10_897 <= 0;
        i_10_898 <= 0;
        i_10_899 <= 0;
        i_10_900 <= 0;
        i_10_901 <= 0;
        i_10_902 <= 0;
        i_10_903 <= 0;
        i_10_904 <= 0;
        i_10_905 <= 0;
        i_10_906 <= 0;
        i_10_907 <= 0;
        i_10_908 <= 0;
        i_10_909 <= 0;
        i_10_910 <= 0;
        i_10_911 <= 0;
        i_10_912 <= 0;
        i_10_913 <= 0;
        i_10_914 <= 0;
        i_10_915 <= 0;
        i_10_916 <= 0;
        i_10_917 <= 0;
        i_10_918 <= 0;
        i_10_919 <= 0;
        i_10_920 <= 0;
        i_10_921 <= 0;
        i_10_922 <= 0;
        i_10_923 <= 0;
        i_10_924 <= 0;
        i_10_925 <= 0;
        i_10_926 <= 0;
        i_10_927 <= 0;
        i_10_928 <= 0;
        i_10_929 <= 0;
        i_10_930 <= 0;
        i_10_931 <= 0;
        i_10_932 <= 0;
        i_10_933 <= 0;
        i_10_934 <= 0;
        i_10_935 <= 0;
        i_10_936 <= 0;
        i_10_937 <= 0;
        i_10_938 <= 0;
        i_10_939 <= 0;
        i_10_940 <= 0;
        i_10_941 <= 0;
        i_10_942 <= 0;
        i_10_943 <= 0;
        i_10_944 <= 0;
        i_10_945 <= 0;
        i_10_946 <= 0;
        i_10_947 <= 0;
        i_10_948 <= 0;
        i_10_949 <= 0;
        i_10_950 <= 0;
        i_10_951 <= 0;
        i_10_952 <= 0;
        i_10_953 <= 0;
        i_10_954 <= 0;
        i_10_955 <= 0;
        i_10_956 <= 0;
        i_10_957 <= 0;
        i_10_958 <= 0;
        i_10_959 <= 0;
        i_10_960 <= 0;
        i_10_961 <= 0;
        i_10_962 <= 0;
        i_10_963 <= 0;
        i_10_964 <= 0;
        i_10_965 <= 0;
        i_10_966 <= 0;
        i_10_967 <= 0;
        i_10_968 <= 0;
        i_10_969 <= 0;
        i_10_970 <= 0;
        i_10_971 <= 0;
        i_10_972 <= 0;
        i_10_973 <= 0;
        i_10_974 <= 0;
        i_10_975 <= 0;
        i_10_976 <= 0;
        i_10_977 <= 0;
        i_10_978 <= 0;
        i_10_979 <= 0;
        i_10_980 <= 0;
        i_10_981 <= 0;
        i_10_982 <= 0;
        i_10_983 <= 0;
        i_10_984 <= 0;
        i_10_985 <= 0;
        i_10_986 <= 0;
        i_10_987 <= 0;
        i_10_988 <= 0;
        i_10_989 <= 0;
        i_10_990 <= 0;
        i_10_991 <= 0;
        i_10_992 <= 0;
        i_10_993 <= 0;
        i_10_994 <= 0;
        i_10_995 <= 0;
        i_10_996 <= 0;
        i_10_997 <= 0;
        i_10_998 <= 0;
        i_10_999 <= 0;
        i_10_1000 <= 0;
        i_10_1001 <= 0;
        i_10_1002 <= 0;
        i_10_1003 <= 0;
        i_10_1004 <= 0;
        i_10_1005 <= 0;
        i_10_1006 <= 0;
        i_10_1007 <= 0;
        i_10_1008 <= 0;
        i_10_1009 <= 0;
        i_10_1010 <= 0;
        i_10_1011 <= 0;
        i_10_1012 <= 0;
        i_10_1013 <= 0;
        i_10_1014 <= 0;
        i_10_1015 <= 0;
        i_10_1016 <= 0;
        i_10_1017 <= 0;
        i_10_1018 <= 0;
        i_10_1019 <= 0;
        i_10_1020 <= 0;
        i_10_1021 <= 0;
        i_10_1022 <= 0;
        i_10_1023 <= 0;
        i_10_1024 <= 0;
        i_10_1025 <= 0;
        i_10_1026 <= 0;
        i_10_1027 <= 0;
        i_10_1028 <= 0;
        i_10_1029 <= 0;
        i_10_1030 <= 0;
        i_10_1031 <= 0;
        i_10_1032 <= 0;
        i_10_1033 <= 0;
        i_10_1034 <= 0;
        i_10_1035 <= 0;
        i_10_1036 <= 0;
        i_10_1037 <= 0;
        i_10_1038 <= 0;
        i_10_1039 <= 0;
        i_10_1040 <= 0;
        i_10_1041 <= 0;
        i_10_1042 <= 0;
        i_10_1043 <= 0;
        i_10_1044 <= 0;
        i_10_1045 <= 0;
        i_10_1046 <= 0;
        i_10_1047 <= 0;
        i_10_1048 <= 0;
        i_10_1049 <= 0;
        i_10_1050 <= 0;
        i_10_1051 <= 0;
        i_10_1052 <= 0;
        i_10_1053 <= 0;
        i_10_1054 <= 0;
        i_10_1055 <= 0;
        i_10_1056 <= 0;
        i_10_1057 <= 0;
        i_10_1058 <= 0;
        i_10_1059 <= 0;
        i_10_1060 <= 0;
        i_10_1061 <= 0;
        i_10_1062 <= 0;
        i_10_1063 <= 0;
        i_10_1064 <= 0;
        i_10_1065 <= 0;
        i_10_1066 <= 0;
        i_10_1067 <= 0;
        i_10_1068 <= 0;
        i_10_1069 <= 0;
        i_10_1070 <= 0;
        i_10_1071 <= 0;
        i_10_1072 <= 0;
        i_10_1073 <= 0;
        i_10_1074 <= 0;
        i_10_1075 <= 0;
        i_10_1076 <= 0;
        i_10_1077 <= 0;
        i_10_1078 <= 0;
        i_10_1079 <= 0;
        i_10_1080 <= 0;
        i_10_1081 <= 0;
        i_10_1082 <= 0;
        i_10_1083 <= 0;
        i_10_1084 <= 0;
        i_10_1085 <= 0;
        i_10_1086 <= 0;
        i_10_1087 <= 0;
        i_10_1088 <= 0;
        i_10_1089 <= 0;
        i_10_1090 <= 0;
        i_10_1091 <= 0;
        i_10_1092 <= 0;
        i_10_1093 <= 0;
        i_10_1094 <= 0;
        i_10_1095 <= 0;
        i_10_1096 <= 0;
        i_10_1097 <= 0;
        i_10_1098 <= 0;
        i_10_1099 <= 0;
        i_10_1100 <= 0;
        i_10_1101 <= 0;
        i_10_1102 <= 0;
        i_10_1103 <= 0;
        i_10_1104 <= 0;
        i_10_1105 <= 0;
        i_10_1106 <= 0;
        i_10_1107 <= 0;
        i_10_1108 <= 0;
        i_10_1109 <= 0;
        i_10_1110 <= 0;
        i_10_1111 <= 0;
        i_10_1112 <= 0;
        i_10_1113 <= 0;
        i_10_1114 <= 0;
        i_10_1115 <= 0;
        i_10_1116 <= 0;
        i_10_1117 <= 0;
        i_10_1118 <= 0;
        i_10_1119 <= 0;
        i_10_1120 <= 0;
        i_10_1121 <= 0;
        i_10_1122 <= 0;
        i_10_1123 <= 0;
        i_10_1124 <= 0;
        i_10_1125 <= 0;
        i_10_1126 <= 0;
        i_10_1127 <= 0;
        i_10_1128 <= 0;
        i_10_1129 <= 0;
        i_10_1130 <= 0;
        i_10_1131 <= 0;
        i_10_1132 <= 0;
        i_10_1133 <= 0;
        i_10_1134 <= 0;
        i_10_1135 <= 0;
        i_10_1136 <= 0;
        i_10_1137 <= 0;
        i_10_1138 <= 0;
        i_10_1139 <= 0;
        i_10_1140 <= 0;
        i_10_1141 <= 0;
        i_10_1142 <= 0;
        i_10_1143 <= 0;
        i_10_1144 <= 0;
        i_10_1145 <= 0;
        i_10_1146 <= 0;
        i_10_1147 <= 0;
        i_10_1148 <= 0;
        i_10_1149 <= 0;
        i_10_1150 <= 0;
        i_10_1151 <= 0;
        i_10_1152 <= 0;
        i_10_1153 <= 0;
        i_10_1154 <= 0;
        i_10_1155 <= 0;
        i_10_1156 <= 0;
        i_10_1157 <= 0;
        i_10_1158 <= 0;
        i_10_1159 <= 0;
        i_10_1160 <= 0;
        i_10_1161 <= 0;
        i_10_1162 <= 0;
        i_10_1163 <= 0;
        i_10_1164 <= 0;
        i_10_1165 <= 0;
        i_10_1166 <= 0;
        i_10_1167 <= 0;
        i_10_1168 <= 0;
        i_10_1169 <= 0;
        i_10_1170 <= 0;
        i_10_1171 <= 0;
        i_10_1172 <= 0;
        i_10_1173 <= 0;
        i_10_1174 <= 0;
        i_10_1175 <= 0;
        i_10_1176 <= 0;
        i_10_1177 <= 0;
        i_10_1178 <= 0;
        i_10_1179 <= 0;
        i_10_1180 <= 0;
        i_10_1181 <= 0;
        i_10_1182 <= 0;
        i_10_1183 <= 0;
        i_10_1184 <= 0;
        i_10_1185 <= 0;
        i_10_1186 <= 0;
        i_10_1187 <= 0;
        i_10_1188 <= 0;
        i_10_1189 <= 0;
        i_10_1190 <= 0;
        i_10_1191 <= 0;
        i_10_1192 <= 0;
        i_10_1193 <= 0;
        i_10_1194 <= 0;
        i_10_1195 <= 0;
        i_10_1196 <= 0;
        i_10_1197 <= 0;
        i_10_1198 <= 0;
        i_10_1199 <= 0;
        i_10_1200 <= 0;
        i_10_1201 <= 0;
        i_10_1202 <= 0;
        i_10_1203 <= 0;
        i_10_1204 <= 0;
        i_10_1205 <= 0;
        i_10_1206 <= 0;
        i_10_1207 <= 0;
        i_10_1208 <= 0;
        i_10_1209 <= 0;
        i_10_1210 <= 0;
        i_10_1211 <= 0;
        i_10_1212 <= 0;
        i_10_1213 <= 0;
        i_10_1214 <= 0;
        i_10_1215 <= 0;
        i_10_1216 <= 0;
        i_10_1217 <= 0;
        i_10_1218 <= 0;
        i_10_1219 <= 0;
        i_10_1220 <= 0;
        i_10_1221 <= 0;
        i_10_1222 <= 0;
        i_10_1223 <= 0;
        i_10_1224 <= 0;
        i_10_1225 <= 0;
        i_10_1226 <= 0;
        i_10_1227 <= 0;
        i_10_1228 <= 0;
        i_10_1229 <= 0;
        i_10_1230 <= 0;
        i_10_1231 <= 0;
        i_10_1232 <= 0;
        i_10_1233 <= 0;
        i_10_1234 <= 0;
        i_10_1235 <= 0;
        i_10_1236 <= 0;
        i_10_1237 <= 0;
        i_10_1238 <= 0;
        i_10_1239 <= 0;
        i_10_1240 <= 0;
        i_10_1241 <= 0;
        i_10_1242 <= 0;
        i_10_1243 <= 0;
        i_10_1244 <= 0;
        i_10_1245 <= 0;
        i_10_1246 <= 0;
        i_10_1247 <= 0;
        i_10_1248 <= 0;
        i_10_1249 <= 0;
        i_10_1250 <= 0;
        i_10_1251 <= 0;
        i_10_1252 <= 0;
        i_10_1253 <= 0;
        i_10_1254 <= 0;
        i_10_1255 <= 0;
        i_10_1256 <= 0;
        i_10_1257 <= 0;
        i_10_1258 <= 0;
        i_10_1259 <= 0;
        i_10_1260 <= 0;
        i_10_1261 <= 0;
        i_10_1262 <= 0;
        i_10_1263 <= 0;
        i_10_1264 <= 0;
        i_10_1265 <= 0;
        i_10_1266 <= 0;
        i_10_1267 <= 0;
        i_10_1268 <= 0;
        i_10_1269 <= 0;
        i_10_1270 <= 0;
        i_10_1271 <= 0;
        i_10_1272 <= 0;
        i_10_1273 <= 0;
        i_10_1274 <= 0;
        i_10_1275 <= 0;
        i_10_1276 <= 0;
        i_10_1277 <= 0;
        i_10_1278 <= 0;
        i_10_1279 <= 0;
        i_10_1280 <= 0;
        i_10_1281 <= 0;
        i_10_1282 <= 0;
        i_10_1283 <= 0;
        i_10_1284 <= 0;
        i_10_1285 <= 0;
        i_10_1286 <= 0;
        i_10_1287 <= 0;
        i_10_1288 <= 0;
        i_10_1289 <= 0;
        i_10_1290 <= 0;
        i_10_1291 <= 0;
        i_10_1292 <= 0;
        i_10_1293 <= 0;
        i_10_1294 <= 0;
        i_10_1295 <= 0;
        i_10_1296 <= 0;
        i_10_1297 <= 0;
        i_10_1298 <= 0;
        i_10_1299 <= 0;
        i_10_1300 <= 0;
        i_10_1301 <= 0;
        i_10_1302 <= 0;
        i_10_1303 <= 0;
        i_10_1304 <= 0;
        i_10_1305 <= 0;
        i_10_1306 <= 0;
        i_10_1307 <= 0;
        i_10_1308 <= 0;
        i_10_1309 <= 0;
        i_10_1310 <= 0;
        i_10_1311 <= 0;
        i_10_1312 <= 0;
        i_10_1313 <= 0;
        i_10_1314 <= 0;
        i_10_1315 <= 0;
        i_10_1316 <= 0;
        i_10_1317 <= 0;
        i_10_1318 <= 0;
        i_10_1319 <= 0;
        i_10_1320 <= 0;
        i_10_1321 <= 0;
        i_10_1322 <= 0;
        i_10_1323 <= 0;
        i_10_1324 <= 0;
        i_10_1325 <= 0;
        i_10_1326 <= 0;
        i_10_1327 <= 0;
        i_10_1328 <= 0;
        i_10_1329 <= 0;
        i_10_1330 <= 0;
        i_10_1331 <= 0;
        i_10_1332 <= 0;
        i_10_1333 <= 0;
        i_10_1334 <= 0;
        i_10_1335 <= 0;
        i_10_1336 <= 0;
        i_10_1337 <= 0;
        i_10_1338 <= 0;
        i_10_1339 <= 0;
        i_10_1340 <= 0;
        i_10_1341 <= 0;
        i_10_1342 <= 0;
        i_10_1343 <= 0;
        i_10_1344 <= 0;
        i_10_1345 <= 0;
        i_10_1346 <= 0;
        i_10_1347 <= 0;
        i_10_1348 <= 0;
        i_10_1349 <= 0;
        i_10_1350 <= 0;
        i_10_1351 <= 0;
        i_10_1352 <= 0;
        i_10_1353 <= 0;
        i_10_1354 <= 0;
        i_10_1355 <= 0;
        i_10_1356 <= 0;
        i_10_1357 <= 0;
        i_10_1358 <= 0;
        i_10_1359 <= 0;
        i_10_1360 <= 0;
        i_10_1361 <= 0;
        i_10_1362 <= 0;
        i_10_1363 <= 0;
        i_10_1364 <= 0;
        i_10_1365 <= 0;
        i_10_1366 <= 0;
        i_10_1367 <= 0;
        i_10_1368 <= 0;
        i_10_1369 <= 0;
        i_10_1370 <= 0;
        i_10_1371 <= 0;
        i_10_1372 <= 0;
        i_10_1373 <= 0;
        i_10_1374 <= 0;
        i_10_1375 <= 0;
        i_10_1376 <= 0;
        i_10_1377 <= 0;
        i_10_1378 <= 0;
        i_10_1379 <= 0;
        i_10_1380 <= 0;
        i_10_1381 <= 0;
        i_10_1382 <= 0;
        i_10_1383 <= 0;
        i_10_1384 <= 0;
        i_10_1385 <= 0;
        i_10_1386 <= 0;
        i_10_1387 <= 0;
        i_10_1388 <= 0;
        i_10_1389 <= 0;
        i_10_1390 <= 0;
        i_10_1391 <= 0;
        i_10_1392 <= 0;
        i_10_1393 <= 0;
        i_10_1394 <= 0;
        i_10_1395 <= 0;
        i_10_1396 <= 0;
        i_10_1397 <= 0;
        i_10_1398 <= 0;
        i_10_1399 <= 0;
        i_10_1400 <= 0;
        i_10_1401 <= 0;
        i_10_1402 <= 0;
        i_10_1403 <= 0;
        i_10_1404 <= 0;
        i_10_1405 <= 0;
        i_10_1406 <= 0;
        i_10_1407 <= 0;
        i_10_1408 <= 0;
        i_10_1409 <= 0;
        i_10_1410 <= 0;
        i_10_1411 <= 0;
        i_10_1412 <= 0;
        i_10_1413 <= 0;
        i_10_1414 <= 0;
        i_10_1415 <= 0;
        i_10_1416 <= 0;
        i_10_1417 <= 0;
        i_10_1418 <= 0;
        i_10_1419 <= 0;
        i_10_1420 <= 0;
        i_10_1421 <= 0;
        i_10_1422 <= 0;
        i_10_1423 <= 0;
        i_10_1424 <= 0;
        i_10_1425 <= 0;
        i_10_1426 <= 0;
        i_10_1427 <= 0;
        i_10_1428 <= 0;
        i_10_1429 <= 0;
        i_10_1430 <= 0;
        i_10_1431 <= 0;
        i_10_1432 <= 0;
        i_10_1433 <= 0;
        i_10_1434 <= 0;
        i_10_1435 <= 0;
        i_10_1436 <= 0;
        i_10_1437 <= 0;
        i_10_1438 <= 0;
        i_10_1439 <= 0;
        i_10_1440 <= 0;
        i_10_1441 <= 0;
        i_10_1442 <= 0;
        i_10_1443 <= 0;
        i_10_1444 <= 0;
        i_10_1445 <= 0;
        i_10_1446 <= 0;
        i_10_1447 <= 0;
        i_10_1448 <= 0;
        i_10_1449 <= 0;
        i_10_1450 <= 0;
        i_10_1451 <= 0;
        i_10_1452 <= 0;
        i_10_1453 <= 0;
        i_10_1454 <= 0;
        i_10_1455 <= 0;
        i_10_1456 <= 0;
        i_10_1457 <= 0;
        i_10_1458 <= 0;
        i_10_1459 <= 0;
        i_10_1460 <= 0;
        i_10_1461 <= 0;
        i_10_1462 <= 0;
        i_10_1463 <= 0;
        i_10_1464 <= 0;
        i_10_1465 <= 0;
        i_10_1466 <= 0;
        i_10_1467 <= 0;
        i_10_1468 <= 0;
        i_10_1469 <= 0;
        i_10_1470 <= 0;
        i_10_1471 <= 0;
        i_10_1472 <= 0;
        i_10_1473 <= 0;
        i_10_1474 <= 0;
        i_10_1475 <= 0;
        i_10_1476 <= 0;
        i_10_1477 <= 0;
        i_10_1478 <= 0;
        i_10_1479 <= 0;
        i_10_1480 <= 0;
        i_10_1481 <= 0;
        i_10_1482 <= 0;
        i_10_1483 <= 0;
        i_10_1484 <= 0;
        i_10_1485 <= 0;
        i_10_1486 <= 0;
        i_10_1487 <= 0;
        i_10_1488 <= 0;
        i_10_1489 <= 0;
        i_10_1490 <= 0;
        i_10_1491 <= 0;
        i_10_1492 <= 0;
        i_10_1493 <= 0;
        i_10_1494 <= 0;
        i_10_1495 <= 0;
        i_10_1496 <= 0;
        i_10_1497 <= 0;
        i_10_1498 <= 0;
        i_10_1499 <= 0;
        i_10_1500 <= 0;
        i_10_1501 <= 0;
        i_10_1502 <= 0;
        i_10_1503 <= 0;
        i_10_1504 <= 0;
        i_10_1505 <= 0;
        i_10_1506 <= 0;
        i_10_1507 <= 0;
        i_10_1508 <= 0;
        i_10_1509 <= 0;
        i_10_1510 <= 0;
        i_10_1511 <= 0;
        i_10_1512 <= 0;
        i_10_1513 <= 0;
        i_10_1514 <= 0;
        i_10_1515 <= 0;
        i_10_1516 <= 0;
        i_10_1517 <= 0;
        i_10_1518 <= 0;
        i_10_1519 <= 0;
        i_10_1520 <= 0;
        i_10_1521 <= 0;
        i_10_1522 <= 0;
        i_10_1523 <= 0;
        i_10_1524 <= 0;
        i_10_1525 <= 0;
        i_10_1526 <= 0;
        i_10_1527 <= 0;
        i_10_1528 <= 0;
        i_10_1529 <= 0;
        i_10_1530 <= 0;
        i_10_1531 <= 0;
        i_10_1532 <= 0;
        i_10_1533 <= 0;
        i_10_1534 <= 0;
        i_10_1535 <= 0;
        i_10_1536 <= 0;
        i_10_1537 <= 0;
        i_10_1538 <= 0;
        i_10_1539 <= 0;
        i_10_1540 <= 0;
        i_10_1541 <= 0;
        i_10_1542 <= 0;
        i_10_1543 <= 0;
        i_10_1544 <= 0;
        i_10_1545 <= 0;
        i_10_1546 <= 0;
        i_10_1547 <= 0;
        i_10_1548 <= 0;
        i_10_1549 <= 0;
        i_10_1550 <= 0;
        i_10_1551 <= 0;
        i_10_1552 <= 0;
        i_10_1553 <= 0;
        i_10_1554 <= 0;
        i_10_1555 <= 0;
        i_10_1556 <= 0;
        i_10_1557 <= 0;
        i_10_1558 <= 0;
        i_10_1559 <= 0;
        i_10_1560 <= 0;
        i_10_1561 <= 0;
        i_10_1562 <= 0;
        i_10_1563 <= 0;
        i_10_1564 <= 0;
        i_10_1565 <= 0;
        i_10_1566 <= 0;
        i_10_1567 <= 0;
        i_10_1568 <= 0;
        i_10_1569 <= 0;
        i_10_1570 <= 0;
        i_10_1571 <= 0;
        i_10_1572 <= 0;
        i_10_1573 <= 0;
        i_10_1574 <= 0;
        i_10_1575 <= 0;
        i_10_1576 <= 0;
        i_10_1577 <= 0;
        i_10_1578 <= 0;
        i_10_1579 <= 0;
        i_10_1580 <= 0;
        i_10_1581 <= 0;
        i_10_1582 <= 0;
        i_10_1583 <= 0;
        i_10_1584 <= 0;
        i_10_1585 <= 0;
        i_10_1586 <= 0;
        i_10_1587 <= 0;
        i_10_1588 <= 0;
        i_10_1589 <= 0;
        i_10_1590 <= 0;
        i_10_1591 <= 0;
        i_10_1592 <= 0;
        i_10_1593 <= 0;
        i_10_1594 <= 0;
        i_10_1595 <= 0;
        i_10_1596 <= 0;
        i_10_1597 <= 0;
        i_10_1598 <= 0;
        i_10_1599 <= 0;
        i_10_1600 <= 0;
        i_10_1601 <= 0;
        i_10_1602 <= 0;
        i_10_1603 <= 0;
        i_10_1604 <= 0;
        i_10_1605 <= 0;
        i_10_1606 <= 0;
        i_10_1607 <= 0;
        i_10_1608 <= 0;
        i_10_1609 <= 0;
        i_10_1610 <= 0;
        i_10_1611 <= 0;
        i_10_1612 <= 0;
        i_10_1613 <= 0;
        i_10_1614 <= 0;
        i_10_1615 <= 0;
        i_10_1616 <= 0;
        i_10_1617 <= 0;
        i_10_1618 <= 0;
        i_10_1619 <= 0;
        i_10_1620 <= 0;
        i_10_1621 <= 0;
        i_10_1622 <= 0;
        i_10_1623 <= 0;
        i_10_1624 <= 0;
        i_10_1625 <= 0;
        i_10_1626 <= 0;
        i_10_1627 <= 0;
        i_10_1628 <= 0;
        i_10_1629 <= 0;
        i_10_1630 <= 0;
        i_10_1631 <= 0;
        i_10_1632 <= 0;
        i_10_1633 <= 0;
        i_10_1634 <= 0;
        i_10_1635 <= 0;
        i_10_1636 <= 0;
        i_10_1637 <= 0;
        i_10_1638 <= 0;
        i_10_1639 <= 0;
        i_10_1640 <= 0;
        i_10_1641 <= 0;
        i_10_1642 <= 0;
        i_10_1643 <= 0;
        i_10_1644 <= 0;
        i_10_1645 <= 0;
        i_10_1646 <= 0;
        i_10_1647 <= 0;
        i_10_1648 <= 0;
        i_10_1649 <= 0;
        i_10_1650 <= 0;
        i_10_1651 <= 0;
        i_10_1652 <= 0;
        i_10_1653 <= 0;
        i_10_1654 <= 0;
        i_10_1655 <= 0;
        i_10_1656 <= 0;
        i_10_1657 <= 0;
        i_10_1658 <= 0;
        i_10_1659 <= 0;
        i_10_1660 <= 0;
        i_10_1661 <= 0;
        i_10_1662 <= 0;
        i_10_1663 <= 0;
        i_10_1664 <= 0;
        i_10_1665 <= 0;
        i_10_1666 <= 0;
        i_10_1667 <= 0;
        i_10_1668 <= 0;
        i_10_1669 <= 0;
        i_10_1670 <= 0;
        i_10_1671 <= 0;
        i_10_1672 <= 0;
        i_10_1673 <= 0;
        i_10_1674 <= 0;
        i_10_1675 <= 0;
        i_10_1676 <= 0;
        i_10_1677 <= 0;
        i_10_1678 <= 0;
        i_10_1679 <= 0;
        i_10_1680 <= 0;
        i_10_1681 <= 0;
        i_10_1682 <= 0;
        i_10_1683 <= 0;
        i_10_1684 <= 0;
        i_10_1685 <= 0;
        i_10_1686 <= 0;
        i_10_1687 <= 0;
        i_10_1688 <= 0;
        i_10_1689 <= 0;
        i_10_1690 <= 0;
        i_10_1691 <= 0;
        i_10_1692 <= 0;
        i_10_1693 <= 0;
        i_10_1694 <= 0;
        i_10_1695 <= 0;
        i_10_1696 <= 0;
        i_10_1697 <= 0;
        i_10_1698 <= 0;
        i_10_1699 <= 0;
        i_10_1700 <= 0;
        i_10_1701 <= 0;
        i_10_1702 <= 0;
        i_10_1703 <= 0;
        i_10_1704 <= 0;
        i_10_1705 <= 0;
        i_10_1706 <= 0;
        i_10_1707 <= 0;
        i_10_1708 <= 0;
        i_10_1709 <= 0;
        i_10_1710 <= 0;
        i_10_1711 <= 0;
        i_10_1712 <= 0;
        i_10_1713 <= 0;
        i_10_1714 <= 0;
        i_10_1715 <= 0;
        i_10_1716 <= 0;
        i_10_1717 <= 0;
        i_10_1718 <= 0;
        i_10_1719 <= 0;
        i_10_1720 <= 0;
        i_10_1721 <= 0;
        i_10_1722 <= 0;
        i_10_1723 <= 0;
        i_10_1724 <= 0;
        i_10_1725 <= 0;
        i_10_1726 <= 0;
        i_10_1727 <= 0;
        i_10_1728 <= 0;
        i_10_1729 <= 0;
        i_10_1730 <= 0;
        i_10_1731 <= 0;
        i_10_1732 <= 0;
        i_10_1733 <= 0;
        i_10_1734 <= 0;
        i_10_1735 <= 0;
        i_10_1736 <= 0;
        i_10_1737 <= 0;
        i_10_1738 <= 0;
        i_10_1739 <= 0;
        i_10_1740 <= 0;
        i_10_1741 <= 0;
        i_10_1742 <= 0;
        i_10_1743 <= 0;
        i_10_1744 <= 0;
        i_10_1745 <= 0;
        i_10_1746 <= 0;
        i_10_1747 <= 0;
        i_10_1748 <= 0;
        i_10_1749 <= 0;
        i_10_1750 <= 0;
        i_10_1751 <= 0;
        i_10_1752 <= 0;
        i_10_1753 <= 0;
        i_10_1754 <= 0;
        i_10_1755 <= 0;
        i_10_1756 <= 0;
        i_10_1757 <= 0;
        i_10_1758 <= 0;
        i_10_1759 <= 0;
        i_10_1760 <= 0;
        i_10_1761 <= 0;
        i_10_1762 <= 0;
        i_10_1763 <= 0;
        i_10_1764 <= 0;
        i_10_1765 <= 0;
        i_10_1766 <= 0;
        i_10_1767 <= 0;
        i_10_1768 <= 0;
        i_10_1769 <= 0;
        i_10_1770 <= 0;
        i_10_1771 <= 0;
        i_10_1772 <= 0;
        i_10_1773 <= 0;
        i_10_1774 <= 0;
        i_10_1775 <= 0;
        i_10_1776 <= 0;
        i_10_1777 <= 0;
        i_10_1778 <= 0;
        i_10_1779 <= 0;
        i_10_1780 <= 0;
        i_10_1781 <= 0;
        i_10_1782 <= 0;
        i_10_1783 <= 0;
        i_10_1784 <= 0;
        i_10_1785 <= 0;
        i_10_1786 <= 0;
        i_10_1787 <= 0;
        i_10_1788 <= 0;
        i_10_1789 <= 0;
        i_10_1790 <= 0;
        i_10_1791 <= 0;
        i_10_1792 <= 0;
        i_10_1793 <= 0;
        i_10_1794 <= 0;
        i_10_1795 <= 0;
        i_10_1796 <= 0;
        i_10_1797 <= 0;
        i_10_1798 <= 0;
        i_10_1799 <= 0;
        i_10_1800 <= 0;
        i_10_1801 <= 0;
        i_10_1802 <= 0;
        i_10_1803 <= 0;
        i_10_1804 <= 0;
        i_10_1805 <= 0;
        i_10_1806 <= 0;
        i_10_1807 <= 0;
        i_10_1808 <= 0;
        i_10_1809 <= 0;
        i_10_1810 <= 0;
        i_10_1811 <= 0;
        i_10_1812 <= 0;
        i_10_1813 <= 0;
        i_10_1814 <= 0;
        i_10_1815 <= 0;
        i_10_1816 <= 0;
        i_10_1817 <= 0;
        i_10_1818 <= 0;
        i_10_1819 <= 0;
        i_10_1820 <= 0;
        i_10_1821 <= 0;
        i_10_1822 <= 0;
        i_10_1823 <= 0;
        i_10_1824 <= 0;
        i_10_1825 <= 0;
        i_10_1826 <= 0;
        i_10_1827 <= 0;
        i_10_1828 <= 0;
        i_10_1829 <= 0;
        i_10_1830 <= 0;
        i_10_1831 <= 0;
        i_10_1832 <= 0;
        i_10_1833 <= 0;
        i_10_1834 <= 0;
        i_10_1835 <= 0;
        i_10_1836 <= 0;
        i_10_1837 <= 0;
        i_10_1838 <= 0;
        i_10_1839 <= 0;
        i_10_1840 <= 0;
        i_10_1841 <= 0;
        i_10_1842 <= 0;
        i_10_1843 <= 0;
        i_10_1844 <= 0;
        i_10_1845 <= 0;
        i_10_1846 <= 0;
        i_10_1847 <= 0;
        i_10_1848 <= 0;
        i_10_1849 <= 0;
        i_10_1850 <= 0;
        i_10_1851 <= 0;
        i_10_1852 <= 0;
        i_10_1853 <= 0;
        i_10_1854 <= 0;
        i_10_1855 <= 0;
        i_10_1856 <= 0;
        i_10_1857 <= 0;
        i_10_1858 <= 0;
        i_10_1859 <= 0;
        i_10_1860 <= 0;
        i_10_1861 <= 0;
        i_10_1862 <= 0;
        i_10_1863 <= 0;
        i_10_1864 <= 0;
        i_10_1865 <= 0;
        i_10_1866 <= 0;
        i_10_1867 <= 0;
        i_10_1868 <= 0;
        i_10_1869 <= 0;
        i_10_1870 <= 0;
        i_10_1871 <= 0;
        i_10_1872 <= 0;
        i_10_1873 <= 0;
        i_10_1874 <= 0;
        i_10_1875 <= 0;
        i_10_1876 <= 0;
        i_10_1877 <= 0;
        i_10_1878 <= 0;
        i_10_1879 <= 0;
        i_10_1880 <= 0;
        i_10_1881 <= 0;
        i_10_1882 <= 0;
        i_10_1883 <= 0;
        i_10_1884 <= 0;
        i_10_1885 <= 0;
        i_10_1886 <= 0;
        i_10_1887 <= 0;
        i_10_1888 <= 0;
        i_10_1889 <= 0;
        i_10_1890 <= 0;
        i_10_1891 <= 0;
        i_10_1892 <= 0;
        i_10_1893 <= 0;
        i_10_1894 <= 0;
        i_10_1895 <= 0;
        i_10_1896 <= 0;
        i_10_1897 <= 0;
        i_10_1898 <= 0;
        i_10_1899 <= 0;
        i_10_1900 <= 0;
        i_10_1901 <= 0;
        i_10_1902 <= 0;
        i_10_1903 <= 0;
        i_10_1904 <= 0;
        i_10_1905 <= 0;
        i_10_1906 <= 0;
        i_10_1907 <= 0;
        i_10_1908 <= 0;
        i_10_1909 <= 0;
        i_10_1910 <= 0;
        i_10_1911 <= 0;
        i_10_1912 <= 0;
        i_10_1913 <= 0;
        i_10_1914 <= 0;
        i_10_1915 <= 0;
        i_10_1916 <= 0;
        i_10_1917 <= 0;
        i_10_1918 <= 0;
        i_10_1919 <= 0;
        i_10_1920 <= 0;
        i_10_1921 <= 0;
        i_10_1922 <= 0;
        i_10_1923 <= 0;
        i_10_1924 <= 0;
        i_10_1925 <= 0;
        i_10_1926 <= 0;
        i_10_1927 <= 0;
        i_10_1928 <= 0;
        i_10_1929 <= 0;
        i_10_1930 <= 0;
        i_10_1931 <= 0;
        i_10_1932 <= 0;
        i_10_1933 <= 0;
        i_10_1934 <= 0;
        i_10_1935 <= 0;
        i_10_1936 <= 0;
        i_10_1937 <= 0;
        i_10_1938 <= 0;
        i_10_1939 <= 0;
        i_10_1940 <= 0;
        i_10_1941 <= 0;
        i_10_1942 <= 0;
        i_10_1943 <= 0;
        i_10_1944 <= 0;
        i_10_1945 <= 0;
        i_10_1946 <= 0;
        i_10_1947 <= 0;
        i_10_1948 <= 0;
        i_10_1949 <= 0;
        i_10_1950 <= 0;
        i_10_1951 <= 0;
        i_10_1952 <= 0;
        i_10_1953 <= 0;
        i_10_1954 <= 0;
        i_10_1955 <= 0;
        i_10_1956 <= 0;
        i_10_1957 <= 0;
        i_10_1958 <= 0;
        i_10_1959 <= 0;
        i_10_1960 <= 0;
        i_10_1961 <= 0;
        i_10_1962 <= 0;
        i_10_1963 <= 0;
        i_10_1964 <= 0;
        i_10_1965 <= 0;
        i_10_1966 <= 0;
        i_10_1967 <= 0;
        i_10_1968 <= 0;
        i_10_1969 <= 0;
        i_10_1970 <= 0;
        i_10_1971 <= 0;
        i_10_1972 <= 0;
        i_10_1973 <= 0;
        i_10_1974 <= 0;
        i_10_1975 <= 0;
        i_10_1976 <= 0;
        i_10_1977 <= 0;
        i_10_1978 <= 0;
        i_10_1979 <= 0;
        i_10_1980 <= 0;
        i_10_1981 <= 0;
        i_10_1982 <= 0;
        i_10_1983 <= 0;
        i_10_1984 <= 0;
        i_10_1985 <= 0;
        i_10_1986 <= 0;
        i_10_1987 <= 0;
        i_10_1988 <= 0;
        i_10_1989 <= 0;
        i_10_1990 <= 0;
        i_10_1991 <= 0;
        i_10_1992 <= 0;
        i_10_1993 <= 0;
        i_10_1994 <= 0;
        i_10_1995 <= 0;
        i_10_1996 <= 0;
        i_10_1997 <= 0;
        i_10_1998 <= 0;
        i_10_1999 <= 0;
        i_10_2000 <= 0;
        i_10_2001 <= 0;
        i_10_2002 <= 0;
        i_10_2003 <= 0;
        i_10_2004 <= 0;
        i_10_2005 <= 0;
        i_10_2006 <= 0;
        i_10_2007 <= 0;
        i_10_2008 <= 0;
        i_10_2009 <= 0;
        i_10_2010 <= 0;
        i_10_2011 <= 0;
        i_10_2012 <= 0;
        i_10_2013 <= 0;
        i_10_2014 <= 0;
        i_10_2015 <= 0;
        i_10_2016 <= 0;
        i_10_2017 <= 0;
        i_10_2018 <= 0;
        i_10_2019 <= 0;
        i_10_2020 <= 0;
        i_10_2021 <= 0;
        i_10_2022 <= 0;
        i_10_2023 <= 0;
        i_10_2024 <= 0;
        i_10_2025 <= 0;
        i_10_2026 <= 0;
        i_10_2027 <= 0;
        i_10_2028 <= 0;
        i_10_2029 <= 0;
        i_10_2030 <= 0;
        i_10_2031 <= 0;
        i_10_2032 <= 0;
        i_10_2033 <= 0;
        i_10_2034 <= 0;
        i_10_2035 <= 0;
        i_10_2036 <= 0;
        i_10_2037 <= 0;
        i_10_2038 <= 0;
        i_10_2039 <= 0;
        i_10_2040 <= 0;
        i_10_2041 <= 0;
        i_10_2042 <= 0;
        i_10_2043 <= 0;
        i_10_2044 <= 0;
        i_10_2045 <= 0;
        i_10_2046 <= 0;
        i_10_2047 <= 0;
        i_10_2048 <= 0;
        i_10_2049 <= 0;
        i_10_2050 <= 0;
        i_10_2051 <= 0;
        i_10_2052 <= 0;
        i_10_2053 <= 0;
        i_10_2054 <= 0;
        i_10_2055 <= 0;
        i_10_2056 <= 0;
        i_10_2057 <= 0;
        i_10_2058 <= 0;
        i_10_2059 <= 0;
        i_10_2060 <= 0;
        i_10_2061 <= 0;
        i_10_2062 <= 0;
        i_10_2063 <= 0;
        i_10_2064 <= 0;
        i_10_2065 <= 0;
        i_10_2066 <= 0;
        i_10_2067 <= 0;
        i_10_2068 <= 0;
        i_10_2069 <= 0;
        i_10_2070 <= 0;
        i_10_2071 <= 0;
        i_10_2072 <= 0;
        i_10_2073 <= 0;
        i_10_2074 <= 0;
        i_10_2075 <= 0;
        i_10_2076 <= 0;
        i_10_2077 <= 0;
        i_10_2078 <= 0;
        i_10_2079 <= 0;
        i_10_2080 <= 0;
        i_10_2081 <= 0;
        i_10_2082 <= 0;
        i_10_2083 <= 0;
        i_10_2084 <= 0;
        i_10_2085 <= 0;
        i_10_2086 <= 0;
        i_10_2087 <= 0;
        i_10_2088 <= 0;
        i_10_2089 <= 0;
        i_10_2090 <= 0;
        i_10_2091 <= 0;
        i_10_2092 <= 0;
        i_10_2093 <= 0;
        i_10_2094 <= 0;
        i_10_2095 <= 0;
        i_10_2096 <= 0;
        i_10_2097 <= 0;
        i_10_2098 <= 0;
        i_10_2099 <= 0;
        i_10_2100 <= 0;
        i_10_2101 <= 0;
        i_10_2102 <= 0;
        i_10_2103 <= 0;
        i_10_2104 <= 0;
        i_10_2105 <= 0;
        i_10_2106 <= 0;
        i_10_2107 <= 0;
        i_10_2108 <= 0;
        i_10_2109 <= 0;
        i_10_2110 <= 0;
        i_10_2111 <= 0;
        i_10_2112 <= 0;
        i_10_2113 <= 0;
        i_10_2114 <= 0;
        i_10_2115 <= 0;
        i_10_2116 <= 0;
        i_10_2117 <= 0;
        i_10_2118 <= 0;
        i_10_2119 <= 0;
        i_10_2120 <= 0;
        i_10_2121 <= 0;
        i_10_2122 <= 0;
        i_10_2123 <= 0;
        i_10_2124 <= 0;
        i_10_2125 <= 0;
        i_10_2126 <= 0;
        i_10_2127 <= 0;
        i_10_2128 <= 0;
        i_10_2129 <= 0;
        i_10_2130 <= 0;
        i_10_2131 <= 0;
        i_10_2132 <= 0;
        i_10_2133 <= 0;
        i_10_2134 <= 0;
        i_10_2135 <= 0;
        i_10_2136 <= 0;
        i_10_2137 <= 0;
        i_10_2138 <= 0;
        i_10_2139 <= 0;
        i_10_2140 <= 0;
        i_10_2141 <= 0;
        i_10_2142 <= 0;
        i_10_2143 <= 0;
        i_10_2144 <= 0;
        i_10_2145 <= 0;
        i_10_2146 <= 0;
        i_10_2147 <= 0;
        i_10_2148 <= 0;
        i_10_2149 <= 0;
        i_10_2150 <= 0;
        i_10_2151 <= 0;
        i_10_2152 <= 0;
        i_10_2153 <= 0;
        i_10_2154 <= 0;
        i_10_2155 <= 0;
        i_10_2156 <= 0;
        i_10_2157 <= 0;
        i_10_2158 <= 0;
        i_10_2159 <= 0;
        i_10_2160 <= 0;
        i_10_2161 <= 0;
        i_10_2162 <= 0;
        i_10_2163 <= 0;
        i_10_2164 <= 0;
        i_10_2165 <= 0;
        i_10_2166 <= 0;
        i_10_2167 <= 0;
        i_10_2168 <= 0;
        i_10_2169 <= 0;
        i_10_2170 <= 0;
        i_10_2171 <= 0;
        i_10_2172 <= 0;
        i_10_2173 <= 0;
        i_10_2174 <= 0;
        i_10_2175 <= 0;
        i_10_2176 <= 0;
        i_10_2177 <= 0;
        i_10_2178 <= 0;
        i_10_2179 <= 0;
        i_10_2180 <= 0;
        i_10_2181 <= 0;
        i_10_2182 <= 0;
        i_10_2183 <= 0;
        i_10_2184 <= 0;
        i_10_2185 <= 0;
        i_10_2186 <= 0;
        i_10_2187 <= 0;
        i_10_2188 <= 0;
        i_10_2189 <= 0;
        i_10_2190 <= 0;
        i_10_2191 <= 0;
        i_10_2192 <= 0;
        i_10_2193 <= 0;
        i_10_2194 <= 0;
        i_10_2195 <= 0;
        i_10_2196 <= 0;
        i_10_2197 <= 0;
        i_10_2198 <= 0;
        i_10_2199 <= 0;
        i_10_2200 <= 0;
        i_10_2201 <= 0;
        i_10_2202 <= 0;
        i_10_2203 <= 0;
        i_10_2204 <= 0;
        i_10_2205 <= 0;
        i_10_2206 <= 0;
        i_10_2207 <= 0;
        i_10_2208 <= 0;
        i_10_2209 <= 0;
        i_10_2210 <= 0;
        i_10_2211 <= 0;
        i_10_2212 <= 0;
        i_10_2213 <= 0;
        i_10_2214 <= 0;
        i_10_2215 <= 0;
        i_10_2216 <= 0;
        i_10_2217 <= 0;
        i_10_2218 <= 0;
        i_10_2219 <= 0;
        i_10_2220 <= 0;
        i_10_2221 <= 0;
        i_10_2222 <= 0;
        i_10_2223 <= 0;
        i_10_2224 <= 0;
        i_10_2225 <= 0;
        i_10_2226 <= 0;
        i_10_2227 <= 0;
        i_10_2228 <= 0;
        i_10_2229 <= 0;
        i_10_2230 <= 0;
        i_10_2231 <= 0;
        i_10_2232 <= 0;
        i_10_2233 <= 0;
        i_10_2234 <= 0;
        i_10_2235 <= 0;
        i_10_2236 <= 0;
        i_10_2237 <= 0;
        i_10_2238 <= 0;
        i_10_2239 <= 0;
        i_10_2240 <= 0;
        i_10_2241 <= 0;
        i_10_2242 <= 0;
        i_10_2243 <= 0;
        i_10_2244 <= 0;
        i_10_2245 <= 0;
        i_10_2246 <= 0;
        i_10_2247 <= 0;
        i_10_2248 <= 0;
        i_10_2249 <= 0;
        i_10_2250 <= 0;
        i_10_2251 <= 0;
        i_10_2252 <= 0;
        i_10_2253 <= 0;
        i_10_2254 <= 0;
        i_10_2255 <= 0;
        i_10_2256 <= 0;
        i_10_2257 <= 0;
        i_10_2258 <= 0;
        i_10_2259 <= 0;
        i_10_2260 <= 0;
        i_10_2261 <= 0;
        i_10_2262 <= 0;
        i_10_2263 <= 0;
        i_10_2264 <= 0;
        i_10_2265 <= 0;
        i_10_2266 <= 0;
        i_10_2267 <= 0;
        i_10_2268 <= 0;
        i_10_2269 <= 0;
        i_10_2270 <= 0;
        i_10_2271 <= 0;
        i_10_2272 <= 0;
        i_10_2273 <= 0;
        i_10_2274 <= 0;
        i_10_2275 <= 0;
        i_10_2276 <= 0;
        i_10_2277 <= 0;
        i_10_2278 <= 0;
        i_10_2279 <= 0;
        i_10_2280 <= 0;
        i_10_2281 <= 0;
        i_10_2282 <= 0;
        i_10_2283 <= 0;
        i_10_2284 <= 0;
        i_10_2285 <= 0;
        i_10_2286 <= 0;
        i_10_2287 <= 0;
        i_10_2288 <= 0;
        i_10_2289 <= 0;
        i_10_2290 <= 0;
        i_10_2291 <= 0;
        i_10_2292 <= 0;
        i_10_2293 <= 0;
        i_10_2294 <= 0;
        i_10_2295 <= 0;
        i_10_2296 <= 0;
        i_10_2297 <= 0;
        i_10_2298 <= 0;
        i_10_2299 <= 0;
        i_10_2300 <= 0;
        i_10_2301 <= 0;
        i_10_2302 <= 0;
        i_10_2303 <= 0;
        i_10_2304 <= 0;
        i_10_2305 <= 0;
        i_10_2306 <= 0;
        i_10_2307 <= 0;
        i_10_2308 <= 0;
        i_10_2309 <= 0;
        i_10_2310 <= 0;
        i_10_2311 <= 0;
        i_10_2312 <= 0;
        i_10_2313 <= 0;
        i_10_2314 <= 0;
        i_10_2315 <= 0;
        i_10_2316 <= 0;
        i_10_2317 <= 0;
        i_10_2318 <= 0;
        i_10_2319 <= 0;
        i_10_2320 <= 0;
        i_10_2321 <= 0;
        i_10_2322 <= 0;
        i_10_2323 <= 0;
        i_10_2324 <= 0;
        i_10_2325 <= 0;
        i_10_2326 <= 0;
        i_10_2327 <= 0;
        i_10_2328 <= 0;
        i_10_2329 <= 0;
        i_10_2330 <= 0;
        i_10_2331 <= 0;
        i_10_2332 <= 0;
        i_10_2333 <= 0;
        i_10_2334 <= 0;
        i_10_2335 <= 0;
        i_10_2336 <= 0;
        i_10_2337 <= 0;
        i_10_2338 <= 0;
        i_10_2339 <= 0;
        i_10_2340 <= 0;
        i_10_2341 <= 0;
        i_10_2342 <= 0;
        i_10_2343 <= 0;
        i_10_2344 <= 0;
        i_10_2345 <= 0;
        i_10_2346 <= 0;
        i_10_2347 <= 0;
        i_10_2348 <= 0;
        i_10_2349 <= 0;
        i_10_2350 <= 0;
        i_10_2351 <= 0;
        i_10_2352 <= 0;
        i_10_2353 <= 0;
        i_10_2354 <= 0;
        i_10_2355 <= 0;
        i_10_2356 <= 0;
        i_10_2357 <= 0;
        i_10_2358 <= 0;
        i_10_2359 <= 0;
        i_10_2360 <= 0;
        i_10_2361 <= 0;
        i_10_2362 <= 0;
        i_10_2363 <= 0;
        i_10_2364 <= 0;
        i_10_2365 <= 0;
        i_10_2366 <= 0;
        i_10_2367 <= 0;
        i_10_2368 <= 0;
        i_10_2369 <= 0;
        i_10_2370 <= 0;
        i_10_2371 <= 0;
        i_10_2372 <= 0;
        i_10_2373 <= 0;
        i_10_2374 <= 0;
        i_10_2375 <= 0;
        i_10_2376 <= 0;
        i_10_2377 <= 0;
        i_10_2378 <= 0;
        i_10_2379 <= 0;
        i_10_2380 <= 0;
        i_10_2381 <= 0;
        i_10_2382 <= 0;
        i_10_2383 <= 0;
        i_10_2384 <= 0;
        i_10_2385 <= 0;
        i_10_2386 <= 0;
        i_10_2387 <= 0;
        i_10_2388 <= 0;
        i_10_2389 <= 0;
        i_10_2390 <= 0;
        i_10_2391 <= 0;
        i_10_2392 <= 0;
        i_10_2393 <= 0;
        i_10_2394 <= 0;
        i_10_2395 <= 0;
        i_10_2396 <= 0;
        i_10_2397 <= 0;
        i_10_2398 <= 0;
        i_10_2399 <= 0;
        i_10_2400 <= 0;
        i_10_2401 <= 0;
        i_10_2402 <= 0;
        i_10_2403 <= 0;
        i_10_2404 <= 0;
        i_10_2405 <= 0;
        i_10_2406 <= 0;
        i_10_2407 <= 0;
        i_10_2408 <= 0;
        i_10_2409 <= 0;
        i_10_2410 <= 0;
        i_10_2411 <= 0;
        i_10_2412 <= 0;
        i_10_2413 <= 0;
        i_10_2414 <= 0;
        i_10_2415 <= 0;
        i_10_2416 <= 0;
        i_10_2417 <= 0;
        i_10_2418 <= 0;
        i_10_2419 <= 0;
        i_10_2420 <= 0;
        i_10_2421 <= 0;
        i_10_2422 <= 0;
        i_10_2423 <= 0;
        i_10_2424 <= 0;
        i_10_2425 <= 0;
        i_10_2426 <= 0;
        i_10_2427 <= 0;
        i_10_2428 <= 0;
        i_10_2429 <= 0;
        i_10_2430 <= 0;
        i_10_2431 <= 0;
        i_10_2432 <= 0;
        i_10_2433 <= 0;
        i_10_2434 <= 0;
        i_10_2435 <= 0;
        i_10_2436 <= 0;
        i_10_2437 <= 0;
        i_10_2438 <= 0;
        i_10_2439 <= 0;
        i_10_2440 <= 0;
        i_10_2441 <= 0;
        i_10_2442 <= 0;
        i_10_2443 <= 0;
        i_10_2444 <= 0;
        i_10_2445 <= 0;
        i_10_2446 <= 0;
        i_10_2447 <= 0;
        i_10_2448 <= 0;
        i_10_2449 <= 0;
        i_10_2450 <= 0;
        i_10_2451 <= 0;
        i_10_2452 <= 0;
        i_10_2453 <= 0;
        i_10_2454 <= 0;
        i_10_2455 <= 0;
        i_10_2456 <= 0;
        i_10_2457 <= 0;
        i_10_2458 <= 0;
        i_10_2459 <= 0;
        i_10_2460 <= 0;
        i_10_2461 <= 0;
        i_10_2462 <= 0;
        i_10_2463 <= 0;
        i_10_2464 <= 0;
        i_10_2465 <= 0;
        i_10_2466 <= 0;
        i_10_2467 <= 0;
        i_10_2468 <= 0;
        i_10_2469 <= 0;
        i_10_2470 <= 0;
        i_10_2471 <= 0;
        i_10_2472 <= 0;
        i_10_2473 <= 0;
        i_10_2474 <= 0;
        i_10_2475 <= 0;
        i_10_2476 <= 0;
        i_10_2477 <= 0;
        i_10_2478 <= 0;
        i_10_2479 <= 0;
        i_10_2480 <= 0;
        i_10_2481 <= 0;
        i_10_2482 <= 0;
        i_10_2483 <= 0;
        i_10_2484 <= 0;
        i_10_2485 <= 0;
        i_10_2486 <= 0;
        i_10_2487 <= 0;
        i_10_2488 <= 0;
        i_10_2489 <= 0;
        i_10_2490 <= 0;
        i_10_2491 <= 0;
        i_10_2492 <= 0;
        i_10_2493 <= 0;
        i_10_2494 <= 0;
        i_10_2495 <= 0;
        i_10_2496 <= 0;
        i_10_2497 <= 0;
        i_10_2498 <= 0;
        i_10_2499 <= 0;
        i_10_2500 <= 0;
        i_10_2501 <= 0;
        i_10_2502 <= 0;
        i_10_2503 <= 0;
        i_10_2504 <= 0;
        i_10_2505 <= 0;
        i_10_2506 <= 0;
        i_10_2507 <= 0;
        i_10_2508 <= 0;
        i_10_2509 <= 0;
        i_10_2510 <= 0;
        i_10_2511 <= 0;
        i_10_2512 <= 0;
        i_10_2513 <= 0;
        i_10_2514 <= 0;
        i_10_2515 <= 0;
        i_10_2516 <= 0;
        i_10_2517 <= 0;
        i_10_2518 <= 0;
        i_10_2519 <= 0;
        i_10_2520 <= 0;
        i_10_2521 <= 0;
        i_10_2522 <= 0;
        i_10_2523 <= 0;
        i_10_2524 <= 0;
        i_10_2525 <= 0;
        i_10_2526 <= 0;
        i_10_2527 <= 0;
        i_10_2528 <= 0;
        i_10_2529 <= 0;
        i_10_2530 <= 0;
        i_10_2531 <= 0;
        i_10_2532 <= 0;
        i_10_2533 <= 0;
        i_10_2534 <= 0;
        i_10_2535 <= 0;
        i_10_2536 <= 0;
        i_10_2537 <= 0;
        i_10_2538 <= 0;
        i_10_2539 <= 0;
        i_10_2540 <= 0;
        i_10_2541 <= 0;
        i_10_2542 <= 0;
        i_10_2543 <= 0;
        i_10_2544 <= 0;
        i_10_2545 <= 0;
        i_10_2546 <= 0;
        i_10_2547 <= 0;
        i_10_2548 <= 0;
        i_10_2549 <= 0;
        i_10_2550 <= 0;
        i_10_2551 <= 0;
        i_10_2552 <= 0;
        i_10_2553 <= 0;
        i_10_2554 <= 0;
        i_10_2555 <= 0;
        i_10_2556 <= 0;
        i_10_2557 <= 0;
        i_10_2558 <= 0;
        i_10_2559 <= 0;
        i_10_2560 <= 0;
        i_10_2561 <= 0;
        i_10_2562 <= 0;
        i_10_2563 <= 0;
        i_10_2564 <= 0;
        i_10_2565 <= 0;
        i_10_2566 <= 0;
        i_10_2567 <= 0;
        i_10_2568 <= 0;
        i_10_2569 <= 0;
        i_10_2570 <= 0;
        i_10_2571 <= 0;
        i_10_2572 <= 0;
        i_10_2573 <= 0;
        i_10_2574 <= 0;
        i_10_2575 <= 0;
        i_10_2576 <= 0;
        i_10_2577 <= 0;
        i_10_2578 <= 0;
        i_10_2579 <= 0;
        i_10_2580 <= 0;
        i_10_2581 <= 0;
        i_10_2582 <= 0;
        i_10_2583 <= 0;
        i_10_2584 <= 0;
        i_10_2585 <= 0;
        i_10_2586 <= 0;
        i_10_2587 <= 0;
        i_10_2588 <= 0;
        i_10_2589 <= 0;
        i_10_2590 <= 0;
        i_10_2591 <= 0;
        i_10_2592 <= 0;
        i_10_2593 <= 0;
        i_10_2594 <= 0;
        i_10_2595 <= 0;
        i_10_2596 <= 0;
        i_10_2597 <= 0;
        i_10_2598 <= 0;
        i_10_2599 <= 0;
        i_10_2600 <= 0;
        i_10_2601 <= 0;
        i_10_2602 <= 0;
        i_10_2603 <= 0;
        i_10_2604 <= 0;
        i_10_2605 <= 0;
        i_10_2606 <= 0;
        i_10_2607 <= 0;
        i_10_2608 <= 0;
        i_10_2609 <= 0;
        i_10_2610 <= 0;
        i_10_2611 <= 0;
        i_10_2612 <= 0;
        i_10_2613 <= 0;
        i_10_2614 <= 0;
        i_10_2615 <= 0;
        i_10_2616 <= 0;
        i_10_2617 <= 0;
        i_10_2618 <= 0;
        i_10_2619 <= 0;
        i_10_2620 <= 0;
        i_10_2621 <= 0;
        i_10_2622 <= 0;
        i_10_2623 <= 0;
        i_10_2624 <= 0;
        i_10_2625 <= 0;
        i_10_2626 <= 0;
        i_10_2627 <= 0;
        i_10_2628 <= 0;
        i_10_2629 <= 0;
        i_10_2630 <= 0;
        i_10_2631 <= 0;
        i_10_2632 <= 0;
        i_10_2633 <= 0;
        i_10_2634 <= 0;
        i_10_2635 <= 0;
        i_10_2636 <= 0;
        i_10_2637 <= 0;
        i_10_2638 <= 0;
        i_10_2639 <= 0;
        i_10_2640 <= 0;
        i_10_2641 <= 0;
        i_10_2642 <= 0;
        i_10_2643 <= 0;
        i_10_2644 <= 0;
        i_10_2645 <= 0;
        i_10_2646 <= 0;
        i_10_2647 <= 0;
        i_10_2648 <= 0;
        i_10_2649 <= 0;
        i_10_2650 <= 0;
        i_10_2651 <= 0;
        i_10_2652 <= 0;
        i_10_2653 <= 0;
        i_10_2654 <= 0;
        i_10_2655 <= 0;
        i_10_2656 <= 0;
        i_10_2657 <= 0;
        i_10_2658 <= 0;
        i_10_2659 <= 0;
        i_10_2660 <= 0;
        i_10_2661 <= 0;
        i_10_2662 <= 0;
        i_10_2663 <= 0;
        i_10_2664 <= 0;
        i_10_2665 <= 0;
        i_10_2666 <= 0;
        i_10_2667 <= 0;
        i_10_2668 <= 0;
        i_10_2669 <= 0;
        i_10_2670 <= 0;
        i_10_2671 <= 0;
        i_10_2672 <= 0;
        i_10_2673 <= 0;
        i_10_2674 <= 0;
        i_10_2675 <= 0;
        i_10_2676 <= 0;
        i_10_2677 <= 0;
        i_10_2678 <= 0;
        i_10_2679 <= 0;
        i_10_2680 <= 0;
        i_10_2681 <= 0;
        i_10_2682 <= 0;
        i_10_2683 <= 0;
        i_10_2684 <= 0;
        i_10_2685 <= 0;
        i_10_2686 <= 0;
        i_10_2687 <= 0;
        i_10_2688 <= 0;
        i_10_2689 <= 0;
        i_10_2690 <= 0;
        i_10_2691 <= 0;
        i_10_2692 <= 0;
        i_10_2693 <= 0;
        i_10_2694 <= 0;
        i_10_2695 <= 0;
        i_10_2696 <= 0;
        i_10_2697 <= 0;
        i_10_2698 <= 0;
        i_10_2699 <= 0;
        i_10_2700 <= 0;
        i_10_2701 <= 0;
        i_10_2702 <= 0;
        i_10_2703 <= 0;
        i_10_2704 <= 0;
        i_10_2705 <= 0;
        i_10_2706 <= 0;
        i_10_2707 <= 0;
        i_10_2708 <= 0;
        i_10_2709 <= 0;
        i_10_2710 <= 0;
        i_10_2711 <= 0;
        i_10_2712 <= 0;
        i_10_2713 <= 0;
        i_10_2714 <= 0;
        i_10_2715 <= 0;
        i_10_2716 <= 0;
        i_10_2717 <= 0;
        i_10_2718 <= 0;
        i_10_2719 <= 0;
        i_10_2720 <= 0;
        i_10_2721 <= 0;
        i_10_2722 <= 0;
        i_10_2723 <= 0;
        i_10_2724 <= 0;
        i_10_2725 <= 0;
        i_10_2726 <= 0;
        i_10_2727 <= 0;
        i_10_2728 <= 0;
        i_10_2729 <= 0;
        i_10_2730 <= 0;
        i_10_2731 <= 0;
        i_10_2732 <= 0;
        i_10_2733 <= 0;
        i_10_2734 <= 0;
        i_10_2735 <= 0;
        i_10_2736 <= 0;
        i_10_2737 <= 0;
        i_10_2738 <= 0;
        i_10_2739 <= 0;
        i_10_2740 <= 0;
        i_10_2741 <= 0;
        i_10_2742 <= 0;
        i_10_2743 <= 0;
        i_10_2744 <= 0;
        i_10_2745 <= 0;
        i_10_2746 <= 0;
        i_10_2747 <= 0;
        i_10_2748 <= 0;
        i_10_2749 <= 0;
        i_10_2750 <= 0;
        i_10_2751 <= 0;
        i_10_2752 <= 0;
        i_10_2753 <= 0;
        i_10_2754 <= 0;
        i_10_2755 <= 0;
        i_10_2756 <= 0;
        i_10_2757 <= 0;
        i_10_2758 <= 0;
        i_10_2759 <= 0;
        i_10_2760 <= 0;
        i_10_2761 <= 0;
        i_10_2762 <= 0;
        i_10_2763 <= 0;
        i_10_2764 <= 0;
        i_10_2765 <= 0;
        i_10_2766 <= 0;
        i_10_2767 <= 0;
        i_10_2768 <= 0;
        i_10_2769 <= 0;
        i_10_2770 <= 0;
        i_10_2771 <= 0;
        i_10_2772 <= 0;
        i_10_2773 <= 0;
        i_10_2774 <= 0;
        i_10_2775 <= 0;
        i_10_2776 <= 0;
        i_10_2777 <= 0;
        i_10_2778 <= 0;
        i_10_2779 <= 0;
        i_10_2780 <= 0;
        i_10_2781 <= 0;
        i_10_2782 <= 0;
        i_10_2783 <= 0;
        i_10_2784 <= 0;
        i_10_2785 <= 0;
        i_10_2786 <= 0;
        i_10_2787 <= 0;
        i_10_2788 <= 0;
        i_10_2789 <= 0;
        i_10_2790 <= 0;
        i_10_2791 <= 0;
        i_10_2792 <= 0;
        i_10_2793 <= 0;
        i_10_2794 <= 0;
        i_10_2795 <= 0;
        i_10_2796 <= 0;
        i_10_2797 <= 0;
        i_10_2798 <= 0;
        i_10_2799 <= 0;
        i_10_2800 <= 0;
        i_10_2801 <= 0;
        i_10_2802 <= 0;
        i_10_2803 <= 0;
        i_10_2804 <= 0;
        i_10_2805 <= 0;
        i_10_2806 <= 0;
        i_10_2807 <= 0;
        i_10_2808 <= 0;
        i_10_2809 <= 0;
        i_10_2810 <= 0;
        i_10_2811 <= 0;
        i_10_2812 <= 0;
        i_10_2813 <= 0;
        i_10_2814 <= 0;
        i_10_2815 <= 0;
        i_10_2816 <= 0;
        i_10_2817 <= 0;
        i_10_2818 <= 0;
        i_10_2819 <= 0;
        i_10_2820 <= 0;
        i_10_2821 <= 0;
        i_10_2822 <= 0;
        i_10_2823 <= 0;
        i_10_2824 <= 0;
        i_10_2825 <= 0;
        i_10_2826 <= 0;
        i_10_2827 <= 0;
        i_10_2828 <= 0;
        i_10_2829 <= 0;
        i_10_2830 <= 0;
        i_10_2831 <= 0;
        i_10_2832 <= 0;
        i_10_2833 <= 0;
        i_10_2834 <= 0;
        i_10_2835 <= 0;
        i_10_2836 <= 0;
        i_10_2837 <= 0;
        i_10_2838 <= 0;
        i_10_2839 <= 0;
        i_10_2840 <= 0;
        i_10_2841 <= 0;
        i_10_2842 <= 0;
        i_10_2843 <= 0;
        i_10_2844 <= 0;
        i_10_2845 <= 0;
        i_10_2846 <= 0;
        i_10_2847 <= 0;
        i_10_2848 <= 0;
        i_10_2849 <= 0;
        i_10_2850 <= 0;
        i_10_2851 <= 0;
        i_10_2852 <= 0;
        i_10_2853 <= 0;
        i_10_2854 <= 0;
        i_10_2855 <= 0;
        i_10_2856 <= 0;
        i_10_2857 <= 0;
        i_10_2858 <= 0;
        i_10_2859 <= 0;
        i_10_2860 <= 0;
        i_10_2861 <= 0;
        i_10_2862 <= 0;
        i_10_2863 <= 0;
        i_10_2864 <= 0;
        i_10_2865 <= 0;
        i_10_2866 <= 0;
        i_10_2867 <= 0;
        i_10_2868 <= 0;
        i_10_2869 <= 0;
        i_10_2870 <= 0;
        i_10_2871 <= 0;
        i_10_2872 <= 0;
        i_10_2873 <= 0;
        i_10_2874 <= 0;
        i_10_2875 <= 0;
        i_10_2876 <= 0;
        i_10_2877 <= 0;
        i_10_2878 <= 0;
        i_10_2879 <= 0;
        i_10_2880 <= 0;
        i_10_2881 <= 0;
        i_10_2882 <= 0;
        i_10_2883 <= 0;
        i_10_2884 <= 0;
        i_10_2885 <= 0;
        i_10_2886 <= 0;
        i_10_2887 <= 0;
        i_10_2888 <= 0;
        i_10_2889 <= 0;
        i_10_2890 <= 0;
        i_10_2891 <= 0;
        i_10_2892 <= 0;
        i_10_2893 <= 0;
        i_10_2894 <= 0;
        i_10_2895 <= 0;
        i_10_2896 <= 0;
        i_10_2897 <= 0;
        i_10_2898 <= 0;
        i_10_2899 <= 0;
        i_10_2900 <= 0;
        i_10_2901 <= 0;
        i_10_2902 <= 0;
        i_10_2903 <= 0;
        i_10_2904 <= 0;
        i_10_2905 <= 0;
        i_10_2906 <= 0;
        i_10_2907 <= 0;
        i_10_2908 <= 0;
        i_10_2909 <= 0;
        i_10_2910 <= 0;
        i_10_2911 <= 0;
        i_10_2912 <= 0;
        i_10_2913 <= 0;
        i_10_2914 <= 0;
        i_10_2915 <= 0;
        i_10_2916 <= 0;
        i_10_2917 <= 0;
        i_10_2918 <= 0;
        i_10_2919 <= 0;
        i_10_2920 <= 0;
        i_10_2921 <= 0;
        i_10_2922 <= 0;
        i_10_2923 <= 0;
        i_10_2924 <= 0;
        i_10_2925 <= 0;
        i_10_2926 <= 0;
        i_10_2927 <= 0;
        i_10_2928 <= 0;
        i_10_2929 <= 0;
        i_10_2930 <= 0;
        i_10_2931 <= 0;
        i_10_2932 <= 0;
        i_10_2933 <= 0;
        i_10_2934 <= 0;
        i_10_2935 <= 0;
        i_10_2936 <= 0;
        i_10_2937 <= 0;
        i_10_2938 <= 0;
        i_10_2939 <= 0;
        i_10_2940 <= 0;
        i_10_2941 <= 0;
        i_10_2942 <= 0;
        i_10_2943 <= 0;
        i_10_2944 <= 0;
        i_10_2945 <= 0;
        i_10_2946 <= 0;
        i_10_2947 <= 0;
        i_10_2948 <= 0;
        i_10_2949 <= 0;
        i_10_2950 <= 0;
        i_10_2951 <= 0;
        i_10_2952 <= 0;
        i_10_2953 <= 0;
        i_10_2954 <= 0;
        i_10_2955 <= 0;
        i_10_2956 <= 0;
        i_10_2957 <= 0;
        i_10_2958 <= 0;
        i_10_2959 <= 0;
        i_10_2960 <= 0;
        i_10_2961 <= 0;
        i_10_2962 <= 0;
        i_10_2963 <= 0;
        i_10_2964 <= 0;
        i_10_2965 <= 0;
        i_10_2966 <= 0;
        i_10_2967 <= 0;
        i_10_2968 <= 0;
        i_10_2969 <= 0;
        i_10_2970 <= 0;
        i_10_2971 <= 0;
        i_10_2972 <= 0;
        i_10_2973 <= 0;
        i_10_2974 <= 0;
        i_10_2975 <= 0;
        i_10_2976 <= 0;
        i_10_2977 <= 0;
        i_10_2978 <= 0;
        i_10_2979 <= 0;
        i_10_2980 <= 0;
        i_10_2981 <= 0;
        i_10_2982 <= 0;
        i_10_2983 <= 0;
        i_10_2984 <= 0;
        i_10_2985 <= 0;
        i_10_2986 <= 0;
        i_10_2987 <= 0;
        i_10_2988 <= 0;
        i_10_2989 <= 0;
        i_10_2990 <= 0;
        i_10_2991 <= 0;
        i_10_2992 <= 0;
        i_10_2993 <= 0;
        i_10_2994 <= 0;
        i_10_2995 <= 0;
        i_10_2996 <= 0;
        i_10_2997 <= 0;
        i_10_2998 <= 0;
        i_10_2999 <= 0;
        i_10_3000 <= 0;
        i_10_3001 <= 0;
        i_10_3002 <= 0;
        i_10_3003 <= 0;
        i_10_3004 <= 0;
        i_10_3005 <= 0;
        i_10_3006 <= 0;
        i_10_3007 <= 0;
        i_10_3008 <= 0;
        i_10_3009 <= 0;
        i_10_3010 <= 0;
        i_10_3011 <= 0;
        i_10_3012 <= 0;
        i_10_3013 <= 0;
        i_10_3014 <= 0;
        i_10_3015 <= 0;
        i_10_3016 <= 0;
        i_10_3017 <= 0;
        i_10_3018 <= 0;
        i_10_3019 <= 0;
        i_10_3020 <= 0;
        i_10_3021 <= 0;
        i_10_3022 <= 0;
        i_10_3023 <= 0;
        i_10_3024 <= 0;
        i_10_3025 <= 0;
        i_10_3026 <= 0;
        i_10_3027 <= 0;
        i_10_3028 <= 0;
        i_10_3029 <= 0;
        i_10_3030 <= 0;
        i_10_3031 <= 0;
        i_10_3032 <= 0;
        i_10_3033 <= 0;
        i_10_3034 <= 0;
        i_10_3035 <= 0;
        i_10_3036 <= 0;
        i_10_3037 <= 0;
        i_10_3038 <= 0;
        i_10_3039 <= 0;
        i_10_3040 <= 0;
        i_10_3041 <= 0;
        i_10_3042 <= 0;
        i_10_3043 <= 0;
        i_10_3044 <= 0;
        i_10_3045 <= 0;
        i_10_3046 <= 0;
        i_10_3047 <= 0;
        i_10_3048 <= 0;
        i_10_3049 <= 0;
        i_10_3050 <= 0;
        i_10_3051 <= 0;
        i_10_3052 <= 0;
        i_10_3053 <= 0;
        i_10_3054 <= 0;
        i_10_3055 <= 0;
        i_10_3056 <= 0;
        i_10_3057 <= 0;
        i_10_3058 <= 0;
        i_10_3059 <= 0;
        i_10_3060 <= 0;
        i_10_3061 <= 0;
        i_10_3062 <= 0;
        i_10_3063 <= 0;
        i_10_3064 <= 0;
        i_10_3065 <= 0;
        i_10_3066 <= 0;
        i_10_3067 <= 0;
        i_10_3068 <= 0;
        i_10_3069 <= 0;
        i_10_3070 <= 0;
        i_10_3071 <= 0;
        i_10_3072 <= 0;
        i_10_3073 <= 0;
        i_10_3074 <= 0;
        i_10_3075 <= 0;
        i_10_3076 <= 0;
        i_10_3077 <= 0;
        i_10_3078 <= 0;
        i_10_3079 <= 0;
        i_10_3080 <= 0;
        i_10_3081 <= 0;
        i_10_3082 <= 0;
        i_10_3083 <= 0;
        i_10_3084 <= 0;
        i_10_3085 <= 0;
        i_10_3086 <= 0;
        i_10_3087 <= 0;
        i_10_3088 <= 0;
        i_10_3089 <= 0;
        i_10_3090 <= 0;
        i_10_3091 <= 0;
        i_10_3092 <= 0;
        i_10_3093 <= 0;
        i_10_3094 <= 0;
        i_10_3095 <= 0;
        i_10_3096 <= 0;
        i_10_3097 <= 0;
        i_10_3098 <= 0;
        i_10_3099 <= 0;
        i_10_3100 <= 0;
        i_10_3101 <= 0;
        i_10_3102 <= 0;
        i_10_3103 <= 0;
        i_10_3104 <= 0;
        i_10_3105 <= 0;
        i_10_3106 <= 0;
        i_10_3107 <= 0;
        i_10_3108 <= 0;
        i_10_3109 <= 0;
        i_10_3110 <= 0;
        i_10_3111 <= 0;
        i_10_3112 <= 0;
        i_10_3113 <= 0;
        i_10_3114 <= 0;
        i_10_3115 <= 0;
        i_10_3116 <= 0;
        i_10_3117 <= 0;
        i_10_3118 <= 0;
        i_10_3119 <= 0;
        i_10_3120 <= 0;
        i_10_3121 <= 0;
        i_10_3122 <= 0;
        i_10_3123 <= 0;
        i_10_3124 <= 0;
        i_10_3125 <= 0;
        i_10_3126 <= 0;
        i_10_3127 <= 0;
        i_10_3128 <= 0;
        i_10_3129 <= 0;
        i_10_3130 <= 0;
        i_10_3131 <= 0;
        i_10_3132 <= 0;
        i_10_3133 <= 0;
        i_10_3134 <= 0;
        i_10_3135 <= 0;
        i_10_3136 <= 0;
        i_10_3137 <= 0;
        i_10_3138 <= 0;
        i_10_3139 <= 0;
        i_10_3140 <= 0;
        i_10_3141 <= 0;
        i_10_3142 <= 0;
        i_10_3143 <= 0;
        i_10_3144 <= 0;
        i_10_3145 <= 0;
        i_10_3146 <= 0;
        i_10_3147 <= 0;
        i_10_3148 <= 0;
        i_10_3149 <= 0;
        i_10_3150 <= 0;
        i_10_3151 <= 0;
        i_10_3152 <= 0;
        i_10_3153 <= 0;
        i_10_3154 <= 0;
        i_10_3155 <= 0;
        i_10_3156 <= 0;
        i_10_3157 <= 0;
        i_10_3158 <= 0;
        i_10_3159 <= 0;
        i_10_3160 <= 0;
        i_10_3161 <= 0;
        i_10_3162 <= 0;
        i_10_3163 <= 0;
        i_10_3164 <= 0;
        i_10_3165 <= 0;
        i_10_3166 <= 0;
        i_10_3167 <= 0;
        i_10_3168 <= 0;
        i_10_3169 <= 0;
        i_10_3170 <= 0;
        i_10_3171 <= 0;
        i_10_3172 <= 0;
        i_10_3173 <= 0;
        i_10_3174 <= 0;
        i_10_3175 <= 0;
        i_10_3176 <= 0;
        i_10_3177 <= 0;
        i_10_3178 <= 0;
        i_10_3179 <= 0;
        i_10_3180 <= 0;
        i_10_3181 <= 0;
        i_10_3182 <= 0;
        i_10_3183 <= 0;
        i_10_3184 <= 0;
        i_10_3185 <= 0;
        i_10_3186 <= 0;
        i_10_3187 <= 0;
        i_10_3188 <= 0;
        i_10_3189 <= 0;
        i_10_3190 <= 0;
        i_10_3191 <= 0;
        i_10_3192 <= 0;
        i_10_3193 <= 0;
        i_10_3194 <= 0;
        i_10_3195 <= 0;
        i_10_3196 <= 0;
        i_10_3197 <= 0;
        i_10_3198 <= 0;
        i_10_3199 <= 0;
        i_10_3200 <= 0;
        i_10_3201 <= 0;
        i_10_3202 <= 0;
        i_10_3203 <= 0;
        i_10_3204 <= 0;
        i_10_3205 <= 0;
        i_10_3206 <= 0;
        i_10_3207 <= 0;
        i_10_3208 <= 0;
        i_10_3209 <= 0;
        i_10_3210 <= 0;
        i_10_3211 <= 0;
        i_10_3212 <= 0;
        i_10_3213 <= 0;
        i_10_3214 <= 0;
        i_10_3215 <= 0;
        i_10_3216 <= 0;
        i_10_3217 <= 0;
        i_10_3218 <= 0;
        i_10_3219 <= 0;
        i_10_3220 <= 0;
        i_10_3221 <= 0;
        i_10_3222 <= 0;
        i_10_3223 <= 0;
        i_10_3224 <= 0;
        i_10_3225 <= 0;
        i_10_3226 <= 0;
        i_10_3227 <= 0;
        i_10_3228 <= 0;
        i_10_3229 <= 0;
        i_10_3230 <= 0;
        i_10_3231 <= 0;
        i_10_3232 <= 0;
        i_10_3233 <= 0;
        i_10_3234 <= 0;
        i_10_3235 <= 0;
        i_10_3236 <= 0;
        i_10_3237 <= 0;
        i_10_3238 <= 0;
        i_10_3239 <= 0;
        i_10_3240 <= 0;
        i_10_3241 <= 0;
        i_10_3242 <= 0;
        i_10_3243 <= 0;
        i_10_3244 <= 0;
        i_10_3245 <= 0;
        i_10_3246 <= 0;
        i_10_3247 <= 0;
        i_10_3248 <= 0;
        i_10_3249 <= 0;
        i_10_3250 <= 0;
        i_10_3251 <= 0;
        i_10_3252 <= 0;
        i_10_3253 <= 0;
        i_10_3254 <= 0;
        i_10_3255 <= 0;
        i_10_3256 <= 0;
        i_10_3257 <= 0;
        i_10_3258 <= 0;
        i_10_3259 <= 0;
        i_10_3260 <= 0;
        i_10_3261 <= 0;
        i_10_3262 <= 0;
        i_10_3263 <= 0;
        i_10_3264 <= 0;
        i_10_3265 <= 0;
        i_10_3266 <= 0;
        i_10_3267 <= 0;
        i_10_3268 <= 0;
        i_10_3269 <= 0;
        i_10_3270 <= 0;
        i_10_3271 <= 0;
        i_10_3272 <= 0;
        i_10_3273 <= 0;
        i_10_3274 <= 0;
        i_10_3275 <= 0;
        i_10_3276 <= 0;
        i_10_3277 <= 0;
        i_10_3278 <= 0;
        i_10_3279 <= 0;
        i_10_3280 <= 0;
        i_10_3281 <= 0;
        i_10_3282 <= 0;
        i_10_3283 <= 0;
        i_10_3284 <= 0;
        i_10_3285 <= 0;
        i_10_3286 <= 0;
        i_10_3287 <= 0;
        i_10_3288 <= 0;
        i_10_3289 <= 0;
        i_10_3290 <= 0;
        i_10_3291 <= 0;
        i_10_3292 <= 0;
        i_10_3293 <= 0;
        i_10_3294 <= 0;
        i_10_3295 <= 0;
        i_10_3296 <= 0;
        i_10_3297 <= 0;
        i_10_3298 <= 0;
        i_10_3299 <= 0;
        i_10_3300 <= 0;
        i_10_3301 <= 0;
        i_10_3302 <= 0;
        i_10_3303 <= 0;
        i_10_3304 <= 0;
        i_10_3305 <= 0;
        i_10_3306 <= 0;
        i_10_3307 <= 0;
        i_10_3308 <= 0;
        i_10_3309 <= 0;
        i_10_3310 <= 0;
        i_10_3311 <= 0;
        i_10_3312 <= 0;
        i_10_3313 <= 0;
        i_10_3314 <= 0;
        i_10_3315 <= 0;
        i_10_3316 <= 0;
        i_10_3317 <= 0;
        i_10_3318 <= 0;
        i_10_3319 <= 0;
        i_10_3320 <= 0;
        i_10_3321 <= 0;
        i_10_3322 <= 0;
        i_10_3323 <= 0;
        i_10_3324 <= 0;
        i_10_3325 <= 0;
        i_10_3326 <= 0;
        i_10_3327 <= 0;
        i_10_3328 <= 0;
        i_10_3329 <= 0;
        i_10_3330 <= 0;
        i_10_3331 <= 0;
        i_10_3332 <= 0;
        i_10_3333 <= 0;
        i_10_3334 <= 0;
        i_10_3335 <= 0;
        i_10_3336 <= 0;
        i_10_3337 <= 0;
        i_10_3338 <= 0;
        i_10_3339 <= 0;
        i_10_3340 <= 0;
        i_10_3341 <= 0;
        i_10_3342 <= 0;
        i_10_3343 <= 0;
        i_10_3344 <= 0;
        i_10_3345 <= 0;
        i_10_3346 <= 0;
        i_10_3347 <= 0;
        i_10_3348 <= 0;
        i_10_3349 <= 0;
        i_10_3350 <= 0;
        i_10_3351 <= 0;
        i_10_3352 <= 0;
        i_10_3353 <= 0;
        i_10_3354 <= 0;
        i_10_3355 <= 0;
        i_10_3356 <= 0;
        i_10_3357 <= 0;
        i_10_3358 <= 0;
        i_10_3359 <= 0;
        i_10_3360 <= 0;
        i_10_3361 <= 0;
        i_10_3362 <= 0;
        i_10_3363 <= 0;
        i_10_3364 <= 0;
        i_10_3365 <= 0;
        i_10_3366 <= 0;
        i_10_3367 <= 0;
        i_10_3368 <= 0;
        i_10_3369 <= 0;
        i_10_3370 <= 0;
        i_10_3371 <= 0;
        i_10_3372 <= 0;
        i_10_3373 <= 0;
        i_10_3374 <= 0;
        i_10_3375 <= 0;
        i_10_3376 <= 0;
        i_10_3377 <= 0;
        i_10_3378 <= 0;
        i_10_3379 <= 0;
        i_10_3380 <= 0;
        i_10_3381 <= 0;
        i_10_3382 <= 0;
        i_10_3383 <= 0;
        i_10_3384 <= 0;
        i_10_3385 <= 0;
        i_10_3386 <= 0;
        i_10_3387 <= 0;
        i_10_3388 <= 0;
        i_10_3389 <= 0;
        i_10_3390 <= 0;
        i_10_3391 <= 0;
        i_10_3392 <= 0;
        i_10_3393 <= 0;
        i_10_3394 <= 0;
        i_10_3395 <= 0;
        i_10_3396 <= 0;
        i_10_3397 <= 0;
        i_10_3398 <= 0;
        i_10_3399 <= 0;
        i_10_3400 <= 0;
        i_10_3401 <= 0;
        i_10_3402 <= 0;
        i_10_3403 <= 0;
        i_10_3404 <= 0;
        i_10_3405 <= 0;
        i_10_3406 <= 0;
        i_10_3407 <= 0;
        i_10_3408 <= 0;
        i_10_3409 <= 0;
        i_10_3410 <= 0;
        i_10_3411 <= 0;
        i_10_3412 <= 0;
        i_10_3413 <= 0;
        i_10_3414 <= 0;
        i_10_3415 <= 0;
        i_10_3416 <= 0;
        i_10_3417 <= 0;
        i_10_3418 <= 0;
        i_10_3419 <= 0;
        i_10_3420 <= 0;
        i_10_3421 <= 0;
        i_10_3422 <= 0;
        i_10_3423 <= 0;
        i_10_3424 <= 0;
        i_10_3425 <= 0;
        i_10_3426 <= 0;
        i_10_3427 <= 0;
        i_10_3428 <= 0;
        i_10_3429 <= 0;
        i_10_3430 <= 0;
        i_10_3431 <= 0;
        i_10_3432 <= 0;
        i_10_3433 <= 0;
        i_10_3434 <= 0;
        i_10_3435 <= 0;
        i_10_3436 <= 0;
        i_10_3437 <= 0;
        i_10_3438 <= 0;
        i_10_3439 <= 0;
        i_10_3440 <= 0;
        i_10_3441 <= 0;
        i_10_3442 <= 0;
        i_10_3443 <= 0;
        i_10_3444 <= 0;
        i_10_3445 <= 0;
        i_10_3446 <= 0;
        i_10_3447 <= 0;
        i_10_3448 <= 0;
        i_10_3449 <= 0;
        i_10_3450 <= 0;
        i_10_3451 <= 0;
        i_10_3452 <= 0;
        i_10_3453 <= 0;
        i_10_3454 <= 0;
        i_10_3455 <= 0;
        i_10_3456 <= 0;
        i_10_3457 <= 0;
        i_10_3458 <= 0;
        i_10_3459 <= 0;
        i_10_3460 <= 0;
        i_10_3461 <= 0;
        i_10_3462 <= 0;
        i_10_3463 <= 0;
        i_10_3464 <= 0;
        i_10_3465 <= 0;
        i_10_3466 <= 0;
        i_10_3467 <= 0;
        i_10_3468 <= 0;
        i_10_3469 <= 0;
        i_10_3470 <= 0;
        i_10_3471 <= 0;
        i_10_3472 <= 0;
        i_10_3473 <= 0;
        i_10_3474 <= 0;
        i_10_3475 <= 0;
        i_10_3476 <= 0;
        i_10_3477 <= 0;
        i_10_3478 <= 0;
        i_10_3479 <= 0;
        i_10_3480 <= 0;
        i_10_3481 <= 0;
        i_10_3482 <= 0;
        i_10_3483 <= 0;
        i_10_3484 <= 0;
        i_10_3485 <= 0;
        i_10_3486 <= 0;
        i_10_3487 <= 0;
        i_10_3488 <= 0;
        i_10_3489 <= 0;
        i_10_3490 <= 0;
        i_10_3491 <= 0;
        i_10_3492 <= 0;
        i_10_3493 <= 0;
        i_10_3494 <= 0;
        i_10_3495 <= 0;
        i_10_3496 <= 0;
        i_10_3497 <= 0;
        i_10_3498 <= 0;
        i_10_3499 <= 0;
        i_10_3500 <= 0;
        i_10_3501 <= 0;
        i_10_3502 <= 0;
        i_10_3503 <= 0;
        i_10_3504 <= 0;
        i_10_3505 <= 0;
        i_10_3506 <= 0;
        i_10_3507 <= 0;
        i_10_3508 <= 0;
        i_10_3509 <= 0;
        i_10_3510 <= 0;
        i_10_3511 <= 0;
        i_10_3512 <= 0;
        i_10_3513 <= 0;
        i_10_3514 <= 0;
        i_10_3515 <= 0;
        i_10_3516 <= 0;
        i_10_3517 <= 0;
        i_10_3518 <= 0;
        i_10_3519 <= 0;
        i_10_3520 <= 0;
        i_10_3521 <= 0;
        i_10_3522 <= 0;
        i_10_3523 <= 0;
        i_10_3524 <= 0;
        i_10_3525 <= 0;
        i_10_3526 <= 0;
        i_10_3527 <= 0;
        i_10_3528 <= 0;
        i_10_3529 <= 0;
        i_10_3530 <= 0;
        i_10_3531 <= 0;
        i_10_3532 <= 0;
        i_10_3533 <= 0;
        i_10_3534 <= 0;
        i_10_3535 <= 0;
        i_10_3536 <= 0;
        i_10_3537 <= 0;
        i_10_3538 <= 0;
        i_10_3539 <= 0;
        i_10_3540 <= 0;
        i_10_3541 <= 0;
        i_10_3542 <= 0;
        i_10_3543 <= 0;
        i_10_3544 <= 0;
        i_10_3545 <= 0;
        i_10_3546 <= 0;
        i_10_3547 <= 0;
        i_10_3548 <= 0;
        i_10_3549 <= 0;
        i_10_3550 <= 0;
        i_10_3551 <= 0;
        i_10_3552 <= 0;
        i_10_3553 <= 0;
        i_10_3554 <= 0;
        i_10_3555 <= 0;
        i_10_3556 <= 0;
        i_10_3557 <= 0;
        i_10_3558 <= 0;
        i_10_3559 <= 0;
        i_10_3560 <= 0;
        i_10_3561 <= 0;
        i_10_3562 <= 0;
        i_10_3563 <= 0;
        i_10_3564 <= 0;
        i_10_3565 <= 0;
        i_10_3566 <= 0;
        i_10_3567 <= 0;
        i_10_3568 <= 0;
        i_10_3569 <= 0;
        i_10_3570 <= 0;
        i_10_3571 <= 0;
        i_10_3572 <= 0;
        i_10_3573 <= 0;
        i_10_3574 <= 0;
        i_10_3575 <= 0;
        i_10_3576 <= 0;
        i_10_3577 <= 0;
        i_10_3578 <= 0;
        i_10_3579 <= 0;
        i_10_3580 <= 0;
        i_10_3581 <= 0;
        i_10_3582 <= 0;
        i_10_3583 <= 0;
        i_10_3584 <= 0;
        i_10_3585 <= 0;
        i_10_3586 <= 0;
        i_10_3587 <= 0;
        i_10_3588 <= 0;
        i_10_3589 <= 0;
        i_10_3590 <= 0;
        i_10_3591 <= 0;
        i_10_3592 <= 0;
        i_10_3593 <= 0;
        i_10_3594 <= 0;
        i_10_3595 <= 0;
        i_10_3596 <= 0;
        i_10_3597 <= 0;
        i_10_3598 <= 0;
        i_10_3599 <= 0;
        i_10_3600 <= 0;
        i_10_3601 <= 0;
        i_10_3602 <= 0;
        i_10_3603 <= 0;
        i_10_3604 <= 0;
        i_10_3605 <= 0;
        i_10_3606 <= 0;
        i_10_3607 <= 0;
        i_10_3608 <= 0;
        i_10_3609 <= 0;
        i_10_3610 <= 0;
        i_10_3611 <= 0;
        i_10_3612 <= 0;
        i_10_3613 <= 0;
        i_10_3614 <= 0;
        i_10_3615 <= 0;
        i_10_3616 <= 0;
        i_10_3617 <= 0;
        i_10_3618 <= 0;
        i_10_3619 <= 0;
        i_10_3620 <= 0;
        i_10_3621 <= 0;
        i_10_3622 <= 0;
        i_10_3623 <= 0;
        i_10_3624 <= 0;
        i_10_3625 <= 0;
        i_10_3626 <= 0;
        i_10_3627 <= 0;
        i_10_3628 <= 0;
        i_10_3629 <= 0;
        i_10_3630 <= 0;
        i_10_3631 <= 0;
        i_10_3632 <= 0;
        i_10_3633 <= 0;
        i_10_3634 <= 0;
        i_10_3635 <= 0;
        i_10_3636 <= 0;
        i_10_3637 <= 0;
        i_10_3638 <= 0;
        i_10_3639 <= 0;
        i_10_3640 <= 0;
        i_10_3641 <= 0;
        i_10_3642 <= 0;
        i_10_3643 <= 0;
        i_10_3644 <= 0;
        i_10_3645 <= 0;
        i_10_3646 <= 0;
        i_10_3647 <= 0;
        i_10_3648 <= 0;
        i_10_3649 <= 0;
        i_10_3650 <= 0;
        i_10_3651 <= 0;
        i_10_3652 <= 0;
        i_10_3653 <= 0;
        i_10_3654 <= 0;
        i_10_3655 <= 0;
        i_10_3656 <= 0;
        i_10_3657 <= 0;
        i_10_3658 <= 0;
        i_10_3659 <= 0;
        i_10_3660 <= 0;
        i_10_3661 <= 0;
        i_10_3662 <= 0;
        i_10_3663 <= 0;
        i_10_3664 <= 0;
        i_10_3665 <= 0;
        i_10_3666 <= 0;
        i_10_3667 <= 0;
        i_10_3668 <= 0;
        i_10_3669 <= 0;
        i_10_3670 <= 0;
        i_10_3671 <= 0;
        i_10_3672 <= 0;
        i_10_3673 <= 0;
        i_10_3674 <= 0;
        i_10_3675 <= 0;
        i_10_3676 <= 0;
        i_10_3677 <= 0;
        i_10_3678 <= 0;
        i_10_3679 <= 0;
        i_10_3680 <= 0;
        i_10_3681 <= 0;
        i_10_3682 <= 0;
        i_10_3683 <= 0;
        i_10_3684 <= 0;
        i_10_3685 <= 0;
        i_10_3686 <= 0;
        i_10_3687 <= 0;
        i_10_3688 <= 0;
        i_10_3689 <= 0;
        i_10_3690 <= 0;
        i_10_3691 <= 0;
        i_10_3692 <= 0;
        i_10_3693 <= 0;
        i_10_3694 <= 0;
        i_10_3695 <= 0;
        i_10_3696 <= 0;
        i_10_3697 <= 0;
        i_10_3698 <= 0;
        i_10_3699 <= 0;
        i_10_3700 <= 0;
        i_10_3701 <= 0;
        i_10_3702 <= 0;
        i_10_3703 <= 0;
        i_10_3704 <= 0;
        i_10_3705 <= 0;
        i_10_3706 <= 0;
        i_10_3707 <= 0;
        i_10_3708 <= 0;
        i_10_3709 <= 0;
        i_10_3710 <= 0;
        i_10_3711 <= 0;
        i_10_3712 <= 0;
        i_10_3713 <= 0;
        i_10_3714 <= 0;
        i_10_3715 <= 0;
        i_10_3716 <= 0;
        i_10_3717 <= 0;
        i_10_3718 <= 0;
        i_10_3719 <= 0;
        i_10_3720 <= 0;
        i_10_3721 <= 0;
        i_10_3722 <= 0;
        i_10_3723 <= 0;
        i_10_3724 <= 0;
        i_10_3725 <= 0;
        i_10_3726 <= 0;
        i_10_3727 <= 0;
        i_10_3728 <= 0;
        i_10_3729 <= 0;
        i_10_3730 <= 0;
        i_10_3731 <= 0;
        i_10_3732 <= 0;
        i_10_3733 <= 0;
        i_10_3734 <= 0;
        i_10_3735 <= 0;
        i_10_3736 <= 0;
        i_10_3737 <= 0;
        i_10_3738 <= 0;
        i_10_3739 <= 0;
        i_10_3740 <= 0;
        i_10_3741 <= 0;
        i_10_3742 <= 0;
        i_10_3743 <= 0;
        i_10_3744 <= 0;
        i_10_3745 <= 0;
        i_10_3746 <= 0;
        i_10_3747 <= 0;
        i_10_3748 <= 0;
        i_10_3749 <= 0;
        i_10_3750 <= 0;
        i_10_3751 <= 0;
        i_10_3752 <= 0;
        i_10_3753 <= 0;
        i_10_3754 <= 0;
        i_10_3755 <= 0;
        i_10_3756 <= 0;
        i_10_3757 <= 0;
        i_10_3758 <= 0;
        i_10_3759 <= 0;
        i_10_3760 <= 0;
        i_10_3761 <= 0;
        i_10_3762 <= 0;
        i_10_3763 <= 0;
        i_10_3764 <= 0;
        i_10_3765 <= 0;
        i_10_3766 <= 0;
        i_10_3767 <= 0;
        i_10_3768 <= 0;
        i_10_3769 <= 0;
        i_10_3770 <= 0;
        i_10_3771 <= 0;
        i_10_3772 <= 0;
        i_10_3773 <= 0;
        i_10_3774 <= 0;
        i_10_3775 <= 0;
        i_10_3776 <= 0;
        i_10_3777 <= 0;
        i_10_3778 <= 0;
        i_10_3779 <= 0;
        i_10_3780 <= 0;
        i_10_3781 <= 0;
        i_10_3782 <= 0;
        i_10_3783 <= 0;
        i_10_3784 <= 0;
        i_10_3785 <= 0;
        i_10_3786 <= 0;
        i_10_3787 <= 0;
        i_10_3788 <= 0;
        i_10_3789 <= 0;
        i_10_3790 <= 0;
        i_10_3791 <= 0;
        i_10_3792 <= 0;
        i_10_3793 <= 0;
        i_10_3794 <= 0;
        i_10_3795 <= 0;
        i_10_3796 <= 0;
        i_10_3797 <= 0;
        i_10_3798 <= 0;
        i_10_3799 <= 0;
        i_10_3800 <= 0;
        i_10_3801 <= 0;
        i_10_3802 <= 0;
        i_10_3803 <= 0;
        i_10_3804 <= 0;
        i_10_3805 <= 0;
        i_10_3806 <= 0;
        i_10_3807 <= 0;
        i_10_3808 <= 0;
        i_10_3809 <= 0;
        i_10_3810 <= 0;
        i_10_3811 <= 0;
        i_10_3812 <= 0;
        i_10_3813 <= 0;
        i_10_3814 <= 0;
        i_10_3815 <= 0;
        i_10_3816 <= 0;
        i_10_3817 <= 0;
        i_10_3818 <= 0;
        i_10_3819 <= 0;
        i_10_3820 <= 0;
        i_10_3821 <= 0;
        i_10_3822 <= 0;
        i_10_3823 <= 0;
        i_10_3824 <= 0;
        i_10_3825 <= 0;
        i_10_3826 <= 0;
        i_10_3827 <= 0;
        i_10_3828 <= 0;
        i_10_3829 <= 0;
        i_10_3830 <= 0;
        i_10_3831 <= 0;
        i_10_3832 <= 0;
        i_10_3833 <= 0;
        i_10_3834 <= 0;
        i_10_3835 <= 0;
        i_10_3836 <= 0;
        i_10_3837 <= 0;
        i_10_3838 <= 0;
        i_10_3839 <= 0;
        i_10_3840 <= 0;
        i_10_3841 <= 0;
        i_10_3842 <= 0;
        i_10_3843 <= 0;
        i_10_3844 <= 0;
        i_10_3845 <= 0;
        i_10_3846 <= 0;
        i_10_3847 <= 0;
        i_10_3848 <= 0;
        i_10_3849 <= 0;
        i_10_3850 <= 0;
        i_10_3851 <= 0;
        i_10_3852 <= 0;
        i_10_3853 <= 0;
        i_10_3854 <= 0;
        i_10_3855 <= 0;
        i_10_3856 <= 0;
        i_10_3857 <= 0;
        i_10_3858 <= 0;
        i_10_3859 <= 0;
        i_10_3860 <= 0;
        i_10_3861 <= 0;
        i_10_3862 <= 0;
        i_10_3863 <= 0;
        i_10_3864 <= 0;
        i_10_3865 <= 0;
        i_10_3866 <= 0;
        i_10_3867 <= 0;
        i_10_3868 <= 0;
        i_10_3869 <= 0;
        i_10_3870 <= 0;
        i_10_3871 <= 0;
        i_10_3872 <= 0;
        i_10_3873 <= 0;
        i_10_3874 <= 0;
        i_10_3875 <= 0;
        i_10_3876 <= 0;
        i_10_3877 <= 0;
        i_10_3878 <= 0;
        i_10_3879 <= 0;
        i_10_3880 <= 0;
        i_10_3881 <= 0;
        i_10_3882 <= 0;
        i_10_3883 <= 0;
        i_10_3884 <= 0;
        i_10_3885 <= 0;
        i_10_3886 <= 0;
        i_10_3887 <= 0;
        i_10_3888 <= 0;
        i_10_3889 <= 0;
        i_10_3890 <= 0;
        i_10_3891 <= 0;
        i_10_3892 <= 0;
        i_10_3893 <= 0;
        i_10_3894 <= 0;
        i_10_3895 <= 0;
        i_10_3896 <= 0;
        i_10_3897 <= 0;
        i_10_3898 <= 0;
        i_10_3899 <= 0;
        i_10_3900 <= 0;
        i_10_3901 <= 0;
        i_10_3902 <= 0;
        i_10_3903 <= 0;
        i_10_3904 <= 0;
        i_10_3905 <= 0;
        i_10_3906 <= 0;
        i_10_3907 <= 0;
        i_10_3908 <= 0;
        i_10_3909 <= 0;
        i_10_3910 <= 0;
        i_10_3911 <= 0;
        i_10_3912 <= 0;
        i_10_3913 <= 0;
        i_10_3914 <= 0;
        i_10_3915 <= 0;
        i_10_3916 <= 0;
        i_10_3917 <= 0;
        i_10_3918 <= 0;
        i_10_3919 <= 0;
        i_10_3920 <= 0;
        i_10_3921 <= 0;
        i_10_3922 <= 0;
        i_10_3923 <= 0;
        i_10_3924 <= 0;
        i_10_3925 <= 0;
        i_10_3926 <= 0;
        i_10_3927 <= 0;
        i_10_3928 <= 0;
        i_10_3929 <= 0;
        i_10_3930 <= 0;
        i_10_3931 <= 0;
        i_10_3932 <= 0;
        i_10_3933 <= 0;
        i_10_3934 <= 0;
        i_10_3935 <= 0;
        i_10_3936 <= 0;
        i_10_3937 <= 0;
        i_10_3938 <= 0;
        i_10_3939 <= 0;
        i_10_3940 <= 0;
        i_10_3941 <= 0;
        i_10_3942 <= 0;
        i_10_3943 <= 0;
        i_10_3944 <= 0;
        i_10_3945 <= 0;
        i_10_3946 <= 0;
        i_10_3947 <= 0;
        i_10_3948 <= 0;
        i_10_3949 <= 0;
        i_10_3950 <= 0;
        i_10_3951 <= 0;
        i_10_3952 <= 0;
        i_10_3953 <= 0;
        i_10_3954 <= 0;
        i_10_3955 <= 0;
        i_10_3956 <= 0;
        i_10_3957 <= 0;
        i_10_3958 <= 0;
        i_10_3959 <= 0;
        i_10_3960 <= 0;
        i_10_3961 <= 0;
        i_10_3962 <= 0;
        i_10_3963 <= 0;
        i_10_3964 <= 0;
        i_10_3965 <= 0;
        i_10_3966 <= 0;
        i_10_3967 <= 0;
        i_10_3968 <= 0;
        i_10_3969 <= 0;
        i_10_3970 <= 0;
        i_10_3971 <= 0;
        i_10_3972 <= 0;
        i_10_3973 <= 0;
        i_10_3974 <= 0;
        i_10_3975 <= 0;
        i_10_3976 <= 0;
        i_10_3977 <= 0;
        i_10_3978 <= 0;
        i_10_3979 <= 0;
        i_10_3980 <= 0;
        i_10_3981 <= 0;
        i_10_3982 <= 0;
        i_10_3983 <= 0;
        i_10_3984 <= 0;
        i_10_3985 <= 0;
        i_10_3986 <= 0;
        i_10_3987 <= 0;
        i_10_3988 <= 0;
        i_10_3989 <= 0;
        i_10_3990 <= 0;
        i_10_3991 <= 0;
        i_10_3992 <= 0;
        i_10_3993 <= 0;
        i_10_3994 <= 0;
        i_10_3995 <= 0;
        i_10_3996 <= 0;
        i_10_3997 <= 0;
        i_10_3998 <= 0;
        i_10_3999 <= 0;
        i_10_4000 <= 0;
        i_10_4001 <= 0;
        i_10_4002 <= 0;
        i_10_4003 <= 0;
        i_10_4004 <= 0;
        i_10_4005 <= 0;
        i_10_4006 <= 0;
        i_10_4007 <= 0;
        i_10_4008 <= 0;
        i_10_4009 <= 0;
        i_10_4010 <= 0;
        i_10_4011 <= 0;
        i_10_4012 <= 0;
        i_10_4013 <= 0;
        i_10_4014 <= 0;
        i_10_4015 <= 0;
        i_10_4016 <= 0;
        i_10_4017 <= 0;
        i_10_4018 <= 0;
        i_10_4019 <= 0;
        i_10_4020 <= 0;
        i_10_4021 <= 0;
        i_10_4022 <= 0;
        i_10_4023 <= 0;
        i_10_4024 <= 0;
        i_10_4025 <= 0;
        i_10_4026 <= 0;
        i_10_4027 <= 0;
        i_10_4028 <= 0;
        i_10_4029 <= 0;
        i_10_4030 <= 0;
        i_10_4031 <= 0;
        i_10_4032 <= 0;
        i_10_4033 <= 0;
        i_10_4034 <= 0;
        i_10_4035 <= 0;
        i_10_4036 <= 0;
        i_10_4037 <= 0;
        i_10_4038 <= 0;
        i_10_4039 <= 0;
        i_10_4040 <= 0;
        i_10_4041 <= 0;
        i_10_4042 <= 0;
        i_10_4043 <= 0;
        i_10_4044 <= 0;
        i_10_4045 <= 0;
        i_10_4046 <= 0;
        i_10_4047 <= 0;
        i_10_4048 <= 0;
        i_10_4049 <= 0;
        i_10_4050 <= 0;
        i_10_4051 <= 0;
        i_10_4052 <= 0;
        i_10_4053 <= 0;
        i_10_4054 <= 0;
        i_10_4055 <= 0;
        i_10_4056 <= 0;
        i_10_4057 <= 0;
        i_10_4058 <= 0;
        i_10_4059 <= 0;
        i_10_4060 <= 0;
        i_10_4061 <= 0;
        i_10_4062 <= 0;
        i_10_4063 <= 0;
        i_10_4064 <= 0;
        i_10_4065 <= 0;
        i_10_4066 <= 0;
        i_10_4067 <= 0;
        i_10_4068 <= 0;
        i_10_4069 <= 0;
        i_10_4070 <= 0;
        i_10_4071 <= 0;
        i_10_4072 <= 0;
        i_10_4073 <= 0;
        i_10_4074 <= 0;
        i_10_4075 <= 0;
        i_10_4076 <= 0;
        i_10_4077 <= 0;
        i_10_4078 <= 0;
        i_10_4079 <= 0;
        i_10_4080 <= 0;
        i_10_4081 <= 0;
        i_10_4082 <= 0;
        i_10_4083 <= 0;
        i_10_4084 <= 0;
        i_10_4085 <= 0;
        i_10_4086 <= 0;
        i_10_4087 <= 0;
        i_10_4088 <= 0;
        i_10_4089 <= 0;
        i_10_4090 <= 0;
        i_10_4091 <= 0;
        i_10_4092 <= 0;
        i_10_4093 <= 0;
        i_10_4094 <= 0;
        i_10_4095 <= 0;
        i_10_4096 <= 0;
        i_10_4097 <= 0;
        i_10_4098 <= 0;
        i_10_4099 <= 0;
        i_10_4100 <= 0;
        i_10_4101 <= 0;
        i_10_4102 <= 0;
        i_10_4103 <= 0;
        i_10_4104 <= 0;
        i_10_4105 <= 0;
        i_10_4106 <= 0;
        i_10_4107 <= 0;
        i_10_4108 <= 0;
        i_10_4109 <= 0;
        i_10_4110 <= 0;
        i_10_4111 <= 0;
        i_10_4112 <= 0;
        i_10_4113 <= 0;
        i_10_4114 <= 0;
        i_10_4115 <= 0;
        i_10_4116 <= 0;
        i_10_4117 <= 0;
        i_10_4118 <= 0;
        i_10_4119 <= 0;
        i_10_4120 <= 0;
        i_10_4121 <= 0;
        i_10_4122 <= 0;
        i_10_4123 <= 0;
        i_10_4124 <= 0;
        i_10_4125 <= 0;
        i_10_4126 <= 0;
        i_10_4127 <= 0;
        i_10_4128 <= 0;
        i_10_4129 <= 0;
        i_10_4130 <= 0;
        i_10_4131 <= 0;
        i_10_4132 <= 0;
        i_10_4133 <= 0;
        i_10_4134 <= 0;
        i_10_4135 <= 0;
        i_10_4136 <= 0;
        i_10_4137 <= 0;
        i_10_4138 <= 0;
        i_10_4139 <= 0;
        i_10_4140 <= 0;
        i_10_4141 <= 0;
        i_10_4142 <= 0;
        i_10_4143 <= 0;
        i_10_4144 <= 0;
        i_10_4145 <= 0;
        i_10_4146 <= 0;
        i_10_4147 <= 0;
        i_10_4148 <= 0;
        i_10_4149 <= 0;
        i_10_4150 <= 0;
        i_10_4151 <= 0;
        i_10_4152 <= 0;
        i_10_4153 <= 0;
        i_10_4154 <= 0;
        i_10_4155 <= 0;
        i_10_4156 <= 0;
        i_10_4157 <= 0;
        i_10_4158 <= 0;
        i_10_4159 <= 0;
        i_10_4160 <= 0;
        i_10_4161 <= 0;
        i_10_4162 <= 0;
        i_10_4163 <= 0;
        i_10_4164 <= 0;
        i_10_4165 <= 0;
        i_10_4166 <= 0;
        i_10_4167 <= 0;
        i_10_4168 <= 0;
        i_10_4169 <= 0;
        i_10_4170 <= 0;
        i_10_4171 <= 0;
        i_10_4172 <= 0;
        i_10_4173 <= 0;
        i_10_4174 <= 0;
        i_10_4175 <= 0;
        i_10_4176 <= 0;
        i_10_4177 <= 0;
        i_10_4178 <= 0;
        i_10_4179 <= 0;
        i_10_4180 <= 0;
        i_10_4181 <= 0;
        i_10_4182 <= 0;
        i_10_4183 <= 0;
        i_10_4184 <= 0;
        i_10_4185 <= 0;
        i_10_4186 <= 0;
        i_10_4187 <= 0;
        i_10_4188 <= 0;
        i_10_4189 <= 0;
        i_10_4190 <= 0;
        i_10_4191 <= 0;
        i_10_4192 <= 0;
        i_10_4193 <= 0;
        i_10_4194 <= 0;
        i_10_4195 <= 0;
        i_10_4196 <= 0;
        i_10_4197 <= 0;
        i_10_4198 <= 0;
        i_10_4199 <= 0;
        i_10_4200 <= 0;
        i_10_4201 <= 0;
        i_10_4202 <= 0;
        i_10_4203 <= 0;
        i_10_4204 <= 0;
        i_10_4205 <= 0;
        i_10_4206 <= 0;
        i_10_4207 <= 0;
        i_10_4208 <= 0;
        i_10_4209 <= 0;
        i_10_4210 <= 0;
        i_10_4211 <= 0;
        i_10_4212 <= 0;
        i_10_4213 <= 0;
        i_10_4214 <= 0;
        i_10_4215 <= 0;
        i_10_4216 <= 0;
        i_10_4217 <= 0;
        i_10_4218 <= 0;
        i_10_4219 <= 0;
        i_10_4220 <= 0;
        i_10_4221 <= 0;
        i_10_4222 <= 0;
        i_10_4223 <= 0;
        i_10_4224 <= 0;
        i_10_4225 <= 0;
        i_10_4226 <= 0;
        i_10_4227 <= 0;
        i_10_4228 <= 0;
        i_10_4229 <= 0;
        i_10_4230 <= 0;
        i_10_4231 <= 0;
        i_10_4232 <= 0;
        i_10_4233 <= 0;
        i_10_4234 <= 0;
        i_10_4235 <= 0;
        i_10_4236 <= 0;
        i_10_4237 <= 0;
        i_10_4238 <= 0;
        i_10_4239 <= 0;
        i_10_4240 <= 0;
        i_10_4241 <= 0;
        i_10_4242 <= 0;
        i_10_4243 <= 0;
        i_10_4244 <= 0;
        i_10_4245 <= 0;
        i_10_4246 <= 0;
        i_10_4247 <= 0;
        i_10_4248 <= 0;
        i_10_4249 <= 0;
        i_10_4250 <= 0;
        i_10_4251 <= 0;
        i_10_4252 <= 0;
        i_10_4253 <= 0;
        i_10_4254 <= 0;
        i_10_4255 <= 0;
        i_10_4256 <= 0;
        i_10_4257 <= 0;
        i_10_4258 <= 0;
        i_10_4259 <= 0;
        i_10_4260 <= 0;
        i_10_4261 <= 0;
        i_10_4262 <= 0;
        i_10_4263 <= 0;
        i_10_4264 <= 0;
        i_10_4265 <= 0;
        i_10_4266 <= 0;
        i_10_4267 <= 0;
        i_10_4268 <= 0;
        i_10_4269 <= 0;
        i_10_4270 <= 0;
        i_10_4271 <= 0;
        i_10_4272 <= 0;
        i_10_4273 <= 0;
        i_10_4274 <= 0;
        i_10_4275 <= 0;
        i_10_4276 <= 0;
        i_10_4277 <= 0;
        i_10_4278 <= 0;
        i_10_4279 <= 0;
        i_10_4280 <= 0;
        i_10_4281 <= 0;
        i_10_4282 <= 0;
        i_10_4283 <= 0;
        i_10_4284 <= 0;
        i_10_4285 <= 0;
        i_10_4286 <= 0;
        i_10_4287 <= 0;
        i_10_4288 <= 0;
        i_10_4289 <= 0;
        i_10_4290 <= 0;
        i_10_4291 <= 0;
        i_10_4292 <= 0;
        i_10_4293 <= 0;
        i_10_4294 <= 0;
        i_10_4295 <= 0;
        i_10_4296 <= 0;
        i_10_4297 <= 0;
        i_10_4298 <= 0;
        i_10_4299 <= 0;
        i_10_4300 <= 0;
        i_10_4301 <= 0;
        i_10_4302 <= 0;
        i_10_4303 <= 0;
        i_10_4304 <= 0;
        i_10_4305 <= 0;
        i_10_4306 <= 0;
        i_10_4307 <= 0;
        i_10_4308 <= 0;
        i_10_4309 <= 0;
        i_10_4310 <= 0;
        i_10_4311 <= 0;
        i_10_4312 <= 0;
        i_10_4313 <= 0;
        i_10_4314 <= 0;
        i_10_4315 <= 0;
        i_10_4316 <= 0;
        i_10_4317 <= 0;
        i_10_4318 <= 0;
        i_10_4319 <= 0;
        i_10_4320 <= 0;
        i_10_4321 <= 0;
        i_10_4322 <= 0;
        i_10_4323 <= 0;
        i_10_4324 <= 0;
        i_10_4325 <= 0;
        i_10_4326 <= 0;
        i_10_4327 <= 0;
        i_10_4328 <= 0;
        i_10_4329 <= 0;
        i_10_4330 <= 0;
        i_10_4331 <= 0;
        i_10_4332 <= 0;
        i_10_4333 <= 0;
        i_10_4334 <= 0;
        i_10_4335 <= 0;
        i_10_4336 <= 0;
        i_10_4337 <= 0;
        i_10_4338 <= 0;
        i_10_4339 <= 0;
        i_10_4340 <= 0;
        i_10_4341 <= 0;
        i_10_4342 <= 0;
        i_10_4343 <= 0;
        i_10_4344 <= 0;
        i_10_4345 <= 0;
        i_10_4346 <= 0;
        i_10_4347 <= 0;
        i_10_4348 <= 0;
        i_10_4349 <= 0;
        i_10_4350 <= 0;
        i_10_4351 <= 0;
        i_10_4352 <= 0;
        i_10_4353 <= 0;
        i_10_4354 <= 0;
        i_10_4355 <= 0;
        i_10_4356 <= 0;
        i_10_4357 <= 0;
        i_10_4358 <= 0;
        i_10_4359 <= 0;
        i_10_4360 <= 0;
        i_10_4361 <= 0;
        i_10_4362 <= 0;
        i_10_4363 <= 0;
        i_10_4364 <= 0;
        i_10_4365 <= 0;
        i_10_4366 <= 0;
        i_10_4367 <= 0;
        i_10_4368 <= 0;
        i_10_4369 <= 0;
        i_10_4370 <= 0;
        i_10_4371 <= 0;
        i_10_4372 <= 0;
        i_10_4373 <= 0;
        i_10_4374 <= 0;
        i_10_4375 <= 0;
        i_10_4376 <= 0;
        i_10_4377 <= 0;
        i_10_4378 <= 0;
        i_10_4379 <= 0;
        i_10_4380 <= 0;
        i_10_4381 <= 0;
        i_10_4382 <= 0;
        i_10_4383 <= 0;
        i_10_4384 <= 0;
        i_10_4385 <= 0;
        i_10_4386 <= 0;
        i_10_4387 <= 0;
        i_10_4388 <= 0;
        i_10_4389 <= 0;
        i_10_4390 <= 0;
        i_10_4391 <= 0;
        i_10_4392 <= 0;
        i_10_4393 <= 0;
        i_10_4394 <= 0;
        i_10_4395 <= 0;
        i_10_4396 <= 0;
        i_10_4397 <= 0;
        i_10_4398 <= 0;
        i_10_4399 <= 0;
        i_10_4400 <= 0;
        i_10_4401 <= 0;
        i_10_4402 <= 0;
        i_10_4403 <= 0;
        i_10_4404 <= 0;
        i_10_4405 <= 0;
        i_10_4406 <= 0;
        i_10_4407 <= 0;
        i_10_4408 <= 0;
        i_10_4409 <= 0;
        i_10_4410 <= 0;
        i_10_4411 <= 0;
        i_10_4412 <= 0;
        i_10_4413 <= 0;
        i_10_4414 <= 0;
        i_10_4415 <= 0;
        i_10_4416 <= 0;
        i_10_4417 <= 0;
        i_10_4418 <= 0;
        i_10_4419 <= 0;
        i_10_4420 <= 0;
        i_10_4421 <= 0;
        i_10_4422 <= 0;
        i_10_4423 <= 0;
        i_10_4424 <= 0;
        i_10_4425 <= 0;
        i_10_4426 <= 0;
        i_10_4427 <= 0;
        i_10_4428 <= 0;
        i_10_4429 <= 0;
        i_10_4430 <= 0;
        i_10_4431 <= 0;
        i_10_4432 <= 0;
        i_10_4433 <= 0;
        i_10_4434 <= 0;
        i_10_4435 <= 0;
        i_10_4436 <= 0;
        i_10_4437 <= 0;
        i_10_4438 <= 0;
        i_10_4439 <= 0;
        i_10_4440 <= 0;
        i_10_4441 <= 0;
        i_10_4442 <= 0;
        i_10_4443 <= 0;
        i_10_4444 <= 0;
        i_10_4445 <= 0;
        i_10_4446 <= 0;
        i_10_4447 <= 0;
        i_10_4448 <= 0;
        i_10_4449 <= 0;
        i_10_4450 <= 0;
        i_10_4451 <= 0;
        i_10_4452 <= 0;
        i_10_4453 <= 0;
        i_10_4454 <= 0;
        i_10_4455 <= 0;
        i_10_4456 <= 0;
        i_10_4457 <= 0;
        i_10_4458 <= 0;
        i_10_4459 <= 0;
        i_10_4460 <= 0;
        i_10_4461 <= 0;
        i_10_4462 <= 0;
        i_10_4463 <= 0;
        i_10_4464 <= 0;
        i_10_4465 <= 0;
        i_10_4466 <= 0;
        i_10_4467 <= 0;
        i_10_4468 <= 0;
        i_10_4469 <= 0;
        i_10_4470 <= 0;
        i_10_4471 <= 0;
        i_10_4472 <= 0;
        i_10_4473 <= 0;
        i_10_4474 <= 0;
        i_10_4475 <= 0;
        i_10_4476 <= 0;
        i_10_4477 <= 0;
        i_10_4478 <= 0;
        i_10_4479 <= 0;
        i_10_4480 <= 0;
        i_10_4481 <= 0;
        i_10_4482 <= 0;
        i_10_4483 <= 0;
        i_10_4484 <= 0;
        i_10_4485 <= 0;
        i_10_4486 <= 0;
        i_10_4487 <= 0;
        i_10_4488 <= 0;
        i_10_4489 <= 0;
        i_10_4490 <= 0;
        i_10_4491 <= 0;
        i_10_4492 <= 0;
        i_10_4493 <= 0;
        i_10_4494 <= 0;
        i_10_4495 <= 0;
        i_10_4496 <= 0;
        i_10_4497 <= 0;
        i_10_4498 <= 0;
        i_10_4499 <= 0;
        i_10_4500 <= 0;
        i_10_4501 <= 0;
        i_10_4502 <= 0;
        i_10_4503 <= 0;
        i_10_4504 <= 0;
        i_10_4505 <= 0;
        i_10_4506 <= 0;
        i_10_4507 <= 0;
        i_10_4508 <= 0;
        i_10_4509 <= 0;
        i_10_4510 <= 0;
        i_10_4511 <= 0;
        i_10_4512 <= 0;
        i_10_4513 <= 0;
        i_10_4514 <= 0;
        i_10_4515 <= 0;
        i_10_4516 <= 0;
        i_10_4517 <= 0;
        i_10_4518 <= 0;
        i_10_4519 <= 0;
        i_10_4520 <= 0;
        i_10_4521 <= 0;
        i_10_4522 <= 0;
        i_10_4523 <= 0;
        i_10_4524 <= 0;
        i_10_4525 <= 0;
        i_10_4526 <= 0;
        i_10_4527 <= 0;
        i_10_4528 <= 0;
        i_10_4529 <= 0;
        i_10_4530 <= 0;
        i_10_4531 <= 0;
        i_10_4532 <= 0;
        i_10_4533 <= 0;
        i_10_4534 <= 0;
        i_10_4535 <= 0;
        i_10_4536 <= 0;
        i_10_4537 <= 0;
        i_10_4538 <= 0;
        i_10_4539 <= 0;
        i_10_4540 <= 0;
        i_10_4541 <= 0;
        i_10_4542 <= 0;
        i_10_4543 <= 0;
        i_10_4544 <= 0;
        i_10_4545 <= 0;
        i_10_4546 <= 0;
        i_10_4547 <= 0;
        i_10_4548 <= 0;
        i_10_4549 <= 0;
        i_10_4550 <= 0;
        i_10_4551 <= 0;
        i_10_4552 <= 0;
        i_10_4553 <= 0;
        i_10_4554 <= 0;
        i_10_4555 <= 0;
        i_10_4556 <= 0;
        i_10_4557 <= 0;
        i_10_4558 <= 0;
        i_10_4559 <= 0;
        i_10_4560 <= 0;
        i_10_4561 <= 0;
        i_10_4562 <= 0;
        i_10_4563 <= 0;
        i_10_4564 <= 0;
        i_10_4565 <= 0;
        i_10_4566 <= 0;
        i_10_4567 <= 0;
        i_10_4568 <= 0;
        i_10_4569 <= 0;
        i_10_4570 <= 0;
        i_10_4571 <= 0;
        i_10_4572 <= 0;
        i_10_4573 <= 0;
        i_10_4574 <= 0;
        i_10_4575 <= 0;
        i_10_4576 <= 0;
        i_10_4577 <= 0;
        i_10_4578 <= 0;
        i_10_4579 <= 0;
        i_10_4580 <= 0;
        i_10_4581 <= 0;
        i_10_4582 <= 0;
        i_10_4583 <= 0;
        i_10_4584 <= 0;
        i_10_4585 <= 0;
        i_10_4586 <= 0;
        i_10_4587 <= 0;
        i_10_4588 <= 0;
        i_10_4589 <= 0;
        i_10_4590 <= 0;
        i_10_4591 <= 0;
        i_10_4592 <= 0;
        i_10_4593 <= 0;
        i_10_4594 <= 0;
        i_10_4595 <= 0;
        i_10_4596 <= 0;
        i_10_4597 <= 0;
        i_10_4598 <= 0;
        i_10_4599 <= 0;
        i_10_4600 <= 0;
        i_10_4601 <= 0;
        i_10_4602 <= 0;
        i_10_4603 <= 0;
        i_10_4604 <= 0;
        i_10_4605 <= 0;
        i_10_4606 <= 0;
        i_10_4607 <= 0;
        dly1 <= 0;
        dly2 <= 0;
      end
    else if (ce)
      begin
        out_reg <= { o_10_511, o_10_510, o_10_509, o_10_508, o_10_507, o_10_506, o_10_505, o_10_504, o_10_503, o_10_502, o_10_501, o_10_500, o_10_499, o_10_498, o_10_497, o_10_496, o_10_495, o_10_494, o_10_493, o_10_492, o_10_491, o_10_490, o_10_489, o_10_488, o_10_487, o_10_486, o_10_485, o_10_484, o_10_483, o_10_482, o_10_481, o_10_480, o_10_479, o_10_478, o_10_477, o_10_476, o_10_475, o_10_474, o_10_473, o_10_472, o_10_471, o_10_470, o_10_469, o_10_468, o_10_467, o_10_466, o_10_465, o_10_464, o_10_463, o_10_462, o_10_461, o_10_460, o_10_459, o_10_458, o_10_457, o_10_456, o_10_455, o_10_454, o_10_453, o_10_452, o_10_451, o_10_450, o_10_449, o_10_448, o_10_447, o_10_446, o_10_445, o_10_444, o_10_443, o_10_442, o_10_441, o_10_440, o_10_439, o_10_438, o_10_437, o_10_436, o_10_435, o_10_434, o_10_433, o_10_432, o_10_431, o_10_430, o_10_429, o_10_428, o_10_427, o_10_426, o_10_425, o_10_424, o_10_423, o_10_422, o_10_421, o_10_420, o_10_419, o_10_418, o_10_417, o_10_416, o_10_415, o_10_414, o_10_413, o_10_412, o_10_411, o_10_410, o_10_409, o_10_408, o_10_407, o_10_406, o_10_405, o_10_404, o_10_403, o_10_402, o_10_401, o_10_400, o_10_399, o_10_398, o_10_397, o_10_396, o_10_395, o_10_394, o_10_393, o_10_392, o_10_391, o_10_390, o_10_389, o_10_388, o_10_387, o_10_386, o_10_385, o_10_384, o_10_383, o_10_382, o_10_381, o_10_380, o_10_379, o_10_378, o_10_377, o_10_376, o_10_375, o_10_374, o_10_373, o_10_372, o_10_371, o_10_370, o_10_369, o_10_368, o_10_367, o_10_366, o_10_365, o_10_364, o_10_363, o_10_362, o_10_361, o_10_360, o_10_359, o_10_358, o_10_357, o_10_356, o_10_355, o_10_354, o_10_353, o_10_352, o_10_351, o_10_350, o_10_349, o_10_348, o_10_347, o_10_346, o_10_345, o_10_344, o_10_343, o_10_342, o_10_341, o_10_340, o_10_339, o_10_338, o_10_337, o_10_336, o_10_335, o_10_334, o_10_333, o_10_332, o_10_331, o_10_330, o_10_329, o_10_328, o_10_327, o_10_326, o_10_325, o_10_324, o_10_323, o_10_322, o_10_321, o_10_320, o_10_319, o_10_318, o_10_317, o_10_316, o_10_315, o_10_314, o_10_313, o_10_312, o_10_311, o_10_310, o_10_309, o_10_308, o_10_307, o_10_306, o_10_305, o_10_304, o_10_303, o_10_302, o_10_301, o_10_300, o_10_299, o_10_298, o_10_297, o_10_296, o_10_295, o_10_294, o_10_293, o_10_292, o_10_291, o_10_290, o_10_289, o_10_288, o_10_287, o_10_286, o_10_285, o_10_284, o_10_283, o_10_282, o_10_281, o_10_280, o_10_279, o_10_278, o_10_277, o_10_276, o_10_275, o_10_274, o_10_273, o_10_272, o_10_271, o_10_270, o_10_269, o_10_268, o_10_267, o_10_266, o_10_265, o_10_264, o_10_263, o_10_262, o_10_261, o_10_260, o_10_259, o_10_258, o_10_257, o_10_256, o_10_255, o_10_254, o_10_253, o_10_252, o_10_251, o_10_250, o_10_249, o_10_248, o_10_247, o_10_246, o_10_245, o_10_244, o_10_243, o_10_242, o_10_241, o_10_240, o_10_239, o_10_238, o_10_237, o_10_236, o_10_235, o_10_234, o_10_233, o_10_232, o_10_231, o_10_230, o_10_229, o_10_228, o_10_227, o_10_226, o_10_225, o_10_224, o_10_223, o_10_222, o_10_221, o_10_220, o_10_219, o_10_218, o_10_217, o_10_216, o_10_215, o_10_214, o_10_213, o_10_212, o_10_211, o_10_210, o_10_209, o_10_208, o_10_207, o_10_206, o_10_205, o_10_204, o_10_203, o_10_202, o_10_201, o_10_200, o_10_199, o_10_198, o_10_197, o_10_196, o_10_195, o_10_194, o_10_193, o_10_192, o_10_191, o_10_190, o_10_189, o_10_188, o_10_187, o_10_186, o_10_185, o_10_184, o_10_183, o_10_182, o_10_181, o_10_180, o_10_179, o_10_178, o_10_177, o_10_176, o_10_175, o_10_174, o_10_173, o_10_172, o_10_171, o_10_170, o_10_169, o_10_168, o_10_167, o_10_166, o_10_165, o_10_164, o_10_163, o_10_162, o_10_161, o_10_160, o_10_159, o_10_158, o_10_157, o_10_156, o_10_155, o_10_154, o_10_153, o_10_152, o_10_151, o_10_150, o_10_149, o_10_148, o_10_147, o_10_146, o_10_145, o_10_144, o_10_143, o_10_142, o_10_141, o_10_140, o_10_139, o_10_138, o_10_137, o_10_136, o_10_135, o_10_134, o_10_133, o_10_132, o_10_131, o_10_130, o_10_129, o_10_128, o_10_127, o_10_126, o_10_125, o_10_124, o_10_123, o_10_122, o_10_121, o_10_120, o_10_119, o_10_118, o_10_117, o_10_116, o_10_115, o_10_114, o_10_113, o_10_112, o_10_111, o_10_110, o_10_109, o_10_108, o_10_107, o_10_106, o_10_105, o_10_104, o_10_103, o_10_102, o_10_101, o_10_100, o_10_99, o_10_98, o_10_97, o_10_96, o_10_95, o_10_94, o_10_93, o_10_92, o_10_91, o_10_90, o_10_89, o_10_88, o_10_87, o_10_86, o_10_85, o_10_84, o_10_83, o_10_82, o_10_81, o_10_80, o_10_79, o_10_78, o_10_77, o_10_76, o_10_75, o_10_74, o_10_73, o_10_72, o_10_71, o_10_70, o_10_69, o_10_68, o_10_67, o_10_66, o_10_65, o_10_64, o_10_63, o_10_62, o_10_61, o_10_60, o_10_59, o_10_58, o_10_57, o_10_56, o_10_55, o_10_54, o_10_53, o_10_52, o_10_51, o_10_50, o_10_49, o_10_48, o_10_47, o_10_46, o_10_45, o_10_44, o_10_43, o_10_42, o_10_41, o_10_40, o_10_39, o_10_38, o_10_37, o_10_36, o_10_35, o_10_34, o_10_33, o_10_32, o_10_31, o_10_30, o_10_29, o_10_28, o_10_27, o_10_26, o_10_25, o_10_24, o_10_23, o_10_22, o_10_21, o_10_20, o_10_19, o_10_18, o_10_17, o_10_16, o_10_15, o_10_14, o_10_13, o_10_12, o_10_11, o_10_10, o_10_9, o_10_8, o_10_7, o_10_6, o_10_5, o_10_4, o_10_3, o_10_2, o_10_1, o_10_0};
        i_10_0 <= in_reg[0];
        i_10_1 <= in_reg[512];
        i_10_2 <= in_reg[1024];
        i_10_3 <= in_reg[1536];
        i_10_4 <= in_reg[2048];
        i_10_5 <= in_reg[2560];
        i_10_6 <= in_reg[3072];
        i_10_7 <= in_reg[3584];
        i_10_8 <= in_reg[4096];
        i_10_9 <= in_reg[1];
        i_10_10 <= in_reg[513];
        i_10_11 <= in_reg[1025];
        i_10_12 <= in_reg[1537];
        i_10_13 <= in_reg[2049];
        i_10_14 <= in_reg[2561];
        i_10_15 <= in_reg[3073];
        i_10_16 <= in_reg[3585];
        i_10_17 <= in_reg[4097];
        i_10_18 <= in_reg[2];
        i_10_19 <= in_reg[514];
        i_10_20 <= in_reg[1026];
        i_10_21 <= in_reg[1538];
        i_10_22 <= in_reg[2050];
        i_10_23 <= in_reg[2562];
        i_10_24 <= in_reg[3074];
        i_10_25 <= in_reg[3586];
        i_10_26 <= in_reg[4098];
        i_10_27 <= in_reg[3];
        i_10_28 <= in_reg[515];
        i_10_29 <= in_reg[1027];
        i_10_30 <= in_reg[1539];
        i_10_31 <= in_reg[2051];
        i_10_32 <= in_reg[2563];
        i_10_33 <= in_reg[3075];
        i_10_34 <= in_reg[3587];
        i_10_35 <= in_reg[4099];
        i_10_36 <= in_reg[4];
        i_10_37 <= in_reg[516];
        i_10_38 <= in_reg[1028];
        i_10_39 <= in_reg[1540];
        i_10_40 <= in_reg[2052];
        i_10_41 <= in_reg[2564];
        i_10_42 <= in_reg[3076];
        i_10_43 <= in_reg[3588];
        i_10_44 <= in_reg[4100];
        i_10_45 <= in_reg[5];
        i_10_46 <= in_reg[517];
        i_10_47 <= in_reg[1029];
        i_10_48 <= in_reg[1541];
        i_10_49 <= in_reg[2053];
        i_10_50 <= in_reg[2565];
        i_10_51 <= in_reg[3077];
        i_10_52 <= in_reg[3589];
        i_10_53 <= in_reg[4101];
        i_10_54 <= in_reg[6];
        i_10_55 <= in_reg[518];
        i_10_56 <= in_reg[1030];
        i_10_57 <= in_reg[1542];
        i_10_58 <= in_reg[2054];
        i_10_59 <= in_reg[2566];
        i_10_60 <= in_reg[3078];
        i_10_61 <= in_reg[3590];
        i_10_62 <= in_reg[4102];
        i_10_63 <= in_reg[7];
        i_10_64 <= in_reg[519];
        i_10_65 <= in_reg[1031];
        i_10_66 <= in_reg[1543];
        i_10_67 <= in_reg[2055];
        i_10_68 <= in_reg[2567];
        i_10_69 <= in_reg[3079];
        i_10_70 <= in_reg[3591];
        i_10_71 <= in_reg[4103];
        i_10_72 <= in_reg[8];
        i_10_73 <= in_reg[520];
        i_10_74 <= in_reg[1032];
        i_10_75 <= in_reg[1544];
        i_10_76 <= in_reg[2056];
        i_10_77 <= in_reg[2568];
        i_10_78 <= in_reg[3080];
        i_10_79 <= in_reg[3592];
        i_10_80 <= in_reg[4104];
        i_10_81 <= in_reg[9];
        i_10_82 <= in_reg[521];
        i_10_83 <= in_reg[1033];
        i_10_84 <= in_reg[1545];
        i_10_85 <= in_reg[2057];
        i_10_86 <= in_reg[2569];
        i_10_87 <= in_reg[3081];
        i_10_88 <= in_reg[3593];
        i_10_89 <= in_reg[4105];
        i_10_90 <= in_reg[10];
        i_10_91 <= in_reg[522];
        i_10_92 <= in_reg[1034];
        i_10_93 <= in_reg[1546];
        i_10_94 <= in_reg[2058];
        i_10_95 <= in_reg[2570];
        i_10_96 <= in_reg[3082];
        i_10_97 <= in_reg[3594];
        i_10_98 <= in_reg[4106];
        i_10_99 <= in_reg[11];
        i_10_100 <= in_reg[523];
        i_10_101 <= in_reg[1035];
        i_10_102 <= in_reg[1547];
        i_10_103 <= in_reg[2059];
        i_10_104 <= in_reg[2571];
        i_10_105 <= in_reg[3083];
        i_10_106 <= in_reg[3595];
        i_10_107 <= in_reg[4107];
        i_10_108 <= in_reg[12];
        i_10_109 <= in_reg[524];
        i_10_110 <= in_reg[1036];
        i_10_111 <= in_reg[1548];
        i_10_112 <= in_reg[2060];
        i_10_113 <= in_reg[2572];
        i_10_114 <= in_reg[3084];
        i_10_115 <= in_reg[3596];
        i_10_116 <= in_reg[4108];
        i_10_117 <= in_reg[13];
        i_10_118 <= in_reg[525];
        i_10_119 <= in_reg[1037];
        i_10_120 <= in_reg[1549];
        i_10_121 <= in_reg[2061];
        i_10_122 <= in_reg[2573];
        i_10_123 <= in_reg[3085];
        i_10_124 <= in_reg[3597];
        i_10_125 <= in_reg[4109];
        i_10_126 <= in_reg[14];
        i_10_127 <= in_reg[526];
        i_10_128 <= in_reg[1038];
        i_10_129 <= in_reg[1550];
        i_10_130 <= in_reg[2062];
        i_10_131 <= in_reg[2574];
        i_10_132 <= in_reg[3086];
        i_10_133 <= in_reg[3598];
        i_10_134 <= in_reg[4110];
        i_10_135 <= in_reg[15];
        i_10_136 <= in_reg[527];
        i_10_137 <= in_reg[1039];
        i_10_138 <= in_reg[1551];
        i_10_139 <= in_reg[2063];
        i_10_140 <= in_reg[2575];
        i_10_141 <= in_reg[3087];
        i_10_142 <= in_reg[3599];
        i_10_143 <= in_reg[4111];
        i_10_144 <= in_reg[16];
        i_10_145 <= in_reg[528];
        i_10_146 <= in_reg[1040];
        i_10_147 <= in_reg[1552];
        i_10_148 <= in_reg[2064];
        i_10_149 <= in_reg[2576];
        i_10_150 <= in_reg[3088];
        i_10_151 <= in_reg[3600];
        i_10_152 <= in_reg[4112];
        i_10_153 <= in_reg[17];
        i_10_154 <= in_reg[529];
        i_10_155 <= in_reg[1041];
        i_10_156 <= in_reg[1553];
        i_10_157 <= in_reg[2065];
        i_10_158 <= in_reg[2577];
        i_10_159 <= in_reg[3089];
        i_10_160 <= in_reg[3601];
        i_10_161 <= in_reg[4113];
        i_10_162 <= in_reg[18];
        i_10_163 <= in_reg[530];
        i_10_164 <= in_reg[1042];
        i_10_165 <= in_reg[1554];
        i_10_166 <= in_reg[2066];
        i_10_167 <= in_reg[2578];
        i_10_168 <= in_reg[3090];
        i_10_169 <= in_reg[3602];
        i_10_170 <= in_reg[4114];
        i_10_171 <= in_reg[19];
        i_10_172 <= in_reg[531];
        i_10_173 <= in_reg[1043];
        i_10_174 <= in_reg[1555];
        i_10_175 <= in_reg[2067];
        i_10_176 <= in_reg[2579];
        i_10_177 <= in_reg[3091];
        i_10_178 <= in_reg[3603];
        i_10_179 <= in_reg[4115];
        i_10_180 <= in_reg[20];
        i_10_181 <= in_reg[532];
        i_10_182 <= in_reg[1044];
        i_10_183 <= in_reg[1556];
        i_10_184 <= in_reg[2068];
        i_10_185 <= in_reg[2580];
        i_10_186 <= in_reg[3092];
        i_10_187 <= in_reg[3604];
        i_10_188 <= in_reg[4116];
        i_10_189 <= in_reg[21];
        i_10_190 <= in_reg[533];
        i_10_191 <= in_reg[1045];
        i_10_192 <= in_reg[1557];
        i_10_193 <= in_reg[2069];
        i_10_194 <= in_reg[2581];
        i_10_195 <= in_reg[3093];
        i_10_196 <= in_reg[3605];
        i_10_197 <= in_reg[4117];
        i_10_198 <= in_reg[22];
        i_10_199 <= in_reg[534];
        i_10_200 <= in_reg[1046];
        i_10_201 <= in_reg[1558];
        i_10_202 <= in_reg[2070];
        i_10_203 <= in_reg[2582];
        i_10_204 <= in_reg[3094];
        i_10_205 <= in_reg[3606];
        i_10_206 <= in_reg[4118];
        i_10_207 <= in_reg[23];
        i_10_208 <= in_reg[535];
        i_10_209 <= in_reg[1047];
        i_10_210 <= in_reg[1559];
        i_10_211 <= in_reg[2071];
        i_10_212 <= in_reg[2583];
        i_10_213 <= in_reg[3095];
        i_10_214 <= in_reg[3607];
        i_10_215 <= in_reg[4119];
        i_10_216 <= in_reg[24];
        i_10_217 <= in_reg[536];
        i_10_218 <= in_reg[1048];
        i_10_219 <= in_reg[1560];
        i_10_220 <= in_reg[2072];
        i_10_221 <= in_reg[2584];
        i_10_222 <= in_reg[3096];
        i_10_223 <= in_reg[3608];
        i_10_224 <= in_reg[4120];
        i_10_225 <= in_reg[25];
        i_10_226 <= in_reg[537];
        i_10_227 <= in_reg[1049];
        i_10_228 <= in_reg[1561];
        i_10_229 <= in_reg[2073];
        i_10_230 <= in_reg[2585];
        i_10_231 <= in_reg[3097];
        i_10_232 <= in_reg[3609];
        i_10_233 <= in_reg[4121];
        i_10_234 <= in_reg[26];
        i_10_235 <= in_reg[538];
        i_10_236 <= in_reg[1050];
        i_10_237 <= in_reg[1562];
        i_10_238 <= in_reg[2074];
        i_10_239 <= in_reg[2586];
        i_10_240 <= in_reg[3098];
        i_10_241 <= in_reg[3610];
        i_10_242 <= in_reg[4122];
        i_10_243 <= in_reg[27];
        i_10_244 <= in_reg[539];
        i_10_245 <= in_reg[1051];
        i_10_246 <= in_reg[1563];
        i_10_247 <= in_reg[2075];
        i_10_248 <= in_reg[2587];
        i_10_249 <= in_reg[3099];
        i_10_250 <= in_reg[3611];
        i_10_251 <= in_reg[4123];
        i_10_252 <= in_reg[28];
        i_10_253 <= in_reg[540];
        i_10_254 <= in_reg[1052];
        i_10_255 <= in_reg[1564];
        i_10_256 <= in_reg[2076];
        i_10_257 <= in_reg[2588];
        i_10_258 <= in_reg[3100];
        i_10_259 <= in_reg[3612];
        i_10_260 <= in_reg[4124];
        i_10_261 <= in_reg[29];
        i_10_262 <= in_reg[541];
        i_10_263 <= in_reg[1053];
        i_10_264 <= in_reg[1565];
        i_10_265 <= in_reg[2077];
        i_10_266 <= in_reg[2589];
        i_10_267 <= in_reg[3101];
        i_10_268 <= in_reg[3613];
        i_10_269 <= in_reg[4125];
        i_10_270 <= in_reg[30];
        i_10_271 <= in_reg[542];
        i_10_272 <= in_reg[1054];
        i_10_273 <= in_reg[1566];
        i_10_274 <= in_reg[2078];
        i_10_275 <= in_reg[2590];
        i_10_276 <= in_reg[3102];
        i_10_277 <= in_reg[3614];
        i_10_278 <= in_reg[4126];
        i_10_279 <= in_reg[31];
        i_10_280 <= in_reg[543];
        i_10_281 <= in_reg[1055];
        i_10_282 <= in_reg[1567];
        i_10_283 <= in_reg[2079];
        i_10_284 <= in_reg[2591];
        i_10_285 <= in_reg[3103];
        i_10_286 <= in_reg[3615];
        i_10_287 <= in_reg[4127];
        i_10_288 <= in_reg[32];
        i_10_289 <= in_reg[544];
        i_10_290 <= in_reg[1056];
        i_10_291 <= in_reg[1568];
        i_10_292 <= in_reg[2080];
        i_10_293 <= in_reg[2592];
        i_10_294 <= in_reg[3104];
        i_10_295 <= in_reg[3616];
        i_10_296 <= in_reg[4128];
        i_10_297 <= in_reg[33];
        i_10_298 <= in_reg[545];
        i_10_299 <= in_reg[1057];
        i_10_300 <= in_reg[1569];
        i_10_301 <= in_reg[2081];
        i_10_302 <= in_reg[2593];
        i_10_303 <= in_reg[3105];
        i_10_304 <= in_reg[3617];
        i_10_305 <= in_reg[4129];
        i_10_306 <= in_reg[34];
        i_10_307 <= in_reg[546];
        i_10_308 <= in_reg[1058];
        i_10_309 <= in_reg[1570];
        i_10_310 <= in_reg[2082];
        i_10_311 <= in_reg[2594];
        i_10_312 <= in_reg[3106];
        i_10_313 <= in_reg[3618];
        i_10_314 <= in_reg[4130];
        i_10_315 <= in_reg[35];
        i_10_316 <= in_reg[547];
        i_10_317 <= in_reg[1059];
        i_10_318 <= in_reg[1571];
        i_10_319 <= in_reg[2083];
        i_10_320 <= in_reg[2595];
        i_10_321 <= in_reg[3107];
        i_10_322 <= in_reg[3619];
        i_10_323 <= in_reg[4131];
        i_10_324 <= in_reg[36];
        i_10_325 <= in_reg[548];
        i_10_326 <= in_reg[1060];
        i_10_327 <= in_reg[1572];
        i_10_328 <= in_reg[2084];
        i_10_329 <= in_reg[2596];
        i_10_330 <= in_reg[3108];
        i_10_331 <= in_reg[3620];
        i_10_332 <= in_reg[4132];
        i_10_333 <= in_reg[37];
        i_10_334 <= in_reg[549];
        i_10_335 <= in_reg[1061];
        i_10_336 <= in_reg[1573];
        i_10_337 <= in_reg[2085];
        i_10_338 <= in_reg[2597];
        i_10_339 <= in_reg[3109];
        i_10_340 <= in_reg[3621];
        i_10_341 <= in_reg[4133];
        i_10_342 <= in_reg[38];
        i_10_343 <= in_reg[550];
        i_10_344 <= in_reg[1062];
        i_10_345 <= in_reg[1574];
        i_10_346 <= in_reg[2086];
        i_10_347 <= in_reg[2598];
        i_10_348 <= in_reg[3110];
        i_10_349 <= in_reg[3622];
        i_10_350 <= in_reg[4134];
        i_10_351 <= in_reg[39];
        i_10_352 <= in_reg[551];
        i_10_353 <= in_reg[1063];
        i_10_354 <= in_reg[1575];
        i_10_355 <= in_reg[2087];
        i_10_356 <= in_reg[2599];
        i_10_357 <= in_reg[3111];
        i_10_358 <= in_reg[3623];
        i_10_359 <= in_reg[4135];
        i_10_360 <= in_reg[40];
        i_10_361 <= in_reg[552];
        i_10_362 <= in_reg[1064];
        i_10_363 <= in_reg[1576];
        i_10_364 <= in_reg[2088];
        i_10_365 <= in_reg[2600];
        i_10_366 <= in_reg[3112];
        i_10_367 <= in_reg[3624];
        i_10_368 <= in_reg[4136];
        i_10_369 <= in_reg[41];
        i_10_370 <= in_reg[553];
        i_10_371 <= in_reg[1065];
        i_10_372 <= in_reg[1577];
        i_10_373 <= in_reg[2089];
        i_10_374 <= in_reg[2601];
        i_10_375 <= in_reg[3113];
        i_10_376 <= in_reg[3625];
        i_10_377 <= in_reg[4137];
        i_10_378 <= in_reg[42];
        i_10_379 <= in_reg[554];
        i_10_380 <= in_reg[1066];
        i_10_381 <= in_reg[1578];
        i_10_382 <= in_reg[2090];
        i_10_383 <= in_reg[2602];
        i_10_384 <= in_reg[3114];
        i_10_385 <= in_reg[3626];
        i_10_386 <= in_reg[4138];
        i_10_387 <= in_reg[43];
        i_10_388 <= in_reg[555];
        i_10_389 <= in_reg[1067];
        i_10_390 <= in_reg[1579];
        i_10_391 <= in_reg[2091];
        i_10_392 <= in_reg[2603];
        i_10_393 <= in_reg[3115];
        i_10_394 <= in_reg[3627];
        i_10_395 <= in_reg[4139];
        i_10_396 <= in_reg[44];
        i_10_397 <= in_reg[556];
        i_10_398 <= in_reg[1068];
        i_10_399 <= in_reg[1580];
        i_10_400 <= in_reg[2092];
        i_10_401 <= in_reg[2604];
        i_10_402 <= in_reg[3116];
        i_10_403 <= in_reg[3628];
        i_10_404 <= in_reg[4140];
        i_10_405 <= in_reg[45];
        i_10_406 <= in_reg[557];
        i_10_407 <= in_reg[1069];
        i_10_408 <= in_reg[1581];
        i_10_409 <= in_reg[2093];
        i_10_410 <= in_reg[2605];
        i_10_411 <= in_reg[3117];
        i_10_412 <= in_reg[3629];
        i_10_413 <= in_reg[4141];
        i_10_414 <= in_reg[46];
        i_10_415 <= in_reg[558];
        i_10_416 <= in_reg[1070];
        i_10_417 <= in_reg[1582];
        i_10_418 <= in_reg[2094];
        i_10_419 <= in_reg[2606];
        i_10_420 <= in_reg[3118];
        i_10_421 <= in_reg[3630];
        i_10_422 <= in_reg[4142];
        i_10_423 <= in_reg[47];
        i_10_424 <= in_reg[559];
        i_10_425 <= in_reg[1071];
        i_10_426 <= in_reg[1583];
        i_10_427 <= in_reg[2095];
        i_10_428 <= in_reg[2607];
        i_10_429 <= in_reg[3119];
        i_10_430 <= in_reg[3631];
        i_10_431 <= in_reg[4143];
        i_10_432 <= in_reg[48];
        i_10_433 <= in_reg[560];
        i_10_434 <= in_reg[1072];
        i_10_435 <= in_reg[1584];
        i_10_436 <= in_reg[2096];
        i_10_437 <= in_reg[2608];
        i_10_438 <= in_reg[3120];
        i_10_439 <= in_reg[3632];
        i_10_440 <= in_reg[4144];
        i_10_441 <= in_reg[49];
        i_10_442 <= in_reg[561];
        i_10_443 <= in_reg[1073];
        i_10_444 <= in_reg[1585];
        i_10_445 <= in_reg[2097];
        i_10_446 <= in_reg[2609];
        i_10_447 <= in_reg[3121];
        i_10_448 <= in_reg[3633];
        i_10_449 <= in_reg[4145];
        i_10_450 <= in_reg[50];
        i_10_451 <= in_reg[562];
        i_10_452 <= in_reg[1074];
        i_10_453 <= in_reg[1586];
        i_10_454 <= in_reg[2098];
        i_10_455 <= in_reg[2610];
        i_10_456 <= in_reg[3122];
        i_10_457 <= in_reg[3634];
        i_10_458 <= in_reg[4146];
        i_10_459 <= in_reg[51];
        i_10_460 <= in_reg[563];
        i_10_461 <= in_reg[1075];
        i_10_462 <= in_reg[1587];
        i_10_463 <= in_reg[2099];
        i_10_464 <= in_reg[2611];
        i_10_465 <= in_reg[3123];
        i_10_466 <= in_reg[3635];
        i_10_467 <= in_reg[4147];
        i_10_468 <= in_reg[52];
        i_10_469 <= in_reg[564];
        i_10_470 <= in_reg[1076];
        i_10_471 <= in_reg[1588];
        i_10_472 <= in_reg[2100];
        i_10_473 <= in_reg[2612];
        i_10_474 <= in_reg[3124];
        i_10_475 <= in_reg[3636];
        i_10_476 <= in_reg[4148];
        i_10_477 <= in_reg[53];
        i_10_478 <= in_reg[565];
        i_10_479 <= in_reg[1077];
        i_10_480 <= in_reg[1589];
        i_10_481 <= in_reg[2101];
        i_10_482 <= in_reg[2613];
        i_10_483 <= in_reg[3125];
        i_10_484 <= in_reg[3637];
        i_10_485 <= in_reg[4149];
        i_10_486 <= in_reg[54];
        i_10_487 <= in_reg[566];
        i_10_488 <= in_reg[1078];
        i_10_489 <= in_reg[1590];
        i_10_490 <= in_reg[2102];
        i_10_491 <= in_reg[2614];
        i_10_492 <= in_reg[3126];
        i_10_493 <= in_reg[3638];
        i_10_494 <= in_reg[4150];
        i_10_495 <= in_reg[55];
        i_10_496 <= in_reg[567];
        i_10_497 <= in_reg[1079];
        i_10_498 <= in_reg[1591];
        i_10_499 <= in_reg[2103];
        i_10_500 <= in_reg[2615];
        i_10_501 <= in_reg[3127];
        i_10_502 <= in_reg[3639];
        i_10_503 <= in_reg[4151];
        i_10_504 <= in_reg[56];
        i_10_505 <= in_reg[568];
        i_10_506 <= in_reg[1080];
        i_10_507 <= in_reg[1592];
        i_10_508 <= in_reg[2104];
        i_10_509 <= in_reg[2616];
        i_10_510 <= in_reg[3128];
        i_10_511 <= in_reg[3640];
        i_10_512 <= in_reg[4152];
        i_10_513 <= in_reg[57];
        i_10_514 <= in_reg[569];
        i_10_515 <= in_reg[1081];
        i_10_516 <= in_reg[1593];
        i_10_517 <= in_reg[2105];
        i_10_518 <= in_reg[2617];
        i_10_519 <= in_reg[3129];
        i_10_520 <= in_reg[3641];
        i_10_521 <= in_reg[4153];
        i_10_522 <= in_reg[58];
        i_10_523 <= in_reg[570];
        i_10_524 <= in_reg[1082];
        i_10_525 <= in_reg[1594];
        i_10_526 <= in_reg[2106];
        i_10_527 <= in_reg[2618];
        i_10_528 <= in_reg[3130];
        i_10_529 <= in_reg[3642];
        i_10_530 <= in_reg[4154];
        i_10_531 <= in_reg[59];
        i_10_532 <= in_reg[571];
        i_10_533 <= in_reg[1083];
        i_10_534 <= in_reg[1595];
        i_10_535 <= in_reg[2107];
        i_10_536 <= in_reg[2619];
        i_10_537 <= in_reg[3131];
        i_10_538 <= in_reg[3643];
        i_10_539 <= in_reg[4155];
        i_10_540 <= in_reg[60];
        i_10_541 <= in_reg[572];
        i_10_542 <= in_reg[1084];
        i_10_543 <= in_reg[1596];
        i_10_544 <= in_reg[2108];
        i_10_545 <= in_reg[2620];
        i_10_546 <= in_reg[3132];
        i_10_547 <= in_reg[3644];
        i_10_548 <= in_reg[4156];
        i_10_549 <= in_reg[61];
        i_10_550 <= in_reg[573];
        i_10_551 <= in_reg[1085];
        i_10_552 <= in_reg[1597];
        i_10_553 <= in_reg[2109];
        i_10_554 <= in_reg[2621];
        i_10_555 <= in_reg[3133];
        i_10_556 <= in_reg[3645];
        i_10_557 <= in_reg[4157];
        i_10_558 <= in_reg[62];
        i_10_559 <= in_reg[574];
        i_10_560 <= in_reg[1086];
        i_10_561 <= in_reg[1598];
        i_10_562 <= in_reg[2110];
        i_10_563 <= in_reg[2622];
        i_10_564 <= in_reg[3134];
        i_10_565 <= in_reg[3646];
        i_10_566 <= in_reg[4158];
        i_10_567 <= in_reg[63];
        i_10_568 <= in_reg[575];
        i_10_569 <= in_reg[1087];
        i_10_570 <= in_reg[1599];
        i_10_571 <= in_reg[2111];
        i_10_572 <= in_reg[2623];
        i_10_573 <= in_reg[3135];
        i_10_574 <= in_reg[3647];
        i_10_575 <= in_reg[4159];
        i_10_576 <= in_reg[64];
        i_10_577 <= in_reg[576];
        i_10_578 <= in_reg[1088];
        i_10_579 <= in_reg[1600];
        i_10_580 <= in_reg[2112];
        i_10_581 <= in_reg[2624];
        i_10_582 <= in_reg[3136];
        i_10_583 <= in_reg[3648];
        i_10_584 <= in_reg[4160];
        i_10_585 <= in_reg[65];
        i_10_586 <= in_reg[577];
        i_10_587 <= in_reg[1089];
        i_10_588 <= in_reg[1601];
        i_10_589 <= in_reg[2113];
        i_10_590 <= in_reg[2625];
        i_10_591 <= in_reg[3137];
        i_10_592 <= in_reg[3649];
        i_10_593 <= in_reg[4161];
        i_10_594 <= in_reg[66];
        i_10_595 <= in_reg[578];
        i_10_596 <= in_reg[1090];
        i_10_597 <= in_reg[1602];
        i_10_598 <= in_reg[2114];
        i_10_599 <= in_reg[2626];
        i_10_600 <= in_reg[3138];
        i_10_601 <= in_reg[3650];
        i_10_602 <= in_reg[4162];
        i_10_603 <= in_reg[67];
        i_10_604 <= in_reg[579];
        i_10_605 <= in_reg[1091];
        i_10_606 <= in_reg[1603];
        i_10_607 <= in_reg[2115];
        i_10_608 <= in_reg[2627];
        i_10_609 <= in_reg[3139];
        i_10_610 <= in_reg[3651];
        i_10_611 <= in_reg[4163];
        i_10_612 <= in_reg[68];
        i_10_613 <= in_reg[580];
        i_10_614 <= in_reg[1092];
        i_10_615 <= in_reg[1604];
        i_10_616 <= in_reg[2116];
        i_10_617 <= in_reg[2628];
        i_10_618 <= in_reg[3140];
        i_10_619 <= in_reg[3652];
        i_10_620 <= in_reg[4164];
        i_10_621 <= in_reg[69];
        i_10_622 <= in_reg[581];
        i_10_623 <= in_reg[1093];
        i_10_624 <= in_reg[1605];
        i_10_625 <= in_reg[2117];
        i_10_626 <= in_reg[2629];
        i_10_627 <= in_reg[3141];
        i_10_628 <= in_reg[3653];
        i_10_629 <= in_reg[4165];
        i_10_630 <= in_reg[70];
        i_10_631 <= in_reg[582];
        i_10_632 <= in_reg[1094];
        i_10_633 <= in_reg[1606];
        i_10_634 <= in_reg[2118];
        i_10_635 <= in_reg[2630];
        i_10_636 <= in_reg[3142];
        i_10_637 <= in_reg[3654];
        i_10_638 <= in_reg[4166];
        i_10_639 <= in_reg[71];
        i_10_640 <= in_reg[583];
        i_10_641 <= in_reg[1095];
        i_10_642 <= in_reg[1607];
        i_10_643 <= in_reg[2119];
        i_10_644 <= in_reg[2631];
        i_10_645 <= in_reg[3143];
        i_10_646 <= in_reg[3655];
        i_10_647 <= in_reg[4167];
        i_10_648 <= in_reg[72];
        i_10_649 <= in_reg[584];
        i_10_650 <= in_reg[1096];
        i_10_651 <= in_reg[1608];
        i_10_652 <= in_reg[2120];
        i_10_653 <= in_reg[2632];
        i_10_654 <= in_reg[3144];
        i_10_655 <= in_reg[3656];
        i_10_656 <= in_reg[4168];
        i_10_657 <= in_reg[73];
        i_10_658 <= in_reg[585];
        i_10_659 <= in_reg[1097];
        i_10_660 <= in_reg[1609];
        i_10_661 <= in_reg[2121];
        i_10_662 <= in_reg[2633];
        i_10_663 <= in_reg[3145];
        i_10_664 <= in_reg[3657];
        i_10_665 <= in_reg[4169];
        i_10_666 <= in_reg[74];
        i_10_667 <= in_reg[586];
        i_10_668 <= in_reg[1098];
        i_10_669 <= in_reg[1610];
        i_10_670 <= in_reg[2122];
        i_10_671 <= in_reg[2634];
        i_10_672 <= in_reg[3146];
        i_10_673 <= in_reg[3658];
        i_10_674 <= in_reg[4170];
        i_10_675 <= in_reg[75];
        i_10_676 <= in_reg[587];
        i_10_677 <= in_reg[1099];
        i_10_678 <= in_reg[1611];
        i_10_679 <= in_reg[2123];
        i_10_680 <= in_reg[2635];
        i_10_681 <= in_reg[3147];
        i_10_682 <= in_reg[3659];
        i_10_683 <= in_reg[4171];
        i_10_684 <= in_reg[76];
        i_10_685 <= in_reg[588];
        i_10_686 <= in_reg[1100];
        i_10_687 <= in_reg[1612];
        i_10_688 <= in_reg[2124];
        i_10_689 <= in_reg[2636];
        i_10_690 <= in_reg[3148];
        i_10_691 <= in_reg[3660];
        i_10_692 <= in_reg[4172];
        i_10_693 <= in_reg[77];
        i_10_694 <= in_reg[589];
        i_10_695 <= in_reg[1101];
        i_10_696 <= in_reg[1613];
        i_10_697 <= in_reg[2125];
        i_10_698 <= in_reg[2637];
        i_10_699 <= in_reg[3149];
        i_10_700 <= in_reg[3661];
        i_10_701 <= in_reg[4173];
        i_10_702 <= in_reg[78];
        i_10_703 <= in_reg[590];
        i_10_704 <= in_reg[1102];
        i_10_705 <= in_reg[1614];
        i_10_706 <= in_reg[2126];
        i_10_707 <= in_reg[2638];
        i_10_708 <= in_reg[3150];
        i_10_709 <= in_reg[3662];
        i_10_710 <= in_reg[4174];
        i_10_711 <= in_reg[79];
        i_10_712 <= in_reg[591];
        i_10_713 <= in_reg[1103];
        i_10_714 <= in_reg[1615];
        i_10_715 <= in_reg[2127];
        i_10_716 <= in_reg[2639];
        i_10_717 <= in_reg[3151];
        i_10_718 <= in_reg[3663];
        i_10_719 <= in_reg[4175];
        i_10_720 <= in_reg[80];
        i_10_721 <= in_reg[592];
        i_10_722 <= in_reg[1104];
        i_10_723 <= in_reg[1616];
        i_10_724 <= in_reg[2128];
        i_10_725 <= in_reg[2640];
        i_10_726 <= in_reg[3152];
        i_10_727 <= in_reg[3664];
        i_10_728 <= in_reg[4176];
        i_10_729 <= in_reg[81];
        i_10_730 <= in_reg[593];
        i_10_731 <= in_reg[1105];
        i_10_732 <= in_reg[1617];
        i_10_733 <= in_reg[2129];
        i_10_734 <= in_reg[2641];
        i_10_735 <= in_reg[3153];
        i_10_736 <= in_reg[3665];
        i_10_737 <= in_reg[4177];
        i_10_738 <= in_reg[82];
        i_10_739 <= in_reg[594];
        i_10_740 <= in_reg[1106];
        i_10_741 <= in_reg[1618];
        i_10_742 <= in_reg[2130];
        i_10_743 <= in_reg[2642];
        i_10_744 <= in_reg[3154];
        i_10_745 <= in_reg[3666];
        i_10_746 <= in_reg[4178];
        i_10_747 <= in_reg[83];
        i_10_748 <= in_reg[595];
        i_10_749 <= in_reg[1107];
        i_10_750 <= in_reg[1619];
        i_10_751 <= in_reg[2131];
        i_10_752 <= in_reg[2643];
        i_10_753 <= in_reg[3155];
        i_10_754 <= in_reg[3667];
        i_10_755 <= in_reg[4179];
        i_10_756 <= in_reg[84];
        i_10_757 <= in_reg[596];
        i_10_758 <= in_reg[1108];
        i_10_759 <= in_reg[1620];
        i_10_760 <= in_reg[2132];
        i_10_761 <= in_reg[2644];
        i_10_762 <= in_reg[3156];
        i_10_763 <= in_reg[3668];
        i_10_764 <= in_reg[4180];
        i_10_765 <= in_reg[85];
        i_10_766 <= in_reg[597];
        i_10_767 <= in_reg[1109];
        i_10_768 <= in_reg[1621];
        i_10_769 <= in_reg[2133];
        i_10_770 <= in_reg[2645];
        i_10_771 <= in_reg[3157];
        i_10_772 <= in_reg[3669];
        i_10_773 <= in_reg[4181];
        i_10_774 <= in_reg[86];
        i_10_775 <= in_reg[598];
        i_10_776 <= in_reg[1110];
        i_10_777 <= in_reg[1622];
        i_10_778 <= in_reg[2134];
        i_10_779 <= in_reg[2646];
        i_10_780 <= in_reg[3158];
        i_10_781 <= in_reg[3670];
        i_10_782 <= in_reg[4182];
        i_10_783 <= in_reg[87];
        i_10_784 <= in_reg[599];
        i_10_785 <= in_reg[1111];
        i_10_786 <= in_reg[1623];
        i_10_787 <= in_reg[2135];
        i_10_788 <= in_reg[2647];
        i_10_789 <= in_reg[3159];
        i_10_790 <= in_reg[3671];
        i_10_791 <= in_reg[4183];
        i_10_792 <= in_reg[88];
        i_10_793 <= in_reg[600];
        i_10_794 <= in_reg[1112];
        i_10_795 <= in_reg[1624];
        i_10_796 <= in_reg[2136];
        i_10_797 <= in_reg[2648];
        i_10_798 <= in_reg[3160];
        i_10_799 <= in_reg[3672];
        i_10_800 <= in_reg[4184];
        i_10_801 <= in_reg[89];
        i_10_802 <= in_reg[601];
        i_10_803 <= in_reg[1113];
        i_10_804 <= in_reg[1625];
        i_10_805 <= in_reg[2137];
        i_10_806 <= in_reg[2649];
        i_10_807 <= in_reg[3161];
        i_10_808 <= in_reg[3673];
        i_10_809 <= in_reg[4185];
        i_10_810 <= in_reg[90];
        i_10_811 <= in_reg[602];
        i_10_812 <= in_reg[1114];
        i_10_813 <= in_reg[1626];
        i_10_814 <= in_reg[2138];
        i_10_815 <= in_reg[2650];
        i_10_816 <= in_reg[3162];
        i_10_817 <= in_reg[3674];
        i_10_818 <= in_reg[4186];
        i_10_819 <= in_reg[91];
        i_10_820 <= in_reg[603];
        i_10_821 <= in_reg[1115];
        i_10_822 <= in_reg[1627];
        i_10_823 <= in_reg[2139];
        i_10_824 <= in_reg[2651];
        i_10_825 <= in_reg[3163];
        i_10_826 <= in_reg[3675];
        i_10_827 <= in_reg[4187];
        i_10_828 <= in_reg[92];
        i_10_829 <= in_reg[604];
        i_10_830 <= in_reg[1116];
        i_10_831 <= in_reg[1628];
        i_10_832 <= in_reg[2140];
        i_10_833 <= in_reg[2652];
        i_10_834 <= in_reg[3164];
        i_10_835 <= in_reg[3676];
        i_10_836 <= in_reg[4188];
        i_10_837 <= in_reg[93];
        i_10_838 <= in_reg[605];
        i_10_839 <= in_reg[1117];
        i_10_840 <= in_reg[1629];
        i_10_841 <= in_reg[2141];
        i_10_842 <= in_reg[2653];
        i_10_843 <= in_reg[3165];
        i_10_844 <= in_reg[3677];
        i_10_845 <= in_reg[4189];
        i_10_846 <= in_reg[94];
        i_10_847 <= in_reg[606];
        i_10_848 <= in_reg[1118];
        i_10_849 <= in_reg[1630];
        i_10_850 <= in_reg[2142];
        i_10_851 <= in_reg[2654];
        i_10_852 <= in_reg[3166];
        i_10_853 <= in_reg[3678];
        i_10_854 <= in_reg[4190];
        i_10_855 <= in_reg[95];
        i_10_856 <= in_reg[607];
        i_10_857 <= in_reg[1119];
        i_10_858 <= in_reg[1631];
        i_10_859 <= in_reg[2143];
        i_10_860 <= in_reg[2655];
        i_10_861 <= in_reg[3167];
        i_10_862 <= in_reg[3679];
        i_10_863 <= in_reg[4191];
        i_10_864 <= in_reg[96];
        i_10_865 <= in_reg[608];
        i_10_866 <= in_reg[1120];
        i_10_867 <= in_reg[1632];
        i_10_868 <= in_reg[2144];
        i_10_869 <= in_reg[2656];
        i_10_870 <= in_reg[3168];
        i_10_871 <= in_reg[3680];
        i_10_872 <= in_reg[4192];
        i_10_873 <= in_reg[97];
        i_10_874 <= in_reg[609];
        i_10_875 <= in_reg[1121];
        i_10_876 <= in_reg[1633];
        i_10_877 <= in_reg[2145];
        i_10_878 <= in_reg[2657];
        i_10_879 <= in_reg[3169];
        i_10_880 <= in_reg[3681];
        i_10_881 <= in_reg[4193];
        i_10_882 <= in_reg[98];
        i_10_883 <= in_reg[610];
        i_10_884 <= in_reg[1122];
        i_10_885 <= in_reg[1634];
        i_10_886 <= in_reg[2146];
        i_10_887 <= in_reg[2658];
        i_10_888 <= in_reg[3170];
        i_10_889 <= in_reg[3682];
        i_10_890 <= in_reg[4194];
        i_10_891 <= in_reg[99];
        i_10_892 <= in_reg[611];
        i_10_893 <= in_reg[1123];
        i_10_894 <= in_reg[1635];
        i_10_895 <= in_reg[2147];
        i_10_896 <= in_reg[2659];
        i_10_897 <= in_reg[3171];
        i_10_898 <= in_reg[3683];
        i_10_899 <= in_reg[4195];
        i_10_900 <= in_reg[100];
        i_10_901 <= in_reg[612];
        i_10_902 <= in_reg[1124];
        i_10_903 <= in_reg[1636];
        i_10_904 <= in_reg[2148];
        i_10_905 <= in_reg[2660];
        i_10_906 <= in_reg[3172];
        i_10_907 <= in_reg[3684];
        i_10_908 <= in_reg[4196];
        i_10_909 <= in_reg[101];
        i_10_910 <= in_reg[613];
        i_10_911 <= in_reg[1125];
        i_10_912 <= in_reg[1637];
        i_10_913 <= in_reg[2149];
        i_10_914 <= in_reg[2661];
        i_10_915 <= in_reg[3173];
        i_10_916 <= in_reg[3685];
        i_10_917 <= in_reg[4197];
        i_10_918 <= in_reg[102];
        i_10_919 <= in_reg[614];
        i_10_920 <= in_reg[1126];
        i_10_921 <= in_reg[1638];
        i_10_922 <= in_reg[2150];
        i_10_923 <= in_reg[2662];
        i_10_924 <= in_reg[3174];
        i_10_925 <= in_reg[3686];
        i_10_926 <= in_reg[4198];
        i_10_927 <= in_reg[103];
        i_10_928 <= in_reg[615];
        i_10_929 <= in_reg[1127];
        i_10_930 <= in_reg[1639];
        i_10_931 <= in_reg[2151];
        i_10_932 <= in_reg[2663];
        i_10_933 <= in_reg[3175];
        i_10_934 <= in_reg[3687];
        i_10_935 <= in_reg[4199];
        i_10_936 <= in_reg[104];
        i_10_937 <= in_reg[616];
        i_10_938 <= in_reg[1128];
        i_10_939 <= in_reg[1640];
        i_10_940 <= in_reg[2152];
        i_10_941 <= in_reg[2664];
        i_10_942 <= in_reg[3176];
        i_10_943 <= in_reg[3688];
        i_10_944 <= in_reg[4200];
        i_10_945 <= in_reg[105];
        i_10_946 <= in_reg[617];
        i_10_947 <= in_reg[1129];
        i_10_948 <= in_reg[1641];
        i_10_949 <= in_reg[2153];
        i_10_950 <= in_reg[2665];
        i_10_951 <= in_reg[3177];
        i_10_952 <= in_reg[3689];
        i_10_953 <= in_reg[4201];
        i_10_954 <= in_reg[106];
        i_10_955 <= in_reg[618];
        i_10_956 <= in_reg[1130];
        i_10_957 <= in_reg[1642];
        i_10_958 <= in_reg[2154];
        i_10_959 <= in_reg[2666];
        i_10_960 <= in_reg[3178];
        i_10_961 <= in_reg[3690];
        i_10_962 <= in_reg[4202];
        i_10_963 <= in_reg[107];
        i_10_964 <= in_reg[619];
        i_10_965 <= in_reg[1131];
        i_10_966 <= in_reg[1643];
        i_10_967 <= in_reg[2155];
        i_10_968 <= in_reg[2667];
        i_10_969 <= in_reg[3179];
        i_10_970 <= in_reg[3691];
        i_10_971 <= in_reg[4203];
        i_10_972 <= in_reg[108];
        i_10_973 <= in_reg[620];
        i_10_974 <= in_reg[1132];
        i_10_975 <= in_reg[1644];
        i_10_976 <= in_reg[2156];
        i_10_977 <= in_reg[2668];
        i_10_978 <= in_reg[3180];
        i_10_979 <= in_reg[3692];
        i_10_980 <= in_reg[4204];
        i_10_981 <= in_reg[109];
        i_10_982 <= in_reg[621];
        i_10_983 <= in_reg[1133];
        i_10_984 <= in_reg[1645];
        i_10_985 <= in_reg[2157];
        i_10_986 <= in_reg[2669];
        i_10_987 <= in_reg[3181];
        i_10_988 <= in_reg[3693];
        i_10_989 <= in_reg[4205];
        i_10_990 <= in_reg[110];
        i_10_991 <= in_reg[622];
        i_10_992 <= in_reg[1134];
        i_10_993 <= in_reg[1646];
        i_10_994 <= in_reg[2158];
        i_10_995 <= in_reg[2670];
        i_10_996 <= in_reg[3182];
        i_10_997 <= in_reg[3694];
        i_10_998 <= in_reg[4206];
        i_10_999 <= in_reg[111];
        i_10_1000 <= in_reg[623];
        i_10_1001 <= in_reg[1135];
        i_10_1002 <= in_reg[1647];
        i_10_1003 <= in_reg[2159];
        i_10_1004 <= in_reg[2671];
        i_10_1005 <= in_reg[3183];
        i_10_1006 <= in_reg[3695];
        i_10_1007 <= in_reg[4207];
        i_10_1008 <= in_reg[112];
        i_10_1009 <= in_reg[624];
        i_10_1010 <= in_reg[1136];
        i_10_1011 <= in_reg[1648];
        i_10_1012 <= in_reg[2160];
        i_10_1013 <= in_reg[2672];
        i_10_1014 <= in_reg[3184];
        i_10_1015 <= in_reg[3696];
        i_10_1016 <= in_reg[4208];
        i_10_1017 <= in_reg[113];
        i_10_1018 <= in_reg[625];
        i_10_1019 <= in_reg[1137];
        i_10_1020 <= in_reg[1649];
        i_10_1021 <= in_reg[2161];
        i_10_1022 <= in_reg[2673];
        i_10_1023 <= in_reg[3185];
        i_10_1024 <= in_reg[3697];
        i_10_1025 <= in_reg[4209];
        i_10_1026 <= in_reg[114];
        i_10_1027 <= in_reg[626];
        i_10_1028 <= in_reg[1138];
        i_10_1029 <= in_reg[1650];
        i_10_1030 <= in_reg[2162];
        i_10_1031 <= in_reg[2674];
        i_10_1032 <= in_reg[3186];
        i_10_1033 <= in_reg[3698];
        i_10_1034 <= in_reg[4210];
        i_10_1035 <= in_reg[115];
        i_10_1036 <= in_reg[627];
        i_10_1037 <= in_reg[1139];
        i_10_1038 <= in_reg[1651];
        i_10_1039 <= in_reg[2163];
        i_10_1040 <= in_reg[2675];
        i_10_1041 <= in_reg[3187];
        i_10_1042 <= in_reg[3699];
        i_10_1043 <= in_reg[4211];
        i_10_1044 <= in_reg[116];
        i_10_1045 <= in_reg[628];
        i_10_1046 <= in_reg[1140];
        i_10_1047 <= in_reg[1652];
        i_10_1048 <= in_reg[2164];
        i_10_1049 <= in_reg[2676];
        i_10_1050 <= in_reg[3188];
        i_10_1051 <= in_reg[3700];
        i_10_1052 <= in_reg[4212];
        i_10_1053 <= in_reg[117];
        i_10_1054 <= in_reg[629];
        i_10_1055 <= in_reg[1141];
        i_10_1056 <= in_reg[1653];
        i_10_1057 <= in_reg[2165];
        i_10_1058 <= in_reg[2677];
        i_10_1059 <= in_reg[3189];
        i_10_1060 <= in_reg[3701];
        i_10_1061 <= in_reg[4213];
        i_10_1062 <= in_reg[118];
        i_10_1063 <= in_reg[630];
        i_10_1064 <= in_reg[1142];
        i_10_1065 <= in_reg[1654];
        i_10_1066 <= in_reg[2166];
        i_10_1067 <= in_reg[2678];
        i_10_1068 <= in_reg[3190];
        i_10_1069 <= in_reg[3702];
        i_10_1070 <= in_reg[4214];
        i_10_1071 <= in_reg[119];
        i_10_1072 <= in_reg[631];
        i_10_1073 <= in_reg[1143];
        i_10_1074 <= in_reg[1655];
        i_10_1075 <= in_reg[2167];
        i_10_1076 <= in_reg[2679];
        i_10_1077 <= in_reg[3191];
        i_10_1078 <= in_reg[3703];
        i_10_1079 <= in_reg[4215];
        i_10_1080 <= in_reg[120];
        i_10_1081 <= in_reg[632];
        i_10_1082 <= in_reg[1144];
        i_10_1083 <= in_reg[1656];
        i_10_1084 <= in_reg[2168];
        i_10_1085 <= in_reg[2680];
        i_10_1086 <= in_reg[3192];
        i_10_1087 <= in_reg[3704];
        i_10_1088 <= in_reg[4216];
        i_10_1089 <= in_reg[121];
        i_10_1090 <= in_reg[633];
        i_10_1091 <= in_reg[1145];
        i_10_1092 <= in_reg[1657];
        i_10_1093 <= in_reg[2169];
        i_10_1094 <= in_reg[2681];
        i_10_1095 <= in_reg[3193];
        i_10_1096 <= in_reg[3705];
        i_10_1097 <= in_reg[4217];
        i_10_1098 <= in_reg[122];
        i_10_1099 <= in_reg[634];
        i_10_1100 <= in_reg[1146];
        i_10_1101 <= in_reg[1658];
        i_10_1102 <= in_reg[2170];
        i_10_1103 <= in_reg[2682];
        i_10_1104 <= in_reg[3194];
        i_10_1105 <= in_reg[3706];
        i_10_1106 <= in_reg[4218];
        i_10_1107 <= in_reg[123];
        i_10_1108 <= in_reg[635];
        i_10_1109 <= in_reg[1147];
        i_10_1110 <= in_reg[1659];
        i_10_1111 <= in_reg[2171];
        i_10_1112 <= in_reg[2683];
        i_10_1113 <= in_reg[3195];
        i_10_1114 <= in_reg[3707];
        i_10_1115 <= in_reg[4219];
        i_10_1116 <= in_reg[124];
        i_10_1117 <= in_reg[636];
        i_10_1118 <= in_reg[1148];
        i_10_1119 <= in_reg[1660];
        i_10_1120 <= in_reg[2172];
        i_10_1121 <= in_reg[2684];
        i_10_1122 <= in_reg[3196];
        i_10_1123 <= in_reg[3708];
        i_10_1124 <= in_reg[4220];
        i_10_1125 <= in_reg[125];
        i_10_1126 <= in_reg[637];
        i_10_1127 <= in_reg[1149];
        i_10_1128 <= in_reg[1661];
        i_10_1129 <= in_reg[2173];
        i_10_1130 <= in_reg[2685];
        i_10_1131 <= in_reg[3197];
        i_10_1132 <= in_reg[3709];
        i_10_1133 <= in_reg[4221];
        i_10_1134 <= in_reg[126];
        i_10_1135 <= in_reg[638];
        i_10_1136 <= in_reg[1150];
        i_10_1137 <= in_reg[1662];
        i_10_1138 <= in_reg[2174];
        i_10_1139 <= in_reg[2686];
        i_10_1140 <= in_reg[3198];
        i_10_1141 <= in_reg[3710];
        i_10_1142 <= in_reg[4222];
        i_10_1143 <= in_reg[127];
        i_10_1144 <= in_reg[639];
        i_10_1145 <= in_reg[1151];
        i_10_1146 <= in_reg[1663];
        i_10_1147 <= in_reg[2175];
        i_10_1148 <= in_reg[2687];
        i_10_1149 <= in_reg[3199];
        i_10_1150 <= in_reg[3711];
        i_10_1151 <= in_reg[4223];
        i_10_1152 <= in_reg[128];
        i_10_1153 <= in_reg[640];
        i_10_1154 <= in_reg[1152];
        i_10_1155 <= in_reg[1664];
        i_10_1156 <= in_reg[2176];
        i_10_1157 <= in_reg[2688];
        i_10_1158 <= in_reg[3200];
        i_10_1159 <= in_reg[3712];
        i_10_1160 <= in_reg[4224];
        i_10_1161 <= in_reg[129];
        i_10_1162 <= in_reg[641];
        i_10_1163 <= in_reg[1153];
        i_10_1164 <= in_reg[1665];
        i_10_1165 <= in_reg[2177];
        i_10_1166 <= in_reg[2689];
        i_10_1167 <= in_reg[3201];
        i_10_1168 <= in_reg[3713];
        i_10_1169 <= in_reg[4225];
        i_10_1170 <= in_reg[130];
        i_10_1171 <= in_reg[642];
        i_10_1172 <= in_reg[1154];
        i_10_1173 <= in_reg[1666];
        i_10_1174 <= in_reg[2178];
        i_10_1175 <= in_reg[2690];
        i_10_1176 <= in_reg[3202];
        i_10_1177 <= in_reg[3714];
        i_10_1178 <= in_reg[4226];
        i_10_1179 <= in_reg[131];
        i_10_1180 <= in_reg[643];
        i_10_1181 <= in_reg[1155];
        i_10_1182 <= in_reg[1667];
        i_10_1183 <= in_reg[2179];
        i_10_1184 <= in_reg[2691];
        i_10_1185 <= in_reg[3203];
        i_10_1186 <= in_reg[3715];
        i_10_1187 <= in_reg[4227];
        i_10_1188 <= in_reg[132];
        i_10_1189 <= in_reg[644];
        i_10_1190 <= in_reg[1156];
        i_10_1191 <= in_reg[1668];
        i_10_1192 <= in_reg[2180];
        i_10_1193 <= in_reg[2692];
        i_10_1194 <= in_reg[3204];
        i_10_1195 <= in_reg[3716];
        i_10_1196 <= in_reg[4228];
        i_10_1197 <= in_reg[133];
        i_10_1198 <= in_reg[645];
        i_10_1199 <= in_reg[1157];
        i_10_1200 <= in_reg[1669];
        i_10_1201 <= in_reg[2181];
        i_10_1202 <= in_reg[2693];
        i_10_1203 <= in_reg[3205];
        i_10_1204 <= in_reg[3717];
        i_10_1205 <= in_reg[4229];
        i_10_1206 <= in_reg[134];
        i_10_1207 <= in_reg[646];
        i_10_1208 <= in_reg[1158];
        i_10_1209 <= in_reg[1670];
        i_10_1210 <= in_reg[2182];
        i_10_1211 <= in_reg[2694];
        i_10_1212 <= in_reg[3206];
        i_10_1213 <= in_reg[3718];
        i_10_1214 <= in_reg[4230];
        i_10_1215 <= in_reg[135];
        i_10_1216 <= in_reg[647];
        i_10_1217 <= in_reg[1159];
        i_10_1218 <= in_reg[1671];
        i_10_1219 <= in_reg[2183];
        i_10_1220 <= in_reg[2695];
        i_10_1221 <= in_reg[3207];
        i_10_1222 <= in_reg[3719];
        i_10_1223 <= in_reg[4231];
        i_10_1224 <= in_reg[136];
        i_10_1225 <= in_reg[648];
        i_10_1226 <= in_reg[1160];
        i_10_1227 <= in_reg[1672];
        i_10_1228 <= in_reg[2184];
        i_10_1229 <= in_reg[2696];
        i_10_1230 <= in_reg[3208];
        i_10_1231 <= in_reg[3720];
        i_10_1232 <= in_reg[4232];
        i_10_1233 <= in_reg[137];
        i_10_1234 <= in_reg[649];
        i_10_1235 <= in_reg[1161];
        i_10_1236 <= in_reg[1673];
        i_10_1237 <= in_reg[2185];
        i_10_1238 <= in_reg[2697];
        i_10_1239 <= in_reg[3209];
        i_10_1240 <= in_reg[3721];
        i_10_1241 <= in_reg[4233];
        i_10_1242 <= in_reg[138];
        i_10_1243 <= in_reg[650];
        i_10_1244 <= in_reg[1162];
        i_10_1245 <= in_reg[1674];
        i_10_1246 <= in_reg[2186];
        i_10_1247 <= in_reg[2698];
        i_10_1248 <= in_reg[3210];
        i_10_1249 <= in_reg[3722];
        i_10_1250 <= in_reg[4234];
        i_10_1251 <= in_reg[139];
        i_10_1252 <= in_reg[651];
        i_10_1253 <= in_reg[1163];
        i_10_1254 <= in_reg[1675];
        i_10_1255 <= in_reg[2187];
        i_10_1256 <= in_reg[2699];
        i_10_1257 <= in_reg[3211];
        i_10_1258 <= in_reg[3723];
        i_10_1259 <= in_reg[4235];
        i_10_1260 <= in_reg[140];
        i_10_1261 <= in_reg[652];
        i_10_1262 <= in_reg[1164];
        i_10_1263 <= in_reg[1676];
        i_10_1264 <= in_reg[2188];
        i_10_1265 <= in_reg[2700];
        i_10_1266 <= in_reg[3212];
        i_10_1267 <= in_reg[3724];
        i_10_1268 <= in_reg[4236];
        i_10_1269 <= in_reg[141];
        i_10_1270 <= in_reg[653];
        i_10_1271 <= in_reg[1165];
        i_10_1272 <= in_reg[1677];
        i_10_1273 <= in_reg[2189];
        i_10_1274 <= in_reg[2701];
        i_10_1275 <= in_reg[3213];
        i_10_1276 <= in_reg[3725];
        i_10_1277 <= in_reg[4237];
        i_10_1278 <= in_reg[142];
        i_10_1279 <= in_reg[654];
        i_10_1280 <= in_reg[1166];
        i_10_1281 <= in_reg[1678];
        i_10_1282 <= in_reg[2190];
        i_10_1283 <= in_reg[2702];
        i_10_1284 <= in_reg[3214];
        i_10_1285 <= in_reg[3726];
        i_10_1286 <= in_reg[4238];
        i_10_1287 <= in_reg[143];
        i_10_1288 <= in_reg[655];
        i_10_1289 <= in_reg[1167];
        i_10_1290 <= in_reg[1679];
        i_10_1291 <= in_reg[2191];
        i_10_1292 <= in_reg[2703];
        i_10_1293 <= in_reg[3215];
        i_10_1294 <= in_reg[3727];
        i_10_1295 <= in_reg[4239];
        i_10_1296 <= in_reg[144];
        i_10_1297 <= in_reg[656];
        i_10_1298 <= in_reg[1168];
        i_10_1299 <= in_reg[1680];
        i_10_1300 <= in_reg[2192];
        i_10_1301 <= in_reg[2704];
        i_10_1302 <= in_reg[3216];
        i_10_1303 <= in_reg[3728];
        i_10_1304 <= in_reg[4240];
        i_10_1305 <= in_reg[145];
        i_10_1306 <= in_reg[657];
        i_10_1307 <= in_reg[1169];
        i_10_1308 <= in_reg[1681];
        i_10_1309 <= in_reg[2193];
        i_10_1310 <= in_reg[2705];
        i_10_1311 <= in_reg[3217];
        i_10_1312 <= in_reg[3729];
        i_10_1313 <= in_reg[4241];
        i_10_1314 <= in_reg[146];
        i_10_1315 <= in_reg[658];
        i_10_1316 <= in_reg[1170];
        i_10_1317 <= in_reg[1682];
        i_10_1318 <= in_reg[2194];
        i_10_1319 <= in_reg[2706];
        i_10_1320 <= in_reg[3218];
        i_10_1321 <= in_reg[3730];
        i_10_1322 <= in_reg[4242];
        i_10_1323 <= in_reg[147];
        i_10_1324 <= in_reg[659];
        i_10_1325 <= in_reg[1171];
        i_10_1326 <= in_reg[1683];
        i_10_1327 <= in_reg[2195];
        i_10_1328 <= in_reg[2707];
        i_10_1329 <= in_reg[3219];
        i_10_1330 <= in_reg[3731];
        i_10_1331 <= in_reg[4243];
        i_10_1332 <= in_reg[148];
        i_10_1333 <= in_reg[660];
        i_10_1334 <= in_reg[1172];
        i_10_1335 <= in_reg[1684];
        i_10_1336 <= in_reg[2196];
        i_10_1337 <= in_reg[2708];
        i_10_1338 <= in_reg[3220];
        i_10_1339 <= in_reg[3732];
        i_10_1340 <= in_reg[4244];
        i_10_1341 <= in_reg[149];
        i_10_1342 <= in_reg[661];
        i_10_1343 <= in_reg[1173];
        i_10_1344 <= in_reg[1685];
        i_10_1345 <= in_reg[2197];
        i_10_1346 <= in_reg[2709];
        i_10_1347 <= in_reg[3221];
        i_10_1348 <= in_reg[3733];
        i_10_1349 <= in_reg[4245];
        i_10_1350 <= in_reg[150];
        i_10_1351 <= in_reg[662];
        i_10_1352 <= in_reg[1174];
        i_10_1353 <= in_reg[1686];
        i_10_1354 <= in_reg[2198];
        i_10_1355 <= in_reg[2710];
        i_10_1356 <= in_reg[3222];
        i_10_1357 <= in_reg[3734];
        i_10_1358 <= in_reg[4246];
        i_10_1359 <= in_reg[151];
        i_10_1360 <= in_reg[663];
        i_10_1361 <= in_reg[1175];
        i_10_1362 <= in_reg[1687];
        i_10_1363 <= in_reg[2199];
        i_10_1364 <= in_reg[2711];
        i_10_1365 <= in_reg[3223];
        i_10_1366 <= in_reg[3735];
        i_10_1367 <= in_reg[4247];
        i_10_1368 <= in_reg[152];
        i_10_1369 <= in_reg[664];
        i_10_1370 <= in_reg[1176];
        i_10_1371 <= in_reg[1688];
        i_10_1372 <= in_reg[2200];
        i_10_1373 <= in_reg[2712];
        i_10_1374 <= in_reg[3224];
        i_10_1375 <= in_reg[3736];
        i_10_1376 <= in_reg[4248];
        i_10_1377 <= in_reg[153];
        i_10_1378 <= in_reg[665];
        i_10_1379 <= in_reg[1177];
        i_10_1380 <= in_reg[1689];
        i_10_1381 <= in_reg[2201];
        i_10_1382 <= in_reg[2713];
        i_10_1383 <= in_reg[3225];
        i_10_1384 <= in_reg[3737];
        i_10_1385 <= in_reg[4249];
        i_10_1386 <= in_reg[154];
        i_10_1387 <= in_reg[666];
        i_10_1388 <= in_reg[1178];
        i_10_1389 <= in_reg[1690];
        i_10_1390 <= in_reg[2202];
        i_10_1391 <= in_reg[2714];
        i_10_1392 <= in_reg[3226];
        i_10_1393 <= in_reg[3738];
        i_10_1394 <= in_reg[4250];
        i_10_1395 <= in_reg[155];
        i_10_1396 <= in_reg[667];
        i_10_1397 <= in_reg[1179];
        i_10_1398 <= in_reg[1691];
        i_10_1399 <= in_reg[2203];
        i_10_1400 <= in_reg[2715];
        i_10_1401 <= in_reg[3227];
        i_10_1402 <= in_reg[3739];
        i_10_1403 <= in_reg[4251];
        i_10_1404 <= in_reg[156];
        i_10_1405 <= in_reg[668];
        i_10_1406 <= in_reg[1180];
        i_10_1407 <= in_reg[1692];
        i_10_1408 <= in_reg[2204];
        i_10_1409 <= in_reg[2716];
        i_10_1410 <= in_reg[3228];
        i_10_1411 <= in_reg[3740];
        i_10_1412 <= in_reg[4252];
        i_10_1413 <= in_reg[157];
        i_10_1414 <= in_reg[669];
        i_10_1415 <= in_reg[1181];
        i_10_1416 <= in_reg[1693];
        i_10_1417 <= in_reg[2205];
        i_10_1418 <= in_reg[2717];
        i_10_1419 <= in_reg[3229];
        i_10_1420 <= in_reg[3741];
        i_10_1421 <= in_reg[4253];
        i_10_1422 <= in_reg[158];
        i_10_1423 <= in_reg[670];
        i_10_1424 <= in_reg[1182];
        i_10_1425 <= in_reg[1694];
        i_10_1426 <= in_reg[2206];
        i_10_1427 <= in_reg[2718];
        i_10_1428 <= in_reg[3230];
        i_10_1429 <= in_reg[3742];
        i_10_1430 <= in_reg[4254];
        i_10_1431 <= in_reg[159];
        i_10_1432 <= in_reg[671];
        i_10_1433 <= in_reg[1183];
        i_10_1434 <= in_reg[1695];
        i_10_1435 <= in_reg[2207];
        i_10_1436 <= in_reg[2719];
        i_10_1437 <= in_reg[3231];
        i_10_1438 <= in_reg[3743];
        i_10_1439 <= in_reg[4255];
        i_10_1440 <= in_reg[160];
        i_10_1441 <= in_reg[672];
        i_10_1442 <= in_reg[1184];
        i_10_1443 <= in_reg[1696];
        i_10_1444 <= in_reg[2208];
        i_10_1445 <= in_reg[2720];
        i_10_1446 <= in_reg[3232];
        i_10_1447 <= in_reg[3744];
        i_10_1448 <= in_reg[4256];
        i_10_1449 <= in_reg[161];
        i_10_1450 <= in_reg[673];
        i_10_1451 <= in_reg[1185];
        i_10_1452 <= in_reg[1697];
        i_10_1453 <= in_reg[2209];
        i_10_1454 <= in_reg[2721];
        i_10_1455 <= in_reg[3233];
        i_10_1456 <= in_reg[3745];
        i_10_1457 <= in_reg[4257];
        i_10_1458 <= in_reg[162];
        i_10_1459 <= in_reg[674];
        i_10_1460 <= in_reg[1186];
        i_10_1461 <= in_reg[1698];
        i_10_1462 <= in_reg[2210];
        i_10_1463 <= in_reg[2722];
        i_10_1464 <= in_reg[3234];
        i_10_1465 <= in_reg[3746];
        i_10_1466 <= in_reg[4258];
        i_10_1467 <= in_reg[163];
        i_10_1468 <= in_reg[675];
        i_10_1469 <= in_reg[1187];
        i_10_1470 <= in_reg[1699];
        i_10_1471 <= in_reg[2211];
        i_10_1472 <= in_reg[2723];
        i_10_1473 <= in_reg[3235];
        i_10_1474 <= in_reg[3747];
        i_10_1475 <= in_reg[4259];
        i_10_1476 <= in_reg[164];
        i_10_1477 <= in_reg[676];
        i_10_1478 <= in_reg[1188];
        i_10_1479 <= in_reg[1700];
        i_10_1480 <= in_reg[2212];
        i_10_1481 <= in_reg[2724];
        i_10_1482 <= in_reg[3236];
        i_10_1483 <= in_reg[3748];
        i_10_1484 <= in_reg[4260];
        i_10_1485 <= in_reg[165];
        i_10_1486 <= in_reg[677];
        i_10_1487 <= in_reg[1189];
        i_10_1488 <= in_reg[1701];
        i_10_1489 <= in_reg[2213];
        i_10_1490 <= in_reg[2725];
        i_10_1491 <= in_reg[3237];
        i_10_1492 <= in_reg[3749];
        i_10_1493 <= in_reg[4261];
        i_10_1494 <= in_reg[166];
        i_10_1495 <= in_reg[678];
        i_10_1496 <= in_reg[1190];
        i_10_1497 <= in_reg[1702];
        i_10_1498 <= in_reg[2214];
        i_10_1499 <= in_reg[2726];
        i_10_1500 <= in_reg[3238];
        i_10_1501 <= in_reg[3750];
        i_10_1502 <= in_reg[4262];
        i_10_1503 <= in_reg[167];
        i_10_1504 <= in_reg[679];
        i_10_1505 <= in_reg[1191];
        i_10_1506 <= in_reg[1703];
        i_10_1507 <= in_reg[2215];
        i_10_1508 <= in_reg[2727];
        i_10_1509 <= in_reg[3239];
        i_10_1510 <= in_reg[3751];
        i_10_1511 <= in_reg[4263];
        i_10_1512 <= in_reg[168];
        i_10_1513 <= in_reg[680];
        i_10_1514 <= in_reg[1192];
        i_10_1515 <= in_reg[1704];
        i_10_1516 <= in_reg[2216];
        i_10_1517 <= in_reg[2728];
        i_10_1518 <= in_reg[3240];
        i_10_1519 <= in_reg[3752];
        i_10_1520 <= in_reg[4264];
        i_10_1521 <= in_reg[169];
        i_10_1522 <= in_reg[681];
        i_10_1523 <= in_reg[1193];
        i_10_1524 <= in_reg[1705];
        i_10_1525 <= in_reg[2217];
        i_10_1526 <= in_reg[2729];
        i_10_1527 <= in_reg[3241];
        i_10_1528 <= in_reg[3753];
        i_10_1529 <= in_reg[4265];
        i_10_1530 <= in_reg[170];
        i_10_1531 <= in_reg[682];
        i_10_1532 <= in_reg[1194];
        i_10_1533 <= in_reg[1706];
        i_10_1534 <= in_reg[2218];
        i_10_1535 <= in_reg[2730];
        i_10_1536 <= in_reg[3242];
        i_10_1537 <= in_reg[3754];
        i_10_1538 <= in_reg[4266];
        i_10_1539 <= in_reg[171];
        i_10_1540 <= in_reg[683];
        i_10_1541 <= in_reg[1195];
        i_10_1542 <= in_reg[1707];
        i_10_1543 <= in_reg[2219];
        i_10_1544 <= in_reg[2731];
        i_10_1545 <= in_reg[3243];
        i_10_1546 <= in_reg[3755];
        i_10_1547 <= in_reg[4267];
        i_10_1548 <= in_reg[172];
        i_10_1549 <= in_reg[684];
        i_10_1550 <= in_reg[1196];
        i_10_1551 <= in_reg[1708];
        i_10_1552 <= in_reg[2220];
        i_10_1553 <= in_reg[2732];
        i_10_1554 <= in_reg[3244];
        i_10_1555 <= in_reg[3756];
        i_10_1556 <= in_reg[4268];
        i_10_1557 <= in_reg[173];
        i_10_1558 <= in_reg[685];
        i_10_1559 <= in_reg[1197];
        i_10_1560 <= in_reg[1709];
        i_10_1561 <= in_reg[2221];
        i_10_1562 <= in_reg[2733];
        i_10_1563 <= in_reg[3245];
        i_10_1564 <= in_reg[3757];
        i_10_1565 <= in_reg[4269];
        i_10_1566 <= in_reg[174];
        i_10_1567 <= in_reg[686];
        i_10_1568 <= in_reg[1198];
        i_10_1569 <= in_reg[1710];
        i_10_1570 <= in_reg[2222];
        i_10_1571 <= in_reg[2734];
        i_10_1572 <= in_reg[3246];
        i_10_1573 <= in_reg[3758];
        i_10_1574 <= in_reg[4270];
        i_10_1575 <= in_reg[175];
        i_10_1576 <= in_reg[687];
        i_10_1577 <= in_reg[1199];
        i_10_1578 <= in_reg[1711];
        i_10_1579 <= in_reg[2223];
        i_10_1580 <= in_reg[2735];
        i_10_1581 <= in_reg[3247];
        i_10_1582 <= in_reg[3759];
        i_10_1583 <= in_reg[4271];
        i_10_1584 <= in_reg[176];
        i_10_1585 <= in_reg[688];
        i_10_1586 <= in_reg[1200];
        i_10_1587 <= in_reg[1712];
        i_10_1588 <= in_reg[2224];
        i_10_1589 <= in_reg[2736];
        i_10_1590 <= in_reg[3248];
        i_10_1591 <= in_reg[3760];
        i_10_1592 <= in_reg[4272];
        i_10_1593 <= in_reg[177];
        i_10_1594 <= in_reg[689];
        i_10_1595 <= in_reg[1201];
        i_10_1596 <= in_reg[1713];
        i_10_1597 <= in_reg[2225];
        i_10_1598 <= in_reg[2737];
        i_10_1599 <= in_reg[3249];
        i_10_1600 <= in_reg[3761];
        i_10_1601 <= in_reg[4273];
        i_10_1602 <= in_reg[178];
        i_10_1603 <= in_reg[690];
        i_10_1604 <= in_reg[1202];
        i_10_1605 <= in_reg[1714];
        i_10_1606 <= in_reg[2226];
        i_10_1607 <= in_reg[2738];
        i_10_1608 <= in_reg[3250];
        i_10_1609 <= in_reg[3762];
        i_10_1610 <= in_reg[4274];
        i_10_1611 <= in_reg[179];
        i_10_1612 <= in_reg[691];
        i_10_1613 <= in_reg[1203];
        i_10_1614 <= in_reg[1715];
        i_10_1615 <= in_reg[2227];
        i_10_1616 <= in_reg[2739];
        i_10_1617 <= in_reg[3251];
        i_10_1618 <= in_reg[3763];
        i_10_1619 <= in_reg[4275];
        i_10_1620 <= in_reg[180];
        i_10_1621 <= in_reg[692];
        i_10_1622 <= in_reg[1204];
        i_10_1623 <= in_reg[1716];
        i_10_1624 <= in_reg[2228];
        i_10_1625 <= in_reg[2740];
        i_10_1626 <= in_reg[3252];
        i_10_1627 <= in_reg[3764];
        i_10_1628 <= in_reg[4276];
        i_10_1629 <= in_reg[181];
        i_10_1630 <= in_reg[693];
        i_10_1631 <= in_reg[1205];
        i_10_1632 <= in_reg[1717];
        i_10_1633 <= in_reg[2229];
        i_10_1634 <= in_reg[2741];
        i_10_1635 <= in_reg[3253];
        i_10_1636 <= in_reg[3765];
        i_10_1637 <= in_reg[4277];
        i_10_1638 <= in_reg[182];
        i_10_1639 <= in_reg[694];
        i_10_1640 <= in_reg[1206];
        i_10_1641 <= in_reg[1718];
        i_10_1642 <= in_reg[2230];
        i_10_1643 <= in_reg[2742];
        i_10_1644 <= in_reg[3254];
        i_10_1645 <= in_reg[3766];
        i_10_1646 <= in_reg[4278];
        i_10_1647 <= in_reg[183];
        i_10_1648 <= in_reg[695];
        i_10_1649 <= in_reg[1207];
        i_10_1650 <= in_reg[1719];
        i_10_1651 <= in_reg[2231];
        i_10_1652 <= in_reg[2743];
        i_10_1653 <= in_reg[3255];
        i_10_1654 <= in_reg[3767];
        i_10_1655 <= in_reg[4279];
        i_10_1656 <= in_reg[184];
        i_10_1657 <= in_reg[696];
        i_10_1658 <= in_reg[1208];
        i_10_1659 <= in_reg[1720];
        i_10_1660 <= in_reg[2232];
        i_10_1661 <= in_reg[2744];
        i_10_1662 <= in_reg[3256];
        i_10_1663 <= in_reg[3768];
        i_10_1664 <= in_reg[4280];
        i_10_1665 <= in_reg[185];
        i_10_1666 <= in_reg[697];
        i_10_1667 <= in_reg[1209];
        i_10_1668 <= in_reg[1721];
        i_10_1669 <= in_reg[2233];
        i_10_1670 <= in_reg[2745];
        i_10_1671 <= in_reg[3257];
        i_10_1672 <= in_reg[3769];
        i_10_1673 <= in_reg[4281];
        i_10_1674 <= in_reg[186];
        i_10_1675 <= in_reg[698];
        i_10_1676 <= in_reg[1210];
        i_10_1677 <= in_reg[1722];
        i_10_1678 <= in_reg[2234];
        i_10_1679 <= in_reg[2746];
        i_10_1680 <= in_reg[3258];
        i_10_1681 <= in_reg[3770];
        i_10_1682 <= in_reg[4282];
        i_10_1683 <= in_reg[187];
        i_10_1684 <= in_reg[699];
        i_10_1685 <= in_reg[1211];
        i_10_1686 <= in_reg[1723];
        i_10_1687 <= in_reg[2235];
        i_10_1688 <= in_reg[2747];
        i_10_1689 <= in_reg[3259];
        i_10_1690 <= in_reg[3771];
        i_10_1691 <= in_reg[4283];
        i_10_1692 <= in_reg[188];
        i_10_1693 <= in_reg[700];
        i_10_1694 <= in_reg[1212];
        i_10_1695 <= in_reg[1724];
        i_10_1696 <= in_reg[2236];
        i_10_1697 <= in_reg[2748];
        i_10_1698 <= in_reg[3260];
        i_10_1699 <= in_reg[3772];
        i_10_1700 <= in_reg[4284];
        i_10_1701 <= in_reg[189];
        i_10_1702 <= in_reg[701];
        i_10_1703 <= in_reg[1213];
        i_10_1704 <= in_reg[1725];
        i_10_1705 <= in_reg[2237];
        i_10_1706 <= in_reg[2749];
        i_10_1707 <= in_reg[3261];
        i_10_1708 <= in_reg[3773];
        i_10_1709 <= in_reg[4285];
        i_10_1710 <= in_reg[190];
        i_10_1711 <= in_reg[702];
        i_10_1712 <= in_reg[1214];
        i_10_1713 <= in_reg[1726];
        i_10_1714 <= in_reg[2238];
        i_10_1715 <= in_reg[2750];
        i_10_1716 <= in_reg[3262];
        i_10_1717 <= in_reg[3774];
        i_10_1718 <= in_reg[4286];
        i_10_1719 <= in_reg[191];
        i_10_1720 <= in_reg[703];
        i_10_1721 <= in_reg[1215];
        i_10_1722 <= in_reg[1727];
        i_10_1723 <= in_reg[2239];
        i_10_1724 <= in_reg[2751];
        i_10_1725 <= in_reg[3263];
        i_10_1726 <= in_reg[3775];
        i_10_1727 <= in_reg[4287];
        i_10_1728 <= in_reg[192];
        i_10_1729 <= in_reg[704];
        i_10_1730 <= in_reg[1216];
        i_10_1731 <= in_reg[1728];
        i_10_1732 <= in_reg[2240];
        i_10_1733 <= in_reg[2752];
        i_10_1734 <= in_reg[3264];
        i_10_1735 <= in_reg[3776];
        i_10_1736 <= in_reg[4288];
        i_10_1737 <= in_reg[193];
        i_10_1738 <= in_reg[705];
        i_10_1739 <= in_reg[1217];
        i_10_1740 <= in_reg[1729];
        i_10_1741 <= in_reg[2241];
        i_10_1742 <= in_reg[2753];
        i_10_1743 <= in_reg[3265];
        i_10_1744 <= in_reg[3777];
        i_10_1745 <= in_reg[4289];
        i_10_1746 <= in_reg[194];
        i_10_1747 <= in_reg[706];
        i_10_1748 <= in_reg[1218];
        i_10_1749 <= in_reg[1730];
        i_10_1750 <= in_reg[2242];
        i_10_1751 <= in_reg[2754];
        i_10_1752 <= in_reg[3266];
        i_10_1753 <= in_reg[3778];
        i_10_1754 <= in_reg[4290];
        i_10_1755 <= in_reg[195];
        i_10_1756 <= in_reg[707];
        i_10_1757 <= in_reg[1219];
        i_10_1758 <= in_reg[1731];
        i_10_1759 <= in_reg[2243];
        i_10_1760 <= in_reg[2755];
        i_10_1761 <= in_reg[3267];
        i_10_1762 <= in_reg[3779];
        i_10_1763 <= in_reg[4291];
        i_10_1764 <= in_reg[196];
        i_10_1765 <= in_reg[708];
        i_10_1766 <= in_reg[1220];
        i_10_1767 <= in_reg[1732];
        i_10_1768 <= in_reg[2244];
        i_10_1769 <= in_reg[2756];
        i_10_1770 <= in_reg[3268];
        i_10_1771 <= in_reg[3780];
        i_10_1772 <= in_reg[4292];
        i_10_1773 <= in_reg[197];
        i_10_1774 <= in_reg[709];
        i_10_1775 <= in_reg[1221];
        i_10_1776 <= in_reg[1733];
        i_10_1777 <= in_reg[2245];
        i_10_1778 <= in_reg[2757];
        i_10_1779 <= in_reg[3269];
        i_10_1780 <= in_reg[3781];
        i_10_1781 <= in_reg[4293];
        i_10_1782 <= in_reg[198];
        i_10_1783 <= in_reg[710];
        i_10_1784 <= in_reg[1222];
        i_10_1785 <= in_reg[1734];
        i_10_1786 <= in_reg[2246];
        i_10_1787 <= in_reg[2758];
        i_10_1788 <= in_reg[3270];
        i_10_1789 <= in_reg[3782];
        i_10_1790 <= in_reg[4294];
        i_10_1791 <= in_reg[199];
        i_10_1792 <= in_reg[711];
        i_10_1793 <= in_reg[1223];
        i_10_1794 <= in_reg[1735];
        i_10_1795 <= in_reg[2247];
        i_10_1796 <= in_reg[2759];
        i_10_1797 <= in_reg[3271];
        i_10_1798 <= in_reg[3783];
        i_10_1799 <= in_reg[4295];
        i_10_1800 <= in_reg[200];
        i_10_1801 <= in_reg[712];
        i_10_1802 <= in_reg[1224];
        i_10_1803 <= in_reg[1736];
        i_10_1804 <= in_reg[2248];
        i_10_1805 <= in_reg[2760];
        i_10_1806 <= in_reg[3272];
        i_10_1807 <= in_reg[3784];
        i_10_1808 <= in_reg[4296];
        i_10_1809 <= in_reg[201];
        i_10_1810 <= in_reg[713];
        i_10_1811 <= in_reg[1225];
        i_10_1812 <= in_reg[1737];
        i_10_1813 <= in_reg[2249];
        i_10_1814 <= in_reg[2761];
        i_10_1815 <= in_reg[3273];
        i_10_1816 <= in_reg[3785];
        i_10_1817 <= in_reg[4297];
        i_10_1818 <= in_reg[202];
        i_10_1819 <= in_reg[714];
        i_10_1820 <= in_reg[1226];
        i_10_1821 <= in_reg[1738];
        i_10_1822 <= in_reg[2250];
        i_10_1823 <= in_reg[2762];
        i_10_1824 <= in_reg[3274];
        i_10_1825 <= in_reg[3786];
        i_10_1826 <= in_reg[4298];
        i_10_1827 <= in_reg[203];
        i_10_1828 <= in_reg[715];
        i_10_1829 <= in_reg[1227];
        i_10_1830 <= in_reg[1739];
        i_10_1831 <= in_reg[2251];
        i_10_1832 <= in_reg[2763];
        i_10_1833 <= in_reg[3275];
        i_10_1834 <= in_reg[3787];
        i_10_1835 <= in_reg[4299];
        i_10_1836 <= in_reg[204];
        i_10_1837 <= in_reg[716];
        i_10_1838 <= in_reg[1228];
        i_10_1839 <= in_reg[1740];
        i_10_1840 <= in_reg[2252];
        i_10_1841 <= in_reg[2764];
        i_10_1842 <= in_reg[3276];
        i_10_1843 <= in_reg[3788];
        i_10_1844 <= in_reg[4300];
        i_10_1845 <= in_reg[205];
        i_10_1846 <= in_reg[717];
        i_10_1847 <= in_reg[1229];
        i_10_1848 <= in_reg[1741];
        i_10_1849 <= in_reg[2253];
        i_10_1850 <= in_reg[2765];
        i_10_1851 <= in_reg[3277];
        i_10_1852 <= in_reg[3789];
        i_10_1853 <= in_reg[4301];
        i_10_1854 <= in_reg[206];
        i_10_1855 <= in_reg[718];
        i_10_1856 <= in_reg[1230];
        i_10_1857 <= in_reg[1742];
        i_10_1858 <= in_reg[2254];
        i_10_1859 <= in_reg[2766];
        i_10_1860 <= in_reg[3278];
        i_10_1861 <= in_reg[3790];
        i_10_1862 <= in_reg[4302];
        i_10_1863 <= in_reg[207];
        i_10_1864 <= in_reg[719];
        i_10_1865 <= in_reg[1231];
        i_10_1866 <= in_reg[1743];
        i_10_1867 <= in_reg[2255];
        i_10_1868 <= in_reg[2767];
        i_10_1869 <= in_reg[3279];
        i_10_1870 <= in_reg[3791];
        i_10_1871 <= in_reg[4303];
        i_10_1872 <= in_reg[208];
        i_10_1873 <= in_reg[720];
        i_10_1874 <= in_reg[1232];
        i_10_1875 <= in_reg[1744];
        i_10_1876 <= in_reg[2256];
        i_10_1877 <= in_reg[2768];
        i_10_1878 <= in_reg[3280];
        i_10_1879 <= in_reg[3792];
        i_10_1880 <= in_reg[4304];
        i_10_1881 <= in_reg[209];
        i_10_1882 <= in_reg[721];
        i_10_1883 <= in_reg[1233];
        i_10_1884 <= in_reg[1745];
        i_10_1885 <= in_reg[2257];
        i_10_1886 <= in_reg[2769];
        i_10_1887 <= in_reg[3281];
        i_10_1888 <= in_reg[3793];
        i_10_1889 <= in_reg[4305];
        i_10_1890 <= in_reg[210];
        i_10_1891 <= in_reg[722];
        i_10_1892 <= in_reg[1234];
        i_10_1893 <= in_reg[1746];
        i_10_1894 <= in_reg[2258];
        i_10_1895 <= in_reg[2770];
        i_10_1896 <= in_reg[3282];
        i_10_1897 <= in_reg[3794];
        i_10_1898 <= in_reg[4306];
        i_10_1899 <= in_reg[211];
        i_10_1900 <= in_reg[723];
        i_10_1901 <= in_reg[1235];
        i_10_1902 <= in_reg[1747];
        i_10_1903 <= in_reg[2259];
        i_10_1904 <= in_reg[2771];
        i_10_1905 <= in_reg[3283];
        i_10_1906 <= in_reg[3795];
        i_10_1907 <= in_reg[4307];
        i_10_1908 <= in_reg[212];
        i_10_1909 <= in_reg[724];
        i_10_1910 <= in_reg[1236];
        i_10_1911 <= in_reg[1748];
        i_10_1912 <= in_reg[2260];
        i_10_1913 <= in_reg[2772];
        i_10_1914 <= in_reg[3284];
        i_10_1915 <= in_reg[3796];
        i_10_1916 <= in_reg[4308];
        i_10_1917 <= in_reg[213];
        i_10_1918 <= in_reg[725];
        i_10_1919 <= in_reg[1237];
        i_10_1920 <= in_reg[1749];
        i_10_1921 <= in_reg[2261];
        i_10_1922 <= in_reg[2773];
        i_10_1923 <= in_reg[3285];
        i_10_1924 <= in_reg[3797];
        i_10_1925 <= in_reg[4309];
        i_10_1926 <= in_reg[214];
        i_10_1927 <= in_reg[726];
        i_10_1928 <= in_reg[1238];
        i_10_1929 <= in_reg[1750];
        i_10_1930 <= in_reg[2262];
        i_10_1931 <= in_reg[2774];
        i_10_1932 <= in_reg[3286];
        i_10_1933 <= in_reg[3798];
        i_10_1934 <= in_reg[4310];
        i_10_1935 <= in_reg[215];
        i_10_1936 <= in_reg[727];
        i_10_1937 <= in_reg[1239];
        i_10_1938 <= in_reg[1751];
        i_10_1939 <= in_reg[2263];
        i_10_1940 <= in_reg[2775];
        i_10_1941 <= in_reg[3287];
        i_10_1942 <= in_reg[3799];
        i_10_1943 <= in_reg[4311];
        i_10_1944 <= in_reg[216];
        i_10_1945 <= in_reg[728];
        i_10_1946 <= in_reg[1240];
        i_10_1947 <= in_reg[1752];
        i_10_1948 <= in_reg[2264];
        i_10_1949 <= in_reg[2776];
        i_10_1950 <= in_reg[3288];
        i_10_1951 <= in_reg[3800];
        i_10_1952 <= in_reg[4312];
        i_10_1953 <= in_reg[217];
        i_10_1954 <= in_reg[729];
        i_10_1955 <= in_reg[1241];
        i_10_1956 <= in_reg[1753];
        i_10_1957 <= in_reg[2265];
        i_10_1958 <= in_reg[2777];
        i_10_1959 <= in_reg[3289];
        i_10_1960 <= in_reg[3801];
        i_10_1961 <= in_reg[4313];
        i_10_1962 <= in_reg[218];
        i_10_1963 <= in_reg[730];
        i_10_1964 <= in_reg[1242];
        i_10_1965 <= in_reg[1754];
        i_10_1966 <= in_reg[2266];
        i_10_1967 <= in_reg[2778];
        i_10_1968 <= in_reg[3290];
        i_10_1969 <= in_reg[3802];
        i_10_1970 <= in_reg[4314];
        i_10_1971 <= in_reg[219];
        i_10_1972 <= in_reg[731];
        i_10_1973 <= in_reg[1243];
        i_10_1974 <= in_reg[1755];
        i_10_1975 <= in_reg[2267];
        i_10_1976 <= in_reg[2779];
        i_10_1977 <= in_reg[3291];
        i_10_1978 <= in_reg[3803];
        i_10_1979 <= in_reg[4315];
        i_10_1980 <= in_reg[220];
        i_10_1981 <= in_reg[732];
        i_10_1982 <= in_reg[1244];
        i_10_1983 <= in_reg[1756];
        i_10_1984 <= in_reg[2268];
        i_10_1985 <= in_reg[2780];
        i_10_1986 <= in_reg[3292];
        i_10_1987 <= in_reg[3804];
        i_10_1988 <= in_reg[4316];
        i_10_1989 <= in_reg[221];
        i_10_1990 <= in_reg[733];
        i_10_1991 <= in_reg[1245];
        i_10_1992 <= in_reg[1757];
        i_10_1993 <= in_reg[2269];
        i_10_1994 <= in_reg[2781];
        i_10_1995 <= in_reg[3293];
        i_10_1996 <= in_reg[3805];
        i_10_1997 <= in_reg[4317];
        i_10_1998 <= in_reg[222];
        i_10_1999 <= in_reg[734];
        i_10_2000 <= in_reg[1246];
        i_10_2001 <= in_reg[1758];
        i_10_2002 <= in_reg[2270];
        i_10_2003 <= in_reg[2782];
        i_10_2004 <= in_reg[3294];
        i_10_2005 <= in_reg[3806];
        i_10_2006 <= in_reg[4318];
        i_10_2007 <= in_reg[223];
        i_10_2008 <= in_reg[735];
        i_10_2009 <= in_reg[1247];
        i_10_2010 <= in_reg[1759];
        i_10_2011 <= in_reg[2271];
        i_10_2012 <= in_reg[2783];
        i_10_2013 <= in_reg[3295];
        i_10_2014 <= in_reg[3807];
        i_10_2015 <= in_reg[4319];
        i_10_2016 <= in_reg[224];
        i_10_2017 <= in_reg[736];
        i_10_2018 <= in_reg[1248];
        i_10_2019 <= in_reg[1760];
        i_10_2020 <= in_reg[2272];
        i_10_2021 <= in_reg[2784];
        i_10_2022 <= in_reg[3296];
        i_10_2023 <= in_reg[3808];
        i_10_2024 <= in_reg[4320];
        i_10_2025 <= in_reg[225];
        i_10_2026 <= in_reg[737];
        i_10_2027 <= in_reg[1249];
        i_10_2028 <= in_reg[1761];
        i_10_2029 <= in_reg[2273];
        i_10_2030 <= in_reg[2785];
        i_10_2031 <= in_reg[3297];
        i_10_2032 <= in_reg[3809];
        i_10_2033 <= in_reg[4321];
        i_10_2034 <= in_reg[226];
        i_10_2035 <= in_reg[738];
        i_10_2036 <= in_reg[1250];
        i_10_2037 <= in_reg[1762];
        i_10_2038 <= in_reg[2274];
        i_10_2039 <= in_reg[2786];
        i_10_2040 <= in_reg[3298];
        i_10_2041 <= in_reg[3810];
        i_10_2042 <= in_reg[4322];
        i_10_2043 <= in_reg[227];
        i_10_2044 <= in_reg[739];
        i_10_2045 <= in_reg[1251];
        i_10_2046 <= in_reg[1763];
        i_10_2047 <= in_reg[2275];
        i_10_2048 <= in_reg[2787];
        i_10_2049 <= in_reg[3299];
        i_10_2050 <= in_reg[3811];
        i_10_2051 <= in_reg[4323];
        i_10_2052 <= in_reg[228];
        i_10_2053 <= in_reg[740];
        i_10_2054 <= in_reg[1252];
        i_10_2055 <= in_reg[1764];
        i_10_2056 <= in_reg[2276];
        i_10_2057 <= in_reg[2788];
        i_10_2058 <= in_reg[3300];
        i_10_2059 <= in_reg[3812];
        i_10_2060 <= in_reg[4324];
        i_10_2061 <= in_reg[229];
        i_10_2062 <= in_reg[741];
        i_10_2063 <= in_reg[1253];
        i_10_2064 <= in_reg[1765];
        i_10_2065 <= in_reg[2277];
        i_10_2066 <= in_reg[2789];
        i_10_2067 <= in_reg[3301];
        i_10_2068 <= in_reg[3813];
        i_10_2069 <= in_reg[4325];
        i_10_2070 <= in_reg[230];
        i_10_2071 <= in_reg[742];
        i_10_2072 <= in_reg[1254];
        i_10_2073 <= in_reg[1766];
        i_10_2074 <= in_reg[2278];
        i_10_2075 <= in_reg[2790];
        i_10_2076 <= in_reg[3302];
        i_10_2077 <= in_reg[3814];
        i_10_2078 <= in_reg[4326];
        i_10_2079 <= in_reg[231];
        i_10_2080 <= in_reg[743];
        i_10_2081 <= in_reg[1255];
        i_10_2082 <= in_reg[1767];
        i_10_2083 <= in_reg[2279];
        i_10_2084 <= in_reg[2791];
        i_10_2085 <= in_reg[3303];
        i_10_2086 <= in_reg[3815];
        i_10_2087 <= in_reg[4327];
        i_10_2088 <= in_reg[232];
        i_10_2089 <= in_reg[744];
        i_10_2090 <= in_reg[1256];
        i_10_2091 <= in_reg[1768];
        i_10_2092 <= in_reg[2280];
        i_10_2093 <= in_reg[2792];
        i_10_2094 <= in_reg[3304];
        i_10_2095 <= in_reg[3816];
        i_10_2096 <= in_reg[4328];
        i_10_2097 <= in_reg[233];
        i_10_2098 <= in_reg[745];
        i_10_2099 <= in_reg[1257];
        i_10_2100 <= in_reg[1769];
        i_10_2101 <= in_reg[2281];
        i_10_2102 <= in_reg[2793];
        i_10_2103 <= in_reg[3305];
        i_10_2104 <= in_reg[3817];
        i_10_2105 <= in_reg[4329];
        i_10_2106 <= in_reg[234];
        i_10_2107 <= in_reg[746];
        i_10_2108 <= in_reg[1258];
        i_10_2109 <= in_reg[1770];
        i_10_2110 <= in_reg[2282];
        i_10_2111 <= in_reg[2794];
        i_10_2112 <= in_reg[3306];
        i_10_2113 <= in_reg[3818];
        i_10_2114 <= in_reg[4330];
        i_10_2115 <= in_reg[235];
        i_10_2116 <= in_reg[747];
        i_10_2117 <= in_reg[1259];
        i_10_2118 <= in_reg[1771];
        i_10_2119 <= in_reg[2283];
        i_10_2120 <= in_reg[2795];
        i_10_2121 <= in_reg[3307];
        i_10_2122 <= in_reg[3819];
        i_10_2123 <= in_reg[4331];
        i_10_2124 <= in_reg[236];
        i_10_2125 <= in_reg[748];
        i_10_2126 <= in_reg[1260];
        i_10_2127 <= in_reg[1772];
        i_10_2128 <= in_reg[2284];
        i_10_2129 <= in_reg[2796];
        i_10_2130 <= in_reg[3308];
        i_10_2131 <= in_reg[3820];
        i_10_2132 <= in_reg[4332];
        i_10_2133 <= in_reg[237];
        i_10_2134 <= in_reg[749];
        i_10_2135 <= in_reg[1261];
        i_10_2136 <= in_reg[1773];
        i_10_2137 <= in_reg[2285];
        i_10_2138 <= in_reg[2797];
        i_10_2139 <= in_reg[3309];
        i_10_2140 <= in_reg[3821];
        i_10_2141 <= in_reg[4333];
        i_10_2142 <= in_reg[238];
        i_10_2143 <= in_reg[750];
        i_10_2144 <= in_reg[1262];
        i_10_2145 <= in_reg[1774];
        i_10_2146 <= in_reg[2286];
        i_10_2147 <= in_reg[2798];
        i_10_2148 <= in_reg[3310];
        i_10_2149 <= in_reg[3822];
        i_10_2150 <= in_reg[4334];
        i_10_2151 <= in_reg[239];
        i_10_2152 <= in_reg[751];
        i_10_2153 <= in_reg[1263];
        i_10_2154 <= in_reg[1775];
        i_10_2155 <= in_reg[2287];
        i_10_2156 <= in_reg[2799];
        i_10_2157 <= in_reg[3311];
        i_10_2158 <= in_reg[3823];
        i_10_2159 <= in_reg[4335];
        i_10_2160 <= in_reg[240];
        i_10_2161 <= in_reg[752];
        i_10_2162 <= in_reg[1264];
        i_10_2163 <= in_reg[1776];
        i_10_2164 <= in_reg[2288];
        i_10_2165 <= in_reg[2800];
        i_10_2166 <= in_reg[3312];
        i_10_2167 <= in_reg[3824];
        i_10_2168 <= in_reg[4336];
        i_10_2169 <= in_reg[241];
        i_10_2170 <= in_reg[753];
        i_10_2171 <= in_reg[1265];
        i_10_2172 <= in_reg[1777];
        i_10_2173 <= in_reg[2289];
        i_10_2174 <= in_reg[2801];
        i_10_2175 <= in_reg[3313];
        i_10_2176 <= in_reg[3825];
        i_10_2177 <= in_reg[4337];
        i_10_2178 <= in_reg[242];
        i_10_2179 <= in_reg[754];
        i_10_2180 <= in_reg[1266];
        i_10_2181 <= in_reg[1778];
        i_10_2182 <= in_reg[2290];
        i_10_2183 <= in_reg[2802];
        i_10_2184 <= in_reg[3314];
        i_10_2185 <= in_reg[3826];
        i_10_2186 <= in_reg[4338];
        i_10_2187 <= in_reg[243];
        i_10_2188 <= in_reg[755];
        i_10_2189 <= in_reg[1267];
        i_10_2190 <= in_reg[1779];
        i_10_2191 <= in_reg[2291];
        i_10_2192 <= in_reg[2803];
        i_10_2193 <= in_reg[3315];
        i_10_2194 <= in_reg[3827];
        i_10_2195 <= in_reg[4339];
        i_10_2196 <= in_reg[244];
        i_10_2197 <= in_reg[756];
        i_10_2198 <= in_reg[1268];
        i_10_2199 <= in_reg[1780];
        i_10_2200 <= in_reg[2292];
        i_10_2201 <= in_reg[2804];
        i_10_2202 <= in_reg[3316];
        i_10_2203 <= in_reg[3828];
        i_10_2204 <= in_reg[4340];
        i_10_2205 <= in_reg[245];
        i_10_2206 <= in_reg[757];
        i_10_2207 <= in_reg[1269];
        i_10_2208 <= in_reg[1781];
        i_10_2209 <= in_reg[2293];
        i_10_2210 <= in_reg[2805];
        i_10_2211 <= in_reg[3317];
        i_10_2212 <= in_reg[3829];
        i_10_2213 <= in_reg[4341];
        i_10_2214 <= in_reg[246];
        i_10_2215 <= in_reg[758];
        i_10_2216 <= in_reg[1270];
        i_10_2217 <= in_reg[1782];
        i_10_2218 <= in_reg[2294];
        i_10_2219 <= in_reg[2806];
        i_10_2220 <= in_reg[3318];
        i_10_2221 <= in_reg[3830];
        i_10_2222 <= in_reg[4342];
        i_10_2223 <= in_reg[247];
        i_10_2224 <= in_reg[759];
        i_10_2225 <= in_reg[1271];
        i_10_2226 <= in_reg[1783];
        i_10_2227 <= in_reg[2295];
        i_10_2228 <= in_reg[2807];
        i_10_2229 <= in_reg[3319];
        i_10_2230 <= in_reg[3831];
        i_10_2231 <= in_reg[4343];
        i_10_2232 <= in_reg[248];
        i_10_2233 <= in_reg[760];
        i_10_2234 <= in_reg[1272];
        i_10_2235 <= in_reg[1784];
        i_10_2236 <= in_reg[2296];
        i_10_2237 <= in_reg[2808];
        i_10_2238 <= in_reg[3320];
        i_10_2239 <= in_reg[3832];
        i_10_2240 <= in_reg[4344];
        i_10_2241 <= in_reg[249];
        i_10_2242 <= in_reg[761];
        i_10_2243 <= in_reg[1273];
        i_10_2244 <= in_reg[1785];
        i_10_2245 <= in_reg[2297];
        i_10_2246 <= in_reg[2809];
        i_10_2247 <= in_reg[3321];
        i_10_2248 <= in_reg[3833];
        i_10_2249 <= in_reg[4345];
        i_10_2250 <= in_reg[250];
        i_10_2251 <= in_reg[762];
        i_10_2252 <= in_reg[1274];
        i_10_2253 <= in_reg[1786];
        i_10_2254 <= in_reg[2298];
        i_10_2255 <= in_reg[2810];
        i_10_2256 <= in_reg[3322];
        i_10_2257 <= in_reg[3834];
        i_10_2258 <= in_reg[4346];
        i_10_2259 <= in_reg[251];
        i_10_2260 <= in_reg[763];
        i_10_2261 <= in_reg[1275];
        i_10_2262 <= in_reg[1787];
        i_10_2263 <= in_reg[2299];
        i_10_2264 <= in_reg[2811];
        i_10_2265 <= in_reg[3323];
        i_10_2266 <= in_reg[3835];
        i_10_2267 <= in_reg[4347];
        i_10_2268 <= in_reg[252];
        i_10_2269 <= in_reg[764];
        i_10_2270 <= in_reg[1276];
        i_10_2271 <= in_reg[1788];
        i_10_2272 <= in_reg[2300];
        i_10_2273 <= in_reg[2812];
        i_10_2274 <= in_reg[3324];
        i_10_2275 <= in_reg[3836];
        i_10_2276 <= in_reg[4348];
        i_10_2277 <= in_reg[253];
        i_10_2278 <= in_reg[765];
        i_10_2279 <= in_reg[1277];
        i_10_2280 <= in_reg[1789];
        i_10_2281 <= in_reg[2301];
        i_10_2282 <= in_reg[2813];
        i_10_2283 <= in_reg[3325];
        i_10_2284 <= in_reg[3837];
        i_10_2285 <= in_reg[4349];
        i_10_2286 <= in_reg[254];
        i_10_2287 <= in_reg[766];
        i_10_2288 <= in_reg[1278];
        i_10_2289 <= in_reg[1790];
        i_10_2290 <= in_reg[2302];
        i_10_2291 <= in_reg[2814];
        i_10_2292 <= in_reg[3326];
        i_10_2293 <= in_reg[3838];
        i_10_2294 <= in_reg[4350];
        i_10_2295 <= in_reg[255];
        i_10_2296 <= in_reg[767];
        i_10_2297 <= in_reg[1279];
        i_10_2298 <= in_reg[1791];
        i_10_2299 <= in_reg[2303];
        i_10_2300 <= in_reg[2815];
        i_10_2301 <= in_reg[3327];
        i_10_2302 <= in_reg[3839];
        i_10_2303 <= in_reg[4351];
        i_10_2304 <= in_reg[256];
        i_10_2305 <= in_reg[768];
        i_10_2306 <= in_reg[1280];
        i_10_2307 <= in_reg[1792];
        i_10_2308 <= in_reg[2304];
        i_10_2309 <= in_reg[2816];
        i_10_2310 <= in_reg[3328];
        i_10_2311 <= in_reg[3840];
        i_10_2312 <= in_reg[4352];
        i_10_2313 <= in_reg[257];
        i_10_2314 <= in_reg[769];
        i_10_2315 <= in_reg[1281];
        i_10_2316 <= in_reg[1793];
        i_10_2317 <= in_reg[2305];
        i_10_2318 <= in_reg[2817];
        i_10_2319 <= in_reg[3329];
        i_10_2320 <= in_reg[3841];
        i_10_2321 <= in_reg[4353];
        i_10_2322 <= in_reg[258];
        i_10_2323 <= in_reg[770];
        i_10_2324 <= in_reg[1282];
        i_10_2325 <= in_reg[1794];
        i_10_2326 <= in_reg[2306];
        i_10_2327 <= in_reg[2818];
        i_10_2328 <= in_reg[3330];
        i_10_2329 <= in_reg[3842];
        i_10_2330 <= in_reg[4354];
        i_10_2331 <= in_reg[259];
        i_10_2332 <= in_reg[771];
        i_10_2333 <= in_reg[1283];
        i_10_2334 <= in_reg[1795];
        i_10_2335 <= in_reg[2307];
        i_10_2336 <= in_reg[2819];
        i_10_2337 <= in_reg[3331];
        i_10_2338 <= in_reg[3843];
        i_10_2339 <= in_reg[4355];
        i_10_2340 <= in_reg[260];
        i_10_2341 <= in_reg[772];
        i_10_2342 <= in_reg[1284];
        i_10_2343 <= in_reg[1796];
        i_10_2344 <= in_reg[2308];
        i_10_2345 <= in_reg[2820];
        i_10_2346 <= in_reg[3332];
        i_10_2347 <= in_reg[3844];
        i_10_2348 <= in_reg[4356];
        i_10_2349 <= in_reg[261];
        i_10_2350 <= in_reg[773];
        i_10_2351 <= in_reg[1285];
        i_10_2352 <= in_reg[1797];
        i_10_2353 <= in_reg[2309];
        i_10_2354 <= in_reg[2821];
        i_10_2355 <= in_reg[3333];
        i_10_2356 <= in_reg[3845];
        i_10_2357 <= in_reg[4357];
        i_10_2358 <= in_reg[262];
        i_10_2359 <= in_reg[774];
        i_10_2360 <= in_reg[1286];
        i_10_2361 <= in_reg[1798];
        i_10_2362 <= in_reg[2310];
        i_10_2363 <= in_reg[2822];
        i_10_2364 <= in_reg[3334];
        i_10_2365 <= in_reg[3846];
        i_10_2366 <= in_reg[4358];
        i_10_2367 <= in_reg[263];
        i_10_2368 <= in_reg[775];
        i_10_2369 <= in_reg[1287];
        i_10_2370 <= in_reg[1799];
        i_10_2371 <= in_reg[2311];
        i_10_2372 <= in_reg[2823];
        i_10_2373 <= in_reg[3335];
        i_10_2374 <= in_reg[3847];
        i_10_2375 <= in_reg[4359];
        i_10_2376 <= in_reg[264];
        i_10_2377 <= in_reg[776];
        i_10_2378 <= in_reg[1288];
        i_10_2379 <= in_reg[1800];
        i_10_2380 <= in_reg[2312];
        i_10_2381 <= in_reg[2824];
        i_10_2382 <= in_reg[3336];
        i_10_2383 <= in_reg[3848];
        i_10_2384 <= in_reg[4360];
        i_10_2385 <= in_reg[265];
        i_10_2386 <= in_reg[777];
        i_10_2387 <= in_reg[1289];
        i_10_2388 <= in_reg[1801];
        i_10_2389 <= in_reg[2313];
        i_10_2390 <= in_reg[2825];
        i_10_2391 <= in_reg[3337];
        i_10_2392 <= in_reg[3849];
        i_10_2393 <= in_reg[4361];
        i_10_2394 <= in_reg[266];
        i_10_2395 <= in_reg[778];
        i_10_2396 <= in_reg[1290];
        i_10_2397 <= in_reg[1802];
        i_10_2398 <= in_reg[2314];
        i_10_2399 <= in_reg[2826];
        i_10_2400 <= in_reg[3338];
        i_10_2401 <= in_reg[3850];
        i_10_2402 <= in_reg[4362];
        i_10_2403 <= in_reg[267];
        i_10_2404 <= in_reg[779];
        i_10_2405 <= in_reg[1291];
        i_10_2406 <= in_reg[1803];
        i_10_2407 <= in_reg[2315];
        i_10_2408 <= in_reg[2827];
        i_10_2409 <= in_reg[3339];
        i_10_2410 <= in_reg[3851];
        i_10_2411 <= in_reg[4363];
        i_10_2412 <= in_reg[268];
        i_10_2413 <= in_reg[780];
        i_10_2414 <= in_reg[1292];
        i_10_2415 <= in_reg[1804];
        i_10_2416 <= in_reg[2316];
        i_10_2417 <= in_reg[2828];
        i_10_2418 <= in_reg[3340];
        i_10_2419 <= in_reg[3852];
        i_10_2420 <= in_reg[4364];
        i_10_2421 <= in_reg[269];
        i_10_2422 <= in_reg[781];
        i_10_2423 <= in_reg[1293];
        i_10_2424 <= in_reg[1805];
        i_10_2425 <= in_reg[2317];
        i_10_2426 <= in_reg[2829];
        i_10_2427 <= in_reg[3341];
        i_10_2428 <= in_reg[3853];
        i_10_2429 <= in_reg[4365];
        i_10_2430 <= in_reg[270];
        i_10_2431 <= in_reg[782];
        i_10_2432 <= in_reg[1294];
        i_10_2433 <= in_reg[1806];
        i_10_2434 <= in_reg[2318];
        i_10_2435 <= in_reg[2830];
        i_10_2436 <= in_reg[3342];
        i_10_2437 <= in_reg[3854];
        i_10_2438 <= in_reg[4366];
        i_10_2439 <= in_reg[271];
        i_10_2440 <= in_reg[783];
        i_10_2441 <= in_reg[1295];
        i_10_2442 <= in_reg[1807];
        i_10_2443 <= in_reg[2319];
        i_10_2444 <= in_reg[2831];
        i_10_2445 <= in_reg[3343];
        i_10_2446 <= in_reg[3855];
        i_10_2447 <= in_reg[4367];
        i_10_2448 <= in_reg[272];
        i_10_2449 <= in_reg[784];
        i_10_2450 <= in_reg[1296];
        i_10_2451 <= in_reg[1808];
        i_10_2452 <= in_reg[2320];
        i_10_2453 <= in_reg[2832];
        i_10_2454 <= in_reg[3344];
        i_10_2455 <= in_reg[3856];
        i_10_2456 <= in_reg[4368];
        i_10_2457 <= in_reg[273];
        i_10_2458 <= in_reg[785];
        i_10_2459 <= in_reg[1297];
        i_10_2460 <= in_reg[1809];
        i_10_2461 <= in_reg[2321];
        i_10_2462 <= in_reg[2833];
        i_10_2463 <= in_reg[3345];
        i_10_2464 <= in_reg[3857];
        i_10_2465 <= in_reg[4369];
        i_10_2466 <= in_reg[274];
        i_10_2467 <= in_reg[786];
        i_10_2468 <= in_reg[1298];
        i_10_2469 <= in_reg[1810];
        i_10_2470 <= in_reg[2322];
        i_10_2471 <= in_reg[2834];
        i_10_2472 <= in_reg[3346];
        i_10_2473 <= in_reg[3858];
        i_10_2474 <= in_reg[4370];
        i_10_2475 <= in_reg[275];
        i_10_2476 <= in_reg[787];
        i_10_2477 <= in_reg[1299];
        i_10_2478 <= in_reg[1811];
        i_10_2479 <= in_reg[2323];
        i_10_2480 <= in_reg[2835];
        i_10_2481 <= in_reg[3347];
        i_10_2482 <= in_reg[3859];
        i_10_2483 <= in_reg[4371];
        i_10_2484 <= in_reg[276];
        i_10_2485 <= in_reg[788];
        i_10_2486 <= in_reg[1300];
        i_10_2487 <= in_reg[1812];
        i_10_2488 <= in_reg[2324];
        i_10_2489 <= in_reg[2836];
        i_10_2490 <= in_reg[3348];
        i_10_2491 <= in_reg[3860];
        i_10_2492 <= in_reg[4372];
        i_10_2493 <= in_reg[277];
        i_10_2494 <= in_reg[789];
        i_10_2495 <= in_reg[1301];
        i_10_2496 <= in_reg[1813];
        i_10_2497 <= in_reg[2325];
        i_10_2498 <= in_reg[2837];
        i_10_2499 <= in_reg[3349];
        i_10_2500 <= in_reg[3861];
        i_10_2501 <= in_reg[4373];
        i_10_2502 <= in_reg[278];
        i_10_2503 <= in_reg[790];
        i_10_2504 <= in_reg[1302];
        i_10_2505 <= in_reg[1814];
        i_10_2506 <= in_reg[2326];
        i_10_2507 <= in_reg[2838];
        i_10_2508 <= in_reg[3350];
        i_10_2509 <= in_reg[3862];
        i_10_2510 <= in_reg[4374];
        i_10_2511 <= in_reg[279];
        i_10_2512 <= in_reg[791];
        i_10_2513 <= in_reg[1303];
        i_10_2514 <= in_reg[1815];
        i_10_2515 <= in_reg[2327];
        i_10_2516 <= in_reg[2839];
        i_10_2517 <= in_reg[3351];
        i_10_2518 <= in_reg[3863];
        i_10_2519 <= in_reg[4375];
        i_10_2520 <= in_reg[280];
        i_10_2521 <= in_reg[792];
        i_10_2522 <= in_reg[1304];
        i_10_2523 <= in_reg[1816];
        i_10_2524 <= in_reg[2328];
        i_10_2525 <= in_reg[2840];
        i_10_2526 <= in_reg[3352];
        i_10_2527 <= in_reg[3864];
        i_10_2528 <= in_reg[4376];
        i_10_2529 <= in_reg[281];
        i_10_2530 <= in_reg[793];
        i_10_2531 <= in_reg[1305];
        i_10_2532 <= in_reg[1817];
        i_10_2533 <= in_reg[2329];
        i_10_2534 <= in_reg[2841];
        i_10_2535 <= in_reg[3353];
        i_10_2536 <= in_reg[3865];
        i_10_2537 <= in_reg[4377];
        i_10_2538 <= in_reg[282];
        i_10_2539 <= in_reg[794];
        i_10_2540 <= in_reg[1306];
        i_10_2541 <= in_reg[1818];
        i_10_2542 <= in_reg[2330];
        i_10_2543 <= in_reg[2842];
        i_10_2544 <= in_reg[3354];
        i_10_2545 <= in_reg[3866];
        i_10_2546 <= in_reg[4378];
        i_10_2547 <= in_reg[283];
        i_10_2548 <= in_reg[795];
        i_10_2549 <= in_reg[1307];
        i_10_2550 <= in_reg[1819];
        i_10_2551 <= in_reg[2331];
        i_10_2552 <= in_reg[2843];
        i_10_2553 <= in_reg[3355];
        i_10_2554 <= in_reg[3867];
        i_10_2555 <= in_reg[4379];
        i_10_2556 <= in_reg[284];
        i_10_2557 <= in_reg[796];
        i_10_2558 <= in_reg[1308];
        i_10_2559 <= in_reg[1820];
        i_10_2560 <= in_reg[2332];
        i_10_2561 <= in_reg[2844];
        i_10_2562 <= in_reg[3356];
        i_10_2563 <= in_reg[3868];
        i_10_2564 <= in_reg[4380];
        i_10_2565 <= in_reg[285];
        i_10_2566 <= in_reg[797];
        i_10_2567 <= in_reg[1309];
        i_10_2568 <= in_reg[1821];
        i_10_2569 <= in_reg[2333];
        i_10_2570 <= in_reg[2845];
        i_10_2571 <= in_reg[3357];
        i_10_2572 <= in_reg[3869];
        i_10_2573 <= in_reg[4381];
        i_10_2574 <= in_reg[286];
        i_10_2575 <= in_reg[798];
        i_10_2576 <= in_reg[1310];
        i_10_2577 <= in_reg[1822];
        i_10_2578 <= in_reg[2334];
        i_10_2579 <= in_reg[2846];
        i_10_2580 <= in_reg[3358];
        i_10_2581 <= in_reg[3870];
        i_10_2582 <= in_reg[4382];
        i_10_2583 <= in_reg[287];
        i_10_2584 <= in_reg[799];
        i_10_2585 <= in_reg[1311];
        i_10_2586 <= in_reg[1823];
        i_10_2587 <= in_reg[2335];
        i_10_2588 <= in_reg[2847];
        i_10_2589 <= in_reg[3359];
        i_10_2590 <= in_reg[3871];
        i_10_2591 <= in_reg[4383];
        i_10_2592 <= in_reg[288];
        i_10_2593 <= in_reg[800];
        i_10_2594 <= in_reg[1312];
        i_10_2595 <= in_reg[1824];
        i_10_2596 <= in_reg[2336];
        i_10_2597 <= in_reg[2848];
        i_10_2598 <= in_reg[3360];
        i_10_2599 <= in_reg[3872];
        i_10_2600 <= in_reg[4384];
        i_10_2601 <= in_reg[289];
        i_10_2602 <= in_reg[801];
        i_10_2603 <= in_reg[1313];
        i_10_2604 <= in_reg[1825];
        i_10_2605 <= in_reg[2337];
        i_10_2606 <= in_reg[2849];
        i_10_2607 <= in_reg[3361];
        i_10_2608 <= in_reg[3873];
        i_10_2609 <= in_reg[4385];
        i_10_2610 <= in_reg[290];
        i_10_2611 <= in_reg[802];
        i_10_2612 <= in_reg[1314];
        i_10_2613 <= in_reg[1826];
        i_10_2614 <= in_reg[2338];
        i_10_2615 <= in_reg[2850];
        i_10_2616 <= in_reg[3362];
        i_10_2617 <= in_reg[3874];
        i_10_2618 <= in_reg[4386];
        i_10_2619 <= in_reg[291];
        i_10_2620 <= in_reg[803];
        i_10_2621 <= in_reg[1315];
        i_10_2622 <= in_reg[1827];
        i_10_2623 <= in_reg[2339];
        i_10_2624 <= in_reg[2851];
        i_10_2625 <= in_reg[3363];
        i_10_2626 <= in_reg[3875];
        i_10_2627 <= in_reg[4387];
        i_10_2628 <= in_reg[292];
        i_10_2629 <= in_reg[804];
        i_10_2630 <= in_reg[1316];
        i_10_2631 <= in_reg[1828];
        i_10_2632 <= in_reg[2340];
        i_10_2633 <= in_reg[2852];
        i_10_2634 <= in_reg[3364];
        i_10_2635 <= in_reg[3876];
        i_10_2636 <= in_reg[4388];
        i_10_2637 <= in_reg[293];
        i_10_2638 <= in_reg[805];
        i_10_2639 <= in_reg[1317];
        i_10_2640 <= in_reg[1829];
        i_10_2641 <= in_reg[2341];
        i_10_2642 <= in_reg[2853];
        i_10_2643 <= in_reg[3365];
        i_10_2644 <= in_reg[3877];
        i_10_2645 <= in_reg[4389];
        i_10_2646 <= in_reg[294];
        i_10_2647 <= in_reg[806];
        i_10_2648 <= in_reg[1318];
        i_10_2649 <= in_reg[1830];
        i_10_2650 <= in_reg[2342];
        i_10_2651 <= in_reg[2854];
        i_10_2652 <= in_reg[3366];
        i_10_2653 <= in_reg[3878];
        i_10_2654 <= in_reg[4390];
        i_10_2655 <= in_reg[295];
        i_10_2656 <= in_reg[807];
        i_10_2657 <= in_reg[1319];
        i_10_2658 <= in_reg[1831];
        i_10_2659 <= in_reg[2343];
        i_10_2660 <= in_reg[2855];
        i_10_2661 <= in_reg[3367];
        i_10_2662 <= in_reg[3879];
        i_10_2663 <= in_reg[4391];
        i_10_2664 <= in_reg[296];
        i_10_2665 <= in_reg[808];
        i_10_2666 <= in_reg[1320];
        i_10_2667 <= in_reg[1832];
        i_10_2668 <= in_reg[2344];
        i_10_2669 <= in_reg[2856];
        i_10_2670 <= in_reg[3368];
        i_10_2671 <= in_reg[3880];
        i_10_2672 <= in_reg[4392];
        i_10_2673 <= in_reg[297];
        i_10_2674 <= in_reg[809];
        i_10_2675 <= in_reg[1321];
        i_10_2676 <= in_reg[1833];
        i_10_2677 <= in_reg[2345];
        i_10_2678 <= in_reg[2857];
        i_10_2679 <= in_reg[3369];
        i_10_2680 <= in_reg[3881];
        i_10_2681 <= in_reg[4393];
        i_10_2682 <= in_reg[298];
        i_10_2683 <= in_reg[810];
        i_10_2684 <= in_reg[1322];
        i_10_2685 <= in_reg[1834];
        i_10_2686 <= in_reg[2346];
        i_10_2687 <= in_reg[2858];
        i_10_2688 <= in_reg[3370];
        i_10_2689 <= in_reg[3882];
        i_10_2690 <= in_reg[4394];
        i_10_2691 <= in_reg[299];
        i_10_2692 <= in_reg[811];
        i_10_2693 <= in_reg[1323];
        i_10_2694 <= in_reg[1835];
        i_10_2695 <= in_reg[2347];
        i_10_2696 <= in_reg[2859];
        i_10_2697 <= in_reg[3371];
        i_10_2698 <= in_reg[3883];
        i_10_2699 <= in_reg[4395];
        i_10_2700 <= in_reg[300];
        i_10_2701 <= in_reg[812];
        i_10_2702 <= in_reg[1324];
        i_10_2703 <= in_reg[1836];
        i_10_2704 <= in_reg[2348];
        i_10_2705 <= in_reg[2860];
        i_10_2706 <= in_reg[3372];
        i_10_2707 <= in_reg[3884];
        i_10_2708 <= in_reg[4396];
        i_10_2709 <= in_reg[301];
        i_10_2710 <= in_reg[813];
        i_10_2711 <= in_reg[1325];
        i_10_2712 <= in_reg[1837];
        i_10_2713 <= in_reg[2349];
        i_10_2714 <= in_reg[2861];
        i_10_2715 <= in_reg[3373];
        i_10_2716 <= in_reg[3885];
        i_10_2717 <= in_reg[4397];
        i_10_2718 <= in_reg[302];
        i_10_2719 <= in_reg[814];
        i_10_2720 <= in_reg[1326];
        i_10_2721 <= in_reg[1838];
        i_10_2722 <= in_reg[2350];
        i_10_2723 <= in_reg[2862];
        i_10_2724 <= in_reg[3374];
        i_10_2725 <= in_reg[3886];
        i_10_2726 <= in_reg[4398];
        i_10_2727 <= in_reg[303];
        i_10_2728 <= in_reg[815];
        i_10_2729 <= in_reg[1327];
        i_10_2730 <= in_reg[1839];
        i_10_2731 <= in_reg[2351];
        i_10_2732 <= in_reg[2863];
        i_10_2733 <= in_reg[3375];
        i_10_2734 <= in_reg[3887];
        i_10_2735 <= in_reg[4399];
        i_10_2736 <= in_reg[304];
        i_10_2737 <= in_reg[816];
        i_10_2738 <= in_reg[1328];
        i_10_2739 <= in_reg[1840];
        i_10_2740 <= in_reg[2352];
        i_10_2741 <= in_reg[2864];
        i_10_2742 <= in_reg[3376];
        i_10_2743 <= in_reg[3888];
        i_10_2744 <= in_reg[4400];
        i_10_2745 <= in_reg[305];
        i_10_2746 <= in_reg[817];
        i_10_2747 <= in_reg[1329];
        i_10_2748 <= in_reg[1841];
        i_10_2749 <= in_reg[2353];
        i_10_2750 <= in_reg[2865];
        i_10_2751 <= in_reg[3377];
        i_10_2752 <= in_reg[3889];
        i_10_2753 <= in_reg[4401];
        i_10_2754 <= in_reg[306];
        i_10_2755 <= in_reg[818];
        i_10_2756 <= in_reg[1330];
        i_10_2757 <= in_reg[1842];
        i_10_2758 <= in_reg[2354];
        i_10_2759 <= in_reg[2866];
        i_10_2760 <= in_reg[3378];
        i_10_2761 <= in_reg[3890];
        i_10_2762 <= in_reg[4402];
        i_10_2763 <= in_reg[307];
        i_10_2764 <= in_reg[819];
        i_10_2765 <= in_reg[1331];
        i_10_2766 <= in_reg[1843];
        i_10_2767 <= in_reg[2355];
        i_10_2768 <= in_reg[2867];
        i_10_2769 <= in_reg[3379];
        i_10_2770 <= in_reg[3891];
        i_10_2771 <= in_reg[4403];
        i_10_2772 <= in_reg[308];
        i_10_2773 <= in_reg[820];
        i_10_2774 <= in_reg[1332];
        i_10_2775 <= in_reg[1844];
        i_10_2776 <= in_reg[2356];
        i_10_2777 <= in_reg[2868];
        i_10_2778 <= in_reg[3380];
        i_10_2779 <= in_reg[3892];
        i_10_2780 <= in_reg[4404];
        i_10_2781 <= in_reg[309];
        i_10_2782 <= in_reg[821];
        i_10_2783 <= in_reg[1333];
        i_10_2784 <= in_reg[1845];
        i_10_2785 <= in_reg[2357];
        i_10_2786 <= in_reg[2869];
        i_10_2787 <= in_reg[3381];
        i_10_2788 <= in_reg[3893];
        i_10_2789 <= in_reg[4405];
        i_10_2790 <= in_reg[310];
        i_10_2791 <= in_reg[822];
        i_10_2792 <= in_reg[1334];
        i_10_2793 <= in_reg[1846];
        i_10_2794 <= in_reg[2358];
        i_10_2795 <= in_reg[2870];
        i_10_2796 <= in_reg[3382];
        i_10_2797 <= in_reg[3894];
        i_10_2798 <= in_reg[4406];
        i_10_2799 <= in_reg[311];
        i_10_2800 <= in_reg[823];
        i_10_2801 <= in_reg[1335];
        i_10_2802 <= in_reg[1847];
        i_10_2803 <= in_reg[2359];
        i_10_2804 <= in_reg[2871];
        i_10_2805 <= in_reg[3383];
        i_10_2806 <= in_reg[3895];
        i_10_2807 <= in_reg[4407];
        i_10_2808 <= in_reg[312];
        i_10_2809 <= in_reg[824];
        i_10_2810 <= in_reg[1336];
        i_10_2811 <= in_reg[1848];
        i_10_2812 <= in_reg[2360];
        i_10_2813 <= in_reg[2872];
        i_10_2814 <= in_reg[3384];
        i_10_2815 <= in_reg[3896];
        i_10_2816 <= in_reg[4408];
        i_10_2817 <= in_reg[313];
        i_10_2818 <= in_reg[825];
        i_10_2819 <= in_reg[1337];
        i_10_2820 <= in_reg[1849];
        i_10_2821 <= in_reg[2361];
        i_10_2822 <= in_reg[2873];
        i_10_2823 <= in_reg[3385];
        i_10_2824 <= in_reg[3897];
        i_10_2825 <= in_reg[4409];
        i_10_2826 <= in_reg[314];
        i_10_2827 <= in_reg[826];
        i_10_2828 <= in_reg[1338];
        i_10_2829 <= in_reg[1850];
        i_10_2830 <= in_reg[2362];
        i_10_2831 <= in_reg[2874];
        i_10_2832 <= in_reg[3386];
        i_10_2833 <= in_reg[3898];
        i_10_2834 <= in_reg[4410];
        i_10_2835 <= in_reg[315];
        i_10_2836 <= in_reg[827];
        i_10_2837 <= in_reg[1339];
        i_10_2838 <= in_reg[1851];
        i_10_2839 <= in_reg[2363];
        i_10_2840 <= in_reg[2875];
        i_10_2841 <= in_reg[3387];
        i_10_2842 <= in_reg[3899];
        i_10_2843 <= in_reg[4411];
        i_10_2844 <= in_reg[316];
        i_10_2845 <= in_reg[828];
        i_10_2846 <= in_reg[1340];
        i_10_2847 <= in_reg[1852];
        i_10_2848 <= in_reg[2364];
        i_10_2849 <= in_reg[2876];
        i_10_2850 <= in_reg[3388];
        i_10_2851 <= in_reg[3900];
        i_10_2852 <= in_reg[4412];
        i_10_2853 <= in_reg[317];
        i_10_2854 <= in_reg[829];
        i_10_2855 <= in_reg[1341];
        i_10_2856 <= in_reg[1853];
        i_10_2857 <= in_reg[2365];
        i_10_2858 <= in_reg[2877];
        i_10_2859 <= in_reg[3389];
        i_10_2860 <= in_reg[3901];
        i_10_2861 <= in_reg[4413];
        i_10_2862 <= in_reg[318];
        i_10_2863 <= in_reg[830];
        i_10_2864 <= in_reg[1342];
        i_10_2865 <= in_reg[1854];
        i_10_2866 <= in_reg[2366];
        i_10_2867 <= in_reg[2878];
        i_10_2868 <= in_reg[3390];
        i_10_2869 <= in_reg[3902];
        i_10_2870 <= in_reg[4414];
        i_10_2871 <= in_reg[319];
        i_10_2872 <= in_reg[831];
        i_10_2873 <= in_reg[1343];
        i_10_2874 <= in_reg[1855];
        i_10_2875 <= in_reg[2367];
        i_10_2876 <= in_reg[2879];
        i_10_2877 <= in_reg[3391];
        i_10_2878 <= in_reg[3903];
        i_10_2879 <= in_reg[4415];
        i_10_2880 <= in_reg[320];
        i_10_2881 <= in_reg[832];
        i_10_2882 <= in_reg[1344];
        i_10_2883 <= in_reg[1856];
        i_10_2884 <= in_reg[2368];
        i_10_2885 <= in_reg[2880];
        i_10_2886 <= in_reg[3392];
        i_10_2887 <= in_reg[3904];
        i_10_2888 <= in_reg[4416];
        i_10_2889 <= in_reg[321];
        i_10_2890 <= in_reg[833];
        i_10_2891 <= in_reg[1345];
        i_10_2892 <= in_reg[1857];
        i_10_2893 <= in_reg[2369];
        i_10_2894 <= in_reg[2881];
        i_10_2895 <= in_reg[3393];
        i_10_2896 <= in_reg[3905];
        i_10_2897 <= in_reg[4417];
        i_10_2898 <= in_reg[322];
        i_10_2899 <= in_reg[834];
        i_10_2900 <= in_reg[1346];
        i_10_2901 <= in_reg[1858];
        i_10_2902 <= in_reg[2370];
        i_10_2903 <= in_reg[2882];
        i_10_2904 <= in_reg[3394];
        i_10_2905 <= in_reg[3906];
        i_10_2906 <= in_reg[4418];
        i_10_2907 <= in_reg[323];
        i_10_2908 <= in_reg[835];
        i_10_2909 <= in_reg[1347];
        i_10_2910 <= in_reg[1859];
        i_10_2911 <= in_reg[2371];
        i_10_2912 <= in_reg[2883];
        i_10_2913 <= in_reg[3395];
        i_10_2914 <= in_reg[3907];
        i_10_2915 <= in_reg[4419];
        i_10_2916 <= in_reg[324];
        i_10_2917 <= in_reg[836];
        i_10_2918 <= in_reg[1348];
        i_10_2919 <= in_reg[1860];
        i_10_2920 <= in_reg[2372];
        i_10_2921 <= in_reg[2884];
        i_10_2922 <= in_reg[3396];
        i_10_2923 <= in_reg[3908];
        i_10_2924 <= in_reg[4420];
        i_10_2925 <= in_reg[325];
        i_10_2926 <= in_reg[837];
        i_10_2927 <= in_reg[1349];
        i_10_2928 <= in_reg[1861];
        i_10_2929 <= in_reg[2373];
        i_10_2930 <= in_reg[2885];
        i_10_2931 <= in_reg[3397];
        i_10_2932 <= in_reg[3909];
        i_10_2933 <= in_reg[4421];
        i_10_2934 <= in_reg[326];
        i_10_2935 <= in_reg[838];
        i_10_2936 <= in_reg[1350];
        i_10_2937 <= in_reg[1862];
        i_10_2938 <= in_reg[2374];
        i_10_2939 <= in_reg[2886];
        i_10_2940 <= in_reg[3398];
        i_10_2941 <= in_reg[3910];
        i_10_2942 <= in_reg[4422];
        i_10_2943 <= in_reg[327];
        i_10_2944 <= in_reg[839];
        i_10_2945 <= in_reg[1351];
        i_10_2946 <= in_reg[1863];
        i_10_2947 <= in_reg[2375];
        i_10_2948 <= in_reg[2887];
        i_10_2949 <= in_reg[3399];
        i_10_2950 <= in_reg[3911];
        i_10_2951 <= in_reg[4423];
        i_10_2952 <= in_reg[328];
        i_10_2953 <= in_reg[840];
        i_10_2954 <= in_reg[1352];
        i_10_2955 <= in_reg[1864];
        i_10_2956 <= in_reg[2376];
        i_10_2957 <= in_reg[2888];
        i_10_2958 <= in_reg[3400];
        i_10_2959 <= in_reg[3912];
        i_10_2960 <= in_reg[4424];
        i_10_2961 <= in_reg[329];
        i_10_2962 <= in_reg[841];
        i_10_2963 <= in_reg[1353];
        i_10_2964 <= in_reg[1865];
        i_10_2965 <= in_reg[2377];
        i_10_2966 <= in_reg[2889];
        i_10_2967 <= in_reg[3401];
        i_10_2968 <= in_reg[3913];
        i_10_2969 <= in_reg[4425];
        i_10_2970 <= in_reg[330];
        i_10_2971 <= in_reg[842];
        i_10_2972 <= in_reg[1354];
        i_10_2973 <= in_reg[1866];
        i_10_2974 <= in_reg[2378];
        i_10_2975 <= in_reg[2890];
        i_10_2976 <= in_reg[3402];
        i_10_2977 <= in_reg[3914];
        i_10_2978 <= in_reg[4426];
        i_10_2979 <= in_reg[331];
        i_10_2980 <= in_reg[843];
        i_10_2981 <= in_reg[1355];
        i_10_2982 <= in_reg[1867];
        i_10_2983 <= in_reg[2379];
        i_10_2984 <= in_reg[2891];
        i_10_2985 <= in_reg[3403];
        i_10_2986 <= in_reg[3915];
        i_10_2987 <= in_reg[4427];
        i_10_2988 <= in_reg[332];
        i_10_2989 <= in_reg[844];
        i_10_2990 <= in_reg[1356];
        i_10_2991 <= in_reg[1868];
        i_10_2992 <= in_reg[2380];
        i_10_2993 <= in_reg[2892];
        i_10_2994 <= in_reg[3404];
        i_10_2995 <= in_reg[3916];
        i_10_2996 <= in_reg[4428];
        i_10_2997 <= in_reg[333];
        i_10_2998 <= in_reg[845];
        i_10_2999 <= in_reg[1357];
        i_10_3000 <= in_reg[1869];
        i_10_3001 <= in_reg[2381];
        i_10_3002 <= in_reg[2893];
        i_10_3003 <= in_reg[3405];
        i_10_3004 <= in_reg[3917];
        i_10_3005 <= in_reg[4429];
        i_10_3006 <= in_reg[334];
        i_10_3007 <= in_reg[846];
        i_10_3008 <= in_reg[1358];
        i_10_3009 <= in_reg[1870];
        i_10_3010 <= in_reg[2382];
        i_10_3011 <= in_reg[2894];
        i_10_3012 <= in_reg[3406];
        i_10_3013 <= in_reg[3918];
        i_10_3014 <= in_reg[4430];
        i_10_3015 <= in_reg[335];
        i_10_3016 <= in_reg[847];
        i_10_3017 <= in_reg[1359];
        i_10_3018 <= in_reg[1871];
        i_10_3019 <= in_reg[2383];
        i_10_3020 <= in_reg[2895];
        i_10_3021 <= in_reg[3407];
        i_10_3022 <= in_reg[3919];
        i_10_3023 <= in_reg[4431];
        i_10_3024 <= in_reg[336];
        i_10_3025 <= in_reg[848];
        i_10_3026 <= in_reg[1360];
        i_10_3027 <= in_reg[1872];
        i_10_3028 <= in_reg[2384];
        i_10_3029 <= in_reg[2896];
        i_10_3030 <= in_reg[3408];
        i_10_3031 <= in_reg[3920];
        i_10_3032 <= in_reg[4432];
        i_10_3033 <= in_reg[337];
        i_10_3034 <= in_reg[849];
        i_10_3035 <= in_reg[1361];
        i_10_3036 <= in_reg[1873];
        i_10_3037 <= in_reg[2385];
        i_10_3038 <= in_reg[2897];
        i_10_3039 <= in_reg[3409];
        i_10_3040 <= in_reg[3921];
        i_10_3041 <= in_reg[4433];
        i_10_3042 <= in_reg[338];
        i_10_3043 <= in_reg[850];
        i_10_3044 <= in_reg[1362];
        i_10_3045 <= in_reg[1874];
        i_10_3046 <= in_reg[2386];
        i_10_3047 <= in_reg[2898];
        i_10_3048 <= in_reg[3410];
        i_10_3049 <= in_reg[3922];
        i_10_3050 <= in_reg[4434];
        i_10_3051 <= in_reg[339];
        i_10_3052 <= in_reg[851];
        i_10_3053 <= in_reg[1363];
        i_10_3054 <= in_reg[1875];
        i_10_3055 <= in_reg[2387];
        i_10_3056 <= in_reg[2899];
        i_10_3057 <= in_reg[3411];
        i_10_3058 <= in_reg[3923];
        i_10_3059 <= in_reg[4435];
        i_10_3060 <= in_reg[340];
        i_10_3061 <= in_reg[852];
        i_10_3062 <= in_reg[1364];
        i_10_3063 <= in_reg[1876];
        i_10_3064 <= in_reg[2388];
        i_10_3065 <= in_reg[2900];
        i_10_3066 <= in_reg[3412];
        i_10_3067 <= in_reg[3924];
        i_10_3068 <= in_reg[4436];
        i_10_3069 <= in_reg[341];
        i_10_3070 <= in_reg[853];
        i_10_3071 <= in_reg[1365];
        i_10_3072 <= in_reg[1877];
        i_10_3073 <= in_reg[2389];
        i_10_3074 <= in_reg[2901];
        i_10_3075 <= in_reg[3413];
        i_10_3076 <= in_reg[3925];
        i_10_3077 <= in_reg[4437];
        i_10_3078 <= in_reg[342];
        i_10_3079 <= in_reg[854];
        i_10_3080 <= in_reg[1366];
        i_10_3081 <= in_reg[1878];
        i_10_3082 <= in_reg[2390];
        i_10_3083 <= in_reg[2902];
        i_10_3084 <= in_reg[3414];
        i_10_3085 <= in_reg[3926];
        i_10_3086 <= in_reg[4438];
        i_10_3087 <= in_reg[343];
        i_10_3088 <= in_reg[855];
        i_10_3089 <= in_reg[1367];
        i_10_3090 <= in_reg[1879];
        i_10_3091 <= in_reg[2391];
        i_10_3092 <= in_reg[2903];
        i_10_3093 <= in_reg[3415];
        i_10_3094 <= in_reg[3927];
        i_10_3095 <= in_reg[4439];
        i_10_3096 <= in_reg[344];
        i_10_3097 <= in_reg[856];
        i_10_3098 <= in_reg[1368];
        i_10_3099 <= in_reg[1880];
        i_10_3100 <= in_reg[2392];
        i_10_3101 <= in_reg[2904];
        i_10_3102 <= in_reg[3416];
        i_10_3103 <= in_reg[3928];
        i_10_3104 <= in_reg[4440];
        i_10_3105 <= in_reg[345];
        i_10_3106 <= in_reg[857];
        i_10_3107 <= in_reg[1369];
        i_10_3108 <= in_reg[1881];
        i_10_3109 <= in_reg[2393];
        i_10_3110 <= in_reg[2905];
        i_10_3111 <= in_reg[3417];
        i_10_3112 <= in_reg[3929];
        i_10_3113 <= in_reg[4441];
        i_10_3114 <= in_reg[346];
        i_10_3115 <= in_reg[858];
        i_10_3116 <= in_reg[1370];
        i_10_3117 <= in_reg[1882];
        i_10_3118 <= in_reg[2394];
        i_10_3119 <= in_reg[2906];
        i_10_3120 <= in_reg[3418];
        i_10_3121 <= in_reg[3930];
        i_10_3122 <= in_reg[4442];
        i_10_3123 <= in_reg[347];
        i_10_3124 <= in_reg[859];
        i_10_3125 <= in_reg[1371];
        i_10_3126 <= in_reg[1883];
        i_10_3127 <= in_reg[2395];
        i_10_3128 <= in_reg[2907];
        i_10_3129 <= in_reg[3419];
        i_10_3130 <= in_reg[3931];
        i_10_3131 <= in_reg[4443];
        i_10_3132 <= in_reg[348];
        i_10_3133 <= in_reg[860];
        i_10_3134 <= in_reg[1372];
        i_10_3135 <= in_reg[1884];
        i_10_3136 <= in_reg[2396];
        i_10_3137 <= in_reg[2908];
        i_10_3138 <= in_reg[3420];
        i_10_3139 <= in_reg[3932];
        i_10_3140 <= in_reg[4444];
        i_10_3141 <= in_reg[349];
        i_10_3142 <= in_reg[861];
        i_10_3143 <= in_reg[1373];
        i_10_3144 <= in_reg[1885];
        i_10_3145 <= in_reg[2397];
        i_10_3146 <= in_reg[2909];
        i_10_3147 <= in_reg[3421];
        i_10_3148 <= in_reg[3933];
        i_10_3149 <= in_reg[4445];
        i_10_3150 <= in_reg[350];
        i_10_3151 <= in_reg[862];
        i_10_3152 <= in_reg[1374];
        i_10_3153 <= in_reg[1886];
        i_10_3154 <= in_reg[2398];
        i_10_3155 <= in_reg[2910];
        i_10_3156 <= in_reg[3422];
        i_10_3157 <= in_reg[3934];
        i_10_3158 <= in_reg[4446];
        i_10_3159 <= in_reg[351];
        i_10_3160 <= in_reg[863];
        i_10_3161 <= in_reg[1375];
        i_10_3162 <= in_reg[1887];
        i_10_3163 <= in_reg[2399];
        i_10_3164 <= in_reg[2911];
        i_10_3165 <= in_reg[3423];
        i_10_3166 <= in_reg[3935];
        i_10_3167 <= in_reg[4447];
        i_10_3168 <= in_reg[352];
        i_10_3169 <= in_reg[864];
        i_10_3170 <= in_reg[1376];
        i_10_3171 <= in_reg[1888];
        i_10_3172 <= in_reg[2400];
        i_10_3173 <= in_reg[2912];
        i_10_3174 <= in_reg[3424];
        i_10_3175 <= in_reg[3936];
        i_10_3176 <= in_reg[4448];
        i_10_3177 <= in_reg[353];
        i_10_3178 <= in_reg[865];
        i_10_3179 <= in_reg[1377];
        i_10_3180 <= in_reg[1889];
        i_10_3181 <= in_reg[2401];
        i_10_3182 <= in_reg[2913];
        i_10_3183 <= in_reg[3425];
        i_10_3184 <= in_reg[3937];
        i_10_3185 <= in_reg[4449];
        i_10_3186 <= in_reg[354];
        i_10_3187 <= in_reg[866];
        i_10_3188 <= in_reg[1378];
        i_10_3189 <= in_reg[1890];
        i_10_3190 <= in_reg[2402];
        i_10_3191 <= in_reg[2914];
        i_10_3192 <= in_reg[3426];
        i_10_3193 <= in_reg[3938];
        i_10_3194 <= in_reg[4450];
        i_10_3195 <= in_reg[355];
        i_10_3196 <= in_reg[867];
        i_10_3197 <= in_reg[1379];
        i_10_3198 <= in_reg[1891];
        i_10_3199 <= in_reg[2403];
        i_10_3200 <= in_reg[2915];
        i_10_3201 <= in_reg[3427];
        i_10_3202 <= in_reg[3939];
        i_10_3203 <= in_reg[4451];
        i_10_3204 <= in_reg[356];
        i_10_3205 <= in_reg[868];
        i_10_3206 <= in_reg[1380];
        i_10_3207 <= in_reg[1892];
        i_10_3208 <= in_reg[2404];
        i_10_3209 <= in_reg[2916];
        i_10_3210 <= in_reg[3428];
        i_10_3211 <= in_reg[3940];
        i_10_3212 <= in_reg[4452];
        i_10_3213 <= in_reg[357];
        i_10_3214 <= in_reg[869];
        i_10_3215 <= in_reg[1381];
        i_10_3216 <= in_reg[1893];
        i_10_3217 <= in_reg[2405];
        i_10_3218 <= in_reg[2917];
        i_10_3219 <= in_reg[3429];
        i_10_3220 <= in_reg[3941];
        i_10_3221 <= in_reg[4453];
        i_10_3222 <= in_reg[358];
        i_10_3223 <= in_reg[870];
        i_10_3224 <= in_reg[1382];
        i_10_3225 <= in_reg[1894];
        i_10_3226 <= in_reg[2406];
        i_10_3227 <= in_reg[2918];
        i_10_3228 <= in_reg[3430];
        i_10_3229 <= in_reg[3942];
        i_10_3230 <= in_reg[4454];
        i_10_3231 <= in_reg[359];
        i_10_3232 <= in_reg[871];
        i_10_3233 <= in_reg[1383];
        i_10_3234 <= in_reg[1895];
        i_10_3235 <= in_reg[2407];
        i_10_3236 <= in_reg[2919];
        i_10_3237 <= in_reg[3431];
        i_10_3238 <= in_reg[3943];
        i_10_3239 <= in_reg[4455];
        i_10_3240 <= in_reg[360];
        i_10_3241 <= in_reg[872];
        i_10_3242 <= in_reg[1384];
        i_10_3243 <= in_reg[1896];
        i_10_3244 <= in_reg[2408];
        i_10_3245 <= in_reg[2920];
        i_10_3246 <= in_reg[3432];
        i_10_3247 <= in_reg[3944];
        i_10_3248 <= in_reg[4456];
        i_10_3249 <= in_reg[361];
        i_10_3250 <= in_reg[873];
        i_10_3251 <= in_reg[1385];
        i_10_3252 <= in_reg[1897];
        i_10_3253 <= in_reg[2409];
        i_10_3254 <= in_reg[2921];
        i_10_3255 <= in_reg[3433];
        i_10_3256 <= in_reg[3945];
        i_10_3257 <= in_reg[4457];
        i_10_3258 <= in_reg[362];
        i_10_3259 <= in_reg[874];
        i_10_3260 <= in_reg[1386];
        i_10_3261 <= in_reg[1898];
        i_10_3262 <= in_reg[2410];
        i_10_3263 <= in_reg[2922];
        i_10_3264 <= in_reg[3434];
        i_10_3265 <= in_reg[3946];
        i_10_3266 <= in_reg[4458];
        i_10_3267 <= in_reg[363];
        i_10_3268 <= in_reg[875];
        i_10_3269 <= in_reg[1387];
        i_10_3270 <= in_reg[1899];
        i_10_3271 <= in_reg[2411];
        i_10_3272 <= in_reg[2923];
        i_10_3273 <= in_reg[3435];
        i_10_3274 <= in_reg[3947];
        i_10_3275 <= in_reg[4459];
        i_10_3276 <= in_reg[364];
        i_10_3277 <= in_reg[876];
        i_10_3278 <= in_reg[1388];
        i_10_3279 <= in_reg[1900];
        i_10_3280 <= in_reg[2412];
        i_10_3281 <= in_reg[2924];
        i_10_3282 <= in_reg[3436];
        i_10_3283 <= in_reg[3948];
        i_10_3284 <= in_reg[4460];
        i_10_3285 <= in_reg[365];
        i_10_3286 <= in_reg[877];
        i_10_3287 <= in_reg[1389];
        i_10_3288 <= in_reg[1901];
        i_10_3289 <= in_reg[2413];
        i_10_3290 <= in_reg[2925];
        i_10_3291 <= in_reg[3437];
        i_10_3292 <= in_reg[3949];
        i_10_3293 <= in_reg[4461];
        i_10_3294 <= in_reg[366];
        i_10_3295 <= in_reg[878];
        i_10_3296 <= in_reg[1390];
        i_10_3297 <= in_reg[1902];
        i_10_3298 <= in_reg[2414];
        i_10_3299 <= in_reg[2926];
        i_10_3300 <= in_reg[3438];
        i_10_3301 <= in_reg[3950];
        i_10_3302 <= in_reg[4462];
        i_10_3303 <= in_reg[367];
        i_10_3304 <= in_reg[879];
        i_10_3305 <= in_reg[1391];
        i_10_3306 <= in_reg[1903];
        i_10_3307 <= in_reg[2415];
        i_10_3308 <= in_reg[2927];
        i_10_3309 <= in_reg[3439];
        i_10_3310 <= in_reg[3951];
        i_10_3311 <= in_reg[4463];
        i_10_3312 <= in_reg[368];
        i_10_3313 <= in_reg[880];
        i_10_3314 <= in_reg[1392];
        i_10_3315 <= in_reg[1904];
        i_10_3316 <= in_reg[2416];
        i_10_3317 <= in_reg[2928];
        i_10_3318 <= in_reg[3440];
        i_10_3319 <= in_reg[3952];
        i_10_3320 <= in_reg[4464];
        i_10_3321 <= in_reg[369];
        i_10_3322 <= in_reg[881];
        i_10_3323 <= in_reg[1393];
        i_10_3324 <= in_reg[1905];
        i_10_3325 <= in_reg[2417];
        i_10_3326 <= in_reg[2929];
        i_10_3327 <= in_reg[3441];
        i_10_3328 <= in_reg[3953];
        i_10_3329 <= in_reg[4465];
        i_10_3330 <= in_reg[370];
        i_10_3331 <= in_reg[882];
        i_10_3332 <= in_reg[1394];
        i_10_3333 <= in_reg[1906];
        i_10_3334 <= in_reg[2418];
        i_10_3335 <= in_reg[2930];
        i_10_3336 <= in_reg[3442];
        i_10_3337 <= in_reg[3954];
        i_10_3338 <= in_reg[4466];
        i_10_3339 <= in_reg[371];
        i_10_3340 <= in_reg[883];
        i_10_3341 <= in_reg[1395];
        i_10_3342 <= in_reg[1907];
        i_10_3343 <= in_reg[2419];
        i_10_3344 <= in_reg[2931];
        i_10_3345 <= in_reg[3443];
        i_10_3346 <= in_reg[3955];
        i_10_3347 <= in_reg[4467];
        i_10_3348 <= in_reg[372];
        i_10_3349 <= in_reg[884];
        i_10_3350 <= in_reg[1396];
        i_10_3351 <= in_reg[1908];
        i_10_3352 <= in_reg[2420];
        i_10_3353 <= in_reg[2932];
        i_10_3354 <= in_reg[3444];
        i_10_3355 <= in_reg[3956];
        i_10_3356 <= in_reg[4468];
        i_10_3357 <= in_reg[373];
        i_10_3358 <= in_reg[885];
        i_10_3359 <= in_reg[1397];
        i_10_3360 <= in_reg[1909];
        i_10_3361 <= in_reg[2421];
        i_10_3362 <= in_reg[2933];
        i_10_3363 <= in_reg[3445];
        i_10_3364 <= in_reg[3957];
        i_10_3365 <= in_reg[4469];
        i_10_3366 <= in_reg[374];
        i_10_3367 <= in_reg[886];
        i_10_3368 <= in_reg[1398];
        i_10_3369 <= in_reg[1910];
        i_10_3370 <= in_reg[2422];
        i_10_3371 <= in_reg[2934];
        i_10_3372 <= in_reg[3446];
        i_10_3373 <= in_reg[3958];
        i_10_3374 <= in_reg[4470];
        i_10_3375 <= in_reg[375];
        i_10_3376 <= in_reg[887];
        i_10_3377 <= in_reg[1399];
        i_10_3378 <= in_reg[1911];
        i_10_3379 <= in_reg[2423];
        i_10_3380 <= in_reg[2935];
        i_10_3381 <= in_reg[3447];
        i_10_3382 <= in_reg[3959];
        i_10_3383 <= in_reg[4471];
        i_10_3384 <= in_reg[376];
        i_10_3385 <= in_reg[888];
        i_10_3386 <= in_reg[1400];
        i_10_3387 <= in_reg[1912];
        i_10_3388 <= in_reg[2424];
        i_10_3389 <= in_reg[2936];
        i_10_3390 <= in_reg[3448];
        i_10_3391 <= in_reg[3960];
        i_10_3392 <= in_reg[4472];
        i_10_3393 <= in_reg[377];
        i_10_3394 <= in_reg[889];
        i_10_3395 <= in_reg[1401];
        i_10_3396 <= in_reg[1913];
        i_10_3397 <= in_reg[2425];
        i_10_3398 <= in_reg[2937];
        i_10_3399 <= in_reg[3449];
        i_10_3400 <= in_reg[3961];
        i_10_3401 <= in_reg[4473];
        i_10_3402 <= in_reg[378];
        i_10_3403 <= in_reg[890];
        i_10_3404 <= in_reg[1402];
        i_10_3405 <= in_reg[1914];
        i_10_3406 <= in_reg[2426];
        i_10_3407 <= in_reg[2938];
        i_10_3408 <= in_reg[3450];
        i_10_3409 <= in_reg[3962];
        i_10_3410 <= in_reg[4474];
        i_10_3411 <= in_reg[379];
        i_10_3412 <= in_reg[891];
        i_10_3413 <= in_reg[1403];
        i_10_3414 <= in_reg[1915];
        i_10_3415 <= in_reg[2427];
        i_10_3416 <= in_reg[2939];
        i_10_3417 <= in_reg[3451];
        i_10_3418 <= in_reg[3963];
        i_10_3419 <= in_reg[4475];
        i_10_3420 <= in_reg[380];
        i_10_3421 <= in_reg[892];
        i_10_3422 <= in_reg[1404];
        i_10_3423 <= in_reg[1916];
        i_10_3424 <= in_reg[2428];
        i_10_3425 <= in_reg[2940];
        i_10_3426 <= in_reg[3452];
        i_10_3427 <= in_reg[3964];
        i_10_3428 <= in_reg[4476];
        i_10_3429 <= in_reg[381];
        i_10_3430 <= in_reg[893];
        i_10_3431 <= in_reg[1405];
        i_10_3432 <= in_reg[1917];
        i_10_3433 <= in_reg[2429];
        i_10_3434 <= in_reg[2941];
        i_10_3435 <= in_reg[3453];
        i_10_3436 <= in_reg[3965];
        i_10_3437 <= in_reg[4477];
        i_10_3438 <= in_reg[382];
        i_10_3439 <= in_reg[894];
        i_10_3440 <= in_reg[1406];
        i_10_3441 <= in_reg[1918];
        i_10_3442 <= in_reg[2430];
        i_10_3443 <= in_reg[2942];
        i_10_3444 <= in_reg[3454];
        i_10_3445 <= in_reg[3966];
        i_10_3446 <= in_reg[4478];
        i_10_3447 <= in_reg[383];
        i_10_3448 <= in_reg[895];
        i_10_3449 <= in_reg[1407];
        i_10_3450 <= in_reg[1919];
        i_10_3451 <= in_reg[2431];
        i_10_3452 <= in_reg[2943];
        i_10_3453 <= in_reg[3455];
        i_10_3454 <= in_reg[3967];
        i_10_3455 <= in_reg[4479];
        i_10_3456 <= in_reg[384];
        i_10_3457 <= in_reg[896];
        i_10_3458 <= in_reg[1408];
        i_10_3459 <= in_reg[1920];
        i_10_3460 <= in_reg[2432];
        i_10_3461 <= in_reg[2944];
        i_10_3462 <= in_reg[3456];
        i_10_3463 <= in_reg[3968];
        i_10_3464 <= in_reg[4480];
        i_10_3465 <= in_reg[385];
        i_10_3466 <= in_reg[897];
        i_10_3467 <= in_reg[1409];
        i_10_3468 <= in_reg[1921];
        i_10_3469 <= in_reg[2433];
        i_10_3470 <= in_reg[2945];
        i_10_3471 <= in_reg[3457];
        i_10_3472 <= in_reg[3969];
        i_10_3473 <= in_reg[4481];
        i_10_3474 <= in_reg[386];
        i_10_3475 <= in_reg[898];
        i_10_3476 <= in_reg[1410];
        i_10_3477 <= in_reg[1922];
        i_10_3478 <= in_reg[2434];
        i_10_3479 <= in_reg[2946];
        i_10_3480 <= in_reg[3458];
        i_10_3481 <= in_reg[3970];
        i_10_3482 <= in_reg[4482];
        i_10_3483 <= in_reg[387];
        i_10_3484 <= in_reg[899];
        i_10_3485 <= in_reg[1411];
        i_10_3486 <= in_reg[1923];
        i_10_3487 <= in_reg[2435];
        i_10_3488 <= in_reg[2947];
        i_10_3489 <= in_reg[3459];
        i_10_3490 <= in_reg[3971];
        i_10_3491 <= in_reg[4483];
        i_10_3492 <= in_reg[388];
        i_10_3493 <= in_reg[900];
        i_10_3494 <= in_reg[1412];
        i_10_3495 <= in_reg[1924];
        i_10_3496 <= in_reg[2436];
        i_10_3497 <= in_reg[2948];
        i_10_3498 <= in_reg[3460];
        i_10_3499 <= in_reg[3972];
        i_10_3500 <= in_reg[4484];
        i_10_3501 <= in_reg[389];
        i_10_3502 <= in_reg[901];
        i_10_3503 <= in_reg[1413];
        i_10_3504 <= in_reg[1925];
        i_10_3505 <= in_reg[2437];
        i_10_3506 <= in_reg[2949];
        i_10_3507 <= in_reg[3461];
        i_10_3508 <= in_reg[3973];
        i_10_3509 <= in_reg[4485];
        i_10_3510 <= in_reg[390];
        i_10_3511 <= in_reg[902];
        i_10_3512 <= in_reg[1414];
        i_10_3513 <= in_reg[1926];
        i_10_3514 <= in_reg[2438];
        i_10_3515 <= in_reg[2950];
        i_10_3516 <= in_reg[3462];
        i_10_3517 <= in_reg[3974];
        i_10_3518 <= in_reg[4486];
        i_10_3519 <= in_reg[391];
        i_10_3520 <= in_reg[903];
        i_10_3521 <= in_reg[1415];
        i_10_3522 <= in_reg[1927];
        i_10_3523 <= in_reg[2439];
        i_10_3524 <= in_reg[2951];
        i_10_3525 <= in_reg[3463];
        i_10_3526 <= in_reg[3975];
        i_10_3527 <= in_reg[4487];
        i_10_3528 <= in_reg[392];
        i_10_3529 <= in_reg[904];
        i_10_3530 <= in_reg[1416];
        i_10_3531 <= in_reg[1928];
        i_10_3532 <= in_reg[2440];
        i_10_3533 <= in_reg[2952];
        i_10_3534 <= in_reg[3464];
        i_10_3535 <= in_reg[3976];
        i_10_3536 <= in_reg[4488];
        i_10_3537 <= in_reg[393];
        i_10_3538 <= in_reg[905];
        i_10_3539 <= in_reg[1417];
        i_10_3540 <= in_reg[1929];
        i_10_3541 <= in_reg[2441];
        i_10_3542 <= in_reg[2953];
        i_10_3543 <= in_reg[3465];
        i_10_3544 <= in_reg[3977];
        i_10_3545 <= in_reg[4489];
        i_10_3546 <= in_reg[394];
        i_10_3547 <= in_reg[906];
        i_10_3548 <= in_reg[1418];
        i_10_3549 <= in_reg[1930];
        i_10_3550 <= in_reg[2442];
        i_10_3551 <= in_reg[2954];
        i_10_3552 <= in_reg[3466];
        i_10_3553 <= in_reg[3978];
        i_10_3554 <= in_reg[4490];
        i_10_3555 <= in_reg[395];
        i_10_3556 <= in_reg[907];
        i_10_3557 <= in_reg[1419];
        i_10_3558 <= in_reg[1931];
        i_10_3559 <= in_reg[2443];
        i_10_3560 <= in_reg[2955];
        i_10_3561 <= in_reg[3467];
        i_10_3562 <= in_reg[3979];
        i_10_3563 <= in_reg[4491];
        i_10_3564 <= in_reg[396];
        i_10_3565 <= in_reg[908];
        i_10_3566 <= in_reg[1420];
        i_10_3567 <= in_reg[1932];
        i_10_3568 <= in_reg[2444];
        i_10_3569 <= in_reg[2956];
        i_10_3570 <= in_reg[3468];
        i_10_3571 <= in_reg[3980];
        i_10_3572 <= in_reg[4492];
        i_10_3573 <= in_reg[397];
        i_10_3574 <= in_reg[909];
        i_10_3575 <= in_reg[1421];
        i_10_3576 <= in_reg[1933];
        i_10_3577 <= in_reg[2445];
        i_10_3578 <= in_reg[2957];
        i_10_3579 <= in_reg[3469];
        i_10_3580 <= in_reg[3981];
        i_10_3581 <= in_reg[4493];
        i_10_3582 <= in_reg[398];
        i_10_3583 <= in_reg[910];
        i_10_3584 <= in_reg[1422];
        i_10_3585 <= in_reg[1934];
        i_10_3586 <= in_reg[2446];
        i_10_3587 <= in_reg[2958];
        i_10_3588 <= in_reg[3470];
        i_10_3589 <= in_reg[3982];
        i_10_3590 <= in_reg[4494];
        i_10_3591 <= in_reg[399];
        i_10_3592 <= in_reg[911];
        i_10_3593 <= in_reg[1423];
        i_10_3594 <= in_reg[1935];
        i_10_3595 <= in_reg[2447];
        i_10_3596 <= in_reg[2959];
        i_10_3597 <= in_reg[3471];
        i_10_3598 <= in_reg[3983];
        i_10_3599 <= in_reg[4495];
        i_10_3600 <= in_reg[400];
        i_10_3601 <= in_reg[912];
        i_10_3602 <= in_reg[1424];
        i_10_3603 <= in_reg[1936];
        i_10_3604 <= in_reg[2448];
        i_10_3605 <= in_reg[2960];
        i_10_3606 <= in_reg[3472];
        i_10_3607 <= in_reg[3984];
        i_10_3608 <= in_reg[4496];
        i_10_3609 <= in_reg[401];
        i_10_3610 <= in_reg[913];
        i_10_3611 <= in_reg[1425];
        i_10_3612 <= in_reg[1937];
        i_10_3613 <= in_reg[2449];
        i_10_3614 <= in_reg[2961];
        i_10_3615 <= in_reg[3473];
        i_10_3616 <= in_reg[3985];
        i_10_3617 <= in_reg[4497];
        i_10_3618 <= in_reg[402];
        i_10_3619 <= in_reg[914];
        i_10_3620 <= in_reg[1426];
        i_10_3621 <= in_reg[1938];
        i_10_3622 <= in_reg[2450];
        i_10_3623 <= in_reg[2962];
        i_10_3624 <= in_reg[3474];
        i_10_3625 <= in_reg[3986];
        i_10_3626 <= in_reg[4498];
        i_10_3627 <= in_reg[403];
        i_10_3628 <= in_reg[915];
        i_10_3629 <= in_reg[1427];
        i_10_3630 <= in_reg[1939];
        i_10_3631 <= in_reg[2451];
        i_10_3632 <= in_reg[2963];
        i_10_3633 <= in_reg[3475];
        i_10_3634 <= in_reg[3987];
        i_10_3635 <= in_reg[4499];
        i_10_3636 <= in_reg[404];
        i_10_3637 <= in_reg[916];
        i_10_3638 <= in_reg[1428];
        i_10_3639 <= in_reg[1940];
        i_10_3640 <= in_reg[2452];
        i_10_3641 <= in_reg[2964];
        i_10_3642 <= in_reg[3476];
        i_10_3643 <= in_reg[3988];
        i_10_3644 <= in_reg[4500];
        i_10_3645 <= in_reg[405];
        i_10_3646 <= in_reg[917];
        i_10_3647 <= in_reg[1429];
        i_10_3648 <= in_reg[1941];
        i_10_3649 <= in_reg[2453];
        i_10_3650 <= in_reg[2965];
        i_10_3651 <= in_reg[3477];
        i_10_3652 <= in_reg[3989];
        i_10_3653 <= in_reg[4501];
        i_10_3654 <= in_reg[406];
        i_10_3655 <= in_reg[918];
        i_10_3656 <= in_reg[1430];
        i_10_3657 <= in_reg[1942];
        i_10_3658 <= in_reg[2454];
        i_10_3659 <= in_reg[2966];
        i_10_3660 <= in_reg[3478];
        i_10_3661 <= in_reg[3990];
        i_10_3662 <= in_reg[4502];
        i_10_3663 <= in_reg[407];
        i_10_3664 <= in_reg[919];
        i_10_3665 <= in_reg[1431];
        i_10_3666 <= in_reg[1943];
        i_10_3667 <= in_reg[2455];
        i_10_3668 <= in_reg[2967];
        i_10_3669 <= in_reg[3479];
        i_10_3670 <= in_reg[3991];
        i_10_3671 <= in_reg[4503];
        i_10_3672 <= in_reg[408];
        i_10_3673 <= in_reg[920];
        i_10_3674 <= in_reg[1432];
        i_10_3675 <= in_reg[1944];
        i_10_3676 <= in_reg[2456];
        i_10_3677 <= in_reg[2968];
        i_10_3678 <= in_reg[3480];
        i_10_3679 <= in_reg[3992];
        i_10_3680 <= in_reg[4504];
        i_10_3681 <= in_reg[409];
        i_10_3682 <= in_reg[921];
        i_10_3683 <= in_reg[1433];
        i_10_3684 <= in_reg[1945];
        i_10_3685 <= in_reg[2457];
        i_10_3686 <= in_reg[2969];
        i_10_3687 <= in_reg[3481];
        i_10_3688 <= in_reg[3993];
        i_10_3689 <= in_reg[4505];
        i_10_3690 <= in_reg[410];
        i_10_3691 <= in_reg[922];
        i_10_3692 <= in_reg[1434];
        i_10_3693 <= in_reg[1946];
        i_10_3694 <= in_reg[2458];
        i_10_3695 <= in_reg[2970];
        i_10_3696 <= in_reg[3482];
        i_10_3697 <= in_reg[3994];
        i_10_3698 <= in_reg[4506];
        i_10_3699 <= in_reg[411];
        i_10_3700 <= in_reg[923];
        i_10_3701 <= in_reg[1435];
        i_10_3702 <= in_reg[1947];
        i_10_3703 <= in_reg[2459];
        i_10_3704 <= in_reg[2971];
        i_10_3705 <= in_reg[3483];
        i_10_3706 <= in_reg[3995];
        i_10_3707 <= in_reg[4507];
        i_10_3708 <= in_reg[412];
        i_10_3709 <= in_reg[924];
        i_10_3710 <= in_reg[1436];
        i_10_3711 <= in_reg[1948];
        i_10_3712 <= in_reg[2460];
        i_10_3713 <= in_reg[2972];
        i_10_3714 <= in_reg[3484];
        i_10_3715 <= in_reg[3996];
        i_10_3716 <= in_reg[4508];
        i_10_3717 <= in_reg[413];
        i_10_3718 <= in_reg[925];
        i_10_3719 <= in_reg[1437];
        i_10_3720 <= in_reg[1949];
        i_10_3721 <= in_reg[2461];
        i_10_3722 <= in_reg[2973];
        i_10_3723 <= in_reg[3485];
        i_10_3724 <= in_reg[3997];
        i_10_3725 <= in_reg[4509];
        i_10_3726 <= in_reg[414];
        i_10_3727 <= in_reg[926];
        i_10_3728 <= in_reg[1438];
        i_10_3729 <= in_reg[1950];
        i_10_3730 <= in_reg[2462];
        i_10_3731 <= in_reg[2974];
        i_10_3732 <= in_reg[3486];
        i_10_3733 <= in_reg[3998];
        i_10_3734 <= in_reg[4510];
        i_10_3735 <= in_reg[415];
        i_10_3736 <= in_reg[927];
        i_10_3737 <= in_reg[1439];
        i_10_3738 <= in_reg[1951];
        i_10_3739 <= in_reg[2463];
        i_10_3740 <= in_reg[2975];
        i_10_3741 <= in_reg[3487];
        i_10_3742 <= in_reg[3999];
        i_10_3743 <= in_reg[4511];
        i_10_3744 <= in_reg[416];
        i_10_3745 <= in_reg[928];
        i_10_3746 <= in_reg[1440];
        i_10_3747 <= in_reg[1952];
        i_10_3748 <= in_reg[2464];
        i_10_3749 <= in_reg[2976];
        i_10_3750 <= in_reg[3488];
        i_10_3751 <= in_reg[4000];
        i_10_3752 <= in_reg[4512];
        i_10_3753 <= in_reg[417];
        i_10_3754 <= in_reg[929];
        i_10_3755 <= in_reg[1441];
        i_10_3756 <= in_reg[1953];
        i_10_3757 <= in_reg[2465];
        i_10_3758 <= in_reg[2977];
        i_10_3759 <= in_reg[3489];
        i_10_3760 <= in_reg[4001];
        i_10_3761 <= in_reg[4513];
        i_10_3762 <= in_reg[418];
        i_10_3763 <= in_reg[930];
        i_10_3764 <= in_reg[1442];
        i_10_3765 <= in_reg[1954];
        i_10_3766 <= in_reg[2466];
        i_10_3767 <= in_reg[2978];
        i_10_3768 <= in_reg[3490];
        i_10_3769 <= in_reg[4002];
        i_10_3770 <= in_reg[4514];
        i_10_3771 <= in_reg[419];
        i_10_3772 <= in_reg[931];
        i_10_3773 <= in_reg[1443];
        i_10_3774 <= in_reg[1955];
        i_10_3775 <= in_reg[2467];
        i_10_3776 <= in_reg[2979];
        i_10_3777 <= in_reg[3491];
        i_10_3778 <= in_reg[4003];
        i_10_3779 <= in_reg[4515];
        i_10_3780 <= in_reg[420];
        i_10_3781 <= in_reg[932];
        i_10_3782 <= in_reg[1444];
        i_10_3783 <= in_reg[1956];
        i_10_3784 <= in_reg[2468];
        i_10_3785 <= in_reg[2980];
        i_10_3786 <= in_reg[3492];
        i_10_3787 <= in_reg[4004];
        i_10_3788 <= in_reg[4516];
        i_10_3789 <= in_reg[421];
        i_10_3790 <= in_reg[933];
        i_10_3791 <= in_reg[1445];
        i_10_3792 <= in_reg[1957];
        i_10_3793 <= in_reg[2469];
        i_10_3794 <= in_reg[2981];
        i_10_3795 <= in_reg[3493];
        i_10_3796 <= in_reg[4005];
        i_10_3797 <= in_reg[4517];
        i_10_3798 <= in_reg[422];
        i_10_3799 <= in_reg[934];
        i_10_3800 <= in_reg[1446];
        i_10_3801 <= in_reg[1958];
        i_10_3802 <= in_reg[2470];
        i_10_3803 <= in_reg[2982];
        i_10_3804 <= in_reg[3494];
        i_10_3805 <= in_reg[4006];
        i_10_3806 <= in_reg[4518];
        i_10_3807 <= in_reg[423];
        i_10_3808 <= in_reg[935];
        i_10_3809 <= in_reg[1447];
        i_10_3810 <= in_reg[1959];
        i_10_3811 <= in_reg[2471];
        i_10_3812 <= in_reg[2983];
        i_10_3813 <= in_reg[3495];
        i_10_3814 <= in_reg[4007];
        i_10_3815 <= in_reg[4519];
        i_10_3816 <= in_reg[424];
        i_10_3817 <= in_reg[936];
        i_10_3818 <= in_reg[1448];
        i_10_3819 <= in_reg[1960];
        i_10_3820 <= in_reg[2472];
        i_10_3821 <= in_reg[2984];
        i_10_3822 <= in_reg[3496];
        i_10_3823 <= in_reg[4008];
        i_10_3824 <= in_reg[4520];
        i_10_3825 <= in_reg[425];
        i_10_3826 <= in_reg[937];
        i_10_3827 <= in_reg[1449];
        i_10_3828 <= in_reg[1961];
        i_10_3829 <= in_reg[2473];
        i_10_3830 <= in_reg[2985];
        i_10_3831 <= in_reg[3497];
        i_10_3832 <= in_reg[4009];
        i_10_3833 <= in_reg[4521];
        i_10_3834 <= in_reg[426];
        i_10_3835 <= in_reg[938];
        i_10_3836 <= in_reg[1450];
        i_10_3837 <= in_reg[1962];
        i_10_3838 <= in_reg[2474];
        i_10_3839 <= in_reg[2986];
        i_10_3840 <= in_reg[3498];
        i_10_3841 <= in_reg[4010];
        i_10_3842 <= in_reg[4522];
        i_10_3843 <= in_reg[427];
        i_10_3844 <= in_reg[939];
        i_10_3845 <= in_reg[1451];
        i_10_3846 <= in_reg[1963];
        i_10_3847 <= in_reg[2475];
        i_10_3848 <= in_reg[2987];
        i_10_3849 <= in_reg[3499];
        i_10_3850 <= in_reg[4011];
        i_10_3851 <= in_reg[4523];
        i_10_3852 <= in_reg[428];
        i_10_3853 <= in_reg[940];
        i_10_3854 <= in_reg[1452];
        i_10_3855 <= in_reg[1964];
        i_10_3856 <= in_reg[2476];
        i_10_3857 <= in_reg[2988];
        i_10_3858 <= in_reg[3500];
        i_10_3859 <= in_reg[4012];
        i_10_3860 <= in_reg[4524];
        i_10_3861 <= in_reg[429];
        i_10_3862 <= in_reg[941];
        i_10_3863 <= in_reg[1453];
        i_10_3864 <= in_reg[1965];
        i_10_3865 <= in_reg[2477];
        i_10_3866 <= in_reg[2989];
        i_10_3867 <= in_reg[3501];
        i_10_3868 <= in_reg[4013];
        i_10_3869 <= in_reg[4525];
        i_10_3870 <= in_reg[430];
        i_10_3871 <= in_reg[942];
        i_10_3872 <= in_reg[1454];
        i_10_3873 <= in_reg[1966];
        i_10_3874 <= in_reg[2478];
        i_10_3875 <= in_reg[2990];
        i_10_3876 <= in_reg[3502];
        i_10_3877 <= in_reg[4014];
        i_10_3878 <= in_reg[4526];
        i_10_3879 <= in_reg[431];
        i_10_3880 <= in_reg[943];
        i_10_3881 <= in_reg[1455];
        i_10_3882 <= in_reg[1967];
        i_10_3883 <= in_reg[2479];
        i_10_3884 <= in_reg[2991];
        i_10_3885 <= in_reg[3503];
        i_10_3886 <= in_reg[4015];
        i_10_3887 <= in_reg[4527];
        i_10_3888 <= in_reg[432];
        i_10_3889 <= in_reg[944];
        i_10_3890 <= in_reg[1456];
        i_10_3891 <= in_reg[1968];
        i_10_3892 <= in_reg[2480];
        i_10_3893 <= in_reg[2992];
        i_10_3894 <= in_reg[3504];
        i_10_3895 <= in_reg[4016];
        i_10_3896 <= in_reg[4528];
        i_10_3897 <= in_reg[433];
        i_10_3898 <= in_reg[945];
        i_10_3899 <= in_reg[1457];
        i_10_3900 <= in_reg[1969];
        i_10_3901 <= in_reg[2481];
        i_10_3902 <= in_reg[2993];
        i_10_3903 <= in_reg[3505];
        i_10_3904 <= in_reg[4017];
        i_10_3905 <= in_reg[4529];
        i_10_3906 <= in_reg[434];
        i_10_3907 <= in_reg[946];
        i_10_3908 <= in_reg[1458];
        i_10_3909 <= in_reg[1970];
        i_10_3910 <= in_reg[2482];
        i_10_3911 <= in_reg[2994];
        i_10_3912 <= in_reg[3506];
        i_10_3913 <= in_reg[4018];
        i_10_3914 <= in_reg[4530];
        i_10_3915 <= in_reg[435];
        i_10_3916 <= in_reg[947];
        i_10_3917 <= in_reg[1459];
        i_10_3918 <= in_reg[1971];
        i_10_3919 <= in_reg[2483];
        i_10_3920 <= in_reg[2995];
        i_10_3921 <= in_reg[3507];
        i_10_3922 <= in_reg[4019];
        i_10_3923 <= in_reg[4531];
        i_10_3924 <= in_reg[436];
        i_10_3925 <= in_reg[948];
        i_10_3926 <= in_reg[1460];
        i_10_3927 <= in_reg[1972];
        i_10_3928 <= in_reg[2484];
        i_10_3929 <= in_reg[2996];
        i_10_3930 <= in_reg[3508];
        i_10_3931 <= in_reg[4020];
        i_10_3932 <= in_reg[4532];
        i_10_3933 <= in_reg[437];
        i_10_3934 <= in_reg[949];
        i_10_3935 <= in_reg[1461];
        i_10_3936 <= in_reg[1973];
        i_10_3937 <= in_reg[2485];
        i_10_3938 <= in_reg[2997];
        i_10_3939 <= in_reg[3509];
        i_10_3940 <= in_reg[4021];
        i_10_3941 <= in_reg[4533];
        i_10_3942 <= in_reg[438];
        i_10_3943 <= in_reg[950];
        i_10_3944 <= in_reg[1462];
        i_10_3945 <= in_reg[1974];
        i_10_3946 <= in_reg[2486];
        i_10_3947 <= in_reg[2998];
        i_10_3948 <= in_reg[3510];
        i_10_3949 <= in_reg[4022];
        i_10_3950 <= in_reg[4534];
        i_10_3951 <= in_reg[439];
        i_10_3952 <= in_reg[951];
        i_10_3953 <= in_reg[1463];
        i_10_3954 <= in_reg[1975];
        i_10_3955 <= in_reg[2487];
        i_10_3956 <= in_reg[2999];
        i_10_3957 <= in_reg[3511];
        i_10_3958 <= in_reg[4023];
        i_10_3959 <= in_reg[4535];
        i_10_3960 <= in_reg[440];
        i_10_3961 <= in_reg[952];
        i_10_3962 <= in_reg[1464];
        i_10_3963 <= in_reg[1976];
        i_10_3964 <= in_reg[2488];
        i_10_3965 <= in_reg[3000];
        i_10_3966 <= in_reg[3512];
        i_10_3967 <= in_reg[4024];
        i_10_3968 <= in_reg[4536];
        i_10_3969 <= in_reg[441];
        i_10_3970 <= in_reg[953];
        i_10_3971 <= in_reg[1465];
        i_10_3972 <= in_reg[1977];
        i_10_3973 <= in_reg[2489];
        i_10_3974 <= in_reg[3001];
        i_10_3975 <= in_reg[3513];
        i_10_3976 <= in_reg[4025];
        i_10_3977 <= in_reg[4537];
        i_10_3978 <= in_reg[442];
        i_10_3979 <= in_reg[954];
        i_10_3980 <= in_reg[1466];
        i_10_3981 <= in_reg[1978];
        i_10_3982 <= in_reg[2490];
        i_10_3983 <= in_reg[3002];
        i_10_3984 <= in_reg[3514];
        i_10_3985 <= in_reg[4026];
        i_10_3986 <= in_reg[4538];
        i_10_3987 <= in_reg[443];
        i_10_3988 <= in_reg[955];
        i_10_3989 <= in_reg[1467];
        i_10_3990 <= in_reg[1979];
        i_10_3991 <= in_reg[2491];
        i_10_3992 <= in_reg[3003];
        i_10_3993 <= in_reg[3515];
        i_10_3994 <= in_reg[4027];
        i_10_3995 <= in_reg[4539];
        i_10_3996 <= in_reg[444];
        i_10_3997 <= in_reg[956];
        i_10_3998 <= in_reg[1468];
        i_10_3999 <= in_reg[1980];
        i_10_4000 <= in_reg[2492];
        i_10_4001 <= in_reg[3004];
        i_10_4002 <= in_reg[3516];
        i_10_4003 <= in_reg[4028];
        i_10_4004 <= in_reg[4540];
        i_10_4005 <= in_reg[445];
        i_10_4006 <= in_reg[957];
        i_10_4007 <= in_reg[1469];
        i_10_4008 <= in_reg[1981];
        i_10_4009 <= in_reg[2493];
        i_10_4010 <= in_reg[3005];
        i_10_4011 <= in_reg[3517];
        i_10_4012 <= in_reg[4029];
        i_10_4013 <= in_reg[4541];
        i_10_4014 <= in_reg[446];
        i_10_4015 <= in_reg[958];
        i_10_4016 <= in_reg[1470];
        i_10_4017 <= in_reg[1982];
        i_10_4018 <= in_reg[2494];
        i_10_4019 <= in_reg[3006];
        i_10_4020 <= in_reg[3518];
        i_10_4021 <= in_reg[4030];
        i_10_4022 <= in_reg[4542];
        i_10_4023 <= in_reg[447];
        i_10_4024 <= in_reg[959];
        i_10_4025 <= in_reg[1471];
        i_10_4026 <= in_reg[1983];
        i_10_4027 <= in_reg[2495];
        i_10_4028 <= in_reg[3007];
        i_10_4029 <= in_reg[3519];
        i_10_4030 <= in_reg[4031];
        i_10_4031 <= in_reg[4543];
        i_10_4032 <= in_reg[448];
        i_10_4033 <= in_reg[960];
        i_10_4034 <= in_reg[1472];
        i_10_4035 <= in_reg[1984];
        i_10_4036 <= in_reg[2496];
        i_10_4037 <= in_reg[3008];
        i_10_4038 <= in_reg[3520];
        i_10_4039 <= in_reg[4032];
        i_10_4040 <= in_reg[4544];
        i_10_4041 <= in_reg[449];
        i_10_4042 <= in_reg[961];
        i_10_4043 <= in_reg[1473];
        i_10_4044 <= in_reg[1985];
        i_10_4045 <= in_reg[2497];
        i_10_4046 <= in_reg[3009];
        i_10_4047 <= in_reg[3521];
        i_10_4048 <= in_reg[4033];
        i_10_4049 <= in_reg[4545];
        i_10_4050 <= in_reg[450];
        i_10_4051 <= in_reg[962];
        i_10_4052 <= in_reg[1474];
        i_10_4053 <= in_reg[1986];
        i_10_4054 <= in_reg[2498];
        i_10_4055 <= in_reg[3010];
        i_10_4056 <= in_reg[3522];
        i_10_4057 <= in_reg[4034];
        i_10_4058 <= in_reg[4546];
        i_10_4059 <= in_reg[451];
        i_10_4060 <= in_reg[963];
        i_10_4061 <= in_reg[1475];
        i_10_4062 <= in_reg[1987];
        i_10_4063 <= in_reg[2499];
        i_10_4064 <= in_reg[3011];
        i_10_4065 <= in_reg[3523];
        i_10_4066 <= in_reg[4035];
        i_10_4067 <= in_reg[4547];
        i_10_4068 <= in_reg[452];
        i_10_4069 <= in_reg[964];
        i_10_4070 <= in_reg[1476];
        i_10_4071 <= in_reg[1988];
        i_10_4072 <= in_reg[2500];
        i_10_4073 <= in_reg[3012];
        i_10_4074 <= in_reg[3524];
        i_10_4075 <= in_reg[4036];
        i_10_4076 <= in_reg[4548];
        i_10_4077 <= in_reg[453];
        i_10_4078 <= in_reg[965];
        i_10_4079 <= in_reg[1477];
        i_10_4080 <= in_reg[1989];
        i_10_4081 <= in_reg[2501];
        i_10_4082 <= in_reg[3013];
        i_10_4083 <= in_reg[3525];
        i_10_4084 <= in_reg[4037];
        i_10_4085 <= in_reg[4549];
        i_10_4086 <= in_reg[454];
        i_10_4087 <= in_reg[966];
        i_10_4088 <= in_reg[1478];
        i_10_4089 <= in_reg[1990];
        i_10_4090 <= in_reg[2502];
        i_10_4091 <= in_reg[3014];
        i_10_4092 <= in_reg[3526];
        i_10_4093 <= in_reg[4038];
        i_10_4094 <= in_reg[4550];
        i_10_4095 <= in_reg[455];
        i_10_4096 <= in_reg[967];
        i_10_4097 <= in_reg[1479];
        i_10_4098 <= in_reg[1991];
        i_10_4099 <= in_reg[2503];
        i_10_4100 <= in_reg[3015];
        i_10_4101 <= in_reg[3527];
        i_10_4102 <= in_reg[4039];
        i_10_4103 <= in_reg[4551];
        i_10_4104 <= in_reg[456];
        i_10_4105 <= in_reg[968];
        i_10_4106 <= in_reg[1480];
        i_10_4107 <= in_reg[1992];
        i_10_4108 <= in_reg[2504];
        i_10_4109 <= in_reg[3016];
        i_10_4110 <= in_reg[3528];
        i_10_4111 <= in_reg[4040];
        i_10_4112 <= in_reg[4552];
        i_10_4113 <= in_reg[457];
        i_10_4114 <= in_reg[969];
        i_10_4115 <= in_reg[1481];
        i_10_4116 <= in_reg[1993];
        i_10_4117 <= in_reg[2505];
        i_10_4118 <= in_reg[3017];
        i_10_4119 <= in_reg[3529];
        i_10_4120 <= in_reg[4041];
        i_10_4121 <= in_reg[4553];
        i_10_4122 <= in_reg[458];
        i_10_4123 <= in_reg[970];
        i_10_4124 <= in_reg[1482];
        i_10_4125 <= in_reg[1994];
        i_10_4126 <= in_reg[2506];
        i_10_4127 <= in_reg[3018];
        i_10_4128 <= in_reg[3530];
        i_10_4129 <= in_reg[4042];
        i_10_4130 <= in_reg[4554];
        i_10_4131 <= in_reg[459];
        i_10_4132 <= in_reg[971];
        i_10_4133 <= in_reg[1483];
        i_10_4134 <= in_reg[1995];
        i_10_4135 <= in_reg[2507];
        i_10_4136 <= in_reg[3019];
        i_10_4137 <= in_reg[3531];
        i_10_4138 <= in_reg[4043];
        i_10_4139 <= in_reg[4555];
        i_10_4140 <= in_reg[460];
        i_10_4141 <= in_reg[972];
        i_10_4142 <= in_reg[1484];
        i_10_4143 <= in_reg[1996];
        i_10_4144 <= in_reg[2508];
        i_10_4145 <= in_reg[3020];
        i_10_4146 <= in_reg[3532];
        i_10_4147 <= in_reg[4044];
        i_10_4148 <= in_reg[4556];
        i_10_4149 <= in_reg[461];
        i_10_4150 <= in_reg[973];
        i_10_4151 <= in_reg[1485];
        i_10_4152 <= in_reg[1997];
        i_10_4153 <= in_reg[2509];
        i_10_4154 <= in_reg[3021];
        i_10_4155 <= in_reg[3533];
        i_10_4156 <= in_reg[4045];
        i_10_4157 <= in_reg[4557];
        i_10_4158 <= in_reg[462];
        i_10_4159 <= in_reg[974];
        i_10_4160 <= in_reg[1486];
        i_10_4161 <= in_reg[1998];
        i_10_4162 <= in_reg[2510];
        i_10_4163 <= in_reg[3022];
        i_10_4164 <= in_reg[3534];
        i_10_4165 <= in_reg[4046];
        i_10_4166 <= in_reg[4558];
        i_10_4167 <= in_reg[463];
        i_10_4168 <= in_reg[975];
        i_10_4169 <= in_reg[1487];
        i_10_4170 <= in_reg[1999];
        i_10_4171 <= in_reg[2511];
        i_10_4172 <= in_reg[3023];
        i_10_4173 <= in_reg[3535];
        i_10_4174 <= in_reg[4047];
        i_10_4175 <= in_reg[4559];
        i_10_4176 <= in_reg[464];
        i_10_4177 <= in_reg[976];
        i_10_4178 <= in_reg[1488];
        i_10_4179 <= in_reg[2000];
        i_10_4180 <= in_reg[2512];
        i_10_4181 <= in_reg[3024];
        i_10_4182 <= in_reg[3536];
        i_10_4183 <= in_reg[4048];
        i_10_4184 <= in_reg[4560];
        i_10_4185 <= in_reg[465];
        i_10_4186 <= in_reg[977];
        i_10_4187 <= in_reg[1489];
        i_10_4188 <= in_reg[2001];
        i_10_4189 <= in_reg[2513];
        i_10_4190 <= in_reg[3025];
        i_10_4191 <= in_reg[3537];
        i_10_4192 <= in_reg[4049];
        i_10_4193 <= in_reg[4561];
        i_10_4194 <= in_reg[466];
        i_10_4195 <= in_reg[978];
        i_10_4196 <= in_reg[1490];
        i_10_4197 <= in_reg[2002];
        i_10_4198 <= in_reg[2514];
        i_10_4199 <= in_reg[3026];
        i_10_4200 <= in_reg[3538];
        i_10_4201 <= in_reg[4050];
        i_10_4202 <= in_reg[4562];
        i_10_4203 <= in_reg[467];
        i_10_4204 <= in_reg[979];
        i_10_4205 <= in_reg[1491];
        i_10_4206 <= in_reg[2003];
        i_10_4207 <= in_reg[2515];
        i_10_4208 <= in_reg[3027];
        i_10_4209 <= in_reg[3539];
        i_10_4210 <= in_reg[4051];
        i_10_4211 <= in_reg[4563];
        i_10_4212 <= in_reg[468];
        i_10_4213 <= in_reg[980];
        i_10_4214 <= in_reg[1492];
        i_10_4215 <= in_reg[2004];
        i_10_4216 <= in_reg[2516];
        i_10_4217 <= in_reg[3028];
        i_10_4218 <= in_reg[3540];
        i_10_4219 <= in_reg[4052];
        i_10_4220 <= in_reg[4564];
        i_10_4221 <= in_reg[469];
        i_10_4222 <= in_reg[981];
        i_10_4223 <= in_reg[1493];
        i_10_4224 <= in_reg[2005];
        i_10_4225 <= in_reg[2517];
        i_10_4226 <= in_reg[3029];
        i_10_4227 <= in_reg[3541];
        i_10_4228 <= in_reg[4053];
        i_10_4229 <= in_reg[4565];
        i_10_4230 <= in_reg[470];
        i_10_4231 <= in_reg[982];
        i_10_4232 <= in_reg[1494];
        i_10_4233 <= in_reg[2006];
        i_10_4234 <= in_reg[2518];
        i_10_4235 <= in_reg[3030];
        i_10_4236 <= in_reg[3542];
        i_10_4237 <= in_reg[4054];
        i_10_4238 <= in_reg[4566];
        i_10_4239 <= in_reg[471];
        i_10_4240 <= in_reg[983];
        i_10_4241 <= in_reg[1495];
        i_10_4242 <= in_reg[2007];
        i_10_4243 <= in_reg[2519];
        i_10_4244 <= in_reg[3031];
        i_10_4245 <= in_reg[3543];
        i_10_4246 <= in_reg[4055];
        i_10_4247 <= in_reg[4567];
        i_10_4248 <= in_reg[472];
        i_10_4249 <= in_reg[984];
        i_10_4250 <= in_reg[1496];
        i_10_4251 <= in_reg[2008];
        i_10_4252 <= in_reg[2520];
        i_10_4253 <= in_reg[3032];
        i_10_4254 <= in_reg[3544];
        i_10_4255 <= in_reg[4056];
        i_10_4256 <= in_reg[4568];
        i_10_4257 <= in_reg[473];
        i_10_4258 <= in_reg[985];
        i_10_4259 <= in_reg[1497];
        i_10_4260 <= in_reg[2009];
        i_10_4261 <= in_reg[2521];
        i_10_4262 <= in_reg[3033];
        i_10_4263 <= in_reg[3545];
        i_10_4264 <= in_reg[4057];
        i_10_4265 <= in_reg[4569];
        i_10_4266 <= in_reg[474];
        i_10_4267 <= in_reg[986];
        i_10_4268 <= in_reg[1498];
        i_10_4269 <= in_reg[2010];
        i_10_4270 <= in_reg[2522];
        i_10_4271 <= in_reg[3034];
        i_10_4272 <= in_reg[3546];
        i_10_4273 <= in_reg[4058];
        i_10_4274 <= in_reg[4570];
        i_10_4275 <= in_reg[475];
        i_10_4276 <= in_reg[987];
        i_10_4277 <= in_reg[1499];
        i_10_4278 <= in_reg[2011];
        i_10_4279 <= in_reg[2523];
        i_10_4280 <= in_reg[3035];
        i_10_4281 <= in_reg[3547];
        i_10_4282 <= in_reg[4059];
        i_10_4283 <= in_reg[4571];
        i_10_4284 <= in_reg[476];
        i_10_4285 <= in_reg[988];
        i_10_4286 <= in_reg[1500];
        i_10_4287 <= in_reg[2012];
        i_10_4288 <= in_reg[2524];
        i_10_4289 <= in_reg[3036];
        i_10_4290 <= in_reg[3548];
        i_10_4291 <= in_reg[4060];
        i_10_4292 <= in_reg[4572];
        i_10_4293 <= in_reg[477];
        i_10_4294 <= in_reg[989];
        i_10_4295 <= in_reg[1501];
        i_10_4296 <= in_reg[2013];
        i_10_4297 <= in_reg[2525];
        i_10_4298 <= in_reg[3037];
        i_10_4299 <= in_reg[3549];
        i_10_4300 <= in_reg[4061];
        i_10_4301 <= in_reg[4573];
        i_10_4302 <= in_reg[478];
        i_10_4303 <= in_reg[990];
        i_10_4304 <= in_reg[1502];
        i_10_4305 <= in_reg[2014];
        i_10_4306 <= in_reg[2526];
        i_10_4307 <= in_reg[3038];
        i_10_4308 <= in_reg[3550];
        i_10_4309 <= in_reg[4062];
        i_10_4310 <= in_reg[4574];
        i_10_4311 <= in_reg[479];
        i_10_4312 <= in_reg[991];
        i_10_4313 <= in_reg[1503];
        i_10_4314 <= in_reg[2015];
        i_10_4315 <= in_reg[2527];
        i_10_4316 <= in_reg[3039];
        i_10_4317 <= in_reg[3551];
        i_10_4318 <= in_reg[4063];
        i_10_4319 <= in_reg[4575];
        i_10_4320 <= in_reg[480];
        i_10_4321 <= in_reg[992];
        i_10_4322 <= in_reg[1504];
        i_10_4323 <= in_reg[2016];
        i_10_4324 <= in_reg[2528];
        i_10_4325 <= in_reg[3040];
        i_10_4326 <= in_reg[3552];
        i_10_4327 <= in_reg[4064];
        i_10_4328 <= in_reg[4576];
        i_10_4329 <= in_reg[481];
        i_10_4330 <= in_reg[993];
        i_10_4331 <= in_reg[1505];
        i_10_4332 <= in_reg[2017];
        i_10_4333 <= in_reg[2529];
        i_10_4334 <= in_reg[3041];
        i_10_4335 <= in_reg[3553];
        i_10_4336 <= in_reg[4065];
        i_10_4337 <= in_reg[4577];
        i_10_4338 <= in_reg[482];
        i_10_4339 <= in_reg[994];
        i_10_4340 <= in_reg[1506];
        i_10_4341 <= in_reg[2018];
        i_10_4342 <= in_reg[2530];
        i_10_4343 <= in_reg[3042];
        i_10_4344 <= in_reg[3554];
        i_10_4345 <= in_reg[4066];
        i_10_4346 <= in_reg[4578];
        i_10_4347 <= in_reg[483];
        i_10_4348 <= in_reg[995];
        i_10_4349 <= in_reg[1507];
        i_10_4350 <= in_reg[2019];
        i_10_4351 <= in_reg[2531];
        i_10_4352 <= in_reg[3043];
        i_10_4353 <= in_reg[3555];
        i_10_4354 <= in_reg[4067];
        i_10_4355 <= in_reg[4579];
        i_10_4356 <= in_reg[484];
        i_10_4357 <= in_reg[996];
        i_10_4358 <= in_reg[1508];
        i_10_4359 <= in_reg[2020];
        i_10_4360 <= in_reg[2532];
        i_10_4361 <= in_reg[3044];
        i_10_4362 <= in_reg[3556];
        i_10_4363 <= in_reg[4068];
        i_10_4364 <= in_reg[4580];
        i_10_4365 <= in_reg[485];
        i_10_4366 <= in_reg[997];
        i_10_4367 <= in_reg[1509];
        i_10_4368 <= in_reg[2021];
        i_10_4369 <= in_reg[2533];
        i_10_4370 <= in_reg[3045];
        i_10_4371 <= in_reg[3557];
        i_10_4372 <= in_reg[4069];
        i_10_4373 <= in_reg[4581];
        i_10_4374 <= in_reg[486];
        i_10_4375 <= in_reg[998];
        i_10_4376 <= in_reg[1510];
        i_10_4377 <= in_reg[2022];
        i_10_4378 <= in_reg[2534];
        i_10_4379 <= in_reg[3046];
        i_10_4380 <= in_reg[3558];
        i_10_4381 <= in_reg[4070];
        i_10_4382 <= in_reg[4582];
        i_10_4383 <= in_reg[487];
        i_10_4384 <= in_reg[999];
        i_10_4385 <= in_reg[1511];
        i_10_4386 <= in_reg[2023];
        i_10_4387 <= in_reg[2535];
        i_10_4388 <= in_reg[3047];
        i_10_4389 <= in_reg[3559];
        i_10_4390 <= in_reg[4071];
        i_10_4391 <= in_reg[4583];
        i_10_4392 <= in_reg[488];
        i_10_4393 <= in_reg[1000];
        i_10_4394 <= in_reg[1512];
        i_10_4395 <= in_reg[2024];
        i_10_4396 <= in_reg[2536];
        i_10_4397 <= in_reg[3048];
        i_10_4398 <= in_reg[3560];
        i_10_4399 <= in_reg[4072];
        i_10_4400 <= in_reg[4584];
        i_10_4401 <= in_reg[489];
        i_10_4402 <= in_reg[1001];
        i_10_4403 <= in_reg[1513];
        i_10_4404 <= in_reg[2025];
        i_10_4405 <= in_reg[2537];
        i_10_4406 <= in_reg[3049];
        i_10_4407 <= in_reg[3561];
        i_10_4408 <= in_reg[4073];
        i_10_4409 <= in_reg[4585];
        i_10_4410 <= in_reg[490];
        i_10_4411 <= in_reg[1002];
        i_10_4412 <= in_reg[1514];
        i_10_4413 <= in_reg[2026];
        i_10_4414 <= in_reg[2538];
        i_10_4415 <= in_reg[3050];
        i_10_4416 <= in_reg[3562];
        i_10_4417 <= in_reg[4074];
        i_10_4418 <= in_reg[4586];
        i_10_4419 <= in_reg[491];
        i_10_4420 <= in_reg[1003];
        i_10_4421 <= in_reg[1515];
        i_10_4422 <= in_reg[2027];
        i_10_4423 <= in_reg[2539];
        i_10_4424 <= in_reg[3051];
        i_10_4425 <= in_reg[3563];
        i_10_4426 <= in_reg[4075];
        i_10_4427 <= in_reg[4587];
        i_10_4428 <= in_reg[492];
        i_10_4429 <= in_reg[1004];
        i_10_4430 <= in_reg[1516];
        i_10_4431 <= in_reg[2028];
        i_10_4432 <= in_reg[2540];
        i_10_4433 <= in_reg[3052];
        i_10_4434 <= in_reg[3564];
        i_10_4435 <= in_reg[4076];
        i_10_4436 <= in_reg[4588];
        i_10_4437 <= in_reg[493];
        i_10_4438 <= in_reg[1005];
        i_10_4439 <= in_reg[1517];
        i_10_4440 <= in_reg[2029];
        i_10_4441 <= in_reg[2541];
        i_10_4442 <= in_reg[3053];
        i_10_4443 <= in_reg[3565];
        i_10_4444 <= in_reg[4077];
        i_10_4445 <= in_reg[4589];
        i_10_4446 <= in_reg[494];
        i_10_4447 <= in_reg[1006];
        i_10_4448 <= in_reg[1518];
        i_10_4449 <= in_reg[2030];
        i_10_4450 <= in_reg[2542];
        i_10_4451 <= in_reg[3054];
        i_10_4452 <= in_reg[3566];
        i_10_4453 <= in_reg[4078];
        i_10_4454 <= in_reg[4590];
        i_10_4455 <= in_reg[495];
        i_10_4456 <= in_reg[1007];
        i_10_4457 <= in_reg[1519];
        i_10_4458 <= in_reg[2031];
        i_10_4459 <= in_reg[2543];
        i_10_4460 <= in_reg[3055];
        i_10_4461 <= in_reg[3567];
        i_10_4462 <= in_reg[4079];
        i_10_4463 <= in_reg[4591];
        i_10_4464 <= in_reg[496];
        i_10_4465 <= in_reg[1008];
        i_10_4466 <= in_reg[1520];
        i_10_4467 <= in_reg[2032];
        i_10_4468 <= in_reg[2544];
        i_10_4469 <= in_reg[3056];
        i_10_4470 <= in_reg[3568];
        i_10_4471 <= in_reg[4080];
        i_10_4472 <= in_reg[4592];
        i_10_4473 <= in_reg[497];
        i_10_4474 <= in_reg[1009];
        i_10_4475 <= in_reg[1521];
        i_10_4476 <= in_reg[2033];
        i_10_4477 <= in_reg[2545];
        i_10_4478 <= in_reg[3057];
        i_10_4479 <= in_reg[3569];
        i_10_4480 <= in_reg[4081];
        i_10_4481 <= in_reg[4593];
        i_10_4482 <= in_reg[498];
        i_10_4483 <= in_reg[1010];
        i_10_4484 <= in_reg[1522];
        i_10_4485 <= in_reg[2034];
        i_10_4486 <= in_reg[2546];
        i_10_4487 <= in_reg[3058];
        i_10_4488 <= in_reg[3570];
        i_10_4489 <= in_reg[4082];
        i_10_4490 <= in_reg[4594];
        i_10_4491 <= in_reg[499];
        i_10_4492 <= in_reg[1011];
        i_10_4493 <= in_reg[1523];
        i_10_4494 <= in_reg[2035];
        i_10_4495 <= in_reg[2547];
        i_10_4496 <= in_reg[3059];
        i_10_4497 <= in_reg[3571];
        i_10_4498 <= in_reg[4083];
        i_10_4499 <= in_reg[4595];
        i_10_4500 <= in_reg[500];
        i_10_4501 <= in_reg[1012];
        i_10_4502 <= in_reg[1524];
        i_10_4503 <= in_reg[2036];
        i_10_4504 <= in_reg[2548];
        i_10_4505 <= in_reg[3060];
        i_10_4506 <= in_reg[3572];
        i_10_4507 <= in_reg[4084];
        i_10_4508 <= in_reg[4596];
        i_10_4509 <= in_reg[501];
        i_10_4510 <= in_reg[1013];
        i_10_4511 <= in_reg[1525];
        i_10_4512 <= in_reg[2037];
        i_10_4513 <= in_reg[2549];
        i_10_4514 <= in_reg[3061];
        i_10_4515 <= in_reg[3573];
        i_10_4516 <= in_reg[4085];
        i_10_4517 <= in_reg[4597];
        i_10_4518 <= in_reg[502];
        i_10_4519 <= in_reg[1014];
        i_10_4520 <= in_reg[1526];
        i_10_4521 <= in_reg[2038];
        i_10_4522 <= in_reg[2550];
        i_10_4523 <= in_reg[3062];
        i_10_4524 <= in_reg[3574];
        i_10_4525 <= in_reg[4086];
        i_10_4526 <= in_reg[4598];
        i_10_4527 <= in_reg[503];
        i_10_4528 <= in_reg[1015];
        i_10_4529 <= in_reg[1527];
        i_10_4530 <= in_reg[2039];
        i_10_4531 <= in_reg[2551];
        i_10_4532 <= in_reg[3063];
        i_10_4533 <= in_reg[3575];
        i_10_4534 <= in_reg[4087];
        i_10_4535 <= in_reg[4599];
        i_10_4536 <= in_reg[504];
        i_10_4537 <= in_reg[1016];
        i_10_4538 <= in_reg[1528];
        i_10_4539 <= in_reg[2040];
        i_10_4540 <= in_reg[2552];
        i_10_4541 <= in_reg[3064];
        i_10_4542 <= in_reg[3576];
        i_10_4543 <= in_reg[4088];
        i_10_4544 <= in_reg[4600];
        i_10_4545 <= in_reg[505];
        i_10_4546 <= in_reg[1017];
        i_10_4547 <= in_reg[1529];
        i_10_4548 <= in_reg[2041];
        i_10_4549 <= in_reg[2553];
        i_10_4550 <= in_reg[3065];
        i_10_4551 <= in_reg[3577];
        i_10_4552 <= in_reg[4089];
        i_10_4553 <= in_reg[4601];
        i_10_4554 <= in_reg[506];
        i_10_4555 <= in_reg[1018];
        i_10_4556 <= in_reg[1530];
        i_10_4557 <= in_reg[2042];
        i_10_4558 <= in_reg[2554];
        i_10_4559 <= in_reg[3066];
        i_10_4560 <= in_reg[3578];
        i_10_4561 <= in_reg[4090];
        i_10_4562 <= in_reg[4602];
        i_10_4563 <= in_reg[507];
        i_10_4564 <= in_reg[1019];
        i_10_4565 <= in_reg[1531];
        i_10_4566 <= in_reg[2043];
        i_10_4567 <= in_reg[2555];
        i_10_4568 <= in_reg[3067];
        i_10_4569 <= in_reg[3579];
        i_10_4570 <= in_reg[4091];
        i_10_4571 <= in_reg[4603];
        i_10_4572 <= in_reg[508];
        i_10_4573 <= in_reg[1020];
        i_10_4574 <= in_reg[1532];
        i_10_4575 <= in_reg[2044];
        i_10_4576 <= in_reg[2556];
        i_10_4577 <= in_reg[3068];
        i_10_4578 <= in_reg[3580];
        i_10_4579 <= in_reg[4092];
        i_10_4580 <= in_reg[4604];
        i_10_4581 <= in_reg[509];
        i_10_4582 <= in_reg[1021];
        i_10_4583 <= in_reg[1533];
        i_10_4584 <= in_reg[2045];
        i_10_4585 <= in_reg[2557];
        i_10_4586 <= in_reg[3069];
        i_10_4587 <= in_reg[3581];
        i_10_4588 <= in_reg[4093];
        i_10_4589 <= in_reg[4605];
        i_10_4590 <= in_reg[510];
        i_10_4591 <= in_reg[1022];
        i_10_4592 <= in_reg[1534];
        i_10_4593 <= in_reg[2046];
        i_10_4594 <= in_reg[2558];
        i_10_4595 <= in_reg[3070];
        i_10_4596 <= in_reg[3582];
        i_10_4597 <= in_reg[4094];
        i_10_4598 <= in_reg[4606];
        i_10_4599 <= in_reg[511];
        i_10_4600 <= in_reg[1023];
        i_10_4601 <= in_reg[1535];
        i_10_4602 <= in_reg[2047];
        i_10_4603 <= in_reg[2559];
        i_10_4604 <= in_reg[3071];
        i_10_4605 <= in_reg[3583];
        i_10_4606 <= in_reg[4095];
        i_10_4607 <= in_reg[4607];
        dly1 <= ap_start;
        dly2 <= dly1;
      end

  assign out_reg_ap_vld = dly2;
  assign ap_ready = dly2;
  assign ap_done = dly2;
  assign ap_idle = ~ap_start;

endmodule
