// Benchmark "kernel_13_0" written by ABC on Sun Jul 19 10:45:26 2020

module kernel_13_0 ( 
    i_13_0_20_0, i_13_0_59_0, i_13_0_74_0, i_13_0_76_0, i_13_0_182_0,
    i_13_0_187_0, i_13_0_232_0, i_13_0_283_0, i_13_0_286_0, i_13_0_338_0,
    i_13_0_445_0, i_13_0_448_0, i_13_0_535_0, i_13_0_548_0, i_13_0_574_0,
    i_13_0_617_0, i_13_0_629_0, i_13_0_643_0, i_13_0_644_0, i_13_0_646_0,
    i_13_0_647_0, i_13_0_652_0, i_13_0_689_0, i_13_0_718_0, i_13_0_781_0,
    i_13_0_782_0, i_13_0_827_0, i_13_0_835_0, i_13_0_895_0, i_13_0_977_0,
    i_13_0_980_0, i_13_0_1120_0, i_13_0_1124_0, i_13_0_1132_0,
    i_13_0_1142_0, i_13_0_1151_0, i_13_0_1231_0, i_13_0_1258_0,
    i_13_0_1277_0, i_13_0_1286_0, i_13_0_1394_0, i_13_0_1411_0,
    i_13_0_1435_0, i_13_0_1465_0, i_13_0_1483_0, i_13_0_1484_0,
    i_13_0_1627_0, i_13_0_1642_0, i_13_0_1646_0, i_13_0_1673_0,
    i_13_0_1753_0, i_13_0_1790_0, i_13_0_1796_0, i_13_0_1799_0,
    i_13_0_1802_0, i_13_0_1804_0, i_13_0_1840_0, i_13_0_1862_0,
    i_13_0_2000_0, i_13_0_2150_0, i_13_0_2168_0, i_13_0_2201_0,
    i_13_0_2239_0, i_13_0_2276_0, i_13_0_2311_0, i_13_0_2383_0,
    i_13_0_2545_0, i_13_0_2570_0, i_13_0_2848_0, i_13_0_2851_0,
    i_13_0_2852_0, i_13_0_2878_0, i_13_0_2879_0, i_13_0_2885_0,
    i_13_0_3028_0, i_13_0_3047_0, i_13_0_3095_0, i_13_0_3122_0,
    i_13_0_3293_0, i_13_0_3356_0, i_13_0_3389_0, i_13_0_3406_0,
    i_13_0_3433_0, i_13_0_3446_0, i_13_0_3482_0, i_13_0_3722_0,
    i_13_0_3734_0, i_13_0_3794_0, i_13_0_3839_0, i_13_0_3887_0,
    i_13_0_3985_0, i_13_0_4012_0, i_13_0_4013_0, i_13_0_4046_0,
    i_13_0_4189_0, i_13_0_4301_0, i_13_0_4315_0, i_13_0_4435_0,
    i_13_0_4481_0, i_13_0_4541_0,
    o_13_0_0_0  );
  input  i_13_0_20_0, i_13_0_59_0, i_13_0_74_0, i_13_0_76_0,
    i_13_0_182_0, i_13_0_187_0, i_13_0_232_0, i_13_0_283_0, i_13_0_286_0,
    i_13_0_338_0, i_13_0_445_0, i_13_0_448_0, i_13_0_535_0, i_13_0_548_0,
    i_13_0_574_0, i_13_0_617_0, i_13_0_629_0, i_13_0_643_0, i_13_0_644_0,
    i_13_0_646_0, i_13_0_647_0, i_13_0_652_0, i_13_0_689_0, i_13_0_718_0,
    i_13_0_781_0, i_13_0_782_0, i_13_0_827_0, i_13_0_835_0, i_13_0_895_0,
    i_13_0_977_0, i_13_0_980_0, i_13_0_1120_0, i_13_0_1124_0,
    i_13_0_1132_0, i_13_0_1142_0, i_13_0_1151_0, i_13_0_1231_0,
    i_13_0_1258_0, i_13_0_1277_0, i_13_0_1286_0, i_13_0_1394_0,
    i_13_0_1411_0, i_13_0_1435_0, i_13_0_1465_0, i_13_0_1483_0,
    i_13_0_1484_0, i_13_0_1627_0, i_13_0_1642_0, i_13_0_1646_0,
    i_13_0_1673_0, i_13_0_1753_0, i_13_0_1790_0, i_13_0_1796_0,
    i_13_0_1799_0, i_13_0_1802_0, i_13_0_1804_0, i_13_0_1840_0,
    i_13_0_1862_0, i_13_0_2000_0, i_13_0_2150_0, i_13_0_2168_0,
    i_13_0_2201_0, i_13_0_2239_0, i_13_0_2276_0, i_13_0_2311_0,
    i_13_0_2383_0, i_13_0_2545_0, i_13_0_2570_0, i_13_0_2848_0,
    i_13_0_2851_0, i_13_0_2852_0, i_13_0_2878_0, i_13_0_2879_0,
    i_13_0_2885_0, i_13_0_3028_0, i_13_0_3047_0, i_13_0_3095_0,
    i_13_0_3122_0, i_13_0_3293_0, i_13_0_3356_0, i_13_0_3389_0,
    i_13_0_3406_0, i_13_0_3433_0, i_13_0_3446_0, i_13_0_3482_0,
    i_13_0_3722_0, i_13_0_3734_0, i_13_0_3794_0, i_13_0_3839_0,
    i_13_0_3887_0, i_13_0_3985_0, i_13_0_4012_0, i_13_0_4013_0,
    i_13_0_4046_0, i_13_0_4189_0, i_13_0_4301_0, i_13_0_4315_0,
    i_13_0_4435_0, i_13_0_4481_0, i_13_0_4541_0;
  output o_13_0_0_0;
  assign o_13_0_0_0 = ~((~i_13_0_1627_0 & ((i_13_0_283_0 & ~i_13_0_535_0 & ~i_13_0_1483_0 & ~i_13_0_1484_0) | (~i_13_0_448_0 & ~i_13_0_4046_0))) | (~i_13_0_895_0 & ~i_13_0_1646_0 & ~i_13_0_2150_0) | (~i_13_0_1753_0 & ~i_13_0_2879_0 & ~i_13_0_4013_0) | (~i_13_0_1142_0 & i_13_0_4315_0));
endmodule



// Benchmark "kernel_13_1" written by ABC on Sun Jul 19 10:45:27 2020

module kernel_13_1 ( 
    i_13_1_40_0, i_13_1_73_0, i_13_1_90_0, i_13_1_91_0, i_13_1_93_0,
    i_13_1_94_0, i_13_1_97_0, i_13_1_111_0, i_13_1_118_0, i_13_1_160_0,
    i_13_1_177_0, i_13_1_273_0, i_13_1_306_0, i_13_1_310_0, i_13_1_364_0,
    i_13_1_411_0, i_13_1_561_0, i_13_1_567_0, i_13_1_568_0, i_13_1_571_0,
    i_13_1_604_0, i_13_1_694_0, i_13_1_697_0, i_13_1_729_0, i_13_1_730_0,
    i_13_1_733_0, i_13_1_793_0, i_13_1_855_0, i_13_1_861_0, i_13_1_863_0,
    i_13_1_942_0, i_13_1_1058_0, i_13_1_1210_0, i_13_1_1405_0,
    i_13_1_1440_0, i_13_1_1486_0, i_13_1_1491_0, i_13_1_1681_0,
    i_13_1_1781_0, i_13_1_1828_0, i_13_1_1836_0, i_13_1_1837_0,
    i_13_1_1862_0, i_13_1_1918_0, i_13_1_2172_0, i_13_1_2173_0,
    i_13_1_2205_0, i_13_1_2206_0, i_13_1_2316_0, i_13_1_2365_0,
    i_13_1_2421_0, i_13_1_2422_0, i_13_1_2433_0, i_13_1_2434_0,
    i_13_1_2437_0, i_13_1_2452_0, i_13_1_2464_0, i_13_1_2551_0,
    i_13_1_2677_0, i_13_1_2888_0, i_13_1_2985_0, i_13_1_3023_0,
    i_13_1_3064_0, i_13_1_3102_0, i_13_1_3149_0, i_13_1_3164_0,
    i_13_1_3166_0, i_13_1_3208_0, i_13_1_3423_0, i_13_1_3424_0,
    i_13_1_3489_0, i_13_1_3490_0, i_13_1_3535_0, i_13_1_3541_0,
    i_13_1_3568_0, i_13_1_3577_0, i_13_1_3682_0, i_13_1_3699_0,
    i_13_1_3762_0, i_13_1_3856_0, i_13_1_3870_0, i_13_1_3871_0,
    i_13_1_3872_0, i_13_1_3877_0, i_13_1_3972_0, i_13_1_3982_0,
    i_13_1_4118_0, i_13_1_4155_0, i_13_1_4278_0, i_13_1_4335_0,
    i_13_1_4350_0, i_13_1_4351_0, i_13_1_4354_0, i_13_1_4378_0,
    i_13_1_4390_0, i_13_1_4425_0, i_13_1_4536_0, i_13_1_4540_0,
    i_13_1_4567_0, i_13_1_4591_0,
    o_13_1_0_0  );
  input  i_13_1_40_0, i_13_1_73_0, i_13_1_90_0, i_13_1_91_0, i_13_1_93_0,
    i_13_1_94_0, i_13_1_97_0, i_13_1_111_0, i_13_1_118_0, i_13_1_160_0,
    i_13_1_177_0, i_13_1_273_0, i_13_1_306_0, i_13_1_310_0, i_13_1_364_0,
    i_13_1_411_0, i_13_1_561_0, i_13_1_567_0, i_13_1_568_0, i_13_1_571_0,
    i_13_1_604_0, i_13_1_694_0, i_13_1_697_0, i_13_1_729_0, i_13_1_730_0,
    i_13_1_733_0, i_13_1_793_0, i_13_1_855_0, i_13_1_861_0, i_13_1_863_0,
    i_13_1_942_0, i_13_1_1058_0, i_13_1_1210_0, i_13_1_1405_0,
    i_13_1_1440_0, i_13_1_1486_0, i_13_1_1491_0, i_13_1_1681_0,
    i_13_1_1781_0, i_13_1_1828_0, i_13_1_1836_0, i_13_1_1837_0,
    i_13_1_1862_0, i_13_1_1918_0, i_13_1_2172_0, i_13_1_2173_0,
    i_13_1_2205_0, i_13_1_2206_0, i_13_1_2316_0, i_13_1_2365_0,
    i_13_1_2421_0, i_13_1_2422_0, i_13_1_2433_0, i_13_1_2434_0,
    i_13_1_2437_0, i_13_1_2452_0, i_13_1_2464_0, i_13_1_2551_0,
    i_13_1_2677_0, i_13_1_2888_0, i_13_1_2985_0, i_13_1_3023_0,
    i_13_1_3064_0, i_13_1_3102_0, i_13_1_3149_0, i_13_1_3164_0,
    i_13_1_3166_0, i_13_1_3208_0, i_13_1_3423_0, i_13_1_3424_0,
    i_13_1_3489_0, i_13_1_3490_0, i_13_1_3535_0, i_13_1_3541_0,
    i_13_1_3568_0, i_13_1_3577_0, i_13_1_3682_0, i_13_1_3699_0,
    i_13_1_3762_0, i_13_1_3856_0, i_13_1_3870_0, i_13_1_3871_0,
    i_13_1_3872_0, i_13_1_3877_0, i_13_1_3972_0, i_13_1_3982_0,
    i_13_1_4118_0, i_13_1_4155_0, i_13_1_4278_0, i_13_1_4335_0,
    i_13_1_4350_0, i_13_1_4351_0, i_13_1_4354_0, i_13_1_4378_0,
    i_13_1_4390_0, i_13_1_4425_0, i_13_1_4536_0, i_13_1_4540_0,
    i_13_1_4567_0, i_13_1_4591_0;
  output o_13_1_0_0;
  assign o_13_1_0_0 = ~(i_13_1_1491_0 | (i_13_1_3568_0 & i_13_1_4378_0) | (~i_13_1_91_0 & ~i_13_1_3423_0) | (~i_13_1_90_0 & ~i_13_1_2173_0) | (~i_13_1_2206_0 & ~i_13_1_3164_0 & ~i_13_1_3762_0 & ~i_13_1_3871_0 & ~i_13_1_4350_0));
endmodule



// Benchmark "kernel_13_2" written by ABC on Sun Jul 19 10:45:27 2020

module kernel_13_2 ( 
    i_13_2_94_0, i_13_2_103_0, i_13_2_104_0, i_13_2_143_0, i_13_2_157_0,
    i_13_2_280_0, i_13_2_316_0, i_13_2_379_0, i_13_2_523_0, i_13_2_586_0,
    i_13_2_604_0, i_13_2_666_0, i_13_2_671_0, i_13_2_696_0, i_13_2_768_0,
    i_13_2_802_0, i_13_2_850_0, i_13_2_959_0, i_13_2_1081_0, i_13_2_1142_0,
    i_13_2_1206_0, i_13_2_1207_0, i_13_2_1274_0, i_13_2_1277_0,
    i_13_2_1300_0, i_13_2_1341_0, i_13_2_1342_0, i_13_2_1343_0,
    i_13_2_1363_0, i_13_2_1403_0, i_13_2_1435_0, i_13_2_1440_0,
    i_13_2_1467_0, i_13_2_1515_0, i_13_2_1594_0, i_13_2_1692_0,
    i_13_2_1714_0, i_13_2_1750_0, i_13_2_1781_0, i_13_2_1802_0,
    i_13_2_1810_0, i_13_2_1840_0, i_13_2_1882_0, i_13_2_1900_0,
    i_13_2_1926_0, i_13_2_1927_0, i_13_2_1939_0, i_13_2_2002_0,
    i_13_2_2011_0, i_13_2_2052_0, i_13_2_2053_0, i_13_2_2054_0,
    i_13_2_2173_0, i_13_2_2189_0, i_13_2_2197_0, i_13_2_2236_0,
    i_13_2_2278_0, i_13_2_2396_0, i_13_2_2423_0, i_13_2_2450_0,
    i_13_2_2548_0, i_13_2_2592_0, i_13_2_2614_0, i_13_2_2615_0,
    i_13_2_2695_0, i_13_2_2710_0, i_13_2_2853_0, i_13_2_2854_0,
    i_13_2_3019_0, i_13_2_3109_0, i_13_2_3329_0, i_13_2_3343_0,
    i_13_2_3366_0, i_13_2_3367_0, i_13_2_3386_0, i_13_2_3398_0,
    i_13_2_3404_0, i_13_2_3439_0, i_13_2_3487_0, i_13_2_3502_0,
    i_13_2_3611_0, i_13_2_3619_0, i_13_2_3650_0, i_13_2_3736_0,
    i_13_2_3910_0, i_13_2_3931_0, i_13_2_3994_0, i_13_2_3995_0,
    i_13_2_4015_0, i_13_2_4087_0, i_13_2_4104_0, i_13_2_4230_0,
    i_13_2_4231_0, i_13_2_4232_0, i_13_2_4267_0, i_13_2_4392_0,
    i_13_2_4393_0, i_13_2_4394_0, i_13_2_4554_0, i_13_2_4559_0,
    o_13_2_0_0  );
  input  i_13_2_94_0, i_13_2_103_0, i_13_2_104_0, i_13_2_143_0,
    i_13_2_157_0, i_13_2_280_0, i_13_2_316_0, i_13_2_379_0, i_13_2_523_0,
    i_13_2_586_0, i_13_2_604_0, i_13_2_666_0, i_13_2_671_0, i_13_2_696_0,
    i_13_2_768_0, i_13_2_802_0, i_13_2_850_0, i_13_2_959_0, i_13_2_1081_0,
    i_13_2_1142_0, i_13_2_1206_0, i_13_2_1207_0, i_13_2_1274_0,
    i_13_2_1277_0, i_13_2_1300_0, i_13_2_1341_0, i_13_2_1342_0,
    i_13_2_1343_0, i_13_2_1363_0, i_13_2_1403_0, i_13_2_1435_0,
    i_13_2_1440_0, i_13_2_1467_0, i_13_2_1515_0, i_13_2_1594_0,
    i_13_2_1692_0, i_13_2_1714_0, i_13_2_1750_0, i_13_2_1781_0,
    i_13_2_1802_0, i_13_2_1810_0, i_13_2_1840_0, i_13_2_1882_0,
    i_13_2_1900_0, i_13_2_1926_0, i_13_2_1927_0, i_13_2_1939_0,
    i_13_2_2002_0, i_13_2_2011_0, i_13_2_2052_0, i_13_2_2053_0,
    i_13_2_2054_0, i_13_2_2173_0, i_13_2_2189_0, i_13_2_2197_0,
    i_13_2_2236_0, i_13_2_2278_0, i_13_2_2396_0, i_13_2_2423_0,
    i_13_2_2450_0, i_13_2_2548_0, i_13_2_2592_0, i_13_2_2614_0,
    i_13_2_2615_0, i_13_2_2695_0, i_13_2_2710_0, i_13_2_2853_0,
    i_13_2_2854_0, i_13_2_3019_0, i_13_2_3109_0, i_13_2_3329_0,
    i_13_2_3343_0, i_13_2_3366_0, i_13_2_3367_0, i_13_2_3386_0,
    i_13_2_3398_0, i_13_2_3404_0, i_13_2_3439_0, i_13_2_3487_0,
    i_13_2_3502_0, i_13_2_3611_0, i_13_2_3619_0, i_13_2_3650_0,
    i_13_2_3736_0, i_13_2_3910_0, i_13_2_3931_0, i_13_2_3994_0,
    i_13_2_3995_0, i_13_2_4015_0, i_13_2_4087_0, i_13_2_4104_0,
    i_13_2_4230_0, i_13_2_4231_0, i_13_2_4232_0, i_13_2_4267_0,
    i_13_2_4392_0, i_13_2_4393_0, i_13_2_4394_0, i_13_2_4554_0,
    i_13_2_4559_0;
  output o_13_2_0_0;
  assign o_13_2_0_0 = ~(~i_13_2_586_0 | (~i_13_2_4267_0 & ~i_13_2_4393_0) | (~i_13_2_1342_0 & ~i_13_2_3109_0));
endmodule



// Benchmark "kernel_13_3" written by ABC on Sun Jul 19 10:45:28 2020

module kernel_13_3 ( 
    i_13_3_46_0, i_13_3_74_0, i_13_3_100_0, i_13_3_108_0, i_13_3_110_0,
    i_13_3_127_0, i_13_3_166_0, i_13_3_280_0, i_13_3_281_0, i_13_3_284_0,
    i_13_3_486_0, i_13_3_677_0, i_13_3_723_0, i_13_3_758_0, i_13_3_760_0,
    i_13_3_794_0, i_13_3_820_0, i_13_3_821_0, i_13_3_856_0, i_13_3_946_0,
    i_13_3_1215_0, i_13_3_1216_0, i_13_3_1217_0, i_13_3_1219_0,
    i_13_3_1317_0, i_13_3_1341_0, i_13_3_1388_0, i_13_3_1422_0,
    i_13_3_1424_0, i_13_3_1486_0, i_13_3_1487_0, i_13_3_1494_0,
    i_13_3_1566_0, i_13_3_1605_0, i_13_3_1630_0, i_13_3_1732_0,
    i_13_3_1774_0, i_13_3_1804_0, i_13_3_1837_0, i_13_3_1838_0,
    i_13_3_1841_0, i_13_3_1883_0, i_13_3_1911_0, i_13_3_1940_0,
    i_13_3_1945_0, i_13_3_1999_0, i_13_3_2000_0, i_13_3_2055_0,
    i_13_3_2146_0, i_13_3_2170_0, i_13_3_2236_0, i_13_3_2263_0,
    i_13_3_2335_0, i_13_3_2422_0, i_13_3_2435_0, i_13_3_2448_0,
    i_13_3_2532_0, i_13_3_2611_0, i_13_3_2612_0, i_13_3_2614_0,
    i_13_3_2709_0, i_13_3_2716_0, i_13_3_2746_0, i_13_3_2767_0,
    i_13_3_2782_0, i_13_3_2882_0, i_13_3_2955_0, i_13_3_2961_0,
    i_13_3_3034_0, i_13_3_3051_0, i_13_3_3145_0, i_13_3_3146_0,
    i_13_3_3379_0, i_13_3_3422_0, i_13_3_3438_0, i_13_3_3452_0,
    i_13_3_3502_0, i_13_3_3503_0, i_13_3_3529_0, i_13_3_3530_0,
    i_13_3_3610_0, i_13_3_3726_0, i_13_3_3729_0, i_13_3_3735_0,
    i_13_3_3736_0, i_13_3_3739_0, i_13_3_3872_0, i_13_3_3889_0,
    i_13_3_3890_0, i_13_3_3980_0, i_13_3_4053_0, i_13_3_4121_0,
    i_13_3_4158_0, i_13_3_4248_0, i_13_3_4252_0, i_13_3_4262_0,
    i_13_3_4322_0, i_13_3_4340_0, i_13_3_4415_0, i_13_3_4557_0,
    o_13_3_0_0  );
  input  i_13_3_46_0, i_13_3_74_0, i_13_3_100_0, i_13_3_108_0,
    i_13_3_110_0, i_13_3_127_0, i_13_3_166_0, i_13_3_280_0, i_13_3_281_0,
    i_13_3_284_0, i_13_3_486_0, i_13_3_677_0, i_13_3_723_0, i_13_3_758_0,
    i_13_3_760_0, i_13_3_794_0, i_13_3_820_0, i_13_3_821_0, i_13_3_856_0,
    i_13_3_946_0, i_13_3_1215_0, i_13_3_1216_0, i_13_3_1217_0,
    i_13_3_1219_0, i_13_3_1317_0, i_13_3_1341_0, i_13_3_1388_0,
    i_13_3_1422_0, i_13_3_1424_0, i_13_3_1486_0, i_13_3_1487_0,
    i_13_3_1494_0, i_13_3_1566_0, i_13_3_1605_0, i_13_3_1630_0,
    i_13_3_1732_0, i_13_3_1774_0, i_13_3_1804_0, i_13_3_1837_0,
    i_13_3_1838_0, i_13_3_1841_0, i_13_3_1883_0, i_13_3_1911_0,
    i_13_3_1940_0, i_13_3_1945_0, i_13_3_1999_0, i_13_3_2000_0,
    i_13_3_2055_0, i_13_3_2146_0, i_13_3_2170_0, i_13_3_2236_0,
    i_13_3_2263_0, i_13_3_2335_0, i_13_3_2422_0, i_13_3_2435_0,
    i_13_3_2448_0, i_13_3_2532_0, i_13_3_2611_0, i_13_3_2612_0,
    i_13_3_2614_0, i_13_3_2709_0, i_13_3_2716_0, i_13_3_2746_0,
    i_13_3_2767_0, i_13_3_2782_0, i_13_3_2882_0, i_13_3_2955_0,
    i_13_3_2961_0, i_13_3_3034_0, i_13_3_3051_0, i_13_3_3145_0,
    i_13_3_3146_0, i_13_3_3379_0, i_13_3_3422_0, i_13_3_3438_0,
    i_13_3_3452_0, i_13_3_3502_0, i_13_3_3503_0, i_13_3_3529_0,
    i_13_3_3530_0, i_13_3_3610_0, i_13_3_3726_0, i_13_3_3729_0,
    i_13_3_3735_0, i_13_3_3736_0, i_13_3_3739_0, i_13_3_3872_0,
    i_13_3_3889_0, i_13_3_3890_0, i_13_3_3980_0, i_13_3_4053_0,
    i_13_3_4121_0, i_13_3_4158_0, i_13_3_4248_0, i_13_3_4252_0,
    i_13_3_4262_0, i_13_3_4322_0, i_13_3_4340_0, i_13_3_4415_0,
    i_13_3_4557_0;
  output o_13_3_0_0;
  assign o_13_3_0_0 = ~((i_13_3_2236_0 & (~i_13_3_2170_0 | (~i_13_3_3739_0 & ~i_13_3_4252_0))) | (~i_13_3_3890_0 & ((~i_13_3_280_0 & ~i_13_3_1217_0 & ~i_13_3_1837_0) | (~i_13_3_1216_0 & i_13_3_2146_0 & ~i_13_3_3530_0))) | (~i_13_3_821_0 & ~i_13_3_1219_0 & ~i_13_3_1732_0) | (~i_13_3_1774_0 & ~i_13_3_3503_0 & ~i_13_3_4415_0));
endmodule



// Benchmark "kernel_13_4" written by ABC on Sun Jul 19 10:45:29 2020

module kernel_13_4 ( 
    i_13_4_192_0, i_13_4_199_0, i_13_4_225_0, i_13_4_324_0, i_13_4_378_0,
    i_13_4_531_0, i_13_4_532_0, i_13_4_573_0, i_13_4_577_0, i_13_4_639_0,
    i_13_4_640_0, i_13_4_658_0, i_13_4_660_0, i_13_4_661_0, i_13_4_714_0,
    i_13_4_768_0, i_13_4_849_0, i_13_4_927_0, i_13_4_945_0, i_13_4_1062_0,
    i_13_4_1080_0, i_13_4_1084_0, i_13_4_1116_0, i_13_4_1188_0,
    i_13_4_1206_0, i_13_4_1254_0, i_13_4_1407_0, i_13_4_1423_0,
    i_13_4_1506_0, i_13_4_1513_0, i_13_4_1539_0, i_13_4_1593_0,
    i_13_4_1594_0, i_13_4_1638_0, i_13_4_1639_0, i_13_4_1710_0,
    i_13_4_1719_0, i_13_4_1782_0, i_13_4_1783_0, i_13_4_1792_0,
    i_13_4_1800_0, i_13_4_1801_0, i_13_4_1881_0, i_13_4_1882_0,
    i_13_4_1929_0, i_13_4_1989_0, i_13_4_1990_0, i_13_4_2055_0,
    i_13_4_2092_0, i_13_4_2100_0, i_13_4_2116_0, i_13_4_2341_0,
    i_13_4_2358_0, i_13_4_2376_0, i_13_4_2424_0, i_13_4_2460_0,
    i_13_4_2524_0, i_13_4_2532_0, i_13_4_2569_0, i_13_4_2673_0,
    i_13_4_2817_0, i_13_4_2844_0, i_13_4_2845_0, i_13_4_2934_0,
    i_13_4_2935_0, i_13_4_3024_0, i_13_4_3114_0, i_13_4_3141_0,
    i_13_4_3258_0, i_13_4_3259_0, i_13_4_3267_0, i_13_4_3285_0,
    i_13_4_3286_0, i_13_4_3381_0, i_13_4_3384_0, i_13_4_3394_0,
    i_13_4_3415_0, i_13_4_3420_0, i_13_4_3421_0, i_13_4_3423_0,
    i_13_4_3424_0, i_13_4_3447_0, i_13_4_3451_0, i_13_4_3472_0,
    i_13_4_3753_0, i_13_4_3790_0, i_13_4_3873_0, i_13_4_3919_0,
    i_13_4_3924_0, i_13_4_3982_0, i_13_4_4008_0, i_13_4_4009_0,
    i_13_4_4018_0, i_13_4_4050_0, i_13_4_4077_0, i_13_4_4078_0,
    i_13_4_4207_0, i_13_4_4249_0, i_13_4_4420_0, i_13_4_4521_0,
    o_13_4_0_0  );
  input  i_13_4_192_0, i_13_4_199_0, i_13_4_225_0, i_13_4_324_0,
    i_13_4_378_0, i_13_4_531_0, i_13_4_532_0, i_13_4_573_0, i_13_4_577_0,
    i_13_4_639_0, i_13_4_640_0, i_13_4_658_0, i_13_4_660_0, i_13_4_661_0,
    i_13_4_714_0, i_13_4_768_0, i_13_4_849_0, i_13_4_927_0, i_13_4_945_0,
    i_13_4_1062_0, i_13_4_1080_0, i_13_4_1084_0, i_13_4_1116_0,
    i_13_4_1188_0, i_13_4_1206_0, i_13_4_1254_0, i_13_4_1407_0,
    i_13_4_1423_0, i_13_4_1506_0, i_13_4_1513_0, i_13_4_1539_0,
    i_13_4_1593_0, i_13_4_1594_0, i_13_4_1638_0, i_13_4_1639_0,
    i_13_4_1710_0, i_13_4_1719_0, i_13_4_1782_0, i_13_4_1783_0,
    i_13_4_1792_0, i_13_4_1800_0, i_13_4_1801_0, i_13_4_1881_0,
    i_13_4_1882_0, i_13_4_1929_0, i_13_4_1989_0, i_13_4_1990_0,
    i_13_4_2055_0, i_13_4_2092_0, i_13_4_2100_0, i_13_4_2116_0,
    i_13_4_2341_0, i_13_4_2358_0, i_13_4_2376_0, i_13_4_2424_0,
    i_13_4_2460_0, i_13_4_2524_0, i_13_4_2532_0, i_13_4_2569_0,
    i_13_4_2673_0, i_13_4_2817_0, i_13_4_2844_0, i_13_4_2845_0,
    i_13_4_2934_0, i_13_4_2935_0, i_13_4_3024_0, i_13_4_3114_0,
    i_13_4_3141_0, i_13_4_3258_0, i_13_4_3259_0, i_13_4_3267_0,
    i_13_4_3285_0, i_13_4_3286_0, i_13_4_3381_0, i_13_4_3384_0,
    i_13_4_3394_0, i_13_4_3415_0, i_13_4_3420_0, i_13_4_3421_0,
    i_13_4_3423_0, i_13_4_3424_0, i_13_4_3447_0, i_13_4_3451_0,
    i_13_4_3472_0, i_13_4_3753_0, i_13_4_3790_0, i_13_4_3873_0,
    i_13_4_3919_0, i_13_4_3924_0, i_13_4_3982_0, i_13_4_4008_0,
    i_13_4_4009_0, i_13_4_4018_0, i_13_4_4050_0, i_13_4_4077_0,
    i_13_4_4078_0, i_13_4_4207_0, i_13_4_4249_0, i_13_4_4420_0,
    i_13_4_4521_0;
  output o_13_4_0_0;
  assign o_13_4_0_0 = ~(~i_13_4_3286_0 | (~i_13_4_531_0 & ~i_13_4_3420_0) | (~i_13_4_2055_0 & ~i_13_4_3285_0));
endmodule



// Benchmark "kernel_13_5" written by ABC on Sun Jul 19 10:45:30 2020

module kernel_13_5 ( 
    i_13_5_71_0, i_13_5_76_0, i_13_5_175_0, i_13_5_178_0, i_13_5_209_0,
    i_13_5_245_0, i_13_5_283_0, i_13_5_284_0, i_13_5_286_0, i_13_5_287_0,
    i_13_5_374_0, i_13_5_410_0, i_13_5_517_0, i_13_5_526_0, i_13_5_527_0,
    i_13_5_625_0, i_13_5_689_0, i_13_5_691_0, i_13_5_800_0, i_13_5_814_0,
    i_13_5_818_0, i_13_5_826_0, i_13_5_851_0, i_13_5_923_0, i_13_5_1073_0,
    i_13_5_1097_0, i_13_5_1147_0, i_13_5_1312_0, i_13_5_1313_0,
    i_13_5_1499_0, i_13_5_1502_0, i_13_5_1543_0, i_13_5_1633_0,
    i_13_5_1634_0, i_13_5_1636_0, i_13_5_1637_0, i_13_5_1678_0,
    i_13_5_1681_0, i_13_5_1696_0, i_13_5_2005_0, i_13_5_2146_0,
    i_13_5_2194_0, i_13_5_2195_0, i_13_5_2291_0, i_13_5_2426_0,
    i_13_5_2438_0, i_13_5_2453_0, i_13_5_2462_0, i_13_5_2465_0,
    i_13_5_2527_0, i_13_5_2543_0, i_13_5_2677_0, i_13_5_2906_0,
    i_13_5_3025_0, i_13_5_3029_0, i_13_5_3050_0, i_13_5_3145_0,
    i_13_5_3146_0, i_13_5_3148_0, i_13_5_3172_0, i_13_5_3175_0,
    i_13_5_3272_0, i_13_5_3274_0, i_13_5_3275_0, i_13_5_3418_0,
    i_13_5_3425_0, i_13_5_3427_0, i_13_5_3428_0, i_13_5_3485_0,
    i_13_5_3490_0, i_13_5_3548_0, i_13_5_3616_0, i_13_5_3730_0,
    i_13_5_3731_0, i_13_5_3733_0, i_13_5_3734_0, i_13_5_3866_0,
    i_13_5_3892_0, i_13_5_3911_0, i_13_5_3913_0, i_13_5_3937_0,
    i_13_5_3995_0, i_13_5_4018_0, i_13_5_4019_0, i_13_5_4021_0,
    i_13_5_4022_0, i_13_5_4252_0, i_13_5_4253_0, i_13_5_4255_0,
    i_13_5_4256_0, i_13_5_4262_0, i_13_5_4264_0, i_13_5_4265_0,
    i_13_5_4342_0, i_13_5_4511_0, i_13_5_4559_0, i_13_5_4561_0,
    i_13_5_4562_0, i_13_5_4565_0, i_13_5_4586_0,
    o_13_5_0_0  );
  input  i_13_5_71_0, i_13_5_76_0, i_13_5_175_0, i_13_5_178_0,
    i_13_5_209_0, i_13_5_245_0, i_13_5_283_0, i_13_5_284_0, i_13_5_286_0,
    i_13_5_287_0, i_13_5_374_0, i_13_5_410_0, i_13_5_517_0, i_13_5_526_0,
    i_13_5_527_0, i_13_5_625_0, i_13_5_689_0, i_13_5_691_0, i_13_5_800_0,
    i_13_5_814_0, i_13_5_818_0, i_13_5_826_0, i_13_5_851_0, i_13_5_923_0,
    i_13_5_1073_0, i_13_5_1097_0, i_13_5_1147_0, i_13_5_1312_0,
    i_13_5_1313_0, i_13_5_1499_0, i_13_5_1502_0, i_13_5_1543_0,
    i_13_5_1633_0, i_13_5_1634_0, i_13_5_1636_0, i_13_5_1637_0,
    i_13_5_1678_0, i_13_5_1681_0, i_13_5_1696_0, i_13_5_2005_0,
    i_13_5_2146_0, i_13_5_2194_0, i_13_5_2195_0, i_13_5_2291_0,
    i_13_5_2426_0, i_13_5_2438_0, i_13_5_2453_0, i_13_5_2462_0,
    i_13_5_2465_0, i_13_5_2527_0, i_13_5_2543_0, i_13_5_2677_0,
    i_13_5_2906_0, i_13_5_3025_0, i_13_5_3029_0, i_13_5_3050_0,
    i_13_5_3145_0, i_13_5_3146_0, i_13_5_3148_0, i_13_5_3172_0,
    i_13_5_3175_0, i_13_5_3272_0, i_13_5_3274_0, i_13_5_3275_0,
    i_13_5_3418_0, i_13_5_3425_0, i_13_5_3427_0, i_13_5_3428_0,
    i_13_5_3485_0, i_13_5_3490_0, i_13_5_3548_0, i_13_5_3616_0,
    i_13_5_3730_0, i_13_5_3731_0, i_13_5_3733_0, i_13_5_3734_0,
    i_13_5_3866_0, i_13_5_3892_0, i_13_5_3911_0, i_13_5_3913_0,
    i_13_5_3937_0, i_13_5_3995_0, i_13_5_4018_0, i_13_5_4019_0,
    i_13_5_4021_0, i_13_5_4022_0, i_13_5_4252_0, i_13_5_4253_0,
    i_13_5_4255_0, i_13_5_4256_0, i_13_5_4262_0, i_13_5_4264_0,
    i_13_5_4265_0, i_13_5_4342_0, i_13_5_4511_0, i_13_5_4559_0,
    i_13_5_4561_0, i_13_5_4562_0, i_13_5_4565_0, i_13_5_4586_0;
  output o_13_5_0_0;
  assign o_13_5_0_0 = ~((~i_13_5_3734_0 & ((~i_13_5_2465_0 & ~i_13_5_3427_0) | (i_13_5_1681_0 & ~i_13_5_4262_0 & ~i_13_5_4561_0))) | (~i_13_5_287_0 & ~i_13_5_4559_0) | (~i_13_5_818_0 & ~i_13_5_3866_0 & ~i_13_5_3892_0 & ~i_13_5_3995_0 & ~i_13_5_4562_0));
endmodule



// Benchmark "kernel_13_6" written by ABC on Sun Jul 19 10:45:31 2020

module kernel_13_6 ( 
    i_13_6_139_0, i_13_6_229_0, i_13_6_280_0, i_13_6_282_0, i_13_6_285_0,
    i_13_6_410_0, i_13_6_418_0, i_13_6_475_0, i_13_6_561_0, i_13_6_562_0,
    i_13_6_574_0, i_13_6_849_0, i_13_6_850_0, i_13_6_853_0, i_13_6_924_0,
    i_13_6_981_0, i_13_6_988_0, i_13_6_1018_0, i_13_6_1021_0,
    i_13_6_1075_0, i_13_6_1219_0, i_13_6_1262_0, i_13_6_1308_0,
    i_13_6_1342_0, i_13_6_1345_0, i_13_6_1488_0, i_13_6_1496_0,
    i_13_6_1498_0, i_13_6_1515_0, i_13_6_1520_0, i_13_6_1630_0,
    i_13_6_1669_0, i_13_6_1678_0, i_13_6_1730_0, i_13_6_1753_0,
    i_13_6_1773_0, i_13_6_1809_0, i_13_6_1829_0, i_13_6_1854_0,
    i_13_6_1857_0, i_13_6_1858_0, i_13_6_1861_0, i_13_6_2002_0,
    i_13_6_2008_0, i_13_6_2028_0, i_13_6_2191_0, i_13_6_2226_0,
    i_13_6_2452_0, i_13_6_2455_0, i_13_6_2461_0, i_13_6_2539_0,
    i_13_6_2542_0, i_13_6_2544_0, i_13_6_2590_0, i_13_6_2722_0,
    i_13_6_2767_0, i_13_6_2857_0, i_13_6_3007_0, i_13_6_3010_0,
    i_13_6_3012_0, i_13_6_3037_0, i_13_6_3061_0, i_13_6_3064_0,
    i_13_6_3111_0, i_13_6_3127_0, i_13_6_3211_0, i_13_6_3235_0,
    i_13_6_3271_0, i_13_6_3442_0, i_13_6_3487_0, i_13_6_3490_0,
    i_13_6_3508_0, i_13_6_3541_0, i_13_6_3577_0, i_13_6_3640_0,
    i_13_6_3645_0, i_13_6_3729_0, i_13_6_3787_0, i_13_6_3817_0,
    i_13_6_3820_0, i_13_6_3838_0, i_13_6_3856_0, i_13_6_3888_0,
    i_13_6_3889_0, i_13_6_3907_0, i_13_6_3909_0, i_13_6_3910_0,
    i_13_6_3912_0, i_13_6_4078_0, i_13_6_4086_0, i_13_6_4250_0,
    i_13_6_4252_0, i_13_6_4254_0, i_13_6_4255_0, i_13_6_4375_0,
    i_13_6_4378_0, i_13_6_4380_0, i_13_6_4420_0, i_13_6_4426_0,
    i_13_6_4531_0,
    o_13_6_0_0  );
  input  i_13_6_139_0, i_13_6_229_0, i_13_6_280_0, i_13_6_282_0,
    i_13_6_285_0, i_13_6_410_0, i_13_6_418_0, i_13_6_475_0, i_13_6_561_0,
    i_13_6_562_0, i_13_6_574_0, i_13_6_849_0, i_13_6_850_0, i_13_6_853_0,
    i_13_6_924_0, i_13_6_981_0, i_13_6_988_0, i_13_6_1018_0, i_13_6_1021_0,
    i_13_6_1075_0, i_13_6_1219_0, i_13_6_1262_0, i_13_6_1308_0,
    i_13_6_1342_0, i_13_6_1345_0, i_13_6_1488_0, i_13_6_1496_0,
    i_13_6_1498_0, i_13_6_1515_0, i_13_6_1520_0, i_13_6_1630_0,
    i_13_6_1669_0, i_13_6_1678_0, i_13_6_1730_0, i_13_6_1753_0,
    i_13_6_1773_0, i_13_6_1809_0, i_13_6_1829_0, i_13_6_1854_0,
    i_13_6_1857_0, i_13_6_1858_0, i_13_6_1861_0, i_13_6_2002_0,
    i_13_6_2008_0, i_13_6_2028_0, i_13_6_2191_0, i_13_6_2226_0,
    i_13_6_2452_0, i_13_6_2455_0, i_13_6_2461_0, i_13_6_2539_0,
    i_13_6_2542_0, i_13_6_2544_0, i_13_6_2590_0, i_13_6_2722_0,
    i_13_6_2767_0, i_13_6_2857_0, i_13_6_3007_0, i_13_6_3010_0,
    i_13_6_3012_0, i_13_6_3037_0, i_13_6_3061_0, i_13_6_3064_0,
    i_13_6_3111_0, i_13_6_3127_0, i_13_6_3211_0, i_13_6_3235_0,
    i_13_6_3271_0, i_13_6_3442_0, i_13_6_3487_0, i_13_6_3490_0,
    i_13_6_3508_0, i_13_6_3541_0, i_13_6_3577_0, i_13_6_3640_0,
    i_13_6_3645_0, i_13_6_3729_0, i_13_6_3787_0, i_13_6_3817_0,
    i_13_6_3820_0, i_13_6_3838_0, i_13_6_3856_0, i_13_6_3888_0,
    i_13_6_3889_0, i_13_6_3907_0, i_13_6_3909_0, i_13_6_3910_0,
    i_13_6_3912_0, i_13_6_4078_0, i_13_6_4086_0, i_13_6_4250_0,
    i_13_6_4252_0, i_13_6_4254_0, i_13_6_4255_0, i_13_6_4375_0,
    i_13_6_4378_0, i_13_6_4380_0, i_13_6_4420_0, i_13_6_4426_0,
    i_13_6_4531_0;
  output o_13_6_0_0;
  assign o_13_6_0_0 = ~((i_13_6_229_0 & ((i_13_6_2539_0 & i_13_6_3541_0 & ~i_13_6_3856_0) | (~i_13_6_981_0 & ~i_13_6_3211_0 & ~i_13_6_4254_0 & ~i_13_6_4378_0 & ~i_13_6_4380_0))) | (~i_13_6_418_0 & ((~i_13_6_1018_0 & ~i_13_6_1854_0 & ~i_13_6_1861_0 & ~i_13_6_4250_0) | (~i_13_6_988_0 & ~i_13_6_1773_0 & ~i_13_6_1829_0 & ~i_13_6_2226_0 & ~i_13_6_3909_0 & i_13_6_4252_0))) | (~i_13_6_981_0 & ((~i_13_6_2226_0 & i_13_6_3037_0 & i_13_6_3442_0) | (i_13_6_1021_0 & ~i_13_6_2002_0 & ~i_13_6_3541_0 & ~i_13_6_3912_0))) | (~i_13_6_2028_0 & ((~i_13_6_2461_0 & i_13_6_3235_0) | (~i_13_6_1753_0 & ~i_13_6_1858_0 & ~i_13_6_3912_0 & ~i_13_6_4078_0))) | (~i_13_6_988_0 & ~i_13_6_1075_0 & i_13_6_3211_0) | (~i_13_6_2461_0 & i_13_6_3442_0) | (~i_13_6_574_0 & ~i_13_6_3907_0 & ~i_13_6_3909_0 & ~i_13_6_4254_0 & ~i_13_6_4378_0));
endmodule



// Benchmark "kernel_13_7" written by ABC on Sun Jul 19 10:45:32 2020

module kernel_13_7 ( 
    i_13_7_20_0, i_13_7_38_0, i_13_7_76_0, i_13_7_77_0, i_13_7_158_0,
    i_13_7_166_0, i_13_7_185_0, i_13_7_334_0, i_13_7_337_0, i_13_7_338_0,
    i_13_7_354_0, i_13_7_379_0, i_13_7_407_0, i_13_7_418_0, i_13_7_516_0,
    i_13_7_532_0, i_13_7_545_0, i_13_7_571_0, i_13_7_596_0, i_13_7_597_0,
    i_13_7_641_0, i_13_7_697_0, i_13_7_698_0, i_13_7_699_0, i_13_7_715_0,
    i_13_7_757_0, i_13_7_778_0, i_13_7_834_0, i_13_7_892_0, i_13_7_911_0,
    i_13_7_1067_0, i_13_7_1120_0, i_13_7_1219_0, i_13_7_1224_0,
    i_13_7_1297_0, i_13_7_1298_0, i_13_7_1301_0, i_13_7_1426_0,
    i_13_7_1499_0, i_13_7_1504_0, i_13_7_1523_0, i_13_7_1550_0,
    i_13_7_1558_0, i_13_7_1623_0, i_13_7_1747_0, i_13_7_1757_0,
    i_13_7_1783_0, i_13_7_1814_0, i_13_7_1840_0, i_13_7_1856_0,
    i_13_7_1904_0, i_13_7_1940_0, i_13_7_2116_0, i_13_7_2165_0,
    i_13_7_2169_0, i_13_7_2207_0, i_13_7_2209_0, i_13_7_2210_0,
    i_13_7_2225_0, i_13_7_2236_0, i_13_7_2261_0, i_13_7_2452_0,
    i_13_7_2458_0, i_13_7_2459_0, i_13_7_2549_0, i_13_7_2585_0,
    i_13_7_2639_0, i_13_7_2884_0, i_13_7_2935_0, i_13_7_2939_0,
    i_13_7_2980_0, i_13_7_2981_0, i_13_7_2985_0, i_13_7_3037_0,
    i_13_7_3170_0, i_13_7_3206_0, i_13_7_3217_0, i_13_7_3241_0,
    i_13_7_3290_0, i_13_7_3308_0, i_13_7_3415_0, i_13_7_3424_0,
    i_13_7_3568_0, i_13_7_3640_0, i_13_7_3700_0, i_13_7_3718_0,
    i_13_7_3755_0, i_13_7_3874_0, i_13_7_3908_0, i_13_7_3925_0,
    i_13_7_3987_0, i_13_7_4009_0, i_13_7_4010_0, i_13_7_4052_0,
    i_13_7_4054_0, i_13_7_4060_0, i_13_7_4261_0, i_13_7_4313_0,
    i_13_7_4333_0, i_13_7_4335_0,
    o_13_7_0_0  );
  input  i_13_7_20_0, i_13_7_38_0, i_13_7_76_0, i_13_7_77_0,
    i_13_7_158_0, i_13_7_166_0, i_13_7_185_0, i_13_7_334_0, i_13_7_337_0,
    i_13_7_338_0, i_13_7_354_0, i_13_7_379_0, i_13_7_407_0, i_13_7_418_0,
    i_13_7_516_0, i_13_7_532_0, i_13_7_545_0, i_13_7_571_0, i_13_7_596_0,
    i_13_7_597_0, i_13_7_641_0, i_13_7_697_0, i_13_7_698_0, i_13_7_699_0,
    i_13_7_715_0, i_13_7_757_0, i_13_7_778_0, i_13_7_834_0, i_13_7_892_0,
    i_13_7_911_0, i_13_7_1067_0, i_13_7_1120_0, i_13_7_1219_0,
    i_13_7_1224_0, i_13_7_1297_0, i_13_7_1298_0, i_13_7_1301_0,
    i_13_7_1426_0, i_13_7_1499_0, i_13_7_1504_0, i_13_7_1523_0,
    i_13_7_1550_0, i_13_7_1558_0, i_13_7_1623_0, i_13_7_1747_0,
    i_13_7_1757_0, i_13_7_1783_0, i_13_7_1814_0, i_13_7_1840_0,
    i_13_7_1856_0, i_13_7_1904_0, i_13_7_1940_0, i_13_7_2116_0,
    i_13_7_2165_0, i_13_7_2169_0, i_13_7_2207_0, i_13_7_2209_0,
    i_13_7_2210_0, i_13_7_2225_0, i_13_7_2236_0, i_13_7_2261_0,
    i_13_7_2452_0, i_13_7_2458_0, i_13_7_2459_0, i_13_7_2549_0,
    i_13_7_2585_0, i_13_7_2639_0, i_13_7_2884_0, i_13_7_2935_0,
    i_13_7_2939_0, i_13_7_2980_0, i_13_7_2981_0, i_13_7_2985_0,
    i_13_7_3037_0, i_13_7_3170_0, i_13_7_3206_0, i_13_7_3217_0,
    i_13_7_3241_0, i_13_7_3290_0, i_13_7_3308_0, i_13_7_3415_0,
    i_13_7_3424_0, i_13_7_3568_0, i_13_7_3640_0, i_13_7_3700_0,
    i_13_7_3718_0, i_13_7_3755_0, i_13_7_3874_0, i_13_7_3908_0,
    i_13_7_3925_0, i_13_7_3987_0, i_13_7_4009_0, i_13_7_4010_0,
    i_13_7_4052_0, i_13_7_4054_0, i_13_7_4060_0, i_13_7_4261_0,
    i_13_7_4313_0, i_13_7_4333_0, i_13_7_4335_0;
  output o_13_7_0_0;
  assign o_13_7_0_0 = ~((~i_13_7_1301_0 & ((~i_13_7_337_0 & ~i_13_7_4060_0) | (~i_13_7_185_0 & ~i_13_7_2458_0 & ~i_13_7_2980_0 & ~i_13_7_4313_0))) | (~i_13_7_1840_0 & ((i_13_7_1426_0 & ~i_13_7_4052_0) | (~i_13_7_3206_0 & ~i_13_7_3217_0 & ~i_13_7_4313_0))) | (~i_13_7_2935_0 & (i_13_7_698_0 | (~i_13_7_1120_0 & i_13_7_2452_0) | (~i_13_7_334_0 & ~i_13_7_1499_0 & ~i_13_7_3290_0))) | (i_13_7_76_0 & ~i_13_7_2209_0 & ~i_13_7_3206_0) | (i_13_7_337_0 & ~i_13_7_2236_0 & i_13_7_2884_0 & i_13_7_3874_0));
endmodule



// Benchmark "kernel_13_8" written by ABC on Sun Jul 19 10:45:32 2020

module kernel_13_8 ( 
    i_13_8_65_0, i_13_8_101_0, i_13_8_207_0, i_13_8_208_0, i_13_8_209_0,
    i_13_8_266_0, i_13_8_273_0, i_13_8_355_0, i_13_8_371_0, i_13_8_415_0,
    i_13_8_416_0, i_13_8_463_0, i_13_8_464_0, i_13_8_567_0, i_13_8_614_0,
    i_13_8_671_0, i_13_8_761_0, i_13_8_948_0, i_13_8_950_0, i_13_8_956_0,
    i_13_8_1081_0, i_13_8_1129_0, i_13_8_1319_0, i_13_8_1372_0,
    i_13_8_1504_0, i_13_8_1522_0, i_13_8_1523_0, i_13_8_1553_0,
    i_13_8_1604_0, i_13_8_1640_0, i_13_8_1687_0, i_13_8_1697_0,
    i_13_8_1786_0, i_13_8_1827_0, i_13_8_1830_0, i_13_8_1840_0,
    i_13_8_1841_0, i_13_8_1846_0, i_13_8_1847_0, i_13_8_1930_0,
    i_13_8_1931_0, i_13_8_1958_0, i_13_8_2056_0, i_13_8_2143_0,
    i_13_8_2200_0, i_13_8_2201_0, i_13_8_2237_0, i_13_8_2297_0,
    i_13_8_2399_0, i_13_8_2403_0, i_13_8_2444_0, i_13_8_2563_0,
    i_13_8_2692_0, i_13_8_2821_0, i_13_8_2822_0, i_13_8_3001_0,
    i_13_8_3045_0, i_13_8_3062_0, i_13_8_3164_0, i_13_8_3234_0,
    i_13_8_3240_0, i_13_8_3241_0, i_13_8_3242_0, i_13_8_3259_0,
    i_13_8_3261_0, i_13_8_3308_0, i_13_8_3343_0, i_13_8_3344_0,
    i_13_8_3388_0, i_13_8_3519_0, i_13_8_3538_0, i_13_8_3618_0,
    i_13_8_3619_0, i_13_8_3620_0, i_13_8_3631_0, i_13_8_3632_0,
    i_13_8_3637_0, i_13_8_3638_0, i_13_8_3857_0, i_13_8_3873_0,
    i_13_8_3904_0, i_13_8_3916_0, i_13_8_3928_0, i_13_8_3935_0,
    i_13_8_3988_0, i_13_8_3989_0, i_13_8_3992_0, i_13_8_4008_0,
    i_13_8_4061_0, i_13_8_4118_0, i_13_8_4205_0, i_13_8_4270_0,
    i_13_8_4271_0, i_13_8_4302_0, i_13_8_4312_0, i_13_8_4313_0,
    i_13_8_4339_0, i_13_8_4378_0, i_13_8_4477_0, i_13_8_4536_0,
    o_13_8_0_0  );
  input  i_13_8_65_0, i_13_8_101_0, i_13_8_207_0, i_13_8_208_0,
    i_13_8_209_0, i_13_8_266_0, i_13_8_273_0, i_13_8_355_0, i_13_8_371_0,
    i_13_8_415_0, i_13_8_416_0, i_13_8_463_0, i_13_8_464_0, i_13_8_567_0,
    i_13_8_614_0, i_13_8_671_0, i_13_8_761_0, i_13_8_948_0, i_13_8_950_0,
    i_13_8_956_0, i_13_8_1081_0, i_13_8_1129_0, i_13_8_1319_0,
    i_13_8_1372_0, i_13_8_1504_0, i_13_8_1522_0, i_13_8_1523_0,
    i_13_8_1553_0, i_13_8_1604_0, i_13_8_1640_0, i_13_8_1687_0,
    i_13_8_1697_0, i_13_8_1786_0, i_13_8_1827_0, i_13_8_1830_0,
    i_13_8_1840_0, i_13_8_1841_0, i_13_8_1846_0, i_13_8_1847_0,
    i_13_8_1930_0, i_13_8_1931_0, i_13_8_1958_0, i_13_8_2056_0,
    i_13_8_2143_0, i_13_8_2200_0, i_13_8_2201_0, i_13_8_2237_0,
    i_13_8_2297_0, i_13_8_2399_0, i_13_8_2403_0, i_13_8_2444_0,
    i_13_8_2563_0, i_13_8_2692_0, i_13_8_2821_0, i_13_8_2822_0,
    i_13_8_3001_0, i_13_8_3045_0, i_13_8_3062_0, i_13_8_3164_0,
    i_13_8_3234_0, i_13_8_3240_0, i_13_8_3241_0, i_13_8_3242_0,
    i_13_8_3259_0, i_13_8_3261_0, i_13_8_3308_0, i_13_8_3343_0,
    i_13_8_3344_0, i_13_8_3388_0, i_13_8_3519_0, i_13_8_3538_0,
    i_13_8_3618_0, i_13_8_3619_0, i_13_8_3620_0, i_13_8_3631_0,
    i_13_8_3632_0, i_13_8_3637_0, i_13_8_3638_0, i_13_8_3857_0,
    i_13_8_3873_0, i_13_8_3904_0, i_13_8_3916_0, i_13_8_3928_0,
    i_13_8_3935_0, i_13_8_3988_0, i_13_8_3989_0, i_13_8_3992_0,
    i_13_8_4008_0, i_13_8_4061_0, i_13_8_4118_0, i_13_8_4205_0,
    i_13_8_4270_0, i_13_8_4271_0, i_13_8_4302_0, i_13_8_4312_0,
    i_13_8_4313_0, i_13_8_4339_0, i_13_8_4378_0, i_13_8_4477_0,
    i_13_8_4536_0;
  output o_13_8_0_0;
  assign o_13_8_0_0 = ~(~i_13_8_2237_0 | ~i_13_8_416_0 | ~i_13_8_1522_0);
endmodule



// Benchmark "kernel_13_9" written by ABC on Sun Jul 19 10:45:33 2020

module kernel_13_9 ( 
    i_13_9_48_0, i_13_9_73_0, i_13_9_94_0, i_13_9_173_0, i_13_9_193_0,
    i_13_9_225_0, i_13_9_280_0, i_13_9_391_0, i_13_9_443_0, i_13_9_451_0,
    i_13_9_515_0, i_13_9_533_0, i_13_9_550_0, i_13_9_551_0, i_13_9_553_0,
    i_13_9_645_0, i_13_9_651_0, i_13_9_652_0, i_13_9_655_0, i_13_9_656_0,
    i_13_9_658_0, i_13_9_668_0, i_13_9_675_0, i_13_9_676_0, i_13_9_685_0,
    i_13_9_688_0, i_13_9_691_0, i_13_9_830_0, i_13_9_841_0, i_13_9_949_0,
    i_13_9_1098_0, i_13_9_1117_0, i_13_9_1144_0, i_13_9_1191_0,
    i_13_9_1267_0, i_13_9_1270_0, i_13_9_1305_0, i_13_9_1347_0,
    i_13_9_1383_0, i_13_9_1384_0, i_13_9_1404_0, i_13_9_1465_0,
    i_13_9_1515_0, i_13_9_1518_0, i_13_9_1773_0, i_13_9_1774_0,
    i_13_9_1777_0, i_13_9_1836_0, i_13_9_1858_0, i_13_9_1909_0,
    i_13_9_2046_0, i_13_9_2049_0, i_13_9_2058_0, i_13_9_2191_0,
    i_13_9_2351_0, i_13_9_2503_0, i_13_9_2511_0, i_13_9_2581_0,
    i_13_9_2627_0, i_13_9_2650_0, i_13_9_2749_0, i_13_9_2857_0,
    i_13_9_2999_0, i_13_9_3000_0, i_13_9_3037_0, i_13_9_3062_0,
    i_13_9_3087_0, i_13_9_3101_0, i_13_9_3214_0, i_13_9_3216_0,
    i_13_9_3235_0, i_13_9_3367_0, i_13_9_3371_0, i_13_9_3418_0,
    i_13_9_3532_0, i_13_9_3646_0, i_13_9_3863_0, i_13_9_3865_0,
    i_13_9_3888_0, i_13_9_3889_0, i_13_9_3890_0, i_13_9_3987_0,
    i_13_9_3988_0, i_13_9_3989_0, i_13_9_4018_0, i_13_9_4051_0,
    i_13_9_4054_0, i_13_9_4117_0, i_13_9_4122_0, i_13_9_4189_0,
    i_13_9_4233_0, i_13_9_4263_0, i_13_9_4305_0, i_13_9_4330_0,
    i_13_9_4366_0, i_13_9_4539_0, i_13_9_4594_0, i_13_9_4600_0,
    i_13_9_4601_0, i_13_9_4603_0,
    o_13_9_0_0  );
  input  i_13_9_48_0, i_13_9_73_0, i_13_9_94_0, i_13_9_173_0,
    i_13_9_193_0, i_13_9_225_0, i_13_9_280_0, i_13_9_391_0, i_13_9_443_0,
    i_13_9_451_0, i_13_9_515_0, i_13_9_533_0, i_13_9_550_0, i_13_9_551_0,
    i_13_9_553_0, i_13_9_645_0, i_13_9_651_0, i_13_9_652_0, i_13_9_655_0,
    i_13_9_656_0, i_13_9_658_0, i_13_9_668_0, i_13_9_675_0, i_13_9_676_0,
    i_13_9_685_0, i_13_9_688_0, i_13_9_691_0, i_13_9_830_0, i_13_9_841_0,
    i_13_9_949_0, i_13_9_1098_0, i_13_9_1117_0, i_13_9_1144_0,
    i_13_9_1191_0, i_13_9_1267_0, i_13_9_1270_0, i_13_9_1305_0,
    i_13_9_1347_0, i_13_9_1383_0, i_13_9_1384_0, i_13_9_1404_0,
    i_13_9_1465_0, i_13_9_1515_0, i_13_9_1518_0, i_13_9_1773_0,
    i_13_9_1774_0, i_13_9_1777_0, i_13_9_1836_0, i_13_9_1858_0,
    i_13_9_1909_0, i_13_9_2046_0, i_13_9_2049_0, i_13_9_2058_0,
    i_13_9_2191_0, i_13_9_2351_0, i_13_9_2503_0, i_13_9_2511_0,
    i_13_9_2581_0, i_13_9_2627_0, i_13_9_2650_0, i_13_9_2749_0,
    i_13_9_2857_0, i_13_9_2999_0, i_13_9_3000_0, i_13_9_3037_0,
    i_13_9_3062_0, i_13_9_3087_0, i_13_9_3101_0, i_13_9_3214_0,
    i_13_9_3216_0, i_13_9_3235_0, i_13_9_3367_0, i_13_9_3371_0,
    i_13_9_3418_0, i_13_9_3532_0, i_13_9_3646_0, i_13_9_3863_0,
    i_13_9_3865_0, i_13_9_3888_0, i_13_9_3889_0, i_13_9_3890_0,
    i_13_9_3987_0, i_13_9_3988_0, i_13_9_3989_0, i_13_9_4018_0,
    i_13_9_4051_0, i_13_9_4054_0, i_13_9_4117_0, i_13_9_4122_0,
    i_13_9_4189_0, i_13_9_4233_0, i_13_9_4263_0, i_13_9_4305_0,
    i_13_9_4330_0, i_13_9_4366_0, i_13_9_4539_0, i_13_9_4594_0,
    i_13_9_4600_0, i_13_9_4601_0, i_13_9_4603_0;
  output o_13_9_0_0;
  assign o_13_9_0_0 = ~((i_13_9_949_0 & i_13_9_4305_0) | (~i_13_9_688_0 & ~i_13_9_3988_0) | (~i_13_9_675_0 & ~i_13_9_676_0 & ~i_13_9_4330_0) | (~i_13_9_652_0 & ~i_13_9_3889_0 & ~i_13_9_3890_0));
endmodule



// Benchmark "kernel_13_10" written by ABC on Sun Jul 19 10:45:34 2020

module kernel_13_10 ( 
    i_13_10_34_0, i_13_10_43_0, i_13_10_69_0, i_13_10_70_0, i_13_10_322_0,
    i_13_10_384_0, i_13_10_411_0, i_13_10_421_0, i_13_10_426_0,
    i_13_10_448_0, i_13_10_463_0, i_13_10_467_0, i_13_10_493_0,
    i_13_10_525_0, i_13_10_538_0, i_13_10_591_0, i_13_10_619_0,
    i_13_10_628_0, i_13_10_646_0, i_13_10_679_0, i_13_10_762_0,
    i_13_10_763_0, i_13_10_931_0, i_13_10_934_0, i_13_10_943_0,
    i_13_10_1021_0, i_13_10_1083_0, i_13_10_1096_0, i_13_10_1104_0,
    i_13_10_1105_0, i_13_10_1123_0, i_13_10_1131_0, i_13_10_1132_0,
    i_13_10_1347_0, i_13_10_1473_0, i_13_10_1510_0, i_13_10_1536_0,
    i_13_10_1537_0, i_13_10_1795_0, i_13_10_1797_0, i_13_10_1798_0,
    i_13_10_1803_0, i_13_10_1912_0, i_13_10_2001_0, i_13_10_2002_0,
    i_13_10_2023_0, i_13_10_2044_0, i_13_10_2048_0, i_13_10_2055_0,
    i_13_10_2231_0, i_13_10_2472_0, i_13_10_2508_0, i_13_10_2551_0,
    i_13_10_2599_0, i_13_10_2680_0, i_13_10_2724_0, i_13_10_2850_0,
    i_13_10_2859_0, i_13_10_2860_0, i_13_10_2904_0, i_13_10_2998_0,
    i_13_10_3030_0, i_13_10_3094_0, i_13_10_3127_0, i_13_10_3131_0,
    i_13_10_3155_0, i_13_10_3262_0, i_13_10_3264_0, i_13_10_3370_0,
    i_13_10_3390_0, i_13_10_3391_0, i_13_10_3417_0, i_13_10_3445_0,
    i_13_10_3558_0, i_13_10_3639_0, i_13_10_3640_0, i_13_10_3643_0,
    i_13_10_3649_0, i_13_10_3652_0, i_13_10_3680_0, i_13_10_3730_0,
    i_13_10_3769_0, i_13_10_3799_0, i_13_10_3847_0, i_13_10_3892_0,
    i_13_10_4021_0, i_13_10_4038_0, i_13_10_4039_0, i_13_10_4057_0,
    i_13_10_4084_0, i_13_10_4117_0, i_13_10_4166_0, i_13_10_4398_0,
    i_13_10_4408_0, i_13_10_4435_0, i_13_10_4541_0, i_13_10_4586_0,
    i_13_10_4596_0, i_13_10_4597_0, i_13_10_4606_0,
    o_13_10_0_0  );
  input  i_13_10_34_0, i_13_10_43_0, i_13_10_69_0, i_13_10_70_0,
    i_13_10_322_0, i_13_10_384_0, i_13_10_411_0, i_13_10_421_0,
    i_13_10_426_0, i_13_10_448_0, i_13_10_463_0, i_13_10_467_0,
    i_13_10_493_0, i_13_10_525_0, i_13_10_538_0, i_13_10_591_0,
    i_13_10_619_0, i_13_10_628_0, i_13_10_646_0, i_13_10_679_0,
    i_13_10_762_0, i_13_10_763_0, i_13_10_931_0, i_13_10_934_0,
    i_13_10_943_0, i_13_10_1021_0, i_13_10_1083_0, i_13_10_1096_0,
    i_13_10_1104_0, i_13_10_1105_0, i_13_10_1123_0, i_13_10_1131_0,
    i_13_10_1132_0, i_13_10_1347_0, i_13_10_1473_0, i_13_10_1510_0,
    i_13_10_1536_0, i_13_10_1537_0, i_13_10_1795_0, i_13_10_1797_0,
    i_13_10_1798_0, i_13_10_1803_0, i_13_10_1912_0, i_13_10_2001_0,
    i_13_10_2002_0, i_13_10_2023_0, i_13_10_2044_0, i_13_10_2048_0,
    i_13_10_2055_0, i_13_10_2231_0, i_13_10_2472_0, i_13_10_2508_0,
    i_13_10_2551_0, i_13_10_2599_0, i_13_10_2680_0, i_13_10_2724_0,
    i_13_10_2850_0, i_13_10_2859_0, i_13_10_2860_0, i_13_10_2904_0,
    i_13_10_2998_0, i_13_10_3030_0, i_13_10_3094_0, i_13_10_3127_0,
    i_13_10_3131_0, i_13_10_3155_0, i_13_10_3262_0, i_13_10_3264_0,
    i_13_10_3370_0, i_13_10_3390_0, i_13_10_3391_0, i_13_10_3417_0,
    i_13_10_3445_0, i_13_10_3558_0, i_13_10_3639_0, i_13_10_3640_0,
    i_13_10_3643_0, i_13_10_3649_0, i_13_10_3652_0, i_13_10_3680_0,
    i_13_10_3730_0, i_13_10_3769_0, i_13_10_3799_0, i_13_10_3847_0,
    i_13_10_3892_0, i_13_10_4021_0, i_13_10_4038_0, i_13_10_4039_0,
    i_13_10_4057_0, i_13_10_4084_0, i_13_10_4117_0, i_13_10_4166_0,
    i_13_10_4398_0, i_13_10_4408_0, i_13_10_4435_0, i_13_10_4541_0,
    i_13_10_4586_0, i_13_10_4596_0, i_13_10_4597_0, i_13_10_4606_0;
  output o_13_10_0_0;
  assign o_13_10_0_0 = ~((i_13_10_931_0 & ~i_13_10_4057_0) | (~i_13_10_3390_0 & ~i_13_10_4039_0) | (~i_13_10_538_0 & ~i_13_10_762_0 & ~i_13_10_1798_0));
endmodule



// Benchmark "kernel_13_11" written by ABC on Sun Jul 19 10:45:35 2020

module kernel_13_11 ( 
    i_13_11_45_0, i_13_11_69_0, i_13_11_76_0, i_13_11_93_0, i_13_11_127_0,
    i_13_11_384_0, i_13_11_385_0, i_13_11_411_0, i_13_11_462_0,
    i_13_11_537_0, i_13_11_564_0, i_13_11_603_0, i_13_11_645_0,
    i_13_11_682_0, i_13_11_825_0, i_13_11_882_0, i_13_11_933_0,
    i_13_11_1080_0, i_13_11_1086_0, i_13_11_1104_0, i_13_11_1341_0,
    i_13_11_1342_0, i_13_11_1401_0, i_13_11_1402_0, i_13_11_1468_0,
    i_13_11_1473_0, i_13_11_1479_0, i_13_11_1509_0, i_13_11_1510_0,
    i_13_11_1599_0, i_13_11_1600_0, i_13_11_1644_0, i_13_11_1657_0,
    i_13_11_1716_0, i_13_11_1717_0, i_13_11_1725_0, i_13_11_1728_0,
    i_13_11_1780_0, i_13_11_1797_0, i_13_11_1941_0, i_13_11_1995_0,
    i_13_11_1996_0, i_13_11_2053_0, i_13_11_2058_0, i_13_11_2176_0,
    i_13_11_2187_0, i_13_11_2188_0, i_13_11_2193_0, i_13_11_2265_0,
    i_13_11_2275_0, i_13_11_2277_0, i_13_11_2278_0, i_13_11_2304_0,
    i_13_11_2305_0, i_13_11_2340_0, i_13_11_2341_0, i_13_11_2424_0,
    i_13_11_2679_0, i_13_11_2725_0, i_13_11_2919_0, i_13_11_3066_0,
    i_13_11_3067_0, i_13_11_3102_0, i_13_11_3103_0, i_13_11_3147_0,
    i_13_11_3234_0, i_13_11_3289_0, i_13_11_3366_0, i_13_11_3394_0,
    i_13_11_3410_0, i_13_11_3441_0, i_13_11_3525_0, i_13_11_3555_0,
    i_13_11_3556_0, i_13_11_3580_0, i_13_11_3687_0, i_13_11_3688_0,
    i_13_11_3729_0, i_13_11_3730_0, i_13_11_3742_0, i_13_11_3786_0,
    i_13_11_3787_0, i_13_11_3796_0, i_13_11_3805_0, i_13_11_3816_0,
    i_13_11_3817_0, i_13_11_3894_0, i_13_11_3930_0, i_13_11_3991_0,
    i_13_11_3993_0, i_13_11_3994_0, i_13_11_4056_0, i_13_11_4057_0,
    i_13_11_4065_0, i_13_11_4093_0, i_13_11_4119_0, i_13_11_4166_0,
    i_13_11_4257_0, i_13_11_4393_0, i_13_11_4399_0,
    o_13_11_0_0  );
  input  i_13_11_45_0, i_13_11_69_0, i_13_11_76_0, i_13_11_93_0,
    i_13_11_127_0, i_13_11_384_0, i_13_11_385_0, i_13_11_411_0,
    i_13_11_462_0, i_13_11_537_0, i_13_11_564_0, i_13_11_603_0,
    i_13_11_645_0, i_13_11_682_0, i_13_11_825_0, i_13_11_882_0,
    i_13_11_933_0, i_13_11_1080_0, i_13_11_1086_0, i_13_11_1104_0,
    i_13_11_1341_0, i_13_11_1342_0, i_13_11_1401_0, i_13_11_1402_0,
    i_13_11_1468_0, i_13_11_1473_0, i_13_11_1479_0, i_13_11_1509_0,
    i_13_11_1510_0, i_13_11_1599_0, i_13_11_1600_0, i_13_11_1644_0,
    i_13_11_1657_0, i_13_11_1716_0, i_13_11_1717_0, i_13_11_1725_0,
    i_13_11_1728_0, i_13_11_1780_0, i_13_11_1797_0, i_13_11_1941_0,
    i_13_11_1995_0, i_13_11_1996_0, i_13_11_2053_0, i_13_11_2058_0,
    i_13_11_2176_0, i_13_11_2187_0, i_13_11_2188_0, i_13_11_2193_0,
    i_13_11_2265_0, i_13_11_2275_0, i_13_11_2277_0, i_13_11_2278_0,
    i_13_11_2304_0, i_13_11_2305_0, i_13_11_2340_0, i_13_11_2341_0,
    i_13_11_2424_0, i_13_11_2679_0, i_13_11_2725_0, i_13_11_2919_0,
    i_13_11_3066_0, i_13_11_3067_0, i_13_11_3102_0, i_13_11_3103_0,
    i_13_11_3147_0, i_13_11_3234_0, i_13_11_3289_0, i_13_11_3366_0,
    i_13_11_3394_0, i_13_11_3410_0, i_13_11_3441_0, i_13_11_3525_0,
    i_13_11_3555_0, i_13_11_3556_0, i_13_11_3580_0, i_13_11_3687_0,
    i_13_11_3688_0, i_13_11_3729_0, i_13_11_3730_0, i_13_11_3742_0,
    i_13_11_3786_0, i_13_11_3787_0, i_13_11_3796_0, i_13_11_3805_0,
    i_13_11_3816_0, i_13_11_3817_0, i_13_11_3894_0, i_13_11_3930_0,
    i_13_11_3991_0, i_13_11_3993_0, i_13_11_3994_0, i_13_11_4056_0,
    i_13_11_4057_0, i_13_11_4065_0, i_13_11_4093_0, i_13_11_4119_0,
    i_13_11_4166_0, i_13_11_4257_0, i_13_11_4393_0, i_13_11_4399_0;
  output o_13_11_0_0;
  assign o_13_11_0_0 = ~((~i_13_11_69_0 & ~i_13_11_3688_0) | (i_13_11_3580_0 & i_13_11_3688_0) | (~i_13_11_3441_0 & ~i_13_11_3525_0 & ~i_13_11_4166_0) | (~i_13_11_1401_0 & ~i_13_11_1510_0 & ~i_13_11_3066_0));
endmodule



// Benchmark "kernel_13_12" written by ABC on Sun Jul 19 10:45:36 2020

module kernel_13_12 ( 
    i_13_12_60_0, i_13_12_90_0, i_13_12_91_0, i_13_12_93_0, i_13_12_94_0,
    i_13_12_97_0, i_13_12_126_0, i_13_12_174_0, i_13_12_175_0,
    i_13_12_184_0, i_13_12_280_0, i_13_12_282_0, i_13_12_307_0,
    i_13_12_310_0, i_13_12_315_0, i_13_12_316_0, i_13_12_328_0,
    i_13_12_516_0, i_13_12_570_0, i_13_12_571_0, i_13_12_599_0,
    i_13_12_616_0, i_13_12_661_0, i_13_12_667_0, i_13_12_697_0,
    i_13_12_759_0, i_13_12_981_0, i_13_12_982_0, i_13_12_1020_0,
    i_13_12_1226_0, i_13_12_1256_0, i_13_12_1305_0, i_13_12_1323_0,
    i_13_12_1404_0, i_13_12_1426_0, i_13_12_1440_0, i_13_12_1441_0,
    i_13_12_1446_0, i_13_12_1494_0, i_13_12_1515_0, i_13_12_1629_0,
    i_13_12_1669_0, i_13_12_1769_0, i_13_12_1777_0, i_13_12_1828_0,
    i_13_12_1848_0, i_13_12_1849_0, i_13_12_1859_0, i_13_12_1885_0,
    i_13_12_1908_0, i_13_12_1921_0, i_13_12_1998_0, i_13_12_2003_0,
    i_13_12_2116_0, i_13_12_2172_0, i_13_12_2173_0, i_13_12_2407_0,
    i_13_12_2421_0, i_13_12_2676_0, i_13_12_2692_0, i_13_12_2875_0,
    i_13_12_2983_0, i_13_12_3026_0, i_13_12_3109_0, i_13_12_3163_0,
    i_13_12_3207_0, i_13_12_3241_0, i_13_12_3263_0, i_13_12_3327_0,
    i_13_12_3420_0, i_13_12_3421_0, i_13_12_3471_0, i_13_12_3478_0,
    i_13_12_3529_0, i_13_12_3556_0, i_13_12_3568_0, i_13_12_3575_0,
    i_13_12_3756_0, i_13_12_3765_0, i_13_12_3766_0, i_13_12_3782_0,
    i_13_12_3817_0, i_13_12_3844_0, i_13_12_3864_0, i_13_12_3871_0,
    i_13_12_3888_0, i_13_12_4037_0, i_13_12_4060_0, i_13_12_4066_0,
    i_13_12_4080_0, i_13_12_4163_0, i_13_12_4252_0, i_13_12_4316_0,
    i_13_12_4350_0, i_13_12_4351_0, i_13_12_4452_0, i_13_12_4469_0,
    i_13_12_4566_0, i_13_12_4567_0, i_13_12_4601_0,
    o_13_12_0_0  );
  input  i_13_12_60_0, i_13_12_90_0, i_13_12_91_0, i_13_12_93_0,
    i_13_12_94_0, i_13_12_97_0, i_13_12_126_0, i_13_12_174_0,
    i_13_12_175_0, i_13_12_184_0, i_13_12_280_0, i_13_12_282_0,
    i_13_12_307_0, i_13_12_310_0, i_13_12_315_0, i_13_12_316_0,
    i_13_12_328_0, i_13_12_516_0, i_13_12_570_0, i_13_12_571_0,
    i_13_12_599_0, i_13_12_616_0, i_13_12_661_0, i_13_12_667_0,
    i_13_12_697_0, i_13_12_759_0, i_13_12_981_0, i_13_12_982_0,
    i_13_12_1020_0, i_13_12_1226_0, i_13_12_1256_0, i_13_12_1305_0,
    i_13_12_1323_0, i_13_12_1404_0, i_13_12_1426_0, i_13_12_1440_0,
    i_13_12_1441_0, i_13_12_1446_0, i_13_12_1494_0, i_13_12_1515_0,
    i_13_12_1629_0, i_13_12_1669_0, i_13_12_1769_0, i_13_12_1777_0,
    i_13_12_1828_0, i_13_12_1848_0, i_13_12_1849_0, i_13_12_1859_0,
    i_13_12_1885_0, i_13_12_1908_0, i_13_12_1921_0, i_13_12_1998_0,
    i_13_12_2003_0, i_13_12_2116_0, i_13_12_2172_0, i_13_12_2173_0,
    i_13_12_2407_0, i_13_12_2421_0, i_13_12_2676_0, i_13_12_2692_0,
    i_13_12_2875_0, i_13_12_2983_0, i_13_12_3026_0, i_13_12_3109_0,
    i_13_12_3163_0, i_13_12_3207_0, i_13_12_3241_0, i_13_12_3263_0,
    i_13_12_3327_0, i_13_12_3420_0, i_13_12_3421_0, i_13_12_3471_0,
    i_13_12_3478_0, i_13_12_3529_0, i_13_12_3556_0, i_13_12_3568_0,
    i_13_12_3575_0, i_13_12_3756_0, i_13_12_3765_0, i_13_12_3766_0,
    i_13_12_3782_0, i_13_12_3817_0, i_13_12_3844_0, i_13_12_3864_0,
    i_13_12_3871_0, i_13_12_3888_0, i_13_12_4037_0, i_13_12_4060_0,
    i_13_12_4066_0, i_13_12_4080_0, i_13_12_4163_0, i_13_12_4252_0,
    i_13_12_4316_0, i_13_12_4350_0, i_13_12_4351_0, i_13_12_4452_0,
    i_13_12_4469_0, i_13_12_4566_0, i_13_12_4567_0, i_13_12_4601_0;
  output o_13_12_0_0;
  assign o_13_12_0_0 = ~(i_13_12_516_0 | (~i_13_12_90_0 & ~i_13_12_3765_0) | (~i_13_12_316_0 & i_13_12_1426_0) | (~i_13_12_981_0 & ~i_13_12_2692_0 & ~i_13_12_3241_0 & ~i_13_12_3817_0));
endmodule



// Benchmark "kernel_13_13" written by ABC on Sun Jul 19 10:45:37 2020

module kernel_13_13 ( 
    i_13_13_48_0, i_13_13_49_0, i_13_13_70_0, i_13_13_76_0, i_13_13_106_0,
    i_13_13_127_0, i_13_13_229_0, i_13_13_270_0, i_13_13_271_0,
    i_13_13_313_0, i_13_13_369_0, i_13_13_411_0, i_13_13_447_0,
    i_13_13_475_0, i_13_13_561_0, i_13_13_564_0, i_13_13_565_0,
    i_13_13_620_0, i_13_13_663_0, i_13_13_673_0, i_13_13_732_0,
    i_13_13_736_0, i_13_13_745_0, i_13_13_834_0, i_13_13_835_0,
    i_13_13_934_0, i_13_13_946_0, i_13_13_952_0, i_13_13_1043_0,
    i_13_13_1087_0, i_13_13_1104_0, i_13_13_1131_0, i_13_13_1150_0,
    i_13_13_1231_0, i_13_13_1232_0, i_13_13_1246_0, i_13_13_1402_0,
    i_13_13_1431_0, i_13_13_1465_0, i_13_13_1468_0, i_13_13_1497_0,
    i_13_13_1537_0, i_13_13_1566_0, i_13_13_1626_0, i_13_13_1657_0,
    i_13_13_1663_0, i_13_13_1729_0, i_13_13_1732_0, i_13_13_1735_0,
    i_13_13_1764_0, i_13_13_1765_0, i_13_13_1767_0, i_13_13_1797_0,
    i_13_13_1798_0, i_13_13_1805_0, i_13_13_1894_0, i_13_13_1947_0,
    i_13_13_2022_0, i_13_13_2029_0, i_13_13_2107_0, i_13_13_2175_0,
    i_13_13_2208_0, i_13_13_2223_0, i_13_13_2224_0, i_13_13_2436_0,
    i_13_13_2564_0, i_13_13_2709_0, i_13_13_2724_0, i_13_13_2754_0,
    i_13_13_2955_0, i_13_13_2968_0, i_13_13_3217_0, i_13_13_3258_0,
    i_13_13_3259_0, i_13_13_3264_0, i_13_13_3283_0, i_13_13_3354_0,
    i_13_13_3370_0, i_13_13_3478_0, i_13_13_3520_0, i_13_13_3536_0,
    i_13_13_3551_0, i_13_13_3757_0, i_13_13_3783_0, i_13_13_3900_0,
    i_13_13_3918_0, i_13_13_3930_0, i_13_13_4038_0, i_13_13_4045_0,
    i_13_13_4083_0, i_13_13_4164_0, i_13_13_4165_0, i_13_13_4189_0,
    i_13_13_4233_0, i_13_13_4269_0, i_13_13_4296_0, i_13_13_4324_0,
    i_13_13_4372_0, i_13_13_4513_0, i_13_13_4606_0,
    o_13_13_0_0  );
  input  i_13_13_48_0, i_13_13_49_0, i_13_13_70_0, i_13_13_76_0,
    i_13_13_106_0, i_13_13_127_0, i_13_13_229_0, i_13_13_270_0,
    i_13_13_271_0, i_13_13_313_0, i_13_13_369_0, i_13_13_411_0,
    i_13_13_447_0, i_13_13_475_0, i_13_13_561_0, i_13_13_564_0,
    i_13_13_565_0, i_13_13_620_0, i_13_13_663_0, i_13_13_673_0,
    i_13_13_732_0, i_13_13_736_0, i_13_13_745_0, i_13_13_834_0,
    i_13_13_835_0, i_13_13_934_0, i_13_13_946_0, i_13_13_952_0,
    i_13_13_1043_0, i_13_13_1087_0, i_13_13_1104_0, i_13_13_1131_0,
    i_13_13_1150_0, i_13_13_1231_0, i_13_13_1232_0, i_13_13_1246_0,
    i_13_13_1402_0, i_13_13_1431_0, i_13_13_1465_0, i_13_13_1468_0,
    i_13_13_1497_0, i_13_13_1537_0, i_13_13_1566_0, i_13_13_1626_0,
    i_13_13_1657_0, i_13_13_1663_0, i_13_13_1729_0, i_13_13_1732_0,
    i_13_13_1735_0, i_13_13_1764_0, i_13_13_1765_0, i_13_13_1767_0,
    i_13_13_1797_0, i_13_13_1798_0, i_13_13_1805_0, i_13_13_1894_0,
    i_13_13_1947_0, i_13_13_2022_0, i_13_13_2029_0, i_13_13_2107_0,
    i_13_13_2175_0, i_13_13_2208_0, i_13_13_2223_0, i_13_13_2224_0,
    i_13_13_2436_0, i_13_13_2564_0, i_13_13_2709_0, i_13_13_2724_0,
    i_13_13_2754_0, i_13_13_2955_0, i_13_13_2968_0, i_13_13_3217_0,
    i_13_13_3258_0, i_13_13_3259_0, i_13_13_3264_0, i_13_13_3283_0,
    i_13_13_3354_0, i_13_13_3370_0, i_13_13_3478_0, i_13_13_3520_0,
    i_13_13_3536_0, i_13_13_3551_0, i_13_13_3757_0, i_13_13_3783_0,
    i_13_13_3900_0, i_13_13_3918_0, i_13_13_3930_0, i_13_13_4038_0,
    i_13_13_4045_0, i_13_13_4083_0, i_13_13_4164_0, i_13_13_4165_0,
    i_13_13_4189_0, i_13_13_4233_0, i_13_13_4269_0, i_13_13_4296_0,
    i_13_13_4324_0, i_13_13_4372_0, i_13_13_4513_0, i_13_13_4606_0;
  output o_13_13_0_0;
  assign o_13_13_0_0 = ~(~i_13_13_4165_0 | (~i_13_13_2175_0 & ~i_13_13_4513_0) | (~i_13_13_4269_0 & ~i_13_13_4324_0) | (~i_13_13_564_0 & ~i_13_13_4164_0));
endmodule



// Benchmark "kernel_13_14" written by ABC on Sun Jul 19 10:45:37 2020

module kernel_13_14 ( 
    i_13_14_51_0, i_13_14_76_0, i_13_14_112_0, i_13_14_123_0,
    i_13_14_124_0, i_13_14_169_0, i_13_14_178_0, i_13_14_186_0,
    i_13_14_187_0, i_13_14_195_0, i_13_14_283_0, i_13_14_339_0,
    i_13_14_520_0, i_13_14_535_0, i_13_14_573_0, i_13_14_574_0,
    i_13_14_618_0, i_13_14_642_0, i_13_14_643_0, i_13_14_644_0,
    i_13_14_646_0, i_13_14_690_0, i_13_14_691_0, i_13_14_697_0,
    i_13_14_717_0, i_13_14_756_0, i_13_14_816_0, i_13_14_859_0,
    i_13_14_932_0, i_13_14_1068_0, i_13_14_1069_0, i_13_14_1123_0,
    i_13_14_1138_0, i_13_14_1258_0, i_13_14_1273_0, i_13_14_1282_0,
    i_13_14_1297_0, i_13_14_1384_0, i_13_14_1407_0, i_13_14_1426_0,
    i_13_14_1461_0, i_13_14_1552_0, i_13_14_1610_0, i_13_14_1642_0,
    i_13_14_1804_0, i_13_14_1839_0, i_13_14_1851_0, i_13_14_1852_0,
    i_13_14_1861_0, i_13_14_1990_0, i_13_14_1993_0, i_13_14_2118_0,
    i_13_14_2128_0, i_13_14_2133_0, i_13_14_2136_0, i_13_14_2149_0,
    i_13_14_2212_0, i_13_14_2227_0, i_13_14_2262_0, i_13_14_2263_0,
    i_13_14_2275_0, i_13_14_2379_0, i_13_14_2410_0, i_13_14_2451_0,
    i_13_14_2536_0, i_13_14_2636_0, i_13_14_2709_0, i_13_14_2847_0,
    i_13_14_2920_0, i_13_14_2986_0, i_13_14_3030_0, i_13_14_3112_0,
    i_13_14_3166_0, i_13_14_3174_0, i_13_14_3211_0, i_13_14_3220_0,
    i_13_14_3303_0, i_13_14_3339_0, i_13_14_3424_0, i_13_14_3426_0,
    i_13_14_3427_0, i_13_14_3541_0, i_13_14_3706_0, i_13_14_3768_0,
    i_13_14_3769_0, i_13_14_3823_0, i_13_14_3918_0, i_13_14_3995_0,
    i_13_14_4011_0, i_13_14_4012_0, i_13_14_4066_0, i_13_14_4081_0,
    i_13_14_4189_0, i_13_14_4282_0, i_13_14_4314_0, i_13_14_4317_0,
    i_13_14_4318_0, i_13_14_4566_0, i_13_14_4569_0, i_13_14_4594_0,
    o_13_14_0_0  );
  input  i_13_14_51_0, i_13_14_76_0, i_13_14_112_0, i_13_14_123_0,
    i_13_14_124_0, i_13_14_169_0, i_13_14_178_0, i_13_14_186_0,
    i_13_14_187_0, i_13_14_195_0, i_13_14_283_0, i_13_14_339_0,
    i_13_14_520_0, i_13_14_535_0, i_13_14_573_0, i_13_14_574_0,
    i_13_14_618_0, i_13_14_642_0, i_13_14_643_0, i_13_14_644_0,
    i_13_14_646_0, i_13_14_690_0, i_13_14_691_0, i_13_14_697_0,
    i_13_14_717_0, i_13_14_756_0, i_13_14_816_0, i_13_14_859_0,
    i_13_14_932_0, i_13_14_1068_0, i_13_14_1069_0, i_13_14_1123_0,
    i_13_14_1138_0, i_13_14_1258_0, i_13_14_1273_0, i_13_14_1282_0,
    i_13_14_1297_0, i_13_14_1384_0, i_13_14_1407_0, i_13_14_1426_0,
    i_13_14_1461_0, i_13_14_1552_0, i_13_14_1610_0, i_13_14_1642_0,
    i_13_14_1804_0, i_13_14_1839_0, i_13_14_1851_0, i_13_14_1852_0,
    i_13_14_1861_0, i_13_14_1990_0, i_13_14_1993_0, i_13_14_2118_0,
    i_13_14_2128_0, i_13_14_2133_0, i_13_14_2136_0, i_13_14_2149_0,
    i_13_14_2212_0, i_13_14_2227_0, i_13_14_2262_0, i_13_14_2263_0,
    i_13_14_2275_0, i_13_14_2379_0, i_13_14_2410_0, i_13_14_2451_0,
    i_13_14_2536_0, i_13_14_2636_0, i_13_14_2709_0, i_13_14_2847_0,
    i_13_14_2920_0, i_13_14_2986_0, i_13_14_3030_0, i_13_14_3112_0,
    i_13_14_3166_0, i_13_14_3174_0, i_13_14_3211_0, i_13_14_3220_0,
    i_13_14_3303_0, i_13_14_3339_0, i_13_14_3424_0, i_13_14_3426_0,
    i_13_14_3427_0, i_13_14_3541_0, i_13_14_3706_0, i_13_14_3768_0,
    i_13_14_3769_0, i_13_14_3823_0, i_13_14_3918_0, i_13_14_3995_0,
    i_13_14_4011_0, i_13_14_4012_0, i_13_14_4066_0, i_13_14_4081_0,
    i_13_14_4189_0, i_13_14_4282_0, i_13_14_4314_0, i_13_14_4317_0,
    i_13_14_4318_0, i_13_14_4566_0, i_13_14_4569_0, i_13_14_4594_0;
  output o_13_14_0_0;
  assign o_13_14_0_0 = ~((i_13_14_3823_0 & ~i_13_14_4189_0) | (i_13_14_1426_0 & ~i_13_14_2536_0) | (~i_13_14_123_0 & ~i_13_14_574_0) | (~i_13_14_1804_0 & ~i_13_14_1861_0 & ~i_13_14_4569_0));
endmodule



// Benchmark "kernel_13_15" written by ABC on Sun Jul 19 10:45:38 2020

module kernel_13_15 ( 
    i_13_15_235_0, i_13_15_328_0, i_13_15_329_0, i_13_15_527_0,
    i_13_15_530_0, i_13_15_599_0, i_13_15_611_0, i_13_15_646_0,
    i_13_15_671_0, i_13_15_676_0, i_13_15_700_0, i_13_15_718_0,
    i_13_15_777_0, i_13_15_799_0, i_13_15_826_0, i_13_15_827_0,
    i_13_15_862_0, i_13_15_863_0, i_13_15_895_0, i_13_15_941_0,
    i_13_15_1024_0, i_13_15_1025_0, i_13_15_1078_0, i_13_15_1079_0,
    i_13_15_1231_0, i_13_15_1258_0, i_13_15_1259_0, i_13_15_1318_0,
    i_13_15_1411_0, i_13_15_1430_0, i_13_15_1486_0, i_13_15_1492_0,
    i_13_15_1493_0, i_13_15_1609_0, i_13_15_1636_0, i_13_15_1651_0,
    i_13_15_1691_0, i_13_15_1736_0, i_13_15_1780_0, i_13_15_1781_0,
    i_13_15_1858_0, i_13_15_1861_0, i_13_15_1862_0, i_13_15_1921_0,
    i_13_15_2021_0, i_13_15_2023_0, i_13_15_2059_0, i_13_15_2194_0,
    i_13_15_2201_0, i_13_15_2239_0, i_13_15_2266_0, i_13_15_2294_0,
    i_13_15_2404_0, i_13_15_2405_0, i_13_15_2455_0, i_13_15_2464_0,
    i_13_15_2465_0, i_13_15_2545_0, i_13_15_2546_0, i_13_15_2617_0,
    i_13_15_2618_0, i_13_15_2633_0, i_13_15_2654_0, i_13_15_2708_0,
    i_13_15_2876_0, i_13_15_3017_0, i_13_15_3172_0, i_13_15_3173_0,
    i_13_15_3175_0, i_13_15_3176_0, i_13_15_3233_0, i_13_15_3367_0,
    i_13_15_3373_0, i_13_15_3464_0, i_13_15_3482_0, i_13_15_3536_0,
    i_13_15_3542_0, i_13_15_3544_0, i_13_15_3563_0, i_13_15_3622_0,
    i_13_15_3788_0, i_13_15_3806_0, i_13_15_3847_0, i_13_15_3859_0,
    i_13_15_3877_0, i_13_15_3890_0, i_13_15_3896_0, i_13_15_3914_0,
    i_13_15_4013_0, i_13_15_4019_0, i_13_15_4100_0, i_13_15_4118_0,
    i_13_15_4126_0, i_13_15_4162_0, i_13_15_4192_0, i_13_15_4262_0,
    i_13_15_4280_0, i_13_15_4373_0, i_13_15_4396_0, i_13_15_4444_0,
    o_13_15_0_0  );
  input  i_13_15_235_0, i_13_15_328_0, i_13_15_329_0, i_13_15_527_0,
    i_13_15_530_0, i_13_15_599_0, i_13_15_611_0, i_13_15_646_0,
    i_13_15_671_0, i_13_15_676_0, i_13_15_700_0, i_13_15_718_0,
    i_13_15_777_0, i_13_15_799_0, i_13_15_826_0, i_13_15_827_0,
    i_13_15_862_0, i_13_15_863_0, i_13_15_895_0, i_13_15_941_0,
    i_13_15_1024_0, i_13_15_1025_0, i_13_15_1078_0, i_13_15_1079_0,
    i_13_15_1231_0, i_13_15_1258_0, i_13_15_1259_0, i_13_15_1318_0,
    i_13_15_1411_0, i_13_15_1430_0, i_13_15_1486_0, i_13_15_1492_0,
    i_13_15_1493_0, i_13_15_1609_0, i_13_15_1636_0, i_13_15_1651_0,
    i_13_15_1691_0, i_13_15_1736_0, i_13_15_1780_0, i_13_15_1781_0,
    i_13_15_1858_0, i_13_15_1861_0, i_13_15_1862_0, i_13_15_1921_0,
    i_13_15_2021_0, i_13_15_2023_0, i_13_15_2059_0, i_13_15_2194_0,
    i_13_15_2201_0, i_13_15_2239_0, i_13_15_2266_0, i_13_15_2294_0,
    i_13_15_2404_0, i_13_15_2405_0, i_13_15_2455_0, i_13_15_2464_0,
    i_13_15_2465_0, i_13_15_2545_0, i_13_15_2546_0, i_13_15_2617_0,
    i_13_15_2618_0, i_13_15_2633_0, i_13_15_2654_0, i_13_15_2708_0,
    i_13_15_2876_0, i_13_15_3017_0, i_13_15_3172_0, i_13_15_3173_0,
    i_13_15_3175_0, i_13_15_3176_0, i_13_15_3233_0, i_13_15_3367_0,
    i_13_15_3373_0, i_13_15_3464_0, i_13_15_3482_0, i_13_15_3536_0,
    i_13_15_3542_0, i_13_15_3544_0, i_13_15_3563_0, i_13_15_3622_0,
    i_13_15_3788_0, i_13_15_3806_0, i_13_15_3847_0, i_13_15_3859_0,
    i_13_15_3877_0, i_13_15_3890_0, i_13_15_3896_0, i_13_15_3914_0,
    i_13_15_4013_0, i_13_15_4019_0, i_13_15_4100_0, i_13_15_4118_0,
    i_13_15_4126_0, i_13_15_4162_0, i_13_15_4192_0, i_13_15_4262_0,
    i_13_15_4280_0, i_13_15_4373_0, i_13_15_4396_0, i_13_15_4444_0;
  output o_13_15_0_0;
  assign o_13_15_0_0 = ~((~i_13_15_329_0 & ~i_13_15_3536_0) | (~i_13_15_1079_0 & ~i_13_15_3176_0) | (~i_13_15_328_0 & ~i_13_15_863_0 & ~i_13_15_3464_0));
endmodule



// Benchmark "kernel_13_16" written by ABC on Sun Jul 19 10:45:39 2020

module kernel_13_16 ( 
    i_13_16_35_0, i_13_16_106_0, i_13_16_178_0, i_13_16_187_0,
    i_13_16_284_0, i_13_16_322_0, i_13_16_325_0, i_13_16_326_0,
    i_13_16_355_0, i_13_16_454_0, i_13_16_480_0, i_13_16_496_0,
    i_13_16_521_0, i_13_16_562_0, i_13_16_574_0, i_13_16_575_0,
    i_13_16_599_0, i_13_16_644_0, i_13_16_646_0, i_13_16_647_0,
    i_13_16_685_0, i_13_16_718_0, i_13_16_849_0, i_13_16_850_0,
    i_13_16_851_0, i_13_16_914_0, i_13_16_1210_0, i_13_16_1229_0,
    i_13_16_1255_0, i_13_16_1282_0, i_13_16_1345_0, i_13_16_1410_0,
    i_13_16_1444_0, i_13_16_1471_0, i_13_16_1552_0, i_13_16_1646_0,
    i_13_16_1678_0, i_13_16_1683_0, i_13_16_1691_0, i_13_16_1740_0,
    i_13_16_1750_0, i_13_16_1753_0, i_13_16_1788_0, i_13_16_1807_0,
    i_13_16_1857_0, i_13_16_1858_0, i_13_16_1859_0, i_13_16_1861_0,
    i_13_16_1862_0, i_13_16_1958_0, i_13_16_1993_0, i_13_16_2050_0,
    i_13_16_2103_0, i_13_16_2141_0, i_13_16_2159_0, i_13_16_2182_0,
    i_13_16_2281_0, i_13_16_2302_0, i_13_16_2311_0, i_13_16_2459_0,
    i_13_16_2463_0, i_13_16_2551_0, i_13_16_2588_0, i_13_16_2653_0,
    i_13_16_2654_0, i_13_16_2722_0, i_13_16_2752_0, i_13_16_2790_0,
    i_13_16_3064_0, i_13_16_3170_0, i_13_16_3172_0, i_13_16_3175_0,
    i_13_16_3209_0, i_13_16_3235_0, i_13_16_3271_0, i_13_16_3272_0,
    i_13_16_3274_0, i_13_16_3275_0, i_13_16_3309_0, i_13_16_3401_0,
    i_13_16_3426_0, i_13_16_3433_0, i_13_16_3562_0, i_13_16_3563_0,
    i_13_16_3847_0, i_13_16_3856_0, i_13_16_3892_0, i_13_16_3911_0,
    i_13_16_3912_0, i_13_16_3913_0, i_13_16_3914_0, i_13_16_4016_0,
    i_13_16_4047_0, i_13_16_4098_0, i_13_16_4149_0, i_13_16_4262_0,
    i_13_16_4378_0, i_13_16_4379_0, i_13_16_4382_0, i_13_16_4581_0,
    o_13_16_0_0  );
  input  i_13_16_35_0, i_13_16_106_0, i_13_16_178_0, i_13_16_187_0,
    i_13_16_284_0, i_13_16_322_0, i_13_16_325_0, i_13_16_326_0,
    i_13_16_355_0, i_13_16_454_0, i_13_16_480_0, i_13_16_496_0,
    i_13_16_521_0, i_13_16_562_0, i_13_16_574_0, i_13_16_575_0,
    i_13_16_599_0, i_13_16_644_0, i_13_16_646_0, i_13_16_647_0,
    i_13_16_685_0, i_13_16_718_0, i_13_16_849_0, i_13_16_850_0,
    i_13_16_851_0, i_13_16_914_0, i_13_16_1210_0, i_13_16_1229_0,
    i_13_16_1255_0, i_13_16_1282_0, i_13_16_1345_0, i_13_16_1410_0,
    i_13_16_1444_0, i_13_16_1471_0, i_13_16_1552_0, i_13_16_1646_0,
    i_13_16_1678_0, i_13_16_1683_0, i_13_16_1691_0, i_13_16_1740_0,
    i_13_16_1750_0, i_13_16_1753_0, i_13_16_1788_0, i_13_16_1807_0,
    i_13_16_1857_0, i_13_16_1858_0, i_13_16_1859_0, i_13_16_1861_0,
    i_13_16_1862_0, i_13_16_1958_0, i_13_16_1993_0, i_13_16_2050_0,
    i_13_16_2103_0, i_13_16_2141_0, i_13_16_2159_0, i_13_16_2182_0,
    i_13_16_2281_0, i_13_16_2302_0, i_13_16_2311_0, i_13_16_2459_0,
    i_13_16_2463_0, i_13_16_2551_0, i_13_16_2588_0, i_13_16_2653_0,
    i_13_16_2654_0, i_13_16_2722_0, i_13_16_2752_0, i_13_16_2790_0,
    i_13_16_3064_0, i_13_16_3170_0, i_13_16_3172_0, i_13_16_3175_0,
    i_13_16_3209_0, i_13_16_3235_0, i_13_16_3271_0, i_13_16_3272_0,
    i_13_16_3274_0, i_13_16_3275_0, i_13_16_3309_0, i_13_16_3401_0,
    i_13_16_3426_0, i_13_16_3433_0, i_13_16_3562_0, i_13_16_3563_0,
    i_13_16_3847_0, i_13_16_3856_0, i_13_16_3892_0, i_13_16_3911_0,
    i_13_16_3912_0, i_13_16_3913_0, i_13_16_3914_0, i_13_16_4016_0,
    i_13_16_4047_0, i_13_16_4098_0, i_13_16_4149_0, i_13_16_4262_0,
    i_13_16_4378_0, i_13_16_4379_0, i_13_16_4382_0, i_13_16_4581_0;
  output o_13_16_0_0;
  assign o_13_16_0_0 = ~((~i_13_16_1858_0 & ((~i_13_16_325_0 & ~i_13_16_521_0 & ~i_13_16_1857_0 & ~i_13_16_1859_0 & ~i_13_16_2141_0 & ~i_13_16_3912_0) | (i_13_16_2182_0 & ~i_13_16_3401_0 & ~i_13_16_3426_0 & ~i_13_16_4382_0))) | (~i_13_16_178_0 & ~i_13_16_1750_0 & ~i_13_16_1859_0 & ~i_13_16_2653_0) | (~i_13_16_187_0 & ~i_13_16_322_0 & ~i_13_16_1862_0 & ~i_13_16_3209_0 & ~i_13_16_3856_0) | (i_13_16_1993_0 & ~i_13_16_3911_0 & ~i_13_16_3913_0) | (~i_13_16_1753_0 & ~i_13_16_2463_0 & i_13_16_3892_0 & ~i_13_16_4262_0) | (~i_13_16_1861_0 & ~i_13_16_3401_0 & ~i_13_16_3892_0 & ~i_13_16_4378_0 & ~i_13_16_4382_0));
endmodule



// Benchmark "kernel_13_17" written by ABC on Sun Jul 19 10:45:40 2020

module kernel_13_17 ( 
    i_13_17_27_0, i_13_17_28_0, i_13_17_31_0, i_13_17_63_0, i_13_17_67_0,
    i_13_17_90_0, i_13_17_100_0, i_13_17_111_0, i_13_17_130_0,
    i_13_17_174_0, i_13_17_196_0, i_13_17_225_0, i_13_17_226_0,
    i_13_17_255_0, i_13_17_306_0, i_13_17_307_0, i_13_17_372_0,
    i_13_17_462_0, i_13_17_612_0, i_13_17_616_0, i_13_17_666_0,
    i_13_17_667_0, i_13_17_670_0, i_13_17_729_0, i_13_17_796_0,
    i_13_17_828_0, i_13_17_853_0, i_13_17_855_0, i_13_17_858_0,
    i_13_17_1075_0, i_13_17_1120_0, i_13_17_1128_0, i_13_17_1200_0,
    i_13_17_1215_0, i_13_17_1225_0, i_13_17_1231_0, i_13_17_1306_0,
    i_13_17_1321_0, i_13_17_1344_0, i_13_17_1398_0, i_13_17_1440_0,
    i_13_17_1480_0, i_13_17_1620_0, i_13_17_1689_0, i_13_17_1696_0,
    i_13_17_1846_0, i_13_17_1927_0, i_13_17_1998_0, i_13_17_1999_0,
    i_13_17_2100_0, i_13_17_2200_0, i_13_17_2205_0, i_13_17_2206_0,
    i_13_17_2422_0, i_13_17_2430_0, i_13_17_2431_0, i_13_17_2538_0,
    i_13_17_2718_0, i_13_17_2719_0, i_13_17_2739_0, i_13_17_2740_0,
    i_13_17_2766_0, i_13_17_2781_0, i_13_17_2796_0, i_13_17_2797_0,
    i_13_17_2880_0, i_13_17_3066_0, i_13_17_3126_0, i_13_17_3133_0,
    i_13_17_3231_0, i_13_17_3240_0, i_13_17_3241_0, i_13_17_3309_0,
    i_13_17_3388_0, i_13_17_3414_0, i_13_17_3420_0, i_13_17_3460_0,
    i_13_17_3619_0, i_13_17_3636_0, i_13_17_3637_0, i_13_17_3682_0,
    i_13_17_3699_0, i_13_17_3717_0, i_13_17_3760_0, i_13_17_3762_0,
    i_13_17_3795_0, i_13_17_3843_0, i_13_17_3844_0, i_13_17_3862_0,
    i_13_17_3870_0, i_13_17_3906_0, i_13_17_3934_0, i_13_17_4050_0,
    i_13_17_4212_0, i_13_17_4326_0, i_13_17_4347_0, i_13_17_4350_0,
    i_13_17_4360_0, i_13_17_4387_0, i_13_17_4470_0,
    o_13_17_0_0  );
  input  i_13_17_27_0, i_13_17_28_0, i_13_17_31_0, i_13_17_63_0,
    i_13_17_67_0, i_13_17_90_0, i_13_17_100_0, i_13_17_111_0,
    i_13_17_130_0, i_13_17_174_0, i_13_17_196_0, i_13_17_225_0,
    i_13_17_226_0, i_13_17_255_0, i_13_17_306_0, i_13_17_307_0,
    i_13_17_372_0, i_13_17_462_0, i_13_17_612_0, i_13_17_616_0,
    i_13_17_666_0, i_13_17_667_0, i_13_17_670_0, i_13_17_729_0,
    i_13_17_796_0, i_13_17_828_0, i_13_17_853_0, i_13_17_855_0,
    i_13_17_858_0, i_13_17_1075_0, i_13_17_1120_0, i_13_17_1128_0,
    i_13_17_1200_0, i_13_17_1215_0, i_13_17_1225_0, i_13_17_1231_0,
    i_13_17_1306_0, i_13_17_1321_0, i_13_17_1344_0, i_13_17_1398_0,
    i_13_17_1440_0, i_13_17_1480_0, i_13_17_1620_0, i_13_17_1689_0,
    i_13_17_1696_0, i_13_17_1846_0, i_13_17_1927_0, i_13_17_1998_0,
    i_13_17_1999_0, i_13_17_2100_0, i_13_17_2200_0, i_13_17_2205_0,
    i_13_17_2206_0, i_13_17_2422_0, i_13_17_2430_0, i_13_17_2431_0,
    i_13_17_2538_0, i_13_17_2718_0, i_13_17_2719_0, i_13_17_2739_0,
    i_13_17_2740_0, i_13_17_2766_0, i_13_17_2781_0, i_13_17_2796_0,
    i_13_17_2797_0, i_13_17_2880_0, i_13_17_3066_0, i_13_17_3126_0,
    i_13_17_3133_0, i_13_17_3231_0, i_13_17_3240_0, i_13_17_3241_0,
    i_13_17_3309_0, i_13_17_3388_0, i_13_17_3414_0, i_13_17_3420_0,
    i_13_17_3460_0, i_13_17_3619_0, i_13_17_3636_0, i_13_17_3637_0,
    i_13_17_3682_0, i_13_17_3699_0, i_13_17_3717_0, i_13_17_3760_0,
    i_13_17_3762_0, i_13_17_3795_0, i_13_17_3843_0, i_13_17_3844_0,
    i_13_17_3862_0, i_13_17_3870_0, i_13_17_3906_0, i_13_17_3934_0,
    i_13_17_4050_0, i_13_17_4212_0, i_13_17_4326_0, i_13_17_4347_0,
    i_13_17_4350_0, i_13_17_4360_0, i_13_17_4387_0, i_13_17_4470_0;
  output o_13_17_0_0;
  assign o_13_17_0_0 = ~((~i_13_17_2431_0 & ~i_13_17_3844_0 & ~i_13_17_4050_0) | (~i_13_17_63_0 & ~i_13_17_90_0 & ~i_13_17_3240_0));
endmodule



// Benchmark "kernel_13_18" written by ABC on Sun Jul 19 10:45:41 2020

module kernel_13_18 ( 
    i_13_18_38_0, i_13_18_41_0, i_13_18_91_0, i_13_18_109_0, i_13_18_210_0,
    i_13_18_227_0, i_13_18_279_0, i_13_18_282_0, i_13_18_405_0,
    i_13_18_459_0, i_13_18_643_0, i_13_18_651_0, i_13_18_686_0,
    i_13_18_734_0, i_13_18_792_0, i_13_18_793_0, i_13_18_847_0,
    i_13_18_855_0, i_13_18_902_0, i_13_18_955_0, i_13_18_1017_0,
    i_13_18_1018_0, i_13_18_1020_0, i_13_18_1021_0, i_13_18_1120_0,
    i_13_18_1200_0, i_13_18_1270_0, i_13_18_1273_0, i_13_18_1308_0,
    i_13_18_1440_0, i_13_18_1459_0, i_13_18_1485_0, i_13_18_1486_0,
    i_13_18_1535_0, i_13_18_1548_0, i_13_18_1603_0, i_13_18_1629_0,
    i_13_18_1630_0, i_13_18_1639_0, i_13_18_1792_0, i_13_18_1813_0,
    i_13_18_1828_0, i_13_18_1832_0, i_13_18_1854_0, i_13_18_1998_0,
    i_13_18_2197_0, i_13_18_2205_0, i_13_18_2421_0, i_13_18_2435_0,
    i_13_18_2457_0, i_13_18_2458_0, i_13_18_2461_0, i_13_18_2467_0,
    i_13_18_2529_0, i_13_18_2538_0, i_13_18_2539_0, i_13_18_2542_0,
    i_13_18_2551_0, i_13_18_2712_0, i_13_18_2848_0, i_13_18_2916_0,
    i_13_18_2917_0, i_13_18_2918_0, i_13_18_3126_0, i_13_18_3160_0,
    i_13_18_3169_0, i_13_18_3268_0, i_13_18_3404_0, i_13_18_3407_0,
    i_13_18_3450_0, i_13_18_3460_0, i_13_18_3537_0, i_13_18_3551_0,
    i_13_18_3577_0, i_13_18_3663_0, i_13_18_3684_0, i_13_18_3726_0,
    i_13_18_3728_0, i_13_18_3754_0, i_13_18_3843_0, i_13_18_3853_0,
    i_13_18_3907_0, i_13_18_3910_0, i_13_18_3928_0, i_13_18_3987_0,
    i_13_18_4015_0, i_13_18_4033_0, i_13_18_4123_0, i_13_18_4186_0,
    i_13_18_4252_0, i_13_18_4322_0, i_13_18_4338_0, i_13_18_4341_0,
    i_13_18_4519_0, i_13_18_4522_0, i_13_18_4534_0, i_13_18_4558_0,
    i_13_18_4559_0, i_13_18_4591_0, i_13_18_4600_0,
    o_13_18_0_0  );
  input  i_13_18_38_0, i_13_18_41_0, i_13_18_91_0, i_13_18_109_0,
    i_13_18_210_0, i_13_18_227_0, i_13_18_279_0, i_13_18_282_0,
    i_13_18_405_0, i_13_18_459_0, i_13_18_643_0, i_13_18_651_0,
    i_13_18_686_0, i_13_18_734_0, i_13_18_792_0, i_13_18_793_0,
    i_13_18_847_0, i_13_18_855_0, i_13_18_902_0, i_13_18_955_0,
    i_13_18_1017_0, i_13_18_1018_0, i_13_18_1020_0, i_13_18_1021_0,
    i_13_18_1120_0, i_13_18_1200_0, i_13_18_1270_0, i_13_18_1273_0,
    i_13_18_1308_0, i_13_18_1440_0, i_13_18_1459_0, i_13_18_1485_0,
    i_13_18_1486_0, i_13_18_1535_0, i_13_18_1548_0, i_13_18_1603_0,
    i_13_18_1629_0, i_13_18_1630_0, i_13_18_1639_0, i_13_18_1792_0,
    i_13_18_1813_0, i_13_18_1828_0, i_13_18_1832_0, i_13_18_1854_0,
    i_13_18_1998_0, i_13_18_2197_0, i_13_18_2205_0, i_13_18_2421_0,
    i_13_18_2435_0, i_13_18_2457_0, i_13_18_2458_0, i_13_18_2461_0,
    i_13_18_2467_0, i_13_18_2529_0, i_13_18_2538_0, i_13_18_2539_0,
    i_13_18_2542_0, i_13_18_2551_0, i_13_18_2712_0, i_13_18_2848_0,
    i_13_18_2916_0, i_13_18_2917_0, i_13_18_2918_0, i_13_18_3126_0,
    i_13_18_3160_0, i_13_18_3169_0, i_13_18_3268_0, i_13_18_3404_0,
    i_13_18_3407_0, i_13_18_3450_0, i_13_18_3460_0, i_13_18_3537_0,
    i_13_18_3551_0, i_13_18_3577_0, i_13_18_3663_0, i_13_18_3684_0,
    i_13_18_3726_0, i_13_18_3728_0, i_13_18_3754_0, i_13_18_3843_0,
    i_13_18_3853_0, i_13_18_3907_0, i_13_18_3910_0, i_13_18_3928_0,
    i_13_18_3987_0, i_13_18_4015_0, i_13_18_4033_0, i_13_18_4123_0,
    i_13_18_4186_0, i_13_18_4252_0, i_13_18_4322_0, i_13_18_4338_0,
    i_13_18_4341_0, i_13_18_4519_0, i_13_18_4522_0, i_13_18_4534_0,
    i_13_18_4558_0, i_13_18_4559_0, i_13_18_4591_0, i_13_18_4600_0;
  output o_13_18_0_0;
  assign o_13_18_0_0 = ~(~i_13_18_2458_0 | (i_13_18_1270_0 & ~i_13_18_3726_0) | (~i_13_18_2529_0 & ~i_13_18_2916_0));
endmodule



// Benchmark "kernel_13_19" written by ABC on Sun Jul 19 10:45:41 2020

module kernel_13_19 ( 
    i_13_19_41_0, i_13_19_59_0, i_13_19_76_0, i_13_19_100_0, i_13_19_106_0,
    i_13_19_136_0, i_13_19_190_0, i_13_19_193_0, i_13_19_218_0,
    i_13_19_256_0, i_13_19_328_0, i_13_19_376_0, i_13_19_416_0,
    i_13_19_428_0, i_13_19_533_0, i_13_19_577_0, i_13_19_599_0,
    i_13_19_614_0, i_13_19_622_0, i_13_19_626_0, i_13_19_628_0,
    i_13_19_629_0, i_13_19_644_0, i_13_19_685_0, i_13_19_715_0,
    i_13_19_725_0, i_13_19_778_0, i_13_19_854_0, i_13_19_884_0,
    i_13_19_892_0, i_13_19_895_0, i_13_19_911_0, i_13_19_980_0,
    i_13_19_1022_0, i_13_19_1096_0, i_13_19_1124_0, i_13_19_1249_0,
    i_13_19_1256_0, i_13_19_1280_0, i_13_19_1391_0, i_13_19_1445_0,
    i_13_19_1462_0, i_13_19_1471_0, i_13_19_1483_0, i_13_19_1484_0,
    i_13_19_1541_0, i_13_19_1597_0, i_13_19_1643_0, i_13_19_1676_0,
    i_13_19_1678_0, i_13_19_1688_0, i_13_19_1691_0, i_13_19_1748_0,
    i_13_19_1757_0, i_13_19_1849_0, i_13_19_1855_0, i_13_19_1856_0,
    i_13_19_1858_0, i_13_19_1862_0, i_13_19_1883_0, i_13_19_2053_0,
    i_13_19_2209_0, i_13_19_2245_0, i_13_19_2434_0, i_13_19_2506_0,
    i_13_19_2507_0, i_13_19_2630_0, i_13_19_2717_0, i_13_19_2818_0,
    i_13_19_2845_0, i_13_19_2848_0, i_13_19_2849_0, i_13_19_2851_0,
    i_13_19_2857_0, i_13_19_2875_0, i_13_19_2878_0, i_13_19_2909_0,
    i_13_19_2911_0, i_13_19_2921_0, i_13_19_3064_0, i_13_19_3065_0,
    i_13_19_3118_0, i_13_19_3170_0, i_13_19_3265_0, i_13_19_3305_0,
    i_13_19_3433_0, i_13_19_3436_0, i_13_19_3766_0, i_13_19_3791_0,
    i_13_19_3818_0, i_13_19_3832_0, i_13_19_3869_0, i_13_19_3884_0,
    i_13_19_4297_0, i_13_19_4328_0, i_13_19_4379_0, i_13_19_4421_0,
    i_13_19_4441_0, i_13_19_4508_0, i_13_19_4607_0,
    o_13_19_0_0  );
  input  i_13_19_41_0, i_13_19_59_0, i_13_19_76_0, i_13_19_100_0,
    i_13_19_106_0, i_13_19_136_0, i_13_19_190_0, i_13_19_193_0,
    i_13_19_218_0, i_13_19_256_0, i_13_19_328_0, i_13_19_376_0,
    i_13_19_416_0, i_13_19_428_0, i_13_19_533_0, i_13_19_577_0,
    i_13_19_599_0, i_13_19_614_0, i_13_19_622_0, i_13_19_626_0,
    i_13_19_628_0, i_13_19_629_0, i_13_19_644_0, i_13_19_685_0,
    i_13_19_715_0, i_13_19_725_0, i_13_19_778_0, i_13_19_854_0,
    i_13_19_884_0, i_13_19_892_0, i_13_19_895_0, i_13_19_911_0,
    i_13_19_980_0, i_13_19_1022_0, i_13_19_1096_0, i_13_19_1124_0,
    i_13_19_1249_0, i_13_19_1256_0, i_13_19_1280_0, i_13_19_1391_0,
    i_13_19_1445_0, i_13_19_1462_0, i_13_19_1471_0, i_13_19_1483_0,
    i_13_19_1484_0, i_13_19_1541_0, i_13_19_1597_0, i_13_19_1643_0,
    i_13_19_1676_0, i_13_19_1678_0, i_13_19_1688_0, i_13_19_1691_0,
    i_13_19_1748_0, i_13_19_1757_0, i_13_19_1849_0, i_13_19_1855_0,
    i_13_19_1856_0, i_13_19_1858_0, i_13_19_1862_0, i_13_19_1883_0,
    i_13_19_2053_0, i_13_19_2209_0, i_13_19_2245_0, i_13_19_2434_0,
    i_13_19_2506_0, i_13_19_2507_0, i_13_19_2630_0, i_13_19_2717_0,
    i_13_19_2818_0, i_13_19_2845_0, i_13_19_2848_0, i_13_19_2849_0,
    i_13_19_2851_0, i_13_19_2857_0, i_13_19_2875_0, i_13_19_2878_0,
    i_13_19_2909_0, i_13_19_2911_0, i_13_19_2921_0, i_13_19_3064_0,
    i_13_19_3065_0, i_13_19_3118_0, i_13_19_3170_0, i_13_19_3265_0,
    i_13_19_3305_0, i_13_19_3433_0, i_13_19_3436_0, i_13_19_3766_0,
    i_13_19_3791_0, i_13_19_3818_0, i_13_19_3832_0, i_13_19_3869_0,
    i_13_19_3884_0, i_13_19_4297_0, i_13_19_4328_0, i_13_19_4379_0,
    i_13_19_4421_0, i_13_19_4441_0, i_13_19_4508_0, i_13_19_4607_0;
  output o_13_19_0_0;
  assign o_13_19_0_0 = ~((~i_13_19_59_0 & (~i_13_19_2245_0 | (i_13_19_1597_0 & ~i_13_19_1643_0 & ~i_13_19_2845_0))) | (~i_13_19_895_0 & ((i_13_19_1597_0 & i_13_19_2845_0) | (~i_13_19_328_0 & ~i_13_19_1484_0 & ~i_13_19_3170_0 & ~i_13_19_4379_0))) | (~i_13_19_2875_0 & (i_13_19_2434_0 | (~i_13_19_1124_0 & ~i_13_19_1856_0))) | (i_13_19_1471_0 & ~i_13_19_1862_0 & ~i_13_19_2851_0 & ~i_13_19_3170_0) | (~i_13_19_2848_0 & ~i_13_19_3869_0 & ~i_13_19_4379_0));
endmodule



// Benchmark "kernel_13_20" written by ABC on Sun Jul 19 10:45:42 2020

module kernel_13_20 ( 
    i_13_20_45_0, i_13_20_75_0, i_13_20_117_0, i_13_20_139_0,
    i_13_20_162_0, i_13_20_167_0, i_13_20_178_0, i_13_20_184_0,
    i_13_20_211_0, i_13_20_336_0, i_13_20_419_0, i_13_20_517_0,
    i_13_20_562_0, i_13_20_571_0, i_13_20_574_0, i_13_20_607_0,
    i_13_20_746_0, i_13_20_814_0, i_13_20_815_0, i_13_20_875_0,
    i_13_20_910_0, i_13_20_955_0, i_13_20_1080_0, i_13_20_1084_0,
    i_13_20_1132_0, i_13_20_1192_0, i_13_20_1219_0, i_13_20_1220_0,
    i_13_20_1345_0, i_13_20_1404_0, i_13_20_1409_0, i_13_20_1465_0,
    i_13_20_1496_0, i_13_20_1525_0, i_13_20_1526_0, i_13_20_1552_0,
    i_13_20_1555_0, i_13_20_1642_0, i_13_20_1699_0, i_13_20_1782_0,
    i_13_20_1800_0, i_13_20_1857_0, i_13_20_1858_0, i_13_20_1886_0,
    i_13_20_1960_0, i_13_20_1961_0, i_13_20_2201_0, i_13_20_2209_0,
    i_13_20_2223_0, i_13_20_2239_0, i_13_20_2240_0, i_13_20_2259_0,
    i_13_20_2277_0, i_13_20_2296_0, i_13_20_2381_0, i_13_20_2407_0,
    i_13_20_2428_0, i_13_20_2508_0, i_13_20_2552_0, i_13_20_2712_0,
    i_13_20_2848_0, i_13_20_2857_0, i_13_20_2898_0, i_13_20_2938_0,
    i_13_20_3100_0, i_13_20_3101_0, i_13_20_3146_0, i_13_20_3169_0,
    i_13_20_3208_0, i_13_20_3244_0, i_13_20_3347_0, i_13_20_3419_0,
    i_13_20_3473_0, i_13_20_3490_0, i_13_20_3505_0, i_13_20_3542_0,
    i_13_20_3555_0, i_13_20_3592_0, i_13_20_3618_0, i_13_20_3641_0,
    i_13_20_3670_0, i_13_20_3739_0, i_13_20_3804_0, i_13_20_3859_0,
    i_13_20_3860_0, i_13_20_3899_0, i_13_20_3909_0, i_13_20_3911_0,
    i_13_20_3913_0, i_13_20_4012_0, i_13_20_4081_0, i_13_20_4096_0,
    i_13_20_4097_0, i_13_20_4147_0, i_13_20_4189_0, i_13_20_4237_0,
    i_13_20_4293_0, i_13_20_4315_0, i_13_20_4322_0, i_13_20_4433_0,
    o_13_20_0_0  );
  input  i_13_20_45_0, i_13_20_75_0, i_13_20_117_0, i_13_20_139_0,
    i_13_20_162_0, i_13_20_167_0, i_13_20_178_0, i_13_20_184_0,
    i_13_20_211_0, i_13_20_336_0, i_13_20_419_0, i_13_20_517_0,
    i_13_20_562_0, i_13_20_571_0, i_13_20_574_0, i_13_20_607_0,
    i_13_20_746_0, i_13_20_814_0, i_13_20_815_0, i_13_20_875_0,
    i_13_20_910_0, i_13_20_955_0, i_13_20_1080_0, i_13_20_1084_0,
    i_13_20_1132_0, i_13_20_1192_0, i_13_20_1219_0, i_13_20_1220_0,
    i_13_20_1345_0, i_13_20_1404_0, i_13_20_1409_0, i_13_20_1465_0,
    i_13_20_1496_0, i_13_20_1525_0, i_13_20_1526_0, i_13_20_1552_0,
    i_13_20_1555_0, i_13_20_1642_0, i_13_20_1699_0, i_13_20_1782_0,
    i_13_20_1800_0, i_13_20_1857_0, i_13_20_1858_0, i_13_20_1886_0,
    i_13_20_1960_0, i_13_20_1961_0, i_13_20_2201_0, i_13_20_2209_0,
    i_13_20_2223_0, i_13_20_2239_0, i_13_20_2240_0, i_13_20_2259_0,
    i_13_20_2277_0, i_13_20_2296_0, i_13_20_2381_0, i_13_20_2407_0,
    i_13_20_2428_0, i_13_20_2508_0, i_13_20_2552_0, i_13_20_2712_0,
    i_13_20_2848_0, i_13_20_2857_0, i_13_20_2898_0, i_13_20_2938_0,
    i_13_20_3100_0, i_13_20_3101_0, i_13_20_3146_0, i_13_20_3169_0,
    i_13_20_3208_0, i_13_20_3244_0, i_13_20_3347_0, i_13_20_3419_0,
    i_13_20_3473_0, i_13_20_3490_0, i_13_20_3505_0, i_13_20_3542_0,
    i_13_20_3555_0, i_13_20_3592_0, i_13_20_3618_0, i_13_20_3641_0,
    i_13_20_3670_0, i_13_20_3739_0, i_13_20_3804_0, i_13_20_3859_0,
    i_13_20_3860_0, i_13_20_3899_0, i_13_20_3909_0, i_13_20_3911_0,
    i_13_20_3913_0, i_13_20_4012_0, i_13_20_4081_0, i_13_20_4096_0,
    i_13_20_4097_0, i_13_20_4147_0, i_13_20_4189_0, i_13_20_4237_0,
    i_13_20_4293_0, i_13_20_4315_0, i_13_20_4322_0, i_13_20_4433_0;
  output o_13_20_0_0;
  assign o_13_20_0_0 = ~((~i_13_20_2239_0 & ((~i_13_20_1409_0 & ~i_13_20_1526_0 & ~i_13_20_1857_0) | (i_13_20_1858_0 & ~i_13_20_3146_0 & ~i_13_20_3860_0 & ~i_13_20_4315_0))) | (~i_13_20_2223_0 & ((~i_13_20_2209_0 & i_13_20_2898_0) | i_13_20_3592_0 | (~i_13_20_419_0 & ~i_13_20_1404_0 & ~i_13_20_1960_0 & ~i_13_20_4012_0))) | (~i_13_20_1555_0 & ~i_13_20_1858_0 & ~i_13_20_3859_0) | (~i_13_20_336_0 & ~i_13_20_1642_0 & i_13_20_4081_0) | (i_13_20_3505_0 & ~i_13_20_3911_0 & ~i_13_20_3913_0 & ~i_13_20_4081_0));
endmodule



// Benchmark "kernel_13_21" written by ABC on Sun Jul 19 10:45:43 2020

module kernel_13_21 ( 
    i_13_21_69_0, i_13_21_70_0, i_13_21_78_0, i_13_21_124_0, i_13_21_286_0,
    i_13_21_313_0, i_13_21_375_0, i_13_21_385_0, i_13_21_411_0,
    i_13_21_448_0, i_13_21_520_0, i_13_21_535_0, i_13_21_588_0,
    i_13_21_646_0, i_13_21_672_0, i_13_21_673_0, i_13_21_682_0,
    i_13_21_699_0, i_13_21_700_0, i_13_21_843_0, i_13_21_844_0,
    i_13_21_886_0, i_13_21_934_0, i_13_21_980_0, i_13_21_1102_0,
    i_13_21_1104_0, i_13_21_1105_0, i_13_21_1122_0, i_13_21_1222_0,
    i_13_21_1275_0, i_13_21_1276_0, i_13_21_1302_0, i_13_21_1311_0,
    i_13_21_1312_0, i_13_21_1402_0, i_13_21_1403_0, i_13_21_1428_0,
    i_13_21_1437_0, i_13_21_1438_0, i_13_21_1510_0, i_13_21_1600_0,
    i_13_21_1663_0, i_13_21_1665_0, i_13_21_1723_0, i_13_21_1725_0,
    i_13_21_1735_0, i_13_21_1777_0, i_13_21_1779_0, i_13_21_1798_0,
    i_13_21_1887_0, i_13_21_1888_0, i_13_21_1933_0, i_13_21_1935_0,
    i_13_21_1936_0, i_13_21_1947_0, i_13_21_1948_0, i_13_21_1995_0,
    i_13_21_1996_0, i_13_21_2004_0, i_13_21_2014_0, i_13_21_2029_0,
    i_13_21_2139_0, i_13_21_2140_0, i_13_21_2379_0, i_13_21_2383_0,
    i_13_21_2480_0, i_13_21_2551_0, i_13_21_2569_0, i_13_21_2599_0,
    i_13_21_2616_0, i_13_21_2650_0, i_13_21_2679_0, i_13_21_2697_0,
    i_13_21_2698_0, i_13_21_2712_0, i_13_21_2770_0, i_13_21_2824_0,
    i_13_21_2851_0, i_13_21_2901_0, i_13_21_2923_0, i_13_21_2958_0,
    i_13_21_3031_0, i_13_21_3208_0, i_13_21_3595_0, i_13_21_3596_0,
    i_13_21_3613_0, i_13_21_3742_0, i_13_21_3787_0, i_13_21_3930_0,
    i_13_21_3931_0, i_13_21_4063_0, i_13_21_4260_0, i_13_21_4302_0,
    i_13_21_4308_0, i_13_21_4309_0, i_13_21_4450_0, i_13_21_4596_0,
    i_13_21_4597_0, i_13_21_4606_0, i_13_21_4607_0,
    o_13_21_0_0  );
  input  i_13_21_69_0, i_13_21_70_0, i_13_21_78_0, i_13_21_124_0,
    i_13_21_286_0, i_13_21_313_0, i_13_21_375_0, i_13_21_385_0,
    i_13_21_411_0, i_13_21_448_0, i_13_21_520_0, i_13_21_535_0,
    i_13_21_588_0, i_13_21_646_0, i_13_21_672_0, i_13_21_673_0,
    i_13_21_682_0, i_13_21_699_0, i_13_21_700_0, i_13_21_843_0,
    i_13_21_844_0, i_13_21_886_0, i_13_21_934_0, i_13_21_980_0,
    i_13_21_1102_0, i_13_21_1104_0, i_13_21_1105_0, i_13_21_1122_0,
    i_13_21_1222_0, i_13_21_1275_0, i_13_21_1276_0, i_13_21_1302_0,
    i_13_21_1311_0, i_13_21_1312_0, i_13_21_1402_0, i_13_21_1403_0,
    i_13_21_1428_0, i_13_21_1437_0, i_13_21_1438_0, i_13_21_1510_0,
    i_13_21_1600_0, i_13_21_1663_0, i_13_21_1665_0, i_13_21_1723_0,
    i_13_21_1725_0, i_13_21_1735_0, i_13_21_1777_0, i_13_21_1779_0,
    i_13_21_1798_0, i_13_21_1887_0, i_13_21_1888_0, i_13_21_1933_0,
    i_13_21_1935_0, i_13_21_1936_0, i_13_21_1947_0, i_13_21_1948_0,
    i_13_21_1995_0, i_13_21_1996_0, i_13_21_2004_0, i_13_21_2014_0,
    i_13_21_2029_0, i_13_21_2139_0, i_13_21_2140_0, i_13_21_2379_0,
    i_13_21_2383_0, i_13_21_2480_0, i_13_21_2551_0, i_13_21_2569_0,
    i_13_21_2599_0, i_13_21_2616_0, i_13_21_2650_0, i_13_21_2679_0,
    i_13_21_2697_0, i_13_21_2698_0, i_13_21_2712_0, i_13_21_2770_0,
    i_13_21_2824_0, i_13_21_2851_0, i_13_21_2901_0, i_13_21_2923_0,
    i_13_21_2958_0, i_13_21_3031_0, i_13_21_3208_0, i_13_21_3595_0,
    i_13_21_3596_0, i_13_21_3613_0, i_13_21_3742_0, i_13_21_3787_0,
    i_13_21_3930_0, i_13_21_3931_0, i_13_21_4063_0, i_13_21_4260_0,
    i_13_21_4302_0, i_13_21_4308_0, i_13_21_4309_0, i_13_21_4450_0,
    i_13_21_4596_0, i_13_21_4597_0, i_13_21_4606_0, i_13_21_4607_0;
  output o_13_21_0_0;
  assign o_13_21_0_0 = ~((~i_13_21_1798_0 & ~i_13_21_2770_0 & ~i_13_21_3930_0) | (~i_13_21_286_0 & ~i_13_21_1402_0 & ~i_13_21_2851_0) | (~i_13_21_70_0 & ~i_13_21_1779_0 & ~i_13_21_2697_0) | (~i_13_21_672_0 & ~i_13_21_1276_0 & ~i_13_21_3931_0 & ~i_13_21_4260_0));
endmodule



// Benchmark "kernel_13_22" written by ABC on Sun Jul 19 10:45:44 2020

module kernel_13_22 ( 
    i_13_22_142_0, i_13_22_169_0, i_13_22_224_0, i_13_22_240_0,
    i_13_22_310_0, i_13_22_327_0, i_13_22_328_0, i_13_22_340_0,
    i_13_22_367_0, i_13_22_472_0, i_13_22_529_0, i_13_22_553_0,
    i_13_22_599_0, i_13_22_607_0, i_13_22_618_0, i_13_22_619_0,
    i_13_22_620_0, i_13_22_670_0, i_13_22_689_0, i_13_22_699_0,
    i_13_22_725_0, i_13_22_780_0, i_13_22_824_0, i_13_22_912_0,
    i_13_22_980_0, i_13_22_1024_0, i_13_22_1078_0, i_13_22_1214_0,
    i_13_22_1259_0, i_13_22_1273_0, i_13_22_1483_0, i_13_22_1636_0,
    i_13_22_1687_0, i_13_22_1726_0, i_13_22_1749_0, i_13_22_1780_0,
    i_13_22_1781_0, i_13_22_1852_0, i_13_22_1888_0, i_13_22_1996_0,
    i_13_22_2020_0, i_13_22_2186_0, i_13_22_2200_0, i_13_22_2293_0,
    i_13_22_2391_0, i_13_22_2455_0, i_13_22_2461_0, i_13_22_2462_0,
    i_13_22_2464_0, i_13_22_2465_0, i_13_22_2470_0, i_13_22_2507_0,
    i_13_22_2509_0, i_13_22_2545_0, i_13_22_2633_0, i_13_22_2789_0,
    i_13_22_3109_0, i_13_22_3172_0, i_13_22_3174_0, i_13_22_3175_0,
    i_13_22_3262_0, i_13_22_3388_0, i_13_22_3409_0, i_13_22_3414_0,
    i_13_22_3415_0, i_13_22_3419_0, i_13_22_3432_0, i_13_22_3463_0,
    i_13_22_3477_0, i_13_22_3482_0, i_13_22_3535_0, i_13_22_3536_0,
    i_13_22_3544_0, i_13_22_3545_0, i_13_22_3562_0, i_13_22_3643_0,
    i_13_22_3666_0, i_13_22_3723_0, i_13_22_3734_0, i_13_22_3766_0,
    i_13_22_3910_0, i_13_22_3913_0, i_13_22_3914_0, i_13_22_3927_0,
    i_13_22_3928_0, i_13_22_4019_0, i_13_22_4099_0, i_13_22_4100_0,
    i_13_22_4126_0, i_13_22_4255_0, i_13_22_4333_0, i_13_22_4354_0,
    i_13_22_4381_0, i_13_22_4391_0, i_13_22_4396_0, i_13_22_4440_0,
    i_13_22_4449_0, i_13_22_4525_0, i_13_22_4534_0, i_13_22_4561_0,
    o_13_22_0_0  );
  input  i_13_22_142_0, i_13_22_169_0, i_13_22_224_0, i_13_22_240_0,
    i_13_22_310_0, i_13_22_327_0, i_13_22_328_0, i_13_22_340_0,
    i_13_22_367_0, i_13_22_472_0, i_13_22_529_0, i_13_22_553_0,
    i_13_22_599_0, i_13_22_607_0, i_13_22_618_0, i_13_22_619_0,
    i_13_22_620_0, i_13_22_670_0, i_13_22_689_0, i_13_22_699_0,
    i_13_22_725_0, i_13_22_780_0, i_13_22_824_0, i_13_22_912_0,
    i_13_22_980_0, i_13_22_1024_0, i_13_22_1078_0, i_13_22_1214_0,
    i_13_22_1259_0, i_13_22_1273_0, i_13_22_1483_0, i_13_22_1636_0,
    i_13_22_1687_0, i_13_22_1726_0, i_13_22_1749_0, i_13_22_1780_0,
    i_13_22_1781_0, i_13_22_1852_0, i_13_22_1888_0, i_13_22_1996_0,
    i_13_22_2020_0, i_13_22_2186_0, i_13_22_2200_0, i_13_22_2293_0,
    i_13_22_2391_0, i_13_22_2455_0, i_13_22_2461_0, i_13_22_2462_0,
    i_13_22_2464_0, i_13_22_2465_0, i_13_22_2470_0, i_13_22_2507_0,
    i_13_22_2509_0, i_13_22_2545_0, i_13_22_2633_0, i_13_22_2789_0,
    i_13_22_3109_0, i_13_22_3172_0, i_13_22_3174_0, i_13_22_3175_0,
    i_13_22_3262_0, i_13_22_3388_0, i_13_22_3409_0, i_13_22_3414_0,
    i_13_22_3415_0, i_13_22_3419_0, i_13_22_3432_0, i_13_22_3463_0,
    i_13_22_3477_0, i_13_22_3482_0, i_13_22_3535_0, i_13_22_3536_0,
    i_13_22_3544_0, i_13_22_3545_0, i_13_22_3562_0, i_13_22_3643_0,
    i_13_22_3666_0, i_13_22_3723_0, i_13_22_3734_0, i_13_22_3766_0,
    i_13_22_3910_0, i_13_22_3913_0, i_13_22_3914_0, i_13_22_3927_0,
    i_13_22_3928_0, i_13_22_4019_0, i_13_22_4099_0, i_13_22_4100_0,
    i_13_22_4126_0, i_13_22_4255_0, i_13_22_4333_0, i_13_22_4354_0,
    i_13_22_4381_0, i_13_22_4391_0, i_13_22_4396_0, i_13_22_4440_0,
    i_13_22_4449_0, i_13_22_4525_0, i_13_22_4534_0, i_13_22_4561_0;
  output o_13_22_0_0;
  assign o_13_22_0_0 = ~((i_13_22_3262_0 & (~i_13_22_3928_0 | (i_13_22_310_0 & ~i_13_22_3544_0 & ~i_13_22_3734_0 & ~i_13_22_3914_0))) | (~i_13_22_4561_0 & ((~i_13_22_328_0 & ~i_13_22_3535_0) | (~i_13_22_619_0 & ~i_13_22_824_0 & ~i_13_22_2465_0 & ~i_13_22_3463_0 & ~i_13_22_3914_0))) | (~i_13_22_340_0 & ~i_13_22_1024_0 & ~i_13_22_2200_0 & i_13_22_3109_0) | (~i_13_22_1780_0 & ~i_13_22_1781_0 & ~i_13_22_3175_0));
endmodule



// Benchmark "kernel_13_23" written by ABC on Sun Jul 19 10:45:45 2020

module kernel_13_23 ( 
    i_13_23_48_0, i_13_23_52_0, i_13_23_53_0, i_13_23_118_0, i_13_23_167_0,
    i_13_23_183_0, i_13_23_287_0, i_13_23_319_0, i_13_23_320_0,
    i_13_23_337_0, i_13_23_518_0, i_13_23_532_0, i_13_23_574_0,
    i_13_23_575_0, i_13_23_602_0, i_13_23_625_0, i_13_23_644_0,
    i_13_23_647_0, i_13_23_651_0, i_13_23_655_0, i_13_23_676_0,
    i_13_23_679_0, i_13_23_680_0, i_13_23_688_0, i_13_23_689_0,
    i_13_23_844_0, i_13_23_981_0, i_13_23_986_0, i_13_23_1048_0,
    i_13_23_1049_0, i_13_23_1070_0, i_13_23_1123_0, i_13_23_1124_0,
    i_13_23_1151_0, i_13_23_1228_0, i_13_23_1256_0, i_13_23_1385_0,
    i_13_23_1441_0, i_13_23_1465_0, i_13_23_1515_0, i_13_23_1519_0,
    i_13_23_1574_0, i_13_23_1712_0, i_13_23_1746_0, i_13_23_1751_0,
    i_13_23_1852_0, i_13_23_1857_0, i_13_23_1862_0, i_13_23_1888_0,
    i_13_23_2009_0, i_13_23_2050_0, i_13_23_2101_0, i_13_23_2136_0,
    i_13_23_2264_0, i_13_23_2267_0, i_13_23_2411_0, i_13_23_2556_0,
    i_13_23_2649_0, i_13_23_2651_0, i_13_23_2653_0, i_13_23_2654_0,
    i_13_23_2677_0, i_13_23_2678_0, i_13_23_2699_0, i_13_23_2722_0,
    i_13_23_2752_0, i_13_23_2753_0, i_13_23_2849_0, i_13_23_2984_0,
    i_13_23_3001_0, i_13_23_3146_0, i_13_23_3214_0, i_13_23_3217_0,
    i_13_23_3259_0, i_13_23_3260_0, i_13_23_3293_0, i_13_23_3398_0,
    i_13_23_3401_0, i_13_23_3437_0, i_13_23_3523_0, i_13_23_3734_0,
    i_13_23_3866_0, i_13_23_3888_0, i_13_23_3893_0, i_13_23_3909_0,
    i_13_23_3914_0, i_13_23_3991_0, i_13_23_3992_0, i_13_23_3995_0,
    i_13_23_4021_0, i_13_23_4067_0, i_13_23_4117_0, i_13_23_4307_0,
    i_13_23_4310_0, i_13_23_4318_0, i_13_23_4319_0, i_13_23_4513_0,
    i_13_23_4514_0, i_13_23_4556_0, i_13_23_4598_0,
    o_13_23_0_0  );
  input  i_13_23_48_0, i_13_23_52_0, i_13_23_53_0, i_13_23_118_0,
    i_13_23_167_0, i_13_23_183_0, i_13_23_287_0, i_13_23_319_0,
    i_13_23_320_0, i_13_23_337_0, i_13_23_518_0, i_13_23_532_0,
    i_13_23_574_0, i_13_23_575_0, i_13_23_602_0, i_13_23_625_0,
    i_13_23_644_0, i_13_23_647_0, i_13_23_651_0, i_13_23_655_0,
    i_13_23_676_0, i_13_23_679_0, i_13_23_680_0, i_13_23_688_0,
    i_13_23_689_0, i_13_23_844_0, i_13_23_981_0, i_13_23_986_0,
    i_13_23_1048_0, i_13_23_1049_0, i_13_23_1070_0, i_13_23_1123_0,
    i_13_23_1124_0, i_13_23_1151_0, i_13_23_1228_0, i_13_23_1256_0,
    i_13_23_1385_0, i_13_23_1441_0, i_13_23_1465_0, i_13_23_1515_0,
    i_13_23_1519_0, i_13_23_1574_0, i_13_23_1712_0, i_13_23_1746_0,
    i_13_23_1751_0, i_13_23_1852_0, i_13_23_1857_0, i_13_23_1862_0,
    i_13_23_1888_0, i_13_23_2009_0, i_13_23_2050_0, i_13_23_2101_0,
    i_13_23_2136_0, i_13_23_2264_0, i_13_23_2267_0, i_13_23_2411_0,
    i_13_23_2556_0, i_13_23_2649_0, i_13_23_2651_0, i_13_23_2653_0,
    i_13_23_2654_0, i_13_23_2677_0, i_13_23_2678_0, i_13_23_2699_0,
    i_13_23_2722_0, i_13_23_2752_0, i_13_23_2753_0, i_13_23_2849_0,
    i_13_23_2984_0, i_13_23_3001_0, i_13_23_3146_0, i_13_23_3214_0,
    i_13_23_3217_0, i_13_23_3259_0, i_13_23_3260_0, i_13_23_3293_0,
    i_13_23_3398_0, i_13_23_3401_0, i_13_23_3437_0, i_13_23_3523_0,
    i_13_23_3734_0, i_13_23_3866_0, i_13_23_3888_0, i_13_23_3893_0,
    i_13_23_3909_0, i_13_23_3914_0, i_13_23_3991_0, i_13_23_3992_0,
    i_13_23_3995_0, i_13_23_4021_0, i_13_23_4067_0, i_13_23_4117_0,
    i_13_23_4307_0, i_13_23_4310_0, i_13_23_4318_0, i_13_23_4319_0,
    i_13_23_4513_0, i_13_23_4514_0, i_13_23_4556_0, i_13_23_4598_0;
  output o_13_23_0_0;
  assign o_13_23_0_0 = ~((~i_13_23_3523_0 & (i_13_23_3909_0 | (~i_13_23_532_0 & ~i_13_23_1852_0))) | (~i_13_23_655_0 & ~i_13_23_679_0 & ~i_13_23_1124_0) | (i_13_23_1256_0 & ~i_13_23_2678_0) | (i_13_23_1228_0 & ~i_13_23_2649_0 & ~i_13_23_2654_0 & ~i_13_23_3214_0) | (~i_13_23_689_0 & ~i_13_23_2653_0 & ~i_13_23_3866_0));
endmodule



// Benchmark "kernel_13_24" written by ABC on Sun Jul 19 10:45:46 2020

module kernel_13_24 ( 
    i_13_24_40_0, i_13_24_52_0, i_13_24_94_0, i_13_24_101_0, i_13_24_241_0,
    i_13_24_251_0, i_13_24_259_0, i_13_24_278_0, i_13_24_310_0,
    i_13_24_334_0, i_13_24_377_0, i_13_24_519_0, i_13_24_607_0,
    i_13_24_619_0, i_13_24_620_0, i_13_24_663_0, i_13_24_700_0,
    i_13_24_701_0, i_13_24_858_0, i_13_24_868_0, i_13_24_871_0,
    i_13_24_886_0, i_13_24_929_0, i_13_24_980_0, i_13_24_1024_0,
    i_13_24_1075_0, i_13_24_1078_0, i_13_24_1079_0, i_13_24_1213_0,
    i_13_24_1214_0, i_13_24_1265_0, i_13_24_1282_0, i_13_24_1283_0,
    i_13_24_1397_0, i_13_24_1408_0, i_13_24_1426_0, i_13_24_1441_0,
    i_13_24_1480_0, i_13_24_1535_0, i_13_24_1561_0, i_13_24_1573_0,
    i_13_24_1609_0, i_13_24_1637_0, i_13_24_1642_0, i_13_24_1715_0,
    i_13_24_1776_0, i_13_24_1921_0, i_13_24_2104_0, i_13_24_2149_0,
    i_13_24_2150_0, i_13_24_2201_0, i_13_24_2260_0, i_13_24_2294_0,
    i_13_24_2455_0, i_13_24_2456_0, i_13_24_2546_0, i_13_24_2596_0,
    i_13_24_2647_0, i_13_24_2707_0, i_13_24_2768_0, i_13_24_2788_0,
    i_13_24_2789_0, i_13_24_2901_0, i_13_24_2959_0, i_13_24_3002_0,
    i_13_24_3005_0, i_13_24_3037_0, i_13_24_3292_0, i_13_24_3410_0,
    i_13_24_3419_0, i_13_24_3435_0, i_13_24_3449_0, i_13_24_3462_0,
    i_13_24_3464_0, i_13_24_3520_0, i_13_24_3559_0, i_13_24_3647_0,
    i_13_24_3650_0, i_13_24_3688_0, i_13_24_3689_0, i_13_24_3712_0,
    i_13_24_3847_0, i_13_24_3904_0, i_13_24_3918_0, i_13_24_3966_0,
    i_13_24_3994_0, i_13_24_4030_0, i_13_24_4090_0, i_13_24_4091_0,
    i_13_24_4157_0, i_13_24_4218_0, i_13_24_4250_0, i_13_24_4256_0,
    i_13_24_4271_0, i_13_24_4354_0, i_13_24_4361_0, i_13_24_4396_0,
    i_13_24_4450_0, i_13_24_4526_0, i_13_24_4541_0,
    o_13_24_0_0  );
  input  i_13_24_40_0, i_13_24_52_0, i_13_24_94_0, i_13_24_101_0,
    i_13_24_241_0, i_13_24_251_0, i_13_24_259_0, i_13_24_278_0,
    i_13_24_310_0, i_13_24_334_0, i_13_24_377_0, i_13_24_519_0,
    i_13_24_607_0, i_13_24_619_0, i_13_24_620_0, i_13_24_663_0,
    i_13_24_700_0, i_13_24_701_0, i_13_24_858_0, i_13_24_868_0,
    i_13_24_871_0, i_13_24_886_0, i_13_24_929_0, i_13_24_980_0,
    i_13_24_1024_0, i_13_24_1075_0, i_13_24_1078_0, i_13_24_1079_0,
    i_13_24_1213_0, i_13_24_1214_0, i_13_24_1265_0, i_13_24_1282_0,
    i_13_24_1283_0, i_13_24_1397_0, i_13_24_1408_0, i_13_24_1426_0,
    i_13_24_1441_0, i_13_24_1480_0, i_13_24_1535_0, i_13_24_1561_0,
    i_13_24_1573_0, i_13_24_1609_0, i_13_24_1637_0, i_13_24_1642_0,
    i_13_24_1715_0, i_13_24_1776_0, i_13_24_1921_0, i_13_24_2104_0,
    i_13_24_2149_0, i_13_24_2150_0, i_13_24_2201_0, i_13_24_2260_0,
    i_13_24_2294_0, i_13_24_2455_0, i_13_24_2456_0, i_13_24_2546_0,
    i_13_24_2596_0, i_13_24_2647_0, i_13_24_2707_0, i_13_24_2768_0,
    i_13_24_2788_0, i_13_24_2789_0, i_13_24_2901_0, i_13_24_2959_0,
    i_13_24_3002_0, i_13_24_3005_0, i_13_24_3037_0, i_13_24_3292_0,
    i_13_24_3410_0, i_13_24_3419_0, i_13_24_3435_0, i_13_24_3449_0,
    i_13_24_3462_0, i_13_24_3464_0, i_13_24_3520_0, i_13_24_3559_0,
    i_13_24_3647_0, i_13_24_3650_0, i_13_24_3688_0, i_13_24_3689_0,
    i_13_24_3712_0, i_13_24_3847_0, i_13_24_3904_0, i_13_24_3918_0,
    i_13_24_3966_0, i_13_24_3994_0, i_13_24_4030_0, i_13_24_4090_0,
    i_13_24_4091_0, i_13_24_4157_0, i_13_24_4218_0, i_13_24_4250_0,
    i_13_24_4256_0, i_13_24_4271_0, i_13_24_4354_0, i_13_24_4361_0,
    i_13_24_4396_0, i_13_24_4450_0, i_13_24_4526_0, i_13_24_4541_0;
  output o_13_24_0_0;
  assign o_13_24_0_0 = ~((~i_13_24_2788_0 & ((~i_13_24_619_0 & ~i_13_24_2455_0 & ~i_13_24_4218_0) | (~i_13_24_1078_0 & ~i_13_24_4450_0))) | (i_13_24_310_0 & ~i_13_24_1024_0 & ~i_13_24_4256_0) | (~i_13_24_3688_0 & i_13_24_4354_0 & i_13_24_4450_0));
endmodule



// Benchmark "kernel_13_25" written by ABC on Sun Jul 19 10:45:46 2020

module kernel_13_25 ( 
    i_13_25_17_0, i_13_25_64_0, i_13_25_111_0, i_13_25_139_0,
    i_13_25_160_0, i_13_25_169_0, i_13_25_170_0, i_13_25_188_0,
    i_13_25_251_0, i_13_25_259_0, i_13_25_310_0, i_13_25_320_0,
    i_13_25_340_0, i_13_25_341_0, i_13_25_457_0, i_13_25_458_0,
    i_13_25_493_0, i_13_25_494_0, i_13_25_619_0, i_13_25_657_0,
    i_13_25_728_0, i_13_25_814_0, i_13_25_817_0, i_13_25_818_0,
    i_13_25_945_0, i_13_25_980_0, i_13_25_1070_0, i_13_25_1079_0,
    i_13_25_1129_0, i_13_25_1142_0, i_13_25_1273_0, i_13_25_1303_0,
    i_13_25_1304_0, i_13_25_1305_0, i_13_25_1349_0, i_13_25_1364_0,
    i_13_25_1440_0, i_13_25_1441_0, i_13_25_1492_0, i_13_25_1565_0,
    i_13_25_1623_0, i_13_25_1640_0, i_13_25_1786_0, i_13_25_1808_0,
    i_13_25_1816_0, i_13_25_1817_0, i_13_25_1831_0, i_13_25_1839_0,
    i_13_25_1943_0, i_13_25_1989_0, i_13_25_1996_0, i_13_25_2123_0,
    i_13_25_2140_0, i_13_25_2150_0, i_13_25_2232_0, i_13_25_2267_0,
    i_13_25_2430_0, i_13_25_2431_0, i_13_25_2470_0, i_13_25_2519_0,
    i_13_25_2719_0, i_13_25_2752_0, i_13_25_2788_0, i_13_25_2789_0,
    i_13_25_2860_0, i_13_25_2941_0, i_13_25_2942_0, i_13_25_2969_0,
    i_13_25_3032_0, i_13_25_3040_0, i_13_25_3112_0, i_13_25_3141_0,
    i_13_25_3162_0, i_13_25_3220_0, i_13_25_3221_0, i_13_25_3428_0,
    i_13_25_3527_0, i_13_25_3541_0, i_13_25_3689_0, i_13_25_3769_0,
    i_13_25_3816_0, i_13_25_3892_0, i_13_25_4049_0, i_13_25_4057_0,
    i_13_25_4058_0, i_13_25_4066_0, i_13_25_4077_0, i_13_25_4081_0,
    i_13_25_4094_0, i_13_25_4237_0, i_13_25_4274_0, i_13_25_4319_0,
    i_13_25_4350_0, i_13_25_4363_0, i_13_25_4391_0, i_13_25_4512_0,
    i_13_25_4519_0, i_13_25_4534_0, i_13_25_4594_0, i_13_25_4604_0,
    o_13_25_0_0  );
  input  i_13_25_17_0, i_13_25_64_0, i_13_25_111_0, i_13_25_139_0,
    i_13_25_160_0, i_13_25_169_0, i_13_25_170_0, i_13_25_188_0,
    i_13_25_251_0, i_13_25_259_0, i_13_25_310_0, i_13_25_320_0,
    i_13_25_340_0, i_13_25_341_0, i_13_25_457_0, i_13_25_458_0,
    i_13_25_493_0, i_13_25_494_0, i_13_25_619_0, i_13_25_657_0,
    i_13_25_728_0, i_13_25_814_0, i_13_25_817_0, i_13_25_818_0,
    i_13_25_945_0, i_13_25_980_0, i_13_25_1070_0, i_13_25_1079_0,
    i_13_25_1129_0, i_13_25_1142_0, i_13_25_1273_0, i_13_25_1303_0,
    i_13_25_1304_0, i_13_25_1305_0, i_13_25_1349_0, i_13_25_1364_0,
    i_13_25_1440_0, i_13_25_1441_0, i_13_25_1492_0, i_13_25_1565_0,
    i_13_25_1623_0, i_13_25_1640_0, i_13_25_1786_0, i_13_25_1808_0,
    i_13_25_1816_0, i_13_25_1817_0, i_13_25_1831_0, i_13_25_1839_0,
    i_13_25_1943_0, i_13_25_1989_0, i_13_25_1996_0, i_13_25_2123_0,
    i_13_25_2140_0, i_13_25_2150_0, i_13_25_2232_0, i_13_25_2267_0,
    i_13_25_2430_0, i_13_25_2431_0, i_13_25_2470_0, i_13_25_2519_0,
    i_13_25_2719_0, i_13_25_2752_0, i_13_25_2788_0, i_13_25_2789_0,
    i_13_25_2860_0, i_13_25_2941_0, i_13_25_2942_0, i_13_25_2969_0,
    i_13_25_3032_0, i_13_25_3040_0, i_13_25_3112_0, i_13_25_3141_0,
    i_13_25_3162_0, i_13_25_3220_0, i_13_25_3221_0, i_13_25_3428_0,
    i_13_25_3527_0, i_13_25_3541_0, i_13_25_3689_0, i_13_25_3769_0,
    i_13_25_3816_0, i_13_25_3892_0, i_13_25_4049_0, i_13_25_4057_0,
    i_13_25_4058_0, i_13_25_4066_0, i_13_25_4077_0, i_13_25_4081_0,
    i_13_25_4094_0, i_13_25_4237_0, i_13_25_4274_0, i_13_25_4319_0,
    i_13_25_4350_0, i_13_25_4363_0, i_13_25_4391_0, i_13_25_4512_0,
    i_13_25_4519_0, i_13_25_4534_0, i_13_25_4594_0, i_13_25_4604_0;
  output o_13_25_0_0;
  assign o_13_25_0_0 = ~((~i_13_25_341_0 & ((~i_13_25_1349_0 & ~i_13_25_2941_0) | (i_13_25_139_0 & ~i_13_25_1808_0 & i_13_25_1831_0 & ~i_13_25_3221_0 & ~i_13_25_4058_0))) | (~i_13_25_1839_0 & ~i_13_25_2140_0 & ~i_13_25_3689_0) | (~i_13_25_1304_0 & ~i_13_25_2788_0 & ~i_13_25_4057_0) | (~i_13_25_4066_0 & i_13_25_4350_0) | (i_13_25_3541_0 & i_13_25_4081_0 & i_13_25_4363_0));
endmodule



// Benchmark "kernel_13_26" written by ABC on Sun Jul 19 10:45:47 2020

module kernel_13_26 ( 
    i_13_26_40_0, i_13_26_45_0, i_13_26_48_0, i_13_26_76_0, i_13_26_90_0,
    i_13_26_91_0, i_13_26_118_0, i_13_26_121_0, i_13_26_163_0,
    i_13_26_333_0, i_13_26_336_0, i_13_26_337_0, i_13_26_374_0,
    i_13_26_377_0, i_13_26_379_0, i_13_26_410_0, i_13_26_450_0,
    i_13_26_567_0, i_13_26_643_0, i_13_26_667_0, i_13_26_688_0,
    i_13_26_694_0, i_13_26_729_0, i_13_26_822_0, i_13_26_823_0,
    i_13_26_850_0, i_13_26_1063_0, i_13_26_1115_0, i_13_26_1120_0,
    i_13_26_1243_0, i_13_26_1267_0, i_13_26_1269_0, i_13_26_1341_0,
    i_13_26_1440_0, i_13_26_1441_0, i_13_26_1498_0, i_13_26_1782_0,
    i_13_26_1845_0, i_13_26_1924_0, i_13_26_1947_0, i_13_26_2116_0,
    i_13_26_2173_0, i_13_26_2197_0, i_13_26_2205_0, i_13_26_2206_0,
    i_13_26_2233_0, i_13_26_2235_0, i_13_26_2317_0, i_13_26_2421_0,
    i_13_26_2424_0, i_13_26_2539_0, i_13_26_2584_0, i_13_26_2613_0,
    i_13_26_2746_0, i_13_26_2781_0, i_13_26_2790_0, i_13_26_2853_0,
    i_13_26_2906_0, i_13_26_2916_0, i_13_26_2935_0, i_13_26_2966_0,
    i_13_26_2969_0, i_13_26_3016_0, i_13_26_3060_0, i_13_26_3108_0,
    i_13_26_3204_0, i_13_26_3213_0, i_13_26_3214_0, i_13_26_3217_0,
    i_13_26_3231_0, i_13_26_3234_0, i_13_26_3239_0, i_13_26_3241_0,
    i_13_26_3367_0, i_13_26_3398_0, i_13_26_3475_0, i_13_26_3477_0,
    i_13_26_3609_0, i_13_26_3717_0, i_13_26_3754_0, i_13_26_3817_0,
    i_13_26_3862_0, i_13_26_3870_0, i_13_26_3873_0, i_13_26_3889_0,
    i_13_26_3925_0, i_13_26_4014_0, i_13_26_4060_0, i_13_26_4158_0,
    i_13_26_4186_0, i_13_26_4189_0, i_13_26_4266_0, i_13_26_4267_0,
    i_13_26_4347_0, i_13_26_4348_0, i_13_26_4423_0, i_13_26_4530_0,
    i_13_26_4588_0, i_13_26_4594_0, i_13_26_4600_0,
    o_13_26_0_0  );
  input  i_13_26_40_0, i_13_26_45_0, i_13_26_48_0, i_13_26_76_0,
    i_13_26_90_0, i_13_26_91_0, i_13_26_118_0, i_13_26_121_0,
    i_13_26_163_0, i_13_26_333_0, i_13_26_336_0, i_13_26_337_0,
    i_13_26_374_0, i_13_26_377_0, i_13_26_379_0, i_13_26_410_0,
    i_13_26_450_0, i_13_26_567_0, i_13_26_643_0, i_13_26_667_0,
    i_13_26_688_0, i_13_26_694_0, i_13_26_729_0, i_13_26_822_0,
    i_13_26_823_0, i_13_26_850_0, i_13_26_1063_0, i_13_26_1115_0,
    i_13_26_1120_0, i_13_26_1243_0, i_13_26_1267_0, i_13_26_1269_0,
    i_13_26_1341_0, i_13_26_1440_0, i_13_26_1441_0, i_13_26_1498_0,
    i_13_26_1782_0, i_13_26_1845_0, i_13_26_1924_0, i_13_26_1947_0,
    i_13_26_2116_0, i_13_26_2173_0, i_13_26_2197_0, i_13_26_2205_0,
    i_13_26_2206_0, i_13_26_2233_0, i_13_26_2235_0, i_13_26_2317_0,
    i_13_26_2421_0, i_13_26_2424_0, i_13_26_2539_0, i_13_26_2584_0,
    i_13_26_2613_0, i_13_26_2746_0, i_13_26_2781_0, i_13_26_2790_0,
    i_13_26_2853_0, i_13_26_2906_0, i_13_26_2916_0, i_13_26_2935_0,
    i_13_26_2966_0, i_13_26_2969_0, i_13_26_3016_0, i_13_26_3060_0,
    i_13_26_3108_0, i_13_26_3204_0, i_13_26_3213_0, i_13_26_3214_0,
    i_13_26_3217_0, i_13_26_3231_0, i_13_26_3234_0, i_13_26_3239_0,
    i_13_26_3241_0, i_13_26_3367_0, i_13_26_3398_0, i_13_26_3475_0,
    i_13_26_3477_0, i_13_26_3609_0, i_13_26_3717_0, i_13_26_3754_0,
    i_13_26_3817_0, i_13_26_3862_0, i_13_26_3870_0, i_13_26_3873_0,
    i_13_26_3889_0, i_13_26_3925_0, i_13_26_4014_0, i_13_26_4060_0,
    i_13_26_4158_0, i_13_26_4186_0, i_13_26_4189_0, i_13_26_4266_0,
    i_13_26_4267_0, i_13_26_4347_0, i_13_26_4348_0, i_13_26_4423_0,
    i_13_26_4530_0, i_13_26_4588_0, i_13_26_4594_0, i_13_26_4600_0;
  output o_13_26_0_0;
  assign o_13_26_0_0 = ~((~i_13_26_3213_0 & (~i_13_26_3214_0 | (i_13_26_823_0 & ~i_13_26_3817_0 & ~i_13_26_3873_0 & ~i_13_26_4347_0))) | (i_13_26_76_0 & i_13_26_3241_0 & i_13_26_3398_0) | (~i_13_26_337_0 & i_13_26_4189_0 & ~i_13_26_4347_0));
endmodule



// Benchmark "kernel_13_27" written by ABC on Sun Jul 19 10:45:48 2020

module kernel_13_27 ( 
    i_13_27_23_0, i_13_27_28_0, i_13_27_29_0, i_13_27_41_0, i_13_27_92_0,
    i_13_27_112_0, i_13_27_244_0, i_13_27_257_0, i_13_27_266_0,
    i_13_27_367_0, i_13_27_370_0, i_13_27_373_0, i_13_27_376_0,
    i_13_27_384_0, i_13_27_391_0, i_13_27_442_0, i_13_27_443_0,
    i_13_27_463_0, i_13_27_483_0, i_13_27_526_0, i_13_27_604_0,
    i_13_27_605_0, i_13_27_608_0, i_13_27_613_0, i_13_27_668_0,
    i_13_27_730_0, i_13_27_797_0, i_13_27_830_0, i_13_27_832_0,
    i_13_27_947_0, i_13_27_1082_0, i_13_27_1085_0, i_13_27_1145_0,
    i_13_27_1226_0, i_13_27_1271_0, i_13_27_1318_0, i_13_27_1423_0,
    i_13_27_1424_0, i_13_27_1473_0, i_13_27_1487_0, i_13_27_1496_0,
    i_13_27_1514_0, i_13_27_1571_0, i_13_27_1621_0, i_13_27_1721_0,
    i_13_27_1730_0, i_13_27_1750_0, i_13_27_1804_0, i_13_27_1837_0,
    i_13_27_1838_0, i_13_27_1840_0, i_13_27_1841_0, i_13_27_1851_0,
    i_13_27_2017_0, i_13_27_2112_0, i_13_27_2137_0, i_13_27_2170_0,
    i_13_27_2171_0, i_13_27_2173_0, i_13_27_2207_0, i_13_27_2380_0,
    i_13_27_2422_0, i_13_27_2423_0, i_13_27_2426_0, i_13_27_2431_0,
    i_13_27_2432_0, i_13_27_2435_0, i_13_27_2471_0, i_13_27_2579_0,
    i_13_27_2938_0, i_13_27_3018_0, i_13_27_3034_0, i_13_27_3127_0,
    i_13_27_3237_0, i_13_27_3260_0, i_13_27_3422_0, i_13_27_3425_0,
    i_13_27_3433_0, i_13_27_3503_0, i_13_27_3547_0, i_13_27_3622_0,
    i_13_27_3667_0, i_13_27_3763_0, i_13_27_3767_0, i_13_27_3871_0,
    i_13_27_3872_0, i_13_27_3875_0, i_13_27_3889_0, i_13_27_3964_0,
    i_13_27_4033_0, i_13_27_4047_0, i_13_27_4079_0, i_13_27_4089_0,
    i_13_27_4118_0, i_13_27_4343_0, i_13_27_4349_0, i_13_27_4351_0,
    i_13_27_4352_0, i_13_27_4541_0, i_13_27_4558_0,
    o_13_27_0_0  );
  input  i_13_27_23_0, i_13_27_28_0, i_13_27_29_0, i_13_27_41_0,
    i_13_27_92_0, i_13_27_112_0, i_13_27_244_0, i_13_27_257_0,
    i_13_27_266_0, i_13_27_367_0, i_13_27_370_0, i_13_27_373_0,
    i_13_27_376_0, i_13_27_384_0, i_13_27_391_0, i_13_27_442_0,
    i_13_27_443_0, i_13_27_463_0, i_13_27_483_0, i_13_27_526_0,
    i_13_27_604_0, i_13_27_605_0, i_13_27_608_0, i_13_27_613_0,
    i_13_27_668_0, i_13_27_730_0, i_13_27_797_0, i_13_27_830_0,
    i_13_27_832_0, i_13_27_947_0, i_13_27_1082_0, i_13_27_1085_0,
    i_13_27_1145_0, i_13_27_1226_0, i_13_27_1271_0, i_13_27_1318_0,
    i_13_27_1423_0, i_13_27_1424_0, i_13_27_1473_0, i_13_27_1487_0,
    i_13_27_1496_0, i_13_27_1514_0, i_13_27_1571_0, i_13_27_1621_0,
    i_13_27_1721_0, i_13_27_1730_0, i_13_27_1750_0, i_13_27_1804_0,
    i_13_27_1837_0, i_13_27_1838_0, i_13_27_1840_0, i_13_27_1841_0,
    i_13_27_1851_0, i_13_27_2017_0, i_13_27_2112_0, i_13_27_2137_0,
    i_13_27_2170_0, i_13_27_2171_0, i_13_27_2173_0, i_13_27_2207_0,
    i_13_27_2380_0, i_13_27_2422_0, i_13_27_2423_0, i_13_27_2426_0,
    i_13_27_2431_0, i_13_27_2432_0, i_13_27_2435_0, i_13_27_2471_0,
    i_13_27_2579_0, i_13_27_2938_0, i_13_27_3018_0, i_13_27_3034_0,
    i_13_27_3127_0, i_13_27_3237_0, i_13_27_3260_0, i_13_27_3422_0,
    i_13_27_3425_0, i_13_27_3433_0, i_13_27_3503_0, i_13_27_3547_0,
    i_13_27_3622_0, i_13_27_3667_0, i_13_27_3763_0, i_13_27_3767_0,
    i_13_27_3871_0, i_13_27_3872_0, i_13_27_3875_0, i_13_27_3889_0,
    i_13_27_3964_0, i_13_27_4033_0, i_13_27_4047_0, i_13_27_4079_0,
    i_13_27_4089_0, i_13_27_4118_0, i_13_27_4343_0, i_13_27_4349_0,
    i_13_27_4351_0, i_13_27_4352_0, i_13_27_4541_0, i_13_27_4558_0;
  output o_13_27_0_0;
  assign o_13_27_0_0 = ~(~i_13_27_2431_0 | ~i_13_27_4352_0);
endmodule



// Benchmark "kernel_13_28" written by ABC on Sun Jul 19 10:45:49 2020

module kernel_13_28 ( 
    i_13_28_72_0, i_13_28_318_0, i_13_28_342_0, i_13_28_406_0,
    i_13_28_433_0, i_13_28_469_0, i_13_28_531_0, i_13_28_532_0,
    i_13_28_536_0, i_13_28_550_0, i_13_28_553_0, i_13_28_562_0,
    i_13_28_651_0, i_13_28_660_0, i_13_28_661_0, i_13_28_666_0,
    i_13_28_669_0, i_13_28_676_0, i_13_28_693_0, i_13_28_694_0,
    i_13_28_696_0, i_13_28_700_0, i_13_28_828_0, i_13_28_843_0,
    i_13_28_885_0, i_13_28_930_0, i_13_28_942_0, i_13_28_1098_0,
    i_13_28_1116_0, i_13_28_1117_0, i_13_28_1144_0, i_13_28_1263_0,
    i_13_28_1269_0, i_13_28_1279_0, i_13_28_1656_0, i_13_28_1657_0,
    i_13_28_1659_0, i_13_28_1660_0, i_13_28_1693_0, i_13_28_1719_0,
    i_13_28_1731_0, i_13_28_1774_0, i_13_28_1791_0, i_13_28_1836_0,
    i_13_28_1915_0, i_13_28_2016_0, i_13_28_2017_0, i_13_28_2339_0,
    i_13_28_2398_0, i_13_28_2413_0, i_13_28_2442_0, i_13_28_2460_0,
    i_13_28_2466_0, i_13_28_2467_0, i_13_28_2692_0, i_13_28_2844_0,
    i_13_28_2845_0, i_13_28_2881_0, i_13_28_2888_0, i_13_28_2925_0,
    i_13_28_2958_0, i_13_28_2983_0, i_13_28_3025_0, i_13_28_3061_0,
    i_13_28_3101_0, i_13_28_3114_0, i_13_28_3153_0, i_13_28_3207_0,
    i_13_28_3216_0, i_13_28_3258_0, i_13_28_3372_0, i_13_28_3531_0,
    i_13_28_3549_0, i_13_28_3579_0, i_13_28_3592_0, i_13_28_3639_0,
    i_13_28_3654_0, i_13_28_3703_0, i_13_28_3738_0, i_13_28_3739_0,
    i_13_28_3862_0, i_13_28_3875_0, i_13_28_3906_0, i_13_28_3987_0,
    i_13_28_4015_0, i_13_28_4077_0, i_13_28_4123_0, i_13_28_4185_0,
    i_13_28_4186_0, i_13_28_4212_0, i_13_28_4279_0, i_13_28_4323_0,
    i_13_28_4329_0, i_13_28_4339_0, i_13_28_4368_0, i_13_28_4512_0,
    i_13_28_4590_0, i_13_28_4599_0, i_13_28_4600_0, i_13_28_4602_0,
    o_13_28_0_0  );
  input  i_13_28_72_0, i_13_28_318_0, i_13_28_342_0, i_13_28_406_0,
    i_13_28_433_0, i_13_28_469_0, i_13_28_531_0, i_13_28_532_0,
    i_13_28_536_0, i_13_28_550_0, i_13_28_553_0, i_13_28_562_0,
    i_13_28_651_0, i_13_28_660_0, i_13_28_661_0, i_13_28_666_0,
    i_13_28_669_0, i_13_28_676_0, i_13_28_693_0, i_13_28_694_0,
    i_13_28_696_0, i_13_28_700_0, i_13_28_828_0, i_13_28_843_0,
    i_13_28_885_0, i_13_28_930_0, i_13_28_942_0, i_13_28_1098_0,
    i_13_28_1116_0, i_13_28_1117_0, i_13_28_1144_0, i_13_28_1263_0,
    i_13_28_1269_0, i_13_28_1279_0, i_13_28_1656_0, i_13_28_1657_0,
    i_13_28_1659_0, i_13_28_1660_0, i_13_28_1693_0, i_13_28_1719_0,
    i_13_28_1731_0, i_13_28_1774_0, i_13_28_1791_0, i_13_28_1836_0,
    i_13_28_1915_0, i_13_28_2016_0, i_13_28_2017_0, i_13_28_2339_0,
    i_13_28_2398_0, i_13_28_2413_0, i_13_28_2442_0, i_13_28_2460_0,
    i_13_28_2466_0, i_13_28_2467_0, i_13_28_2692_0, i_13_28_2844_0,
    i_13_28_2845_0, i_13_28_2881_0, i_13_28_2888_0, i_13_28_2925_0,
    i_13_28_2958_0, i_13_28_2983_0, i_13_28_3025_0, i_13_28_3061_0,
    i_13_28_3101_0, i_13_28_3114_0, i_13_28_3153_0, i_13_28_3207_0,
    i_13_28_3216_0, i_13_28_3258_0, i_13_28_3372_0, i_13_28_3531_0,
    i_13_28_3549_0, i_13_28_3579_0, i_13_28_3592_0, i_13_28_3639_0,
    i_13_28_3654_0, i_13_28_3703_0, i_13_28_3738_0, i_13_28_3739_0,
    i_13_28_3862_0, i_13_28_3875_0, i_13_28_3906_0, i_13_28_3987_0,
    i_13_28_4015_0, i_13_28_4077_0, i_13_28_4123_0, i_13_28_4185_0,
    i_13_28_4186_0, i_13_28_4212_0, i_13_28_4279_0, i_13_28_4323_0,
    i_13_28_4329_0, i_13_28_4339_0, i_13_28_4368_0, i_13_28_4512_0,
    i_13_28_4590_0, i_13_28_4599_0, i_13_28_4600_0, i_13_28_4602_0;
  output o_13_28_0_0;
  assign o_13_28_0_0 = ~((~i_13_28_3739_0 & ~i_13_28_4512_0) | (~i_13_28_2016_0 & ~i_13_28_4212_0) | (~i_13_28_3258_0 & ~i_13_28_4186_0) | (~i_13_28_1659_0 & ~i_13_28_2844_0 & ~i_13_28_2881_0 & ~i_13_28_3987_0));
endmodule



// Benchmark "kernel_13_29" written by ABC on Sun Jul 19 10:45:50 2020

module kernel_13_29 ( 
    i_13_29_49_0, i_13_29_69_0, i_13_29_94_0, i_13_29_282_0, i_13_29_321_0,
    i_13_29_327_0, i_13_29_328_0, i_13_29_375_0, i_13_29_411_0,
    i_13_29_529_0, i_13_29_547_0, i_13_29_598_0, i_13_29_624_0,
    i_13_29_717_0, i_13_29_745_0, i_13_29_780_0, i_13_29_796_0,
    i_13_29_825_0, i_13_29_826_0, i_13_29_861_0, i_13_29_862_0,
    i_13_29_894_0, i_13_29_912_0, i_13_29_922_0, i_13_29_1023_0,
    i_13_29_1077_0, i_13_29_1257_0, i_13_29_1258_0, i_13_29_1320_0,
    i_13_29_1321_0, i_13_29_1383_0, i_13_29_1410_0, i_13_29_1491_0,
    i_13_29_1501_0, i_13_29_1608_0, i_13_29_1635_0, i_13_29_1643_0,
    i_13_29_1762_0, i_13_29_1770_0, i_13_29_1777_0, i_13_29_1861_0,
    i_13_29_2032_0, i_13_29_2059_0, i_13_29_2060_0, i_13_29_2139_0,
    i_13_29_2185_0, i_13_29_2240_0, i_13_29_2310_0, i_13_29_2427_0,
    i_13_29_2454_0, i_13_29_2461_0, i_13_29_2613_0, i_13_29_2632_0,
    i_13_29_2653_0, i_13_29_2654_0, i_13_29_2679_0, i_13_29_2749_0,
    i_13_29_2762_0, i_13_29_2848_0, i_13_29_2883_0, i_13_29_2886_0,
    i_13_29_2966_0, i_13_29_3056_0, i_13_29_3145_0, i_13_29_3174_0,
    i_13_29_3175_0, i_13_29_3219_0, i_13_29_3347_0, i_13_29_3392_0,
    i_13_29_3417_0, i_13_29_3418_0, i_13_29_3432_0, i_13_29_3450_0,
    i_13_29_3463_0, i_13_29_3490_0, i_13_29_3535_0, i_13_29_3550_0,
    i_13_29_3562_0, i_13_29_3571_0, i_13_29_3579_0, i_13_29_3640_0,
    i_13_29_3702_0, i_13_29_3723_0, i_13_29_3733_0, i_13_29_3786_0,
    i_13_29_3793_0, i_13_29_3846_0, i_13_29_3876_0, i_13_29_3912_0,
    i_13_29_3913_0, i_13_29_3948_0, i_13_29_4012_0, i_13_29_4238_0,
    i_13_29_4274_0, i_13_29_4380_0, i_13_29_4381_0, i_13_29_4443_0,
    i_13_29_4560_0, i_13_29_4561_0, i_13_29_4597_0,
    o_13_29_0_0  );
  input  i_13_29_49_0, i_13_29_69_0, i_13_29_94_0, i_13_29_282_0,
    i_13_29_321_0, i_13_29_327_0, i_13_29_328_0, i_13_29_375_0,
    i_13_29_411_0, i_13_29_529_0, i_13_29_547_0, i_13_29_598_0,
    i_13_29_624_0, i_13_29_717_0, i_13_29_745_0, i_13_29_780_0,
    i_13_29_796_0, i_13_29_825_0, i_13_29_826_0, i_13_29_861_0,
    i_13_29_862_0, i_13_29_894_0, i_13_29_912_0, i_13_29_922_0,
    i_13_29_1023_0, i_13_29_1077_0, i_13_29_1257_0, i_13_29_1258_0,
    i_13_29_1320_0, i_13_29_1321_0, i_13_29_1383_0, i_13_29_1410_0,
    i_13_29_1491_0, i_13_29_1501_0, i_13_29_1608_0, i_13_29_1635_0,
    i_13_29_1643_0, i_13_29_1762_0, i_13_29_1770_0, i_13_29_1777_0,
    i_13_29_1861_0, i_13_29_2032_0, i_13_29_2059_0, i_13_29_2060_0,
    i_13_29_2139_0, i_13_29_2185_0, i_13_29_2240_0, i_13_29_2310_0,
    i_13_29_2427_0, i_13_29_2454_0, i_13_29_2461_0, i_13_29_2613_0,
    i_13_29_2632_0, i_13_29_2653_0, i_13_29_2654_0, i_13_29_2679_0,
    i_13_29_2749_0, i_13_29_2762_0, i_13_29_2848_0, i_13_29_2883_0,
    i_13_29_2886_0, i_13_29_2966_0, i_13_29_3056_0, i_13_29_3145_0,
    i_13_29_3174_0, i_13_29_3175_0, i_13_29_3219_0, i_13_29_3347_0,
    i_13_29_3392_0, i_13_29_3417_0, i_13_29_3418_0, i_13_29_3432_0,
    i_13_29_3450_0, i_13_29_3463_0, i_13_29_3490_0, i_13_29_3535_0,
    i_13_29_3550_0, i_13_29_3562_0, i_13_29_3571_0, i_13_29_3579_0,
    i_13_29_3640_0, i_13_29_3702_0, i_13_29_3723_0, i_13_29_3733_0,
    i_13_29_3786_0, i_13_29_3793_0, i_13_29_3846_0, i_13_29_3876_0,
    i_13_29_3912_0, i_13_29_3913_0, i_13_29_3948_0, i_13_29_4012_0,
    i_13_29_4238_0, i_13_29_4274_0, i_13_29_4380_0, i_13_29_4381_0,
    i_13_29_4443_0, i_13_29_4560_0, i_13_29_4561_0, i_13_29_4597_0;
  output o_13_29_0_0;
  assign o_13_29_0_0 = ~(i_13_29_2185_0 | ~i_13_29_3174_0);
endmodule



// Benchmark "kernel_13_30" written by ABC on Sun Jul 19 10:45:51 2020

module kernel_13_30 ( 
    i_13_30_108_0, i_13_30_121_0, i_13_30_274_0, i_13_30_275_0,
    i_13_30_309_0, i_13_30_310_0, i_13_30_337_0, i_13_30_357_0,
    i_13_30_454_0, i_13_30_558_0, i_13_30_559_0, i_13_30_562_0,
    i_13_30_618_0, i_13_30_633_0, i_13_30_658_0, i_13_30_850_0,
    i_13_30_851_0, i_13_30_1064_0, i_13_30_1081_0, i_13_30_1085_0,
    i_13_30_1228_0, i_13_30_1266_0, i_13_30_1309_0, i_13_30_1336_0,
    i_13_30_1396_0, i_13_30_1407_0, i_13_30_1471_0, i_13_30_1525_0,
    i_13_30_1549_0, i_13_30_1597_0, i_13_30_1621_0, i_13_30_1624_0,
    i_13_30_1629_0, i_13_30_1678_0, i_13_30_1719_0, i_13_30_1783_0,
    i_13_30_1787_0, i_13_30_1813_0, i_13_30_1841_0, i_13_30_1858_0,
    i_13_30_1914_0, i_13_30_1929_0, i_13_30_1936_0, i_13_30_1937_0,
    i_13_30_2110_0, i_13_30_2170_0, i_13_30_2202_0, i_13_30_2431_0,
    i_13_30_2542_0, i_13_30_2563_0, i_13_30_2564_0, i_13_30_2592_0,
    i_13_30_2709_0, i_13_30_2712_0, i_13_30_2768_0, i_13_30_2855_0,
    i_13_30_2859_0, i_13_30_2903_0, i_13_30_2916_0, i_13_30_2984_0,
    i_13_30_3061_0, i_13_30_3062_0, i_13_30_3096_0, i_13_30_3097_0,
    i_13_30_3100_0, i_13_30_3106_0, i_13_30_3153_0, i_13_30_3160_0,
    i_13_30_3217_0, i_13_30_3231_0, i_13_30_3232_0, i_13_30_3234_0,
    i_13_30_3235_0, i_13_30_3276_0, i_13_30_3285_0, i_13_30_3450_0,
    i_13_30_3496_0, i_13_30_3520_0, i_13_30_3537_0, i_13_30_3538_0,
    i_13_30_3600_0, i_13_30_3614_0, i_13_30_3682_0, i_13_30_3684_0,
    i_13_30_3685_0, i_13_30_3720_0, i_13_30_3753_0, i_13_30_3865_0,
    i_13_30_3878_0, i_13_30_3904_0, i_13_30_3937_0, i_13_30_4090_0,
    i_13_30_4091_0, i_13_30_4189_0, i_13_30_4249_0, i_13_30_4302_0,
    i_13_30_4351_0, i_13_30_4385_0, i_13_30_4517_0, i_13_30_4554_0,
    o_13_30_0_0  );
  input  i_13_30_108_0, i_13_30_121_0, i_13_30_274_0, i_13_30_275_0,
    i_13_30_309_0, i_13_30_310_0, i_13_30_337_0, i_13_30_357_0,
    i_13_30_454_0, i_13_30_558_0, i_13_30_559_0, i_13_30_562_0,
    i_13_30_618_0, i_13_30_633_0, i_13_30_658_0, i_13_30_850_0,
    i_13_30_851_0, i_13_30_1064_0, i_13_30_1081_0, i_13_30_1085_0,
    i_13_30_1228_0, i_13_30_1266_0, i_13_30_1309_0, i_13_30_1336_0,
    i_13_30_1396_0, i_13_30_1407_0, i_13_30_1471_0, i_13_30_1525_0,
    i_13_30_1549_0, i_13_30_1597_0, i_13_30_1621_0, i_13_30_1624_0,
    i_13_30_1629_0, i_13_30_1678_0, i_13_30_1719_0, i_13_30_1783_0,
    i_13_30_1787_0, i_13_30_1813_0, i_13_30_1841_0, i_13_30_1858_0,
    i_13_30_1914_0, i_13_30_1929_0, i_13_30_1936_0, i_13_30_1937_0,
    i_13_30_2110_0, i_13_30_2170_0, i_13_30_2202_0, i_13_30_2431_0,
    i_13_30_2542_0, i_13_30_2563_0, i_13_30_2564_0, i_13_30_2592_0,
    i_13_30_2709_0, i_13_30_2712_0, i_13_30_2768_0, i_13_30_2855_0,
    i_13_30_2859_0, i_13_30_2903_0, i_13_30_2916_0, i_13_30_2984_0,
    i_13_30_3061_0, i_13_30_3062_0, i_13_30_3096_0, i_13_30_3097_0,
    i_13_30_3100_0, i_13_30_3106_0, i_13_30_3153_0, i_13_30_3160_0,
    i_13_30_3217_0, i_13_30_3231_0, i_13_30_3232_0, i_13_30_3234_0,
    i_13_30_3235_0, i_13_30_3276_0, i_13_30_3285_0, i_13_30_3450_0,
    i_13_30_3496_0, i_13_30_3520_0, i_13_30_3537_0, i_13_30_3538_0,
    i_13_30_3600_0, i_13_30_3614_0, i_13_30_3682_0, i_13_30_3684_0,
    i_13_30_3685_0, i_13_30_3720_0, i_13_30_3753_0, i_13_30_3865_0,
    i_13_30_3878_0, i_13_30_3904_0, i_13_30_3937_0, i_13_30_4090_0,
    i_13_30_4091_0, i_13_30_4189_0, i_13_30_4249_0, i_13_30_4302_0,
    i_13_30_4351_0, i_13_30_4385_0, i_13_30_4517_0, i_13_30_4554_0;
  output o_13_30_0_0;
  assign o_13_30_0_0 = ~((~i_13_30_274_0 & (~i_13_30_3685_0 | i_13_30_3904_0)) | (i_13_30_310_0 & ~i_13_30_558_0) | (~i_13_30_275_0 & ~i_13_30_2431_0 & ~i_13_30_3682_0) | (i_13_30_3904_0 & ~i_13_30_4351_0) | (~i_13_30_559_0 & ~i_13_30_3904_0 & ~i_13_30_4554_0));
endmodule



// Benchmark "kernel_13_31" written by ABC on Sun Jul 19 10:45:51 2020

module kernel_13_31 ( 
    i_13_31_34_0, i_13_31_44_0, i_13_31_71_0, i_13_31_79_0, i_13_31_114_0,
    i_13_31_138_0, i_13_31_142_0, i_13_31_231_0, i_13_31_232_0,
    i_13_31_411_0, i_13_31_447_0, i_13_31_448_0, i_13_31_480_0,
    i_13_31_537_0, i_13_31_538_0, i_13_31_556_0, i_13_31_584_0,
    i_13_31_589_0, i_13_31_593_0, i_13_31_600_0, i_13_31_606_0,
    i_13_31_609_0, i_13_31_610_0, i_13_31_646_0, i_13_31_660_0,
    i_13_31_673_0, i_13_31_681_0, i_13_31_682_0, i_13_31_688_0,
    i_13_31_760_0, i_13_31_763_0, i_13_31_952_0, i_13_31_1119_0,
    i_13_31_1150_0, i_13_31_1275_0, i_13_31_1308_0, i_13_31_1311_0,
    i_13_31_1312_0, i_13_31_1344_0, i_13_31_1402_0, i_13_31_1428_0,
    i_13_31_1510_0, i_13_31_1626_0, i_13_31_1663_0, i_13_31_1672_0,
    i_13_31_1713_0, i_13_31_1725_0, i_13_31_1726_0, i_13_31_1734_0,
    i_13_31_1780_0, i_13_31_1798_0, i_13_31_1887_0, i_13_31_1911_0,
    i_13_31_1912_0, i_13_31_1923_0, i_13_31_1934_0, i_13_31_1947_0,
    i_13_31_1948_0, i_13_31_2175_0, i_13_31_2321_0, i_13_31_2379_0,
    i_13_31_2552_0, i_13_31_2598_0, i_13_31_2599_0, i_13_31_2679_0,
    i_13_31_2712_0, i_13_31_2752_0, i_13_31_2847_0, i_13_31_2850_0,
    i_13_31_2851_0, i_13_31_2856_0, i_13_31_2877_0, i_13_31_2923_0,
    i_13_31_3046_0, i_13_31_3067_0, i_13_31_3103_0, i_13_31_3129_0,
    i_13_31_3370_0, i_13_31_3371_0, i_13_31_3652_0, i_13_31_3668_0,
    i_13_31_3786_0, i_13_31_3930_0, i_13_31_3931_0, i_13_31_3940_0,
    i_13_31_4154_0, i_13_31_4188_0, i_13_31_4189_0, i_13_31_4219_0,
    i_13_31_4296_0, i_13_31_4297_0, i_13_31_4306_0, i_13_31_4308_0,
    i_13_31_4325_0, i_13_31_4336_0, i_13_31_4435_0, i_13_31_4450_0,
    i_13_31_4539_0, i_13_31_4596_0, i_13_31_4597_0,
    o_13_31_0_0  );
  input  i_13_31_34_0, i_13_31_44_0, i_13_31_71_0, i_13_31_79_0,
    i_13_31_114_0, i_13_31_138_0, i_13_31_142_0, i_13_31_231_0,
    i_13_31_232_0, i_13_31_411_0, i_13_31_447_0, i_13_31_448_0,
    i_13_31_480_0, i_13_31_537_0, i_13_31_538_0, i_13_31_556_0,
    i_13_31_584_0, i_13_31_589_0, i_13_31_593_0, i_13_31_600_0,
    i_13_31_606_0, i_13_31_609_0, i_13_31_610_0, i_13_31_646_0,
    i_13_31_660_0, i_13_31_673_0, i_13_31_681_0, i_13_31_682_0,
    i_13_31_688_0, i_13_31_760_0, i_13_31_763_0, i_13_31_952_0,
    i_13_31_1119_0, i_13_31_1150_0, i_13_31_1275_0, i_13_31_1308_0,
    i_13_31_1311_0, i_13_31_1312_0, i_13_31_1344_0, i_13_31_1402_0,
    i_13_31_1428_0, i_13_31_1510_0, i_13_31_1626_0, i_13_31_1663_0,
    i_13_31_1672_0, i_13_31_1713_0, i_13_31_1725_0, i_13_31_1726_0,
    i_13_31_1734_0, i_13_31_1780_0, i_13_31_1798_0, i_13_31_1887_0,
    i_13_31_1911_0, i_13_31_1912_0, i_13_31_1923_0, i_13_31_1934_0,
    i_13_31_1947_0, i_13_31_1948_0, i_13_31_2175_0, i_13_31_2321_0,
    i_13_31_2379_0, i_13_31_2552_0, i_13_31_2598_0, i_13_31_2599_0,
    i_13_31_2679_0, i_13_31_2712_0, i_13_31_2752_0, i_13_31_2847_0,
    i_13_31_2850_0, i_13_31_2851_0, i_13_31_2856_0, i_13_31_2877_0,
    i_13_31_2923_0, i_13_31_3046_0, i_13_31_3067_0, i_13_31_3103_0,
    i_13_31_3129_0, i_13_31_3370_0, i_13_31_3371_0, i_13_31_3652_0,
    i_13_31_3668_0, i_13_31_3786_0, i_13_31_3930_0, i_13_31_3931_0,
    i_13_31_3940_0, i_13_31_4154_0, i_13_31_4188_0, i_13_31_4189_0,
    i_13_31_4219_0, i_13_31_4296_0, i_13_31_4297_0, i_13_31_4306_0,
    i_13_31_4308_0, i_13_31_4325_0, i_13_31_4336_0, i_13_31_4435_0,
    i_13_31_4450_0, i_13_31_4539_0, i_13_31_4596_0, i_13_31_4597_0;
  output o_13_31_0_0;
  assign o_13_31_0_0 = ~((i_13_31_593_0 & i_13_31_4306_0 & ~i_13_31_4435_0) | (~i_13_31_1312_0 & ~i_13_31_2851_0 & i_13_31_4154_0 & ~i_13_31_4219_0) | (~i_13_31_79_0 & ~i_13_31_538_0 & ~i_13_31_1311_0 & ~i_13_31_3103_0) | (~i_13_31_447_0 & ~i_13_31_448_0 & ~i_13_31_537_0 & ~i_13_31_1150_0) | (~i_13_31_34_0 & ~i_13_31_231_0 & ~i_13_31_1663_0 & ~i_13_31_1948_0 & ~i_13_31_3652_0 & ~i_13_31_3931_0));
endmodule



// Benchmark "kernel_13_32" written by ABC on Sun Jul 19 10:45:52 2020

module kernel_13_32 ( 
    i_13_32_258_0, i_13_32_259_0, i_13_32_276_0, i_13_32_382_0,
    i_13_32_515_0, i_13_32_516_0, i_13_32_519_0, i_13_32_526_0,
    i_13_32_546_0, i_13_32_551_0, i_13_32_578_0, i_13_32_580_0,
    i_13_32_627_0, i_13_32_640_0, i_13_32_663_0, i_13_32_797_0,
    i_13_32_838_0, i_13_32_843_0, i_13_32_844_0, i_13_32_885_0,
    i_13_32_888_0, i_13_32_932_0, i_13_32_939_0, i_13_32_942_0,
    i_13_32_1077_0, i_13_32_1111_0, i_13_32_1119_0, i_13_32_1149_0,
    i_13_32_1222_0, i_13_32_1224_0, i_13_32_1230_0, i_13_32_1323_0,
    i_13_32_1404_0, i_13_32_1444_0, i_13_32_1464_0, i_13_32_1469_0,
    i_13_32_1483_0, i_13_32_1516_0, i_13_32_1552_0, i_13_32_1660_0,
    i_13_32_1677_0, i_13_32_1732_0, i_13_32_1734_0, i_13_32_1744_0,
    i_13_32_1745_0, i_13_32_1770_0, i_13_32_1830_0, i_13_32_1914_0,
    i_13_32_1915_0, i_13_32_1923_0, i_13_32_1947_0, i_13_32_1959_0,
    i_13_32_2002_0, i_13_32_2004_0, i_13_32_2019_0, i_13_32_2020_0,
    i_13_32_2022_0, i_13_32_2025_0, i_13_32_2197_0, i_13_32_2209_0,
    i_13_32_2320_0, i_13_32_2425_0, i_13_32_2722_0, i_13_32_2742_0,
    i_13_32_2860_0, i_13_32_2898_0, i_13_32_2938_0, i_13_32_2959_0,
    i_13_32_3030_0, i_13_32_3117_0, i_13_32_3156_0, i_13_32_3315_0,
    i_13_32_3351_0, i_13_32_3354_0, i_13_32_3355_0, i_13_32_3412_0,
    i_13_32_3418_0, i_13_32_3478_0, i_13_32_3525_0, i_13_32_3570_0,
    i_13_32_3684_0, i_13_32_3759_0, i_13_32_3763_0, i_13_32_3822_0,
    i_13_32_3864_0, i_13_32_3901_0, i_13_32_4029_0, i_13_32_4054_0,
    i_13_32_4063_0, i_13_32_4124_0, i_13_32_4161_0, i_13_32_4165_0,
    i_13_32_4230_0, i_13_32_4300_0, i_13_32_4303_0, i_13_32_4362_0,
    i_13_32_4567_0, i_13_32_4602_0, i_13_32_4605_0, i_13_32_4606_0,
    o_13_32_0_0  );
  input  i_13_32_258_0, i_13_32_259_0, i_13_32_276_0, i_13_32_382_0,
    i_13_32_515_0, i_13_32_516_0, i_13_32_519_0, i_13_32_526_0,
    i_13_32_546_0, i_13_32_551_0, i_13_32_578_0, i_13_32_580_0,
    i_13_32_627_0, i_13_32_640_0, i_13_32_663_0, i_13_32_797_0,
    i_13_32_838_0, i_13_32_843_0, i_13_32_844_0, i_13_32_885_0,
    i_13_32_888_0, i_13_32_932_0, i_13_32_939_0, i_13_32_942_0,
    i_13_32_1077_0, i_13_32_1111_0, i_13_32_1119_0, i_13_32_1149_0,
    i_13_32_1222_0, i_13_32_1224_0, i_13_32_1230_0, i_13_32_1323_0,
    i_13_32_1404_0, i_13_32_1444_0, i_13_32_1464_0, i_13_32_1469_0,
    i_13_32_1483_0, i_13_32_1516_0, i_13_32_1552_0, i_13_32_1660_0,
    i_13_32_1677_0, i_13_32_1732_0, i_13_32_1734_0, i_13_32_1744_0,
    i_13_32_1745_0, i_13_32_1770_0, i_13_32_1830_0, i_13_32_1914_0,
    i_13_32_1915_0, i_13_32_1923_0, i_13_32_1947_0, i_13_32_1959_0,
    i_13_32_2002_0, i_13_32_2004_0, i_13_32_2019_0, i_13_32_2020_0,
    i_13_32_2022_0, i_13_32_2025_0, i_13_32_2197_0, i_13_32_2209_0,
    i_13_32_2320_0, i_13_32_2425_0, i_13_32_2722_0, i_13_32_2742_0,
    i_13_32_2860_0, i_13_32_2898_0, i_13_32_2938_0, i_13_32_2959_0,
    i_13_32_3030_0, i_13_32_3117_0, i_13_32_3156_0, i_13_32_3315_0,
    i_13_32_3351_0, i_13_32_3354_0, i_13_32_3355_0, i_13_32_3412_0,
    i_13_32_3418_0, i_13_32_3478_0, i_13_32_3525_0, i_13_32_3570_0,
    i_13_32_3684_0, i_13_32_3759_0, i_13_32_3763_0, i_13_32_3822_0,
    i_13_32_3864_0, i_13_32_3901_0, i_13_32_4029_0, i_13_32_4054_0,
    i_13_32_4063_0, i_13_32_4124_0, i_13_32_4161_0, i_13_32_4165_0,
    i_13_32_4230_0, i_13_32_4300_0, i_13_32_4303_0, i_13_32_4362_0,
    i_13_32_4567_0, i_13_32_4602_0, i_13_32_4605_0, i_13_32_4606_0;
  output o_13_32_0_0;
  assign o_13_32_0_0 = ~((~i_13_32_843_0 & ((~i_13_32_516_0 & ~i_13_32_939_0 & ~i_13_32_3684_0 & ~i_13_32_3759_0) | (i_13_32_1552_0 & ~i_13_32_2025_0 & ~i_13_32_2742_0 & ~i_13_32_3822_0))) | (~i_13_32_3315_0 & ((~i_13_32_2019_0 & ~i_13_32_2020_0) | (i_13_32_2938_0 & ~i_13_32_3759_0))) | (~i_13_32_1734_0 & i_13_32_2004_0) | (i_13_32_2002_0 & ~i_13_32_3570_0 & ~i_13_32_4567_0));
endmodule



// Benchmark "kernel_13_33" written by ABC on Sun Jul 19 10:45:53 2020

module kernel_13_33 ( 
    i_13_33_45_0, i_13_33_67_0, i_13_33_117_0, i_13_33_135_0,
    i_13_33_136_0, i_13_33_138_0, i_13_33_192_0, i_13_33_228_0,
    i_13_33_333_0, i_13_33_418_0, i_13_33_534_0, i_13_33_535_0,
    i_13_33_604_0, i_13_33_607_0, i_13_33_612_0, i_13_33_624_0,
    i_13_33_625_0, i_13_33_642_0, i_13_33_643_0, i_13_33_676_0,
    i_13_33_822_0, i_13_33_894_0, i_13_33_976_0, i_13_33_1116_0,
    i_13_33_1119_0, i_13_33_1120_0, i_13_33_1147_0, i_13_33_1272_0,
    i_13_33_1273_0, i_13_33_1390_0, i_13_33_1479_0, i_13_33_1642_0,
    i_13_33_1648_0, i_13_33_1669_0, i_13_33_1777_0, i_13_33_1795_0,
    i_13_33_1885_0, i_13_33_1886_0, i_13_33_1903_0, i_13_33_1944_0,
    i_13_33_1993_0, i_13_33_2230_0, i_13_33_2313_0, i_13_33_2361_0,
    i_13_33_2376_0, i_13_33_2379_0, i_13_33_2380_0, i_13_33_2397_0,
    i_13_33_2400_0, i_13_33_2401_0, i_13_33_2541_0, i_13_33_2578_0,
    i_13_33_2646_0, i_13_33_2647_0, i_13_33_2782_0, i_13_33_2847_0,
    i_13_33_2848_0, i_13_33_2874_0, i_13_33_2878_0, i_13_33_2898_0,
    i_13_33_2899_0, i_13_33_3036_0, i_13_33_3090_0, i_13_33_3091_0,
    i_13_33_3103_0, i_13_33_3117_0, i_13_33_3126_0, i_13_33_3250_0,
    i_13_33_3256_0, i_13_33_3261_0, i_13_33_3262_0, i_13_33_3352_0,
    i_13_33_3367_0, i_13_33_3384_0, i_13_33_3388_0, i_13_33_3508_0,
    i_13_33_3546_0, i_13_33_3547_0, i_13_33_3729_0, i_13_33_3730_0,
    i_13_33_3738_0, i_13_33_3835_0, i_13_33_3889_0, i_13_33_3919_0,
    i_13_33_4018_0, i_13_33_4060_0, i_13_33_4063_0, i_13_33_4185_0,
    i_13_33_4186_0, i_13_33_4209_0, i_13_33_4210_0, i_13_33_4293_0,
    i_13_33_4294_0, i_13_33_4320_0, i_13_33_4351_0, i_13_33_4480_0,
    i_13_33_4500_0, i_13_33_4537_0, i_13_33_4567_0, i_13_33_4594_0,
    o_13_33_0_0  );
  input  i_13_33_45_0, i_13_33_67_0, i_13_33_117_0, i_13_33_135_0,
    i_13_33_136_0, i_13_33_138_0, i_13_33_192_0, i_13_33_228_0,
    i_13_33_333_0, i_13_33_418_0, i_13_33_534_0, i_13_33_535_0,
    i_13_33_604_0, i_13_33_607_0, i_13_33_612_0, i_13_33_624_0,
    i_13_33_625_0, i_13_33_642_0, i_13_33_643_0, i_13_33_676_0,
    i_13_33_822_0, i_13_33_894_0, i_13_33_976_0, i_13_33_1116_0,
    i_13_33_1119_0, i_13_33_1120_0, i_13_33_1147_0, i_13_33_1272_0,
    i_13_33_1273_0, i_13_33_1390_0, i_13_33_1479_0, i_13_33_1642_0,
    i_13_33_1648_0, i_13_33_1669_0, i_13_33_1777_0, i_13_33_1795_0,
    i_13_33_1885_0, i_13_33_1886_0, i_13_33_1903_0, i_13_33_1944_0,
    i_13_33_1993_0, i_13_33_2230_0, i_13_33_2313_0, i_13_33_2361_0,
    i_13_33_2376_0, i_13_33_2379_0, i_13_33_2380_0, i_13_33_2397_0,
    i_13_33_2400_0, i_13_33_2401_0, i_13_33_2541_0, i_13_33_2578_0,
    i_13_33_2646_0, i_13_33_2647_0, i_13_33_2782_0, i_13_33_2847_0,
    i_13_33_2848_0, i_13_33_2874_0, i_13_33_2878_0, i_13_33_2898_0,
    i_13_33_2899_0, i_13_33_3036_0, i_13_33_3090_0, i_13_33_3091_0,
    i_13_33_3103_0, i_13_33_3117_0, i_13_33_3126_0, i_13_33_3250_0,
    i_13_33_3256_0, i_13_33_3261_0, i_13_33_3262_0, i_13_33_3352_0,
    i_13_33_3367_0, i_13_33_3384_0, i_13_33_3388_0, i_13_33_3508_0,
    i_13_33_3546_0, i_13_33_3547_0, i_13_33_3729_0, i_13_33_3730_0,
    i_13_33_3738_0, i_13_33_3835_0, i_13_33_3889_0, i_13_33_3919_0,
    i_13_33_4018_0, i_13_33_4060_0, i_13_33_4063_0, i_13_33_4185_0,
    i_13_33_4186_0, i_13_33_4209_0, i_13_33_4210_0, i_13_33_4293_0,
    i_13_33_4294_0, i_13_33_4320_0, i_13_33_4351_0, i_13_33_4480_0,
    i_13_33_4500_0, i_13_33_4537_0, i_13_33_4567_0, i_13_33_4594_0;
  output o_13_33_0_0;
  assign o_13_33_0_0 = ~(~i_13_33_2848_0 | i_13_33_3103_0 | ~i_13_33_2379_0 | (i_13_33_3919_0 & ~i_13_33_4186_0) | (i_13_33_418_0 & ~i_13_33_4185_0));
endmodule



// Benchmark "kernel_13_34" written by ABC on Sun Jul 19 10:45:54 2020

module kernel_13_34 ( 
    i_13_34_53_0, i_13_34_76_0, i_13_34_121_0, i_13_34_134_0,
    i_13_34_184_0, i_13_34_232_0, i_13_34_251_0, i_13_34_286_0,
    i_13_34_357_0, i_13_34_358_0, i_13_34_359_0, i_13_34_466_0,
    i_13_34_467_0, i_13_34_468_0, i_13_34_592_0, i_13_34_680_0,
    i_13_34_745_0, i_13_34_842_0, i_13_34_916_0, i_13_34_1021_0,
    i_13_34_1025_0, i_13_34_1348_0, i_13_34_1349_0, i_13_34_1400_0,
    i_13_34_1501_0, i_13_34_1507_0, i_13_34_1516_0, i_13_34_1637_0,
    i_13_34_1644_0, i_13_34_1671_0, i_13_34_1727_0, i_13_34_1768_0,
    i_13_34_1816_0, i_13_34_1844_0, i_13_34_1951_0, i_13_34_1952_0,
    i_13_34_1961_0, i_13_34_2032_0, i_13_34_2033_0, i_13_34_2059_0,
    i_13_34_2060_0, i_13_34_2113_0, i_13_34_2203_0, i_13_34_2204_0,
    i_13_34_2284_0, i_13_34_2285_0, i_13_34_2321_0, i_13_34_2382_0,
    i_13_34_2398_0, i_13_34_2399_0, i_13_34_2509_0, i_13_34_2515_0,
    i_13_34_2554_0, i_13_34_2555_0, i_13_34_2570_0, i_13_34_2691_0,
    i_13_34_2752_0, i_13_34_2753_0, i_13_34_2902_0, i_13_34_2923_0,
    i_13_34_2924_0, i_13_34_2959_0, i_13_34_3013_0, i_13_34_3040_0,
    i_13_34_3131_0, i_13_34_3155_0, i_13_34_3163_0, i_13_34_3266_0,
    i_13_34_3373_0, i_13_34_3374_0, i_13_34_3392_0, i_13_34_3419_0,
    i_13_34_3580_0, i_13_34_3581_0, i_13_34_3598_0, i_13_34_3599_0,
    i_13_34_3622_0, i_13_34_3623_0, i_13_34_3634_0, i_13_34_3725_0,
    i_13_34_3787_0, i_13_34_3874_0, i_13_34_3877_0, i_13_34_3915_0,
    i_13_34_3923_0, i_13_34_3968_0, i_13_34_3991_0, i_13_34_3992_0,
    i_13_34_4175_0, i_13_34_4216_0, i_13_34_4256_0, i_13_34_4265_0,
    i_13_34_4316_0, i_13_34_4333_0, i_13_34_4334_0, i_13_34_4433_0,
    i_13_34_4453_0, i_13_34_4454_0, i_13_34_4507_0, i_13_34_4589_0,
    o_13_34_0_0  );
  input  i_13_34_53_0, i_13_34_76_0, i_13_34_121_0, i_13_34_134_0,
    i_13_34_184_0, i_13_34_232_0, i_13_34_251_0, i_13_34_286_0,
    i_13_34_357_0, i_13_34_358_0, i_13_34_359_0, i_13_34_466_0,
    i_13_34_467_0, i_13_34_468_0, i_13_34_592_0, i_13_34_680_0,
    i_13_34_745_0, i_13_34_842_0, i_13_34_916_0, i_13_34_1021_0,
    i_13_34_1025_0, i_13_34_1348_0, i_13_34_1349_0, i_13_34_1400_0,
    i_13_34_1501_0, i_13_34_1507_0, i_13_34_1516_0, i_13_34_1637_0,
    i_13_34_1644_0, i_13_34_1671_0, i_13_34_1727_0, i_13_34_1768_0,
    i_13_34_1816_0, i_13_34_1844_0, i_13_34_1951_0, i_13_34_1952_0,
    i_13_34_1961_0, i_13_34_2032_0, i_13_34_2033_0, i_13_34_2059_0,
    i_13_34_2060_0, i_13_34_2113_0, i_13_34_2203_0, i_13_34_2204_0,
    i_13_34_2284_0, i_13_34_2285_0, i_13_34_2321_0, i_13_34_2382_0,
    i_13_34_2398_0, i_13_34_2399_0, i_13_34_2509_0, i_13_34_2515_0,
    i_13_34_2554_0, i_13_34_2555_0, i_13_34_2570_0, i_13_34_2691_0,
    i_13_34_2752_0, i_13_34_2753_0, i_13_34_2902_0, i_13_34_2923_0,
    i_13_34_2924_0, i_13_34_2959_0, i_13_34_3013_0, i_13_34_3040_0,
    i_13_34_3131_0, i_13_34_3155_0, i_13_34_3163_0, i_13_34_3266_0,
    i_13_34_3373_0, i_13_34_3374_0, i_13_34_3392_0, i_13_34_3419_0,
    i_13_34_3580_0, i_13_34_3581_0, i_13_34_3598_0, i_13_34_3599_0,
    i_13_34_3622_0, i_13_34_3623_0, i_13_34_3634_0, i_13_34_3725_0,
    i_13_34_3787_0, i_13_34_3874_0, i_13_34_3877_0, i_13_34_3915_0,
    i_13_34_3923_0, i_13_34_3968_0, i_13_34_3991_0, i_13_34_3992_0,
    i_13_34_4175_0, i_13_34_4216_0, i_13_34_4256_0, i_13_34_4265_0,
    i_13_34_4316_0, i_13_34_4333_0, i_13_34_4334_0, i_13_34_4433_0,
    i_13_34_4453_0, i_13_34_4454_0, i_13_34_4507_0, i_13_34_4589_0;
  output o_13_34_0_0;
  assign o_13_34_0_0 = ~(~i_13_34_1951_0 & (~i_13_34_466_0 | (~i_13_34_2554_0 & ~i_13_34_4433_0)));
endmodule



// Benchmark "kernel_13_35" written by ABC on Sun Jul 19 10:45:54 2020

module kernel_13_35 ( 
    i_13_35_16_0, i_13_35_43_0, i_13_35_133_0, i_13_35_141_0,
    i_13_35_168_0, i_13_35_186_0, i_13_35_231_0, i_13_35_258_0,
    i_13_35_472_0, i_13_35_531_0, i_13_35_537_0, i_13_35_618_0,
    i_13_35_642_0, i_13_35_643_0, i_13_35_645_0, i_13_35_646_0,
    i_13_35_681_0, i_13_35_688_0, i_13_35_690_0, i_13_35_780_0,
    i_13_35_816_0, i_13_35_817_0, i_13_35_823_0, i_13_35_847_0,
    i_13_35_897_0, i_13_35_979_0, i_13_35_1122_0, i_13_35_1123_0,
    i_13_35_1128_0, i_13_35_1225_0, i_13_35_1275_0, i_13_35_1276_0,
    i_13_35_1464_0, i_13_35_1470_0, i_13_35_1552_0, i_13_35_1600_0,
    i_13_35_1645_0, i_13_35_1723_0, i_13_35_1725_0, i_13_35_1734_0,
    i_13_35_1780_0, i_13_35_1851_0, i_13_35_1887_0, i_13_35_1995_0,
    i_13_35_1996_0, i_13_35_2136_0, i_13_35_2196_0, i_13_35_2262_0,
    i_13_35_2266_0, i_13_35_2379_0, i_13_35_2382_0, i_13_35_2407_0,
    i_13_35_2409_0, i_13_35_2410_0, i_13_35_2422_0, i_13_35_2434_0,
    i_13_35_2542_0, i_13_35_2550_0, i_13_35_2587_0, i_13_35_2616_0,
    i_13_35_2650_0, i_13_35_2653_0, i_13_35_2698_0, i_13_35_2751_0,
    i_13_35_2760_0, i_13_35_2797_0, i_13_35_2877_0, i_13_35_2940_0,
    i_13_35_2941_0, i_13_35_3030_0, i_13_35_3039_0, i_13_35_3067_0,
    i_13_35_3112_0, i_13_35_3291_0, i_13_35_3423_0, i_13_35_3438_0,
    i_13_35_3484_0, i_13_35_3487_0, i_13_35_3526_0, i_13_35_3534_0,
    i_13_35_3724_0, i_13_35_3834_0, i_13_35_3874_0, i_13_35_3921_0,
    i_13_35_3994_0, i_13_35_4015_0, i_13_35_4099_0, i_13_35_4146_0,
    i_13_35_4216_0, i_13_35_4308_0, i_13_35_4309_0, i_13_35_4317_0,
    i_13_35_4318_0, i_13_35_4344_0, i_13_35_4354_0, i_13_35_4375_0,
    i_13_35_4432_0, i_13_35_4554_0, i_13_35_4563_0, i_13_35_4597_0,
    o_13_35_0_0  );
  input  i_13_35_16_0, i_13_35_43_0, i_13_35_133_0, i_13_35_141_0,
    i_13_35_168_0, i_13_35_186_0, i_13_35_231_0, i_13_35_258_0,
    i_13_35_472_0, i_13_35_531_0, i_13_35_537_0, i_13_35_618_0,
    i_13_35_642_0, i_13_35_643_0, i_13_35_645_0, i_13_35_646_0,
    i_13_35_681_0, i_13_35_688_0, i_13_35_690_0, i_13_35_780_0,
    i_13_35_816_0, i_13_35_817_0, i_13_35_823_0, i_13_35_847_0,
    i_13_35_897_0, i_13_35_979_0, i_13_35_1122_0, i_13_35_1123_0,
    i_13_35_1128_0, i_13_35_1225_0, i_13_35_1275_0, i_13_35_1276_0,
    i_13_35_1464_0, i_13_35_1470_0, i_13_35_1552_0, i_13_35_1600_0,
    i_13_35_1645_0, i_13_35_1723_0, i_13_35_1725_0, i_13_35_1734_0,
    i_13_35_1780_0, i_13_35_1851_0, i_13_35_1887_0, i_13_35_1995_0,
    i_13_35_1996_0, i_13_35_2136_0, i_13_35_2196_0, i_13_35_2262_0,
    i_13_35_2266_0, i_13_35_2379_0, i_13_35_2382_0, i_13_35_2407_0,
    i_13_35_2409_0, i_13_35_2410_0, i_13_35_2422_0, i_13_35_2434_0,
    i_13_35_2542_0, i_13_35_2550_0, i_13_35_2587_0, i_13_35_2616_0,
    i_13_35_2650_0, i_13_35_2653_0, i_13_35_2698_0, i_13_35_2751_0,
    i_13_35_2760_0, i_13_35_2797_0, i_13_35_2877_0, i_13_35_2940_0,
    i_13_35_2941_0, i_13_35_3030_0, i_13_35_3039_0, i_13_35_3067_0,
    i_13_35_3112_0, i_13_35_3291_0, i_13_35_3423_0, i_13_35_3438_0,
    i_13_35_3484_0, i_13_35_3487_0, i_13_35_3526_0, i_13_35_3534_0,
    i_13_35_3724_0, i_13_35_3834_0, i_13_35_3874_0, i_13_35_3921_0,
    i_13_35_3994_0, i_13_35_4015_0, i_13_35_4099_0, i_13_35_4146_0,
    i_13_35_4216_0, i_13_35_4308_0, i_13_35_4309_0, i_13_35_4317_0,
    i_13_35_4318_0, i_13_35_4344_0, i_13_35_4354_0, i_13_35_4375_0,
    i_13_35_4432_0, i_13_35_4554_0, i_13_35_4563_0, i_13_35_4597_0;
  output o_13_35_0_0;
  assign o_13_35_0_0 = ~((~i_13_35_897_0 & ((~i_13_35_2698_0 & ~i_13_35_3921_0) | (~i_13_35_1780_0 & ~i_13_35_4317_0))) | (~i_13_35_1734_0 & ~i_13_35_3291_0));
endmodule



// Benchmark "kernel_13_36" written by ABC on Sun Jul 19 10:45:55 2020

module kernel_13_36 ( 
    i_13_36_96_0, i_13_36_105_0, i_13_36_115_0, i_13_36_160_0,
    i_13_36_286_0, i_13_36_453_0, i_13_36_551_0, i_13_36_575_0,
    i_13_36_591_0, i_13_36_592_0, i_13_36_673_0, i_13_36_692_0,
    i_13_36_717_0, i_13_36_832_0, i_13_36_863_0, i_13_36_871_0,
    i_13_36_959_0, i_13_36_1024_0, i_13_36_1084_0, i_13_36_1132_0,
    i_13_36_1150_0, i_13_36_1232_0, i_13_36_1302_0, i_13_36_1303_0,
    i_13_36_1320_0, i_13_36_1464_0, i_13_36_1501_0, i_13_36_1556_0,
    i_13_36_1641_0, i_13_36_1732_0, i_13_36_1754_0, i_13_36_1759_0,
    i_13_36_1768_0, i_13_36_1772_0, i_13_36_1806_0, i_13_36_1807_0,
    i_13_36_1815_0, i_13_36_1816_0, i_13_36_1859_0, i_13_36_1886_0,
    i_13_36_1905_0, i_13_36_1961_0, i_13_36_2059_0, i_13_36_2103_0,
    i_13_36_2123_0, i_13_36_2139_0, i_13_36_2140_0, i_13_36_2141_0,
    i_13_36_2202_0, i_13_36_2284_0, i_13_36_2310_0, i_13_36_2366_0,
    i_13_36_2445_0, i_13_36_2446_0, i_13_36_2470_0, i_13_36_2545_0,
    i_13_36_2617_0, i_13_36_2640_0, i_13_36_2652_0, i_13_36_2654_0,
    i_13_36_2660_0, i_13_36_2663_0, i_13_36_2704_0, i_13_36_2711_0,
    i_13_36_2823_0, i_13_36_2824_0, i_13_36_2858_0, i_13_36_2910_0,
    i_13_36_2941_0, i_13_36_3049_0, i_13_36_3209_0, i_13_36_3219_0,
    i_13_36_3273_0, i_13_36_3374_0, i_13_36_3390_0, i_13_36_3391_0,
    i_13_36_3621_0, i_13_36_3622_0, i_13_36_3633_0, i_13_36_3661_0,
    i_13_36_3740_0, i_13_36_3786_0, i_13_36_3805_0, i_13_36_3868_0,
    i_13_36_3914_0, i_13_36_3991_0, i_13_36_4049_0, i_13_36_4057_0,
    i_13_36_4162_0, i_13_36_4233_0, i_13_36_4236_0, i_13_36_4371_0,
    i_13_36_4372_0, i_13_36_4380_0, i_13_36_4381_0, i_13_36_4382_0,
    i_13_36_4398_0, i_13_36_4399_0, i_13_36_4443_0, i_13_36_4452_0,
    o_13_36_0_0  );
  input  i_13_36_96_0, i_13_36_105_0, i_13_36_115_0, i_13_36_160_0,
    i_13_36_286_0, i_13_36_453_0, i_13_36_551_0, i_13_36_575_0,
    i_13_36_591_0, i_13_36_592_0, i_13_36_673_0, i_13_36_692_0,
    i_13_36_717_0, i_13_36_832_0, i_13_36_863_0, i_13_36_871_0,
    i_13_36_959_0, i_13_36_1024_0, i_13_36_1084_0, i_13_36_1132_0,
    i_13_36_1150_0, i_13_36_1232_0, i_13_36_1302_0, i_13_36_1303_0,
    i_13_36_1320_0, i_13_36_1464_0, i_13_36_1501_0, i_13_36_1556_0,
    i_13_36_1641_0, i_13_36_1732_0, i_13_36_1754_0, i_13_36_1759_0,
    i_13_36_1768_0, i_13_36_1772_0, i_13_36_1806_0, i_13_36_1807_0,
    i_13_36_1815_0, i_13_36_1816_0, i_13_36_1859_0, i_13_36_1886_0,
    i_13_36_1905_0, i_13_36_1961_0, i_13_36_2059_0, i_13_36_2103_0,
    i_13_36_2123_0, i_13_36_2139_0, i_13_36_2140_0, i_13_36_2141_0,
    i_13_36_2202_0, i_13_36_2284_0, i_13_36_2310_0, i_13_36_2366_0,
    i_13_36_2445_0, i_13_36_2446_0, i_13_36_2470_0, i_13_36_2545_0,
    i_13_36_2617_0, i_13_36_2640_0, i_13_36_2652_0, i_13_36_2654_0,
    i_13_36_2660_0, i_13_36_2663_0, i_13_36_2704_0, i_13_36_2711_0,
    i_13_36_2823_0, i_13_36_2824_0, i_13_36_2858_0, i_13_36_2910_0,
    i_13_36_2941_0, i_13_36_3049_0, i_13_36_3209_0, i_13_36_3219_0,
    i_13_36_3273_0, i_13_36_3374_0, i_13_36_3390_0, i_13_36_3391_0,
    i_13_36_3621_0, i_13_36_3622_0, i_13_36_3633_0, i_13_36_3661_0,
    i_13_36_3740_0, i_13_36_3786_0, i_13_36_3805_0, i_13_36_3868_0,
    i_13_36_3914_0, i_13_36_3991_0, i_13_36_4049_0, i_13_36_4057_0,
    i_13_36_4162_0, i_13_36_4233_0, i_13_36_4236_0, i_13_36_4371_0,
    i_13_36_4372_0, i_13_36_4380_0, i_13_36_4381_0, i_13_36_4382_0,
    i_13_36_4398_0, i_13_36_4399_0, i_13_36_4443_0, i_13_36_4452_0;
  output o_13_36_0_0;
  assign o_13_36_0_0 = ~((~i_13_36_105_0 & ((i_13_36_1641_0 & i_13_36_1768_0) | (i_13_36_673_0 & ~i_13_36_1320_0 & ~i_13_36_1859_0 & ~i_13_36_2284_0))) | (~i_13_36_592_0 & i_13_36_832_0 & ~i_13_36_3868_0) | (~i_13_36_1806_0 & ~i_13_36_1807_0 & ~i_13_36_1815_0 & ~i_13_36_3622_0 & ~i_13_36_3914_0) | (i_13_36_1150_0 & ~i_13_36_2059_0 & ~i_13_36_3786_0 & i_13_36_4233_0) | (~i_13_36_1303_0 & ~i_13_36_1641_0 & ~i_13_36_2141_0 & ~i_13_36_2941_0 & ~i_13_36_4452_0));
endmodule



// Benchmark "kernel_13_37" written by ABC on Sun Jul 19 10:45:56 2020

module kernel_13_37 ( 
    i_13_37_30_0, i_13_37_37_0, i_13_37_116_0, i_13_37_120_0,
    i_13_37_126_0, i_13_37_133_0, i_13_37_135_0, i_13_37_136_0,
    i_13_37_324_0, i_13_37_327_0, i_13_37_454_0, i_13_37_487_0,
    i_13_37_544_0, i_13_37_570_0, i_13_37_576_0, i_13_37_594_0,
    i_13_37_595_0, i_13_37_597_0, i_13_37_616_0, i_13_37_684_0,
    i_13_37_714_0, i_13_37_777_0, i_13_37_828_0, i_13_37_891_0,
    i_13_37_910_0, i_13_37_1092_0, i_13_37_1246_0, i_13_37_1296_0,
    i_13_37_1300_0, i_13_37_1306_0, i_13_37_1369_0, i_13_37_1380_0,
    i_13_37_1461_0, i_13_37_1479_0, i_13_37_1480_0, i_13_37_1495_0,
    i_13_37_1552_0, i_13_37_1693_0, i_13_37_1710_0, i_13_37_1723_0,
    i_13_37_1746_0, i_13_37_1756_0, i_13_37_1782_0, i_13_37_1804_0,
    i_13_37_1869_0, i_13_37_1881_0, i_13_37_1903_0, i_13_37_1938_0,
    i_13_37_1939_0, i_13_37_2058_0, i_13_37_2136_0, i_13_37_2289_0,
    i_13_37_2307_0, i_13_37_2316_0, i_13_37_2317_0, i_13_37_2358_0,
    i_13_37_2454_0, i_13_37_2457_0, i_13_37_2458_0, i_13_37_2506_0,
    i_13_37_2596_0, i_13_37_2629_0, i_13_37_2646_0, i_13_37_2649_0,
    i_13_37_2748_0, i_13_37_2755_0, i_13_37_2820_0, i_13_37_2848_0,
    i_13_37_2907_0, i_13_37_2908_0, i_13_37_3010_0, i_13_37_3012_0,
    i_13_37_3013_0, i_13_37_3142_0, i_13_37_3171_0, i_13_37_3205_0,
    i_13_37_3216_0, i_13_37_3217_0, i_13_37_3234_0, i_13_37_3388_0,
    i_13_37_3406_0, i_13_37_3415_0, i_13_37_3429_0, i_13_37_3555_0,
    i_13_37_3556_0, i_13_37_3559_0, i_13_37_3610_0, i_13_37_3790_0,
    i_13_37_3910_0, i_13_37_3918_0, i_13_37_3988_0, i_13_37_4008_0,
    i_13_37_4009_0, i_13_37_4054_0, i_13_37_4078_0, i_13_37_4261_0,
    i_13_37_4263_0, i_13_37_4410_0, i_13_37_4440_0, i_13_37_4584_0,
    o_13_37_0_0  );
  input  i_13_37_30_0, i_13_37_37_0, i_13_37_116_0, i_13_37_120_0,
    i_13_37_126_0, i_13_37_133_0, i_13_37_135_0, i_13_37_136_0,
    i_13_37_324_0, i_13_37_327_0, i_13_37_454_0, i_13_37_487_0,
    i_13_37_544_0, i_13_37_570_0, i_13_37_576_0, i_13_37_594_0,
    i_13_37_595_0, i_13_37_597_0, i_13_37_616_0, i_13_37_684_0,
    i_13_37_714_0, i_13_37_777_0, i_13_37_828_0, i_13_37_891_0,
    i_13_37_910_0, i_13_37_1092_0, i_13_37_1246_0, i_13_37_1296_0,
    i_13_37_1300_0, i_13_37_1306_0, i_13_37_1369_0, i_13_37_1380_0,
    i_13_37_1461_0, i_13_37_1479_0, i_13_37_1480_0, i_13_37_1495_0,
    i_13_37_1552_0, i_13_37_1693_0, i_13_37_1710_0, i_13_37_1723_0,
    i_13_37_1746_0, i_13_37_1756_0, i_13_37_1782_0, i_13_37_1804_0,
    i_13_37_1869_0, i_13_37_1881_0, i_13_37_1903_0, i_13_37_1938_0,
    i_13_37_1939_0, i_13_37_2058_0, i_13_37_2136_0, i_13_37_2289_0,
    i_13_37_2307_0, i_13_37_2316_0, i_13_37_2317_0, i_13_37_2358_0,
    i_13_37_2454_0, i_13_37_2457_0, i_13_37_2458_0, i_13_37_2506_0,
    i_13_37_2596_0, i_13_37_2629_0, i_13_37_2646_0, i_13_37_2649_0,
    i_13_37_2748_0, i_13_37_2755_0, i_13_37_2820_0, i_13_37_2848_0,
    i_13_37_2907_0, i_13_37_2908_0, i_13_37_3010_0, i_13_37_3012_0,
    i_13_37_3013_0, i_13_37_3142_0, i_13_37_3171_0, i_13_37_3205_0,
    i_13_37_3216_0, i_13_37_3217_0, i_13_37_3234_0, i_13_37_3388_0,
    i_13_37_3406_0, i_13_37_3415_0, i_13_37_3429_0, i_13_37_3555_0,
    i_13_37_3556_0, i_13_37_3559_0, i_13_37_3610_0, i_13_37_3790_0,
    i_13_37_3910_0, i_13_37_3918_0, i_13_37_3988_0, i_13_37_4008_0,
    i_13_37_4009_0, i_13_37_4054_0, i_13_37_4078_0, i_13_37_4261_0,
    i_13_37_4263_0, i_13_37_4410_0, i_13_37_4440_0, i_13_37_4584_0;
  output o_13_37_0_0;
  assign o_13_37_0_0 = ~((~i_13_37_4078_0 & (~i_13_37_2848_0 | ~i_13_37_4009_0)) | ~i_13_37_2136_0 | (~i_13_37_891_0 & i_13_37_3610_0));
endmodule



// Benchmark "kernel_13_38" written by ABC on Sun Jul 19 10:45:57 2020

module kernel_13_38 ( 
    i_13_38_52_0, i_13_38_53_0, i_13_38_163_0, i_13_38_170_0,
    i_13_38_175_0, i_13_38_176_0, i_13_38_178_0, i_13_38_179_0,
    i_13_38_188_0, i_13_38_283_0, i_13_38_284_0, i_13_38_286_0,
    i_13_38_287_0, i_13_38_319_0, i_13_38_529_0, i_13_38_572_0,
    i_13_38_574_0, i_13_38_575_0, i_13_38_613_0, i_13_38_692_0,
    i_13_38_718_0, i_13_38_797_0, i_13_38_812_0, i_13_38_826_0,
    i_13_38_827_0, i_13_38_859_0, i_13_38_887_0, i_13_38_955_0,
    i_13_38_1019_0, i_13_38_1067_0, i_13_38_1070_0, i_13_38_1072_0,
    i_13_38_1252_0, i_13_38_1310_0, i_13_38_1313_0, i_13_38_1316_0,
    i_13_38_1447_0, i_13_38_1499_0, i_13_38_1501_0, i_13_38_1502_0,
    i_13_38_1523_0, i_13_38_1634_0, i_13_38_1636_0, i_13_38_1673_0,
    i_13_38_1676_0, i_13_38_1808_0, i_13_38_1849_0, i_13_38_1855_0,
    i_13_38_1861_0, i_13_38_2242_0, i_13_38_2263_0, i_13_38_2297_0,
    i_13_38_2410_0, i_13_38_2411_0, i_13_38_2428_0, i_13_38_2429_0,
    i_13_38_2465_0, i_13_38_2555_0, i_13_38_2612_0, i_13_38_2677_0,
    i_13_38_2681_0, i_13_38_2695_0, i_13_38_3110_0, i_13_38_3113_0,
    i_13_38_3209_0, i_13_38_3245_0, i_13_38_3272_0, i_13_38_3274_0,
    i_13_38_3275_0, i_13_38_3424_0, i_13_38_3425_0, i_13_38_3427_0,
    i_13_38_3428_0, i_13_38_3458_0, i_13_38_3485_0, i_13_38_3731_0,
    i_13_38_3733_0, i_13_38_3734_0, i_13_38_3770_0, i_13_38_3821_0,
    i_13_38_3838_0, i_13_38_3853_0, i_13_38_3854_0, i_13_38_3857_0,
    i_13_38_3875_0, i_13_38_3992_0, i_13_38_4018_0, i_13_38_4019_0,
    i_13_38_4021_0, i_13_38_4022_0, i_13_38_4085_0, i_13_38_4090_0,
    i_13_38_4253_0, i_13_38_4256_0, i_13_38_4264_0, i_13_38_4354_0,
    i_13_38_4510_0, i_13_38_4561_0, i_13_38_4562_0, i_13_38_4598_0,
    o_13_38_0_0  );
  input  i_13_38_52_0, i_13_38_53_0, i_13_38_163_0, i_13_38_170_0,
    i_13_38_175_0, i_13_38_176_0, i_13_38_178_0, i_13_38_179_0,
    i_13_38_188_0, i_13_38_283_0, i_13_38_284_0, i_13_38_286_0,
    i_13_38_287_0, i_13_38_319_0, i_13_38_529_0, i_13_38_572_0,
    i_13_38_574_0, i_13_38_575_0, i_13_38_613_0, i_13_38_692_0,
    i_13_38_718_0, i_13_38_797_0, i_13_38_812_0, i_13_38_826_0,
    i_13_38_827_0, i_13_38_859_0, i_13_38_887_0, i_13_38_955_0,
    i_13_38_1019_0, i_13_38_1067_0, i_13_38_1070_0, i_13_38_1072_0,
    i_13_38_1252_0, i_13_38_1310_0, i_13_38_1313_0, i_13_38_1316_0,
    i_13_38_1447_0, i_13_38_1499_0, i_13_38_1501_0, i_13_38_1502_0,
    i_13_38_1523_0, i_13_38_1634_0, i_13_38_1636_0, i_13_38_1673_0,
    i_13_38_1676_0, i_13_38_1808_0, i_13_38_1849_0, i_13_38_1855_0,
    i_13_38_1861_0, i_13_38_2242_0, i_13_38_2263_0, i_13_38_2297_0,
    i_13_38_2410_0, i_13_38_2411_0, i_13_38_2428_0, i_13_38_2429_0,
    i_13_38_2465_0, i_13_38_2555_0, i_13_38_2612_0, i_13_38_2677_0,
    i_13_38_2681_0, i_13_38_2695_0, i_13_38_3110_0, i_13_38_3113_0,
    i_13_38_3209_0, i_13_38_3245_0, i_13_38_3272_0, i_13_38_3274_0,
    i_13_38_3275_0, i_13_38_3424_0, i_13_38_3425_0, i_13_38_3427_0,
    i_13_38_3428_0, i_13_38_3458_0, i_13_38_3485_0, i_13_38_3731_0,
    i_13_38_3733_0, i_13_38_3734_0, i_13_38_3770_0, i_13_38_3821_0,
    i_13_38_3838_0, i_13_38_3853_0, i_13_38_3854_0, i_13_38_3857_0,
    i_13_38_3875_0, i_13_38_3992_0, i_13_38_4018_0, i_13_38_4019_0,
    i_13_38_4021_0, i_13_38_4022_0, i_13_38_4085_0, i_13_38_4090_0,
    i_13_38_4253_0, i_13_38_4256_0, i_13_38_4264_0, i_13_38_4354_0,
    i_13_38_4510_0, i_13_38_4561_0, i_13_38_4562_0, i_13_38_4598_0;
  output o_13_38_0_0;
  assign o_13_38_0_0 = ~((~i_13_38_1070_0 & ((~i_13_38_284_0 & ~i_13_38_574_0 & ~i_13_38_2465_0 & ~i_13_38_3821_0) | (~i_13_38_2429_0 & ~i_13_38_4256_0 & ~i_13_38_4562_0))) | (~i_13_38_1310_0 & ~i_13_38_2681_0 & ~i_13_38_2695_0 & ~i_13_38_3113_0) | (~i_13_38_178_0 & ~i_13_38_3733_0 & ~i_13_38_3734_0) | (~i_13_38_179_0 & ~i_13_38_3209_0 & ~i_13_38_4090_0));
endmodule



// Benchmark "kernel_13_39" written by ABC on Sun Jul 19 10:45:58 2020

module kernel_13_39 ( 
    i_13_39_62_0, i_13_39_76_0, i_13_39_77_0, i_13_39_326_0, i_13_39_416_0,
    i_13_39_562_0, i_13_39_571_0, i_13_39_622_0, i_13_39_688_0,
    i_13_39_697_0, i_13_39_707_0, i_13_39_719_0, i_13_39_827_0,
    i_13_39_841_0, i_13_39_863_0, i_13_39_925_0, i_13_39_938_0,
    i_13_39_958_0, i_13_39_1022_0, i_13_39_1072_0, i_13_39_1073_0,
    i_13_39_1077_0, i_13_39_1219_0, i_13_39_1225_0, i_13_39_1228_0,
    i_13_39_1256_0, i_13_39_1259_0, i_13_39_1262_0, i_13_39_1280_0,
    i_13_39_1300_0, i_13_39_1315_0, i_13_39_1318_0, i_13_39_1319_0,
    i_13_39_1444_0, i_13_39_1445_0, i_13_39_1465_0, i_13_39_1553_0,
    i_13_39_1589_0, i_13_39_1606_0, i_13_39_1679_0, i_13_39_1774_0,
    i_13_39_1775_0, i_13_39_1778_0, i_13_39_1855_0, i_13_39_1858_0,
    i_13_39_1859_0, i_13_39_1914_0, i_13_39_1922_0, i_13_39_1982_0,
    i_13_39_1989_0, i_13_39_2000_0, i_13_39_2002_0, i_13_39_2056_0,
    i_13_39_2159_0, i_13_39_2173_0, i_13_39_2270_0, i_13_39_2461_0,
    i_13_39_2540_0, i_13_39_2630_0, i_13_39_2657_0, i_13_39_2677_0,
    i_13_39_2705_0, i_13_39_2774_0, i_13_39_2858_0, i_13_39_3010_0,
    i_13_39_3064_0, i_13_39_3091_0, i_13_39_3145_0, i_13_39_3173_0,
    i_13_39_3269_0, i_13_39_3308_0, i_13_39_3416_0, i_13_39_3449_0,
    i_13_39_3484_0, i_13_39_3487_0, i_13_39_3507_0, i_13_39_3541_0,
    i_13_39_3542_0, i_13_39_3544_0, i_13_39_3578_0, i_13_39_3634_0,
    i_13_39_3761_0, i_13_39_3803_0, i_13_39_3814_0, i_13_39_3863_0,
    i_13_39_4013_0, i_13_39_4018_0, i_13_39_4054_0, i_13_39_4253_0,
    i_13_39_4279_0, i_13_39_4333_0, i_13_39_4351_0, i_13_39_4370_0,
    i_13_39_4372_0, i_13_39_4376_0, i_13_39_4378_0, i_13_39_4379_0,
    i_13_39_4519_0, i_13_39_4520_0, i_13_39_4567_0,
    o_13_39_0_0  );
  input  i_13_39_62_0, i_13_39_76_0, i_13_39_77_0, i_13_39_326_0,
    i_13_39_416_0, i_13_39_562_0, i_13_39_571_0, i_13_39_622_0,
    i_13_39_688_0, i_13_39_697_0, i_13_39_707_0, i_13_39_719_0,
    i_13_39_827_0, i_13_39_841_0, i_13_39_863_0, i_13_39_925_0,
    i_13_39_938_0, i_13_39_958_0, i_13_39_1022_0, i_13_39_1072_0,
    i_13_39_1073_0, i_13_39_1077_0, i_13_39_1219_0, i_13_39_1225_0,
    i_13_39_1228_0, i_13_39_1256_0, i_13_39_1259_0, i_13_39_1262_0,
    i_13_39_1280_0, i_13_39_1300_0, i_13_39_1315_0, i_13_39_1318_0,
    i_13_39_1319_0, i_13_39_1444_0, i_13_39_1445_0, i_13_39_1465_0,
    i_13_39_1553_0, i_13_39_1589_0, i_13_39_1606_0, i_13_39_1679_0,
    i_13_39_1774_0, i_13_39_1775_0, i_13_39_1778_0, i_13_39_1855_0,
    i_13_39_1858_0, i_13_39_1859_0, i_13_39_1914_0, i_13_39_1922_0,
    i_13_39_1982_0, i_13_39_1989_0, i_13_39_2000_0, i_13_39_2002_0,
    i_13_39_2056_0, i_13_39_2159_0, i_13_39_2173_0, i_13_39_2270_0,
    i_13_39_2461_0, i_13_39_2540_0, i_13_39_2630_0, i_13_39_2657_0,
    i_13_39_2677_0, i_13_39_2705_0, i_13_39_2774_0, i_13_39_2858_0,
    i_13_39_3010_0, i_13_39_3064_0, i_13_39_3091_0, i_13_39_3145_0,
    i_13_39_3173_0, i_13_39_3269_0, i_13_39_3308_0, i_13_39_3416_0,
    i_13_39_3449_0, i_13_39_3484_0, i_13_39_3487_0, i_13_39_3507_0,
    i_13_39_3541_0, i_13_39_3542_0, i_13_39_3544_0, i_13_39_3578_0,
    i_13_39_3634_0, i_13_39_3761_0, i_13_39_3803_0, i_13_39_3814_0,
    i_13_39_3863_0, i_13_39_4013_0, i_13_39_4018_0, i_13_39_4054_0,
    i_13_39_4253_0, i_13_39_4279_0, i_13_39_4333_0, i_13_39_4351_0,
    i_13_39_4370_0, i_13_39_4372_0, i_13_39_4376_0, i_13_39_4378_0,
    i_13_39_4379_0, i_13_39_4519_0, i_13_39_4520_0, i_13_39_4567_0;
  output o_13_39_0_0;
  assign o_13_39_0_0 = ~((~i_13_39_1259_0 & ((~i_13_39_76_0 & i_13_39_841_0 & ~i_13_39_1315_0 & ~i_13_39_1858_0) | (~i_13_39_1300_0 & ~i_13_39_2540_0 & ~i_13_39_3761_0 & ~i_13_39_4054_0 & ~i_13_39_4333_0))) | (~i_13_39_2000_0 & ((i_13_39_562_0 & ~i_13_39_1219_0 & ~i_13_39_3010_0) | (~i_13_39_2540_0 & ~i_13_39_3173_0 & ~i_13_39_3484_0 & ~i_13_39_3541_0 & ~i_13_39_4567_0))) | ~i_13_39_1319_0 | (~i_13_39_1022_0 & ~i_13_39_1315_0 & ~i_13_39_1775_0));
endmodule



// Benchmark "kernel_13_40" written by ABC on Sun Jul 19 10:45:58 2020

module kernel_13_40 ( 
    i_13_40_31_0, i_13_40_44_0, i_13_40_77_0, i_13_40_103_0, i_13_40_275_0,
    i_13_40_469_0, i_13_40_497_0, i_13_40_527_0, i_13_40_557_0,
    i_13_40_562_0, i_13_40_563_0, i_13_40_611_0, i_13_40_664_0,
    i_13_40_827_0, i_13_40_941_0, i_13_40_953_0, i_13_40_1021_0,
    i_13_40_1022_0, i_13_40_1025_0, i_13_40_1060_0, i_13_40_1075_0,
    i_13_40_1076_0, i_13_40_1139_0, i_13_40_1151_0, i_13_40_1256_0,
    i_13_40_1259_0, i_13_40_1270_0, i_13_40_1313_0, i_13_40_1318_0,
    i_13_40_1319_0, i_13_40_1333_0, i_13_40_1339_0, i_13_40_1372_0,
    i_13_40_1377_0, i_13_40_1553_0, i_13_40_1634_0, i_13_40_1691_0,
    i_13_40_1717_0, i_13_40_1723_0, i_13_40_1786_0, i_13_40_1804_0,
    i_13_40_1858_0, i_13_40_1861_0, i_13_40_1862_0, i_13_40_1942_0,
    i_13_40_1958_0, i_13_40_2026_0, i_13_40_2158_0, i_13_40_2197_0,
    i_13_40_2455_0, i_13_40_2476_0, i_13_40_2552_0, i_13_40_2618_0,
    i_13_40_2702_0, i_13_40_2744_0, i_13_40_2750_0, i_13_40_2921_0,
    i_13_40_2966_0, i_13_40_3010_0, i_13_40_3011_0, i_13_40_3014_0,
    i_13_40_3037_0, i_13_40_3163_0, i_13_40_3173_0, i_13_40_3226_0,
    i_13_40_3235_0, i_13_40_3245_0, i_13_40_3272_0, i_13_40_3443_0,
    i_13_40_3461_0, i_13_40_3479_0, i_13_40_3482_0, i_13_40_3487_0,
    i_13_40_3488_0, i_13_40_3491_0, i_13_40_3541_0, i_13_40_3542_0,
    i_13_40_3569_0, i_13_40_3571_0, i_13_40_3572_0, i_13_40_3574_0,
    i_13_40_3577_0, i_13_40_3578_0, i_13_40_3784_0, i_13_40_3785_0,
    i_13_40_3859_0, i_13_40_3895_0, i_13_40_3911_0, i_13_40_3960_0,
    i_13_40_4252_0, i_13_40_4253_0, i_13_40_4256_0, i_13_40_4258_0,
    i_13_40_4261_0, i_13_40_4262_0, i_13_40_4351_0, i_13_40_4372_0,
    i_13_40_4378_0, i_13_40_4447_0, i_13_40_4567_0,
    o_13_40_0_0  );
  input  i_13_40_31_0, i_13_40_44_0, i_13_40_77_0, i_13_40_103_0,
    i_13_40_275_0, i_13_40_469_0, i_13_40_497_0, i_13_40_527_0,
    i_13_40_557_0, i_13_40_562_0, i_13_40_563_0, i_13_40_611_0,
    i_13_40_664_0, i_13_40_827_0, i_13_40_941_0, i_13_40_953_0,
    i_13_40_1021_0, i_13_40_1022_0, i_13_40_1025_0, i_13_40_1060_0,
    i_13_40_1075_0, i_13_40_1076_0, i_13_40_1139_0, i_13_40_1151_0,
    i_13_40_1256_0, i_13_40_1259_0, i_13_40_1270_0, i_13_40_1313_0,
    i_13_40_1318_0, i_13_40_1319_0, i_13_40_1333_0, i_13_40_1339_0,
    i_13_40_1372_0, i_13_40_1377_0, i_13_40_1553_0, i_13_40_1634_0,
    i_13_40_1691_0, i_13_40_1717_0, i_13_40_1723_0, i_13_40_1786_0,
    i_13_40_1804_0, i_13_40_1858_0, i_13_40_1861_0, i_13_40_1862_0,
    i_13_40_1942_0, i_13_40_1958_0, i_13_40_2026_0, i_13_40_2158_0,
    i_13_40_2197_0, i_13_40_2455_0, i_13_40_2476_0, i_13_40_2552_0,
    i_13_40_2618_0, i_13_40_2702_0, i_13_40_2744_0, i_13_40_2750_0,
    i_13_40_2921_0, i_13_40_2966_0, i_13_40_3010_0, i_13_40_3011_0,
    i_13_40_3014_0, i_13_40_3037_0, i_13_40_3163_0, i_13_40_3173_0,
    i_13_40_3226_0, i_13_40_3235_0, i_13_40_3245_0, i_13_40_3272_0,
    i_13_40_3443_0, i_13_40_3461_0, i_13_40_3479_0, i_13_40_3482_0,
    i_13_40_3487_0, i_13_40_3488_0, i_13_40_3491_0, i_13_40_3541_0,
    i_13_40_3542_0, i_13_40_3569_0, i_13_40_3571_0, i_13_40_3572_0,
    i_13_40_3574_0, i_13_40_3577_0, i_13_40_3578_0, i_13_40_3784_0,
    i_13_40_3785_0, i_13_40_3859_0, i_13_40_3895_0, i_13_40_3911_0,
    i_13_40_3960_0, i_13_40_4252_0, i_13_40_4253_0, i_13_40_4256_0,
    i_13_40_4258_0, i_13_40_4261_0, i_13_40_4262_0, i_13_40_4351_0,
    i_13_40_4372_0, i_13_40_4378_0, i_13_40_4447_0, i_13_40_4567_0;
  output o_13_40_0_0;
  assign o_13_40_0_0 = ~(i_13_40_1270_0 | ~i_13_40_3542_0 | (~i_13_40_1858_0 & ~i_13_40_4372_0) | (~i_13_40_2744_0 & ~i_13_40_3578_0 & ~i_13_40_4378_0));
endmodule



// Benchmark "kernel_13_41" written by ABC on Sun Jul 19 10:46:00 2020

module kernel_13_41 ( 
    i_13_41_27_0, i_13_41_105_0, i_13_41_183_0, i_13_41_185_0,
    i_13_41_186_0, i_13_41_187_0, i_13_41_205_0, i_13_41_229_0,
    i_13_41_256_0, i_13_41_376_0, i_13_41_382_0, i_13_41_388_0,
    i_13_41_439_0, i_13_41_526_0, i_13_41_550_0, i_13_41_589_0,
    i_13_41_600_0, i_13_41_610_0, i_13_41_624_0, i_13_41_625_0,
    i_13_41_658_0, i_13_41_669_0, i_13_41_673_0, i_13_41_676_0,
    i_13_41_681_0, i_13_41_765_0, i_13_41_796_0, i_13_41_887_0,
    i_13_41_1111_0, i_13_41_1123_0, i_13_41_1144_0, i_13_41_1150_0,
    i_13_41_1195_0, i_13_41_1201_0, i_13_41_1270_0, i_13_41_1326_0,
    i_13_41_1327_0, i_13_41_1363_0, i_13_41_1404_0, i_13_41_1497_0,
    i_13_41_1503_0, i_13_41_1515_0, i_13_41_1516_0, i_13_41_1653_0,
    i_13_41_1677_0, i_13_41_1678_0, i_13_41_1680_0, i_13_41_1714_0,
    i_13_41_1729_0, i_13_41_1733_0, i_13_41_1741_0, i_13_41_1834_0,
    i_13_41_1839_0, i_13_41_1857_0, i_13_41_1860_0, i_13_41_1909_0,
    i_13_41_1911_0, i_13_41_1912_0, i_13_41_1999_0, i_13_41_2001_0,
    i_13_41_2002_0, i_13_41_2020_0, i_13_41_2175_0, i_13_41_2176_0,
    i_13_41_2200_0, i_13_41_2363_0, i_13_41_2556_0, i_13_41_2616_0,
    i_13_41_2722_0, i_13_41_2727_0, i_13_41_2760_0, i_13_41_2793_0,
    i_13_41_2857_0, i_13_41_2860_0, i_13_41_2973_0, i_13_41_3000_0,
    i_13_41_3028_0, i_13_41_3087_0, i_13_41_3090_0, i_13_41_3121_0,
    i_13_41_3382_0, i_13_41_3460_0, i_13_41_3522_0, i_13_41_3546_0,
    i_13_41_3552_0, i_13_41_3685_0, i_13_41_3730_0, i_13_41_3766_0,
    i_13_41_3864_0, i_13_41_3925_0, i_13_41_4054_0, i_13_41_4080_0,
    i_13_41_4186_0, i_13_41_4200_0, i_13_41_4393_0, i_13_41_4480_0,
    i_13_41_4567_0, i_13_41_4581_0, i_13_41_4600_0, i_13_41_4602_0,
    o_13_41_0_0  );
  input  i_13_41_27_0, i_13_41_105_0, i_13_41_183_0, i_13_41_185_0,
    i_13_41_186_0, i_13_41_187_0, i_13_41_205_0, i_13_41_229_0,
    i_13_41_256_0, i_13_41_376_0, i_13_41_382_0, i_13_41_388_0,
    i_13_41_439_0, i_13_41_526_0, i_13_41_550_0, i_13_41_589_0,
    i_13_41_600_0, i_13_41_610_0, i_13_41_624_0, i_13_41_625_0,
    i_13_41_658_0, i_13_41_669_0, i_13_41_673_0, i_13_41_676_0,
    i_13_41_681_0, i_13_41_765_0, i_13_41_796_0, i_13_41_887_0,
    i_13_41_1111_0, i_13_41_1123_0, i_13_41_1144_0, i_13_41_1150_0,
    i_13_41_1195_0, i_13_41_1201_0, i_13_41_1270_0, i_13_41_1326_0,
    i_13_41_1327_0, i_13_41_1363_0, i_13_41_1404_0, i_13_41_1497_0,
    i_13_41_1503_0, i_13_41_1515_0, i_13_41_1516_0, i_13_41_1653_0,
    i_13_41_1677_0, i_13_41_1678_0, i_13_41_1680_0, i_13_41_1714_0,
    i_13_41_1729_0, i_13_41_1733_0, i_13_41_1741_0, i_13_41_1834_0,
    i_13_41_1839_0, i_13_41_1857_0, i_13_41_1860_0, i_13_41_1909_0,
    i_13_41_1911_0, i_13_41_1912_0, i_13_41_1999_0, i_13_41_2001_0,
    i_13_41_2002_0, i_13_41_2020_0, i_13_41_2175_0, i_13_41_2176_0,
    i_13_41_2200_0, i_13_41_2363_0, i_13_41_2556_0, i_13_41_2616_0,
    i_13_41_2722_0, i_13_41_2727_0, i_13_41_2760_0, i_13_41_2793_0,
    i_13_41_2857_0, i_13_41_2860_0, i_13_41_2973_0, i_13_41_3000_0,
    i_13_41_3028_0, i_13_41_3087_0, i_13_41_3090_0, i_13_41_3121_0,
    i_13_41_3382_0, i_13_41_3460_0, i_13_41_3522_0, i_13_41_3546_0,
    i_13_41_3552_0, i_13_41_3685_0, i_13_41_3730_0, i_13_41_3766_0,
    i_13_41_3864_0, i_13_41_3925_0, i_13_41_4054_0, i_13_41_4080_0,
    i_13_41_4186_0, i_13_41_4200_0, i_13_41_4393_0, i_13_41_4480_0,
    i_13_41_4567_0, i_13_41_4581_0, i_13_41_4600_0, i_13_41_4602_0;
  output o_13_41_0_0;
  assign o_13_41_0_0 = ~(~i_13_41_3864_0 | (i_13_41_673_0 & ~i_13_41_4567_0) | (~i_13_41_3522_0 & ~i_13_41_4080_0) | (i_13_41_526_0 & i_13_41_3685_0) | (~i_13_41_187_0 & ~i_13_41_1326_0));
endmodule



// Benchmark "kernel_13_42" written by ABC on Sun Jul 19 10:46:00 2020

module kernel_13_42 ( 
    i_13_42_40_0, i_13_42_90_0, i_13_42_129_0, i_13_42_130_0,
    i_13_42_156_0, i_13_42_190_0, i_13_42_270_0, i_13_42_273_0,
    i_13_42_336_0, i_13_42_418_0, i_13_42_453_0, i_13_42_468_0,
    i_13_42_490_0, i_13_42_526_0, i_13_42_558_0, i_13_42_561_0,
    i_13_42_562_0, i_13_42_633_0, i_13_42_657_0, i_13_42_724_0,
    i_13_42_732_0, i_13_42_742_0, i_13_42_823_0, i_13_42_838_0,
    i_13_42_945_0, i_13_42_1083_0, i_13_42_1084_0, i_13_42_1143_0,
    i_13_42_1147_0, i_13_42_1242_0, i_13_42_1350_0, i_13_42_1470_0,
    i_13_42_1620_0, i_13_42_1650_0, i_13_42_1768_0, i_13_42_1785_0,
    i_13_42_1812_0, i_13_42_1840_0, i_13_42_1857_0, i_13_42_1936_0,
    i_13_42_2001_0, i_13_42_2205_0, i_13_42_2430_0, i_13_42_2497_0,
    i_13_42_2529_0, i_13_42_2546_0, i_13_42_2649_0, i_13_42_2650_0,
    i_13_42_2664_0, i_13_42_2709_0, i_13_42_2784_0, i_13_42_2982_0,
    i_13_42_3019_0, i_13_42_3043_0, i_13_42_3046_0, i_13_42_3070_0,
    i_13_42_3097_0, i_13_42_3099_0, i_13_42_3100_0, i_13_42_3135_0,
    i_13_42_3141_0, i_13_42_3213_0, i_13_42_3231_0, i_13_42_3234_0,
    i_13_42_3252_0, i_13_42_3351_0, i_13_42_3388_0, i_13_42_3415_0,
    i_13_42_3487_0, i_13_42_3541_0, i_13_42_3549_0, i_13_42_3603_0,
    i_13_42_3636_0, i_13_42_3640_0, i_13_42_3655_0, i_13_42_3682_0,
    i_13_42_3685_0, i_13_42_3699_0, i_13_42_3730_0, i_13_42_3747_0,
    i_13_42_3762_0, i_13_42_3870_0, i_13_42_3897_0, i_13_42_3909_0,
    i_13_42_3979_0, i_13_42_3981_0, i_13_42_3982_0, i_13_42_4158_0,
    i_13_42_4159_0, i_13_42_4161_0, i_13_42_4162_0, i_13_42_4164_0,
    i_13_42_4177_0, i_13_42_4194_0, i_13_42_4195_0, i_13_42_4269_0,
    i_13_42_4321_0, i_13_42_4324_0, i_13_42_4428_0, i_13_42_4539_0,
    o_13_42_0_0  );
  input  i_13_42_40_0, i_13_42_90_0, i_13_42_129_0, i_13_42_130_0,
    i_13_42_156_0, i_13_42_190_0, i_13_42_270_0, i_13_42_273_0,
    i_13_42_336_0, i_13_42_418_0, i_13_42_453_0, i_13_42_468_0,
    i_13_42_490_0, i_13_42_526_0, i_13_42_558_0, i_13_42_561_0,
    i_13_42_562_0, i_13_42_633_0, i_13_42_657_0, i_13_42_724_0,
    i_13_42_732_0, i_13_42_742_0, i_13_42_823_0, i_13_42_838_0,
    i_13_42_945_0, i_13_42_1083_0, i_13_42_1084_0, i_13_42_1143_0,
    i_13_42_1147_0, i_13_42_1242_0, i_13_42_1350_0, i_13_42_1470_0,
    i_13_42_1620_0, i_13_42_1650_0, i_13_42_1768_0, i_13_42_1785_0,
    i_13_42_1812_0, i_13_42_1840_0, i_13_42_1857_0, i_13_42_1936_0,
    i_13_42_2001_0, i_13_42_2205_0, i_13_42_2430_0, i_13_42_2497_0,
    i_13_42_2529_0, i_13_42_2546_0, i_13_42_2649_0, i_13_42_2650_0,
    i_13_42_2664_0, i_13_42_2709_0, i_13_42_2784_0, i_13_42_2982_0,
    i_13_42_3019_0, i_13_42_3043_0, i_13_42_3046_0, i_13_42_3070_0,
    i_13_42_3097_0, i_13_42_3099_0, i_13_42_3100_0, i_13_42_3135_0,
    i_13_42_3141_0, i_13_42_3213_0, i_13_42_3231_0, i_13_42_3234_0,
    i_13_42_3252_0, i_13_42_3351_0, i_13_42_3388_0, i_13_42_3415_0,
    i_13_42_3487_0, i_13_42_3541_0, i_13_42_3549_0, i_13_42_3603_0,
    i_13_42_3636_0, i_13_42_3640_0, i_13_42_3655_0, i_13_42_3682_0,
    i_13_42_3685_0, i_13_42_3699_0, i_13_42_3730_0, i_13_42_3747_0,
    i_13_42_3762_0, i_13_42_3870_0, i_13_42_3897_0, i_13_42_3909_0,
    i_13_42_3979_0, i_13_42_3981_0, i_13_42_3982_0, i_13_42_4158_0,
    i_13_42_4159_0, i_13_42_4161_0, i_13_42_4162_0, i_13_42_4164_0,
    i_13_42_4177_0, i_13_42_4194_0, i_13_42_4195_0, i_13_42_4269_0,
    i_13_42_4321_0, i_13_42_4324_0, i_13_42_4428_0, i_13_42_4539_0;
  output o_13_42_0_0;
  assign o_13_42_0_0 = ~((~i_13_42_1084_0 & (~i_13_42_3549_0 | (i_13_42_823_0 & ~i_13_42_4159_0))) | (~i_13_42_3099_0 & ((~i_13_42_561_0 & ~i_13_42_1147_0) | (~i_13_42_1768_0 & ~i_13_42_3100_0 & i_13_42_3603_0) | (~i_13_42_270_0 & ~i_13_42_2529_0 & ~i_13_42_2982_0 & ~i_13_42_4164_0))) | (i_13_42_3909_0 & ~i_13_42_3981_0 & ~i_13_42_4269_0) | (~i_13_42_562_0 & ~i_13_42_3897_0 & ~i_13_42_4324_0));
endmodule



// Benchmark "kernel_13_43" written by ABC on Sun Jul 19 10:46:01 2020

module kernel_13_43 ( 
    i_13_43_31_0, i_13_43_49_0, i_13_43_63_0, i_13_43_66_0, i_13_43_67_0,
    i_13_43_136_0, i_13_43_140_0, i_13_43_211_0, i_13_43_227_0,
    i_13_43_228_0, i_13_43_285_0, i_13_43_409_0, i_13_43_447_0,
    i_13_43_490_0, i_13_43_537_0, i_13_43_609_0, i_13_43_612_0,
    i_13_43_614_0, i_13_43_645_0, i_13_43_649_0, i_13_43_672_0,
    i_13_43_684_0, i_13_43_686_0, i_13_43_699_0, i_13_43_771_0,
    i_13_43_814_0, i_13_43_820_0, i_13_43_982_0, i_13_43_1066_0,
    i_13_43_1116_0, i_13_43_1117_0, i_13_43_1118_0, i_13_43_1119_0,
    i_13_43_1225_0, i_13_43_1226_0, i_13_43_1270_0, i_13_43_1274_0,
    i_13_43_1307_0, i_13_43_1327_0, i_13_43_1388_0, i_13_43_1411_0,
    i_13_43_1427_0, i_13_43_1489_0, i_13_43_1513_0, i_13_43_1539_0,
    i_13_43_1570_0, i_13_43_1639_0, i_13_43_1672_0, i_13_43_1723_0,
    i_13_43_1732_0, i_13_43_1793_0, i_13_43_1795_0, i_13_43_1801_0,
    i_13_43_1849_0, i_13_43_1885_0, i_13_43_1909_0, i_13_43_2056_0,
    i_13_43_2128_0, i_13_43_2135_0, i_13_43_2297_0, i_13_43_2407_0,
    i_13_43_2408_0, i_13_43_2423_0, i_13_43_2433_0, i_13_43_2434_0,
    i_13_43_2635_0, i_13_43_2719_0, i_13_43_2722_0, i_13_43_2847_0,
    i_13_43_2848_0, i_13_43_2850_0, i_13_43_2875_0, i_13_43_3037_0,
    i_13_43_3093_0, i_13_43_3165_0, i_13_43_3268_0, i_13_43_3387_0,
    i_13_43_3400_0, i_13_43_3520_0, i_13_43_3537_0, i_13_43_3539_0,
    i_13_43_3577_0, i_13_43_3741_0, i_13_43_3766_0, i_13_43_3793_0,
    i_13_43_3836_0, i_13_43_3837_0, i_13_43_3894_0, i_13_43_3924_0,
    i_13_43_3965_0, i_13_43_4033_0, i_13_43_4043_0, i_13_43_4053_0,
    i_13_43_4078_0, i_13_43_4216_0, i_13_43_4294_0, i_13_43_4295_0,
    i_13_43_4296_0, i_13_43_4297_0, i_13_43_4376_0,
    o_13_43_0_0  );
  input  i_13_43_31_0, i_13_43_49_0, i_13_43_63_0, i_13_43_66_0,
    i_13_43_67_0, i_13_43_136_0, i_13_43_140_0, i_13_43_211_0,
    i_13_43_227_0, i_13_43_228_0, i_13_43_285_0, i_13_43_409_0,
    i_13_43_447_0, i_13_43_490_0, i_13_43_537_0, i_13_43_609_0,
    i_13_43_612_0, i_13_43_614_0, i_13_43_645_0, i_13_43_649_0,
    i_13_43_672_0, i_13_43_684_0, i_13_43_686_0, i_13_43_699_0,
    i_13_43_771_0, i_13_43_814_0, i_13_43_820_0, i_13_43_982_0,
    i_13_43_1066_0, i_13_43_1116_0, i_13_43_1117_0, i_13_43_1118_0,
    i_13_43_1119_0, i_13_43_1225_0, i_13_43_1226_0, i_13_43_1270_0,
    i_13_43_1274_0, i_13_43_1307_0, i_13_43_1327_0, i_13_43_1388_0,
    i_13_43_1411_0, i_13_43_1427_0, i_13_43_1489_0, i_13_43_1513_0,
    i_13_43_1539_0, i_13_43_1570_0, i_13_43_1639_0, i_13_43_1672_0,
    i_13_43_1723_0, i_13_43_1732_0, i_13_43_1793_0, i_13_43_1795_0,
    i_13_43_1801_0, i_13_43_1849_0, i_13_43_1885_0, i_13_43_1909_0,
    i_13_43_2056_0, i_13_43_2128_0, i_13_43_2135_0, i_13_43_2297_0,
    i_13_43_2407_0, i_13_43_2408_0, i_13_43_2423_0, i_13_43_2433_0,
    i_13_43_2434_0, i_13_43_2635_0, i_13_43_2719_0, i_13_43_2722_0,
    i_13_43_2847_0, i_13_43_2848_0, i_13_43_2850_0, i_13_43_2875_0,
    i_13_43_3037_0, i_13_43_3093_0, i_13_43_3165_0, i_13_43_3268_0,
    i_13_43_3387_0, i_13_43_3400_0, i_13_43_3520_0, i_13_43_3537_0,
    i_13_43_3539_0, i_13_43_3577_0, i_13_43_3741_0, i_13_43_3766_0,
    i_13_43_3793_0, i_13_43_3836_0, i_13_43_3837_0, i_13_43_3894_0,
    i_13_43_3924_0, i_13_43_3965_0, i_13_43_4033_0, i_13_43_4043_0,
    i_13_43_4053_0, i_13_43_4078_0, i_13_43_4216_0, i_13_43_4294_0,
    i_13_43_4295_0, i_13_43_4296_0, i_13_43_4297_0, i_13_43_4376_0;
  output o_13_43_0_0;
  assign o_13_43_0_0 = ~((~i_13_43_4078_0 & ((~i_13_43_537_0 & ~i_13_43_1793_0 & ~i_13_43_2848_0 & ~i_13_43_3924_0) | (~i_13_43_31_0 & ~i_13_43_67_0 & i_13_43_2434_0 & ~i_13_43_2847_0 & i_13_43_4216_0))) | (i_13_43_63_0 & ~i_13_43_66_0 & i_13_43_67_0 & ~i_13_43_1801_0) | (i_13_43_1795_0 & i_13_43_2408_0) | (~i_13_43_820_0 & ~i_13_43_1489_0 & ~i_13_43_1795_0 & ~i_13_43_2433_0) | (i_13_43_490_0 & i_13_43_1732_0 & ~i_13_43_2719_0) | (i_13_43_285_0 & ~i_13_43_1732_0 & ~i_13_43_2850_0) | (~i_13_43_649_0 & ~i_13_43_672_0 & ~i_13_43_1117_0 & ~i_13_43_1411_0 & ~i_13_43_3520_0) | (~i_13_43_228_0 & ~i_13_43_614_0 & i_13_43_1327_0 & ~i_13_43_3537_0));
endmodule



// Benchmark "kernel_13_44" written by ABC on Sun Jul 19 10:46:02 2020

module kernel_13_44 ( 
    i_13_44_31_0, i_13_44_61_0, i_13_44_99_0, i_13_44_116_0, i_13_44_184_0,
    i_13_44_186_0, i_13_44_187_0, i_13_44_229_0, i_13_44_258_0,
    i_13_44_259_0, i_13_44_426_0, i_13_44_431_0, i_13_44_526_0,
    i_13_44_601_0, i_13_44_618_0, i_13_44_619_0, i_13_44_620_0,
    i_13_44_628_0, i_13_44_670_0, i_13_44_691_0, i_13_44_756_0,
    i_13_44_799_0, i_13_44_800_0, i_13_44_840_0, i_13_44_962_0,
    i_13_44_1024_0, i_13_44_1077_0, i_13_44_1079_0, i_13_44_1123_0,
    i_13_44_1184_0, i_13_44_1187_0, i_13_44_1411_0, i_13_44_1444_0,
    i_13_44_1457_0, i_13_44_1482_0, i_13_44_1483_0, i_13_44_1519_0,
    i_13_44_1529_0, i_13_44_1573_0, i_13_44_1637_0, i_13_44_1677_0,
    i_13_44_1681_0, i_13_44_1747_0, i_13_44_1753_0, i_13_44_1771_0,
    i_13_44_1806_0, i_13_44_1807_0, i_13_44_1817_0, i_13_44_1861_0,
    i_13_44_1908_0, i_13_44_1912_0, i_13_44_1930_0, i_13_44_2001_0,
    i_13_44_2002_0, i_13_44_2003_0, i_13_44_2005_0, i_13_44_2024_0,
    i_13_44_2139_0, i_13_44_2140_0, i_13_44_2223_0, i_13_44_2224_0,
    i_13_44_2248_0, i_13_44_2259_0, i_13_44_2425_0, i_13_44_2446_0,
    i_13_44_2482_0, i_13_44_2653_0, i_13_44_2722_0, i_13_44_2743_0,
    i_13_44_2745_0, i_13_44_2751_0, i_13_44_2789_0, i_13_44_2798_0,
    i_13_44_2807_0, i_13_44_2857_0, i_13_44_3030_0, i_13_44_3122_0,
    i_13_44_3221_0, i_13_44_3244_0, i_13_44_3291_0, i_13_44_3293_0,
    i_13_44_3405_0, i_13_44_3439_0, i_13_44_3464_0, i_13_44_3525_0,
    i_13_44_3532_0, i_13_44_3552_0, i_13_44_3553_0, i_13_44_3759_0,
    i_13_44_3869_0, i_13_44_3905_0, i_13_44_4044_0, i_13_44_4054_0,
    i_13_44_4094_0, i_13_44_4152_0, i_13_44_4189_0, i_13_44_4317_0,
    i_13_44_4363_0, i_13_44_4387_0, i_13_44_4390_0,
    o_13_44_0_0  );
  input  i_13_44_31_0, i_13_44_61_0, i_13_44_99_0, i_13_44_116_0,
    i_13_44_184_0, i_13_44_186_0, i_13_44_187_0, i_13_44_229_0,
    i_13_44_258_0, i_13_44_259_0, i_13_44_426_0, i_13_44_431_0,
    i_13_44_526_0, i_13_44_601_0, i_13_44_618_0, i_13_44_619_0,
    i_13_44_620_0, i_13_44_628_0, i_13_44_670_0, i_13_44_691_0,
    i_13_44_756_0, i_13_44_799_0, i_13_44_800_0, i_13_44_840_0,
    i_13_44_962_0, i_13_44_1024_0, i_13_44_1077_0, i_13_44_1079_0,
    i_13_44_1123_0, i_13_44_1184_0, i_13_44_1187_0, i_13_44_1411_0,
    i_13_44_1444_0, i_13_44_1457_0, i_13_44_1482_0, i_13_44_1483_0,
    i_13_44_1519_0, i_13_44_1529_0, i_13_44_1573_0, i_13_44_1637_0,
    i_13_44_1677_0, i_13_44_1681_0, i_13_44_1747_0, i_13_44_1753_0,
    i_13_44_1771_0, i_13_44_1806_0, i_13_44_1807_0, i_13_44_1817_0,
    i_13_44_1861_0, i_13_44_1908_0, i_13_44_1912_0, i_13_44_1930_0,
    i_13_44_2001_0, i_13_44_2002_0, i_13_44_2003_0, i_13_44_2005_0,
    i_13_44_2024_0, i_13_44_2139_0, i_13_44_2140_0, i_13_44_2223_0,
    i_13_44_2224_0, i_13_44_2248_0, i_13_44_2259_0, i_13_44_2425_0,
    i_13_44_2446_0, i_13_44_2482_0, i_13_44_2653_0, i_13_44_2722_0,
    i_13_44_2743_0, i_13_44_2745_0, i_13_44_2751_0, i_13_44_2789_0,
    i_13_44_2798_0, i_13_44_2807_0, i_13_44_2857_0, i_13_44_3030_0,
    i_13_44_3122_0, i_13_44_3221_0, i_13_44_3244_0, i_13_44_3291_0,
    i_13_44_3293_0, i_13_44_3405_0, i_13_44_3439_0, i_13_44_3464_0,
    i_13_44_3525_0, i_13_44_3532_0, i_13_44_3552_0, i_13_44_3553_0,
    i_13_44_3759_0, i_13_44_3869_0, i_13_44_3905_0, i_13_44_4044_0,
    i_13_44_4054_0, i_13_44_4094_0, i_13_44_4152_0, i_13_44_4189_0,
    i_13_44_4317_0, i_13_44_4363_0, i_13_44_4387_0, i_13_44_4390_0;
  output o_13_44_0_0;
  assign o_13_44_0_0 = ~((~i_13_44_1483_0 & (i_13_44_2003_0 | (i_13_44_2002_0 & ~i_13_44_4189_0))) | (~i_13_44_619_0 & ~i_13_44_1411_0 & i_13_44_2002_0 & ~i_13_44_3464_0 & ~i_13_44_3759_0) | (~i_13_44_1079_0 & ~i_13_44_2024_0 & ~i_13_44_4152_0) | (~i_13_44_3293_0 & ~i_13_44_3525_0 & ~i_13_44_4363_0));
endmodule



// Benchmark "kernel_13_45" written by ABC on Sun Jul 19 10:46:03 2020

module kernel_13_45 ( 
    i_13_45_36_0, i_13_45_37_0, i_13_45_80_0, i_13_45_179_0, i_13_45_314_0,
    i_13_45_324_0, i_13_45_431_0, i_13_45_525_0, i_13_45_531_0,
    i_13_45_544_0, i_13_45_553_0, i_13_45_554_0, i_13_45_557_0,
    i_13_45_570_0, i_13_45_576_0, i_13_45_595_0, i_13_45_611_0,
    i_13_45_662_0, i_13_45_682_0, i_13_45_683_0, i_13_45_701_0,
    i_13_45_714_0, i_13_45_724_0, i_13_45_777_0, i_13_45_845_0,
    i_13_45_891_0, i_13_45_895_0, i_13_45_927_0, i_13_45_1041_0,
    i_13_45_1092_0, i_13_45_1151_0, i_13_45_1214_0, i_13_45_1369_0,
    i_13_45_1380_0, i_13_45_1399_0, i_13_45_1430_0, i_13_45_1461_0,
    i_13_45_1479_0, i_13_45_1480_0, i_13_45_1484_0, i_13_45_1596_0,
    i_13_45_1634_0, i_13_45_1710_0, i_13_45_1719_0, i_13_45_1720_0,
    i_13_45_1736_0, i_13_45_1767_0, i_13_45_1781_0, i_13_45_1782_0,
    i_13_45_1792_0, i_13_45_1881_0, i_13_45_1882_0, i_13_45_1952_0,
    i_13_45_2048_0, i_13_45_2129_0, i_13_45_2164_0, i_13_45_2210_0,
    i_13_45_2224_0, i_13_45_2236_0, i_13_45_2277_0, i_13_45_2307_0,
    i_13_45_2457_0, i_13_45_2600_0, i_13_45_2610_0, i_13_45_2629_0,
    i_13_45_2646_0, i_13_45_2649_0, i_13_45_2726_0, i_13_45_2820_0,
    i_13_45_2844_0, i_13_45_2845_0, i_13_45_2871_0, i_13_45_2885_0,
    i_13_45_3216_0, i_13_45_3420_0, i_13_45_3429_0, i_13_45_3448_0,
    i_13_45_3599_0, i_13_45_3743_0, i_13_45_3758_0, i_13_45_3784_0,
    i_13_45_3790_0, i_13_45_3866_0, i_13_45_3902_0, i_13_45_3924_0,
    i_13_45_3941_0, i_13_45_4014_0, i_13_45_4077_0, i_13_45_4114_0,
    i_13_45_4257_0, i_13_45_4265_0, i_13_45_4337_0, i_13_45_4360_0,
    i_13_45_4361_0, i_13_45_4436_0, i_13_45_4440_0, i_13_45_4540_0,
    i_13_45_4594_0, i_13_45_4598_0, i_13_45_4607_0,
    o_13_45_0_0  );
  input  i_13_45_36_0, i_13_45_37_0, i_13_45_80_0, i_13_45_179_0,
    i_13_45_314_0, i_13_45_324_0, i_13_45_431_0, i_13_45_525_0,
    i_13_45_531_0, i_13_45_544_0, i_13_45_553_0, i_13_45_554_0,
    i_13_45_557_0, i_13_45_570_0, i_13_45_576_0, i_13_45_595_0,
    i_13_45_611_0, i_13_45_662_0, i_13_45_682_0, i_13_45_683_0,
    i_13_45_701_0, i_13_45_714_0, i_13_45_724_0, i_13_45_777_0,
    i_13_45_845_0, i_13_45_891_0, i_13_45_895_0, i_13_45_927_0,
    i_13_45_1041_0, i_13_45_1092_0, i_13_45_1151_0, i_13_45_1214_0,
    i_13_45_1369_0, i_13_45_1380_0, i_13_45_1399_0, i_13_45_1430_0,
    i_13_45_1461_0, i_13_45_1479_0, i_13_45_1480_0, i_13_45_1484_0,
    i_13_45_1596_0, i_13_45_1634_0, i_13_45_1710_0, i_13_45_1719_0,
    i_13_45_1720_0, i_13_45_1736_0, i_13_45_1767_0, i_13_45_1781_0,
    i_13_45_1782_0, i_13_45_1792_0, i_13_45_1881_0, i_13_45_1882_0,
    i_13_45_1952_0, i_13_45_2048_0, i_13_45_2129_0, i_13_45_2164_0,
    i_13_45_2210_0, i_13_45_2224_0, i_13_45_2236_0, i_13_45_2277_0,
    i_13_45_2307_0, i_13_45_2457_0, i_13_45_2600_0, i_13_45_2610_0,
    i_13_45_2629_0, i_13_45_2646_0, i_13_45_2649_0, i_13_45_2726_0,
    i_13_45_2820_0, i_13_45_2844_0, i_13_45_2845_0, i_13_45_2871_0,
    i_13_45_2885_0, i_13_45_3216_0, i_13_45_3420_0, i_13_45_3429_0,
    i_13_45_3448_0, i_13_45_3599_0, i_13_45_3743_0, i_13_45_3758_0,
    i_13_45_3784_0, i_13_45_3790_0, i_13_45_3866_0, i_13_45_3902_0,
    i_13_45_3924_0, i_13_45_3941_0, i_13_45_4014_0, i_13_45_4077_0,
    i_13_45_4114_0, i_13_45_4257_0, i_13_45_4265_0, i_13_45_4337_0,
    i_13_45_4360_0, i_13_45_4361_0, i_13_45_4436_0, i_13_45_4440_0,
    i_13_45_4540_0, i_13_45_4594_0, i_13_45_4598_0, i_13_45_4607_0;
  output o_13_45_0_0;
  assign o_13_45_0_0 = ~((~i_13_45_3448_0 & (~i_13_45_1767_0 | (i_13_45_1596_0 & ~i_13_45_2457_0 & ~i_13_45_4077_0))) | (~i_13_45_4360_0 & (~i_13_45_4077_0 | (~i_13_45_2610_0 & ~i_13_45_3216_0))) | (~i_13_45_324_0 & ~i_13_45_927_0 & ~i_13_45_2649_0 & ~i_13_45_2845_0) | (~i_13_45_2224_0 & ~i_13_45_2871_0 & i_13_45_3448_0) | (~i_13_45_531_0 & ~i_13_45_3784_0) | (~i_13_45_1480_0 & i_13_45_4361_0));
endmodule



// Benchmark "kernel_13_46" written by ABC on Sun Jul 19 10:46:04 2020

module kernel_13_46 ( 
    i_13_46_114_0, i_13_46_127_0, i_13_46_159_0, i_13_46_160_0,
    i_13_46_166_0, i_13_46_211_0, i_13_46_241_0, i_13_46_247_0,
    i_13_46_268_0, i_13_46_269_0, i_13_46_275_0, i_13_46_319_0,
    i_13_46_340_0, i_13_46_357_0, i_13_46_375_0, i_13_46_443_0,
    i_13_46_465_0, i_13_46_466_0, i_13_46_519_0, i_13_46_520_0,
    i_13_46_536_0, i_13_46_643_0, i_13_46_699_0, i_13_46_714_0,
    i_13_46_744_0, i_13_46_745_0, i_13_46_762_0, i_13_46_862_0,
    i_13_46_947_0, i_13_46_1123_0, i_13_46_1212_0, i_13_46_1213_0,
    i_13_46_1255_0, i_13_46_1303_0, i_13_46_1347_0, i_13_46_1400_0,
    i_13_46_1411_0, i_13_46_1428_0, i_13_46_1456_0, i_13_46_1482_0,
    i_13_46_1483_0, i_13_46_1774_0, i_13_46_1775_0, i_13_46_1813_0,
    i_13_46_1816_0, i_13_46_1945_0, i_13_46_1946_0, i_13_46_2059_0,
    i_13_46_2132_0, i_13_46_2181_0, i_13_46_2202_0, i_13_46_2283_0,
    i_13_46_2284_0, i_13_46_2285_0, i_13_46_2354_0, i_13_46_2417_0,
    i_13_46_2496_0, i_13_46_2715_0, i_13_46_2724_0, i_13_46_2725_0,
    i_13_46_2770_0, i_13_46_2771_0, i_13_46_2788_0, i_13_46_2792_0,
    i_13_46_2938_0, i_13_46_3048_0, i_13_46_3056_0, i_13_46_3063_0,
    i_13_46_3068_0, i_13_46_3122_0, i_13_46_3144_0, i_13_46_3220_0,
    i_13_46_3235_0, i_13_46_3271_0, i_13_46_3373_0, i_13_46_3419_0,
    i_13_46_3441_0, i_13_46_3453_0, i_13_46_3523_0, i_13_46_3530_0,
    i_13_46_3597_0, i_13_46_3598_0, i_13_46_3617_0, i_13_46_3621_0,
    i_13_46_3635_0, i_13_46_3666_0, i_13_46_3685_0, i_13_46_3824_0,
    i_13_46_3875_0, i_13_46_3922_0, i_13_46_4057_0, i_13_46_4081_0,
    i_13_46_4093_0, i_13_46_4184_0, i_13_46_4197_0, i_13_46_4261_0,
    i_13_46_4272_0, i_13_46_4273_0, i_13_46_4274_0, i_13_46_4399_0,
    o_13_46_0_0  );
  input  i_13_46_114_0, i_13_46_127_0, i_13_46_159_0, i_13_46_160_0,
    i_13_46_166_0, i_13_46_211_0, i_13_46_241_0, i_13_46_247_0,
    i_13_46_268_0, i_13_46_269_0, i_13_46_275_0, i_13_46_319_0,
    i_13_46_340_0, i_13_46_357_0, i_13_46_375_0, i_13_46_443_0,
    i_13_46_465_0, i_13_46_466_0, i_13_46_519_0, i_13_46_520_0,
    i_13_46_536_0, i_13_46_643_0, i_13_46_699_0, i_13_46_714_0,
    i_13_46_744_0, i_13_46_745_0, i_13_46_762_0, i_13_46_862_0,
    i_13_46_947_0, i_13_46_1123_0, i_13_46_1212_0, i_13_46_1213_0,
    i_13_46_1255_0, i_13_46_1303_0, i_13_46_1347_0, i_13_46_1400_0,
    i_13_46_1411_0, i_13_46_1428_0, i_13_46_1456_0, i_13_46_1482_0,
    i_13_46_1483_0, i_13_46_1774_0, i_13_46_1775_0, i_13_46_1813_0,
    i_13_46_1816_0, i_13_46_1945_0, i_13_46_1946_0, i_13_46_2059_0,
    i_13_46_2132_0, i_13_46_2181_0, i_13_46_2202_0, i_13_46_2283_0,
    i_13_46_2284_0, i_13_46_2285_0, i_13_46_2354_0, i_13_46_2417_0,
    i_13_46_2496_0, i_13_46_2715_0, i_13_46_2724_0, i_13_46_2725_0,
    i_13_46_2770_0, i_13_46_2771_0, i_13_46_2788_0, i_13_46_2792_0,
    i_13_46_2938_0, i_13_46_3048_0, i_13_46_3056_0, i_13_46_3063_0,
    i_13_46_3068_0, i_13_46_3122_0, i_13_46_3144_0, i_13_46_3220_0,
    i_13_46_3235_0, i_13_46_3271_0, i_13_46_3373_0, i_13_46_3419_0,
    i_13_46_3441_0, i_13_46_3453_0, i_13_46_3523_0, i_13_46_3530_0,
    i_13_46_3597_0, i_13_46_3598_0, i_13_46_3617_0, i_13_46_3621_0,
    i_13_46_3635_0, i_13_46_3666_0, i_13_46_3685_0, i_13_46_3824_0,
    i_13_46_3875_0, i_13_46_3922_0, i_13_46_4057_0, i_13_46_4081_0,
    i_13_46_4093_0, i_13_46_4184_0, i_13_46_4197_0, i_13_46_4261_0,
    i_13_46_4272_0, i_13_46_4273_0, i_13_46_4274_0, i_13_46_4399_0;
  output o_13_46_0_0;
  assign o_13_46_0_0 = ~((~i_13_46_762_0 & ~i_13_46_3235_0 & ~i_13_46_3685_0) | (~i_13_46_241_0 & ~i_13_46_466_0 & ~i_13_46_519_0 & ~i_13_46_3597_0 & ~i_13_46_4093_0));
endmodule



// Benchmark "kernel_13_47" written by ABC on Sun Jul 19 10:46:04 2020

module kernel_13_47 ( 
    i_13_47_63_0, i_13_47_97_0, i_13_47_124_0, i_13_47_125_0,
    i_13_47_140_0, i_13_47_187_0, i_13_47_188_0, i_13_47_196_0,
    i_13_47_328_0, i_13_47_374_0, i_13_47_520_0, i_13_47_536_0,
    i_13_47_552_0, i_13_47_574_0, i_13_47_577_0, i_13_47_580_0,
    i_13_47_583_0, i_13_47_592_0, i_13_47_603_0, i_13_47_641_0,
    i_13_47_664_0, i_13_47_715_0, i_13_47_718_0, i_13_47_729_0,
    i_13_47_745_0, i_13_47_781_0, i_13_47_793_0, i_13_47_800_0,
    i_13_47_862_0, i_13_47_863_0, i_13_47_886_0, i_13_47_989_0,
    i_13_47_1025_0, i_13_47_1135_0, i_13_47_1193_0, i_13_47_1258_0,
    i_13_47_1411_0, i_13_47_1447_0, i_13_47_1457_0, i_13_47_1493_0,
    i_13_47_1502_0, i_13_47_1573_0, i_13_47_1627_0, i_13_47_1636_0,
    i_13_47_1744_0, i_13_47_1751_0, i_13_47_1787_0, i_13_47_1831_0,
    i_13_47_1836_0, i_13_47_1859_0, i_13_47_1871_0, i_13_47_1885_0,
    i_13_47_1952_0, i_13_47_2015_0, i_13_47_2029_0, i_13_47_2168_0,
    i_13_47_2177_0, i_13_47_2267_0, i_13_47_2362_0, i_13_47_2383_0,
    i_13_47_2428_0, i_13_47_2465_0, i_13_47_2503_0, i_13_47_2536_0,
    i_13_47_2537_0, i_13_47_2633_0, i_13_47_2770_0, i_13_47_2825_0,
    i_13_47_2984_0, i_13_47_3004_0, i_13_47_3040_0, i_13_47_3159_0,
    i_13_47_3167_0, i_13_47_3175_0, i_13_47_3246_0, i_13_47_3290_0,
    i_13_47_3322_0, i_13_47_3323_0, i_13_47_3427_0, i_13_47_3428_0,
    i_13_47_3466_0, i_13_47_3581_0, i_13_47_3617_0, i_13_47_3699_0,
    i_13_47_3748_0, i_13_47_3787_0, i_13_47_3794_0, i_13_47_3806_0,
    i_13_47_3839_0, i_13_47_3877_0, i_13_47_3914_0, i_13_47_3922_0,
    i_13_47_4012_0, i_13_47_4013_0, i_13_47_4081_0, i_13_47_4171_0,
    i_13_47_4522_0, i_13_47_4566_0, i_13_47_4586_0, i_13_47_4588_0,
    o_13_47_0_0  );
  input  i_13_47_63_0, i_13_47_97_0, i_13_47_124_0, i_13_47_125_0,
    i_13_47_140_0, i_13_47_187_0, i_13_47_188_0, i_13_47_196_0,
    i_13_47_328_0, i_13_47_374_0, i_13_47_520_0, i_13_47_536_0,
    i_13_47_552_0, i_13_47_574_0, i_13_47_577_0, i_13_47_580_0,
    i_13_47_583_0, i_13_47_592_0, i_13_47_603_0, i_13_47_641_0,
    i_13_47_664_0, i_13_47_715_0, i_13_47_718_0, i_13_47_729_0,
    i_13_47_745_0, i_13_47_781_0, i_13_47_793_0, i_13_47_800_0,
    i_13_47_862_0, i_13_47_863_0, i_13_47_886_0, i_13_47_989_0,
    i_13_47_1025_0, i_13_47_1135_0, i_13_47_1193_0, i_13_47_1258_0,
    i_13_47_1411_0, i_13_47_1447_0, i_13_47_1457_0, i_13_47_1493_0,
    i_13_47_1502_0, i_13_47_1573_0, i_13_47_1627_0, i_13_47_1636_0,
    i_13_47_1744_0, i_13_47_1751_0, i_13_47_1787_0, i_13_47_1831_0,
    i_13_47_1836_0, i_13_47_1859_0, i_13_47_1871_0, i_13_47_1885_0,
    i_13_47_1952_0, i_13_47_2015_0, i_13_47_2029_0, i_13_47_2168_0,
    i_13_47_2177_0, i_13_47_2267_0, i_13_47_2362_0, i_13_47_2383_0,
    i_13_47_2428_0, i_13_47_2465_0, i_13_47_2503_0, i_13_47_2536_0,
    i_13_47_2537_0, i_13_47_2633_0, i_13_47_2770_0, i_13_47_2825_0,
    i_13_47_2984_0, i_13_47_3004_0, i_13_47_3040_0, i_13_47_3159_0,
    i_13_47_3167_0, i_13_47_3175_0, i_13_47_3246_0, i_13_47_3290_0,
    i_13_47_3322_0, i_13_47_3323_0, i_13_47_3427_0, i_13_47_3428_0,
    i_13_47_3466_0, i_13_47_3581_0, i_13_47_3617_0, i_13_47_3699_0,
    i_13_47_3748_0, i_13_47_3787_0, i_13_47_3794_0, i_13_47_3806_0,
    i_13_47_3839_0, i_13_47_3877_0, i_13_47_3914_0, i_13_47_3922_0,
    i_13_47_4012_0, i_13_47_4013_0, i_13_47_4081_0, i_13_47_4171_0,
    i_13_47_4522_0, i_13_47_4566_0, i_13_47_4586_0, i_13_47_4588_0;
  output o_13_47_0_0;
  assign o_13_47_0_0 = 0;
endmodule



// Benchmark "kernel_13_48" written by ABC on Sun Jul 19 10:46:05 2020

module kernel_13_48 ( 
    i_13_48_37_0, i_13_48_59_0, i_13_48_136_0, i_13_48_167_0,
    i_13_48_230_0, i_13_48_260_0, i_13_48_283_0, i_13_48_308_0,
    i_13_48_545_0, i_13_48_577_0, i_13_48_596_0, i_13_48_617_0,
    i_13_48_625_0, i_13_48_626_0, i_13_48_646_0, i_13_48_671_0,
    i_13_48_717_0, i_13_48_728_0, i_13_48_778_0, i_13_48_779_0,
    i_13_48_838_0, i_13_48_839_0, i_13_48_852_0, i_13_48_865_0,
    i_13_48_911_0, i_13_48_956_0, i_13_48_1022_0, i_13_48_1094_0,
    i_13_48_1097_0, i_13_48_1118_0, i_13_48_1121_0, i_13_48_1146_0,
    i_13_48_1228_0, i_13_48_1281_0, i_13_48_1301_0, i_13_48_1318_0,
    i_13_48_1462_0, i_13_48_1464_0, i_13_48_1480_0, i_13_48_1481_0,
    i_13_48_1484_0, i_13_48_1522_0, i_13_48_1643_0, i_13_48_1675_0,
    i_13_48_1678_0, i_13_48_1688_0, i_13_48_1691_0, i_13_48_1721_0,
    i_13_48_1747_0, i_13_48_1750_0, i_13_48_1757_0, i_13_48_1768_0,
    i_13_48_1804_0, i_13_48_1805_0, i_13_48_1857_0, i_13_48_1858_0,
    i_13_48_1860_0, i_13_48_2002_0, i_13_48_2120_0, i_13_48_2138_0,
    i_13_48_2139_0, i_13_48_2165_0, i_13_48_2225_0, i_13_48_2308_0,
    i_13_48_2380_0, i_13_48_2425_0, i_13_48_2443_0, i_13_48_2444_0,
    i_13_48_2446_0, i_13_48_2447_0, i_13_48_2647_0, i_13_48_2650_0,
    i_13_48_2692_0, i_13_48_2693_0, i_13_48_2822_0, i_13_48_2999_0,
    i_13_48_3012_0, i_13_48_3076_0, i_13_48_3094_0, i_13_48_3110_0,
    i_13_48_3197_0, i_13_48_3290_0, i_13_48_3320_0, i_13_48_3353_0,
    i_13_48_3430_0, i_13_48_3560_0, i_13_48_3741_0, i_13_48_3911_0,
    i_13_48_3989_0, i_13_48_4115_0, i_13_48_4187_0, i_13_48_4189_0,
    i_13_48_4235_0, i_13_48_4263_0, i_13_48_4300_0, i_13_48_4351_0,
    i_13_48_4352_0, i_13_48_4379_0, i_13_48_4396_0, i_13_48_4441_0,
    o_13_48_0_0  );
  input  i_13_48_37_0, i_13_48_59_0, i_13_48_136_0, i_13_48_167_0,
    i_13_48_230_0, i_13_48_260_0, i_13_48_283_0, i_13_48_308_0,
    i_13_48_545_0, i_13_48_577_0, i_13_48_596_0, i_13_48_617_0,
    i_13_48_625_0, i_13_48_626_0, i_13_48_646_0, i_13_48_671_0,
    i_13_48_717_0, i_13_48_728_0, i_13_48_778_0, i_13_48_779_0,
    i_13_48_838_0, i_13_48_839_0, i_13_48_852_0, i_13_48_865_0,
    i_13_48_911_0, i_13_48_956_0, i_13_48_1022_0, i_13_48_1094_0,
    i_13_48_1097_0, i_13_48_1118_0, i_13_48_1121_0, i_13_48_1146_0,
    i_13_48_1228_0, i_13_48_1281_0, i_13_48_1301_0, i_13_48_1318_0,
    i_13_48_1462_0, i_13_48_1464_0, i_13_48_1480_0, i_13_48_1481_0,
    i_13_48_1484_0, i_13_48_1522_0, i_13_48_1643_0, i_13_48_1675_0,
    i_13_48_1678_0, i_13_48_1688_0, i_13_48_1691_0, i_13_48_1721_0,
    i_13_48_1747_0, i_13_48_1750_0, i_13_48_1757_0, i_13_48_1768_0,
    i_13_48_1804_0, i_13_48_1805_0, i_13_48_1857_0, i_13_48_1858_0,
    i_13_48_1860_0, i_13_48_2002_0, i_13_48_2120_0, i_13_48_2138_0,
    i_13_48_2139_0, i_13_48_2165_0, i_13_48_2225_0, i_13_48_2308_0,
    i_13_48_2380_0, i_13_48_2425_0, i_13_48_2443_0, i_13_48_2444_0,
    i_13_48_2446_0, i_13_48_2447_0, i_13_48_2647_0, i_13_48_2650_0,
    i_13_48_2692_0, i_13_48_2693_0, i_13_48_2822_0, i_13_48_2999_0,
    i_13_48_3012_0, i_13_48_3076_0, i_13_48_3094_0, i_13_48_3110_0,
    i_13_48_3197_0, i_13_48_3290_0, i_13_48_3320_0, i_13_48_3353_0,
    i_13_48_3430_0, i_13_48_3560_0, i_13_48_3741_0, i_13_48_3911_0,
    i_13_48_3989_0, i_13_48_4115_0, i_13_48_4187_0, i_13_48_4189_0,
    i_13_48_4235_0, i_13_48_4263_0, i_13_48_4300_0, i_13_48_4351_0,
    i_13_48_4352_0, i_13_48_4379_0, i_13_48_4396_0, i_13_48_4441_0;
  output o_13_48_0_0;
  assign o_13_48_0_0 = 0;
endmodule



// Benchmark "kernel_13_49" written by ABC on Sun Jul 19 10:46:06 2020

module kernel_13_49 ( 
    i_13_49_22_0, i_13_49_61_0, i_13_49_79_0, i_13_49_94_0, i_13_49_95_0,
    i_13_49_259_0, i_13_49_261_0, i_13_49_319_0, i_13_49_322_0,
    i_13_49_336_0, i_13_49_492_0, i_13_49_521_0, i_13_49_619_0,
    i_13_49_697_0, i_13_49_700_0, i_13_49_745_0, i_13_49_823_0,
    i_13_49_835_0, i_13_49_837_0, i_13_49_870_0, i_13_49_960_0,
    i_13_49_970_0, i_13_49_978_0, i_13_49_979_0, i_13_49_980_0,
    i_13_49_1025_0, i_13_49_1075_0, i_13_49_1076_0, i_13_49_1095_0,
    i_13_49_1213_0, i_13_49_1281_0, i_13_49_1283_0, i_13_49_1302_0,
    i_13_49_1320_0, i_13_49_1321_0, i_13_49_1364_0, i_13_49_1384_0,
    i_13_49_1434_0, i_13_49_1438_0, i_13_49_1444_0, i_13_49_1464_0,
    i_13_49_1483_0, i_13_49_1568_0, i_13_49_1658_0, i_13_49_1813_0,
    i_13_49_1816_0, i_13_49_1817_0, i_13_49_1830_0, i_13_49_1870_0,
    i_13_49_1921_0, i_13_49_1943_0, i_13_49_1951_0, i_13_49_2082_0,
    i_13_49_2176_0, i_13_49_2209_0, i_13_49_2248_0, i_13_49_2425_0,
    i_13_49_2445_0, i_13_49_2446_0, i_13_49_2447_0, i_13_49_2460_0,
    i_13_49_2511_0, i_13_49_2516_0, i_13_49_2542_0, i_13_49_2554_0,
    i_13_49_2619_0, i_13_49_2923_0, i_13_49_3004_0, i_13_49_3056_0,
    i_13_49_3077_0, i_13_49_3094_0, i_13_49_3130_0, i_13_49_3220_0,
    i_13_49_3306_0, i_13_49_3418_0, i_13_49_3419_0, i_13_49_3433_0,
    i_13_49_3444_0, i_13_49_3482_0, i_13_49_3490_0, i_13_49_3550_0,
    i_13_49_3598_0, i_13_49_3737_0, i_13_49_3821_0, i_13_49_3874_0,
    i_13_49_3888_0, i_13_49_3992_0, i_13_49_4004_0, i_13_49_4018_0,
    i_13_49_4087_0, i_13_49_4188_0, i_13_49_4273_0, i_13_49_4333_0,
    i_13_49_4347_0, i_13_49_4351_0, i_13_49_4354_0, i_13_49_4381_0,
    i_13_49_4382_0, i_13_49_4390_0, i_13_49_4586_0,
    o_13_49_0_0  );
  input  i_13_49_22_0, i_13_49_61_0, i_13_49_79_0, i_13_49_94_0,
    i_13_49_95_0, i_13_49_259_0, i_13_49_261_0, i_13_49_319_0,
    i_13_49_322_0, i_13_49_336_0, i_13_49_492_0, i_13_49_521_0,
    i_13_49_619_0, i_13_49_697_0, i_13_49_700_0, i_13_49_745_0,
    i_13_49_823_0, i_13_49_835_0, i_13_49_837_0, i_13_49_870_0,
    i_13_49_960_0, i_13_49_970_0, i_13_49_978_0, i_13_49_979_0,
    i_13_49_980_0, i_13_49_1025_0, i_13_49_1075_0, i_13_49_1076_0,
    i_13_49_1095_0, i_13_49_1213_0, i_13_49_1281_0, i_13_49_1283_0,
    i_13_49_1302_0, i_13_49_1320_0, i_13_49_1321_0, i_13_49_1364_0,
    i_13_49_1384_0, i_13_49_1434_0, i_13_49_1438_0, i_13_49_1444_0,
    i_13_49_1464_0, i_13_49_1483_0, i_13_49_1568_0, i_13_49_1658_0,
    i_13_49_1813_0, i_13_49_1816_0, i_13_49_1817_0, i_13_49_1830_0,
    i_13_49_1870_0, i_13_49_1921_0, i_13_49_1943_0, i_13_49_1951_0,
    i_13_49_2082_0, i_13_49_2176_0, i_13_49_2209_0, i_13_49_2248_0,
    i_13_49_2425_0, i_13_49_2445_0, i_13_49_2446_0, i_13_49_2447_0,
    i_13_49_2460_0, i_13_49_2511_0, i_13_49_2516_0, i_13_49_2542_0,
    i_13_49_2554_0, i_13_49_2619_0, i_13_49_2923_0, i_13_49_3004_0,
    i_13_49_3056_0, i_13_49_3077_0, i_13_49_3094_0, i_13_49_3130_0,
    i_13_49_3220_0, i_13_49_3306_0, i_13_49_3418_0, i_13_49_3419_0,
    i_13_49_3433_0, i_13_49_3444_0, i_13_49_3482_0, i_13_49_3490_0,
    i_13_49_3550_0, i_13_49_3598_0, i_13_49_3737_0, i_13_49_3821_0,
    i_13_49_3874_0, i_13_49_3888_0, i_13_49_3992_0, i_13_49_4004_0,
    i_13_49_4018_0, i_13_49_4087_0, i_13_49_4188_0, i_13_49_4273_0,
    i_13_49_4333_0, i_13_49_4347_0, i_13_49_4351_0, i_13_49_4354_0,
    i_13_49_4381_0, i_13_49_4382_0, i_13_49_4390_0, i_13_49_4586_0;
  output o_13_49_0_0;
  assign o_13_49_0_0 = ~((~i_13_49_2446_0 & (~i_13_49_3220_0 | (~i_13_49_79_0 & ~i_13_49_3821_0))) | (~i_13_49_4354_0 & (~i_13_49_1321_0 | (~i_13_49_1483_0 & i_13_49_2176_0))) | (i_13_49_94_0 & ~i_13_49_697_0) | (~i_13_49_1213_0 & i_13_49_3821_0));
endmodule



// Benchmark "kernel_13_50" written by ABC on Sun Jul 19 10:46:07 2020

module kernel_13_50 ( 
    i_13_50_72_0, i_13_50_75_0, i_13_50_78_0, i_13_50_112_0, i_13_50_141_0,
    i_13_50_240_0, i_13_50_250_0, i_13_50_258_0, i_13_50_282_0,
    i_13_50_310_0, i_13_50_372_0, i_13_50_559_0, i_13_50_579_0,
    i_13_50_618_0, i_13_50_619_0, i_13_50_697_0, i_13_50_699_0,
    i_13_50_816_0, i_13_50_843_0, i_13_50_931_0, i_13_50_1023_0,
    i_13_50_1024_0, i_13_50_1077_0, i_13_50_1078_0, i_13_50_1084_0,
    i_13_50_1143_0, i_13_50_1204_0, i_13_50_1212_0, i_13_50_1255_0,
    i_13_50_1273_0, i_13_50_1284_0, i_13_50_1317_0, i_13_50_1332_0,
    i_13_50_1348_0, i_13_50_1427_0, i_13_50_1468_0, i_13_50_1513_0,
    i_13_50_1521_0, i_13_50_1572_0, i_13_50_1573_0, i_13_50_1597_0,
    i_13_50_1609_0, i_13_50_1633_0, i_13_50_1635_0, i_13_50_1725_0,
    i_13_50_1812_0, i_13_50_1843_0, i_13_50_1849_0, i_13_50_1881_0,
    i_13_50_1888_0, i_13_50_2103_0, i_13_50_2198_0, i_13_50_2278_0,
    i_13_50_2404_0, i_13_50_2442_0, i_13_50_2454_0, i_13_50_2563_0,
    i_13_50_2710_0, i_13_50_2712_0, i_13_50_2715_0, i_13_50_2742_0,
    i_13_50_2887_0, i_13_50_2955_0, i_13_50_2958_0, i_13_50_3036_0,
    i_13_50_3169_0, i_13_50_3204_0, i_13_50_3208_0, i_13_50_3241_0,
    i_13_50_3244_0, i_13_50_3291_0, i_13_50_3379_0, i_13_50_3412_0,
    i_13_50_3450_0, i_13_50_3451_0, i_13_50_3453_0, i_13_50_3454_0,
    i_13_50_3462_0, i_13_50_3525_0, i_13_50_3532_0, i_13_50_3570_0,
    i_13_50_3571_0, i_13_50_3649_0, i_13_50_3684_0, i_13_50_3685_0,
    i_13_50_3687_0, i_13_50_3688_0, i_13_50_3708_0, i_13_50_3756_0,
    i_13_50_3757_0, i_13_50_3781_0, i_13_50_3982_0, i_13_50_4020_0,
    i_13_50_4188_0, i_13_50_4233_0, i_13_50_4260_0, i_13_50_4312_0,
    i_13_50_4393_0, i_13_50_4497_0, i_13_50_4509_0,
    o_13_50_0_0  );
  input  i_13_50_72_0, i_13_50_75_0, i_13_50_78_0, i_13_50_112_0,
    i_13_50_141_0, i_13_50_240_0, i_13_50_250_0, i_13_50_258_0,
    i_13_50_282_0, i_13_50_310_0, i_13_50_372_0, i_13_50_559_0,
    i_13_50_579_0, i_13_50_618_0, i_13_50_619_0, i_13_50_697_0,
    i_13_50_699_0, i_13_50_816_0, i_13_50_843_0, i_13_50_931_0,
    i_13_50_1023_0, i_13_50_1024_0, i_13_50_1077_0, i_13_50_1078_0,
    i_13_50_1084_0, i_13_50_1143_0, i_13_50_1204_0, i_13_50_1212_0,
    i_13_50_1255_0, i_13_50_1273_0, i_13_50_1284_0, i_13_50_1317_0,
    i_13_50_1332_0, i_13_50_1348_0, i_13_50_1427_0, i_13_50_1468_0,
    i_13_50_1513_0, i_13_50_1521_0, i_13_50_1572_0, i_13_50_1573_0,
    i_13_50_1597_0, i_13_50_1609_0, i_13_50_1633_0, i_13_50_1635_0,
    i_13_50_1725_0, i_13_50_1812_0, i_13_50_1843_0, i_13_50_1849_0,
    i_13_50_1881_0, i_13_50_1888_0, i_13_50_2103_0, i_13_50_2198_0,
    i_13_50_2278_0, i_13_50_2404_0, i_13_50_2442_0, i_13_50_2454_0,
    i_13_50_2563_0, i_13_50_2710_0, i_13_50_2712_0, i_13_50_2715_0,
    i_13_50_2742_0, i_13_50_2887_0, i_13_50_2955_0, i_13_50_2958_0,
    i_13_50_3036_0, i_13_50_3169_0, i_13_50_3204_0, i_13_50_3208_0,
    i_13_50_3241_0, i_13_50_3244_0, i_13_50_3291_0, i_13_50_3379_0,
    i_13_50_3412_0, i_13_50_3450_0, i_13_50_3451_0, i_13_50_3453_0,
    i_13_50_3454_0, i_13_50_3462_0, i_13_50_3525_0, i_13_50_3532_0,
    i_13_50_3570_0, i_13_50_3571_0, i_13_50_3649_0, i_13_50_3684_0,
    i_13_50_3685_0, i_13_50_3687_0, i_13_50_3688_0, i_13_50_3708_0,
    i_13_50_3756_0, i_13_50_3757_0, i_13_50_3781_0, i_13_50_3982_0,
    i_13_50_4020_0, i_13_50_4188_0, i_13_50_4233_0, i_13_50_4260_0,
    i_13_50_4312_0, i_13_50_4393_0, i_13_50_4497_0, i_13_50_4509_0;
  output o_13_50_0_0;
  assign o_13_50_0_0 = ~(~i_13_50_618_0 | ~i_13_50_3685_0);
endmodule



// Benchmark "kernel_13_51" written by ABC on Sun Jul 19 10:46:07 2020

module kernel_13_51 ( 
    i_13_51_35_0, i_13_51_76_0, i_13_51_94_0, i_13_51_121_0, i_13_51_184_0,
    i_13_51_193_0, i_13_51_241_0, i_13_51_251_0, i_13_51_260_0,
    i_13_51_278_0, i_13_51_358_0, i_13_51_361_0, i_13_51_521_0,
    i_13_51_527_0, i_13_51_535_0, i_13_51_616_0, i_13_51_652_0,
    i_13_51_664_0, i_13_51_715_0, i_13_51_896_0, i_13_51_898_0,
    i_13_51_1024_0, i_13_51_1025_0, i_13_51_1078_0, i_13_51_1079_0,
    i_13_51_1211_0, i_13_51_1213_0, i_13_51_1244_0, i_13_51_1259_0,
    i_13_51_1286_0, i_13_51_1331_0, i_13_51_1349_0, i_13_51_1400_0,
    i_13_51_1408_0, i_13_51_1424_0, i_13_51_1427_0, i_13_51_1430_0,
    i_13_51_1483_0, i_13_51_1501_0, i_13_51_1502_0, i_13_51_1508_0,
    i_13_51_1609_0, i_13_51_1637_0, i_13_51_1696_0, i_13_51_1817_0,
    i_13_51_1835_0, i_13_51_1841_0, i_13_51_1921_0, i_13_51_1943_0,
    i_13_51_1961_0, i_13_51_2005_0, i_13_51_2006_0, i_13_51_2033_0,
    i_13_51_2131_0, i_13_51_2201_0, i_13_51_2315_0, i_13_51_2360_0,
    i_13_51_2455_0, i_13_51_2456_0, i_13_51_2471_0, i_13_51_2546_0,
    i_13_51_2573_0, i_13_51_2651_0, i_13_51_2716_0, i_13_51_2717_0,
    i_13_51_2726_0, i_13_51_2768_0, i_13_51_2923_0, i_13_51_2924_0,
    i_13_51_2959_0, i_13_51_2965_0, i_13_51_3163_0, i_13_51_3373_0,
    i_13_51_3374_0, i_13_51_3419_0, i_13_51_3565_0, i_13_51_3580_0,
    i_13_51_3599_0, i_13_51_3650_0, i_13_51_3731_0, i_13_51_3733_0,
    i_13_51_3734_0, i_13_51_3787_0, i_13_51_3905_0, i_13_51_3910_0,
    i_13_51_3919_0, i_13_51_3923_0, i_13_51_3985_0, i_13_51_4253_0,
    i_13_51_4255_0, i_13_51_4256_0, i_13_51_4262_0, i_13_51_4265_0,
    i_13_51_4453_0, i_13_51_4454_0, i_13_51_4526_0, i_13_51_4541_0,
    i_13_51_4558_0, i_13_51_4559_0, i_13_51_4561_0,
    o_13_51_0_0  );
  input  i_13_51_35_0, i_13_51_76_0, i_13_51_94_0, i_13_51_121_0,
    i_13_51_184_0, i_13_51_193_0, i_13_51_241_0, i_13_51_251_0,
    i_13_51_260_0, i_13_51_278_0, i_13_51_358_0, i_13_51_361_0,
    i_13_51_521_0, i_13_51_527_0, i_13_51_535_0, i_13_51_616_0,
    i_13_51_652_0, i_13_51_664_0, i_13_51_715_0, i_13_51_896_0,
    i_13_51_898_0, i_13_51_1024_0, i_13_51_1025_0, i_13_51_1078_0,
    i_13_51_1079_0, i_13_51_1211_0, i_13_51_1213_0, i_13_51_1244_0,
    i_13_51_1259_0, i_13_51_1286_0, i_13_51_1331_0, i_13_51_1349_0,
    i_13_51_1400_0, i_13_51_1408_0, i_13_51_1424_0, i_13_51_1427_0,
    i_13_51_1430_0, i_13_51_1483_0, i_13_51_1501_0, i_13_51_1502_0,
    i_13_51_1508_0, i_13_51_1609_0, i_13_51_1637_0, i_13_51_1696_0,
    i_13_51_1817_0, i_13_51_1835_0, i_13_51_1841_0, i_13_51_1921_0,
    i_13_51_1943_0, i_13_51_1961_0, i_13_51_2005_0, i_13_51_2006_0,
    i_13_51_2033_0, i_13_51_2131_0, i_13_51_2201_0, i_13_51_2315_0,
    i_13_51_2360_0, i_13_51_2455_0, i_13_51_2456_0, i_13_51_2471_0,
    i_13_51_2546_0, i_13_51_2573_0, i_13_51_2651_0, i_13_51_2716_0,
    i_13_51_2717_0, i_13_51_2726_0, i_13_51_2768_0, i_13_51_2923_0,
    i_13_51_2924_0, i_13_51_2959_0, i_13_51_2965_0, i_13_51_3163_0,
    i_13_51_3373_0, i_13_51_3374_0, i_13_51_3419_0, i_13_51_3565_0,
    i_13_51_3580_0, i_13_51_3599_0, i_13_51_3650_0, i_13_51_3731_0,
    i_13_51_3733_0, i_13_51_3734_0, i_13_51_3787_0, i_13_51_3905_0,
    i_13_51_3910_0, i_13_51_3919_0, i_13_51_3923_0, i_13_51_3985_0,
    i_13_51_4253_0, i_13_51_4255_0, i_13_51_4256_0, i_13_51_4262_0,
    i_13_51_4265_0, i_13_51_4453_0, i_13_51_4454_0, i_13_51_4526_0,
    i_13_51_4541_0, i_13_51_4558_0, i_13_51_4559_0, i_13_51_4561_0;
  output o_13_51_0_0;
  assign o_13_51_0_0 = ~((~i_13_51_3923_0 & ~i_13_51_4559_0) | (~i_13_51_2546_0 & ~i_13_51_4454_0));
endmodule



// Benchmark "kernel_13_52" written by ABC on Sun Jul 19 10:46:08 2020

module kernel_13_52 ( 
    i_13_52_2_0, i_13_52_78_0, i_13_52_180_0, i_13_52_184_0, i_13_52_185_0,
    i_13_52_187_0, i_13_52_189_0, i_13_52_192_0, i_13_52_193_0,
    i_13_52_283_0, i_13_52_324_0, i_13_52_370_0, i_13_52_509_0,
    i_13_52_517_0, i_13_52_533_0, i_13_52_570_0, i_13_52_571_0,
    i_13_52_594_0, i_13_52_640_0, i_13_52_641_0, i_13_52_714_0,
    i_13_52_715_0, i_13_52_718_0, i_13_52_798_0, i_13_52_858_0,
    i_13_52_887_0, i_13_52_939_0, i_13_52_958_0, i_13_52_1116_0,
    i_13_52_1193_0, i_13_52_1219_0, i_13_52_1228_0, i_13_52_1229_0,
    i_13_52_1254_0, i_13_52_1299_0, i_13_52_1314_0, i_13_52_1407_0,
    i_13_52_1408_0, i_13_52_1435_0, i_13_52_1464_0, i_13_52_1479_0,
    i_13_52_1530_0, i_13_52_1597_0, i_13_52_1639_0, i_13_52_1674_0,
    i_13_52_1713_0, i_13_52_1732_0, i_13_52_1741_0, i_13_52_1761_0,
    i_13_52_1762_0, i_13_52_1764_0, i_13_52_1769_0, i_13_52_1782_0,
    i_13_52_1785_0, i_13_52_1786_0, i_13_52_1801_0, i_13_52_1804_0,
    i_13_52_1957_0, i_13_52_2017_0, i_13_52_2055_0, i_13_52_2210_0,
    i_13_52_2280_0, i_13_52_2365_0, i_13_52_2397_0, i_13_52_2502_0,
    i_13_52_2567_0, i_13_52_2619_0, i_13_52_2693_0, i_13_52_2713_0,
    i_13_52_2857_0, i_13_52_3025_0, i_13_52_3030_0, i_13_52_3034_0,
    i_13_52_3045_0, i_13_52_3046_0, i_13_52_3163_0, i_13_52_3168_0,
    i_13_52_3259_0, i_13_52_3265_0, i_13_52_3286_0, i_13_52_3287_0,
    i_13_52_3352_0, i_13_52_3403_0, i_13_52_3423_0, i_13_52_3424_0,
    i_13_52_3754_0, i_13_52_3756_0, i_13_52_3759_0, i_13_52_3972_0,
    i_13_52_3979_0, i_13_52_3981_0, i_13_52_3984_0, i_13_52_4042_0,
    i_13_52_4086_0, i_13_52_4187_0, i_13_52_4199_0, i_13_52_4363_0,
    i_13_52_4434_0, i_13_52_4537_0, i_13_52_4565_0,
    o_13_52_0_0  );
  input  i_13_52_2_0, i_13_52_78_0, i_13_52_180_0, i_13_52_184_0,
    i_13_52_185_0, i_13_52_187_0, i_13_52_189_0, i_13_52_192_0,
    i_13_52_193_0, i_13_52_283_0, i_13_52_324_0, i_13_52_370_0,
    i_13_52_509_0, i_13_52_517_0, i_13_52_533_0, i_13_52_570_0,
    i_13_52_571_0, i_13_52_594_0, i_13_52_640_0, i_13_52_641_0,
    i_13_52_714_0, i_13_52_715_0, i_13_52_718_0, i_13_52_798_0,
    i_13_52_858_0, i_13_52_887_0, i_13_52_939_0, i_13_52_958_0,
    i_13_52_1116_0, i_13_52_1193_0, i_13_52_1219_0, i_13_52_1228_0,
    i_13_52_1229_0, i_13_52_1254_0, i_13_52_1299_0, i_13_52_1314_0,
    i_13_52_1407_0, i_13_52_1408_0, i_13_52_1435_0, i_13_52_1464_0,
    i_13_52_1479_0, i_13_52_1530_0, i_13_52_1597_0, i_13_52_1639_0,
    i_13_52_1674_0, i_13_52_1713_0, i_13_52_1732_0, i_13_52_1741_0,
    i_13_52_1761_0, i_13_52_1762_0, i_13_52_1764_0, i_13_52_1769_0,
    i_13_52_1782_0, i_13_52_1785_0, i_13_52_1786_0, i_13_52_1801_0,
    i_13_52_1804_0, i_13_52_1957_0, i_13_52_2017_0, i_13_52_2055_0,
    i_13_52_2210_0, i_13_52_2280_0, i_13_52_2365_0, i_13_52_2397_0,
    i_13_52_2502_0, i_13_52_2567_0, i_13_52_2619_0, i_13_52_2693_0,
    i_13_52_2713_0, i_13_52_2857_0, i_13_52_3025_0, i_13_52_3030_0,
    i_13_52_3034_0, i_13_52_3045_0, i_13_52_3046_0, i_13_52_3163_0,
    i_13_52_3168_0, i_13_52_3259_0, i_13_52_3265_0, i_13_52_3286_0,
    i_13_52_3287_0, i_13_52_3352_0, i_13_52_3403_0, i_13_52_3423_0,
    i_13_52_3424_0, i_13_52_3754_0, i_13_52_3756_0, i_13_52_3759_0,
    i_13_52_3972_0, i_13_52_3979_0, i_13_52_3981_0, i_13_52_3984_0,
    i_13_52_4042_0, i_13_52_4086_0, i_13_52_4187_0, i_13_52_4199_0,
    i_13_52_4363_0, i_13_52_4434_0, i_13_52_4537_0, i_13_52_4565_0;
  output o_13_52_0_0;
  assign o_13_52_0_0 = ~((~i_13_52_3981_0 & (~i_13_52_1408_0 | (~i_13_52_1732_0 & i_13_52_3984_0))) | (~i_13_52_1408_0 & ((i_13_52_858_0 & ~i_13_52_4042_0) | (~i_13_52_1254_0 & i_13_52_4363_0))) | (~i_13_52_858_0 & i_13_52_1597_0 & i_13_52_2713_0) | (~i_13_52_1479_0 & ~i_13_52_3423_0 & ~i_13_52_3424_0) | (~i_13_52_1314_0 & ~i_13_52_1769_0 & ~i_13_52_3979_0 & ~i_13_52_3984_0) | (~i_13_52_192_0 & ~i_13_52_3287_0 & ~i_13_52_4565_0));
endmodule



// Benchmark "kernel_13_53" written by ABC on Sun Jul 19 10:46:09 2020

module kernel_13_53 ( 
    i_13_53_172_0, i_13_53_192_0, i_13_53_199_0, i_13_53_280_0,
    i_13_53_324_0, i_13_53_361_0, i_13_53_378_0, i_13_53_525_0,
    i_13_53_570_0, i_13_53_576_0, i_13_53_639_0, i_13_53_640_0,
    i_13_53_685_0, i_13_53_714_0, i_13_53_777_0, i_13_53_810_0,
    i_13_53_858_0, i_13_53_891_0, i_13_53_927_0, i_13_53_948_0,
    i_13_53_954_0, i_13_53_1020_0, i_13_53_1026_0, i_13_53_1059_0,
    i_13_53_1063_0, i_13_53_1098_0, i_13_53_1209_0, i_13_53_1224_0,
    i_13_53_1225_0, i_13_53_1227_0, i_13_53_1254_0, i_13_53_1263_0,
    i_13_53_1296_0, i_13_53_1297_0, i_13_53_1407_0, i_13_53_1443_0,
    i_13_53_1498_0, i_13_53_1539_0, i_13_53_1594_0, i_13_53_1632_0,
    i_13_53_1710_0, i_13_53_1719_0, i_13_53_1747_0, i_13_53_1767_0,
    i_13_53_1782_0, i_13_53_1792_0, i_13_53_1800_0, i_13_53_1801_0,
    i_13_53_1857_0, i_13_53_1881_0, i_13_53_1926_0, i_13_53_1990_0,
    i_13_53_2011_0, i_13_53_2100_0, i_13_53_2116_0, i_13_53_2259_0,
    i_13_53_2358_0, i_13_53_2403_0, i_13_53_2460_0, i_13_53_2514_0,
    i_13_53_2532_0, i_13_53_2629_0, i_13_53_2646_0, i_13_53_2844_0,
    i_13_53_2853_0, i_13_53_2899_0, i_13_53_2934_0, i_13_53_2980_0,
    i_13_53_3105_0, i_13_53_3171_0, i_13_53_3241_0, i_13_53_3259_0,
    i_13_53_3267_0, i_13_53_3268_0, i_13_53_3285_0, i_13_53_3286_0,
    i_13_53_3325_0, i_13_53_3420_0, i_13_53_3421_0, i_13_53_3423_0,
    i_13_53_3447_0, i_13_53_3790_0, i_13_53_3873_0, i_13_53_3970_0,
    i_13_53_3991_0, i_13_53_4008_0, i_13_53_4009_0, i_13_53_4041_0,
    i_13_53_4042_0, i_13_53_4077_0, i_13_53_4086_0, i_13_53_4087_0,
    i_13_53_4153_0, i_13_53_4231_0, i_13_53_4248_0, i_13_53_4267_0,
    i_13_53_4278_0, i_13_53_4293_0, i_13_53_4410_0, i_13_53_4584_0,
    o_13_53_0_0  );
  input  i_13_53_172_0, i_13_53_192_0, i_13_53_199_0, i_13_53_280_0,
    i_13_53_324_0, i_13_53_361_0, i_13_53_378_0, i_13_53_525_0,
    i_13_53_570_0, i_13_53_576_0, i_13_53_639_0, i_13_53_640_0,
    i_13_53_685_0, i_13_53_714_0, i_13_53_777_0, i_13_53_810_0,
    i_13_53_858_0, i_13_53_891_0, i_13_53_927_0, i_13_53_948_0,
    i_13_53_954_0, i_13_53_1020_0, i_13_53_1026_0, i_13_53_1059_0,
    i_13_53_1063_0, i_13_53_1098_0, i_13_53_1209_0, i_13_53_1224_0,
    i_13_53_1225_0, i_13_53_1227_0, i_13_53_1254_0, i_13_53_1263_0,
    i_13_53_1296_0, i_13_53_1297_0, i_13_53_1407_0, i_13_53_1443_0,
    i_13_53_1498_0, i_13_53_1539_0, i_13_53_1594_0, i_13_53_1632_0,
    i_13_53_1710_0, i_13_53_1719_0, i_13_53_1747_0, i_13_53_1767_0,
    i_13_53_1782_0, i_13_53_1792_0, i_13_53_1800_0, i_13_53_1801_0,
    i_13_53_1857_0, i_13_53_1881_0, i_13_53_1926_0, i_13_53_1990_0,
    i_13_53_2011_0, i_13_53_2100_0, i_13_53_2116_0, i_13_53_2259_0,
    i_13_53_2358_0, i_13_53_2403_0, i_13_53_2460_0, i_13_53_2514_0,
    i_13_53_2532_0, i_13_53_2629_0, i_13_53_2646_0, i_13_53_2844_0,
    i_13_53_2853_0, i_13_53_2899_0, i_13_53_2934_0, i_13_53_2980_0,
    i_13_53_3105_0, i_13_53_3171_0, i_13_53_3241_0, i_13_53_3259_0,
    i_13_53_3267_0, i_13_53_3268_0, i_13_53_3285_0, i_13_53_3286_0,
    i_13_53_3325_0, i_13_53_3420_0, i_13_53_3421_0, i_13_53_3423_0,
    i_13_53_3447_0, i_13_53_3790_0, i_13_53_3873_0, i_13_53_3970_0,
    i_13_53_3991_0, i_13_53_4008_0, i_13_53_4009_0, i_13_53_4041_0,
    i_13_53_4042_0, i_13_53_4077_0, i_13_53_4086_0, i_13_53_4087_0,
    i_13_53_4153_0, i_13_53_4231_0, i_13_53_4248_0, i_13_53_4267_0,
    i_13_53_4278_0, i_13_53_4293_0, i_13_53_4410_0, i_13_53_4584_0;
  output o_13_53_0_0;
  assign o_13_53_0_0 = ~((~i_13_53_685_0 & ~i_13_53_1926_0) | (~i_13_53_1407_0 & i_13_53_1857_0 & ~i_13_53_3421_0) | (~i_13_53_378_0 & ~i_13_53_891_0 & ~i_13_53_3241_0 & ~i_13_53_4248_0) | (~i_13_53_1254_0 & ~i_13_53_3420_0 & ~i_13_53_4086_0 & ~i_13_53_4267_0 & ~i_13_53_4410_0) | (~i_13_53_1800_0 & ~i_13_53_2403_0 & ~i_13_53_3285_0 & ~i_13_53_3873_0 & ~i_13_53_4009_0));
endmodule



// Benchmark "kernel_13_54" written by ABC on Sun Jul 19 10:46:10 2020

module kernel_13_54 ( 
    i_13_54_31_0, i_13_54_58_0, i_13_54_67_0, i_13_54_130_0, i_13_54_139_0,
    i_13_54_183_0, i_13_54_184_0, i_13_54_192_0, i_13_54_219_0,
    i_13_54_255_0, i_13_54_361_0, i_13_54_373_0, i_13_54_382_0,
    i_13_54_390_0, i_13_54_549_0, i_13_54_624_0, i_13_54_685_0,
    i_13_54_717_0, i_13_54_777_0, i_13_54_822_0, i_13_54_891_0,
    i_13_54_894_0, i_13_54_897_0, i_13_54_975_0, i_13_54_976_0,
    i_13_54_1093_0, i_13_54_1108_0, i_13_54_1116_0, i_13_54_1120_0,
    i_13_54_1145_0, i_13_54_1308_0, i_13_54_1314_0, i_13_54_1345_0,
    i_13_54_1380_0, i_13_54_1386_0, i_13_54_1387_0, i_13_54_1393_0,
    i_13_54_1407_0, i_13_54_1461_0, i_13_54_1476_0, i_13_54_1479_0,
    i_13_54_1480_0, i_13_54_1487_0, i_13_54_1498_0, i_13_54_1513_0,
    i_13_54_1526_0, i_13_54_1585_0, i_13_54_1597_0, i_13_54_1669_0,
    i_13_54_1674_0, i_13_54_1677_0, i_13_54_1690_0, i_13_54_1731_0,
    i_13_54_1749_0, i_13_54_1752_0, i_13_54_1756_0, i_13_54_1803_0,
    i_13_54_1956_0, i_13_54_2017_0, i_13_54_2190_0, i_13_54_2191_0,
    i_13_54_2442_0, i_13_54_2443_0, i_13_54_2449_0, i_13_54_2461_0,
    i_13_54_2479_0, i_13_54_2539_0, i_13_54_2559_0, i_13_54_2632_0,
    i_13_54_2676_0, i_13_54_2686_0, i_13_54_2739_0, i_13_54_2751_0,
    i_13_54_2895_0, i_13_54_2967_0, i_13_54_2997_0, i_13_54_3001_0,
    i_13_54_3114_0, i_13_54_3199_0, i_13_54_3261_0, i_13_54_3348_0,
    i_13_54_3352_0, i_13_54_3433_0, i_13_54_3468_0, i_13_54_3478_0,
    i_13_54_3520_0, i_13_54_3522_0, i_13_54_3525_0, i_13_54_3561_0,
    i_13_54_3567_0, i_13_54_3756_0, i_13_54_3865_0, i_13_54_3981_0,
    i_13_54_4294_0, i_13_54_4348_0, i_13_54_4351_0, i_13_54_4363_0,
    i_13_54_4413_0, i_13_54_4532_0, i_13_54_4591_0,
    o_13_54_0_0  );
  input  i_13_54_31_0, i_13_54_58_0, i_13_54_67_0, i_13_54_130_0,
    i_13_54_139_0, i_13_54_183_0, i_13_54_184_0, i_13_54_192_0,
    i_13_54_219_0, i_13_54_255_0, i_13_54_361_0, i_13_54_373_0,
    i_13_54_382_0, i_13_54_390_0, i_13_54_549_0, i_13_54_624_0,
    i_13_54_685_0, i_13_54_717_0, i_13_54_777_0, i_13_54_822_0,
    i_13_54_891_0, i_13_54_894_0, i_13_54_897_0, i_13_54_975_0,
    i_13_54_976_0, i_13_54_1093_0, i_13_54_1108_0, i_13_54_1116_0,
    i_13_54_1120_0, i_13_54_1145_0, i_13_54_1308_0, i_13_54_1314_0,
    i_13_54_1345_0, i_13_54_1380_0, i_13_54_1386_0, i_13_54_1387_0,
    i_13_54_1393_0, i_13_54_1407_0, i_13_54_1461_0, i_13_54_1476_0,
    i_13_54_1479_0, i_13_54_1480_0, i_13_54_1487_0, i_13_54_1498_0,
    i_13_54_1513_0, i_13_54_1526_0, i_13_54_1585_0, i_13_54_1597_0,
    i_13_54_1669_0, i_13_54_1674_0, i_13_54_1677_0, i_13_54_1690_0,
    i_13_54_1731_0, i_13_54_1749_0, i_13_54_1752_0, i_13_54_1756_0,
    i_13_54_1803_0, i_13_54_1956_0, i_13_54_2017_0, i_13_54_2190_0,
    i_13_54_2191_0, i_13_54_2442_0, i_13_54_2443_0, i_13_54_2449_0,
    i_13_54_2461_0, i_13_54_2479_0, i_13_54_2539_0, i_13_54_2559_0,
    i_13_54_2632_0, i_13_54_2676_0, i_13_54_2686_0, i_13_54_2739_0,
    i_13_54_2751_0, i_13_54_2895_0, i_13_54_2967_0, i_13_54_2997_0,
    i_13_54_3001_0, i_13_54_3114_0, i_13_54_3199_0, i_13_54_3261_0,
    i_13_54_3348_0, i_13_54_3352_0, i_13_54_3433_0, i_13_54_3468_0,
    i_13_54_3478_0, i_13_54_3520_0, i_13_54_3522_0, i_13_54_3525_0,
    i_13_54_3561_0, i_13_54_3567_0, i_13_54_3756_0, i_13_54_3865_0,
    i_13_54_3981_0, i_13_54_4294_0, i_13_54_4348_0, i_13_54_4351_0,
    i_13_54_4363_0, i_13_54_4413_0, i_13_54_4532_0, i_13_54_4591_0;
  output o_13_54_0_0;
  assign o_13_54_0_0 = ~((~i_13_54_822_0 & ((~i_13_54_1345_0 & ~i_13_54_1677_0) | (i_13_54_2461_0 & i_13_54_4413_0))) | (~i_13_54_1479_0 & (~i_13_54_2017_0 | ~i_13_54_3522_0)) | (i_13_54_4351_0 & ((~i_13_54_1674_0 & ~i_13_54_1803_0) | (~i_13_54_3520_0 & ~i_13_54_3567_0 & ~i_13_54_4363_0))) | (~i_13_54_255_0 & ~i_13_54_1308_0 & ~i_13_54_2676_0) | (~i_13_54_891_0 & ~i_13_54_897_0 & ~i_13_54_2539_0 & ~i_13_54_3522_0));
endmodule



// Benchmark "kernel_13_55" written by ABC on Sun Jul 19 10:46:11 2020

module kernel_13_55 ( 
    i_13_55_47_0, i_13_55_92_0, i_13_55_94_0, i_13_55_95_0, i_13_55_139_0,
    i_13_55_170_0, i_13_55_173_0, i_13_55_175_0, i_13_55_178_0,
    i_13_55_214_0, i_13_55_215_0, i_13_55_311_0, i_13_55_362_0,
    i_13_55_441_0, i_13_55_452_0, i_13_55_535_0, i_13_55_555_0,
    i_13_55_569_0, i_13_55_571_0, i_13_55_572_0, i_13_55_609_0,
    i_13_55_659_0, i_13_55_662_0, i_13_55_686_0, i_13_55_847_0,
    i_13_55_851_0, i_13_55_854_0, i_13_55_951_0, i_13_55_956_0,
    i_13_55_986_0, i_13_55_1120_0, i_13_55_1229_0, i_13_55_1250_0,
    i_13_55_1260_0, i_13_55_1307_0, i_13_55_1311_0, i_13_55_1408_0,
    i_13_55_1422_0, i_13_55_1513_0, i_13_55_1514_0, i_13_55_1527_0,
    i_13_55_1540_0, i_13_55_1567_0, i_13_55_1723_0, i_13_55_1766_0,
    i_13_55_1791_0, i_13_55_1802_0, i_13_55_1829_0, i_13_55_1832_0,
    i_13_55_1847_0, i_13_55_1850_0, i_13_55_1858_0, i_13_55_1885_0,
    i_13_55_2108_0, i_13_55_2150_0, i_13_55_2227_0, i_13_55_2234_0,
    i_13_55_2297_0, i_13_55_2410_0, i_13_55_2467_0, i_13_55_2677_0,
    i_13_55_2680_0, i_13_55_2696_0, i_13_55_2713_0, i_13_55_2740_0,
    i_13_55_2934_0, i_13_55_2980_0, i_13_55_2985_0, i_13_55_3007_0,
    i_13_55_3011_0, i_13_55_3012_0, i_13_55_3025_0, i_13_55_3026_0,
    i_13_55_3064_0, i_13_55_3109_0, i_13_55_3110_0, i_13_55_3113_0,
    i_13_55_3208_0, i_13_55_3217_0, i_13_55_3268_0, i_13_55_3269_0,
    i_13_55_3386_0, i_13_55_3519_0, i_13_55_3739_0, i_13_55_3755_0,
    i_13_55_3764_0, i_13_55_3818_0, i_13_55_3879_0, i_13_55_3987_0,
    i_13_55_4061_0, i_13_55_4064_0, i_13_55_4371_0, i_13_55_4375_0,
    i_13_55_4432_0, i_13_55_4472_0, i_13_55_4514_0, i_13_55_4565_0,
    i_13_55_4568_0, i_13_55_4569_0, i_13_55_4591_0,
    o_13_55_0_0  );
  input  i_13_55_47_0, i_13_55_92_0, i_13_55_94_0, i_13_55_95_0,
    i_13_55_139_0, i_13_55_170_0, i_13_55_173_0, i_13_55_175_0,
    i_13_55_178_0, i_13_55_214_0, i_13_55_215_0, i_13_55_311_0,
    i_13_55_362_0, i_13_55_441_0, i_13_55_452_0, i_13_55_535_0,
    i_13_55_555_0, i_13_55_569_0, i_13_55_571_0, i_13_55_572_0,
    i_13_55_609_0, i_13_55_659_0, i_13_55_662_0, i_13_55_686_0,
    i_13_55_847_0, i_13_55_851_0, i_13_55_854_0, i_13_55_951_0,
    i_13_55_956_0, i_13_55_986_0, i_13_55_1120_0, i_13_55_1229_0,
    i_13_55_1250_0, i_13_55_1260_0, i_13_55_1307_0, i_13_55_1311_0,
    i_13_55_1408_0, i_13_55_1422_0, i_13_55_1513_0, i_13_55_1514_0,
    i_13_55_1527_0, i_13_55_1540_0, i_13_55_1567_0, i_13_55_1723_0,
    i_13_55_1766_0, i_13_55_1791_0, i_13_55_1802_0, i_13_55_1829_0,
    i_13_55_1832_0, i_13_55_1847_0, i_13_55_1850_0, i_13_55_1858_0,
    i_13_55_1885_0, i_13_55_2108_0, i_13_55_2150_0, i_13_55_2227_0,
    i_13_55_2234_0, i_13_55_2297_0, i_13_55_2410_0, i_13_55_2467_0,
    i_13_55_2677_0, i_13_55_2680_0, i_13_55_2696_0, i_13_55_2713_0,
    i_13_55_2740_0, i_13_55_2934_0, i_13_55_2980_0, i_13_55_2985_0,
    i_13_55_3007_0, i_13_55_3011_0, i_13_55_3012_0, i_13_55_3025_0,
    i_13_55_3026_0, i_13_55_3064_0, i_13_55_3109_0, i_13_55_3110_0,
    i_13_55_3113_0, i_13_55_3208_0, i_13_55_3217_0, i_13_55_3268_0,
    i_13_55_3269_0, i_13_55_3386_0, i_13_55_3519_0, i_13_55_3739_0,
    i_13_55_3755_0, i_13_55_3764_0, i_13_55_3818_0, i_13_55_3879_0,
    i_13_55_3987_0, i_13_55_4061_0, i_13_55_4064_0, i_13_55_4371_0,
    i_13_55_4375_0, i_13_55_4432_0, i_13_55_4472_0, i_13_55_4514_0,
    i_13_55_4565_0, i_13_55_4568_0, i_13_55_4569_0, i_13_55_4591_0;
  output o_13_55_0_0;
  assign o_13_55_0_0 = ~(~i_13_55_173_0 | (~i_13_55_2980_0 & ~i_13_55_3755_0) | (i_13_55_94_0 & ~i_13_55_1567_0 & ~i_13_55_3109_0 & ~i_13_55_4064_0));
endmodule



// Benchmark "kernel_13_56" written by ABC on Sun Jul 19 10:46:12 2020

module kernel_13_56 ( 
    i_13_56_40_0, i_13_56_76_0, i_13_56_133_0, i_13_56_192_0,
    i_13_56_251_0, i_13_56_283_0, i_13_56_318_0, i_13_56_334_0,
    i_13_56_336_0, i_13_56_358_0, i_13_56_457_0, i_13_56_492_0,
    i_13_56_493_0, i_13_56_620_0, i_13_56_715_0, i_13_56_758_0,
    i_13_56_813_0, i_13_56_829_0, i_13_56_876_0, i_13_56_956_0,
    i_13_56_1025_0, i_13_56_1100_0, i_13_56_1102_0, i_13_56_1230_0,
    i_13_56_1257_0, i_13_56_1300_0, i_13_56_1303_0, i_13_56_1327_0,
    i_13_56_1405_0, i_13_56_1446_0, i_13_56_1447_0, i_13_56_1502_0,
    i_13_56_1525_0, i_13_56_1640_0, i_13_56_1641_0, i_13_56_1698_0,
    i_13_56_1722_0, i_13_56_1723_0, i_13_56_1742_0, i_13_56_1785_0,
    i_13_56_1793_0, i_13_56_1794_0, i_13_56_1835_0, i_13_56_1937_0,
    i_13_56_2014_0, i_13_56_2056_0, i_13_56_2060_0, i_13_56_2103_0,
    i_13_56_2118_0, i_13_56_2146_0, i_13_56_2185_0, i_13_56_2236_0,
    i_13_56_2237_0, i_13_56_2239_0, i_13_56_2365_0, i_13_56_2407_0,
    i_13_56_2427_0, i_13_56_2445_0, i_13_56_2452_0, i_13_56_2535_0,
    i_13_56_2587_0, i_13_56_2617_0, i_13_56_2721_0, i_13_56_2922_0,
    i_13_56_2924_0, i_13_56_2937_0, i_13_56_3032_0, i_13_56_3036_0,
    i_13_56_3217_0, i_13_56_3219_0, i_13_56_3220_0, i_13_56_3234_0,
    i_13_56_3243_0, i_13_56_3244_0, i_13_56_3343_0, i_13_56_3424_0,
    i_13_56_3480_0, i_13_56_3550_0, i_13_56_3639_0, i_13_56_3649_0,
    i_13_56_3700_0, i_13_56_3702_0, i_13_56_3757_0, i_13_56_3766_0,
    i_13_56_3846_0, i_13_56_3865_0, i_13_56_3878_0, i_13_56_3889_0,
    i_13_56_3984_0, i_13_56_3985_0, i_13_56_4054_0, i_13_56_4213_0,
    i_13_56_4237_0, i_13_56_4273_0, i_13_56_4315_0, i_13_56_4400_0,
    i_13_56_4510_0, i_13_56_4513_0, i_13_56_4561_0, i_13_56_4587_0,
    o_13_56_0_0  );
  input  i_13_56_40_0, i_13_56_76_0, i_13_56_133_0, i_13_56_192_0,
    i_13_56_251_0, i_13_56_283_0, i_13_56_318_0, i_13_56_334_0,
    i_13_56_336_0, i_13_56_358_0, i_13_56_457_0, i_13_56_492_0,
    i_13_56_493_0, i_13_56_620_0, i_13_56_715_0, i_13_56_758_0,
    i_13_56_813_0, i_13_56_829_0, i_13_56_876_0, i_13_56_956_0,
    i_13_56_1025_0, i_13_56_1100_0, i_13_56_1102_0, i_13_56_1230_0,
    i_13_56_1257_0, i_13_56_1300_0, i_13_56_1303_0, i_13_56_1327_0,
    i_13_56_1405_0, i_13_56_1446_0, i_13_56_1447_0, i_13_56_1502_0,
    i_13_56_1525_0, i_13_56_1640_0, i_13_56_1641_0, i_13_56_1698_0,
    i_13_56_1722_0, i_13_56_1723_0, i_13_56_1742_0, i_13_56_1785_0,
    i_13_56_1793_0, i_13_56_1794_0, i_13_56_1835_0, i_13_56_1937_0,
    i_13_56_2014_0, i_13_56_2056_0, i_13_56_2060_0, i_13_56_2103_0,
    i_13_56_2118_0, i_13_56_2146_0, i_13_56_2185_0, i_13_56_2236_0,
    i_13_56_2237_0, i_13_56_2239_0, i_13_56_2365_0, i_13_56_2407_0,
    i_13_56_2427_0, i_13_56_2445_0, i_13_56_2452_0, i_13_56_2535_0,
    i_13_56_2587_0, i_13_56_2617_0, i_13_56_2721_0, i_13_56_2922_0,
    i_13_56_2924_0, i_13_56_2937_0, i_13_56_3032_0, i_13_56_3036_0,
    i_13_56_3217_0, i_13_56_3219_0, i_13_56_3220_0, i_13_56_3234_0,
    i_13_56_3243_0, i_13_56_3244_0, i_13_56_3343_0, i_13_56_3424_0,
    i_13_56_3480_0, i_13_56_3550_0, i_13_56_3639_0, i_13_56_3649_0,
    i_13_56_3700_0, i_13_56_3702_0, i_13_56_3757_0, i_13_56_3766_0,
    i_13_56_3846_0, i_13_56_3865_0, i_13_56_3878_0, i_13_56_3889_0,
    i_13_56_3984_0, i_13_56_3985_0, i_13_56_4054_0, i_13_56_4213_0,
    i_13_56_4237_0, i_13_56_4273_0, i_13_56_4315_0, i_13_56_4400_0,
    i_13_56_4510_0, i_13_56_4513_0, i_13_56_4561_0, i_13_56_4587_0;
  output o_13_56_0_0;
  assign o_13_56_0_0 = ~((~i_13_56_3984_0 & ((~i_13_56_2427_0 & ((~i_13_56_3550_0 & ~i_13_56_3757_0) | (~i_13_56_620_0 & ~i_13_56_2445_0 & ~i_13_56_2924_0 & ~i_13_56_3878_0))) | (i_13_56_283_0 & ~i_13_56_4315_0))) | (~i_13_56_1300_0 & ~i_13_56_1525_0 & i_13_56_2185_0) | ~i_13_56_3985_0 | (i_13_56_2237_0 & i_13_56_4561_0));
endmodule



// Benchmark "kernel_13_57" written by ABC on Sun Jul 19 10:46:12 2020

module kernel_13_57 ( 
    i_13_57_63_0, i_13_57_76_0, i_13_57_136_0, i_13_57_339_0,
    i_13_57_340_0, i_13_57_357_0, i_13_57_358_0, i_13_57_534_0,
    i_13_57_535_0, i_13_57_546_0, i_13_57_579_0, i_13_57_645_0,
    i_13_57_687_0, i_13_57_690_0, i_13_57_697_0, i_13_57_825_0,
    i_13_57_915_0, i_13_57_1066_0, i_13_57_1213_0, i_13_57_1303_0,
    i_13_57_1306_0, i_13_57_1321_0, i_13_57_1347_0, i_13_57_1383_0,
    i_13_57_1446_0, i_13_57_1465_0, i_13_57_1501_0, i_13_57_1518_0,
    i_13_57_1642_0, i_13_57_1722_0, i_13_57_1723_0, i_13_57_1740_0,
    i_13_57_1815_0, i_13_57_1845_0, i_13_57_1950_0, i_13_57_1951_0,
    i_13_57_1960_0, i_13_57_2005_0, i_13_57_2023_0, i_13_57_2032_0,
    i_13_57_2058_0, i_13_57_2106_0, i_13_57_2110_0, i_13_57_2320_0,
    i_13_57_2428_0, i_13_57_2446_0, i_13_57_2514_0, i_13_57_2554_0,
    i_13_57_2640_0, i_13_57_2644_0, i_13_57_2649_0, i_13_57_2652_0,
    i_13_57_2677_0, i_13_57_2692_0, i_13_57_2751_0, i_13_57_2763_0,
    i_13_57_2847_0, i_13_57_2848_0, i_13_57_2913_0, i_13_57_2920_0,
    i_13_57_2922_0, i_13_57_2923_0, i_13_57_2958_0, i_13_57_2962_0,
    i_13_57_3028_0, i_13_57_3144_0, i_13_57_3219_0, i_13_57_3372_0,
    i_13_57_3373_0, i_13_57_3391_0, i_13_57_3393_0, i_13_57_3418_0,
    i_13_57_3444_0, i_13_57_3577_0, i_13_57_3595_0, i_13_57_3597_0,
    i_13_57_3598_0, i_13_57_3621_0, i_13_57_3669_0, i_13_57_3721_0,
    i_13_57_3741_0, i_13_57_3787_0, i_13_57_3793_0, i_13_57_3928_0,
    i_13_57_3990_0, i_13_57_3991_0, i_13_57_4021_0, i_13_57_4191_0,
    i_13_57_4237_0, i_13_57_4263_0, i_13_57_4264_0, i_13_57_4315_0,
    i_13_57_4332_0, i_13_57_4333_0, i_13_57_4350_0, i_13_57_4381_0,
    i_13_57_4398_0, i_13_57_4435_0, i_13_57_4452_0, i_13_57_4453_0,
    o_13_57_0_0  );
  input  i_13_57_63_0, i_13_57_76_0, i_13_57_136_0, i_13_57_339_0,
    i_13_57_340_0, i_13_57_357_0, i_13_57_358_0, i_13_57_534_0,
    i_13_57_535_0, i_13_57_546_0, i_13_57_579_0, i_13_57_645_0,
    i_13_57_687_0, i_13_57_690_0, i_13_57_697_0, i_13_57_825_0,
    i_13_57_915_0, i_13_57_1066_0, i_13_57_1213_0, i_13_57_1303_0,
    i_13_57_1306_0, i_13_57_1321_0, i_13_57_1347_0, i_13_57_1383_0,
    i_13_57_1446_0, i_13_57_1465_0, i_13_57_1501_0, i_13_57_1518_0,
    i_13_57_1642_0, i_13_57_1722_0, i_13_57_1723_0, i_13_57_1740_0,
    i_13_57_1815_0, i_13_57_1845_0, i_13_57_1950_0, i_13_57_1951_0,
    i_13_57_1960_0, i_13_57_2005_0, i_13_57_2023_0, i_13_57_2032_0,
    i_13_57_2058_0, i_13_57_2106_0, i_13_57_2110_0, i_13_57_2320_0,
    i_13_57_2428_0, i_13_57_2446_0, i_13_57_2514_0, i_13_57_2554_0,
    i_13_57_2640_0, i_13_57_2644_0, i_13_57_2649_0, i_13_57_2652_0,
    i_13_57_2677_0, i_13_57_2692_0, i_13_57_2751_0, i_13_57_2763_0,
    i_13_57_2847_0, i_13_57_2848_0, i_13_57_2913_0, i_13_57_2920_0,
    i_13_57_2922_0, i_13_57_2923_0, i_13_57_2958_0, i_13_57_2962_0,
    i_13_57_3028_0, i_13_57_3144_0, i_13_57_3219_0, i_13_57_3372_0,
    i_13_57_3373_0, i_13_57_3391_0, i_13_57_3393_0, i_13_57_3418_0,
    i_13_57_3444_0, i_13_57_3577_0, i_13_57_3595_0, i_13_57_3597_0,
    i_13_57_3598_0, i_13_57_3621_0, i_13_57_3669_0, i_13_57_3721_0,
    i_13_57_3741_0, i_13_57_3787_0, i_13_57_3793_0, i_13_57_3928_0,
    i_13_57_3990_0, i_13_57_3991_0, i_13_57_4021_0, i_13_57_4191_0,
    i_13_57_4237_0, i_13_57_4263_0, i_13_57_4264_0, i_13_57_4315_0,
    i_13_57_4332_0, i_13_57_4333_0, i_13_57_4350_0, i_13_57_4381_0,
    i_13_57_4398_0, i_13_57_4435_0, i_13_57_4452_0, i_13_57_4453_0;
  output o_13_57_0_0;
  assign o_13_57_0_0 = ~((i_13_57_3595_0 & ~i_13_57_4237_0) | (i_13_57_2110_0 & ~i_13_57_3597_0) | (~i_13_57_690_0 & ~i_13_57_1951_0 & ~i_13_57_4452_0) | (~i_13_57_535_0 & ~i_13_57_1960_0 & ~i_13_57_4315_0));
endmodule



// Benchmark "kernel_13_58" written by ABC on Sun Jul 19 10:46:13 2020

module kernel_13_58 ( 
    i_13_58_42_0, i_13_58_78_0, i_13_58_111_0, i_13_58_194_0,
    i_13_58_199_0, i_13_58_276_0, i_13_58_282_0, i_13_58_285_0,
    i_13_58_310_0, i_13_58_384_0, i_13_58_417_0, i_13_58_418_0,
    i_13_58_448_0, i_13_58_519_0, i_13_58_520_0, i_13_58_535_0,
    i_13_58_553_0, i_13_58_643_0, i_13_58_670_0, i_13_58_838_0,
    i_13_58_873_0, i_13_58_935_0, i_13_58_952_0, i_13_58_1020_0,
    i_13_58_1021_0, i_13_58_1023_0, i_13_58_1024_0, i_13_58_1075_0,
    i_13_58_1203_0, i_13_58_1254_0, i_13_58_1317_0, i_13_58_1390_0,
    i_13_58_1428_0, i_13_58_1429_0, i_13_58_1600_0, i_13_58_1605_0,
    i_13_58_1626_0, i_13_58_1632_0, i_13_58_1642_0, i_13_58_1777_0,
    i_13_58_1779_0, i_13_58_1780_0, i_13_58_1807_0, i_13_58_1813_0,
    i_13_58_1933_0, i_13_58_1940_0, i_13_58_2159_0, i_13_58_2199_0,
    i_13_58_2356_0, i_13_58_2454_0, i_13_58_2464_0, i_13_58_2541_0,
    i_13_58_2542_0, i_13_58_2575_0, i_13_58_2583_0, i_13_58_2617_0,
    i_13_58_2708_0, i_13_58_2769_0, i_13_58_2770_0, i_13_58_2847_0,
    i_13_58_2904_0, i_13_58_2919_0, i_13_58_2920_0, i_13_58_3031_0,
    i_13_58_3045_0, i_13_58_3246_0, i_13_58_3261_0, i_13_58_3353_0,
    i_13_58_3415_0, i_13_58_3453_0, i_13_58_3454_0, i_13_58_3456_0,
    i_13_58_3457_0, i_13_58_3459_0, i_13_58_3460_0, i_13_58_3462_0,
    i_13_58_3463_0, i_13_58_3534_0, i_13_58_3535_0, i_13_58_3541_0,
    i_13_58_3544_0, i_13_58_3558_0, i_13_58_3576_0, i_13_58_3619_0,
    i_13_58_3739_0, i_13_58_3783_0, i_13_58_3822_0, i_13_58_3868_0,
    i_13_58_3927_0, i_13_58_3975_0, i_13_58_3999_0, i_13_58_4080_0,
    i_13_58_4081_0, i_13_58_4252_0, i_13_58_4254_0, i_13_58_4255_0,
    i_13_58_4371_0, i_13_58_4449_0, i_13_58_4450_0, i_13_58_4602_0,
    o_13_58_0_0  );
  input  i_13_58_42_0, i_13_58_78_0, i_13_58_111_0, i_13_58_194_0,
    i_13_58_199_0, i_13_58_276_0, i_13_58_282_0, i_13_58_285_0,
    i_13_58_310_0, i_13_58_384_0, i_13_58_417_0, i_13_58_418_0,
    i_13_58_448_0, i_13_58_519_0, i_13_58_520_0, i_13_58_535_0,
    i_13_58_553_0, i_13_58_643_0, i_13_58_670_0, i_13_58_838_0,
    i_13_58_873_0, i_13_58_935_0, i_13_58_952_0, i_13_58_1020_0,
    i_13_58_1021_0, i_13_58_1023_0, i_13_58_1024_0, i_13_58_1075_0,
    i_13_58_1203_0, i_13_58_1254_0, i_13_58_1317_0, i_13_58_1390_0,
    i_13_58_1428_0, i_13_58_1429_0, i_13_58_1600_0, i_13_58_1605_0,
    i_13_58_1626_0, i_13_58_1632_0, i_13_58_1642_0, i_13_58_1777_0,
    i_13_58_1779_0, i_13_58_1780_0, i_13_58_1807_0, i_13_58_1813_0,
    i_13_58_1933_0, i_13_58_1940_0, i_13_58_2159_0, i_13_58_2199_0,
    i_13_58_2356_0, i_13_58_2454_0, i_13_58_2464_0, i_13_58_2541_0,
    i_13_58_2542_0, i_13_58_2575_0, i_13_58_2583_0, i_13_58_2617_0,
    i_13_58_2708_0, i_13_58_2769_0, i_13_58_2770_0, i_13_58_2847_0,
    i_13_58_2904_0, i_13_58_2919_0, i_13_58_2920_0, i_13_58_3031_0,
    i_13_58_3045_0, i_13_58_3246_0, i_13_58_3261_0, i_13_58_3353_0,
    i_13_58_3415_0, i_13_58_3453_0, i_13_58_3454_0, i_13_58_3456_0,
    i_13_58_3457_0, i_13_58_3459_0, i_13_58_3460_0, i_13_58_3462_0,
    i_13_58_3463_0, i_13_58_3534_0, i_13_58_3535_0, i_13_58_3541_0,
    i_13_58_3544_0, i_13_58_3558_0, i_13_58_3576_0, i_13_58_3619_0,
    i_13_58_3739_0, i_13_58_3783_0, i_13_58_3822_0, i_13_58_3868_0,
    i_13_58_3927_0, i_13_58_3975_0, i_13_58_3999_0, i_13_58_4080_0,
    i_13_58_4081_0, i_13_58_4252_0, i_13_58_4254_0, i_13_58_4255_0,
    i_13_58_4371_0, i_13_58_4449_0, i_13_58_4450_0, i_13_58_4602_0;
  output o_13_58_0_0;
  assign o_13_58_0_0 = ~((~i_13_58_3535_0 & ~i_13_58_3822_0) | (~i_13_58_1024_0 & ~i_13_58_1428_0) | (~i_13_58_78_0 & ~i_13_58_520_0 & ~i_13_58_4449_0) | (~i_13_58_276_0 & ~i_13_58_1642_0 & ~i_13_58_3783_0));
endmodule



// Benchmark "kernel_13_59" written by ABC on Sun Jul 19 10:46:14 2020

module kernel_13_59 ( 
    i_13_59_33_0, i_13_59_61_0, i_13_59_192_0, i_13_59_195_0,
    i_13_59_205_0, i_13_59_253_0, i_13_59_260_0, i_13_59_282_0,
    i_13_59_309_0, i_13_59_310_0, i_13_59_375_0, i_13_59_382_0,
    i_13_59_463_0, i_13_59_466_0, i_13_59_578_0, i_13_59_589_0,
    i_13_59_617_0, i_13_59_618_0, i_13_59_619_0, i_13_59_624_0,
    i_13_59_625_0, i_13_59_672_0, i_13_59_673_0, i_13_59_760_0,
    i_13_59_768_0, i_13_59_816_0, i_13_59_942_0, i_13_59_976_0,
    i_13_59_979_0, i_13_59_1023_0, i_13_59_1081_0, i_13_59_1082_0,
    i_13_59_1087_0, i_13_59_1088_0, i_13_59_1096_0, i_13_59_1106_0,
    i_13_59_1147_0, i_13_59_1214_0, i_13_59_1270_0, i_13_59_1282_0,
    i_13_59_1309_0, i_13_59_1411_0, i_13_59_1514_0, i_13_59_1518_0,
    i_13_59_1561_0, i_13_59_1597_0, i_13_59_1680_0, i_13_59_1734_0,
    i_13_59_1741_0, i_13_59_1780_0, i_13_59_1849_0, i_13_59_1860_0,
    i_13_59_2002_0, i_13_59_2056_0, i_13_59_2191_0, i_13_59_2225_0,
    i_13_59_2383_0, i_13_59_2622_0, i_13_59_2769_0, i_13_59_2851_0,
    i_13_59_2878_0, i_13_59_2887_0, i_13_59_2907_0, i_13_59_2959_0,
    i_13_59_3028_0, i_13_59_3049_0, i_13_59_3113_0, i_13_59_3118_0,
    i_13_59_3156_0, i_13_59_3349_0, i_13_59_3352_0, i_13_59_3355_0,
    i_13_59_3382_0, i_13_59_3464_0, i_13_59_3534_0, i_13_59_3552_0,
    i_13_59_3571_0, i_13_59_3667_0, i_13_59_3730_0, i_13_59_3742_0,
    i_13_59_3984_0, i_13_59_3994_0, i_13_59_4063_0, i_13_59_4070_0,
    i_13_59_4108_0, i_13_59_4128_0, i_13_59_4155_0, i_13_59_4162_0,
    i_13_59_4165_0, i_13_59_4187_0, i_13_59_4299_0, i_13_59_4325_0,
    i_13_59_4335_0, i_13_59_4363_0, i_13_59_4369_0, i_13_59_4372_0,
    i_13_59_4418_0, i_13_59_4434_0, i_13_59_4532_0, i_13_59_4539_0,
    o_13_59_0_0  );
  input  i_13_59_33_0, i_13_59_61_0, i_13_59_192_0, i_13_59_195_0,
    i_13_59_205_0, i_13_59_253_0, i_13_59_260_0, i_13_59_282_0,
    i_13_59_309_0, i_13_59_310_0, i_13_59_375_0, i_13_59_382_0,
    i_13_59_463_0, i_13_59_466_0, i_13_59_578_0, i_13_59_589_0,
    i_13_59_617_0, i_13_59_618_0, i_13_59_619_0, i_13_59_624_0,
    i_13_59_625_0, i_13_59_672_0, i_13_59_673_0, i_13_59_760_0,
    i_13_59_768_0, i_13_59_816_0, i_13_59_942_0, i_13_59_976_0,
    i_13_59_979_0, i_13_59_1023_0, i_13_59_1081_0, i_13_59_1082_0,
    i_13_59_1087_0, i_13_59_1088_0, i_13_59_1096_0, i_13_59_1106_0,
    i_13_59_1147_0, i_13_59_1214_0, i_13_59_1270_0, i_13_59_1282_0,
    i_13_59_1309_0, i_13_59_1411_0, i_13_59_1514_0, i_13_59_1518_0,
    i_13_59_1561_0, i_13_59_1597_0, i_13_59_1680_0, i_13_59_1734_0,
    i_13_59_1741_0, i_13_59_1780_0, i_13_59_1849_0, i_13_59_1860_0,
    i_13_59_2002_0, i_13_59_2056_0, i_13_59_2191_0, i_13_59_2225_0,
    i_13_59_2383_0, i_13_59_2622_0, i_13_59_2769_0, i_13_59_2851_0,
    i_13_59_2878_0, i_13_59_2887_0, i_13_59_2907_0, i_13_59_2959_0,
    i_13_59_3028_0, i_13_59_3049_0, i_13_59_3113_0, i_13_59_3118_0,
    i_13_59_3156_0, i_13_59_3349_0, i_13_59_3352_0, i_13_59_3355_0,
    i_13_59_3382_0, i_13_59_3464_0, i_13_59_3534_0, i_13_59_3552_0,
    i_13_59_3571_0, i_13_59_3667_0, i_13_59_3730_0, i_13_59_3742_0,
    i_13_59_3984_0, i_13_59_3994_0, i_13_59_4063_0, i_13_59_4070_0,
    i_13_59_4108_0, i_13_59_4128_0, i_13_59_4155_0, i_13_59_4162_0,
    i_13_59_4165_0, i_13_59_4187_0, i_13_59_4299_0, i_13_59_4325_0,
    i_13_59_4335_0, i_13_59_4363_0, i_13_59_4369_0, i_13_59_4372_0,
    i_13_59_4418_0, i_13_59_4434_0, i_13_59_4532_0, i_13_59_4539_0;
  output o_13_59_0_0;
  assign o_13_59_0_0 = ~((i_13_59_1597_0 & (i_13_59_463_0 | (~i_13_59_1734_0 & ~i_13_59_2887_0 & ~i_13_59_3571_0))) | (~i_13_59_4165_0 & ((~i_13_59_192_0 & ~i_13_59_1214_0 & ~i_13_59_3464_0 & ~i_13_59_3571_0 & ~i_13_59_4187_0) | (i_13_59_1309_0 & ~i_13_59_4372_0))) | (i_13_59_192_0 & ~i_13_59_1081_0 & i_13_59_1270_0) | (~i_13_59_1087_0 & ~i_13_59_1860_0 & ~i_13_59_2851_0 & ~i_13_59_4162_0) | (~i_13_59_619_0 & i_13_59_760_0 & ~i_13_59_4363_0) | (i_13_59_2056_0 & ~i_13_59_4369_0));
endmodule



// Benchmark "kernel_13_60" written by ABC on Sun Jul 19 10:46:15 2020

module kernel_13_60 ( 
    i_13_60_48_0, i_13_60_70_0, i_13_60_76_0, i_13_60_177_0, i_13_60_193_0,
    i_13_60_197_0, i_13_60_204_0, i_13_60_411_0, i_13_60_445_0,
    i_13_60_482_0, i_13_60_570_0, i_13_60_610_0, i_13_60_628_0,
    i_13_60_660_0, i_13_60_663_0, i_13_60_672_0, i_13_60_682_0,
    i_13_60_853_0, i_13_60_939_0, i_13_60_980_0, i_13_60_989_0,
    i_13_60_1084_0, i_13_60_1105_0, i_13_60_1224_0, i_13_60_1227_0,
    i_13_60_1228_0, i_13_60_1231_0, i_13_60_1232_0, i_13_60_1246_0,
    i_13_60_1275_0, i_13_60_1317_0, i_13_60_1385_0, i_13_60_1483_0,
    i_13_60_1515_0, i_13_60_1525_0, i_13_60_1626_0, i_13_60_1645_0,
    i_13_60_1677_0, i_13_60_1727_0, i_13_60_1732_0, i_13_60_1764_0,
    i_13_60_1767_0, i_13_60_1768_0, i_13_60_1830_0, i_13_60_1894_0,
    i_13_60_1914_0, i_13_60_1929_0, i_13_60_1933_0, i_13_60_1936_0,
    i_13_60_2022_0, i_13_60_2137_0, i_13_60_2199_0, i_13_60_2298_0,
    i_13_60_2301_0, i_13_60_2366_0, i_13_60_2473_0, i_13_60_2518_0,
    i_13_60_2707_0, i_13_60_2851_0, i_13_60_3031_0, i_13_60_3117_0,
    i_13_60_3135_0, i_13_60_3176_0, i_13_60_3264_0, i_13_60_3274_0,
    i_13_60_3354_0, i_13_60_3426_0, i_13_60_3483_0, i_13_60_3486_0,
    i_13_60_3489_0, i_13_60_3549_0, i_13_60_3576_0, i_13_60_3577_0,
    i_13_60_3651_0, i_13_60_3729_0, i_13_60_3730_0, i_13_60_3756_0,
    i_13_60_3785_0, i_13_60_3822_0, i_13_60_3869_0, i_13_60_3900_0,
    i_13_60_3901_0, i_13_60_3932_0, i_13_60_3981_0, i_13_60_3994_0,
    i_13_60_4017_0, i_13_60_4164_0, i_13_60_4297_0, i_13_60_4321_0,
    i_13_60_4324_0, i_13_60_4336_0, i_13_60_4368_0, i_13_60_4371_0,
    i_13_60_4372_0, i_13_60_4379_0, i_13_60_4435_0, i_13_60_4506_0,
    i_13_60_4540_0, i_13_60_4566_0, i_13_60_4606_0,
    o_13_60_0_0  );
  input  i_13_60_48_0, i_13_60_70_0, i_13_60_76_0, i_13_60_177_0,
    i_13_60_193_0, i_13_60_197_0, i_13_60_204_0, i_13_60_411_0,
    i_13_60_445_0, i_13_60_482_0, i_13_60_570_0, i_13_60_610_0,
    i_13_60_628_0, i_13_60_660_0, i_13_60_663_0, i_13_60_672_0,
    i_13_60_682_0, i_13_60_853_0, i_13_60_939_0, i_13_60_980_0,
    i_13_60_989_0, i_13_60_1084_0, i_13_60_1105_0, i_13_60_1224_0,
    i_13_60_1227_0, i_13_60_1228_0, i_13_60_1231_0, i_13_60_1232_0,
    i_13_60_1246_0, i_13_60_1275_0, i_13_60_1317_0, i_13_60_1385_0,
    i_13_60_1483_0, i_13_60_1515_0, i_13_60_1525_0, i_13_60_1626_0,
    i_13_60_1645_0, i_13_60_1677_0, i_13_60_1727_0, i_13_60_1732_0,
    i_13_60_1764_0, i_13_60_1767_0, i_13_60_1768_0, i_13_60_1830_0,
    i_13_60_1894_0, i_13_60_1914_0, i_13_60_1929_0, i_13_60_1933_0,
    i_13_60_1936_0, i_13_60_2022_0, i_13_60_2137_0, i_13_60_2199_0,
    i_13_60_2298_0, i_13_60_2301_0, i_13_60_2366_0, i_13_60_2473_0,
    i_13_60_2518_0, i_13_60_2707_0, i_13_60_2851_0, i_13_60_3031_0,
    i_13_60_3117_0, i_13_60_3135_0, i_13_60_3176_0, i_13_60_3264_0,
    i_13_60_3274_0, i_13_60_3354_0, i_13_60_3426_0, i_13_60_3483_0,
    i_13_60_3486_0, i_13_60_3489_0, i_13_60_3549_0, i_13_60_3576_0,
    i_13_60_3577_0, i_13_60_3651_0, i_13_60_3729_0, i_13_60_3730_0,
    i_13_60_3756_0, i_13_60_3785_0, i_13_60_3822_0, i_13_60_3869_0,
    i_13_60_3900_0, i_13_60_3901_0, i_13_60_3932_0, i_13_60_3981_0,
    i_13_60_3994_0, i_13_60_4017_0, i_13_60_4164_0, i_13_60_4297_0,
    i_13_60_4321_0, i_13_60_4324_0, i_13_60_4336_0, i_13_60_4368_0,
    i_13_60_4371_0, i_13_60_4372_0, i_13_60_4379_0, i_13_60_4435_0,
    i_13_60_4506_0, i_13_60_4540_0, i_13_60_4566_0, i_13_60_4606_0;
  output o_13_60_0_0;
  assign o_13_60_0_0 = 0;
endmodule



// Benchmark "kernel_13_61" written by ABC on Sun Jul 19 10:46:16 2020

module kernel_13_61 ( 
    i_13_61_91_0, i_13_61_92_0, i_13_61_94_0, i_13_61_175_0, i_13_61_176_0,
    i_13_61_186_0, i_13_61_231_0, i_13_61_238_0, i_13_61_256_0,
    i_13_61_308_0, i_13_61_316_0, i_13_61_317_0, i_13_61_375_0,
    i_13_61_381_0, i_13_61_382_0, i_13_61_558_0, i_13_61_572_0,
    i_13_61_582_0, i_13_61_604_0, i_13_61_605_0, i_13_61_607_0,
    i_13_61_609_0, i_13_61_613_0, i_13_61_641_0, i_13_61_644_0,
    i_13_61_658_0, i_13_61_659_0, i_13_61_668_0, i_13_61_689_0,
    i_13_61_743_0, i_13_61_758_0, i_13_61_829_0, i_13_61_986_0,
    i_13_61_1060_0, i_13_61_1100_0, i_13_61_1119_0, i_13_61_1226_0,
    i_13_61_1228_0, i_13_61_1273_0, i_13_61_1391_0, i_13_61_1398_0,
    i_13_61_1399_0, i_13_61_1408_0, i_13_61_1442_0, i_13_61_1518_0,
    i_13_61_1568_0, i_13_61_1595_0, i_13_61_1638_0, i_13_61_1639_0,
    i_13_61_1765_0, i_13_61_1805_0, i_13_61_1813_0, i_13_61_1828_0,
    i_13_61_1831_0, i_13_61_1840_0, i_13_61_1918_0, i_13_61_2012_0,
    i_13_61_2128_0, i_13_61_2173_0, i_13_61_2281_0, i_13_61_2423_0,
    i_13_61_2431_0, i_13_61_2677_0, i_13_61_2767_0, i_13_61_3047_0,
    i_13_61_3107_0, i_13_61_3164_0, i_13_61_3235_0, i_13_61_3241_0,
    i_13_61_3291_0, i_13_61_3416_0, i_13_61_3423_0, i_13_61_3426_0,
    i_13_61_3451_0, i_13_61_3547_0, i_13_61_3631_0, i_13_61_3686_0,
    i_13_61_3709_0, i_13_61_3754_0, i_13_61_3767_0, i_13_61_3817_0,
    i_13_61_3872_0, i_13_61_3893_0, i_13_61_3919_0, i_13_61_3928_0,
    i_13_61_3992_0, i_13_61_4164_0, i_13_61_4186_0, i_13_61_4273_0,
    i_13_61_4376_0, i_13_61_4396_0, i_13_61_4430_0, i_13_61_4487_0,
    i_13_61_4511_0, i_13_61_4523_0, i_13_61_4538_0, i_13_61_4566_0,
    i_13_61_4567_0, i_13_61_4568_0, i_13_61_4591_0,
    o_13_61_0_0  );
  input  i_13_61_91_0, i_13_61_92_0, i_13_61_94_0, i_13_61_175_0,
    i_13_61_176_0, i_13_61_186_0, i_13_61_231_0, i_13_61_238_0,
    i_13_61_256_0, i_13_61_308_0, i_13_61_316_0, i_13_61_317_0,
    i_13_61_375_0, i_13_61_381_0, i_13_61_382_0, i_13_61_558_0,
    i_13_61_572_0, i_13_61_582_0, i_13_61_604_0, i_13_61_605_0,
    i_13_61_607_0, i_13_61_609_0, i_13_61_613_0, i_13_61_641_0,
    i_13_61_644_0, i_13_61_658_0, i_13_61_659_0, i_13_61_668_0,
    i_13_61_689_0, i_13_61_743_0, i_13_61_758_0, i_13_61_829_0,
    i_13_61_986_0, i_13_61_1060_0, i_13_61_1100_0, i_13_61_1119_0,
    i_13_61_1226_0, i_13_61_1228_0, i_13_61_1273_0, i_13_61_1391_0,
    i_13_61_1398_0, i_13_61_1399_0, i_13_61_1408_0, i_13_61_1442_0,
    i_13_61_1518_0, i_13_61_1568_0, i_13_61_1595_0, i_13_61_1638_0,
    i_13_61_1639_0, i_13_61_1765_0, i_13_61_1805_0, i_13_61_1813_0,
    i_13_61_1828_0, i_13_61_1831_0, i_13_61_1840_0, i_13_61_1918_0,
    i_13_61_2012_0, i_13_61_2128_0, i_13_61_2173_0, i_13_61_2281_0,
    i_13_61_2423_0, i_13_61_2431_0, i_13_61_2677_0, i_13_61_2767_0,
    i_13_61_3047_0, i_13_61_3107_0, i_13_61_3164_0, i_13_61_3235_0,
    i_13_61_3241_0, i_13_61_3291_0, i_13_61_3416_0, i_13_61_3423_0,
    i_13_61_3426_0, i_13_61_3451_0, i_13_61_3547_0, i_13_61_3631_0,
    i_13_61_3686_0, i_13_61_3709_0, i_13_61_3754_0, i_13_61_3767_0,
    i_13_61_3817_0, i_13_61_3872_0, i_13_61_3893_0, i_13_61_3919_0,
    i_13_61_3928_0, i_13_61_3992_0, i_13_61_4164_0, i_13_61_4186_0,
    i_13_61_4273_0, i_13_61_4376_0, i_13_61_4396_0, i_13_61_4430_0,
    i_13_61_4487_0, i_13_61_4511_0, i_13_61_4523_0, i_13_61_4538_0,
    i_13_61_4566_0, i_13_61_4567_0, i_13_61_4568_0, i_13_61_4591_0;
  output o_13_61_0_0;
  assign o_13_61_0_0 = ~((~i_13_61_1408_0 & ((~i_13_61_176_0 & ~i_13_61_1765_0 & i_13_61_2767_0 & i_13_61_3235_0 & ~i_13_61_3872_0 & ~i_13_61_3992_0) | (~i_13_61_91_0 & ~i_13_61_1638_0 & ~i_13_61_1828_0 & ~i_13_61_2677_0 & ~i_13_61_3423_0 & ~i_13_61_3893_0 & ~i_13_61_4511_0))) | (~i_13_61_176_0 & ((~i_13_61_2677_0 & i_13_61_3235_0 & ~i_13_61_4430_0) | (~i_13_61_1595_0 & i_13_61_3919_0 & ~i_13_61_4186_0 & i_13_61_4396_0 & ~i_13_61_4567_0))) | (i_13_61_1813_0 & ((~i_13_61_1226_0 & ~i_13_61_1831_0 & ~i_13_61_3919_0) | (i_13_61_1805_0 & i_13_61_3686_0 & ~i_13_61_4568_0))) | (i_13_61_3423_0 & ((~i_13_61_2677_0 & i_13_61_3451_0) | (~i_13_61_1828_0 & ~i_13_61_2431_0 & ~i_13_61_3426_0 & ~i_13_61_3928_0 & ~i_13_61_4273_0))) | (i_13_61_231_0 & ~i_13_61_1831_0 & ~i_13_61_3426_0) | (~i_13_61_689_0 & ~i_13_61_1119_0 & ~i_13_61_2173_0 & ~i_13_61_3754_0 & ~i_13_61_3893_0) | (~i_13_61_175_0 & i_13_61_2767_0 & i_13_61_4396_0) | (~i_13_61_94_0 & i_13_61_238_0 & ~i_13_61_1805_0 & ~i_13_61_4568_0));
endmodule



// Benchmark "kernel_13_62" written by ABC on Sun Jul 19 10:46:17 2020

module kernel_13_62 ( 
    i_13_62_41_0, i_13_62_113_0, i_13_62_115_0, i_13_62_137_0,
    i_13_62_166_0, i_13_62_167_0, i_13_62_189_0, i_13_62_227_0,
    i_13_62_266_0, i_13_62_279_0, i_13_62_367_0, i_13_62_390_0,
    i_13_62_534_0, i_13_62_572_0, i_13_62_606_0, i_13_62_608_0,
    i_13_62_660_0, i_13_62_679_0, i_13_62_811_0, i_13_62_814_0,
    i_13_62_856_0, i_13_62_947_0, i_13_62_1084_0, i_13_62_1085_0,
    i_13_62_1094_0, i_13_62_1211_0, i_13_62_1217_0, i_13_62_1219_0,
    i_13_62_1352_0, i_13_62_1427_0, i_13_62_1462_0, i_13_62_1621_0,
    i_13_62_1622_0, i_13_62_1634_0, i_13_62_1640_0, i_13_62_1778_0,
    i_13_62_1788_0, i_13_62_1837_0, i_13_62_1838_0, i_13_62_1840_0,
    i_13_62_1841_0, i_13_62_1849_0, i_13_62_1939_0, i_13_62_1998_0,
    i_13_62_2021_0, i_13_62_2128_0, i_13_62_2135_0, i_13_62_2170_0,
    i_13_62_2172_0, i_13_62_2173_0, i_13_62_2209_0, i_13_62_2264_0,
    i_13_62_2404_0, i_13_62_2405_0, i_13_62_2407_0, i_13_62_2408_0,
    i_13_62_2421_0, i_13_62_2426_0, i_13_62_2432_0, i_13_62_2435_0,
    i_13_62_2448_0, i_13_62_2458_0, i_13_62_2495_0, i_13_62_2498_0,
    i_13_62_2564_0, i_13_62_2713_0, i_13_62_2714_0, i_13_62_2791_0,
    i_13_62_2846_0, i_13_62_2880_0, i_13_62_2907_0, i_13_62_2920_0,
    i_13_62_3044_0, i_13_62_3128_0, i_13_62_3141_0, i_13_62_3145_0,
    i_13_62_3146_0, i_13_62_3149_0, i_13_62_3407_0, i_13_62_3451_0,
    i_13_62_3452_0, i_13_62_3505_0, i_13_62_3509_0, i_13_62_3515_0,
    i_13_62_3529_0, i_13_62_3605_0, i_13_62_3613_0, i_13_62_3699_0,
    i_13_62_3737_0, i_13_62_3739_0, i_13_62_3763_0, i_13_62_3891_0,
    i_13_62_3892_0, i_13_62_4007_0, i_13_62_4160_0, i_13_62_4315_0,
    i_13_62_4325_0, i_13_62_4542_0, i_13_62_4555_0, i_13_62_4559_0,
    o_13_62_0_0  );
  input  i_13_62_41_0, i_13_62_113_0, i_13_62_115_0, i_13_62_137_0,
    i_13_62_166_0, i_13_62_167_0, i_13_62_189_0, i_13_62_227_0,
    i_13_62_266_0, i_13_62_279_0, i_13_62_367_0, i_13_62_390_0,
    i_13_62_534_0, i_13_62_572_0, i_13_62_606_0, i_13_62_608_0,
    i_13_62_660_0, i_13_62_679_0, i_13_62_811_0, i_13_62_814_0,
    i_13_62_856_0, i_13_62_947_0, i_13_62_1084_0, i_13_62_1085_0,
    i_13_62_1094_0, i_13_62_1211_0, i_13_62_1217_0, i_13_62_1219_0,
    i_13_62_1352_0, i_13_62_1427_0, i_13_62_1462_0, i_13_62_1621_0,
    i_13_62_1622_0, i_13_62_1634_0, i_13_62_1640_0, i_13_62_1778_0,
    i_13_62_1788_0, i_13_62_1837_0, i_13_62_1838_0, i_13_62_1840_0,
    i_13_62_1841_0, i_13_62_1849_0, i_13_62_1939_0, i_13_62_1998_0,
    i_13_62_2021_0, i_13_62_2128_0, i_13_62_2135_0, i_13_62_2170_0,
    i_13_62_2172_0, i_13_62_2173_0, i_13_62_2209_0, i_13_62_2264_0,
    i_13_62_2404_0, i_13_62_2405_0, i_13_62_2407_0, i_13_62_2408_0,
    i_13_62_2421_0, i_13_62_2426_0, i_13_62_2432_0, i_13_62_2435_0,
    i_13_62_2448_0, i_13_62_2458_0, i_13_62_2495_0, i_13_62_2498_0,
    i_13_62_2564_0, i_13_62_2713_0, i_13_62_2714_0, i_13_62_2791_0,
    i_13_62_2846_0, i_13_62_2880_0, i_13_62_2907_0, i_13_62_2920_0,
    i_13_62_3044_0, i_13_62_3128_0, i_13_62_3141_0, i_13_62_3145_0,
    i_13_62_3146_0, i_13_62_3149_0, i_13_62_3407_0, i_13_62_3451_0,
    i_13_62_3452_0, i_13_62_3505_0, i_13_62_3509_0, i_13_62_3515_0,
    i_13_62_3529_0, i_13_62_3605_0, i_13_62_3613_0, i_13_62_3699_0,
    i_13_62_3737_0, i_13_62_3739_0, i_13_62_3763_0, i_13_62_3891_0,
    i_13_62_3892_0, i_13_62_4007_0, i_13_62_4160_0, i_13_62_4315_0,
    i_13_62_4325_0, i_13_62_4542_0, i_13_62_4555_0, i_13_62_4559_0;
  output o_13_62_0_0;
  assign o_13_62_0_0 = ~((~i_13_62_1084_0 & ((~i_13_62_811_0 & ~i_13_62_1085_0 & ~i_13_62_1998_0 & ~i_13_62_2170_0 & ~i_13_62_2713_0 & ~i_13_62_3452_0) | (~i_13_62_2432_0 & ~i_13_62_2458_0 & ~i_13_62_3141_0 & ~i_13_62_3149_0 & ~i_13_62_4007_0))) | (~i_13_62_2880_0 & ((~i_13_62_1219_0 & ~i_13_62_1427_0 & ~i_13_62_1998_0 & ~i_13_62_2421_0 & ~i_13_62_4160_0) | (i_13_62_2404_0 & ~i_13_62_4325_0))) | (~i_13_62_4559_0 & (i_13_62_2408_0 | (i_13_62_3892_0 & ~i_13_62_4555_0))) | (~i_13_62_113_0 & ~i_13_62_2021_0 & ~i_13_62_2448_0 & ~i_13_62_2458_0) | (~i_13_62_115_0 & ~i_13_62_1838_0 & ~i_13_62_2172_0 & ~i_13_62_3451_0 & ~i_13_62_4007_0) | (i_13_62_2405_0 & ~i_13_62_4325_0));
endmodule



// Benchmark "kernel_13_63" written by ABC on Sun Jul 19 10:46:17 2020

module kernel_13_63 ( 
    i_13_63_49_0, i_13_63_67_0, i_13_63_71_0, i_13_63_77_0, i_13_63_183_0,
    i_13_63_314_0, i_13_63_319_0, i_13_63_412_0, i_13_63_439_0,
    i_13_63_445_0, i_13_63_456_0, i_13_63_459_0, i_13_63_611_0,
    i_13_63_616_0, i_13_63_619_0, i_13_63_661_0, i_13_63_664_0,
    i_13_63_683_0, i_13_63_760_0, i_13_63_761_0, i_13_63_763_0,
    i_13_63_833_0, i_13_63_846_0, i_13_63_912_0, i_13_63_934_0,
    i_13_63_935_0, i_13_63_1096_0, i_13_63_1097_0, i_13_63_1102_0,
    i_13_63_1105_0, i_13_63_1132_0, i_13_63_1133_0, i_13_63_1155_0,
    i_13_63_1247_0, i_13_63_1258_0, i_13_63_1409_0, i_13_63_1483_0,
    i_13_63_1511_0, i_13_63_1525_0, i_13_63_1597_0, i_13_63_1645_0,
    i_13_63_1679_0, i_13_63_1733_0, i_13_63_1736_0, i_13_63_1754_0,
    i_13_63_1768_0, i_13_63_1771_0, i_13_63_1798_0, i_13_63_1799_0,
    i_13_63_1808_0, i_13_63_1885_0, i_13_63_1915_0, i_13_63_2023_0,
    i_13_63_2024_0, i_13_63_2029_0, i_13_63_2056_0, i_13_63_2149_0,
    i_13_63_2473_0, i_13_63_2474_0, i_13_63_2677_0, i_13_63_2708_0,
    i_13_63_2744_0, i_13_63_2857_0, i_13_63_2898_0, i_13_63_2902_0,
    i_13_63_2941_0, i_13_63_3031_0, i_13_63_3032_0, i_13_63_3077_0,
    i_13_63_3121_0, i_13_63_3231_0, i_13_63_3246_0, i_13_63_3265_0,
    i_13_63_3266_0, i_13_63_3346_0, i_13_63_3356_0, i_13_63_3397_0,
    i_13_63_3436_0, i_13_63_3461_0, i_13_63_3550_0, i_13_63_3551_0,
    i_13_63_3702_0, i_13_63_3739_0, i_13_63_3760_0, i_13_63_3784_0,
    i_13_63_3823_0, i_13_63_3847_0, i_13_63_3902_0, i_13_63_3911_0,
    i_13_63_3928_0, i_13_63_4085_0, i_13_63_4165_0, i_13_63_4245_0,
    i_13_63_4274_0, i_13_63_4325_0, i_13_63_4374_0, i_13_63_4397_0,
    i_13_63_4558_0, i_13_63_4606_0, i_13_63_4607_0,
    o_13_63_0_0  );
  input  i_13_63_49_0, i_13_63_67_0, i_13_63_71_0, i_13_63_77_0,
    i_13_63_183_0, i_13_63_314_0, i_13_63_319_0, i_13_63_412_0,
    i_13_63_439_0, i_13_63_445_0, i_13_63_456_0, i_13_63_459_0,
    i_13_63_611_0, i_13_63_616_0, i_13_63_619_0, i_13_63_661_0,
    i_13_63_664_0, i_13_63_683_0, i_13_63_760_0, i_13_63_761_0,
    i_13_63_763_0, i_13_63_833_0, i_13_63_846_0, i_13_63_912_0,
    i_13_63_934_0, i_13_63_935_0, i_13_63_1096_0, i_13_63_1097_0,
    i_13_63_1102_0, i_13_63_1105_0, i_13_63_1132_0, i_13_63_1133_0,
    i_13_63_1155_0, i_13_63_1247_0, i_13_63_1258_0, i_13_63_1409_0,
    i_13_63_1483_0, i_13_63_1511_0, i_13_63_1525_0, i_13_63_1597_0,
    i_13_63_1645_0, i_13_63_1679_0, i_13_63_1733_0, i_13_63_1736_0,
    i_13_63_1754_0, i_13_63_1768_0, i_13_63_1771_0, i_13_63_1798_0,
    i_13_63_1799_0, i_13_63_1808_0, i_13_63_1885_0, i_13_63_1915_0,
    i_13_63_2023_0, i_13_63_2024_0, i_13_63_2029_0, i_13_63_2056_0,
    i_13_63_2149_0, i_13_63_2473_0, i_13_63_2474_0, i_13_63_2677_0,
    i_13_63_2708_0, i_13_63_2744_0, i_13_63_2857_0, i_13_63_2898_0,
    i_13_63_2902_0, i_13_63_2941_0, i_13_63_3031_0, i_13_63_3032_0,
    i_13_63_3077_0, i_13_63_3121_0, i_13_63_3231_0, i_13_63_3246_0,
    i_13_63_3265_0, i_13_63_3266_0, i_13_63_3346_0, i_13_63_3356_0,
    i_13_63_3397_0, i_13_63_3436_0, i_13_63_3461_0, i_13_63_3550_0,
    i_13_63_3551_0, i_13_63_3702_0, i_13_63_3739_0, i_13_63_3760_0,
    i_13_63_3784_0, i_13_63_3823_0, i_13_63_3847_0, i_13_63_3902_0,
    i_13_63_3911_0, i_13_63_3928_0, i_13_63_4085_0, i_13_63_4165_0,
    i_13_63_4245_0, i_13_63_4274_0, i_13_63_4325_0, i_13_63_4374_0,
    i_13_63_4397_0, i_13_63_4558_0, i_13_63_4606_0, i_13_63_4607_0;
  output o_13_63_0_0;
  assign o_13_63_0_0 = ~((~i_13_63_934_0 & ((i_13_63_1597_0 & ~i_13_63_2023_0) | (~i_13_63_3784_0 & ~i_13_63_3911_0 & ~i_13_63_4085_0))) | (i_13_63_4374_0 & (i_13_63_1885_0 | ~i_13_63_2029_0)) | (~i_13_63_3265_0 & (i_13_63_616_0 | (~i_13_63_2149_0 & i_13_63_3397_0) | (~i_13_63_459_0 & ~i_13_63_1679_0 & ~i_13_63_4274_0))) | (~i_13_63_4274_0 & ((i_13_63_445_0 & i_13_63_2677_0) | (~i_13_63_1525_0 & ~i_13_63_3550_0 & i_13_63_3928_0 & ~i_13_63_4085_0))) | (i_13_63_319_0 & ~i_13_63_3346_0) | (i_13_63_761_0 & ~i_13_63_4165_0) | (~i_13_63_77_0 & ~i_13_63_683_0 & ~i_13_63_2941_0 & ~i_13_63_3847_0 & ~i_13_63_4374_0));
endmodule



// Benchmark "kernel_13_64" written by ABC on Sun Jul 19 10:46:18 2020

module kernel_13_64 ( 
    i_13_64_46_0, i_13_64_48_0, i_13_64_166_0, i_13_64_506_0,
    i_13_64_551_0, i_13_64_837_0, i_13_64_840_0, i_13_64_870_0,
    i_13_64_936_0, i_13_64_1058_0, i_13_64_1066_0, i_13_64_1119_0,
    i_13_64_1188_0, i_13_64_1189_0, i_13_64_1219_0, i_13_64_1245_0,
    i_13_64_1262_0, i_13_64_1323_0, i_13_64_1324_0, i_13_64_1326_0,
    i_13_64_1327_0, i_13_64_1405_0, i_13_64_1458_0, i_13_64_1512_0,
    i_13_64_1527_0, i_13_64_1628_0, i_13_64_1664_0, i_13_64_1777_0,
    i_13_64_1803_0, i_13_64_1805_0, i_13_64_1828_0, i_13_64_1831_0,
    i_13_64_1848_0, i_13_64_1849_0, i_13_64_1850_0, i_13_64_1855_0,
    i_13_64_1884_0, i_13_64_1885_0, i_13_64_1892_0, i_13_64_1896_0,
    i_13_64_2009_0, i_13_64_2043_0, i_13_64_2107_0, i_13_64_2145_0,
    i_13_64_2262_0, i_13_64_2299_0, i_13_64_2302_0, i_13_64_2351_0,
    i_13_64_2403_0, i_13_64_2469_0, i_13_64_2470_0, i_13_64_2472_0,
    i_13_64_2694_0, i_13_64_2697_0, i_13_64_2735_0, i_13_64_2740_0,
    i_13_64_2745_0, i_13_64_2980_0, i_13_64_2981_0, i_13_64_2982_0,
    i_13_64_2985_0, i_13_64_3028_0, i_13_64_3029_0, i_13_64_3055_0,
    i_13_64_3068_0, i_13_64_3105_0, i_13_64_3107_0, i_13_64_3108_0,
    i_13_64_3126_0, i_13_64_3211_0, i_13_64_3343_0, i_13_64_3503_0,
    i_13_64_3512_0, i_13_64_3523_0, i_13_64_3547_0, i_13_64_3548_0,
    i_13_64_3549_0, i_13_64_3604_0, i_13_64_3739_0, i_13_64_3763_0,
    i_13_64_3785_0, i_13_64_3816_0, i_13_64_3817_0, i_13_64_3820_0,
    i_13_64_3908_0, i_13_64_3930_0, i_13_64_4045_0, i_13_64_4059_0,
    i_13_64_4062_0, i_13_64_4063_0, i_13_64_4126_0, i_13_64_4162_0,
    i_13_64_4218_0, i_13_64_4315_0, i_13_64_4322_0, i_13_64_4376_0,
    i_13_64_4441_0, i_13_64_4497_0, i_13_64_4563_0, i_13_64_4567_0,
    o_13_64_0_0  );
  input  i_13_64_46_0, i_13_64_48_0, i_13_64_166_0, i_13_64_506_0,
    i_13_64_551_0, i_13_64_837_0, i_13_64_840_0, i_13_64_870_0,
    i_13_64_936_0, i_13_64_1058_0, i_13_64_1066_0, i_13_64_1119_0,
    i_13_64_1188_0, i_13_64_1189_0, i_13_64_1219_0, i_13_64_1245_0,
    i_13_64_1262_0, i_13_64_1323_0, i_13_64_1324_0, i_13_64_1326_0,
    i_13_64_1327_0, i_13_64_1405_0, i_13_64_1458_0, i_13_64_1512_0,
    i_13_64_1527_0, i_13_64_1628_0, i_13_64_1664_0, i_13_64_1777_0,
    i_13_64_1803_0, i_13_64_1805_0, i_13_64_1828_0, i_13_64_1831_0,
    i_13_64_1848_0, i_13_64_1849_0, i_13_64_1850_0, i_13_64_1855_0,
    i_13_64_1884_0, i_13_64_1885_0, i_13_64_1892_0, i_13_64_1896_0,
    i_13_64_2009_0, i_13_64_2043_0, i_13_64_2107_0, i_13_64_2145_0,
    i_13_64_2262_0, i_13_64_2299_0, i_13_64_2302_0, i_13_64_2351_0,
    i_13_64_2403_0, i_13_64_2469_0, i_13_64_2470_0, i_13_64_2472_0,
    i_13_64_2694_0, i_13_64_2697_0, i_13_64_2735_0, i_13_64_2740_0,
    i_13_64_2745_0, i_13_64_2980_0, i_13_64_2981_0, i_13_64_2982_0,
    i_13_64_2985_0, i_13_64_3028_0, i_13_64_3029_0, i_13_64_3055_0,
    i_13_64_3068_0, i_13_64_3105_0, i_13_64_3107_0, i_13_64_3108_0,
    i_13_64_3126_0, i_13_64_3211_0, i_13_64_3343_0, i_13_64_3503_0,
    i_13_64_3512_0, i_13_64_3523_0, i_13_64_3547_0, i_13_64_3548_0,
    i_13_64_3549_0, i_13_64_3604_0, i_13_64_3739_0, i_13_64_3763_0,
    i_13_64_3785_0, i_13_64_3816_0, i_13_64_3817_0, i_13_64_3820_0,
    i_13_64_3908_0, i_13_64_3930_0, i_13_64_4045_0, i_13_64_4059_0,
    i_13_64_4062_0, i_13_64_4063_0, i_13_64_4126_0, i_13_64_4162_0,
    i_13_64_4218_0, i_13_64_4315_0, i_13_64_4322_0, i_13_64_4376_0,
    i_13_64_4441_0, i_13_64_4497_0, i_13_64_4563_0, i_13_64_4567_0;
  output o_13_64_0_0;
  assign o_13_64_0_0 = ~((~i_13_64_48_0 & ((~i_13_64_936_0 & ~i_13_64_1324_0 & ~i_13_64_1848_0 & ~i_13_64_3930_0) | (~i_13_64_46_0 & ~i_13_64_2145_0 & ~i_13_64_4315_0 & ~i_13_64_4563_0))) | (~i_13_64_3820_0 & ((~i_13_64_1323_0 & ~i_13_64_1828_0 & ~i_13_64_2694_0) | (~i_13_64_2982_0 & ~i_13_64_3604_0 & ~i_13_64_3817_0 & ~i_13_64_4563_0))) | (~i_13_64_1855_0 & i_13_64_1885_0 & ~i_13_64_3343_0 & ~i_13_64_4563_0) | (i_13_64_1219_0 & ~i_13_64_2740_0 & i_13_64_3604_0) | (~i_13_64_1066_0 & i_13_64_3785_0) | (~i_13_64_1848_0 & ~i_13_64_2145_0 & ~i_13_64_2299_0 & ~i_13_64_4376_0) | (~i_13_64_1831_0 & ~i_13_64_4567_0));
endmodule



// Benchmark "kernel_13_65" written by ABC on Sun Jul 19 10:46:19 2020

module kernel_13_65 ( 
    i_13_65_137_0, i_13_65_164_0, i_13_65_166_0, i_13_65_167_0,
    i_13_65_169_0, i_13_65_172_0, i_13_65_229_0, i_13_65_263_0,
    i_13_65_266_0, i_13_65_281_0, i_13_65_380_0, i_13_65_460_0,
    i_13_65_530_0, i_13_65_607_0, i_13_65_640_0, i_13_65_676_0,
    i_13_65_688_0, i_13_65_794_0, i_13_65_811_0, i_13_65_814_0,
    i_13_65_815_0, i_13_65_821_0, i_13_65_823_0, i_13_65_824_0,
    i_13_65_913_0, i_13_65_961_0, i_13_65_982_0, i_13_65_1063_0,
    i_13_65_1064_0, i_13_65_1249_0, i_13_65_1324_0, i_13_65_1332_0,
    i_13_65_1495_0, i_13_65_1499_0, i_13_65_1502_0, i_13_65_1655_0,
    i_13_65_1846_0, i_13_65_1847_0, i_13_65_1849_0, i_13_65_1850_0,
    i_13_65_1852_0, i_13_65_1909_0, i_13_65_1958_0, i_13_65_1962_0,
    i_13_65_2107_0, i_13_65_2108_0, i_13_65_2116_0, i_13_65_2117_0,
    i_13_65_2134_0, i_13_65_2146_0, i_13_65_2227_0, i_13_65_2234_0,
    i_13_65_2247_0, i_13_65_2260_0, i_13_65_2261_0, i_13_65_2404_0,
    i_13_65_2405_0, i_13_65_2407_0, i_13_65_2408_0, i_13_65_2419_0,
    i_13_65_2449_0, i_13_65_2674_0, i_13_65_2678_0, i_13_65_2753_0,
    i_13_65_2848_0, i_13_65_2935_0, i_13_65_2936_0, i_13_65_3011_0,
    i_13_65_3148_0, i_13_65_3268_0, i_13_65_3374_0, i_13_65_3394_0,
    i_13_65_3438_0, i_13_65_3503_0, i_13_65_3505_0, i_13_65_3523_0,
    i_13_65_3595_0, i_13_65_3641_0, i_13_65_3739_0, i_13_65_3762_0,
    i_13_65_3817_0, i_13_65_3818_0, i_13_65_3862_0, i_13_65_3977_0,
    i_13_65_4015_0, i_13_65_4042_0, i_13_65_4060_0, i_13_65_4061_0,
    i_13_65_4063_0, i_13_65_4064_0, i_13_65_4123_0, i_13_65_4268_0,
    i_13_65_4303_0, i_13_65_4304_0, i_13_65_4315_0, i_13_65_4316_0,
    i_13_65_4319_0, i_13_65_4335_0, i_13_65_4405_0, i_13_65_4466_0,
    o_13_65_0_0  );
  input  i_13_65_137_0, i_13_65_164_0, i_13_65_166_0, i_13_65_167_0,
    i_13_65_169_0, i_13_65_172_0, i_13_65_229_0, i_13_65_263_0,
    i_13_65_266_0, i_13_65_281_0, i_13_65_380_0, i_13_65_460_0,
    i_13_65_530_0, i_13_65_607_0, i_13_65_640_0, i_13_65_676_0,
    i_13_65_688_0, i_13_65_794_0, i_13_65_811_0, i_13_65_814_0,
    i_13_65_815_0, i_13_65_821_0, i_13_65_823_0, i_13_65_824_0,
    i_13_65_913_0, i_13_65_961_0, i_13_65_982_0, i_13_65_1063_0,
    i_13_65_1064_0, i_13_65_1249_0, i_13_65_1324_0, i_13_65_1332_0,
    i_13_65_1495_0, i_13_65_1499_0, i_13_65_1502_0, i_13_65_1655_0,
    i_13_65_1846_0, i_13_65_1847_0, i_13_65_1849_0, i_13_65_1850_0,
    i_13_65_1852_0, i_13_65_1909_0, i_13_65_1958_0, i_13_65_1962_0,
    i_13_65_2107_0, i_13_65_2108_0, i_13_65_2116_0, i_13_65_2117_0,
    i_13_65_2134_0, i_13_65_2146_0, i_13_65_2227_0, i_13_65_2234_0,
    i_13_65_2247_0, i_13_65_2260_0, i_13_65_2261_0, i_13_65_2404_0,
    i_13_65_2405_0, i_13_65_2407_0, i_13_65_2408_0, i_13_65_2419_0,
    i_13_65_2449_0, i_13_65_2674_0, i_13_65_2678_0, i_13_65_2753_0,
    i_13_65_2848_0, i_13_65_2935_0, i_13_65_2936_0, i_13_65_3011_0,
    i_13_65_3148_0, i_13_65_3268_0, i_13_65_3374_0, i_13_65_3394_0,
    i_13_65_3438_0, i_13_65_3503_0, i_13_65_3505_0, i_13_65_3523_0,
    i_13_65_3595_0, i_13_65_3641_0, i_13_65_3739_0, i_13_65_3762_0,
    i_13_65_3817_0, i_13_65_3818_0, i_13_65_3862_0, i_13_65_3977_0,
    i_13_65_4015_0, i_13_65_4042_0, i_13_65_4060_0, i_13_65_4061_0,
    i_13_65_4063_0, i_13_65_4064_0, i_13_65_4123_0, i_13_65_4268_0,
    i_13_65_4303_0, i_13_65_4304_0, i_13_65_4315_0, i_13_65_4316_0,
    i_13_65_4319_0, i_13_65_4335_0, i_13_65_4405_0, i_13_65_4466_0;
  output o_13_65_0_0;
  assign o_13_65_0_0 = ~((~i_13_65_1063_0 & ~i_13_65_4316_0) | (i_13_65_3438_0 & ~i_13_65_4315_0) | (~i_13_65_982_0 & ~i_13_65_4303_0) | (i_13_65_3762_0 & i_13_65_4303_0) | (~i_13_65_1846_0 & ~i_13_65_2405_0 & ~i_13_65_3438_0));
endmodule



// Benchmark "kernel_13_66" written by ABC on Sun Jul 19 10:46:20 2020

module kernel_13_66 ( 
    i_13_66_40_0, i_13_66_59_0, i_13_66_121_0, i_13_66_139_0,
    i_13_66_192_0, i_13_66_229_0, i_13_66_236_0, i_13_66_383_0,
    i_13_66_398_0, i_13_66_576_0, i_13_66_589_0, i_13_66_658_0,
    i_13_66_660_0, i_13_66_661_0, i_13_66_829_0, i_13_66_832_0,
    i_13_66_886_0, i_13_66_928_0, i_13_66_939_0, i_13_66_1000_0,
    i_13_66_1063_0, i_13_66_1098_0, i_13_66_1117_0, i_13_66_1118_0,
    i_13_66_1147_0, i_13_66_1225_0, i_13_66_1226_0, i_13_66_1227_0,
    i_13_66_1228_0, i_13_66_1244_0, i_13_66_1407_0, i_13_66_1408_0,
    i_13_66_1410_0, i_13_66_1479_0, i_13_66_1481_0, i_13_66_1513_0,
    i_13_66_1539_0, i_13_66_1552_0, i_13_66_1596_0, i_13_66_1652_0,
    i_13_66_1657_0, i_13_66_1675_0, i_13_66_1678_0, i_13_66_1733_0,
    i_13_66_1764_0, i_13_66_1765_0, i_13_66_1801_0, i_13_66_1802_0,
    i_13_66_1892_0, i_13_66_1927_0, i_13_66_1999_0, i_13_66_2002_0,
    i_13_66_2016_0, i_13_66_2296_0, i_13_66_2359_0, i_13_66_2443_0,
    i_13_66_2467_0, i_13_66_2569_0, i_13_66_2702_0, i_13_66_2705_0,
    i_13_66_2835_0, i_13_66_2857_0, i_13_66_2859_0, i_13_66_2874_0,
    i_13_66_2907_0, i_13_66_2980_0, i_13_66_2982_0, i_13_66_3017_0,
    i_13_66_3109_0, i_13_66_3133_0, i_13_66_3145_0, i_13_66_3371_0,
    i_13_66_3421_0, i_13_66_3475_0, i_13_66_3476_0, i_13_66_3486_0,
    i_13_66_3546_0, i_13_66_3547_0, i_13_66_3667_0, i_13_66_3730_0,
    i_13_66_3754_0, i_13_66_3757_0, i_13_66_3862_0, i_13_66_3979_0,
    i_13_66_3980_0, i_13_66_4086_0, i_13_66_4162_0, i_13_66_4186_0,
    i_13_66_4195_0, i_13_66_4295_0, i_13_66_4369_0, i_13_66_4393_0,
    i_13_66_4396_0, i_13_66_4428_0, i_13_66_4510_0, i_13_66_4511_0,
    i_13_66_4538_0, i_13_66_4599_0, i_13_66_4600_0, i_13_66_4603_0,
    o_13_66_0_0  );
  input  i_13_66_40_0, i_13_66_59_0, i_13_66_121_0, i_13_66_139_0,
    i_13_66_192_0, i_13_66_229_0, i_13_66_236_0, i_13_66_383_0,
    i_13_66_398_0, i_13_66_576_0, i_13_66_589_0, i_13_66_658_0,
    i_13_66_660_0, i_13_66_661_0, i_13_66_829_0, i_13_66_832_0,
    i_13_66_886_0, i_13_66_928_0, i_13_66_939_0, i_13_66_1000_0,
    i_13_66_1063_0, i_13_66_1098_0, i_13_66_1117_0, i_13_66_1118_0,
    i_13_66_1147_0, i_13_66_1225_0, i_13_66_1226_0, i_13_66_1227_0,
    i_13_66_1228_0, i_13_66_1244_0, i_13_66_1407_0, i_13_66_1408_0,
    i_13_66_1410_0, i_13_66_1479_0, i_13_66_1481_0, i_13_66_1513_0,
    i_13_66_1539_0, i_13_66_1552_0, i_13_66_1596_0, i_13_66_1652_0,
    i_13_66_1657_0, i_13_66_1675_0, i_13_66_1678_0, i_13_66_1733_0,
    i_13_66_1764_0, i_13_66_1765_0, i_13_66_1801_0, i_13_66_1802_0,
    i_13_66_1892_0, i_13_66_1927_0, i_13_66_1999_0, i_13_66_2002_0,
    i_13_66_2016_0, i_13_66_2296_0, i_13_66_2359_0, i_13_66_2443_0,
    i_13_66_2467_0, i_13_66_2569_0, i_13_66_2702_0, i_13_66_2705_0,
    i_13_66_2835_0, i_13_66_2857_0, i_13_66_2859_0, i_13_66_2874_0,
    i_13_66_2907_0, i_13_66_2980_0, i_13_66_2982_0, i_13_66_3017_0,
    i_13_66_3109_0, i_13_66_3133_0, i_13_66_3145_0, i_13_66_3371_0,
    i_13_66_3421_0, i_13_66_3475_0, i_13_66_3476_0, i_13_66_3486_0,
    i_13_66_3546_0, i_13_66_3547_0, i_13_66_3667_0, i_13_66_3730_0,
    i_13_66_3754_0, i_13_66_3757_0, i_13_66_3862_0, i_13_66_3979_0,
    i_13_66_3980_0, i_13_66_4086_0, i_13_66_4162_0, i_13_66_4186_0,
    i_13_66_4195_0, i_13_66_4295_0, i_13_66_4369_0, i_13_66_4393_0,
    i_13_66_4396_0, i_13_66_4428_0, i_13_66_4510_0, i_13_66_4511_0,
    i_13_66_4538_0, i_13_66_4599_0, i_13_66_4600_0, i_13_66_4603_0;
  output o_13_66_0_0;
  assign o_13_66_0_0 = ~((~i_13_66_1764_0 & ((~i_13_66_1801_0 & ~i_13_66_4086_0) | (~i_13_66_1765_0 & ~i_13_66_4162_0))) | (~i_13_66_3754_0 & (~i_13_66_3546_0 | ~i_13_66_3979_0)) | (~i_13_66_3980_0 & (~i_13_66_886_0 | (i_13_66_2002_0 & ~i_13_66_4428_0))) | ~i_13_66_1147_0 | (i_13_66_928_0 & ~i_13_66_3979_0));
endmodule



// Benchmark "kernel_13_67" written by ABC on Sun Jul 19 10:46:21 2020

module kernel_13_67 ( 
    i_13_67_64_0, i_13_67_90_0, i_13_67_91_0, i_13_67_139_0, i_13_67_174_0,
    i_13_67_175_0, i_13_67_204_0, i_13_67_228_0, i_13_67_229_0,
    i_13_67_282_0, i_13_67_283_0, i_13_67_284_0, i_13_67_336_0,
    i_13_67_337_0, i_13_67_341_0, i_13_67_393_0, i_13_67_414_0,
    i_13_67_417_0, i_13_67_450_0, i_13_67_522_0, i_13_67_535_0,
    i_13_67_567_0, i_13_67_657_0, i_13_67_661_0, i_13_67_733_0,
    i_13_67_796_0, i_13_67_823_0, i_13_67_824_0, i_13_67_846_0,
    i_13_67_847_0, i_13_67_849_0, i_13_67_850_0, i_13_67_981_0,
    i_13_67_985_0, i_13_67_1219_0, i_13_67_1224_0, i_13_67_1252_0,
    i_13_67_1263_0, i_13_67_1309_0, i_13_67_1312_0, i_13_67_1317_0,
    i_13_67_1462_0, i_13_67_1485_0, i_13_67_1549_0, i_13_67_1551_0,
    i_13_67_1552_0, i_13_67_1624_0, i_13_67_1644_0, i_13_67_1710_0,
    i_13_67_1803_0, i_13_67_1857_0, i_13_67_1858_0, i_13_67_1860_0,
    i_13_67_2197_0, i_13_67_2431_0, i_13_67_2452_0, i_13_67_2454_0,
    i_13_67_2517_0, i_13_67_2566_0, i_13_67_3006_0, i_13_67_3009_0,
    i_13_67_3012_0, i_13_67_3037_0, i_13_67_3061_0, i_13_67_3099_0,
    i_13_67_3100_0, i_13_67_3108_0, i_13_67_3168_0, i_13_67_3173_0,
    i_13_67_3217_0, i_13_67_3274_0, i_13_67_3343_0, i_13_67_3403_0,
    i_13_67_3456_0, i_13_67_3486_0, i_13_67_3487_0, i_13_67_3537_0,
    i_13_67_3540_0, i_13_67_3541_0, i_13_67_3574_0, i_13_67_3763_0,
    i_13_67_3799_0, i_13_67_3855_0, i_13_67_3856_0, i_13_67_3864_0,
    i_13_67_3867_0, i_13_67_3892_0, i_13_67_3937_0, i_13_67_4116_0,
    i_13_67_4200_0, i_13_67_4252_0, i_13_67_4254_0, i_13_67_4255_0,
    i_13_67_4257_0, i_13_67_4258_0, i_13_67_4260_0, i_13_67_4377_0,
    i_13_67_4378_0, i_13_67_4557_0, i_13_67_4560_0,
    o_13_67_0_0  );
  input  i_13_67_64_0, i_13_67_90_0, i_13_67_91_0, i_13_67_139_0,
    i_13_67_174_0, i_13_67_175_0, i_13_67_204_0, i_13_67_228_0,
    i_13_67_229_0, i_13_67_282_0, i_13_67_283_0, i_13_67_284_0,
    i_13_67_336_0, i_13_67_337_0, i_13_67_341_0, i_13_67_393_0,
    i_13_67_414_0, i_13_67_417_0, i_13_67_450_0, i_13_67_522_0,
    i_13_67_535_0, i_13_67_567_0, i_13_67_657_0, i_13_67_661_0,
    i_13_67_733_0, i_13_67_796_0, i_13_67_823_0, i_13_67_824_0,
    i_13_67_846_0, i_13_67_847_0, i_13_67_849_0, i_13_67_850_0,
    i_13_67_981_0, i_13_67_985_0, i_13_67_1219_0, i_13_67_1224_0,
    i_13_67_1252_0, i_13_67_1263_0, i_13_67_1309_0, i_13_67_1312_0,
    i_13_67_1317_0, i_13_67_1462_0, i_13_67_1485_0, i_13_67_1549_0,
    i_13_67_1551_0, i_13_67_1552_0, i_13_67_1624_0, i_13_67_1644_0,
    i_13_67_1710_0, i_13_67_1803_0, i_13_67_1857_0, i_13_67_1858_0,
    i_13_67_1860_0, i_13_67_2197_0, i_13_67_2431_0, i_13_67_2452_0,
    i_13_67_2454_0, i_13_67_2517_0, i_13_67_2566_0, i_13_67_3006_0,
    i_13_67_3009_0, i_13_67_3012_0, i_13_67_3037_0, i_13_67_3061_0,
    i_13_67_3099_0, i_13_67_3100_0, i_13_67_3108_0, i_13_67_3168_0,
    i_13_67_3173_0, i_13_67_3217_0, i_13_67_3274_0, i_13_67_3343_0,
    i_13_67_3403_0, i_13_67_3456_0, i_13_67_3486_0, i_13_67_3487_0,
    i_13_67_3537_0, i_13_67_3540_0, i_13_67_3541_0, i_13_67_3574_0,
    i_13_67_3763_0, i_13_67_3799_0, i_13_67_3855_0, i_13_67_3856_0,
    i_13_67_3864_0, i_13_67_3867_0, i_13_67_3892_0, i_13_67_3937_0,
    i_13_67_4116_0, i_13_67_4200_0, i_13_67_4252_0, i_13_67_4254_0,
    i_13_67_4255_0, i_13_67_4257_0, i_13_67_4258_0, i_13_67_4260_0,
    i_13_67_4377_0, i_13_67_4378_0, i_13_67_4557_0, i_13_67_4560_0;
  output o_13_67_0_0;
  assign o_13_67_0_0 = ~((~i_13_67_1857_0 & ((~i_13_67_3009_0 & ~i_13_67_3856_0) | (~i_13_67_3168_0 & ~i_13_67_3173_0 & ~i_13_67_3864_0 & ~i_13_67_4378_0 & ~i_13_67_4560_0))) | (i_13_67_733_0 & i_13_67_3173_0) | (~i_13_67_414_0 & ~i_13_67_3012_0 & ~i_13_67_3108_0 & ~i_13_67_3892_0) | (i_13_67_1219_0 & ~i_13_67_4257_0) | (~i_13_67_1263_0 & ~i_13_67_4255_0 & ~i_13_67_4258_0) | (~i_13_67_282_0 & ~i_13_67_522_0 & ~i_13_67_1549_0 & i_13_67_3217_0 & ~i_13_67_4377_0));
endmodule



// Benchmark "kernel_13_68" written by ABC on Sun Jul 19 10:46:21 2020

module kernel_13_68 ( 
    i_13_68_28_0, i_13_68_48_0, i_13_68_63_0, i_13_68_64_0, i_13_68_73_0,
    i_13_68_142_0, i_13_68_144_0, i_13_68_226_0, i_13_68_279_0,
    i_13_68_282_0, i_13_68_307_0, i_13_68_315_0, i_13_68_316_0,
    i_13_68_405_0, i_13_68_532_0, i_13_68_550_0, i_13_68_604_0,
    i_13_68_639_0, i_13_68_651_0, i_13_68_666_0, i_13_68_667_0,
    i_13_68_675_0, i_13_68_676_0, i_13_68_688_0, i_13_68_757_0,
    i_13_68_868_0, i_13_68_875_0, i_13_68_931_0, i_13_68_940_0,
    i_13_68_947_0, i_13_68_1021_0, i_13_68_1099_0, i_13_68_1116_0,
    i_13_68_1207_0, i_13_68_1216_0, i_13_68_1278_0, i_13_68_1319_0,
    i_13_68_1467_0, i_13_68_1504_0, i_13_68_1522_0, i_13_68_1593_0,
    i_13_68_1594_0, i_13_68_1595_0, i_13_68_1602_0, i_13_68_1711_0,
    i_13_68_1839_0, i_13_68_1881_0, i_13_68_1990_0, i_13_68_2052_0,
    i_13_68_2053_0, i_13_68_2127_0, i_13_68_2169_0, i_13_68_2209_0,
    i_13_68_2260_0, i_13_68_2264_0, i_13_68_2277_0, i_13_68_2278_0,
    i_13_68_2380_0, i_13_68_2467_0, i_13_68_2470_0, i_13_68_2505_0,
    i_13_68_2578_0, i_13_68_2630_0, i_13_68_2674_0, i_13_68_2844_0,
    i_13_68_2845_0, i_13_68_2853_0, i_13_68_2908_0, i_13_68_2938_0,
    i_13_68_3001_0, i_13_68_3087_0, i_13_68_3096_0, i_13_68_3097_0,
    i_13_68_3108_0, i_13_68_3142_0, i_13_68_3260_0, i_13_68_3343_0,
    i_13_68_3349_0, i_13_68_3385_0, i_13_68_3501_0, i_13_68_3502_0,
    i_13_68_3525_0, i_13_68_3532_0, i_13_68_3646_0, i_13_68_3765_0,
    i_13_68_3767_0, i_13_68_3817_0, i_13_68_3888_0, i_13_68_3898_0,
    i_13_68_3907_0, i_13_68_3910_0, i_13_68_3925_0, i_13_68_4006_0,
    i_13_68_4033_0, i_13_68_4077_0, i_13_68_4107_0, i_13_68_4159_0,
    i_13_68_4186_0, i_13_68_4591_0, i_13_68_4600_0,
    o_13_68_0_0  );
  input  i_13_68_28_0, i_13_68_48_0, i_13_68_63_0, i_13_68_64_0,
    i_13_68_73_0, i_13_68_142_0, i_13_68_144_0, i_13_68_226_0,
    i_13_68_279_0, i_13_68_282_0, i_13_68_307_0, i_13_68_315_0,
    i_13_68_316_0, i_13_68_405_0, i_13_68_532_0, i_13_68_550_0,
    i_13_68_604_0, i_13_68_639_0, i_13_68_651_0, i_13_68_666_0,
    i_13_68_667_0, i_13_68_675_0, i_13_68_676_0, i_13_68_688_0,
    i_13_68_757_0, i_13_68_868_0, i_13_68_875_0, i_13_68_931_0,
    i_13_68_940_0, i_13_68_947_0, i_13_68_1021_0, i_13_68_1099_0,
    i_13_68_1116_0, i_13_68_1207_0, i_13_68_1216_0, i_13_68_1278_0,
    i_13_68_1319_0, i_13_68_1467_0, i_13_68_1504_0, i_13_68_1522_0,
    i_13_68_1593_0, i_13_68_1594_0, i_13_68_1595_0, i_13_68_1602_0,
    i_13_68_1711_0, i_13_68_1839_0, i_13_68_1881_0, i_13_68_1990_0,
    i_13_68_2052_0, i_13_68_2053_0, i_13_68_2127_0, i_13_68_2169_0,
    i_13_68_2209_0, i_13_68_2260_0, i_13_68_2264_0, i_13_68_2277_0,
    i_13_68_2278_0, i_13_68_2380_0, i_13_68_2467_0, i_13_68_2470_0,
    i_13_68_2505_0, i_13_68_2578_0, i_13_68_2630_0, i_13_68_2674_0,
    i_13_68_2844_0, i_13_68_2845_0, i_13_68_2853_0, i_13_68_2908_0,
    i_13_68_2938_0, i_13_68_3001_0, i_13_68_3087_0, i_13_68_3096_0,
    i_13_68_3097_0, i_13_68_3108_0, i_13_68_3142_0, i_13_68_3260_0,
    i_13_68_3343_0, i_13_68_3349_0, i_13_68_3385_0, i_13_68_3501_0,
    i_13_68_3502_0, i_13_68_3525_0, i_13_68_3532_0, i_13_68_3646_0,
    i_13_68_3765_0, i_13_68_3767_0, i_13_68_3817_0, i_13_68_3888_0,
    i_13_68_3898_0, i_13_68_3907_0, i_13_68_3910_0, i_13_68_3925_0,
    i_13_68_4006_0, i_13_68_4033_0, i_13_68_4077_0, i_13_68_4107_0,
    i_13_68_4159_0, i_13_68_4186_0, i_13_68_4591_0, i_13_68_4600_0;
  output o_13_68_0_0;
  assign o_13_68_0_0 = ~(i_13_68_3767_0 | (~i_13_68_2380_0 & ~i_13_68_4077_0) | (~i_13_68_1116_0 & ~i_13_68_3097_0) | (~i_13_68_2278_0 & ~i_13_68_2853_0 & ~i_13_68_3646_0 & ~i_13_68_3817_0));
endmodule



// Benchmark "kernel_13_69" written by ABC on Sun Jul 19 10:46:22 2020

module kernel_13_69 ( 
    i_13_69_48_0, i_13_69_52_0, i_13_69_75_0, i_13_69_158_0, i_13_69_182_0,
    i_13_69_213_0, i_13_69_214_0, i_13_69_277_0, i_13_69_286_0,
    i_13_69_383_0, i_13_69_526_0, i_13_69_577_0, i_13_69_578_0,
    i_13_69_582_0, i_13_69_599_0, i_13_69_618_0, i_13_69_619_0,
    i_13_69_661_0, i_13_69_697_0, i_13_69_715_0, i_13_69_792_0,
    i_13_69_937_0, i_13_69_949_0, i_13_69_1022_0, i_13_69_1076_0,
    i_13_69_1085_0, i_13_69_1141_0, i_13_69_1302_0, i_13_69_1304_0,
    i_13_69_1330_0, i_13_69_1362_0, i_13_69_1404_0, i_13_69_1492_0,
    i_13_69_1498_0, i_13_69_1500_0, i_13_69_1572_0, i_13_69_1623_0,
    i_13_69_1636_0, i_13_69_1807_0, i_13_69_1816_0, i_13_69_1817_0,
    i_13_69_2023_0, i_13_69_2107_0, i_13_69_2128_0, i_13_69_2141_0,
    i_13_69_2173_0, i_13_69_2284_0, i_13_69_2428_0, i_13_69_2440_0,
    i_13_69_2449_0, i_13_69_2452_0, i_13_69_2455_0, i_13_69_2459_0,
    i_13_69_2462_0, i_13_69_2668_0, i_13_69_2716_0, i_13_69_2753_0,
    i_13_69_2785_0, i_13_69_2787_0, i_13_69_2940_0, i_13_69_2958_0,
    i_13_69_3020_0, i_13_69_3105_0, i_13_69_3110_0, i_13_69_3143_0,
    i_13_69_3148_0, i_13_69_3231_0, i_13_69_3327_0, i_13_69_3428_0,
    i_13_69_3444_0, i_13_69_3454_0, i_13_69_3522_0, i_13_69_3523_0,
    i_13_69_3527_0, i_13_69_3553_0, i_13_69_3687_0, i_13_69_3688_0,
    i_13_69_3730_0, i_13_69_3733_0, i_13_69_3734_0, i_13_69_3757_0,
    i_13_69_3876_0, i_13_69_3911_0, i_13_69_4019_0, i_13_69_4020_0,
    i_13_69_4021_0, i_13_69_4047_0, i_13_69_4090_0, i_13_69_4093_0,
    i_13_69_4130_0, i_13_69_4254_0, i_13_69_4255_0, i_13_69_4270_0,
    i_13_69_4307_0, i_13_69_4416_0, i_13_69_4526_0, i_13_69_4539_0,
    i_13_69_4557_0, i_13_69_4559_0, i_13_69_4561_0,
    o_13_69_0_0  );
  input  i_13_69_48_0, i_13_69_52_0, i_13_69_75_0, i_13_69_158_0,
    i_13_69_182_0, i_13_69_213_0, i_13_69_214_0, i_13_69_277_0,
    i_13_69_286_0, i_13_69_383_0, i_13_69_526_0, i_13_69_577_0,
    i_13_69_578_0, i_13_69_582_0, i_13_69_599_0, i_13_69_618_0,
    i_13_69_619_0, i_13_69_661_0, i_13_69_697_0, i_13_69_715_0,
    i_13_69_792_0, i_13_69_937_0, i_13_69_949_0, i_13_69_1022_0,
    i_13_69_1076_0, i_13_69_1085_0, i_13_69_1141_0, i_13_69_1302_0,
    i_13_69_1304_0, i_13_69_1330_0, i_13_69_1362_0, i_13_69_1404_0,
    i_13_69_1492_0, i_13_69_1498_0, i_13_69_1500_0, i_13_69_1572_0,
    i_13_69_1623_0, i_13_69_1636_0, i_13_69_1807_0, i_13_69_1816_0,
    i_13_69_1817_0, i_13_69_2023_0, i_13_69_2107_0, i_13_69_2128_0,
    i_13_69_2141_0, i_13_69_2173_0, i_13_69_2284_0, i_13_69_2428_0,
    i_13_69_2440_0, i_13_69_2449_0, i_13_69_2452_0, i_13_69_2455_0,
    i_13_69_2459_0, i_13_69_2462_0, i_13_69_2668_0, i_13_69_2716_0,
    i_13_69_2753_0, i_13_69_2785_0, i_13_69_2787_0, i_13_69_2940_0,
    i_13_69_2958_0, i_13_69_3020_0, i_13_69_3105_0, i_13_69_3110_0,
    i_13_69_3143_0, i_13_69_3148_0, i_13_69_3231_0, i_13_69_3327_0,
    i_13_69_3428_0, i_13_69_3444_0, i_13_69_3454_0, i_13_69_3522_0,
    i_13_69_3523_0, i_13_69_3527_0, i_13_69_3553_0, i_13_69_3687_0,
    i_13_69_3688_0, i_13_69_3730_0, i_13_69_3733_0, i_13_69_3734_0,
    i_13_69_3757_0, i_13_69_3876_0, i_13_69_3911_0, i_13_69_4019_0,
    i_13_69_4020_0, i_13_69_4021_0, i_13_69_4047_0, i_13_69_4090_0,
    i_13_69_4093_0, i_13_69_4130_0, i_13_69_4254_0, i_13_69_4255_0,
    i_13_69_4270_0, i_13_69_4307_0, i_13_69_4416_0, i_13_69_4526_0,
    i_13_69_4539_0, i_13_69_4557_0, i_13_69_4559_0, i_13_69_4561_0;
  output o_13_69_0_0;
  assign o_13_69_0_0 = 0;
endmodule



// Benchmark "kernel_13_70" written by ABC on Sun Jul 19 10:46:23 2020

module kernel_13_70 ( 
    i_13_70_31_0, i_13_70_51_0, i_13_70_52_0, i_13_70_78_0, i_13_70_105_0,
    i_13_70_129_0, i_13_70_173_0, i_13_70_177_0, i_13_70_279_0,
    i_13_70_280_0, i_13_70_281_0, i_13_70_282_0, i_13_70_283_0,
    i_13_70_316_0, i_13_70_445_0, i_13_70_490_0, i_13_70_514_0,
    i_13_70_562_0, i_13_70_577_0, i_13_70_600_0, i_13_70_676_0,
    i_13_70_724_0, i_13_70_757_0, i_13_70_823_0, i_13_70_856_0,
    i_13_70_1018_0, i_13_70_1019_0, i_13_70_1022_0, i_13_70_1063_0,
    i_13_70_1082_0, i_13_70_1093_0, i_13_70_1143_0, i_13_70_1147_0,
    i_13_70_1526_0, i_13_70_1631_0, i_13_70_1634_0, i_13_70_1653_0,
    i_13_70_1654_0, i_13_70_1691_0, i_13_70_1786_0, i_13_70_1851_0,
    i_13_70_1940_0, i_13_70_2053_0, i_13_70_2055_0, i_13_70_2108_0,
    i_13_70_2116_0, i_13_70_2134_0, i_13_70_2198_0, i_13_70_2234_0,
    i_13_70_2236_0, i_13_70_2260_0, i_13_70_2335_0, i_13_70_2408_0,
    i_13_70_2443_0, i_13_70_2444_0, i_13_70_2506_0, i_13_70_2532_0,
    i_13_70_2543_0, i_13_70_2748_0, i_13_70_2752_0, i_13_70_3025_0,
    i_13_70_3093_0, i_13_70_3152_0, i_13_70_3165_0, i_13_70_3166_0,
    i_13_70_3175_0, i_13_70_3210_0, i_13_70_3262_0, i_13_70_3291_0,
    i_13_70_3461_0, i_13_70_3525_0, i_13_70_3539_0, i_13_70_3665_0,
    i_13_70_3727_0, i_13_70_3729_0, i_13_70_3731_0, i_13_70_3768_0,
    i_13_70_3817_0, i_13_70_3841_0, i_13_70_3854_0, i_13_70_3877_0,
    i_13_70_3889_0, i_13_70_3890_0, i_13_70_3910_0, i_13_70_3911_0,
    i_13_70_3971_0, i_13_70_3982_0, i_13_70_4015_0, i_13_70_4016_0,
    i_13_70_4063_0, i_13_70_4065_0, i_13_70_4216_0, i_13_70_4237_0,
    i_13_70_4258_0, i_13_70_4259_0, i_13_70_4297_0, i_13_70_4351_0,
    i_13_70_4375_0, i_13_70_4417_0, i_13_70_4524_0,
    o_13_70_0_0  );
  input  i_13_70_31_0, i_13_70_51_0, i_13_70_52_0, i_13_70_78_0,
    i_13_70_105_0, i_13_70_129_0, i_13_70_173_0, i_13_70_177_0,
    i_13_70_279_0, i_13_70_280_0, i_13_70_281_0, i_13_70_282_0,
    i_13_70_283_0, i_13_70_316_0, i_13_70_445_0, i_13_70_490_0,
    i_13_70_514_0, i_13_70_562_0, i_13_70_577_0, i_13_70_600_0,
    i_13_70_676_0, i_13_70_724_0, i_13_70_757_0, i_13_70_823_0,
    i_13_70_856_0, i_13_70_1018_0, i_13_70_1019_0, i_13_70_1022_0,
    i_13_70_1063_0, i_13_70_1082_0, i_13_70_1093_0, i_13_70_1143_0,
    i_13_70_1147_0, i_13_70_1526_0, i_13_70_1631_0, i_13_70_1634_0,
    i_13_70_1653_0, i_13_70_1654_0, i_13_70_1691_0, i_13_70_1786_0,
    i_13_70_1851_0, i_13_70_1940_0, i_13_70_2053_0, i_13_70_2055_0,
    i_13_70_2108_0, i_13_70_2116_0, i_13_70_2134_0, i_13_70_2198_0,
    i_13_70_2234_0, i_13_70_2236_0, i_13_70_2260_0, i_13_70_2335_0,
    i_13_70_2408_0, i_13_70_2443_0, i_13_70_2444_0, i_13_70_2506_0,
    i_13_70_2532_0, i_13_70_2543_0, i_13_70_2748_0, i_13_70_2752_0,
    i_13_70_3025_0, i_13_70_3093_0, i_13_70_3152_0, i_13_70_3165_0,
    i_13_70_3166_0, i_13_70_3175_0, i_13_70_3210_0, i_13_70_3262_0,
    i_13_70_3291_0, i_13_70_3461_0, i_13_70_3525_0, i_13_70_3539_0,
    i_13_70_3665_0, i_13_70_3727_0, i_13_70_3729_0, i_13_70_3731_0,
    i_13_70_3768_0, i_13_70_3817_0, i_13_70_3841_0, i_13_70_3854_0,
    i_13_70_3877_0, i_13_70_3889_0, i_13_70_3890_0, i_13_70_3910_0,
    i_13_70_3911_0, i_13_70_3971_0, i_13_70_3982_0, i_13_70_4015_0,
    i_13_70_4016_0, i_13_70_4063_0, i_13_70_4065_0, i_13_70_4216_0,
    i_13_70_4237_0, i_13_70_4258_0, i_13_70_4259_0, i_13_70_4297_0,
    i_13_70_4351_0, i_13_70_4375_0, i_13_70_4417_0, i_13_70_4524_0;
  output o_13_70_0_0;
  assign o_13_70_0_0 = ~((~i_13_70_3731_0 & ((~i_13_70_280_0 & ~i_13_70_4063_0) | (i_13_70_3982_0 & ~i_13_70_4375_0))) | (~i_13_70_757_0 & ~i_13_70_3817_0 & ~i_13_70_3889_0) | (i_13_70_3262_0 & ~i_13_70_4259_0));
endmodule



// Benchmark "kernel_13_71" written by ABC on Sun Jul 19 10:46:24 2020

module kernel_13_71 ( 
    i_13_71_51_0, i_13_71_52_0, i_13_71_107_0, i_13_71_111_0,
    i_13_71_117_0, i_13_71_277_0, i_13_71_340_0, i_13_71_418_0,
    i_13_71_511_0, i_13_71_561_0, i_13_71_565_0, i_13_71_618_0,
    i_13_71_628_0, i_13_71_651_0, i_13_71_745_0, i_13_71_835_0,
    i_13_71_855_0, i_13_71_915_0, i_13_71_1069_0, i_13_71_1083_0,
    i_13_71_1086_0, i_13_71_1120_0, i_13_71_1231_0, i_13_71_1335_0,
    i_13_71_1347_0, i_13_71_1363_0, i_13_71_1412_0, i_13_71_1467_0,
    i_13_71_1491_0, i_13_71_1492_0, i_13_71_1525_0, i_13_71_1572_0,
    i_13_71_1573_0, i_13_71_1623_0, i_13_71_1642_0, i_13_71_1654_0,
    i_13_71_1672_0, i_13_71_1785_0, i_13_71_1795_0, i_13_71_1806_0,
    i_13_71_1815_0, i_13_71_1906_0, i_13_71_1950_0, i_13_71_2008_0,
    i_13_71_2058_0, i_13_71_2059_0, i_13_71_2184_0, i_13_71_2283_0,
    i_13_71_2341_0, i_13_71_2353_0, i_13_71_2707_0, i_13_71_2712_0,
    i_13_71_2713_0, i_13_71_2715_0, i_13_71_2716_0, i_13_71_2787_0,
    i_13_71_2958_0, i_13_71_3010_0, i_13_71_3019_0, i_13_71_3063_0,
    i_13_71_3066_0, i_13_71_3099_0, i_13_71_3100_0, i_13_71_3156_0,
    i_13_71_3160_0, i_13_71_3165_0, i_13_71_3219_0, i_13_71_3220_0,
    i_13_71_3237_0, i_13_71_3238_0, i_13_71_3273_0, i_13_71_3291_0,
    i_13_71_3328_0, i_13_71_3346_0, i_13_71_3489_0, i_13_71_3525_0,
    i_13_71_3526_0, i_13_71_3540_0, i_13_71_3550_0, i_13_71_3552_0,
    i_13_71_3553_0, i_13_71_3598_0, i_13_71_3684_0, i_13_71_3687_0,
    i_13_71_3688_0, i_13_71_3922_0, i_13_71_4021_0, i_13_71_4047_0,
    i_13_71_4057_0, i_13_71_4065_0, i_13_71_4119_0, i_13_71_4120_0,
    i_13_71_4206_0, i_13_71_4216_0, i_13_71_4273_0, i_13_71_4387_0,
    i_13_71_4416_0, i_13_71_4452_0, i_13_71_4521_0, i_13_71_4560_0,
    o_13_71_0_0  );
  input  i_13_71_51_0, i_13_71_52_0, i_13_71_107_0, i_13_71_111_0,
    i_13_71_117_0, i_13_71_277_0, i_13_71_340_0, i_13_71_418_0,
    i_13_71_511_0, i_13_71_561_0, i_13_71_565_0, i_13_71_618_0,
    i_13_71_628_0, i_13_71_651_0, i_13_71_745_0, i_13_71_835_0,
    i_13_71_855_0, i_13_71_915_0, i_13_71_1069_0, i_13_71_1083_0,
    i_13_71_1086_0, i_13_71_1120_0, i_13_71_1231_0, i_13_71_1335_0,
    i_13_71_1347_0, i_13_71_1363_0, i_13_71_1412_0, i_13_71_1467_0,
    i_13_71_1491_0, i_13_71_1492_0, i_13_71_1525_0, i_13_71_1572_0,
    i_13_71_1573_0, i_13_71_1623_0, i_13_71_1642_0, i_13_71_1654_0,
    i_13_71_1672_0, i_13_71_1785_0, i_13_71_1795_0, i_13_71_1806_0,
    i_13_71_1815_0, i_13_71_1906_0, i_13_71_1950_0, i_13_71_2008_0,
    i_13_71_2058_0, i_13_71_2059_0, i_13_71_2184_0, i_13_71_2283_0,
    i_13_71_2341_0, i_13_71_2353_0, i_13_71_2707_0, i_13_71_2712_0,
    i_13_71_2713_0, i_13_71_2715_0, i_13_71_2716_0, i_13_71_2787_0,
    i_13_71_2958_0, i_13_71_3010_0, i_13_71_3019_0, i_13_71_3063_0,
    i_13_71_3066_0, i_13_71_3099_0, i_13_71_3100_0, i_13_71_3156_0,
    i_13_71_3160_0, i_13_71_3165_0, i_13_71_3219_0, i_13_71_3220_0,
    i_13_71_3237_0, i_13_71_3238_0, i_13_71_3273_0, i_13_71_3291_0,
    i_13_71_3328_0, i_13_71_3346_0, i_13_71_3489_0, i_13_71_3525_0,
    i_13_71_3526_0, i_13_71_3540_0, i_13_71_3550_0, i_13_71_3552_0,
    i_13_71_3553_0, i_13_71_3598_0, i_13_71_3684_0, i_13_71_3687_0,
    i_13_71_3688_0, i_13_71_3922_0, i_13_71_4021_0, i_13_71_4047_0,
    i_13_71_4057_0, i_13_71_4065_0, i_13_71_4119_0, i_13_71_4120_0,
    i_13_71_4206_0, i_13_71_4216_0, i_13_71_4273_0, i_13_71_4387_0,
    i_13_71_4416_0, i_13_71_4452_0, i_13_71_4521_0, i_13_71_4560_0;
  output o_13_71_0_0;
  assign o_13_71_0_0 = ~((~i_13_71_3165_0 & i_13_71_4216_0) | (~i_13_71_340_0 & ~i_13_71_3688_0) | (~i_13_71_1572_0 & ~i_13_71_2715_0));
endmodule



// Benchmark "kernel_13_72" written by ABC on Sun Jul 19 10:46:25 2020

module kernel_13_72 ( 
    i_13_72_68_0, i_13_72_134_0, i_13_72_138_0, i_13_72_283_0,
    i_13_72_358_0, i_13_72_359_0, i_13_72_363_0, i_13_72_400_0,
    i_13_72_472_0, i_13_72_529_0, i_13_72_661_0, i_13_72_662_0,
    i_13_72_664_0, i_13_72_665_0, i_13_72_745_0, i_13_72_827_0,
    i_13_72_835_0, i_13_72_842_0, i_13_72_854_0, i_13_72_887_0,
    i_13_72_943_0, i_13_72_949_0, i_13_72_959_0, i_13_72_1098_0,
    i_13_72_1123_0, i_13_72_1222_0, i_13_72_1229_0, i_13_72_1232_0,
    i_13_72_1259_0, i_13_72_1447_0, i_13_72_1501_0, i_13_72_1502_0,
    i_13_72_1508_0, i_13_72_1726_0, i_13_72_1745_0, i_13_72_1754_0,
    i_13_72_1951_0, i_13_72_1961_0, i_13_72_2002_0, i_13_72_2006_0,
    i_13_72_2020_0, i_13_72_2024_0, i_13_72_2033_0, i_13_72_2060_0,
    i_13_72_2104_0, i_13_72_2146_0, i_13_72_2181_0, i_13_72_2203_0,
    i_13_72_2240_0, i_13_72_2258_0, i_13_72_2284_0, i_13_72_2285_0,
    i_13_72_2344_0, i_13_72_2429_0, i_13_72_2447_0, i_13_72_2455_0,
    i_13_72_2515_0, i_13_72_2555_0, i_13_72_2696_0, i_13_72_2860_0,
    i_13_72_2885_0, i_13_72_2891_0, i_13_72_2920_0, i_13_72_3004_0,
    i_13_72_3013_0, i_13_72_3076_0, i_13_72_3172_0, i_13_72_3272_0,
    i_13_72_3404_0, i_13_72_3419_0, i_13_72_3490_0, i_13_72_3491_0,
    i_13_72_3580_0, i_13_72_3598_0, i_13_72_3599_0, i_13_72_3623_0,
    i_13_72_3757_0, i_13_72_3758_0, i_13_72_3787_0, i_13_72_3919_0,
    i_13_72_3959_0, i_13_72_3991_0, i_13_72_4122_0, i_13_72_4165_0,
    i_13_72_4166_0, i_13_72_4264_0, i_13_72_4265_0, i_13_72_4273_0,
    i_13_72_4333_0, i_13_72_4345_0, i_13_72_4382_0, i_13_72_4405_0,
    i_13_72_4433_0, i_13_72_4453_0, i_13_72_4454_0, i_13_72_4513_0,
    i_13_72_4571_0, i_13_72_4595_0, i_13_72_4597_0, i_13_72_4604_0,
    o_13_72_0_0  );
  input  i_13_72_68_0, i_13_72_134_0, i_13_72_138_0, i_13_72_283_0,
    i_13_72_358_0, i_13_72_359_0, i_13_72_363_0, i_13_72_400_0,
    i_13_72_472_0, i_13_72_529_0, i_13_72_661_0, i_13_72_662_0,
    i_13_72_664_0, i_13_72_665_0, i_13_72_745_0, i_13_72_827_0,
    i_13_72_835_0, i_13_72_842_0, i_13_72_854_0, i_13_72_887_0,
    i_13_72_943_0, i_13_72_949_0, i_13_72_959_0, i_13_72_1098_0,
    i_13_72_1123_0, i_13_72_1222_0, i_13_72_1229_0, i_13_72_1232_0,
    i_13_72_1259_0, i_13_72_1447_0, i_13_72_1501_0, i_13_72_1502_0,
    i_13_72_1508_0, i_13_72_1726_0, i_13_72_1745_0, i_13_72_1754_0,
    i_13_72_1951_0, i_13_72_1961_0, i_13_72_2002_0, i_13_72_2006_0,
    i_13_72_2020_0, i_13_72_2024_0, i_13_72_2033_0, i_13_72_2060_0,
    i_13_72_2104_0, i_13_72_2146_0, i_13_72_2181_0, i_13_72_2203_0,
    i_13_72_2240_0, i_13_72_2258_0, i_13_72_2284_0, i_13_72_2285_0,
    i_13_72_2344_0, i_13_72_2429_0, i_13_72_2447_0, i_13_72_2455_0,
    i_13_72_2515_0, i_13_72_2555_0, i_13_72_2696_0, i_13_72_2860_0,
    i_13_72_2885_0, i_13_72_2891_0, i_13_72_2920_0, i_13_72_3004_0,
    i_13_72_3013_0, i_13_72_3076_0, i_13_72_3172_0, i_13_72_3272_0,
    i_13_72_3404_0, i_13_72_3419_0, i_13_72_3490_0, i_13_72_3491_0,
    i_13_72_3580_0, i_13_72_3598_0, i_13_72_3599_0, i_13_72_3623_0,
    i_13_72_3757_0, i_13_72_3758_0, i_13_72_3787_0, i_13_72_3919_0,
    i_13_72_3959_0, i_13_72_3991_0, i_13_72_4122_0, i_13_72_4165_0,
    i_13_72_4166_0, i_13_72_4264_0, i_13_72_4265_0, i_13_72_4273_0,
    i_13_72_4333_0, i_13_72_4345_0, i_13_72_4382_0, i_13_72_4405_0,
    i_13_72_4433_0, i_13_72_4453_0, i_13_72_4454_0, i_13_72_4513_0,
    i_13_72_4571_0, i_13_72_4595_0, i_13_72_4597_0, i_13_72_4604_0;
  output o_13_72_0_0;
  assign o_13_72_0_0 = ~((~i_13_72_2696_0 & ((i_13_72_3757_0 & ~i_13_72_3758_0) | (~i_13_72_1123_0 & ~i_13_72_1754_0 & ~i_13_72_4433_0))) | (~i_13_72_4273_0 & (~i_13_72_3490_0 | (~i_13_72_1501_0 & i_13_72_2006_0 & ~i_13_72_3758_0))) | (~i_13_72_359_0 & ~i_13_72_2024_0 & ~i_13_72_2447_0 & ~i_13_72_4453_0));
endmodule



// Benchmark "kernel_13_73" written by ABC on Sun Jul 19 10:46:26 2020

module kernel_13_73 ( 
    i_13_73_33_0, i_13_73_34_0, i_13_73_40_0, i_13_73_67_0, i_13_73_138_0,
    i_13_73_139_0, i_13_73_228_0, i_13_73_232_0, i_13_73_447_0,
    i_13_73_448_0, i_13_73_457_0, i_13_73_511_0, i_13_73_529_0,
    i_13_73_535_0, i_13_73_591_0, i_13_73_615_0, i_13_73_678_0,
    i_13_73_679_0, i_13_73_695_0, i_13_73_867_0, i_13_73_872_0,
    i_13_73_985_0, i_13_73_1110_0, i_13_73_1201_0, i_13_73_1301_0,
    i_13_73_1303_0, i_13_73_1348_0, i_13_73_1409_0, i_13_73_1435_0,
    i_13_73_1438_0, i_13_73_1447_0, i_13_73_1471_0, i_13_73_1714_0,
    i_13_73_1715_0, i_13_73_1717_0, i_13_73_1723_0, i_13_73_1725_0,
    i_13_73_1740_0, i_13_73_1783_0, i_13_73_1816_0, i_13_73_1832_0,
    i_13_73_1852_0, i_13_73_1888_0, i_13_73_1889_0, i_13_73_1928_0,
    i_13_73_1938_0, i_13_73_2044_0, i_13_73_2209_0, i_13_73_2228_0,
    i_13_73_2239_0, i_13_73_2361_0, i_13_73_2380_0, i_13_73_2427_0,
    i_13_73_2938_0, i_13_73_2949_0, i_13_73_2983_0, i_13_73_3001_0,
    i_13_73_3036_0, i_13_73_3039_0, i_13_73_3104_0, i_13_73_3109_0,
    i_13_73_3111_0, i_13_73_3112_0, i_13_73_3211_0, i_13_73_3217_0,
    i_13_73_3347_0, i_13_73_3388_0, i_13_73_3390_0, i_13_73_3391_0,
    i_13_73_3598_0, i_13_73_3612_0, i_13_73_3640_0, i_13_73_3683_0,
    i_13_73_3687_0, i_13_73_3703_0, i_13_73_3741_0, i_13_73_3746_0,
    i_13_73_3766_0, i_13_73_3793_0, i_13_73_3820_0, i_13_73_3836_0,
    i_13_73_3838_0, i_13_73_3847_0, i_13_73_3848_0, i_13_73_3984_0,
    i_13_73_4038_0, i_13_73_4054_0, i_13_73_4055_0, i_13_73_4110_0,
    i_13_73_4236_0, i_13_73_4237_0, i_13_73_4318_0, i_13_73_4352_0,
    i_13_73_4369_0, i_13_73_4397_0, i_13_73_4398_0, i_13_73_4399_0,
    i_13_73_4502_0, i_13_73_4536_0, i_13_73_4567_0,
    o_13_73_0_0  );
  input  i_13_73_33_0, i_13_73_34_0, i_13_73_40_0, i_13_73_67_0,
    i_13_73_138_0, i_13_73_139_0, i_13_73_228_0, i_13_73_232_0,
    i_13_73_447_0, i_13_73_448_0, i_13_73_457_0, i_13_73_511_0,
    i_13_73_529_0, i_13_73_535_0, i_13_73_591_0, i_13_73_615_0,
    i_13_73_678_0, i_13_73_679_0, i_13_73_695_0, i_13_73_867_0,
    i_13_73_872_0, i_13_73_985_0, i_13_73_1110_0, i_13_73_1201_0,
    i_13_73_1301_0, i_13_73_1303_0, i_13_73_1348_0, i_13_73_1409_0,
    i_13_73_1435_0, i_13_73_1438_0, i_13_73_1447_0, i_13_73_1471_0,
    i_13_73_1714_0, i_13_73_1715_0, i_13_73_1717_0, i_13_73_1723_0,
    i_13_73_1725_0, i_13_73_1740_0, i_13_73_1783_0, i_13_73_1816_0,
    i_13_73_1832_0, i_13_73_1852_0, i_13_73_1888_0, i_13_73_1889_0,
    i_13_73_1928_0, i_13_73_1938_0, i_13_73_2044_0, i_13_73_2209_0,
    i_13_73_2228_0, i_13_73_2239_0, i_13_73_2361_0, i_13_73_2380_0,
    i_13_73_2427_0, i_13_73_2938_0, i_13_73_2949_0, i_13_73_2983_0,
    i_13_73_3001_0, i_13_73_3036_0, i_13_73_3039_0, i_13_73_3104_0,
    i_13_73_3109_0, i_13_73_3111_0, i_13_73_3112_0, i_13_73_3211_0,
    i_13_73_3217_0, i_13_73_3347_0, i_13_73_3388_0, i_13_73_3390_0,
    i_13_73_3391_0, i_13_73_3598_0, i_13_73_3612_0, i_13_73_3640_0,
    i_13_73_3683_0, i_13_73_3687_0, i_13_73_3703_0, i_13_73_3741_0,
    i_13_73_3746_0, i_13_73_3766_0, i_13_73_3793_0, i_13_73_3820_0,
    i_13_73_3836_0, i_13_73_3838_0, i_13_73_3847_0, i_13_73_3848_0,
    i_13_73_3984_0, i_13_73_4038_0, i_13_73_4054_0, i_13_73_4055_0,
    i_13_73_4110_0, i_13_73_4236_0, i_13_73_4237_0, i_13_73_4318_0,
    i_13_73_4352_0, i_13_73_4369_0, i_13_73_4397_0, i_13_73_4398_0,
    i_13_73_4399_0, i_13_73_4502_0, i_13_73_4536_0, i_13_73_4567_0;
  output o_13_73_0_0;
  assign o_13_73_0_0 = ~((i_13_73_985_0 & ~i_13_73_4398_0 & (~i_13_73_138_0 | ~i_13_73_4237_0)) | (~i_13_73_1717_0 & i_13_73_1832_0) | (~i_13_73_34_0 & ~i_13_73_1348_0 & ~i_13_73_1888_0) | (~i_13_73_67_0 & ~i_13_73_2239_0) | (i_13_73_2228_0 & ~i_13_73_3388_0));
endmodule



// Benchmark "kernel_13_74" written by ABC on Sun Jul 19 10:46:27 2020

module kernel_13_74 ( 
    i_13_74_64_0, i_13_74_120_0, i_13_74_192_0, i_13_74_199_0,
    i_13_74_324_0, i_13_74_361_0, i_13_74_378_0, i_13_74_379_0,
    i_13_74_441_0, i_13_74_517_0, i_13_74_531_0, i_13_74_532_0,
    i_13_74_570_0, i_13_74_571_0, i_13_74_575_0, i_13_74_576_0,
    i_13_74_588_0, i_13_74_615_0, i_13_74_639_0, i_13_74_640_0,
    i_13_74_676_0, i_13_74_678_0, i_13_74_697_0, i_13_74_698_0,
    i_13_74_714_0, i_13_74_756_0, i_13_74_820_0, i_13_74_891_0,
    i_13_74_927_0, i_13_74_928_0, i_13_74_930_0, i_13_74_931_0,
    i_13_74_1063_0, i_13_74_1080_0, i_13_74_1098_0, i_13_74_1099_0,
    i_13_74_1101_0, i_13_74_1227_0, i_13_74_1257_0, i_13_74_1270_0,
    i_13_74_1407_0, i_13_74_1503_0, i_13_74_1504_0, i_13_74_1596_0,
    i_13_74_1597_0, i_13_74_1638_0, i_13_74_1719_0, i_13_74_1746_0,
    i_13_74_1747_0, i_13_74_1782_0, i_13_74_1792_0, i_13_74_1795_0,
    i_13_74_1800_0, i_13_74_1881_0, i_13_74_1989_0, i_13_74_1990_0,
    i_13_74_2011_0, i_13_74_2116_0, i_13_74_2118_0, i_13_74_2191_0,
    i_13_74_2259_0, i_13_74_2260_0, i_13_74_2358_0, i_13_74_2458_0,
    i_13_74_2466_0, i_13_74_2505_0, i_13_74_2609_0, i_13_74_2722_0,
    i_13_74_2848_0, i_13_74_2881_0, i_13_74_2901_0, i_13_74_2934_0,
    i_13_74_3000_0, i_13_74_3024_0, i_13_74_3027_0, i_13_74_3060_0,
    i_13_74_3114_0, i_13_74_3204_0, i_13_74_3259_0, i_13_74_3286_0,
    i_13_74_3420_0, i_13_74_3421_0, i_13_74_3448_0, i_13_74_3537_0,
    i_13_74_3753_0, i_13_74_3781_0, i_13_74_3790_0, i_13_74_3808_0,
    i_13_74_3811_0, i_13_74_3873_0, i_13_74_3924_0, i_13_74_3925_0,
    i_13_74_3928_0, i_13_74_3936_0, i_13_74_4008_0, i_13_74_4009_0,
    i_13_74_4077_0, i_13_74_4078_0, i_13_74_4086_0, i_13_74_4231_0,
    o_13_74_0_0  );
  input  i_13_74_64_0, i_13_74_120_0, i_13_74_192_0, i_13_74_199_0,
    i_13_74_324_0, i_13_74_361_0, i_13_74_378_0, i_13_74_379_0,
    i_13_74_441_0, i_13_74_517_0, i_13_74_531_0, i_13_74_532_0,
    i_13_74_570_0, i_13_74_571_0, i_13_74_575_0, i_13_74_576_0,
    i_13_74_588_0, i_13_74_615_0, i_13_74_639_0, i_13_74_640_0,
    i_13_74_676_0, i_13_74_678_0, i_13_74_697_0, i_13_74_698_0,
    i_13_74_714_0, i_13_74_756_0, i_13_74_820_0, i_13_74_891_0,
    i_13_74_927_0, i_13_74_928_0, i_13_74_930_0, i_13_74_931_0,
    i_13_74_1063_0, i_13_74_1080_0, i_13_74_1098_0, i_13_74_1099_0,
    i_13_74_1101_0, i_13_74_1227_0, i_13_74_1257_0, i_13_74_1270_0,
    i_13_74_1407_0, i_13_74_1503_0, i_13_74_1504_0, i_13_74_1596_0,
    i_13_74_1597_0, i_13_74_1638_0, i_13_74_1719_0, i_13_74_1746_0,
    i_13_74_1747_0, i_13_74_1782_0, i_13_74_1792_0, i_13_74_1795_0,
    i_13_74_1800_0, i_13_74_1881_0, i_13_74_1989_0, i_13_74_1990_0,
    i_13_74_2011_0, i_13_74_2116_0, i_13_74_2118_0, i_13_74_2191_0,
    i_13_74_2259_0, i_13_74_2260_0, i_13_74_2358_0, i_13_74_2458_0,
    i_13_74_2466_0, i_13_74_2505_0, i_13_74_2609_0, i_13_74_2722_0,
    i_13_74_2848_0, i_13_74_2881_0, i_13_74_2901_0, i_13_74_2934_0,
    i_13_74_3000_0, i_13_74_3024_0, i_13_74_3027_0, i_13_74_3060_0,
    i_13_74_3114_0, i_13_74_3204_0, i_13_74_3259_0, i_13_74_3286_0,
    i_13_74_3420_0, i_13_74_3421_0, i_13_74_3448_0, i_13_74_3537_0,
    i_13_74_3753_0, i_13_74_3781_0, i_13_74_3790_0, i_13_74_3808_0,
    i_13_74_3811_0, i_13_74_3873_0, i_13_74_3924_0, i_13_74_3925_0,
    i_13_74_3928_0, i_13_74_3936_0, i_13_74_4008_0, i_13_74_4009_0,
    i_13_74_4077_0, i_13_74_4078_0, i_13_74_4086_0, i_13_74_4231_0;
  output o_13_74_0_0;
  assign o_13_74_0_0 = ~((~i_13_74_4077_0 & (i_13_74_697_0 | ~i_13_74_3259_0 | (~i_13_74_1792_0 & ~i_13_74_3448_0))) | (i_13_74_1597_0 & ~i_13_74_1746_0 & ~i_13_74_2934_0) | (~i_13_74_379_0 & ~i_13_74_927_0 & ~i_13_74_2848_0 & ~i_13_74_3928_0));
endmodule



// Benchmark "kernel_13_75" written by ABC on Sun Jul 19 10:46:28 2020

module kernel_13_75 ( 
    i_13_75_49_0, i_13_75_166_0, i_13_75_245_0, i_13_75_262_0,
    i_13_75_266_0, i_13_75_375_0, i_13_75_382_0, i_13_75_417_0,
    i_13_75_446_0, i_13_75_464_0, i_13_75_490_0, i_13_75_571_0,
    i_13_75_589_0, i_13_75_607_0, i_13_75_760_0, i_13_75_761_0,
    i_13_75_771_0, i_13_75_812_0, i_13_75_814_0, i_13_75_823_0,
    i_13_75_862_0, i_13_75_987_0, i_13_75_1066_0, i_13_75_1137_0,
    i_13_75_1147_0, i_13_75_1196_0, i_13_75_1228_0, i_13_75_1343_0,
    i_13_75_1489_0, i_13_75_1502_0, i_13_75_1558_0, i_13_75_1598_0,
    i_13_75_1760_0, i_13_75_1840_0, i_13_75_1841_0, i_13_75_1849_0,
    i_13_75_1853_0, i_13_75_1859_0, i_13_75_1931_0, i_13_75_1994_0,
    i_13_75_2137_0, i_13_75_2149_0, i_13_75_2179_0, i_13_75_2183_0,
    i_13_75_2192_0, i_13_75_2207_0, i_13_75_2263_0, i_13_75_2266_0,
    i_13_75_2346_0, i_13_75_2380_0, i_13_75_2396_0, i_13_75_2400_0,
    i_13_75_2408_0, i_13_75_2411_0, i_13_75_2469_0, i_13_75_2533_0,
    i_13_75_2696_0, i_13_75_2722_0, i_13_75_2749_0, i_13_75_2760_0,
    i_13_75_2769_0, i_13_75_2786_0, i_13_75_2857_0, i_13_75_2884_0,
    i_13_75_2938_0, i_13_75_2941_0, i_13_75_3028_0, i_13_75_3034_0,
    i_13_75_3047_0, i_13_75_3068_0, i_13_75_3218_0, i_13_75_3262_0,
    i_13_75_3316_0, i_13_75_3341_0, i_13_75_3343_0, i_13_75_3371_0,
    i_13_75_3394_0, i_13_75_3413_0, i_13_75_3442_0, i_13_75_3475_0,
    i_13_75_3506_0, i_13_75_3542_0, i_13_75_3630_0, i_13_75_3664_0,
    i_13_75_3667_0, i_13_75_3668_0, i_13_75_3750_0, i_13_75_3920_0,
    i_13_75_4009_0, i_13_75_4015_0, i_13_75_4061_0, i_13_75_4063_0,
    i_13_75_4162_0, i_13_75_4171_0, i_13_75_4315_0, i_13_75_4316_0,
    i_13_75_4317_0, i_13_75_4318_0, i_13_75_4369_0, i_13_75_4396_0,
    o_13_75_0_0  );
  input  i_13_75_49_0, i_13_75_166_0, i_13_75_245_0, i_13_75_262_0,
    i_13_75_266_0, i_13_75_375_0, i_13_75_382_0, i_13_75_417_0,
    i_13_75_446_0, i_13_75_464_0, i_13_75_490_0, i_13_75_571_0,
    i_13_75_589_0, i_13_75_607_0, i_13_75_760_0, i_13_75_761_0,
    i_13_75_771_0, i_13_75_812_0, i_13_75_814_0, i_13_75_823_0,
    i_13_75_862_0, i_13_75_987_0, i_13_75_1066_0, i_13_75_1137_0,
    i_13_75_1147_0, i_13_75_1196_0, i_13_75_1228_0, i_13_75_1343_0,
    i_13_75_1489_0, i_13_75_1502_0, i_13_75_1558_0, i_13_75_1598_0,
    i_13_75_1760_0, i_13_75_1840_0, i_13_75_1841_0, i_13_75_1849_0,
    i_13_75_1853_0, i_13_75_1859_0, i_13_75_1931_0, i_13_75_1994_0,
    i_13_75_2137_0, i_13_75_2149_0, i_13_75_2179_0, i_13_75_2183_0,
    i_13_75_2192_0, i_13_75_2207_0, i_13_75_2263_0, i_13_75_2266_0,
    i_13_75_2346_0, i_13_75_2380_0, i_13_75_2396_0, i_13_75_2400_0,
    i_13_75_2408_0, i_13_75_2411_0, i_13_75_2469_0, i_13_75_2533_0,
    i_13_75_2696_0, i_13_75_2722_0, i_13_75_2749_0, i_13_75_2760_0,
    i_13_75_2769_0, i_13_75_2786_0, i_13_75_2857_0, i_13_75_2884_0,
    i_13_75_2938_0, i_13_75_2941_0, i_13_75_3028_0, i_13_75_3034_0,
    i_13_75_3047_0, i_13_75_3068_0, i_13_75_3218_0, i_13_75_3262_0,
    i_13_75_3316_0, i_13_75_3341_0, i_13_75_3343_0, i_13_75_3371_0,
    i_13_75_3394_0, i_13_75_3413_0, i_13_75_3442_0, i_13_75_3475_0,
    i_13_75_3506_0, i_13_75_3542_0, i_13_75_3630_0, i_13_75_3664_0,
    i_13_75_3667_0, i_13_75_3668_0, i_13_75_3750_0, i_13_75_3920_0,
    i_13_75_4009_0, i_13_75_4015_0, i_13_75_4061_0, i_13_75_4063_0,
    i_13_75_4162_0, i_13_75_4171_0, i_13_75_4315_0, i_13_75_4316_0,
    i_13_75_4317_0, i_13_75_4318_0, i_13_75_4369_0, i_13_75_4396_0;
  output o_13_75_0_0;
  assign o_13_75_0_0 = ~((~i_13_75_382_0 & ((i_13_75_1228_0 & ~i_13_75_2137_0 & ~i_13_75_2941_0) | (i_13_75_3506_0 & ~i_13_75_4315_0))) | (i_13_75_862_0 & ~i_13_75_2857_0 & ~i_13_75_2941_0 & i_13_75_3506_0) | (i_13_75_1147_0 & ~i_13_75_2380_0 & i_13_75_3394_0) | (~i_13_75_49_0 & ~i_13_75_812_0 & i_13_75_823_0 & ~i_13_75_2411_0 & ~i_13_75_3316_0 & ~i_13_75_3920_0) | (~i_13_75_862_0 & ~i_13_75_4063_0) | (~i_13_75_2696_0 & i_13_75_3262_0 & ~i_13_75_4162_0));
endmodule



// Benchmark "kernel_13_76" written by ABC on Sun Jul 19 10:46:28 2020

module kernel_13_76 ( 
    i_13_76_19_0, i_13_76_80_0, i_13_76_111_0, i_13_76_113_0,
    i_13_76_125_0, i_13_76_241_0, i_13_76_242_0, i_13_76_277_0,
    i_13_76_278_0, i_13_76_336_0, i_13_76_386_0, i_13_76_418_0,
    i_13_76_558_0, i_13_76_619_0, i_13_76_643_0, i_13_76_696_0,
    i_13_76_718_0, i_13_76_741_0, i_13_76_779_0, i_13_76_855_0,
    i_13_76_910_0, i_13_76_1017_0, i_13_76_1083_0, i_13_76_1084_0,
    i_13_76_1085_0, i_13_76_1087_0, i_13_76_1092_0, i_13_76_1381_0,
    i_13_76_1569_0, i_13_76_1620_0, i_13_76_1623_0, i_13_76_1624_0,
    i_13_76_1637_0, i_13_76_1642_0, i_13_76_1710_0, i_13_76_1774_0,
    i_13_76_1817_0, i_13_76_1840_0, i_13_76_1918_0, i_13_76_1952_0,
    i_13_76_1990_0, i_13_76_2174_0, i_13_76_2185_0, i_13_76_2348_0,
    i_13_76_2358_0, i_13_76_2433_0, i_13_76_2497_0, i_13_76_2548_0,
    i_13_76_2610_0, i_13_76_2712_0, i_13_76_2713_0, i_13_76_2716_0,
    i_13_76_2717_0, i_13_76_2739_0, i_13_76_2788_0, i_13_76_2921_0,
    i_13_76_2959_0, i_13_76_3047_0, i_13_76_3067_0, i_13_76_3097_0,
    i_13_76_3100_0, i_13_76_3101_0, i_13_76_3141_0, i_13_76_3145_0,
    i_13_76_3167_0, i_13_76_3221_0, i_13_76_3302_0, i_13_76_3312_0,
    i_13_76_3329_0, i_13_76_3374_0, i_13_76_3450_0, i_13_76_3454_0,
    i_13_76_3484_0, i_13_76_3486_0, i_13_76_3549_0, i_13_76_3553_0,
    i_13_76_3576_0, i_13_76_3684_0, i_13_76_3685_0, i_13_76_3688_0,
    i_13_76_3689_0, i_13_76_3736_0, i_13_76_3738_0, i_13_76_3878_0,
    i_13_76_3913_0, i_13_76_4022_0, i_13_76_4036_0, i_13_76_4050_0,
    i_13_76_4066_0, i_13_76_4081_0, i_13_76_4174_0, i_13_76_4269_0,
    i_13_76_4274_0, i_13_76_4328_0, i_13_76_4356_0, i_13_76_4363_0,
    i_13_76_4417_0, i_13_76_4522_0, i_13_76_4526_0, i_13_76_4536_0,
    o_13_76_0_0  );
  input  i_13_76_19_0, i_13_76_80_0, i_13_76_111_0, i_13_76_113_0,
    i_13_76_125_0, i_13_76_241_0, i_13_76_242_0, i_13_76_277_0,
    i_13_76_278_0, i_13_76_336_0, i_13_76_386_0, i_13_76_418_0,
    i_13_76_558_0, i_13_76_619_0, i_13_76_643_0, i_13_76_696_0,
    i_13_76_718_0, i_13_76_741_0, i_13_76_779_0, i_13_76_855_0,
    i_13_76_910_0, i_13_76_1017_0, i_13_76_1083_0, i_13_76_1084_0,
    i_13_76_1085_0, i_13_76_1087_0, i_13_76_1092_0, i_13_76_1381_0,
    i_13_76_1569_0, i_13_76_1620_0, i_13_76_1623_0, i_13_76_1624_0,
    i_13_76_1637_0, i_13_76_1642_0, i_13_76_1710_0, i_13_76_1774_0,
    i_13_76_1817_0, i_13_76_1840_0, i_13_76_1918_0, i_13_76_1952_0,
    i_13_76_1990_0, i_13_76_2174_0, i_13_76_2185_0, i_13_76_2348_0,
    i_13_76_2358_0, i_13_76_2433_0, i_13_76_2497_0, i_13_76_2548_0,
    i_13_76_2610_0, i_13_76_2712_0, i_13_76_2713_0, i_13_76_2716_0,
    i_13_76_2717_0, i_13_76_2739_0, i_13_76_2788_0, i_13_76_2921_0,
    i_13_76_2959_0, i_13_76_3047_0, i_13_76_3067_0, i_13_76_3097_0,
    i_13_76_3100_0, i_13_76_3101_0, i_13_76_3141_0, i_13_76_3145_0,
    i_13_76_3167_0, i_13_76_3221_0, i_13_76_3302_0, i_13_76_3312_0,
    i_13_76_3329_0, i_13_76_3374_0, i_13_76_3450_0, i_13_76_3454_0,
    i_13_76_3484_0, i_13_76_3486_0, i_13_76_3549_0, i_13_76_3553_0,
    i_13_76_3576_0, i_13_76_3684_0, i_13_76_3685_0, i_13_76_3688_0,
    i_13_76_3689_0, i_13_76_3736_0, i_13_76_3738_0, i_13_76_3878_0,
    i_13_76_3913_0, i_13_76_4022_0, i_13_76_4036_0, i_13_76_4050_0,
    i_13_76_4066_0, i_13_76_4081_0, i_13_76_4174_0, i_13_76_4269_0,
    i_13_76_4274_0, i_13_76_4328_0, i_13_76_4356_0, i_13_76_4363_0,
    i_13_76_4417_0, i_13_76_4522_0, i_13_76_4526_0, i_13_76_4536_0;
  output o_13_76_0_0;
  assign o_13_76_0_0 = 0;
endmodule



// Benchmark "kernel_13_77" written by ABC on Sun Jul 19 10:46:29 2020

module kernel_13_77 ( 
    i_13_77_43_0, i_13_77_49_0, i_13_77_80_0, i_13_77_115_0, i_13_77_196_0,
    i_13_77_265_0, i_13_77_277_0, i_13_77_278_0, i_13_77_310_0,
    i_13_77_352_0, i_13_77_377_0, i_13_77_405_0, i_13_77_454_0,
    i_13_77_476_0, i_13_77_520_0, i_13_77_562_0, i_13_77_563_0,
    i_13_77_578_0, i_13_77_582_0, i_13_77_661_0, i_13_77_664_0,
    i_13_77_665_0, i_13_77_673_0, i_13_77_741_0, i_13_77_823_0,
    i_13_77_833_0, i_13_77_850_0, i_13_77_935_0, i_13_77_1145_0,
    i_13_77_1327_0, i_13_77_1333_0, i_13_77_1364_0, i_13_77_1473_0,
    i_13_77_1508_0, i_13_77_1552_0, i_13_77_1627_0, i_13_77_1730_0,
    i_13_77_1732_0, i_13_77_1735_0, i_13_77_1754_0, i_13_77_1768_0,
    i_13_77_1841_0, i_13_77_1844_0, i_13_77_1864_0, i_13_77_2003_0,
    i_13_77_2018_0, i_13_77_2019_0, i_13_77_2020_0, i_13_77_2024_0,
    i_13_77_2098_0, i_13_77_2149_0, i_13_77_2265_0, i_13_77_2300_0,
    i_13_77_2452_0, i_13_77_2471_0, i_13_77_2519_0, i_13_77_2653_0,
    i_13_77_2708_0, i_13_77_2712_0, i_13_77_2743_0, i_13_77_2744_0,
    i_13_77_2898_0, i_13_77_2955_0, i_13_77_3007_0, i_13_77_3050_0,
    i_13_77_3100_0, i_13_77_3118_0, i_13_77_3234_0, i_13_77_3266_0,
    i_13_77_3316_0, i_13_77_3351_0, i_13_77_3418_0, i_13_77_3453_0,
    i_13_77_3464_0, i_13_77_3479_0, i_13_77_3553_0, i_13_77_3571_0,
    i_13_77_3604_0, i_13_77_3730_0, i_13_77_3757_0, i_13_77_3781_0,
    i_13_77_3799_0, i_13_77_3823_0, i_13_77_3904_0, i_13_77_3905_0,
    i_13_77_3972_0, i_13_77_4056_0, i_13_77_4122_0, i_13_77_4130_0,
    i_13_77_4162_0, i_13_77_4163_0, i_13_77_4165_0, i_13_77_4166_0,
    i_13_77_4237_0, i_13_77_4370_0, i_13_77_4432_0, i_13_77_4513_0,
    i_13_77_4517_0, i_13_77_4555_0, i_13_77_4607_0,
    o_13_77_0_0  );
  input  i_13_77_43_0, i_13_77_49_0, i_13_77_80_0, i_13_77_115_0,
    i_13_77_196_0, i_13_77_265_0, i_13_77_277_0, i_13_77_278_0,
    i_13_77_310_0, i_13_77_352_0, i_13_77_377_0, i_13_77_405_0,
    i_13_77_454_0, i_13_77_476_0, i_13_77_520_0, i_13_77_562_0,
    i_13_77_563_0, i_13_77_578_0, i_13_77_582_0, i_13_77_661_0,
    i_13_77_664_0, i_13_77_665_0, i_13_77_673_0, i_13_77_741_0,
    i_13_77_823_0, i_13_77_833_0, i_13_77_850_0, i_13_77_935_0,
    i_13_77_1145_0, i_13_77_1327_0, i_13_77_1333_0, i_13_77_1364_0,
    i_13_77_1473_0, i_13_77_1508_0, i_13_77_1552_0, i_13_77_1627_0,
    i_13_77_1730_0, i_13_77_1732_0, i_13_77_1735_0, i_13_77_1754_0,
    i_13_77_1768_0, i_13_77_1841_0, i_13_77_1844_0, i_13_77_1864_0,
    i_13_77_2003_0, i_13_77_2018_0, i_13_77_2019_0, i_13_77_2020_0,
    i_13_77_2024_0, i_13_77_2098_0, i_13_77_2149_0, i_13_77_2265_0,
    i_13_77_2300_0, i_13_77_2452_0, i_13_77_2471_0, i_13_77_2519_0,
    i_13_77_2653_0, i_13_77_2708_0, i_13_77_2712_0, i_13_77_2743_0,
    i_13_77_2744_0, i_13_77_2898_0, i_13_77_2955_0, i_13_77_3007_0,
    i_13_77_3050_0, i_13_77_3100_0, i_13_77_3118_0, i_13_77_3234_0,
    i_13_77_3266_0, i_13_77_3316_0, i_13_77_3351_0, i_13_77_3418_0,
    i_13_77_3453_0, i_13_77_3464_0, i_13_77_3479_0, i_13_77_3553_0,
    i_13_77_3571_0, i_13_77_3604_0, i_13_77_3730_0, i_13_77_3757_0,
    i_13_77_3781_0, i_13_77_3799_0, i_13_77_3823_0, i_13_77_3904_0,
    i_13_77_3905_0, i_13_77_3972_0, i_13_77_4056_0, i_13_77_4122_0,
    i_13_77_4130_0, i_13_77_4162_0, i_13_77_4163_0, i_13_77_4165_0,
    i_13_77_4166_0, i_13_77_4237_0, i_13_77_4370_0, i_13_77_4432_0,
    i_13_77_4513_0, i_13_77_4517_0, i_13_77_4555_0, i_13_77_4607_0;
  output o_13_77_0_0;
  assign o_13_77_0_0 = ~((~i_13_77_3905_0 & ((~i_13_77_935_0 & ~i_13_77_1145_0 & ~i_13_77_4165_0) | (~i_13_77_80_0 & ~i_13_77_520_0 & ~i_13_77_4370_0 & ~i_13_77_4432_0))) | (i_13_77_4555_0 & (~i_13_77_1768_0 | (i_13_77_3730_0 & ~i_13_77_4513_0))) | (~i_13_77_1732_0 & ~i_13_77_1735_0) | (~i_13_77_2020_0 & ~i_13_77_2744_0 & ~i_13_77_3100_0) | (~i_13_77_115_0 & ~i_13_77_3553_0 & ~i_13_77_3604_0) | (~i_13_77_277_0 & ~i_13_77_1627_0 & ~i_13_77_2300_0 & ~i_13_77_3904_0));
endmodule



// Benchmark "kernel_13_78" written by ABC on Sun Jul 19 10:46:30 2020

module kernel_13_78 ( 
    i_13_78_39_0, i_13_78_49_0, i_13_78_79_0, i_13_78_285_0, i_13_78_327_0,
    i_13_78_340_0, i_13_78_528_0, i_13_78_530_0, i_13_78_672_0,
    i_13_78_673_0, i_13_78_717_0, i_13_78_797_0, i_13_78_825_0,
    i_13_78_862_0, i_13_78_894_0, i_13_78_1023_0, i_13_78_1024_0,
    i_13_78_1029_0, i_13_78_1258_0, i_13_78_1300_0, i_13_78_1320_0,
    i_13_78_1321_0, i_13_78_1383_0, i_13_78_1489_0, i_13_78_1500_0,
    i_13_78_1543_0, i_13_78_1552_0, i_13_78_1732_0, i_13_78_1743_0,
    i_13_78_1857_0, i_13_78_1884_0, i_13_78_1933_0, i_13_78_1947_0,
    i_13_78_1960_0, i_13_78_2014_0, i_13_78_2015_0, i_13_78_2032_0,
    i_13_78_2136_0, i_13_78_2139_0, i_13_78_2190_0, i_13_78_2204_0,
    i_13_78_2229_0, i_13_78_2460_0, i_13_78_2461_0, i_13_78_2463_0,
    i_13_78_2464_0, i_13_78_2595_0, i_13_78_2613_0, i_13_78_2652_0,
    i_13_78_2824_0, i_13_78_2874_0, i_13_78_2922_0, i_13_78_2923_0,
    i_13_78_2983_0, i_13_78_3174_0, i_13_78_3321_0, i_13_78_3322_0,
    i_13_78_3406_0, i_13_78_3417_0, i_13_78_3418_0, i_13_78_3432_0,
    i_13_78_3498_0, i_13_78_3522_0, i_13_78_3540_0, i_13_78_3541_0,
    i_13_78_3543_0, i_13_78_3550_0, i_13_78_3579_0, i_13_78_3613_0,
    i_13_78_3730_0, i_13_78_3731_0, i_13_78_3732_0, i_13_78_3733_0,
    i_13_78_3768_0, i_13_78_3769_0, i_13_78_3786_0, i_13_78_3787_0,
    i_13_78_3805_0, i_13_78_3831_0, i_13_78_3858_0, i_13_78_3912_0,
    i_13_78_3913_0, i_13_78_3931_0, i_13_78_3994_0, i_13_78_4117_0,
    i_13_78_4161_0, i_13_78_4188_0, i_13_78_4237_0, i_13_78_4255_0,
    i_13_78_4263_0, i_13_78_4296_0, i_13_78_4341_0, i_13_78_4380_0,
    i_13_78_4381_0, i_13_78_4414_0, i_13_78_4443_0, i_13_78_4567_0,
    i_13_78_4587_0, i_13_78_4597_0, i_13_78_4602_0,
    o_13_78_0_0  );
  input  i_13_78_39_0, i_13_78_49_0, i_13_78_79_0, i_13_78_285_0,
    i_13_78_327_0, i_13_78_340_0, i_13_78_528_0, i_13_78_530_0,
    i_13_78_672_0, i_13_78_673_0, i_13_78_717_0, i_13_78_797_0,
    i_13_78_825_0, i_13_78_862_0, i_13_78_894_0, i_13_78_1023_0,
    i_13_78_1024_0, i_13_78_1029_0, i_13_78_1258_0, i_13_78_1300_0,
    i_13_78_1320_0, i_13_78_1321_0, i_13_78_1383_0, i_13_78_1489_0,
    i_13_78_1500_0, i_13_78_1543_0, i_13_78_1552_0, i_13_78_1732_0,
    i_13_78_1743_0, i_13_78_1857_0, i_13_78_1884_0, i_13_78_1933_0,
    i_13_78_1947_0, i_13_78_1960_0, i_13_78_2014_0, i_13_78_2015_0,
    i_13_78_2032_0, i_13_78_2136_0, i_13_78_2139_0, i_13_78_2190_0,
    i_13_78_2204_0, i_13_78_2229_0, i_13_78_2460_0, i_13_78_2461_0,
    i_13_78_2463_0, i_13_78_2464_0, i_13_78_2595_0, i_13_78_2613_0,
    i_13_78_2652_0, i_13_78_2824_0, i_13_78_2874_0, i_13_78_2922_0,
    i_13_78_2923_0, i_13_78_2983_0, i_13_78_3174_0, i_13_78_3321_0,
    i_13_78_3322_0, i_13_78_3406_0, i_13_78_3417_0, i_13_78_3418_0,
    i_13_78_3432_0, i_13_78_3498_0, i_13_78_3522_0, i_13_78_3540_0,
    i_13_78_3541_0, i_13_78_3543_0, i_13_78_3550_0, i_13_78_3579_0,
    i_13_78_3613_0, i_13_78_3730_0, i_13_78_3731_0, i_13_78_3732_0,
    i_13_78_3733_0, i_13_78_3768_0, i_13_78_3769_0, i_13_78_3786_0,
    i_13_78_3787_0, i_13_78_3805_0, i_13_78_3831_0, i_13_78_3858_0,
    i_13_78_3912_0, i_13_78_3913_0, i_13_78_3931_0, i_13_78_3994_0,
    i_13_78_4117_0, i_13_78_4161_0, i_13_78_4188_0, i_13_78_4237_0,
    i_13_78_4255_0, i_13_78_4263_0, i_13_78_4296_0, i_13_78_4341_0,
    i_13_78_4380_0, i_13_78_4381_0, i_13_78_4414_0, i_13_78_4443_0,
    i_13_78_4567_0, i_13_78_4587_0, i_13_78_4597_0, i_13_78_4602_0;
  output o_13_78_0_0;
  assign o_13_78_0_0 = ~(~i_13_78_1321_0 | (~i_13_78_3913_0 & i_13_78_4161_0) | (~i_13_78_3858_0 & ~i_13_78_4263_0 & ~i_13_78_4380_0));
endmodule



// Benchmark "kernel_13_79" written by ABC on Sun Jul 19 10:46:31 2020

module kernel_13_79 ( 
    i_13_79_94_0, i_13_79_95_0, i_13_79_98_0, i_13_79_106_0, i_13_79_107_0,
    i_13_79_179_0, i_13_79_187_0, i_13_79_278_0, i_13_79_283_0,
    i_13_79_310_0, i_13_79_311_0, i_13_79_313_0, i_13_79_314_0,
    i_13_79_316_0, i_13_79_318_0, i_13_79_319_0, i_13_79_320_0,
    i_13_79_323_0, i_13_79_508_0, i_13_79_554_0, i_13_79_567_0,
    i_13_79_575_0, i_13_79_607_0, i_13_79_647_0, i_13_79_689_0,
    i_13_79_692_0, i_13_79_707_0, i_13_79_821_0, i_13_79_837_0,
    i_13_79_973_0, i_13_79_981_0, i_13_79_982_0, i_13_79_1024_0,
    i_13_79_1070_0, i_13_79_1101_0, i_13_79_1115_0, i_13_79_1123_0,
    i_13_79_1124_0, i_13_79_1184_0, i_13_79_1327_0, i_13_79_1394_0,
    i_13_79_1408_0, i_13_79_1471_0, i_13_79_1574_0, i_13_79_1609_0,
    i_13_79_1754_0, i_13_79_1773_0, i_13_79_1796_0, i_13_79_1859_0,
    i_13_79_1889_0, i_13_79_1931_0, i_13_79_1992_0, i_13_79_2123_0,
    i_13_79_2266_0, i_13_79_2267_0, i_13_79_2277_0, i_13_79_2403_0,
    i_13_79_2411_0, i_13_79_2494_0, i_13_79_2503_0, i_13_79_2545_0,
    i_13_79_2614_0, i_13_79_2680_0, i_13_79_2681_0, i_13_79_2699_0,
    i_13_79_2768_0, i_13_79_2824_0, i_13_79_2986_0, i_13_79_3065_0,
    i_13_79_3068_0, i_13_79_3130_0, i_13_79_3157_0, i_13_79_3167_0,
    i_13_79_3211_0, i_13_79_3212_0, i_13_79_3275_0, i_13_79_3339_0,
    i_13_79_3347_0, i_13_79_3392_0, i_13_79_3410_0, i_13_79_3416_0,
    i_13_79_3460_0, i_13_79_3544_0, i_13_79_3646_0, i_13_79_3685_0,
    i_13_79_3689_0, i_13_79_3799_0, i_13_79_3928_0, i_13_79_3931_0,
    i_13_79_4037_0, i_13_79_4080_0, i_13_79_4085_0, i_13_79_4270_0,
    i_13_79_4309_0, i_13_79_4342_0, i_13_79_4354_0, i_13_79_4369_0,
    i_13_79_4534_0, i_13_79_4570_0, i_13_79_4598_0,
    o_13_79_0_0  );
  input  i_13_79_94_0, i_13_79_95_0, i_13_79_98_0, i_13_79_106_0,
    i_13_79_107_0, i_13_79_179_0, i_13_79_187_0, i_13_79_278_0,
    i_13_79_283_0, i_13_79_310_0, i_13_79_311_0, i_13_79_313_0,
    i_13_79_314_0, i_13_79_316_0, i_13_79_318_0, i_13_79_319_0,
    i_13_79_320_0, i_13_79_323_0, i_13_79_508_0, i_13_79_554_0,
    i_13_79_567_0, i_13_79_575_0, i_13_79_607_0, i_13_79_647_0,
    i_13_79_689_0, i_13_79_692_0, i_13_79_707_0, i_13_79_821_0,
    i_13_79_837_0, i_13_79_973_0, i_13_79_981_0, i_13_79_982_0,
    i_13_79_1024_0, i_13_79_1070_0, i_13_79_1101_0, i_13_79_1115_0,
    i_13_79_1123_0, i_13_79_1124_0, i_13_79_1184_0, i_13_79_1327_0,
    i_13_79_1394_0, i_13_79_1408_0, i_13_79_1471_0, i_13_79_1574_0,
    i_13_79_1609_0, i_13_79_1754_0, i_13_79_1773_0, i_13_79_1796_0,
    i_13_79_1859_0, i_13_79_1889_0, i_13_79_1931_0, i_13_79_1992_0,
    i_13_79_2123_0, i_13_79_2266_0, i_13_79_2267_0, i_13_79_2277_0,
    i_13_79_2403_0, i_13_79_2411_0, i_13_79_2494_0, i_13_79_2503_0,
    i_13_79_2545_0, i_13_79_2614_0, i_13_79_2680_0, i_13_79_2681_0,
    i_13_79_2699_0, i_13_79_2768_0, i_13_79_2824_0, i_13_79_2986_0,
    i_13_79_3065_0, i_13_79_3068_0, i_13_79_3130_0, i_13_79_3157_0,
    i_13_79_3167_0, i_13_79_3211_0, i_13_79_3212_0, i_13_79_3275_0,
    i_13_79_3339_0, i_13_79_3347_0, i_13_79_3392_0, i_13_79_3410_0,
    i_13_79_3416_0, i_13_79_3460_0, i_13_79_3544_0, i_13_79_3646_0,
    i_13_79_3685_0, i_13_79_3689_0, i_13_79_3799_0, i_13_79_3928_0,
    i_13_79_3931_0, i_13_79_4037_0, i_13_79_4080_0, i_13_79_4085_0,
    i_13_79_4270_0, i_13_79_4309_0, i_13_79_4342_0, i_13_79_4354_0,
    i_13_79_4369_0, i_13_79_4534_0, i_13_79_4570_0, i_13_79_4598_0;
  output o_13_79_0_0;
  assign o_13_79_0_0 = ~((~i_13_79_313_0 & ((~i_13_79_821_0 & i_13_79_2614_0 & ~i_13_79_2681_0 & ~i_13_79_3931_0) | (~i_13_79_982_0 & ~i_13_79_3167_0 & i_13_79_4270_0))) | (~i_13_79_323_0 & ((~i_13_79_310_0 & ~i_13_79_1754_0 & ~i_13_79_2986_0) | (i_13_79_1574_0 & ~i_13_79_4570_0))) | (~i_13_79_1992_0 & ((~i_13_79_319_0 & ~i_13_79_320_0 & ~i_13_79_2681_0) | (~i_13_79_95_0 & ~i_13_79_187_0 & ~i_13_79_4085_0 & ~i_13_79_4354_0))) | (~i_13_79_2986_0 & (i_13_79_278_0 | i_13_79_1574_0)) | (~i_13_79_1859_0 & ~i_13_79_3167_0 & ~i_13_79_3931_0 & i_13_79_4270_0) | (~i_13_79_1408_0 & i_13_79_1992_0 & i_13_79_4570_0));
endmodule



// Benchmark "kernel_13_80" written by ABC on Sun Jul 19 10:46:32 2020

module kernel_13_80 ( 
    i_13_80_93_0, i_13_80_94_0, i_13_80_170_0, i_13_80_179_0,
    i_13_80_188_0, i_13_80_258_0, i_13_80_307_0, i_13_80_310_0,
    i_13_80_319_0, i_13_80_451_0, i_13_80_575_0, i_13_80_670_0,
    i_13_80_697_0, i_13_80_812_0, i_13_80_822_0, i_13_80_979_0,
    i_13_80_1020_0, i_13_80_1021_0, i_13_80_1023_0, i_13_80_1024_0,
    i_13_80_1077_0, i_13_80_1078_0, i_13_80_1138_0, i_13_80_1179_0,
    i_13_80_1219_0, i_13_80_1228_0, i_13_80_1273_0, i_13_80_1317_0,
    i_13_80_1318_0, i_13_80_1320_0, i_13_80_1429_0, i_13_80_1438_0,
    i_13_80_1608_0, i_13_80_1631_0, i_13_80_1633_0, i_13_80_1779_0,
    i_13_80_1780_0, i_13_80_1840_0, i_13_80_1853_0, i_13_80_1857_0,
    i_13_80_1920_0, i_13_80_2026_0, i_13_80_2136_0, i_13_80_2172_0,
    i_13_80_2200_0, i_13_80_2213_0, i_13_80_2245_0, i_13_80_2267_0,
    i_13_80_2399_0, i_13_80_2434_0, i_13_80_2454_0, i_13_80_2509_0,
    i_13_80_2571_0, i_13_80_2616_0, i_13_80_2617_0, i_13_80_2707_0,
    i_13_80_2749_0, i_13_80_2767_0, i_13_80_2787_0, i_13_80_2912_0,
    i_13_80_2983_0, i_13_80_3002_0, i_13_80_3094_0, i_13_80_3113_0,
    i_13_80_3171_0, i_13_80_3172_0, i_13_80_3209_0, i_13_80_3271_0,
    i_13_80_3326_0, i_13_80_3460_0, i_13_80_3463_0, i_13_80_3464_0,
    i_13_80_3534_0, i_13_80_3541_0, i_13_80_3544_0, i_13_80_3576_0,
    i_13_80_3664_0, i_13_80_3784_0, i_13_80_3821_0, i_13_80_3850_0,
    i_13_80_3855_0, i_13_80_3877_0, i_13_80_3894_0, i_13_80_3913_0,
    i_13_80_3927_0, i_13_80_4036_0, i_13_80_4067_0, i_13_80_4099_0,
    i_13_80_4178_0, i_13_80_4219_0, i_13_80_4255_0, i_13_80_4351_0,
    i_13_80_4353_0, i_13_80_4354_0, i_13_80_4381_0, i_13_80_4395_0,
    i_13_80_4431_0, i_13_80_4450_0, i_13_80_4556_0, i_13_80_4567_0,
    o_13_80_0_0  );
  input  i_13_80_93_0, i_13_80_94_0, i_13_80_170_0, i_13_80_179_0,
    i_13_80_188_0, i_13_80_258_0, i_13_80_307_0, i_13_80_310_0,
    i_13_80_319_0, i_13_80_451_0, i_13_80_575_0, i_13_80_670_0,
    i_13_80_697_0, i_13_80_812_0, i_13_80_822_0, i_13_80_979_0,
    i_13_80_1020_0, i_13_80_1021_0, i_13_80_1023_0, i_13_80_1024_0,
    i_13_80_1077_0, i_13_80_1078_0, i_13_80_1138_0, i_13_80_1179_0,
    i_13_80_1219_0, i_13_80_1228_0, i_13_80_1273_0, i_13_80_1317_0,
    i_13_80_1318_0, i_13_80_1320_0, i_13_80_1429_0, i_13_80_1438_0,
    i_13_80_1608_0, i_13_80_1631_0, i_13_80_1633_0, i_13_80_1779_0,
    i_13_80_1780_0, i_13_80_1840_0, i_13_80_1853_0, i_13_80_1857_0,
    i_13_80_1920_0, i_13_80_2026_0, i_13_80_2136_0, i_13_80_2172_0,
    i_13_80_2200_0, i_13_80_2213_0, i_13_80_2245_0, i_13_80_2267_0,
    i_13_80_2399_0, i_13_80_2434_0, i_13_80_2454_0, i_13_80_2509_0,
    i_13_80_2571_0, i_13_80_2616_0, i_13_80_2617_0, i_13_80_2707_0,
    i_13_80_2749_0, i_13_80_2767_0, i_13_80_2787_0, i_13_80_2912_0,
    i_13_80_2983_0, i_13_80_3002_0, i_13_80_3094_0, i_13_80_3113_0,
    i_13_80_3171_0, i_13_80_3172_0, i_13_80_3209_0, i_13_80_3271_0,
    i_13_80_3326_0, i_13_80_3460_0, i_13_80_3463_0, i_13_80_3464_0,
    i_13_80_3534_0, i_13_80_3541_0, i_13_80_3544_0, i_13_80_3576_0,
    i_13_80_3664_0, i_13_80_3784_0, i_13_80_3821_0, i_13_80_3850_0,
    i_13_80_3855_0, i_13_80_3877_0, i_13_80_3894_0, i_13_80_3913_0,
    i_13_80_3927_0, i_13_80_4036_0, i_13_80_4067_0, i_13_80_4099_0,
    i_13_80_4178_0, i_13_80_4219_0, i_13_80_4255_0, i_13_80_4351_0,
    i_13_80_4353_0, i_13_80_4354_0, i_13_80_4381_0, i_13_80_4395_0,
    i_13_80_4431_0, i_13_80_4450_0, i_13_80_4556_0, i_13_80_4567_0;
  output o_13_80_0_0;
  assign o_13_80_0_0 = ~((~i_13_80_3172_0 & i_13_80_4067_0) | (~i_13_80_1320_0 & ~i_13_80_3463_0) | (~i_13_80_2200_0 & ~i_13_80_2616_0) | (~i_13_80_179_0 & i_13_80_3464_0 & i_13_80_4381_0) | (~i_13_80_1317_0 & ~i_13_80_2767_0 & ~i_13_80_3113_0 & ~i_13_80_4381_0));
endmodule



// Benchmark "kernel_13_81" written by ABC on Sun Jul 19 10:46:33 2020

module kernel_13_81 ( 
    i_13_81_51_0, i_13_81_52_0, i_13_81_75_0, i_13_81_120_0, i_13_81_121_0,
    i_13_81_138_0, i_13_81_183_0, i_13_81_240_0, i_13_81_250_0,
    i_13_81_338_0, i_13_81_339_0, i_13_81_357_0, i_13_81_373_0,
    i_13_81_392_0, i_13_81_465_0, i_13_81_529_0, i_13_81_561_0,
    i_13_81_596_0, i_13_81_655_0, i_13_81_663_0, i_13_81_714_0,
    i_13_81_743_0, i_13_81_937_0, i_13_81_941_0, i_13_81_942_0,
    i_13_81_1077_0, i_13_81_1100_0, i_13_81_1211_0, i_13_81_1212_0,
    i_13_81_1397_0, i_13_81_1407_0, i_13_81_1408_0, i_13_81_1424_0,
    i_13_81_1469_0, i_13_81_1500_0, i_13_81_1501_0, i_13_81_1507_0,
    i_13_81_1523_0, i_13_81_1572_0, i_13_81_1608_0, i_13_81_1635_0,
    i_13_81_1636_0, i_13_81_1695_0, i_13_81_1722_0, i_13_81_1730_0,
    i_13_81_1775_0, i_13_81_1920_0, i_13_81_1951_0, i_13_81_1992_0,
    i_13_81_2031_0, i_13_81_2032_0, i_13_81_2058_0, i_13_81_2117_0,
    i_13_81_2169_0, i_13_81_2284_0, i_13_81_2343_0, i_13_81_2425_0,
    i_13_81_2455_0, i_13_81_2545_0, i_13_81_2724_0, i_13_81_2767_0,
    i_13_81_2787_0, i_13_81_2882_0, i_13_81_2923_0, i_13_81_2958_0,
    i_13_81_3061_0, i_13_81_3087_0, i_13_81_3088_0, i_13_81_3291_0,
    i_13_81_3372_0, i_13_81_3373_0, i_13_81_3417_0, i_13_81_3418_0,
    i_13_81_3427_0, i_13_81_3448_0, i_13_81_3463_0, i_13_81_3469_0,
    i_13_81_3489_0, i_13_81_3579_0, i_13_81_3597_0, i_13_81_3598_0,
    i_13_81_3633_0, i_13_81_3647_0, i_13_81_3649_0, i_13_81_3682_0,
    i_13_81_3687_0, i_13_81_3733_0, i_13_81_3767_0, i_13_81_3903_0,
    i_13_81_3990_0, i_13_81_4191_0, i_13_81_4249_0, i_13_81_4250_0,
    i_13_81_4263_0, i_13_81_4264_0, i_13_81_4412_0, i_13_81_4430_0,
    i_13_81_4452_0, i_13_81_4453_0, i_13_81_4541_0,
    o_13_81_0_0  );
  input  i_13_81_51_0, i_13_81_52_0, i_13_81_75_0, i_13_81_120_0,
    i_13_81_121_0, i_13_81_138_0, i_13_81_183_0, i_13_81_240_0,
    i_13_81_250_0, i_13_81_338_0, i_13_81_339_0, i_13_81_357_0,
    i_13_81_373_0, i_13_81_392_0, i_13_81_465_0, i_13_81_529_0,
    i_13_81_561_0, i_13_81_596_0, i_13_81_655_0, i_13_81_663_0,
    i_13_81_714_0, i_13_81_743_0, i_13_81_937_0, i_13_81_941_0,
    i_13_81_942_0, i_13_81_1077_0, i_13_81_1100_0, i_13_81_1211_0,
    i_13_81_1212_0, i_13_81_1397_0, i_13_81_1407_0, i_13_81_1408_0,
    i_13_81_1424_0, i_13_81_1469_0, i_13_81_1500_0, i_13_81_1501_0,
    i_13_81_1507_0, i_13_81_1523_0, i_13_81_1572_0, i_13_81_1608_0,
    i_13_81_1635_0, i_13_81_1636_0, i_13_81_1695_0, i_13_81_1722_0,
    i_13_81_1730_0, i_13_81_1775_0, i_13_81_1920_0, i_13_81_1951_0,
    i_13_81_1992_0, i_13_81_2031_0, i_13_81_2032_0, i_13_81_2058_0,
    i_13_81_2117_0, i_13_81_2169_0, i_13_81_2284_0, i_13_81_2343_0,
    i_13_81_2425_0, i_13_81_2455_0, i_13_81_2545_0, i_13_81_2724_0,
    i_13_81_2767_0, i_13_81_2787_0, i_13_81_2882_0, i_13_81_2923_0,
    i_13_81_2958_0, i_13_81_3061_0, i_13_81_3087_0, i_13_81_3088_0,
    i_13_81_3291_0, i_13_81_3372_0, i_13_81_3373_0, i_13_81_3417_0,
    i_13_81_3418_0, i_13_81_3427_0, i_13_81_3448_0, i_13_81_3463_0,
    i_13_81_3469_0, i_13_81_3489_0, i_13_81_3579_0, i_13_81_3597_0,
    i_13_81_3598_0, i_13_81_3633_0, i_13_81_3647_0, i_13_81_3649_0,
    i_13_81_3682_0, i_13_81_3687_0, i_13_81_3733_0, i_13_81_3767_0,
    i_13_81_3903_0, i_13_81_3990_0, i_13_81_4191_0, i_13_81_4249_0,
    i_13_81_4250_0, i_13_81_4263_0, i_13_81_4264_0, i_13_81_4412_0,
    i_13_81_4430_0, i_13_81_4452_0, i_13_81_4453_0, i_13_81_4541_0;
  output o_13_81_0_0;
  assign o_13_81_0_0 = 0;
endmodule



// Benchmark "kernel_13_82" written by ABC on Sun Jul 19 10:46:34 2020

module kernel_13_82 ( 
    i_13_82_40_0, i_13_82_46_0, i_13_82_76_0, i_13_82_172_0, i_13_82_264_0,
    i_13_82_279_0, i_13_82_282_0, i_13_82_283_0, i_13_82_337_0,
    i_13_82_378_0, i_13_82_525_0, i_13_82_693_0, i_13_82_697_0,
    i_13_82_1021_0, i_13_82_1066_0, i_13_82_1081_0, i_13_82_1082_0,
    i_13_82_1120_0, i_13_82_1224_0, i_13_82_1270_0, i_13_82_1306_0,
    i_13_82_1323_0, i_13_82_1401_0, i_13_82_1444_0, i_13_82_1495_0,
    i_13_82_1497_0, i_13_82_1498_0, i_13_82_1541_0, i_13_82_1566_0,
    i_13_82_1569_0, i_13_82_1633_0, i_13_82_1634_0, i_13_82_1783_0,
    i_13_82_1802_0, i_13_82_1916_0, i_13_82_1921_0, i_13_82_1927_0,
    i_13_82_1984_0, i_13_82_1990_0, i_13_82_1991_0, i_13_82_2001_0,
    i_13_82_2034_0, i_13_82_2037_0, i_13_82_2092_0, i_13_82_2117_0,
    i_13_82_2128_0, i_13_82_2177_0, i_13_82_2363_0, i_13_82_2424_0,
    i_13_82_2425_0, i_13_82_2430_0, i_13_82_2431_0, i_13_82_2449_0,
    i_13_82_2461_0, i_13_82_2548_0, i_13_82_2551_0, i_13_82_2601_0,
    i_13_82_2660_0, i_13_82_2674_0, i_13_82_2675_0, i_13_82_2934_0,
    i_13_82_2936_0, i_13_82_3004_0, i_13_82_3127_0, i_13_82_3142_0,
    i_13_82_3268_0, i_13_82_3269_0, i_13_82_3272_0, i_13_82_3393_0,
    i_13_82_3406_0, i_13_82_3421_0, i_13_82_3424_0, i_13_82_3582_0,
    i_13_82_3647_0, i_13_82_3727_0, i_13_82_3728_0, i_13_82_3730_0,
    i_13_82_3872_0, i_13_82_3987_0, i_13_82_4010_0, i_13_82_4014_0,
    i_13_82_4015_0, i_13_82_4016_0, i_13_82_4051_0, i_13_82_4087_0,
    i_13_82_4088_0, i_13_82_4120_0, i_13_82_4171_0, i_13_82_4224_0,
    i_13_82_4225_0, i_13_82_4249_0, i_13_82_4252_0, i_13_82_4261_0,
    i_13_82_4268_0, i_13_82_4297_0, i_13_82_4305_0, i_13_82_4393_0,
    i_13_82_4404_0, i_13_82_4475_0, i_13_82_4558_0,
    o_13_82_0_0  );
  input  i_13_82_40_0, i_13_82_46_0, i_13_82_76_0, i_13_82_172_0,
    i_13_82_264_0, i_13_82_279_0, i_13_82_282_0, i_13_82_283_0,
    i_13_82_337_0, i_13_82_378_0, i_13_82_525_0, i_13_82_693_0,
    i_13_82_697_0, i_13_82_1021_0, i_13_82_1066_0, i_13_82_1081_0,
    i_13_82_1082_0, i_13_82_1120_0, i_13_82_1224_0, i_13_82_1270_0,
    i_13_82_1306_0, i_13_82_1323_0, i_13_82_1401_0, i_13_82_1444_0,
    i_13_82_1495_0, i_13_82_1497_0, i_13_82_1498_0, i_13_82_1541_0,
    i_13_82_1566_0, i_13_82_1569_0, i_13_82_1633_0, i_13_82_1634_0,
    i_13_82_1783_0, i_13_82_1802_0, i_13_82_1916_0, i_13_82_1921_0,
    i_13_82_1927_0, i_13_82_1984_0, i_13_82_1990_0, i_13_82_1991_0,
    i_13_82_2001_0, i_13_82_2034_0, i_13_82_2037_0, i_13_82_2092_0,
    i_13_82_2117_0, i_13_82_2128_0, i_13_82_2177_0, i_13_82_2363_0,
    i_13_82_2424_0, i_13_82_2425_0, i_13_82_2430_0, i_13_82_2431_0,
    i_13_82_2449_0, i_13_82_2461_0, i_13_82_2548_0, i_13_82_2551_0,
    i_13_82_2601_0, i_13_82_2660_0, i_13_82_2674_0, i_13_82_2675_0,
    i_13_82_2934_0, i_13_82_2936_0, i_13_82_3004_0, i_13_82_3127_0,
    i_13_82_3142_0, i_13_82_3268_0, i_13_82_3269_0, i_13_82_3272_0,
    i_13_82_3393_0, i_13_82_3406_0, i_13_82_3421_0, i_13_82_3424_0,
    i_13_82_3582_0, i_13_82_3647_0, i_13_82_3727_0, i_13_82_3728_0,
    i_13_82_3730_0, i_13_82_3872_0, i_13_82_3987_0, i_13_82_4010_0,
    i_13_82_4014_0, i_13_82_4015_0, i_13_82_4016_0, i_13_82_4051_0,
    i_13_82_4087_0, i_13_82_4088_0, i_13_82_4120_0, i_13_82_4171_0,
    i_13_82_4224_0, i_13_82_4225_0, i_13_82_4249_0, i_13_82_4252_0,
    i_13_82_4261_0, i_13_82_4268_0, i_13_82_4297_0, i_13_82_4305_0,
    i_13_82_4393_0, i_13_82_4404_0, i_13_82_4475_0, i_13_82_4558_0;
  output o_13_82_0_0;
  assign o_13_82_0_0 = ~((~i_13_82_697_0 & ((~i_13_82_1306_0 & ~i_13_82_2001_0 & ~i_13_82_3142_0) | (~i_13_82_1802_0 & ~i_13_82_2424_0 & ~i_13_82_3872_0 & ~i_13_82_4087_0 & ~i_13_82_4088_0 & ~i_13_82_4249_0 & ~i_13_82_4268_0))) | (~i_13_82_1497_0 & ((~i_13_82_3142_0 & ~i_13_82_3727_0 & ~i_13_82_4010_0) | (i_13_82_697_0 & ~i_13_82_2936_0 & ~i_13_82_4249_0))) | (~i_13_82_2425_0 & ((i_13_82_1082_0 & ~i_13_82_3142_0) | (~i_13_82_1990_0 & ~i_13_82_3730_0))) | (~i_13_82_2449_0 & ((~i_13_82_1991_0 & i_13_82_2551_0) | (~i_13_82_282_0 & ~i_13_82_378_0 & i_13_82_2425_0 & ~i_13_82_2674_0))) | (~i_13_82_1224_0 & ~i_13_82_1495_0 & i_13_82_2128_0 & ~i_13_82_2675_0) | (i_13_82_1066_0 & ~i_13_82_3727_0 & ~i_13_82_3987_0) | (~i_13_82_172_0 & ~i_13_82_1498_0 & ~i_13_82_4249_0 & ~i_13_82_4558_0));
endmodule



// Benchmark "kernel_13_83" written by ABC on Sun Jul 19 10:46:35 2020

module kernel_13_83 ( 
    i_13_83_73_0, i_13_83_74_0, i_13_83_76_0, i_13_83_104_0, i_13_83_109_0,
    i_13_83_110_0, i_13_83_112_0, i_13_83_116_0, i_13_83_122_0,
    i_13_83_193_0, i_13_83_284_0, i_13_83_287_0, i_13_83_320_0,
    i_13_83_368_0, i_13_83_376_0, i_13_83_407_0, i_13_83_559_0,
    i_13_83_586_0, i_13_83_589_0, i_13_83_605_0, i_13_83_652_0,
    i_13_83_757_0, i_13_83_856_0, i_13_83_859_0, i_13_83_1021_0,
    i_13_83_1076_0, i_13_83_1086_0, i_13_83_1087_0, i_13_83_1217_0,
    i_13_83_1219_0, i_13_83_1273_0, i_13_83_1274_0, i_13_83_1474_0,
    i_13_83_1486_0, i_13_83_1567_0, i_13_83_1574_0, i_13_83_1630_0,
    i_13_83_1634_0, i_13_83_1678_0, i_13_83_1719_0, i_13_83_1775_0,
    i_13_83_1778_0, i_13_83_1837_0, i_13_83_1841_0, i_13_83_1849_0,
    i_13_83_1945_0, i_13_83_2137_0, i_13_83_2175_0, i_13_83_2192_0,
    i_13_83_2263_0, i_13_83_2423_0, i_13_83_2434_0, i_13_83_2435_0,
    i_13_83_2437_0, i_13_83_2438_0, i_13_83_2462_0, i_13_83_2465_0,
    i_13_83_2501_0, i_13_83_2535_0, i_13_83_2542_0, i_13_83_2716_0,
    i_13_83_2722_0, i_13_83_2920_0, i_13_83_3098_0, i_13_83_3101_0,
    i_13_83_3102_0, i_13_83_3143_0, i_13_83_3145_0, i_13_83_3146_0,
    i_13_83_3167_0, i_13_83_3290_0, i_13_83_3385_0, i_13_83_3452_0,
    i_13_83_3453_0, i_13_83_3478_0, i_13_83_3530_0, i_13_83_3532_0,
    i_13_83_3570_0, i_13_83_3578_0, i_13_83_3734_0, i_13_83_3764_0,
    i_13_83_3874_0, i_13_83_3938_0, i_13_83_4021_0, i_13_83_4036_0,
    i_13_83_4051_0, i_13_83_4093_0, i_13_83_4120_0, i_13_83_4121_0,
    i_13_83_4254_0, i_13_83_4255_0, i_13_83_4282_0, i_13_83_4283_0,
    i_13_83_4325_0, i_13_83_4366_0, i_13_83_4379_0, i_13_83_4524_0,
    i_13_83_4541_0, i_13_83_4559_0, i_13_83_4562_0,
    o_13_83_0_0  );
  input  i_13_83_73_0, i_13_83_74_0, i_13_83_76_0, i_13_83_104_0,
    i_13_83_109_0, i_13_83_110_0, i_13_83_112_0, i_13_83_116_0,
    i_13_83_122_0, i_13_83_193_0, i_13_83_284_0, i_13_83_287_0,
    i_13_83_320_0, i_13_83_368_0, i_13_83_376_0, i_13_83_407_0,
    i_13_83_559_0, i_13_83_586_0, i_13_83_589_0, i_13_83_605_0,
    i_13_83_652_0, i_13_83_757_0, i_13_83_856_0, i_13_83_859_0,
    i_13_83_1021_0, i_13_83_1076_0, i_13_83_1086_0, i_13_83_1087_0,
    i_13_83_1217_0, i_13_83_1219_0, i_13_83_1273_0, i_13_83_1274_0,
    i_13_83_1474_0, i_13_83_1486_0, i_13_83_1567_0, i_13_83_1574_0,
    i_13_83_1630_0, i_13_83_1634_0, i_13_83_1678_0, i_13_83_1719_0,
    i_13_83_1775_0, i_13_83_1778_0, i_13_83_1837_0, i_13_83_1841_0,
    i_13_83_1849_0, i_13_83_1945_0, i_13_83_2137_0, i_13_83_2175_0,
    i_13_83_2192_0, i_13_83_2263_0, i_13_83_2423_0, i_13_83_2434_0,
    i_13_83_2435_0, i_13_83_2437_0, i_13_83_2438_0, i_13_83_2462_0,
    i_13_83_2465_0, i_13_83_2501_0, i_13_83_2535_0, i_13_83_2542_0,
    i_13_83_2716_0, i_13_83_2722_0, i_13_83_2920_0, i_13_83_3098_0,
    i_13_83_3101_0, i_13_83_3102_0, i_13_83_3143_0, i_13_83_3145_0,
    i_13_83_3146_0, i_13_83_3167_0, i_13_83_3290_0, i_13_83_3385_0,
    i_13_83_3452_0, i_13_83_3453_0, i_13_83_3478_0, i_13_83_3530_0,
    i_13_83_3532_0, i_13_83_3570_0, i_13_83_3578_0, i_13_83_3734_0,
    i_13_83_3764_0, i_13_83_3874_0, i_13_83_3938_0, i_13_83_4021_0,
    i_13_83_4036_0, i_13_83_4051_0, i_13_83_4093_0, i_13_83_4120_0,
    i_13_83_4121_0, i_13_83_4254_0, i_13_83_4255_0, i_13_83_4282_0,
    i_13_83_4283_0, i_13_83_4325_0, i_13_83_4366_0, i_13_83_4379_0,
    i_13_83_4524_0, i_13_83_4541_0, i_13_83_4559_0, i_13_83_4562_0;
  output o_13_83_0_0;
  assign o_13_83_0_0 = ~((~i_13_83_110_0 & ((~i_13_83_284_0 & ~i_13_83_1219_0) | (~i_13_83_2542_0 & ~i_13_83_3578_0 & ~i_13_83_3734_0))) | (~i_13_83_3764_0 & (i_13_83_586_0 | (~i_13_83_3167_0 & ~i_13_83_3578_0 & ~i_13_83_4255_0 & ~i_13_83_4366_0))) | (~i_13_83_4562_0 & ((i_13_83_193_0 & i_13_83_1273_0) | (~i_13_83_73_0 & i_13_83_589_0 & ~i_13_83_2423_0 & ~i_13_83_3385_0 & ~i_13_83_3874_0))) | (~i_13_83_112_0 & i_13_83_1849_0 & ~i_13_83_4036_0) | (~i_13_83_1021_0 & ~i_13_83_4093_0 & i_13_83_4562_0));
endmodule



// Benchmark "kernel_13_84" written by ABC on Sun Jul 19 10:46:36 2020

module kernel_13_84 ( 
    i_13_84_35_0, i_13_84_171_0, i_13_84_192_0, i_13_84_193_0,
    i_13_84_199_0, i_13_84_256_0, i_13_84_382_0, i_13_84_450_0,
    i_13_84_567_0, i_13_84_585_0, i_13_84_626_0, i_13_84_639_0,
    i_13_84_640_0, i_13_84_660_0, i_13_84_927_0, i_13_84_939_0,
    i_13_84_955_0, i_13_84_1062_0, i_13_84_1116_0, i_13_84_1121_0,
    i_13_84_1147_0, i_13_84_1192_0, i_13_84_1224_0, i_13_84_1225_0,
    i_13_84_1227_0, i_13_84_1228_0, i_13_84_1255_0, i_13_84_1314_0,
    i_13_84_1341_0, i_13_84_1407_0, i_13_84_1488_0, i_13_84_1494_0,
    i_13_84_1512_0, i_13_84_1521_0, i_13_84_1534_0, i_13_84_1552_0,
    i_13_84_1567_0, i_13_84_1570_0, i_13_84_1677_0, i_13_84_1724_0,
    i_13_84_1764_0, i_13_84_1765_0, i_13_84_1767_0, i_13_84_1801_0,
    i_13_84_1890_0, i_13_84_1891_0, i_13_84_1926_0, i_13_84_1956_0,
    i_13_84_1990_0, i_13_84_2044_0, i_13_84_2055_0, i_13_84_2056_0,
    i_13_84_2092_0, i_13_84_2240_0, i_13_84_2300_0, i_13_84_2568_0,
    i_13_84_2614_0, i_13_84_2646_0, i_13_84_2691_0, i_13_84_2781_0,
    i_13_84_2899_0, i_13_84_2934_0, i_13_84_2935_0, i_13_84_3006_0,
    i_13_84_3025_0, i_13_84_3118_0, i_13_84_3136_0, i_13_84_3144_0,
    i_13_84_3164_0, i_13_84_3214_0, i_13_84_3230_0, i_13_84_3267_0,
    i_13_84_3285_0, i_13_84_3286_0, i_13_84_3312_0, i_13_84_3339_0,
    i_13_84_3420_0, i_13_84_3421_0, i_13_84_3478_0, i_13_84_3531_0,
    i_13_84_3537_0, i_13_84_3901_0, i_13_84_3918_0, i_13_84_3978_0,
    i_13_84_3986_0, i_13_84_4009_0, i_13_84_4042_0, i_13_84_4077_0,
    i_13_84_4086_0, i_13_84_4087_0, i_13_84_4185_0, i_13_84_4248_0,
    i_13_84_4266_0, i_13_84_4267_0, i_13_84_4293_0, i_13_84_4302_0,
    i_13_84_4351_0, i_13_84_4368_0, i_13_84_4375_0, i_13_84_4468_0,
    o_13_84_0_0  );
  input  i_13_84_35_0, i_13_84_171_0, i_13_84_192_0, i_13_84_193_0,
    i_13_84_199_0, i_13_84_256_0, i_13_84_382_0, i_13_84_450_0,
    i_13_84_567_0, i_13_84_585_0, i_13_84_626_0, i_13_84_639_0,
    i_13_84_640_0, i_13_84_660_0, i_13_84_927_0, i_13_84_939_0,
    i_13_84_955_0, i_13_84_1062_0, i_13_84_1116_0, i_13_84_1121_0,
    i_13_84_1147_0, i_13_84_1192_0, i_13_84_1224_0, i_13_84_1225_0,
    i_13_84_1227_0, i_13_84_1228_0, i_13_84_1255_0, i_13_84_1314_0,
    i_13_84_1341_0, i_13_84_1407_0, i_13_84_1488_0, i_13_84_1494_0,
    i_13_84_1512_0, i_13_84_1521_0, i_13_84_1534_0, i_13_84_1552_0,
    i_13_84_1567_0, i_13_84_1570_0, i_13_84_1677_0, i_13_84_1724_0,
    i_13_84_1764_0, i_13_84_1765_0, i_13_84_1767_0, i_13_84_1801_0,
    i_13_84_1890_0, i_13_84_1891_0, i_13_84_1926_0, i_13_84_1956_0,
    i_13_84_1990_0, i_13_84_2044_0, i_13_84_2055_0, i_13_84_2056_0,
    i_13_84_2092_0, i_13_84_2240_0, i_13_84_2300_0, i_13_84_2568_0,
    i_13_84_2614_0, i_13_84_2646_0, i_13_84_2691_0, i_13_84_2781_0,
    i_13_84_2899_0, i_13_84_2934_0, i_13_84_2935_0, i_13_84_3006_0,
    i_13_84_3025_0, i_13_84_3118_0, i_13_84_3136_0, i_13_84_3144_0,
    i_13_84_3164_0, i_13_84_3214_0, i_13_84_3230_0, i_13_84_3267_0,
    i_13_84_3285_0, i_13_84_3286_0, i_13_84_3312_0, i_13_84_3339_0,
    i_13_84_3420_0, i_13_84_3421_0, i_13_84_3478_0, i_13_84_3531_0,
    i_13_84_3537_0, i_13_84_3901_0, i_13_84_3918_0, i_13_84_3978_0,
    i_13_84_3986_0, i_13_84_4009_0, i_13_84_4042_0, i_13_84_4077_0,
    i_13_84_4086_0, i_13_84_4087_0, i_13_84_4185_0, i_13_84_4248_0,
    i_13_84_4266_0, i_13_84_4267_0, i_13_84_4293_0, i_13_84_4302_0,
    i_13_84_4351_0, i_13_84_4368_0, i_13_84_4375_0, i_13_84_4468_0;
  output o_13_84_0_0;
  assign o_13_84_0_0 = ~((~i_13_84_2646_0 & ~i_13_84_4302_0) | (~i_13_84_1801_0 & ~i_13_84_4042_0) | (~i_13_84_192_0 & ~i_13_84_3537_0));
endmodule



// Benchmark "kernel_13_85" written by ABC on Sun Jul 19 10:46:37 2020

module kernel_13_85 ( 
    i_13_85_67_0, i_13_85_282_0, i_13_85_285_0, i_13_85_384_0,
    i_13_85_385_0, i_13_85_448_0, i_13_85_456_0, i_13_85_625_0,
    i_13_85_669_0, i_13_85_745_0, i_13_85_796_0, i_13_85_816_0,
    i_13_85_852_0, i_13_85_865_0, i_13_85_889_0, i_13_85_948_0,
    i_13_85_1068_0, i_13_85_1101_0, i_13_85_1120_0, i_13_85_1259_0,
    i_13_85_1272_0, i_13_85_1273_0, i_13_85_1302_0, i_13_85_1303_0,
    i_13_85_1312_0, i_13_85_1390_0, i_13_85_1402_0, i_13_85_1484_0,
    i_13_85_1507_0, i_13_85_1573_0, i_13_85_1632_0, i_13_85_1642_0,
    i_13_85_1768_0, i_13_85_1777_0, i_13_85_1794_0, i_13_85_1795_0,
    i_13_85_1851_0, i_13_85_1933_0, i_13_85_1995_0, i_13_85_1996_0,
    i_13_85_2001_0, i_13_85_2014_0, i_13_85_2122_0, i_13_85_2211_0,
    i_13_85_2256_0, i_13_85_2266_0, i_13_85_2380_0, i_13_85_2427_0,
    i_13_85_2433_0, i_13_85_2434_0, i_13_85_2461_0, i_13_85_2463_0,
    i_13_85_2464_0, i_13_85_2470_0, i_13_85_2541_0, i_13_85_2754_0,
    i_13_85_2796_0, i_13_85_2884_0, i_13_85_2905_0, i_13_85_2916_0,
    i_13_85_2919_0, i_13_85_2940_0, i_13_85_2941_0, i_13_85_3021_0,
    i_13_85_3022_0, i_13_85_3039_0, i_13_85_3127_0, i_13_85_3273_0,
    i_13_85_3291_0, i_13_85_3307_0, i_13_85_3345_0, i_13_85_3399_0,
    i_13_85_3418_0, i_13_85_3427_0, i_13_85_3453_0, i_13_85_3454_0,
    i_13_85_3526_0, i_13_85_3534_0, i_13_85_3729_0, i_13_85_3730_0,
    i_13_85_3780_0, i_13_85_3788_0, i_13_85_3874_0, i_13_85_3927_0,
    i_13_85_3967_0, i_13_85_3990_0, i_13_85_4036_0, i_13_85_4065_0,
    i_13_85_4092_0, i_13_85_4189_0, i_13_85_4273_0, i_13_85_4297_0,
    i_13_85_4318_0, i_13_85_4341_0, i_13_85_4525_0, i_13_85_4560_0,
    i_13_85_4561_0, i_13_85_4567_0, i_13_85_4594_0, i_13_85_4603_0,
    o_13_85_0_0  );
  input  i_13_85_67_0, i_13_85_282_0, i_13_85_285_0, i_13_85_384_0,
    i_13_85_385_0, i_13_85_448_0, i_13_85_456_0, i_13_85_625_0,
    i_13_85_669_0, i_13_85_745_0, i_13_85_796_0, i_13_85_816_0,
    i_13_85_852_0, i_13_85_865_0, i_13_85_889_0, i_13_85_948_0,
    i_13_85_1068_0, i_13_85_1101_0, i_13_85_1120_0, i_13_85_1259_0,
    i_13_85_1272_0, i_13_85_1273_0, i_13_85_1302_0, i_13_85_1303_0,
    i_13_85_1312_0, i_13_85_1390_0, i_13_85_1402_0, i_13_85_1484_0,
    i_13_85_1507_0, i_13_85_1573_0, i_13_85_1632_0, i_13_85_1642_0,
    i_13_85_1768_0, i_13_85_1777_0, i_13_85_1794_0, i_13_85_1795_0,
    i_13_85_1851_0, i_13_85_1933_0, i_13_85_1995_0, i_13_85_1996_0,
    i_13_85_2001_0, i_13_85_2014_0, i_13_85_2122_0, i_13_85_2211_0,
    i_13_85_2256_0, i_13_85_2266_0, i_13_85_2380_0, i_13_85_2427_0,
    i_13_85_2433_0, i_13_85_2434_0, i_13_85_2461_0, i_13_85_2463_0,
    i_13_85_2464_0, i_13_85_2470_0, i_13_85_2541_0, i_13_85_2754_0,
    i_13_85_2796_0, i_13_85_2884_0, i_13_85_2905_0, i_13_85_2916_0,
    i_13_85_2919_0, i_13_85_2940_0, i_13_85_2941_0, i_13_85_3021_0,
    i_13_85_3022_0, i_13_85_3039_0, i_13_85_3127_0, i_13_85_3273_0,
    i_13_85_3291_0, i_13_85_3307_0, i_13_85_3345_0, i_13_85_3399_0,
    i_13_85_3418_0, i_13_85_3427_0, i_13_85_3453_0, i_13_85_3454_0,
    i_13_85_3526_0, i_13_85_3534_0, i_13_85_3729_0, i_13_85_3730_0,
    i_13_85_3780_0, i_13_85_3788_0, i_13_85_3874_0, i_13_85_3927_0,
    i_13_85_3967_0, i_13_85_3990_0, i_13_85_4036_0, i_13_85_4065_0,
    i_13_85_4092_0, i_13_85_4189_0, i_13_85_4273_0, i_13_85_4297_0,
    i_13_85_4318_0, i_13_85_4341_0, i_13_85_4525_0, i_13_85_4560_0,
    i_13_85_4561_0, i_13_85_4567_0, i_13_85_4594_0, i_13_85_4603_0;
  output o_13_85_0_0;
  assign o_13_85_0_0 = ~(~i_13_85_2461_0 | (i_13_85_1642_0 & ~i_13_85_4560_0) | (~i_13_85_384_0 & ~i_13_85_2463_0));
endmodule



// Benchmark "kernel_13_86" written by ABC on Sun Jul 19 10:46:38 2020

module kernel_13_86 ( 
    i_13_86_51_0, i_13_86_52_0, i_13_86_66_0, i_13_86_75_0, i_13_86_76_0,
    i_13_86_110_0, i_13_86_111_0, i_13_86_119_0, i_13_86_123_0,
    i_13_86_182_0, i_13_86_183_0, i_13_86_250_0, i_13_86_277_0,
    i_13_86_451_0, i_13_86_507_0, i_13_86_528_0, i_13_86_554_0,
    i_13_86_559_0, i_13_86_561_0, i_13_86_562_0, i_13_86_563_0,
    i_13_86_605_0, i_13_86_618_0, i_13_86_655_0, i_13_86_679_0,
    i_13_86_697_0, i_13_86_699_0, i_13_86_730_0, i_13_86_942_0,
    i_13_86_1078_0, i_13_86_1081_0, i_13_86_1082_0, i_13_86_1084_0,
    i_13_86_1147_0, i_13_86_1210_0, i_13_86_1213_0, i_13_86_1284_0,
    i_13_86_1495_0, i_13_86_1573_0, i_13_86_1622_0, i_13_86_1645_0,
    i_13_86_1659_0, i_13_86_1660_0, i_13_86_1783_0, i_13_86_1784_0,
    i_13_86_1858_0, i_13_86_1920_0, i_13_86_1938_0, i_13_86_2002_0,
    i_13_86_2023_0, i_13_86_2170_0, i_13_86_2234_0, i_13_86_2320_0,
    i_13_86_2423_0, i_13_86_2436_0, i_13_86_2454_0, i_13_86_2455_0,
    i_13_86_2545_0, i_13_86_2616_0, i_13_86_2715_0, i_13_86_2752_0,
    i_13_86_2886_0, i_13_86_2887_0, i_13_86_2958_0, i_13_86_2959_0,
    i_13_86_3035_0, i_13_86_3062_0, i_13_86_3112_0, i_13_86_3129_0,
    i_13_86_3207_0, i_13_86_3214_0, i_13_86_3291_0, i_13_86_3372_0,
    i_13_86_3373_0, i_13_86_3390_0, i_13_86_3405_0, i_13_86_3417_0,
    i_13_86_3418_0, i_13_86_3454_0, i_13_86_3521_0, i_13_86_3526_0,
    i_13_86_3552_0, i_13_86_3571_0, i_13_86_3598_0, i_13_86_3649_0,
    i_13_86_3682_0, i_13_86_3687_0, i_13_86_3700_0, i_13_86_3769_0,
    i_13_86_3903_0, i_13_86_3904_0, i_13_86_3910_0, i_13_86_4332_0,
    i_13_86_4348_0, i_13_86_4349_0, i_13_86_4362_0, i_13_86_4371_0,
    i_13_86_4454_0, i_13_86_4538_0, i_13_86_4603_0,
    o_13_86_0_0  );
  input  i_13_86_51_0, i_13_86_52_0, i_13_86_66_0, i_13_86_75_0,
    i_13_86_76_0, i_13_86_110_0, i_13_86_111_0, i_13_86_119_0,
    i_13_86_123_0, i_13_86_182_0, i_13_86_183_0, i_13_86_250_0,
    i_13_86_277_0, i_13_86_451_0, i_13_86_507_0, i_13_86_528_0,
    i_13_86_554_0, i_13_86_559_0, i_13_86_561_0, i_13_86_562_0,
    i_13_86_563_0, i_13_86_605_0, i_13_86_618_0, i_13_86_655_0,
    i_13_86_679_0, i_13_86_697_0, i_13_86_699_0, i_13_86_730_0,
    i_13_86_942_0, i_13_86_1078_0, i_13_86_1081_0, i_13_86_1082_0,
    i_13_86_1084_0, i_13_86_1147_0, i_13_86_1210_0, i_13_86_1213_0,
    i_13_86_1284_0, i_13_86_1495_0, i_13_86_1573_0, i_13_86_1622_0,
    i_13_86_1645_0, i_13_86_1659_0, i_13_86_1660_0, i_13_86_1783_0,
    i_13_86_1784_0, i_13_86_1858_0, i_13_86_1920_0, i_13_86_1938_0,
    i_13_86_2002_0, i_13_86_2023_0, i_13_86_2170_0, i_13_86_2234_0,
    i_13_86_2320_0, i_13_86_2423_0, i_13_86_2436_0, i_13_86_2454_0,
    i_13_86_2455_0, i_13_86_2545_0, i_13_86_2616_0, i_13_86_2715_0,
    i_13_86_2752_0, i_13_86_2886_0, i_13_86_2887_0, i_13_86_2958_0,
    i_13_86_2959_0, i_13_86_3035_0, i_13_86_3062_0, i_13_86_3112_0,
    i_13_86_3129_0, i_13_86_3207_0, i_13_86_3214_0, i_13_86_3291_0,
    i_13_86_3372_0, i_13_86_3373_0, i_13_86_3390_0, i_13_86_3405_0,
    i_13_86_3417_0, i_13_86_3418_0, i_13_86_3454_0, i_13_86_3521_0,
    i_13_86_3526_0, i_13_86_3552_0, i_13_86_3571_0, i_13_86_3598_0,
    i_13_86_3649_0, i_13_86_3682_0, i_13_86_3687_0, i_13_86_3700_0,
    i_13_86_3769_0, i_13_86_3903_0, i_13_86_3904_0, i_13_86_3910_0,
    i_13_86_4332_0, i_13_86_4348_0, i_13_86_4349_0, i_13_86_4362_0,
    i_13_86_4371_0, i_13_86_4454_0, i_13_86_4538_0, i_13_86_4603_0;
  output o_13_86_0_0;
  assign o_13_86_0_0 = ~((~i_13_86_4362_0 & ~i_13_86_4454_0) | (~i_13_86_1084_0 & ~i_13_86_4371_0));
endmodule



// Benchmark "kernel_13_87" written by ABC on Sun Jul 19 10:46:38 2020

module kernel_13_87 ( 
    i_13_87_51_0, i_13_87_52_0, i_13_87_62_0, i_13_87_79_0, i_13_87_105_0,
    i_13_87_114_0, i_13_87_139_0, i_13_87_143_0, i_13_87_169_0,
    i_13_87_229_0, i_13_87_268_0, i_13_87_269_0, i_13_87_281_0,
    i_13_87_285_0, i_13_87_339_0, i_13_87_340_0, i_13_87_462_0,
    i_13_87_573_0, i_13_87_574_0, i_13_87_610_0, i_13_87_679_0,
    i_13_87_690_0, i_13_87_759_0, i_13_87_813_0, i_13_87_816_0,
    i_13_87_817_0, i_13_87_821_0, i_13_87_984_0, i_13_87_985_0,
    i_13_87_1142_0, i_13_87_1147_0, i_13_87_1274_0, i_13_87_1326_0,
    i_13_87_1476_0, i_13_87_1492_0, i_13_87_1599_0, i_13_87_1626_0,
    i_13_87_1749_0, i_13_87_1780_0, i_13_87_1807_0, i_13_87_1851_0,
    i_13_87_1852_0, i_13_87_1911_0, i_13_87_1950_0, i_13_87_2055_0,
    i_13_87_2058_0, i_13_87_2059_0, i_13_87_2110_0, i_13_87_2119_0,
    i_13_87_2139_0, i_13_87_2184_0, i_13_87_2283_0, i_13_87_2284_0,
    i_13_87_2409_0, i_13_87_2410_0, i_13_87_2579_0, i_13_87_2652_0,
    i_13_87_2696_0, i_13_87_2714_0, i_13_87_2752_0, i_13_87_2859_0,
    i_13_87_2879_0, i_13_87_2940_0, i_13_87_3049_0, i_13_87_3144_0,
    i_13_87_3211_0, i_13_87_3266_0, i_13_87_3291_0, i_13_87_3372_0,
    i_13_87_3373_0, i_13_87_3452_0, i_13_87_3480_0, i_13_87_3505_0,
    i_13_87_3535_0, i_13_87_3563_0, i_13_87_3646_0, i_13_87_3732_0,
    i_13_87_3820_0, i_13_87_3912_0, i_13_87_4018_0, i_13_87_4020_0,
    i_13_87_4045_0, i_13_87_4047_0, i_13_87_4062_0, i_13_87_4065_0,
    i_13_87_4066_0, i_13_87_4116_0, i_13_87_4117_0, i_13_87_4234_0,
    i_13_87_4262_0, i_13_87_4263_0, i_13_87_4296_0, i_13_87_4297_0,
    i_13_87_4309_0, i_13_87_4318_0, i_13_87_4380_0, i_13_87_4391_0,
    i_13_87_4453_0, i_13_87_4560_0, i_13_87_4564_0,
    o_13_87_0_0  );
  input  i_13_87_51_0, i_13_87_52_0, i_13_87_62_0, i_13_87_79_0,
    i_13_87_105_0, i_13_87_114_0, i_13_87_139_0, i_13_87_143_0,
    i_13_87_169_0, i_13_87_229_0, i_13_87_268_0, i_13_87_269_0,
    i_13_87_281_0, i_13_87_285_0, i_13_87_339_0, i_13_87_340_0,
    i_13_87_462_0, i_13_87_573_0, i_13_87_574_0, i_13_87_610_0,
    i_13_87_679_0, i_13_87_690_0, i_13_87_759_0, i_13_87_813_0,
    i_13_87_816_0, i_13_87_817_0, i_13_87_821_0, i_13_87_984_0,
    i_13_87_985_0, i_13_87_1142_0, i_13_87_1147_0, i_13_87_1274_0,
    i_13_87_1326_0, i_13_87_1476_0, i_13_87_1492_0, i_13_87_1599_0,
    i_13_87_1626_0, i_13_87_1749_0, i_13_87_1780_0, i_13_87_1807_0,
    i_13_87_1851_0, i_13_87_1852_0, i_13_87_1911_0, i_13_87_1950_0,
    i_13_87_2055_0, i_13_87_2058_0, i_13_87_2059_0, i_13_87_2110_0,
    i_13_87_2119_0, i_13_87_2139_0, i_13_87_2184_0, i_13_87_2283_0,
    i_13_87_2284_0, i_13_87_2409_0, i_13_87_2410_0, i_13_87_2579_0,
    i_13_87_2652_0, i_13_87_2696_0, i_13_87_2714_0, i_13_87_2752_0,
    i_13_87_2859_0, i_13_87_2879_0, i_13_87_2940_0, i_13_87_3049_0,
    i_13_87_3144_0, i_13_87_3211_0, i_13_87_3266_0, i_13_87_3291_0,
    i_13_87_3372_0, i_13_87_3373_0, i_13_87_3452_0, i_13_87_3480_0,
    i_13_87_3505_0, i_13_87_3535_0, i_13_87_3563_0, i_13_87_3646_0,
    i_13_87_3732_0, i_13_87_3820_0, i_13_87_3912_0, i_13_87_4018_0,
    i_13_87_4020_0, i_13_87_4045_0, i_13_87_4047_0, i_13_87_4062_0,
    i_13_87_4065_0, i_13_87_4066_0, i_13_87_4116_0, i_13_87_4117_0,
    i_13_87_4234_0, i_13_87_4262_0, i_13_87_4263_0, i_13_87_4296_0,
    i_13_87_4297_0, i_13_87_4309_0, i_13_87_4318_0, i_13_87_4380_0,
    i_13_87_4391_0, i_13_87_4453_0, i_13_87_4560_0, i_13_87_4564_0;
  output o_13_87_0_0;
  assign o_13_87_0_0 = ~(i_13_87_62_0 | (~i_13_87_679_0 & ~i_13_87_813_0) | (~i_13_87_2283_0 & ~i_13_87_2410_0 & ~i_13_87_4263_0));
endmodule



// Benchmark "kernel_13_88" written by ABC on Sun Jul 19 10:46:39 2020

module kernel_13_88 ( 
    i_13_88_35_0, i_13_88_66_0, i_13_88_130_0, i_13_88_133_0,
    i_13_88_177_0, i_13_88_236_0, i_13_88_253_0, i_13_88_357_0,
    i_13_88_444_0, i_13_88_455_0, i_13_88_465_0, i_13_88_466_0,
    i_13_88_528_0, i_13_88_582_0, i_13_88_606_0, i_13_88_720_0,
    i_13_88_744_0, i_13_88_915_0, i_13_88_1085_0, i_13_88_1276_0,
    i_13_88_1321_0, i_13_88_1329_0, i_13_88_1363_0, i_13_88_1396_0,
    i_13_88_1444_0, i_13_88_1446_0, i_13_88_1492_0, i_13_88_1500_0,
    i_13_88_1501_0, i_13_88_1507_0, i_13_88_1554_0, i_13_88_1555_0,
    i_13_88_1573_0, i_13_88_1604_0, i_13_88_1641_0, i_13_88_1644_0,
    i_13_88_1699_0, i_13_88_1700_0, i_13_88_1802_0, i_13_88_1848_0,
    i_13_88_1849_0, i_13_88_1929_0, i_13_88_2028_0, i_13_88_2032_0,
    i_13_88_2103_0, i_13_88_2143_0, i_13_88_2202_0, i_13_88_2203_0,
    i_13_88_2297_0, i_13_88_2346_0, i_13_88_2424_0, i_13_88_2425_0,
    i_13_88_2427_0, i_13_88_2468_0, i_13_88_2498_0, i_13_88_2499_0,
    i_13_88_2524_0, i_13_88_2559_0, i_13_88_2569_0, i_13_88_2720_0,
    i_13_88_2755_0, i_13_88_2767_0, i_13_88_2796_0, i_13_88_2887_0,
    i_13_88_2938_0, i_13_88_3027_0, i_13_88_3136_0, i_13_88_3232_0,
    i_13_88_3242_0, i_13_88_3243_0, i_13_88_3244_0, i_13_88_3470_0,
    i_13_88_3507_0, i_13_88_3541_0, i_13_88_3548_0, i_13_88_3596_0,
    i_13_88_3597_0, i_13_88_3613_0, i_13_88_3621_0, i_13_88_3633_0,
    i_13_88_3794_0, i_13_88_3840_0, i_13_88_3847_0, i_13_88_3849_0,
    i_13_88_3859_0, i_13_88_3994_0, i_13_88_4061_0, i_13_88_4063_0,
    i_13_88_4092_0, i_13_88_4125_0, i_13_88_4254_0, i_13_88_4265_0,
    i_13_88_4297_0, i_13_88_4315_0, i_13_88_4325_0, i_13_88_4398_0,
    i_13_88_4471_0, i_13_88_4512_0, i_13_88_4557_0, i_13_88_4603_0,
    o_13_88_0_0  );
  input  i_13_88_35_0, i_13_88_66_0, i_13_88_130_0, i_13_88_133_0,
    i_13_88_177_0, i_13_88_236_0, i_13_88_253_0, i_13_88_357_0,
    i_13_88_444_0, i_13_88_455_0, i_13_88_465_0, i_13_88_466_0,
    i_13_88_528_0, i_13_88_582_0, i_13_88_606_0, i_13_88_720_0,
    i_13_88_744_0, i_13_88_915_0, i_13_88_1085_0, i_13_88_1276_0,
    i_13_88_1321_0, i_13_88_1329_0, i_13_88_1363_0, i_13_88_1396_0,
    i_13_88_1444_0, i_13_88_1446_0, i_13_88_1492_0, i_13_88_1500_0,
    i_13_88_1501_0, i_13_88_1507_0, i_13_88_1554_0, i_13_88_1555_0,
    i_13_88_1573_0, i_13_88_1604_0, i_13_88_1641_0, i_13_88_1644_0,
    i_13_88_1699_0, i_13_88_1700_0, i_13_88_1802_0, i_13_88_1848_0,
    i_13_88_1849_0, i_13_88_1929_0, i_13_88_2028_0, i_13_88_2032_0,
    i_13_88_2103_0, i_13_88_2143_0, i_13_88_2202_0, i_13_88_2203_0,
    i_13_88_2297_0, i_13_88_2346_0, i_13_88_2424_0, i_13_88_2425_0,
    i_13_88_2427_0, i_13_88_2468_0, i_13_88_2498_0, i_13_88_2499_0,
    i_13_88_2524_0, i_13_88_2559_0, i_13_88_2569_0, i_13_88_2720_0,
    i_13_88_2755_0, i_13_88_2767_0, i_13_88_2796_0, i_13_88_2887_0,
    i_13_88_2938_0, i_13_88_3027_0, i_13_88_3136_0, i_13_88_3232_0,
    i_13_88_3242_0, i_13_88_3243_0, i_13_88_3244_0, i_13_88_3470_0,
    i_13_88_3507_0, i_13_88_3541_0, i_13_88_3548_0, i_13_88_3596_0,
    i_13_88_3597_0, i_13_88_3613_0, i_13_88_3621_0, i_13_88_3633_0,
    i_13_88_3794_0, i_13_88_3840_0, i_13_88_3847_0, i_13_88_3849_0,
    i_13_88_3859_0, i_13_88_3994_0, i_13_88_4061_0, i_13_88_4063_0,
    i_13_88_4092_0, i_13_88_4125_0, i_13_88_4254_0, i_13_88_4265_0,
    i_13_88_4297_0, i_13_88_4315_0, i_13_88_4325_0, i_13_88_4398_0,
    i_13_88_4471_0, i_13_88_4512_0, i_13_88_4557_0, i_13_88_4603_0;
  output o_13_88_0_0;
  assign o_13_88_0_0 = ~(i_13_88_4325_0 | (~i_13_88_3859_0 & ~i_13_88_4398_0) | (~i_13_88_35_0 & ~i_13_88_1848_0));
endmodule



// Benchmark "kernel_13_89" written by ABC on Sun Jul 19 10:46:40 2020

module kernel_13_89 ( 
    i_13_89_95_0, i_13_89_121_0, i_13_89_139_0, i_13_89_140_0,
    i_13_89_335_0, i_13_89_362_0, i_13_89_370_0, i_13_89_380_0,
    i_13_89_461_0, i_13_89_586_0, i_13_89_587_0, i_13_89_659_0,
    i_13_89_685_0, i_13_89_812_0, i_13_89_856_0, i_13_89_1063_0,
    i_13_89_1064_0, i_13_89_1082_0, i_13_89_1090_0, i_13_89_1189_0,
    i_13_89_1217_0, i_13_89_1252_0, i_13_89_1273_0, i_13_89_1277_0,
    i_13_89_1298_0, i_13_89_1342_0, i_13_89_1343_0, i_13_89_1441_0,
    i_13_89_1468_0, i_13_89_1487_0, i_13_89_1568_0, i_13_89_1598_0,
    i_13_89_1678_0, i_13_89_1712_0, i_13_89_1778_0, i_13_89_1802_0,
    i_13_89_1811_0, i_13_89_1859_0, i_13_89_1928_0, i_13_89_1954_0,
    i_13_89_1958_0, i_13_89_1990_0, i_13_89_1994_0, i_13_89_2003_0,
    i_13_89_2053_0, i_13_89_2056_0, i_13_89_2189_0, i_13_89_2207_0,
    i_13_89_2260_0, i_13_89_2278_0, i_13_89_2279_0, i_13_89_2377_0,
    i_13_89_2404_0, i_13_89_2494_0, i_13_89_2548_0, i_13_89_2611_0,
    i_13_89_2612_0, i_13_89_2615_0, i_13_89_2633_0, i_13_89_2709_0,
    i_13_89_2710_0, i_13_89_2711_0, i_13_89_2746_0, i_13_89_2794_0,
    i_13_89_2855_0, i_13_89_2984_0, i_13_89_3110_0, i_13_89_3125_0,
    i_13_89_3136_0, i_13_89_3206_0, i_13_89_3217_0, i_13_89_3341_0,
    i_13_89_3367_0, i_13_89_3379_0, i_13_89_3385_0, i_13_89_3386_0,
    i_13_89_3407_0, i_13_89_3415_0, i_13_89_3416_0, i_13_89_3461_0,
    i_13_89_3476_0, i_13_89_3478_0, i_13_89_3532_0, i_13_89_3652_0,
    i_13_89_3664_0, i_13_89_3682_0, i_13_89_3703_0, i_13_89_3704_0,
    i_13_89_3818_0, i_13_89_3862_0, i_13_89_4051_0, i_13_89_4052_0,
    i_13_89_4097_0, i_13_89_4231_0, i_13_89_4268_0, i_13_89_4315_0,
    i_13_89_4393_0, i_13_89_4394_0, i_13_89_4405_0, i_13_89_4411_0,
    o_13_89_0_0  );
  input  i_13_89_95_0, i_13_89_121_0, i_13_89_139_0, i_13_89_140_0,
    i_13_89_335_0, i_13_89_362_0, i_13_89_370_0, i_13_89_380_0,
    i_13_89_461_0, i_13_89_586_0, i_13_89_587_0, i_13_89_659_0,
    i_13_89_685_0, i_13_89_812_0, i_13_89_856_0, i_13_89_1063_0,
    i_13_89_1064_0, i_13_89_1082_0, i_13_89_1090_0, i_13_89_1189_0,
    i_13_89_1217_0, i_13_89_1252_0, i_13_89_1273_0, i_13_89_1277_0,
    i_13_89_1298_0, i_13_89_1342_0, i_13_89_1343_0, i_13_89_1441_0,
    i_13_89_1468_0, i_13_89_1487_0, i_13_89_1568_0, i_13_89_1598_0,
    i_13_89_1678_0, i_13_89_1712_0, i_13_89_1778_0, i_13_89_1802_0,
    i_13_89_1811_0, i_13_89_1859_0, i_13_89_1928_0, i_13_89_1954_0,
    i_13_89_1958_0, i_13_89_1990_0, i_13_89_1994_0, i_13_89_2003_0,
    i_13_89_2053_0, i_13_89_2056_0, i_13_89_2189_0, i_13_89_2207_0,
    i_13_89_2260_0, i_13_89_2278_0, i_13_89_2279_0, i_13_89_2377_0,
    i_13_89_2404_0, i_13_89_2494_0, i_13_89_2548_0, i_13_89_2611_0,
    i_13_89_2612_0, i_13_89_2615_0, i_13_89_2633_0, i_13_89_2709_0,
    i_13_89_2710_0, i_13_89_2711_0, i_13_89_2746_0, i_13_89_2794_0,
    i_13_89_2855_0, i_13_89_2984_0, i_13_89_3110_0, i_13_89_3125_0,
    i_13_89_3136_0, i_13_89_3206_0, i_13_89_3217_0, i_13_89_3341_0,
    i_13_89_3367_0, i_13_89_3379_0, i_13_89_3385_0, i_13_89_3386_0,
    i_13_89_3407_0, i_13_89_3415_0, i_13_89_3416_0, i_13_89_3461_0,
    i_13_89_3476_0, i_13_89_3478_0, i_13_89_3532_0, i_13_89_3652_0,
    i_13_89_3664_0, i_13_89_3682_0, i_13_89_3703_0, i_13_89_3704_0,
    i_13_89_3818_0, i_13_89_3862_0, i_13_89_4051_0, i_13_89_4052_0,
    i_13_89_4097_0, i_13_89_4231_0, i_13_89_4268_0, i_13_89_4315_0,
    i_13_89_4393_0, i_13_89_4394_0, i_13_89_4405_0, i_13_89_4411_0;
  output o_13_89_0_0;
  assign o_13_89_0_0 = ~((~i_13_89_4315_0 & ((~i_13_89_2709_0 & ~i_13_89_3386_0) | (~i_13_89_1273_0 & i_13_89_2278_0 & ~i_13_89_4268_0))) | (~i_13_89_4394_0 & ((~i_13_89_380_0 & ~i_13_89_1342_0 & ~i_13_89_2711_0) | (~i_13_89_2056_0 & ~i_13_89_4411_0))) | (~i_13_89_3682_0 & ~i_13_89_4052_0 & ~i_13_89_4411_0));
endmodule



// Benchmark "kernel_13_90" written by ABC on Sun Jul 19 10:46:41 2020

module kernel_13_90 ( 
    i_13_90_40_0, i_13_90_49_0, i_13_90_95_0, i_13_90_96_0, i_13_90_274_0,
    i_13_90_279_0, i_13_90_443_0, i_13_90_446_0, i_13_90_454_0,
    i_13_90_497_0, i_13_90_536_0, i_13_90_562_0, i_13_90_565_0,
    i_13_90_697_0, i_13_90_910_0, i_13_90_931_0, i_13_90_949_0,
    i_13_90_1067_0, i_13_90_1069_0, i_13_90_1214_0, i_13_90_1273_0,
    i_13_90_1391_0, i_13_90_1426_0, i_13_90_1480_0, i_13_90_1499_0,
    i_13_90_1532_0, i_13_90_1624_0, i_13_90_1636_0, i_13_90_1637_0,
    i_13_90_1642_0, i_13_90_1752_0, i_13_90_1783_0, i_13_90_1784_0,
    i_13_90_1840_0, i_13_90_1885_0, i_13_90_1932_0, i_13_90_2137_0,
    i_13_90_2170_0, i_13_90_2174_0, i_13_90_2209_0, i_13_90_2211_0,
    i_13_90_2233_0, i_13_90_2288_0, i_13_90_2434_0, i_13_90_2437_0,
    i_13_90_2438_0, i_13_90_2446_0, i_13_90_2486_0, i_13_90_2544_0,
    i_13_90_2545_0, i_13_90_2576_0, i_13_90_2650_0, i_13_90_2713_0,
    i_13_90_2716_0, i_13_90_2764_0, i_13_90_3020_0, i_13_90_3064_0,
    i_13_90_3091_0, i_13_90_3093_0, i_13_90_3109_0, i_13_90_3110_0,
    i_13_90_3143_0, i_13_90_3145_0, i_13_90_3164_0, i_13_90_3218_0,
    i_13_90_3271_0, i_13_90_3308_0, i_13_90_3371_0, i_13_90_3394_0,
    i_13_90_3424_0, i_13_90_3425_0, i_13_90_3692_0, i_13_90_3721_0,
    i_13_90_3750_0, i_13_90_3766_0, i_13_90_3767_0, i_13_90_3821_0,
    i_13_90_3856_0, i_13_90_3874_0, i_13_90_3875_0, i_13_90_3878_0,
    i_13_90_3905_0, i_13_90_4018_0, i_13_90_4019_0, i_13_90_4066_0,
    i_13_90_4087_0, i_13_90_4090_0, i_13_90_4091_0, i_13_90_4162_0,
    i_13_90_4205_0, i_13_90_4253_0, i_13_90_4271_0, i_13_90_4351_0,
    i_13_90_4352_0, i_13_90_4354_0, i_13_90_4361_0, i_13_90_4526_0,
    i_13_90_4561_0, i_13_90_4562_0, i_13_90_4567_0,
    o_13_90_0_0  );
  input  i_13_90_40_0, i_13_90_49_0, i_13_90_95_0, i_13_90_96_0,
    i_13_90_274_0, i_13_90_279_0, i_13_90_443_0, i_13_90_446_0,
    i_13_90_454_0, i_13_90_497_0, i_13_90_536_0, i_13_90_562_0,
    i_13_90_565_0, i_13_90_697_0, i_13_90_910_0, i_13_90_931_0,
    i_13_90_949_0, i_13_90_1067_0, i_13_90_1069_0, i_13_90_1214_0,
    i_13_90_1273_0, i_13_90_1391_0, i_13_90_1426_0, i_13_90_1480_0,
    i_13_90_1499_0, i_13_90_1532_0, i_13_90_1624_0, i_13_90_1636_0,
    i_13_90_1637_0, i_13_90_1642_0, i_13_90_1752_0, i_13_90_1783_0,
    i_13_90_1784_0, i_13_90_1840_0, i_13_90_1885_0, i_13_90_1932_0,
    i_13_90_2137_0, i_13_90_2170_0, i_13_90_2174_0, i_13_90_2209_0,
    i_13_90_2211_0, i_13_90_2233_0, i_13_90_2288_0, i_13_90_2434_0,
    i_13_90_2437_0, i_13_90_2438_0, i_13_90_2446_0, i_13_90_2486_0,
    i_13_90_2544_0, i_13_90_2545_0, i_13_90_2576_0, i_13_90_2650_0,
    i_13_90_2713_0, i_13_90_2716_0, i_13_90_2764_0, i_13_90_3020_0,
    i_13_90_3064_0, i_13_90_3091_0, i_13_90_3093_0, i_13_90_3109_0,
    i_13_90_3110_0, i_13_90_3143_0, i_13_90_3145_0, i_13_90_3164_0,
    i_13_90_3218_0, i_13_90_3271_0, i_13_90_3308_0, i_13_90_3371_0,
    i_13_90_3394_0, i_13_90_3424_0, i_13_90_3425_0, i_13_90_3692_0,
    i_13_90_3721_0, i_13_90_3750_0, i_13_90_3766_0, i_13_90_3767_0,
    i_13_90_3821_0, i_13_90_3856_0, i_13_90_3874_0, i_13_90_3875_0,
    i_13_90_3878_0, i_13_90_3905_0, i_13_90_4018_0, i_13_90_4019_0,
    i_13_90_4066_0, i_13_90_4087_0, i_13_90_4090_0, i_13_90_4091_0,
    i_13_90_4162_0, i_13_90_4205_0, i_13_90_4253_0, i_13_90_4271_0,
    i_13_90_4351_0, i_13_90_4352_0, i_13_90_4354_0, i_13_90_4361_0,
    i_13_90_4526_0, i_13_90_4561_0, i_13_90_4562_0, i_13_90_4567_0;
  output o_13_90_0_0;
  assign o_13_90_0_0 = ~((~i_13_90_4087_0 & ((~i_13_90_1069_0 & ~i_13_90_3874_0 & ~i_13_90_4271_0) | (i_13_90_1480_0 & ~i_13_90_4567_0))) | (~i_13_90_3164_0 & ~i_13_90_3218_0) | (~i_13_90_562_0 & ~i_13_90_3875_0) | (~i_13_90_2174_0 & ~i_13_90_4090_0));
endmodule



// Benchmark "kernel_13_91" written by ABC on Sun Jul 19 10:46:42 2020

module kernel_13_91 ( 
    i_13_91_51_0, i_13_91_52_0, i_13_91_53_0, i_13_91_94_0, i_13_91_106_0,
    i_13_91_125_0, i_13_91_149_0, i_13_91_166_0, i_13_91_168_0,
    i_13_91_169_0, i_13_91_188_0, i_13_91_241_0, i_13_91_251_0,
    i_13_91_261_0, i_13_91_264_0, i_13_91_340_0, i_13_91_370_0,
    i_13_91_374_0, i_13_91_418_0, i_13_91_459_0, i_13_91_531_0,
    i_13_91_574_0, i_13_91_619_0, i_13_91_620_0, i_13_91_679_0,
    i_13_91_680_0, i_13_91_772_0, i_13_91_842_0, i_13_91_889_0,
    i_13_91_895_0, i_13_91_952_0, i_13_91_976_0, i_13_91_980_0,
    i_13_91_1024_0, i_13_91_1048_0, i_13_91_1078_0, i_13_91_1079_0,
    i_13_91_1092_0, i_13_91_1142_0, i_13_91_1204_0, i_13_91_1255_0,
    i_13_91_1318_0, i_13_91_1465_0, i_13_91_1479_0, i_13_91_1502_0,
    i_13_91_1573_0, i_13_91_1574_0, i_13_91_1589_0, i_13_91_1609_0,
    i_13_91_1636_0, i_13_91_1637_0, i_13_91_1710_0, i_13_91_1749_0,
    i_13_91_1750_0, i_13_91_1751_0, i_13_91_1761_0, i_13_91_1808_0,
    i_13_91_1817_0, i_13_91_2033_0, i_13_91_2050_0, i_13_91_2411_0,
    i_13_91_2447_0, i_13_91_2722_0, i_13_91_2736_0, i_13_91_2752_0,
    i_13_91_2753_0, i_13_91_2788_0, i_13_91_2941_0, i_13_91_2942_0,
    i_13_91_2959_0, i_13_91_3220_0, i_13_91_3221_0, i_13_91_3373_0,
    i_13_91_3374_0, i_13_91_3418_0, i_13_91_3419_0, i_13_91_3423_0,
    i_13_91_3452_0, i_13_91_3550_0, i_13_91_3554_0, i_13_91_3559_0,
    i_13_91_3652_0, i_13_91_3653_0, i_13_91_3688_0, i_13_91_3719_0,
    i_13_91_3847_0, i_13_91_3965_0, i_13_91_3991_0, i_13_91_4000_0,
    i_13_91_4009_0, i_13_91_4021_0, i_13_91_4048_0, i_13_91_4066_0,
    i_13_91_4094_0, i_13_91_4318_0, i_13_91_4319_0, i_13_91_4364_0,
    i_13_91_4382_0, i_13_91_4391_0, i_13_91_4525_0,
    o_13_91_0_0  );
  input  i_13_91_51_0, i_13_91_52_0, i_13_91_53_0, i_13_91_94_0,
    i_13_91_106_0, i_13_91_125_0, i_13_91_149_0, i_13_91_166_0,
    i_13_91_168_0, i_13_91_169_0, i_13_91_188_0, i_13_91_241_0,
    i_13_91_251_0, i_13_91_261_0, i_13_91_264_0, i_13_91_340_0,
    i_13_91_370_0, i_13_91_374_0, i_13_91_418_0, i_13_91_459_0,
    i_13_91_531_0, i_13_91_574_0, i_13_91_619_0, i_13_91_620_0,
    i_13_91_679_0, i_13_91_680_0, i_13_91_772_0, i_13_91_842_0,
    i_13_91_889_0, i_13_91_895_0, i_13_91_952_0, i_13_91_976_0,
    i_13_91_980_0, i_13_91_1024_0, i_13_91_1048_0, i_13_91_1078_0,
    i_13_91_1079_0, i_13_91_1092_0, i_13_91_1142_0, i_13_91_1204_0,
    i_13_91_1255_0, i_13_91_1318_0, i_13_91_1465_0, i_13_91_1479_0,
    i_13_91_1502_0, i_13_91_1573_0, i_13_91_1574_0, i_13_91_1589_0,
    i_13_91_1609_0, i_13_91_1636_0, i_13_91_1637_0, i_13_91_1710_0,
    i_13_91_1749_0, i_13_91_1750_0, i_13_91_1751_0, i_13_91_1761_0,
    i_13_91_1808_0, i_13_91_1817_0, i_13_91_2033_0, i_13_91_2050_0,
    i_13_91_2411_0, i_13_91_2447_0, i_13_91_2722_0, i_13_91_2736_0,
    i_13_91_2752_0, i_13_91_2753_0, i_13_91_2788_0, i_13_91_2941_0,
    i_13_91_2942_0, i_13_91_2959_0, i_13_91_3220_0, i_13_91_3221_0,
    i_13_91_3373_0, i_13_91_3374_0, i_13_91_3418_0, i_13_91_3419_0,
    i_13_91_3423_0, i_13_91_3452_0, i_13_91_3550_0, i_13_91_3554_0,
    i_13_91_3559_0, i_13_91_3652_0, i_13_91_3653_0, i_13_91_3688_0,
    i_13_91_3719_0, i_13_91_3847_0, i_13_91_3965_0, i_13_91_3991_0,
    i_13_91_4000_0, i_13_91_4009_0, i_13_91_4021_0, i_13_91_4048_0,
    i_13_91_4066_0, i_13_91_4094_0, i_13_91_4318_0, i_13_91_4319_0,
    i_13_91_4364_0, i_13_91_4382_0, i_13_91_4391_0, i_13_91_4525_0;
  output o_13_91_0_0;
  assign o_13_91_0_0 = ~((~i_13_91_1609_0 & ((~i_13_91_1808_0 & ~i_13_91_4048_0) | (~i_13_91_52_0 & ~i_13_91_3221_0 & ~i_13_91_4318_0))) | (~i_13_91_2942_0 & ((i_13_91_418_0 & ~i_13_91_619_0 & ~i_13_91_895_0) | (~i_13_91_340_0 & ~i_13_91_1078_0))) | (~i_13_91_1574_0 & i_13_91_3652_0 & ~i_13_91_3991_0));
endmodule



// Benchmark "kernel_13_92" written by ABC on Sun Jul 19 10:46:43 2020

module kernel_13_92 ( 
    i_13_92_31_0, i_13_92_45_0, i_13_92_49_0, i_13_92_139_0, i_13_92_160_0,
    i_13_92_175_0, i_13_92_214_0, i_13_92_514_0, i_13_92_550_0,
    i_13_92_617_0, i_13_92_648_0, i_13_92_654_0, i_13_92_656_0,
    i_13_92_659_0, i_13_92_679_0, i_13_92_683_0, i_13_92_823_0,
    i_13_92_847_0, i_13_92_850_0, i_13_92_981_0, i_13_92_984_0,
    i_13_92_985_0, i_13_92_1115_0, i_13_92_1148_0, i_13_92_1326_0,
    i_13_92_1327_0, i_13_92_1331_0, i_13_92_1456_0, i_13_92_1516_0,
    i_13_92_1517_0, i_13_92_1519_0, i_13_92_1573_0, i_13_92_1660_0,
    i_13_92_1749_0, i_13_92_1807_0, i_13_92_1885_0, i_13_92_2021_0,
    i_13_92_2024_0, i_13_92_2059_0, i_13_92_2091_0, i_13_92_2097_0,
    i_13_92_2107_0, i_13_92_2185_0, i_13_92_2195_0, i_13_92_2230_0,
    i_13_92_2277_0, i_13_92_2469_0, i_13_92_2470_0, i_13_92_2473_0,
    i_13_92_2474_0, i_13_92_2519_0, i_13_92_2556_0, i_13_92_2642_0,
    i_13_92_2691_0, i_13_92_2699_0, i_13_92_2722_0, i_13_92_2749_0,
    i_13_92_2766_0, i_13_92_2889_0, i_13_92_3009_0, i_13_92_3031_0,
    i_13_92_3032_0, i_13_92_3037_0, i_13_92_3077_0, i_13_92_3112_0,
    i_13_92_3113_0, i_13_92_3138_0, i_13_92_3274_0, i_13_92_3378_0,
    i_13_92_3388_0, i_13_92_3474_0, i_13_92_3483_0, i_13_92_3522_0,
    i_13_92_3547_0, i_13_92_3558_0, i_13_92_3649_0, i_13_92_3662_0,
    i_13_92_3781_0, i_13_92_3819_0, i_13_92_3820_0, i_13_92_3823_0,
    i_13_92_3861_0, i_13_92_3973_0, i_13_92_3978_0, i_13_92_4055_0,
    i_13_92_4120_0, i_13_92_4123_0, i_13_92_4162_0, i_13_92_4165_0,
    i_13_92_4166_0, i_13_92_4365_0, i_13_92_4366_0, i_13_92_4370_0,
    i_13_92_4396_0, i_13_92_4557_0, i_13_92_4564_0, i_13_92_4567_0,
    i_13_92_4597_0, i_13_92_4600_0, i_13_92_4603_0,
    o_13_92_0_0  );
  input  i_13_92_31_0, i_13_92_45_0, i_13_92_49_0, i_13_92_139_0,
    i_13_92_160_0, i_13_92_175_0, i_13_92_214_0, i_13_92_514_0,
    i_13_92_550_0, i_13_92_617_0, i_13_92_648_0, i_13_92_654_0,
    i_13_92_656_0, i_13_92_659_0, i_13_92_679_0, i_13_92_683_0,
    i_13_92_823_0, i_13_92_847_0, i_13_92_850_0, i_13_92_981_0,
    i_13_92_984_0, i_13_92_985_0, i_13_92_1115_0, i_13_92_1148_0,
    i_13_92_1326_0, i_13_92_1327_0, i_13_92_1331_0, i_13_92_1456_0,
    i_13_92_1516_0, i_13_92_1517_0, i_13_92_1519_0, i_13_92_1573_0,
    i_13_92_1660_0, i_13_92_1749_0, i_13_92_1807_0, i_13_92_1885_0,
    i_13_92_2021_0, i_13_92_2024_0, i_13_92_2059_0, i_13_92_2091_0,
    i_13_92_2097_0, i_13_92_2107_0, i_13_92_2185_0, i_13_92_2195_0,
    i_13_92_2230_0, i_13_92_2277_0, i_13_92_2469_0, i_13_92_2470_0,
    i_13_92_2473_0, i_13_92_2474_0, i_13_92_2519_0, i_13_92_2556_0,
    i_13_92_2642_0, i_13_92_2691_0, i_13_92_2699_0, i_13_92_2722_0,
    i_13_92_2749_0, i_13_92_2766_0, i_13_92_2889_0, i_13_92_3009_0,
    i_13_92_3031_0, i_13_92_3032_0, i_13_92_3037_0, i_13_92_3077_0,
    i_13_92_3112_0, i_13_92_3113_0, i_13_92_3138_0, i_13_92_3274_0,
    i_13_92_3378_0, i_13_92_3388_0, i_13_92_3474_0, i_13_92_3483_0,
    i_13_92_3522_0, i_13_92_3547_0, i_13_92_3558_0, i_13_92_3649_0,
    i_13_92_3662_0, i_13_92_3781_0, i_13_92_3819_0, i_13_92_3820_0,
    i_13_92_3823_0, i_13_92_3861_0, i_13_92_3973_0, i_13_92_3978_0,
    i_13_92_4055_0, i_13_92_4120_0, i_13_92_4123_0, i_13_92_4162_0,
    i_13_92_4165_0, i_13_92_4166_0, i_13_92_4365_0, i_13_92_4366_0,
    i_13_92_4370_0, i_13_92_4396_0, i_13_92_4557_0, i_13_92_4564_0,
    i_13_92_4567_0, i_13_92_4597_0, i_13_92_4600_0, i_13_92_4603_0;
  output o_13_92_0_0;
  assign o_13_92_0_0 = ~((~i_13_92_3823_0 & ((~i_13_92_985_0 & ~i_13_92_1326_0) | (~i_13_92_45_0 & ~i_13_92_679_0 & ~i_13_92_1327_0 & ~i_13_92_3112_0 & ~i_13_92_3483_0 & ~i_13_92_3978_0 & ~i_13_92_4370_0))) | (i_13_92_3037_0 & ~i_13_92_3522_0 & ~i_13_92_4162_0) | (~i_13_92_1331_0 & ~i_13_92_1749_0 & ~i_13_92_2107_0 & ~i_13_92_2766_0 & ~i_13_92_3820_0 & ~i_13_92_4165_0 & ~i_13_92_4166_0 & ~i_13_92_4366_0));
endmodule



// Benchmark "kernel_13_93" written by ABC on Sun Jul 19 10:46:43 2020

module kernel_13_93 ( 
    i_13_93_78_0, i_13_93_92_0, i_13_93_157_0, i_13_93_166_0,
    i_13_93_176_0, i_13_93_317_0, i_13_93_382_0, i_13_93_383_0,
    i_13_93_449_0, i_13_93_536_0, i_13_93_551_0, i_13_93_605_0,
    i_13_93_644_0, i_13_93_652_0, i_13_93_653_0, i_13_93_659_0,
    i_13_93_668_0, i_13_93_676_0, i_13_93_679_0, i_13_93_683_0,
    i_13_93_689_0, i_13_93_699_0, i_13_93_701_0, i_13_93_841_0,
    i_13_93_842_0, i_13_93_910_0, i_13_93_1106_0, i_13_93_1120_0,
    i_13_93_1121_0, i_13_93_1145_0, i_13_93_1207_0, i_13_93_1208_0,
    i_13_93_1310_0, i_13_93_1330_0, i_13_93_1423_0, i_13_93_1507_0,
    i_13_93_1516_0, i_13_93_1517_0, i_13_93_1570_0, i_13_93_1571_0,
    i_13_93_1664_0, i_13_93_1733_0, i_13_93_1742_0, i_13_93_1749_0,
    i_13_93_1924_0, i_13_93_1925_0, i_13_93_1937_0, i_13_93_2021_0,
    i_13_93_2054_0, i_13_93_2092_0, i_13_93_2208_0, i_13_93_2209_0,
    i_13_93_2318_0, i_13_93_2398_0, i_13_93_2468_0, i_13_93_2549_0,
    i_13_93_2552_0, i_13_93_2567_0, i_13_93_2582_0, i_13_93_2693_0,
    i_13_93_2699_0, i_13_93_3044_0, i_13_93_3077_0, i_13_93_3089_0,
    i_13_93_3101_0, i_13_93_3214_0, i_13_93_3217_0, i_13_93_3269_0,
    i_13_93_3532_0, i_13_93_3536_0, i_13_93_3559_0, i_13_93_3568_0,
    i_13_93_3569_0, i_13_93_3730_0, i_13_93_3731_0, i_13_93_3857_0,
    i_13_93_3863_0, i_13_93_3866_0, i_13_93_3874_0, i_13_93_3928_0,
    i_13_93_3991_0, i_13_93_3995_0, i_13_93_4033_0, i_13_93_4187_0,
    i_13_93_4190_0, i_13_93_4276_0, i_13_93_4280_0, i_13_93_4307_0,
    i_13_93_4335_0, i_13_93_4364_0, i_13_93_4435_0, i_13_93_4531_0,
    i_13_93_4565_0, i_13_93_4568_0, i_13_93_4585_0, i_13_93_4591_0,
    i_13_93_4592_0, i_13_93_4595_0, i_13_93_4600_0, i_13_93_4601_0,
    o_13_93_0_0  );
  input  i_13_93_78_0, i_13_93_92_0, i_13_93_157_0, i_13_93_166_0,
    i_13_93_176_0, i_13_93_317_0, i_13_93_382_0, i_13_93_383_0,
    i_13_93_449_0, i_13_93_536_0, i_13_93_551_0, i_13_93_605_0,
    i_13_93_644_0, i_13_93_652_0, i_13_93_653_0, i_13_93_659_0,
    i_13_93_668_0, i_13_93_676_0, i_13_93_679_0, i_13_93_683_0,
    i_13_93_689_0, i_13_93_699_0, i_13_93_701_0, i_13_93_841_0,
    i_13_93_842_0, i_13_93_910_0, i_13_93_1106_0, i_13_93_1120_0,
    i_13_93_1121_0, i_13_93_1145_0, i_13_93_1207_0, i_13_93_1208_0,
    i_13_93_1310_0, i_13_93_1330_0, i_13_93_1423_0, i_13_93_1507_0,
    i_13_93_1516_0, i_13_93_1517_0, i_13_93_1570_0, i_13_93_1571_0,
    i_13_93_1664_0, i_13_93_1733_0, i_13_93_1742_0, i_13_93_1749_0,
    i_13_93_1924_0, i_13_93_1925_0, i_13_93_1937_0, i_13_93_2021_0,
    i_13_93_2054_0, i_13_93_2092_0, i_13_93_2208_0, i_13_93_2209_0,
    i_13_93_2318_0, i_13_93_2398_0, i_13_93_2468_0, i_13_93_2549_0,
    i_13_93_2552_0, i_13_93_2567_0, i_13_93_2582_0, i_13_93_2693_0,
    i_13_93_2699_0, i_13_93_3044_0, i_13_93_3077_0, i_13_93_3089_0,
    i_13_93_3101_0, i_13_93_3214_0, i_13_93_3217_0, i_13_93_3269_0,
    i_13_93_3532_0, i_13_93_3536_0, i_13_93_3559_0, i_13_93_3568_0,
    i_13_93_3569_0, i_13_93_3730_0, i_13_93_3731_0, i_13_93_3857_0,
    i_13_93_3863_0, i_13_93_3866_0, i_13_93_3874_0, i_13_93_3928_0,
    i_13_93_3991_0, i_13_93_3995_0, i_13_93_4033_0, i_13_93_4187_0,
    i_13_93_4190_0, i_13_93_4276_0, i_13_93_4280_0, i_13_93_4307_0,
    i_13_93_4335_0, i_13_93_4364_0, i_13_93_4435_0, i_13_93_4531_0,
    i_13_93_4565_0, i_13_93_4568_0, i_13_93_4585_0, i_13_93_4591_0,
    i_13_93_4592_0, i_13_93_4595_0, i_13_93_4600_0, i_13_93_4601_0;
  output o_13_93_0_0;
  assign o_13_93_0_0 = ~((~i_13_93_4033_0 & ~i_13_93_4190_0) | (~i_13_93_2021_0 & ~i_13_93_2054_0 & ~i_13_93_4565_0) | (i_13_93_3532_0 & ~i_13_93_3928_0 & ~i_13_93_4435_0) | (~i_13_93_652_0 & ~i_13_93_683_0 & ~i_13_93_4187_0) | (~i_13_93_679_0 & ~i_13_93_3568_0 & ~i_13_93_3863_0));
endmodule



// Benchmark "kernel_13_94" written by ABC on Sun Jul 19 10:46:44 2020

module kernel_13_94 ( 
    i_13_94_80_0, i_13_94_176_0, i_13_94_263_0, i_13_94_280_0,
    i_13_94_310_0, i_13_94_311_0, i_13_94_316_0, i_13_94_317_0,
    i_13_94_320_0, i_13_94_338_0, i_13_94_355_0, i_13_94_425_0,
    i_13_94_454_0, i_13_94_490_0, i_13_94_550_0, i_13_94_569_0,
    i_13_94_640_0, i_13_94_641_0, i_13_94_644_0, i_13_94_655_0,
    i_13_94_670_0, i_13_94_671_0, i_13_94_685_0, i_13_94_686_0,
    i_13_94_688_0, i_13_94_689_0, i_13_94_820_0, i_13_94_841_0,
    i_13_94_848_0, i_13_94_949_0, i_13_94_1072_0, i_13_94_1120_0,
    i_13_94_1121_0, i_13_94_1123_0, i_13_94_1136_0, i_13_94_1228_0,
    i_13_94_1273_0, i_13_94_1274_0, i_13_94_1276_0, i_13_94_1328_0,
    i_13_94_1361_0, i_13_94_1598_0, i_13_94_1661_0, i_13_94_1739_0,
    i_13_94_1786_0, i_13_94_1940_0, i_13_94_2027_0, i_13_94_2053_0,
    i_13_94_2054_0, i_13_94_2057_0, i_13_94_2173_0, i_13_94_2264_0,
    i_13_94_2345_0, i_13_94_2377_0, i_13_94_2398_0, i_13_94_2405_0,
    i_13_94_2453_0, i_13_94_2462_0, i_13_94_2507_0, i_13_94_2548_0,
    i_13_94_2549_0, i_13_94_2570_0, i_13_94_2579_0, i_13_94_2599_0,
    i_13_94_2651_0, i_13_94_2677_0, i_13_94_2693_0, i_13_94_2695_0,
    i_13_94_2696_0, i_13_94_2699_0, i_13_94_2747_0, i_13_94_3004_0,
    i_13_94_3008_0, i_13_94_3217_0, i_13_94_3340_0, i_13_94_3479_0,
    i_13_94_3538_0, i_13_94_3592_0, i_13_94_3721_0, i_13_94_3782_0,
    i_13_94_3862_0, i_13_94_3875_0, i_13_94_3893_0, i_13_94_3931_0,
    i_13_94_3982_0, i_13_94_3991_0, i_13_94_3992_0, i_13_94_3994_0,
    i_13_94_4019_0, i_13_94_4033_0, i_13_94_4186_0, i_13_94_4258_0,
    i_13_94_4259_0, i_13_94_4262_0, i_13_94_4375_0, i_13_94_4540_0,
    i_13_94_4565_0, i_13_94_4592_0, i_13_94_4595_0, i_13_94_4601_0,
    o_13_94_0_0  );
  input  i_13_94_80_0, i_13_94_176_0, i_13_94_263_0, i_13_94_280_0,
    i_13_94_310_0, i_13_94_311_0, i_13_94_316_0, i_13_94_317_0,
    i_13_94_320_0, i_13_94_338_0, i_13_94_355_0, i_13_94_425_0,
    i_13_94_454_0, i_13_94_490_0, i_13_94_550_0, i_13_94_569_0,
    i_13_94_640_0, i_13_94_641_0, i_13_94_644_0, i_13_94_655_0,
    i_13_94_670_0, i_13_94_671_0, i_13_94_685_0, i_13_94_686_0,
    i_13_94_688_0, i_13_94_689_0, i_13_94_820_0, i_13_94_841_0,
    i_13_94_848_0, i_13_94_949_0, i_13_94_1072_0, i_13_94_1120_0,
    i_13_94_1121_0, i_13_94_1123_0, i_13_94_1136_0, i_13_94_1228_0,
    i_13_94_1273_0, i_13_94_1274_0, i_13_94_1276_0, i_13_94_1328_0,
    i_13_94_1361_0, i_13_94_1598_0, i_13_94_1661_0, i_13_94_1739_0,
    i_13_94_1786_0, i_13_94_1940_0, i_13_94_2027_0, i_13_94_2053_0,
    i_13_94_2054_0, i_13_94_2057_0, i_13_94_2173_0, i_13_94_2264_0,
    i_13_94_2345_0, i_13_94_2377_0, i_13_94_2398_0, i_13_94_2405_0,
    i_13_94_2453_0, i_13_94_2462_0, i_13_94_2507_0, i_13_94_2548_0,
    i_13_94_2549_0, i_13_94_2570_0, i_13_94_2579_0, i_13_94_2599_0,
    i_13_94_2651_0, i_13_94_2677_0, i_13_94_2693_0, i_13_94_2695_0,
    i_13_94_2696_0, i_13_94_2699_0, i_13_94_2747_0, i_13_94_3004_0,
    i_13_94_3008_0, i_13_94_3217_0, i_13_94_3340_0, i_13_94_3479_0,
    i_13_94_3538_0, i_13_94_3592_0, i_13_94_3721_0, i_13_94_3782_0,
    i_13_94_3862_0, i_13_94_3875_0, i_13_94_3893_0, i_13_94_3931_0,
    i_13_94_3982_0, i_13_94_3991_0, i_13_94_3992_0, i_13_94_3994_0,
    i_13_94_4019_0, i_13_94_4033_0, i_13_94_4186_0, i_13_94_4258_0,
    i_13_94_4259_0, i_13_94_4262_0, i_13_94_4375_0, i_13_94_4540_0,
    i_13_94_4565_0, i_13_94_4592_0, i_13_94_4595_0, i_13_94_4601_0;
  output o_13_94_0_0;
  assign o_13_94_0_0 = ~((~i_13_94_1121_0 & ~i_13_94_2696_0) | (i_13_94_355_0 & ~i_13_94_2057_0) | (~i_13_94_3994_0 & ~i_13_94_4033_0 & ~i_13_94_4258_0) | (~i_13_94_2377_0 & ~i_13_94_3008_0 & ~i_13_94_3893_0) | (~i_13_94_1136_0 & ~i_13_94_1228_0 & ~i_13_94_1276_0));
endmodule



// Benchmark "kernel_13_95" written by ABC on Sun Jul 19 10:46:45 2020

module kernel_13_95 ( 
    i_13_95_48_0, i_13_95_53_0, i_13_95_93_0, i_13_95_188_0, i_13_95_316_0,
    i_13_95_351_0, i_13_95_444_0, i_13_95_454_0, i_13_95_549_0,
    i_13_95_550_0, i_13_95_612_0, i_13_95_620_0, i_13_95_640_0,
    i_13_95_643_0, i_13_95_651_0, i_13_95_652_0, i_13_95_667_0,
    i_13_95_675_0, i_13_95_676_0, i_13_95_692_0, i_13_95_742_0,
    i_13_95_839_0, i_13_95_844_0, i_13_95_981_0, i_13_95_982_0,
    i_13_95_985_0, i_13_95_1117_0, i_13_95_1179_0, i_13_95_1181_0,
    i_13_95_1210_0, i_13_95_1498_0, i_13_95_1513_0, i_13_95_1515_0,
    i_13_95_1516_0, i_13_95_1519_0, i_13_95_1574_0, i_13_95_1641_0,
    i_13_95_1747_0, i_13_95_1792_0, i_13_95_1808_0, i_13_95_1810_0,
    i_13_95_1852_0, i_13_95_1853_0, i_13_95_1912_0, i_13_95_2003_0,
    i_13_95_2017_0, i_13_95_2050_0, i_13_95_2060_0, i_13_95_2169_0,
    i_13_95_2170_0, i_13_95_2243_0, i_13_95_2278_0, i_13_95_2348_0,
    i_13_95_2467_0, i_13_95_2511_0, i_13_95_2614_0, i_13_95_2674_0,
    i_13_95_2857_0, i_13_95_2935_0, i_13_95_2980_0, i_13_95_3208_0,
    i_13_95_3212_0, i_13_95_3214_0, i_13_95_3367_0, i_13_95_3369_0,
    i_13_95_3374_0, i_13_95_3401_0, i_13_95_3413_0, i_13_95_3416_0,
    i_13_95_3428_0, i_13_95_3491_0, i_13_95_3532_0, i_13_95_3541_0,
    i_13_95_3550_0, i_13_95_3554_0, i_13_95_3592_0, i_13_95_3645_0,
    i_13_95_3727_0, i_13_95_3730_0, i_13_95_3736_0, i_13_95_3765_0,
    i_13_95_3770_0, i_13_95_3862_0, i_13_95_3866_0, i_13_95_3888_0,
    i_13_95_3889_0, i_13_95_3890_0, i_13_95_3925_0, i_13_95_3987_0,
    i_13_95_3988_0, i_13_95_4049_0, i_13_95_4123_0, i_13_95_4265_0,
    i_13_95_4361_0, i_13_95_4544_0, i_13_95_4564_0, i_13_95_4566_0,
    i_13_95_4591_0, i_13_95_4599_0, i_13_95_4600_0,
    o_13_95_0_0  );
  input  i_13_95_48_0, i_13_95_53_0, i_13_95_93_0, i_13_95_188_0,
    i_13_95_316_0, i_13_95_351_0, i_13_95_444_0, i_13_95_454_0,
    i_13_95_549_0, i_13_95_550_0, i_13_95_612_0, i_13_95_620_0,
    i_13_95_640_0, i_13_95_643_0, i_13_95_651_0, i_13_95_652_0,
    i_13_95_667_0, i_13_95_675_0, i_13_95_676_0, i_13_95_692_0,
    i_13_95_742_0, i_13_95_839_0, i_13_95_844_0, i_13_95_981_0,
    i_13_95_982_0, i_13_95_985_0, i_13_95_1117_0, i_13_95_1179_0,
    i_13_95_1181_0, i_13_95_1210_0, i_13_95_1498_0, i_13_95_1513_0,
    i_13_95_1515_0, i_13_95_1516_0, i_13_95_1519_0, i_13_95_1574_0,
    i_13_95_1641_0, i_13_95_1747_0, i_13_95_1792_0, i_13_95_1808_0,
    i_13_95_1810_0, i_13_95_1852_0, i_13_95_1853_0, i_13_95_1912_0,
    i_13_95_2003_0, i_13_95_2017_0, i_13_95_2050_0, i_13_95_2060_0,
    i_13_95_2169_0, i_13_95_2170_0, i_13_95_2243_0, i_13_95_2278_0,
    i_13_95_2348_0, i_13_95_2467_0, i_13_95_2511_0, i_13_95_2614_0,
    i_13_95_2674_0, i_13_95_2857_0, i_13_95_2935_0, i_13_95_2980_0,
    i_13_95_3208_0, i_13_95_3212_0, i_13_95_3214_0, i_13_95_3367_0,
    i_13_95_3369_0, i_13_95_3374_0, i_13_95_3401_0, i_13_95_3413_0,
    i_13_95_3416_0, i_13_95_3428_0, i_13_95_3491_0, i_13_95_3532_0,
    i_13_95_3541_0, i_13_95_3550_0, i_13_95_3554_0, i_13_95_3592_0,
    i_13_95_3645_0, i_13_95_3727_0, i_13_95_3730_0, i_13_95_3736_0,
    i_13_95_3765_0, i_13_95_3770_0, i_13_95_3862_0, i_13_95_3866_0,
    i_13_95_3888_0, i_13_95_3889_0, i_13_95_3890_0, i_13_95_3925_0,
    i_13_95_3987_0, i_13_95_3988_0, i_13_95_4049_0, i_13_95_4123_0,
    i_13_95_4265_0, i_13_95_4361_0, i_13_95_4544_0, i_13_95_4564_0,
    i_13_95_4566_0, i_13_95_4591_0, i_13_95_4599_0, i_13_95_4600_0;
  output o_13_95_0_0;
  assign o_13_95_0_0 = ~(~i_13_95_3862_0 | (~i_13_95_316_0 & i_13_95_2614_0) | (~i_13_95_676_0 & ~i_13_95_1747_0));
endmodule



// Benchmark "kernel_13_96" written by ABC on Sun Jul 19 10:46:46 2020

module kernel_13_96 ( 
    i_13_96_33_0, i_13_96_40_0, i_13_96_61_0, i_13_96_105_0, i_13_96_142_0,
    i_13_96_184_0, i_13_96_186_0, i_13_96_187_0, i_13_96_231_0,
    i_13_96_237_0, i_13_96_274_0, i_13_96_282_0, i_13_96_310_0,
    i_13_96_313_0, i_13_96_318_0, i_13_96_319_0, i_13_96_445_0,
    i_13_96_453_0, i_13_96_537_0, i_13_96_564_0, i_13_96_573_0,
    i_13_96_574_0, i_13_96_601_0, i_13_96_643_0, i_13_96_645_0,
    i_13_96_646_0, i_13_96_688_0, i_13_96_690_0, i_13_96_691_0,
    i_13_96_700_0, i_13_96_714_0, i_13_96_823_0, i_13_96_897_0,
    i_13_96_898_0, i_13_96_940_0, i_13_96_1069_0, i_13_96_1119_0,
    i_13_96_1123_0, i_13_96_1221_0, i_13_96_1275_0, i_13_96_1276_0,
    i_13_96_1383_0, i_13_96_1498_0, i_13_96_1635_0, i_13_96_1641_0,
    i_13_96_1642_0, i_13_96_1671_0, i_13_96_1716_0, i_13_96_1745_0,
    i_13_96_1852_0, i_13_96_1862_0, i_13_96_2047_0, i_13_96_2103_0,
    i_13_96_2140_0, i_13_96_2239_0, i_13_96_2299_0, i_13_96_2316_0,
    i_13_96_2321_0, i_13_96_2407_0, i_13_96_2509_0, i_13_96_2514_0,
    i_13_96_2635_0, i_13_96_2650_0, i_13_96_2652_0, i_13_96_2653_0,
    i_13_96_2679_0, i_13_96_2698_0, i_13_96_2722_0, i_13_96_2767_0,
    i_13_96_2770_0, i_13_96_2847_0, i_13_96_2848_0, i_13_96_2851_0,
    i_13_96_2984_0, i_13_96_3129_0, i_13_96_3210_0, i_13_96_3274_0,
    i_13_96_3292_0, i_13_96_3387_0, i_13_96_3390_0, i_13_96_3391_0,
    i_13_96_3408_0, i_13_96_3426_0, i_13_96_3460_0, i_13_96_3487_0,
    i_13_96_3606_0, i_13_96_3838_0, i_13_96_3892_0, i_13_96_3921_0,
    i_13_96_3927_0, i_13_96_3930_0, i_13_96_4018_0, i_13_96_4080_0,
    i_13_96_4084_0, i_13_96_4201_0, i_13_96_4344_0, i_13_96_4372_0,
    i_13_96_4570_0, i_13_96_4584_0, i_13_96_4597_0,
    o_13_96_0_0  );
  input  i_13_96_33_0, i_13_96_40_0, i_13_96_61_0, i_13_96_105_0,
    i_13_96_142_0, i_13_96_184_0, i_13_96_186_0, i_13_96_187_0,
    i_13_96_231_0, i_13_96_237_0, i_13_96_274_0, i_13_96_282_0,
    i_13_96_310_0, i_13_96_313_0, i_13_96_318_0, i_13_96_319_0,
    i_13_96_445_0, i_13_96_453_0, i_13_96_537_0, i_13_96_564_0,
    i_13_96_573_0, i_13_96_574_0, i_13_96_601_0, i_13_96_643_0,
    i_13_96_645_0, i_13_96_646_0, i_13_96_688_0, i_13_96_690_0,
    i_13_96_691_0, i_13_96_700_0, i_13_96_714_0, i_13_96_823_0,
    i_13_96_897_0, i_13_96_898_0, i_13_96_940_0, i_13_96_1069_0,
    i_13_96_1119_0, i_13_96_1123_0, i_13_96_1221_0, i_13_96_1275_0,
    i_13_96_1276_0, i_13_96_1383_0, i_13_96_1498_0, i_13_96_1635_0,
    i_13_96_1641_0, i_13_96_1642_0, i_13_96_1671_0, i_13_96_1716_0,
    i_13_96_1745_0, i_13_96_1852_0, i_13_96_1862_0, i_13_96_2047_0,
    i_13_96_2103_0, i_13_96_2140_0, i_13_96_2239_0, i_13_96_2299_0,
    i_13_96_2316_0, i_13_96_2321_0, i_13_96_2407_0, i_13_96_2509_0,
    i_13_96_2514_0, i_13_96_2635_0, i_13_96_2650_0, i_13_96_2652_0,
    i_13_96_2653_0, i_13_96_2679_0, i_13_96_2698_0, i_13_96_2722_0,
    i_13_96_2767_0, i_13_96_2770_0, i_13_96_2847_0, i_13_96_2848_0,
    i_13_96_2851_0, i_13_96_2984_0, i_13_96_3129_0, i_13_96_3210_0,
    i_13_96_3274_0, i_13_96_3292_0, i_13_96_3387_0, i_13_96_3390_0,
    i_13_96_3391_0, i_13_96_3408_0, i_13_96_3426_0, i_13_96_3460_0,
    i_13_96_3487_0, i_13_96_3606_0, i_13_96_3838_0, i_13_96_3892_0,
    i_13_96_3921_0, i_13_96_3927_0, i_13_96_3930_0, i_13_96_4018_0,
    i_13_96_4080_0, i_13_96_4084_0, i_13_96_4201_0, i_13_96_4344_0,
    i_13_96_4372_0, i_13_96_4570_0, i_13_96_4584_0, i_13_96_4597_0;
  output o_13_96_0_0;
  assign o_13_96_0_0 = ~((~i_13_96_897_0 & ((~i_13_96_690_0 & ~i_13_96_1276_0) | (~i_13_96_1716_0 & ~i_13_96_4570_0))) | (~i_13_96_1642_0 & ~i_13_96_3210_0) | (~i_13_96_186_0 & i_13_96_3487_0) | (i_13_96_3892_0 & ~i_13_96_4084_0));
endmodule



// Benchmark "kernel_13_97" written by ABC on Sun Jul 19 10:46:47 2020

module kernel_13_97 ( 
    i_13_97_52_0, i_13_97_103_0, i_13_97_106_0, i_13_97_107_0,
    i_13_97_158_0, i_13_97_166_0, i_13_97_233_0, i_13_97_287_0,
    i_13_97_310_0, i_13_97_337_0, i_13_97_454_0, i_13_97_470_0,
    i_13_97_537_0, i_13_97_553_0, i_13_97_584_0, i_13_97_607_0,
    i_13_97_608_0, i_13_97_646_0, i_13_97_647_0, i_13_97_679_0,
    i_13_97_688_0, i_13_97_691_0, i_13_97_692_0, i_13_97_843_0,
    i_13_97_844_0, i_13_97_1070_0, i_13_97_1086_0, i_13_97_1087_0,
    i_13_97_1106_0, i_13_97_1123_0, i_13_97_1131_0, i_13_97_1300_0,
    i_13_97_1331_0, i_13_97_1519_0, i_13_97_1554_0, i_13_97_1572_0,
    i_13_97_1573_0, i_13_97_1780_0, i_13_97_1804_0, i_13_97_1840_0,
    i_13_97_1915_0, i_13_97_1930_0, i_13_97_2024_0, i_13_97_2059_0,
    i_13_97_2060_0, i_13_97_2172_0, i_13_97_2173_0, i_13_97_2194_0,
    i_13_97_2284_0, i_13_97_2316_0, i_13_97_2380_0, i_13_97_2455_0,
    i_13_97_2624_0, i_13_97_2680_0, i_13_97_2698_0, i_13_97_2715_0,
    i_13_97_2798_0, i_13_97_2852_0, i_13_97_2902_0, i_13_97_2923_0,
    i_13_97_2938_0, i_13_97_3046_0, i_13_97_3066_0, i_13_97_3067_0,
    i_13_97_3103_0, i_13_97_3147_0, i_13_97_3148_0, i_13_97_3209_0,
    i_13_97_3289_0, i_13_97_3346_0, i_13_97_3383_0, i_13_97_3391_0,
    i_13_97_3392_0, i_13_97_3397_0, i_13_97_3446_0, i_13_97_3526_0,
    i_13_97_3530_0, i_13_97_3535_0, i_13_97_3544_0, i_13_97_3687_0,
    i_13_97_3742_0, i_13_97_3748_0, i_13_97_3865_0, i_13_97_3930_0,
    i_13_97_4020_0, i_13_97_4021_0, i_13_97_4048_0, i_13_97_4085_0,
    i_13_97_4119_0, i_13_97_4120_0, i_13_97_4121_0, i_13_97_4214_0,
    i_13_97_4308_0, i_13_97_4417_0, i_13_97_4450_0, i_13_97_4568_0,
    i_13_97_4570_0, i_13_97_4597_0, i_13_97_4598_0, i_13_97_4604_0,
    o_13_97_0_0  );
  input  i_13_97_52_0, i_13_97_103_0, i_13_97_106_0, i_13_97_107_0,
    i_13_97_158_0, i_13_97_166_0, i_13_97_233_0, i_13_97_287_0,
    i_13_97_310_0, i_13_97_337_0, i_13_97_454_0, i_13_97_470_0,
    i_13_97_537_0, i_13_97_553_0, i_13_97_584_0, i_13_97_607_0,
    i_13_97_608_0, i_13_97_646_0, i_13_97_647_0, i_13_97_679_0,
    i_13_97_688_0, i_13_97_691_0, i_13_97_692_0, i_13_97_843_0,
    i_13_97_844_0, i_13_97_1070_0, i_13_97_1086_0, i_13_97_1087_0,
    i_13_97_1106_0, i_13_97_1123_0, i_13_97_1131_0, i_13_97_1300_0,
    i_13_97_1331_0, i_13_97_1519_0, i_13_97_1554_0, i_13_97_1572_0,
    i_13_97_1573_0, i_13_97_1780_0, i_13_97_1804_0, i_13_97_1840_0,
    i_13_97_1915_0, i_13_97_1930_0, i_13_97_2024_0, i_13_97_2059_0,
    i_13_97_2060_0, i_13_97_2172_0, i_13_97_2173_0, i_13_97_2194_0,
    i_13_97_2284_0, i_13_97_2316_0, i_13_97_2380_0, i_13_97_2455_0,
    i_13_97_2624_0, i_13_97_2680_0, i_13_97_2698_0, i_13_97_2715_0,
    i_13_97_2798_0, i_13_97_2852_0, i_13_97_2902_0, i_13_97_2923_0,
    i_13_97_2938_0, i_13_97_3046_0, i_13_97_3066_0, i_13_97_3067_0,
    i_13_97_3103_0, i_13_97_3147_0, i_13_97_3148_0, i_13_97_3209_0,
    i_13_97_3289_0, i_13_97_3346_0, i_13_97_3383_0, i_13_97_3391_0,
    i_13_97_3392_0, i_13_97_3397_0, i_13_97_3446_0, i_13_97_3526_0,
    i_13_97_3530_0, i_13_97_3535_0, i_13_97_3544_0, i_13_97_3687_0,
    i_13_97_3742_0, i_13_97_3748_0, i_13_97_3865_0, i_13_97_3930_0,
    i_13_97_4020_0, i_13_97_4021_0, i_13_97_4048_0, i_13_97_4085_0,
    i_13_97_4119_0, i_13_97_4120_0, i_13_97_4121_0, i_13_97_4214_0,
    i_13_97_4308_0, i_13_97_4417_0, i_13_97_4450_0, i_13_97_4568_0,
    i_13_97_4570_0, i_13_97_4597_0, i_13_97_4598_0, i_13_97_4604_0;
  output o_13_97_0_0;
  assign o_13_97_0_0 = ~((~i_13_97_3147_0 & ((i_13_97_337_0 & ~i_13_97_1070_0) | (~i_13_97_106_0 & ~i_13_97_3067_0))) | (i_13_97_103_0 & ~i_13_97_2059_0 & ~i_13_97_3526_0) | (~i_13_97_1087_0 & i_13_97_3535_0) | (i_13_97_3544_0 & ~i_13_97_3742_0));
endmodule



// Benchmark "kernel_13_98" written by ABC on Sun Jul 19 10:46:47 2020

module kernel_13_98 ( 
    i_13_98_67_0, i_13_98_122_0, i_13_98_162_0, i_13_98_185_0,
    i_13_98_193_0, i_13_98_277_0, i_13_98_333_0, i_13_98_363_0,
    i_13_98_367_0, i_13_98_412_0, i_13_98_444_0, i_13_98_457_0,
    i_13_98_493_0, i_13_98_565_0, i_13_98_571_0, i_13_98_572_0,
    i_13_98_608_0, i_13_98_661_0, i_13_98_715_0, i_13_98_760_0,
    i_13_98_935_0, i_13_98_949_0, i_13_98_952_0, i_13_98_953_0,
    i_13_98_1210_0, i_13_98_1232_0, i_13_98_1267_0, i_13_98_1408_0,
    i_13_98_1443_0, i_13_98_1507_0, i_13_98_1625_0, i_13_98_1627_0,
    i_13_98_1628_0, i_13_98_1634_0, i_13_98_1637_0, i_13_98_1717_0,
    i_13_98_1736_0, i_13_98_1768_0, i_13_98_1771_0, i_13_98_1789_0,
    i_13_98_1790_0, i_13_98_1805_0, i_13_98_1808_0, i_13_98_1832_0,
    i_13_98_1912_0, i_13_98_1921_0, i_13_98_1940_0, i_13_98_2003_0,
    i_13_98_2012_0, i_13_98_2056_0, i_13_98_2123_0, i_13_98_2209_0,
    i_13_98_2240_0, i_13_98_2314_0, i_13_98_2426_0, i_13_98_2437_0,
    i_13_98_2533_0, i_13_98_2534_0, i_13_98_2538_0, i_13_98_2620_0,
    i_13_98_2987_0, i_13_98_3023_0, i_13_98_3032_0, i_13_98_3047_0,
    i_13_98_3104_0, i_13_98_3105_0, i_13_98_3166_0, i_13_98_3167_0,
    i_13_98_3231_0, i_13_98_3253_0, i_13_98_3265_0, i_13_98_3329_0,
    i_13_98_3397_0, i_13_98_3416_0, i_13_98_3420_0, i_13_98_3527_0,
    i_13_98_3550_0, i_13_98_3616_0, i_13_98_3681_0, i_13_98_3703_0,
    i_13_98_3847_0, i_13_98_3870_0, i_13_98_3874_0, i_13_98_3875_0,
    i_13_98_3878_0, i_13_98_3892_0, i_13_98_3982_0, i_13_98_3985_0,
    i_13_98_3986_0, i_13_98_4009_0, i_13_98_4198_0, i_13_98_4248_0,
    i_13_98_4311_0, i_13_98_4325_0, i_13_98_4327_0, i_13_98_4347_0,
    i_13_98_4351_0, i_13_98_4509_0, i_13_98_4514_0, i_13_98_4541_0,
    o_13_98_0_0  );
  input  i_13_98_67_0, i_13_98_122_0, i_13_98_162_0, i_13_98_185_0,
    i_13_98_193_0, i_13_98_277_0, i_13_98_333_0, i_13_98_363_0,
    i_13_98_367_0, i_13_98_412_0, i_13_98_444_0, i_13_98_457_0,
    i_13_98_493_0, i_13_98_565_0, i_13_98_571_0, i_13_98_572_0,
    i_13_98_608_0, i_13_98_661_0, i_13_98_715_0, i_13_98_760_0,
    i_13_98_935_0, i_13_98_949_0, i_13_98_952_0, i_13_98_953_0,
    i_13_98_1210_0, i_13_98_1232_0, i_13_98_1267_0, i_13_98_1408_0,
    i_13_98_1443_0, i_13_98_1507_0, i_13_98_1625_0, i_13_98_1627_0,
    i_13_98_1628_0, i_13_98_1634_0, i_13_98_1637_0, i_13_98_1717_0,
    i_13_98_1736_0, i_13_98_1768_0, i_13_98_1771_0, i_13_98_1789_0,
    i_13_98_1790_0, i_13_98_1805_0, i_13_98_1808_0, i_13_98_1832_0,
    i_13_98_1912_0, i_13_98_1921_0, i_13_98_1940_0, i_13_98_2003_0,
    i_13_98_2012_0, i_13_98_2056_0, i_13_98_2123_0, i_13_98_2209_0,
    i_13_98_2240_0, i_13_98_2314_0, i_13_98_2426_0, i_13_98_2437_0,
    i_13_98_2533_0, i_13_98_2534_0, i_13_98_2538_0, i_13_98_2620_0,
    i_13_98_2987_0, i_13_98_3023_0, i_13_98_3032_0, i_13_98_3047_0,
    i_13_98_3104_0, i_13_98_3105_0, i_13_98_3166_0, i_13_98_3167_0,
    i_13_98_3231_0, i_13_98_3253_0, i_13_98_3265_0, i_13_98_3329_0,
    i_13_98_3397_0, i_13_98_3416_0, i_13_98_3420_0, i_13_98_3527_0,
    i_13_98_3550_0, i_13_98_3616_0, i_13_98_3681_0, i_13_98_3703_0,
    i_13_98_3847_0, i_13_98_3870_0, i_13_98_3874_0, i_13_98_3875_0,
    i_13_98_3878_0, i_13_98_3892_0, i_13_98_3982_0, i_13_98_3985_0,
    i_13_98_3986_0, i_13_98_4009_0, i_13_98_4198_0, i_13_98_4248_0,
    i_13_98_4311_0, i_13_98_4325_0, i_13_98_4327_0, i_13_98_4347_0,
    i_13_98_4351_0, i_13_98_4509_0, i_13_98_4514_0, i_13_98_4541_0;
  output o_13_98_0_0;
  assign o_13_98_0_0 = ~((~i_13_98_2534_0 & ((~i_13_98_1408_0 & ~i_13_98_1627_0 & ~i_13_98_3982_0) | (~i_13_98_1736_0 & ~i_13_98_2437_0 & ~i_13_98_3875_0 & ~i_13_98_4347_0))) | ~i_13_98_193_0 | (~i_13_98_2209_0 & ~i_13_98_3982_0 & ~i_13_98_3986_0) | (~i_13_98_122_0 & ~i_13_98_4009_0) | (~i_13_98_185_0 & i_13_98_3397_0 & ~i_13_98_4514_0));
endmodule



// Benchmark "kernel_13_99" written by ABC on Sun Jul 19 10:46:48 2020

module kernel_13_99 ( 
    i_13_99_31_0, i_13_99_67_0, i_13_99_94_0, i_13_99_229_0, i_13_99_258_0,
    i_13_99_276_0, i_13_99_310_0, i_13_99_311_0, i_13_99_319_0,
    i_13_99_320_0, i_13_99_418_0, i_13_99_425_0, i_13_99_515_0,
    i_13_99_517_0, i_13_99_520_0, i_13_99_628_0, i_13_99_662_0,
    i_13_99_688_0, i_13_99_868_0, i_13_99_915_0, i_13_99_941_0,
    i_13_99_980_0, i_13_99_1021_0, i_13_99_1077_0, i_13_99_1202_0,
    i_13_99_1330_0, i_13_99_1331_0, i_13_99_1424_0, i_13_99_1444_0,
    i_13_99_1596_0, i_13_99_1598_0, i_13_99_1642_0, i_13_99_1663_0,
    i_13_99_1723_0, i_13_99_1734_0, i_13_99_1745_0, i_13_99_1824_0,
    i_13_99_1832_0, i_13_99_2008_0, i_13_99_2027_0, i_13_99_2132_0,
    i_13_99_2272_0, i_13_99_2317_0, i_13_99_2374_0, i_13_99_2450_0,
    i_13_99_2453_0, i_13_99_2497_0, i_13_99_2541_0, i_13_99_2542_0,
    i_13_99_2593_0, i_13_99_2666_0, i_13_99_2677_0, i_13_99_2740_0,
    i_13_99_2743_0, i_13_99_2744_0, i_13_99_2904_0, i_13_99_2915_0,
    i_13_99_2920_0, i_13_99_2968_0, i_13_99_3002_0, i_13_99_3121_0,
    i_13_99_3139_0, i_13_99_3176_0, i_13_99_3245_0, i_13_99_3312_0,
    i_13_99_3316_0, i_13_99_3414_0, i_13_99_3454_0, i_13_99_3455_0,
    i_13_99_3460_0, i_13_99_3463_0, i_13_99_3464_0, i_13_99_3479_0,
    i_13_99_3486_0, i_13_99_3488_0, i_13_99_3523_0, i_13_99_3569_0,
    i_13_99_3570_0, i_13_99_3571_0, i_13_99_3572_0, i_13_99_3577_0,
    i_13_99_3578_0, i_13_99_3593_0, i_13_99_3767_0, i_13_99_3831_0,
    i_13_99_3866_0, i_13_99_3942_0, i_13_99_4054_0, i_13_99_4094_0,
    i_13_99_4153_0, i_13_99_4164_0, i_13_99_4255_0, i_13_99_4256_0,
    i_13_99_4336_0, i_13_99_4352_0, i_13_99_4368_0, i_13_99_4372_0,
    i_13_99_4373_0, i_13_99_4517_0, i_13_99_4557_0,
    o_13_99_0_0  );
  input  i_13_99_31_0, i_13_99_67_0, i_13_99_94_0, i_13_99_229_0,
    i_13_99_258_0, i_13_99_276_0, i_13_99_310_0, i_13_99_311_0,
    i_13_99_319_0, i_13_99_320_0, i_13_99_418_0, i_13_99_425_0,
    i_13_99_515_0, i_13_99_517_0, i_13_99_520_0, i_13_99_628_0,
    i_13_99_662_0, i_13_99_688_0, i_13_99_868_0, i_13_99_915_0,
    i_13_99_941_0, i_13_99_980_0, i_13_99_1021_0, i_13_99_1077_0,
    i_13_99_1202_0, i_13_99_1330_0, i_13_99_1331_0, i_13_99_1424_0,
    i_13_99_1444_0, i_13_99_1596_0, i_13_99_1598_0, i_13_99_1642_0,
    i_13_99_1663_0, i_13_99_1723_0, i_13_99_1734_0, i_13_99_1745_0,
    i_13_99_1824_0, i_13_99_1832_0, i_13_99_2008_0, i_13_99_2027_0,
    i_13_99_2132_0, i_13_99_2272_0, i_13_99_2317_0, i_13_99_2374_0,
    i_13_99_2450_0, i_13_99_2453_0, i_13_99_2497_0, i_13_99_2541_0,
    i_13_99_2542_0, i_13_99_2593_0, i_13_99_2666_0, i_13_99_2677_0,
    i_13_99_2740_0, i_13_99_2743_0, i_13_99_2744_0, i_13_99_2904_0,
    i_13_99_2915_0, i_13_99_2920_0, i_13_99_2968_0, i_13_99_3002_0,
    i_13_99_3121_0, i_13_99_3139_0, i_13_99_3176_0, i_13_99_3245_0,
    i_13_99_3312_0, i_13_99_3316_0, i_13_99_3414_0, i_13_99_3454_0,
    i_13_99_3455_0, i_13_99_3460_0, i_13_99_3463_0, i_13_99_3464_0,
    i_13_99_3479_0, i_13_99_3486_0, i_13_99_3488_0, i_13_99_3523_0,
    i_13_99_3569_0, i_13_99_3570_0, i_13_99_3571_0, i_13_99_3572_0,
    i_13_99_3577_0, i_13_99_3578_0, i_13_99_3593_0, i_13_99_3767_0,
    i_13_99_3831_0, i_13_99_3866_0, i_13_99_3942_0, i_13_99_4054_0,
    i_13_99_4094_0, i_13_99_4153_0, i_13_99_4164_0, i_13_99_4255_0,
    i_13_99_4256_0, i_13_99_4336_0, i_13_99_4352_0, i_13_99_4368_0,
    i_13_99_4372_0, i_13_99_4373_0, i_13_99_4517_0, i_13_99_4557_0;
  output o_13_99_0_0;
  assign o_13_99_0_0 = ~((~i_13_99_3316_0 & (i_13_99_67_0 | (~i_13_99_3488_0 & i_13_99_3593_0))) | (~i_13_99_2542_0 & i_13_99_2677_0 & ~i_13_99_3455_0) | (~i_13_99_276_0 & ~i_13_99_2453_0 & ~i_13_99_3571_0) | (~i_13_99_2740_0 & ~i_13_99_3577_0 & ~i_13_99_3578_0) | (i_13_99_688_0 & i_13_99_1077_0 & ~i_13_99_4372_0));
endmodule



// Benchmark "kernel_13_100" written by ABC on Sun Jul 19 10:46:49 2020

module kernel_13_100 ( 
    i_13_100_48_0, i_13_100_49_0, i_13_100_70_0, i_13_100_163_0,
    i_13_100_175_0, i_13_100_258_0, i_13_100_259_0, i_13_100_266_0,
    i_13_100_285_0, i_13_100_310_0, i_13_100_336_0, i_13_100_373_0,
    i_13_100_448_0, i_13_100_474_0, i_13_100_616_0, i_13_100_625_0,
    i_13_100_669_0, i_13_100_697_0, i_13_100_834_0, i_13_100_930_0,
    i_13_100_933_0, i_13_100_1071_0, i_13_100_1104_0, i_13_100_1105_0,
    i_13_100_1402_0, i_13_100_1648_0, i_13_100_1726_0, i_13_100_1735_0,
    i_13_100_1780_0, i_13_100_1797_0, i_13_100_1798_0, i_13_100_1804_0,
    i_13_100_1816_0, i_13_100_1818_0, i_13_100_1950_0, i_13_100_1995_0,
    i_13_100_1996_0, i_13_100_2004_0, i_13_100_2022_0, i_13_100_2148_0,
    i_13_100_2212_0, i_13_100_2356_0, i_13_100_2407_0, i_13_100_2409_0,
    i_13_100_2472_0, i_13_100_2473_0, i_13_100_2501_0, i_13_100_2617_0,
    i_13_100_2652_0, i_13_100_2673_0, i_13_100_2907_0, i_13_100_2915_0,
    i_13_100_2940_0, i_13_100_2941_0, i_13_100_2987_0, i_13_100_2997_0,
    i_13_100_3000_0, i_13_100_3030_0, i_13_100_3031_0, i_13_100_3127_0,
    i_13_100_3129_0, i_13_100_3130_0, i_13_100_3135_0, i_13_100_3217_0,
    i_13_100_3220_0, i_13_100_3265_0, i_13_100_3291_0, i_13_100_3312_0,
    i_13_100_3315_0, i_13_100_3376_0, i_13_100_3399_0, i_13_100_3417_0,
    i_13_100_3453_0, i_13_100_3639_0, i_13_100_3702_0, i_13_100_3741_0,
    i_13_100_3822_0, i_13_100_3834_0, i_13_100_3892_0, i_13_100_3940_0,
    i_13_100_3994_0, i_13_100_4045_0, i_13_100_4056_0, i_13_100_4057_0,
    i_13_100_4065_0, i_13_100_4083_0, i_13_100_4094_0, i_13_100_4153_0,
    i_13_100_4164_0, i_13_100_4188_0, i_13_100_4234_0, i_13_100_4251_0,
    i_13_100_4269_0, i_13_100_4273_0, i_13_100_4274_0, i_13_100_4324_0,
    i_13_100_4360_0, i_13_100_4526_0, i_13_100_4533_0, i_13_100_4606_0,
    o_13_100_0_0  );
  input  i_13_100_48_0, i_13_100_49_0, i_13_100_70_0, i_13_100_163_0,
    i_13_100_175_0, i_13_100_258_0, i_13_100_259_0, i_13_100_266_0,
    i_13_100_285_0, i_13_100_310_0, i_13_100_336_0, i_13_100_373_0,
    i_13_100_448_0, i_13_100_474_0, i_13_100_616_0, i_13_100_625_0,
    i_13_100_669_0, i_13_100_697_0, i_13_100_834_0, i_13_100_930_0,
    i_13_100_933_0, i_13_100_1071_0, i_13_100_1104_0, i_13_100_1105_0,
    i_13_100_1402_0, i_13_100_1648_0, i_13_100_1726_0, i_13_100_1735_0,
    i_13_100_1780_0, i_13_100_1797_0, i_13_100_1798_0, i_13_100_1804_0,
    i_13_100_1816_0, i_13_100_1818_0, i_13_100_1950_0, i_13_100_1995_0,
    i_13_100_1996_0, i_13_100_2004_0, i_13_100_2022_0, i_13_100_2148_0,
    i_13_100_2212_0, i_13_100_2356_0, i_13_100_2407_0, i_13_100_2409_0,
    i_13_100_2472_0, i_13_100_2473_0, i_13_100_2501_0, i_13_100_2617_0,
    i_13_100_2652_0, i_13_100_2673_0, i_13_100_2907_0, i_13_100_2915_0,
    i_13_100_2940_0, i_13_100_2941_0, i_13_100_2987_0, i_13_100_2997_0,
    i_13_100_3000_0, i_13_100_3030_0, i_13_100_3031_0, i_13_100_3127_0,
    i_13_100_3129_0, i_13_100_3130_0, i_13_100_3135_0, i_13_100_3217_0,
    i_13_100_3220_0, i_13_100_3265_0, i_13_100_3291_0, i_13_100_3312_0,
    i_13_100_3315_0, i_13_100_3376_0, i_13_100_3399_0, i_13_100_3417_0,
    i_13_100_3453_0, i_13_100_3639_0, i_13_100_3702_0, i_13_100_3741_0,
    i_13_100_3822_0, i_13_100_3834_0, i_13_100_3892_0, i_13_100_3940_0,
    i_13_100_3994_0, i_13_100_4045_0, i_13_100_4056_0, i_13_100_4057_0,
    i_13_100_4065_0, i_13_100_4083_0, i_13_100_4094_0, i_13_100_4153_0,
    i_13_100_4164_0, i_13_100_4188_0, i_13_100_4234_0, i_13_100_4251_0,
    i_13_100_4269_0, i_13_100_4273_0, i_13_100_4274_0, i_13_100_4324_0,
    i_13_100_4360_0, i_13_100_4526_0, i_13_100_4533_0, i_13_100_4606_0;
  output o_13_100_0_0;
  assign o_13_100_0_0 = ~((~i_13_100_616_0 & ((i_13_100_310_0 & i_13_100_4057_0 & ~i_13_100_4083_0) | (~i_13_100_1735_0 & ~i_13_100_2987_0 & i_13_100_4094_0))) | (i_13_100_259_0 & ~i_13_100_1780_0 & i_13_100_4057_0) | (~i_13_100_474_0 & ~i_13_100_1996_0 & ~i_13_100_4083_0) | (~i_13_100_448_0 & ~i_13_100_2940_0) | (~i_13_100_4188_0 & i_13_100_4269_0 & ~i_13_100_4273_0) | (~i_13_100_48_0 & ~i_13_100_697_0 & ~i_13_100_1402_0 & ~i_13_100_2004_0 & ~i_13_100_3741_0 & ~i_13_100_4251_0 & ~i_13_100_4274_0));
endmodule



// Benchmark "kernel_13_101" written by ABC on Sun Jul 19 10:46:50 2020

module kernel_13_101 ( 
    i_13_101_51_0, i_13_101_52_0, i_13_101_105_0, i_13_101_106_0,
    i_13_101_312_0, i_13_101_381_0, i_13_101_508_0, i_13_101_537_0,
    i_13_101_552_0, i_13_101_553_0, i_13_101_655_0, i_13_101_679_0,
    i_13_101_691_0, i_13_101_817_0, i_13_101_843_0, i_13_101_983_0,
    i_13_101_984_0, i_13_101_985_0, i_13_101_1068_0, i_13_101_1069_0,
    i_13_101_1258_0, i_13_101_1300_0, i_13_101_1326_0, i_13_101_1329_0,
    i_13_101_1330_0, i_13_101_1345_0, i_13_101_1429_0, i_13_101_1492_0,
    i_13_101_1511_0, i_13_101_1516_0, i_13_101_1518_0, i_13_101_1519_0,
    i_13_101_1572_0, i_13_101_1573_0, i_13_101_1714_0, i_13_101_1778_0,
    i_13_101_1779_0, i_13_101_1803_0, i_13_101_1861_0, i_13_101_1885_0,
    i_13_101_1906_0, i_13_101_1911_0, i_13_101_1912_0, i_13_101_2002_0,
    i_13_101_2049_0, i_13_101_2059_0, i_13_101_2109_0, i_13_101_2175_0,
    i_13_101_2242_0, i_13_101_2243_0, i_13_101_2361_0, i_13_101_2409_0,
    i_13_101_2410_0, i_13_101_2464_0, i_13_101_2469_0, i_13_101_2470_0,
    i_13_101_2472_0, i_13_101_2533_0, i_13_101_2617_0, i_13_101_2693_0,
    i_13_101_2698_0, i_13_101_2725_0, i_13_101_2901_0, i_13_101_2919_0,
    i_13_101_2920_0, i_13_101_2982_0, i_13_101_2983_0, i_13_101_3030_0,
    i_13_101_3099_0, i_13_101_3111_0, i_13_101_3118_0, i_13_101_3130_0,
    i_13_101_3209_0, i_13_101_3346_0, i_13_101_3417_0, i_13_101_3418_0,
    i_13_101_3490_0, i_13_101_3525_0, i_13_101_3526_0, i_13_101_3535_0,
    i_13_101_3729_0, i_13_101_3769_0, i_13_101_3822_0, i_13_101_3864_0,
    i_13_101_3865_0, i_13_101_3891_0, i_13_101_3999_0, i_13_101_4038_0,
    i_13_101_4047_0, i_13_101_4048_0, i_13_101_4066_0, i_13_101_4119_0,
    i_13_101_4125_0, i_13_101_4126_0, i_13_101_4270_0, i_13_101_4323_0,
    i_13_101_4332_0, i_13_101_4353_0, i_13_101_4530_0, i_13_101_4569_0,
    o_13_101_0_0  );
  input  i_13_101_51_0, i_13_101_52_0, i_13_101_105_0, i_13_101_106_0,
    i_13_101_312_0, i_13_101_381_0, i_13_101_508_0, i_13_101_537_0,
    i_13_101_552_0, i_13_101_553_0, i_13_101_655_0, i_13_101_679_0,
    i_13_101_691_0, i_13_101_817_0, i_13_101_843_0, i_13_101_983_0,
    i_13_101_984_0, i_13_101_985_0, i_13_101_1068_0, i_13_101_1069_0,
    i_13_101_1258_0, i_13_101_1300_0, i_13_101_1326_0, i_13_101_1329_0,
    i_13_101_1330_0, i_13_101_1345_0, i_13_101_1429_0, i_13_101_1492_0,
    i_13_101_1511_0, i_13_101_1516_0, i_13_101_1518_0, i_13_101_1519_0,
    i_13_101_1572_0, i_13_101_1573_0, i_13_101_1714_0, i_13_101_1778_0,
    i_13_101_1779_0, i_13_101_1803_0, i_13_101_1861_0, i_13_101_1885_0,
    i_13_101_1906_0, i_13_101_1911_0, i_13_101_1912_0, i_13_101_2002_0,
    i_13_101_2049_0, i_13_101_2059_0, i_13_101_2109_0, i_13_101_2175_0,
    i_13_101_2242_0, i_13_101_2243_0, i_13_101_2361_0, i_13_101_2409_0,
    i_13_101_2410_0, i_13_101_2464_0, i_13_101_2469_0, i_13_101_2470_0,
    i_13_101_2472_0, i_13_101_2533_0, i_13_101_2617_0, i_13_101_2693_0,
    i_13_101_2698_0, i_13_101_2725_0, i_13_101_2901_0, i_13_101_2919_0,
    i_13_101_2920_0, i_13_101_2982_0, i_13_101_2983_0, i_13_101_3030_0,
    i_13_101_3099_0, i_13_101_3111_0, i_13_101_3118_0, i_13_101_3130_0,
    i_13_101_3209_0, i_13_101_3346_0, i_13_101_3417_0, i_13_101_3418_0,
    i_13_101_3490_0, i_13_101_3525_0, i_13_101_3526_0, i_13_101_3535_0,
    i_13_101_3729_0, i_13_101_3769_0, i_13_101_3822_0, i_13_101_3864_0,
    i_13_101_3865_0, i_13_101_3891_0, i_13_101_3999_0, i_13_101_4038_0,
    i_13_101_4047_0, i_13_101_4048_0, i_13_101_4066_0, i_13_101_4119_0,
    i_13_101_4125_0, i_13_101_4126_0, i_13_101_4270_0, i_13_101_4323_0,
    i_13_101_4332_0, i_13_101_4353_0, i_13_101_4530_0, i_13_101_4569_0;
  output o_13_101_0_0;
  assign o_13_101_0_0 = ~((i_13_101_1778_0 & i_13_101_3490_0) | (~i_13_101_52_0 & ~i_13_101_3111_0) | (~i_13_101_679_0 & i_13_101_2617_0));
endmodule



// Benchmark "kernel_13_102" written by ABC on Sun Jul 19 10:46:51 2020

module kernel_13_102 ( 
    i_13_102_48_0, i_13_102_79_0, i_13_102_251_0, i_13_102_277_0,
    i_13_102_310_0, i_13_102_319_0, i_13_102_340_0, i_13_102_409_0,
    i_13_102_597_0, i_13_102_643_0, i_13_102_664_0, i_13_102_745_0,
    i_13_102_760_0, i_13_102_1023_0, i_13_102_1024_0, i_13_102_1075_0,
    i_13_102_1096_0, i_13_102_1120_0, i_13_102_1140_0, i_13_102_1213_0,
    i_13_102_1266_0, i_13_102_1329_0, i_13_102_1403_0, i_13_102_1429_0,
    i_13_102_1430_0, i_13_102_1437_0, i_13_102_1482_0, i_13_102_1507_0,
    i_13_102_1573_0, i_13_102_1597_0, i_13_102_1626_0, i_13_102_1627_0,
    i_13_102_1634_0, i_13_102_1642_0, i_13_102_1686_0, i_13_102_1726_0,
    i_13_102_1780_0, i_13_102_1795_0, i_13_102_1844_0, i_13_102_2030_0,
    i_13_102_2106_0, i_13_102_2200_0, i_13_102_2272_0, i_13_102_2451_0,
    i_13_102_2454_0, i_13_102_2455_0, i_13_102_2541_0, i_13_102_2542_0,
    i_13_102_2545_0, i_13_102_2650_0, i_13_102_2708_0, i_13_102_2715_0,
    i_13_102_2716_0, i_13_102_2743_0, i_13_102_2770_0, i_13_102_2794_0,
    i_13_102_2904_0, i_13_102_2914_0, i_13_102_2919_0, i_13_102_2920_0,
    i_13_102_2921_0, i_13_102_3030_0, i_13_102_3105_0, i_13_102_3145_0,
    i_13_102_3244_0, i_13_102_3383_0, i_13_102_3388_0, i_13_102_3411_0,
    i_13_102_3412_0, i_13_102_3417_0, i_13_102_3418_0, i_13_102_3454_0,
    i_13_102_3463_0, i_13_102_3490_0, i_13_102_3535_0, i_13_102_3559_0,
    i_13_102_3568_0, i_13_102_3572_0, i_13_102_3574_0, i_13_102_3577_0,
    i_13_102_3688_0, i_13_102_3699_0, i_13_102_3877_0, i_13_102_3922_0,
    i_13_102_3928_0, i_13_102_3937_0, i_13_102_4036_0, i_13_102_4063_0,
    i_13_102_4255_0, i_13_102_4338_0, i_13_102_4352_0, i_13_102_4372_0,
    i_13_102_4373_0, i_13_102_4449_0, i_13_102_4522_0, i_13_102_4523_0,
    i_13_102_4525_0, i_13_102_4540_0, i_13_102_4558_0, i_13_102_4561_0,
    o_13_102_0_0  );
  input  i_13_102_48_0, i_13_102_79_0, i_13_102_251_0, i_13_102_277_0,
    i_13_102_310_0, i_13_102_319_0, i_13_102_340_0, i_13_102_409_0,
    i_13_102_597_0, i_13_102_643_0, i_13_102_664_0, i_13_102_745_0,
    i_13_102_760_0, i_13_102_1023_0, i_13_102_1024_0, i_13_102_1075_0,
    i_13_102_1096_0, i_13_102_1120_0, i_13_102_1140_0, i_13_102_1213_0,
    i_13_102_1266_0, i_13_102_1329_0, i_13_102_1403_0, i_13_102_1429_0,
    i_13_102_1430_0, i_13_102_1437_0, i_13_102_1482_0, i_13_102_1507_0,
    i_13_102_1573_0, i_13_102_1597_0, i_13_102_1626_0, i_13_102_1627_0,
    i_13_102_1634_0, i_13_102_1642_0, i_13_102_1686_0, i_13_102_1726_0,
    i_13_102_1780_0, i_13_102_1795_0, i_13_102_1844_0, i_13_102_2030_0,
    i_13_102_2106_0, i_13_102_2200_0, i_13_102_2272_0, i_13_102_2451_0,
    i_13_102_2454_0, i_13_102_2455_0, i_13_102_2541_0, i_13_102_2542_0,
    i_13_102_2545_0, i_13_102_2650_0, i_13_102_2708_0, i_13_102_2715_0,
    i_13_102_2716_0, i_13_102_2743_0, i_13_102_2770_0, i_13_102_2794_0,
    i_13_102_2904_0, i_13_102_2914_0, i_13_102_2919_0, i_13_102_2920_0,
    i_13_102_2921_0, i_13_102_3030_0, i_13_102_3105_0, i_13_102_3145_0,
    i_13_102_3244_0, i_13_102_3383_0, i_13_102_3388_0, i_13_102_3411_0,
    i_13_102_3412_0, i_13_102_3417_0, i_13_102_3418_0, i_13_102_3454_0,
    i_13_102_3463_0, i_13_102_3490_0, i_13_102_3535_0, i_13_102_3559_0,
    i_13_102_3568_0, i_13_102_3572_0, i_13_102_3574_0, i_13_102_3577_0,
    i_13_102_3688_0, i_13_102_3699_0, i_13_102_3877_0, i_13_102_3922_0,
    i_13_102_3928_0, i_13_102_3937_0, i_13_102_4036_0, i_13_102_4063_0,
    i_13_102_4255_0, i_13_102_4338_0, i_13_102_4352_0, i_13_102_4372_0,
    i_13_102_4373_0, i_13_102_4449_0, i_13_102_4522_0, i_13_102_4523_0,
    i_13_102_4525_0, i_13_102_4540_0, i_13_102_4558_0, i_13_102_4561_0;
  output o_13_102_0_0;
  assign o_13_102_0_0 = ~((~i_13_102_3922_0 & ((~i_13_102_79_0 & ~i_13_102_2200_0) | (~i_13_102_1780_0 & i_13_102_3244_0))) | (~i_13_102_2716_0 & ~i_13_102_2743_0 & ~i_13_102_3463_0) | (i_13_102_1597_0 & ~i_13_102_2919_0 & ~i_13_102_3568_0));
endmodule



// Benchmark "kernel_13_103" written by ABC on Sun Jul 19 10:46:52 2020

module kernel_13_103 ( 
    i_13_103_23_0, i_13_103_49_0, i_13_103_50_0, i_13_103_73_0,
    i_13_103_74_0, i_13_103_118_0, i_13_103_163_0, i_13_103_198_0,
    i_13_103_230_0, i_13_103_248_0, i_13_103_275_0, i_13_103_338_0,
    i_13_103_515_0, i_13_103_518_0, i_13_103_535_0, i_13_103_578_0,
    i_13_103_676_0, i_13_103_695_0, i_13_103_712_0, i_13_103_742_0,
    i_13_103_839_0, i_13_103_977_0, i_13_103_1082_0, i_13_103_1208_0,
    i_13_103_1210_0, i_13_103_1243_0, i_13_103_1262_0, i_13_103_1307_0,
    i_13_103_1397_0, i_13_103_1424_0, i_13_103_1505_0, i_13_103_1570_0,
    i_13_103_1658_0, i_13_103_1900_0, i_13_103_1918_0, i_13_103_1919_0,
    i_13_103_1928_0, i_13_103_1936_0, i_13_103_1954_0, i_13_103_1991_0,
    i_13_103_2030_0, i_13_103_2057_0, i_13_103_2173_0, i_13_103_2187_0,
    i_13_103_2261_0, i_13_103_2362_0, i_13_103_2395_0, i_13_103_2450_0,
    i_13_103_2452_0, i_13_103_2453_0, i_13_103_2512_0, i_13_103_2531_0,
    i_13_103_2549_0, i_13_103_2552_0, i_13_103_2576_0, i_13_103_2711_0,
    i_13_103_2741_0, i_13_103_2749_0, i_13_103_2764_0, i_13_103_2765_0,
    i_13_103_2785_0, i_13_103_2956_0, i_13_103_2963_0, i_13_103_3026_0,
    i_13_103_3061_0, i_13_103_3062_0, i_13_103_3128_0, i_13_103_3313_0,
    i_13_103_3370_0, i_13_103_3371_0, i_13_103_3376_0, i_13_103_3377_0,
    i_13_103_3415_0, i_13_103_3416_0, i_13_103_3475_0, i_13_103_3506_0,
    i_13_103_3533_0, i_13_103_3596_0, i_13_103_3613_0, i_13_103_3646_0,
    i_13_103_3647_0, i_13_103_3656_0, i_13_103_3671_0, i_13_103_3710_0,
    i_13_103_3719_0, i_13_103_3793_0, i_13_103_3872_0, i_13_103_3902_0,
    i_13_103_3920_0, i_13_103_4086_0, i_13_103_4123_0, i_13_103_4262_0,
    i_13_103_4331_0, i_13_103_4351_0, i_13_103_4367_0, i_13_103_4430_0,
    i_13_103_4450_0, i_13_103_4451_0, i_13_103_4557_0, i_13_103_4591_0,
    o_13_103_0_0  );
  input  i_13_103_23_0, i_13_103_49_0, i_13_103_50_0, i_13_103_73_0,
    i_13_103_74_0, i_13_103_118_0, i_13_103_163_0, i_13_103_198_0,
    i_13_103_230_0, i_13_103_248_0, i_13_103_275_0, i_13_103_338_0,
    i_13_103_515_0, i_13_103_518_0, i_13_103_535_0, i_13_103_578_0,
    i_13_103_676_0, i_13_103_695_0, i_13_103_712_0, i_13_103_742_0,
    i_13_103_839_0, i_13_103_977_0, i_13_103_1082_0, i_13_103_1208_0,
    i_13_103_1210_0, i_13_103_1243_0, i_13_103_1262_0, i_13_103_1307_0,
    i_13_103_1397_0, i_13_103_1424_0, i_13_103_1505_0, i_13_103_1570_0,
    i_13_103_1658_0, i_13_103_1900_0, i_13_103_1918_0, i_13_103_1919_0,
    i_13_103_1928_0, i_13_103_1936_0, i_13_103_1954_0, i_13_103_1991_0,
    i_13_103_2030_0, i_13_103_2057_0, i_13_103_2173_0, i_13_103_2187_0,
    i_13_103_2261_0, i_13_103_2362_0, i_13_103_2395_0, i_13_103_2450_0,
    i_13_103_2452_0, i_13_103_2453_0, i_13_103_2512_0, i_13_103_2531_0,
    i_13_103_2549_0, i_13_103_2552_0, i_13_103_2576_0, i_13_103_2711_0,
    i_13_103_2741_0, i_13_103_2749_0, i_13_103_2764_0, i_13_103_2765_0,
    i_13_103_2785_0, i_13_103_2956_0, i_13_103_2963_0, i_13_103_3026_0,
    i_13_103_3061_0, i_13_103_3062_0, i_13_103_3128_0, i_13_103_3313_0,
    i_13_103_3370_0, i_13_103_3371_0, i_13_103_3376_0, i_13_103_3377_0,
    i_13_103_3415_0, i_13_103_3416_0, i_13_103_3475_0, i_13_103_3506_0,
    i_13_103_3533_0, i_13_103_3596_0, i_13_103_3613_0, i_13_103_3646_0,
    i_13_103_3647_0, i_13_103_3656_0, i_13_103_3671_0, i_13_103_3710_0,
    i_13_103_3719_0, i_13_103_3793_0, i_13_103_3872_0, i_13_103_3902_0,
    i_13_103_3920_0, i_13_103_4086_0, i_13_103_4123_0, i_13_103_4262_0,
    i_13_103_4331_0, i_13_103_4351_0, i_13_103_4367_0, i_13_103_4430_0,
    i_13_103_4450_0, i_13_103_4451_0, i_13_103_4557_0, i_13_103_4591_0;
  output o_13_103_0_0;
  assign o_13_103_0_0 = ~(i_13_103_1954_0 | (~i_13_103_1424_0 & ~i_13_103_2765_0) | (~i_13_103_50_0 & ~i_13_103_1658_0 & ~i_13_103_2030_0));
endmodule



// Benchmark "kernel_13_104" written by ABC on Sun Jul 19 10:46:52 2020

module kernel_13_104 ( 
    i_13_104_49_0, i_13_104_52_0, i_13_104_53_0, i_13_104_94_0,
    i_13_104_95_0, i_13_104_98_0, i_13_104_106_0, i_13_104_107_0,
    i_13_104_139_0, i_13_104_166_0, i_13_104_179_0, i_13_104_283_0,
    i_13_104_311_0, i_13_104_319_0, i_13_104_337_0, i_13_104_367_0,
    i_13_104_512_0, i_13_104_554_0, i_13_104_575_0, i_13_104_655_0,
    i_13_104_656_0, i_13_104_670_0, i_13_104_671_0, i_13_104_679_0,
    i_13_104_680_0, i_13_104_688_0, i_13_104_691_0, i_13_104_692_0,
    i_13_104_823_0, i_13_104_844_0, i_13_104_845_0, i_13_104_889_0,
    i_13_104_962_0, i_13_104_974_0, i_13_104_985_0, i_13_104_986_0,
    i_13_104_1052_0, i_13_104_1222_0, i_13_104_1331_0, i_13_104_1519_0,
    i_13_104_1520_0, i_13_104_1627_0, i_13_104_1636_0, i_13_104_1697_0,
    i_13_104_1789_0, i_13_104_1839_0, i_13_104_1861_0, i_13_104_1942_0,
    i_13_104_2032_0, i_13_104_2173_0, i_13_104_2182_0, i_13_104_2438_0,
    i_13_104_2618_0, i_13_104_2680_0, i_13_104_2725_0, i_13_104_2753_0,
    i_13_104_2905_0, i_13_104_2938_0, i_13_104_3002_0, i_13_104_3028_0,
    i_13_104_3112_0, i_13_104_3130_0, i_13_104_3155_0, i_13_104_3166_0,
    i_13_104_3167_0, i_13_104_3217_0, i_13_104_3218_0, i_13_104_3227_0,
    i_13_104_3280_0, i_13_104_3374_0, i_13_104_3418_0, i_13_104_3479_0,
    i_13_104_3505_0, i_13_104_3526_0, i_13_104_3536_0, i_13_104_3685_0,
    i_13_104_3719_0, i_13_104_3739_0, i_13_104_3769_0, i_13_104_3770_0,
    i_13_104_3865_0, i_13_104_3866_0, i_13_104_3892_0, i_13_104_3893_0,
    i_13_104_4021_0, i_13_104_4022_0, i_13_104_4049_0, i_13_104_4120_0,
    i_13_104_4121_0, i_13_104_4126_0, i_13_104_4127_0, i_13_104_4265_0,
    i_13_104_4270_0, i_13_104_4339_0, i_13_104_4340_0, i_13_104_4354_0,
    i_13_104_4534_0, i_13_104_4561_0, i_13_104_4570_0, i_13_104_4571_0,
    o_13_104_0_0  );
  input  i_13_104_49_0, i_13_104_52_0, i_13_104_53_0, i_13_104_94_0,
    i_13_104_95_0, i_13_104_98_0, i_13_104_106_0, i_13_104_107_0,
    i_13_104_139_0, i_13_104_166_0, i_13_104_179_0, i_13_104_283_0,
    i_13_104_311_0, i_13_104_319_0, i_13_104_337_0, i_13_104_367_0,
    i_13_104_512_0, i_13_104_554_0, i_13_104_575_0, i_13_104_655_0,
    i_13_104_656_0, i_13_104_670_0, i_13_104_671_0, i_13_104_679_0,
    i_13_104_680_0, i_13_104_688_0, i_13_104_691_0, i_13_104_692_0,
    i_13_104_823_0, i_13_104_844_0, i_13_104_845_0, i_13_104_889_0,
    i_13_104_962_0, i_13_104_974_0, i_13_104_985_0, i_13_104_986_0,
    i_13_104_1052_0, i_13_104_1222_0, i_13_104_1331_0, i_13_104_1519_0,
    i_13_104_1520_0, i_13_104_1627_0, i_13_104_1636_0, i_13_104_1697_0,
    i_13_104_1789_0, i_13_104_1839_0, i_13_104_1861_0, i_13_104_1942_0,
    i_13_104_2032_0, i_13_104_2173_0, i_13_104_2182_0, i_13_104_2438_0,
    i_13_104_2618_0, i_13_104_2680_0, i_13_104_2725_0, i_13_104_2753_0,
    i_13_104_2905_0, i_13_104_2938_0, i_13_104_3002_0, i_13_104_3028_0,
    i_13_104_3112_0, i_13_104_3130_0, i_13_104_3155_0, i_13_104_3166_0,
    i_13_104_3167_0, i_13_104_3217_0, i_13_104_3218_0, i_13_104_3227_0,
    i_13_104_3280_0, i_13_104_3374_0, i_13_104_3418_0, i_13_104_3479_0,
    i_13_104_3505_0, i_13_104_3526_0, i_13_104_3536_0, i_13_104_3685_0,
    i_13_104_3719_0, i_13_104_3739_0, i_13_104_3769_0, i_13_104_3770_0,
    i_13_104_3865_0, i_13_104_3866_0, i_13_104_3892_0, i_13_104_3893_0,
    i_13_104_4021_0, i_13_104_4022_0, i_13_104_4049_0, i_13_104_4120_0,
    i_13_104_4121_0, i_13_104_4126_0, i_13_104_4127_0, i_13_104_4265_0,
    i_13_104_4270_0, i_13_104_4339_0, i_13_104_4340_0, i_13_104_4354_0,
    i_13_104_4534_0, i_13_104_4561_0, i_13_104_4570_0, i_13_104_4571_0;
  output o_13_104_0_0;
  assign o_13_104_0_0 = ~((~i_13_104_3893_0 & i_13_104_4571_0) | (~i_13_104_4049_0 & ~i_13_104_4354_0) | (~i_13_104_671_0 & ~i_13_104_679_0 & ~i_13_104_4265_0) | (~i_13_104_53_0 & ~i_13_104_575_0 & ~i_13_104_3112_0));
endmodule



// Benchmark "kernel_13_105" written by ABC on Sun Jul 19 10:46:53 2020

module kernel_13_105 ( 
    i_13_105_31_0, i_13_105_33_0, i_13_105_38_0, i_13_105_67_0,
    i_13_105_76_0, i_13_105_121_0, i_13_105_138_0, i_13_105_139_0,
    i_13_105_165_0, i_13_105_184_0, i_13_105_229_0, i_13_105_230_0,
    i_13_105_254_0, i_13_105_284_0, i_13_105_382_0, i_13_105_401_0,
    i_13_105_415_0, i_13_105_443_0, i_13_105_474_0, i_13_105_516_0,
    i_13_105_535_0, i_13_105_537_0, i_13_105_571_0, i_13_105_578_0,
    i_13_105_636_0, i_13_105_661_0, i_13_105_673_0, i_13_105_677_0,
    i_13_105_698_0, i_13_105_704_0, i_13_105_760_0, i_13_105_797_0,
    i_13_105_822_0, i_13_105_850_0, i_13_105_884_0, i_13_105_944_0,
    i_13_105_950_0, i_13_105_959_0, i_13_105_1042_0, i_13_105_1135_0,
    i_13_105_1218_0, i_13_105_1286_0, i_13_105_1339_0, i_13_105_1394_0,
    i_13_105_1472_0, i_13_105_1723_0, i_13_105_1725_0, i_13_105_1734_0,
    i_13_105_1794_0, i_13_105_1858_0, i_13_105_1943_0, i_13_105_1993_0,
    i_13_105_1994_0, i_13_105_1999_0, i_13_105_2000_0, i_13_105_2012_0,
    i_13_105_2060_0, i_13_105_2170_0, i_13_105_2407_0, i_13_105_2418_0,
    i_13_105_2434_0, i_13_105_2501_0, i_13_105_2509_0, i_13_105_2668_0,
    i_13_105_2679_0, i_13_105_2722_0, i_13_105_2749_0, i_13_105_2805_0,
    i_13_105_2858_0, i_13_105_2872_0, i_13_105_2897_0, i_13_105_3036_0,
    i_13_105_3064_0, i_13_105_3108_0, i_13_105_3109_0, i_13_105_3329_0,
    i_13_105_3374_0, i_13_105_3395_0, i_13_105_3444_0, i_13_105_3604_0,
    i_13_105_3622_0, i_13_105_3637_0, i_13_105_3651_0, i_13_105_3786_0,
    i_13_105_3794_0, i_13_105_3894_0, i_13_105_3974_0, i_13_105_3984_0,
    i_13_105_3988_0, i_13_105_4050_0, i_13_105_4064_0, i_13_105_4078_0,
    i_13_105_4094_0, i_13_105_4121_0, i_13_105_4195_0, i_13_105_4265_0,
    i_13_105_4336_0, i_13_105_4370_0, i_13_105_4454_0, i_13_105_4567_0,
    o_13_105_0_0  );
  input  i_13_105_31_0, i_13_105_33_0, i_13_105_38_0, i_13_105_67_0,
    i_13_105_76_0, i_13_105_121_0, i_13_105_138_0, i_13_105_139_0,
    i_13_105_165_0, i_13_105_184_0, i_13_105_229_0, i_13_105_230_0,
    i_13_105_254_0, i_13_105_284_0, i_13_105_382_0, i_13_105_401_0,
    i_13_105_415_0, i_13_105_443_0, i_13_105_474_0, i_13_105_516_0,
    i_13_105_535_0, i_13_105_537_0, i_13_105_571_0, i_13_105_578_0,
    i_13_105_636_0, i_13_105_661_0, i_13_105_673_0, i_13_105_677_0,
    i_13_105_698_0, i_13_105_704_0, i_13_105_760_0, i_13_105_797_0,
    i_13_105_822_0, i_13_105_850_0, i_13_105_884_0, i_13_105_944_0,
    i_13_105_950_0, i_13_105_959_0, i_13_105_1042_0, i_13_105_1135_0,
    i_13_105_1218_0, i_13_105_1286_0, i_13_105_1339_0, i_13_105_1394_0,
    i_13_105_1472_0, i_13_105_1723_0, i_13_105_1725_0, i_13_105_1734_0,
    i_13_105_1794_0, i_13_105_1858_0, i_13_105_1943_0, i_13_105_1993_0,
    i_13_105_1994_0, i_13_105_1999_0, i_13_105_2000_0, i_13_105_2012_0,
    i_13_105_2060_0, i_13_105_2170_0, i_13_105_2407_0, i_13_105_2418_0,
    i_13_105_2434_0, i_13_105_2501_0, i_13_105_2509_0, i_13_105_2668_0,
    i_13_105_2679_0, i_13_105_2722_0, i_13_105_2749_0, i_13_105_2805_0,
    i_13_105_2858_0, i_13_105_2872_0, i_13_105_2897_0, i_13_105_3036_0,
    i_13_105_3064_0, i_13_105_3108_0, i_13_105_3109_0, i_13_105_3329_0,
    i_13_105_3374_0, i_13_105_3395_0, i_13_105_3444_0, i_13_105_3604_0,
    i_13_105_3622_0, i_13_105_3637_0, i_13_105_3651_0, i_13_105_3786_0,
    i_13_105_3794_0, i_13_105_3894_0, i_13_105_3974_0, i_13_105_3984_0,
    i_13_105_3988_0, i_13_105_4050_0, i_13_105_4064_0, i_13_105_4078_0,
    i_13_105_4094_0, i_13_105_4121_0, i_13_105_4195_0, i_13_105_4265_0,
    i_13_105_4336_0, i_13_105_4370_0, i_13_105_4454_0, i_13_105_4567_0;
  output o_13_105_0_0;
  assign o_13_105_0_0 = 0;
endmodule



// Benchmark "kernel_13_106" written by ABC on Sun Jul 19 10:46:54 2020

module kernel_13_106 ( 
    i_13_106_45_0, i_13_106_48_0, i_13_106_121_0, i_13_106_172_0,
    i_13_106_226_0, i_13_106_234_0, i_13_106_279_0, i_13_106_333_0,
    i_13_106_414_0, i_13_106_553_0, i_13_106_607_0, i_13_106_612_0,
    i_13_106_613_0, i_13_106_640_0, i_13_106_643_0, i_13_106_657_0,
    i_13_106_658_0, i_13_106_660_0, i_13_106_666_0, i_13_106_684_0,
    i_13_106_685_0, i_13_106_711_0, i_13_106_760_0, i_13_106_828_0,
    i_13_106_939_0, i_13_106_955_0, i_13_106_1071_0, i_13_106_1072_0,
    i_13_106_1116_0, i_13_106_1117_0, i_13_106_1225_0, i_13_106_1228_0,
    i_13_106_1232_0, i_13_106_1286_0, i_13_106_1390_0, i_13_106_1440_0,
    i_13_106_1493_0, i_13_106_1521_0, i_13_106_1522_0, i_13_106_1554_0,
    i_13_106_1638_0, i_13_106_1639_0, i_13_106_1696_0, i_13_106_1729_0,
    i_13_106_1736_0, i_13_106_1764_0, i_13_106_1792_0, i_13_106_1795_0,
    i_13_106_1801_0, i_13_106_1891_0, i_13_106_1926_0, i_13_106_1927_0,
    i_13_106_1944_0, i_13_106_2100_0, i_13_106_2115_0, i_13_106_2142_0,
    i_13_106_2211_0, i_13_106_2254_0, i_13_106_2299_0, i_13_106_2303_0,
    i_13_106_2313_0, i_13_106_2340_0, i_13_106_2376_0, i_13_106_2461_0,
    i_13_106_2595_0, i_13_106_2676_0, i_13_106_2677_0, i_13_106_2678_0,
    i_13_106_2721_0, i_13_106_2847_0, i_13_106_2848_0, i_13_106_2880_0,
    i_13_106_2881_0, i_13_106_3114_0, i_13_106_3261_0, i_13_106_3267_0,
    i_13_106_3367_0, i_13_106_3420_0, i_13_106_3421_0, i_13_106_3423_0,
    i_13_106_3546_0, i_13_106_3555_0, i_13_106_3564_0, i_13_106_3636_0,
    i_13_106_3753_0, i_13_106_3754_0, i_13_106_3892_0, i_13_106_3910_0,
    i_13_106_3924_0, i_13_106_4063_0, i_13_106_4186_0, i_13_106_4266_0,
    i_13_106_4280_0, i_13_106_4293_0, i_13_106_4294_0, i_13_106_4311_0,
    i_13_106_4467_0, i_13_106_4509_0, i_13_106_4593_0, i_13_106_4594_0,
    o_13_106_0_0  );
  input  i_13_106_45_0, i_13_106_48_0, i_13_106_121_0, i_13_106_172_0,
    i_13_106_226_0, i_13_106_234_0, i_13_106_279_0, i_13_106_333_0,
    i_13_106_414_0, i_13_106_553_0, i_13_106_607_0, i_13_106_612_0,
    i_13_106_613_0, i_13_106_640_0, i_13_106_643_0, i_13_106_657_0,
    i_13_106_658_0, i_13_106_660_0, i_13_106_666_0, i_13_106_684_0,
    i_13_106_685_0, i_13_106_711_0, i_13_106_760_0, i_13_106_828_0,
    i_13_106_939_0, i_13_106_955_0, i_13_106_1071_0, i_13_106_1072_0,
    i_13_106_1116_0, i_13_106_1117_0, i_13_106_1225_0, i_13_106_1228_0,
    i_13_106_1232_0, i_13_106_1286_0, i_13_106_1390_0, i_13_106_1440_0,
    i_13_106_1493_0, i_13_106_1521_0, i_13_106_1522_0, i_13_106_1554_0,
    i_13_106_1638_0, i_13_106_1639_0, i_13_106_1696_0, i_13_106_1729_0,
    i_13_106_1736_0, i_13_106_1764_0, i_13_106_1792_0, i_13_106_1795_0,
    i_13_106_1801_0, i_13_106_1891_0, i_13_106_1926_0, i_13_106_1927_0,
    i_13_106_1944_0, i_13_106_2100_0, i_13_106_2115_0, i_13_106_2142_0,
    i_13_106_2211_0, i_13_106_2254_0, i_13_106_2299_0, i_13_106_2303_0,
    i_13_106_2313_0, i_13_106_2340_0, i_13_106_2376_0, i_13_106_2461_0,
    i_13_106_2595_0, i_13_106_2676_0, i_13_106_2677_0, i_13_106_2678_0,
    i_13_106_2721_0, i_13_106_2847_0, i_13_106_2848_0, i_13_106_2880_0,
    i_13_106_2881_0, i_13_106_3114_0, i_13_106_3261_0, i_13_106_3267_0,
    i_13_106_3367_0, i_13_106_3420_0, i_13_106_3421_0, i_13_106_3423_0,
    i_13_106_3546_0, i_13_106_3555_0, i_13_106_3564_0, i_13_106_3636_0,
    i_13_106_3753_0, i_13_106_3754_0, i_13_106_3892_0, i_13_106_3910_0,
    i_13_106_3924_0, i_13_106_4063_0, i_13_106_4186_0, i_13_106_4266_0,
    i_13_106_4280_0, i_13_106_4293_0, i_13_106_4294_0, i_13_106_4311_0,
    i_13_106_4467_0, i_13_106_4509_0, i_13_106_4593_0, i_13_106_4594_0;
  output o_13_106_0_0;
  assign o_13_106_0_0 = ~((~i_13_106_4509_0 & (~i_13_106_1764_0 | ~i_13_106_4311_0)) | ~i_13_106_3753_0 | (i_13_106_279_0 & ~i_13_106_414_0 & ~i_13_106_1071_0 & i_13_106_3910_0));
endmodule



// Benchmark "kernel_13_107" written by ABC on Sun Jul 19 10:46:55 2020

module kernel_13_107 ( 
    i_13_107_46_0, i_13_107_64_0, i_13_107_172_0, i_13_107_279_0,
    i_13_107_355_0, i_13_107_516_0, i_13_107_522_0, i_13_107_523_0,
    i_13_107_626_0, i_13_107_657_0, i_13_107_658_0, i_13_107_667_0,
    i_13_107_723_0, i_13_107_724_0, i_13_107_793_0, i_13_107_847_0,
    i_13_107_930_0, i_13_107_937_0, i_13_107_938_0, i_13_107_1017_0,
    i_13_107_1018_0, i_13_107_1071_0, i_13_107_1072_0, i_13_107_1093_0,
    i_13_107_1094_0, i_13_107_1099_0, i_13_107_1201_0, i_13_107_1225_0,
    i_13_107_1226_0, i_13_107_1279_0, i_13_107_1282_0, i_13_107_1315_0,
    i_13_107_1389_0, i_13_107_1423_0, i_13_107_1480_0, i_13_107_1486_0,
    i_13_107_1495_0, i_13_107_1523_0, i_13_107_1549_0, i_13_107_1630_0,
    i_13_107_1639_0, i_13_107_1792_0, i_13_107_1855_0, i_13_107_1884_0,
    i_13_107_1937_0, i_13_107_1955_0, i_13_107_2019_0, i_13_107_2020_0,
    i_13_107_2026_0, i_13_107_2127_0, i_13_107_2196_0, i_13_107_2197_0,
    i_13_107_2287_0, i_13_107_2317_0, i_13_107_2449_0, i_13_107_2452_0,
    i_13_107_2498_0, i_13_107_2539_0, i_13_107_2540_0, i_13_107_2592_0,
    i_13_107_2746_0, i_13_107_2917_0, i_13_107_2918_0, i_13_107_3029_0,
    i_13_107_3127_0, i_13_107_3241_0, i_13_107_3421_0, i_13_107_3422_0,
    i_13_107_3457_0, i_13_107_3458_0, i_13_107_3479_0, i_13_107_3483_0,
    i_13_107_3484_0, i_13_107_3485_0, i_13_107_3538_0, i_13_107_3574_0,
    i_13_107_3575_0, i_13_107_3595_0, i_13_107_3648_0, i_13_107_3738_0,
    i_13_107_3780_0, i_13_107_3781_0, i_13_107_3782_0, i_13_107_3820_0,
    i_13_107_3837_0, i_13_107_3918_0, i_13_107_4249_0, i_13_107_4250_0,
    i_13_107_4252_0, i_13_107_4257_0, i_13_107_4259_0, i_13_107_4321_0,
    i_13_107_4356_0, i_13_107_4366_0, i_13_107_4376_0, i_13_107_4446_0,
    i_13_107_4448_0, i_13_107_4450_0, i_13_107_4555_0, i_13_107_4604_0,
    o_13_107_0_0  );
  input  i_13_107_46_0, i_13_107_64_0, i_13_107_172_0, i_13_107_279_0,
    i_13_107_355_0, i_13_107_516_0, i_13_107_522_0, i_13_107_523_0,
    i_13_107_626_0, i_13_107_657_0, i_13_107_658_0, i_13_107_667_0,
    i_13_107_723_0, i_13_107_724_0, i_13_107_793_0, i_13_107_847_0,
    i_13_107_930_0, i_13_107_937_0, i_13_107_938_0, i_13_107_1017_0,
    i_13_107_1018_0, i_13_107_1071_0, i_13_107_1072_0, i_13_107_1093_0,
    i_13_107_1094_0, i_13_107_1099_0, i_13_107_1201_0, i_13_107_1225_0,
    i_13_107_1226_0, i_13_107_1279_0, i_13_107_1282_0, i_13_107_1315_0,
    i_13_107_1389_0, i_13_107_1423_0, i_13_107_1480_0, i_13_107_1486_0,
    i_13_107_1495_0, i_13_107_1523_0, i_13_107_1549_0, i_13_107_1630_0,
    i_13_107_1639_0, i_13_107_1792_0, i_13_107_1855_0, i_13_107_1884_0,
    i_13_107_1937_0, i_13_107_1955_0, i_13_107_2019_0, i_13_107_2020_0,
    i_13_107_2026_0, i_13_107_2127_0, i_13_107_2196_0, i_13_107_2197_0,
    i_13_107_2287_0, i_13_107_2317_0, i_13_107_2449_0, i_13_107_2452_0,
    i_13_107_2498_0, i_13_107_2539_0, i_13_107_2540_0, i_13_107_2592_0,
    i_13_107_2746_0, i_13_107_2917_0, i_13_107_2918_0, i_13_107_3029_0,
    i_13_107_3127_0, i_13_107_3241_0, i_13_107_3421_0, i_13_107_3422_0,
    i_13_107_3457_0, i_13_107_3458_0, i_13_107_3479_0, i_13_107_3483_0,
    i_13_107_3484_0, i_13_107_3485_0, i_13_107_3538_0, i_13_107_3574_0,
    i_13_107_3575_0, i_13_107_3595_0, i_13_107_3648_0, i_13_107_3738_0,
    i_13_107_3780_0, i_13_107_3781_0, i_13_107_3782_0, i_13_107_3820_0,
    i_13_107_3837_0, i_13_107_3918_0, i_13_107_4249_0, i_13_107_4250_0,
    i_13_107_4252_0, i_13_107_4257_0, i_13_107_4259_0, i_13_107_4321_0,
    i_13_107_4356_0, i_13_107_4366_0, i_13_107_4376_0, i_13_107_4446_0,
    i_13_107_4448_0, i_13_107_4450_0, i_13_107_4555_0, i_13_107_4604_0;
  output o_13_107_0_0;
  assign o_13_107_0_0 = ~(~i_13_107_4252_0 | (~i_13_107_938_0 & ~i_13_107_4376_0));
endmodule



// Benchmark "kernel_13_108" written by ABC on Sun Jul 19 10:46:56 2020

module kernel_13_108 ( 
    i_13_108_25_0, i_13_108_34_0, i_13_108_156_0, i_13_108_160_0,
    i_13_108_224_0, i_13_108_228_0, i_13_108_231_0, i_13_108_273_0,
    i_13_108_278_0, i_13_108_328_0, i_13_108_382_0, i_13_108_411_0,
    i_13_108_417_0, i_13_108_534_0, i_13_108_565_0, i_13_108_603_0,
    i_13_108_604_0, i_13_108_665_0, i_13_108_688_0, i_13_108_732_0,
    i_13_108_741_0, i_13_108_933_0, i_13_108_945_0, i_13_108_946_0,
    i_13_108_1083_0, i_13_108_1084_0, i_13_108_1120_0, i_13_108_1218_0,
    i_13_108_1269_0, i_13_108_1344_0, i_13_108_1354_0, i_13_108_1443_0,
    i_13_108_1444_0, i_13_108_1473_0, i_13_108_1569_0, i_13_108_1605_0,
    i_13_108_1620_0, i_13_108_1687_0, i_13_108_1769_0, i_13_108_1836_0,
    i_13_108_1857_0, i_13_108_1957_0, i_13_108_2001_0, i_13_108_2047_0,
    i_13_108_2056_0, i_13_108_2150_0, i_13_108_2275_0, i_13_108_2280_0,
    i_13_108_2421_0, i_13_108_2424_0, i_13_108_2430_0, i_13_108_2497_0,
    i_13_108_2584_0, i_13_108_2712_0, i_13_108_2721_0, i_13_108_2722_0,
    i_13_108_2725_0, i_13_108_2784_0, i_13_108_2786_0, i_13_108_2856_0,
    i_13_108_2857_0, i_13_108_2859_0, i_13_108_2860_0, i_13_108_3010_0,
    i_13_108_3063_0, i_13_108_3064_0, i_13_108_3066_0, i_13_108_3097_0,
    i_13_108_3100_0, i_13_108_3103_0, i_13_108_3213_0, i_13_108_3234_0,
    i_13_108_3238_0, i_13_108_3255_0, i_13_108_3334_0, i_13_108_3428_0,
    i_13_108_3442_0, i_13_108_3487_0, i_13_108_3541_0, i_13_108_3554_0,
    i_13_108_3684_0, i_13_108_3691_0, i_13_108_3702_0, i_13_108_3717_0,
    i_13_108_3865_0, i_13_108_3871_0, i_13_108_3931_0, i_13_108_3977_0,
    i_13_108_4020_0, i_13_108_4252_0, i_13_108_4270_0, i_13_108_4328_0,
    i_13_108_4337_0, i_13_108_4350_0, i_13_108_4351_0, i_13_108_4395_0,
    i_13_108_4398_0, i_13_108_4413_0, i_13_108_4517_0, i_13_108_4593_0,
    o_13_108_0_0  );
  input  i_13_108_25_0, i_13_108_34_0, i_13_108_156_0, i_13_108_160_0,
    i_13_108_224_0, i_13_108_228_0, i_13_108_231_0, i_13_108_273_0,
    i_13_108_278_0, i_13_108_328_0, i_13_108_382_0, i_13_108_411_0,
    i_13_108_417_0, i_13_108_534_0, i_13_108_565_0, i_13_108_603_0,
    i_13_108_604_0, i_13_108_665_0, i_13_108_688_0, i_13_108_732_0,
    i_13_108_741_0, i_13_108_933_0, i_13_108_945_0, i_13_108_946_0,
    i_13_108_1083_0, i_13_108_1084_0, i_13_108_1120_0, i_13_108_1218_0,
    i_13_108_1269_0, i_13_108_1344_0, i_13_108_1354_0, i_13_108_1443_0,
    i_13_108_1444_0, i_13_108_1473_0, i_13_108_1569_0, i_13_108_1605_0,
    i_13_108_1620_0, i_13_108_1687_0, i_13_108_1769_0, i_13_108_1836_0,
    i_13_108_1857_0, i_13_108_1957_0, i_13_108_2001_0, i_13_108_2047_0,
    i_13_108_2056_0, i_13_108_2150_0, i_13_108_2275_0, i_13_108_2280_0,
    i_13_108_2421_0, i_13_108_2424_0, i_13_108_2430_0, i_13_108_2497_0,
    i_13_108_2584_0, i_13_108_2712_0, i_13_108_2721_0, i_13_108_2722_0,
    i_13_108_2725_0, i_13_108_2784_0, i_13_108_2786_0, i_13_108_2856_0,
    i_13_108_2857_0, i_13_108_2859_0, i_13_108_2860_0, i_13_108_3010_0,
    i_13_108_3063_0, i_13_108_3064_0, i_13_108_3066_0, i_13_108_3097_0,
    i_13_108_3100_0, i_13_108_3103_0, i_13_108_3213_0, i_13_108_3234_0,
    i_13_108_3238_0, i_13_108_3255_0, i_13_108_3334_0, i_13_108_3428_0,
    i_13_108_3442_0, i_13_108_3487_0, i_13_108_3541_0, i_13_108_3554_0,
    i_13_108_3684_0, i_13_108_3691_0, i_13_108_3702_0, i_13_108_3717_0,
    i_13_108_3865_0, i_13_108_3871_0, i_13_108_3931_0, i_13_108_3977_0,
    i_13_108_4020_0, i_13_108_4252_0, i_13_108_4270_0, i_13_108_4328_0,
    i_13_108_4337_0, i_13_108_4350_0, i_13_108_4351_0, i_13_108_4395_0,
    i_13_108_4398_0, i_13_108_4413_0, i_13_108_4517_0, i_13_108_4593_0;
  output o_13_108_0_0;
  assign o_13_108_0_0 = ~((i_13_108_3487_0 & (~i_13_108_3234_0 | (~i_13_108_3063_0 & ~i_13_108_4351_0))) | (~i_13_108_3684_0 & ((~i_13_108_3931_0 & ~i_13_108_4351_0) | (~i_13_108_1605_0 & ~i_13_108_3066_0 & ~i_13_108_4413_0))) | (~i_13_108_382_0 & ~i_13_108_1620_0 & ~i_13_108_3238_0) | (~i_13_108_534_0 & ~i_13_108_2056_0 & ~i_13_108_4351_0 & ~i_13_108_4398_0));
endmodule



// Benchmark "kernel_13_109" written by ABC on Sun Jul 19 10:46:56 2020

module kernel_13_109 ( 
    i_13_109_118_0, i_13_109_127_0, i_13_109_181_0, i_13_109_182_0,
    i_13_109_260_0, i_13_109_280_0, i_13_109_281_0, i_13_109_283_0,
    i_13_109_325_0, i_13_109_355_0, i_13_109_535_0, i_13_109_569_0,
    i_13_109_596_0, i_13_109_598_0, i_13_109_599_0, i_13_109_667_0,
    i_13_109_697_0, i_13_109_712_0, i_13_109_728_0, i_13_109_742_0,
    i_13_109_745_0, i_13_109_778_0, i_13_109_821_0, i_13_109_847_0,
    i_13_109_853_0, i_13_109_856_0, i_13_109_863_0, i_13_109_898_0,
    i_13_109_946_0, i_13_109_986_0, i_13_109_1082_0, i_13_109_1094_0,
    i_13_109_1279_0, i_13_109_1280_0, i_13_109_1486_0, i_13_109_1487_0,
    i_13_109_1507_0, i_13_109_1669_0, i_13_109_1688_0, i_13_109_1724_0,
    i_13_109_1747_0, i_13_109_1751_0, i_13_109_1787_0, i_13_109_1808_0,
    i_13_109_1855_0, i_13_109_1856_0, i_13_109_1921_0, i_13_109_1940_0,
    i_13_109_1955_0, i_13_109_2056_0, i_13_109_2120_0, i_13_109_2146_0,
    i_13_109_2227_0, i_13_109_2305_0, i_13_109_2308_0, i_13_109_2314_0,
    i_13_109_2363_0, i_13_109_2425_0, i_13_109_2458_0, i_13_109_2459_0,
    i_13_109_2462_0, i_13_109_2467_0, i_13_109_2539_0, i_13_109_2540_0,
    i_13_109_2611_0, i_13_109_2612_0, i_13_109_2630_0, i_13_109_2765_0,
    i_13_109_2824_0, i_13_109_2882_0, i_13_109_2942_0, i_13_109_2981_0,
    i_13_109_3014_0, i_13_109_3020_0, i_13_109_3146_0, i_13_109_3148_0,
    i_13_109_3164_0, i_13_109_3169_0, i_13_109_3170_0, i_13_109_3173_0,
    i_13_109_3268_0, i_13_109_3290_0, i_13_109_3313_0, i_13_109_3370_0,
    i_13_109_3380_0, i_13_109_3425_0, i_13_109_3529_0, i_13_109_3782_0,
    i_13_109_3854_0, i_13_109_3871_0, i_13_109_3872_0, i_13_109_3875_0,
    i_13_109_3907_0, i_13_109_3908_0, i_13_109_3911_0, i_13_109_3941_0,
    i_13_109_4015_0, i_13_109_4261_0, i_13_109_4441_0, i_13_109_4519_0,
    o_13_109_0_0  );
  input  i_13_109_118_0, i_13_109_127_0, i_13_109_181_0, i_13_109_182_0,
    i_13_109_260_0, i_13_109_280_0, i_13_109_281_0, i_13_109_283_0,
    i_13_109_325_0, i_13_109_355_0, i_13_109_535_0, i_13_109_569_0,
    i_13_109_596_0, i_13_109_598_0, i_13_109_599_0, i_13_109_667_0,
    i_13_109_697_0, i_13_109_712_0, i_13_109_728_0, i_13_109_742_0,
    i_13_109_745_0, i_13_109_778_0, i_13_109_821_0, i_13_109_847_0,
    i_13_109_853_0, i_13_109_856_0, i_13_109_863_0, i_13_109_898_0,
    i_13_109_946_0, i_13_109_986_0, i_13_109_1082_0, i_13_109_1094_0,
    i_13_109_1279_0, i_13_109_1280_0, i_13_109_1486_0, i_13_109_1487_0,
    i_13_109_1507_0, i_13_109_1669_0, i_13_109_1688_0, i_13_109_1724_0,
    i_13_109_1747_0, i_13_109_1751_0, i_13_109_1787_0, i_13_109_1808_0,
    i_13_109_1855_0, i_13_109_1856_0, i_13_109_1921_0, i_13_109_1940_0,
    i_13_109_1955_0, i_13_109_2056_0, i_13_109_2120_0, i_13_109_2146_0,
    i_13_109_2227_0, i_13_109_2305_0, i_13_109_2308_0, i_13_109_2314_0,
    i_13_109_2363_0, i_13_109_2425_0, i_13_109_2458_0, i_13_109_2459_0,
    i_13_109_2462_0, i_13_109_2467_0, i_13_109_2539_0, i_13_109_2540_0,
    i_13_109_2611_0, i_13_109_2612_0, i_13_109_2630_0, i_13_109_2765_0,
    i_13_109_2824_0, i_13_109_2882_0, i_13_109_2942_0, i_13_109_2981_0,
    i_13_109_3014_0, i_13_109_3020_0, i_13_109_3146_0, i_13_109_3148_0,
    i_13_109_3164_0, i_13_109_3169_0, i_13_109_3170_0, i_13_109_3173_0,
    i_13_109_3268_0, i_13_109_3290_0, i_13_109_3313_0, i_13_109_3370_0,
    i_13_109_3380_0, i_13_109_3425_0, i_13_109_3529_0, i_13_109_3782_0,
    i_13_109_3854_0, i_13_109_3871_0, i_13_109_3872_0, i_13_109_3875_0,
    i_13_109_3907_0, i_13_109_3908_0, i_13_109_3911_0, i_13_109_3941_0,
    i_13_109_4015_0, i_13_109_4261_0, i_13_109_4441_0, i_13_109_4519_0;
  output o_13_109_0_0;
  assign o_13_109_0_0 = ~((~i_13_109_1856_0 & (~i_13_109_1486_0 | (~i_13_109_1487_0 & ~i_13_109_1747_0))) | (~i_13_109_1955_0 & ((i_13_109_667_0 & i_13_109_2146_0) | (~i_13_109_3164_0 & i_13_109_3911_0))) | (~i_13_109_2458_0 & ~i_13_109_3782_0) | (~i_13_109_3170_0 & ~i_13_109_3871_0 & ~i_13_109_3911_0));
endmodule



// Benchmark "kernel_13_110" written by ABC on Sun Jul 19 10:46:57 2020

module kernel_13_110 ( 
    i_13_110_31_0, i_13_110_34_0, i_13_110_35_0, i_13_110_39_0,
    i_13_110_64_0, i_13_110_67_0, i_13_110_122_0, i_13_110_134_0,
    i_13_110_161_0, i_13_110_225_0, i_13_110_232_0, i_13_110_233_0,
    i_13_110_272_0, i_13_110_306_0, i_13_110_386_0, i_13_110_449_0,
    i_13_110_490_0, i_13_110_493_0, i_13_110_538_0, i_13_110_607_0,
    i_13_110_612_0, i_13_110_648_0, i_13_110_746_0, i_13_110_759_0,
    i_13_110_762_0, i_13_110_763_0, i_13_110_764_0, i_13_110_868_0,
    i_13_110_1078_0, i_13_110_1128_0, i_13_110_1132_0, i_13_110_1186_0,
    i_13_110_1230_0, i_13_110_1303_0, i_13_110_1349_0, i_13_110_1444_0,
    i_13_110_1445_0, i_13_110_1447_0, i_13_110_1609_0, i_13_110_1700_0,
    i_13_110_1723_0, i_13_110_1724_0, i_13_110_1799_0, i_13_110_1817_0,
    i_13_110_1844_0, i_13_110_1912_0, i_13_110_1934_0, i_13_110_2142_0,
    i_13_110_2177_0, i_13_110_2194_0, i_13_110_2240_0, i_13_110_2318_0,
    i_13_110_2399_0, i_13_110_2430_0, i_13_110_2560_0, i_13_110_2681_0,
    i_13_110_2721_0, i_13_110_2722_0, i_13_110_2723_0, i_13_110_2726_0,
    i_13_110_2762_0, i_13_110_2825_0, i_13_110_2856_0, i_13_110_2860_0,
    i_13_110_2861_0, i_13_110_3002_0, i_13_110_3037_0, i_13_110_3130_0,
    i_13_110_3139_0, i_13_110_3213_0, i_13_110_3233_0, i_13_110_3366_0,
    i_13_110_3392_0, i_13_110_3415_0, i_13_110_3418_0, i_13_110_3438_0,
    i_13_110_3443_0, i_13_110_3618_0, i_13_110_3636_0, i_13_110_3637_0,
    i_13_110_3641_0, i_13_110_3650_0, i_13_110_3683_0, i_13_110_3686_0,
    i_13_110_3719_0, i_13_110_3725_0, i_13_110_3731_0, i_13_110_3843_0,
    i_13_110_3847_0, i_13_110_3848_0, i_13_110_3892_0, i_13_110_3991_0,
    i_13_110_4039_0, i_13_110_4040_0, i_13_110_4054_0, i_13_110_4237_0,
    i_13_110_4273_0, i_13_110_4347_0, i_13_110_4399_0, i_13_110_4400_0,
    o_13_110_0_0  );
  input  i_13_110_31_0, i_13_110_34_0, i_13_110_35_0, i_13_110_39_0,
    i_13_110_64_0, i_13_110_67_0, i_13_110_122_0, i_13_110_134_0,
    i_13_110_161_0, i_13_110_225_0, i_13_110_232_0, i_13_110_233_0,
    i_13_110_272_0, i_13_110_306_0, i_13_110_386_0, i_13_110_449_0,
    i_13_110_490_0, i_13_110_493_0, i_13_110_538_0, i_13_110_607_0,
    i_13_110_612_0, i_13_110_648_0, i_13_110_746_0, i_13_110_759_0,
    i_13_110_762_0, i_13_110_763_0, i_13_110_764_0, i_13_110_868_0,
    i_13_110_1078_0, i_13_110_1128_0, i_13_110_1132_0, i_13_110_1186_0,
    i_13_110_1230_0, i_13_110_1303_0, i_13_110_1349_0, i_13_110_1444_0,
    i_13_110_1445_0, i_13_110_1447_0, i_13_110_1609_0, i_13_110_1700_0,
    i_13_110_1723_0, i_13_110_1724_0, i_13_110_1799_0, i_13_110_1817_0,
    i_13_110_1844_0, i_13_110_1912_0, i_13_110_1934_0, i_13_110_2142_0,
    i_13_110_2177_0, i_13_110_2194_0, i_13_110_2240_0, i_13_110_2318_0,
    i_13_110_2399_0, i_13_110_2430_0, i_13_110_2560_0, i_13_110_2681_0,
    i_13_110_2721_0, i_13_110_2722_0, i_13_110_2723_0, i_13_110_2726_0,
    i_13_110_2762_0, i_13_110_2825_0, i_13_110_2856_0, i_13_110_2860_0,
    i_13_110_2861_0, i_13_110_3002_0, i_13_110_3037_0, i_13_110_3130_0,
    i_13_110_3139_0, i_13_110_3213_0, i_13_110_3233_0, i_13_110_3366_0,
    i_13_110_3392_0, i_13_110_3415_0, i_13_110_3418_0, i_13_110_3438_0,
    i_13_110_3443_0, i_13_110_3618_0, i_13_110_3636_0, i_13_110_3637_0,
    i_13_110_3641_0, i_13_110_3650_0, i_13_110_3683_0, i_13_110_3686_0,
    i_13_110_3719_0, i_13_110_3725_0, i_13_110_3731_0, i_13_110_3843_0,
    i_13_110_3847_0, i_13_110_3848_0, i_13_110_3892_0, i_13_110_3991_0,
    i_13_110_4039_0, i_13_110_4040_0, i_13_110_4054_0, i_13_110_4237_0,
    i_13_110_4273_0, i_13_110_4347_0, i_13_110_4399_0, i_13_110_4400_0;
  output o_13_110_0_0;
  assign o_13_110_0_0 = ~((~i_13_110_449_0 & ~i_13_110_4273_0) | (~i_13_110_35_0 & ~i_13_110_67_0) | (~i_13_110_2681_0 & ~i_13_110_3443_0 & ~i_13_110_3686_0 & ~i_13_110_3731_0));
endmodule



// Benchmark "kernel_13_111" written by ABC on Sun Jul 19 10:46:58 2020

module kernel_13_111 ( 
    i_13_111_38_0, i_13_111_103_0, i_13_111_112_0, i_13_111_185_0,
    i_13_111_280_0, i_13_111_281_0, i_13_111_284_0, i_13_111_320_0,
    i_13_111_338_0, i_13_111_373_0, i_13_111_376_0, i_13_111_454_0,
    i_13_111_533_0, i_13_111_571_0, i_13_111_590_0, i_13_111_596_0,
    i_13_111_598_0, i_13_111_599_0, i_13_111_641_0, i_13_111_677_0,
    i_13_111_685_0, i_13_111_686_0, i_13_111_715_0, i_13_111_761_0,
    i_13_111_814_0, i_13_111_815_0, i_13_111_820_0, i_13_111_821_0,
    i_13_111_832_0, i_13_111_896_0, i_13_111_1067_0, i_13_111_1076_0,
    i_13_111_1084_0, i_13_111_1129_0, i_13_111_1381_0, i_13_111_1438_0,
    i_13_111_1694_0, i_13_111_1714_0, i_13_111_1747_0, i_13_111_1748_0,
    i_13_111_1814_0, i_13_111_1856_0, i_13_111_1859_0, i_13_111_1909_0,
    i_13_111_1991_0, i_13_111_2138_0, i_13_111_2308_0, i_13_111_2366_0,
    i_13_111_2407_0, i_13_111_2458_0, i_13_111_2459_0, i_13_111_2461_0,
    i_13_111_2479_0, i_13_111_2506_0, i_13_111_2615_0, i_13_111_2633_0,
    i_13_111_2647_0, i_13_111_2650_0, i_13_111_2651_0, i_13_111_2722_0,
    i_13_111_2732_0, i_13_111_2749_0, i_13_111_2876_0, i_13_111_2938_0,
    i_13_111_2981_0, i_13_111_3142_0, i_13_111_3169_0, i_13_111_3206_0,
    i_13_111_3290_0, i_13_111_3376_0, i_13_111_3398_0, i_13_111_3415_0,
    i_13_111_3422_0, i_13_111_3524_0, i_13_111_3647_0, i_13_111_3692_0,
    i_13_111_3791_0, i_13_111_3844_0, i_13_111_3889_0, i_13_111_3890_0,
    i_13_111_3910_0, i_13_111_3911_0, i_13_111_3937_0, i_13_111_3989_0,
    i_13_111_3992_0, i_13_111_4015_0, i_13_111_4019_0, i_13_111_4036_0,
    i_13_111_4045_0, i_13_111_4052_0, i_13_111_4064_0, i_13_111_4078_0,
    i_13_111_4090_0, i_13_111_4097_0, i_13_111_4217_0, i_13_111_4259_0,
    i_13_111_4369_0, i_13_111_4559_0, i_13_111_4594_0, i_13_111_4603_0,
    o_13_111_0_0  );
  input  i_13_111_38_0, i_13_111_103_0, i_13_111_112_0, i_13_111_185_0,
    i_13_111_280_0, i_13_111_281_0, i_13_111_284_0, i_13_111_320_0,
    i_13_111_338_0, i_13_111_373_0, i_13_111_376_0, i_13_111_454_0,
    i_13_111_533_0, i_13_111_571_0, i_13_111_590_0, i_13_111_596_0,
    i_13_111_598_0, i_13_111_599_0, i_13_111_641_0, i_13_111_677_0,
    i_13_111_685_0, i_13_111_686_0, i_13_111_715_0, i_13_111_761_0,
    i_13_111_814_0, i_13_111_815_0, i_13_111_820_0, i_13_111_821_0,
    i_13_111_832_0, i_13_111_896_0, i_13_111_1067_0, i_13_111_1076_0,
    i_13_111_1084_0, i_13_111_1129_0, i_13_111_1381_0, i_13_111_1438_0,
    i_13_111_1694_0, i_13_111_1714_0, i_13_111_1747_0, i_13_111_1748_0,
    i_13_111_1814_0, i_13_111_1856_0, i_13_111_1859_0, i_13_111_1909_0,
    i_13_111_1991_0, i_13_111_2138_0, i_13_111_2308_0, i_13_111_2366_0,
    i_13_111_2407_0, i_13_111_2458_0, i_13_111_2459_0, i_13_111_2461_0,
    i_13_111_2479_0, i_13_111_2506_0, i_13_111_2615_0, i_13_111_2633_0,
    i_13_111_2647_0, i_13_111_2650_0, i_13_111_2651_0, i_13_111_2722_0,
    i_13_111_2732_0, i_13_111_2749_0, i_13_111_2876_0, i_13_111_2938_0,
    i_13_111_2981_0, i_13_111_3142_0, i_13_111_3169_0, i_13_111_3206_0,
    i_13_111_3290_0, i_13_111_3376_0, i_13_111_3398_0, i_13_111_3415_0,
    i_13_111_3422_0, i_13_111_3524_0, i_13_111_3647_0, i_13_111_3692_0,
    i_13_111_3791_0, i_13_111_3844_0, i_13_111_3889_0, i_13_111_3890_0,
    i_13_111_3910_0, i_13_111_3911_0, i_13_111_3937_0, i_13_111_3989_0,
    i_13_111_3992_0, i_13_111_4015_0, i_13_111_4019_0, i_13_111_4036_0,
    i_13_111_4045_0, i_13_111_4052_0, i_13_111_4064_0, i_13_111_4078_0,
    i_13_111_4090_0, i_13_111_4097_0, i_13_111_4217_0, i_13_111_4259_0,
    i_13_111_4369_0, i_13_111_4559_0, i_13_111_4594_0, i_13_111_4603_0;
  output o_13_111_0_0;
  assign o_13_111_0_0 = ~(~i_13_111_1859_0 | (~i_13_111_533_0 & ~i_13_111_677_0 & ~i_13_111_2647_0));
endmodule



// Benchmark "kernel_13_112" written by ABC on Sun Jul 19 10:46:59 2020

module kernel_13_112 ( 
    i_13_112_3_0, i_13_112_37_0, i_13_112_180_0, i_13_112_181_0,
    i_13_112_183_0, i_13_112_185_0, i_13_112_187_0, i_13_112_193_0,
    i_13_112_210_0, i_13_112_244_0, i_13_112_255_0, i_13_112_360_0,
    i_13_112_382_0, i_13_112_446_0, i_13_112_526_0, i_13_112_550_0,
    i_13_112_596_0, i_13_112_597_0, i_13_112_625_0, i_13_112_640_0,
    i_13_112_642_0, i_13_112_643_0, i_13_112_646_0, i_13_112_647_0,
    i_13_112_685_0, i_13_112_692_0, i_13_112_851_0, i_13_112_894_0,
    i_13_112_898_0, i_13_112_975_0, i_13_112_1021_0, i_13_112_1093_0,
    i_13_112_1119_0, i_13_112_1120_0, i_13_112_1124_0, i_13_112_1276_0,
    i_13_112_1277_0, i_13_112_1391_0, i_13_112_1394_0, i_13_112_1407_0,
    i_13_112_1408_0, i_13_112_1461_0, i_13_112_1479_0, i_13_112_1488_0,
    i_13_112_1516_0, i_13_112_1643_0, i_13_112_1646_0, i_13_112_1668_0,
    i_13_112_1673_0, i_13_112_1813_0, i_13_112_1871_0, i_13_112_1990_0,
    i_13_112_2002_0, i_13_112_2046_0, i_13_112_2231_0, i_13_112_2361_0,
    i_13_112_2442_0, i_13_112_2542_0, i_13_112_2570_0, i_13_112_2676_0,
    i_13_112_2696_0, i_13_112_2767_0, i_13_112_2848_0, i_13_112_2852_0,
    i_13_112_2874_0, i_13_112_2920_0, i_13_112_2923_0, i_13_112_3092_0,
    i_13_112_3200_0, i_13_112_3291_0, i_13_112_3352_0, i_13_112_3419_0,
    i_13_112_3519_0, i_13_112_3523_0, i_13_112_3532_0, i_13_112_3541_0,
    i_13_112_3622_0, i_13_112_3730_0, i_13_112_3796_0, i_13_112_3900_0,
    i_13_112_3909_0, i_13_112_3918_0, i_13_112_3927_0, i_13_112_3928_0,
    i_13_112_3931_0, i_13_112_3993_0, i_13_112_3995_0, i_13_112_4083_0,
    i_13_112_4186_0, i_13_112_4189_0, i_13_112_4190_0, i_13_112_4192_0,
    i_13_112_4270_0, i_13_112_4297_0, i_13_112_4298_0, i_13_112_4341_0,
    i_13_112_4417_0, i_13_112_4596_0, i_13_112_4598_0, i_13_112_4599_0,
    o_13_112_0_0  );
  input  i_13_112_3_0, i_13_112_37_0, i_13_112_180_0, i_13_112_181_0,
    i_13_112_183_0, i_13_112_185_0, i_13_112_187_0, i_13_112_193_0,
    i_13_112_210_0, i_13_112_244_0, i_13_112_255_0, i_13_112_360_0,
    i_13_112_382_0, i_13_112_446_0, i_13_112_526_0, i_13_112_550_0,
    i_13_112_596_0, i_13_112_597_0, i_13_112_625_0, i_13_112_640_0,
    i_13_112_642_0, i_13_112_643_0, i_13_112_646_0, i_13_112_647_0,
    i_13_112_685_0, i_13_112_692_0, i_13_112_851_0, i_13_112_894_0,
    i_13_112_898_0, i_13_112_975_0, i_13_112_1021_0, i_13_112_1093_0,
    i_13_112_1119_0, i_13_112_1120_0, i_13_112_1124_0, i_13_112_1276_0,
    i_13_112_1277_0, i_13_112_1391_0, i_13_112_1394_0, i_13_112_1407_0,
    i_13_112_1408_0, i_13_112_1461_0, i_13_112_1479_0, i_13_112_1488_0,
    i_13_112_1516_0, i_13_112_1643_0, i_13_112_1646_0, i_13_112_1668_0,
    i_13_112_1673_0, i_13_112_1813_0, i_13_112_1871_0, i_13_112_1990_0,
    i_13_112_2002_0, i_13_112_2046_0, i_13_112_2231_0, i_13_112_2361_0,
    i_13_112_2442_0, i_13_112_2542_0, i_13_112_2570_0, i_13_112_2676_0,
    i_13_112_2696_0, i_13_112_2767_0, i_13_112_2848_0, i_13_112_2852_0,
    i_13_112_2874_0, i_13_112_2920_0, i_13_112_2923_0, i_13_112_3092_0,
    i_13_112_3200_0, i_13_112_3291_0, i_13_112_3352_0, i_13_112_3419_0,
    i_13_112_3519_0, i_13_112_3523_0, i_13_112_3532_0, i_13_112_3541_0,
    i_13_112_3622_0, i_13_112_3730_0, i_13_112_3796_0, i_13_112_3900_0,
    i_13_112_3909_0, i_13_112_3918_0, i_13_112_3927_0, i_13_112_3928_0,
    i_13_112_3931_0, i_13_112_3993_0, i_13_112_3995_0, i_13_112_4083_0,
    i_13_112_4186_0, i_13_112_4189_0, i_13_112_4190_0, i_13_112_4192_0,
    i_13_112_4270_0, i_13_112_4297_0, i_13_112_4298_0, i_13_112_4341_0,
    i_13_112_4417_0, i_13_112_4596_0, i_13_112_4598_0, i_13_112_4599_0;
  output o_13_112_0_0;
  assign o_13_112_0_0 = ~((i_13_112_526_0 & ((~i_13_112_1120_0 & ((~i_13_112_898_0 & ~i_13_112_1643_0 & ~i_13_112_3993_0) | (i_13_112_3541_0 & i_13_112_4186_0))) | (i_13_112_185_0 & i_13_112_1813_0 & i_13_112_4186_0))) | (i_13_112_2002_0 & ((i_13_112_244_0 & ~i_13_112_446_0 & ~i_13_112_2874_0 & ~i_13_112_3928_0) | (~i_13_112_1276_0 & ~i_13_112_2848_0 & ~i_13_112_3927_0 & ~i_13_112_3995_0))) | (~i_13_112_187_0 & ~i_13_112_685_0 & ~i_13_112_692_0 & ~i_13_112_3900_0 & ~i_13_112_3931_0 & ~i_13_112_4189_0) | (~i_13_112_1408_0 & ~i_13_112_1479_0 & i_13_112_2920_0 & ~i_13_112_4190_0) | (~i_13_112_2874_0 & i_13_112_3532_0 & ~i_13_112_3622_0 & ~i_13_112_4186_0 & i_13_112_4270_0));
endmodule



// Benchmark "kernel_13_113" written by ABC on Sun Jul 19 10:46:59 2020

module kernel_13_113 ( 
    i_13_113_26_0, i_13_113_52_0, i_13_113_167_0, i_13_113_170_0,
    i_13_113_248_0, i_13_113_263_0, i_13_113_278_0, i_13_113_320_0,
    i_13_113_340_0, i_13_113_376_0, i_13_113_452_0, i_13_113_454_0,
    i_13_113_460_0, i_13_113_607_0, i_13_113_732_0, i_13_113_811_0,
    i_13_113_815_0, i_13_113_1078_0, i_13_113_1079_0, i_13_113_1217_0,
    i_13_113_1304_0, i_13_113_1313_0, i_13_113_1343_0, i_13_113_1346_0,
    i_13_113_1402_0, i_13_113_1403_0, i_13_113_1408_0, i_13_113_1468_0,
    i_13_113_1529_0, i_13_113_1781_0, i_13_113_1805_0, i_13_113_1814_0,
    i_13_113_1835_0, i_13_113_1851_0, i_13_113_1852_0, i_13_113_1853_0,
    i_13_113_1912_0, i_13_113_1957_0, i_13_113_2006_0, i_13_113_2111_0,
    i_13_113_2128_0, i_13_113_2150_0, i_13_113_2174_0, i_13_113_2201_0,
    i_13_113_2234_0, i_13_113_2278_0, i_13_113_2279_0, i_13_113_2303_0,
    i_13_113_2318_0, i_13_113_2453_0, i_13_113_2618_0, i_13_113_2746_0,
    i_13_113_2765_0, i_13_113_2767_0, i_13_113_2788_0, i_13_113_2789_0,
    i_13_113_2848_0, i_13_113_2858_0, i_13_113_2872_0, i_13_113_3001_0,
    i_13_113_3002_0, i_13_113_3020_0, i_13_113_3091_0, i_13_113_3124_0,
    i_13_113_3131_0, i_13_113_3154_0, i_13_113_3215_0, i_13_113_3218_0,
    i_13_113_3232_0, i_13_113_3238_0, i_13_113_3305_0, i_13_113_3371_0,
    i_13_113_3442_0, i_13_113_3464_0, i_13_113_3505_0, i_13_113_3532_0,
    i_13_113_3545_0, i_13_113_3613_0, i_13_113_3616_0, i_13_113_3644_0,
    i_13_113_3689_0, i_13_113_3706_0, i_13_113_3712_0, i_13_113_3739_0,
    i_13_113_3892_0, i_13_113_3904_0, i_13_113_3961_0, i_13_113_4063_0,
    i_13_113_4231_0, i_13_113_4268_0, i_13_113_4271_0, i_13_113_4316_0,
    i_13_113_4367_0, i_13_113_4384_0, i_13_113_4393_0, i_13_113_4413_0,
    i_13_113_4450_0, i_13_113_4523_0, i_13_113_4532_0, i_13_113_4595_0,
    o_13_113_0_0  );
  input  i_13_113_26_0, i_13_113_52_0, i_13_113_167_0, i_13_113_170_0,
    i_13_113_248_0, i_13_113_263_0, i_13_113_278_0, i_13_113_320_0,
    i_13_113_340_0, i_13_113_376_0, i_13_113_452_0, i_13_113_454_0,
    i_13_113_460_0, i_13_113_607_0, i_13_113_732_0, i_13_113_811_0,
    i_13_113_815_0, i_13_113_1078_0, i_13_113_1079_0, i_13_113_1217_0,
    i_13_113_1304_0, i_13_113_1313_0, i_13_113_1343_0, i_13_113_1346_0,
    i_13_113_1402_0, i_13_113_1403_0, i_13_113_1408_0, i_13_113_1468_0,
    i_13_113_1529_0, i_13_113_1781_0, i_13_113_1805_0, i_13_113_1814_0,
    i_13_113_1835_0, i_13_113_1851_0, i_13_113_1852_0, i_13_113_1853_0,
    i_13_113_1912_0, i_13_113_1957_0, i_13_113_2006_0, i_13_113_2111_0,
    i_13_113_2128_0, i_13_113_2150_0, i_13_113_2174_0, i_13_113_2201_0,
    i_13_113_2234_0, i_13_113_2278_0, i_13_113_2279_0, i_13_113_2303_0,
    i_13_113_2318_0, i_13_113_2453_0, i_13_113_2618_0, i_13_113_2746_0,
    i_13_113_2765_0, i_13_113_2767_0, i_13_113_2788_0, i_13_113_2789_0,
    i_13_113_2848_0, i_13_113_2858_0, i_13_113_2872_0, i_13_113_3001_0,
    i_13_113_3002_0, i_13_113_3020_0, i_13_113_3091_0, i_13_113_3124_0,
    i_13_113_3131_0, i_13_113_3154_0, i_13_113_3215_0, i_13_113_3218_0,
    i_13_113_3232_0, i_13_113_3238_0, i_13_113_3305_0, i_13_113_3371_0,
    i_13_113_3442_0, i_13_113_3464_0, i_13_113_3505_0, i_13_113_3532_0,
    i_13_113_3545_0, i_13_113_3613_0, i_13_113_3616_0, i_13_113_3644_0,
    i_13_113_3689_0, i_13_113_3706_0, i_13_113_3712_0, i_13_113_3739_0,
    i_13_113_3892_0, i_13_113_3904_0, i_13_113_3961_0, i_13_113_4063_0,
    i_13_113_4231_0, i_13_113_4268_0, i_13_113_4271_0, i_13_113_4316_0,
    i_13_113_4367_0, i_13_113_4384_0, i_13_113_4393_0, i_13_113_4413_0,
    i_13_113_4450_0, i_13_113_4523_0, i_13_113_4532_0, i_13_113_4595_0;
  output o_13_113_0_0;
  assign o_13_113_0_0 = ~(~i_13_113_3238_0 | ~i_13_113_3442_0 | i_13_113_3091_0 | ~i_13_113_1529_0 | ~i_13_113_1853_0);
endmodule



// Benchmark "kernel_13_114" written by ABC on Sun Jul 19 10:47:00 2020

module kernel_13_114 ( 
    i_13_114_67_0, i_13_114_68_0, i_13_114_76_0, i_13_114_100_0,
    i_13_114_115_0, i_13_114_121_0, i_13_114_135_0, i_13_114_136_0,
    i_13_114_372_0, i_13_114_550_0, i_13_114_553_0, i_13_114_587_0,
    i_13_114_598_0, i_13_114_604_0, i_13_114_625_0, i_13_114_643_0,
    i_13_114_658_0, i_13_114_667_0, i_13_114_679_0, i_13_114_685_0,
    i_13_114_694_0, i_13_114_703_0, i_13_114_711_0, i_13_114_760_0,
    i_13_114_819_0, i_13_114_825_0, i_13_114_1116_0, i_13_114_1117_0,
    i_13_114_1153_0, i_13_114_1206_0, i_13_114_1207_0, i_13_114_1211_0,
    i_13_114_1273_0, i_13_114_1314_0, i_13_114_1390_0, i_13_114_1440_0,
    i_13_114_1507_0, i_13_114_1660_0, i_13_114_1668_0, i_13_114_1725_0,
    i_13_114_1729_0, i_13_114_1732_0, i_13_114_1735_0, i_13_114_1742_0,
    i_13_114_1774_0, i_13_114_1795_0, i_13_114_1796_0, i_13_114_1831_0,
    i_13_114_1944_0, i_13_114_1945_0, i_13_114_1999_0, i_13_114_2115_0,
    i_13_114_2201_0, i_13_114_2377_0, i_13_114_2380_0, i_13_114_2381_0,
    i_13_114_2422_0, i_13_114_2461_0, i_13_114_2548_0, i_13_114_2584_0,
    i_13_114_2646_0, i_13_114_2676_0, i_13_114_2718_0, i_13_114_2749_0,
    i_13_114_2847_0, i_13_114_2848_0, i_13_114_2881_0, i_13_114_2962_0,
    i_13_114_3090_0, i_13_114_3092_0, i_13_114_3094_0, i_13_114_3153_0,
    i_13_114_3352_0, i_13_114_3367_0, i_13_114_3414_0, i_13_114_3445_0,
    i_13_114_3637_0, i_13_114_3649_0, i_13_114_3865_0, i_13_114_3892_0,
    i_13_114_3893_0, i_13_114_3910_0, i_13_114_3927_0, i_13_114_3928_0,
    i_13_114_3990_0, i_13_114_4060_0, i_13_114_4063_0, i_13_114_4186_0,
    i_13_114_4192_0, i_13_114_4216_0, i_13_114_4293_0, i_13_114_4295_0,
    i_13_114_4297_0, i_13_114_4303_0, i_13_114_4305_0, i_13_114_4329_0,
    i_13_114_4432_0, i_13_114_4447_0, i_13_114_4558_0, i_13_114_4593_0,
    o_13_114_0_0  );
  input  i_13_114_67_0, i_13_114_68_0, i_13_114_76_0, i_13_114_100_0,
    i_13_114_115_0, i_13_114_121_0, i_13_114_135_0, i_13_114_136_0,
    i_13_114_372_0, i_13_114_550_0, i_13_114_553_0, i_13_114_587_0,
    i_13_114_598_0, i_13_114_604_0, i_13_114_625_0, i_13_114_643_0,
    i_13_114_658_0, i_13_114_667_0, i_13_114_679_0, i_13_114_685_0,
    i_13_114_694_0, i_13_114_703_0, i_13_114_711_0, i_13_114_760_0,
    i_13_114_819_0, i_13_114_825_0, i_13_114_1116_0, i_13_114_1117_0,
    i_13_114_1153_0, i_13_114_1206_0, i_13_114_1207_0, i_13_114_1211_0,
    i_13_114_1273_0, i_13_114_1314_0, i_13_114_1390_0, i_13_114_1440_0,
    i_13_114_1507_0, i_13_114_1660_0, i_13_114_1668_0, i_13_114_1725_0,
    i_13_114_1729_0, i_13_114_1732_0, i_13_114_1735_0, i_13_114_1742_0,
    i_13_114_1774_0, i_13_114_1795_0, i_13_114_1796_0, i_13_114_1831_0,
    i_13_114_1944_0, i_13_114_1945_0, i_13_114_1999_0, i_13_114_2115_0,
    i_13_114_2201_0, i_13_114_2377_0, i_13_114_2380_0, i_13_114_2381_0,
    i_13_114_2422_0, i_13_114_2461_0, i_13_114_2548_0, i_13_114_2584_0,
    i_13_114_2646_0, i_13_114_2676_0, i_13_114_2718_0, i_13_114_2749_0,
    i_13_114_2847_0, i_13_114_2848_0, i_13_114_2881_0, i_13_114_2962_0,
    i_13_114_3090_0, i_13_114_3092_0, i_13_114_3094_0, i_13_114_3153_0,
    i_13_114_3352_0, i_13_114_3367_0, i_13_114_3414_0, i_13_114_3445_0,
    i_13_114_3637_0, i_13_114_3649_0, i_13_114_3865_0, i_13_114_3892_0,
    i_13_114_3893_0, i_13_114_3910_0, i_13_114_3927_0, i_13_114_3928_0,
    i_13_114_3990_0, i_13_114_4060_0, i_13_114_4063_0, i_13_114_4186_0,
    i_13_114_4192_0, i_13_114_4216_0, i_13_114_4293_0, i_13_114_4295_0,
    i_13_114_4297_0, i_13_114_4303_0, i_13_114_4305_0, i_13_114_4329_0,
    i_13_114_4432_0, i_13_114_4447_0, i_13_114_4558_0, i_13_114_4593_0;
  output o_13_114_0_0;
  assign o_13_114_0_0 = ~((~i_13_114_1314_0 & ((i_13_114_760_0 & ~i_13_114_2380_0) | (~i_13_114_667_0 & ~i_13_114_1211_0 & ~i_13_114_2646_0 & ~i_13_114_3649_0))) | (~i_13_114_1729_0 & ((i_13_114_1116_0 & i_13_114_2676_0 & ~i_13_114_3892_0) | (~i_13_114_1206_0 & ~i_13_114_3865_0 & ~i_13_114_4432_0))) | (~i_13_114_4329_0 & ((~i_13_114_685_0 & ~i_13_114_2847_0) | (~i_13_114_1507_0 & ~i_13_114_3927_0))) | (~i_13_114_2676_0 & ~i_13_114_3649_0 & ~i_13_114_3910_0 & ~i_13_114_4303_0));
endmodule



// Benchmark "kernel_13_115" written by ABC on Sun Jul 19 10:47:01 2020

module kernel_13_115 ( 
    i_13_115_45_0, i_13_115_50_0, i_13_115_174_0, i_13_115_251_0,
    i_13_115_279_0, i_13_115_280_0, i_13_115_282_0, i_13_115_285_0,
    i_13_115_286_0, i_13_115_373_0, i_13_115_516_0, i_13_115_531_0,
    i_13_115_665_0, i_13_115_670_0, i_13_115_688_0, i_13_115_762_0,
    i_13_115_769_0, i_13_115_851_0, i_13_115_1020_0, i_13_115_1021_0,
    i_13_115_1024_0, i_13_115_1071_0, i_13_115_1272_0, i_13_115_1273_0,
    i_13_115_1425_0, i_13_115_1529_0, i_13_115_1601_0, i_13_115_1632_0,
    i_13_115_1633_0, i_13_115_1635_0, i_13_115_1636_0, i_13_115_1637_0,
    i_13_115_1693_0, i_13_115_1780_0, i_13_115_1932_0, i_13_115_2001_0,
    i_13_115_2034_0, i_13_115_2352_0, i_13_115_2380_0, i_13_115_2448_0,
    i_13_115_2449_0, i_13_115_2454_0, i_13_115_2455_0, i_13_115_2461_0,
    i_13_115_2464_0, i_13_115_2475_0, i_13_115_2545_0, i_13_115_2617_0,
    i_13_115_2641_0, i_13_115_2677_0, i_13_115_2762_0, i_13_115_2839_0,
    i_13_115_2844_0, i_13_115_2961_0, i_13_115_3105_0, i_13_115_3118_0,
    i_13_115_3129_0, i_13_115_3167_0, i_13_115_3198_0, i_13_115_3417_0,
    i_13_115_3421_0, i_13_115_3424_0, i_13_115_3447_0, i_13_115_3450_0,
    i_13_115_3460_0, i_13_115_3535_0, i_13_115_3612_0, i_13_115_3727_0,
    i_13_115_3729_0, i_13_115_3730_0, i_13_115_3731_0, i_13_115_3733_0,
    i_13_115_3793_0, i_13_115_3838_0, i_13_115_3909_0, i_13_115_3913_0,
    i_13_115_4014_0, i_13_115_4017_0, i_13_115_4018_0, i_13_115_4248_0,
    i_13_115_4251_0, i_13_115_4252_0, i_13_115_4253_0, i_13_115_4255_0,
    i_13_115_4256_0, i_13_115_4258_0, i_13_115_4260_0, i_13_115_4350_0,
    i_13_115_4407_0, i_13_115_4461_0, i_13_115_4513_0, i_13_115_4524_0,
    i_13_115_4554_0, i_13_115_4555_0, i_13_115_4557_0, i_13_115_4558_0,
    i_13_115_4560_0, i_13_115_4561_0, i_13_115_4562_0, i_13_115_4579_0,
    o_13_115_0_0  );
  input  i_13_115_45_0, i_13_115_50_0, i_13_115_174_0, i_13_115_251_0,
    i_13_115_279_0, i_13_115_280_0, i_13_115_282_0, i_13_115_285_0,
    i_13_115_286_0, i_13_115_373_0, i_13_115_516_0, i_13_115_531_0,
    i_13_115_665_0, i_13_115_670_0, i_13_115_688_0, i_13_115_762_0,
    i_13_115_769_0, i_13_115_851_0, i_13_115_1020_0, i_13_115_1021_0,
    i_13_115_1024_0, i_13_115_1071_0, i_13_115_1272_0, i_13_115_1273_0,
    i_13_115_1425_0, i_13_115_1529_0, i_13_115_1601_0, i_13_115_1632_0,
    i_13_115_1633_0, i_13_115_1635_0, i_13_115_1636_0, i_13_115_1637_0,
    i_13_115_1693_0, i_13_115_1780_0, i_13_115_1932_0, i_13_115_2001_0,
    i_13_115_2034_0, i_13_115_2352_0, i_13_115_2380_0, i_13_115_2448_0,
    i_13_115_2449_0, i_13_115_2454_0, i_13_115_2455_0, i_13_115_2461_0,
    i_13_115_2464_0, i_13_115_2475_0, i_13_115_2545_0, i_13_115_2617_0,
    i_13_115_2641_0, i_13_115_2677_0, i_13_115_2762_0, i_13_115_2839_0,
    i_13_115_2844_0, i_13_115_2961_0, i_13_115_3105_0, i_13_115_3118_0,
    i_13_115_3129_0, i_13_115_3167_0, i_13_115_3198_0, i_13_115_3417_0,
    i_13_115_3421_0, i_13_115_3424_0, i_13_115_3447_0, i_13_115_3450_0,
    i_13_115_3460_0, i_13_115_3535_0, i_13_115_3612_0, i_13_115_3727_0,
    i_13_115_3729_0, i_13_115_3730_0, i_13_115_3731_0, i_13_115_3733_0,
    i_13_115_3793_0, i_13_115_3838_0, i_13_115_3909_0, i_13_115_3913_0,
    i_13_115_4014_0, i_13_115_4017_0, i_13_115_4018_0, i_13_115_4248_0,
    i_13_115_4251_0, i_13_115_4252_0, i_13_115_4253_0, i_13_115_4255_0,
    i_13_115_4256_0, i_13_115_4258_0, i_13_115_4260_0, i_13_115_4350_0,
    i_13_115_4407_0, i_13_115_4461_0, i_13_115_4513_0, i_13_115_4524_0,
    i_13_115_4554_0, i_13_115_4555_0, i_13_115_4557_0, i_13_115_4558_0,
    i_13_115_4560_0, i_13_115_4561_0, i_13_115_4562_0, i_13_115_4579_0;
  output o_13_115_0_0;
  assign o_13_115_0_0 = ~((~i_13_115_3733_0 & ((~i_13_115_282_0 & i_13_115_1273_0) | (i_13_115_174_0 & ~i_13_115_531_0 & ~i_13_115_2464_0 & ~i_13_115_4555_0))) | (i_13_115_3421_0 & ~i_13_115_3909_0) | (~i_13_115_1020_0 & ~i_13_115_2454_0 & ~i_13_115_4248_0 & ~i_13_115_4260_0));
endmodule



// Benchmark "kernel_13_116" written by ABC on Sun Jul 19 10:47:02 2020

module kernel_13_116 ( 
    i_13_116_56_0, i_13_116_128_0, i_13_116_139_0, i_13_116_168_0,
    i_13_116_173_0, i_13_116_175_0, i_13_116_176_0, i_13_116_193_0,
    i_13_116_317_0, i_13_116_355_0, i_13_116_418_0, i_13_116_420_0,
    i_13_116_454_0, i_13_116_515_0, i_13_116_571_0, i_13_116_572_0,
    i_13_116_608_0, i_13_116_647_0, i_13_116_812_0, i_13_116_947_0,
    i_13_116_959_0, i_13_116_986_0, i_13_116_988_0, i_13_116_1216_0,
    i_13_116_1300_0, i_13_116_1345_0, i_13_116_1399_0, i_13_116_1405_0,
    i_13_116_1410_0, i_13_116_1453_0, i_13_116_1516_0, i_13_116_1552_0,
    i_13_116_1602_0, i_13_116_1714_0, i_13_116_1765_0, i_13_116_1767_0,
    i_13_116_1777_0, i_13_116_1793_0, i_13_116_1804_0, i_13_116_1828_0,
    i_13_116_1829_0, i_13_116_1831_0, i_13_116_1833_0, i_13_116_1885_0,
    i_13_116_2018_0, i_13_116_2019_0, i_13_116_2108_0, i_13_116_2146_0,
    i_13_116_2300_0, i_13_116_2335_0, i_13_116_2408_0, i_13_116_2470_0,
    i_13_116_2472_0, i_13_116_2474_0, i_13_116_2697_0, i_13_116_2705_0,
    i_13_116_2713_0, i_13_116_2746_0, i_13_116_2857_0, i_13_116_2858_0,
    i_13_116_2952_0, i_13_116_2980_0, i_13_116_2981_0, i_13_116_2982_0,
    i_13_116_2983_0, i_13_116_2985_0, i_13_116_3007_0, i_13_116_3027_0,
    i_13_116_3110_0, i_13_116_3154_0, i_13_116_3160_0, i_13_116_3211_0,
    i_13_116_3233_0, i_13_116_3386_0, i_13_116_3451_0, i_13_116_3549_0,
    i_13_116_3619_0, i_13_116_3710_0, i_13_116_3739_0, i_13_116_3763_0,
    i_13_116_3782_0, i_13_116_3817_0, i_13_116_3818_0, i_13_116_3872_0,
    i_13_116_4018_0, i_13_116_4054_0, i_13_116_4079_0, i_13_116_4084_0,
    i_13_116_4198_0, i_13_116_4258_0, i_13_116_4259_0, i_13_116_4376_0,
    i_13_116_4396_0, i_13_116_4511_0, i_13_116_4513_0, i_13_116_4522_0,
    i_13_116_4564_0, i_13_116_4565_0, i_13_116_4567_0, i_13_116_4570_0,
    o_13_116_0_0  );
  input  i_13_116_56_0, i_13_116_128_0, i_13_116_139_0, i_13_116_168_0,
    i_13_116_173_0, i_13_116_175_0, i_13_116_176_0, i_13_116_193_0,
    i_13_116_317_0, i_13_116_355_0, i_13_116_418_0, i_13_116_420_0,
    i_13_116_454_0, i_13_116_515_0, i_13_116_571_0, i_13_116_572_0,
    i_13_116_608_0, i_13_116_647_0, i_13_116_812_0, i_13_116_947_0,
    i_13_116_959_0, i_13_116_986_0, i_13_116_988_0, i_13_116_1216_0,
    i_13_116_1300_0, i_13_116_1345_0, i_13_116_1399_0, i_13_116_1405_0,
    i_13_116_1410_0, i_13_116_1453_0, i_13_116_1516_0, i_13_116_1552_0,
    i_13_116_1602_0, i_13_116_1714_0, i_13_116_1765_0, i_13_116_1767_0,
    i_13_116_1777_0, i_13_116_1793_0, i_13_116_1804_0, i_13_116_1828_0,
    i_13_116_1829_0, i_13_116_1831_0, i_13_116_1833_0, i_13_116_1885_0,
    i_13_116_2018_0, i_13_116_2019_0, i_13_116_2108_0, i_13_116_2146_0,
    i_13_116_2300_0, i_13_116_2335_0, i_13_116_2408_0, i_13_116_2470_0,
    i_13_116_2472_0, i_13_116_2474_0, i_13_116_2697_0, i_13_116_2705_0,
    i_13_116_2713_0, i_13_116_2746_0, i_13_116_2857_0, i_13_116_2858_0,
    i_13_116_2952_0, i_13_116_2980_0, i_13_116_2981_0, i_13_116_2982_0,
    i_13_116_2983_0, i_13_116_2985_0, i_13_116_3007_0, i_13_116_3027_0,
    i_13_116_3110_0, i_13_116_3154_0, i_13_116_3160_0, i_13_116_3211_0,
    i_13_116_3233_0, i_13_116_3386_0, i_13_116_3451_0, i_13_116_3549_0,
    i_13_116_3619_0, i_13_116_3710_0, i_13_116_3739_0, i_13_116_3763_0,
    i_13_116_3782_0, i_13_116_3817_0, i_13_116_3818_0, i_13_116_3872_0,
    i_13_116_4018_0, i_13_116_4054_0, i_13_116_4079_0, i_13_116_4084_0,
    i_13_116_4198_0, i_13_116_4258_0, i_13_116_4259_0, i_13_116_4376_0,
    i_13_116_4396_0, i_13_116_4511_0, i_13_116_4513_0, i_13_116_4522_0,
    i_13_116_4564_0, i_13_116_4565_0, i_13_116_4567_0, i_13_116_4570_0;
  output o_13_116_0_0;
  assign o_13_116_0_0 = ~((i_13_116_139_0 & ((~i_13_116_1399_0 & ~i_13_116_2981_0 & ~i_13_116_4376_0) | (i_13_116_3549_0 & i_13_116_4513_0))) | (~i_13_116_2980_0 & ((~i_13_116_2018_0 & ~i_13_116_2981_0 & ~i_13_116_4376_0) | (~i_13_116_193_0 & ~i_13_116_4565_0))) | (i_13_116_1552_0 & i_13_116_2857_0 & ~i_13_116_2981_0) | (~i_13_116_2108_0 & ~i_13_116_2982_0 & ~i_13_116_3872_0 & ~i_13_116_4565_0) | (~i_13_116_1552_0 & ~i_13_116_4513_0 & ~i_13_116_4567_0));
endmodule



// Benchmark "kernel_13_117" written by ABC on Sun Jul 19 10:47:03 2020

module kernel_13_117 ( 
    i_13_117_70_0, i_13_117_71_0, i_13_117_80_0, i_13_117_260_0,
    i_13_117_262_0, i_13_117_377_0, i_13_117_386_0, i_13_117_448_0,
    i_13_117_449_0, i_13_117_464_0, i_13_117_523_0, i_13_117_527_0,
    i_13_117_592_0, i_13_117_674_0, i_13_117_687_0, i_13_117_701_0,
    i_13_117_763_0, i_13_117_845_0, i_13_117_887_0, i_13_117_935_0,
    i_13_117_979_0, i_13_117_1070_0, i_13_117_1214_0, i_13_117_1346_0,
    i_13_117_1402_0, i_13_117_1403_0, i_13_117_1430_0, i_13_117_1439_0,
    i_13_117_1492_0, i_13_117_1538_0, i_13_117_1600_0, i_13_117_1601_0,
    i_13_117_1645_0, i_13_117_1722_0, i_13_117_1727_0, i_13_117_1731_0,
    i_13_117_1733_0, i_13_117_1736_0, i_13_117_1781_0, i_13_117_1798_0,
    i_13_117_1799_0, i_13_117_1810_0, i_13_117_1889_0, i_13_117_1934_0,
    i_13_117_1948_0, i_13_117_1993_0, i_13_117_2001_0, i_13_117_2002_0,
    i_13_117_2020_0, i_13_117_2030_0, i_13_117_2059_0, i_13_117_2177_0,
    i_13_117_2194_0, i_13_117_2197_0, i_13_117_2285_0, i_13_117_2376_0,
    i_13_117_2381_0, i_13_117_2384_0, i_13_117_2507_0, i_13_117_2552_0,
    i_13_117_2680_0, i_13_117_2699_0, i_13_117_2723_0, i_13_117_2726_0,
    i_13_117_2744_0, i_13_117_2770_0, i_13_117_2771_0, i_13_117_2888_0,
    i_13_117_2916_0, i_13_117_2917_0, i_13_117_2973_0, i_13_117_3032_0,
    i_13_117_3064_0, i_13_117_3140_0, i_13_117_3262_0, i_13_117_3367_0,
    i_13_117_3371_0, i_13_117_3418_0, i_13_117_3438_0, i_13_117_3442_0,
    i_13_117_3536_0, i_13_117_3596_0, i_13_117_3639_0, i_13_117_3641_0,
    i_13_117_3684_0, i_13_117_3689_0, i_13_117_3780_0, i_13_117_3842_0,
    i_13_117_3896_0, i_13_117_3928_0, i_13_117_3994_0, i_13_117_3995_0,
    i_13_117_4058_0, i_13_117_4096_0, i_13_117_4392_0, i_13_117_4429_0,
    i_13_117_4451_0, i_13_117_4501_0, i_13_117_4598_0, i_13_117_4599_0,
    o_13_117_0_0  );
  input  i_13_117_70_0, i_13_117_71_0, i_13_117_80_0, i_13_117_260_0,
    i_13_117_262_0, i_13_117_377_0, i_13_117_386_0, i_13_117_448_0,
    i_13_117_449_0, i_13_117_464_0, i_13_117_523_0, i_13_117_527_0,
    i_13_117_592_0, i_13_117_674_0, i_13_117_687_0, i_13_117_701_0,
    i_13_117_763_0, i_13_117_845_0, i_13_117_887_0, i_13_117_935_0,
    i_13_117_979_0, i_13_117_1070_0, i_13_117_1214_0, i_13_117_1346_0,
    i_13_117_1402_0, i_13_117_1403_0, i_13_117_1430_0, i_13_117_1439_0,
    i_13_117_1492_0, i_13_117_1538_0, i_13_117_1600_0, i_13_117_1601_0,
    i_13_117_1645_0, i_13_117_1722_0, i_13_117_1727_0, i_13_117_1731_0,
    i_13_117_1733_0, i_13_117_1736_0, i_13_117_1781_0, i_13_117_1798_0,
    i_13_117_1799_0, i_13_117_1810_0, i_13_117_1889_0, i_13_117_1934_0,
    i_13_117_1948_0, i_13_117_1993_0, i_13_117_2001_0, i_13_117_2002_0,
    i_13_117_2020_0, i_13_117_2030_0, i_13_117_2059_0, i_13_117_2177_0,
    i_13_117_2194_0, i_13_117_2197_0, i_13_117_2285_0, i_13_117_2376_0,
    i_13_117_2381_0, i_13_117_2384_0, i_13_117_2507_0, i_13_117_2552_0,
    i_13_117_2680_0, i_13_117_2699_0, i_13_117_2723_0, i_13_117_2726_0,
    i_13_117_2744_0, i_13_117_2770_0, i_13_117_2771_0, i_13_117_2888_0,
    i_13_117_2916_0, i_13_117_2917_0, i_13_117_2973_0, i_13_117_3032_0,
    i_13_117_3064_0, i_13_117_3140_0, i_13_117_3262_0, i_13_117_3367_0,
    i_13_117_3371_0, i_13_117_3418_0, i_13_117_3438_0, i_13_117_3442_0,
    i_13_117_3536_0, i_13_117_3596_0, i_13_117_3639_0, i_13_117_3641_0,
    i_13_117_3684_0, i_13_117_3689_0, i_13_117_3780_0, i_13_117_3842_0,
    i_13_117_3896_0, i_13_117_3928_0, i_13_117_3994_0, i_13_117_3995_0,
    i_13_117_4058_0, i_13_117_4096_0, i_13_117_4392_0, i_13_117_4429_0,
    i_13_117_4451_0, i_13_117_4501_0, i_13_117_4598_0, i_13_117_4599_0;
  output o_13_117_0_0;
  assign o_13_117_0_0 = ~((~i_13_117_1799_0 & ~i_13_117_4058_0) | (~i_13_117_71_0 & ~i_13_117_2744_0));
endmodule



// Benchmark "kernel_13_118" written by ABC on Sun Jul 19 10:47:04 2020

module kernel_13_118 ( 
    i_13_118_14_0, i_13_118_31_0, i_13_118_32_0, i_13_118_62_0,
    i_13_118_67_0, i_13_118_100_0, i_13_118_187_0, i_13_118_193_0,
    i_13_118_196_0, i_13_118_224_0, i_13_118_240_0, i_13_118_258_0,
    i_13_118_259_0, i_13_118_260_0, i_13_118_263_0, i_13_118_276_0,
    i_13_118_310_0, i_13_118_311_0, i_13_118_377_0, i_13_118_618_0,
    i_13_118_620_0, i_13_118_622_0, i_13_118_626_0, i_13_118_628_0,
    i_13_118_629_0, i_13_118_778_0, i_13_118_781_0, i_13_118_782_0,
    i_13_118_895_0, i_13_118_979_0, i_13_118_980_0, i_13_118_1077_0,
    i_13_118_1096_0, i_13_118_1112_0, i_13_118_1124_0, i_13_118_1140_0,
    i_13_118_1255_0, i_13_118_1256_0, i_13_118_1318_0, i_13_118_1391_0,
    i_13_118_1411_0, i_13_118_1469_0, i_13_118_1480_0, i_13_118_1483_0,
    i_13_118_1484_0, i_13_118_1558_0, i_13_118_1565_0, i_13_118_1643_0,
    i_13_118_1678_0, i_13_118_1688_0, i_13_118_1691_0, i_13_118_1745_0,
    i_13_118_1771_0, i_13_118_1805_0, i_13_118_1862_0, i_13_118_1991_0,
    i_13_118_2002_0, i_13_118_2120_0, i_13_118_2150_0, i_13_118_2291_0,
    i_13_118_2314_0, i_13_118_2365_0, i_13_118_2400_0, i_13_118_2425_0,
    i_13_118_2446_0, i_13_118_2447_0, i_13_118_2454_0, i_13_118_2677_0,
    i_13_118_2743_0, i_13_118_2857_0, i_13_118_2858_0, i_13_118_3005_0,
    i_13_118_3040_0, i_13_118_3131_0, i_13_118_3156_0, i_13_118_3292_0,
    i_13_118_3299_0, i_13_118_3356_0, i_13_118_3380_0, i_13_118_3383_0,
    i_13_118_3413_0, i_13_118_3419_0, i_13_118_3482_0, i_13_118_3523_0,
    i_13_118_3525_0, i_13_118_3526_0, i_13_118_3553_0, i_13_118_3554_0,
    i_13_118_3562_0, i_13_118_3570_0, i_13_118_3571_0, i_13_118_3642_0,
    i_13_118_4022_0, i_13_118_4254_0, i_13_118_4261_0, i_13_118_4364_0,
    i_13_118_4379_0, i_13_118_4391_0, i_13_118_4412_0, i_13_118_4508_0,
    o_13_118_0_0  );
  input  i_13_118_14_0, i_13_118_31_0, i_13_118_32_0, i_13_118_62_0,
    i_13_118_67_0, i_13_118_100_0, i_13_118_187_0, i_13_118_193_0,
    i_13_118_196_0, i_13_118_224_0, i_13_118_240_0, i_13_118_258_0,
    i_13_118_259_0, i_13_118_260_0, i_13_118_263_0, i_13_118_276_0,
    i_13_118_310_0, i_13_118_311_0, i_13_118_377_0, i_13_118_618_0,
    i_13_118_620_0, i_13_118_622_0, i_13_118_626_0, i_13_118_628_0,
    i_13_118_629_0, i_13_118_778_0, i_13_118_781_0, i_13_118_782_0,
    i_13_118_895_0, i_13_118_979_0, i_13_118_980_0, i_13_118_1077_0,
    i_13_118_1096_0, i_13_118_1112_0, i_13_118_1124_0, i_13_118_1140_0,
    i_13_118_1255_0, i_13_118_1256_0, i_13_118_1318_0, i_13_118_1391_0,
    i_13_118_1411_0, i_13_118_1469_0, i_13_118_1480_0, i_13_118_1483_0,
    i_13_118_1484_0, i_13_118_1558_0, i_13_118_1565_0, i_13_118_1643_0,
    i_13_118_1678_0, i_13_118_1688_0, i_13_118_1691_0, i_13_118_1745_0,
    i_13_118_1771_0, i_13_118_1805_0, i_13_118_1862_0, i_13_118_1991_0,
    i_13_118_2002_0, i_13_118_2120_0, i_13_118_2150_0, i_13_118_2291_0,
    i_13_118_2314_0, i_13_118_2365_0, i_13_118_2400_0, i_13_118_2425_0,
    i_13_118_2446_0, i_13_118_2447_0, i_13_118_2454_0, i_13_118_2677_0,
    i_13_118_2743_0, i_13_118_2857_0, i_13_118_2858_0, i_13_118_3005_0,
    i_13_118_3040_0, i_13_118_3131_0, i_13_118_3156_0, i_13_118_3292_0,
    i_13_118_3299_0, i_13_118_3356_0, i_13_118_3380_0, i_13_118_3383_0,
    i_13_118_3413_0, i_13_118_3419_0, i_13_118_3482_0, i_13_118_3523_0,
    i_13_118_3525_0, i_13_118_3526_0, i_13_118_3553_0, i_13_118_3554_0,
    i_13_118_3562_0, i_13_118_3570_0, i_13_118_3571_0, i_13_118_3642_0,
    i_13_118_4022_0, i_13_118_4254_0, i_13_118_4261_0, i_13_118_4364_0,
    i_13_118_4379_0, i_13_118_4391_0, i_13_118_4412_0, i_13_118_4508_0;
  output o_13_118_0_0;
  assign o_13_118_0_0 = ~((~i_13_118_2446_0 & ~i_13_118_2447_0 & ~i_13_118_2743_0) | (~i_13_118_618_0 & i_13_118_2002_0 & ~i_13_118_3571_0 & ~i_13_118_4364_0));
endmodule



// Benchmark "kernel_13_119" written by ABC on Sun Jul 19 10:47:04 2020

module kernel_13_119 ( 
    i_13_119_76_0, i_13_119_249_0, i_13_119_258_0, i_13_119_324_0,
    i_13_119_372_0, i_13_119_531_0, i_13_119_576_0, i_13_119_580_0,
    i_13_119_595_0, i_13_119_670_0, i_13_119_699_0, i_13_119_714_0,
    i_13_119_718_0, i_13_119_719_0, i_13_119_777_0, i_13_119_781_0,
    i_13_119_811_0, i_13_119_838_0, i_13_119_843_0, i_13_119_891_0,
    i_13_119_942_0, i_13_119_1036_0, i_13_119_1092_0, i_13_119_1098_0,
    i_13_119_1116_0, i_13_119_1192_0, i_13_119_1321_0, i_13_119_1380_0,
    i_13_119_1461_0, i_13_119_1462_0, i_13_119_1479_0, i_13_119_1500_0,
    i_13_119_1664_0, i_13_119_1710_0, i_13_119_1743_0, i_13_119_1746_0,
    i_13_119_1756_0, i_13_119_1884_0, i_13_119_1887_0, i_13_119_1979_0,
    i_13_119_2140_0, i_13_119_2223_0, i_13_119_2224_0, i_13_119_2388_0,
    i_13_119_2404_0, i_13_119_2442_0, i_13_119_2452_0, i_13_119_2457_0,
    i_13_119_2499_0, i_13_119_2502_0, i_13_119_2565_0, i_13_119_2616_0,
    i_13_119_2633_0, i_13_119_2646_0, i_13_119_2667_0, i_13_119_2752_0,
    i_13_119_2820_0, i_13_119_2821_0, i_13_119_2824_0, i_13_119_3034_0,
    i_13_119_3046_0, i_13_119_3108_0, i_13_119_3171_0, i_13_119_3172_0,
    i_13_119_3216_0, i_13_119_3286_0, i_13_119_3289_0, i_13_119_3294_0,
    i_13_119_3306_0, i_13_119_3324_0, i_13_119_3372_0, i_13_119_3379_0,
    i_13_119_3433_0, i_13_119_3447_0, i_13_119_3462_0, i_13_119_3525_0,
    i_13_119_3559_0, i_13_119_3613_0, i_13_119_3639_0, i_13_119_3733_0,
    i_13_119_3790_0, i_13_119_3794_0, i_13_119_3798_0, i_13_119_3873_0,
    i_13_119_3913_0, i_13_119_3988_0, i_13_119_3992_0, i_13_119_4008_0,
    i_13_119_4212_0, i_13_119_4238_0, i_13_119_4377_0, i_13_119_4382_0,
    i_13_119_4387_0, i_13_119_4389_0, i_13_119_4410_0, i_13_119_4411_0,
    i_13_119_4440_0, i_13_119_4518_0, i_13_119_4557_0, i_13_119_4561_0,
    o_13_119_0_0  );
  input  i_13_119_76_0, i_13_119_249_0, i_13_119_258_0, i_13_119_324_0,
    i_13_119_372_0, i_13_119_531_0, i_13_119_576_0, i_13_119_580_0,
    i_13_119_595_0, i_13_119_670_0, i_13_119_699_0, i_13_119_714_0,
    i_13_119_718_0, i_13_119_719_0, i_13_119_777_0, i_13_119_781_0,
    i_13_119_811_0, i_13_119_838_0, i_13_119_843_0, i_13_119_891_0,
    i_13_119_942_0, i_13_119_1036_0, i_13_119_1092_0, i_13_119_1098_0,
    i_13_119_1116_0, i_13_119_1192_0, i_13_119_1321_0, i_13_119_1380_0,
    i_13_119_1461_0, i_13_119_1462_0, i_13_119_1479_0, i_13_119_1500_0,
    i_13_119_1664_0, i_13_119_1710_0, i_13_119_1743_0, i_13_119_1746_0,
    i_13_119_1756_0, i_13_119_1884_0, i_13_119_1887_0, i_13_119_1979_0,
    i_13_119_2140_0, i_13_119_2223_0, i_13_119_2224_0, i_13_119_2388_0,
    i_13_119_2404_0, i_13_119_2442_0, i_13_119_2452_0, i_13_119_2457_0,
    i_13_119_2499_0, i_13_119_2502_0, i_13_119_2565_0, i_13_119_2616_0,
    i_13_119_2633_0, i_13_119_2646_0, i_13_119_2667_0, i_13_119_2752_0,
    i_13_119_2820_0, i_13_119_2821_0, i_13_119_2824_0, i_13_119_3034_0,
    i_13_119_3046_0, i_13_119_3108_0, i_13_119_3171_0, i_13_119_3172_0,
    i_13_119_3216_0, i_13_119_3286_0, i_13_119_3289_0, i_13_119_3294_0,
    i_13_119_3306_0, i_13_119_3324_0, i_13_119_3372_0, i_13_119_3379_0,
    i_13_119_3433_0, i_13_119_3447_0, i_13_119_3462_0, i_13_119_3525_0,
    i_13_119_3559_0, i_13_119_3613_0, i_13_119_3639_0, i_13_119_3733_0,
    i_13_119_3790_0, i_13_119_3794_0, i_13_119_3798_0, i_13_119_3873_0,
    i_13_119_3913_0, i_13_119_3988_0, i_13_119_3992_0, i_13_119_4008_0,
    i_13_119_4212_0, i_13_119_4238_0, i_13_119_4377_0, i_13_119_4382_0,
    i_13_119_4387_0, i_13_119_4389_0, i_13_119_4410_0, i_13_119_4411_0,
    i_13_119_4440_0, i_13_119_4518_0, i_13_119_4557_0, i_13_119_4561_0;
  output o_13_119_0_0;
  assign o_13_119_0_0 = ~(~i_13_119_891_0 | ~i_13_119_3286_0);
endmodule



// Benchmark "kernel_13_120" written by ABC on Sun Jul 19 10:47:05 2020

module kernel_13_120 ( 
    i_13_120_49_0, i_13_120_70_0, i_13_120_142_0, i_13_120_187_0,
    i_13_120_428_0, i_13_120_447_0, i_13_120_448_0, i_13_120_571_0,
    i_13_120_612_0, i_13_120_639_0, i_13_120_646_0, i_13_120_672_0,
    i_13_120_682_0, i_13_120_683_0, i_13_120_688_0, i_13_120_701_0,
    i_13_120_818_0, i_13_120_823_0, i_13_120_843_0, i_13_120_1105_0,
    i_13_120_1116_0, i_13_120_1123_0, i_13_120_1124_0, i_13_120_1269_0,
    i_13_120_1276_0, i_13_120_1277_0, i_13_120_1313_0, i_13_120_1374_0,
    i_13_120_1403_0, i_13_120_1474_0, i_13_120_1510_0, i_13_120_1511_0,
    i_13_120_1599_0, i_13_120_1600_0, i_13_120_1601_0, i_13_120_1638_0,
    i_13_120_1644_0, i_13_120_1645_0, i_13_120_1672_0, i_13_120_1726_0,
    i_13_120_1727_0, i_13_120_1736_0, i_13_120_1798_0, i_13_120_1925_0,
    i_13_120_1933_0, i_13_120_1996_0, i_13_120_2005_0, i_13_120_2052_0,
    i_13_120_2057_0, i_13_120_2107_0, i_13_120_2116_0, i_13_120_2133_0,
    i_13_120_2194_0, i_13_120_2266_0, i_13_120_2278_0, i_13_120_2403_0,
    i_13_120_2455_0, i_13_120_2456_0, i_13_120_2614_0, i_13_120_2679_0,
    i_13_120_2680_0, i_13_120_2697_0, i_13_120_2698_0, i_13_120_2699_0,
    i_13_120_2746_0, i_13_120_2887_0, i_13_120_2934_0, i_13_120_2940_0,
    i_13_120_3024_0, i_13_120_3113_0, i_13_120_3285_0, i_13_120_3393_0,
    i_13_120_3519_0, i_13_120_3595_0, i_13_120_3596_0, i_13_120_3652_0,
    i_13_120_3653_0, i_13_120_3733_0, i_13_120_3753_0, i_13_120_3797_0,
    i_13_120_3930_0, i_13_120_3940_0, i_13_120_3994_0, i_13_120_3995_0,
    i_13_120_4018_0, i_13_120_4019_0, i_13_120_4039_0, i_13_120_4085_0,
    i_13_120_4121_0, i_13_120_4252_0, i_13_120_4255_0, i_13_120_4262_0,
    i_13_120_4309_0, i_13_120_4310_0, i_13_120_4311_0, i_13_120_4318_0,
    i_13_120_4396_0, i_13_120_4559_0, i_13_120_4597_0, i_13_120_4598_0,
    o_13_120_0_0  );
  input  i_13_120_49_0, i_13_120_70_0, i_13_120_142_0, i_13_120_187_0,
    i_13_120_428_0, i_13_120_447_0, i_13_120_448_0, i_13_120_571_0,
    i_13_120_612_0, i_13_120_639_0, i_13_120_646_0, i_13_120_672_0,
    i_13_120_682_0, i_13_120_683_0, i_13_120_688_0, i_13_120_701_0,
    i_13_120_818_0, i_13_120_823_0, i_13_120_843_0, i_13_120_1105_0,
    i_13_120_1116_0, i_13_120_1123_0, i_13_120_1124_0, i_13_120_1269_0,
    i_13_120_1276_0, i_13_120_1277_0, i_13_120_1313_0, i_13_120_1374_0,
    i_13_120_1403_0, i_13_120_1474_0, i_13_120_1510_0, i_13_120_1511_0,
    i_13_120_1599_0, i_13_120_1600_0, i_13_120_1601_0, i_13_120_1638_0,
    i_13_120_1644_0, i_13_120_1645_0, i_13_120_1672_0, i_13_120_1726_0,
    i_13_120_1727_0, i_13_120_1736_0, i_13_120_1798_0, i_13_120_1925_0,
    i_13_120_1933_0, i_13_120_1996_0, i_13_120_2005_0, i_13_120_2052_0,
    i_13_120_2057_0, i_13_120_2107_0, i_13_120_2116_0, i_13_120_2133_0,
    i_13_120_2194_0, i_13_120_2266_0, i_13_120_2278_0, i_13_120_2403_0,
    i_13_120_2455_0, i_13_120_2456_0, i_13_120_2614_0, i_13_120_2679_0,
    i_13_120_2680_0, i_13_120_2697_0, i_13_120_2698_0, i_13_120_2699_0,
    i_13_120_2746_0, i_13_120_2887_0, i_13_120_2934_0, i_13_120_2940_0,
    i_13_120_3024_0, i_13_120_3113_0, i_13_120_3285_0, i_13_120_3393_0,
    i_13_120_3519_0, i_13_120_3595_0, i_13_120_3596_0, i_13_120_3652_0,
    i_13_120_3653_0, i_13_120_3733_0, i_13_120_3753_0, i_13_120_3797_0,
    i_13_120_3930_0, i_13_120_3940_0, i_13_120_3994_0, i_13_120_3995_0,
    i_13_120_4018_0, i_13_120_4019_0, i_13_120_4039_0, i_13_120_4085_0,
    i_13_120_4121_0, i_13_120_4252_0, i_13_120_4255_0, i_13_120_4262_0,
    i_13_120_4309_0, i_13_120_4310_0, i_13_120_4311_0, i_13_120_4318_0,
    i_13_120_4396_0, i_13_120_4559_0, i_13_120_4597_0, i_13_120_4598_0;
  output o_13_120_0_0;
  assign o_13_120_0_0 = ~((~i_13_120_1798_0 & ((~i_13_120_1276_0 & ~i_13_120_2456_0 & ~i_13_120_3653_0 & ~i_13_120_4255_0) | (~i_13_120_1511_0 & ~i_13_120_3930_0 & ~i_13_120_4310_0))) | (~i_13_120_823_0 & i_13_120_2614_0 & ~i_13_120_3652_0 & ~i_13_120_3733_0) | (~i_13_120_70_0 & i_13_120_1474_0 & ~i_13_120_4318_0));
endmodule



// Benchmark "kernel_13_121" written by ABC on Sun Jul 19 10:47:06 2020

module kernel_13_121 ( 
    i_13_121_1_0, i_13_121_31_0, i_13_121_36_0, i_13_121_37_0,
    i_13_121_76_0, i_13_121_99_0, i_13_121_163_0, i_13_121_165_0,
    i_13_121_167_0, i_13_121_168_0, i_13_121_183_0, i_13_121_184_0,
    i_13_121_217_0, i_13_121_336_0, i_13_121_372_0, i_13_121_526_0,
    i_13_121_532_0, i_13_121_570_0, i_13_121_676_0, i_13_121_686_0,
    i_13_121_714_0, i_13_121_718_0, i_13_121_813_0, i_13_121_814_0,
    i_13_121_1027_0, i_13_121_1067_0, i_13_121_1210_0, i_13_121_1272_0,
    i_13_121_1426_0, i_13_121_1495_0, i_13_121_1515_0, i_13_121_1525_0,
    i_13_121_1597_0, i_13_121_1677_0, i_13_121_1683_0, i_13_121_1731_0,
    i_13_121_1746_0, i_13_121_1747_0, i_13_121_1749_0, i_13_121_1756_0,
    i_13_121_1782_0, i_13_121_1801_0, i_13_121_1804_0, i_13_121_1805_0,
    i_13_121_1831_0, i_13_121_1832_0, i_13_121_1909_0, i_13_121_1911_0,
    i_13_121_2043_0, i_13_121_2046_0, i_13_121_2115_0, i_13_121_2116_0,
    i_13_121_2233_0, i_13_121_2263_0, i_13_121_2277_0, i_13_121_2407_0,
    i_13_121_2434_0, i_13_121_2476_0, i_13_121_2556_0, i_13_121_2722_0,
    i_13_121_2736_0, i_13_121_2748_0, i_13_121_2857_0, i_13_121_2889_0,
    i_13_121_2937_0, i_13_121_2980_0, i_13_121_3024_0, i_13_121_3027_0,
    i_13_121_3091_0, i_13_121_3126_0, i_13_121_3142_0, i_13_121_3196_0,
    i_13_121_3205_0, i_13_121_3216_0, i_13_121_3249_0, i_13_121_3289_0,
    i_13_121_3414_0, i_13_121_3444_0, i_13_121_3445_0, i_13_121_3472_0,
    i_13_121_3519_0, i_13_121_3549_0, i_13_121_3607_0, i_13_121_3661_0,
    i_13_121_3720_0, i_13_121_3739_0, i_13_121_3817_0, i_13_121_3918_0,
    i_13_121_3919_0, i_13_121_3988_0, i_13_121_4036_0, i_13_121_4044_0,
    i_13_121_4045_0, i_13_121_4059_0, i_13_121_4404_0, i_13_121_4413_0,
    i_13_121_4425_0, i_13_121_4497_0, i_13_121_4521_0, i_13_121_4593_0,
    o_13_121_0_0  );
  input  i_13_121_1_0, i_13_121_31_0, i_13_121_36_0, i_13_121_37_0,
    i_13_121_76_0, i_13_121_99_0, i_13_121_163_0, i_13_121_165_0,
    i_13_121_167_0, i_13_121_168_0, i_13_121_183_0, i_13_121_184_0,
    i_13_121_217_0, i_13_121_336_0, i_13_121_372_0, i_13_121_526_0,
    i_13_121_532_0, i_13_121_570_0, i_13_121_676_0, i_13_121_686_0,
    i_13_121_714_0, i_13_121_718_0, i_13_121_813_0, i_13_121_814_0,
    i_13_121_1027_0, i_13_121_1067_0, i_13_121_1210_0, i_13_121_1272_0,
    i_13_121_1426_0, i_13_121_1495_0, i_13_121_1515_0, i_13_121_1525_0,
    i_13_121_1597_0, i_13_121_1677_0, i_13_121_1683_0, i_13_121_1731_0,
    i_13_121_1746_0, i_13_121_1747_0, i_13_121_1749_0, i_13_121_1756_0,
    i_13_121_1782_0, i_13_121_1801_0, i_13_121_1804_0, i_13_121_1805_0,
    i_13_121_1831_0, i_13_121_1832_0, i_13_121_1909_0, i_13_121_1911_0,
    i_13_121_2043_0, i_13_121_2046_0, i_13_121_2115_0, i_13_121_2116_0,
    i_13_121_2233_0, i_13_121_2263_0, i_13_121_2277_0, i_13_121_2407_0,
    i_13_121_2434_0, i_13_121_2476_0, i_13_121_2556_0, i_13_121_2722_0,
    i_13_121_2736_0, i_13_121_2748_0, i_13_121_2857_0, i_13_121_2889_0,
    i_13_121_2937_0, i_13_121_2980_0, i_13_121_3024_0, i_13_121_3027_0,
    i_13_121_3091_0, i_13_121_3126_0, i_13_121_3142_0, i_13_121_3196_0,
    i_13_121_3205_0, i_13_121_3216_0, i_13_121_3249_0, i_13_121_3289_0,
    i_13_121_3414_0, i_13_121_3444_0, i_13_121_3445_0, i_13_121_3472_0,
    i_13_121_3519_0, i_13_121_3549_0, i_13_121_3607_0, i_13_121_3661_0,
    i_13_121_3720_0, i_13_121_3739_0, i_13_121_3817_0, i_13_121_3918_0,
    i_13_121_3919_0, i_13_121_3988_0, i_13_121_4036_0, i_13_121_4044_0,
    i_13_121_4045_0, i_13_121_4059_0, i_13_121_4404_0, i_13_121_4413_0,
    i_13_121_4425_0, i_13_121_4497_0, i_13_121_4521_0, i_13_121_4593_0;
  output o_13_121_0_0;
  assign o_13_121_0_0 = ~((i_13_121_1426_0 & ((~i_13_121_183_0 & ~i_13_121_1747_0 & ~i_13_121_1801_0 & ~i_13_121_2736_0) | (~i_13_121_2407_0 & ~i_13_121_3988_0))) | (~i_13_121_1677_0 & ((i_13_121_1597_0 & i_13_121_2857_0 & ~i_13_121_2980_0) | (~i_13_121_1747_0 & ~i_13_121_4059_0 & ~i_13_121_4413_0))) | (~i_13_121_2980_0 & ((~i_13_121_570_0 & ~i_13_121_1597_0 & ~i_13_121_1831_0) | (i_13_121_526_0 & i_13_121_1832_0))) | (~i_13_121_4036_0 & ((~i_13_121_1731_0 & i_13_121_3918_0) | (~i_13_121_1747_0 & ~i_13_121_1749_0 & ~i_13_121_3445_0 & ~i_13_121_4059_0))) | (i_13_121_1067_0 & ~i_13_121_3988_0) | (~i_13_121_813_0 & ~i_13_121_1525_0 & i_13_121_1831_0 & ~i_13_121_3216_0 & i_13_121_4036_0 & ~i_13_121_4045_0));
endmodule



// Benchmark "kernel_13_122" written by ABC on Sun Jul 19 10:47:07 2020

module kernel_13_122 ( 
    i_13_122_40_0, i_13_122_50_0, i_13_122_112_0, i_13_122_115_0,
    i_13_122_121_0, i_13_122_192_0, i_13_122_251_0, i_13_122_274_0,
    i_13_122_277_0, i_13_122_415_0, i_13_122_457_0, i_13_122_561_0,
    i_13_122_562_0, i_13_122_607_0, i_13_122_616_0, i_13_122_688_0,
    i_13_122_928_0, i_13_122_951_0, i_13_122_952_0, i_13_122_1084_0,
    i_13_122_1085_0, i_13_122_1134_0, i_13_122_1141_0, i_13_122_1163_0,
    i_13_122_1273_0, i_13_122_1318_0, i_13_122_1444_0, i_13_122_1502_0,
    i_13_122_1573_0, i_13_122_1624_0, i_13_122_1633_0, i_13_122_1636_0,
    i_13_122_1642_0, i_13_122_1669_0, i_13_122_1678_0, i_13_122_1750_0,
    i_13_122_1839_0, i_13_122_1840_0, i_13_122_1858_0, i_13_122_1885_0,
    i_13_122_1930_0, i_13_122_2116_0, i_13_122_2175_0, i_13_122_2206_0,
    i_13_122_2233_0, i_13_122_2380_0, i_13_122_2433_0, i_13_122_2434_0,
    i_13_122_2435_0, i_13_122_2437_0, i_13_122_2438_0, i_13_122_2465_0,
    i_13_122_2505_0, i_13_122_2541_0, i_13_122_2590_0, i_13_122_2650_0,
    i_13_122_2716_0, i_13_122_2875_0, i_13_122_3004_0, i_13_122_3016_0,
    i_13_122_3047_0, i_13_122_3098_0, i_13_122_3101_0, i_13_122_3145_0,
    i_13_122_3146_0, i_13_122_3160_0, i_13_122_3162_0, i_13_122_3163_0,
    i_13_122_3166_0, i_13_122_3379_0, i_13_122_3455_0, i_13_122_3473_0,
    i_13_122_3527_0, i_13_122_3541_0, i_13_122_3604_0, i_13_122_3686_0,
    i_13_122_3688_0, i_13_122_3689_0, i_13_122_3784_0, i_13_122_3871_0,
    i_13_122_3872_0, i_13_122_3874_0, i_13_122_3904_0, i_13_122_3938_0,
    i_13_122_3991_0, i_13_122_4036_0, i_13_122_4057_0, i_13_122_4094_0,
    i_13_122_4158_0, i_13_122_4207_0, i_13_122_4253_0, i_13_122_4324_0,
    i_13_122_4350_0, i_13_122_4351_0, i_13_122_4352_0, i_13_122_4378_0,
    i_13_122_4379_0, i_13_122_4429_0, i_13_122_4468_0, i_13_122_4593_0,
    o_13_122_0_0  );
  input  i_13_122_40_0, i_13_122_50_0, i_13_122_112_0, i_13_122_115_0,
    i_13_122_121_0, i_13_122_192_0, i_13_122_251_0, i_13_122_274_0,
    i_13_122_277_0, i_13_122_415_0, i_13_122_457_0, i_13_122_561_0,
    i_13_122_562_0, i_13_122_607_0, i_13_122_616_0, i_13_122_688_0,
    i_13_122_928_0, i_13_122_951_0, i_13_122_952_0, i_13_122_1084_0,
    i_13_122_1085_0, i_13_122_1134_0, i_13_122_1141_0, i_13_122_1163_0,
    i_13_122_1273_0, i_13_122_1318_0, i_13_122_1444_0, i_13_122_1502_0,
    i_13_122_1573_0, i_13_122_1624_0, i_13_122_1633_0, i_13_122_1636_0,
    i_13_122_1642_0, i_13_122_1669_0, i_13_122_1678_0, i_13_122_1750_0,
    i_13_122_1839_0, i_13_122_1840_0, i_13_122_1858_0, i_13_122_1885_0,
    i_13_122_1930_0, i_13_122_2116_0, i_13_122_2175_0, i_13_122_2206_0,
    i_13_122_2233_0, i_13_122_2380_0, i_13_122_2433_0, i_13_122_2434_0,
    i_13_122_2435_0, i_13_122_2437_0, i_13_122_2438_0, i_13_122_2465_0,
    i_13_122_2505_0, i_13_122_2541_0, i_13_122_2590_0, i_13_122_2650_0,
    i_13_122_2716_0, i_13_122_2875_0, i_13_122_3004_0, i_13_122_3016_0,
    i_13_122_3047_0, i_13_122_3098_0, i_13_122_3101_0, i_13_122_3145_0,
    i_13_122_3146_0, i_13_122_3160_0, i_13_122_3162_0, i_13_122_3163_0,
    i_13_122_3166_0, i_13_122_3379_0, i_13_122_3455_0, i_13_122_3473_0,
    i_13_122_3527_0, i_13_122_3541_0, i_13_122_3604_0, i_13_122_3686_0,
    i_13_122_3688_0, i_13_122_3689_0, i_13_122_3784_0, i_13_122_3871_0,
    i_13_122_3872_0, i_13_122_3874_0, i_13_122_3904_0, i_13_122_3938_0,
    i_13_122_3991_0, i_13_122_4036_0, i_13_122_4057_0, i_13_122_4094_0,
    i_13_122_4158_0, i_13_122_4207_0, i_13_122_4253_0, i_13_122_4324_0,
    i_13_122_4350_0, i_13_122_4351_0, i_13_122_4352_0, i_13_122_4378_0,
    i_13_122_4379_0, i_13_122_4429_0, i_13_122_4468_0, i_13_122_4593_0;
  output o_13_122_0_0;
  assign o_13_122_0_0 = ~((~i_13_122_3604_0 & ((~i_13_122_1839_0 & ~i_13_122_2716_0 & ~i_13_122_3101_0) | (~i_13_122_1502_0 & ~i_13_122_3098_0 & ~i_13_122_3162_0 & ~i_13_122_3689_0 & ~i_13_122_3904_0))) | (~i_13_122_561_0 & ~i_13_122_1085_0 & i_13_122_2380_0) | (~i_13_122_115_0 & ~i_13_122_277_0 & ~i_13_122_1624_0 & i_13_122_4036_0 & ~i_13_122_4352_0));
endmodule



// Benchmark "kernel_13_123" written by ABC on Sun Jul 19 10:47:08 2020

module kernel_13_123 ( 
    i_13_123_46_0, i_13_123_91_0, i_13_123_100_0, i_13_123_121_0,
    i_13_123_167_0, i_13_123_169_0, i_13_123_219_0, i_13_123_280_0,
    i_13_123_284_0, i_13_123_379_0, i_13_123_380_0, i_13_123_425_0,
    i_13_123_523_0, i_13_123_535_0, i_13_123_571_0, i_13_123_697_0,
    i_13_123_730_0, i_13_123_731_0, i_13_123_928_0, i_13_123_949_0,
    i_13_123_954_0, i_13_123_1063_0, i_13_123_1064_0, i_13_123_1093_0,
    i_13_123_1156_0, i_13_123_1297_0, i_13_123_1323_0, i_13_123_1324_0,
    i_13_123_1381_0, i_13_123_1441_0, i_13_123_1443_0, i_13_123_1471_0,
    i_13_123_1495_0, i_13_123_1525_0, i_13_123_1783_0, i_13_123_1800_0,
    i_13_123_1810_0, i_13_123_1828_0, i_13_123_1829_0, i_13_123_1846_0,
    i_13_123_1848_0, i_13_123_1849_0, i_13_123_1850_0, i_13_123_1928_0,
    i_13_123_2053_0, i_13_123_2107_0, i_13_123_2108_0, i_13_123_2116_0,
    i_13_123_2133_0, i_13_123_2134_0, i_13_123_2205_0, i_13_123_2232_0,
    i_13_123_2233_0, i_13_123_2234_0, i_13_123_2342_0, i_13_123_2404_0,
    i_13_123_2544_0, i_13_123_2746_0, i_13_123_2793_0, i_13_123_2848_0,
    i_13_123_2854_0, i_13_123_2872_0, i_13_123_2925_0, i_13_123_2935_0,
    i_13_123_3007_0, i_13_123_3053_0, i_13_123_3091_0, i_13_123_3108_0,
    i_13_123_3109_0, i_13_123_3110_0, i_13_123_3232_0, i_13_123_3242_0,
    i_13_123_3244_0, i_13_123_3306_0, i_13_123_3386_0, i_13_123_3394_0,
    i_13_123_3431_0, i_13_123_3612_0, i_13_123_3613_0, i_13_123_3739_0,
    i_13_123_3762_0, i_13_123_3765_0, i_13_123_3769_0, i_13_123_3817_0,
    i_13_123_3818_0, i_13_123_3820_0, i_13_123_3996_0, i_13_123_4015_0,
    i_13_123_4016_0, i_13_123_4042_0, i_13_123_4060_0, i_13_123_4061_0,
    i_13_123_4063_0, i_13_123_4064_0, i_13_123_4231_0, i_13_123_4249_0,
    i_13_123_4250_0, i_13_123_4267_0, i_13_123_4268_0, i_13_123_4567_0,
    o_13_123_0_0  );
  input  i_13_123_46_0, i_13_123_91_0, i_13_123_100_0, i_13_123_121_0,
    i_13_123_167_0, i_13_123_169_0, i_13_123_219_0, i_13_123_280_0,
    i_13_123_284_0, i_13_123_379_0, i_13_123_380_0, i_13_123_425_0,
    i_13_123_523_0, i_13_123_535_0, i_13_123_571_0, i_13_123_697_0,
    i_13_123_730_0, i_13_123_731_0, i_13_123_928_0, i_13_123_949_0,
    i_13_123_954_0, i_13_123_1063_0, i_13_123_1064_0, i_13_123_1093_0,
    i_13_123_1156_0, i_13_123_1297_0, i_13_123_1323_0, i_13_123_1324_0,
    i_13_123_1381_0, i_13_123_1441_0, i_13_123_1443_0, i_13_123_1471_0,
    i_13_123_1495_0, i_13_123_1525_0, i_13_123_1783_0, i_13_123_1800_0,
    i_13_123_1810_0, i_13_123_1828_0, i_13_123_1829_0, i_13_123_1846_0,
    i_13_123_1848_0, i_13_123_1849_0, i_13_123_1850_0, i_13_123_1928_0,
    i_13_123_2053_0, i_13_123_2107_0, i_13_123_2108_0, i_13_123_2116_0,
    i_13_123_2133_0, i_13_123_2134_0, i_13_123_2205_0, i_13_123_2232_0,
    i_13_123_2233_0, i_13_123_2234_0, i_13_123_2342_0, i_13_123_2404_0,
    i_13_123_2544_0, i_13_123_2746_0, i_13_123_2793_0, i_13_123_2848_0,
    i_13_123_2854_0, i_13_123_2872_0, i_13_123_2925_0, i_13_123_2935_0,
    i_13_123_3007_0, i_13_123_3053_0, i_13_123_3091_0, i_13_123_3108_0,
    i_13_123_3109_0, i_13_123_3110_0, i_13_123_3232_0, i_13_123_3242_0,
    i_13_123_3244_0, i_13_123_3306_0, i_13_123_3386_0, i_13_123_3394_0,
    i_13_123_3431_0, i_13_123_3612_0, i_13_123_3613_0, i_13_123_3739_0,
    i_13_123_3762_0, i_13_123_3765_0, i_13_123_3769_0, i_13_123_3817_0,
    i_13_123_3818_0, i_13_123_3820_0, i_13_123_3996_0, i_13_123_4015_0,
    i_13_123_4016_0, i_13_123_4042_0, i_13_123_4060_0, i_13_123_4061_0,
    i_13_123_4063_0, i_13_123_4064_0, i_13_123_4231_0, i_13_123_4249_0,
    i_13_123_4250_0, i_13_123_4267_0, i_13_123_4268_0, i_13_123_4567_0;
  output o_13_123_0_0;
  assign o_13_123_0_0 = ~((~i_13_123_2233_0 & ~i_13_123_3818_0) | (~i_13_123_3232_0 & i_13_123_3765_0));
endmodule



// Benchmark "kernel_13_124" written by ABC on Sun Jul 19 10:47:09 2020

module kernel_13_124 ( 
    i_13_124_63_0, i_13_124_64_0, i_13_124_73_0, i_13_124_130_0,
    i_13_124_139_0, i_13_124_175_0, i_13_124_191_0, i_13_124_283_0,
    i_13_124_354_0, i_13_124_355_0, i_13_124_356_0, i_13_124_357_0,
    i_13_124_450_0, i_13_124_468_0, i_13_124_469_0, i_13_124_470_0,
    i_13_124_485_0, i_13_124_507_0, i_13_124_668_0, i_13_124_694_0,
    i_13_124_831_0, i_13_124_883_0, i_13_124_946_0, i_13_124_947_0,
    i_13_124_1099_0, i_13_124_1208_0, i_13_124_1219_0, i_13_124_1337_0,
    i_13_124_1393_0, i_13_124_1395_0, i_13_124_1396_0, i_13_124_1517_0,
    i_13_124_1554_0, i_13_124_1696_0, i_13_124_1719_0, i_13_124_1721_0,
    i_13_124_1729_0, i_13_124_1730_0, i_13_124_1774_0, i_13_124_1777_0,
    i_13_124_1838_0, i_13_124_1846_0, i_13_124_1927_0, i_13_124_2143_0,
    i_13_124_2202_0, i_13_124_2230_0, i_13_124_2231_0, i_13_124_2366_0,
    i_13_124_2426_0, i_13_124_2430_0, i_13_124_2443_0, i_13_124_2444_0,
    i_13_124_2461_0, i_13_124_2466_0, i_13_124_2477_0, i_13_124_2511_0,
    i_13_124_2512_0, i_13_124_2538_0, i_13_124_2608_0, i_13_124_2692_0,
    i_13_124_2719_0, i_13_124_2755_0, i_13_124_2845_0, i_13_124_2881_0,
    i_13_124_2882_0, i_13_124_2920_0, i_13_124_2921_0, i_13_124_2938_0,
    i_13_124_3012_0, i_13_124_3087_0, i_13_124_3128_0, i_13_124_3133_0,
    i_13_124_3208_0, i_13_124_3370_0, i_13_124_3375_0, i_13_124_3532_0,
    i_13_124_3547_0, i_13_124_3595_0, i_13_124_3596_0, i_13_124_3619_0,
    i_13_124_3620_0, i_13_124_3632_0, i_13_124_3754_0, i_13_124_3781_0,
    i_13_124_3793_0, i_13_124_3924_0, i_13_124_3935_0, i_13_124_3982_0,
    i_13_124_3987_0, i_13_124_4162_0, i_13_124_4213_0, i_13_124_4214_0,
    i_13_124_4312_0, i_13_124_4329_0, i_13_124_4330_0, i_13_124_4331_0,
    i_13_124_4429_0, i_13_124_4450_0, i_13_124_4513_0, i_13_124_4540_0,
    o_13_124_0_0  );
  input  i_13_124_63_0, i_13_124_64_0, i_13_124_73_0, i_13_124_130_0,
    i_13_124_139_0, i_13_124_175_0, i_13_124_191_0, i_13_124_283_0,
    i_13_124_354_0, i_13_124_355_0, i_13_124_356_0, i_13_124_357_0,
    i_13_124_450_0, i_13_124_468_0, i_13_124_469_0, i_13_124_470_0,
    i_13_124_485_0, i_13_124_507_0, i_13_124_668_0, i_13_124_694_0,
    i_13_124_831_0, i_13_124_883_0, i_13_124_946_0, i_13_124_947_0,
    i_13_124_1099_0, i_13_124_1208_0, i_13_124_1219_0, i_13_124_1337_0,
    i_13_124_1393_0, i_13_124_1395_0, i_13_124_1396_0, i_13_124_1517_0,
    i_13_124_1554_0, i_13_124_1696_0, i_13_124_1719_0, i_13_124_1721_0,
    i_13_124_1729_0, i_13_124_1730_0, i_13_124_1774_0, i_13_124_1777_0,
    i_13_124_1838_0, i_13_124_1846_0, i_13_124_1927_0, i_13_124_2143_0,
    i_13_124_2202_0, i_13_124_2230_0, i_13_124_2231_0, i_13_124_2366_0,
    i_13_124_2426_0, i_13_124_2430_0, i_13_124_2443_0, i_13_124_2444_0,
    i_13_124_2461_0, i_13_124_2466_0, i_13_124_2477_0, i_13_124_2511_0,
    i_13_124_2512_0, i_13_124_2538_0, i_13_124_2608_0, i_13_124_2692_0,
    i_13_124_2719_0, i_13_124_2755_0, i_13_124_2845_0, i_13_124_2881_0,
    i_13_124_2882_0, i_13_124_2920_0, i_13_124_2921_0, i_13_124_2938_0,
    i_13_124_3012_0, i_13_124_3087_0, i_13_124_3128_0, i_13_124_3133_0,
    i_13_124_3208_0, i_13_124_3370_0, i_13_124_3375_0, i_13_124_3532_0,
    i_13_124_3547_0, i_13_124_3595_0, i_13_124_3596_0, i_13_124_3619_0,
    i_13_124_3620_0, i_13_124_3632_0, i_13_124_3754_0, i_13_124_3781_0,
    i_13_124_3793_0, i_13_124_3924_0, i_13_124_3935_0, i_13_124_3982_0,
    i_13_124_3987_0, i_13_124_4162_0, i_13_124_4213_0, i_13_124_4214_0,
    i_13_124_4312_0, i_13_124_4329_0, i_13_124_4330_0, i_13_124_4331_0,
    i_13_124_4429_0, i_13_124_4450_0, i_13_124_4513_0, i_13_124_4540_0;
  output o_13_124_0_0;
  assign o_13_124_0_0 = ~(~i_13_124_4429_0 & (i_13_124_2430_0 | (~i_13_124_694_0 & i_13_124_4329_0) | (~i_13_124_4312_0 & ~i_13_124_4329_0) | (i_13_124_3532_0 & ~i_13_124_4331_0) | (i_13_124_2538_0 & ~i_13_124_4513_0)));
endmodule



// Benchmark "kernel_13_125" written by ABC on Sun Jul 19 10:47:10 2020

module kernel_13_125 ( 
    i_13_125_52_0, i_13_125_71_0, i_13_125_80_0, i_13_125_140_0,
    i_13_125_232_0, i_13_125_323_0, i_13_125_419_0, i_13_125_448_0,
    i_13_125_521_0, i_13_125_526_0, i_13_125_539_0, i_13_125_557_0,
    i_13_125_629_0, i_13_125_646_0, i_13_125_647_0, i_13_125_681_0,
    i_13_125_683_0, i_13_125_698_0, i_13_125_718_0, i_13_125_745_0,
    i_13_125_814_0, i_13_125_823_0, i_13_125_827_0, i_13_125_871_0,
    i_13_125_872_0, i_13_125_985_0, i_13_125_1066_0, i_13_125_1075_0,
    i_13_125_1103_0, i_13_125_1133_0, i_13_125_1214_0, i_13_125_1219_0,
    i_13_125_1398_0, i_13_125_1430_0, i_13_125_1454_0, i_13_125_1510_0,
    i_13_125_1511_0, i_13_125_1529_0, i_13_125_1538_0, i_13_125_1664_0,
    i_13_125_1668_0, i_13_125_1673_0, i_13_125_1736_0, i_13_125_1750_0,
    i_13_125_1798_0, i_13_125_1799_0, i_13_125_1835_0, i_13_125_1889_0,
    i_13_125_1898_0, i_13_125_1912_0, i_13_125_1948_0, i_13_125_2046_0,
    i_13_125_2110_0, i_13_125_2181_0, i_13_125_2236_0, i_13_125_2555_0,
    i_13_125_2561_0, i_13_125_2680_0, i_13_125_2725_0, i_13_125_2726_0,
    i_13_125_2748_0, i_13_125_2851_0, i_13_125_2852_0, i_13_125_2884_0,
    i_13_125_2885_0, i_13_125_2938_0, i_13_125_3094_0, i_13_125_3243_0,
    i_13_125_3265_0, i_13_125_3381_0, i_13_125_3392_0, i_13_125_3541_0,
    i_13_125_3597_0, i_13_125_3742_0, i_13_125_3743_0, i_13_125_3759_0,
    i_13_125_3797_0, i_13_125_3821_0, i_13_125_3895_0, i_13_125_3896_0,
    i_13_125_3931_0, i_13_125_3994_0, i_13_125_4040_0, i_13_125_4063_0,
    i_13_125_4084_0, i_13_125_4190_0, i_13_125_4193_0, i_13_125_4219_0,
    i_13_125_4297_0, i_13_125_4298_0, i_13_125_4301_0, i_13_125_4325_0,
    i_13_125_4342_0, i_13_125_4377_0, i_13_125_4399_0, i_13_125_4400_0,
    i_13_125_4436_0, i_13_125_4597_0, i_13_125_4598_0, i_13_125_4607_0,
    o_13_125_0_0  );
  input  i_13_125_52_0, i_13_125_71_0, i_13_125_80_0, i_13_125_140_0,
    i_13_125_232_0, i_13_125_323_0, i_13_125_419_0, i_13_125_448_0,
    i_13_125_521_0, i_13_125_526_0, i_13_125_539_0, i_13_125_557_0,
    i_13_125_629_0, i_13_125_646_0, i_13_125_647_0, i_13_125_681_0,
    i_13_125_683_0, i_13_125_698_0, i_13_125_718_0, i_13_125_745_0,
    i_13_125_814_0, i_13_125_823_0, i_13_125_827_0, i_13_125_871_0,
    i_13_125_872_0, i_13_125_985_0, i_13_125_1066_0, i_13_125_1075_0,
    i_13_125_1103_0, i_13_125_1133_0, i_13_125_1214_0, i_13_125_1219_0,
    i_13_125_1398_0, i_13_125_1430_0, i_13_125_1454_0, i_13_125_1510_0,
    i_13_125_1511_0, i_13_125_1529_0, i_13_125_1538_0, i_13_125_1664_0,
    i_13_125_1668_0, i_13_125_1673_0, i_13_125_1736_0, i_13_125_1750_0,
    i_13_125_1798_0, i_13_125_1799_0, i_13_125_1835_0, i_13_125_1889_0,
    i_13_125_1898_0, i_13_125_1912_0, i_13_125_1948_0, i_13_125_2046_0,
    i_13_125_2110_0, i_13_125_2181_0, i_13_125_2236_0, i_13_125_2555_0,
    i_13_125_2561_0, i_13_125_2680_0, i_13_125_2725_0, i_13_125_2726_0,
    i_13_125_2748_0, i_13_125_2851_0, i_13_125_2852_0, i_13_125_2884_0,
    i_13_125_2885_0, i_13_125_2938_0, i_13_125_3094_0, i_13_125_3243_0,
    i_13_125_3265_0, i_13_125_3381_0, i_13_125_3392_0, i_13_125_3541_0,
    i_13_125_3597_0, i_13_125_3742_0, i_13_125_3743_0, i_13_125_3759_0,
    i_13_125_3797_0, i_13_125_3821_0, i_13_125_3895_0, i_13_125_3896_0,
    i_13_125_3931_0, i_13_125_3994_0, i_13_125_4040_0, i_13_125_4063_0,
    i_13_125_4084_0, i_13_125_4190_0, i_13_125_4193_0, i_13_125_4219_0,
    i_13_125_4297_0, i_13_125_4298_0, i_13_125_4301_0, i_13_125_4325_0,
    i_13_125_4342_0, i_13_125_4377_0, i_13_125_4399_0, i_13_125_4400_0,
    i_13_125_4436_0, i_13_125_4597_0, i_13_125_4598_0, i_13_125_4607_0;
  output o_13_125_0_0;
  assign o_13_125_0_0 = ~((~i_13_125_4399_0 & ((~i_13_125_232_0 & ~i_13_125_323_0 & ~i_13_125_1219_0) | (~i_13_125_2726_0 & ~i_13_125_2884_0))) | i_13_125_2181_0 | (~i_13_125_3094_0 & ~i_13_125_3742_0) | (i_13_125_3243_0 & ~i_13_125_4219_0));
endmodule



// Benchmark "kernel_13_126" written by ABC on Sun Jul 19 10:47:10 2020

module kernel_13_126 ( 
    i_13_126_34_0, i_13_126_121_0, i_13_126_126_0, i_13_126_191_0,
    i_13_126_205_0, i_13_126_231_0, i_13_126_324_0, i_13_126_416_0,
    i_13_126_493_0, i_13_126_494_0, i_13_126_529_0, i_13_126_534_0,
    i_13_126_538_0, i_13_126_576_0, i_13_126_602_0, i_13_126_715_0,
    i_13_126_728_0, i_13_126_782_0, i_13_126_832_0, i_13_126_841_0,
    i_13_126_930_0, i_13_126_1074_0, i_13_126_1096_0, i_13_126_1097_0,
    i_13_126_1204_0, i_13_126_1220_0, i_13_126_1304_0, i_13_126_1309_0,
    i_13_126_1474_0, i_13_126_1508_0, i_13_126_1627_0, i_13_126_1674_0,
    i_13_126_1723_0, i_13_126_1726_0, i_13_126_1727_0, i_13_126_1772_0,
    i_13_126_1784_0, i_13_126_1785_0, i_13_126_1786_0, i_13_126_1787_0,
    i_13_126_1790_0, i_13_126_1930_0, i_13_126_2056_0, i_13_126_2119_0,
    i_13_126_2123_0, i_13_126_2239_0, i_13_126_2248_0, i_13_126_2312_0,
    i_13_126_2340_0, i_13_126_2365_0, i_13_126_2461_0, i_13_126_2467_0,
    i_13_126_2501_0, i_13_126_2547_0, i_13_126_2646_0, i_13_126_2717_0,
    i_13_126_2898_0, i_13_126_2941_0, i_13_126_2942_0, i_13_126_3019_0,
    i_13_126_3023_0, i_13_126_3027_0, i_13_126_3034_0, i_13_126_3036_0,
    i_13_126_3104_0, i_13_126_3159_0, i_13_126_3160_0, i_13_126_3215_0,
    i_13_126_3254_0, i_13_126_3396_0, i_13_126_3409_0, i_13_126_3416_0,
    i_13_126_3506_0, i_13_126_3535_0, i_13_126_3616_0, i_13_126_3687_0,
    i_13_126_3703_0, i_13_126_3769_0, i_13_126_3794_0, i_13_126_3910_0,
    i_13_126_3951_0, i_13_126_3986_0, i_13_126_4008_0, i_13_126_4009_0,
    i_13_126_4036_0, i_13_126_4057_0, i_13_126_4063_0, i_13_126_4109_0,
    i_13_126_4193_0, i_13_126_4238_0, i_13_126_4261_0, i_13_126_4310_0,
    i_13_126_4328_0, i_13_126_4408_0, i_13_126_4416_0, i_13_126_4518_0,
    i_13_126_4519_0, i_13_126_4522_0, i_13_126_4523_0, i_13_126_4594_0,
    o_13_126_0_0  );
  input  i_13_126_34_0, i_13_126_121_0, i_13_126_126_0, i_13_126_191_0,
    i_13_126_205_0, i_13_126_231_0, i_13_126_324_0, i_13_126_416_0,
    i_13_126_493_0, i_13_126_494_0, i_13_126_529_0, i_13_126_534_0,
    i_13_126_538_0, i_13_126_576_0, i_13_126_602_0, i_13_126_715_0,
    i_13_126_728_0, i_13_126_782_0, i_13_126_832_0, i_13_126_841_0,
    i_13_126_930_0, i_13_126_1074_0, i_13_126_1096_0, i_13_126_1097_0,
    i_13_126_1204_0, i_13_126_1220_0, i_13_126_1304_0, i_13_126_1309_0,
    i_13_126_1474_0, i_13_126_1508_0, i_13_126_1627_0, i_13_126_1674_0,
    i_13_126_1723_0, i_13_126_1726_0, i_13_126_1727_0, i_13_126_1772_0,
    i_13_126_1784_0, i_13_126_1785_0, i_13_126_1786_0, i_13_126_1787_0,
    i_13_126_1790_0, i_13_126_1930_0, i_13_126_2056_0, i_13_126_2119_0,
    i_13_126_2123_0, i_13_126_2239_0, i_13_126_2248_0, i_13_126_2312_0,
    i_13_126_2340_0, i_13_126_2365_0, i_13_126_2461_0, i_13_126_2467_0,
    i_13_126_2501_0, i_13_126_2547_0, i_13_126_2646_0, i_13_126_2717_0,
    i_13_126_2898_0, i_13_126_2941_0, i_13_126_2942_0, i_13_126_3019_0,
    i_13_126_3023_0, i_13_126_3027_0, i_13_126_3034_0, i_13_126_3036_0,
    i_13_126_3104_0, i_13_126_3159_0, i_13_126_3160_0, i_13_126_3215_0,
    i_13_126_3254_0, i_13_126_3396_0, i_13_126_3409_0, i_13_126_3416_0,
    i_13_126_3506_0, i_13_126_3535_0, i_13_126_3616_0, i_13_126_3687_0,
    i_13_126_3703_0, i_13_126_3769_0, i_13_126_3794_0, i_13_126_3910_0,
    i_13_126_3951_0, i_13_126_3986_0, i_13_126_4008_0, i_13_126_4009_0,
    i_13_126_4036_0, i_13_126_4057_0, i_13_126_4063_0, i_13_126_4109_0,
    i_13_126_4193_0, i_13_126_4238_0, i_13_126_4261_0, i_13_126_4310_0,
    i_13_126_4328_0, i_13_126_4408_0, i_13_126_4416_0, i_13_126_4518_0,
    i_13_126_4519_0, i_13_126_4522_0, i_13_126_4523_0, i_13_126_4594_0;
  output o_13_126_0_0;
  assign o_13_126_0_0 = ~((~i_13_126_4057_0 & (i_13_126_4261_0 | (~i_13_126_2646_0 & ~i_13_126_2941_0))) | (~i_13_126_4328_0 & ((i_13_126_529_0 & ~i_13_126_538_0) | (~i_13_126_3535_0 & i_13_126_4036_0))) | (~i_13_126_494_0 & ~i_13_126_930_0 & ~i_13_126_3396_0 & ~i_13_126_4416_0));
endmodule



// Benchmark "kernel_13_127" written by ABC on Sun Jul 19 10:47:11 2020

module kernel_13_127 ( 
    i_13_127_4_0, i_13_127_38_0, i_13_127_64_0, i_13_127_65_0,
    i_13_127_73_0, i_13_127_74_0, i_13_127_76_0, i_13_127_208_0,
    i_13_127_226_0, i_13_127_229_0, i_13_127_308_0, i_13_127_355_0,
    i_13_127_356_0, i_13_127_469_0, i_13_127_470_0, i_13_127_509_0,
    i_13_127_533_0, i_13_127_541_0, i_13_127_668_0, i_13_127_676_0,
    i_13_127_677_0, i_13_127_829_0, i_13_127_839_0, i_13_127_887_0,
    i_13_127_1100_0, i_13_127_1144_0, i_13_127_1145_0, i_13_127_1192_0,
    i_13_127_1246_0, i_13_127_1279_0, i_13_127_1307_0, i_13_127_1397_0,
    i_13_127_1400_0, i_13_127_1408_0, i_13_127_1445_0, i_13_127_1505_0,
    i_13_127_1621_0, i_13_127_1720_0, i_13_127_1721_0, i_13_127_1724_0,
    i_13_127_1730_0, i_13_127_1777_0, i_13_127_1778_0, i_13_127_1792_0,
    i_13_127_1909_0, i_13_127_1919_0, i_13_127_1928_0, i_13_127_2027_0,
    i_13_127_2056_0, i_13_127_2057_0, i_13_127_2237_0, i_13_127_2281_0,
    i_13_127_2282_0, i_13_127_2318_0, i_13_127_2354_0, i_13_127_2378_0,
    i_13_127_2468_0, i_13_127_2512_0, i_13_127_2534_0, i_13_127_2639_0,
    i_13_127_2656_0, i_13_127_2674_0, i_13_127_2692_0, i_13_127_2693_0,
    i_13_127_2720_0, i_13_127_2875_0, i_13_127_2882_0, i_13_127_2908_0,
    i_13_127_2974_0, i_13_127_3025_0, i_13_127_3034_0, i_13_127_3062_0,
    i_13_127_3136_0, i_13_127_3242_0, i_13_127_3251_0, i_13_127_3254_0,
    i_13_127_3371_0, i_13_127_3529_0, i_13_127_3532_0, i_13_127_3533_0,
    i_13_127_3593_0, i_13_127_3596_0, i_13_127_3619_0, i_13_127_3620_0,
    i_13_127_3631_0, i_13_127_3794_0, i_13_127_3935_0, i_13_127_3965_0,
    i_13_127_3988_0, i_13_127_3989_0, i_13_127_4034_0, i_13_127_4124_0,
    i_13_127_4187_0, i_13_127_4213_0, i_13_127_4214_0, i_13_127_4330_0,
    i_13_127_4331_0, i_13_127_4405_0, i_13_127_4430_0, i_13_127_4591_0,
    o_13_127_0_0  );
  input  i_13_127_4_0, i_13_127_38_0, i_13_127_64_0, i_13_127_65_0,
    i_13_127_73_0, i_13_127_74_0, i_13_127_76_0, i_13_127_208_0,
    i_13_127_226_0, i_13_127_229_0, i_13_127_308_0, i_13_127_355_0,
    i_13_127_356_0, i_13_127_469_0, i_13_127_470_0, i_13_127_509_0,
    i_13_127_533_0, i_13_127_541_0, i_13_127_668_0, i_13_127_676_0,
    i_13_127_677_0, i_13_127_829_0, i_13_127_839_0, i_13_127_887_0,
    i_13_127_1100_0, i_13_127_1144_0, i_13_127_1145_0, i_13_127_1192_0,
    i_13_127_1246_0, i_13_127_1279_0, i_13_127_1307_0, i_13_127_1397_0,
    i_13_127_1400_0, i_13_127_1408_0, i_13_127_1445_0, i_13_127_1505_0,
    i_13_127_1621_0, i_13_127_1720_0, i_13_127_1721_0, i_13_127_1724_0,
    i_13_127_1730_0, i_13_127_1777_0, i_13_127_1778_0, i_13_127_1792_0,
    i_13_127_1909_0, i_13_127_1919_0, i_13_127_1928_0, i_13_127_2027_0,
    i_13_127_2056_0, i_13_127_2057_0, i_13_127_2237_0, i_13_127_2281_0,
    i_13_127_2282_0, i_13_127_2318_0, i_13_127_2354_0, i_13_127_2378_0,
    i_13_127_2468_0, i_13_127_2512_0, i_13_127_2534_0, i_13_127_2639_0,
    i_13_127_2656_0, i_13_127_2674_0, i_13_127_2692_0, i_13_127_2693_0,
    i_13_127_2720_0, i_13_127_2875_0, i_13_127_2882_0, i_13_127_2908_0,
    i_13_127_2974_0, i_13_127_3025_0, i_13_127_3034_0, i_13_127_3062_0,
    i_13_127_3136_0, i_13_127_3242_0, i_13_127_3251_0, i_13_127_3254_0,
    i_13_127_3371_0, i_13_127_3529_0, i_13_127_3532_0, i_13_127_3533_0,
    i_13_127_3593_0, i_13_127_3596_0, i_13_127_3619_0, i_13_127_3620_0,
    i_13_127_3631_0, i_13_127_3794_0, i_13_127_3935_0, i_13_127_3965_0,
    i_13_127_3988_0, i_13_127_3989_0, i_13_127_4034_0, i_13_127_4124_0,
    i_13_127_4187_0, i_13_127_4213_0, i_13_127_4214_0, i_13_127_4330_0,
    i_13_127_4331_0, i_13_127_4405_0, i_13_127_4430_0, i_13_127_4591_0;
  output o_13_127_0_0;
  assign o_13_127_0_0 = ~(~i_13_127_469_0 | (~i_13_127_1397_0 & ~i_13_127_2693_0));
endmodule



// Benchmark "kernel_13_128" written by ABC on Sun Jul 19 10:47:12 2020

module kernel_13_128 ( 
    i_13_128_101_0, i_13_128_196_0, i_13_128_340_0, i_13_128_379_0,
    i_13_128_380_0, i_13_128_452_0, i_13_128_454_0, i_13_128_504_0,
    i_13_128_553_0, i_13_128_623_0, i_13_128_825_0, i_13_128_928_0,
    i_13_128_985_0, i_13_128_1063_0, i_13_128_1081_0, i_13_128_1082_0,
    i_13_128_1232_0, i_13_128_1297_0, i_13_128_1298_0, i_13_128_1320_0,
    i_13_128_1342_0, i_13_128_1410_0, i_13_128_1411_0, i_13_128_1412_0,
    i_13_128_1489_0, i_13_128_1491_0, i_13_128_1499_0, i_13_128_1502_0,
    i_13_128_1516_0, i_13_128_1517_0, i_13_128_1553_0, i_13_128_1554_0,
    i_13_128_1566_0, i_13_128_1627_0, i_13_128_1637_0, i_13_128_1801_0,
    i_13_128_1810_0, i_13_128_1926_0, i_13_128_1959_0, i_13_128_1990_0,
    i_13_128_2002_0, i_13_128_2107_0, i_13_128_2116_0, i_13_128_2134_0,
    i_13_128_2135_0, i_13_128_2201_0, i_13_128_2233_0, i_13_128_2234_0,
    i_13_128_2237_0, i_13_128_2294_0, i_13_128_2401_0, i_13_128_2461_0,
    i_13_128_2463_0, i_13_128_2515_0, i_13_128_2535_0, i_13_128_2572_0,
    i_13_128_2618_0, i_13_128_2934_0, i_13_128_2935_0, i_13_128_2936_0,
    i_13_128_2939_0, i_13_128_2977_0, i_13_128_3039_0, i_13_128_3172_0,
    i_13_128_3174_0, i_13_128_3218_0, i_13_128_3259_0, i_13_128_3285_0,
    i_13_128_3287_0, i_13_128_3339_0, i_13_128_3340_0, i_13_128_3341_0,
    i_13_128_3385_0, i_13_128_3421_0, i_13_128_3464_0, i_13_128_3521_0,
    i_13_128_3536_0, i_13_128_3579_0, i_13_128_3865_0, i_13_128_3877_0,
    i_13_128_3905_0, i_13_128_3912_0, i_13_128_4012_0, i_13_128_4013_0,
    i_13_128_4043_0, i_13_128_4051_0, i_13_128_4087_0, i_13_128_4162_0,
    i_13_128_4189_0, i_13_128_4266_0, i_13_128_4267_0, i_13_128_4271_0,
    i_13_128_4362_0, i_13_128_4393_0, i_13_128_4394_0, i_13_128_4396_0,
    i_13_128_4414_0, i_13_128_4443_0, i_13_128_4531_0, i_13_128_4594_0,
    o_13_128_0_0  );
  input  i_13_128_101_0, i_13_128_196_0, i_13_128_340_0, i_13_128_379_0,
    i_13_128_380_0, i_13_128_452_0, i_13_128_454_0, i_13_128_504_0,
    i_13_128_553_0, i_13_128_623_0, i_13_128_825_0, i_13_128_928_0,
    i_13_128_985_0, i_13_128_1063_0, i_13_128_1081_0, i_13_128_1082_0,
    i_13_128_1232_0, i_13_128_1297_0, i_13_128_1298_0, i_13_128_1320_0,
    i_13_128_1342_0, i_13_128_1410_0, i_13_128_1411_0, i_13_128_1412_0,
    i_13_128_1489_0, i_13_128_1491_0, i_13_128_1499_0, i_13_128_1502_0,
    i_13_128_1516_0, i_13_128_1517_0, i_13_128_1553_0, i_13_128_1554_0,
    i_13_128_1566_0, i_13_128_1627_0, i_13_128_1637_0, i_13_128_1801_0,
    i_13_128_1810_0, i_13_128_1926_0, i_13_128_1959_0, i_13_128_1990_0,
    i_13_128_2002_0, i_13_128_2107_0, i_13_128_2116_0, i_13_128_2134_0,
    i_13_128_2135_0, i_13_128_2201_0, i_13_128_2233_0, i_13_128_2234_0,
    i_13_128_2237_0, i_13_128_2294_0, i_13_128_2401_0, i_13_128_2461_0,
    i_13_128_2463_0, i_13_128_2515_0, i_13_128_2535_0, i_13_128_2572_0,
    i_13_128_2618_0, i_13_128_2934_0, i_13_128_2935_0, i_13_128_2936_0,
    i_13_128_2939_0, i_13_128_2977_0, i_13_128_3039_0, i_13_128_3172_0,
    i_13_128_3174_0, i_13_128_3218_0, i_13_128_3259_0, i_13_128_3285_0,
    i_13_128_3287_0, i_13_128_3339_0, i_13_128_3340_0, i_13_128_3341_0,
    i_13_128_3385_0, i_13_128_3421_0, i_13_128_3464_0, i_13_128_3521_0,
    i_13_128_3536_0, i_13_128_3579_0, i_13_128_3865_0, i_13_128_3877_0,
    i_13_128_3905_0, i_13_128_3912_0, i_13_128_4012_0, i_13_128_4013_0,
    i_13_128_4043_0, i_13_128_4051_0, i_13_128_4087_0, i_13_128_4162_0,
    i_13_128_4189_0, i_13_128_4266_0, i_13_128_4267_0, i_13_128_4271_0,
    i_13_128_4362_0, i_13_128_4393_0, i_13_128_4394_0, i_13_128_4396_0,
    i_13_128_4414_0, i_13_128_4443_0, i_13_128_4531_0, i_13_128_4594_0;
  output o_13_128_0_0;
  assign o_13_128_0_0 = ~((i_13_128_3865_0 & ((~i_13_128_3340_0 & ~i_13_128_3341_0 & ~i_13_128_4267_0) | (~i_13_128_2233_0 & ~i_13_128_4043_0 & ~i_13_128_4271_0))) | (~i_13_128_1297_0 & ~i_13_128_4271_0) | (~i_13_128_1990_0 & ~i_13_128_2936_0) | (~i_13_128_928_0 & i_13_128_4414_0));
endmodule



// Benchmark "kernel_13_129" written by ABC on Sun Jul 19 10:47:13 2020

module kernel_13_129 ( 
    i_13_129_116_0, i_13_129_121_0, i_13_129_122_0, i_13_129_139_0,
    i_13_129_173_0, i_13_129_175_0, i_13_129_226_0, i_13_129_229_0,
    i_13_129_280_0, i_13_129_281_0, i_13_129_311_0, i_13_129_319_0,
    i_13_129_337_0, i_13_129_373_0, i_13_129_416_0, i_13_129_523_0,
    i_13_129_526_0, i_13_129_563_0, i_13_129_590_0, i_13_129_658_0,
    i_13_129_733_0, i_13_129_847_0, i_13_129_848_0, i_13_129_850_0,
    i_13_129_851_0, i_13_129_938_0, i_13_129_986_0, i_13_129_1073_0,
    i_13_129_1201_0, i_13_129_1225_0, i_13_129_1280_0, i_13_129_1306_0,
    i_13_129_1345_0, i_13_129_1471_0, i_13_129_1549_0, i_13_129_1550_0,
    i_13_129_1712_0, i_13_129_1723_0, i_13_129_1751_0, i_13_129_1783_0,
    i_13_129_1855_0, i_13_129_1857_0, i_13_129_1858_0, i_13_129_1859_0,
    i_13_129_1901_0, i_13_129_1928_0, i_13_129_2125_0, i_13_129_2126_0,
    i_13_129_2169_0, i_13_129_2209_0, i_13_129_2238_0, i_13_129_2468_0,
    i_13_129_2510_0, i_13_129_2570_0, i_13_129_2692_0, i_13_129_2713_0,
    i_13_129_3001_0, i_13_129_3007_0, i_13_129_3008_0, i_13_129_3010_0,
    i_13_129_3037_0, i_13_129_3128_0, i_13_129_3133_0, i_13_129_3196_0,
    i_13_129_3217_0, i_13_129_3262_0, i_13_129_3269_0, i_13_129_3394_0,
    i_13_129_3412_0, i_13_129_3439_0, i_13_129_3442_0, i_13_129_3484_0,
    i_13_129_3485_0, i_13_129_3538_0, i_13_129_3539_0, i_13_129_3575_0,
    i_13_129_3685_0, i_13_129_3686_0, i_13_129_3820_0, i_13_129_3854_0,
    i_13_129_3862_0, i_13_129_3863_0, i_13_129_3868_0, i_13_129_3890_0,
    i_13_129_3908_0, i_13_129_4045_0, i_13_129_4106_0, i_13_129_4250_0,
    i_13_129_4253_0, i_13_129_4259_0, i_13_129_4276_0, i_13_129_4352_0,
    i_13_129_4369_0, i_13_129_4376_0, i_13_129_4379_0, i_13_129_4411_0,
    i_13_129_4522_0, i_13_129_4523_0, i_13_129_4531_0, i_13_129_4595_0,
    o_13_129_0_0  );
  input  i_13_129_116_0, i_13_129_121_0, i_13_129_122_0, i_13_129_139_0,
    i_13_129_173_0, i_13_129_175_0, i_13_129_226_0, i_13_129_229_0,
    i_13_129_280_0, i_13_129_281_0, i_13_129_311_0, i_13_129_319_0,
    i_13_129_337_0, i_13_129_373_0, i_13_129_416_0, i_13_129_523_0,
    i_13_129_526_0, i_13_129_563_0, i_13_129_590_0, i_13_129_658_0,
    i_13_129_733_0, i_13_129_847_0, i_13_129_848_0, i_13_129_850_0,
    i_13_129_851_0, i_13_129_938_0, i_13_129_986_0, i_13_129_1073_0,
    i_13_129_1201_0, i_13_129_1225_0, i_13_129_1280_0, i_13_129_1306_0,
    i_13_129_1345_0, i_13_129_1471_0, i_13_129_1549_0, i_13_129_1550_0,
    i_13_129_1712_0, i_13_129_1723_0, i_13_129_1751_0, i_13_129_1783_0,
    i_13_129_1855_0, i_13_129_1857_0, i_13_129_1858_0, i_13_129_1859_0,
    i_13_129_1901_0, i_13_129_1928_0, i_13_129_2125_0, i_13_129_2126_0,
    i_13_129_2169_0, i_13_129_2209_0, i_13_129_2238_0, i_13_129_2468_0,
    i_13_129_2510_0, i_13_129_2570_0, i_13_129_2692_0, i_13_129_2713_0,
    i_13_129_3001_0, i_13_129_3007_0, i_13_129_3008_0, i_13_129_3010_0,
    i_13_129_3037_0, i_13_129_3128_0, i_13_129_3133_0, i_13_129_3196_0,
    i_13_129_3217_0, i_13_129_3262_0, i_13_129_3269_0, i_13_129_3394_0,
    i_13_129_3412_0, i_13_129_3439_0, i_13_129_3442_0, i_13_129_3484_0,
    i_13_129_3485_0, i_13_129_3538_0, i_13_129_3539_0, i_13_129_3575_0,
    i_13_129_3685_0, i_13_129_3686_0, i_13_129_3820_0, i_13_129_3854_0,
    i_13_129_3862_0, i_13_129_3863_0, i_13_129_3868_0, i_13_129_3890_0,
    i_13_129_3908_0, i_13_129_4045_0, i_13_129_4106_0, i_13_129_4250_0,
    i_13_129_4253_0, i_13_129_4259_0, i_13_129_4276_0, i_13_129_4352_0,
    i_13_129_4369_0, i_13_129_4376_0, i_13_129_4379_0, i_13_129_4411_0,
    i_13_129_4522_0, i_13_129_4523_0, i_13_129_4531_0, i_13_129_4595_0;
  output o_13_129_0_0;
  assign o_13_129_0_0 = ~(~i_13_129_3010_0 | (~i_13_129_3538_0 & ~i_13_129_3890_0 & ~i_13_129_4376_0) | (i_13_129_121_0 & i_13_129_229_0 & ~i_13_129_4253_0) | (i_13_129_1471_0 & ~i_13_129_3539_0 & ~i_13_129_4045_0) | (~i_13_129_1858_0 & ~i_13_129_2126_0 & ~i_13_129_3854_0));
endmodule



// Benchmark "kernel_13_130" written by ABC on Sun Jul 19 10:47:14 2020

module kernel_13_130 ( 
    i_13_130_73_0, i_13_130_77_0, i_13_130_95_0, i_13_130_121_0,
    i_13_130_122_0, i_13_130_126_0, i_13_130_184_0, i_13_130_207_0,
    i_13_130_208_0, i_13_130_238_0, i_13_130_243_0, i_13_130_297_0,
    i_13_130_415_0, i_13_130_418_0, i_13_130_473_0, i_13_130_516_0,
    i_13_130_517_0, i_13_130_520_0, i_13_130_697_0, i_13_130_721_0,
    i_13_130_850_0, i_13_130_853_0, i_13_130_855_0, i_13_130_933_0,
    i_13_130_936_0, i_13_130_937_0, i_13_130_949_0, i_13_130_985_0,
    i_13_130_990_0, i_13_130_1071_0, i_13_130_1080_0, i_13_130_1128_0,
    i_13_130_1203_0, i_13_130_1209_0, i_13_130_1222_0, i_13_130_1252_0,
    i_13_130_1305_0, i_13_130_1317_0, i_13_130_1404_0, i_13_130_1521_0,
    i_13_130_1522_0, i_13_130_1548_0, i_13_130_1549_0, i_13_130_1552_0,
    i_13_130_1553_0, i_13_130_1602_0, i_13_130_1603_0, i_13_130_1699_0,
    i_13_130_1700_0, i_13_130_1711_0, i_13_130_1719_0, i_13_130_1723_0,
    i_13_130_1750_0, i_13_130_1786_0, i_13_130_1840_0, i_13_130_1843_0,
    i_13_130_1943_0, i_13_130_1957_0, i_13_130_1962_0, i_13_130_2033_0,
    i_13_130_2101_0, i_13_130_2113_0, i_13_130_2124_0, i_13_130_2125_0,
    i_13_130_2244_0, i_13_130_2248_0, i_13_130_2263_0, i_13_130_2333_0,
    i_13_130_2365_0, i_13_130_2442_0, i_13_130_2539_0, i_13_130_2581_0,
    i_13_130_2969_0, i_13_130_3007_0, i_13_130_3009_0, i_13_130_3040_0,
    i_13_130_3163_0, i_13_130_3268_0, i_13_130_3456_0, i_13_130_3461_0,
    i_13_130_3541_0, i_13_130_3577_0, i_13_130_3635_0, i_13_130_3739_0,
    i_13_130_3791_0, i_13_130_3796_0, i_13_130_3854_0, i_13_130_3898_0,
    i_13_130_3919_0, i_13_130_3921_0, i_13_130_3971_0, i_13_130_4078_0,
    i_13_130_4101_0, i_13_130_4261_0, i_13_130_4321_0, i_13_130_4334_0,
    i_13_130_4363_0, i_13_130_4380_0, i_13_130_4472_0, i_13_130_4509_0,
    o_13_130_0_0  );
  input  i_13_130_73_0, i_13_130_77_0, i_13_130_95_0, i_13_130_121_0,
    i_13_130_122_0, i_13_130_126_0, i_13_130_184_0, i_13_130_207_0,
    i_13_130_208_0, i_13_130_238_0, i_13_130_243_0, i_13_130_297_0,
    i_13_130_415_0, i_13_130_418_0, i_13_130_473_0, i_13_130_516_0,
    i_13_130_517_0, i_13_130_520_0, i_13_130_697_0, i_13_130_721_0,
    i_13_130_850_0, i_13_130_853_0, i_13_130_855_0, i_13_130_933_0,
    i_13_130_936_0, i_13_130_937_0, i_13_130_949_0, i_13_130_985_0,
    i_13_130_990_0, i_13_130_1071_0, i_13_130_1080_0, i_13_130_1128_0,
    i_13_130_1203_0, i_13_130_1209_0, i_13_130_1222_0, i_13_130_1252_0,
    i_13_130_1305_0, i_13_130_1317_0, i_13_130_1404_0, i_13_130_1521_0,
    i_13_130_1522_0, i_13_130_1548_0, i_13_130_1549_0, i_13_130_1552_0,
    i_13_130_1553_0, i_13_130_1602_0, i_13_130_1603_0, i_13_130_1699_0,
    i_13_130_1700_0, i_13_130_1711_0, i_13_130_1719_0, i_13_130_1723_0,
    i_13_130_1750_0, i_13_130_1786_0, i_13_130_1840_0, i_13_130_1843_0,
    i_13_130_1943_0, i_13_130_1957_0, i_13_130_1962_0, i_13_130_2033_0,
    i_13_130_2101_0, i_13_130_2113_0, i_13_130_2124_0, i_13_130_2125_0,
    i_13_130_2244_0, i_13_130_2248_0, i_13_130_2263_0, i_13_130_2333_0,
    i_13_130_2365_0, i_13_130_2442_0, i_13_130_2539_0, i_13_130_2581_0,
    i_13_130_2969_0, i_13_130_3007_0, i_13_130_3009_0, i_13_130_3040_0,
    i_13_130_3163_0, i_13_130_3268_0, i_13_130_3456_0, i_13_130_3461_0,
    i_13_130_3541_0, i_13_130_3577_0, i_13_130_3635_0, i_13_130_3739_0,
    i_13_130_3791_0, i_13_130_3796_0, i_13_130_3854_0, i_13_130_3898_0,
    i_13_130_3919_0, i_13_130_3921_0, i_13_130_3971_0, i_13_130_4078_0,
    i_13_130_4101_0, i_13_130_4261_0, i_13_130_4321_0, i_13_130_4334_0,
    i_13_130_4363_0, i_13_130_4380_0, i_13_130_4472_0, i_13_130_4509_0;
  output o_13_130_0_0;
  assign o_13_130_0_0 = ~((~i_13_130_517_0 & ((~i_13_130_1252_0 & ~i_13_130_1602_0 & ~i_13_130_2125_0) | (~i_13_130_1548_0 & ~i_13_130_4261_0))) | ~i_13_130_1549_0 | (~i_13_130_73_0 & i_13_130_1553_0 & ~i_13_130_1750_0 & ~i_13_130_3007_0));
endmodule



// Benchmark "kernel_13_131" written by ABC on Sun Jul 19 10:47:15 2020

module kernel_13_131 ( 
    i_13_131_37_0, i_13_131_91_0, i_13_131_92_0, i_13_131_94_0,
    i_13_131_95_0, i_13_131_112_0, i_13_131_230_0, i_13_131_238_0,
    i_13_131_256_0, i_13_131_260_0, i_13_131_263_0, i_13_131_274_0,
    i_13_131_277_0, i_13_131_315_0, i_13_131_316_0, i_13_131_326_0,
    i_13_131_364_0, i_13_131_374_0, i_13_131_518_0, i_13_131_607_0,
    i_13_131_670_0, i_13_131_694_0, i_13_131_697_0, i_13_131_698_0,
    i_13_131_778_0, i_13_131_832_0, i_13_131_943_0, i_13_131_976_0,
    i_13_131_977_0, i_13_131_979_0, i_13_131_1076_0, i_13_131_1082_0,
    i_13_131_1231_0, i_13_131_1262_0, i_13_131_1315_0, i_13_131_1336_0,
    i_13_131_1427_0, i_13_131_1433_0, i_13_131_1444_0, i_13_131_1468_0,
    i_13_131_1469_0, i_13_131_1512_0, i_13_131_1516_0, i_13_131_1669_0,
    i_13_131_1840_0, i_13_131_1861_0, i_13_131_1862_0, i_13_131_1886_0,
    i_13_131_1918_0, i_13_131_2140_0, i_13_131_2147_0, i_13_131_2198_0,
    i_13_131_2245_0, i_13_131_2298_0, i_13_131_2434_0, i_13_131_2521_0,
    i_13_131_2647_0, i_13_131_2651_0, i_13_131_2677_0, i_13_131_2702_0,
    i_13_131_2734_0, i_13_131_2735_0, i_13_131_2740_0, i_13_131_2899_0,
    i_13_131_2983_0, i_13_131_3143_0, i_13_131_3172_0, i_13_131_3208_0,
    i_13_131_3313_0, i_13_131_3341_0, i_13_131_3370_0, i_13_131_3373_0,
    i_13_131_3430_0, i_13_131_3448_0, i_13_131_3452_0, i_13_131_3593_0,
    i_13_131_3763_0, i_13_131_3806_0, i_13_131_3871_0, i_13_131_3907_0,
    i_13_131_4097_0, i_13_131_4118_0, i_13_131_4162_0, i_13_131_4177_0,
    i_13_131_4185_0, i_13_131_4278_0, i_13_131_4307_0, i_13_131_4351_0,
    i_13_131_4379_0, i_13_131_4387_0, i_13_131_4388_0, i_13_131_4390_0,
    i_13_131_4393_0, i_13_131_4441_0, i_13_131_4447_0, i_13_131_4448_0,
    i_13_131_4451_0, i_13_131_4518_0, i_13_131_4523_0, i_13_131_4567_0,
    o_13_131_0_0  );
  input  i_13_131_37_0, i_13_131_91_0, i_13_131_92_0, i_13_131_94_0,
    i_13_131_95_0, i_13_131_112_0, i_13_131_230_0, i_13_131_238_0,
    i_13_131_256_0, i_13_131_260_0, i_13_131_263_0, i_13_131_274_0,
    i_13_131_277_0, i_13_131_315_0, i_13_131_316_0, i_13_131_326_0,
    i_13_131_364_0, i_13_131_374_0, i_13_131_518_0, i_13_131_607_0,
    i_13_131_670_0, i_13_131_694_0, i_13_131_697_0, i_13_131_698_0,
    i_13_131_778_0, i_13_131_832_0, i_13_131_943_0, i_13_131_976_0,
    i_13_131_977_0, i_13_131_979_0, i_13_131_1076_0, i_13_131_1082_0,
    i_13_131_1231_0, i_13_131_1262_0, i_13_131_1315_0, i_13_131_1336_0,
    i_13_131_1427_0, i_13_131_1433_0, i_13_131_1444_0, i_13_131_1468_0,
    i_13_131_1469_0, i_13_131_1512_0, i_13_131_1516_0, i_13_131_1669_0,
    i_13_131_1840_0, i_13_131_1861_0, i_13_131_1862_0, i_13_131_1886_0,
    i_13_131_1918_0, i_13_131_2140_0, i_13_131_2147_0, i_13_131_2198_0,
    i_13_131_2245_0, i_13_131_2298_0, i_13_131_2434_0, i_13_131_2521_0,
    i_13_131_2647_0, i_13_131_2651_0, i_13_131_2677_0, i_13_131_2702_0,
    i_13_131_2734_0, i_13_131_2735_0, i_13_131_2740_0, i_13_131_2899_0,
    i_13_131_2983_0, i_13_131_3143_0, i_13_131_3172_0, i_13_131_3208_0,
    i_13_131_3313_0, i_13_131_3341_0, i_13_131_3370_0, i_13_131_3373_0,
    i_13_131_3430_0, i_13_131_3448_0, i_13_131_3452_0, i_13_131_3593_0,
    i_13_131_3763_0, i_13_131_3806_0, i_13_131_3871_0, i_13_131_3907_0,
    i_13_131_4097_0, i_13_131_4118_0, i_13_131_4162_0, i_13_131_4177_0,
    i_13_131_4185_0, i_13_131_4278_0, i_13_131_4307_0, i_13_131_4351_0,
    i_13_131_4379_0, i_13_131_4387_0, i_13_131_4388_0, i_13_131_4390_0,
    i_13_131_4393_0, i_13_131_4441_0, i_13_131_4447_0, i_13_131_4448_0,
    i_13_131_4451_0, i_13_131_4518_0, i_13_131_4523_0, i_13_131_4567_0;
  output o_13_131_0_0;
  assign o_13_131_0_0 = ~((~i_13_131_256_0 & ((~i_13_131_2740_0 & i_13_131_3208_0) | (~i_13_131_698_0 & ~i_13_131_1886_0 & ~i_13_131_4448_0))) | (~i_13_131_274_0 & ((~i_13_131_1076_0 & ~i_13_131_1427_0 & ~i_13_131_2647_0 & i_13_131_2677_0) | (~i_13_131_1468_0 & i_13_131_3208_0 & ~i_13_131_3452_0))) | (~i_13_131_1262_0 & ((i_13_131_1840_0 & ~i_13_131_3452_0) | (~i_13_131_230_0 & ~i_13_131_1468_0 & ~i_13_131_4379_0))) | (i_13_131_2140_0 & i_13_131_2434_0) | (~i_13_131_698_0 & i_13_131_4351_0) | (~i_13_131_238_0 & i_13_131_2677_0 & ~i_13_131_3313_0 & ~i_13_131_3341_0 & ~i_13_131_4307_0 & ~i_13_131_4393_0) | (i_13_131_112_0 & ~i_13_131_2147_0 & ~i_13_131_2647_0 & ~i_13_131_3448_0 & ~i_13_131_4448_0) | (i_13_131_274_0 & ~i_13_131_694_0 & i_13_131_4185_0 & i_13_131_4567_0));
endmodule



// Benchmark "kernel_13_132" written by ABC on Sun Jul 19 10:47:16 2020

module kernel_13_132 ( 
    i_13_132_46_0, i_13_132_78_0, i_13_132_103_0, i_13_132_154_0,
    i_13_132_245_0, i_13_132_379_0, i_13_132_411_0, i_13_132_421_0,
    i_13_132_443_0, i_13_132_450_0, i_13_132_451_0, i_13_132_460_0,
    i_13_132_461_0, i_13_132_552_0, i_13_132_658_0, i_13_132_661_0,
    i_13_132_698_0, i_13_132_820_0, i_13_132_897_0, i_13_132_940_0,
    i_13_132_1193_0, i_13_132_1251_0, i_13_132_1285_0, i_13_132_1297_0,
    i_13_132_1331_0, i_13_132_1342_0, i_13_132_1422_0, i_13_132_1432_0,
    i_13_132_1441_0, i_13_132_1442_0, i_13_132_1495_0, i_13_132_1567_0,
    i_13_132_1568_0, i_13_132_1601_0, i_13_132_1632_0, i_13_132_1633_0,
    i_13_132_1786_0, i_13_132_1801_0, i_13_132_1835_0, i_13_132_1858_0,
    i_13_132_1921_0, i_13_132_1928_0, i_13_132_1944_0, i_13_132_1945_0,
    i_13_132_1957_0, i_13_132_1959_0, i_13_132_2002_0, i_13_132_2098_0,
    i_13_132_2134_0, i_13_132_2135_0, i_13_132_2150_0, i_13_132_2197_0,
    i_13_132_2198_0, i_13_132_2278_0, i_13_132_2302_0, i_13_132_2316_0,
    i_13_132_2357_0, i_13_132_2380_0, i_13_132_2381_0, i_13_132_2405_0,
    i_13_132_2452_0, i_13_132_2544_0, i_13_132_2579_0, i_13_132_2614_0,
    i_13_132_2821_0, i_13_132_2983_0, i_13_132_2987_0, i_13_132_3010_0,
    i_13_132_3014_0, i_13_132_3017_0, i_13_132_3212_0, i_13_132_3268_0,
    i_13_132_3269_0, i_13_132_3341_0, i_13_132_3366_0, i_13_132_3375_0,
    i_13_132_3422_0, i_13_132_3485_0, i_13_132_3593_0, i_13_132_3727_0,
    i_13_132_3817_0, i_13_132_4015_0, i_13_132_4051_0, i_13_132_4086_0,
    i_13_132_4087_0, i_13_132_4208_0, i_13_132_4230_0, i_13_132_4231_0,
    i_13_132_4234_0, i_13_132_4249_0, i_13_132_4251_0, i_13_132_4252_0,
    i_13_132_4259_0, i_13_132_4261_0, i_13_132_4267_0, i_13_132_4268_0,
    i_13_132_4274_0, i_13_132_4393_0, i_13_132_4414_0, i_13_132_4447_0,
    o_13_132_0_0  );
  input  i_13_132_46_0, i_13_132_78_0, i_13_132_103_0, i_13_132_154_0,
    i_13_132_245_0, i_13_132_379_0, i_13_132_411_0, i_13_132_421_0,
    i_13_132_443_0, i_13_132_450_0, i_13_132_451_0, i_13_132_460_0,
    i_13_132_461_0, i_13_132_552_0, i_13_132_658_0, i_13_132_661_0,
    i_13_132_698_0, i_13_132_820_0, i_13_132_897_0, i_13_132_940_0,
    i_13_132_1193_0, i_13_132_1251_0, i_13_132_1285_0, i_13_132_1297_0,
    i_13_132_1331_0, i_13_132_1342_0, i_13_132_1422_0, i_13_132_1432_0,
    i_13_132_1441_0, i_13_132_1442_0, i_13_132_1495_0, i_13_132_1567_0,
    i_13_132_1568_0, i_13_132_1601_0, i_13_132_1632_0, i_13_132_1633_0,
    i_13_132_1786_0, i_13_132_1801_0, i_13_132_1835_0, i_13_132_1858_0,
    i_13_132_1921_0, i_13_132_1928_0, i_13_132_1944_0, i_13_132_1945_0,
    i_13_132_1957_0, i_13_132_1959_0, i_13_132_2002_0, i_13_132_2098_0,
    i_13_132_2134_0, i_13_132_2135_0, i_13_132_2150_0, i_13_132_2197_0,
    i_13_132_2198_0, i_13_132_2278_0, i_13_132_2302_0, i_13_132_2316_0,
    i_13_132_2357_0, i_13_132_2380_0, i_13_132_2381_0, i_13_132_2405_0,
    i_13_132_2452_0, i_13_132_2544_0, i_13_132_2579_0, i_13_132_2614_0,
    i_13_132_2821_0, i_13_132_2983_0, i_13_132_2987_0, i_13_132_3010_0,
    i_13_132_3014_0, i_13_132_3017_0, i_13_132_3212_0, i_13_132_3268_0,
    i_13_132_3269_0, i_13_132_3341_0, i_13_132_3366_0, i_13_132_3375_0,
    i_13_132_3422_0, i_13_132_3485_0, i_13_132_3593_0, i_13_132_3727_0,
    i_13_132_3817_0, i_13_132_4015_0, i_13_132_4051_0, i_13_132_4086_0,
    i_13_132_4087_0, i_13_132_4208_0, i_13_132_4230_0, i_13_132_4231_0,
    i_13_132_4234_0, i_13_132_4249_0, i_13_132_4251_0, i_13_132_4252_0,
    i_13_132_4259_0, i_13_132_4261_0, i_13_132_4267_0, i_13_132_4268_0,
    i_13_132_4274_0, i_13_132_4393_0, i_13_132_4414_0, i_13_132_4447_0;
  output o_13_132_0_0;
  assign o_13_132_0_0 = ~((~i_13_132_2614_0 & ~i_13_132_4268_0) | (~i_13_132_1567_0 & ~i_13_132_2198_0 & ~i_13_132_3817_0 & ~i_13_132_4447_0));
endmodule



// Benchmark "kernel_13_133" written by ABC on Sun Jul 19 10:47:16 2020

module kernel_13_133 ( 
    i_13_133_25_0, i_13_133_168_0, i_13_133_229_0, i_13_133_318_0,
    i_13_133_463_0, i_13_133_517_0, i_13_133_523_0, i_13_133_526_0,
    i_13_133_535_0, i_13_133_538_0, i_13_133_571_0, i_13_133_601_0,
    i_13_133_717_0, i_13_133_759_0, i_13_133_850_0, i_13_133_895_0,
    i_13_133_1018_0, i_13_133_1120_0, i_13_133_1144_0, i_13_133_1210_0,
    i_13_133_1219_0, i_13_133_1273_0, i_13_133_1279_0, i_13_133_1426_0,
    i_13_133_1495_0, i_13_133_1497_0, i_13_133_1498_0, i_13_133_1528_0,
    i_13_133_1549_0, i_13_133_1606_0, i_13_133_1630_0, i_13_133_1631_0,
    i_13_133_1632_0, i_13_133_2001_0, i_13_133_2197_0, i_13_133_2198_0,
    i_13_133_2200_0, i_13_133_2365_0, i_13_133_2384_0, i_13_133_2457_0,
    i_13_133_2538_0, i_13_133_2541_0, i_13_133_2542_0, i_13_133_2764_0,
    i_13_133_2765_0, i_13_133_2767_0, i_13_133_2919_0, i_13_133_2935_0,
    i_13_133_3010_0, i_13_133_3037_0, i_13_133_3052_0, i_13_133_3100_0,
    i_13_133_3108_0, i_13_133_3119_0, i_13_133_3122_0, i_13_133_3141_0,
    i_13_133_3163_0, i_13_133_3169_0, i_13_133_3247_0, i_13_133_3262_0,
    i_13_133_3342_0, i_13_133_3459_0, i_13_133_3460_0, i_13_133_3540_0,
    i_13_133_3541_0, i_13_133_3612_0, i_13_133_3666_0, i_13_133_3722_0,
    i_13_133_3726_0, i_13_133_3727_0, i_13_133_3729_0, i_13_133_3730_0,
    i_13_133_3731_0, i_13_133_3838_0, i_13_133_3855_0, i_13_133_3859_0,
    i_13_133_3907_0, i_13_133_3916_0, i_13_133_3996_0, i_13_133_4014_0,
    i_13_133_4059_0, i_13_133_4060_0, i_13_133_4081_0, i_13_133_4162_0,
    i_13_133_4189_0, i_13_133_4207_0, i_13_133_4208_0, i_13_133_4251_0,
    i_13_133_4252_0, i_13_133_4255_0, i_13_133_4260_0, i_13_133_4266_0,
    i_13_133_4311_0, i_13_133_4341_0, i_13_133_4353_0, i_13_133_4465_0,
    i_13_133_4530_0, i_13_133_4555_0, i_13_133_4600_0, i_13_133_4603_0,
    o_13_133_0_0  );
  input  i_13_133_25_0, i_13_133_168_0, i_13_133_229_0, i_13_133_318_0,
    i_13_133_463_0, i_13_133_517_0, i_13_133_523_0, i_13_133_526_0,
    i_13_133_535_0, i_13_133_538_0, i_13_133_571_0, i_13_133_601_0,
    i_13_133_717_0, i_13_133_759_0, i_13_133_850_0, i_13_133_895_0,
    i_13_133_1018_0, i_13_133_1120_0, i_13_133_1144_0, i_13_133_1210_0,
    i_13_133_1219_0, i_13_133_1273_0, i_13_133_1279_0, i_13_133_1426_0,
    i_13_133_1495_0, i_13_133_1497_0, i_13_133_1498_0, i_13_133_1528_0,
    i_13_133_1549_0, i_13_133_1606_0, i_13_133_1630_0, i_13_133_1631_0,
    i_13_133_1632_0, i_13_133_2001_0, i_13_133_2197_0, i_13_133_2198_0,
    i_13_133_2200_0, i_13_133_2365_0, i_13_133_2384_0, i_13_133_2457_0,
    i_13_133_2538_0, i_13_133_2541_0, i_13_133_2542_0, i_13_133_2764_0,
    i_13_133_2765_0, i_13_133_2767_0, i_13_133_2919_0, i_13_133_2935_0,
    i_13_133_3010_0, i_13_133_3037_0, i_13_133_3052_0, i_13_133_3100_0,
    i_13_133_3108_0, i_13_133_3119_0, i_13_133_3122_0, i_13_133_3141_0,
    i_13_133_3163_0, i_13_133_3169_0, i_13_133_3247_0, i_13_133_3262_0,
    i_13_133_3342_0, i_13_133_3459_0, i_13_133_3460_0, i_13_133_3540_0,
    i_13_133_3541_0, i_13_133_3612_0, i_13_133_3666_0, i_13_133_3722_0,
    i_13_133_3726_0, i_13_133_3727_0, i_13_133_3729_0, i_13_133_3730_0,
    i_13_133_3731_0, i_13_133_3838_0, i_13_133_3855_0, i_13_133_3859_0,
    i_13_133_3907_0, i_13_133_3916_0, i_13_133_3996_0, i_13_133_4014_0,
    i_13_133_4059_0, i_13_133_4060_0, i_13_133_4081_0, i_13_133_4162_0,
    i_13_133_4189_0, i_13_133_4207_0, i_13_133_4208_0, i_13_133_4251_0,
    i_13_133_4252_0, i_13_133_4255_0, i_13_133_4260_0, i_13_133_4266_0,
    i_13_133_4311_0, i_13_133_4341_0, i_13_133_4353_0, i_13_133_4465_0,
    i_13_133_4530_0, i_13_133_4555_0, i_13_133_4600_0, i_13_133_4603_0;
  output o_13_133_0_0;
  assign o_13_133_0_0 = ~((~i_13_133_3731_0 & ((~i_13_133_2200_0 & ~i_13_133_3729_0) | (~i_13_133_3108_0 & ~i_13_133_3459_0 & ~i_13_133_4311_0))) | (i_13_133_4255_0 & (~i_13_133_2767_0 | (i_13_133_3731_0 & ~i_13_133_4252_0))) | (i_13_133_1120_0 & ~i_13_133_1497_0) | (~i_13_133_523_0 & ~i_13_133_3247_0 & ~i_13_133_3855_0 & ~i_13_133_3859_0 & ~i_13_133_3916_0) | (i_13_133_1273_0 & ~i_13_133_2198_0 & ~i_13_133_3342_0 & ~i_13_133_4266_0) | (~i_13_133_517_0 & ~i_13_133_3460_0 & ~i_13_133_3541_0 & ~i_13_133_4311_0));
endmodule



// Benchmark "kernel_13_134" written by ABC on Sun Jul 19 10:47:17 2020

module kernel_13_134 ( 
    i_13_134_65_0, i_13_134_94_0, i_13_134_95_0, i_13_134_173_0,
    i_13_134_175_0, i_13_134_176_0, i_13_134_202_0, i_13_134_235_0,
    i_13_134_307_0, i_13_134_308_0, i_13_134_442_0, i_13_134_443_0,
    i_13_134_485_0, i_13_134_572_0, i_13_134_604_0, i_13_134_605_0,
    i_13_134_658_0, i_13_134_662_0, i_13_134_667_0, i_13_134_668_0,
    i_13_134_676_0, i_13_134_677_0, i_13_134_698_0, i_13_134_934_0,
    i_13_134_946_0, i_13_134_1066_0, i_13_134_1217_0, i_13_134_1267_0,
    i_13_134_1306_0, i_13_134_1310_0, i_13_134_1388_0, i_13_134_1499_0,
    i_13_134_1504_0, i_13_134_1505_0, i_13_134_1561_0, i_13_134_1621_0,
    i_13_134_1630_0, i_13_134_1670_0, i_13_134_1720_0, i_13_134_1730_0,
    i_13_134_1802_0, i_13_134_1837_0, i_13_134_1838_0, i_13_134_1840_0,
    i_13_134_1841_0, i_13_134_1904_0, i_13_134_2170_0, i_13_134_2173_0,
    i_13_134_2230_0, i_13_134_2422_0, i_13_134_2423_0, i_13_134_2424_0,
    i_13_134_2425_0, i_13_134_2426_0, i_13_134_2431_0, i_13_134_2432_0,
    i_13_134_2435_0, i_13_134_2503_0, i_13_134_2593_0, i_13_134_2674_0,
    i_13_134_2675_0, i_13_134_2677_0, i_13_134_2678_0, i_13_134_2702_0,
    i_13_134_2912_0, i_13_134_2950_0, i_13_134_2951_0, i_13_134_3142_0,
    i_13_134_3143_0, i_13_134_3145_0, i_13_134_3242_0, i_13_134_3260_0,
    i_13_134_3269_0, i_13_134_3304_0, i_13_134_3305_0, i_13_134_3421_0,
    i_13_134_3422_0, i_13_134_3424_0, i_13_134_3425_0, i_13_134_3446_0,
    i_13_134_3529_0, i_13_134_3592_0, i_13_134_3726_0, i_13_134_3871_0,
    i_13_134_4016_0, i_13_134_4018_0, i_13_134_4019_0, i_13_134_4078_0,
    i_13_134_4079_0, i_13_134_4249_0, i_13_134_4253_0, i_13_134_4258_0,
    i_13_134_4351_0, i_13_134_4430_0, i_13_134_4447_0, i_13_134_4541_0,
    i_13_134_4555_0, i_13_134_4556_0, i_13_134_4559_0, i_13_134_4591_0,
    o_13_134_0_0  );
  input  i_13_134_65_0, i_13_134_94_0, i_13_134_95_0, i_13_134_173_0,
    i_13_134_175_0, i_13_134_176_0, i_13_134_202_0, i_13_134_235_0,
    i_13_134_307_0, i_13_134_308_0, i_13_134_442_0, i_13_134_443_0,
    i_13_134_485_0, i_13_134_572_0, i_13_134_604_0, i_13_134_605_0,
    i_13_134_658_0, i_13_134_662_0, i_13_134_667_0, i_13_134_668_0,
    i_13_134_676_0, i_13_134_677_0, i_13_134_698_0, i_13_134_934_0,
    i_13_134_946_0, i_13_134_1066_0, i_13_134_1217_0, i_13_134_1267_0,
    i_13_134_1306_0, i_13_134_1310_0, i_13_134_1388_0, i_13_134_1499_0,
    i_13_134_1504_0, i_13_134_1505_0, i_13_134_1561_0, i_13_134_1621_0,
    i_13_134_1630_0, i_13_134_1670_0, i_13_134_1720_0, i_13_134_1730_0,
    i_13_134_1802_0, i_13_134_1837_0, i_13_134_1838_0, i_13_134_1840_0,
    i_13_134_1841_0, i_13_134_1904_0, i_13_134_2170_0, i_13_134_2173_0,
    i_13_134_2230_0, i_13_134_2422_0, i_13_134_2423_0, i_13_134_2424_0,
    i_13_134_2425_0, i_13_134_2426_0, i_13_134_2431_0, i_13_134_2432_0,
    i_13_134_2435_0, i_13_134_2503_0, i_13_134_2593_0, i_13_134_2674_0,
    i_13_134_2675_0, i_13_134_2677_0, i_13_134_2678_0, i_13_134_2702_0,
    i_13_134_2912_0, i_13_134_2950_0, i_13_134_2951_0, i_13_134_3142_0,
    i_13_134_3143_0, i_13_134_3145_0, i_13_134_3242_0, i_13_134_3260_0,
    i_13_134_3269_0, i_13_134_3304_0, i_13_134_3305_0, i_13_134_3421_0,
    i_13_134_3422_0, i_13_134_3424_0, i_13_134_3425_0, i_13_134_3446_0,
    i_13_134_3529_0, i_13_134_3592_0, i_13_134_3726_0, i_13_134_3871_0,
    i_13_134_4016_0, i_13_134_4018_0, i_13_134_4019_0, i_13_134_4078_0,
    i_13_134_4079_0, i_13_134_4249_0, i_13_134_4253_0, i_13_134_4258_0,
    i_13_134_4351_0, i_13_134_4430_0, i_13_134_4447_0, i_13_134_4541_0,
    i_13_134_4555_0, i_13_134_4556_0, i_13_134_4559_0, i_13_134_4591_0;
  output o_13_134_0_0;
  assign o_13_134_0_0 = ~((~i_13_134_307_0 & ((~i_13_134_308_0 & ~i_13_134_667_0 & ~i_13_134_1838_0 & ~i_13_134_3260_0) | (~i_13_134_2424_0 & ~i_13_134_2675_0 & ~i_13_134_2678_0 & ~i_13_134_4555_0))) | (~i_13_134_2678_0 & ~i_13_134_4555_0 & ~i_13_134_442_0 & ~i_13_134_2424_0) | (~i_13_134_676_0 & i_13_134_1499_0 & ~i_13_134_2426_0 & ~i_13_134_2431_0) | (~i_13_134_668_0 & ~i_13_134_2425_0 & i_13_134_3421_0 & ~i_13_134_3424_0) | (~i_13_134_95_0 & ~i_13_134_1837_0 & ~i_13_134_3422_0 & ~i_13_134_3871_0));
endmodule



// Benchmark "kernel_13_135" written by ABC on Sun Jul 19 10:47:18 2020

module kernel_13_135 ( 
    i_13_135_90_0, i_13_135_91_0, i_13_135_94_0, i_13_135_117_0,
    i_13_135_118_0, i_13_135_165_0, i_13_135_168_0, i_13_135_180_0,
    i_13_135_181_0, i_13_135_183_0, i_13_135_201_0, i_13_135_306_0,
    i_13_135_561_0, i_13_135_567_0, i_13_135_685_0, i_13_135_694_0,
    i_13_135_697_0, i_13_135_729_0, i_13_135_732_0, i_13_135_822_0,
    i_13_135_855_0, i_13_135_945_0, i_13_135_949_0, i_13_135_1065_0,
    i_13_135_1075_0, i_13_135_1251_0, i_13_135_1263_0, i_13_135_1297_0,
    i_13_135_1341_0, i_13_135_1344_0, i_13_135_1363_0, i_13_135_1404_0,
    i_13_135_1405_0, i_13_135_1440_0, i_13_135_1485_0, i_13_135_1515_0,
    i_13_135_1620_0, i_13_135_1624_0, i_13_135_1629_0, i_13_135_1633_0,
    i_13_135_1828_0, i_13_135_1836_0, i_13_135_1885_0, i_13_135_1888_0,
    i_13_135_1917_0, i_13_135_1921_0, i_13_135_1936_0, i_13_135_2004_0,
    i_13_135_2107_0, i_13_135_2170_0, i_13_135_2172_0, i_13_135_2205_0,
    i_13_135_2208_0, i_13_135_2233_0, i_13_135_2421_0, i_13_135_2424_0,
    i_13_135_2433_0, i_13_135_2452_0, i_13_135_2467_0, i_13_135_2614_0,
    i_13_135_2676_0, i_13_135_2725_0, i_13_135_2910_0, i_13_135_3019_0,
    i_13_135_3034_0, i_13_135_3063_0, i_13_135_3099_0, i_13_135_3106_0,
    i_13_135_3108_0, i_13_135_3126_0, i_13_135_3144_0, i_13_135_3162_0,
    i_13_135_3163_0, i_13_135_3172_0, i_13_135_3207_0, i_13_135_3208_0,
    i_13_135_3213_0, i_13_135_3240_0, i_13_135_3396_0, i_13_135_3414_0,
    i_13_135_3415_0, i_13_135_3486_0, i_13_135_3699_0, i_13_135_3717_0,
    i_13_135_3762_0, i_13_135_3783_0, i_13_135_3834_0, i_13_135_3843_0,
    i_13_135_3870_0, i_13_135_3871_0, i_13_135_4005_0, i_13_135_4006_0,
    i_13_135_4044_0, i_13_135_4117_0, i_13_135_4350_0, i_13_135_4374_0,
    i_13_135_4401_0, i_13_135_4440_0, i_13_135_4452_0, i_13_135_4564_0,
    o_13_135_0_0  );
  input  i_13_135_90_0, i_13_135_91_0, i_13_135_94_0, i_13_135_117_0,
    i_13_135_118_0, i_13_135_165_0, i_13_135_168_0, i_13_135_180_0,
    i_13_135_181_0, i_13_135_183_0, i_13_135_201_0, i_13_135_306_0,
    i_13_135_561_0, i_13_135_567_0, i_13_135_685_0, i_13_135_694_0,
    i_13_135_697_0, i_13_135_729_0, i_13_135_732_0, i_13_135_822_0,
    i_13_135_855_0, i_13_135_945_0, i_13_135_949_0, i_13_135_1065_0,
    i_13_135_1075_0, i_13_135_1251_0, i_13_135_1263_0, i_13_135_1297_0,
    i_13_135_1341_0, i_13_135_1344_0, i_13_135_1363_0, i_13_135_1404_0,
    i_13_135_1405_0, i_13_135_1440_0, i_13_135_1485_0, i_13_135_1515_0,
    i_13_135_1620_0, i_13_135_1624_0, i_13_135_1629_0, i_13_135_1633_0,
    i_13_135_1828_0, i_13_135_1836_0, i_13_135_1885_0, i_13_135_1888_0,
    i_13_135_1917_0, i_13_135_1921_0, i_13_135_1936_0, i_13_135_2004_0,
    i_13_135_2107_0, i_13_135_2170_0, i_13_135_2172_0, i_13_135_2205_0,
    i_13_135_2208_0, i_13_135_2233_0, i_13_135_2421_0, i_13_135_2424_0,
    i_13_135_2433_0, i_13_135_2452_0, i_13_135_2467_0, i_13_135_2614_0,
    i_13_135_2676_0, i_13_135_2725_0, i_13_135_2910_0, i_13_135_3019_0,
    i_13_135_3034_0, i_13_135_3063_0, i_13_135_3099_0, i_13_135_3106_0,
    i_13_135_3108_0, i_13_135_3126_0, i_13_135_3144_0, i_13_135_3162_0,
    i_13_135_3163_0, i_13_135_3172_0, i_13_135_3207_0, i_13_135_3208_0,
    i_13_135_3213_0, i_13_135_3240_0, i_13_135_3396_0, i_13_135_3414_0,
    i_13_135_3415_0, i_13_135_3486_0, i_13_135_3699_0, i_13_135_3717_0,
    i_13_135_3762_0, i_13_135_3783_0, i_13_135_3834_0, i_13_135_3843_0,
    i_13_135_3870_0, i_13_135_3871_0, i_13_135_4005_0, i_13_135_4006_0,
    i_13_135_4044_0, i_13_135_4117_0, i_13_135_4350_0, i_13_135_4374_0,
    i_13_135_4401_0, i_13_135_4440_0, i_13_135_4452_0, i_13_135_4564_0;
  output o_13_135_0_0;
  assign o_13_135_0_0 = ~((~i_13_135_4005_0 & ((~i_13_135_1065_0 & ~i_13_135_3099_0 & ~i_13_135_3108_0) | (~i_13_135_90_0 & ~i_13_135_3240_0 & ~i_13_135_4374_0))) | (~i_13_135_1405_0 & ~i_13_135_1485_0 & ~i_13_135_4044_0));
endmodule



// Benchmark "kernel_13_136" written by ABC on Sun Jul 19 10:47:19 2020

module kernel_13_136 ( 
    i_13_136_49_0, i_13_136_73_0, i_13_136_76_0, i_13_136_157_0,
    i_13_136_228_0, i_13_136_229_0, i_13_136_282_0, i_13_136_283_0,
    i_13_136_515_0, i_13_136_517_0, i_13_136_535_0, i_13_136_657_0,
    i_13_136_659_0, i_13_136_660_0, i_13_136_724_0, i_13_136_821_0,
    i_13_136_850_0, i_13_136_1017_0, i_13_136_1019_0, i_13_136_1053_0,
    i_13_136_1074_0, i_13_136_1075_0, i_13_136_1286_0, i_13_136_1422_0,
    i_13_136_1425_0, i_13_136_1426_0, i_13_136_1570_0, i_13_136_1632_0,
    i_13_136_1633_0, i_13_136_1634_0, i_13_136_1635_0, i_13_136_1773_0,
    i_13_136_1786_0, i_13_136_1795_0, i_13_136_1841_0, i_13_136_2026_0,
    i_13_136_2029_0, i_13_136_2209_0, i_13_136_2236_0, i_13_136_2396_0,
    i_13_136_2426_0, i_13_136_2448_0, i_13_136_2449_0, i_13_136_2451_0,
    i_13_136_2452_0, i_13_136_2453_0, i_13_136_2454_0, i_13_136_2707_0,
    i_13_136_2722_0, i_13_136_3009_0, i_13_136_3010_0, i_13_136_3037_0,
    i_13_136_3269_0, i_13_136_3388_0, i_13_136_3450_0, i_13_136_3459_0,
    i_13_136_3460_0, i_13_136_3467_0, i_13_136_3484_0, i_13_136_3551_0,
    i_13_136_3567_0, i_13_136_3568_0, i_13_136_3573_0, i_13_136_3576_0,
    i_13_136_3577_0, i_13_136_3636_0, i_13_136_3645_0, i_13_136_3646_0,
    i_13_136_3647_0, i_13_136_3648_0, i_13_136_3684_0, i_13_136_3702_0,
    i_13_136_3729_0, i_13_136_3730_0, i_13_136_3838_0, i_13_136_3852_0,
    i_13_136_3862_0, i_13_136_3889_0, i_13_136_3890_0, i_13_136_3893_0,
    i_13_136_3988_0, i_13_136_4015_0, i_13_136_4017_0, i_13_136_4018_0,
    i_13_136_4079_0, i_13_136_4189_0, i_13_136_4251_0, i_13_136_4252_0,
    i_13_136_4253_0, i_13_136_4261_0, i_13_136_4262_0, i_13_136_4305_0,
    i_13_136_4358_0, i_13_136_4361_0, i_13_136_4513_0, i_13_136_4556_0,
    i_13_136_4557_0, i_13_136_4558_0, i_13_136_4559_0, i_13_136_4591_0,
    o_13_136_0_0  );
  input  i_13_136_49_0, i_13_136_73_0, i_13_136_76_0, i_13_136_157_0,
    i_13_136_228_0, i_13_136_229_0, i_13_136_282_0, i_13_136_283_0,
    i_13_136_515_0, i_13_136_517_0, i_13_136_535_0, i_13_136_657_0,
    i_13_136_659_0, i_13_136_660_0, i_13_136_724_0, i_13_136_821_0,
    i_13_136_850_0, i_13_136_1017_0, i_13_136_1019_0, i_13_136_1053_0,
    i_13_136_1074_0, i_13_136_1075_0, i_13_136_1286_0, i_13_136_1422_0,
    i_13_136_1425_0, i_13_136_1426_0, i_13_136_1570_0, i_13_136_1632_0,
    i_13_136_1633_0, i_13_136_1634_0, i_13_136_1635_0, i_13_136_1773_0,
    i_13_136_1786_0, i_13_136_1795_0, i_13_136_1841_0, i_13_136_2026_0,
    i_13_136_2029_0, i_13_136_2209_0, i_13_136_2236_0, i_13_136_2396_0,
    i_13_136_2426_0, i_13_136_2448_0, i_13_136_2449_0, i_13_136_2451_0,
    i_13_136_2452_0, i_13_136_2453_0, i_13_136_2454_0, i_13_136_2707_0,
    i_13_136_2722_0, i_13_136_3009_0, i_13_136_3010_0, i_13_136_3037_0,
    i_13_136_3269_0, i_13_136_3388_0, i_13_136_3450_0, i_13_136_3459_0,
    i_13_136_3460_0, i_13_136_3467_0, i_13_136_3484_0, i_13_136_3551_0,
    i_13_136_3567_0, i_13_136_3568_0, i_13_136_3573_0, i_13_136_3576_0,
    i_13_136_3577_0, i_13_136_3636_0, i_13_136_3645_0, i_13_136_3646_0,
    i_13_136_3647_0, i_13_136_3648_0, i_13_136_3684_0, i_13_136_3702_0,
    i_13_136_3729_0, i_13_136_3730_0, i_13_136_3838_0, i_13_136_3852_0,
    i_13_136_3862_0, i_13_136_3889_0, i_13_136_3890_0, i_13_136_3893_0,
    i_13_136_3988_0, i_13_136_4015_0, i_13_136_4017_0, i_13_136_4018_0,
    i_13_136_4079_0, i_13_136_4189_0, i_13_136_4251_0, i_13_136_4252_0,
    i_13_136_4253_0, i_13_136_4261_0, i_13_136_4262_0, i_13_136_4305_0,
    i_13_136_4358_0, i_13_136_4361_0, i_13_136_4513_0, i_13_136_4556_0,
    i_13_136_4557_0, i_13_136_4558_0, i_13_136_4559_0, i_13_136_4591_0;
  output o_13_136_0_0;
  assign o_13_136_0_0 = ~((~i_13_136_517_0 & ((~i_13_136_1425_0 & ~i_13_136_3647_0) | (~i_13_136_1019_0 & ~i_13_136_2454_0 & ~i_13_136_3459_0 & ~i_13_136_3645_0 & ~i_13_136_3852_0 & ~i_13_136_4358_0))) | (i_13_136_535_0 & ~i_13_136_3460_0) | (~i_13_136_3576_0 & ~i_13_136_3729_0 & ~i_13_136_3852_0 & ~i_13_136_3889_0) | (i_13_136_3388_0 & ~i_13_136_4252_0) | (i_13_136_229_0 & ~i_13_136_1570_0 & ~i_13_136_1773_0 & ~i_13_136_4261_0) | (~i_13_136_2026_0 & ~i_13_136_4361_0 & ~i_13_136_4557_0));
endmodule



// Benchmark "kernel_13_137" written by ABC on Sun Jul 19 10:47:20 2020

module kernel_13_137 ( 
    i_13_137_31_0, i_13_137_48_0, i_13_137_55_0, i_13_137_75_0,
    i_13_137_139_0, i_13_137_205_0, i_13_137_210_0, i_13_137_214_0,
    i_13_137_228_0, i_13_137_229_0, i_13_137_230_0, i_13_137_379_0,
    i_13_137_422_0, i_13_137_514_0, i_13_137_517_0, i_13_137_520_0,
    i_13_137_572_0, i_13_137_625_0, i_13_137_659_0, i_13_137_705_0,
    i_13_137_710_0, i_13_137_813_0, i_13_137_848_0, i_13_137_850_0,
    i_13_137_856_0, i_13_137_865_0, i_13_137_949_0, i_13_137_981_0,
    i_13_137_985_0, i_13_137_1018_0, i_13_137_1200_0, i_13_137_1219_0,
    i_13_137_1300_0, i_13_137_1327_0, i_13_137_1334_0, i_13_137_1438_0,
    i_13_137_1569_0, i_13_137_1570_0, i_13_137_1630_0, i_13_137_1678_0,
    i_13_137_1682_0, i_13_137_1831_0, i_13_137_1840_0, i_13_137_1853_0,
    i_13_137_1861_0, i_13_137_1908_0, i_13_137_1909_0, i_13_137_1923_0,
    i_13_137_2027_0, i_13_137_2107_0, i_13_137_2197_0, i_13_137_2239_0,
    i_13_137_2406_0, i_13_137_2407_0, i_13_137_2452_0, i_13_137_2455_0,
    i_13_137_2698_0, i_13_137_2699_0, i_13_137_2721_0, i_13_137_2722_0,
    i_13_137_2753_0, i_13_137_2794_0, i_13_137_2942_0, i_13_137_3010_0,
    i_13_137_3011_0, i_13_137_3014_0, i_13_137_3027_0, i_13_137_3037_0,
    i_13_137_3109_0, i_13_137_3288_0, i_13_137_3397_0, i_13_137_3403_0,
    i_13_137_3464_0, i_13_137_3488_0, i_13_137_3526_0, i_13_137_3546_0,
    i_13_137_3646_0, i_13_137_3763_0, i_13_137_3764_0, i_13_137_3788_0,
    i_13_137_3864_0, i_13_137_3865_0, i_13_137_3888_0, i_13_137_3907_0,
    i_13_137_3910_0, i_13_137_3914_0, i_13_137_4009_0, i_13_137_4018_0,
    i_13_137_4022_0, i_13_137_4157_0, i_13_137_4249_0, i_13_137_4252_0,
    i_13_137_4255_0, i_13_137_4265_0, i_13_137_4382_0, i_13_137_4432_0,
    i_13_137_4557_0, i_13_137_4561_0, i_13_137_4562_0, i_13_137_4589_0,
    o_13_137_0_0  );
  input  i_13_137_31_0, i_13_137_48_0, i_13_137_55_0, i_13_137_75_0,
    i_13_137_139_0, i_13_137_205_0, i_13_137_210_0, i_13_137_214_0,
    i_13_137_228_0, i_13_137_229_0, i_13_137_230_0, i_13_137_379_0,
    i_13_137_422_0, i_13_137_514_0, i_13_137_517_0, i_13_137_520_0,
    i_13_137_572_0, i_13_137_625_0, i_13_137_659_0, i_13_137_705_0,
    i_13_137_710_0, i_13_137_813_0, i_13_137_848_0, i_13_137_850_0,
    i_13_137_856_0, i_13_137_865_0, i_13_137_949_0, i_13_137_981_0,
    i_13_137_985_0, i_13_137_1018_0, i_13_137_1200_0, i_13_137_1219_0,
    i_13_137_1300_0, i_13_137_1327_0, i_13_137_1334_0, i_13_137_1438_0,
    i_13_137_1569_0, i_13_137_1570_0, i_13_137_1630_0, i_13_137_1678_0,
    i_13_137_1682_0, i_13_137_1831_0, i_13_137_1840_0, i_13_137_1853_0,
    i_13_137_1861_0, i_13_137_1908_0, i_13_137_1909_0, i_13_137_1923_0,
    i_13_137_2027_0, i_13_137_2107_0, i_13_137_2197_0, i_13_137_2239_0,
    i_13_137_2406_0, i_13_137_2407_0, i_13_137_2452_0, i_13_137_2455_0,
    i_13_137_2698_0, i_13_137_2699_0, i_13_137_2721_0, i_13_137_2722_0,
    i_13_137_2753_0, i_13_137_2794_0, i_13_137_2942_0, i_13_137_3010_0,
    i_13_137_3011_0, i_13_137_3014_0, i_13_137_3027_0, i_13_137_3037_0,
    i_13_137_3109_0, i_13_137_3288_0, i_13_137_3397_0, i_13_137_3403_0,
    i_13_137_3464_0, i_13_137_3488_0, i_13_137_3526_0, i_13_137_3546_0,
    i_13_137_3646_0, i_13_137_3763_0, i_13_137_3764_0, i_13_137_3788_0,
    i_13_137_3864_0, i_13_137_3865_0, i_13_137_3888_0, i_13_137_3907_0,
    i_13_137_3910_0, i_13_137_3914_0, i_13_137_4009_0, i_13_137_4018_0,
    i_13_137_4022_0, i_13_137_4157_0, i_13_137_4249_0, i_13_137_4252_0,
    i_13_137_4255_0, i_13_137_4265_0, i_13_137_4382_0, i_13_137_4432_0,
    i_13_137_4557_0, i_13_137_4561_0, i_13_137_4562_0, i_13_137_4589_0;
  output o_13_137_0_0;
  assign o_13_137_0_0 = ~((~i_13_137_48_0 & ((i_13_137_139_0 & ~i_13_137_3010_0 & ~i_13_137_3788_0) | (i_13_137_229_0 & ~i_13_137_3546_0 & i_13_137_4252_0))) | (i_13_137_139_0 & ((~i_13_137_3397_0 & i_13_137_3764_0) | (~i_13_137_1569_0 & ~i_13_137_2455_0 & ~i_13_137_3646_0 & ~i_13_137_3864_0))) | (~i_13_137_2406_0 & ((i_13_137_1300_0 & ~i_13_137_1327_0 & ~i_13_137_3864_0) | (~i_13_137_1018_0 & ~i_13_137_1682_0 & ~i_13_137_3526_0 & ~i_13_137_3763_0 & ~i_13_137_3764_0 & ~i_13_137_4561_0))) | (~i_13_137_3763_0 & ((i_13_137_949_0 & ~i_13_137_3109_0) | (~i_13_137_139_0 & ~i_13_137_2107_0 & i_13_137_3109_0 & ~i_13_137_3526_0 & ~i_13_137_3888_0 & ~i_13_137_4561_0))) | (i_13_137_1840_0 & i_13_137_4432_0 & ~i_13_137_4557_0) | (~i_13_137_520_0 & ~i_13_137_981_0 & ~i_13_137_1570_0 & ~i_13_137_1678_0 & ~i_13_137_4562_0));
endmodule



// Benchmark "kernel_13_138" written by ABC on Sun Jul 19 10:47:21 2020

module kernel_13_138 ( 
    i_13_138_40_0, i_13_138_76_0, i_13_138_121_0, i_13_138_122_0,
    i_13_138_226_0, i_13_138_372_0, i_13_138_442_0, i_13_138_456_0,
    i_13_138_490_0, i_13_138_517_0, i_13_138_531_0, i_13_138_532_0,
    i_13_138_533_0, i_13_138_572_0, i_13_138_715_0, i_13_138_722_0,
    i_13_138_930_0, i_13_138_948_0, i_13_138_951_0, i_13_138_1099_0,
    i_13_138_1100_0, i_13_138_1280_0, i_13_138_1303_0, i_13_138_1327_0,
    i_13_138_1408_0, i_13_138_1426_0, i_13_138_1433_0, i_13_138_1446_0,
    i_13_138_1468_0, i_13_138_1623_0, i_13_138_1666_0, i_13_138_1720_0,
    i_13_138_1723_0, i_13_138_1758_0, i_13_138_1783_0, i_13_138_1785_0,
    i_13_138_1786_0, i_13_138_1787_0, i_13_138_1837_0, i_13_138_1904_0,
    i_13_138_1940_0, i_13_138_2014_0, i_13_138_2103_0, i_13_138_2207_0,
    i_13_138_2209_0, i_13_138_2225_0, i_13_138_2236_0, i_13_138_2238_0,
    i_13_138_2242_0, i_13_138_2243_0, i_13_138_2343_0, i_13_138_2358_0,
    i_13_138_2425_0, i_13_138_2428_0, i_13_138_2533_0, i_13_138_2677_0,
    i_13_138_2695_0, i_13_138_2845_0, i_13_138_3018_0, i_13_138_3037_0,
    i_13_138_3038_0, i_13_138_3163_0, i_13_138_3164_0, i_13_138_3217_0,
    i_13_138_3218_0, i_13_138_3219_0, i_13_138_3259_0, i_13_138_3281_0,
    i_13_138_3286_0, i_13_138_3287_0, i_13_138_3322_0, i_13_138_3422_0,
    i_13_138_3426_0, i_13_138_3649_0, i_13_138_3739_0, i_13_138_3754_0,
    i_13_138_3791_0, i_13_138_3873_0, i_13_138_3874_0, i_13_138_3875_0,
    i_13_138_3876_0, i_13_138_3919_0, i_13_138_3925_0, i_13_138_3984_0,
    i_13_138_3985_0, i_13_138_3998_0, i_13_138_4009_0, i_13_138_4010_0,
    i_13_138_4051_0, i_13_138_4078_0, i_13_138_4079_0, i_13_138_4106_0,
    i_13_138_4162_0, i_13_138_4213_0, i_13_138_4261_0, i_13_138_4519_0,
    i_13_138_4524_0, i_13_138_4531_0, i_13_138_4540_0, i_13_138_4558_0,
    o_13_138_0_0  );
  input  i_13_138_40_0, i_13_138_76_0, i_13_138_121_0, i_13_138_122_0,
    i_13_138_226_0, i_13_138_372_0, i_13_138_442_0, i_13_138_456_0,
    i_13_138_490_0, i_13_138_517_0, i_13_138_531_0, i_13_138_532_0,
    i_13_138_533_0, i_13_138_572_0, i_13_138_715_0, i_13_138_722_0,
    i_13_138_930_0, i_13_138_948_0, i_13_138_951_0, i_13_138_1099_0,
    i_13_138_1100_0, i_13_138_1280_0, i_13_138_1303_0, i_13_138_1327_0,
    i_13_138_1408_0, i_13_138_1426_0, i_13_138_1433_0, i_13_138_1446_0,
    i_13_138_1468_0, i_13_138_1623_0, i_13_138_1666_0, i_13_138_1720_0,
    i_13_138_1723_0, i_13_138_1758_0, i_13_138_1783_0, i_13_138_1785_0,
    i_13_138_1786_0, i_13_138_1787_0, i_13_138_1837_0, i_13_138_1904_0,
    i_13_138_1940_0, i_13_138_2014_0, i_13_138_2103_0, i_13_138_2207_0,
    i_13_138_2209_0, i_13_138_2225_0, i_13_138_2236_0, i_13_138_2238_0,
    i_13_138_2242_0, i_13_138_2243_0, i_13_138_2343_0, i_13_138_2358_0,
    i_13_138_2425_0, i_13_138_2428_0, i_13_138_2533_0, i_13_138_2677_0,
    i_13_138_2695_0, i_13_138_2845_0, i_13_138_3018_0, i_13_138_3037_0,
    i_13_138_3038_0, i_13_138_3163_0, i_13_138_3164_0, i_13_138_3217_0,
    i_13_138_3218_0, i_13_138_3219_0, i_13_138_3259_0, i_13_138_3281_0,
    i_13_138_3286_0, i_13_138_3287_0, i_13_138_3322_0, i_13_138_3422_0,
    i_13_138_3426_0, i_13_138_3649_0, i_13_138_3739_0, i_13_138_3754_0,
    i_13_138_3791_0, i_13_138_3873_0, i_13_138_3874_0, i_13_138_3875_0,
    i_13_138_3876_0, i_13_138_3919_0, i_13_138_3925_0, i_13_138_3984_0,
    i_13_138_3985_0, i_13_138_3998_0, i_13_138_4009_0, i_13_138_4010_0,
    i_13_138_4051_0, i_13_138_4078_0, i_13_138_4079_0, i_13_138_4106_0,
    i_13_138_4162_0, i_13_138_4213_0, i_13_138_4261_0, i_13_138_4519_0,
    i_13_138_4524_0, i_13_138_4531_0, i_13_138_4540_0, i_13_138_4558_0;
  output o_13_138_0_0;
  assign o_13_138_0_0 = ~((~i_13_138_3422_0 & ((i_13_138_2677_0 & ~i_13_138_3925_0) | (~i_13_138_3219_0 & ~i_13_138_4078_0))) | (i_13_138_1426_0 & ~i_13_138_2533_0) | (~i_13_138_2428_0 & i_13_138_3985_0) | (~i_13_138_3874_0 & ~i_13_138_4010_0) | (~i_13_138_3426_0 & ~i_13_138_3876_0 & ~i_13_138_4051_0 & i_13_138_4558_0));
endmodule



// Benchmark "kernel_13_139" written by ABC on Sun Jul 19 10:47:22 2020

module kernel_13_139 ( 
    i_13_139_135_0, i_13_139_136_0, i_13_139_181_0, i_13_139_255_0,
    i_13_139_264_0, i_13_139_418_0, i_13_139_517_0, i_13_139_535_0,
    i_13_139_577_0, i_13_139_624_0, i_13_139_640_0, i_13_139_643_0,
    i_13_139_685_0, i_13_139_689_0, i_13_139_696_0, i_13_139_718_0,
    i_13_139_777_0, i_13_139_778_0, i_13_139_891_0, i_13_139_894_0,
    i_13_139_928_0, i_13_139_975_0, i_13_139_976_0, i_13_139_1079_0,
    i_13_139_1120_0, i_13_139_1152_0, i_13_139_1210_0, i_13_139_1257_0,
    i_13_139_1269_0, i_13_139_1277_0, i_13_139_1359_0, i_13_139_1386_0,
    i_13_139_1387_0, i_13_139_1390_0, i_13_139_1407_0, i_13_139_1412_0,
    i_13_139_1462_0, i_13_139_1465_0, i_13_139_1479_0, i_13_139_1480_0,
    i_13_139_1484_0, i_13_139_1669_0, i_13_139_1677_0, i_13_139_1683_0,
    i_13_139_1687_0, i_13_139_1711_0, i_13_139_1756_0, i_13_139_1792_0,
    i_13_139_1800_0, i_13_139_1858_0, i_13_139_1861_0, i_13_139_1907_0,
    i_13_139_2191_0, i_13_139_2379_0, i_13_139_2404_0, i_13_139_2442_0,
    i_13_139_2503_0, i_13_139_2542_0, i_13_139_2586_0, i_13_139_2646_0,
    i_13_139_2647_0, i_13_139_2687_0, i_13_139_2718_0, i_13_139_2746_0,
    i_13_139_2844_0, i_13_139_2845_0, i_13_139_2872_0, i_13_139_2874_0,
    i_13_139_2875_0, i_13_139_2884_0, i_13_139_3224_0, i_13_139_3343_0,
    i_13_139_3352_0, i_13_139_3384_0, i_13_139_3392_0, i_13_139_3402_0,
    i_13_139_3415_0, i_13_139_3429_0, i_13_139_3558_0, i_13_139_3567_0,
    i_13_139_3735_0, i_13_139_3766_0, i_13_139_3790_0, i_13_139_3791_0,
    i_13_139_3836_0, i_13_139_3933_0, i_13_139_4063_0, i_13_139_4077_0,
    i_13_139_4086_0, i_13_139_4097_0, i_13_139_4185_0, i_13_139_4186_0,
    i_13_139_4216_0, i_13_139_4294_0, i_13_139_4296_0, i_13_139_4306_0,
    i_13_139_4375_0, i_13_139_4433_0, i_13_139_4444_0, i_13_139_4599_0,
    o_13_139_0_0  );
  input  i_13_139_135_0, i_13_139_136_0, i_13_139_181_0, i_13_139_255_0,
    i_13_139_264_0, i_13_139_418_0, i_13_139_517_0, i_13_139_535_0,
    i_13_139_577_0, i_13_139_624_0, i_13_139_640_0, i_13_139_643_0,
    i_13_139_685_0, i_13_139_689_0, i_13_139_696_0, i_13_139_718_0,
    i_13_139_777_0, i_13_139_778_0, i_13_139_891_0, i_13_139_894_0,
    i_13_139_928_0, i_13_139_975_0, i_13_139_976_0, i_13_139_1079_0,
    i_13_139_1120_0, i_13_139_1152_0, i_13_139_1210_0, i_13_139_1257_0,
    i_13_139_1269_0, i_13_139_1277_0, i_13_139_1359_0, i_13_139_1386_0,
    i_13_139_1387_0, i_13_139_1390_0, i_13_139_1407_0, i_13_139_1412_0,
    i_13_139_1462_0, i_13_139_1465_0, i_13_139_1479_0, i_13_139_1480_0,
    i_13_139_1484_0, i_13_139_1669_0, i_13_139_1677_0, i_13_139_1683_0,
    i_13_139_1687_0, i_13_139_1711_0, i_13_139_1756_0, i_13_139_1792_0,
    i_13_139_1800_0, i_13_139_1858_0, i_13_139_1861_0, i_13_139_1907_0,
    i_13_139_2191_0, i_13_139_2379_0, i_13_139_2404_0, i_13_139_2442_0,
    i_13_139_2503_0, i_13_139_2542_0, i_13_139_2586_0, i_13_139_2646_0,
    i_13_139_2647_0, i_13_139_2687_0, i_13_139_2718_0, i_13_139_2746_0,
    i_13_139_2844_0, i_13_139_2845_0, i_13_139_2872_0, i_13_139_2874_0,
    i_13_139_2875_0, i_13_139_2884_0, i_13_139_3224_0, i_13_139_3343_0,
    i_13_139_3352_0, i_13_139_3384_0, i_13_139_3392_0, i_13_139_3402_0,
    i_13_139_3415_0, i_13_139_3429_0, i_13_139_3558_0, i_13_139_3567_0,
    i_13_139_3735_0, i_13_139_3766_0, i_13_139_3790_0, i_13_139_3791_0,
    i_13_139_3836_0, i_13_139_3933_0, i_13_139_4063_0, i_13_139_4077_0,
    i_13_139_4086_0, i_13_139_4097_0, i_13_139_4185_0, i_13_139_4186_0,
    i_13_139_4216_0, i_13_139_4294_0, i_13_139_4296_0, i_13_139_4306_0,
    i_13_139_4375_0, i_13_139_4433_0, i_13_139_4444_0, i_13_139_4599_0;
  output o_13_139_0_0;
  assign o_13_139_0_0 = ~(~i_13_139_4185_0 | (~i_13_139_2844_0 & i_13_139_3766_0) | (~i_13_139_135_0 & ~i_13_139_2874_0) | (~i_13_139_1800_0 & ~i_13_139_2872_0));
endmodule



// Benchmark "kernel_13_140" written by ABC on Sun Jul 19 10:47:23 2020

module kernel_13_140 ( 
    i_13_140_39_0, i_13_140_80_0, i_13_140_105_0, i_13_140_159_0,
    i_13_140_169_0, i_13_140_247_0, i_13_140_268_0, i_13_140_337_0,
    i_13_140_339_0, i_13_140_340_0, i_13_140_373_0, i_13_140_386_0,
    i_13_140_466_0, i_13_140_490_0, i_13_140_607_0, i_13_140_610_0,
    i_13_140_618_0, i_13_140_661_0, i_13_140_780_0, i_13_140_816_0,
    i_13_140_817_0, i_13_140_886_0, i_13_140_931_0, i_13_140_979_0,
    i_13_140_1084_0, i_13_140_1147_0, i_13_140_1150_0, i_13_140_1185_0,
    i_13_140_1210_0, i_13_140_1248_0, i_13_140_1255_0, i_13_140_1265_0,
    i_13_140_1302_0, i_13_140_1303_0, i_13_140_1304_0, i_13_140_1313_0,
    i_13_140_1464_0, i_13_140_1600_0, i_13_140_1725_0, i_13_140_1750_0,
    i_13_140_1763_0, i_13_140_1806_0, i_13_140_1807_0, i_13_140_1815_0,
    i_13_140_1816_0, i_13_140_1934_0, i_13_140_2106_0, i_13_140_2130_0,
    i_13_140_2139_0, i_13_140_2140_0, i_13_140_2141_0, i_13_140_2266_0,
    i_13_140_2267_0, i_13_140_2410_0, i_13_140_2446_0, i_13_140_2463_0,
    i_13_140_2484_0, i_13_140_2657_0, i_13_140_2705_0, i_13_140_2752_0,
    i_13_140_2759_0, i_13_140_2824_0, i_13_140_2859_0, i_13_140_2918_0,
    i_13_140_2941_0, i_13_140_3001_0, i_13_140_3219_0, i_13_140_3220_0,
    i_13_140_3250_0, i_13_140_3272_0, i_13_140_3292_0, i_13_140_3308_0,
    i_13_140_3392_0, i_13_140_3416_0, i_13_140_3476_0, i_13_140_3479_0,
    i_13_140_3482_0, i_13_140_3505_0, i_13_140_3733_0, i_13_140_3874_0,
    i_13_140_3910_0, i_13_140_3913_0, i_13_140_3931_0, i_13_140_3991_0,
    i_13_140_4015_0, i_13_140_4016_0, i_13_140_4066_0, i_13_140_4136_0,
    i_13_140_4162_0, i_13_140_4232_0, i_13_140_4237_0, i_13_140_4273_0,
    i_13_140_4309_0, i_13_140_4310_0, i_13_140_4317_0, i_13_140_4319_0,
    i_13_140_4371_0, i_13_140_4372_0, i_13_140_4381_0, i_13_140_4497_0,
    o_13_140_0_0  );
  input  i_13_140_39_0, i_13_140_80_0, i_13_140_105_0, i_13_140_159_0,
    i_13_140_169_0, i_13_140_247_0, i_13_140_268_0, i_13_140_337_0,
    i_13_140_339_0, i_13_140_340_0, i_13_140_373_0, i_13_140_386_0,
    i_13_140_466_0, i_13_140_490_0, i_13_140_607_0, i_13_140_610_0,
    i_13_140_618_0, i_13_140_661_0, i_13_140_780_0, i_13_140_816_0,
    i_13_140_817_0, i_13_140_886_0, i_13_140_931_0, i_13_140_979_0,
    i_13_140_1084_0, i_13_140_1147_0, i_13_140_1150_0, i_13_140_1185_0,
    i_13_140_1210_0, i_13_140_1248_0, i_13_140_1255_0, i_13_140_1265_0,
    i_13_140_1302_0, i_13_140_1303_0, i_13_140_1304_0, i_13_140_1313_0,
    i_13_140_1464_0, i_13_140_1600_0, i_13_140_1725_0, i_13_140_1750_0,
    i_13_140_1763_0, i_13_140_1806_0, i_13_140_1807_0, i_13_140_1815_0,
    i_13_140_1816_0, i_13_140_1934_0, i_13_140_2106_0, i_13_140_2130_0,
    i_13_140_2139_0, i_13_140_2140_0, i_13_140_2141_0, i_13_140_2266_0,
    i_13_140_2267_0, i_13_140_2410_0, i_13_140_2446_0, i_13_140_2463_0,
    i_13_140_2484_0, i_13_140_2657_0, i_13_140_2705_0, i_13_140_2752_0,
    i_13_140_2759_0, i_13_140_2824_0, i_13_140_2859_0, i_13_140_2918_0,
    i_13_140_2941_0, i_13_140_3001_0, i_13_140_3219_0, i_13_140_3220_0,
    i_13_140_3250_0, i_13_140_3272_0, i_13_140_3292_0, i_13_140_3308_0,
    i_13_140_3392_0, i_13_140_3416_0, i_13_140_3476_0, i_13_140_3479_0,
    i_13_140_3482_0, i_13_140_3505_0, i_13_140_3733_0, i_13_140_3874_0,
    i_13_140_3910_0, i_13_140_3913_0, i_13_140_3931_0, i_13_140_3991_0,
    i_13_140_4015_0, i_13_140_4016_0, i_13_140_4066_0, i_13_140_4136_0,
    i_13_140_4162_0, i_13_140_4232_0, i_13_140_4237_0, i_13_140_4273_0,
    i_13_140_4309_0, i_13_140_4310_0, i_13_140_4317_0, i_13_140_4319_0,
    i_13_140_4371_0, i_13_140_4372_0, i_13_140_4381_0, i_13_140_4497_0;
  output o_13_140_0_0;
  assign o_13_140_0_0 = ~((~i_13_140_2140_0 & ((~i_13_140_340_0 & ~i_13_140_1816_0 & ~i_13_140_2410_0) | (~i_13_140_2139_0 & ~i_13_140_3292_0))) | (i_13_140_1084_0 & i_13_140_1147_0) | (~i_13_140_386_0 & ~i_13_140_3219_0 & i_13_140_3505_0 & i_13_140_4162_0));
endmodule



// Benchmark "kernel_13_141" written by ABC on Sun Jul 19 10:47:24 2020

module kernel_13_141 ( 
    i_13_141_45_0, i_13_141_91_0, i_13_141_95_0, i_13_141_116_0,
    i_13_141_139_0, i_13_141_164_0, i_13_141_165_0, i_13_141_167_0,
    i_13_141_175_0, i_13_141_180_0, i_13_141_185_0, i_13_141_310_0,
    i_13_141_319_0, i_13_141_412_0, i_13_141_455_0, i_13_141_568_0,
    i_13_141_648_0, i_13_141_696_0, i_13_141_697_0, i_13_141_698_0,
    i_13_141_743_0, i_13_141_763_0, i_13_141_813_0, i_13_141_853_0,
    i_13_141_858_0, i_13_141_898_0, i_13_141_961_0, i_13_141_978_0,
    i_13_141_981_0, i_13_141_982_0, i_13_141_984_0, i_13_141_1065_0,
    i_13_141_1067_0, i_13_141_1133_0, i_13_141_1219_0, i_13_141_1360_0,
    i_13_141_1394_0, i_13_141_1405_0, i_13_141_1408_0, i_13_141_1515_0,
    i_13_141_1517_0, i_13_141_1526_0, i_13_141_1664_0, i_13_141_1695_0,
    i_13_141_1777_0, i_13_141_1790_0, i_13_141_1831_0, i_13_141_1832_0,
    i_13_141_1849_0, i_13_141_1852_0, i_13_141_1885_0, i_13_141_2046_0,
    i_13_141_2097_0, i_13_141_2246_0, i_13_141_2265_0, i_13_141_2356_0,
    i_13_141_2404_0, i_13_141_2407_0, i_13_141_2437_0, i_13_141_2469_0,
    i_13_141_2473_0, i_13_141_2532_0, i_13_141_2544_0, i_13_141_2691_0,
    i_13_141_2921_0, i_13_141_2982_0, i_13_141_2983_0, i_13_141_2984_0,
    i_13_141_3000_0, i_13_141_3006_0, i_13_141_3059_0, i_13_141_3108_0,
    i_13_141_3110_0, i_13_141_3145_0, i_13_141_3159_0, i_13_141_3205_0,
    i_13_141_3207_0, i_13_141_3208_0, i_13_141_3209_0, i_13_141_3210_0,
    i_13_141_3211_0, i_13_141_3343_0, i_13_141_3355_0, i_13_141_3406_0,
    i_13_141_3428_0, i_13_141_3511_0, i_13_141_3764_0, i_13_141_3793_0,
    i_13_141_3819_0, i_13_141_3907_0, i_13_141_3911_0, i_13_141_3931_0,
    i_13_141_3995_0, i_13_141_4063_0, i_13_141_4066_0, i_13_141_4182_0,
    i_13_141_4375_0, i_13_141_4519_0, i_13_141_4564_0, i_13_141_4567_0,
    o_13_141_0_0  );
  input  i_13_141_45_0, i_13_141_91_0, i_13_141_95_0, i_13_141_116_0,
    i_13_141_139_0, i_13_141_164_0, i_13_141_165_0, i_13_141_167_0,
    i_13_141_175_0, i_13_141_180_0, i_13_141_185_0, i_13_141_310_0,
    i_13_141_319_0, i_13_141_412_0, i_13_141_455_0, i_13_141_568_0,
    i_13_141_648_0, i_13_141_696_0, i_13_141_697_0, i_13_141_698_0,
    i_13_141_743_0, i_13_141_763_0, i_13_141_813_0, i_13_141_853_0,
    i_13_141_858_0, i_13_141_898_0, i_13_141_961_0, i_13_141_978_0,
    i_13_141_981_0, i_13_141_982_0, i_13_141_984_0, i_13_141_1065_0,
    i_13_141_1067_0, i_13_141_1133_0, i_13_141_1219_0, i_13_141_1360_0,
    i_13_141_1394_0, i_13_141_1405_0, i_13_141_1408_0, i_13_141_1515_0,
    i_13_141_1517_0, i_13_141_1526_0, i_13_141_1664_0, i_13_141_1695_0,
    i_13_141_1777_0, i_13_141_1790_0, i_13_141_1831_0, i_13_141_1832_0,
    i_13_141_1849_0, i_13_141_1852_0, i_13_141_1885_0, i_13_141_2046_0,
    i_13_141_2097_0, i_13_141_2246_0, i_13_141_2265_0, i_13_141_2356_0,
    i_13_141_2404_0, i_13_141_2407_0, i_13_141_2437_0, i_13_141_2469_0,
    i_13_141_2473_0, i_13_141_2532_0, i_13_141_2544_0, i_13_141_2691_0,
    i_13_141_2921_0, i_13_141_2982_0, i_13_141_2983_0, i_13_141_2984_0,
    i_13_141_3000_0, i_13_141_3006_0, i_13_141_3059_0, i_13_141_3108_0,
    i_13_141_3110_0, i_13_141_3145_0, i_13_141_3159_0, i_13_141_3205_0,
    i_13_141_3207_0, i_13_141_3208_0, i_13_141_3209_0, i_13_141_3210_0,
    i_13_141_3211_0, i_13_141_3343_0, i_13_141_3355_0, i_13_141_3406_0,
    i_13_141_3428_0, i_13_141_3511_0, i_13_141_3764_0, i_13_141_3793_0,
    i_13_141_3819_0, i_13_141_3907_0, i_13_141_3911_0, i_13_141_3931_0,
    i_13_141_3995_0, i_13_141_4063_0, i_13_141_4066_0, i_13_141_4182_0,
    i_13_141_4375_0, i_13_141_4519_0, i_13_141_4564_0, i_13_141_4567_0;
  output o_13_141_0_0;
  assign o_13_141_0_0 = ~((i_13_141_1777_0 & ((i_13_141_3108_0 & ~i_13_141_3208_0) | (i_13_141_858_0 & ~i_13_141_2983_0 & ~i_13_141_4063_0 & ~i_13_141_4567_0))) | (~i_13_141_2407_0 & ((i_13_141_696_0 & i_13_141_697_0 & i_13_141_3931_0) | (~i_13_141_982_0 & ~i_13_141_1408_0 & ~i_13_141_2404_0 & ~i_13_141_3995_0 & ~i_13_141_4063_0))) | (~i_13_141_648_0 & ~i_13_141_2984_0 & ~i_13_141_3208_0 & ~i_13_141_3210_0 & ~i_13_141_4063_0) | (~i_13_141_319_0 & ~i_13_141_984_0 & ~i_13_141_1526_0 & ~i_13_141_3995_0 & ~i_13_141_4066_0 & ~i_13_141_4567_0));
endmodule



// Benchmark "kernel_13_142" written by ABC on Sun Jul 19 10:47:24 2020

module kernel_13_142 ( 
    i_13_142_106_0, i_13_142_107_0, i_13_142_112_0, i_13_142_124_0,
    i_13_142_367_0, i_13_142_607_0, i_13_142_624_0, i_13_142_625_0,
    i_13_142_858_0, i_13_142_870_0, i_13_142_948_0, i_13_142_1069_0,
    i_13_142_1070_0, i_13_142_1075_0, i_13_142_1086_0, i_13_142_1087_0,
    i_13_142_1203_0, i_13_142_1348_0, i_13_142_1473_0, i_13_142_1474_0,
    i_13_142_1518_0, i_13_142_1519_0, i_13_142_1571_0, i_13_142_1572_0,
    i_13_142_1573_0, i_13_142_1574_0, i_13_142_1623_0, i_13_142_1632_0,
    i_13_142_1642_0, i_13_142_1780_0, i_13_142_1789_0, i_13_142_1795_0,
    i_13_142_1804_0, i_13_142_1840_0, i_13_142_1843_0, i_13_142_1869_0,
    i_13_142_1993_0, i_13_142_2024_0, i_13_142_2059_0, i_13_142_2060_0,
    i_13_142_2120_0, i_13_142_2137_0, i_13_142_2173_0, i_13_142_2191_0,
    i_13_142_2267_0, i_13_142_2348_0, i_13_142_2380_0, i_13_142_2407_0,
    i_13_142_2417_0, i_13_142_2429_0, i_13_142_2434_0, i_13_142_2437_0,
    i_13_142_2536_0, i_13_142_2563_0, i_13_142_2705_0, i_13_142_2715_0,
    i_13_142_2716_0, i_13_142_2767_0, i_13_142_2986_0, i_13_142_2998_0,
    i_13_142_3103_0, i_13_142_3126_0, i_13_142_3145_0, i_13_142_3147_0,
    i_13_142_3148_0, i_13_142_3166_0, i_13_142_3238_0, i_13_142_3274_0,
    i_13_142_3343_0, i_13_142_3346_0, i_13_142_3373_0, i_13_142_3378_0,
    i_13_142_3392_0, i_13_142_3418_0, i_13_142_3419_0, i_13_142_3423_0,
    i_13_142_3427_0, i_13_142_3454_0, i_13_142_3527_0, i_13_142_3544_0,
    i_13_142_3554_0, i_13_142_3561_0, i_13_142_3767_0, i_13_142_3874_0,
    i_13_142_3937_0, i_13_142_3994_0, i_13_142_4021_0, i_13_142_4045_0,
    i_13_142_4048_0, i_13_142_4093_0, i_13_142_4119_0, i_13_142_4120_0,
    i_13_142_4237_0, i_13_142_4328_0, i_13_142_4342_0, i_13_142_4353_0,
    i_13_142_4399_0, i_13_142_4417_0, i_13_142_4544_0, i_13_142_4561_0,
    o_13_142_0_0  );
  input  i_13_142_106_0, i_13_142_107_0, i_13_142_112_0, i_13_142_124_0,
    i_13_142_367_0, i_13_142_607_0, i_13_142_624_0, i_13_142_625_0,
    i_13_142_858_0, i_13_142_870_0, i_13_142_948_0, i_13_142_1069_0,
    i_13_142_1070_0, i_13_142_1075_0, i_13_142_1086_0, i_13_142_1087_0,
    i_13_142_1203_0, i_13_142_1348_0, i_13_142_1473_0, i_13_142_1474_0,
    i_13_142_1518_0, i_13_142_1519_0, i_13_142_1571_0, i_13_142_1572_0,
    i_13_142_1573_0, i_13_142_1574_0, i_13_142_1623_0, i_13_142_1632_0,
    i_13_142_1642_0, i_13_142_1780_0, i_13_142_1789_0, i_13_142_1795_0,
    i_13_142_1804_0, i_13_142_1840_0, i_13_142_1843_0, i_13_142_1869_0,
    i_13_142_1993_0, i_13_142_2024_0, i_13_142_2059_0, i_13_142_2060_0,
    i_13_142_2120_0, i_13_142_2137_0, i_13_142_2173_0, i_13_142_2191_0,
    i_13_142_2267_0, i_13_142_2348_0, i_13_142_2380_0, i_13_142_2407_0,
    i_13_142_2417_0, i_13_142_2429_0, i_13_142_2434_0, i_13_142_2437_0,
    i_13_142_2536_0, i_13_142_2563_0, i_13_142_2705_0, i_13_142_2715_0,
    i_13_142_2716_0, i_13_142_2767_0, i_13_142_2986_0, i_13_142_2998_0,
    i_13_142_3103_0, i_13_142_3126_0, i_13_142_3145_0, i_13_142_3147_0,
    i_13_142_3148_0, i_13_142_3166_0, i_13_142_3238_0, i_13_142_3274_0,
    i_13_142_3343_0, i_13_142_3346_0, i_13_142_3373_0, i_13_142_3378_0,
    i_13_142_3392_0, i_13_142_3418_0, i_13_142_3419_0, i_13_142_3423_0,
    i_13_142_3427_0, i_13_142_3454_0, i_13_142_3527_0, i_13_142_3544_0,
    i_13_142_3554_0, i_13_142_3561_0, i_13_142_3767_0, i_13_142_3874_0,
    i_13_142_3937_0, i_13_142_3994_0, i_13_142_4021_0, i_13_142_4045_0,
    i_13_142_4048_0, i_13_142_4093_0, i_13_142_4119_0, i_13_142_4120_0,
    i_13_142_4237_0, i_13_142_4328_0, i_13_142_4342_0, i_13_142_4353_0,
    i_13_142_4399_0, i_13_142_4417_0, i_13_142_4544_0, i_13_142_4561_0;
  output o_13_142_0_0;
  assign o_13_142_0_0 = ~(~i_13_142_2173_0 | (~i_13_142_1348_0 & ~i_13_142_2060_0 & ~i_13_142_4353_0) | (~i_13_142_1070_0 & ~i_13_142_1086_0 & ~i_13_142_1572_0 & ~i_13_142_4328_0));
endmodule



// Benchmark "kernel_13_143" written by ABC on Sun Jul 19 10:47:25 2020

module kernel_13_143 ( 
    i_13_143_41_0, i_13_143_52_0, i_13_143_53_0, i_13_143_142_0,
    i_13_143_194_0, i_13_143_196_0, i_13_143_283_0, i_13_143_314_0,
    i_13_143_319_0, i_13_143_320_0, i_13_143_325_0, i_13_143_326_0,
    i_13_143_463_0, i_13_143_464_0, i_13_143_580_0, i_13_143_592_0,
    i_13_143_647_0, i_13_143_661_0, i_13_143_688_0, i_13_143_689_0,
    i_13_143_691_0, i_13_143_692_0, i_13_143_707_0, i_13_143_817_0,
    i_13_143_818_0, i_13_143_826_0, i_13_143_844_0, i_13_143_848_0,
    i_13_143_862_0, i_13_143_1019_0, i_13_143_1124_0, i_13_143_1255_0,
    i_13_143_1316_0, i_13_143_1358_0, i_13_143_1445_0, i_13_143_1471_0,
    i_13_143_1489_0, i_13_143_1492_0, i_13_143_1574_0, i_13_143_1600_0,
    i_13_143_1672_0, i_13_143_1852_0, i_13_143_1876_0, i_13_143_1955_0,
    i_13_143_1997_0, i_13_143_2173_0, i_13_143_2177_0, i_13_143_2185_0,
    i_13_143_2195_0, i_13_143_2264_0, i_13_143_2266_0, i_13_143_2267_0,
    i_13_143_2383_0, i_13_143_2408_0, i_13_143_2410_0, i_13_143_2411_0,
    i_13_143_2591_0, i_13_143_2600_0, i_13_143_2653_0, i_13_143_2654_0,
    i_13_143_2699_0, i_13_143_2860_0, i_13_143_2914_0, i_13_143_2918_0,
    i_13_143_2941_0, i_13_143_3067_0, i_13_143_3068_0, i_13_143_3077_0,
    i_13_143_3145_0, i_13_143_3146_0, i_13_143_3292_0, i_13_143_3373_0,
    i_13_143_3374_0, i_13_143_3392_0, i_13_143_3479_0, i_13_143_3527_0,
    i_13_143_3541_0, i_13_143_3595_0, i_13_143_3722_0, i_13_143_3733_0,
    i_13_143_3770_0, i_13_143_3781_0, i_13_143_3821_0, i_13_143_3982_0,
    i_13_143_3985_0, i_13_143_3995_0, i_13_143_4021_0, i_13_143_4022_0,
    i_13_143_4066_0, i_13_143_4067_0, i_13_143_4171_0, i_13_143_4318_0,
    i_13_143_4319_0, i_13_143_4369_0, i_13_143_4372_0, i_13_143_4448_0,
    i_13_143_4513_0, i_13_143_4540_0, i_13_143_4559_0, i_13_143_4598_0,
    o_13_143_0_0  );
  input  i_13_143_41_0, i_13_143_52_0, i_13_143_53_0, i_13_143_142_0,
    i_13_143_194_0, i_13_143_196_0, i_13_143_283_0, i_13_143_314_0,
    i_13_143_319_0, i_13_143_320_0, i_13_143_325_0, i_13_143_326_0,
    i_13_143_463_0, i_13_143_464_0, i_13_143_580_0, i_13_143_592_0,
    i_13_143_647_0, i_13_143_661_0, i_13_143_688_0, i_13_143_689_0,
    i_13_143_691_0, i_13_143_692_0, i_13_143_707_0, i_13_143_817_0,
    i_13_143_818_0, i_13_143_826_0, i_13_143_844_0, i_13_143_848_0,
    i_13_143_862_0, i_13_143_1019_0, i_13_143_1124_0, i_13_143_1255_0,
    i_13_143_1316_0, i_13_143_1358_0, i_13_143_1445_0, i_13_143_1471_0,
    i_13_143_1489_0, i_13_143_1492_0, i_13_143_1574_0, i_13_143_1600_0,
    i_13_143_1672_0, i_13_143_1852_0, i_13_143_1876_0, i_13_143_1955_0,
    i_13_143_1997_0, i_13_143_2173_0, i_13_143_2177_0, i_13_143_2185_0,
    i_13_143_2195_0, i_13_143_2264_0, i_13_143_2266_0, i_13_143_2267_0,
    i_13_143_2383_0, i_13_143_2408_0, i_13_143_2410_0, i_13_143_2411_0,
    i_13_143_2591_0, i_13_143_2600_0, i_13_143_2653_0, i_13_143_2654_0,
    i_13_143_2699_0, i_13_143_2860_0, i_13_143_2914_0, i_13_143_2918_0,
    i_13_143_2941_0, i_13_143_3067_0, i_13_143_3068_0, i_13_143_3077_0,
    i_13_143_3145_0, i_13_143_3146_0, i_13_143_3292_0, i_13_143_3373_0,
    i_13_143_3374_0, i_13_143_3392_0, i_13_143_3479_0, i_13_143_3527_0,
    i_13_143_3541_0, i_13_143_3595_0, i_13_143_3722_0, i_13_143_3733_0,
    i_13_143_3770_0, i_13_143_3781_0, i_13_143_3821_0, i_13_143_3982_0,
    i_13_143_3985_0, i_13_143_3995_0, i_13_143_4021_0, i_13_143_4022_0,
    i_13_143_4066_0, i_13_143_4067_0, i_13_143_4171_0, i_13_143_4318_0,
    i_13_143_4319_0, i_13_143_4369_0, i_13_143_4372_0, i_13_143_4448_0,
    i_13_143_4513_0, i_13_143_4540_0, i_13_143_4559_0, i_13_143_4598_0;
  output o_13_143_0_0;
  assign o_13_143_0_0 = ~((~i_13_143_2410_0 & ~i_13_143_3068_0) | (~i_13_143_692_0 & ~i_13_143_2411_0));
endmodule



// Benchmark "kernel_13_144" written by ABC on Sun Jul 19 10:47:26 2020

module kernel_13_144 ( 
    i_13_144_20_0, i_13_144_77_0, i_13_144_78_0, i_13_144_107_0,
    i_13_144_113_0, i_13_144_174_0, i_13_144_195_0, i_13_144_368_0,
    i_13_144_386_0, i_13_144_454_0, i_13_144_460_0, i_13_144_502_0,
    i_13_144_528_0, i_13_144_725_0, i_13_144_814_0, i_13_144_859_0,
    i_13_144_949_0, i_13_144_1087_0, i_13_144_1088_0, i_13_144_1148_0,
    i_13_144_1211_0, i_13_144_1219_0, i_13_144_1348_0, i_13_144_1394_0,
    i_13_144_1399_0, i_13_144_1410_0, i_13_144_1426_0, i_13_144_1474_0,
    i_13_144_1509_0, i_13_144_1570_0, i_13_144_1573_0, i_13_144_1622_0,
    i_13_144_1624_0, i_13_144_1633_0, i_13_144_1741_0, i_13_144_1789_0,
    i_13_144_1804_0, i_13_144_1840_0, i_13_144_1841_0, i_13_144_1844_0,
    i_13_144_1942_0, i_13_144_2001_0, i_13_144_2024_0, i_13_144_2059_0,
    i_13_144_2123_0, i_13_144_2128_0, i_13_144_2137_0, i_13_144_2230_0,
    i_13_144_2283_0, i_13_144_2284_0, i_13_144_2317_0, i_13_144_2348_0,
    i_13_144_2383_0, i_13_144_2399_0, i_13_144_2435_0, i_13_144_2437_0,
    i_13_144_2438_0, i_13_144_2501_0, i_13_144_2716_0, i_13_144_2717_0,
    i_13_144_2749_0, i_13_144_2856_0, i_13_144_3023_0, i_13_144_3066_0,
    i_13_144_3067_0, i_13_144_3127_0, i_13_144_3137_0, i_13_144_3144_0,
    i_13_144_3147_0, i_13_144_3148_0, i_13_144_3149_0, i_13_144_3166_0,
    i_13_144_3167_0, i_13_144_3329_0, i_13_144_3343_0, i_13_144_3374_0,
    i_13_144_3392_0, i_13_144_3413_0, i_13_144_3428_0, i_13_144_3432_0,
    i_13_144_3455_0, i_13_144_3553_0, i_13_144_3599_0, i_13_144_3923_0,
    i_13_144_4111_0, i_13_144_4120_0, i_13_144_4121_0, i_13_144_4192_0,
    i_13_144_4256_0, i_13_144_4263_0, i_13_144_4264_0, i_13_144_4328_0,
    i_13_144_4333_0, i_13_144_4400_0, i_13_144_4417_0, i_13_144_4418_0,
    i_13_144_4469_0, i_13_144_4526_0, i_13_144_4544_0, i_13_144_4596_0,
    o_13_144_0_0  );
  input  i_13_144_20_0, i_13_144_77_0, i_13_144_78_0, i_13_144_107_0,
    i_13_144_113_0, i_13_144_174_0, i_13_144_195_0, i_13_144_368_0,
    i_13_144_386_0, i_13_144_454_0, i_13_144_460_0, i_13_144_502_0,
    i_13_144_528_0, i_13_144_725_0, i_13_144_814_0, i_13_144_859_0,
    i_13_144_949_0, i_13_144_1087_0, i_13_144_1088_0, i_13_144_1148_0,
    i_13_144_1211_0, i_13_144_1219_0, i_13_144_1348_0, i_13_144_1394_0,
    i_13_144_1399_0, i_13_144_1410_0, i_13_144_1426_0, i_13_144_1474_0,
    i_13_144_1509_0, i_13_144_1570_0, i_13_144_1573_0, i_13_144_1622_0,
    i_13_144_1624_0, i_13_144_1633_0, i_13_144_1741_0, i_13_144_1789_0,
    i_13_144_1804_0, i_13_144_1840_0, i_13_144_1841_0, i_13_144_1844_0,
    i_13_144_1942_0, i_13_144_2001_0, i_13_144_2024_0, i_13_144_2059_0,
    i_13_144_2123_0, i_13_144_2128_0, i_13_144_2137_0, i_13_144_2230_0,
    i_13_144_2283_0, i_13_144_2284_0, i_13_144_2317_0, i_13_144_2348_0,
    i_13_144_2383_0, i_13_144_2399_0, i_13_144_2435_0, i_13_144_2437_0,
    i_13_144_2438_0, i_13_144_2501_0, i_13_144_2716_0, i_13_144_2717_0,
    i_13_144_2749_0, i_13_144_2856_0, i_13_144_3023_0, i_13_144_3066_0,
    i_13_144_3067_0, i_13_144_3127_0, i_13_144_3137_0, i_13_144_3144_0,
    i_13_144_3147_0, i_13_144_3148_0, i_13_144_3149_0, i_13_144_3166_0,
    i_13_144_3167_0, i_13_144_3329_0, i_13_144_3343_0, i_13_144_3374_0,
    i_13_144_3392_0, i_13_144_3413_0, i_13_144_3428_0, i_13_144_3432_0,
    i_13_144_3455_0, i_13_144_3553_0, i_13_144_3599_0, i_13_144_3923_0,
    i_13_144_4111_0, i_13_144_4120_0, i_13_144_4121_0, i_13_144_4192_0,
    i_13_144_4256_0, i_13_144_4263_0, i_13_144_4264_0, i_13_144_4328_0,
    i_13_144_4333_0, i_13_144_4400_0, i_13_144_4417_0, i_13_144_4418_0,
    i_13_144_4469_0, i_13_144_4526_0, i_13_144_4544_0, i_13_144_4596_0;
  output o_13_144_0_0;
  assign o_13_144_0_0 = ~((~i_13_144_3148_0 & ~i_13_144_3149_0) | (~i_13_144_1509_0 & ~i_13_144_1624_0 & ~i_13_144_2435_0));
endmodule



// Benchmark "kernel_13_145" written by ABC on Sun Jul 19 10:47:27 2020

module kernel_13_145 ( 
    i_13_145_106_0, i_13_145_187_0, i_13_145_284_0, i_13_145_337_0,
    i_13_145_339_0, i_13_145_427_0, i_13_145_454_0, i_13_145_513_0,
    i_13_145_526_0, i_13_145_553_0, i_13_145_589_0, i_13_145_607_0,
    i_13_145_646_0, i_13_145_651_0, i_13_145_673_0, i_13_145_679_0,
    i_13_145_688_0, i_13_145_691_0, i_13_145_694_0, i_13_145_699_0,
    i_13_145_733_0, i_13_145_823_0, i_13_145_840_0, i_13_145_898_0,
    i_13_145_925_0, i_13_145_1033_0, i_13_145_1101_0, i_13_145_1123_0,
    i_13_145_1144_0, i_13_145_1148_0, i_13_145_1179_0, i_13_145_1180_0,
    i_13_145_1226_0, i_13_145_1270_0, i_13_145_1272_0, i_13_145_1273_0,
    i_13_145_1318_0, i_13_145_1345_0, i_13_145_1384_0, i_13_145_1449_0,
    i_13_145_1519_0, i_13_145_1570_0, i_13_145_1633_0, i_13_145_1656_0,
    i_13_145_1657_0, i_13_145_1750_0, i_13_145_1840_0, i_13_145_1858_0,
    i_13_145_1915_0, i_13_145_1930_0, i_13_145_1933_0, i_13_145_1935_0,
    i_13_145_2002_0, i_13_145_2029_0, i_13_145_2088_0, i_13_145_2200_0,
    i_13_145_2209_0, i_13_145_2461_0, i_13_145_2494_0, i_13_145_2496_0,
    i_13_145_2542_0, i_13_145_2600_0, i_13_145_2653_0, i_13_145_2736_0,
    i_13_145_2767_0, i_13_145_2770_0, i_13_145_2845_0, i_13_145_2848_0,
    i_13_145_2886_0, i_13_145_3055_0, i_13_145_3145_0, i_13_145_3151_0,
    i_13_145_3258_0, i_13_145_3316_0, i_13_145_3370_0, i_13_145_3378_0,
    i_13_145_3382_0, i_13_145_3418_0, i_13_145_3431_0, i_13_145_3505_0,
    i_13_145_3535_0, i_13_145_3561_0, i_13_145_3730_0, i_13_145_3736_0,
    i_13_145_3739_0, i_13_145_3756_0, i_13_145_3846_0, i_13_145_3892_0,
    i_13_145_3927_0, i_13_145_4021_0, i_13_145_4036_0, i_13_145_4081_0,
    i_13_145_4158_0, i_13_145_4188_0, i_13_145_4189_0, i_13_145_4315_0,
    i_13_145_4417_0, i_13_145_4578_0, i_13_145_4594_0, i_13_145_4602_0,
    o_13_145_0_0  );
  input  i_13_145_106_0, i_13_145_187_0, i_13_145_284_0, i_13_145_337_0,
    i_13_145_339_0, i_13_145_427_0, i_13_145_454_0, i_13_145_513_0,
    i_13_145_526_0, i_13_145_553_0, i_13_145_589_0, i_13_145_607_0,
    i_13_145_646_0, i_13_145_651_0, i_13_145_673_0, i_13_145_679_0,
    i_13_145_688_0, i_13_145_691_0, i_13_145_694_0, i_13_145_699_0,
    i_13_145_733_0, i_13_145_823_0, i_13_145_840_0, i_13_145_898_0,
    i_13_145_925_0, i_13_145_1033_0, i_13_145_1101_0, i_13_145_1123_0,
    i_13_145_1144_0, i_13_145_1148_0, i_13_145_1179_0, i_13_145_1180_0,
    i_13_145_1226_0, i_13_145_1270_0, i_13_145_1272_0, i_13_145_1273_0,
    i_13_145_1318_0, i_13_145_1345_0, i_13_145_1384_0, i_13_145_1449_0,
    i_13_145_1519_0, i_13_145_1570_0, i_13_145_1633_0, i_13_145_1656_0,
    i_13_145_1657_0, i_13_145_1750_0, i_13_145_1840_0, i_13_145_1858_0,
    i_13_145_1915_0, i_13_145_1930_0, i_13_145_1933_0, i_13_145_1935_0,
    i_13_145_2002_0, i_13_145_2029_0, i_13_145_2088_0, i_13_145_2200_0,
    i_13_145_2209_0, i_13_145_2461_0, i_13_145_2494_0, i_13_145_2496_0,
    i_13_145_2542_0, i_13_145_2600_0, i_13_145_2653_0, i_13_145_2736_0,
    i_13_145_2767_0, i_13_145_2770_0, i_13_145_2845_0, i_13_145_2848_0,
    i_13_145_2886_0, i_13_145_3055_0, i_13_145_3145_0, i_13_145_3151_0,
    i_13_145_3258_0, i_13_145_3316_0, i_13_145_3370_0, i_13_145_3378_0,
    i_13_145_3382_0, i_13_145_3418_0, i_13_145_3431_0, i_13_145_3505_0,
    i_13_145_3535_0, i_13_145_3561_0, i_13_145_3730_0, i_13_145_3736_0,
    i_13_145_3739_0, i_13_145_3756_0, i_13_145_3846_0, i_13_145_3892_0,
    i_13_145_3927_0, i_13_145_4021_0, i_13_145_4036_0, i_13_145_4081_0,
    i_13_145_4158_0, i_13_145_4188_0, i_13_145_4189_0, i_13_145_4315_0,
    i_13_145_4417_0, i_13_145_4578_0, i_13_145_4594_0, i_13_145_4602_0;
  output o_13_145_0_0;
  assign o_13_145_0_0 = ~((~i_13_145_823_0 & ((~i_13_145_284_0 & ~i_13_145_1840_0 & i_13_145_3739_0) | (i_13_145_337_0 & ~i_13_145_4188_0))) | (~i_13_145_898_0 & ~i_13_145_1144_0 & ((i_13_145_589_0 & ~i_13_145_673_0 & ~i_13_145_3892_0 & ~i_13_145_3927_0) | (~i_13_145_4081_0 & ~i_13_145_4189_0))) | (~i_13_145_2848_0 & ((~i_13_145_2653_0 & ((i_13_145_688_0 & ~i_13_145_3258_0) | (i_13_145_2209_0 & ~i_13_145_2736_0 & ~i_13_145_4417_0))) | (i_13_145_1345_0 & i_13_145_2767_0))) | (i_13_145_526_0 & ~i_13_145_1123_0 & ~i_13_145_1656_0));
endmodule



// Benchmark "kernel_13_146" written by ABC on Sun Jul 19 10:47:27 2020

module kernel_13_146 ( 
    i_13_146_28_0, i_13_146_32_0, i_13_146_46_0, i_13_146_49_0,
    i_13_146_65_0, i_13_146_91_0, i_13_146_92_0, i_13_146_118_0,
    i_13_146_122_0, i_13_146_157_0, i_13_146_163_0, i_13_146_317_0,
    i_13_146_320_0, i_13_146_454_0, i_13_146_562_0, i_13_146_568_0,
    i_13_146_671_0, i_13_146_676_0, i_13_146_697_0, i_13_146_722_0,
    i_13_146_730_0, i_13_146_758_0, i_13_146_946_0, i_13_146_1075_0,
    i_13_146_1076_0, i_13_146_1381_0, i_13_146_1405_0, i_13_146_1442_0,
    i_13_146_1454_0, i_13_146_1526_0, i_13_146_1606_0, i_13_146_1621_0,
    i_13_146_1630_0, i_13_146_1633_0, i_13_146_1837_0, i_13_146_1846_0,
    i_13_146_1955_0, i_13_146_1999_0, i_13_146_2000_0, i_13_146_2173_0,
    i_13_146_2174_0, i_13_146_2206_0, i_13_146_2207_0, i_13_146_2422_0,
    i_13_146_2431_0, i_13_146_2432_0, i_13_146_2452_0, i_13_146_2548_0,
    i_13_146_2559_0, i_13_146_2719_0, i_13_146_2750_0, i_13_146_2793_0,
    i_13_146_2846_0, i_13_146_2884_0, i_13_146_3019_0, i_13_146_3034_0,
    i_13_146_3035_0, i_13_146_3126_0, i_13_146_3127_0, i_13_146_3161_0,
    i_13_146_3164_0, i_13_146_3214_0, i_13_146_3242_0, i_13_146_3272_0,
    i_13_146_3415_0, i_13_146_3421_0, i_13_146_3422_0, i_13_146_3434_0,
    i_13_146_3449_0, i_13_146_3477_0, i_13_146_3528_0, i_13_146_3530_0,
    i_13_146_3637_0, i_13_146_3638_0, i_13_146_3646_0, i_13_146_3647_0,
    i_13_146_3699_0, i_13_146_3700_0, i_13_146_3718_0, i_13_146_3837_0,
    i_13_146_3843_0, i_13_146_3844_0, i_13_146_3857_0, i_13_146_3871_0,
    i_13_146_3872_0, i_13_146_3889_0, i_13_146_3901_0, i_13_146_4006_0,
    i_13_146_4007_0, i_13_146_4042_0, i_13_146_4043_0, i_13_146_4105_0,
    i_13_146_4177_0, i_13_146_4304_0, i_13_146_4312_0, i_13_146_4348_0,
    i_13_146_4349_0, i_13_146_4351_0, i_13_146_4387_0, i_13_146_4510_0,
    o_13_146_0_0  );
  input  i_13_146_28_0, i_13_146_32_0, i_13_146_46_0, i_13_146_49_0,
    i_13_146_65_0, i_13_146_91_0, i_13_146_92_0, i_13_146_118_0,
    i_13_146_122_0, i_13_146_157_0, i_13_146_163_0, i_13_146_317_0,
    i_13_146_320_0, i_13_146_454_0, i_13_146_562_0, i_13_146_568_0,
    i_13_146_671_0, i_13_146_676_0, i_13_146_697_0, i_13_146_722_0,
    i_13_146_730_0, i_13_146_758_0, i_13_146_946_0, i_13_146_1075_0,
    i_13_146_1076_0, i_13_146_1381_0, i_13_146_1405_0, i_13_146_1442_0,
    i_13_146_1454_0, i_13_146_1526_0, i_13_146_1606_0, i_13_146_1621_0,
    i_13_146_1630_0, i_13_146_1633_0, i_13_146_1837_0, i_13_146_1846_0,
    i_13_146_1955_0, i_13_146_1999_0, i_13_146_2000_0, i_13_146_2173_0,
    i_13_146_2174_0, i_13_146_2206_0, i_13_146_2207_0, i_13_146_2422_0,
    i_13_146_2431_0, i_13_146_2432_0, i_13_146_2452_0, i_13_146_2548_0,
    i_13_146_2559_0, i_13_146_2719_0, i_13_146_2750_0, i_13_146_2793_0,
    i_13_146_2846_0, i_13_146_2884_0, i_13_146_3019_0, i_13_146_3034_0,
    i_13_146_3035_0, i_13_146_3126_0, i_13_146_3127_0, i_13_146_3161_0,
    i_13_146_3164_0, i_13_146_3214_0, i_13_146_3242_0, i_13_146_3272_0,
    i_13_146_3415_0, i_13_146_3421_0, i_13_146_3422_0, i_13_146_3434_0,
    i_13_146_3449_0, i_13_146_3477_0, i_13_146_3528_0, i_13_146_3530_0,
    i_13_146_3637_0, i_13_146_3638_0, i_13_146_3646_0, i_13_146_3647_0,
    i_13_146_3699_0, i_13_146_3700_0, i_13_146_3718_0, i_13_146_3837_0,
    i_13_146_3843_0, i_13_146_3844_0, i_13_146_3857_0, i_13_146_3871_0,
    i_13_146_3872_0, i_13_146_3889_0, i_13_146_3901_0, i_13_146_4006_0,
    i_13_146_4007_0, i_13_146_4042_0, i_13_146_4043_0, i_13_146_4105_0,
    i_13_146_4177_0, i_13_146_4304_0, i_13_146_4312_0, i_13_146_4348_0,
    i_13_146_4349_0, i_13_146_4351_0, i_13_146_4387_0, i_13_146_4510_0;
  output o_13_146_0_0;
  assign o_13_146_0_0 = ~((~i_13_146_32_0 & ((~i_13_146_1846_0 & ~i_13_146_2422_0) | (i_13_146_1606_0 & ~i_13_146_3857_0))) | (~i_13_146_4348_0 & (i_13_146_697_0 | (~i_13_146_3034_0 & ~i_13_146_3214_0 & ~i_13_146_4304_0))) | (~i_13_146_46_0 & ~i_13_146_4006_0 & ~i_13_146_4312_0));
endmodule



// Benchmark "kernel_13_147" written by ABC on Sun Jul 19 10:47:28 2020

module kernel_13_147 ( 
    i_13_147_26_0, i_13_147_34_0, i_13_147_76_0, i_13_147_79_0,
    i_13_147_102_0, i_13_147_115_0, i_13_147_127_0, i_13_147_128_0,
    i_13_147_140_0, i_13_147_142_0, i_13_147_230_0, i_13_147_232_0,
    i_13_147_233_0, i_13_147_268_0, i_13_147_362_0, i_13_147_538_0,
    i_13_147_539_0, i_13_147_573_0, i_13_147_620_0, i_13_147_690_0,
    i_13_147_691_0, i_13_147_696_0, i_13_147_697_0, i_13_147_699_0,
    i_13_147_700_0, i_13_147_768_0, i_13_147_814_0, i_13_147_826_0,
    i_13_147_827_0, i_13_147_857_0, i_13_147_885_0, i_13_147_1066_0,
    i_13_147_1123_0, i_13_147_1219_0, i_13_147_1220_0, i_13_147_1222_0,
    i_13_147_1275_0, i_13_147_1391_0, i_13_147_1440_0, i_13_147_1629_0,
    i_13_147_1714_0, i_13_147_1718_0, i_13_147_1726_0, i_13_147_1777_0,
    i_13_147_1795_0, i_13_147_1804_0, i_13_147_1807_0, i_13_147_1843_0,
    i_13_147_1888_0, i_13_147_2006_0, i_13_147_2101_0, i_13_147_2119_0,
    i_13_147_2317_0, i_13_147_2342_0, i_13_147_2410_0, i_13_147_2434_0,
    i_13_147_2469_0, i_13_147_2472_0, i_13_147_2654_0, i_13_147_2657_0,
    i_13_147_2713_0, i_13_147_2722_0, i_13_147_2726_0, i_13_147_2851_0,
    i_13_147_3028_0, i_13_147_3038_0, i_13_147_3067_0, i_13_147_3100_0,
    i_13_147_3145_0, i_13_147_3146_0, i_13_147_3148_0, i_13_147_3208_0,
    i_13_147_3211_0, i_13_147_3313_0, i_13_147_3419_0, i_13_147_3443_0,
    i_13_147_3490_0, i_13_147_3501_0, i_13_147_3505_0, i_13_147_3506_0,
    i_13_147_3557_0, i_13_147_3571_0, i_13_147_3572_0, i_13_147_3685_0,
    i_13_147_3741_0, i_13_147_3742_0, i_13_147_3743_0, i_13_147_4063_0,
    i_13_147_4084_0, i_13_147_4092_0, i_13_147_4208_0, i_13_147_4256_0,
    i_13_147_4269_0, i_13_147_4297_0, i_13_147_4298_0, i_13_147_4316_0,
    i_13_147_4367_0, i_13_147_4399_0, i_13_147_4513_0, i_13_147_4538_0,
    o_13_147_0_0  );
  input  i_13_147_26_0, i_13_147_34_0, i_13_147_76_0, i_13_147_79_0,
    i_13_147_102_0, i_13_147_115_0, i_13_147_127_0, i_13_147_128_0,
    i_13_147_140_0, i_13_147_142_0, i_13_147_230_0, i_13_147_232_0,
    i_13_147_233_0, i_13_147_268_0, i_13_147_362_0, i_13_147_538_0,
    i_13_147_539_0, i_13_147_573_0, i_13_147_620_0, i_13_147_690_0,
    i_13_147_691_0, i_13_147_696_0, i_13_147_697_0, i_13_147_699_0,
    i_13_147_700_0, i_13_147_768_0, i_13_147_814_0, i_13_147_826_0,
    i_13_147_827_0, i_13_147_857_0, i_13_147_885_0, i_13_147_1066_0,
    i_13_147_1123_0, i_13_147_1219_0, i_13_147_1220_0, i_13_147_1222_0,
    i_13_147_1275_0, i_13_147_1391_0, i_13_147_1440_0, i_13_147_1629_0,
    i_13_147_1714_0, i_13_147_1718_0, i_13_147_1726_0, i_13_147_1777_0,
    i_13_147_1795_0, i_13_147_1804_0, i_13_147_1807_0, i_13_147_1843_0,
    i_13_147_1888_0, i_13_147_2006_0, i_13_147_2101_0, i_13_147_2119_0,
    i_13_147_2317_0, i_13_147_2342_0, i_13_147_2410_0, i_13_147_2434_0,
    i_13_147_2469_0, i_13_147_2472_0, i_13_147_2654_0, i_13_147_2657_0,
    i_13_147_2713_0, i_13_147_2722_0, i_13_147_2726_0, i_13_147_2851_0,
    i_13_147_3028_0, i_13_147_3038_0, i_13_147_3067_0, i_13_147_3100_0,
    i_13_147_3145_0, i_13_147_3146_0, i_13_147_3148_0, i_13_147_3208_0,
    i_13_147_3211_0, i_13_147_3313_0, i_13_147_3419_0, i_13_147_3443_0,
    i_13_147_3490_0, i_13_147_3501_0, i_13_147_3505_0, i_13_147_3506_0,
    i_13_147_3557_0, i_13_147_3571_0, i_13_147_3572_0, i_13_147_3685_0,
    i_13_147_3741_0, i_13_147_3742_0, i_13_147_3743_0, i_13_147_4063_0,
    i_13_147_4084_0, i_13_147_4092_0, i_13_147_4208_0, i_13_147_4256_0,
    i_13_147_4269_0, i_13_147_4297_0, i_13_147_4298_0, i_13_147_4316_0,
    i_13_147_4367_0, i_13_147_4399_0, i_13_147_4513_0, i_13_147_4538_0;
  output o_13_147_0_0;
  assign o_13_147_0_0 = ~((~i_13_147_115_0 & (~i_13_147_1888_0 | ~i_13_147_2851_0)) | (~i_13_147_4399_0 & ((~i_13_147_697_0 & ((~i_13_147_539_0 & i_13_147_3208_0) | (~i_13_147_233_0 & ~i_13_147_2713_0 & i_13_147_3211_0))) | (~i_13_147_3506_0 & ~i_13_147_4092_0 & ~i_13_147_4269_0))) | (~i_13_147_539_0 & ((i_13_147_233_0 & ~i_13_147_691_0) | (~i_13_147_2713_0 & i_13_147_3146_0 & ~i_13_147_4256_0))) | (~i_13_147_700_0 & ~i_13_147_3742_0));
endmodule



// Benchmark "kernel_13_148" written by ABC on Sun Jul 19 10:47:29 2020

module kernel_13_148 ( 
    i_13_148_61_0, i_13_148_71_0, i_13_148_179_0, i_13_148_274_0,
    i_13_148_275_0, i_13_148_280_0, i_13_148_286_0, i_13_148_493_0,
    i_13_148_529_0, i_13_148_530_0, i_13_148_553_0, i_13_148_562_0,
    i_13_148_599_0, i_13_148_673_0, i_13_148_797_0, i_13_148_841_0,
    i_13_148_853_0, i_13_148_854_0, i_13_148_965_0, i_13_148_1025_0,
    i_13_148_1075_0, i_13_148_1147_0, i_13_148_1282_0, i_13_148_1303_0,
    i_13_148_1304_0, i_13_148_1321_0, i_13_148_1327_0, i_13_148_1490_0,
    i_13_148_1502_0, i_13_148_1516_0, i_13_148_1552_0, i_13_148_1553_0,
    i_13_148_1660_0, i_13_148_1700_0, i_13_148_1817_0, i_13_148_1858_0,
    i_13_148_2002_0, i_13_148_2003_0, i_13_148_2020_0, i_13_148_2021_0,
    i_13_148_2050_0, i_13_148_2201_0, i_13_148_2240_0, i_13_148_2263_0,
    i_13_148_2275_0, i_13_148_2366_0, i_13_148_2461_0, i_13_148_2462_0,
    i_13_148_2470_0, i_13_148_2471_0, i_13_148_2509_0, i_13_148_2543_0,
    i_13_148_2551_0, i_13_148_2615_0, i_13_148_2653_0, i_13_148_2824_0,
    i_13_148_2825_0, i_13_148_2860_0, i_13_148_2920_0, i_13_148_2984_0,
    i_13_148_3173_0, i_13_148_3274_0, i_13_148_3347_0, i_13_148_3418_0,
    i_13_148_3424_0, i_13_148_3428_0, i_13_148_3482_0, i_13_148_3533_0,
    i_13_148_3541_0, i_13_148_3542_0, i_13_148_3544_0, i_13_148_3545_0,
    i_13_148_3580_0, i_13_148_3614_0, i_13_148_3622_0, i_13_148_3634_0,
    i_13_148_3730_0, i_13_148_3731_0, i_13_148_3743_0, i_13_148_3787_0,
    i_13_148_3788_0, i_13_148_3910_0, i_13_148_3911_0, i_13_148_3913_0,
    i_13_148_3914_0, i_13_148_4118_0, i_13_148_4126_0, i_13_148_4162_0,
    i_13_148_4189_0, i_13_148_4237_0, i_13_148_4238_0, i_13_148_4256_0,
    i_13_148_4282_0, i_13_148_4378_0, i_13_148_4381_0, i_13_148_4382_0,
    i_13_148_4400_0, i_13_148_4567_0, i_13_148_4594_0, i_13_148_4604_0,
    o_13_148_0_0  );
  input  i_13_148_61_0, i_13_148_71_0, i_13_148_179_0, i_13_148_274_0,
    i_13_148_275_0, i_13_148_280_0, i_13_148_286_0, i_13_148_493_0,
    i_13_148_529_0, i_13_148_530_0, i_13_148_553_0, i_13_148_562_0,
    i_13_148_599_0, i_13_148_673_0, i_13_148_797_0, i_13_148_841_0,
    i_13_148_853_0, i_13_148_854_0, i_13_148_965_0, i_13_148_1025_0,
    i_13_148_1075_0, i_13_148_1147_0, i_13_148_1282_0, i_13_148_1303_0,
    i_13_148_1304_0, i_13_148_1321_0, i_13_148_1327_0, i_13_148_1490_0,
    i_13_148_1502_0, i_13_148_1516_0, i_13_148_1552_0, i_13_148_1553_0,
    i_13_148_1660_0, i_13_148_1700_0, i_13_148_1817_0, i_13_148_1858_0,
    i_13_148_2002_0, i_13_148_2003_0, i_13_148_2020_0, i_13_148_2021_0,
    i_13_148_2050_0, i_13_148_2201_0, i_13_148_2240_0, i_13_148_2263_0,
    i_13_148_2275_0, i_13_148_2366_0, i_13_148_2461_0, i_13_148_2462_0,
    i_13_148_2470_0, i_13_148_2471_0, i_13_148_2509_0, i_13_148_2543_0,
    i_13_148_2551_0, i_13_148_2615_0, i_13_148_2653_0, i_13_148_2824_0,
    i_13_148_2825_0, i_13_148_2860_0, i_13_148_2920_0, i_13_148_2984_0,
    i_13_148_3173_0, i_13_148_3274_0, i_13_148_3347_0, i_13_148_3418_0,
    i_13_148_3424_0, i_13_148_3428_0, i_13_148_3482_0, i_13_148_3533_0,
    i_13_148_3541_0, i_13_148_3542_0, i_13_148_3544_0, i_13_148_3545_0,
    i_13_148_3580_0, i_13_148_3614_0, i_13_148_3622_0, i_13_148_3634_0,
    i_13_148_3730_0, i_13_148_3731_0, i_13_148_3743_0, i_13_148_3787_0,
    i_13_148_3788_0, i_13_148_3910_0, i_13_148_3911_0, i_13_148_3913_0,
    i_13_148_3914_0, i_13_148_4118_0, i_13_148_4126_0, i_13_148_4162_0,
    i_13_148_4189_0, i_13_148_4237_0, i_13_148_4238_0, i_13_148_4256_0,
    i_13_148_4282_0, i_13_148_4378_0, i_13_148_4381_0, i_13_148_4382_0,
    i_13_148_4400_0, i_13_148_4567_0, i_13_148_4594_0, i_13_148_4604_0;
  output o_13_148_0_0;
  assign o_13_148_0_0 = ~((~i_13_148_493_0 & ~i_13_148_1490_0) | (~i_13_148_3347_0 & ~i_13_148_3544_0 & ~i_13_148_4382_0) | (i_13_148_841_0 & i_13_148_2275_0 & ~i_13_148_3545_0 & ~i_13_148_3731_0 & ~i_13_148_3914_0));
endmodule



// Benchmark "kernel_13_149" written by ABC on Sun Jul 19 10:47:30 2020

module kernel_13_149 ( 
    i_13_149_63_0, i_13_149_207_0, i_13_149_265_0, i_13_149_306_0,
    i_13_149_354_0, i_13_149_370_0, i_13_149_372_0, i_13_149_381_0,
    i_13_149_409_0, i_13_149_414_0, i_13_149_462_0, i_13_149_463_0,
    i_13_149_466_0, i_13_149_467_0, i_13_149_588_0, i_13_149_589_0,
    i_13_149_595_0, i_13_149_660_0, i_13_149_666_0, i_13_149_670_0,
    i_13_149_697_0, i_13_149_759_0, i_13_149_948_0, i_13_149_1179_0,
    i_13_149_1344_0, i_13_149_1349_0, i_13_149_1549_0, i_13_149_1569_0,
    i_13_149_1594_0, i_13_149_1603_0, i_13_149_1767_0, i_13_149_1845_0,
    i_13_149_1846_0, i_13_149_1854_0, i_13_149_1947_0, i_13_149_1959_0,
    i_13_149_1993_0, i_13_149_2028_0, i_13_149_2029_0, i_13_149_2100_0,
    i_13_149_2137_0, i_13_149_2142_0, i_13_149_2199_0, i_13_149_2200_0,
    i_13_149_2204_0, i_13_149_2263_0, i_13_149_2280_0, i_13_149_2434_0,
    i_13_149_2457_0, i_13_149_2503_0, i_13_149_2506_0, i_13_149_2511_0,
    i_13_149_2554_0, i_13_149_2559_0, i_13_149_2820_0, i_13_149_2821_0,
    i_13_149_2856_0, i_13_149_2880_0, i_13_149_2982_0, i_13_149_3000_0,
    i_13_149_3001_0, i_13_149_3046_0, i_13_149_3130_0, i_13_149_3144_0,
    i_13_149_3213_0, i_13_149_3240_0, i_13_149_3241_0, i_13_149_3343_0,
    i_13_149_3387_0, i_13_149_3392_0, i_13_149_3411_0, i_13_149_3412_0,
    i_13_149_3480_0, i_13_149_3537_0, i_13_149_3538_0, i_13_149_3567_0,
    i_13_149_3592_0, i_13_149_3594_0, i_13_149_3595_0, i_13_149_3618_0,
    i_13_149_3619_0, i_13_149_3630_0, i_13_149_3631_0, i_13_149_3634_0,
    i_13_149_3636_0, i_13_149_3637_0, i_13_149_3666_0, i_13_149_3670_0,
    i_13_149_3766_0, i_13_149_3846_0, i_13_149_3906_0, i_13_149_3915_0,
    i_13_149_4060_0, i_13_149_4162_0, i_13_149_4269_0, i_13_149_4316_0,
    i_13_149_4324_0, i_13_149_4327_0, i_13_149_4368_0, i_13_149_4443_0,
    o_13_149_0_0  );
  input  i_13_149_63_0, i_13_149_207_0, i_13_149_265_0, i_13_149_306_0,
    i_13_149_354_0, i_13_149_370_0, i_13_149_372_0, i_13_149_381_0,
    i_13_149_409_0, i_13_149_414_0, i_13_149_462_0, i_13_149_463_0,
    i_13_149_466_0, i_13_149_467_0, i_13_149_588_0, i_13_149_589_0,
    i_13_149_595_0, i_13_149_660_0, i_13_149_666_0, i_13_149_670_0,
    i_13_149_697_0, i_13_149_759_0, i_13_149_948_0, i_13_149_1179_0,
    i_13_149_1344_0, i_13_149_1349_0, i_13_149_1549_0, i_13_149_1569_0,
    i_13_149_1594_0, i_13_149_1603_0, i_13_149_1767_0, i_13_149_1845_0,
    i_13_149_1846_0, i_13_149_1854_0, i_13_149_1947_0, i_13_149_1959_0,
    i_13_149_1993_0, i_13_149_2028_0, i_13_149_2029_0, i_13_149_2100_0,
    i_13_149_2137_0, i_13_149_2142_0, i_13_149_2199_0, i_13_149_2200_0,
    i_13_149_2204_0, i_13_149_2263_0, i_13_149_2280_0, i_13_149_2434_0,
    i_13_149_2457_0, i_13_149_2503_0, i_13_149_2506_0, i_13_149_2511_0,
    i_13_149_2554_0, i_13_149_2559_0, i_13_149_2820_0, i_13_149_2821_0,
    i_13_149_2856_0, i_13_149_2880_0, i_13_149_2982_0, i_13_149_3000_0,
    i_13_149_3001_0, i_13_149_3046_0, i_13_149_3130_0, i_13_149_3144_0,
    i_13_149_3213_0, i_13_149_3240_0, i_13_149_3241_0, i_13_149_3343_0,
    i_13_149_3387_0, i_13_149_3392_0, i_13_149_3411_0, i_13_149_3412_0,
    i_13_149_3480_0, i_13_149_3537_0, i_13_149_3538_0, i_13_149_3567_0,
    i_13_149_3592_0, i_13_149_3594_0, i_13_149_3595_0, i_13_149_3618_0,
    i_13_149_3619_0, i_13_149_3630_0, i_13_149_3631_0, i_13_149_3634_0,
    i_13_149_3636_0, i_13_149_3637_0, i_13_149_3666_0, i_13_149_3670_0,
    i_13_149_3766_0, i_13_149_3846_0, i_13_149_3906_0, i_13_149_3915_0,
    i_13_149_4060_0, i_13_149_4162_0, i_13_149_4269_0, i_13_149_4316_0,
    i_13_149_4324_0, i_13_149_4327_0, i_13_149_4368_0, i_13_149_4443_0;
  output o_13_149_0_0;
  assign o_13_149_0_0 = ~((~i_13_149_2856_0 & ~i_13_149_3537_0) | (~i_13_149_1846_0 & ~i_13_149_1947_0 & ~i_13_149_2200_0));
endmodule



// Benchmark "kernel_13_150" written by ABC on Sun Jul 19 10:47:31 2020

module kernel_13_150 ( 
    i_13_150_136_0, i_13_150_139_0, i_13_150_166_0, i_13_150_190_0,
    i_13_150_229_0, i_13_150_251_0, i_13_150_374_0, i_13_150_419_0,
    i_13_150_508_0, i_13_150_536_0, i_13_150_545_0, i_13_150_556_0,
    i_13_150_613_0, i_13_150_614_0, i_13_150_622_0, i_13_150_646_0,
    i_13_150_665_0, i_13_150_695_0, i_13_150_698_0, i_13_150_713_0,
    i_13_150_793_0, i_13_150_814_0, i_13_150_895_0, i_13_150_939_0,
    i_13_150_952_0, i_13_150_979_0, i_13_150_1021_0, i_13_150_1094_0,
    i_13_150_1117_0, i_13_150_1120_0, i_13_150_1130_0, i_13_150_1228_0,
    i_13_150_1249_0, i_13_150_1252_0, i_13_150_1273_0, i_13_150_1390_0,
    i_13_150_1467_0, i_13_150_1480_0, i_13_150_1484_0, i_13_150_1502_0,
    i_13_150_1642_0, i_13_150_1670_0, i_13_150_1675_0, i_13_150_1757_0,
    i_13_150_1759_0, i_13_150_1778_0, i_13_150_1795_0, i_13_150_1796_0,
    i_13_150_1825_0, i_13_150_1947_0, i_13_150_1960_0, i_13_150_2004_0,
    i_13_150_2030_0, i_13_150_2111_0, i_13_150_2245_0, i_13_150_2288_0,
    i_13_150_2380_0, i_13_150_2407_0, i_13_150_2408_0, i_13_150_2464_0,
    i_13_150_2552_0, i_13_150_2615_0, i_13_150_2747_0, i_13_150_2750_0,
    i_13_150_2767_0, i_13_150_2848_0, i_13_150_2849_0, i_13_150_2850_0,
    i_13_150_2851_0, i_13_150_2875_0, i_13_150_2882_0, i_13_150_2976_0,
    i_13_150_3088_0, i_13_150_3092_0, i_13_150_3116_0, i_13_150_3256_0,
    i_13_150_3368_0, i_13_150_3371_0, i_13_150_3460_0, i_13_150_3556_0,
    i_13_150_3638_0, i_13_150_3730_0, i_13_150_3794_0, i_13_150_3839_0,
    i_13_150_3929_0, i_13_150_3997_0, i_13_150_4055_0, i_13_150_4064_0,
    i_13_150_4117_0, i_13_150_4138_0, i_13_150_4186_0, i_13_150_4189_0,
    i_13_150_4190_0, i_13_150_4197_0, i_13_150_4294_0, i_13_150_4296_0,
    i_13_150_4297_0, i_13_150_4337_0, i_13_150_4344_0, i_13_150_4515_0,
    o_13_150_0_0  );
  input  i_13_150_136_0, i_13_150_139_0, i_13_150_166_0, i_13_150_190_0,
    i_13_150_229_0, i_13_150_251_0, i_13_150_374_0, i_13_150_419_0,
    i_13_150_508_0, i_13_150_536_0, i_13_150_545_0, i_13_150_556_0,
    i_13_150_613_0, i_13_150_614_0, i_13_150_622_0, i_13_150_646_0,
    i_13_150_665_0, i_13_150_695_0, i_13_150_698_0, i_13_150_713_0,
    i_13_150_793_0, i_13_150_814_0, i_13_150_895_0, i_13_150_939_0,
    i_13_150_952_0, i_13_150_979_0, i_13_150_1021_0, i_13_150_1094_0,
    i_13_150_1117_0, i_13_150_1120_0, i_13_150_1130_0, i_13_150_1228_0,
    i_13_150_1249_0, i_13_150_1252_0, i_13_150_1273_0, i_13_150_1390_0,
    i_13_150_1467_0, i_13_150_1480_0, i_13_150_1484_0, i_13_150_1502_0,
    i_13_150_1642_0, i_13_150_1670_0, i_13_150_1675_0, i_13_150_1757_0,
    i_13_150_1759_0, i_13_150_1778_0, i_13_150_1795_0, i_13_150_1796_0,
    i_13_150_1825_0, i_13_150_1947_0, i_13_150_1960_0, i_13_150_2004_0,
    i_13_150_2030_0, i_13_150_2111_0, i_13_150_2245_0, i_13_150_2288_0,
    i_13_150_2380_0, i_13_150_2407_0, i_13_150_2408_0, i_13_150_2464_0,
    i_13_150_2552_0, i_13_150_2615_0, i_13_150_2747_0, i_13_150_2750_0,
    i_13_150_2767_0, i_13_150_2848_0, i_13_150_2849_0, i_13_150_2850_0,
    i_13_150_2851_0, i_13_150_2875_0, i_13_150_2882_0, i_13_150_2976_0,
    i_13_150_3088_0, i_13_150_3092_0, i_13_150_3116_0, i_13_150_3256_0,
    i_13_150_3368_0, i_13_150_3371_0, i_13_150_3460_0, i_13_150_3556_0,
    i_13_150_3638_0, i_13_150_3730_0, i_13_150_3794_0, i_13_150_3839_0,
    i_13_150_3929_0, i_13_150_3997_0, i_13_150_4055_0, i_13_150_4064_0,
    i_13_150_4117_0, i_13_150_4138_0, i_13_150_4186_0, i_13_150_4189_0,
    i_13_150_4190_0, i_13_150_4197_0, i_13_150_4294_0, i_13_150_4296_0,
    i_13_150_4297_0, i_13_150_4337_0, i_13_150_4344_0, i_13_150_4515_0;
  output o_13_150_0_0;
  assign o_13_150_0_0 = ~((~i_13_150_698_0 & (~i_13_150_4186_0 | (~i_13_150_4055_0 & ~i_13_150_4190_0))) | (~i_13_150_4190_0 & ((~i_13_150_536_0 & ~i_13_150_695_0) | i_13_150_1252_0 | ~i_13_150_3088_0)) | i_13_150_814_0 | (~i_13_150_614_0 & ~i_13_150_1795_0) | (~i_13_150_613_0 & ~i_13_150_2851_0 & ~i_13_150_4064_0));
endmodule



// Benchmark "kernel_13_151" written by ABC on Sun Jul 19 10:47:31 2020

module kernel_13_151 ( 
    i_13_151_113_0, i_13_151_121_0, i_13_151_137_0, i_13_151_138_0,
    i_13_151_139_0, i_13_151_140_0, i_13_151_143_0, i_13_151_175_0,
    i_13_151_229_0, i_13_151_231_0, i_13_151_260_0, i_13_151_340_0,
    i_13_151_380_0, i_13_151_473_0, i_13_151_535_0, i_13_151_536_0,
    i_13_151_537_0, i_13_151_573_0, i_13_151_574_0, i_13_151_725_0,
    i_13_151_832_0, i_13_151_850_0, i_13_151_853_0, i_13_151_868_0,
    i_13_151_869_0, i_13_151_985_0, i_13_151_1216_0, i_13_151_1219_0,
    i_13_151_1228_0, i_13_151_1470_0, i_13_151_1475_0, i_13_151_1540_0,
    i_13_151_1546_0, i_13_151_1547_0, i_13_151_1552_0, i_13_151_1667_0,
    i_13_151_1711_0, i_13_151_1714_0, i_13_151_1715_0, i_13_151_1723_0,
    i_13_151_1724_0, i_13_151_1725_0, i_13_151_1726_0, i_13_151_1734_0,
    i_13_151_1787_0, i_13_151_1831_0, i_13_151_1840_0, i_13_151_1841_0,
    i_13_151_1849_0, i_13_151_1858_0, i_13_151_1940_0, i_13_151_1993_0,
    i_13_151_2128_0, i_13_151_2156_0, i_13_151_2158_0, i_13_151_2345_0,
    i_13_151_2467_0, i_13_151_2570_0, i_13_151_2692_0, i_13_151_2695_0,
    i_13_151_2701_0, i_13_151_2712_0, i_13_151_2845_0, i_13_151_2848_0,
    i_13_151_3010_0, i_13_151_3011_0, i_13_151_3037_0, i_13_151_3064_0,
    i_13_151_3065_0, i_13_151_3066_0, i_13_151_3109_0, i_13_151_3146_0,
    i_13_151_3174_0, i_13_151_3229_0, i_13_151_3293_0, i_13_151_3444_0,
    i_13_151_3452_0, i_13_151_3478_0, i_13_151_3487_0, i_13_151_3524_0,
    i_13_151_3541_0, i_13_151_3570_0, i_13_151_3686_0, i_13_151_3688_0,
    i_13_151_3701_0, i_13_151_3739_0, i_13_151_3799_0, i_13_151_3836_0,
    i_13_151_4054_0, i_13_151_4058_0, i_13_151_4063_0, i_13_151_4151_0,
    i_13_151_4193_0, i_13_151_4234_0, i_13_151_4369_0, i_13_151_4378_0,
    i_13_151_4394_0, i_13_151_4411_0, i_13_151_4415_0, i_13_151_4523_0,
    o_13_151_0_0  );
  input  i_13_151_113_0, i_13_151_121_0, i_13_151_137_0, i_13_151_138_0,
    i_13_151_139_0, i_13_151_140_0, i_13_151_143_0, i_13_151_175_0,
    i_13_151_229_0, i_13_151_231_0, i_13_151_260_0, i_13_151_340_0,
    i_13_151_380_0, i_13_151_473_0, i_13_151_535_0, i_13_151_536_0,
    i_13_151_537_0, i_13_151_573_0, i_13_151_574_0, i_13_151_725_0,
    i_13_151_832_0, i_13_151_850_0, i_13_151_853_0, i_13_151_868_0,
    i_13_151_869_0, i_13_151_985_0, i_13_151_1216_0, i_13_151_1219_0,
    i_13_151_1228_0, i_13_151_1470_0, i_13_151_1475_0, i_13_151_1540_0,
    i_13_151_1546_0, i_13_151_1547_0, i_13_151_1552_0, i_13_151_1667_0,
    i_13_151_1711_0, i_13_151_1714_0, i_13_151_1715_0, i_13_151_1723_0,
    i_13_151_1724_0, i_13_151_1725_0, i_13_151_1726_0, i_13_151_1734_0,
    i_13_151_1787_0, i_13_151_1831_0, i_13_151_1840_0, i_13_151_1841_0,
    i_13_151_1849_0, i_13_151_1858_0, i_13_151_1940_0, i_13_151_1993_0,
    i_13_151_2128_0, i_13_151_2156_0, i_13_151_2158_0, i_13_151_2345_0,
    i_13_151_2467_0, i_13_151_2570_0, i_13_151_2692_0, i_13_151_2695_0,
    i_13_151_2701_0, i_13_151_2712_0, i_13_151_2845_0, i_13_151_2848_0,
    i_13_151_3010_0, i_13_151_3011_0, i_13_151_3037_0, i_13_151_3064_0,
    i_13_151_3065_0, i_13_151_3066_0, i_13_151_3109_0, i_13_151_3146_0,
    i_13_151_3174_0, i_13_151_3229_0, i_13_151_3293_0, i_13_151_3444_0,
    i_13_151_3452_0, i_13_151_3478_0, i_13_151_3487_0, i_13_151_3524_0,
    i_13_151_3541_0, i_13_151_3570_0, i_13_151_3686_0, i_13_151_3688_0,
    i_13_151_3701_0, i_13_151_3739_0, i_13_151_3799_0, i_13_151_3836_0,
    i_13_151_4054_0, i_13_151_4058_0, i_13_151_4063_0, i_13_151_4151_0,
    i_13_151_4193_0, i_13_151_4234_0, i_13_151_4369_0, i_13_151_4378_0,
    i_13_151_4394_0, i_13_151_4411_0, i_13_151_4415_0, i_13_151_4523_0;
  output o_13_151_0_0;
  assign o_13_151_0_0 = ~((i_13_151_138_0 & i_13_151_4378_0 & (~i_13_151_1993_0 | (i_13_151_535_0 & ~i_13_151_1831_0))) | (~i_13_151_537_0 & ~i_13_151_4411_0 & ((~i_13_151_143_0 & ((~i_13_151_140_0 & ~i_13_151_573_0 & ~i_13_151_3064_0) | (~i_13_151_1216_0 & ~i_13_151_1714_0 & ~i_13_151_3686_0))) | (~i_13_151_113_0 & i_13_151_175_0 & i_13_151_2695_0 & ~i_13_151_2845_0 & ~i_13_151_4415_0))) | (~i_13_151_2845_0 & ((~i_13_151_3065_0 & ~i_13_151_3452_0 & i_13_151_3487_0) | (i_13_151_3011_0 & i_13_151_4151_0))) | (~i_13_151_3688_0 & (~i_13_151_139_0 | (~i_13_151_1216_0 & i_13_151_3037_0 & ~i_13_151_3444_0 & ~i_13_151_4378_0 & ~i_13_151_4415_0))) | (~i_13_151_536_0 & i_13_151_1552_0 & i_13_151_1831_0 & ~i_13_151_4394_0) | (~i_13_151_1219_0 & ~i_13_151_3524_0 & i_13_151_4411_0));
endmodule



// Benchmark "kernel_13_152" written by ABC on Sun Jul 19 10:47:33 2020

module kernel_13_152 ( 
    i_13_152_50_0, i_13_152_73_0, i_13_152_102_0, i_13_152_137_0,
    i_13_152_189_0, i_13_152_252_0, i_13_152_280_0, i_13_152_407_0,
    i_13_152_434_0, i_13_152_441_0, i_13_152_515_0, i_13_152_559_0,
    i_13_152_617_0, i_13_152_623_0, i_13_152_659_0, i_13_152_661_0,
    i_13_152_666_0, i_13_152_693_0, i_13_152_694_0, i_13_152_695_0,
    i_13_152_696_0, i_13_152_838_0, i_13_152_839_0, i_13_152_921_0,
    i_13_152_975_0, i_13_152_1072_0, i_13_152_1073_0, i_13_152_1109_0,
    i_13_152_1116_0, i_13_152_1117_0, i_13_152_1118_0, i_13_152_1145_0,
    i_13_152_1270_0, i_13_152_1423_0, i_13_152_1424_0, i_13_152_1427_0,
    i_13_152_1657_0, i_13_152_1658_0, i_13_152_1730_0, i_13_152_1742_0,
    i_13_152_1791_0, i_13_152_1858_0, i_13_152_2016_0, i_13_152_2017_0,
    i_13_152_2020_0, i_13_152_2021_0, i_13_152_2207_0, i_13_152_2209_0,
    i_13_152_2324_0, i_13_152_2344_0, i_13_152_2443_0, i_13_152_2452_0,
    i_13_152_2453_0, i_13_152_2461_0, i_13_152_2467_0, i_13_152_2512_0,
    i_13_152_2513_0, i_13_152_2551_0, i_13_152_2552_0, i_13_152_2718_0,
    i_13_152_2741_0, i_13_152_2880_0, i_13_152_2881_0, i_13_152_2882_0,
    i_13_152_2883_0, i_13_152_2956_0, i_13_152_3001_0, i_13_152_3074_0,
    i_13_152_3089_0, i_13_152_3091_0, i_13_152_3107_0, i_13_152_3269_0,
    i_13_152_3371_0, i_13_152_3416_0, i_13_152_3424_0, i_13_152_3476_0,
    i_13_152_3487_0, i_13_152_3532_0, i_13_152_3547_0, i_13_152_3646_0,
    i_13_152_3740_0, i_13_152_3820_0, i_13_152_3862_0, i_13_152_3919_0,
    i_13_152_3987_0, i_13_152_3989_0, i_13_152_4252_0, i_13_152_4293_0,
    i_13_152_4315_0, i_13_152_4324_0, i_13_152_4330_0, i_13_152_4331_0,
    i_13_152_4429_0, i_13_152_4450_0, i_13_152_4451_0, i_13_152_4455_0,
    i_13_152_4591_0, i_13_152_4592_0, i_13_152_4600_0, i_13_152_4601_0,
    o_13_152_0_0  );
  input  i_13_152_50_0, i_13_152_73_0, i_13_152_102_0, i_13_152_137_0,
    i_13_152_189_0, i_13_152_252_0, i_13_152_280_0, i_13_152_407_0,
    i_13_152_434_0, i_13_152_441_0, i_13_152_515_0, i_13_152_559_0,
    i_13_152_617_0, i_13_152_623_0, i_13_152_659_0, i_13_152_661_0,
    i_13_152_666_0, i_13_152_693_0, i_13_152_694_0, i_13_152_695_0,
    i_13_152_696_0, i_13_152_838_0, i_13_152_839_0, i_13_152_921_0,
    i_13_152_975_0, i_13_152_1072_0, i_13_152_1073_0, i_13_152_1109_0,
    i_13_152_1116_0, i_13_152_1117_0, i_13_152_1118_0, i_13_152_1145_0,
    i_13_152_1270_0, i_13_152_1423_0, i_13_152_1424_0, i_13_152_1427_0,
    i_13_152_1657_0, i_13_152_1658_0, i_13_152_1730_0, i_13_152_1742_0,
    i_13_152_1791_0, i_13_152_1858_0, i_13_152_2016_0, i_13_152_2017_0,
    i_13_152_2020_0, i_13_152_2021_0, i_13_152_2207_0, i_13_152_2209_0,
    i_13_152_2324_0, i_13_152_2344_0, i_13_152_2443_0, i_13_152_2452_0,
    i_13_152_2453_0, i_13_152_2461_0, i_13_152_2467_0, i_13_152_2512_0,
    i_13_152_2513_0, i_13_152_2551_0, i_13_152_2552_0, i_13_152_2718_0,
    i_13_152_2741_0, i_13_152_2880_0, i_13_152_2881_0, i_13_152_2882_0,
    i_13_152_2883_0, i_13_152_2956_0, i_13_152_3001_0, i_13_152_3074_0,
    i_13_152_3089_0, i_13_152_3091_0, i_13_152_3107_0, i_13_152_3269_0,
    i_13_152_3371_0, i_13_152_3416_0, i_13_152_3424_0, i_13_152_3476_0,
    i_13_152_3487_0, i_13_152_3532_0, i_13_152_3547_0, i_13_152_3646_0,
    i_13_152_3740_0, i_13_152_3820_0, i_13_152_3862_0, i_13_152_3919_0,
    i_13_152_3987_0, i_13_152_3989_0, i_13_152_4252_0, i_13_152_4293_0,
    i_13_152_4315_0, i_13_152_4324_0, i_13_152_4330_0, i_13_152_4331_0,
    i_13_152_4429_0, i_13_152_4450_0, i_13_152_4451_0, i_13_152_4455_0,
    i_13_152_4591_0, i_13_152_4592_0, i_13_152_4600_0, i_13_152_4601_0;
  output o_13_152_0_0;
  assign o_13_152_0_0 = ~((~i_13_152_694_0 & ((~i_13_152_1145_0 & i_13_152_3532_0) | (~i_13_152_693_0 & ~i_13_152_1424_0 & ~i_13_152_1658_0 & ~i_13_152_3989_0))) | i_13_152_4315_0 | (~i_13_152_1730_0 & ~i_13_152_3547_0 & ~i_13_152_4330_0));
endmodule



// Benchmark "kernel_13_153" written by ABC on Sun Jul 19 10:47:33 2020

module kernel_13_153 ( 
    i_13_153_138_0, i_13_153_139_0, i_13_153_184_0, i_13_153_226_0,
    i_13_153_280_0, i_13_153_380_0, i_13_153_415_0, i_13_153_524_0,
    i_13_153_585_0, i_13_153_651_0, i_13_153_675_0, i_13_153_832_0,
    i_13_153_1074_0, i_13_153_1182_0, i_13_153_1200_0, i_13_153_1206_0,
    i_13_153_1207_0, i_13_153_1252_0, i_13_153_1296_0, i_13_153_1297_0,
    i_13_153_1341_0, i_13_153_1342_0, i_13_153_1468_0, i_13_153_1515_0,
    i_13_153_1516_0, i_13_153_1711_0, i_13_153_1712_0, i_13_153_1720_0,
    i_13_153_1722_0, i_13_153_1723_0, i_13_153_1777_0, i_13_153_1778_0,
    i_13_153_1881_0, i_13_153_1882_0, i_13_153_1884_0, i_13_153_1923_0,
    i_13_153_1924_0, i_13_153_1926_0, i_13_153_1989_0, i_13_153_1990_0,
    i_13_153_1999_0, i_13_153_2001_0, i_13_153_2020_0, i_13_153_2052_0,
    i_13_153_2133_0, i_13_153_2134_0, i_13_153_2169_0, i_13_153_2277_0,
    i_13_153_2377_0, i_13_153_2470_0, i_13_153_2548_0, i_13_153_2646_0,
    i_13_153_2647_0, i_13_153_2676_0, i_13_153_2694_0, i_13_153_2710_0,
    i_13_153_2787_0, i_13_153_2853_0, i_13_153_2872_0, i_13_153_2934_0,
    i_13_153_2983_0, i_13_153_3037_0, i_13_153_3132_0, i_13_153_3208_0,
    i_13_153_3343_0, i_13_153_3384_0, i_13_153_3414_0, i_13_153_3415_0,
    i_13_153_3438_0, i_13_153_3445_0, i_13_153_3447_0, i_13_153_3448_0,
    i_13_153_3474_0, i_13_153_3475_0, i_13_153_3547_0, i_13_153_3592_0,
    i_13_153_3615_0, i_13_153_3616_0, i_13_153_3645_0, i_13_153_3646_0,
    i_13_153_3663_0, i_13_153_3684_0, i_13_153_3736_0, i_13_153_3820_0,
    i_13_153_3987_0, i_13_153_3988_0, i_13_153_4050_0, i_13_153_4053_0,
    i_13_153_4077_0, i_13_153_4117_0, i_13_153_4159_0, i_13_153_4203_0,
    i_13_153_4270_0, i_13_153_4338_0, i_13_153_4392_0, i_13_153_4393_0,
    i_13_153_4410_0, i_13_153_4411_0, i_13_153_4554_0, i_13_153_4567_0,
    o_13_153_0_0  );
  input  i_13_153_138_0, i_13_153_139_0, i_13_153_184_0, i_13_153_226_0,
    i_13_153_280_0, i_13_153_380_0, i_13_153_415_0, i_13_153_524_0,
    i_13_153_585_0, i_13_153_651_0, i_13_153_675_0, i_13_153_832_0,
    i_13_153_1074_0, i_13_153_1182_0, i_13_153_1200_0, i_13_153_1206_0,
    i_13_153_1207_0, i_13_153_1252_0, i_13_153_1296_0, i_13_153_1297_0,
    i_13_153_1341_0, i_13_153_1342_0, i_13_153_1468_0, i_13_153_1515_0,
    i_13_153_1516_0, i_13_153_1711_0, i_13_153_1712_0, i_13_153_1720_0,
    i_13_153_1722_0, i_13_153_1723_0, i_13_153_1777_0, i_13_153_1778_0,
    i_13_153_1881_0, i_13_153_1882_0, i_13_153_1884_0, i_13_153_1923_0,
    i_13_153_1924_0, i_13_153_1926_0, i_13_153_1989_0, i_13_153_1990_0,
    i_13_153_1999_0, i_13_153_2001_0, i_13_153_2020_0, i_13_153_2052_0,
    i_13_153_2133_0, i_13_153_2134_0, i_13_153_2169_0, i_13_153_2277_0,
    i_13_153_2377_0, i_13_153_2470_0, i_13_153_2548_0, i_13_153_2646_0,
    i_13_153_2647_0, i_13_153_2676_0, i_13_153_2694_0, i_13_153_2710_0,
    i_13_153_2787_0, i_13_153_2853_0, i_13_153_2872_0, i_13_153_2934_0,
    i_13_153_2983_0, i_13_153_3037_0, i_13_153_3132_0, i_13_153_3208_0,
    i_13_153_3343_0, i_13_153_3384_0, i_13_153_3414_0, i_13_153_3415_0,
    i_13_153_3438_0, i_13_153_3445_0, i_13_153_3447_0, i_13_153_3448_0,
    i_13_153_3474_0, i_13_153_3475_0, i_13_153_3547_0, i_13_153_3592_0,
    i_13_153_3615_0, i_13_153_3616_0, i_13_153_3645_0, i_13_153_3646_0,
    i_13_153_3663_0, i_13_153_3684_0, i_13_153_3736_0, i_13_153_3820_0,
    i_13_153_3987_0, i_13_153_3988_0, i_13_153_4050_0, i_13_153_4053_0,
    i_13_153_4077_0, i_13_153_4117_0, i_13_153_4159_0, i_13_153_4203_0,
    i_13_153_4270_0, i_13_153_4338_0, i_13_153_4392_0, i_13_153_4393_0,
    i_13_153_4410_0, i_13_153_4411_0, i_13_153_4554_0, i_13_153_4567_0;
  output o_13_153_0_0;
  assign o_13_153_0_0 = ~((~i_13_153_2646_0 & (~i_13_153_4393_0 | (~i_13_153_1206_0 & ~i_13_153_1712_0 & ~i_13_153_3438_0))) | (~i_13_153_280_0 & ~i_13_153_3438_0 & ~i_13_153_4392_0) | (~i_13_153_4053_0 & ~i_13_153_4411_0) | (~i_13_153_2277_0 & i_13_153_4567_0));
endmodule



// Benchmark "kernel_13_154" written by ABC on Sun Jul 19 10:47:34 2020

module kernel_13_154 ( 
    i_13_154_34_0, i_13_154_67_0, i_13_154_78_0, i_13_154_114_0,
    i_13_154_135_0, i_13_154_138_0, i_13_154_141_0, i_13_154_156_0,
    i_13_154_178_0, i_13_154_189_0, i_13_154_192_0, i_13_154_282_0,
    i_13_154_285_0, i_13_154_373_0, i_13_154_381_0, i_13_154_385_0,
    i_13_154_508_0, i_13_154_585_0, i_13_154_588_0, i_13_154_589_0,
    i_13_154_1119_0, i_13_154_1209_0, i_13_154_1281_0, i_13_154_1300_0,
    i_13_154_1312_0, i_13_154_1344_0, i_13_154_1399_0, i_13_154_1402_0,
    i_13_154_1407_0, i_13_154_1429_0, i_13_154_1443_0, i_13_154_1482_0,
    i_13_154_1515_0, i_13_154_1725_0, i_13_154_1770_0, i_13_154_1771_0,
    i_13_154_1778_0, i_13_154_1779_0, i_13_154_1812_0, i_13_154_1813_0,
    i_13_154_1884_0, i_13_154_1885_0, i_13_154_1888_0, i_13_154_1903_0,
    i_13_154_1924_0, i_13_154_1992_0, i_13_154_1995_0, i_13_154_2002_0,
    i_13_154_2004_0, i_13_154_2005_0, i_13_154_2020_0, i_13_154_2055_0,
    i_13_154_2118_0, i_13_154_2190_0, i_13_154_2193_0, i_13_154_2199_0,
    i_13_154_2235_0, i_13_154_2280_0, i_13_154_2281_0, i_13_154_2454_0,
    i_13_154_2595_0, i_13_154_2712_0, i_13_154_2721_0, i_13_154_2725_0,
    i_13_154_2726_0, i_13_154_2856_0, i_13_154_2857_0, i_13_154_2860_0,
    i_13_154_2899_0, i_13_154_2937_0, i_13_154_2959_0, i_13_154_3236_0,
    i_13_154_3274_0, i_13_154_3417_0, i_13_154_3418_0, i_13_154_3441_0,
    i_13_154_3453_0, i_13_154_3466_0, i_13_154_3477_0, i_13_154_3478_0,
    i_13_154_3481_0, i_13_154_3523_0, i_13_154_3595_0, i_13_154_3613_0,
    i_13_154_3666_0, i_13_154_3721_0, i_13_154_3729_0, i_13_154_3758_0,
    i_13_154_3769_0, i_13_154_3860_0, i_13_154_3897_0, i_13_154_3986_0,
    i_13_154_4017_0, i_13_154_4054_0, i_13_154_4217_0, i_13_154_4233_0,
    i_13_154_4395_0, i_13_154_4396_0, i_13_154_4399_0, i_13_154_4567_0,
    o_13_154_0_0  );
  input  i_13_154_34_0, i_13_154_67_0, i_13_154_78_0, i_13_154_114_0,
    i_13_154_135_0, i_13_154_138_0, i_13_154_141_0, i_13_154_156_0,
    i_13_154_178_0, i_13_154_189_0, i_13_154_192_0, i_13_154_282_0,
    i_13_154_285_0, i_13_154_373_0, i_13_154_381_0, i_13_154_385_0,
    i_13_154_508_0, i_13_154_585_0, i_13_154_588_0, i_13_154_589_0,
    i_13_154_1119_0, i_13_154_1209_0, i_13_154_1281_0, i_13_154_1300_0,
    i_13_154_1312_0, i_13_154_1344_0, i_13_154_1399_0, i_13_154_1402_0,
    i_13_154_1407_0, i_13_154_1429_0, i_13_154_1443_0, i_13_154_1482_0,
    i_13_154_1515_0, i_13_154_1725_0, i_13_154_1770_0, i_13_154_1771_0,
    i_13_154_1778_0, i_13_154_1779_0, i_13_154_1812_0, i_13_154_1813_0,
    i_13_154_1884_0, i_13_154_1885_0, i_13_154_1888_0, i_13_154_1903_0,
    i_13_154_1924_0, i_13_154_1992_0, i_13_154_1995_0, i_13_154_2002_0,
    i_13_154_2004_0, i_13_154_2005_0, i_13_154_2020_0, i_13_154_2055_0,
    i_13_154_2118_0, i_13_154_2190_0, i_13_154_2193_0, i_13_154_2199_0,
    i_13_154_2235_0, i_13_154_2280_0, i_13_154_2281_0, i_13_154_2454_0,
    i_13_154_2595_0, i_13_154_2712_0, i_13_154_2721_0, i_13_154_2725_0,
    i_13_154_2726_0, i_13_154_2856_0, i_13_154_2857_0, i_13_154_2860_0,
    i_13_154_2899_0, i_13_154_2937_0, i_13_154_2959_0, i_13_154_3236_0,
    i_13_154_3274_0, i_13_154_3417_0, i_13_154_3418_0, i_13_154_3441_0,
    i_13_154_3453_0, i_13_154_3466_0, i_13_154_3477_0, i_13_154_3478_0,
    i_13_154_3481_0, i_13_154_3523_0, i_13_154_3595_0, i_13_154_3613_0,
    i_13_154_3666_0, i_13_154_3721_0, i_13_154_3729_0, i_13_154_3758_0,
    i_13_154_3769_0, i_13_154_3860_0, i_13_154_3897_0, i_13_154_3986_0,
    i_13_154_4017_0, i_13_154_4054_0, i_13_154_4217_0, i_13_154_4233_0,
    i_13_154_4395_0, i_13_154_4396_0, i_13_154_4399_0, i_13_154_4567_0;
  output o_13_154_0_0;
  assign o_13_154_0_0 = ~(i_13_154_192_0 | (~i_13_154_2280_0 & ~i_13_154_4399_0) | (i_13_154_3523_0 & ~i_13_154_4395_0) | (~i_13_154_1300_0 & ~i_13_154_2004_0) | (~i_13_154_1813_0 & ~i_13_154_2937_0 & ~i_13_154_4396_0));
endmodule



// Benchmark "kernel_13_155" written by ABC on Sun Jul 19 10:47:35 2020

module kernel_13_155 ( 
    i_13_155_44_0, i_13_155_67_0, i_13_155_70_0, i_13_155_75_0,
    i_13_155_95_0, i_13_155_124_0, i_13_155_269_0, i_13_155_271_0,
    i_13_155_310_0, i_13_155_314_0, i_13_155_322_0, i_13_155_346_0,
    i_13_155_361_0, i_13_155_410_0, i_13_155_412_0, i_13_155_445_0,
    i_13_155_466_0, i_13_155_590_0, i_13_155_592_0, i_13_155_593_0,
    i_13_155_622_0, i_13_155_646_0, i_13_155_647_0, i_13_155_657_0,
    i_13_155_688_0, i_13_155_689_0, i_13_155_700_0, i_13_155_763_0,
    i_13_155_764_0, i_13_155_811_0, i_13_155_842_0, i_13_155_955_0,
    i_13_155_1120_0, i_13_155_1124_0, i_13_155_1132_0, i_13_155_1207_0,
    i_13_155_1261_0, i_13_155_1283_0, i_13_155_1285_0, i_13_155_1286_0,
    i_13_155_1312_0, i_13_155_1349_0, i_13_155_1511_0, i_13_155_1513_0,
    i_13_155_1601_0, i_13_155_1636_0, i_13_155_1728_0, i_13_155_1741_0,
    i_13_155_1754_0, i_13_155_1781_0, i_13_155_1799_0, i_13_155_1807_0,
    i_13_155_1997_0, i_13_155_2056_0, i_13_155_2057_0, i_13_155_2059_0,
    i_13_155_2060_0, i_13_155_2104_0, i_13_155_2123_0, i_13_155_2141_0,
    i_13_155_2195_0, i_13_155_2266_0, i_13_155_2267_0, i_13_155_2272_0,
    i_13_155_2377_0, i_13_155_2384_0, i_13_155_2426_0, i_13_155_2455_0,
    i_13_155_2512_0, i_13_155_2545_0, i_13_155_2555_0, i_13_155_2653_0,
    i_13_155_2680_0, i_13_155_2851_0, i_13_155_2939_0, i_13_155_3043_0,
    i_13_155_3175_0, i_13_155_3274_0, i_13_155_3346_0, i_13_155_3347_0,
    i_13_155_3391_0, i_13_155_3392_0, i_13_155_3640_0, i_13_155_3641_0,
    i_13_155_3722_0, i_13_155_3877_0, i_13_155_3905_0, i_13_155_3940_0,
    i_13_155_3994_0, i_13_155_4036_0, i_13_155_4037_0, i_13_155_4039_0,
    i_13_155_4040_0, i_13_155_4085_0, i_13_155_4144_0, i_13_155_4342_0,
    i_13_155_4382_0, i_13_155_4595_0, i_13_155_4597_0, i_13_155_4598_0,
    o_13_155_0_0  );
  input  i_13_155_44_0, i_13_155_67_0, i_13_155_70_0, i_13_155_75_0,
    i_13_155_95_0, i_13_155_124_0, i_13_155_269_0, i_13_155_271_0,
    i_13_155_310_0, i_13_155_314_0, i_13_155_322_0, i_13_155_346_0,
    i_13_155_361_0, i_13_155_410_0, i_13_155_412_0, i_13_155_445_0,
    i_13_155_466_0, i_13_155_590_0, i_13_155_592_0, i_13_155_593_0,
    i_13_155_622_0, i_13_155_646_0, i_13_155_647_0, i_13_155_657_0,
    i_13_155_688_0, i_13_155_689_0, i_13_155_700_0, i_13_155_763_0,
    i_13_155_764_0, i_13_155_811_0, i_13_155_842_0, i_13_155_955_0,
    i_13_155_1120_0, i_13_155_1124_0, i_13_155_1132_0, i_13_155_1207_0,
    i_13_155_1261_0, i_13_155_1283_0, i_13_155_1285_0, i_13_155_1286_0,
    i_13_155_1312_0, i_13_155_1349_0, i_13_155_1511_0, i_13_155_1513_0,
    i_13_155_1601_0, i_13_155_1636_0, i_13_155_1728_0, i_13_155_1741_0,
    i_13_155_1754_0, i_13_155_1781_0, i_13_155_1799_0, i_13_155_1807_0,
    i_13_155_1997_0, i_13_155_2056_0, i_13_155_2057_0, i_13_155_2059_0,
    i_13_155_2060_0, i_13_155_2104_0, i_13_155_2123_0, i_13_155_2141_0,
    i_13_155_2195_0, i_13_155_2266_0, i_13_155_2267_0, i_13_155_2272_0,
    i_13_155_2377_0, i_13_155_2384_0, i_13_155_2426_0, i_13_155_2455_0,
    i_13_155_2512_0, i_13_155_2545_0, i_13_155_2555_0, i_13_155_2653_0,
    i_13_155_2680_0, i_13_155_2851_0, i_13_155_2939_0, i_13_155_3043_0,
    i_13_155_3175_0, i_13_155_3274_0, i_13_155_3346_0, i_13_155_3347_0,
    i_13_155_3391_0, i_13_155_3392_0, i_13_155_3640_0, i_13_155_3641_0,
    i_13_155_3722_0, i_13_155_3877_0, i_13_155_3905_0, i_13_155_3940_0,
    i_13_155_3994_0, i_13_155_4036_0, i_13_155_4037_0, i_13_155_4039_0,
    i_13_155_4040_0, i_13_155_4085_0, i_13_155_4144_0, i_13_155_4342_0,
    i_13_155_4382_0, i_13_155_4595_0, i_13_155_4597_0, i_13_155_4598_0;
  output o_13_155_0_0;
  assign o_13_155_0_0 = ~((~i_13_155_592_0 & ~i_13_155_3391_0 & ((i_13_155_2056_0 & ~i_13_155_2272_0) | (~i_13_155_322_0 & ~i_13_155_4039_0))) | (~i_13_155_689_0 & ~i_13_155_2272_0 & i_13_155_3877_0) | (~i_13_155_763_0 & ~i_13_155_1511_0 & i_13_155_2272_0 & ~i_13_155_3347_0 & ~i_13_155_4085_0));
endmodule



// Benchmark "kernel_13_156" written by ABC on Sun Jul 19 10:47:36 2020

module kernel_13_156 ( 
    i_13_156_73_0, i_13_156_103_0, i_13_156_109_0, i_13_156_184_0,
    i_13_156_193_0, i_13_156_248_0, i_13_156_379_0, i_13_156_446_0,
    i_13_156_454_0, i_13_156_524_0, i_13_156_554_0, i_13_156_571_0,
    i_13_156_572_0, i_13_156_589_0, i_13_156_590_0, i_13_156_715_0,
    i_13_156_742_0, i_13_156_743_0, i_13_156_859_0, i_13_156_946_0,
    i_13_156_947_0, i_13_156_1021_0, i_13_156_1085_0, i_13_156_1140_0,
    i_13_156_1209_0, i_13_156_1228_0, i_13_156_1248_0, i_13_156_1255_0,
    i_13_156_1286_0, i_13_156_1345_0, i_13_156_1346_0, i_13_156_1397_0,
    i_13_156_1408_0, i_13_156_1427_0, i_13_156_1444_0, i_13_156_1571_0,
    i_13_156_1597_0, i_13_156_1607_0, i_13_156_1629_0, i_13_156_1678_0,
    i_13_156_1750_0, i_13_156_1777_0, i_13_156_1831_0, i_13_156_1858_0,
    i_13_156_1918_0, i_13_156_1930_0, i_13_156_1931_0, i_13_156_1940_0,
    i_13_156_1941_0, i_13_156_1948_0, i_13_156_1954_0, i_13_156_2002_0,
    i_13_156_2056_0, i_13_156_2057_0, i_13_156_2188_0, i_13_156_2281_0,
    i_13_156_2282_0, i_13_156_2299_0, i_13_156_2506_0, i_13_156_2512_0,
    i_13_156_2515_0, i_13_156_2614_0, i_13_156_2710_0, i_13_156_2713_0,
    i_13_156_2714_0, i_13_156_2719_0, i_13_156_2720_0, i_13_156_2723_0,
    i_13_156_2750_0, i_13_156_2768_0, i_13_156_2784_0, i_13_156_2785_0,
    i_13_156_2857_0, i_13_156_2858_0, i_13_156_2916_0, i_13_156_3065_0,
    i_13_156_3145_0, i_13_156_3154_0, i_13_156_3344_0, i_13_156_3370_0,
    i_13_156_3439_0, i_13_156_3596_0, i_13_156_3616_0, i_13_156_3617_0,
    i_13_156_3631_0, i_13_156_3681_0, i_13_156_3683_0, i_13_156_3685_0,
    i_13_156_3727_0, i_13_156_3920_0, i_13_156_3956_0, i_13_156_4037_0,
    i_13_156_4046_0, i_13_156_4091_0, i_13_156_4280_0, i_13_156_4330_0,
    i_13_156_4385_0, i_13_156_4396_0, i_13_156_4426_0, i_13_156_4555_0,
    o_13_156_0_0  );
  input  i_13_156_73_0, i_13_156_103_0, i_13_156_109_0, i_13_156_184_0,
    i_13_156_193_0, i_13_156_248_0, i_13_156_379_0, i_13_156_446_0,
    i_13_156_454_0, i_13_156_524_0, i_13_156_554_0, i_13_156_571_0,
    i_13_156_572_0, i_13_156_589_0, i_13_156_590_0, i_13_156_715_0,
    i_13_156_742_0, i_13_156_743_0, i_13_156_859_0, i_13_156_946_0,
    i_13_156_947_0, i_13_156_1021_0, i_13_156_1085_0, i_13_156_1140_0,
    i_13_156_1209_0, i_13_156_1228_0, i_13_156_1248_0, i_13_156_1255_0,
    i_13_156_1286_0, i_13_156_1345_0, i_13_156_1346_0, i_13_156_1397_0,
    i_13_156_1408_0, i_13_156_1427_0, i_13_156_1444_0, i_13_156_1571_0,
    i_13_156_1597_0, i_13_156_1607_0, i_13_156_1629_0, i_13_156_1678_0,
    i_13_156_1750_0, i_13_156_1777_0, i_13_156_1831_0, i_13_156_1858_0,
    i_13_156_1918_0, i_13_156_1930_0, i_13_156_1931_0, i_13_156_1940_0,
    i_13_156_1941_0, i_13_156_1948_0, i_13_156_1954_0, i_13_156_2002_0,
    i_13_156_2056_0, i_13_156_2057_0, i_13_156_2188_0, i_13_156_2281_0,
    i_13_156_2282_0, i_13_156_2299_0, i_13_156_2506_0, i_13_156_2512_0,
    i_13_156_2515_0, i_13_156_2614_0, i_13_156_2710_0, i_13_156_2713_0,
    i_13_156_2714_0, i_13_156_2719_0, i_13_156_2720_0, i_13_156_2723_0,
    i_13_156_2750_0, i_13_156_2768_0, i_13_156_2784_0, i_13_156_2785_0,
    i_13_156_2857_0, i_13_156_2858_0, i_13_156_2916_0, i_13_156_3065_0,
    i_13_156_3145_0, i_13_156_3154_0, i_13_156_3344_0, i_13_156_3370_0,
    i_13_156_3439_0, i_13_156_3596_0, i_13_156_3616_0, i_13_156_3617_0,
    i_13_156_3631_0, i_13_156_3681_0, i_13_156_3683_0, i_13_156_3685_0,
    i_13_156_3727_0, i_13_156_3920_0, i_13_156_3956_0, i_13_156_4037_0,
    i_13_156_4046_0, i_13_156_4091_0, i_13_156_4280_0, i_13_156_4330_0,
    i_13_156_4385_0, i_13_156_4396_0, i_13_156_4426_0, i_13_156_4555_0;
  output o_13_156_0_0;
  assign o_13_156_0_0 = ~((~i_13_156_3683_0 & ((~i_13_156_379_0 & ~i_13_156_2056_0) | (~i_13_156_524_0 & ~i_13_156_2858_0))) | (~i_13_156_4396_0 & (~i_13_156_3920_0 | (~i_13_156_2713_0 & ~i_13_156_2714_0 & ~i_13_156_3145_0))));
endmodule



// Benchmark "kernel_13_157" written by ABC on Sun Jul 19 10:47:36 2020

module kernel_13_157 ( 
    i_13_157_40_0, i_13_157_51_0, i_13_157_74_0, i_13_157_91_0,
    i_13_157_94_0, i_13_157_139_0, i_13_157_142_0, i_13_157_164_0,
    i_13_157_172_0, i_13_157_241_0, i_13_157_248_0, i_13_157_251_0,
    i_13_157_338_0, i_13_157_365_0, i_13_157_371_0, i_13_157_420_0,
    i_13_157_480_0, i_13_157_533_0, i_13_157_580_0, i_13_157_581_0,
    i_13_157_620_0, i_13_157_640_0, i_13_157_641_0, i_13_157_663_0,
    i_13_157_677_0, i_13_157_699_0, i_13_157_861_0, i_13_157_977_0,
    i_13_157_979_0, i_13_157_985_0, i_13_157_1098_0, i_13_157_1281_0,
    i_13_157_1284_0, i_13_157_1428_0, i_13_157_1462_0, i_13_157_1468_0,
    i_13_157_1487_0, i_13_157_1499_0, i_13_157_1553_0, i_13_157_1633_0,
    i_13_157_1634_0, i_13_157_1658_0, i_13_157_1720_0, i_13_157_1775_0,
    i_13_157_1885_0, i_13_157_1918_0, i_13_157_1990_0, i_13_157_1994_0,
    i_13_157_2050_0, i_13_157_2174_0, i_13_157_2348_0, i_13_157_2457_0,
    i_13_157_2507_0, i_13_157_2544_0, i_13_157_2552_0, i_13_157_2650_0,
    i_13_157_2788_0, i_13_157_2845_0, i_13_157_2846_0, i_13_157_2885_0,
    i_13_157_2888_0, i_13_157_2910_0, i_13_157_2924_0, i_13_157_2936_0,
    i_13_157_2949_0, i_13_157_2956_0, i_13_157_3208_0, i_13_157_3448_0,
    i_13_157_3449_0, i_13_157_3511_0, i_13_157_3524_0, i_13_157_3568_0,
    i_13_157_3572_0, i_13_157_3581_0, i_13_157_3638_0, i_13_157_3647_0,
    i_13_157_3652_0, i_13_157_3685_0, i_13_157_3686_0, i_13_157_3689_0,
    i_13_157_3736_0, i_13_157_3769_0, i_13_157_3847_0, i_13_157_3853_0,
    i_13_157_3905_0, i_13_157_3917_0, i_13_157_3988_0, i_13_157_4021_0,
    i_13_157_4036_0, i_13_157_4079_0, i_13_157_4088_0, i_13_157_4117_0,
    i_13_157_4260_0, i_13_157_4351_0, i_13_157_4352_0, i_13_157_4371_0,
    i_13_157_4391_0, i_13_157_4568_0, i_13_157_4576_0, i_13_157_4601_0,
    o_13_157_0_0  );
  input  i_13_157_40_0, i_13_157_51_0, i_13_157_74_0, i_13_157_91_0,
    i_13_157_94_0, i_13_157_139_0, i_13_157_142_0, i_13_157_164_0,
    i_13_157_172_0, i_13_157_241_0, i_13_157_248_0, i_13_157_251_0,
    i_13_157_338_0, i_13_157_365_0, i_13_157_371_0, i_13_157_420_0,
    i_13_157_480_0, i_13_157_533_0, i_13_157_580_0, i_13_157_581_0,
    i_13_157_620_0, i_13_157_640_0, i_13_157_641_0, i_13_157_663_0,
    i_13_157_677_0, i_13_157_699_0, i_13_157_861_0, i_13_157_977_0,
    i_13_157_979_0, i_13_157_985_0, i_13_157_1098_0, i_13_157_1281_0,
    i_13_157_1284_0, i_13_157_1428_0, i_13_157_1462_0, i_13_157_1468_0,
    i_13_157_1487_0, i_13_157_1499_0, i_13_157_1553_0, i_13_157_1633_0,
    i_13_157_1634_0, i_13_157_1658_0, i_13_157_1720_0, i_13_157_1775_0,
    i_13_157_1885_0, i_13_157_1918_0, i_13_157_1990_0, i_13_157_1994_0,
    i_13_157_2050_0, i_13_157_2174_0, i_13_157_2348_0, i_13_157_2457_0,
    i_13_157_2507_0, i_13_157_2544_0, i_13_157_2552_0, i_13_157_2650_0,
    i_13_157_2788_0, i_13_157_2845_0, i_13_157_2846_0, i_13_157_2885_0,
    i_13_157_2888_0, i_13_157_2910_0, i_13_157_2924_0, i_13_157_2936_0,
    i_13_157_2949_0, i_13_157_2956_0, i_13_157_3208_0, i_13_157_3448_0,
    i_13_157_3449_0, i_13_157_3511_0, i_13_157_3524_0, i_13_157_3568_0,
    i_13_157_3572_0, i_13_157_3581_0, i_13_157_3638_0, i_13_157_3647_0,
    i_13_157_3652_0, i_13_157_3685_0, i_13_157_3686_0, i_13_157_3689_0,
    i_13_157_3736_0, i_13_157_3769_0, i_13_157_3847_0, i_13_157_3853_0,
    i_13_157_3905_0, i_13_157_3917_0, i_13_157_3988_0, i_13_157_4021_0,
    i_13_157_4036_0, i_13_157_4079_0, i_13_157_4088_0, i_13_157_4117_0,
    i_13_157_4260_0, i_13_157_4351_0, i_13_157_4352_0, i_13_157_4371_0,
    i_13_157_4391_0, i_13_157_4568_0, i_13_157_4576_0, i_13_157_4601_0;
  output o_13_157_0_0;
  assign o_13_157_0_0 = ~((~i_13_157_4079_0 & ((~i_13_157_2845_0 & ~i_13_157_2885_0) | (~i_13_157_3685_0 & ~i_13_157_3736_0 & i_13_157_3847_0))) | (i_13_157_1553_0 & i_13_157_2174_0) | (i_13_157_2457_0 & i_13_157_3208_0) | (~i_13_157_620_0 & ~i_13_157_2457_0 & ~i_13_157_2846_0 & ~i_13_157_3449_0) | (~i_13_157_1885_0 & ~i_13_157_4088_0));
endmodule



// Benchmark "kernel_13_158" written by ABC on Sun Jul 19 10:47:37 2020

module kernel_13_158 ( 
    i_13_158_28_0, i_13_158_36_0, i_13_158_37_0, i_13_158_138_0,
    i_13_158_171_0, i_13_158_174_0, i_13_158_280_0, i_13_158_313_0,
    i_13_158_333_0, i_13_158_562_0, i_13_158_639_0, i_13_158_642_0,
    i_13_158_643_0, i_13_158_646_0, i_13_158_675_0, i_13_158_679_0,
    i_13_158_684_0, i_13_158_685_0, i_13_158_687_0, i_13_158_688_0,
    i_13_158_778_0, i_13_158_820_0, i_13_158_823_0, i_13_158_849_0,
    i_13_158_1119_0, i_13_158_1224_0, i_13_158_1269_0, i_13_158_1273_0,
    i_13_158_1305_0, i_13_158_1461_0, i_13_158_1521_0, i_13_158_1636_0,
    i_13_158_1668_0, i_13_158_1713_0, i_13_158_1749_0, i_13_158_1839_0,
    i_13_158_1855_0, i_13_158_1858_0, i_13_158_1881_0, i_13_158_1882_0,
    i_13_158_1884_0, i_13_158_2424_0, i_13_158_2457_0, i_13_158_2505_0,
    i_13_158_2559_0, i_13_158_2584_0, i_13_158_2646_0, i_13_158_2649_0,
    i_13_158_2650_0, i_13_158_2673_0, i_13_158_2677_0, i_13_158_2694_0,
    i_13_158_2730_0, i_13_158_2844_0, i_13_158_2847_0, i_13_158_2848_0,
    i_13_158_2874_0, i_13_158_2919_0, i_13_158_3088_0, i_13_158_3093_0,
    i_13_158_3094_0, i_13_158_3144_0, i_13_158_3234_0, i_13_158_3261_0,
    i_13_158_3270_0, i_13_158_3271_0, i_13_158_3304_0, i_13_158_3378_0,
    i_13_158_3387_0, i_13_158_3388_0, i_13_158_3420_0, i_13_158_3421_0,
    i_13_158_3423_0, i_13_158_3424_0, i_13_158_3429_0, i_13_158_3523_0,
    i_13_158_3561_0, i_13_158_3648_0, i_13_158_3721_0, i_13_158_3738_0,
    i_13_158_3798_0, i_13_158_3819_0, i_13_158_3924_0, i_13_158_3930_0,
    i_13_158_3987_0, i_13_158_4017_0, i_13_158_4036_0, i_13_158_4077_0,
    i_13_158_4080_0, i_13_158_4081_0, i_13_158_4185_0, i_13_158_4186_0,
    i_13_158_4257_0, i_13_158_4293_0, i_13_158_4339_0, i_13_158_4350_0,
    i_13_158_4465_0, i_13_158_4593_0, i_13_158_4594_0, i_13_158_4597_0,
    o_13_158_0_0  );
  input  i_13_158_28_0, i_13_158_36_0, i_13_158_37_0, i_13_158_138_0,
    i_13_158_171_0, i_13_158_174_0, i_13_158_280_0, i_13_158_313_0,
    i_13_158_333_0, i_13_158_562_0, i_13_158_639_0, i_13_158_642_0,
    i_13_158_643_0, i_13_158_646_0, i_13_158_675_0, i_13_158_679_0,
    i_13_158_684_0, i_13_158_685_0, i_13_158_687_0, i_13_158_688_0,
    i_13_158_778_0, i_13_158_820_0, i_13_158_823_0, i_13_158_849_0,
    i_13_158_1119_0, i_13_158_1224_0, i_13_158_1269_0, i_13_158_1273_0,
    i_13_158_1305_0, i_13_158_1461_0, i_13_158_1521_0, i_13_158_1636_0,
    i_13_158_1668_0, i_13_158_1713_0, i_13_158_1749_0, i_13_158_1839_0,
    i_13_158_1855_0, i_13_158_1858_0, i_13_158_1881_0, i_13_158_1882_0,
    i_13_158_1884_0, i_13_158_2424_0, i_13_158_2457_0, i_13_158_2505_0,
    i_13_158_2559_0, i_13_158_2584_0, i_13_158_2646_0, i_13_158_2649_0,
    i_13_158_2650_0, i_13_158_2673_0, i_13_158_2677_0, i_13_158_2694_0,
    i_13_158_2730_0, i_13_158_2844_0, i_13_158_2847_0, i_13_158_2848_0,
    i_13_158_2874_0, i_13_158_2919_0, i_13_158_3088_0, i_13_158_3093_0,
    i_13_158_3094_0, i_13_158_3144_0, i_13_158_3234_0, i_13_158_3261_0,
    i_13_158_3270_0, i_13_158_3271_0, i_13_158_3304_0, i_13_158_3378_0,
    i_13_158_3387_0, i_13_158_3388_0, i_13_158_3420_0, i_13_158_3421_0,
    i_13_158_3423_0, i_13_158_3424_0, i_13_158_3429_0, i_13_158_3523_0,
    i_13_158_3561_0, i_13_158_3648_0, i_13_158_3721_0, i_13_158_3738_0,
    i_13_158_3798_0, i_13_158_3819_0, i_13_158_3924_0, i_13_158_3930_0,
    i_13_158_3987_0, i_13_158_4017_0, i_13_158_4036_0, i_13_158_4077_0,
    i_13_158_4080_0, i_13_158_4081_0, i_13_158_4185_0, i_13_158_4186_0,
    i_13_158_4257_0, i_13_158_4293_0, i_13_158_4339_0, i_13_158_4350_0,
    i_13_158_4465_0, i_13_158_4593_0, i_13_158_4594_0, i_13_158_4597_0;
  output o_13_158_0_0;
  assign o_13_158_0_0 = ~((~i_13_158_685_0 & ~i_13_158_2649_0 & ~i_13_158_3930_0) | (~i_13_158_675_0 & ~i_13_158_1884_0 & ~i_13_158_3819_0));
endmodule



// Benchmark "kernel_13_159" written by ABC on Sun Jul 19 10:47:38 2020

module kernel_13_159 ( 
    i_13_159_67_0, i_13_159_74_0, i_13_159_121_0, i_13_159_122_0,
    i_13_159_140_0, i_13_159_281_0, i_13_159_325_0, i_13_159_373_0,
    i_13_159_379_0, i_13_159_406_0, i_13_159_442_0, i_13_159_443_0,
    i_13_159_463_0, i_13_159_532_0, i_13_159_589_0, i_13_159_622_0,
    i_13_159_641_0, i_13_159_677_0, i_13_159_715_0, i_13_159_742_0,
    i_13_159_760_0, i_13_159_769_0, i_13_159_814_0, i_13_159_820_0,
    i_13_159_821_0, i_13_159_824_0, i_13_159_859_0, i_13_159_860_0,
    i_13_159_919_0, i_13_159_928_0, i_13_159_929_0, i_13_159_959_0,
    i_13_159_1030_0, i_13_159_1066_0, i_13_159_1082_0, i_13_159_1100_0,
    i_13_159_1129_0, i_13_159_1196_0, i_13_159_1226_0, i_13_159_1250_0,
    i_13_159_1256_0, i_13_159_1301_0, i_13_159_1331_0, i_13_159_1489_0,
    i_13_159_1490_0, i_13_159_1642_0, i_13_159_1712_0, i_13_159_1751_0,
    i_13_159_1793_0, i_13_159_1804_0, i_13_159_1883_0, i_13_159_1942_0,
    i_13_159_1990_0, i_13_159_1991_0, i_13_159_2012_0, i_13_159_2056_0,
    i_13_159_2117_0, i_13_159_2260_0, i_13_159_2263_0, i_13_159_2344_0,
    i_13_159_2380_0, i_13_159_2470_0, i_13_159_2542_0, i_13_159_2611_0,
    i_13_159_2675_0, i_13_159_2767_0, i_13_159_2768_0, i_13_159_2846_0,
    i_13_159_2920_0, i_13_159_2983_0, i_13_159_3004_0, i_13_159_3019_0,
    i_13_159_3110_0, i_13_159_3164_0, i_13_159_3259_0, i_13_159_3286_0,
    i_13_159_3287_0, i_13_159_3343_0, i_13_159_3386_0, i_13_159_3416_0,
    i_13_159_3421_0, i_13_159_3422_0, i_13_159_3430_0, i_13_159_3434_0,
    i_13_159_3502_0, i_13_159_3503_0, i_13_159_3731_0, i_13_159_3736_0,
    i_13_159_3740_0, i_13_159_3794_0, i_13_159_3802_0, i_13_159_3874_0,
    i_13_159_3890_0, i_13_159_3892_0, i_13_159_3898_0, i_13_159_3919_0,
    i_13_159_4078_0, i_13_159_4079_0, i_13_159_4270_0, i_13_159_4595_0,
    o_13_159_0_0  );
  input  i_13_159_67_0, i_13_159_74_0, i_13_159_121_0, i_13_159_122_0,
    i_13_159_140_0, i_13_159_281_0, i_13_159_325_0, i_13_159_373_0,
    i_13_159_379_0, i_13_159_406_0, i_13_159_442_0, i_13_159_443_0,
    i_13_159_463_0, i_13_159_532_0, i_13_159_589_0, i_13_159_622_0,
    i_13_159_641_0, i_13_159_677_0, i_13_159_715_0, i_13_159_742_0,
    i_13_159_760_0, i_13_159_769_0, i_13_159_814_0, i_13_159_820_0,
    i_13_159_821_0, i_13_159_824_0, i_13_159_859_0, i_13_159_860_0,
    i_13_159_919_0, i_13_159_928_0, i_13_159_929_0, i_13_159_959_0,
    i_13_159_1030_0, i_13_159_1066_0, i_13_159_1082_0, i_13_159_1100_0,
    i_13_159_1129_0, i_13_159_1196_0, i_13_159_1226_0, i_13_159_1250_0,
    i_13_159_1256_0, i_13_159_1301_0, i_13_159_1331_0, i_13_159_1489_0,
    i_13_159_1490_0, i_13_159_1642_0, i_13_159_1712_0, i_13_159_1751_0,
    i_13_159_1793_0, i_13_159_1804_0, i_13_159_1883_0, i_13_159_1942_0,
    i_13_159_1990_0, i_13_159_1991_0, i_13_159_2012_0, i_13_159_2056_0,
    i_13_159_2117_0, i_13_159_2260_0, i_13_159_2263_0, i_13_159_2344_0,
    i_13_159_2380_0, i_13_159_2470_0, i_13_159_2542_0, i_13_159_2611_0,
    i_13_159_2675_0, i_13_159_2767_0, i_13_159_2768_0, i_13_159_2846_0,
    i_13_159_2920_0, i_13_159_2983_0, i_13_159_3004_0, i_13_159_3019_0,
    i_13_159_3110_0, i_13_159_3164_0, i_13_159_3259_0, i_13_159_3286_0,
    i_13_159_3287_0, i_13_159_3343_0, i_13_159_3386_0, i_13_159_3416_0,
    i_13_159_3421_0, i_13_159_3422_0, i_13_159_3430_0, i_13_159_3434_0,
    i_13_159_3502_0, i_13_159_3503_0, i_13_159_3731_0, i_13_159_3736_0,
    i_13_159_3740_0, i_13_159_3794_0, i_13_159_3802_0, i_13_159_3874_0,
    i_13_159_3890_0, i_13_159_3892_0, i_13_159_3898_0, i_13_159_3919_0,
    i_13_159_4078_0, i_13_159_4079_0, i_13_159_4270_0, i_13_159_4595_0;
  output o_13_159_0_0;
  assign o_13_159_0_0 = ~((~i_13_159_4079_0 & ((~i_13_159_1883_0 & ~i_13_159_3110_0) | (~i_13_159_3422_0 & i_13_159_4270_0))) | (~i_13_159_677_0 & ~i_13_159_929_0 & ~i_13_159_1712_0 & ~i_13_159_2846_0 & ~i_13_159_3731_0) | (~i_13_159_325_0 & ~i_13_159_928_0 & ~i_13_159_3736_0));
endmodule



// Benchmark "kernel_13_160" written by ABC on Sun Jul 19 10:47:39 2020

module kernel_13_160 ( 
    i_13_160_38_0, i_13_160_71_0, i_13_160_95_0, i_13_160_201_0,
    i_13_160_233_0, i_13_160_263_0, i_13_160_308_0, i_13_160_337_0,
    i_13_160_344_0, i_13_160_412_0, i_13_160_527_0, i_13_160_533_0,
    i_13_160_556_0, i_13_160_628_0, i_13_160_643_0, i_13_160_646_0,
    i_13_160_653_0, i_13_160_666_0, i_13_160_683_0, i_13_160_712_0,
    i_13_160_827_0, i_13_160_845_0, i_13_160_897_0, i_13_160_956_0,
    i_13_160_979_0, i_13_160_1120_0, i_13_160_1123_0, i_13_160_1155_0,
    i_13_160_1275_0, i_13_160_1276_0, i_13_160_1312_0, i_13_160_1333_0,
    i_13_160_1381_0, i_13_160_1390_0, i_13_160_1447_0, i_13_160_1462_0,
    i_13_160_1482_0, i_13_160_1499_0, i_13_160_1561_0, i_13_160_1570_0,
    i_13_160_1600_0, i_13_160_1645_0, i_13_160_1646_0, i_13_160_1664_0,
    i_13_160_1670_0, i_13_160_1678_0, i_13_160_1727_0, i_13_160_1753_0,
    i_13_160_1797_0, i_13_160_1882_0, i_13_160_1953_0, i_13_160_2040_0,
    i_13_160_2074_0, i_13_160_2231_0, i_13_160_2277_0, i_13_160_2310_0,
    i_13_160_2315_0, i_13_160_2378_0, i_13_160_2381_0, i_13_160_2384_0,
    i_13_160_2434_0, i_13_160_2548_0, i_13_160_2549_0, i_13_160_2570_0,
    i_13_160_2616_0, i_13_160_2634_0, i_13_160_2686_0, i_13_160_2687_0,
    i_13_160_2887_0, i_13_160_3082_0, i_13_160_3087_0, i_13_160_3197_0,
    i_13_160_3214_0, i_13_160_3241_0, i_13_160_3296_0, i_13_160_3355_0,
    i_13_160_3435_0, i_13_160_3597_0, i_13_160_3652_0, i_13_160_3739_0,
    i_13_160_3743_0, i_13_160_3781_0, i_13_160_3786_0, i_13_160_3838_0,
    i_13_160_3994_0, i_13_160_4063_0, i_13_160_4083_0, i_13_160_4097_0,
    i_13_160_4187_0, i_13_160_4296_0, i_13_160_4351_0, i_13_160_4369_0,
    i_13_160_4381_0, i_13_160_4418_0, i_13_160_4502_0, i_13_160_4558_0,
    i_13_160_4590_0, i_13_160_4595_0, i_13_160_4601_0, i_13_160_4605_0,
    o_13_160_0_0  );
  input  i_13_160_38_0, i_13_160_71_0, i_13_160_95_0, i_13_160_201_0,
    i_13_160_233_0, i_13_160_263_0, i_13_160_308_0, i_13_160_337_0,
    i_13_160_344_0, i_13_160_412_0, i_13_160_527_0, i_13_160_533_0,
    i_13_160_556_0, i_13_160_628_0, i_13_160_643_0, i_13_160_646_0,
    i_13_160_653_0, i_13_160_666_0, i_13_160_683_0, i_13_160_712_0,
    i_13_160_827_0, i_13_160_845_0, i_13_160_897_0, i_13_160_956_0,
    i_13_160_979_0, i_13_160_1120_0, i_13_160_1123_0, i_13_160_1155_0,
    i_13_160_1275_0, i_13_160_1276_0, i_13_160_1312_0, i_13_160_1333_0,
    i_13_160_1381_0, i_13_160_1390_0, i_13_160_1447_0, i_13_160_1462_0,
    i_13_160_1482_0, i_13_160_1499_0, i_13_160_1561_0, i_13_160_1570_0,
    i_13_160_1600_0, i_13_160_1645_0, i_13_160_1646_0, i_13_160_1664_0,
    i_13_160_1670_0, i_13_160_1678_0, i_13_160_1727_0, i_13_160_1753_0,
    i_13_160_1797_0, i_13_160_1882_0, i_13_160_1953_0, i_13_160_2040_0,
    i_13_160_2074_0, i_13_160_2231_0, i_13_160_2277_0, i_13_160_2310_0,
    i_13_160_2315_0, i_13_160_2378_0, i_13_160_2381_0, i_13_160_2384_0,
    i_13_160_2434_0, i_13_160_2548_0, i_13_160_2549_0, i_13_160_2570_0,
    i_13_160_2616_0, i_13_160_2634_0, i_13_160_2686_0, i_13_160_2687_0,
    i_13_160_2887_0, i_13_160_3082_0, i_13_160_3087_0, i_13_160_3197_0,
    i_13_160_3214_0, i_13_160_3241_0, i_13_160_3296_0, i_13_160_3355_0,
    i_13_160_3435_0, i_13_160_3597_0, i_13_160_3652_0, i_13_160_3739_0,
    i_13_160_3743_0, i_13_160_3781_0, i_13_160_3786_0, i_13_160_3838_0,
    i_13_160_3994_0, i_13_160_4063_0, i_13_160_4083_0, i_13_160_4097_0,
    i_13_160_4187_0, i_13_160_4296_0, i_13_160_4351_0, i_13_160_4369_0,
    i_13_160_4381_0, i_13_160_4418_0, i_13_160_4502_0, i_13_160_4558_0,
    i_13_160_4590_0, i_13_160_4595_0, i_13_160_4601_0, i_13_160_4605_0;
  output o_13_160_0_0;
  assign o_13_160_0_0 = 0;
endmodule



// Benchmark "kernel_13_161" written by ABC on Sun Jul 19 10:47:40 2020

module kernel_13_161 ( 
    i_13_161_57_0, i_13_161_76_0, i_13_161_79_0, i_13_161_111_0,
    i_13_161_177_0, i_13_161_243_0, i_13_161_265_0, i_13_161_411_0,
    i_13_161_606_0, i_13_161_607_0, i_13_161_609_0, i_13_161_628_0,
    i_13_161_657_0, i_13_161_660_0, i_13_161_661_0, i_13_161_663_0,
    i_13_161_669_0, i_13_161_850_0, i_13_161_915_0, i_13_161_942_0,
    i_13_161_947_0, i_13_161_1018_0, i_13_161_1020_0, i_13_161_1023_0,
    i_13_161_1060_0, i_13_161_1075_0, i_13_161_1134_0, i_13_161_1150_0,
    i_13_161_1213_0, i_13_161_1317_0, i_13_161_1425_0, i_13_161_1426_0,
    i_13_161_1428_0, i_13_161_1429_0, i_13_161_1571_0, i_13_161_1597_0,
    i_13_161_1632_0, i_13_161_1732_0, i_13_161_1849_0, i_13_161_1857_0,
    i_13_161_1858_0, i_13_161_2022_0, i_13_161_2023_0, i_13_161_2373_0,
    i_13_161_2407_0, i_13_161_2451_0, i_13_161_2454_0, i_13_161_2455_0,
    i_13_161_2498_0, i_13_161_2572_0, i_13_161_2740_0, i_13_161_2908_0,
    i_13_161_2938_0, i_13_161_3009_0, i_13_161_3012_0, i_13_161_3016_0,
    i_13_161_3124_0, i_13_161_3145_0, i_13_161_3148_0, i_13_161_3175_0,
    i_13_161_3250_0, i_13_161_3264_0, i_13_161_3273_0, i_13_161_3321_0,
    i_13_161_3403_0, i_13_161_3459_0, i_13_161_3486_0, i_13_161_3487_0,
    i_13_161_3530_0, i_13_161_3570_0, i_13_161_3640_0, i_13_161_3706_0,
    i_13_161_3783_0, i_13_161_3790_0, i_13_161_3864_0, i_13_161_3865_0,
    i_13_161_3894_0, i_13_161_3990_0, i_13_161_4021_0, i_13_161_4054_0,
    i_13_161_4057_0, i_13_161_4083_0, i_13_161_4095_0, i_13_161_4117_0,
    i_13_161_4119_0, i_13_161_4189_0, i_13_161_4252_0, i_13_161_4254_0,
    i_13_161_4255_0, i_13_161_4261_0, i_13_161_4263_0, i_13_161_4327_0,
    i_13_161_4368_0, i_13_161_4369_0, i_13_161_4370_0, i_13_161_4371_0,
    i_13_161_4471_0, i_13_161_4557_0, i_13_161_4560_0, i_13_161_4596_0,
    o_13_161_0_0  );
  input  i_13_161_57_0, i_13_161_76_0, i_13_161_79_0, i_13_161_111_0,
    i_13_161_177_0, i_13_161_243_0, i_13_161_265_0, i_13_161_411_0,
    i_13_161_606_0, i_13_161_607_0, i_13_161_609_0, i_13_161_628_0,
    i_13_161_657_0, i_13_161_660_0, i_13_161_661_0, i_13_161_663_0,
    i_13_161_669_0, i_13_161_850_0, i_13_161_915_0, i_13_161_942_0,
    i_13_161_947_0, i_13_161_1018_0, i_13_161_1020_0, i_13_161_1023_0,
    i_13_161_1060_0, i_13_161_1075_0, i_13_161_1134_0, i_13_161_1150_0,
    i_13_161_1213_0, i_13_161_1317_0, i_13_161_1425_0, i_13_161_1426_0,
    i_13_161_1428_0, i_13_161_1429_0, i_13_161_1571_0, i_13_161_1597_0,
    i_13_161_1632_0, i_13_161_1732_0, i_13_161_1849_0, i_13_161_1857_0,
    i_13_161_1858_0, i_13_161_2022_0, i_13_161_2023_0, i_13_161_2373_0,
    i_13_161_2407_0, i_13_161_2451_0, i_13_161_2454_0, i_13_161_2455_0,
    i_13_161_2498_0, i_13_161_2572_0, i_13_161_2740_0, i_13_161_2908_0,
    i_13_161_2938_0, i_13_161_3009_0, i_13_161_3012_0, i_13_161_3016_0,
    i_13_161_3124_0, i_13_161_3145_0, i_13_161_3148_0, i_13_161_3175_0,
    i_13_161_3250_0, i_13_161_3264_0, i_13_161_3273_0, i_13_161_3321_0,
    i_13_161_3403_0, i_13_161_3459_0, i_13_161_3486_0, i_13_161_3487_0,
    i_13_161_3530_0, i_13_161_3570_0, i_13_161_3640_0, i_13_161_3706_0,
    i_13_161_3783_0, i_13_161_3790_0, i_13_161_3864_0, i_13_161_3865_0,
    i_13_161_3894_0, i_13_161_3990_0, i_13_161_4021_0, i_13_161_4054_0,
    i_13_161_4057_0, i_13_161_4083_0, i_13_161_4095_0, i_13_161_4117_0,
    i_13_161_4119_0, i_13_161_4189_0, i_13_161_4252_0, i_13_161_4254_0,
    i_13_161_4255_0, i_13_161_4261_0, i_13_161_4263_0, i_13_161_4327_0,
    i_13_161_4368_0, i_13_161_4369_0, i_13_161_4370_0, i_13_161_4371_0,
    i_13_161_4471_0, i_13_161_4557_0, i_13_161_4560_0, i_13_161_4596_0;
  output o_13_161_0_0;
  assign o_13_161_0_0 = ~((~i_13_161_1213_0 & ~i_13_161_4255_0) | (~i_13_161_3148_0 & ~i_13_161_4368_0 & ~i_13_161_4371_0) | (~i_13_161_3459_0 & ~i_13_161_3570_0 & ~i_13_161_3783_0));
endmodule



// Benchmark "kernel_13_162" written by ABC on Sun Jul 19 10:47:41 2020

module kernel_13_162 ( 
    i_13_162_91_0, i_13_162_92_0, i_13_162_94_0, i_13_162_95_0,
    i_13_162_102_0, i_13_162_120_0, i_13_162_185_0, i_13_162_200_0,
    i_13_162_308_0, i_13_162_316_0, i_13_162_317_0, i_13_162_335_0,
    i_13_162_571_0, i_13_162_572_0, i_13_162_617_0, i_13_162_651_0,
    i_13_162_668_0, i_13_162_671_0, i_13_162_730_0, i_13_162_794_0,
    i_13_162_947_0, i_13_162_950_0, i_13_162_1064_0, i_13_162_1067_0,
    i_13_162_1093_0, i_13_162_1202_0, i_13_162_1210_0, i_13_162_1211_0,
    i_13_162_1229_0, i_13_162_1307_0, i_13_162_1318_0, i_13_162_1324_0,
    i_13_162_1325_0, i_13_162_1405_0, i_13_162_1426_0, i_13_162_1497_0,
    i_13_162_1514_0, i_13_162_1526_0, i_13_162_1595_0, i_13_162_1631_0,
    i_13_162_1642_0, i_13_162_1730_0, i_13_162_1757_0, i_13_162_1765_0,
    i_13_162_1802_0, i_13_162_1812_0, i_13_162_1828_0, i_13_162_1829_0,
    i_13_162_1850_0, i_13_162_1885_0, i_13_162_2108_0, i_13_162_2117_0,
    i_13_162_2128_0, i_13_162_2136_0, i_13_162_2206_0, i_13_162_2234_0,
    i_13_162_2261_0, i_13_162_2264_0, i_13_162_2444_0, i_13_162_2506_0,
    i_13_162_2539_0, i_13_162_2674_0, i_13_162_2919_0, i_13_162_3109_0,
    i_13_162_3110_0, i_13_162_3116_0, i_13_162_3164_0, i_13_162_3208_0,
    i_13_162_3209_0, i_13_162_3242_0, i_13_162_3258_0, i_13_162_3286_0,
    i_13_162_3395_0, i_13_162_3407_0, i_13_162_3415_0, i_13_162_3416_0,
    i_13_162_3422_0, i_13_162_3530_0, i_13_162_3766_0, i_13_162_3767_0,
    i_13_162_3783_0, i_13_162_3785_0, i_13_162_3817_0, i_13_162_3818_0,
    i_13_162_3872_0, i_13_162_3924_0, i_13_162_3925_0, i_13_162_3987_0,
    i_13_162_3988_0, i_13_162_4061_0, i_13_162_4132_0, i_13_162_4280_0,
    i_13_162_4339_0, i_13_162_4342_0, i_13_162_4351_0, i_13_162_4352_0,
    i_13_162_4379_0, i_13_162_4567_0, i_13_162_4568_0, i_13_162_4591_0,
    o_13_162_0_0  );
  input  i_13_162_91_0, i_13_162_92_0, i_13_162_94_0, i_13_162_95_0,
    i_13_162_102_0, i_13_162_120_0, i_13_162_185_0, i_13_162_200_0,
    i_13_162_308_0, i_13_162_316_0, i_13_162_317_0, i_13_162_335_0,
    i_13_162_571_0, i_13_162_572_0, i_13_162_617_0, i_13_162_651_0,
    i_13_162_668_0, i_13_162_671_0, i_13_162_730_0, i_13_162_794_0,
    i_13_162_947_0, i_13_162_950_0, i_13_162_1064_0, i_13_162_1067_0,
    i_13_162_1093_0, i_13_162_1202_0, i_13_162_1210_0, i_13_162_1211_0,
    i_13_162_1229_0, i_13_162_1307_0, i_13_162_1318_0, i_13_162_1324_0,
    i_13_162_1325_0, i_13_162_1405_0, i_13_162_1426_0, i_13_162_1497_0,
    i_13_162_1514_0, i_13_162_1526_0, i_13_162_1595_0, i_13_162_1631_0,
    i_13_162_1642_0, i_13_162_1730_0, i_13_162_1757_0, i_13_162_1765_0,
    i_13_162_1802_0, i_13_162_1812_0, i_13_162_1828_0, i_13_162_1829_0,
    i_13_162_1850_0, i_13_162_1885_0, i_13_162_2108_0, i_13_162_2117_0,
    i_13_162_2128_0, i_13_162_2136_0, i_13_162_2206_0, i_13_162_2234_0,
    i_13_162_2261_0, i_13_162_2264_0, i_13_162_2444_0, i_13_162_2506_0,
    i_13_162_2539_0, i_13_162_2674_0, i_13_162_2919_0, i_13_162_3109_0,
    i_13_162_3110_0, i_13_162_3116_0, i_13_162_3164_0, i_13_162_3208_0,
    i_13_162_3209_0, i_13_162_3242_0, i_13_162_3258_0, i_13_162_3286_0,
    i_13_162_3395_0, i_13_162_3407_0, i_13_162_3415_0, i_13_162_3416_0,
    i_13_162_3422_0, i_13_162_3530_0, i_13_162_3766_0, i_13_162_3767_0,
    i_13_162_3783_0, i_13_162_3785_0, i_13_162_3817_0, i_13_162_3818_0,
    i_13_162_3872_0, i_13_162_3924_0, i_13_162_3925_0, i_13_162_3987_0,
    i_13_162_3988_0, i_13_162_4061_0, i_13_162_4132_0, i_13_162_4280_0,
    i_13_162_4339_0, i_13_162_4342_0, i_13_162_4351_0, i_13_162_4352_0,
    i_13_162_4379_0, i_13_162_4567_0, i_13_162_4568_0, i_13_162_4591_0;
  output o_13_162_0_0;
  assign o_13_162_0_0 = ~((~i_13_162_4352_0 & ~i_13_162_4568_0) | (i_13_162_617_0 & ~i_13_162_3422_0) | (~i_13_162_92_0 & ~i_13_162_3242_0 & ~i_13_162_4280_0));
endmodule



// Benchmark "kernel_13_163" written by ABC on Sun Jul 19 10:47:42 2020

module kernel_13_163 ( 
    i_13_163_48_0, i_13_163_69_0, i_13_163_71_0, i_13_163_79_0,
    i_13_163_176_0, i_13_163_181_0, i_13_163_258_0, i_13_163_411_0,
    i_13_163_452_0, i_13_163_535_0, i_13_163_609_0, i_13_163_628_0,
    i_13_163_642_0, i_13_163_650_0, i_13_163_660_0, i_13_163_663_0,
    i_13_163_682_0, i_13_163_690_0, i_13_163_745_0, i_13_163_760_0,
    i_13_163_762_0, i_13_163_812_0, i_13_163_850_0, i_13_163_979_0,
    i_13_163_1067_0, i_13_163_1119_0, i_13_163_1121_0, i_13_163_1122_0,
    i_13_163_1132_0, i_13_163_1136_0, i_13_163_1149_0, i_13_163_1271_0,
    i_13_163_1275_0, i_13_163_1276_0, i_13_163_1311_0, i_13_163_1316_0,
    i_13_163_1402_0, i_13_163_1506_0, i_13_163_1510_0, i_13_163_1514_0,
    i_13_163_1516_0, i_13_163_1551_0, i_13_163_1563_0, i_13_163_1572_0,
    i_13_163_1596_0, i_13_163_1597_0, i_13_163_1676_0, i_13_163_1714_0,
    i_13_163_1797_0, i_13_163_1798_0, i_13_163_1807_0, i_13_163_2028_0,
    i_13_163_2057_0, i_13_163_2194_0, i_13_163_2199_0, i_13_163_2425_0,
    i_13_163_2454_0, i_13_163_2676_0, i_13_163_2678_0, i_13_163_2679_0,
    i_13_163_2697_0, i_13_163_2724_0, i_13_163_2742_0, i_13_163_2940_0,
    i_13_163_2953_0, i_13_163_2967_0, i_13_163_2976_0, i_13_163_3094_0,
    i_13_163_3118_0, i_13_163_3209_0, i_13_163_3264_0, i_13_163_3273_0,
    i_13_163_3354_0, i_13_163_3368_0, i_13_163_3399_0, i_13_163_3459_0,
    i_13_163_3487_0, i_13_163_3549_0, i_13_163_3651_0, i_13_163_3652_0,
    i_13_163_3697_0, i_13_163_3759_0, i_13_163_3764_0, i_13_163_3822_0,
    i_13_163_3864_0, i_13_163_3930_0, i_13_163_3939_0, i_13_163_4018_0,
    i_13_163_4037_0, i_13_163_4082_0, i_13_163_4255_0, i_13_163_4272_0,
    i_13_163_4300_0, i_13_163_4306_0, i_13_163_4335_0, i_13_163_4377_0,
    i_13_163_4447_0, i_13_163_4515_0, i_13_163_4565_0, i_13_163_4606_0,
    o_13_163_0_0  );
  input  i_13_163_48_0, i_13_163_69_0, i_13_163_71_0, i_13_163_79_0,
    i_13_163_176_0, i_13_163_181_0, i_13_163_258_0, i_13_163_411_0,
    i_13_163_452_0, i_13_163_535_0, i_13_163_609_0, i_13_163_628_0,
    i_13_163_642_0, i_13_163_650_0, i_13_163_660_0, i_13_163_663_0,
    i_13_163_682_0, i_13_163_690_0, i_13_163_745_0, i_13_163_760_0,
    i_13_163_762_0, i_13_163_812_0, i_13_163_850_0, i_13_163_979_0,
    i_13_163_1067_0, i_13_163_1119_0, i_13_163_1121_0, i_13_163_1122_0,
    i_13_163_1132_0, i_13_163_1136_0, i_13_163_1149_0, i_13_163_1271_0,
    i_13_163_1275_0, i_13_163_1276_0, i_13_163_1311_0, i_13_163_1316_0,
    i_13_163_1402_0, i_13_163_1506_0, i_13_163_1510_0, i_13_163_1514_0,
    i_13_163_1516_0, i_13_163_1551_0, i_13_163_1563_0, i_13_163_1572_0,
    i_13_163_1596_0, i_13_163_1597_0, i_13_163_1676_0, i_13_163_1714_0,
    i_13_163_1797_0, i_13_163_1798_0, i_13_163_1807_0, i_13_163_2028_0,
    i_13_163_2057_0, i_13_163_2194_0, i_13_163_2199_0, i_13_163_2425_0,
    i_13_163_2454_0, i_13_163_2676_0, i_13_163_2678_0, i_13_163_2679_0,
    i_13_163_2697_0, i_13_163_2724_0, i_13_163_2742_0, i_13_163_2940_0,
    i_13_163_2953_0, i_13_163_2967_0, i_13_163_2976_0, i_13_163_3094_0,
    i_13_163_3118_0, i_13_163_3209_0, i_13_163_3264_0, i_13_163_3273_0,
    i_13_163_3354_0, i_13_163_3368_0, i_13_163_3399_0, i_13_163_3459_0,
    i_13_163_3487_0, i_13_163_3549_0, i_13_163_3651_0, i_13_163_3652_0,
    i_13_163_3697_0, i_13_163_3759_0, i_13_163_3764_0, i_13_163_3822_0,
    i_13_163_3864_0, i_13_163_3930_0, i_13_163_3939_0, i_13_163_4018_0,
    i_13_163_4037_0, i_13_163_4082_0, i_13_163_4255_0, i_13_163_4272_0,
    i_13_163_4300_0, i_13_163_4306_0, i_13_163_4335_0, i_13_163_4377_0,
    i_13_163_4447_0, i_13_163_4515_0, i_13_163_4565_0, i_13_163_4606_0;
  output o_13_163_0_0;
  assign o_13_163_0_0 = ~(~i_13_163_4515_0 | ~i_13_163_1122_0 | i_13_163_4306_0);
endmodule



// Benchmark "kernel_13_164" written by ABC on Sun Jul 19 10:47:42 2020

module kernel_13_164 ( 
    i_13_164_3_0, i_13_164_40_0, i_13_164_62_0, i_13_164_94_0,
    i_13_164_112_0, i_13_164_115_0, i_13_164_127_0, i_13_164_184_0,
    i_13_164_187_0, i_13_164_207_0, i_13_164_225_0, i_13_164_234_0,
    i_13_164_244_0, i_13_164_266_0, i_13_164_268_0, i_13_164_333_0,
    i_13_164_538_0, i_13_164_607_0, i_13_164_670_0, i_13_164_769_0,
    i_13_164_814_0, i_13_164_1084_0, i_13_164_1191_0, i_13_164_1205_0,
    i_13_164_1219_0, i_13_164_1274_0, i_13_164_1321_0, i_13_164_1482_0,
    i_13_164_1489_0, i_13_164_1538_0, i_13_164_1680_0, i_13_164_1749_0,
    i_13_164_1750_0, i_13_164_1752_0, i_13_164_1804_0, i_13_164_1807_0,
    i_13_164_1840_0, i_13_164_1843_0, i_13_164_1845_0, i_13_164_1995_0,
    i_13_164_1996_0, i_13_164_2128_0, i_13_164_2138_0, i_13_164_2140_0,
    i_13_164_2142_0, i_13_164_2173_0, i_13_164_2176_0, i_13_164_2304_0,
    i_13_164_2407_0, i_13_164_2409_0, i_13_164_2425_0, i_13_164_2434_0,
    i_13_164_2446_0, i_13_164_2494_0, i_13_164_2506_0, i_13_164_2576_0,
    i_13_164_2581_0, i_13_164_2694_0, i_13_164_2742_0, i_13_164_2745_0,
    i_13_164_2749_0, i_13_164_2940_0, i_13_164_2965_0, i_13_164_3030_0,
    i_13_164_3031_0, i_13_164_3100_0, i_13_164_3120_0, i_13_164_3123_0,
    i_13_164_3135_0, i_13_164_3145_0, i_13_164_3148_0, i_13_164_3163_0,
    i_13_164_3273_0, i_13_164_3343_0, i_13_164_3373_0, i_13_164_3402_0,
    i_13_164_3418_0, i_13_164_3504_0, i_13_164_3505_0, i_13_164_3537_0,
    i_13_164_3569_0, i_13_164_3637_0, i_13_164_3669_0, i_13_164_3739_0,
    i_13_164_3746_0, i_13_164_3874_0, i_13_164_3878_0, i_13_164_3892_0,
    i_13_164_3909_0, i_13_164_3912_0, i_13_164_3991_0, i_13_164_4104_0,
    i_13_164_4120_0, i_13_164_4341_0, i_13_164_4354_0, i_13_164_4378_0,
    i_13_164_4380_0, i_13_164_4390_0, i_13_164_4461_0, i_13_164_4583_0,
    o_13_164_0_0  );
  input  i_13_164_3_0, i_13_164_40_0, i_13_164_62_0, i_13_164_94_0,
    i_13_164_112_0, i_13_164_115_0, i_13_164_127_0, i_13_164_184_0,
    i_13_164_187_0, i_13_164_207_0, i_13_164_225_0, i_13_164_234_0,
    i_13_164_244_0, i_13_164_266_0, i_13_164_268_0, i_13_164_333_0,
    i_13_164_538_0, i_13_164_607_0, i_13_164_670_0, i_13_164_769_0,
    i_13_164_814_0, i_13_164_1084_0, i_13_164_1191_0, i_13_164_1205_0,
    i_13_164_1219_0, i_13_164_1274_0, i_13_164_1321_0, i_13_164_1482_0,
    i_13_164_1489_0, i_13_164_1538_0, i_13_164_1680_0, i_13_164_1749_0,
    i_13_164_1750_0, i_13_164_1752_0, i_13_164_1804_0, i_13_164_1807_0,
    i_13_164_1840_0, i_13_164_1843_0, i_13_164_1845_0, i_13_164_1995_0,
    i_13_164_1996_0, i_13_164_2128_0, i_13_164_2138_0, i_13_164_2140_0,
    i_13_164_2142_0, i_13_164_2173_0, i_13_164_2176_0, i_13_164_2304_0,
    i_13_164_2407_0, i_13_164_2409_0, i_13_164_2425_0, i_13_164_2434_0,
    i_13_164_2446_0, i_13_164_2494_0, i_13_164_2506_0, i_13_164_2576_0,
    i_13_164_2581_0, i_13_164_2694_0, i_13_164_2742_0, i_13_164_2745_0,
    i_13_164_2749_0, i_13_164_2940_0, i_13_164_2965_0, i_13_164_3030_0,
    i_13_164_3031_0, i_13_164_3100_0, i_13_164_3120_0, i_13_164_3123_0,
    i_13_164_3135_0, i_13_164_3145_0, i_13_164_3148_0, i_13_164_3163_0,
    i_13_164_3273_0, i_13_164_3343_0, i_13_164_3373_0, i_13_164_3402_0,
    i_13_164_3418_0, i_13_164_3504_0, i_13_164_3505_0, i_13_164_3537_0,
    i_13_164_3569_0, i_13_164_3637_0, i_13_164_3669_0, i_13_164_3739_0,
    i_13_164_3746_0, i_13_164_3874_0, i_13_164_3878_0, i_13_164_3892_0,
    i_13_164_3909_0, i_13_164_3912_0, i_13_164_3991_0, i_13_164_4104_0,
    i_13_164_4120_0, i_13_164_4341_0, i_13_164_4354_0, i_13_164_4378_0,
    i_13_164_4380_0, i_13_164_4390_0, i_13_164_4461_0, i_13_164_4583_0;
  output o_13_164_0_0;
  assign o_13_164_0_0 = ~((~i_13_164_1749_0 & ((i_13_164_2173_0 & i_13_164_2434_0 & ~i_13_164_2446_0) | (~i_13_164_1807_0 & i_13_164_3505_0))) | (~i_13_164_1845_0 & ((~i_13_164_184_0 & ~i_13_164_2140_0 & ~i_13_164_2407_0) | (~i_13_164_1996_0 & ~i_13_164_3991_0 & ~i_13_164_4378_0))) | (~i_13_164_2694_0 & ((i_13_164_94_0 & i_13_164_3739_0) | (~i_13_164_1321_0 & ~i_13_164_2940_0 & ~i_13_164_3537_0 & ~i_13_164_3746_0 & ~i_13_164_4354_0))) | i_13_164_112_0 | (~i_13_164_1750_0 & i_13_164_3505_0 & i_13_164_3537_0) | (~i_13_164_1804_0 & ~i_13_164_2140_0 & i_13_164_3991_0));
endmodule



// Benchmark "kernel_13_165" written by ABC on Sun Jul 19 10:47:43 2020

module kernel_13_165 ( 
    i_13_165_51_0, i_13_165_76_0, i_13_165_96_0, i_13_165_129_0,
    i_13_165_157_0, i_13_165_159_0, i_13_165_164_0, i_13_165_167_0,
    i_13_165_169_0, i_13_165_170_0, i_13_165_266_0, i_13_165_282_0,
    i_13_165_375_0, i_13_165_377_0, i_13_165_384_0, i_13_165_568_0,
    i_13_165_598_0, i_13_165_683_0, i_13_165_697_0, i_13_165_714_0,
    i_13_165_814_0, i_13_165_816_0, i_13_165_817_0, i_13_165_844_0,
    i_13_165_858_0, i_13_165_984_0, i_13_165_1068_0, i_13_165_1106_0,
    i_13_165_1301_0, i_13_165_1511_0, i_13_165_1570_0, i_13_165_1749_0,
    i_13_165_1777_0, i_13_165_1795_0, i_13_165_1807_0, i_13_165_1829_0,
    i_13_165_1851_0, i_13_165_1852_0, i_13_165_1857_0, i_13_165_1912_0,
    i_13_165_1924_0, i_13_165_2108_0, i_13_165_2110_0, i_13_165_2122_0,
    i_13_165_2139_0, i_13_165_2208_0, i_13_165_2241_0, i_13_165_2264_0,
    i_13_165_2266_0, i_13_165_2407_0, i_13_165_2425_0, i_13_165_2437_0,
    i_13_165_2497_0, i_13_165_2554_0, i_13_165_2567_0, i_13_165_2570_0,
    i_13_165_2679_0, i_13_165_2698_0, i_13_165_2797_0, i_13_165_2848_0,
    i_13_165_2884_0, i_13_165_2921_0, i_13_165_2940_0, i_13_165_2941_0,
    i_13_165_2983_0, i_13_165_3030_0, i_13_165_3031_0, i_13_165_3038_0,
    i_13_165_3110_0, i_13_165_3116_0, i_13_165_3147_0, i_13_165_3208_0,
    i_13_165_3210_0, i_13_165_3212_0, i_13_165_3239_0, i_13_165_3327_0,
    i_13_165_3345_0, i_13_165_3400_0, i_13_165_3408_0, i_13_165_3505_0,
    i_13_165_3732_0, i_13_165_3739_0, i_13_165_3741_0, i_13_165_3767_0,
    i_13_165_3820_0, i_13_165_3941_0, i_13_165_3994_0, i_13_165_4045_0,
    i_13_165_4048_0, i_13_165_4061_0, i_13_165_4063_0, i_13_165_4064_0,
    i_13_165_4066_0, i_13_165_4080_0, i_13_165_4119_0, i_13_165_4309_0,
    i_13_165_4318_0, i_13_165_4333_0, i_13_165_4397_0, i_13_165_4607_0,
    o_13_165_0_0  );
  input  i_13_165_51_0, i_13_165_76_0, i_13_165_96_0, i_13_165_129_0,
    i_13_165_157_0, i_13_165_159_0, i_13_165_164_0, i_13_165_167_0,
    i_13_165_169_0, i_13_165_170_0, i_13_165_266_0, i_13_165_282_0,
    i_13_165_375_0, i_13_165_377_0, i_13_165_384_0, i_13_165_568_0,
    i_13_165_598_0, i_13_165_683_0, i_13_165_697_0, i_13_165_714_0,
    i_13_165_814_0, i_13_165_816_0, i_13_165_817_0, i_13_165_844_0,
    i_13_165_858_0, i_13_165_984_0, i_13_165_1068_0, i_13_165_1106_0,
    i_13_165_1301_0, i_13_165_1511_0, i_13_165_1570_0, i_13_165_1749_0,
    i_13_165_1777_0, i_13_165_1795_0, i_13_165_1807_0, i_13_165_1829_0,
    i_13_165_1851_0, i_13_165_1852_0, i_13_165_1857_0, i_13_165_1912_0,
    i_13_165_1924_0, i_13_165_2108_0, i_13_165_2110_0, i_13_165_2122_0,
    i_13_165_2139_0, i_13_165_2208_0, i_13_165_2241_0, i_13_165_2264_0,
    i_13_165_2266_0, i_13_165_2407_0, i_13_165_2425_0, i_13_165_2437_0,
    i_13_165_2497_0, i_13_165_2554_0, i_13_165_2567_0, i_13_165_2570_0,
    i_13_165_2679_0, i_13_165_2698_0, i_13_165_2797_0, i_13_165_2848_0,
    i_13_165_2884_0, i_13_165_2921_0, i_13_165_2940_0, i_13_165_2941_0,
    i_13_165_2983_0, i_13_165_3030_0, i_13_165_3031_0, i_13_165_3038_0,
    i_13_165_3110_0, i_13_165_3116_0, i_13_165_3147_0, i_13_165_3208_0,
    i_13_165_3210_0, i_13_165_3212_0, i_13_165_3239_0, i_13_165_3327_0,
    i_13_165_3345_0, i_13_165_3400_0, i_13_165_3408_0, i_13_165_3505_0,
    i_13_165_3732_0, i_13_165_3739_0, i_13_165_3741_0, i_13_165_3767_0,
    i_13_165_3820_0, i_13_165_3941_0, i_13_165_3994_0, i_13_165_4045_0,
    i_13_165_4048_0, i_13_165_4061_0, i_13_165_4063_0, i_13_165_4064_0,
    i_13_165_4066_0, i_13_165_4080_0, i_13_165_4119_0, i_13_165_4309_0,
    i_13_165_4318_0, i_13_165_4333_0, i_13_165_4397_0, i_13_165_4607_0;
  output o_13_165_0_0;
  assign o_13_165_0_0 = ~((~i_13_165_1301_0 & ((~i_13_165_1807_0 & ~i_13_165_1851_0 & i_13_165_3505_0 & ~i_13_165_4064_0 & ~i_13_165_4066_0) | (~i_13_165_2983_0 & ~i_13_165_4309_0 & ~i_13_165_4318_0))) | (~i_13_165_2407_0 & ((i_13_165_2884_0 & i_13_165_2921_0 & i_13_165_3505_0) | (~i_13_165_1511_0 & ~i_13_165_1852_0 & ~i_13_165_2139_0 & ~i_13_165_2698_0 & ~i_13_165_4061_0 & ~i_13_165_4066_0))) | (~i_13_165_2921_0 & i_13_165_4061_0 & (~i_13_165_4064_0 | (~i_13_165_2110_0 & ~i_13_165_4063_0))) | (~i_13_165_2208_0 & ~i_13_165_3110_0 & i_13_165_3505_0 & ~i_13_165_3767_0) | (i_13_165_697_0 & ~i_13_165_4080_0));
endmodule



// Benchmark "kernel_13_166" written by ABC on Sun Jul 19 10:47:44 2020

module kernel_13_166 ( 
    i_13_166_235_0, i_13_166_238_0, i_13_166_414_0, i_13_166_415_0,
    i_13_166_416_0, i_13_166_432_0, i_13_166_446_0, i_13_166_507_0,
    i_13_166_523_0, i_13_166_526_0, i_13_166_535_0, i_13_166_562_0,
    i_13_166_568_0, i_13_166_694_0, i_13_166_797_0, i_13_166_823_0,
    i_13_166_841_0, i_13_166_842_0, i_13_166_946_0, i_13_166_1018_0,
    i_13_166_1073_0, i_13_166_1076_0, i_13_166_1129_0, i_13_166_1132_0,
    i_13_166_1190_0, i_13_166_1193_0, i_13_166_1214_0, i_13_166_1228_0,
    i_13_166_1252_0, i_13_166_1256_0, i_13_166_1268_0, i_13_166_1400_0,
    i_13_166_1411_0, i_13_166_1531_0, i_13_166_1548_0, i_13_166_1549_0,
    i_13_166_1550_0, i_13_166_1552_0, i_13_166_1553_0, i_13_166_1603_0,
    i_13_166_1696_0, i_13_166_1846_0, i_13_166_1934_0, i_13_166_1957_0,
    i_13_166_1958_0, i_13_166_2043_0, i_13_166_2109_0, i_13_166_2203_0,
    i_13_166_2289_0, i_13_166_2334_0, i_13_166_2380_0, i_13_166_2449_0,
    i_13_166_2539_0, i_13_166_2555_0, i_13_166_2611_0, i_13_166_2713_0,
    i_13_166_2754_0, i_13_166_2900_0, i_13_166_3010_0, i_13_166_3013_0,
    i_13_166_3014_0, i_13_166_3064_0, i_13_166_3065_0, i_13_166_3070_0,
    i_13_166_3101_0, i_13_166_3172_0, i_13_166_3272_0, i_13_166_3382_0,
    i_13_166_3416_0, i_13_166_3451_0, i_13_166_3461_0, i_13_166_3484_0,
    i_13_166_3487_0, i_13_166_3488_0, i_13_166_3523_0, i_13_166_3537_0,
    i_13_166_3538_0, i_13_166_3539_0, i_13_166_3541_0, i_13_166_3542_0,
    i_13_166_3544_0, i_13_166_3545_0, i_13_166_3686_0, i_13_166_3730_0,
    i_13_166_3766_0, i_13_166_3852_0, i_13_166_3856_0, i_13_166_3857_0,
    i_13_166_3880_0, i_13_166_3895_0, i_13_166_3908_0, i_13_166_3915_0,
    i_13_166_3916_0, i_13_166_4252_0, i_13_166_4256_0, i_13_166_4369_0,
    i_13_166_4378_0, i_13_166_4379_0, i_13_166_4382_0, i_13_166_4536_0,
    o_13_166_0_0  );
  input  i_13_166_235_0, i_13_166_238_0, i_13_166_414_0, i_13_166_415_0,
    i_13_166_416_0, i_13_166_432_0, i_13_166_446_0, i_13_166_507_0,
    i_13_166_523_0, i_13_166_526_0, i_13_166_535_0, i_13_166_562_0,
    i_13_166_568_0, i_13_166_694_0, i_13_166_797_0, i_13_166_823_0,
    i_13_166_841_0, i_13_166_842_0, i_13_166_946_0, i_13_166_1018_0,
    i_13_166_1073_0, i_13_166_1076_0, i_13_166_1129_0, i_13_166_1132_0,
    i_13_166_1190_0, i_13_166_1193_0, i_13_166_1214_0, i_13_166_1228_0,
    i_13_166_1252_0, i_13_166_1256_0, i_13_166_1268_0, i_13_166_1400_0,
    i_13_166_1411_0, i_13_166_1531_0, i_13_166_1548_0, i_13_166_1549_0,
    i_13_166_1550_0, i_13_166_1552_0, i_13_166_1553_0, i_13_166_1603_0,
    i_13_166_1696_0, i_13_166_1846_0, i_13_166_1934_0, i_13_166_1957_0,
    i_13_166_1958_0, i_13_166_2043_0, i_13_166_2109_0, i_13_166_2203_0,
    i_13_166_2289_0, i_13_166_2334_0, i_13_166_2380_0, i_13_166_2449_0,
    i_13_166_2539_0, i_13_166_2555_0, i_13_166_2611_0, i_13_166_2713_0,
    i_13_166_2754_0, i_13_166_2900_0, i_13_166_3010_0, i_13_166_3013_0,
    i_13_166_3014_0, i_13_166_3064_0, i_13_166_3065_0, i_13_166_3070_0,
    i_13_166_3101_0, i_13_166_3172_0, i_13_166_3272_0, i_13_166_3382_0,
    i_13_166_3416_0, i_13_166_3451_0, i_13_166_3461_0, i_13_166_3484_0,
    i_13_166_3487_0, i_13_166_3488_0, i_13_166_3523_0, i_13_166_3537_0,
    i_13_166_3538_0, i_13_166_3539_0, i_13_166_3541_0, i_13_166_3542_0,
    i_13_166_3544_0, i_13_166_3545_0, i_13_166_3686_0, i_13_166_3730_0,
    i_13_166_3766_0, i_13_166_3852_0, i_13_166_3856_0, i_13_166_3857_0,
    i_13_166_3880_0, i_13_166_3895_0, i_13_166_3908_0, i_13_166_3915_0,
    i_13_166_3916_0, i_13_166_4252_0, i_13_166_4256_0, i_13_166_4369_0,
    i_13_166_4378_0, i_13_166_4379_0, i_13_166_4382_0, i_13_166_4536_0;
  output o_13_166_0_0;
  assign o_13_166_0_0 = ~((~i_13_166_3010_0 & ((~i_13_166_694_0 & i_13_166_3857_0) | (~i_13_166_3539_0 & ~i_13_166_4379_0))) | (i_13_166_841_0 & ~i_13_166_1018_0) | (~i_13_166_415_0 & ~i_13_166_1252_0 & ~i_13_166_1256_0) | (~i_13_166_1549_0 & ~i_13_166_1603_0 & ~i_13_166_3539_0 & ~i_13_166_3541_0));
endmodule



// Benchmark "kernel_13_167" written by ABC on Sun Jul 19 10:47:45 2020

module kernel_13_167 ( 
    i_13_167_80_0, i_13_167_139_0, i_13_167_232_0, i_13_167_283_0,
    i_13_167_332_0, i_13_167_358_0, i_13_167_376_0, i_13_167_428_0,
    i_13_167_447_0, i_13_167_457_0, i_13_167_538_0, i_13_167_599_0,
    i_13_167_607_0, i_13_167_646_0, i_13_167_647_0, i_13_167_688_0,
    i_13_167_689_0, i_13_167_691_0, i_13_167_692_0, i_13_167_718_0,
    i_13_167_728_0, i_13_167_940_0, i_13_167_979_0, i_13_167_1120_0,
    i_13_167_1204_0, i_13_167_1263_0, i_13_167_1275_0, i_13_167_1276_0,
    i_13_167_1277_0, i_13_167_1348_0, i_13_167_1393_0, i_13_167_1484_0,
    i_13_167_1493_0, i_13_167_1570_0, i_13_167_1642_0, i_13_167_1645_0,
    i_13_167_1646_0, i_13_167_1672_0, i_13_167_1673_0, i_13_167_1691_0,
    i_13_167_1713_0, i_13_167_1723_0, i_13_167_1726_0, i_13_167_1727_0,
    i_13_167_1741_0, i_13_167_1780_0, i_13_167_1781_0, i_13_167_1885_0,
    i_13_167_1888_0, i_13_167_1933_0, i_13_167_1996_0, i_13_167_2113_0,
    i_13_167_2137_0, i_13_167_2150_0, i_13_167_2191_0, i_13_167_2194_0,
    i_13_167_2282_0, i_13_167_2379_0, i_13_167_2383_0, i_13_167_2533_0,
    i_13_167_2542_0, i_13_167_2552_0, i_13_167_2617_0, i_13_167_2649_0,
    i_13_167_2650_0, i_13_167_2651_0, i_13_167_2653_0, i_13_167_2654_0,
    i_13_167_2661_0, i_13_167_2671_0, i_13_167_2690_0, i_13_167_2742_0,
    i_13_167_2751_0, i_13_167_2847_0, i_13_167_2848_0, i_13_167_2851_0,
    i_13_167_2852_0, i_13_167_2875_0, i_13_167_2878_0, i_13_167_3139_0,
    i_13_167_3392_0, i_13_167_3535_0, i_13_167_3581_0, i_13_167_3760_0,
    i_13_167_3797_0, i_13_167_3874_0, i_13_167_3995_0, i_13_167_4045_0,
    i_13_167_4162_0, i_13_167_4190_0, i_13_167_4193_0, i_13_167_4219_0,
    i_13_167_4234_0, i_13_167_4354_0, i_13_167_4377_0, i_13_167_4423_0,
    i_13_167_4432_0, i_13_167_4444_0, i_13_167_4597_0, i_13_167_4598_0,
    o_13_167_0_0  );
  input  i_13_167_80_0, i_13_167_139_0, i_13_167_232_0, i_13_167_283_0,
    i_13_167_332_0, i_13_167_358_0, i_13_167_376_0, i_13_167_428_0,
    i_13_167_447_0, i_13_167_457_0, i_13_167_538_0, i_13_167_599_0,
    i_13_167_607_0, i_13_167_646_0, i_13_167_647_0, i_13_167_688_0,
    i_13_167_689_0, i_13_167_691_0, i_13_167_692_0, i_13_167_718_0,
    i_13_167_728_0, i_13_167_940_0, i_13_167_979_0, i_13_167_1120_0,
    i_13_167_1204_0, i_13_167_1263_0, i_13_167_1275_0, i_13_167_1276_0,
    i_13_167_1277_0, i_13_167_1348_0, i_13_167_1393_0, i_13_167_1484_0,
    i_13_167_1493_0, i_13_167_1570_0, i_13_167_1642_0, i_13_167_1645_0,
    i_13_167_1646_0, i_13_167_1672_0, i_13_167_1673_0, i_13_167_1691_0,
    i_13_167_1713_0, i_13_167_1723_0, i_13_167_1726_0, i_13_167_1727_0,
    i_13_167_1741_0, i_13_167_1780_0, i_13_167_1781_0, i_13_167_1885_0,
    i_13_167_1888_0, i_13_167_1933_0, i_13_167_1996_0, i_13_167_2113_0,
    i_13_167_2137_0, i_13_167_2150_0, i_13_167_2191_0, i_13_167_2194_0,
    i_13_167_2282_0, i_13_167_2379_0, i_13_167_2383_0, i_13_167_2533_0,
    i_13_167_2542_0, i_13_167_2552_0, i_13_167_2617_0, i_13_167_2649_0,
    i_13_167_2650_0, i_13_167_2651_0, i_13_167_2653_0, i_13_167_2654_0,
    i_13_167_2661_0, i_13_167_2671_0, i_13_167_2690_0, i_13_167_2742_0,
    i_13_167_2751_0, i_13_167_2847_0, i_13_167_2848_0, i_13_167_2851_0,
    i_13_167_2852_0, i_13_167_2875_0, i_13_167_2878_0, i_13_167_3139_0,
    i_13_167_3392_0, i_13_167_3535_0, i_13_167_3581_0, i_13_167_3760_0,
    i_13_167_3797_0, i_13_167_3874_0, i_13_167_3995_0, i_13_167_4045_0,
    i_13_167_4162_0, i_13_167_4190_0, i_13_167_4193_0, i_13_167_4219_0,
    i_13_167_4234_0, i_13_167_4354_0, i_13_167_4377_0, i_13_167_4423_0,
    i_13_167_4432_0, i_13_167_4444_0, i_13_167_4597_0, i_13_167_4598_0;
  output o_13_167_0_0;
  assign o_13_167_0_0 = ~(~i_13_167_2878_0 | (~i_13_167_1277_0 & ~i_13_167_2851_0) | (~i_13_167_283_0 & ~i_13_167_2651_0));
endmodule



// Benchmark "kernel_13_168" written by ABC on Sun Jul 19 10:47:46 2020

module kernel_13_168 ( 
    i_13_168_52_0, i_13_168_116_0, i_13_168_167_0, i_13_168_185_0,
    i_13_168_199_0, i_13_168_251_0, i_13_168_286_0, i_13_168_287_0,
    i_13_168_418_0, i_13_168_441_0, i_13_168_517_0, i_13_168_556_0,
    i_13_168_559_0, i_13_168_576_0, i_13_168_619_0, i_13_168_620_0,
    i_13_168_655_0, i_13_168_675_0, i_13_168_715_0, i_13_168_928_0,
    i_13_168_929_0, i_13_168_944_0, i_13_168_1018_0, i_13_168_1085_0,
    i_13_168_1098_0, i_13_168_1310_0, i_13_168_1364_0, i_13_168_1397_0,
    i_13_168_1426_0, i_13_168_1471_0, i_13_168_1498_0, i_13_168_1501_0,
    i_13_168_1502_0, i_13_168_1505_0, i_13_168_1606_0, i_13_168_1609_0,
    i_13_168_1633_0, i_13_168_1634_0, i_13_168_1636_0, i_13_168_1637_0,
    i_13_168_1731_0, i_13_168_1735_0, i_13_168_1754_0, i_13_168_1917_0,
    i_13_168_1949_0, i_13_168_2171_0, i_13_168_2276_0, i_13_168_2342_0,
    i_13_168_2369_0, i_13_168_2455_0, i_13_168_2492_0, i_13_168_2545_0,
    i_13_168_2581_0, i_13_168_2673_0, i_13_168_2708_0, i_13_168_2714_0,
    i_13_168_2753_0, i_13_168_2788_0, i_13_168_2888_0, i_13_168_2922_0,
    i_13_168_2923_0, i_13_168_2956_0, i_13_168_2959_0, i_13_168_3130_0,
    i_13_168_3145_0, i_13_168_3146_0, i_13_168_3149_0, i_13_168_3253_0,
    i_13_168_3373_0, i_13_168_3409_0, i_13_168_3418_0, i_13_168_3419_0,
    i_13_168_3447_0, i_13_168_3464_0, i_13_168_3486_0, i_13_168_3581_0,
    i_13_168_3599_0, i_13_168_3647_0, i_13_168_3650_0, i_13_168_3724_0,
    i_13_168_3734_0, i_13_168_3765_0, i_13_168_3770_0, i_13_168_3787_0,
    i_13_168_3816_0, i_13_168_3904_0, i_13_168_3905_0, i_13_168_4015_0,
    i_13_168_4019_0, i_13_168_4077_0, i_13_168_4087_0, i_13_168_4088_0,
    i_13_168_4253_0, i_13_168_4255_0, i_13_168_4256_0, i_13_168_4391_0,
    i_13_168_4531_0, i_13_168_4562_0, i_13_168_4567_0, i_13_168_4590_0,
    o_13_168_0_0  );
  input  i_13_168_52_0, i_13_168_116_0, i_13_168_167_0, i_13_168_185_0,
    i_13_168_199_0, i_13_168_251_0, i_13_168_286_0, i_13_168_287_0,
    i_13_168_418_0, i_13_168_441_0, i_13_168_517_0, i_13_168_556_0,
    i_13_168_559_0, i_13_168_576_0, i_13_168_619_0, i_13_168_620_0,
    i_13_168_655_0, i_13_168_675_0, i_13_168_715_0, i_13_168_928_0,
    i_13_168_929_0, i_13_168_944_0, i_13_168_1018_0, i_13_168_1085_0,
    i_13_168_1098_0, i_13_168_1310_0, i_13_168_1364_0, i_13_168_1397_0,
    i_13_168_1426_0, i_13_168_1471_0, i_13_168_1498_0, i_13_168_1501_0,
    i_13_168_1502_0, i_13_168_1505_0, i_13_168_1606_0, i_13_168_1609_0,
    i_13_168_1633_0, i_13_168_1634_0, i_13_168_1636_0, i_13_168_1637_0,
    i_13_168_1731_0, i_13_168_1735_0, i_13_168_1754_0, i_13_168_1917_0,
    i_13_168_1949_0, i_13_168_2171_0, i_13_168_2276_0, i_13_168_2342_0,
    i_13_168_2369_0, i_13_168_2455_0, i_13_168_2492_0, i_13_168_2545_0,
    i_13_168_2581_0, i_13_168_2673_0, i_13_168_2708_0, i_13_168_2714_0,
    i_13_168_2753_0, i_13_168_2788_0, i_13_168_2888_0, i_13_168_2922_0,
    i_13_168_2923_0, i_13_168_2956_0, i_13_168_2959_0, i_13_168_3130_0,
    i_13_168_3145_0, i_13_168_3146_0, i_13_168_3149_0, i_13_168_3253_0,
    i_13_168_3373_0, i_13_168_3409_0, i_13_168_3418_0, i_13_168_3419_0,
    i_13_168_3447_0, i_13_168_3464_0, i_13_168_3486_0, i_13_168_3581_0,
    i_13_168_3599_0, i_13_168_3647_0, i_13_168_3650_0, i_13_168_3724_0,
    i_13_168_3734_0, i_13_168_3765_0, i_13_168_3770_0, i_13_168_3787_0,
    i_13_168_3816_0, i_13_168_3904_0, i_13_168_3905_0, i_13_168_4015_0,
    i_13_168_4019_0, i_13_168_4077_0, i_13_168_4087_0, i_13_168_4088_0,
    i_13_168_4253_0, i_13_168_4255_0, i_13_168_4256_0, i_13_168_4391_0,
    i_13_168_4531_0, i_13_168_4562_0, i_13_168_4567_0, i_13_168_4590_0;
  output o_13_168_0_0;
  assign o_13_168_0_0 = ~(~i_13_168_3770_0 | (~i_13_168_2923_0 & ~i_13_168_4562_0) | (~i_13_168_1502_0 & ~i_13_168_4253_0) | (~i_13_168_3145_0 & i_13_168_3146_0));
endmodule



// Benchmark "kernel_13_169" written by ABC on Sun Jul 19 10:47:47 2020

module kernel_13_169 ( 
    i_13_169_112_0, i_13_169_136_0, i_13_169_158_0, i_13_169_163_0,
    i_13_169_226_0, i_13_169_229_0, i_13_169_336_0, i_13_169_380_0,
    i_13_169_382_0, i_13_169_418_0, i_13_169_445_0, i_13_169_453_0,
    i_13_169_517_0, i_13_169_569_0, i_13_169_571_0, i_13_169_577_0,
    i_13_169_596_0, i_13_169_614_0, i_13_169_641_0, i_13_169_652_0,
    i_13_169_686_0, i_13_169_715_0, i_13_169_733_0, i_13_169_778_0,
    i_13_169_779_0, i_13_169_841_0, i_13_169_873_0, i_13_169_1101_0,
    i_13_169_1300_0, i_13_169_1327_0, i_13_169_1444_0, i_13_169_1462_0,
    i_13_169_1503_0, i_13_169_1517_0, i_13_169_1521_0, i_13_169_1625_0,
    i_13_169_1711_0, i_13_169_1713_0, i_13_169_1720_0, i_13_169_1721_0,
    i_13_169_1730_0, i_13_169_1783_0, i_13_169_1786_0, i_13_169_1787_0,
    i_13_169_1802_0, i_13_169_1811_0, i_13_169_1882_0, i_13_169_1884_0,
    i_13_169_1999_0, i_13_169_2018_0, i_13_169_2097_0, i_13_169_2120_0,
    i_13_169_2170_0, i_13_169_2192_0, i_13_169_2210_0, i_13_169_2260_0,
    i_13_169_2425_0, i_13_169_2458_0, i_13_169_2541_0, i_13_169_2647_0,
    i_13_169_2712_0, i_13_169_2722_0, i_13_169_2845_0, i_13_169_2935_0,
    i_13_169_2939_0, i_13_169_3015_0, i_13_169_3020_0, i_13_169_3033_0,
    i_13_169_3034_0, i_13_169_3036_0, i_13_169_3037_0, i_13_169_3124_0,
    i_13_169_3142_0, i_13_169_3143_0, i_13_169_3164_0, i_13_169_3213_0,
    i_13_169_3270_0, i_13_169_3290_0, i_13_169_3421_0, i_13_169_3422_0,
    i_13_169_3424_0, i_13_169_3425_0, i_13_169_3430_0, i_13_169_3449_0,
    i_13_169_3547_0, i_13_169_3568_0, i_13_169_3791_0, i_13_169_3862_0,
    i_13_169_3865_0, i_13_169_3983_0, i_13_169_4009_0, i_13_169_4010_0,
    i_13_169_4015_0, i_13_169_4016_0, i_13_169_4054_0, i_13_169_4086_0,
    i_13_169_4234_0, i_13_169_4306_0, i_13_169_4311_0, i_13_169_4369_0,
    o_13_169_0_0  );
  input  i_13_169_112_0, i_13_169_136_0, i_13_169_158_0, i_13_169_163_0,
    i_13_169_226_0, i_13_169_229_0, i_13_169_336_0, i_13_169_380_0,
    i_13_169_382_0, i_13_169_418_0, i_13_169_445_0, i_13_169_453_0,
    i_13_169_517_0, i_13_169_569_0, i_13_169_571_0, i_13_169_577_0,
    i_13_169_596_0, i_13_169_614_0, i_13_169_641_0, i_13_169_652_0,
    i_13_169_686_0, i_13_169_715_0, i_13_169_733_0, i_13_169_778_0,
    i_13_169_779_0, i_13_169_841_0, i_13_169_873_0, i_13_169_1101_0,
    i_13_169_1300_0, i_13_169_1327_0, i_13_169_1444_0, i_13_169_1462_0,
    i_13_169_1503_0, i_13_169_1517_0, i_13_169_1521_0, i_13_169_1625_0,
    i_13_169_1711_0, i_13_169_1713_0, i_13_169_1720_0, i_13_169_1721_0,
    i_13_169_1730_0, i_13_169_1783_0, i_13_169_1786_0, i_13_169_1787_0,
    i_13_169_1802_0, i_13_169_1811_0, i_13_169_1882_0, i_13_169_1884_0,
    i_13_169_1999_0, i_13_169_2018_0, i_13_169_2097_0, i_13_169_2120_0,
    i_13_169_2170_0, i_13_169_2192_0, i_13_169_2210_0, i_13_169_2260_0,
    i_13_169_2425_0, i_13_169_2458_0, i_13_169_2541_0, i_13_169_2647_0,
    i_13_169_2712_0, i_13_169_2722_0, i_13_169_2845_0, i_13_169_2935_0,
    i_13_169_2939_0, i_13_169_3015_0, i_13_169_3020_0, i_13_169_3033_0,
    i_13_169_3034_0, i_13_169_3036_0, i_13_169_3037_0, i_13_169_3124_0,
    i_13_169_3142_0, i_13_169_3143_0, i_13_169_3164_0, i_13_169_3213_0,
    i_13_169_3270_0, i_13_169_3290_0, i_13_169_3421_0, i_13_169_3422_0,
    i_13_169_3424_0, i_13_169_3425_0, i_13_169_3430_0, i_13_169_3449_0,
    i_13_169_3547_0, i_13_169_3568_0, i_13_169_3791_0, i_13_169_3862_0,
    i_13_169_3865_0, i_13_169_3983_0, i_13_169_4009_0, i_13_169_4010_0,
    i_13_169_4015_0, i_13_169_4016_0, i_13_169_4054_0, i_13_169_4086_0,
    i_13_169_4234_0, i_13_169_4306_0, i_13_169_4311_0, i_13_169_4369_0;
  output o_13_169_0_0;
  assign o_13_169_0_0 = ~((~i_13_169_382_0 & ((i_13_169_841_0 & ~i_13_169_1711_0 & ~i_13_169_1811_0 & i_13_169_3865_0) | (~i_13_169_445_0 & ~i_13_169_2458_0 & ~i_13_169_2712_0 & i_13_169_4234_0 & ~i_13_169_4306_0))) | (~i_13_169_2210_0 & ~i_13_169_2425_0 & ((~i_13_169_226_0 & ~i_13_169_569_0 & ~i_13_169_1884_0) | (~i_13_169_380_0 & ~i_13_169_652_0 & ~i_13_169_2845_0 & ~i_13_169_3033_0 & ~i_13_169_3164_0 & ~i_13_169_3213_0 & ~i_13_169_4009_0))) | (~i_13_169_3421_0 & (i_13_169_418_0 | (~i_13_169_571_0 & ~i_13_169_2712_0 & ~i_13_169_2845_0 & ~i_13_169_3983_0))) | (~i_13_169_136_0 & ~i_13_169_1300_0 & ~i_13_169_3425_0) | (~i_13_169_1882_0 & ~i_13_169_3164_0 & ~i_13_169_3422_0 & i_13_169_3865_0) | (i_13_169_2712_0 & ~i_13_169_3547_0 & ~i_13_169_4234_0));
endmodule



// Benchmark "kernel_13_170" written by ABC on Sun Jul 19 10:47:47 2020

module kernel_13_170 ( 
    i_13_170_48_0, i_13_170_136_0, i_13_170_144_0, i_13_170_211_0,
    i_13_170_229_0, i_13_170_271_0, i_13_170_283_0, i_13_170_300_0,
    i_13_170_382_0, i_13_170_517_0, i_13_170_571_0, i_13_170_585_0,
    i_13_170_639_0, i_13_170_705_0, i_13_170_711_0, i_13_170_738_0,
    i_13_170_796_0, i_13_170_940_0, i_13_170_999_0, i_13_170_1044_0,
    i_13_170_1101_0, i_13_170_1344_0, i_13_170_1377_0, i_13_170_1390_0,
    i_13_170_1399_0, i_13_170_1408_0, i_13_170_1432_0, i_13_170_1513_0,
    i_13_170_1632_0, i_13_170_1633_0, i_13_170_1639_0, i_13_170_1768_0,
    i_13_170_1776_0, i_13_170_1795_0, i_13_170_1848_0, i_13_170_1893_0,
    i_13_170_1936_0, i_13_170_1945_0, i_13_170_2029_0, i_13_170_2030_0,
    i_13_170_2053_0, i_13_170_2250_0, i_13_170_2251_0, i_13_170_2253_0,
    i_13_170_2278_0, i_13_170_2413_0, i_13_170_2424_0, i_13_170_2433_0,
    i_13_170_2497_0, i_13_170_2515_0, i_13_170_2542_0, i_13_170_2547_0,
    i_13_170_2614_0, i_13_170_2668_0, i_13_170_2674_0, i_13_170_2712_0,
    i_13_170_2713_0, i_13_170_2755_0, i_13_170_2953_0, i_13_170_2980_0,
    i_13_170_3051_0, i_13_170_3123_0, i_13_170_3235_0, i_13_170_3250_0,
    i_13_170_3334_0, i_13_170_3352_0, i_13_170_3487_0, i_13_170_3574_0,
    i_13_170_3592_0, i_13_170_3595_0, i_13_170_3684_0, i_13_170_3700_0,
    i_13_170_3729_0, i_13_170_3730_0, i_13_170_3816_0, i_13_170_3856_0,
    i_13_170_3901_0, i_13_170_3927_0, i_13_170_3928_0, i_13_170_3982_0,
    i_13_170_4009_0, i_13_170_4018_0, i_13_170_4045_0, i_13_170_4054_0,
    i_13_170_4081_0, i_13_170_4090_0, i_13_170_4096_0, i_13_170_4189_0,
    i_13_170_4215_0, i_13_170_4230_0, i_13_170_4234_0, i_13_170_4251_0,
    i_13_170_4252_0, i_13_170_4267_0, i_13_170_4296_0, i_13_170_4297_0,
    i_13_170_4405_0, i_13_170_4432_0, i_13_170_4558_0, i_13_170_4590_0,
    o_13_170_0_0  );
  input  i_13_170_48_0, i_13_170_136_0, i_13_170_144_0, i_13_170_211_0,
    i_13_170_229_0, i_13_170_271_0, i_13_170_283_0, i_13_170_300_0,
    i_13_170_382_0, i_13_170_517_0, i_13_170_571_0, i_13_170_585_0,
    i_13_170_639_0, i_13_170_705_0, i_13_170_711_0, i_13_170_738_0,
    i_13_170_796_0, i_13_170_940_0, i_13_170_999_0, i_13_170_1044_0,
    i_13_170_1101_0, i_13_170_1344_0, i_13_170_1377_0, i_13_170_1390_0,
    i_13_170_1399_0, i_13_170_1408_0, i_13_170_1432_0, i_13_170_1513_0,
    i_13_170_1632_0, i_13_170_1633_0, i_13_170_1639_0, i_13_170_1768_0,
    i_13_170_1776_0, i_13_170_1795_0, i_13_170_1848_0, i_13_170_1893_0,
    i_13_170_1936_0, i_13_170_1945_0, i_13_170_2029_0, i_13_170_2030_0,
    i_13_170_2053_0, i_13_170_2250_0, i_13_170_2251_0, i_13_170_2253_0,
    i_13_170_2278_0, i_13_170_2413_0, i_13_170_2424_0, i_13_170_2433_0,
    i_13_170_2497_0, i_13_170_2515_0, i_13_170_2542_0, i_13_170_2547_0,
    i_13_170_2614_0, i_13_170_2668_0, i_13_170_2674_0, i_13_170_2712_0,
    i_13_170_2713_0, i_13_170_2755_0, i_13_170_2953_0, i_13_170_2980_0,
    i_13_170_3051_0, i_13_170_3123_0, i_13_170_3235_0, i_13_170_3250_0,
    i_13_170_3334_0, i_13_170_3352_0, i_13_170_3487_0, i_13_170_3574_0,
    i_13_170_3592_0, i_13_170_3595_0, i_13_170_3684_0, i_13_170_3700_0,
    i_13_170_3729_0, i_13_170_3730_0, i_13_170_3816_0, i_13_170_3856_0,
    i_13_170_3901_0, i_13_170_3927_0, i_13_170_3928_0, i_13_170_3982_0,
    i_13_170_4009_0, i_13_170_4018_0, i_13_170_4045_0, i_13_170_4054_0,
    i_13_170_4081_0, i_13_170_4090_0, i_13_170_4096_0, i_13_170_4189_0,
    i_13_170_4215_0, i_13_170_4230_0, i_13_170_4234_0, i_13_170_4251_0,
    i_13_170_4252_0, i_13_170_4267_0, i_13_170_4296_0, i_13_170_4297_0,
    i_13_170_4405_0, i_13_170_4432_0, i_13_170_4558_0, i_13_170_4590_0;
  output o_13_170_0_0;
  assign o_13_170_0_0 = 0;
endmodule



// Benchmark "kernel_13_171" written by ABC on Sun Jul 19 10:47:48 2020

module kernel_13_171 ( 
    i_13_171_48_0, i_13_171_63_0, i_13_171_64_0, i_13_171_71_0,
    i_13_171_158_0, i_13_171_172_0, i_13_171_176_0, i_13_171_207_0,
    i_13_171_209_0, i_13_171_227_0, i_13_171_245_0, i_13_171_256_0,
    i_13_171_304_0, i_13_171_415_0, i_13_171_526_0, i_13_171_605_0,
    i_13_171_612_0, i_13_171_613_0, i_13_171_616_0, i_13_171_764_0,
    i_13_171_828_0, i_13_171_838_0, i_13_171_854_0, i_13_171_1075_0,
    i_13_171_1132_0, i_13_171_1227_0, i_13_171_1304_0, i_13_171_1305_0,
    i_13_171_1309_0, i_13_171_1360_0, i_13_171_1441_0, i_13_171_1443_0,
    i_13_171_1495_0, i_13_171_1521_0, i_13_171_1522_0, i_13_171_1523_0,
    i_13_171_1525_0, i_13_171_1548_0, i_13_171_1549_0, i_13_171_1593_0,
    i_13_171_1604_0, i_13_171_1638_0, i_13_171_1639_0, i_13_171_1696_0,
    i_13_171_1721_0, i_13_171_1728_0, i_13_171_1730_0, i_13_171_1799_0,
    i_13_171_1846_0, i_13_171_1926_0, i_13_171_1930_0, i_13_171_1931_0,
    i_13_171_2142_0, i_13_171_2182_0, i_13_171_2199_0, i_13_171_2243_0,
    i_13_171_2297_0, i_13_171_2407_0, i_13_171_2421_0, i_13_171_2430_0,
    i_13_171_2505_0, i_13_171_2554_0, i_13_171_2673_0, i_13_171_2675_0,
    i_13_171_2722_0, i_13_171_2748_0, i_13_171_2881_0, i_13_171_2883_0,
    i_13_171_3240_0, i_13_171_3241_0, i_13_171_3288_0, i_13_171_3367_0,
    i_13_171_3395_0, i_13_171_3414_0, i_13_171_3420_0, i_13_171_3538_0,
    i_13_171_3539_0, i_13_171_3548_0, i_13_171_3636_0, i_13_171_3637_0,
    i_13_171_3638_0, i_13_171_3640_0, i_13_171_3758_0, i_13_171_3766_0,
    i_13_171_3843_0, i_13_171_3845_0, i_13_171_3889_0, i_13_171_3898_0,
    i_13_171_3913_0, i_13_171_3916_0, i_13_171_3934_0, i_13_171_4217_0,
    i_13_171_4312_0, i_13_171_4322_0, i_13_171_4472_0, i_13_171_4509_0,
    i_13_171_4511_0, i_13_171_4522_0, i_13_171_4590_0, i_13_171_4607_0,
    o_13_171_0_0  );
  input  i_13_171_48_0, i_13_171_63_0, i_13_171_64_0, i_13_171_71_0,
    i_13_171_158_0, i_13_171_172_0, i_13_171_176_0, i_13_171_207_0,
    i_13_171_209_0, i_13_171_227_0, i_13_171_245_0, i_13_171_256_0,
    i_13_171_304_0, i_13_171_415_0, i_13_171_526_0, i_13_171_605_0,
    i_13_171_612_0, i_13_171_613_0, i_13_171_616_0, i_13_171_764_0,
    i_13_171_828_0, i_13_171_838_0, i_13_171_854_0, i_13_171_1075_0,
    i_13_171_1132_0, i_13_171_1227_0, i_13_171_1304_0, i_13_171_1305_0,
    i_13_171_1309_0, i_13_171_1360_0, i_13_171_1441_0, i_13_171_1443_0,
    i_13_171_1495_0, i_13_171_1521_0, i_13_171_1522_0, i_13_171_1523_0,
    i_13_171_1525_0, i_13_171_1548_0, i_13_171_1549_0, i_13_171_1593_0,
    i_13_171_1604_0, i_13_171_1638_0, i_13_171_1639_0, i_13_171_1696_0,
    i_13_171_1721_0, i_13_171_1728_0, i_13_171_1730_0, i_13_171_1799_0,
    i_13_171_1846_0, i_13_171_1926_0, i_13_171_1930_0, i_13_171_1931_0,
    i_13_171_2142_0, i_13_171_2182_0, i_13_171_2199_0, i_13_171_2243_0,
    i_13_171_2297_0, i_13_171_2407_0, i_13_171_2421_0, i_13_171_2430_0,
    i_13_171_2505_0, i_13_171_2554_0, i_13_171_2673_0, i_13_171_2675_0,
    i_13_171_2722_0, i_13_171_2748_0, i_13_171_2881_0, i_13_171_2883_0,
    i_13_171_3240_0, i_13_171_3241_0, i_13_171_3288_0, i_13_171_3367_0,
    i_13_171_3395_0, i_13_171_3414_0, i_13_171_3420_0, i_13_171_3538_0,
    i_13_171_3539_0, i_13_171_3548_0, i_13_171_3636_0, i_13_171_3637_0,
    i_13_171_3638_0, i_13_171_3640_0, i_13_171_3758_0, i_13_171_3766_0,
    i_13_171_3843_0, i_13_171_3845_0, i_13_171_3889_0, i_13_171_3898_0,
    i_13_171_3913_0, i_13_171_3916_0, i_13_171_3934_0, i_13_171_4217_0,
    i_13_171_4312_0, i_13_171_4322_0, i_13_171_4472_0, i_13_171_4509_0,
    i_13_171_4511_0, i_13_171_4522_0, i_13_171_4590_0, i_13_171_4607_0;
  output o_13_171_0_0;
  assign o_13_171_0_0 = ~((~i_13_171_1522_0 & ((~i_13_171_3843_0 & i_13_171_4509_0) | (~i_13_171_1523_0 & i_13_171_1525_0 & ~i_13_171_4509_0))) | (~i_13_171_1728_0 & ((~i_13_171_2881_0 & ~i_13_171_4312_0) | (~i_13_171_1305_0 & ~i_13_171_2297_0 & ~i_13_171_4509_0))) | (~i_13_171_4509_0 & ((~i_13_171_3241_0 & i_13_171_3766_0) | (~i_13_171_838_0 & ~i_13_171_3898_0))) | (i_13_171_1075_0 & ~i_13_171_3538_0));
endmodule



// Benchmark "kernel_13_172" written by ABC on Sun Jul 19 10:47:49 2020

module kernel_13_172 ( 
    i_13_172_35_0, i_13_172_52_0, i_13_172_69_0, i_13_172_70_0,
    i_13_172_71_0, i_13_172_78_0, i_13_172_90_0, i_13_172_127_0,
    i_13_172_314_0, i_13_172_402_0, i_13_172_449_0, i_13_172_537_0,
    i_13_172_565_0, i_13_172_641_0, i_13_172_673_0, i_13_172_679_0,
    i_13_172_737_0, i_13_172_763_0, i_13_172_823_0, i_13_172_843_0,
    i_13_172_933_0, i_13_172_1021_0, i_13_172_1101_0, i_13_172_1102_0,
    i_13_172_1105_0, i_13_172_1106_0, i_13_172_1151_0, i_13_172_1228_0,
    i_13_172_1263_0, i_13_172_1276_0, i_13_172_1345_0, i_13_172_1363_0,
    i_13_172_1401_0, i_13_172_1402_0, i_13_172_1519_0, i_13_172_1599_0,
    i_13_172_1627_0, i_13_172_1644_0, i_13_172_1725_0, i_13_172_1726_0,
    i_13_172_1777_0, i_13_172_1780_0, i_13_172_1781_0, i_13_172_1797_0,
    i_13_172_1799_0, i_13_172_1827_0, i_13_172_1853_0, i_13_172_1858_0,
    i_13_172_1925_0, i_13_172_1948_0, i_13_172_1995_0, i_13_172_2054_0,
    i_13_172_2176_0, i_13_172_2208_0, i_13_172_2312_0, i_13_172_2617_0,
    i_13_172_2638_0, i_13_172_2695_0, i_13_172_2698_0, i_13_172_2715_0,
    i_13_172_2725_0, i_13_172_2752_0, i_13_172_2760_0, i_13_172_2770_0,
    i_13_172_2851_0, i_13_172_2878_0, i_13_172_2901_0, i_13_172_2905_0,
    i_13_172_3039_0, i_13_172_3067_0, i_13_172_3128_0, i_13_172_3367_0,
    i_13_172_3370_0, i_13_172_3417_0, i_13_172_3418_0, i_13_172_3441_0,
    i_13_172_3534_0, i_13_172_3580_0, i_13_172_3595_0, i_13_172_3640_0,
    i_13_172_3648_0, i_13_172_3684_0, i_13_172_3685_0, i_13_172_3739_0,
    i_13_172_3757_0, i_13_172_3767_0, i_13_172_3787_0, i_13_172_3796_0,
    i_13_172_3869_0, i_13_172_3895_0, i_13_172_3913_0, i_13_172_3928_0,
    i_13_172_3931_0, i_13_172_3991_0, i_13_172_3994_0, i_13_172_4264_0,
    i_13_172_4335_0, i_13_172_4434_0, i_13_172_4450_0, i_13_172_4451_0,
    o_13_172_0_0  );
  input  i_13_172_35_0, i_13_172_52_0, i_13_172_69_0, i_13_172_70_0,
    i_13_172_71_0, i_13_172_78_0, i_13_172_90_0, i_13_172_127_0,
    i_13_172_314_0, i_13_172_402_0, i_13_172_449_0, i_13_172_537_0,
    i_13_172_565_0, i_13_172_641_0, i_13_172_673_0, i_13_172_679_0,
    i_13_172_737_0, i_13_172_763_0, i_13_172_823_0, i_13_172_843_0,
    i_13_172_933_0, i_13_172_1021_0, i_13_172_1101_0, i_13_172_1102_0,
    i_13_172_1105_0, i_13_172_1106_0, i_13_172_1151_0, i_13_172_1228_0,
    i_13_172_1263_0, i_13_172_1276_0, i_13_172_1345_0, i_13_172_1363_0,
    i_13_172_1401_0, i_13_172_1402_0, i_13_172_1519_0, i_13_172_1599_0,
    i_13_172_1627_0, i_13_172_1644_0, i_13_172_1725_0, i_13_172_1726_0,
    i_13_172_1777_0, i_13_172_1780_0, i_13_172_1781_0, i_13_172_1797_0,
    i_13_172_1799_0, i_13_172_1827_0, i_13_172_1853_0, i_13_172_1858_0,
    i_13_172_1925_0, i_13_172_1948_0, i_13_172_1995_0, i_13_172_2054_0,
    i_13_172_2176_0, i_13_172_2208_0, i_13_172_2312_0, i_13_172_2617_0,
    i_13_172_2638_0, i_13_172_2695_0, i_13_172_2698_0, i_13_172_2715_0,
    i_13_172_2725_0, i_13_172_2752_0, i_13_172_2760_0, i_13_172_2770_0,
    i_13_172_2851_0, i_13_172_2878_0, i_13_172_2901_0, i_13_172_2905_0,
    i_13_172_3039_0, i_13_172_3067_0, i_13_172_3128_0, i_13_172_3367_0,
    i_13_172_3370_0, i_13_172_3417_0, i_13_172_3418_0, i_13_172_3441_0,
    i_13_172_3534_0, i_13_172_3580_0, i_13_172_3595_0, i_13_172_3640_0,
    i_13_172_3648_0, i_13_172_3684_0, i_13_172_3685_0, i_13_172_3739_0,
    i_13_172_3757_0, i_13_172_3767_0, i_13_172_3787_0, i_13_172_3796_0,
    i_13_172_3869_0, i_13_172_3895_0, i_13_172_3913_0, i_13_172_3928_0,
    i_13_172_3931_0, i_13_172_3991_0, i_13_172_3994_0, i_13_172_4264_0,
    i_13_172_4335_0, i_13_172_4434_0, i_13_172_4450_0, i_13_172_4451_0;
  output o_13_172_0_0;
  assign o_13_172_0_0 = ~((~i_13_172_1948_0 & ((~i_13_172_763_0 & ~i_13_172_3441_0) | (~i_13_172_1401_0 & i_13_172_2695_0 & ~i_13_172_3931_0))) | (~i_13_172_537_0 & ~i_13_172_673_0 & ~i_13_172_1402_0) | (~i_13_172_2176_0 & i_13_172_3991_0));
endmodule



// Benchmark "kernel_13_173" written by ABC on Sun Jul 19 10:47:50 2020

module kernel_13_173 ( 
    i_13_173_41_0, i_13_173_74_0, i_13_173_104_0, i_13_173_109_0,
    i_13_173_110_0, i_13_173_280_0, i_13_173_283_0, i_13_173_320_0,
    i_13_173_406_0, i_13_173_452_0, i_13_173_506_0, i_13_173_553_0,
    i_13_173_581_0, i_13_173_599_0, i_13_173_604_0, i_13_173_622_0,
    i_13_173_677_0, i_13_173_680_0, i_13_173_794_0, i_13_173_856_0,
    i_13_173_859_0, i_13_173_946_0, i_13_173_947_0, i_13_173_1019_0,
    i_13_173_1022_0, i_13_173_1084_0, i_13_173_1282_0, i_13_173_1424_0,
    i_13_173_1436_0, i_13_173_1444_0, i_13_173_1472_0, i_13_173_1486_0,
    i_13_173_1487_0, i_13_173_1543_0, i_13_173_1553_0, i_13_173_1621_0,
    i_13_173_1630_0, i_13_173_1670_0, i_13_173_1838_0, i_13_173_1841_0,
    i_13_173_1856_0, i_13_173_1927_0, i_13_173_1999_0, i_13_173_2047_0,
    i_13_173_2053_0, i_13_173_2146_0, i_13_173_2263_0, i_13_173_2314_0,
    i_13_173_2396_0, i_13_173_2432_0, i_13_173_2435_0, i_13_173_2458_0,
    i_13_173_2459_0, i_13_173_2462_0, i_13_173_2501_0, i_13_173_2503_0,
    i_13_173_2504_0, i_13_173_2506_0, i_13_173_2507_0, i_13_173_2521_0,
    i_13_173_2529_0, i_13_173_2539_0, i_13_173_2540_0, i_13_173_2611_0,
    i_13_173_2612_0, i_13_173_2714_0, i_13_173_2746_0, i_13_173_2911_0,
    i_13_173_2920_0, i_13_173_3071_0, i_13_173_3124_0, i_13_173_3143_0,
    i_13_173_3145_0, i_13_173_3146_0, i_13_173_3154_0, i_13_173_3340_0,
    i_13_173_3422_0, i_13_173_3523_0, i_13_173_3529_0, i_13_173_3530_0,
    i_13_173_3542_0, i_13_173_3577_0, i_13_173_3661_0, i_13_173_3757_0,
    i_13_173_3844_0, i_13_173_3871_0, i_13_173_3889_0, i_13_173_3890_0,
    i_13_173_3928_0, i_13_173_4046_0, i_13_173_4063_0, i_13_173_4223_0,
    i_13_173_4252_0, i_13_173_4253_0, i_13_173_4325_0, i_13_173_4366_0,
    i_13_173_4424_0, i_13_173_4519_0, i_13_173_4520_0, i_13_173_4556_0,
    o_13_173_0_0  );
  input  i_13_173_41_0, i_13_173_74_0, i_13_173_104_0, i_13_173_109_0,
    i_13_173_110_0, i_13_173_280_0, i_13_173_283_0, i_13_173_320_0,
    i_13_173_406_0, i_13_173_452_0, i_13_173_506_0, i_13_173_553_0,
    i_13_173_581_0, i_13_173_599_0, i_13_173_604_0, i_13_173_622_0,
    i_13_173_677_0, i_13_173_680_0, i_13_173_794_0, i_13_173_856_0,
    i_13_173_859_0, i_13_173_946_0, i_13_173_947_0, i_13_173_1019_0,
    i_13_173_1022_0, i_13_173_1084_0, i_13_173_1282_0, i_13_173_1424_0,
    i_13_173_1436_0, i_13_173_1444_0, i_13_173_1472_0, i_13_173_1486_0,
    i_13_173_1487_0, i_13_173_1543_0, i_13_173_1553_0, i_13_173_1621_0,
    i_13_173_1630_0, i_13_173_1670_0, i_13_173_1838_0, i_13_173_1841_0,
    i_13_173_1856_0, i_13_173_1927_0, i_13_173_1999_0, i_13_173_2047_0,
    i_13_173_2053_0, i_13_173_2146_0, i_13_173_2263_0, i_13_173_2314_0,
    i_13_173_2396_0, i_13_173_2432_0, i_13_173_2435_0, i_13_173_2458_0,
    i_13_173_2459_0, i_13_173_2462_0, i_13_173_2501_0, i_13_173_2503_0,
    i_13_173_2504_0, i_13_173_2506_0, i_13_173_2507_0, i_13_173_2521_0,
    i_13_173_2529_0, i_13_173_2539_0, i_13_173_2540_0, i_13_173_2611_0,
    i_13_173_2612_0, i_13_173_2714_0, i_13_173_2746_0, i_13_173_2911_0,
    i_13_173_2920_0, i_13_173_3071_0, i_13_173_3124_0, i_13_173_3143_0,
    i_13_173_3145_0, i_13_173_3146_0, i_13_173_3154_0, i_13_173_3340_0,
    i_13_173_3422_0, i_13_173_3523_0, i_13_173_3529_0, i_13_173_3530_0,
    i_13_173_3542_0, i_13_173_3577_0, i_13_173_3661_0, i_13_173_3757_0,
    i_13_173_3844_0, i_13_173_3871_0, i_13_173_3889_0, i_13_173_3890_0,
    i_13_173_3928_0, i_13_173_4046_0, i_13_173_4063_0, i_13_173_4223_0,
    i_13_173_4252_0, i_13_173_4253_0, i_13_173_4325_0, i_13_173_4366_0,
    i_13_173_4424_0, i_13_173_4519_0, i_13_173_4520_0, i_13_173_4556_0;
  output o_13_173_0_0;
  assign o_13_173_0_0 = ~((~i_13_173_3530_0 & ~i_13_173_4325_0) | (~i_13_173_110_0 & ~i_13_173_1486_0));
endmodule



// Benchmark "kernel_13_174" written by ABC on Sun Jul 19 10:47:50 2020

module kernel_13_174 ( 
    i_13_174_67_0, i_13_174_106_0, i_13_174_123_0, i_13_174_138_0,
    i_13_174_139_0, i_13_174_161_0, i_13_174_166_0, i_13_174_232_0,
    i_13_174_247_0, i_13_174_310_0, i_13_174_327_0, i_13_174_328_0,
    i_13_174_430_0, i_13_174_526_0, i_13_174_537_0, i_13_174_571_0,
    i_13_174_598_0, i_13_174_670_0, i_13_174_717_0, i_13_174_780_0,
    i_13_174_825_0, i_13_174_832_0, i_13_174_841_0, i_13_174_861_0,
    i_13_174_890_0, i_13_174_894_0, i_13_174_1023_0, i_13_174_1024_0,
    i_13_174_1095_0, i_13_174_1096_0, i_13_174_1111_0, i_13_174_1281_0,
    i_13_174_1299_0, i_13_174_1303_0, i_13_174_1326_0, i_13_174_1464_0,
    i_13_174_1488_0, i_13_174_1489_0, i_13_174_1490_0, i_13_174_1515_0,
    i_13_174_1777_0, i_13_174_1785_0, i_13_174_1786_0, i_13_174_1788_0,
    i_13_174_1857_0, i_13_174_1858_0, i_13_174_1884_0, i_13_174_1887_0,
    i_13_174_1930_0, i_13_174_2056_0, i_13_174_2146_0, i_13_174_2175_0,
    i_13_174_2190_0, i_13_174_2263_0, i_13_174_2309_0, i_13_174_2310_0,
    i_13_174_2311_0, i_13_174_2316_0, i_13_174_2460_0, i_13_174_2461_0,
    i_13_174_2462_0, i_13_174_2464_0, i_13_174_2500_0, i_13_174_2506_0,
    i_13_174_2532_0, i_13_174_2565_0, i_13_174_2566_0, i_13_174_2613_0,
    i_13_174_2632_0, i_13_174_2885_0, i_13_174_2941_0, i_13_174_3087_0,
    i_13_174_3148_0, i_13_174_3171_0, i_13_174_3173_0, i_13_174_3174_0,
    i_13_174_3348_0, i_13_174_3432_0, i_13_174_3481_0, i_13_174_3532_0,
    i_13_174_3534_0, i_13_174_3535_0, i_13_174_3661_0, i_13_174_3732_0,
    i_13_174_3741_0, i_13_174_3783_0, i_13_174_3797_0, i_13_174_3820_0,
    i_13_174_3913_0, i_13_174_3923_0, i_13_174_3932_0, i_13_174_4012_0,
    i_13_174_4210_0, i_13_174_4237_0, i_13_174_4341_0, i_13_174_4443_0,
    i_13_174_4514_0, i_13_174_4521_0, i_13_174_4522_0, i_13_174_4567_0,
    o_13_174_0_0  );
  input  i_13_174_67_0, i_13_174_106_0, i_13_174_123_0, i_13_174_138_0,
    i_13_174_139_0, i_13_174_161_0, i_13_174_166_0, i_13_174_232_0,
    i_13_174_247_0, i_13_174_310_0, i_13_174_327_0, i_13_174_328_0,
    i_13_174_430_0, i_13_174_526_0, i_13_174_537_0, i_13_174_571_0,
    i_13_174_598_0, i_13_174_670_0, i_13_174_717_0, i_13_174_780_0,
    i_13_174_825_0, i_13_174_832_0, i_13_174_841_0, i_13_174_861_0,
    i_13_174_890_0, i_13_174_894_0, i_13_174_1023_0, i_13_174_1024_0,
    i_13_174_1095_0, i_13_174_1096_0, i_13_174_1111_0, i_13_174_1281_0,
    i_13_174_1299_0, i_13_174_1303_0, i_13_174_1326_0, i_13_174_1464_0,
    i_13_174_1488_0, i_13_174_1489_0, i_13_174_1490_0, i_13_174_1515_0,
    i_13_174_1777_0, i_13_174_1785_0, i_13_174_1786_0, i_13_174_1788_0,
    i_13_174_1857_0, i_13_174_1858_0, i_13_174_1884_0, i_13_174_1887_0,
    i_13_174_1930_0, i_13_174_2056_0, i_13_174_2146_0, i_13_174_2175_0,
    i_13_174_2190_0, i_13_174_2263_0, i_13_174_2309_0, i_13_174_2310_0,
    i_13_174_2311_0, i_13_174_2316_0, i_13_174_2460_0, i_13_174_2461_0,
    i_13_174_2462_0, i_13_174_2464_0, i_13_174_2500_0, i_13_174_2506_0,
    i_13_174_2532_0, i_13_174_2565_0, i_13_174_2566_0, i_13_174_2613_0,
    i_13_174_2632_0, i_13_174_2885_0, i_13_174_2941_0, i_13_174_3087_0,
    i_13_174_3148_0, i_13_174_3171_0, i_13_174_3173_0, i_13_174_3174_0,
    i_13_174_3348_0, i_13_174_3432_0, i_13_174_3481_0, i_13_174_3532_0,
    i_13_174_3534_0, i_13_174_3535_0, i_13_174_3661_0, i_13_174_3732_0,
    i_13_174_3741_0, i_13_174_3783_0, i_13_174_3797_0, i_13_174_3820_0,
    i_13_174_3913_0, i_13_174_3923_0, i_13_174_3932_0, i_13_174_4012_0,
    i_13_174_4210_0, i_13_174_4237_0, i_13_174_4341_0, i_13_174_4443_0,
    i_13_174_4514_0, i_13_174_4521_0, i_13_174_4522_0, i_13_174_4567_0;
  output o_13_174_0_0;
  assign o_13_174_0_0 = ~((~i_13_174_3534_0 & (~i_13_174_537_0 | (i_13_174_526_0 & ~i_13_174_3535_0))) | ~i_13_174_3171_0 | (~i_13_174_3148_0 & ~i_13_174_3174_0) | (~i_13_174_1857_0 & i_13_174_3783_0) | (~i_13_174_1887_0 & i_13_174_4237_0));
endmodule



// Benchmark "kernel_13_175" written by ABC on Sun Jul 19 10:47:51 2020

module kernel_13_175 ( 
    i_13_175_76_0, i_13_175_77_0, i_13_175_88_0, i_13_175_94_0,
    i_13_175_130_0, i_13_175_134_0, i_13_175_256_0, i_13_175_269_0,
    i_13_175_332_0, i_13_175_358_0, i_13_175_359_0, i_13_175_370_0,
    i_13_175_371_0, i_13_175_400_0, i_13_175_458_0, i_13_175_520_0,
    i_13_175_571_0, i_13_175_611_0, i_13_175_617_0, i_13_175_667_0,
    i_13_175_671_0, i_13_175_823_0, i_13_175_842_0, i_13_175_980_0,
    i_13_175_1091_0, i_13_175_1115_0, i_13_175_1213_0, i_13_175_1282_0,
    i_13_175_1348_0, i_13_175_1400_0, i_13_175_1402_0, i_13_175_1403_0,
    i_13_175_1508_0, i_13_175_1519_0, i_13_175_1660_0, i_13_175_1750_0,
    i_13_175_1763_0, i_13_175_1778_0, i_13_175_1951_0, i_13_175_1952_0,
    i_13_175_2032_0, i_13_175_2033_0, i_13_175_2059_0, i_13_175_2060_0,
    i_13_175_2141_0, i_13_175_2191_0, i_13_175_2203_0, i_13_175_2240_0,
    i_13_175_2284_0, i_13_175_2285_0, i_13_175_2321_0, i_13_175_2348_0,
    i_13_175_2408_0, i_13_175_2410_0, i_13_175_2447_0, i_13_175_2497_0,
    i_13_175_2503_0, i_13_175_2510_0, i_13_175_2515_0, i_13_175_2516_0,
    i_13_175_2555_0, i_13_175_2590_0, i_13_175_2696_0, i_13_175_2705_0,
    i_13_175_2902_0, i_13_175_2920_0, i_13_175_2923_0, i_13_175_2924_0,
    i_13_175_2959_0, i_13_175_3013_0, i_13_175_3073_0, i_13_175_3218_0,
    i_13_175_3373_0, i_13_175_3374_0, i_13_175_3419_0, i_13_175_3580_0,
    i_13_175_3581_0, i_13_175_3598_0, i_13_175_3599_0, i_13_175_3622_0,
    i_13_175_3623_0, i_13_175_3634_0, i_13_175_3635_0, i_13_175_3784_0,
    i_13_175_3788_0, i_13_175_3988_0, i_13_175_3991_0, i_13_175_4076_0,
    i_13_175_4190_0, i_13_175_4208_0, i_13_175_4216_0, i_13_175_4237_0,
    i_13_175_4264_0, i_13_175_4265_0, i_13_175_4333_0, i_13_175_4334_0,
    i_13_175_4378_0, i_13_175_4433_0, i_13_175_4453_0, i_13_175_4454_0,
    o_13_175_0_0  );
  input  i_13_175_76_0, i_13_175_77_0, i_13_175_88_0, i_13_175_94_0,
    i_13_175_130_0, i_13_175_134_0, i_13_175_256_0, i_13_175_269_0,
    i_13_175_332_0, i_13_175_358_0, i_13_175_359_0, i_13_175_370_0,
    i_13_175_371_0, i_13_175_400_0, i_13_175_458_0, i_13_175_520_0,
    i_13_175_571_0, i_13_175_611_0, i_13_175_617_0, i_13_175_667_0,
    i_13_175_671_0, i_13_175_823_0, i_13_175_842_0, i_13_175_980_0,
    i_13_175_1091_0, i_13_175_1115_0, i_13_175_1213_0, i_13_175_1282_0,
    i_13_175_1348_0, i_13_175_1400_0, i_13_175_1402_0, i_13_175_1403_0,
    i_13_175_1508_0, i_13_175_1519_0, i_13_175_1660_0, i_13_175_1750_0,
    i_13_175_1763_0, i_13_175_1778_0, i_13_175_1951_0, i_13_175_1952_0,
    i_13_175_2032_0, i_13_175_2033_0, i_13_175_2059_0, i_13_175_2060_0,
    i_13_175_2141_0, i_13_175_2191_0, i_13_175_2203_0, i_13_175_2240_0,
    i_13_175_2284_0, i_13_175_2285_0, i_13_175_2321_0, i_13_175_2348_0,
    i_13_175_2408_0, i_13_175_2410_0, i_13_175_2447_0, i_13_175_2497_0,
    i_13_175_2503_0, i_13_175_2510_0, i_13_175_2515_0, i_13_175_2516_0,
    i_13_175_2555_0, i_13_175_2590_0, i_13_175_2696_0, i_13_175_2705_0,
    i_13_175_2902_0, i_13_175_2920_0, i_13_175_2923_0, i_13_175_2924_0,
    i_13_175_2959_0, i_13_175_3013_0, i_13_175_3073_0, i_13_175_3218_0,
    i_13_175_3373_0, i_13_175_3374_0, i_13_175_3419_0, i_13_175_3580_0,
    i_13_175_3581_0, i_13_175_3598_0, i_13_175_3599_0, i_13_175_3622_0,
    i_13_175_3623_0, i_13_175_3634_0, i_13_175_3635_0, i_13_175_3784_0,
    i_13_175_3788_0, i_13_175_3988_0, i_13_175_3991_0, i_13_175_4076_0,
    i_13_175_4190_0, i_13_175_4208_0, i_13_175_4216_0, i_13_175_4237_0,
    i_13_175_4264_0, i_13_175_4265_0, i_13_175_4333_0, i_13_175_4334_0,
    i_13_175_4378_0, i_13_175_4433_0, i_13_175_4453_0, i_13_175_4454_0;
  output o_13_175_0_0;
  assign o_13_175_0_0 = ~(~i_13_175_2033_0 | ~i_13_175_4454_0);
endmodule



// Benchmark "kernel_13_176" written by ABC on Sun Jul 19 10:47:52 2020

module kernel_13_176 ( 
    i_13_176_68_0, i_13_176_94_0, i_13_176_112_0, i_13_176_139_0,
    i_13_176_140_0, i_13_176_237_0, i_13_176_320_0, i_13_176_380_0,
    i_13_176_445_0, i_13_176_524_0, i_13_176_553_0, i_13_176_586_0,
    i_13_176_587_0, i_13_176_607_0, i_13_176_614_0, i_13_176_686_0,
    i_13_176_696_0, i_13_176_698_0, i_13_176_739_0, i_13_176_796_0,
    i_13_176_883_0, i_13_176_1075_0, i_13_176_1103_0, i_13_176_1117_0,
    i_13_176_1208_0, i_13_176_1268_0, i_13_176_1273_0, i_13_176_1274_0,
    i_13_176_1298_0, i_13_176_1342_0, i_13_176_1343_0, i_13_176_1400_0,
    i_13_176_1441_0, i_13_176_1442_0, i_13_176_1468_0, i_13_176_1507_0,
    i_13_176_1516_0, i_13_176_1568_0, i_13_176_1598_0, i_13_176_1712_0,
    i_13_176_1775_0, i_13_176_1778_0, i_13_176_1810_0, i_13_176_1811_0,
    i_13_176_1921_0, i_13_176_1928_0, i_13_176_1945_0, i_13_176_1990_0,
    i_13_176_1991_0, i_13_176_2053_0, i_13_176_2054_0, i_13_176_2189_0,
    i_13_176_2197_0, i_13_176_2236_0, i_13_176_2260_0, i_13_176_2278_0,
    i_13_176_2279_0, i_13_176_2320_0, i_13_176_2377_0, i_13_176_2503_0,
    i_13_176_2593_0, i_13_176_2647_0, i_13_176_2675_0, i_13_176_2696_0,
    i_13_176_2710_0, i_13_176_2720_0, i_13_176_2723_0, i_13_176_2782_0,
    i_13_176_2899_0, i_13_176_2921_0, i_13_176_2998_0, i_13_176_3001_0,
    i_13_176_3058_0, i_13_176_3059_0, i_13_176_3061_0, i_13_176_3064_0,
    i_13_176_3065_0, i_13_176_3136_0, i_13_176_3208_0, i_13_176_3367_0,
    i_13_176_3368_0, i_13_176_3386_0, i_13_176_3415_0, i_13_176_3439_0,
    i_13_176_3593_0, i_13_176_3650_0, i_13_176_3856_0, i_13_176_4096_0,
    i_13_176_4187_0, i_13_176_4231_0, i_13_176_4258_0, i_13_176_4259_0,
    i_13_176_4268_0, i_13_176_4339_0, i_13_176_4393_0, i_13_176_4394_0,
    i_13_176_4405_0, i_13_176_4429_0, i_13_176_4447_0, i_13_176_4448_0,
    o_13_176_0_0  );
  input  i_13_176_68_0, i_13_176_94_0, i_13_176_112_0, i_13_176_139_0,
    i_13_176_140_0, i_13_176_237_0, i_13_176_320_0, i_13_176_380_0,
    i_13_176_445_0, i_13_176_524_0, i_13_176_553_0, i_13_176_586_0,
    i_13_176_587_0, i_13_176_607_0, i_13_176_614_0, i_13_176_686_0,
    i_13_176_696_0, i_13_176_698_0, i_13_176_739_0, i_13_176_796_0,
    i_13_176_883_0, i_13_176_1075_0, i_13_176_1103_0, i_13_176_1117_0,
    i_13_176_1208_0, i_13_176_1268_0, i_13_176_1273_0, i_13_176_1274_0,
    i_13_176_1298_0, i_13_176_1342_0, i_13_176_1343_0, i_13_176_1400_0,
    i_13_176_1441_0, i_13_176_1442_0, i_13_176_1468_0, i_13_176_1507_0,
    i_13_176_1516_0, i_13_176_1568_0, i_13_176_1598_0, i_13_176_1712_0,
    i_13_176_1775_0, i_13_176_1778_0, i_13_176_1810_0, i_13_176_1811_0,
    i_13_176_1921_0, i_13_176_1928_0, i_13_176_1945_0, i_13_176_1990_0,
    i_13_176_1991_0, i_13_176_2053_0, i_13_176_2054_0, i_13_176_2189_0,
    i_13_176_2197_0, i_13_176_2236_0, i_13_176_2260_0, i_13_176_2278_0,
    i_13_176_2279_0, i_13_176_2320_0, i_13_176_2377_0, i_13_176_2503_0,
    i_13_176_2593_0, i_13_176_2647_0, i_13_176_2675_0, i_13_176_2696_0,
    i_13_176_2710_0, i_13_176_2720_0, i_13_176_2723_0, i_13_176_2782_0,
    i_13_176_2899_0, i_13_176_2921_0, i_13_176_2998_0, i_13_176_3001_0,
    i_13_176_3058_0, i_13_176_3059_0, i_13_176_3061_0, i_13_176_3064_0,
    i_13_176_3065_0, i_13_176_3136_0, i_13_176_3208_0, i_13_176_3367_0,
    i_13_176_3368_0, i_13_176_3386_0, i_13_176_3415_0, i_13_176_3439_0,
    i_13_176_3593_0, i_13_176_3650_0, i_13_176_3856_0, i_13_176_4096_0,
    i_13_176_4187_0, i_13_176_4231_0, i_13_176_4258_0, i_13_176_4259_0,
    i_13_176_4268_0, i_13_176_4339_0, i_13_176_4393_0, i_13_176_4394_0,
    i_13_176_4405_0, i_13_176_4429_0, i_13_176_4447_0, i_13_176_4448_0;
  output o_13_176_0_0;
  assign o_13_176_0_0 = 0;
endmodule



// Benchmark "kernel_13_177" written by ABC on Sun Jul 19 10:47:53 2020

module kernel_13_177 ( 
    i_13_177_52_0, i_13_177_73_0, i_13_177_76_0, i_13_177_121_0,
    i_13_177_158_0, i_13_177_205_0, i_13_177_259_0, i_13_177_275_0,
    i_13_177_277_0, i_13_177_310_0, i_13_177_355_0, i_13_177_450_0,
    i_13_177_451_0, i_13_177_452_0, i_13_177_454_0, i_13_177_661_0,
    i_13_177_665_0, i_13_177_674_0, i_13_177_716_0, i_13_177_874_0,
    i_13_177_929_0, i_13_177_952_0, i_13_177_1063_0, i_13_177_1139_0,
    i_13_177_1151_0, i_13_177_1228_0, i_13_177_1229_0, i_13_177_1256_0,
    i_13_177_1258_0, i_13_177_1408_0, i_13_177_1411_0, i_13_177_1412_0,
    i_13_177_1469_0, i_13_177_1516_0, i_13_177_1528_0, i_13_177_1679_0,
    i_13_177_1681_0, i_13_177_1732_0, i_13_177_1736_0, i_13_177_1768_0,
    i_13_177_1769_0, i_13_177_1781_0, i_13_177_1805_0, i_13_177_1895_0,
    i_13_177_2021_0, i_13_177_2056_0, i_13_177_2111_0, i_13_177_2149_0,
    i_13_177_2284_0, i_13_177_2299_0, i_13_177_2300_0, i_13_177_2354_0,
    i_13_177_2572_0, i_13_177_2596_0, i_13_177_2597_0, i_13_177_2614_0,
    i_13_177_2615_0, i_13_177_2617_0, i_13_177_2665_0, i_13_177_2708_0,
    i_13_177_2782_0, i_13_177_2891_0, i_13_177_2900_0, i_13_177_2983_0,
    i_13_177_2987_0, i_13_177_3029_0, i_13_177_3032_0, i_13_177_3114_0,
    i_13_177_3130_0, i_13_177_3157_0, i_13_177_3215_0, i_13_177_3218_0,
    i_13_177_3287_0, i_13_177_3313_0, i_13_177_3355_0, i_13_177_3461_0,
    i_13_177_3467_0, i_13_177_3488_0, i_13_177_3521_0, i_13_177_3598_0,
    i_13_177_3687_0, i_13_177_3730_0, i_13_177_3757_0, i_13_177_3784_0,
    i_13_177_3875_0, i_13_177_3979_0, i_13_177_4055_0, i_13_177_4073_0,
    i_13_177_4088_0, i_13_177_4102_0, i_13_177_4162_0, i_13_177_4163_0,
    i_13_177_4228_0, i_13_177_4237_0, i_13_177_4268_0, i_13_177_4372_0,
    i_13_177_4448_0, i_13_177_4517_0, i_13_177_4559_0, i_13_177_4607_0,
    o_13_177_0_0  );
  input  i_13_177_52_0, i_13_177_73_0, i_13_177_76_0, i_13_177_121_0,
    i_13_177_158_0, i_13_177_205_0, i_13_177_259_0, i_13_177_275_0,
    i_13_177_277_0, i_13_177_310_0, i_13_177_355_0, i_13_177_450_0,
    i_13_177_451_0, i_13_177_452_0, i_13_177_454_0, i_13_177_661_0,
    i_13_177_665_0, i_13_177_674_0, i_13_177_716_0, i_13_177_874_0,
    i_13_177_929_0, i_13_177_952_0, i_13_177_1063_0, i_13_177_1139_0,
    i_13_177_1151_0, i_13_177_1228_0, i_13_177_1229_0, i_13_177_1256_0,
    i_13_177_1258_0, i_13_177_1408_0, i_13_177_1411_0, i_13_177_1412_0,
    i_13_177_1469_0, i_13_177_1516_0, i_13_177_1528_0, i_13_177_1679_0,
    i_13_177_1681_0, i_13_177_1732_0, i_13_177_1736_0, i_13_177_1768_0,
    i_13_177_1769_0, i_13_177_1781_0, i_13_177_1805_0, i_13_177_1895_0,
    i_13_177_2021_0, i_13_177_2056_0, i_13_177_2111_0, i_13_177_2149_0,
    i_13_177_2284_0, i_13_177_2299_0, i_13_177_2300_0, i_13_177_2354_0,
    i_13_177_2572_0, i_13_177_2596_0, i_13_177_2597_0, i_13_177_2614_0,
    i_13_177_2615_0, i_13_177_2617_0, i_13_177_2665_0, i_13_177_2708_0,
    i_13_177_2782_0, i_13_177_2891_0, i_13_177_2900_0, i_13_177_2983_0,
    i_13_177_2987_0, i_13_177_3029_0, i_13_177_3032_0, i_13_177_3114_0,
    i_13_177_3130_0, i_13_177_3157_0, i_13_177_3215_0, i_13_177_3218_0,
    i_13_177_3287_0, i_13_177_3313_0, i_13_177_3355_0, i_13_177_3461_0,
    i_13_177_3467_0, i_13_177_3488_0, i_13_177_3521_0, i_13_177_3598_0,
    i_13_177_3687_0, i_13_177_3730_0, i_13_177_3757_0, i_13_177_3784_0,
    i_13_177_3875_0, i_13_177_3979_0, i_13_177_4055_0, i_13_177_4073_0,
    i_13_177_4088_0, i_13_177_4102_0, i_13_177_4162_0, i_13_177_4163_0,
    i_13_177_4228_0, i_13_177_4237_0, i_13_177_4268_0, i_13_177_4372_0,
    i_13_177_4448_0, i_13_177_4517_0, i_13_177_4559_0, i_13_177_4607_0;
  output o_13_177_0_0;
  assign o_13_177_0_0 = ~(~i_13_177_1151_0 | (~i_13_177_1411_0 & ~i_13_177_4372_0) | (~i_13_177_1768_0 & ~i_13_177_2983_0) | (~i_13_177_1412_0 & ~i_13_177_2111_0 & ~i_13_177_3218_0) | (~i_13_177_1769_0 & i_13_177_2983_0 & ~i_13_177_3784_0 & ~i_13_177_4162_0));
endmodule



// Benchmark "kernel_13_178" written by ABC on Sun Jul 19 10:47:53 2020

module kernel_13_178 ( 
    i_13_178_40_0, i_13_178_109_0, i_13_178_113_0, i_13_178_116_0,
    i_13_178_129_0, i_13_178_162_0, i_13_178_286_0, i_13_178_322_0,
    i_13_178_325_0, i_13_178_535_0, i_13_178_571_0, i_13_178_687_0,
    i_13_178_691_0, i_13_178_855_0, i_13_178_946_0, i_13_178_1012_0,
    i_13_178_1080_0, i_13_178_1081_0, i_13_178_1087_0, i_13_178_1120_0,
    i_13_178_1220_0, i_13_178_1395_0, i_13_178_1423_0, i_13_178_1424_0,
    i_13_178_1494_0, i_13_178_1569_0, i_13_178_1574_0, i_13_178_1629_0,
    i_13_178_1630_0, i_13_178_1632_0, i_13_178_1633_0, i_13_178_1634_0,
    i_13_178_1637_0, i_13_178_1773_0, i_13_178_1795_0, i_13_178_1938_0,
    i_13_178_1998_0, i_13_178_2059_0, i_13_178_2080_0, i_13_178_2081_0,
    i_13_178_2237_0, i_13_178_2342_0, i_13_178_2433_0, i_13_178_2438_0,
    i_13_178_2452_0, i_13_178_2462_0, i_13_178_2464_0, i_13_178_2498_0,
    i_13_178_2539_0, i_13_178_2541_0, i_13_178_2545_0, i_13_178_2546_0,
    i_13_178_2716_0, i_13_178_2905_0, i_13_178_2917_0, i_13_178_2920_0,
    i_13_178_2921_0, i_13_178_2955_0, i_13_178_3064_0, i_13_178_3065_0,
    i_13_178_3141_0, i_13_178_3143_0, i_13_178_3145_0, i_13_178_3146_0,
    i_13_178_3148_0, i_13_178_3338_0, i_13_178_3454_0, i_13_178_3455_0,
    i_13_178_3463_0, i_13_178_3464_0, i_13_178_3466_0, i_13_178_3688_0,
    i_13_178_3689_0, i_13_178_3727_0, i_13_178_3730_0, i_13_178_3734_0,
    i_13_178_3767_0, i_13_178_3770_0, i_13_178_3919_0, i_13_178_3968_0,
    i_13_178_3995_0, i_13_178_4018_0, i_13_178_4021_0, i_13_178_4022_0,
    i_13_178_4036_0, i_13_178_4049_0, i_13_178_4091_0, i_13_178_4253_0,
    i_13_178_4255_0, i_13_178_4256_0, i_13_178_4309_0, i_13_178_4354_0,
    i_13_178_4469_0, i_13_178_4513_0, i_13_178_4522_0, i_13_178_4523_0,
    i_13_178_4526_0, i_13_178_4558_0, i_13_178_4561_0, i_13_178_4562_0,
    o_13_178_0_0  );
  input  i_13_178_40_0, i_13_178_109_0, i_13_178_113_0, i_13_178_116_0,
    i_13_178_129_0, i_13_178_162_0, i_13_178_286_0, i_13_178_322_0,
    i_13_178_325_0, i_13_178_535_0, i_13_178_571_0, i_13_178_687_0,
    i_13_178_691_0, i_13_178_855_0, i_13_178_946_0, i_13_178_1012_0,
    i_13_178_1080_0, i_13_178_1081_0, i_13_178_1087_0, i_13_178_1120_0,
    i_13_178_1220_0, i_13_178_1395_0, i_13_178_1423_0, i_13_178_1424_0,
    i_13_178_1494_0, i_13_178_1569_0, i_13_178_1574_0, i_13_178_1629_0,
    i_13_178_1630_0, i_13_178_1632_0, i_13_178_1633_0, i_13_178_1634_0,
    i_13_178_1637_0, i_13_178_1773_0, i_13_178_1795_0, i_13_178_1938_0,
    i_13_178_1998_0, i_13_178_2059_0, i_13_178_2080_0, i_13_178_2081_0,
    i_13_178_2237_0, i_13_178_2342_0, i_13_178_2433_0, i_13_178_2438_0,
    i_13_178_2452_0, i_13_178_2462_0, i_13_178_2464_0, i_13_178_2498_0,
    i_13_178_2539_0, i_13_178_2541_0, i_13_178_2545_0, i_13_178_2546_0,
    i_13_178_2716_0, i_13_178_2905_0, i_13_178_2917_0, i_13_178_2920_0,
    i_13_178_2921_0, i_13_178_2955_0, i_13_178_3064_0, i_13_178_3065_0,
    i_13_178_3141_0, i_13_178_3143_0, i_13_178_3145_0, i_13_178_3146_0,
    i_13_178_3148_0, i_13_178_3338_0, i_13_178_3454_0, i_13_178_3455_0,
    i_13_178_3463_0, i_13_178_3464_0, i_13_178_3466_0, i_13_178_3688_0,
    i_13_178_3689_0, i_13_178_3727_0, i_13_178_3730_0, i_13_178_3734_0,
    i_13_178_3767_0, i_13_178_3770_0, i_13_178_3919_0, i_13_178_3968_0,
    i_13_178_3995_0, i_13_178_4018_0, i_13_178_4021_0, i_13_178_4022_0,
    i_13_178_4036_0, i_13_178_4049_0, i_13_178_4091_0, i_13_178_4253_0,
    i_13_178_4255_0, i_13_178_4256_0, i_13_178_4309_0, i_13_178_4354_0,
    i_13_178_4469_0, i_13_178_4513_0, i_13_178_4522_0, i_13_178_4523_0,
    i_13_178_4526_0, i_13_178_4558_0, i_13_178_4561_0, i_13_178_4562_0;
  output o_13_178_0_0;
  assign o_13_178_0_0 = ~((~i_13_178_3689_0 & ~i_13_178_4562_0) | (~i_13_178_3767_0 & ~i_13_178_3770_0));
endmodule



// Benchmark "kernel_13_179" written by ABC on Sun Jul 19 10:47:54 2020

module kernel_13_179 ( 
    i_13_179_31_0, i_13_179_79_0, i_13_179_111_0, i_13_179_112_0,
    i_13_179_114_0, i_13_179_166_0, i_13_179_168_0, i_13_179_169_0,
    i_13_179_229_0, i_13_179_318_0, i_13_179_327_0, i_13_179_490_0,
    i_13_179_525_0, i_13_179_526_0, i_13_179_564_0, i_13_179_643_0,
    i_13_179_822_0, i_13_179_850_0, i_13_179_858_0, i_13_179_862_0,
    i_13_179_924_0, i_13_179_940_0, i_13_179_960_0, i_13_179_1021_0,
    i_13_179_1075_0, i_13_179_1077_0, i_13_179_1200_0, i_13_179_1281_0,
    i_13_179_1419_0, i_13_179_1426_0, i_13_179_1428_0, i_13_179_1488_0,
    i_13_179_1498_0, i_13_179_1552_0, i_13_179_1632_0, i_13_179_1633_0,
    i_13_179_1642_0, i_13_179_1645_0, i_13_179_1704_0, i_13_179_1731_0,
    i_13_179_1831_0, i_13_179_1843_0, i_13_179_1950_0, i_13_179_1957_0,
    i_13_179_1986_0, i_13_179_2004_0, i_13_179_2026_0, i_13_179_2029_0,
    i_13_179_2193_0, i_13_179_2211_0, i_13_179_2271_0, i_13_179_2370_0,
    i_13_179_2452_0, i_13_179_2454_0, i_13_179_2455_0, i_13_179_2463_0,
    i_13_179_2541_0, i_13_179_2613_0, i_13_179_2707_0, i_13_179_2766_0,
    i_13_179_2778_0, i_13_179_2919_0, i_13_179_2920_0, i_13_179_2973_0,
    i_13_179_3030_0, i_13_179_3037_0, i_13_179_3090_0, i_13_179_3117_0,
    i_13_179_3148_0, i_13_179_3172_0, i_13_179_3180_0, i_13_179_3414_0,
    i_13_179_3453_0, i_13_179_3454_0, i_13_179_3459_0, i_13_179_3460_0,
    i_13_179_3462_0, i_13_179_3481_0, i_13_179_3483_0, i_13_179_3505_0,
    i_13_179_3540_0, i_13_179_3541_0, i_13_179_3561_0, i_13_179_3567_0,
    i_13_179_3574_0, i_13_179_3721_0, i_13_179_3867_0, i_13_179_3892_0,
    i_13_179_3936_0, i_13_179_4018_0, i_13_179_4063_0, i_13_179_4071_0,
    i_13_179_4164_0, i_13_179_4251_0, i_13_179_4255_0, i_13_179_4324_0,
    i_13_179_4341_0, i_13_179_4372_0, i_13_179_4378_0, i_13_179_4558_0,
    o_13_179_0_0  );
  input  i_13_179_31_0, i_13_179_79_0, i_13_179_111_0, i_13_179_112_0,
    i_13_179_114_0, i_13_179_166_0, i_13_179_168_0, i_13_179_169_0,
    i_13_179_229_0, i_13_179_318_0, i_13_179_327_0, i_13_179_490_0,
    i_13_179_525_0, i_13_179_526_0, i_13_179_564_0, i_13_179_643_0,
    i_13_179_822_0, i_13_179_850_0, i_13_179_858_0, i_13_179_862_0,
    i_13_179_924_0, i_13_179_940_0, i_13_179_960_0, i_13_179_1021_0,
    i_13_179_1075_0, i_13_179_1077_0, i_13_179_1200_0, i_13_179_1281_0,
    i_13_179_1419_0, i_13_179_1426_0, i_13_179_1428_0, i_13_179_1488_0,
    i_13_179_1498_0, i_13_179_1552_0, i_13_179_1632_0, i_13_179_1633_0,
    i_13_179_1642_0, i_13_179_1645_0, i_13_179_1704_0, i_13_179_1731_0,
    i_13_179_1831_0, i_13_179_1843_0, i_13_179_1950_0, i_13_179_1957_0,
    i_13_179_1986_0, i_13_179_2004_0, i_13_179_2026_0, i_13_179_2029_0,
    i_13_179_2193_0, i_13_179_2211_0, i_13_179_2271_0, i_13_179_2370_0,
    i_13_179_2452_0, i_13_179_2454_0, i_13_179_2455_0, i_13_179_2463_0,
    i_13_179_2541_0, i_13_179_2613_0, i_13_179_2707_0, i_13_179_2766_0,
    i_13_179_2778_0, i_13_179_2919_0, i_13_179_2920_0, i_13_179_2973_0,
    i_13_179_3030_0, i_13_179_3037_0, i_13_179_3090_0, i_13_179_3117_0,
    i_13_179_3148_0, i_13_179_3172_0, i_13_179_3180_0, i_13_179_3414_0,
    i_13_179_3453_0, i_13_179_3454_0, i_13_179_3459_0, i_13_179_3460_0,
    i_13_179_3462_0, i_13_179_3481_0, i_13_179_3483_0, i_13_179_3505_0,
    i_13_179_3540_0, i_13_179_3541_0, i_13_179_3561_0, i_13_179_3567_0,
    i_13_179_3574_0, i_13_179_3721_0, i_13_179_3867_0, i_13_179_3892_0,
    i_13_179_3936_0, i_13_179_4018_0, i_13_179_4063_0, i_13_179_4071_0,
    i_13_179_4164_0, i_13_179_4251_0, i_13_179_4255_0, i_13_179_4324_0,
    i_13_179_4341_0, i_13_179_4372_0, i_13_179_4378_0, i_13_179_4558_0;
  output o_13_179_0_0;
  assign o_13_179_0_0 = 0;
endmodule



// Benchmark "kernel_13_180" written by ABC on Sun Jul 19 10:47:55 2020

module kernel_13_180 ( 
    i_13_180_49_0, i_13_180_50_0, i_13_180_104_0, i_13_180_164_0,
    i_13_180_268_0, i_13_180_308_0, i_13_180_316_0, i_13_180_317_0,
    i_13_180_334_0, i_13_180_373_0, i_13_180_374_0, i_13_180_376_0,
    i_13_180_445_0, i_13_180_533_0, i_13_180_551_0, i_13_180_605_0,
    i_13_180_641_0, i_13_180_652_0, i_13_180_668_0, i_13_180_676_0,
    i_13_180_677_0, i_13_180_689_0, i_13_180_698_0, i_13_180_757_0,
    i_13_180_772_0, i_13_180_896_0, i_13_180_982_0, i_13_180_983_0,
    i_13_180_1121_0, i_13_180_1148_0, i_13_180_1250_0, i_13_180_1348_0,
    i_13_180_1412_0, i_13_180_1442_0, i_13_180_1516_0, i_13_180_1573_0,
    i_13_180_1648_0, i_13_180_1721_0, i_13_180_1750_0, i_13_180_1760_0,
    i_13_180_1789_0, i_13_180_1814_0, i_13_180_1832_0, i_13_180_1885_0,
    i_13_180_1909_0, i_13_180_1934_0, i_13_180_1957_0, i_13_180_2018_0,
    i_13_180_2032_0, i_13_180_2053_0, i_13_180_2113_0, i_13_180_2170_0,
    i_13_180_2281_0, i_13_180_2320_0, i_13_180_2348_0, i_13_180_2363_0,
    i_13_180_2468_0, i_13_180_2506_0, i_13_180_2507_0, i_13_180_2555_0,
    i_13_180_2716_0, i_13_180_2999_0, i_13_180_3047_0, i_13_180_3139_0,
    i_13_180_3215_0, i_13_180_3328_0, i_13_180_3352_0, i_13_180_3370_0,
    i_13_180_3376_0, i_13_180_3433_0, i_13_180_3437_0, i_13_180_3524_0,
    i_13_180_3533_0, i_13_180_3541_0, i_13_180_3565_0, i_13_180_3646_0,
    i_13_180_3686_0, i_13_180_3767_0, i_13_180_3865_0, i_13_180_3889_0,
    i_13_180_3890_0, i_13_180_3983_0, i_13_180_3988_0, i_13_180_4018_0,
    i_13_180_4019_0, i_13_180_4033_0, i_13_180_4046_0, i_13_180_4048_0,
    i_13_180_4079_0, i_13_180_4121_0, i_13_180_4124_0, i_13_180_4178_0,
    i_13_180_4447_0, i_13_180_4459_0, i_13_180_4471_0, i_13_180_4544_0,
    i_13_180_4591_0, i_13_180_4592_0, i_13_180_4600_0, i_13_180_4601_0,
    o_13_180_0_0  );
  input  i_13_180_49_0, i_13_180_50_0, i_13_180_104_0, i_13_180_164_0,
    i_13_180_268_0, i_13_180_308_0, i_13_180_316_0, i_13_180_317_0,
    i_13_180_334_0, i_13_180_373_0, i_13_180_374_0, i_13_180_376_0,
    i_13_180_445_0, i_13_180_533_0, i_13_180_551_0, i_13_180_605_0,
    i_13_180_641_0, i_13_180_652_0, i_13_180_668_0, i_13_180_676_0,
    i_13_180_677_0, i_13_180_689_0, i_13_180_698_0, i_13_180_757_0,
    i_13_180_772_0, i_13_180_896_0, i_13_180_982_0, i_13_180_983_0,
    i_13_180_1121_0, i_13_180_1148_0, i_13_180_1250_0, i_13_180_1348_0,
    i_13_180_1412_0, i_13_180_1442_0, i_13_180_1516_0, i_13_180_1573_0,
    i_13_180_1648_0, i_13_180_1721_0, i_13_180_1750_0, i_13_180_1760_0,
    i_13_180_1789_0, i_13_180_1814_0, i_13_180_1832_0, i_13_180_1885_0,
    i_13_180_1909_0, i_13_180_1934_0, i_13_180_1957_0, i_13_180_2018_0,
    i_13_180_2032_0, i_13_180_2053_0, i_13_180_2113_0, i_13_180_2170_0,
    i_13_180_2281_0, i_13_180_2320_0, i_13_180_2348_0, i_13_180_2363_0,
    i_13_180_2468_0, i_13_180_2506_0, i_13_180_2507_0, i_13_180_2555_0,
    i_13_180_2716_0, i_13_180_2999_0, i_13_180_3047_0, i_13_180_3139_0,
    i_13_180_3215_0, i_13_180_3328_0, i_13_180_3352_0, i_13_180_3370_0,
    i_13_180_3376_0, i_13_180_3433_0, i_13_180_3437_0, i_13_180_3524_0,
    i_13_180_3533_0, i_13_180_3541_0, i_13_180_3565_0, i_13_180_3646_0,
    i_13_180_3686_0, i_13_180_3767_0, i_13_180_3865_0, i_13_180_3889_0,
    i_13_180_3890_0, i_13_180_3983_0, i_13_180_3988_0, i_13_180_4018_0,
    i_13_180_4019_0, i_13_180_4033_0, i_13_180_4046_0, i_13_180_4048_0,
    i_13_180_4079_0, i_13_180_4121_0, i_13_180_4124_0, i_13_180_4178_0,
    i_13_180_4447_0, i_13_180_4459_0, i_13_180_4471_0, i_13_180_4544_0,
    i_13_180_4591_0, i_13_180_4592_0, i_13_180_4600_0, i_13_180_4601_0;
  output o_13_180_0_0;
  assign o_13_180_0_0 = ~(~i_13_180_689_0 | i_13_180_4048_0 | (~i_13_180_1814_0 & ~i_13_180_4079_0) | (i_13_180_1832_0 & ~i_13_180_1885_0 & ~i_13_180_4033_0) | (~i_13_180_676_0 & ~i_13_180_1412_0 & ~i_13_180_2113_0));
endmodule



// Benchmark "kernel_13_181" written by ABC on Sun Jul 19 10:47:56 2020

module kernel_13_181 ( 
    i_13_181_76_0, i_13_181_93_0, i_13_181_117_0, i_13_181_180_0,
    i_13_181_181_0, i_13_181_226_0, i_13_181_228_0, i_13_181_394_0,
    i_13_181_517_0, i_13_181_534_0, i_13_181_594_0, i_13_181_680_0,
    i_13_181_696_0, i_13_181_711_0, i_13_181_728_0, i_13_181_732_0,
    i_13_181_737_0, i_13_181_861_0, i_13_181_894_0, i_13_181_1075_0,
    i_13_181_1121_0, i_13_181_1207_0, i_13_181_1209_0, i_13_181_1252_0,
    i_13_181_1299_0, i_13_181_1408_0, i_13_181_1495_0, i_13_181_1507_0,
    i_13_181_1602_0, i_13_181_1632_0, i_13_181_1640_0, i_13_181_1700_0,
    i_13_181_1721_0, i_13_181_1723_0, i_13_181_1747_0, i_13_181_1782_0,
    i_13_181_1783_0, i_13_181_1785_0, i_13_181_1786_0, i_13_181_1921_0,
    i_13_181_1949_0, i_13_181_1955_0, i_13_181_1991_0, i_13_181_2055_0,
    i_13_181_2056_0, i_13_181_2096_0, i_13_181_2119_0, i_13_181_2182_0,
    i_13_181_2201_0, i_13_181_2204_0, i_13_181_2205_0, i_13_181_2208_0,
    i_13_181_2209_0, i_13_181_2235_0, i_13_181_2361_0, i_13_181_2452_0,
    i_13_181_2465_0, i_13_181_2560_0, i_13_181_2641_0, i_13_181_2789_0,
    i_13_181_2938_0, i_13_181_3019_0, i_13_181_3037_0, i_13_181_3062_0,
    i_13_181_3162_0, i_13_181_3163_0, i_13_181_3176_0, i_13_181_3204_0,
    i_13_181_3213_0, i_13_181_3285_0, i_13_181_3289_0, i_13_181_3353_0,
    i_13_181_3420_0, i_13_181_3423_0, i_13_181_3424_0, i_13_181_3531_0,
    i_13_181_3596_0, i_13_181_3620_0, i_13_181_3766_0, i_13_181_3782_0,
    i_13_181_3794_0, i_13_181_3870_0, i_13_181_3871_0, i_13_181_3981_0,
    i_13_181_4006_0, i_13_181_4008_0, i_13_181_4014_0, i_13_181_4022_0,
    i_13_181_4050_0, i_13_181_4058_0, i_13_181_4184_0, i_13_181_4214_0,
    i_13_181_4238_0, i_13_181_4261_0, i_13_181_4302_0, i_13_181_4397_0,
    i_13_181_4413_0, i_13_181_4451_0, i_13_181_4518_0, i_13_181_4540_0,
    o_13_181_0_0  );
  input  i_13_181_76_0, i_13_181_93_0, i_13_181_117_0, i_13_181_180_0,
    i_13_181_181_0, i_13_181_226_0, i_13_181_228_0, i_13_181_394_0,
    i_13_181_517_0, i_13_181_534_0, i_13_181_594_0, i_13_181_680_0,
    i_13_181_696_0, i_13_181_711_0, i_13_181_728_0, i_13_181_732_0,
    i_13_181_737_0, i_13_181_861_0, i_13_181_894_0, i_13_181_1075_0,
    i_13_181_1121_0, i_13_181_1207_0, i_13_181_1209_0, i_13_181_1252_0,
    i_13_181_1299_0, i_13_181_1408_0, i_13_181_1495_0, i_13_181_1507_0,
    i_13_181_1602_0, i_13_181_1632_0, i_13_181_1640_0, i_13_181_1700_0,
    i_13_181_1721_0, i_13_181_1723_0, i_13_181_1747_0, i_13_181_1782_0,
    i_13_181_1783_0, i_13_181_1785_0, i_13_181_1786_0, i_13_181_1921_0,
    i_13_181_1949_0, i_13_181_1955_0, i_13_181_1991_0, i_13_181_2055_0,
    i_13_181_2056_0, i_13_181_2096_0, i_13_181_2119_0, i_13_181_2182_0,
    i_13_181_2201_0, i_13_181_2204_0, i_13_181_2205_0, i_13_181_2208_0,
    i_13_181_2209_0, i_13_181_2235_0, i_13_181_2361_0, i_13_181_2452_0,
    i_13_181_2465_0, i_13_181_2560_0, i_13_181_2641_0, i_13_181_2789_0,
    i_13_181_2938_0, i_13_181_3019_0, i_13_181_3037_0, i_13_181_3062_0,
    i_13_181_3162_0, i_13_181_3163_0, i_13_181_3176_0, i_13_181_3204_0,
    i_13_181_3213_0, i_13_181_3285_0, i_13_181_3289_0, i_13_181_3353_0,
    i_13_181_3420_0, i_13_181_3423_0, i_13_181_3424_0, i_13_181_3531_0,
    i_13_181_3596_0, i_13_181_3620_0, i_13_181_3766_0, i_13_181_3782_0,
    i_13_181_3794_0, i_13_181_3870_0, i_13_181_3871_0, i_13_181_3981_0,
    i_13_181_4006_0, i_13_181_4008_0, i_13_181_4014_0, i_13_181_4022_0,
    i_13_181_4050_0, i_13_181_4058_0, i_13_181_4184_0, i_13_181_4214_0,
    i_13_181_4238_0, i_13_181_4261_0, i_13_181_4302_0, i_13_181_4397_0,
    i_13_181_4413_0, i_13_181_4451_0, i_13_181_4518_0, i_13_181_4540_0;
  output o_13_181_0_0;
  assign o_13_181_0_0 = ~((~i_13_181_3981_0 & (i_13_181_2452_0 | (~i_13_181_2208_0 & ~i_13_181_3163_0))) | (i_13_181_1075_0 & ~i_13_181_1299_0) | (~i_13_181_2209_0 & ~i_13_181_3870_0) | (~i_13_181_534_0 & ~i_13_181_2235_0 & ~i_13_181_4008_0 & ~i_13_181_4413_0));
endmodule



// Benchmark "kernel_13_182" written by ABC on Sun Jul 19 10:47:57 2020

module kernel_13_182 ( 
    i_13_182_45_0, i_13_182_48_0, i_13_182_76_0, i_13_182_94_0,
    i_13_182_247_0, i_13_182_411_0, i_13_182_450_0, i_13_182_534_0,
    i_13_182_556_0, i_13_182_601_0, i_13_182_625_0, i_13_182_626_0,
    i_13_182_660_0, i_13_182_661_0, i_13_182_812_0, i_13_182_834_0,
    i_13_182_835_0, i_13_182_850_0, i_13_182_909_0, i_13_182_940_0,
    i_13_182_1075_0, i_13_182_1147_0, i_13_182_1204_0, i_13_182_1227_0,
    i_13_182_1228_0, i_13_182_1230_0, i_13_182_1255_0, i_13_182_1271_0,
    i_13_182_1305_0, i_13_182_1314_0, i_13_182_1329_0, i_13_182_1345_0,
    i_13_182_1404_0, i_13_182_1463_0, i_13_182_1480_0, i_13_182_1497_0,
    i_13_182_1515_0, i_13_182_1522_0, i_13_182_1551_0, i_13_182_1647_0,
    i_13_182_1732_0, i_13_182_1744_0, i_13_182_1757_0, i_13_182_1767_0,
    i_13_182_1768_0, i_13_182_1803_0, i_13_182_1804_0, i_13_182_1884_0,
    i_13_182_1885_0, i_13_182_1944_0, i_13_182_1954_0, i_13_182_2001_0,
    i_13_182_2002_0, i_13_182_2100_0, i_13_182_2135_0, i_13_182_2145_0,
    i_13_182_2148_0, i_13_182_2199_0, i_13_182_2244_0, i_13_182_2469_0,
    i_13_182_2470_0, i_13_182_2472_0, i_13_182_2571_0, i_13_182_2625_0,
    i_13_182_2679_0, i_13_182_2854_0, i_13_182_2857_0, i_13_182_2896_0,
    i_13_182_2911_0, i_13_182_2968_0, i_13_182_2982_0, i_13_182_2985_0,
    i_13_182_3013_0, i_13_182_3031_0, i_13_182_3145_0, i_13_182_3258_0,
    i_13_182_3399_0, i_13_182_3423_0, i_13_182_3486_0, i_13_182_3549_0,
    i_13_182_3739_0, i_13_182_3803_0, i_13_182_3819_0, i_13_182_3850_0,
    i_13_182_3864_0, i_13_182_3868_0, i_13_182_3981_0, i_13_182_4126_0,
    i_13_182_4164_0, i_13_182_4252_0, i_13_182_4267_0, i_13_182_4269_0,
    i_13_182_4295_0, i_13_182_4369_0, i_13_182_4455_0, i_13_182_4467_0,
    i_13_182_4512_0, i_13_182_4513_0, i_13_182_4539_0, i_13_182_4566_0,
    o_13_182_0_0  );
  input  i_13_182_45_0, i_13_182_48_0, i_13_182_76_0, i_13_182_94_0,
    i_13_182_247_0, i_13_182_411_0, i_13_182_450_0, i_13_182_534_0,
    i_13_182_556_0, i_13_182_601_0, i_13_182_625_0, i_13_182_626_0,
    i_13_182_660_0, i_13_182_661_0, i_13_182_812_0, i_13_182_834_0,
    i_13_182_835_0, i_13_182_850_0, i_13_182_909_0, i_13_182_940_0,
    i_13_182_1075_0, i_13_182_1147_0, i_13_182_1204_0, i_13_182_1227_0,
    i_13_182_1228_0, i_13_182_1230_0, i_13_182_1255_0, i_13_182_1271_0,
    i_13_182_1305_0, i_13_182_1314_0, i_13_182_1329_0, i_13_182_1345_0,
    i_13_182_1404_0, i_13_182_1463_0, i_13_182_1480_0, i_13_182_1497_0,
    i_13_182_1515_0, i_13_182_1522_0, i_13_182_1551_0, i_13_182_1647_0,
    i_13_182_1732_0, i_13_182_1744_0, i_13_182_1757_0, i_13_182_1767_0,
    i_13_182_1768_0, i_13_182_1803_0, i_13_182_1804_0, i_13_182_1884_0,
    i_13_182_1885_0, i_13_182_1944_0, i_13_182_1954_0, i_13_182_2001_0,
    i_13_182_2002_0, i_13_182_2100_0, i_13_182_2135_0, i_13_182_2145_0,
    i_13_182_2148_0, i_13_182_2199_0, i_13_182_2244_0, i_13_182_2469_0,
    i_13_182_2470_0, i_13_182_2472_0, i_13_182_2571_0, i_13_182_2625_0,
    i_13_182_2679_0, i_13_182_2854_0, i_13_182_2857_0, i_13_182_2896_0,
    i_13_182_2911_0, i_13_182_2968_0, i_13_182_2982_0, i_13_182_2985_0,
    i_13_182_3013_0, i_13_182_3031_0, i_13_182_3145_0, i_13_182_3258_0,
    i_13_182_3399_0, i_13_182_3423_0, i_13_182_3486_0, i_13_182_3549_0,
    i_13_182_3739_0, i_13_182_3803_0, i_13_182_3819_0, i_13_182_3850_0,
    i_13_182_3864_0, i_13_182_3868_0, i_13_182_3981_0, i_13_182_4126_0,
    i_13_182_4164_0, i_13_182_4252_0, i_13_182_4267_0, i_13_182_4269_0,
    i_13_182_4295_0, i_13_182_4369_0, i_13_182_4455_0, i_13_182_4467_0,
    i_13_182_4512_0, i_13_182_4513_0, i_13_182_4539_0, i_13_182_4566_0;
  output o_13_182_0_0;
  assign o_13_182_0_0 = 0;
endmodule



// Benchmark "kernel_13_183" written by ABC on Sun Jul 19 10:47:57 2020

module kernel_13_183 ( 
    i_13_183_39_0, i_13_183_40_0, i_13_183_46_0, i_13_183_154_0,
    i_13_183_156_0, i_13_183_229_0, i_13_183_238_0, i_13_183_274_0,
    i_13_183_275_0, i_13_183_280_0, i_13_183_306_0, i_13_183_310_0,
    i_13_183_311_0, i_13_183_319_0, i_13_183_335_0, i_13_183_351_0,
    i_13_183_362_0, i_13_183_409_0, i_13_183_451_0, i_13_183_452_0,
    i_13_183_517_0, i_13_183_567_0, i_13_183_568_0, i_13_183_644_0,
    i_13_183_739_0, i_13_183_837_0, i_13_183_928_0, i_13_183_929_0,
    i_13_183_937_0, i_13_183_1082_0, i_13_183_1368_0, i_13_183_1432_0,
    i_13_183_1469_0, i_13_183_1496_0, i_13_183_1661_0, i_13_183_1765_0,
    i_13_183_1766_0, i_13_183_1829_0, i_13_183_1892_0, i_13_183_1945_0,
    i_13_183_2098_0, i_13_183_2227_0, i_13_183_2233_0, i_13_183_2234_0,
    i_13_183_2297_0, i_13_183_2434_0, i_13_183_2452_0, i_13_183_2542_0,
    i_13_183_2650_0, i_13_183_2677_0, i_13_183_2744_0, i_13_183_2746_0,
    i_13_183_2765_0, i_13_183_2767_0, i_13_183_2875_0, i_13_183_2981_0,
    i_13_183_3017_0, i_13_183_3029_0, i_13_183_3056_0, i_13_183_3107_0,
    i_13_183_3164_0, i_13_183_3214_0, i_13_183_3218_0, i_13_183_3232_0,
    i_13_183_3235_0, i_13_183_3286_0, i_13_183_3312_0, i_13_183_3313_0,
    i_13_183_3485_0, i_13_183_3487_0, i_13_183_3488_0, i_13_183_3523_0,
    i_13_183_3684_0, i_13_183_3698_0, i_13_183_3764_0, i_13_183_3766_0,
    i_13_183_3869_0, i_13_183_3898_0, i_13_183_3899_0, i_13_183_3901_0,
    i_13_183_4041_0, i_13_183_4063_0, i_13_183_4087_0, i_13_183_4088_0,
    i_13_183_4159_0, i_13_183_4162_0, i_13_183_4231_0, i_13_183_4250_0,
    i_13_183_4253_0, i_13_183_4267_0, i_13_183_4268_0, i_13_183_4270_0,
    i_13_183_4325_0, i_13_183_4359_0, i_13_183_4369_0, i_13_183_4370_0,
    i_13_183_4392_0, i_13_183_4447_0, i_13_183_4448_0, i_13_183_4559_0,
    o_13_183_0_0  );
  input  i_13_183_39_0, i_13_183_40_0, i_13_183_46_0, i_13_183_154_0,
    i_13_183_156_0, i_13_183_229_0, i_13_183_238_0, i_13_183_274_0,
    i_13_183_275_0, i_13_183_280_0, i_13_183_306_0, i_13_183_310_0,
    i_13_183_311_0, i_13_183_319_0, i_13_183_335_0, i_13_183_351_0,
    i_13_183_362_0, i_13_183_409_0, i_13_183_451_0, i_13_183_452_0,
    i_13_183_517_0, i_13_183_567_0, i_13_183_568_0, i_13_183_644_0,
    i_13_183_739_0, i_13_183_837_0, i_13_183_928_0, i_13_183_929_0,
    i_13_183_937_0, i_13_183_1082_0, i_13_183_1368_0, i_13_183_1432_0,
    i_13_183_1469_0, i_13_183_1496_0, i_13_183_1661_0, i_13_183_1765_0,
    i_13_183_1766_0, i_13_183_1829_0, i_13_183_1892_0, i_13_183_1945_0,
    i_13_183_2098_0, i_13_183_2227_0, i_13_183_2233_0, i_13_183_2234_0,
    i_13_183_2297_0, i_13_183_2434_0, i_13_183_2452_0, i_13_183_2542_0,
    i_13_183_2650_0, i_13_183_2677_0, i_13_183_2744_0, i_13_183_2746_0,
    i_13_183_2765_0, i_13_183_2767_0, i_13_183_2875_0, i_13_183_2981_0,
    i_13_183_3017_0, i_13_183_3029_0, i_13_183_3056_0, i_13_183_3107_0,
    i_13_183_3164_0, i_13_183_3214_0, i_13_183_3218_0, i_13_183_3232_0,
    i_13_183_3235_0, i_13_183_3286_0, i_13_183_3312_0, i_13_183_3313_0,
    i_13_183_3485_0, i_13_183_3487_0, i_13_183_3488_0, i_13_183_3523_0,
    i_13_183_3684_0, i_13_183_3698_0, i_13_183_3764_0, i_13_183_3766_0,
    i_13_183_3869_0, i_13_183_3898_0, i_13_183_3899_0, i_13_183_3901_0,
    i_13_183_4041_0, i_13_183_4063_0, i_13_183_4087_0, i_13_183_4088_0,
    i_13_183_4159_0, i_13_183_4162_0, i_13_183_4231_0, i_13_183_4250_0,
    i_13_183_4253_0, i_13_183_4267_0, i_13_183_4268_0, i_13_183_4270_0,
    i_13_183_4325_0, i_13_183_4359_0, i_13_183_4369_0, i_13_183_4370_0,
    i_13_183_4392_0, i_13_183_4447_0, i_13_183_4448_0, i_13_183_4559_0;
  output o_13_183_0_0;
  assign o_13_183_0_0 = ~((~i_13_183_3313_0 & ~i_13_183_4231_0) | (~i_13_183_46_0 & ~i_13_183_3901_0 & ~i_13_183_4369_0) | (i_13_183_229_0 & i_13_183_567_0 & ~i_13_183_3232_0) | (~i_13_183_2434_0 & ~i_13_183_3286_0 & ~i_13_183_4087_0 & ~i_13_183_4448_0) | (~i_13_183_928_0 & ~i_13_183_3898_0 & ~i_13_183_4088_0 & ~i_13_183_4267_0));
endmodule



// Benchmark "kernel_13_184" written by ABC on Sun Jul 19 10:47:58 2020

module kernel_13_184 ( 
    i_13_184_19_0, i_13_184_40_0, i_13_184_55_0, i_13_184_73_0,
    i_13_184_94_0, i_13_184_103_0, i_13_184_157_0, i_13_184_211_0,
    i_13_184_280_0, i_13_184_425_0, i_13_184_451_0, i_13_184_463_0,
    i_13_184_524_0, i_13_184_586_0, i_13_184_697_0, i_13_184_715_0,
    i_13_184_824_0, i_13_184_868_0, i_13_184_928_0, i_13_184_1017_0,
    i_13_184_1021_0, i_13_184_1066_0, i_13_184_1075_0, i_13_184_1204_0,
    i_13_184_1205_0, i_13_184_1207_0, i_13_184_1228_0, i_13_184_1274_0,
    i_13_184_1297_0, i_13_184_1342_0, i_13_184_1343_0, i_13_184_1405_0,
    i_13_184_1426_0, i_13_184_1427_0, i_13_184_1435_0, i_13_184_1468_0,
    i_13_184_1568_0, i_13_184_1634_0, i_13_184_1642_0, i_13_184_1711_0,
    i_13_184_1777_0, i_13_184_1811_0, i_13_184_1831_0, i_13_184_1882_0,
    i_13_184_1918_0, i_13_184_1940_0, i_13_184_1990_0, i_13_184_2004_0,
    i_13_184_2053_0, i_13_184_2110_0, i_13_184_2197_0, i_13_184_2236_0,
    i_13_184_2311_0, i_13_184_2362_0, i_13_184_2376_0, i_13_184_2452_0,
    i_13_184_2453_0, i_13_184_2504_0, i_13_184_2542_0, i_13_184_2549_0,
    i_13_184_2615_0, i_13_184_2710_0, i_13_184_2749_0, i_13_184_2854_0,
    i_13_184_2855_0, i_13_184_2912_0, i_13_184_2917_0, i_13_184_2918_0,
    i_13_184_3142_0, i_13_184_3143_0, i_13_184_3163_0, i_13_184_3208_0,
    i_13_184_3343_0, i_13_184_3441_0, i_13_184_3460_0, i_13_184_3467_0,
    i_13_184_3502_0, i_13_184_3503_0, i_13_184_3576_0, i_13_184_3637_0,
    i_13_184_3646_0, i_13_184_3764_0, i_13_184_3966_0, i_13_184_3982_0,
    i_13_184_4087_0, i_13_184_4088_0, i_13_184_4231_0, i_13_184_4258_0,
    i_13_184_4259_0, i_13_184_4392_0, i_13_184_4393_0, i_13_184_4394_0,
    i_13_184_4446_0, i_13_184_4447_0, i_13_184_4448_0, i_13_184_4511_0,
    i_13_184_4513_0, i_13_184_4555_0, i_13_184_4559_0, i_13_184_4564_0,
    o_13_184_0_0  );
  input  i_13_184_19_0, i_13_184_40_0, i_13_184_55_0, i_13_184_73_0,
    i_13_184_94_0, i_13_184_103_0, i_13_184_157_0, i_13_184_211_0,
    i_13_184_280_0, i_13_184_425_0, i_13_184_451_0, i_13_184_463_0,
    i_13_184_524_0, i_13_184_586_0, i_13_184_697_0, i_13_184_715_0,
    i_13_184_824_0, i_13_184_868_0, i_13_184_928_0, i_13_184_1017_0,
    i_13_184_1021_0, i_13_184_1066_0, i_13_184_1075_0, i_13_184_1204_0,
    i_13_184_1205_0, i_13_184_1207_0, i_13_184_1228_0, i_13_184_1274_0,
    i_13_184_1297_0, i_13_184_1342_0, i_13_184_1343_0, i_13_184_1405_0,
    i_13_184_1426_0, i_13_184_1427_0, i_13_184_1435_0, i_13_184_1468_0,
    i_13_184_1568_0, i_13_184_1634_0, i_13_184_1642_0, i_13_184_1711_0,
    i_13_184_1777_0, i_13_184_1811_0, i_13_184_1831_0, i_13_184_1882_0,
    i_13_184_1918_0, i_13_184_1940_0, i_13_184_1990_0, i_13_184_2004_0,
    i_13_184_2053_0, i_13_184_2110_0, i_13_184_2197_0, i_13_184_2236_0,
    i_13_184_2311_0, i_13_184_2362_0, i_13_184_2376_0, i_13_184_2452_0,
    i_13_184_2453_0, i_13_184_2504_0, i_13_184_2542_0, i_13_184_2549_0,
    i_13_184_2615_0, i_13_184_2710_0, i_13_184_2749_0, i_13_184_2854_0,
    i_13_184_2855_0, i_13_184_2912_0, i_13_184_2917_0, i_13_184_2918_0,
    i_13_184_3142_0, i_13_184_3143_0, i_13_184_3163_0, i_13_184_3208_0,
    i_13_184_3343_0, i_13_184_3441_0, i_13_184_3460_0, i_13_184_3467_0,
    i_13_184_3502_0, i_13_184_3503_0, i_13_184_3576_0, i_13_184_3637_0,
    i_13_184_3646_0, i_13_184_3764_0, i_13_184_3966_0, i_13_184_3982_0,
    i_13_184_4087_0, i_13_184_4088_0, i_13_184_4231_0, i_13_184_4258_0,
    i_13_184_4259_0, i_13_184_4392_0, i_13_184_4393_0, i_13_184_4394_0,
    i_13_184_4446_0, i_13_184_4447_0, i_13_184_4448_0, i_13_184_4511_0,
    i_13_184_4513_0, i_13_184_4555_0, i_13_184_4559_0, i_13_184_4564_0;
  output o_13_184_0_0;
  assign o_13_184_0_0 = ~((~i_13_184_4448_0 & ((~i_13_184_1274_0 & ~i_13_184_3646_0 & ~i_13_184_4258_0) | (~i_13_184_4088_0 & ~i_13_184_4393_0 & ~i_13_184_4555_0))) | (~i_13_184_1405_0 & ~i_13_184_1468_0 & i_13_184_1831_0) | (i_13_184_1468_0 & ~i_13_184_4231_0 & ~i_13_184_4259_0) | (~i_13_184_2855_0 & ~i_13_184_2918_0 & ~i_13_184_3460_0 & ~i_13_184_4394_0 & ~i_13_184_4446_0) | (i_13_184_1017_0 & ~i_13_184_1075_0 & i_13_184_4513_0));
endmodule



// Benchmark "kernel_13_185" written by ABC on Sun Jul 19 10:47:59 2020

module kernel_13_185 ( 
    i_13_185_27_0, i_13_185_49_0, i_13_185_64_0, i_13_185_67_0,
    i_13_185_120_0, i_13_185_121_0, i_13_185_192_0, i_13_185_193_0,
    i_13_185_201_0, i_13_185_225_0, i_13_185_270_0, i_13_185_324_0,
    i_13_185_378_0, i_13_185_379_0, i_13_185_441_0, i_13_185_507_0,
    i_13_185_553_0, i_13_185_570_0, i_13_185_571_0, i_13_185_576_0,
    i_13_185_694_0, i_13_185_697_0, i_13_185_714_0, i_13_185_715_0,
    i_13_185_717_0, i_13_185_768_0, i_13_185_858_0, i_13_185_948_0,
    i_13_185_1120_0, i_13_185_1200_0, i_13_185_1228_0, i_13_185_1372_0,
    i_13_185_1407_0, i_13_185_1426_0, i_13_185_1443_0, i_13_185_1467_0,
    i_13_185_1507_0, i_13_185_1516_0, i_13_185_1552_0, i_13_185_1623_0,
    i_13_185_1782_0, i_13_185_1783_0, i_13_185_1800_0, i_13_185_1801_0,
    i_13_185_1990_0, i_13_185_2011_0, i_13_185_2055_0, i_13_185_2056_0,
    i_13_185_2116_0, i_13_185_2128_0, i_13_185_2134_0, i_13_185_2206_0,
    i_13_185_2208_0, i_13_185_2209_0, i_13_185_2260_0, i_13_185_2358_0,
    i_13_185_2404_0, i_13_185_2424_0, i_13_185_2430_0, i_13_185_2452_0,
    i_13_185_2532_0, i_13_185_2589_0, i_13_185_2593_0, i_13_185_2710_0,
    i_13_185_2718_0, i_13_185_2934_0, i_13_185_2935_0, i_13_185_3015_0,
    i_13_185_3016_0, i_13_185_3151_0, i_13_185_3171_0, i_13_185_3208_0,
    i_13_185_3214_0, i_13_185_3241_0, i_13_185_3258_0, i_13_185_3267_0,
    i_13_185_3286_0, i_13_185_3342_0, i_13_185_3415_0, i_13_185_3420_0,
    i_13_185_3421_0, i_13_185_3423_0, i_13_185_3424_0, i_13_185_3532_0,
    i_13_185_3610_0, i_13_185_3846_0, i_13_185_3847_0, i_13_185_3871_0,
    i_13_185_3873_0, i_13_185_3874_0, i_13_185_3981_0, i_13_185_4009_0,
    i_13_185_4050_0, i_13_185_4051_0, i_13_185_4123_0, i_13_185_4150_0,
    i_13_185_4188_0, i_13_185_4404_0, i_13_185_4410_0, i_13_185_4594_0,
    o_13_185_0_0  );
  input  i_13_185_27_0, i_13_185_49_0, i_13_185_64_0, i_13_185_67_0,
    i_13_185_120_0, i_13_185_121_0, i_13_185_192_0, i_13_185_193_0,
    i_13_185_201_0, i_13_185_225_0, i_13_185_270_0, i_13_185_324_0,
    i_13_185_378_0, i_13_185_379_0, i_13_185_441_0, i_13_185_507_0,
    i_13_185_553_0, i_13_185_570_0, i_13_185_571_0, i_13_185_576_0,
    i_13_185_694_0, i_13_185_697_0, i_13_185_714_0, i_13_185_715_0,
    i_13_185_717_0, i_13_185_768_0, i_13_185_858_0, i_13_185_948_0,
    i_13_185_1120_0, i_13_185_1200_0, i_13_185_1228_0, i_13_185_1372_0,
    i_13_185_1407_0, i_13_185_1426_0, i_13_185_1443_0, i_13_185_1467_0,
    i_13_185_1507_0, i_13_185_1516_0, i_13_185_1552_0, i_13_185_1623_0,
    i_13_185_1782_0, i_13_185_1783_0, i_13_185_1800_0, i_13_185_1801_0,
    i_13_185_1990_0, i_13_185_2011_0, i_13_185_2055_0, i_13_185_2056_0,
    i_13_185_2116_0, i_13_185_2128_0, i_13_185_2134_0, i_13_185_2206_0,
    i_13_185_2208_0, i_13_185_2209_0, i_13_185_2260_0, i_13_185_2358_0,
    i_13_185_2404_0, i_13_185_2424_0, i_13_185_2430_0, i_13_185_2452_0,
    i_13_185_2532_0, i_13_185_2589_0, i_13_185_2593_0, i_13_185_2710_0,
    i_13_185_2718_0, i_13_185_2934_0, i_13_185_2935_0, i_13_185_3015_0,
    i_13_185_3016_0, i_13_185_3151_0, i_13_185_3171_0, i_13_185_3208_0,
    i_13_185_3214_0, i_13_185_3241_0, i_13_185_3258_0, i_13_185_3267_0,
    i_13_185_3286_0, i_13_185_3342_0, i_13_185_3415_0, i_13_185_3420_0,
    i_13_185_3421_0, i_13_185_3423_0, i_13_185_3424_0, i_13_185_3532_0,
    i_13_185_3610_0, i_13_185_3846_0, i_13_185_3847_0, i_13_185_3871_0,
    i_13_185_3873_0, i_13_185_3874_0, i_13_185_3981_0, i_13_185_4009_0,
    i_13_185_4050_0, i_13_185_4051_0, i_13_185_4123_0, i_13_185_4150_0,
    i_13_185_4188_0, i_13_185_4404_0, i_13_185_4410_0, i_13_185_4594_0;
  output o_13_185_0_0;
  assign o_13_185_0_0 = ~((~i_13_185_1407_0 & ((i_13_185_1507_0 & ~i_13_185_1800_0 & ~i_13_185_2424_0) | (i_13_185_2056_0 & ~i_13_185_3420_0) | (i_13_185_697_0 & ~i_13_185_2710_0 & ~i_13_185_3214_0 & ~i_13_185_3981_0))) | (~i_13_185_2935_0 & ~i_13_185_3423_0 & ~i_13_185_3846_0) | (~i_13_185_120_0 & ~i_13_185_2430_0 & ~i_13_185_3874_0 & ~i_13_185_4050_0));
endmodule



// Benchmark "kernel_13_186" written by ABC on Sun Jul 19 10:48:00 2020

module kernel_13_186 ( 
    i_13_186_78_0, i_13_186_96_0, i_13_186_106_0, i_13_186_327_0,
    i_13_186_529_0, i_13_186_598_0, i_13_186_627_0, i_13_186_672_0,
    i_13_186_673_0, i_13_186_717_0, i_13_186_727_0, i_13_186_780_0,
    i_13_186_781_0, i_13_186_815_0, i_13_186_825_0, i_13_186_841_0,
    i_13_186_850_0, i_13_186_894_0, i_13_186_949_0, i_13_186_979_0,
    i_13_186_1095_0, i_13_186_1141_0, i_13_186_1259_0, i_13_186_1302_0,
    i_13_186_1303_0, i_13_186_1320_0, i_13_186_1327_0, i_13_186_1383_0,
    i_13_186_1464_0, i_13_186_1465_0, i_13_186_1466_0, i_13_186_1482_0,
    i_13_186_1483_0, i_13_186_1484_0, i_13_186_1643_0, i_13_186_1751_0,
    i_13_186_1759_0, i_13_186_1789_0, i_13_186_1806_0, i_13_186_1807_0,
    i_13_186_1808_0, i_13_186_1815_0, i_13_186_1885_0, i_13_186_1887_0,
    i_13_186_1905_0, i_13_186_1906_0, i_13_186_2033_0, i_13_186_2122_0,
    i_13_186_2123_0, i_13_186_2139_0, i_13_186_2140_0, i_13_186_2167_0,
    i_13_186_2177_0, i_13_186_2247_0, i_13_186_2310_0, i_13_186_2380_0,
    i_13_186_2445_0, i_13_186_2446_0, i_13_186_2470_0, i_13_186_2474_0,
    i_13_186_2652_0, i_13_186_2698_0, i_13_186_2751_0, i_13_186_2823_0,
    i_13_186_2824_0, i_13_186_2861_0, i_13_186_3009_0, i_13_186_3112_0,
    i_13_186_3174_0, i_13_186_3219_0, i_13_186_3220_0, i_13_186_3293_0,
    i_13_186_3391_0, i_13_186_3398_0, i_13_186_3432_0, i_13_186_3451_0,
    i_13_186_3452_0, i_13_186_3564_0, i_13_186_3577_0, i_13_186_3579_0,
    i_13_186_3734_0, i_13_186_3793_0, i_13_186_3820_0, i_13_186_3855_0,
    i_13_186_3874_0, i_13_186_3883_0, i_13_186_3927_0, i_13_186_3929_0,
    i_13_186_3991_0, i_13_186_3992_0, i_13_186_4049_0, i_13_186_4237_0,
    i_13_186_4308_0, i_13_186_4318_0, i_13_186_4365_0, i_13_186_4380_0,
    i_13_186_4414_0, i_13_186_4443_0, i_13_186_4453_0, i_13_186_4521_0,
    o_13_186_0_0  );
  input  i_13_186_78_0, i_13_186_96_0, i_13_186_106_0, i_13_186_327_0,
    i_13_186_529_0, i_13_186_598_0, i_13_186_627_0, i_13_186_672_0,
    i_13_186_673_0, i_13_186_717_0, i_13_186_727_0, i_13_186_780_0,
    i_13_186_781_0, i_13_186_815_0, i_13_186_825_0, i_13_186_841_0,
    i_13_186_850_0, i_13_186_894_0, i_13_186_949_0, i_13_186_979_0,
    i_13_186_1095_0, i_13_186_1141_0, i_13_186_1259_0, i_13_186_1302_0,
    i_13_186_1303_0, i_13_186_1320_0, i_13_186_1327_0, i_13_186_1383_0,
    i_13_186_1464_0, i_13_186_1465_0, i_13_186_1466_0, i_13_186_1482_0,
    i_13_186_1483_0, i_13_186_1484_0, i_13_186_1643_0, i_13_186_1751_0,
    i_13_186_1759_0, i_13_186_1789_0, i_13_186_1806_0, i_13_186_1807_0,
    i_13_186_1808_0, i_13_186_1815_0, i_13_186_1885_0, i_13_186_1887_0,
    i_13_186_1905_0, i_13_186_1906_0, i_13_186_2033_0, i_13_186_2122_0,
    i_13_186_2123_0, i_13_186_2139_0, i_13_186_2140_0, i_13_186_2167_0,
    i_13_186_2177_0, i_13_186_2247_0, i_13_186_2310_0, i_13_186_2380_0,
    i_13_186_2445_0, i_13_186_2446_0, i_13_186_2470_0, i_13_186_2474_0,
    i_13_186_2652_0, i_13_186_2698_0, i_13_186_2751_0, i_13_186_2823_0,
    i_13_186_2824_0, i_13_186_2861_0, i_13_186_3009_0, i_13_186_3112_0,
    i_13_186_3174_0, i_13_186_3219_0, i_13_186_3220_0, i_13_186_3293_0,
    i_13_186_3391_0, i_13_186_3398_0, i_13_186_3432_0, i_13_186_3451_0,
    i_13_186_3452_0, i_13_186_3564_0, i_13_186_3577_0, i_13_186_3579_0,
    i_13_186_3734_0, i_13_186_3793_0, i_13_186_3820_0, i_13_186_3855_0,
    i_13_186_3874_0, i_13_186_3883_0, i_13_186_3927_0, i_13_186_3929_0,
    i_13_186_3991_0, i_13_186_3992_0, i_13_186_4049_0, i_13_186_4237_0,
    i_13_186_4308_0, i_13_186_4318_0, i_13_186_4365_0, i_13_186_4380_0,
    i_13_186_4414_0, i_13_186_4443_0, i_13_186_4453_0, i_13_186_4521_0;
  output o_13_186_0_0;
  assign o_13_186_0_0 = ~((~i_13_186_2446_0 & ~i_13_186_4453_0) | (i_13_186_3112_0 & i_13_186_3452_0) | (i_13_186_673_0 & ~i_13_186_3220_0 & ~i_13_186_3734_0 & ~i_13_186_3927_0));
endmodule



// Benchmark "kernel_13_187" written by ABC on Sun Jul 19 10:48:01 2020

module kernel_13_187 ( 
    i_13_187_31_0, i_13_187_101_0, i_13_187_235_0, i_13_187_238_0,
    i_13_187_248_0, i_13_187_251_0, i_13_187_256_0, i_13_187_263_0,
    i_13_187_275_0, i_13_187_278_0, i_13_187_338_0, i_13_187_407_0,
    i_13_187_411_0, i_13_187_447_0, i_13_187_451_0, i_13_187_485_0,
    i_13_187_535_0, i_13_187_559_0, i_13_187_563_0, i_13_187_577_0,
    i_13_187_578_0, i_13_187_616_0, i_13_187_619_0, i_13_187_620_0,
    i_13_187_644_0, i_13_187_793_0, i_13_187_813_0, i_13_187_832_0,
    i_13_187_841_0, i_13_187_941_0, i_13_187_942_0, i_13_187_977_0,
    i_13_187_979_0, i_13_187_1095_0, i_13_187_1112_0, i_13_187_1262_0,
    i_13_187_1333_0, i_13_187_1342_0, i_13_187_1396_0, i_13_187_1397_0,
    i_13_187_1477_0, i_13_187_1494_0, i_13_187_1541_0, i_13_187_1570_0,
    i_13_187_1647_0, i_13_187_1658_0, i_13_187_1722_0, i_13_187_1729_0,
    i_13_187_1814_0, i_13_187_1835_0, i_13_187_1842_0, i_13_187_1858_0,
    i_13_187_1920_0, i_13_187_1947_0, i_13_187_2106_0, i_13_187_2108_0,
    i_13_187_2113_0, i_13_187_2230_0, i_13_187_2233_0, i_13_187_2261_0,
    i_13_187_2280_0, i_13_187_2445_0, i_13_187_2713_0, i_13_187_2721_0,
    i_13_187_2737_0, i_13_187_2740_0, i_13_187_2765_0, i_13_187_2785_0,
    i_13_187_2888_0, i_13_187_2951_0, i_13_187_3018_0, i_13_187_3056_0,
    i_13_187_3115_0, i_13_187_3135_0, i_13_187_3152_0, i_13_187_3208_0,
    i_13_187_3217_0, i_13_187_3218_0, i_13_187_3313_0, i_13_187_3316_0,
    i_13_187_3403_0, i_13_187_3412_0, i_13_187_3435_0, i_13_187_3461_0,
    i_13_187_3601_0, i_13_187_3602_0, i_13_187_3616_0, i_13_187_3617_0,
    i_13_187_3709_0, i_13_187_3764_0, i_13_187_3858_0, i_13_187_3901_0,
    i_13_187_3902_0, i_13_187_4124_0, i_13_187_4178_0, i_13_187_4207_0,
    i_13_187_4268_0, i_13_187_4360_0, i_13_187_4391_0, i_13_187_4483_0,
    o_13_187_0_0  );
  input  i_13_187_31_0, i_13_187_101_0, i_13_187_235_0, i_13_187_238_0,
    i_13_187_248_0, i_13_187_251_0, i_13_187_256_0, i_13_187_263_0,
    i_13_187_275_0, i_13_187_278_0, i_13_187_338_0, i_13_187_407_0,
    i_13_187_411_0, i_13_187_447_0, i_13_187_451_0, i_13_187_485_0,
    i_13_187_535_0, i_13_187_559_0, i_13_187_563_0, i_13_187_577_0,
    i_13_187_578_0, i_13_187_616_0, i_13_187_619_0, i_13_187_620_0,
    i_13_187_644_0, i_13_187_793_0, i_13_187_813_0, i_13_187_832_0,
    i_13_187_841_0, i_13_187_941_0, i_13_187_942_0, i_13_187_977_0,
    i_13_187_979_0, i_13_187_1095_0, i_13_187_1112_0, i_13_187_1262_0,
    i_13_187_1333_0, i_13_187_1342_0, i_13_187_1396_0, i_13_187_1397_0,
    i_13_187_1477_0, i_13_187_1494_0, i_13_187_1541_0, i_13_187_1570_0,
    i_13_187_1647_0, i_13_187_1658_0, i_13_187_1722_0, i_13_187_1729_0,
    i_13_187_1814_0, i_13_187_1835_0, i_13_187_1842_0, i_13_187_1858_0,
    i_13_187_1920_0, i_13_187_1947_0, i_13_187_2106_0, i_13_187_2108_0,
    i_13_187_2113_0, i_13_187_2230_0, i_13_187_2233_0, i_13_187_2261_0,
    i_13_187_2280_0, i_13_187_2445_0, i_13_187_2713_0, i_13_187_2721_0,
    i_13_187_2737_0, i_13_187_2740_0, i_13_187_2765_0, i_13_187_2785_0,
    i_13_187_2888_0, i_13_187_2951_0, i_13_187_3018_0, i_13_187_3056_0,
    i_13_187_3115_0, i_13_187_3135_0, i_13_187_3152_0, i_13_187_3208_0,
    i_13_187_3217_0, i_13_187_3218_0, i_13_187_3313_0, i_13_187_3316_0,
    i_13_187_3403_0, i_13_187_3412_0, i_13_187_3435_0, i_13_187_3461_0,
    i_13_187_3601_0, i_13_187_3602_0, i_13_187_3616_0, i_13_187_3617_0,
    i_13_187_3709_0, i_13_187_3764_0, i_13_187_3858_0, i_13_187_3901_0,
    i_13_187_3902_0, i_13_187_4124_0, i_13_187_4178_0, i_13_187_4207_0,
    i_13_187_4268_0, i_13_187_4360_0, i_13_187_4391_0, i_13_187_4483_0;
  output o_13_187_0_0;
  assign o_13_187_0_0 = ~((~i_13_187_275_0 & ~i_13_187_3901_0) | (~i_13_187_1397_0 & ~i_13_187_3602_0));
endmodule



// Benchmark "kernel_13_188" written by ABC on Sun Jul 19 10:48:02 2020

module kernel_13_188 ( 
    i_13_188_44_0, i_13_188_91_0, i_13_188_98_0, i_13_188_175_0,
    i_13_188_176_0, i_13_188_179_0, i_13_188_181_0, i_13_188_229_0,
    i_13_188_280_0, i_13_188_283_0, i_13_188_308_0, i_13_188_309_0,
    i_13_188_313_0, i_13_188_314_0, i_13_188_317_0, i_13_188_320_0,
    i_13_188_549_0, i_13_188_554_0, i_13_188_571_0, i_13_188_657_0,
    i_13_188_697_0, i_13_188_710_0, i_13_188_758_0, i_13_188_846_0,
    i_13_188_847_0, i_13_188_855_0, i_13_188_981_0, i_13_188_985_0,
    i_13_188_986_0, i_13_188_1105_0, i_13_188_1106_0, i_13_188_1260_0,
    i_13_188_1327_0, i_13_188_1471_0, i_13_188_1486_0, i_13_188_1511_0,
    i_13_188_1532_0, i_13_188_1714_0, i_13_188_1799_0, i_13_188_1832_0,
    i_13_188_1852_0, i_13_188_1853_0, i_13_188_1858_0, i_13_188_1859_0,
    i_13_188_1861_0, i_13_188_1996_0, i_13_188_2096_0, i_13_188_2406_0,
    i_13_188_2411_0, i_13_188_2447_0, i_13_188_2452_0, i_13_188_2460_0,
    i_13_188_2473_0, i_13_188_2475_0, i_13_188_2565_0, i_13_188_2676_0,
    i_13_188_2699_0, i_13_188_2798_0, i_13_188_2849_0, i_13_188_2983_0,
    i_13_188_3006_0, i_13_188_3008_0, i_13_188_3009_0, i_13_188_3032_0,
    i_13_188_3061_0, i_13_188_3108_0, i_13_188_3109_0, i_13_188_3112_0,
    i_13_188_3141_0, i_13_188_3204_0, i_13_188_3205_0, i_13_188_3208_0,
    i_13_188_3211_0, i_13_188_3212_0, i_13_188_3335_0, i_13_188_3343_0,
    i_13_188_3382_0, i_13_188_3397_0, i_13_188_3405_0, i_13_188_3765_0,
    i_13_188_3766_0, i_13_188_3816_0, i_13_188_3817_0, i_13_188_3818_0,
    i_13_188_3823_0, i_13_188_3865_0, i_13_188_3866_0, i_13_188_3910_0,
    i_13_188_4043_0, i_13_188_4063_0, i_13_188_4067_0, i_13_188_4084_0,
    i_13_188_4085_0, i_13_188_4304_0, i_13_188_4350_0, i_13_188_4379_0,
    i_13_188_4414_0, i_13_188_4522_0, i_13_188_4581_0, i_13_188_4598_0,
    o_13_188_0_0  );
  input  i_13_188_44_0, i_13_188_91_0, i_13_188_98_0, i_13_188_175_0,
    i_13_188_176_0, i_13_188_179_0, i_13_188_181_0, i_13_188_229_0,
    i_13_188_280_0, i_13_188_283_0, i_13_188_308_0, i_13_188_309_0,
    i_13_188_313_0, i_13_188_314_0, i_13_188_317_0, i_13_188_320_0,
    i_13_188_549_0, i_13_188_554_0, i_13_188_571_0, i_13_188_657_0,
    i_13_188_697_0, i_13_188_710_0, i_13_188_758_0, i_13_188_846_0,
    i_13_188_847_0, i_13_188_855_0, i_13_188_981_0, i_13_188_985_0,
    i_13_188_986_0, i_13_188_1105_0, i_13_188_1106_0, i_13_188_1260_0,
    i_13_188_1327_0, i_13_188_1471_0, i_13_188_1486_0, i_13_188_1511_0,
    i_13_188_1532_0, i_13_188_1714_0, i_13_188_1799_0, i_13_188_1832_0,
    i_13_188_1852_0, i_13_188_1853_0, i_13_188_1858_0, i_13_188_1859_0,
    i_13_188_1861_0, i_13_188_1996_0, i_13_188_2096_0, i_13_188_2406_0,
    i_13_188_2411_0, i_13_188_2447_0, i_13_188_2452_0, i_13_188_2460_0,
    i_13_188_2473_0, i_13_188_2475_0, i_13_188_2565_0, i_13_188_2676_0,
    i_13_188_2699_0, i_13_188_2798_0, i_13_188_2849_0, i_13_188_2983_0,
    i_13_188_3006_0, i_13_188_3008_0, i_13_188_3009_0, i_13_188_3032_0,
    i_13_188_3061_0, i_13_188_3108_0, i_13_188_3109_0, i_13_188_3112_0,
    i_13_188_3141_0, i_13_188_3204_0, i_13_188_3205_0, i_13_188_3208_0,
    i_13_188_3211_0, i_13_188_3212_0, i_13_188_3335_0, i_13_188_3343_0,
    i_13_188_3382_0, i_13_188_3397_0, i_13_188_3405_0, i_13_188_3765_0,
    i_13_188_3766_0, i_13_188_3816_0, i_13_188_3817_0, i_13_188_3818_0,
    i_13_188_3823_0, i_13_188_3865_0, i_13_188_3866_0, i_13_188_3910_0,
    i_13_188_4043_0, i_13_188_4063_0, i_13_188_4067_0, i_13_188_4084_0,
    i_13_188_4085_0, i_13_188_4304_0, i_13_188_4350_0, i_13_188_4379_0,
    i_13_188_4414_0, i_13_188_4522_0, i_13_188_4581_0, i_13_188_4598_0;
  output o_13_188_0_0;
  assign o_13_188_0_0 = ~(i_13_188_4304_0 | (~i_13_188_1486_0 & ~i_13_188_4085_0) | (~i_13_188_3817_0 & ~i_13_188_3823_0 & ~i_13_188_4067_0) | (~i_13_188_1799_0 & ~i_13_188_2411_0 & ~i_13_188_3008_0));
endmodule



// Benchmark "kernel_13_189" written by ABC on Sun Jul 19 10:48:03 2020

module kernel_13_189 ( 
    i_13_189_29_0, i_13_189_36_0, i_13_189_37_0, i_13_189_46_0,
    i_13_189_64_0, i_13_189_121_0, i_13_189_136_0, i_13_189_311_0,
    i_13_189_334_0, i_13_189_370_0, i_13_189_412_0, i_13_189_414_0,
    i_13_189_415_0, i_13_189_585_0, i_13_189_612_0, i_13_189_613_0,
    i_13_189_654_0, i_13_189_684_0, i_13_189_685_0, i_13_189_693_0,
    i_13_189_694_0, i_13_189_760_0, i_13_189_837_0, i_13_189_838_0,
    i_13_189_841_0, i_13_189_889_0, i_13_189_955_0, i_13_189_1071_0,
    i_13_189_1072_0, i_13_189_1081_0, i_13_189_1117_0, i_13_189_1121_0,
    i_13_189_1270_0, i_13_189_1285_0, i_13_189_1299_0, i_13_189_1317_0,
    i_13_189_1360_0, i_13_189_1390_0, i_13_189_1516_0, i_13_189_1521_0,
    i_13_189_1522_0, i_13_189_1534_0, i_13_189_1633_0, i_13_189_1639_0,
    i_13_189_1668_0, i_13_189_1750_0, i_13_189_1756_0, i_13_189_1792_0,
    i_13_189_1885_0, i_13_189_1914_0, i_13_189_2125_0, i_13_189_2191_0,
    i_13_189_2244_0, i_13_189_2379_0, i_13_189_2380_0, i_13_189_2434_0,
    i_13_189_2457_0, i_13_189_2541_0, i_13_189_2646_0, i_13_189_2647_0,
    i_13_189_2650_0, i_13_189_2820_0, i_13_189_2821_0, i_13_189_2847_0,
    i_13_189_2848_0, i_13_189_3091_0, i_13_189_3109_0, i_13_189_3269_0,
    i_13_189_3306_0, i_13_189_3307_0, i_13_189_3372_0, i_13_189_3387_0,
    i_13_189_3388_0, i_13_189_3429_0, i_13_189_3451_0, i_13_189_3538_0,
    i_13_189_3547_0, i_13_189_3555_0, i_13_189_3636_0, i_13_189_3637_0,
    i_13_189_3766_0, i_13_189_3836_0, i_13_189_3889_0, i_13_189_3906_0,
    i_13_189_3910_0, i_13_189_3934_0, i_13_189_3936_0, i_13_189_3988_0,
    i_13_189_4017_0, i_13_189_4032_0, i_13_189_4033_0, i_13_189_4036_0,
    i_13_189_4164_0, i_13_189_4269_0, i_13_189_4294_0, i_13_189_4327_0,
    i_13_189_4378_0, i_13_189_4396_0, i_13_189_4510_0, i_13_189_4593_0,
    o_13_189_0_0  );
  input  i_13_189_29_0, i_13_189_36_0, i_13_189_37_0, i_13_189_46_0,
    i_13_189_64_0, i_13_189_121_0, i_13_189_136_0, i_13_189_311_0,
    i_13_189_334_0, i_13_189_370_0, i_13_189_412_0, i_13_189_414_0,
    i_13_189_415_0, i_13_189_585_0, i_13_189_612_0, i_13_189_613_0,
    i_13_189_654_0, i_13_189_684_0, i_13_189_685_0, i_13_189_693_0,
    i_13_189_694_0, i_13_189_760_0, i_13_189_837_0, i_13_189_838_0,
    i_13_189_841_0, i_13_189_889_0, i_13_189_955_0, i_13_189_1071_0,
    i_13_189_1072_0, i_13_189_1081_0, i_13_189_1117_0, i_13_189_1121_0,
    i_13_189_1270_0, i_13_189_1285_0, i_13_189_1299_0, i_13_189_1317_0,
    i_13_189_1360_0, i_13_189_1390_0, i_13_189_1516_0, i_13_189_1521_0,
    i_13_189_1522_0, i_13_189_1534_0, i_13_189_1633_0, i_13_189_1639_0,
    i_13_189_1668_0, i_13_189_1750_0, i_13_189_1756_0, i_13_189_1792_0,
    i_13_189_1885_0, i_13_189_1914_0, i_13_189_2125_0, i_13_189_2191_0,
    i_13_189_2244_0, i_13_189_2379_0, i_13_189_2380_0, i_13_189_2434_0,
    i_13_189_2457_0, i_13_189_2541_0, i_13_189_2646_0, i_13_189_2647_0,
    i_13_189_2650_0, i_13_189_2820_0, i_13_189_2821_0, i_13_189_2847_0,
    i_13_189_2848_0, i_13_189_3091_0, i_13_189_3109_0, i_13_189_3269_0,
    i_13_189_3306_0, i_13_189_3307_0, i_13_189_3372_0, i_13_189_3387_0,
    i_13_189_3388_0, i_13_189_3429_0, i_13_189_3451_0, i_13_189_3538_0,
    i_13_189_3547_0, i_13_189_3555_0, i_13_189_3636_0, i_13_189_3637_0,
    i_13_189_3766_0, i_13_189_3836_0, i_13_189_3889_0, i_13_189_3906_0,
    i_13_189_3910_0, i_13_189_3934_0, i_13_189_3936_0, i_13_189_3988_0,
    i_13_189_4017_0, i_13_189_4032_0, i_13_189_4033_0, i_13_189_4036_0,
    i_13_189_4164_0, i_13_189_4269_0, i_13_189_4294_0, i_13_189_4327_0,
    i_13_189_4378_0, i_13_189_4396_0, i_13_189_4510_0, i_13_189_4593_0;
  output o_13_189_0_0;
  assign o_13_189_0_0 = ~((~i_13_189_46_0 & ((i_13_189_685_0 & ~i_13_189_1792_0 & ~i_13_189_3906_0) | (~i_13_189_334_0 & ~i_13_189_4032_0))) | (~i_13_189_2646_0 & (i_13_189_3766_0 | (~i_13_189_1270_0 & ~i_13_189_4032_0))) | (i_13_189_311_0 & ~i_13_189_838_0) | (i_13_189_29_0 & ~i_13_189_1750_0 & ~i_13_189_1792_0) | (i_13_189_334_0 & i_13_189_694_0 & i_13_189_2848_0 & ~i_13_189_3387_0 & ~i_13_189_3451_0) | (~i_13_189_694_0 & ~i_13_189_3388_0 & ~i_13_189_3906_0) | (~i_13_189_1117_0 & ~i_13_189_4269_0));
endmodule



// Benchmark "kernel_13_190" written by ABC on Sun Jul 19 10:48:04 2020

module kernel_13_190 ( 
    i_13_190_76_0, i_13_190_184_0, i_13_190_189_0, i_13_190_229_0,
    i_13_190_408_0, i_13_190_415_0, i_13_190_418_0, i_13_190_517_0,
    i_13_190_549_0, i_13_190_571_0, i_13_190_604_0, i_13_190_657_0,
    i_13_190_658_0, i_13_190_665_0, i_13_190_761_0, i_13_190_793_0,
    i_13_190_847_0, i_13_190_855_0, i_13_190_856_0, i_13_190_885_0,
    i_13_190_936_0, i_13_190_937_0, i_13_190_1129_0, i_13_190_1144_0,
    i_13_190_1266_0, i_13_190_1420_0, i_13_190_1513_0, i_13_190_1518_0,
    i_13_190_1710_0, i_13_190_1711_0, i_13_190_1741_0, i_13_190_1742_0,
    i_13_190_1885_0, i_13_190_2019_0, i_13_190_2020_0, i_13_190_2024_0,
    i_13_190_2159_0, i_13_190_2224_0, i_13_190_2263_0, i_13_190_2321_0,
    i_13_190_2442_0, i_13_190_2448_0, i_13_190_2462_0, i_13_190_2466_0,
    i_13_190_2467_0, i_13_190_2470_0, i_13_190_2501_0, i_13_190_2512_0,
    i_13_190_2514_0, i_13_190_2538_0, i_13_190_2595_0, i_13_190_2611_0,
    i_13_190_2647_0, i_13_190_2692_0, i_13_190_2708_0, i_13_190_2730_0,
    i_13_190_2734_0, i_13_190_2881_0, i_13_190_2907_0, i_13_190_2908_0,
    i_13_190_2938_0, i_13_190_3037_0, i_13_190_3105_0, i_13_190_3325_0,
    i_13_190_3478_0, i_13_190_3483_0, i_13_190_3484_0, i_13_190_3486_0,
    i_13_190_3487_0, i_13_190_3565_0, i_13_190_3639_0, i_13_190_3640_0,
    i_13_190_3763_0, i_13_190_3861_0, i_13_190_3865_0, i_13_190_3868_0,
    i_13_190_3965_0, i_13_190_3992_0, i_13_190_4008_0, i_13_190_4009_0,
    i_13_190_4018_0, i_13_190_4098_0, i_13_190_4116_0, i_13_190_4127_0,
    i_13_190_4158_0, i_13_190_4159_0, i_13_190_4161_0, i_13_190_4198_0,
    i_13_190_4321_0, i_13_190_4324_0, i_13_190_4330_0, i_13_190_4333_0,
    i_13_190_4335_0, i_13_190_4365_0, i_13_190_4366_0, i_13_190_4369_0,
    i_13_190_4454_0, i_13_190_4458_0, i_13_190_4535_0, i_13_190_4599_0,
    o_13_190_0_0  );
  input  i_13_190_76_0, i_13_190_184_0, i_13_190_189_0, i_13_190_229_0,
    i_13_190_408_0, i_13_190_415_0, i_13_190_418_0, i_13_190_517_0,
    i_13_190_549_0, i_13_190_571_0, i_13_190_604_0, i_13_190_657_0,
    i_13_190_658_0, i_13_190_665_0, i_13_190_761_0, i_13_190_793_0,
    i_13_190_847_0, i_13_190_855_0, i_13_190_856_0, i_13_190_885_0,
    i_13_190_936_0, i_13_190_937_0, i_13_190_1129_0, i_13_190_1144_0,
    i_13_190_1266_0, i_13_190_1420_0, i_13_190_1513_0, i_13_190_1518_0,
    i_13_190_1710_0, i_13_190_1711_0, i_13_190_1741_0, i_13_190_1742_0,
    i_13_190_1885_0, i_13_190_2019_0, i_13_190_2020_0, i_13_190_2024_0,
    i_13_190_2159_0, i_13_190_2224_0, i_13_190_2263_0, i_13_190_2321_0,
    i_13_190_2442_0, i_13_190_2448_0, i_13_190_2462_0, i_13_190_2466_0,
    i_13_190_2467_0, i_13_190_2470_0, i_13_190_2501_0, i_13_190_2512_0,
    i_13_190_2514_0, i_13_190_2538_0, i_13_190_2595_0, i_13_190_2611_0,
    i_13_190_2647_0, i_13_190_2692_0, i_13_190_2708_0, i_13_190_2730_0,
    i_13_190_2734_0, i_13_190_2881_0, i_13_190_2907_0, i_13_190_2908_0,
    i_13_190_2938_0, i_13_190_3037_0, i_13_190_3105_0, i_13_190_3325_0,
    i_13_190_3478_0, i_13_190_3483_0, i_13_190_3484_0, i_13_190_3486_0,
    i_13_190_3487_0, i_13_190_3565_0, i_13_190_3639_0, i_13_190_3640_0,
    i_13_190_3763_0, i_13_190_3861_0, i_13_190_3865_0, i_13_190_3868_0,
    i_13_190_3965_0, i_13_190_3992_0, i_13_190_4008_0, i_13_190_4009_0,
    i_13_190_4018_0, i_13_190_4098_0, i_13_190_4116_0, i_13_190_4127_0,
    i_13_190_4158_0, i_13_190_4159_0, i_13_190_4161_0, i_13_190_4198_0,
    i_13_190_4321_0, i_13_190_4324_0, i_13_190_4330_0, i_13_190_4333_0,
    i_13_190_4335_0, i_13_190_4365_0, i_13_190_4366_0, i_13_190_4369_0,
    i_13_190_4454_0, i_13_190_4458_0, i_13_190_4535_0, i_13_190_4599_0;
  output o_13_190_0_0;
  assign o_13_190_0_0 = ~((~i_13_190_2448_0 & ((~i_13_190_517_0 & ~i_13_190_3565_0 & ~i_13_190_4159_0 & ~i_13_190_4365_0) | (~i_13_190_189_0 & ~i_13_190_3484_0 & ~i_13_190_4161_0 & ~i_13_190_4366_0))) | (i_13_190_184_0 & i_13_190_1266_0) | (i_13_190_229_0 & ~i_13_190_3565_0 & ~i_13_190_3861_0 & ~i_13_190_4365_0) | (~i_13_190_855_0 & ~i_13_190_3865_0 & ~i_13_190_4369_0));
endmodule



// Benchmark "kernel_13_191" written by ABC on Sun Jul 19 10:48:05 2020

module kernel_13_191 ( 
    i_13_191_46_0, i_13_191_47_0, i_13_191_66_0, i_13_191_100_0,
    i_13_191_262_0, i_13_191_567_0, i_13_191_585_0, i_13_191_587_0,
    i_13_191_639_0, i_13_191_640_0, i_13_191_675_0, i_13_191_689_0,
    i_13_191_946_0, i_13_191_1063_0, i_13_191_1064_0, i_13_191_1207_0,
    i_13_191_1260_0, i_13_191_1272_0, i_13_191_1282_0, i_13_191_1323_0,
    i_13_191_1343_0, i_13_191_1435_0, i_13_191_1468_0, i_13_191_1505_0,
    i_13_191_1507_0, i_13_191_1567_0, i_13_191_1568_0, i_13_191_1596_0,
    i_13_191_1597_0, i_13_191_1802_0, i_13_191_1810_0, i_13_191_1855_0,
    i_13_191_1927_0, i_13_191_1935_0, i_13_191_1945_0, i_13_191_1992_0,
    i_13_191_2017_0, i_13_191_2053_0, i_13_191_2054_0, i_13_191_2107_0,
    i_13_191_2117_0, i_13_191_2135_0, i_13_191_2146_0, i_13_191_2153_0,
    i_13_191_2189_0, i_13_191_2244_0, i_13_191_2261_0, i_13_191_2278_0,
    i_13_191_2279_0, i_13_191_2351_0, i_13_191_2404_0, i_13_191_2405_0,
    i_13_191_2417_0, i_13_191_2585_0, i_13_191_2611_0, i_13_191_2615_0,
    i_13_191_2694_0, i_13_191_2713_0, i_13_191_2745_0, i_13_191_2746_0,
    i_13_191_2782_0, i_13_191_2898_0, i_13_191_2934_0, i_13_191_2935_0,
    i_13_191_3025_0, i_13_191_3054_0, i_13_191_3145_0, i_13_191_3313_0,
    i_13_191_3339_0, i_13_191_3340_0, i_13_191_3341_0, i_13_191_3367_0,
    i_13_191_3368_0, i_13_191_3385_0, i_13_191_3386_0, i_13_191_3414_0,
    i_13_191_3415_0, i_13_191_3456_0, i_13_191_3481_0, i_13_191_3529_0,
    i_13_191_3548_0, i_13_191_3592_0, i_13_191_3627_0, i_13_191_3754_0,
    i_13_191_3817_0, i_13_191_3818_0, i_13_191_3889_0, i_13_191_3901_0,
    i_13_191_3909_0, i_13_191_3936_0, i_13_191_4041_0, i_13_191_4042_0,
    i_13_191_4230_0, i_13_191_4231_0, i_13_191_4232_0, i_13_191_4258_0,
    i_13_191_4268_0, i_13_191_4304_0, i_13_191_4324_0, i_13_191_4394_0,
    o_13_191_0_0  );
  input  i_13_191_46_0, i_13_191_47_0, i_13_191_66_0, i_13_191_100_0,
    i_13_191_262_0, i_13_191_567_0, i_13_191_585_0, i_13_191_587_0,
    i_13_191_639_0, i_13_191_640_0, i_13_191_675_0, i_13_191_689_0,
    i_13_191_946_0, i_13_191_1063_0, i_13_191_1064_0, i_13_191_1207_0,
    i_13_191_1260_0, i_13_191_1272_0, i_13_191_1282_0, i_13_191_1323_0,
    i_13_191_1343_0, i_13_191_1435_0, i_13_191_1468_0, i_13_191_1505_0,
    i_13_191_1507_0, i_13_191_1567_0, i_13_191_1568_0, i_13_191_1596_0,
    i_13_191_1597_0, i_13_191_1802_0, i_13_191_1810_0, i_13_191_1855_0,
    i_13_191_1927_0, i_13_191_1935_0, i_13_191_1945_0, i_13_191_1992_0,
    i_13_191_2017_0, i_13_191_2053_0, i_13_191_2054_0, i_13_191_2107_0,
    i_13_191_2117_0, i_13_191_2135_0, i_13_191_2146_0, i_13_191_2153_0,
    i_13_191_2189_0, i_13_191_2244_0, i_13_191_2261_0, i_13_191_2278_0,
    i_13_191_2279_0, i_13_191_2351_0, i_13_191_2404_0, i_13_191_2405_0,
    i_13_191_2417_0, i_13_191_2585_0, i_13_191_2611_0, i_13_191_2615_0,
    i_13_191_2694_0, i_13_191_2713_0, i_13_191_2745_0, i_13_191_2746_0,
    i_13_191_2782_0, i_13_191_2898_0, i_13_191_2934_0, i_13_191_2935_0,
    i_13_191_3025_0, i_13_191_3054_0, i_13_191_3145_0, i_13_191_3313_0,
    i_13_191_3339_0, i_13_191_3340_0, i_13_191_3341_0, i_13_191_3367_0,
    i_13_191_3368_0, i_13_191_3385_0, i_13_191_3386_0, i_13_191_3414_0,
    i_13_191_3415_0, i_13_191_3456_0, i_13_191_3481_0, i_13_191_3529_0,
    i_13_191_3548_0, i_13_191_3592_0, i_13_191_3627_0, i_13_191_3754_0,
    i_13_191_3817_0, i_13_191_3818_0, i_13_191_3889_0, i_13_191_3901_0,
    i_13_191_3909_0, i_13_191_3936_0, i_13_191_4041_0, i_13_191_4042_0,
    i_13_191_4230_0, i_13_191_4231_0, i_13_191_4232_0, i_13_191_4258_0,
    i_13_191_4268_0, i_13_191_4304_0, i_13_191_4324_0, i_13_191_4394_0;
  output o_13_191_0_0;
  assign o_13_191_0_0 = ~((~i_13_191_4230_0 & ((~i_13_191_2782_0 & (i_13_191_946_0 | (~i_13_191_587_0 & i_13_191_1597_0))) | (i_13_191_1855_0 & ~i_13_191_3754_0))) | (~i_13_191_2278_0 & ~i_13_191_2404_0 & ~i_13_191_3313_0) | (~i_13_191_2017_0 & ~i_13_191_3592_0));
endmodule



// Benchmark "kernel_13_192" written by ABC on Sun Jul 19 10:48:05 2020

module kernel_13_192 ( 
    i_13_192_45_0, i_13_192_112_0, i_13_192_138_0, i_13_192_139_0,
    i_13_192_172_0, i_13_192_174_0, i_13_192_279_0, i_13_192_405_0,
    i_13_192_406_0, i_13_192_414_0, i_13_192_441_0, i_13_192_505_0,
    i_13_192_567_0, i_13_192_633_0, i_13_192_657_0, i_13_192_658_0,
    i_13_192_660_0, i_13_192_666_0, i_13_192_667_0, i_13_192_669_0,
    i_13_192_828_0, i_13_192_831_0, i_13_192_940_0, i_13_192_945_0,
    i_13_192_1071_0, i_13_192_1072_0, i_13_192_1081_0, i_13_192_1147_0,
    i_13_192_1228_0, i_13_192_1284_0, i_13_192_1305_0, i_13_192_1306_0,
    i_13_192_1326_0, i_13_192_1423_0, i_13_192_1494_0, i_13_192_1497_0,
    i_13_192_1498_0, i_13_192_1504_0, i_13_192_1522_0, i_13_192_1548_0,
    i_13_192_1593_0, i_13_192_1620_0, i_13_192_1633_0, i_13_192_1684_0,
    i_13_192_1695_0, i_13_192_1729_0, i_13_192_1737_0, i_13_192_1764_0,
    i_13_192_1777_0, i_13_192_1837_0, i_13_192_1858_0, i_13_192_1926_0,
    i_13_192_1938_0, i_13_192_2019_0, i_13_192_2020_0, i_13_192_2296_0,
    i_13_192_2316_0, i_13_192_2344_0, i_13_192_2395_0, i_13_192_2430_0,
    i_13_192_2431_0, i_13_192_2448_0, i_13_192_2469_0, i_13_192_2511_0,
    i_13_192_2610_0, i_13_192_2637_0, i_13_192_2719_0, i_13_192_2757_0,
    i_13_192_2781_0, i_13_192_3070_0, i_13_192_3108_0, i_13_192_3126_0,
    i_13_192_3172_0, i_13_192_3241_0, i_13_192_3258_0, i_13_192_3261_0,
    i_13_192_3268_0, i_13_192_3271_0, i_13_192_3406_0, i_13_192_3420_0,
    i_13_192_3423_0, i_13_192_3546_0, i_13_192_3637_0, i_13_192_3640_0,
    i_13_192_3667_0, i_13_192_3897_0, i_13_192_3910_0, i_13_192_4035_0,
    i_13_192_4051_0, i_13_192_4086_0, i_13_192_4248_0, i_13_192_4251_0,
    i_13_192_4252_0, i_13_192_4260_0, i_13_192_4321_0, i_13_192_4429_0,
    i_13_192_4458_0, i_13_192_4503_0, i_13_192_4564_0, i_13_192_4593_0,
    o_13_192_0_0  );
  input  i_13_192_45_0, i_13_192_112_0, i_13_192_138_0, i_13_192_139_0,
    i_13_192_172_0, i_13_192_174_0, i_13_192_279_0, i_13_192_405_0,
    i_13_192_406_0, i_13_192_414_0, i_13_192_441_0, i_13_192_505_0,
    i_13_192_567_0, i_13_192_633_0, i_13_192_657_0, i_13_192_658_0,
    i_13_192_660_0, i_13_192_666_0, i_13_192_667_0, i_13_192_669_0,
    i_13_192_828_0, i_13_192_831_0, i_13_192_940_0, i_13_192_945_0,
    i_13_192_1071_0, i_13_192_1072_0, i_13_192_1081_0, i_13_192_1147_0,
    i_13_192_1228_0, i_13_192_1284_0, i_13_192_1305_0, i_13_192_1306_0,
    i_13_192_1326_0, i_13_192_1423_0, i_13_192_1494_0, i_13_192_1497_0,
    i_13_192_1498_0, i_13_192_1504_0, i_13_192_1522_0, i_13_192_1548_0,
    i_13_192_1593_0, i_13_192_1620_0, i_13_192_1633_0, i_13_192_1684_0,
    i_13_192_1695_0, i_13_192_1729_0, i_13_192_1737_0, i_13_192_1764_0,
    i_13_192_1777_0, i_13_192_1837_0, i_13_192_1858_0, i_13_192_1926_0,
    i_13_192_1938_0, i_13_192_2019_0, i_13_192_2020_0, i_13_192_2296_0,
    i_13_192_2316_0, i_13_192_2344_0, i_13_192_2395_0, i_13_192_2430_0,
    i_13_192_2431_0, i_13_192_2448_0, i_13_192_2469_0, i_13_192_2511_0,
    i_13_192_2610_0, i_13_192_2637_0, i_13_192_2719_0, i_13_192_2757_0,
    i_13_192_2781_0, i_13_192_3070_0, i_13_192_3108_0, i_13_192_3126_0,
    i_13_192_3172_0, i_13_192_3241_0, i_13_192_3258_0, i_13_192_3261_0,
    i_13_192_3268_0, i_13_192_3271_0, i_13_192_3406_0, i_13_192_3420_0,
    i_13_192_3423_0, i_13_192_3546_0, i_13_192_3637_0, i_13_192_3640_0,
    i_13_192_3667_0, i_13_192_3897_0, i_13_192_3910_0, i_13_192_4035_0,
    i_13_192_4051_0, i_13_192_4086_0, i_13_192_4248_0, i_13_192_4251_0,
    i_13_192_4252_0, i_13_192_4260_0, i_13_192_4321_0, i_13_192_4429_0,
    i_13_192_4458_0, i_13_192_4503_0, i_13_192_4564_0, i_13_192_4593_0;
  output o_13_192_0_0;
  assign o_13_192_0_0 = ~((~i_13_192_1326_0 & ~i_13_192_1593_0) | (~i_13_192_828_0 & ~i_13_192_1522_0));
endmodule



// Benchmark "kernel_13_193" written by ABC on Sun Jul 19 10:48:06 2020

module kernel_13_193 ( 
    i_13_193_28_0, i_13_193_91_0, i_13_193_92_0, i_13_193_176_0,
    i_13_193_181_0, i_13_193_256_0, i_13_193_274_0, i_13_193_307_0,
    i_13_193_308_0, i_13_193_310_0, i_13_193_315_0, i_13_193_316_0,
    i_13_193_317_0, i_13_193_337_0, i_13_193_371_0, i_13_193_379_0,
    i_13_193_407_0, i_13_193_408_0, i_13_193_551_0, i_13_193_589_0,
    i_13_193_604_0, i_13_193_639_0, i_13_193_640_0, i_13_193_666_0,
    i_13_193_668_0, i_13_193_670_0, i_13_193_676_0, i_13_193_723_0,
    i_13_193_757_0, i_13_193_769_0, i_13_193_842_0, i_13_193_867_0,
    i_13_193_875_0, i_13_193_981_0, i_13_193_1021_0, i_13_193_1063_0,
    i_13_193_1093_0, i_13_193_1218_0, i_13_193_1300_0, i_13_193_1318_0,
    i_13_193_1324_0, i_13_193_1325_0, i_13_193_1480_0, i_13_193_1595_0,
    i_13_193_1602_0, i_13_193_1699_0, i_13_193_1828_0, i_13_193_1840_0,
    i_13_193_1909_0, i_13_193_1926_0, i_13_193_2116_0, i_13_193_2245_0,
    i_13_193_2260_0, i_13_193_2280_0, i_13_193_2407_0, i_13_193_2511_0,
    i_13_193_2648_0, i_13_193_2660_0, i_13_193_2673_0, i_13_193_2675_0,
    i_13_193_2678_0, i_13_193_2767_0, i_13_193_2781_0, i_13_193_2785_0,
    i_13_193_2981_0, i_13_193_3100_0, i_13_193_3128_0, i_13_193_3416_0,
    i_13_193_3469_0, i_13_193_3479_0, i_13_193_3482_0, i_13_193_3529_0,
    i_13_193_3541_0, i_13_193_3631_0, i_13_193_3682_0, i_13_193_3738_0,
    i_13_193_3766_0, i_13_193_3767_0, i_13_193_3817_0, i_13_193_3818_0,
    i_13_193_3889_0, i_13_193_3925_0, i_13_193_3991_0, i_13_193_3992_0,
    i_13_193_4033_0, i_13_193_4034_0, i_13_193_4041_0, i_13_193_4078_0,
    i_13_193_4086_0, i_13_193_4234_0, i_13_193_4252_0, i_13_193_4262_0,
    i_13_193_4270_0, i_13_193_4305_0, i_13_193_4351_0, i_13_193_4519_0,
    i_13_193_4522_0, i_13_193_4565_0, i_13_193_4567_0, i_13_193_4591_0,
    o_13_193_0_0  );
  input  i_13_193_28_0, i_13_193_91_0, i_13_193_92_0, i_13_193_176_0,
    i_13_193_181_0, i_13_193_256_0, i_13_193_274_0, i_13_193_307_0,
    i_13_193_308_0, i_13_193_310_0, i_13_193_315_0, i_13_193_316_0,
    i_13_193_317_0, i_13_193_337_0, i_13_193_371_0, i_13_193_379_0,
    i_13_193_407_0, i_13_193_408_0, i_13_193_551_0, i_13_193_589_0,
    i_13_193_604_0, i_13_193_639_0, i_13_193_640_0, i_13_193_666_0,
    i_13_193_668_0, i_13_193_670_0, i_13_193_676_0, i_13_193_723_0,
    i_13_193_757_0, i_13_193_769_0, i_13_193_842_0, i_13_193_867_0,
    i_13_193_875_0, i_13_193_981_0, i_13_193_1021_0, i_13_193_1063_0,
    i_13_193_1093_0, i_13_193_1218_0, i_13_193_1300_0, i_13_193_1318_0,
    i_13_193_1324_0, i_13_193_1325_0, i_13_193_1480_0, i_13_193_1595_0,
    i_13_193_1602_0, i_13_193_1699_0, i_13_193_1828_0, i_13_193_1840_0,
    i_13_193_1909_0, i_13_193_1926_0, i_13_193_2116_0, i_13_193_2245_0,
    i_13_193_2260_0, i_13_193_2280_0, i_13_193_2407_0, i_13_193_2511_0,
    i_13_193_2648_0, i_13_193_2660_0, i_13_193_2673_0, i_13_193_2675_0,
    i_13_193_2678_0, i_13_193_2767_0, i_13_193_2781_0, i_13_193_2785_0,
    i_13_193_2981_0, i_13_193_3100_0, i_13_193_3128_0, i_13_193_3416_0,
    i_13_193_3469_0, i_13_193_3479_0, i_13_193_3482_0, i_13_193_3529_0,
    i_13_193_3541_0, i_13_193_3631_0, i_13_193_3682_0, i_13_193_3738_0,
    i_13_193_3766_0, i_13_193_3767_0, i_13_193_3817_0, i_13_193_3818_0,
    i_13_193_3889_0, i_13_193_3925_0, i_13_193_3991_0, i_13_193_3992_0,
    i_13_193_4033_0, i_13_193_4034_0, i_13_193_4041_0, i_13_193_4078_0,
    i_13_193_4086_0, i_13_193_4234_0, i_13_193_4252_0, i_13_193_4262_0,
    i_13_193_4270_0, i_13_193_4305_0, i_13_193_4351_0, i_13_193_4519_0,
    i_13_193_4522_0, i_13_193_4565_0, i_13_193_4567_0, i_13_193_4591_0;
  output o_13_193_0_0;
  assign o_13_193_0_0 = ~((~i_13_193_316_0 & ~i_13_193_842_0 & ((~i_13_193_181_0 & i_13_193_1480_0) | (~i_13_193_4034_0 & ~i_13_193_4567_0))) | (~i_13_193_315_0 & ~i_13_193_317_0 & ~i_13_193_666_0 & ~i_13_193_668_0) | (~i_13_193_1325_0 & ~i_13_193_4078_0 & ~i_13_193_4351_0) | (~i_13_193_91_0 & ~i_13_193_176_0 & i_13_193_1828_0 & ~i_13_193_4565_0));
endmodule



// Benchmark "kernel_13_194" written by ABC on Sun Jul 19 10:48:07 2020

module kernel_13_194 ( 
    i_13_194_51_0, i_13_194_123_0, i_13_194_124_0, i_13_194_141_0,
    i_13_194_169_0, i_13_194_240_0, i_13_194_241_0, i_13_194_250_0,
    i_13_194_375_0, i_13_194_456_0, i_13_194_467_0, i_13_194_588_0,
    i_13_194_618_0, i_13_194_619_0, i_13_194_654_0, i_13_194_682_0,
    i_13_194_699_0, i_13_194_763_0, i_13_194_850_0, i_13_194_931_0,
    i_13_194_943_0, i_13_194_979_0, i_13_194_980_0, i_13_194_1033_0,
    i_13_194_1058_0, i_13_194_1059_0, i_13_194_1077_0, i_13_194_1078_0,
    i_13_194_1079_0, i_13_194_1084_0, i_13_194_1401_0, i_13_194_1448_0,
    i_13_194_1470_0, i_13_194_1501_0, i_13_194_1502_0, i_13_194_1507_0,
    i_13_194_1525_0, i_13_194_1528_0, i_13_194_1599_0, i_13_194_1608_0,
    i_13_194_1609_0, i_13_194_1635_0, i_13_194_1636_0, i_13_194_1637_0,
    i_13_194_1777_0, i_13_194_1815_0, i_13_194_2002_0, i_13_194_2014_0,
    i_13_194_2140_0, i_13_194_2211_0, i_13_194_2226_0, i_13_194_2284_0,
    i_13_194_2294_0, i_13_194_2319_0, i_13_194_2454_0, i_13_194_2544_0,
    i_13_194_2616_0, i_13_194_2787_0, i_13_194_2788_0, i_13_194_2887_0,
    i_13_194_2922_0, i_13_194_2923_0, i_13_194_2959_0, i_13_194_3003_0,
    i_13_194_3023_0, i_13_194_3219_0, i_13_194_3220_0, i_13_194_3372_0,
    i_13_194_3382_0, i_13_194_3406_0, i_13_194_3417_0, i_13_194_3418_0,
    i_13_194_3428_0, i_13_194_3463_0, i_13_194_3464_0, i_13_194_3471_0,
    i_13_194_3541_0, i_13_194_3553_0, i_13_194_3569_0, i_13_194_3577_0,
    i_13_194_3643_0, i_13_194_3723_0, i_13_194_3730_0, i_13_194_3769_0,
    i_13_194_3788_0, i_13_194_3877_0, i_13_194_3903_0, i_13_194_3904_0,
    i_13_194_4011_0, i_13_194_4012_0, i_13_194_4020_0, i_13_194_4082_0,
    i_13_194_4089_0, i_13_194_4091_0, i_13_194_4389_0, i_13_194_4396_0,
    i_13_194_4418_0, i_13_194_4533_0, i_13_194_4557_0, i_13_194_4589_0,
    o_13_194_0_0  );
  input  i_13_194_51_0, i_13_194_123_0, i_13_194_124_0, i_13_194_141_0,
    i_13_194_169_0, i_13_194_240_0, i_13_194_241_0, i_13_194_250_0,
    i_13_194_375_0, i_13_194_456_0, i_13_194_467_0, i_13_194_588_0,
    i_13_194_618_0, i_13_194_619_0, i_13_194_654_0, i_13_194_682_0,
    i_13_194_699_0, i_13_194_763_0, i_13_194_850_0, i_13_194_931_0,
    i_13_194_943_0, i_13_194_979_0, i_13_194_980_0, i_13_194_1033_0,
    i_13_194_1058_0, i_13_194_1059_0, i_13_194_1077_0, i_13_194_1078_0,
    i_13_194_1079_0, i_13_194_1084_0, i_13_194_1401_0, i_13_194_1448_0,
    i_13_194_1470_0, i_13_194_1501_0, i_13_194_1502_0, i_13_194_1507_0,
    i_13_194_1525_0, i_13_194_1528_0, i_13_194_1599_0, i_13_194_1608_0,
    i_13_194_1609_0, i_13_194_1635_0, i_13_194_1636_0, i_13_194_1637_0,
    i_13_194_1777_0, i_13_194_1815_0, i_13_194_2002_0, i_13_194_2014_0,
    i_13_194_2140_0, i_13_194_2211_0, i_13_194_2226_0, i_13_194_2284_0,
    i_13_194_2294_0, i_13_194_2319_0, i_13_194_2454_0, i_13_194_2544_0,
    i_13_194_2616_0, i_13_194_2787_0, i_13_194_2788_0, i_13_194_2887_0,
    i_13_194_2922_0, i_13_194_2923_0, i_13_194_2959_0, i_13_194_3003_0,
    i_13_194_3023_0, i_13_194_3219_0, i_13_194_3220_0, i_13_194_3372_0,
    i_13_194_3382_0, i_13_194_3406_0, i_13_194_3417_0, i_13_194_3418_0,
    i_13_194_3428_0, i_13_194_3463_0, i_13_194_3464_0, i_13_194_3471_0,
    i_13_194_3541_0, i_13_194_3553_0, i_13_194_3569_0, i_13_194_3577_0,
    i_13_194_3643_0, i_13_194_3723_0, i_13_194_3730_0, i_13_194_3769_0,
    i_13_194_3788_0, i_13_194_3877_0, i_13_194_3903_0, i_13_194_3904_0,
    i_13_194_4011_0, i_13_194_4012_0, i_13_194_4020_0, i_13_194_4082_0,
    i_13_194_4089_0, i_13_194_4091_0, i_13_194_4389_0, i_13_194_4396_0,
    i_13_194_4418_0, i_13_194_4533_0, i_13_194_4557_0, i_13_194_4589_0;
  output o_13_194_0_0;
  assign o_13_194_0_0 = ~((i_13_194_4418_0 & (~i_13_194_2788_0 | (~i_13_194_1501_0 & ~i_13_194_4091_0))) | (~i_13_194_619_0 & ~i_13_194_3903_0) | (~i_13_194_1608_0 & ~i_13_194_2923_0 & ~i_13_194_4089_0) | (~i_13_194_943_0 & ~i_13_194_4082_0 & i_13_194_4091_0));
endmodule



// Benchmark "kernel_13_195" written by ABC on Sun Jul 19 10:48:08 2020

module kernel_13_195 ( 
    i_13_195_64_0, i_13_195_65_0, i_13_195_76_0, i_13_195_131_0,
    i_13_195_158_0, i_13_195_160_0, i_13_195_163_0, i_13_195_164_0,
    i_13_195_307_0, i_13_195_355_0, i_13_195_358_0, i_13_195_463_0,
    i_13_195_465_0, i_13_195_466_0, i_13_195_469_0, i_13_195_490_0,
    i_13_195_492_0, i_13_195_537_0, i_13_195_564_0, i_13_195_580_0,
    i_13_195_697_0, i_13_195_812_0, i_13_195_829_0, i_13_195_831_0,
    i_13_195_839_0, i_13_195_1100_0, i_13_195_1121_0, i_13_195_1131_0,
    i_13_195_1302_0, i_13_195_1307_0, i_13_195_1345_0, i_13_195_1389_0,
    i_13_195_1396_0, i_13_195_1397_0, i_13_195_1400_0, i_13_195_1434_0,
    i_13_195_1471_0, i_13_195_1504_0, i_13_195_1594_0, i_13_195_1609_0,
    i_13_195_1696_0, i_13_195_1697_0, i_13_195_1783_0, i_13_195_1784_0,
    i_13_195_1793_0, i_13_195_1794_0, i_13_195_1840_0, i_13_195_1846_0,
    i_13_195_1847_0, i_13_195_1859_0, i_13_195_1928_0, i_13_195_1990_0,
    i_13_195_1995_0, i_13_195_2032_0, i_13_195_2101_0, i_13_195_2108_0,
    i_13_195_2111_0, i_13_195_2143_0, i_13_195_2187_0, i_13_195_2200_0,
    i_13_195_2202_0, i_13_195_2203_0, i_13_195_2206_0, i_13_195_2237_0,
    i_13_195_2297_0, i_13_195_2379_0, i_13_195_2404_0, i_13_195_2405_0,
    i_13_195_2506_0, i_13_195_2585_0, i_13_195_2692_0, i_13_195_2881_0,
    i_13_195_2884_0, i_13_195_2936_0, i_13_195_3165_0, i_13_195_3241_0,
    i_13_195_3242_0, i_13_195_3309_0, i_13_195_3380_0, i_13_195_3415_0,
    i_13_195_3422_0, i_13_195_3539_0, i_13_195_3568_0, i_13_195_3596_0,
    i_13_195_3597_0, i_13_195_3598_0, i_13_195_3619_0, i_13_195_3631_0,
    i_13_195_3633_0, i_13_195_3638_0, i_13_195_3686_0, i_13_195_3845_0,
    i_13_195_3856_0, i_13_195_3912_0, i_13_195_4060_0, i_13_195_4189_0,
    i_13_195_4313_0, i_13_195_4416_0, i_13_195_4453_0, i_13_195_4510_0,
    o_13_195_0_0  );
  input  i_13_195_64_0, i_13_195_65_0, i_13_195_76_0, i_13_195_131_0,
    i_13_195_158_0, i_13_195_160_0, i_13_195_163_0, i_13_195_164_0,
    i_13_195_307_0, i_13_195_355_0, i_13_195_358_0, i_13_195_463_0,
    i_13_195_465_0, i_13_195_466_0, i_13_195_469_0, i_13_195_490_0,
    i_13_195_492_0, i_13_195_537_0, i_13_195_564_0, i_13_195_580_0,
    i_13_195_697_0, i_13_195_812_0, i_13_195_829_0, i_13_195_831_0,
    i_13_195_839_0, i_13_195_1100_0, i_13_195_1121_0, i_13_195_1131_0,
    i_13_195_1302_0, i_13_195_1307_0, i_13_195_1345_0, i_13_195_1389_0,
    i_13_195_1396_0, i_13_195_1397_0, i_13_195_1400_0, i_13_195_1434_0,
    i_13_195_1471_0, i_13_195_1504_0, i_13_195_1594_0, i_13_195_1609_0,
    i_13_195_1696_0, i_13_195_1697_0, i_13_195_1783_0, i_13_195_1784_0,
    i_13_195_1793_0, i_13_195_1794_0, i_13_195_1840_0, i_13_195_1846_0,
    i_13_195_1847_0, i_13_195_1859_0, i_13_195_1928_0, i_13_195_1990_0,
    i_13_195_1995_0, i_13_195_2032_0, i_13_195_2101_0, i_13_195_2108_0,
    i_13_195_2111_0, i_13_195_2143_0, i_13_195_2187_0, i_13_195_2200_0,
    i_13_195_2202_0, i_13_195_2203_0, i_13_195_2206_0, i_13_195_2237_0,
    i_13_195_2297_0, i_13_195_2379_0, i_13_195_2404_0, i_13_195_2405_0,
    i_13_195_2506_0, i_13_195_2585_0, i_13_195_2692_0, i_13_195_2881_0,
    i_13_195_2884_0, i_13_195_2936_0, i_13_195_3165_0, i_13_195_3241_0,
    i_13_195_3242_0, i_13_195_3309_0, i_13_195_3380_0, i_13_195_3415_0,
    i_13_195_3422_0, i_13_195_3539_0, i_13_195_3568_0, i_13_195_3596_0,
    i_13_195_3597_0, i_13_195_3598_0, i_13_195_3619_0, i_13_195_3631_0,
    i_13_195_3633_0, i_13_195_3638_0, i_13_195_3686_0, i_13_195_3845_0,
    i_13_195_3856_0, i_13_195_3912_0, i_13_195_4060_0, i_13_195_4189_0,
    i_13_195_4313_0, i_13_195_4416_0, i_13_195_4453_0, i_13_195_4510_0;
  output o_13_195_0_0;
  assign o_13_195_0_0 = ~((~i_13_195_2143_0 & ~i_13_195_3856_0) | (i_13_195_2884_0 & ~i_13_195_3619_0) | (~i_13_195_64_0 & ~i_13_195_1847_0 & ~i_13_195_2936_0));
endmodule



// Benchmark "kernel_13_196" written by ABC on Sun Jul 19 10:48:08 2020

module kernel_13_196 ( 
    i_13_196_64_0, i_13_196_77_0, i_13_196_121_0, i_13_196_179_0,
    i_13_196_184_0, i_13_196_229_0, i_13_196_232_0, i_13_196_358_0,
    i_13_196_374_0, i_13_196_415_0, i_13_196_527_0, i_13_196_530_0,
    i_13_196_557_0, i_13_196_599_0, i_13_196_608_0, i_13_196_611_0,
    i_13_196_661_0, i_13_196_662_0, i_13_196_664_0, i_13_196_665_0,
    i_13_196_800_0, i_13_196_829_0, i_13_196_832_0, i_13_196_833_0,
    i_13_196_850_0, i_13_196_895_0, i_13_196_1066_0, i_13_196_1121_0,
    i_13_196_1213_0, i_13_196_1228_0, i_13_196_1229_0, i_13_196_1307_0,
    i_13_196_1309_0, i_13_196_1310_0, i_13_196_1313_0, i_13_196_1427_0,
    i_13_196_1430_0, i_13_196_1498_0, i_13_196_1499_0, i_13_196_1505_0,
    i_13_196_1553_0, i_13_196_1556_0, i_13_196_1568_0, i_13_196_1726_0,
    i_13_196_1811_0, i_13_196_1919_0, i_13_196_1922_0, i_13_196_1930_0,
    i_13_196_1961_0, i_13_196_1991_0, i_13_196_1993_0, i_13_196_2033_0,
    i_13_196_2297_0, i_13_196_2399_0, i_13_196_2452_0, i_13_196_2456_0,
    i_13_196_2467_0, i_13_196_2678_0, i_13_196_2693_0, i_13_196_2708_0,
    i_13_196_2768_0, i_13_196_2924_0, i_13_196_3010_0, i_13_196_3013_0,
    i_13_196_3037_0, i_13_196_3061_0, i_13_196_3062_0, i_13_196_3149_0,
    i_13_196_3217_0, i_13_196_3242_0, i_13_196_3260_0, i_13_196_3269_0,
    i_13_196_3289_0, i_13_196_3307_0, i_13_196_3394_0, i_13_196_3406_0,
    i_13_196_3461_0, i_13_196_3490_0, i_13_196_3523_0, i_13_196_3541_0,
    i_13_196_3542_0, i_13_196_3545_0, i_13_196_3580_0, i_13_196_3581_0,
    i_13_196_3734_0, i_13_196_3788_0, i_13_196_3806_0, i_13_196_3859_0,
    i_13_196_3860_0, i_13_196_3892_0, i_13_196_3895_0, i_13_196_3919_0,
    i_13_196_3983_0, i_13_196_4253_0, i_13_196_4256_0, i_13_196_4265_0,
    i_13_196_4430_0, i_13_196_4558_0, i_13_196_4559_0, i_13_196_4580_0,
    o_13_196_0_0  );
  input  i_13_196_64_0, i_13_196_77_0, i_13_196_121_0, i_13_196_179_0,
    i_13_196_184_0, i_13_196_229_0, i_13_196_232_0, i_13_196_358_0,
    i_13_196_374_0, i_13_196_415_0, i_13_196_527_0, i_13_196_530_0,
    i_13_196_557_0, i_13_196_599_0, i_13_196_608_0, i_13_196_611_0,
    i_13_196_661_0, i_13_196_662_0, i_13_196_664_0, i_13_196_665_0,
    i_13_196_800_0, i_13_196_829_0, i_13_196_832_0, i_13_196_833_0,
    i_13_196_850_0, i_13_196_895_0, i_13_196_1066_0, i_13_196_1121_0,
    i_13_196_1213_0, i_13_196_1228_0, i_13_196_1229_0, i_13_196_1307_0,
    i_13_196_1309_0, i_13_196_1310_0, i_13_196_1313_0, i_13_196_1427_0,
    i_13_196_1430_0, i_13_196_1498_0, i_13_196_1499_0, i_13_196_1505_0,
    i_13_196_1553_0, i_13_196_1556_0, i_13_196_1568_0, i_13_196_1726_0,
    i_13_196_1811_0, i_13_196_1919_0, i_13_196_1922_0, i_13_196_1930_0,
    i_13_196_1961_0, i_13_196_1991_0, i_13_196_1993_0, i_13_196_2033_0,
    i_13_196_2297_0, i_13_196_2399_0, i_13_196_2452_0, i_13_196_2456_0,
    i_13_196_2467_0, i_13_196_2678_0, i_13_196_2693_0, i_13_196_2708_0,
    i_13_196_2768_0, i_13_196_2924_0, i_13_196_3010_0, i_13_196_3013_0,
    i_13_196_3037_0, i_13_196_3061_0, i_13_196_3062_0, i_13_196_3149_0,
    i_13_196_3217_0, i_13_196_3242_0, i_13_196_3260_0, i_13_196_3269_0,
    i_13_196_3289_0, i_13_196_3307_0, i_13_196_3394_0, i_13_196_3406_0,
    i_13_196_3461_0, i_13_196_3490_0, i_13_196_3523_0, i_13_196_3541_0,
    i_13_196_3542_0, i_13_196_3545_0, i_13_196_3580_0, i_13_196_3581_0,
    i_13_196_3734_0, i_13_196_3788_0, i_13_196_3806_0, i_13_196_3859_0,
    i_13_196_3860_0, i_13_196_3892_0, i_13_196_3895_0, i_13_196_3919_0,
    i_13_196_3983_0, i_13_196_4253_0, i_13_196_4256_0, i_13_196_4265_0,
    i_13_196_4430_0, i_13_196_4558_0, i_13_196_4559_0, i_13_196_4580_0;
  output o_13_196_0_0;
  assign o_13_196_0_0 = ~((~i_13_196_3788_0 & (~i_13_196_1310_0 | (i_13_196_1228_0 & ~i_13_196_2452_0 & ~i_13_196_3541_0))) | (~i_13_196_4430_0 & ((~i_13_196_833_0 & ~i_13_196_3581_0 & ~i_13_196_3895_0) | (~i_13_196_1553_0 & ~i_13_196_3013_0 & ~i_13_196_4265_0))) | (i_13_196_1307_0 & i_13_196_3289_0 & ~i_13_196_3542_0) | (i_13_196_1811_0 & ~i_13_196_3983_0) | (~i_13_196_1991_0 & ~i_13_196_2924_0 & ~i_13_196_4253_0));
endmodule



// Benchmark "kernel_13_197" written by ABC on Sun Jul 19 10:48:09 2020

module kernel_13_197 ( 
    i_13_197_41_0, i_13_197_71_0, i_13_197_138_0, i_13_197_139_0,
    i_13_197_141_0, i_13_197_142_0, i_13_197_231_0, i_13_197_232_0,
    i_13_197_310_0, i_13_197_418_0, i_13_197_471_0, i_13_197_472_0,
    i_13_197_517_0, i_13_197_537_0, i_13_197_538_0, i_13_197_764_0,
    i_13_197_826_0, i_13_197_832_0, i_13_197_1029_0, i_13_197_1086_0,
    i_13_197_1214_0, i_13_197_1218_0, i_13_197_1219_0, i_13_197_1221_0,
    i_13_197_1222_0, i_13_197_1266_0, i_13_197_1276_0, i_13_197_1362_0,
    i_13_197_1392_0, i_13_197_1426_0, i_13_197_1473_0, i_13_197_1722_0,
    i_13_197_1725_0, i_13_197_1726_0, i_13_197_1734_0, i_13_197_1785_0,
    i_13_197_1788_0, i_13_197_1789_0, i_13_197_1842_0, i_13_197_1849_0,
    i_13_197_1857_0, i_13_197_1883_0, i_13_197_1884_0, i_13_197_1887_0,
    i_13_197_1889_0, i_13_197_2004_0, i_13_197_2122_0, i_13_197_2145_0,
    i_13_197_2146_0, i_13_197_2175_0, i_13_197_2231_0, i_13_197_2299_0,
    i_13_197_2464_0, i_13_197_2543_0, i_13_197_2616_0, i_13_197_2649_0,
    i_13_197_2650_0, i_13_197_2695_0, i_13_197_2766_0, i_13_197_2847_0,
    i_13_197_2851_0, i_13_197_2861_0, i_13_197_2877_0, i_13_197_3039_0,
    i_13_197_3067_0, i_13_197_3095_0, i_13_197_3103_0, i_13_197_3129_0,
    i_13_197_3148_0, i_13_197_3165_0, i_13_197_3173_0, i_13_197_3292_0,
    i_13_197_3391_0, i_13_197_3423_0, i_13_197_3427_0, i_13_197_3432_0,
    i_13_197_3472_0, i_13_197_3507_0, i_13_197_3534_0, i_13_197_3607_0,
    i_13_197_3688_0, i_13_197_3706_0, i_13_197_3796_0, i_13_197_3852_0,
    i_13_197_3869_0, i_13_197_3912_0, i_13_197_4017_0, i_13_197_4063_0,
    i_13_197_4094_0, i_13_197_4110_0, i_13_197_4188_0, i_13_197_4220_0,
    i_13_197_4256_0, i_13_197_4309_0, i_13_197_4315_0, i_13_197_4333_0,
    i_13_197_4381_0, i_13_197_4417_0, i_13_197_4593_0, i_13_197_4597_0,
    o_13_197_0_0  );
  input  i_13_197_41_0, i_13_197_71_0, i_13_197_138_0, i_13_197_139_0,
    i_13_197_141_0, i_13_197_142_0, i_13_197_231_0, i_13_197_232_0,
    i_13_197_310_0, i_13_197_418_0, i_13_197_471_0, i_13_197_472_0,
    i_13_197_517_0, i_13_197_537_0, i_13_197_538_0, i_13_197_764_0,
    i_13_197_826_0, i_13_197_832_0, i_13_197_1029_0, i_13_197_1086_0,
    i_13_197_1214_0, i_13_197_1218_0, i_13_197_1219_0, i_13_197_1221_0,
    i_13_197_1222_0, i_13_197_1266_0, i_13_197_1276_0, i_13_197_1362_0,
    i_13_197_1392_0, i_13_197_1426_0, i_13_197_1473_0, i_13_197_1722_0,
    i_13_197_1725_0, i_13_197_1726_0, i_13_197_1734_0, i_13_197_1785_0,
    i_13_197_1788_0, i_13_197_1789_0, i_13_197_1842_0, i_13_197_1849_0,
    i_13_197_1857_0, i_13_197_1883_0, i_13_197_1884_0, i_13_197_1887_0,
    i_13_197_1889_0, i_13_197_2004_0, i_13_197_2122_0, i_13_197_2145_0,
    i_13_197_2146_0, i_13_197_2175_0, i_13_197_2231_0, i_13_197_2299_0,
    i_13_197_2464_0, i_13_197_2543_0, i_13_197_2616_0, i_13_197_2649_0,
    i_13_197_2650_0, i_13_197_2695_0, i_13_197_2766_0, i_13_197_2847_0,
    i_13_197_2851_0, i_13_197_2861_0, i_13_197_2877_0, i_13_197_3039_0,
    i_13_197_3067_0, i_13_197_3095_0, i_13_197_3103_0, i_13_197_3129_0,
    i_13_197_3148_0, i_13_197_3165_0, i_13_197_3173_0, i_13_197_3292_0,
    i_13_197_3391_0, i_13_197_3423_0, i_13_197_3427_0, i_13_197_3432_0,
    i_13_197_3472_0, i_13_197_3507_0, i_13_197_3534_0, i_13_197_3607_0,
    i_13_197_3688_0, i_13_197_3706_0, i_13_197_3796_0, i_13_197_3852_0,
    i_13_197_3869_0, i_13_197_3912_0, i_13_197_4017_0, i_13_197_4063_0,
    i_13_197_4094_0, i_13_197_4110_0, i_13_197_4188_0, i_13_197_4220_0,
    i_13_197_4256_0, i_13_197_4309_0, i_13_197_4315_0, i_13_197_4333_0,
    i_13_197_4381_0, i_13_197_4417_0, i_13_197_4593_0, i_13_197_4597_0;
  output o_13_197_0_0;
  assign o_13_197_0_0 = ~((~i_13_197_538_0 & ((~i_13_197_1086_0 & ~i_13_197_1276_0) | (~i_13_197_141_0 & ~i_13_197_231_0 & ~i_13_197_1218_0 & ~i_13_197_4381_0))) | (~i_13_197_142_0 & ~i_13_197_537_0 & ~i_13_197_2616_0) | (i_13_197_2695_0 & ~i_13_197_3391_0 & i_13_197_4315_0 & i_13_197_4417_0) | (~i_13_197_1222_0 & ~i_13_197_1426_0 & ~i_13_197_1887_0 & ~i_13_197_4417_0));
endmodule



// Benchmark "kernel_13_198" written by ABC on Sun Jul 19 10:48:10 2020

module kernel_13_198 ( 
    i_13_198_79_0, i_13_198_95_0, i_13_198_140_0, i_13_198_187_0,
    i_13_198_275_0, i_13_198_322_0, i_13_198_328_0, i_13_198_329_0,
    i_13_198_365_0, i_13_198_370_0, i_13_198_431_0, i_13_198_445_0,
    i_13_198_511_0, i_13_198_562_0, i_13_198_599_0, i_13_198_602_0,
    i_13_198_610_0, i_13_198_674_0, i_13_198_718_0, i_13_198_728_0,
    i_13_198_781_0, i_13_198_832_0, i_13_198_861_0, i_13_198_862_0,
    i_13_198_895_0, i_13_198_1023_0, i_13_198_1078_0, i_13_198_1096_0,
    i_13_198_1195_0, i_13_198_1258_0, i_13_198_1321_0, i_13_198_1343_0,
    i_13_198_1384_0, i_13_198_1516_0, i_13_198_1637_0, i_13_198_1687_0,
    i_13_198_1726_0, i_13_198_1751_0, i_13_198_1768_0, i_13_198_1849_0,
    i_13_198_1859_0, i_13_198_1886_0, i_13_198_1888_0, i_13_198_1907_0,
    i_13_198_1913_0, i_13_198_1954_0, i_13_198_2101_0, i_13_198_2123_0,
    i_13_198_2168_0, i_13_198_2290_0, i_13_198_2311_0, i_13_198_2399_0,
    i_13_198_2428_0, i_13_198_2462_0, i_13_198_2492_0, i_13_198_2633_0,
    i_13_198_2650_0, i_13_198_2651_0, i_13_198_2653_0, i_13_198_2654_0,
    i_13_198_2722_0, i_13_198_2852_0, i_13_198_2884_0, i_13_198_2887_0,
    i_13_198_2922_0, i_13_198_2941_0, i_13_198_2942_0, i_13_198_2983_0,
    i_13_198_3023_0, i_13_198_3056_0, i_13_198_3127_0, i_13_198_3146_0,
    i_13_198_3154_0, i_13_198_3172_0, i_13_198_3173_0, i_13_198_3175_0,
    i_13_198_3176_0, i_13_198_3235_0, i_13_198_3238_0, i_13_198_3392_0,
    i_13_198_3433_0, i_13_198_3544_0, i_13_198_3563_0, i_13_198_3732_0,
    i_13_198_3785_0, i_13_198_3794_0, i_13_198_3847_0, i_13_198_3876_0,
    i_13_198_3913_0, i_13_198_3914_0, i_13_198_3965_0, i_13_198_4021_0,
    i_13_198_4100_0, i_13_198_4162_0, i_13_198_4238_0, i_13_198_4342_0,
    i_13_198_4382_0, i_13_198_4409_0, i_13_198_4444_0, i_13_198_4513_0,
    o_13_198_0_0  );
  input  i_13_198_79_0, i_13_198_95_0, i_13_198_140_0, i_13_198_187_0,
    i_13_198_275_0, i_13_198_322_0, i_13_198_328_0, i_13_198_329_0,
    i_13_198_365_0, i_13_198_370_0, i_13_198_431_0, i_13_198_445_0,
    i_13_198_511_0, i_13_198_562_0, i_13_198_599_0, i_13_198_602_0,
    i_13_198_610_0, i_13_198_674_0, i_13_198_718_0, i_13_198_728_0,
    i_13_198_781_0, i_13_198_832_0, i_13_198_861_0, i_13_198_862_0,
    i_13_198_895_0, i_13_198_1023_0, i_13_198_1078_0, i_13_198_1096_0,
    i_13_198_1195_0, i_13_198_1258_0, i_13_198_1321_0, i_13_198_1343_0,
    i_13_198_1384_0, i_13_198_1516_0, i_13_198_1637_0, i_13_198_1687_0,
    i_13_198_1726_0, i_13_198_1751_0, i_13_198_1768_0, i_13_198_1849_0,
    i_13_198_1859_0, i_13_198_1886_0, i_13_198_1888_0, i_13_198_1907_0,
    i_13_198_1913_0, i_13_198_1954_0, i_13_198_2101_0, i_13_198_2123_0,
    i_13_198_2168_0, i_13_198_2290_0, i_13_198_2311_0, i_13_198_2399_0,
    i_13_198_2428_0, i_13_198_2462_0, i_13_198_2492_0, i_13_198_2633_0,
    i_13_198_2650_0, i_13_198_2651_0, i_13_198_2653_0, i_13_198_2654_0,
    i_13_198_2722_0, i_13_198_2852_0, i_13_198_2884_0, i_13_198_2887_0,
    i_13_198_2922_0, i_13_198_2941_0, i_13_198_2942_0, i_13_198_2983_0,
    i_13_198_3023_0, i_13_198_3056_0, i_13_198_3127_0, i_13_198_3146_0,
    i_13_198_3154_0, i_13_198_3172_0, i_13_198_3173_0, i_13_198_3175_0,
    i_13_198_3176_0, i_13_198_3235_0, i_13_198_3238_0, i_13_198_3392_0,
    i_13_198_3433_0, i_13_198_3544_0, i_13_198_3563_0, i_13_198_3732_0,
    i_13_198_3785_0, i_13_198_3794_0, i_13_198_3847_0, i_13_198_3876_0,
    i_13_198_3913_0, i_13_198_3914_0, i_13_198_3965_0, i_13_198_4021_0,
    i_13_198_4100_0, i_13_198_4162_0, i_13_198_4238_0, i_13_198_4342_0,
    i_13_198_4382_0, i_13_198_4409_0, i_13_198_4444_0, i_13_198_4513_0;
  output o_13_198_0_0;
  assign o_13_198_0_0 = ~((~i_13_198_895_0 & (i_13_198_2887_0 | (~i_13_198_3176_0 & i_13_198_3847_0))) | (~i_13_198_1078_0 & ~i_13_198_2942_0) | (~i_13_198_2651_0 & ~i_13_198_3175_0) | (~i_13_198_2653_0 & ~i_13_198_3914_0));
endmodule



// Benchmark "kernel_13_199" written by ABC on Sun Jul 19 10:48:11 2020

module kernel_13_199 ( 
    i_13_199_74_0, i_13_199_121_0, i_13_199_122_0, i_13_199_125_0,
    i_13_199_142_0, i_13_199_175_0, i_13_199_176_0, i_13_199_227_0,
    i_13_199_229_0, i_13_199_311_0, i_13_199_338_0, i_13_199_341_0,
    i_13_199_517_0, i_13_199_524_0, i_13_199_533_0, i_13_199_535_0,
    i_13_199_536_0, i_13_199_596_0, i_13_199_599_0, i_13_199_617_0,
    i_13_199_766_0, i_13_199_830_0, i_13_199_850_0, i_13_199_911_0,
    i_13_199_977_0, i_13_199_1084_0, i_13_199_1085_0, i_13_199_1093_0,
    i_13_199_1139_0, i_13_199_1216_0, i_13_199_1433_0, i_13_199_1469_0,
    i_13_199_1496_0, i_13_199_1597_0, i_13_199_1598_0, i_13_199_1622_0,
    i_13_199_1721_0, i_13_199_1741_0, i_13_199_1757_0, i_13_199_1783_0,
    i_13_199_1784_0, i_13_199_1814_0, i_13_199_1817_0, i_13_199_1958_0,
    i_13_199_2012_0, i_13_199_2021_0, i_13_199_2120_0, i_13_199_2168_0,
    i_13_199_2210_0, i_13_199_2225_0, i_13_199_2309_0, i_13_199_2341_0,
    i_13_199_2432_0, i_13_199_2458_0, i_13_199_2462_0, i_13_199_2465_0,
    i_13_199_2500_0, i_13_199_2612_0, i_13_199_2630_0, i_13_199_2657_0,
    i_13_199_2714_0, i_13_199_2738_0, i_13_199_2818_0, i_13_199_2824_0,
    i_13_199_2885_0, i_13_199_3010_0, i_13_199_3019_0, i_13_199_3035_0,
    i_13_199_3037_0, i_13_199_3044_0, i_13_199_3128_0, i_13_199_3143_0,
    i_13_199_3169_0, i_13_199_3215_0, i_13_199_3217_0, i_13_199_3218_0,
    i_13_199_3221_0, i_13_199_3290_0, i_13_199_3413_0, i_13_199_3416_0,
    i_13_199_3449_0, i_13_199_3452_0, i_13_199_3524_0, i_13_199_3527_0,
    i_13_199_3737_0, i_13_199_3854_0, i_13_199_3865_0, i_13_199_3884_0,
    i_13_199_3998_0, i_13_199_4036_0, i_13_199_4055_0, i_13_199_4097_0,
    i_13_199_4238_0, i_13_199_4391_0, i_13_199_4414_0, i_13_199_4415_0,
    i_13_199_4519_0, i_13_199_4520_0, i_13_199_4523_0, i_13_199_4538_0,
    o_13_199_0_0  );
  input  i_13_199_74_0, i_13_199_121_0, i_13_199_122_0, i_13_199_125_0,
    i_13_199_142_0, i_13_199_175_0, i_13_199_176_0, i_13_199_227_0,
    i_13_199_229_0, i_13_199_311_0, i_13_199_338_0, i_13_199_341_0,
    i_13_199_517_0, i_13_199_524_0, i_13_199_533_0, i_13_199_535_0,
    i_13_199_536_0, i_13_199_596_0, i_13_199_599_0, i_13_199_617_0,
    i_13_199_766_0, i_13_199_830_0, i_13_199_850_0, i_13_199_911_0,
    i_13_199_977_0, i_13_199_1084_0, i_13_199_1085_0, i_13_199_1093_0,
    i_13_199_1139_0, i_13_199_1216_0, i_13_199_1433_0, i_13_199_1469_0,
    i_13_199_1496_0, i_13_199_1597_0, i_13_199_1598_0, i_13_199_1622_0,
    i_13_199_1721_0, i_13_199_1741_0, i_13_199_1757_0, i_13_199_1783_0,
    i_13_199_1784_0, i_13_199_1814_0, i_13_199_1817_0, i_13_199_1958_0,
    i_13_199_2012_0, i_13_199_2021_0, i_13_199_2120_0, i_13_199_2168_0,
    i_13_199_2210_0, i_13_199_2225_0, i_13_199_2309_0, i_13_199_2341_0,
    i_13_199_2432_0, i_13_199_2458_0, i_13_199_2462_0, i_13_199_2465_0,
    i_13_199_2500_0, i_13_199_2612_0, i_13_199_2630_0, i_13_199_2657_0,
    i_13_199_2714_0, i_13_199_2738_0, i_13_199_2818_0, i_13_199_2824_0,
    i_13_199_2885_0, i_13_199_3010_0, i_13_199_3019_0, i_13_199_3035_0,
    i_13_199_3037_0, i_13_199_3044_0, i_13_199_3128_0, i_13_199_3143_0,
    i_13_199_3169_0, i_13_199_3215_0, i_13_199_3217_0, i_13_199_3218_0,
    i_13_199_3221_0, i_13_199_3290_0, i_13_199_3413_0, i_13_199_3416_0,
    i_13_199_3449_0, i_13_199_3452_0, i_13_199_3524_0, i_13_199_3527_0,
    i_13_199_3737_0, i_13_199_3854_0, i_13_199_3865_0, i_13_199_3884_0,
    i_13_199_3998_0, i_13_199_4036_0, i_13_199_4055_0, i_13_199_4097_0,
    i_13_199_4238_0, i_13_199_4391_0, i_13_199_4414_0, i_13_199_4415_0,
    i_13_199_4519_0, i_13_199_4520_0, i_13_199_4523_0, i_13_199_4538_0;
  output o_13_199_0_0;
  assign o_13_199_0_0 = ~((~i_13_199_533_0 & (~i_13_199_3218_0 | (~i_13_199_1814_0 & ~i_13_199_2738_0 & ~i_13_199_4415_0))) | (i_13_199_311_0 & ~i_13_199_338_0) | (~i_13_199_1469_0 & ~i_13_199_2738_0 & i_13_199_3010_0) | (i_13_199_176_0 & ~i_13_199_1085_0 & ~i_13_199_3169_0 & ~i_13_199_3215_0) | (~i_13_199_1622_0 & ~i_13_199_2885_0 & ~i_13_199_3143_0 & i_13_199_4036_0) | (~i_13_199_122_0 & ~i_13_199_4414_0));
endmodule



// Benchmark "kernel_13_200" written by ABC on Sun Jul 19 10:48:12 2020

module kernel_13_200 ( 
    i_13_200_31_0, i_13_200_271_0, i_13_200_273_0, i_13_200_274_0,
    i_13_200_275_0, i_13_200_279_0, i_13_200_310_0, i_13_200_322_0,
    i_13_200_426_0, i_13_200_442_0, i_13_200_450_0, i_13_200_451_0,
    i_13_200_589_0, i_13_200_592_0, i_13_200_643_0, i_13_200_657_0,
    i_13_200_660_0, i_13_200_760_0, i_13_200_831_0, i_13_200_838_0,
    i_13_200_858_0, i_13_200_867_0, i_13_200_868_0, i_13_200_894_0,
    i_13_200_928_0, i_13_200_939_0, i_13_200_940_0, i_13_200_944_0,
    i_13_200_1017_0, i_13_200_1080_0, i_13_200_1081_0, i_13_200_1148_0,
    i_13_200_1150_0, i_13_200_1444_0, i_13_200_1470_0, i_13_200_1492_0,
    i_13_200_1497_0, i_13_200_1597_0, i_13_200_1632_0, i_13_200_1642_0,
    i_13_200_1733_0, i_13_200_1750_0, i_13_200_1765_0, i_13_200_1854_0,
    i_13_200_1947_0, i_13_200_2011_0, i_13_200_2140_0, i_13_200_2191_0,
    i_13_200_2226_0, i_13_200_2233_0, i_13_200_2380_0, i_13_200_2421_0,
    i_13_200_2449_0, i_13_200_2451_0, i_13_200_2467_0, i_13_200_2506_0,
    i_13_200_2541_0, i_13_200_2542_0, i_13_200_2544_0, i_13_200_2545_0,
    i_13_200_2568_0, i_13_200_2857_0, i_13_200_2884_0, i_13_200_2924_0,
    i_13_200_2955_0, i_13_200_3109_0, i_13_200_3142_0, i_13_200_3388_0,
    i_13_200_3414_0, i_13_200_3415_0, i_13_200_3451_0, i_13_200_3459_0,
    i_13_200_3460_0, i_13_200_3463_0, i_13_200_3475_0, i_13_200_3477_0,
    i_13_200_3486_0, i_13_200_3549_0, i_13_200_3567_0, i_13_200_3570_0,
    i_13_200_3576_0, i_13_200_3627_0, i_13_200_3900_0, i_13_200_3919_0,
    i_13_200_3928_0, i_13_200_3991_0, i_13_200_4054_0, i_13_200_4086_0,
    i_13_200_4162_0, i_13_200_4166_0, i_13_200_4265_0, i_13_200_4266_0,
    i_13_200_4368_0, i_13_200_4369_0, i_13_200_4433_0, i_13_200_4514_0,
    i_13_200_4537_0, i_13_200_4554_0, i_13_200_4555_0, i_13_200_4593_0,
    o_13_200_0_0  );
  input  i_13_200_31_0, i_13_200_271_0, i_13_200_273_0, i_13_200_274_0,
    i_13_200_275_0, i_13_200_279_0, i_13_200_310_0, i_13_200_322_0,
    i_13_200_426_0, i_13_200_442_0, i_13_200_450_0, i_13_200_451_0,
    i_13_200_589_0, i_13_200_592_0, i_13_200_643_0, i_13_200_657_0,
    i_13_200_660_0, i_13_200_760_0, i_13_200_831_0, i_13_200_838_0,
    i_13_200_858_0, i_13_200_867_0, i_13_200_868_0, i_13_200_894_0,
    i_13_200_928_0, i_13_200_939_0, i_13_200_940_0, i_13_200_944_0,
    i_13_200_1017_0, i_13_200_1080_0, i_13_200_1081_0, i_13_200_1148_0,
    i_13_200_1150_0, i_13_200_1444_0, i_13_200_1470_0, i_13_200_1492_0,
    i_13_200_1497_0, i_13_200_1597_0, i_13_200_1632_0, i_13_200_1642_0,
    i_13_200_1733_0, i_13_200_1750_0, i_13_200_1765_0, i_13_200_1854_0,
    i_13_200_1947_0, i_13_200_2011_0, i_13_200_2140_0, i_13_200_2191_0,
    i_13_200_2226_0, i_13_200_2233_0, i_13_200_2380_0, i_13_200_2421_0,
    i_13_200_2449_0, i_13_200_2451_0, i_13_200_2467_0, i_13_200_2506_0,
    i_13_200_2541_0, i_13_200_2542_0, i_13_200_2544_0, i_13_200_2545_0,
    i_13_200_2568_0, i_13_200_2857_0, i_13_200_2884_0, i_13_200_2924_0,
    i_13_200_2955_0, i_13_200_3109_0, i_13_200_3142_0, i_13_200_3388_0,
    i_13_200_3414_0, i_13_200_3415_0, i_13_200_3451_0, i_13_200_3459_0,
    i_13_200_3460_0, i_13_200_3463_0, i_13_200_3475_0, i_13_200_3477_0,
    i_13_200_3486_0, i_13_200_3549_0, i_13_200_3567_0, i_13_200_3570_0,
    i_13_200_3576_0, i_13_200_3627_0, i_13_200_3900_0, i_13_200_3919_0,
    i_13_200_3928_0, i_13_200_3991_0, i_13_200_4054_0, i_13_200_4086_0,
    i_13_200_4162_0, i_13_200_4166_0, i_13_200_4265_0, i_13_200_4266_0,
    i_13_200_4368_0, i_13_200_4369_0, i_13_200_4433_0, i_13_200_4514_0,
    i_13_200_4537_0, i_13_200_4554_0, i_13_200_4555_0, i_13_200_4593_0;
  output o_13_200_0_0;
  assign o_13_200_0_0 = ~((~i_13_200_940_0 & ((~i_13_200_3460_0 & ~i_13_200_3486_0 & ~i_13_200_3549_0) | (~i_13_200_944_0 & ~i_13_200_1080_0 & ~i_13_200_1854_0 & ~i_13_200_3570_0))) | (i_13_200_4514_0 & (~i_13_200_274_0 | (~i_13_200_275_0 & i_13_200_1642_0) | (i_13_200_592_0 & i_13_200_2380_0))) | (~i_13_200_2542_0 & ~i_13_200_2545_0 & ~i_13_200_4086_0) | (~i_13_200_271_0 & ~i_13_200_2924_0 & i_13_200_4433_0) | (i_13_200_275_0 & ~i_13_200_4162_0 & ~i_13_200_4514_0));
endmodule



// Benchmark "kernel_13_201" written by ABC on Sun Jul 19 10:48:13 2020

module kernel_13_201 ( 
    i_13_201_38_0, i_13_201_92_0, i_13_201_95_0, i_13_201_107_0,
    i_13_201_113_0, i_13_201_118_0, i_13_201_274_0, i_13_201_361_0,
    i_13_201_406_0, i_13_201_407_0, i_13_201_446_0, i_13_201_448_0,
    i_13_201_449_0, i_13_201_562_0, i_13_201_565_0, i_13_201_572_0,
    i_13_201_607_0, i_13_201_608_0, i_13_201_610_0, i_13_201_733_0,
    i_13_201_796_0, i_13_201_797_0, i_13_201_895_0, i_13_201_949_0,
    i_13_201_950_0, i_13_201_952_0, i_13_201_1034_0, i_13_201_1084_0,
    i_13_201_1087_0, i_13_201_1096_0, i_13_201_1186_0, i_13_201_1244_0,
    i_13_201_1253_0, i_13_201_1262_0, i_13_201_1409_0, i_13_201_1432_0,
    i_13_201_1441_0, i_13_201_1510_0, i_13_201_1541_0, i_13_201_1589_0,
    i_13_201_1633_0, i_13_201_1730_0, i_13_201_1750_0, i_13_201_1765_0,
    i_13_201_1787_0, i_13_201_1832_0, i_13_201_1841_0, i_13_201_1885_0,
    i_13_201_1954_0, i_13_201_2003_0, i_13_201_2120_0, i_13_201_2137_0,
    i_13_201_2173_0, i_13_201_2174_0, i_13_201_2177_0, i_13_201_2209_0,
    i_13_201_2435_0, i_13_201_2498_0, i_13_201_2564_0, i_13_201_2702_0,
    i_13_201_2875_0, i_13_201_2939_0, i_13_201_3035_0, i_13_201_3044_0,
    i_13_201_3047_0, i_13_201_3101_0, i_13_201_3104_0, i_13_201_3161_0,
    i_13_201_3163_0, i_13_201_3164_0, i_13_201_3209_0, i_13_201_3235_0,
    i_13_201_3344_0, i_13_201_3511_0, i_13_201_3703_0, i_13_201_3764_0,
    i_13_201_3803_0, i_13_201_3844_0, i_13_201_3847_0, i_13_201_3871_0,
    i_13_201_3872_0, i_13_201_3874_0, i_13_201_3875_0, i_13_201_3979_0,
    i_13_201_3980_0, i_13_201_4010_0, i_13_201_4081_0, i_13_201_4090_0,
    i_13_201_4118_0, i_13_201_4120_0, i_13_201_4121_0, i_13_201_4162_0,
    i_13_201_4163_0, i_13_201_4349_0, i_13_201_4351_0, i_13_201_4352_0,
    i_13_201_4354_0, i_13_201_4541_0, i_13_201_4568_0, i_13_201_4598_0,
    o_13_201_0_0  );
  input  i_13_201_38_0, i_13_201_92_0, i_13_201_95_0, i_13_201_107_0,
    i_13_201_113_0, i_13_201_118_0, i_13_201_274_0, i_13_201_361_0,
    i_13_201_406_0, i_13_201_407_0, i_13_201_446_0, i_13_201_448_0,
    i_13_201_449_0, i_13_201_562_0, i_13_201_565_0, i_13_201_572_0,
    i_13_201_607_0, i_13_201_608_0, i_13_201_610_0, i_13_201_733_0,
    i_13_201_796_0, i_13_201_797_0, i_13_201_895_0, i_13_201_949_0,
    i_13_201_950_0, i_13_201_952_0, i_13_201_1034_0, i_13_201_1084_0,
    i_13_201_1087_0, i_13_201_1096_0, i_13_201_1186_0, i_13_201_1244_0,
    i_13_201_1253_0, i_13_201_1262_0, i_13_201_1409_0, i_13_201_1432_0,
    i_13_201_1441_0, i_13_201_1510_0, i_13_201_1541_0, i_13_201_1589_0,
    i_13_201_1633_0, i_13_201_1730_0, i_13_201_1750_0, i_13_201_1765_0,
    i_13_201_1787_0, i_13_201_1832_0, i_13_201_1841_0, i_13_201_1885_0,
    i_13_201_1954_0, i_13_201_2003_0, i_13_201_2120_0, i_13_201_2137_0,
    i_13_201_2173_0, i_13_201_2174_0, i_13_201_2177_0, i_13_201_2209_0,
    i_13_201_2435_0, i_13_201_2498_0, i_13_201_2564_0, i_13_201_2702_0,
    i_13_201_2875_0, i_13_201_2939_0, i_13_201_3035_0, i_13_201_3044_0,
    i_13_201_3047_0, i_13_201_3101_0, i_13_201_3104_0, i_13_201_3161_0,
    i_13_201_3163_0, i_13_201_3164_0, i_13_201_3209_0, i_13_201_3235_0,
    i_13_201_3344_0, i_13_201_3511_0, i_13_201_3703_0, i_13_201_3764_0,
    i_13_201_3803_0, i_13_201_3844_0, i_13_201_3847_0, i_13_201_3871_0,
    i_13_201_3872_0, i_13_201_3874_0, i_13_201_3875_0, i_13_201_3979_0,
    i_13_201_3980_0, i_13_201_4010_0, i_13_201_4081_0, i_13_201_4090_0,
    i_13_201_4118_0, i_13_201_4120_0, i_13_201_4121_0, i_13_201_4162_0,
    i_13_201_4163_0, i_13_201_4349_0, i_13_201_4351_0, i_13_201_4352_0,
    i_13_201_4354_0, i_13_201_4541_0, i_13_201_4568_0, i_13_201_4598_0;
  output o_13_201_0_0;
  assign o_13_201_0_0 = ~((~i_13_201_3161_0 & (i_13_201_895_0 | (~i_13_201_1885_0 & ~i_13_201_3104_0 & ~i_13_201_3163_0 & ~i_13_201_3874_0))) | (~i_13_201_95_0 & ~i_13_201_3101_0) | (~i_13_201_113_0 & ~i_13_201_274_0 & ~i_13_201_4349_0) | (~i_13_201_4163_0 & ~i_13_201_4352_0) | (~i_13_201_2003_0 & ~i_13_201_2177_0 & ~i_13_201_3235_0 & i_13_201_4354_0));
endmodule



// Benchmark "kernel_13_202" written by ABC on Sun Jul 19 10:48:14 2020

module kernel_13_202 ( 
    i_13_202_112_0, i_13_202_131_0, i_13_202_133_0, i_13_202_134_0,
    i_13_202_160_0, i_13_202_169_0, i_13_202_170_0, i_13_202_358_0,
    i_13_202_457_0, i_13_202_466_0, i_13_202_664_0, i_13_202_799_0,
    i_13_202_831_0, i_13_202_853_0, i_13_202_956_0, i_13_202_959_0,
    i_13_202_1078_0, i_13_202_1132_0, i_13_202_1231_0, i_13_202_1303_0,
    i_13_202_1310_0, i_13_202_1364_0, i_13_202_1400_0, i_13_202_1407_0,
    i_13_202_1446_0, i_13_202_1447_0, i_13_202_1471_0, i_13_202_1501_0,
    i_13_202_1507_0, i_13_202_1555_0, i_13_202_1556_0, i_13_202_1639_0,
    i_13_202_1699_0, i_13_202_1847_0, i_13_202_1849_0, i_13_202_1850_0,
    i_13_202_1896_0, i_13_202_1930_0, i_13_202_1961_0, i_13_202_2103_0,
    i_13_202_2104_0, i_13_202_2111_0, i_13_202_2143_0, i_13_202_2145_0,
    i_13_202_2146_0, i_13_202_2156_0, i_13_202_2202_0, i_13_202_2203_0,
    i_13_202_2204_0, i_13_202_2209_0, i_13_202_2237_0, i_13_202_2398_0,
    i_13_202_2407_0, i_13_202_2428_0, i_13_202_2429_0, i_13_202_2595_0,
    i_13_202_2681_0, i_13_202_2882_0, i_13_202_2936_0, i_13_202_2938_0,
    i_13_202_2939_0, i_13_202_2986_0, i_13_202_3028_0, i_13_202_3101_0,
    i_13_202_3146_0, i_13_202_3232_0, i_13_202_3242_0, i_13_202_3244_0,
    i_13_202_3245_0, i_13_202_3341_0, i_13_202_3406_0, i_13_202_3410_0,
    i_13_202_3637_0, i_13_202_3638_0, i_13_202_3644_0, i_13_202_3739_0,
    i_13_202_3755_0, i_13_202_3757_0, i_13_202_3758_0, i_13_202_3805_0,
    i_13_202_3812_0, i_13_202_3859_0, i_13_202_3860_0, i_13_202_3919_0,
    i_13_202_3935_0, i_13_202_4054_0, i_13_202_4061_0, i_13_202_4063_0,
    i_13_202_4214_0, i_13_202_4220_0, i_13_202_4270_0, i_13_202_4273_0,
    i_13_202_4313_0, i_13_202_4316_0, i_13_202_4423_0, i_13_202_4432_0,
    i_13_202_4453_0, i_13_202_4481_0, i_13_202_4510_0, i_13_202_4512_0,
    o_13_202_0_0  );
  input  i_13_202_112_0, i_13_202_131_0, i_13_202_133_0, i_13_202_134_0,
    i_13_202_160_0, i_13_202_169_0, i_13_202_170_0, i_13_202_358_0,
    i_13_202_457_0, i_13_202_466_0, i_13_202_664_0, i_13_202_799_0,
    i_13_202_831_0, i_13_202_853_0, i_13_202_956_0, i_13_202_959_0,
    i_13_202_1078_0, i_13_202_1132_0, i_13_202_1231_0, i_13_202_1303_0,
    i_13_202_1310_0, i_13_202_1364_0, i_13_202_1400_0, i_13_202_1407_0,
    i_13_202_1446_0, i_13_202_1447_0, i_13_202_1471_0, i_13_202_1501_0,
    i_13_202_1507_0, i_13_202_1555_0, i_13_202_1556_0, i_13_202_1639_0,
    i_13_202_1699_0, i_13_202_1847_0, i_13_202_1849_0, i_13_202_1850_0,
    i_13_202_1896_0, i_13_202_1930_0, i_13_202_1961_0, i_13_202_2103_0,
    i_13_202_2104_0, i_13_202_2111_0, i_13_202_2143_0, i_13_202_2145_0,
    i_13_202_2146_0, i_13_202_2156_0, i_13_202_2202_0, i_13_202_2203_0,
    i_13_202_2204_0, i_13_202_2209_0, i_13_202_2237_0, i_13_202_2398_0,
    i_13_202_2407_0, i_13_202_2428_0, i_13_202_2429_0, i_13_202_2595_0,
    i_13_202_2681_0, i_13_202_2882_0, i_13_202_2936_0, i_13_202_2938_0,
    i_13_202_2939_0, i_13_202_2986_0, i_13_202_3028_0, i_13_202_3101_0,
    i_13_202_3146_0, i_13_202_3232_0, i_13_202_3242_0, i_13_202_3244_0,
    i_13_202_3245_0, i_13_202_3341_0, i_13_202_3406_0, i_13_202_3410_0,
    i_13_202_3637_0, i_13_202_3638_0, i_13_202_3644_0, i_13_202_3739_0,
    i_13_202_3755_0, i_13_202_3757_0, i_13_202_3758_0, i_13_202_3805_0,
    i_13_202_3812_0, i_13_202_3859_0, i_13_202_3860_0, i_13_202_3919_0,
    i_13_202_3935_0, i_13_202_4054_0, i_13_202_4061_0, i_13_202_4063_0,
    i_13_202_4214_0, i_13_202_4220_0, i_13_202_4270_0, i_13_202_4273_0,
    i_13_202_4313_0, i_13_202_4316_0, i_13_202_4423_0, i_13_202_4432_0,
    i_13_202_4453_0, i_13_202_4481_0, i_13_202_4510_0, i_13_202_4512_0;
  output o_13_202_0_0;
  assign o_13_202_0_0 = ~((~i_13_202_358_0 & ~i_13_202_4316_0) | (~i_13_202_466_0 & ~i_13_202_3245_0 & ~i_13_202_4313_0) | (~i_13_202_1556_0 & ~i_13_202_2204_0 & ~i_13_202_2938_0));
endmodule



// Benchmark "kernel_13_203" written by ABC on Sun Jul 19 10:48:14 2020

module kernel_13_203 ( 
    i_13_203_28_0, i_13_203_64_0, i_13_203_65_0, i_13_203_74_0,
    i_13_203_308_0, i_13_203_355_0, i_13_203_442_0, i_13_203_443_0,
    i_13_203_445_0, i_13_203_446_0, i_13_203_667_0, i_13_203_668_0,
    i_13_203_676_0, i_13_203_677_0, i_13_203_743_0, i_13_203_829_0,
    i_13_203_931_0, i_13_203_947_0, i_13_203_1081_0, i_13_203_1099_0,
    i_13_203_1100_0, i_13_203_1102_0, i_13_203_1274_0, i_13_203_1279_0,
    i_13_203_1306_0, i_13_203_1307_0, i_13_203_1397_0, i_13_203_1424_0,
    i_13_203_1435_0, i_13_203_1444_0, i_13_203_1499_0, i_13_203_1504_0,
    i_13_203_1505_0, i_13_203_1594_0, i_13_203_1595_0, i_13_203_1621_0,
    i_13_203_1634_0, i_13_203_1639_0, i_13_203_1642_0, i_13_203_1723_0,
    i_13_203_1768_0, i_13_203_1773_0, i_13_203_1774_0, i_13_203_1783_0,
    i_13_203_1793_0, i_13_203_1838_0, i_13_203_1847_0, i_13_203_1903_0,
    i_13_203_1921_0, i_13_203_1957_0, i_13_203_1958_0, i_13_203_1993_0,
    i_13_203_2002_0, i_13_203_2030_0, i_13_203_2200_0, i_13_203_2209_0,
    i_13_203_2317_0, i_13_203_2468_0, i_13_203_2512_0, i_13_203_2567_0,
    i_13_203_2656_0, i_13_203_2673_0, i_13_203_2675_0, i_13_203_2999_0,
    i_13_203_3061_0, i_13_203_3065_0, i_13_203_3073_0, i_13_203_3089_0,
    i_13_203_3109_0, i_13_203_3127_0, i_13_203_3128_0, i_13_203_3242_0,
    i_13_203_3397_0, i_13_203_3448_0, i_13_203_3449_0, i_13_203_3524_0,
    i_13_203_3551_0, i_13_203_3574_0, i_13_203_3595_0, i_13_203_3596_0,
    i_13_203_3619_0, i_13_203_3646_0, i_13_203_3781_0, i_13_203_3782_0,
    i_13_203_3857_0, i_13_203_3863_0, i_13_203_3890_0, i_13_203_3924_0,
    i_13_203_3925_0, i_13_203_3988_0, i_13_203_4061_0, i_13_203_4078_0,
    i_13_203_4087_0, i_13_203_4330_0, i_13_203_4342_0, i_13_203_4430_0,
    i_13_203_4433_0, i_13_203_4447_0, i_13_203_4520_0, i_13_203_4556_0,
    o_13_203_0_0  );
  input  i_13_203_28_0, i_13_203_64_0, i_13_203_65_0, i_13_203_74_0,
    i_13_203_308_0, i_13_203_355_0, i_13_203_442_0, i_13_203_443_0,
    i_13_203_445_0, i_13_203_446_0, i_13_203_667_0, i_13_203_668_0,
    i_13_203_676_0, i_13_203_677_0, i_13_203_743_0, i_13_203_829_0,
    i_13_203_931_0, i_13_203_947_0, i_13_203_1081_0, i_13_203_1099_0,
    i_13_203_1100_0, i_13_203_1102_0, i_13_203_1274_0, i_13_203_1279_0,
    i_13_203_1306_0, i_13_203_1307_0, i_13_203_1397_0, i_13_203_1424_0,
    i_13_203_1435_0, i_13_203_1444_0, i_13_203_1499_0, i_13_203_1504_0,
    i_13_203_1505_0, i_13_203_1594_0, i_13_203_1595_0, i_13_203_1621_0,
    i_13_203_1634_0, i_13_203_1639_0, i_13_203_1642_0, i_13_203_1723_0,
    i_13_203_1768_0, i_13_203_1773_0, i_13_203_1774_0, i_13_203_1783_0,
    i_13_203_1793_0, i_13_203_1838_0, i_13_203_1847_0, i_13_203_1903_0,
    i_13_203_1921_0, i_13_203_1957_0, i_13_203_1958_0, i_13_203_1993_0,
    i_13_203_2002_0, i_13_203_2030_0, i_13_203_2200_0, i_13_203_2209_0,
    i_13_203_2317_0, i_13_203_2468_0, i_13_203_2512_0, i_13_203_2567_0,
    i_13_203_2656_0, i_13_203_2673_0, i_13_203_2675_0, i_13_203_2999_0,
    i_13_203_3061_0, i_13_203_3065_0, i_13_203_3073_0, i_13_203_3089_0,
    i_13_203_3109_0, i_13_203_3127_0, i_13_203_3128_0, i_13_203_3242_0,
    i_13_203_3397_0, i_13_203_3448_0, i_13_203_3449_0, i_13_203_3524_0,
    i_13_203_3551_0, i_13_203_3574_0, i_13_203_3595_0, i_13_203_3596_0,
    i_13_203_3619_0, i_13_203_3646_0, i_13_203_3781_0, i_13_203_3782_0,
    i_13_203_3857_0, i_13_203_3863_0, i_13_203_3890_0, i_13_203_3924_0,
    i_13_203_3925_0, i_13_203_3988_0, i_13_203_4061_0, i_13_203_4078_0,
    i_13_203_4087_0, i_13_203_4330_0, i_13_203_4342_0, i_13_203_4430_0,
    i_13_203_4433_0, i_13_203_4447_0, i_13_203_4520_0, i_13_203_4556_0;
  output o_13_203_0_0;
  assign o_13_203_0_0 = ~((i_13_203_445_0 & ((~i_13_203_2675_0 & ~i_13_203_3061_0) | (~i_13_203_2002_0 & ~i_13_203_4430_0))) | (~i_13_203_65_0 & ~i_13_203_677_0 & ~i_13_203_1504_0) | (~i_13_203_1595_0 & ~i_13_203_3619_0) | (i_13_203_1274_0 & ~i_13_203_1847_0 & ~i_13_203_4556_0));
endmodule



// Benchmark "kernel_13_204" written by ABC on Sun Jul 19 10:48:15 2020

module kernel_13_204 ( 
    i_13_204_163_0, i_13_204_173_0, i_13_204_175_0, i_13_204_176_0,
    i_13_204_177_0, i_13_204_178_0, i_13_204_280_0, i_13_204_307_0,
    i_13_204_379_0, i_13_204_380_0, i_13_204_452_0, i_13_204_526_0,
    i_13_204_527_0, i_13_204_617_0, i_13_204_625_0, i_13_204_735_0,
    i_13_204_742_0, i_13_204_766_0, i_13_204_797_0, i_13_204_814_0,
    i_13_204_817_0, i_13_204_829_0, i_13_204_976_0, i_13_204_977_0,
    i_13_204_1063_0, i_13_204_1076_0, i_13_204_1093_0, i_13_204_1094_0,
    i_13_204_1204_0, i_13_204_1297_0, i_13_204_1309_0, i_13_204_1319_0,
    i_13_204_1327_0, i_13_204_1442_0, i_13_204_1445_0, i_13_204_1446_0,
    i_13_204_1460_0, i_13_204_1498_0, i_13_204_1499_0, i_13_204_1502_0,
    i_13_204_1594_0, i_13_204_1595_0, i_13_204_1601_0, i_13_204_1687_0,
    i_13_204_1732_0, i_13_204_1846_0, i_13_204_1850_0, i_13_204_1927_0,
    i_13_204_1931_0, i_13_204_1990_0, i_13_204_2020_0, i_13_204_2119_0,
    i_13_204_2135_0, i_13_204_2191_0, i_13_204_2246_0, i_13_204_2264_0,
    i_13_204_2405_0, i_13_204_2413_0, i_13_204_2425_0, i_13_204_2431_0,
    i_13_204_2505_0, i_13_204_2578_0, i_13_204_2849_0, i_13_204_2875_0,
    i_13_204_2935_0, i_13_204_2938_0, i_13_204_3011_0, i_13_204_3053_0,
    i_13_204_3109_0, i_13_204_3110_0, i_13_204_3130_0, i_13_204_3244_0,
    i_13_204_3373_0, i_13_204_3399_0, i_13_204_3416_0, i_13_204_3421_0,
    i_13_204_3423_0, i_13_204_3425_0, i_13_204_3428_0, i_13_204_3437_0,
    i_13_204_3523_0, i_13_204_3649_0, i_13_204_3728_0, i_13_204_3731_0,
    i_13_204_3794_0, i_13_204_3865_0, i_13_204_4018_0, i_13_204_4019_0,
    i_13_204_4051_0, i_13_204_4060_0, i_13_204_4061_0, i_13_204_4063_0,
    i_13_204_4136_0, i_13_204_4267_0, i_13_204_4268_0, i_13_204_4306_0,
    i_13_204_4312_0, i_13_204_4314_0, i_13_204_4342_0, i_13_204_4568_0,
    o_13_204_0_0  );
  input  i_13_204_163_0, i_13_204_173_0, i_13_204_175_0, i_13_204_176_0,
    i_13_204_177_0, i_13_204_178_0, i_13_204_280_0, i_13_204_307_0,
    i_13_204_379_0, i_13_204_380_0, i_13_204_452_0, i_13_204_526_0,
    i_13_204_527_0, i_13_204_617_0, i_13_204_625_0, i_13_204_735_0,
    i_13_204_742_0, i_13_204_766_0, i_13_204_797_0, i_13_204_814_0,
    i_13_204_817_0, i_13_204_829_0, i_13_204_976_0, i_13_204_977_0,
    i_13_204_1063_0, i_13_204_1076_0, i_13_204_1093_0, i_13_204_1094_0,
    i_13_204_1204_0, i_13_204_1297_0, i_13_204_1309_0, i_13_204_1319_0,
    i_13_204_1327_0, i_13_204_1442_0, i_13_204_1445_0, i_13_204_1446_0,
    i_13_204_1460_0, i_13_204_1498_0, i_13_204_1499_0, i_13_204_1502_0,
    i_13_204_1594_0, i_13_204_1595_0, i_13_204_1601_0, i_13_204_1687_0,
    i_13_204_1732_0, i_13_204_1846_0, i_13_204_1850_0, i_13_204_1927_0,
    i_13_204_1931_0, i_13_204_1990_0, i_13_204_2020_0, i_13_204_2119_0,
    i_13_204_2135_0, i_13_204_2191_0, i_13_204_2246_0, i_13_204_2264_0,
    i_13_204_2405_0, i_13_204_2413_0, i_13_204_2425_0, i_13_204_2431_0,
    i_13_204_2505_0, i_13_204_2578_0, i_13_204_2849_0, i_13_204_2875_0,
    i_13_204_2935_0, i_13_204_2938_0, i_13_204_3011_0, i_13_204_3053_0,
    i_13_204_3109_0, i_13_204_3110_0, i_13_204_3130_0, i_13_204_3244_0,
    i_13_204_3373_0, i_13_204_3399_0, i_13_204_3416_0, i_13_204_3421_0,
    i_13_204_3423_0, i_13_204_3425_0, i_13_204_3428_0, i_13_204_3437_0,
    i_13_204_3523_0, i_13_204_3649_0, i_13_204_3728_0, i_13_204_3731_0,
    i_13_204_3794_0, i_13_204_3865_0, i_13_204_4018_0, i_13_204_4019_0,
    i_13_204_4051_0, i_13_204_4060_0, i_13_204_4061_0, i_13_204_4063_0,
    i_13_204_4136_0, i_13_204_4267_0, i_13_204_4268_0, i_13_204_4306_0,
    i_13_204_4312_0, i_13_204_4314_0, i_13_204_4342_0, i_13_204_4568_0;
  output o_13_204_0_0;
  assign o_13_204_0_0 = ~((~i_13_204_4061_0 & ((~i_13_204_280_0 & i_13_204_3523_0) | (~i_13_204_1063_0 & ~i_13_204_3731_0))) | (~i_13_204_4268_0 & ((i_13_204_617_0 & ~i_13_204_817_0) | (i_13_204_1319_0 & ~i_13_204_1846_0 & ~i_13_204_3011_0))) | (i_13_204_176_0 & i_13_204_1076_0 & ~i_13_204_2425_0 & ~i_13_204_4051_0) | (~i_13_204_1595_0 & ~i_13_204_4063_0) | (~i_13_204_3244_0 & i_13_204_4314_0));
endmodule



// Benchmark "kernel_13_205" written by ABC on Sun Jul 19 10:48:16 2020

module kernel_13_205 ( 
    i_13_205_31_0, i_13_205_184_0, i_13_205_196_0, i_13_205_259_0,
    i_13_205_325_0, i_13_205_327_0, i_13_205_328_0, i_13_205_382_0,
    i_13_205_526_0, i_13_205_624_0, i_13_205_660_0, i_13_205_661_0,
    i_13_205_742_0, i_13_205_820_0, i_13_205_840_0, i_13_205_850_0,
    i_13_205_852_0, i_13_205_854_0, i_13_205_858_0, i_13_205_861_0,
    i_13_205_1020_0, i_13_205_1074_0, i_13_205_1093_0, i_13_205_1097_0,
    i_13_205_1227_0, i_13_205_1228_0, i_13_205_1229_0, i_13_205_1254_0,
    i_13_205_1255_0, i_13_205_1256_0, i_13_205_1258_0, i_13_205_1314_0,
    i_13_205_1317_0, i_13_205_1383_0, i_13_205_1428_0, i_13_205_1443_0,
    i_13_205_1444_0, i_13_205_1447_0, i_13_205_1483_0, i_13_205_1488_0,
    i_13_205_1645_0, i_13_205_1675_0, i_13_205_1691_0, i_13_205_1753_0,
    i_13_205_1848_0, i_13_205_1849_0, i_13_205_1854_0, i_13_205_1857_0,
    i_13_205_1858_0, i_13_205_1861_0, i_13_205_1953_0, i_13_205_1957_0,
    i_13_205_1993_0, i_13_205_2042_0, i_13_205_2247_0, i_13_205_2248_0,
    i_13_205_2281_0, i_13_205_2394_0, i_13_205_2407_0, i_13_205_2412_0,
    i_13_205_2434_0, i_13_205_2488_0, i_13_205_2614_0, i_13_205_2617_0,
    i_13_205_2701_0, i_13_205_2712_0, i_13_205_2857_0, i_13_205_2878_0,
    i_13_205_2978_0, i_13_205_3064_0, i_13_205_3118_0, i_13_205_3122_0,
    i_13_205_3153_0, i_13_205_3172_0, i_13_205_3307_0, i_13_205_3338_0,
    i_13_205_3355_0, i_13_205_3418_0, i_13_205_3436_0, i_13_205_3456_0,
    i_13_205_3460_0, i_13_205_3478_0, i_13_205_3484_0, i_13_205_3486_0,
    i_13_205_3487_0, i_13_205_3489_0, i_13_205_3537_0, i_13_205_3562_0,
    i_13_205_3689_0, i_13_205_3783_0, i_13_205_3802_0, i_13_205_3868_0,
    i_13_205_3907_0, i_13_205_4063_0, i_13_205_4351_0, i_13_205_4365_0,
    i_13_205_4372_0, i_13_205_4378_0, i_13_205_4396_0, i_13_205_4518_0,
    o_13_205_0_0  );
  input  i_13_205_31_0, i_13_205_184_0, i_13_205_196_0, i_13_205_259_0,
    i_13_205_325_0, i_13_205_327_0, i_13_205_328_0, i_13_205_382_0,
    i_13_205_526_0, i_13_205_624_0, i_13_205_660_0, i_13_205_661_0,
    i_13_205_742_0, i_13_205_820_0, i_13_205_840_0, i_13_205_850_0,
    i_13_205_852_0, i_13_205_854_0, i_13_205_858_0, i_13_205_861_0,
    i_13_205_1020_0, i_13_205_1074_0, i_13_205_1093_0, i_13_205_1097_0,
    i_13_205_1227_0, i_13_205_1228_0, i_13_205_1229_0, i_13_205_1254_0,
    i_13_205_1255_0, i_13_205_1256_0, i_13_205_1258_0, i_13_205_1314_0,
    i_13_205_1317_0, i_13_205_1383_0, i_13_205_1428_0, i_13_205_1443_0,
    i_13_205_1444_0, i_13_205_1447_0, i_13_205_1483_0, i_13_205_1488_0,
    i_13_205_1645_0, i_13_205_1675_0, i_13_205_1691_0, i_13_205_1753_0,
    i_13_205_1848_0, i_13_205_1849_0, i_13_205_1854_0, i_13_205_1857_0,
    i_13_205_1858_0, i_13_205_1861_0, i_13_205_1953_0, i_13_205_1957_0,
    i_13_205_1993_0, i_13_205_2042_0, i_13_205_2247_0, i_13_205_2248_0,
    i_13_205_2281_0, i_13_205_2394_0, i_13_205_2407_0, i_13_205_2412_0,
    i_13_205_2434_0, i_13_205_2488_0, i_13_205_2614_0, i_13_205_2617_0,
    i_13_205_2701_0, i_13_205_2712_0, i_13_205_2857_0, i_13_205_2878_0,
    i_13_205_2978_0, i_13_205_3064_0, i_13_205_3118_0, i_13_205_3122_0,
    i_13_205_3153_0, i_13_205_3172_0, i_13_205_3307_0, i_13_205_3338_0,
    i_13_205_3355_0, i_13_205_3418_0, i_13_205_3436_0, i_13_205_3456_0,
    i_13_205_3460_0, i_13_205_3478_0, i_13_205_3484_0, i_13_205_3486_0,
    i_13_205_3487_0, i_13_205_3489_0, i_13_205_3537_0, i_13_205_3562_0,
    i_13_205_3689_0, i_13_205_3783_0, i_13_205_3802_0, i_13_205_3868_0,
    i_13_205_3907_0, i_13_205_4063_0, i_13_205_4351_0, i_13_205_4365_0,
    i_13_205_4372_0, i_13_205_4378_0, i_13_205_4396_0, i_13_205_4518_0;
  output o_13_205_0_0;
  assign o_13_205_0_0 = ~((~i_13_205_1753_0 & ~i_13_205_1857_0 & ((~i_13_205_1254_0 & i_13_205_1993_0) | (~i_13_205_1953_0 & ~i_13_205_4372_0))) | (~i_13_205_325_0 & ~i_13_205_1258_0 & ~i_13_205_1488_0 & ~i_13_205_4372_0) | (~i_13_205_1255_0 & ~i_13_205_2248_0));
endmodule



// Benchmark "kernel_13_206" written by ABC on Sun Jul 19 10:48:17 2020

module kernel_13_206 ( 
    i_13_206_13_0, i_13_206_28_0, i_13_206_31_0, i_13_206_43_0,
    i_13_206_64_0, i_13_206_66_0, i_13_206_173_0, i_13_206_310_0,
    i_13_206_399_0, i_13_206_575_0, i_13_206_598_0, i_13_206_604_0,
    i_13_206_607_0, i_13_206_641_0, i_13_206_661_0, i_13_206_670_0,
    i_13_206_672_0, i_13_206_676_0, i_13_206_772_0, i_13_206_814_0,
    i_13_206_829_0, i_13_206_830_0, i_13_206_832_0, i_13_206_833_0,
    i_13_206_851_0, i_13_206_885_0, i_13_206_1066_0, i_13_206_1102_0,
    i_13_206_1113_0, i_13_206_1225_0, i_13_206_1232_0, i_13_206_1259_0,
    i_13_206_1306_0, i_13_206_1307_0, i_13_206_1309_0, i_13_206_1385_0,
    i_13_206_1442_0, i_13_206_1466_0, i_13_206_1491_0, i_13_206_1523_0,
    i_13_206_1549_0, i_13_206_1554_0, i_13_206_1639_0, i_13_206_1697_0,
    i_13_206_1729_0, i_13_206_1795_0, i_13_206_1927_0, i_13_206_1928_0,
    i_13_206_1965_0, i_13_206_2103_0, i_13_206_2135_0, i_13_206_2229_0,
    i_13_206_2297_0, i_13_206_2298_0, i_13_206_2381_0, i_13_206_2535_0,
    i_13_206_2552_0, i_13_206_2677_0, i_13_206_2720_0, i_13_206_2721_0,
    i_13_206_2740_0, i_13_206_2749_0, i_13_206_2802_0, i_13_206_2806_0,
    i_13_206_2879_0, i_13_206_2882_0, i_13_206_2963_0, i_13_206_3000_0,
    i_13_206_3047_0, i_13_206_3255_0, i_13_206_3308_0, i_13_206_3367_0,
    i_13_206_3368_0, i_13_206_3479_0, i_13_206_3537_0, i_13_206_3539_0,
    i_13_206_3544_0, i_13_206_3545_0, i_13_206_3556_0, i_13_206_3637_0,
    i_13_206_3730_0, i_13_206_3754_0, i_13_206_3755_0, i_13_206_3894_0,
    i_13_206_3910_0, i_13_206_3921_0, i_13_206_3935_0, i_13_206_4036_0,
    i_13_206_4063_0, i_13_206_4249_0, i_13_206_4294_0, i_13_206_4313_0,
    i_13_206_4342_0, i_13_206_4349_0, i_13_206_4371_0, i_13_206_4406_0,
    i_13_206_4414_0, i_13_206_4432_0, i_13_206_4592_0, i_13_206_4594_0,
    o_13_206_0_0  );
  input  i_13_206_13_0, i_13_206_28_0, i_13_206_31_0, i_13_206_43_0,
    i_13_206_64_0, i_13_206_66_0, i_13_206_173_0, i_13_206_310_0,
    i_13_206_399_0, i_13_206_575_0, i_13_206_598_0, i_13_206_604_0,
    i_13_206_607_0, i_13_206_641_0, i_13_206_661_0, i_13_206_670_0,
    i_13_206_672_0, i_13_206_676_0, i_13_206_772_0, i_13_206_814_0,
    i_13_206_829_0, i_13_206_830_0, i_13_206_832_0, i_13_206_833_0,
    i_13_206_851_0, i_13_206_885_0, i_13_206_1066_0, i_13_206_1102_0,
    i_13_206_1113_0, i_13_206_1225_0, i_13_206_1232_0, i_13_206_1259_0,
    i_13_206_1306_0, i_13_206_1307_0, i_13_206_1309_0, i_13_206_1385_0,
    i_13_206_1442_0, i_13_206_1466_0, i_13_206_1491_0, i_13_206_1523_0,
    i_13_206_1549_0, i_13_206_1554_0, i_13_206_1639_0, i_13_206_1697_0,
    i_13_206_1729_0, i_13_206_1795_0, i_13_206_1927_0, i_13_206_1928_0,
    i_13_206_1965_0, i_13_206_2103_0, i_13_206_2135_0, i_13_206_2229_0,
    i_13_206_2297_0, i_13_206_2298_0, i_13_206_2381_0, i_13_206_2535_0,
    i_13_206_2552_0, i_13_206_2677_0, i_13_206_2720_0, i_13_206_2721_0,
    i_13_206_2740_0, i_13_206_2749_0, i_13_206_2802_0, i_13_206_2806_0,
    i_13_206_2879_0, i_13_206_2882_0, i_13_206_2963_0, i_13_206_3000_0,
    i_13_206_3047_0, i_13_206_3255_0, i_13_206_3308_0, i_13_206_3367_0,
    i_13_206_3368_0, i_13_206_3479_0, i_13_206_3537_0, i_13_206_3539_0,
    i_13_206_3544_0, i_13_206_3545_0, i_13_206_3556_0, i_13_206_3637_0,
    i_13_206_3730_0, i_13_206_3754_0, i_13_206_3755_0, i_13_206_3894_0,
    i_13_206_3910_0, i_13_206_3921_0, i_13_206_3935_0, i_13_206_4036_0,
    i_13_206_4063_0, i_13_206_4249_0, i_13_206_4294_0, i_13_206_4313_0,
    i_13_206_4342_0, i_13_206_4349_0, i_13_206_4371_0, i_13_206_4406_0,
    i_13_206_4414_0, i_13_206_4432_0, i_13_206_4592_0, i_13_206_4594_0;
  output o_13_206_0_0;
  assign o_13_206_0_0 = ~((~i_13_206_1729_0 & ((~i_13_206_1306_0 & i_13_206_2882_0) | (~i_13_206_885_0 & ~i_13_206_2882_0))) | (~i_13_206_3537_0 & ((~i_13_206_28_0 & ~i_13_206_31_0 & ~i_13_206_2882_0) | (~i_13_206_66_0 & ~i_13_206_2135_0 & ~i_13_206_2298_0 & ~i_13_206_3755_0 & ~i_13_206_4249_0))) | ~i_13_206_1309_0 | (~i_13_206_64_0 & i_13_206_3730_0) | (i_13_206_2677_0 & i_13_206_3537_0 & i_13_206_3910_0) | (~i_13_206_1549_0 & i_13_206_4414_0));
endmodule



// Benchmark "kernel_13_207" written by ABC on Sun Jul 19 10:48:18 2020

module kernel_13_207 ( 
    i_13_207_112_0, i_13_207_143_0, i_13_207_205_0, i_13_207_210_0,
    i_13_207_223_0, i_13_207_251_0, i_13_207_277_0, i_13_207_278_0,
    i_13_207_287_0, i_13_207_322_0, i_13_207_340_0, i_13_207_341_0,
    i_13_207_386_0, i_13_207_447_0, i_13_207_457_0, i_13_207_512_0,
    i_13_207_562_0, i_13_207_563_0, i_13_207_619_0, i_13_207_746_0,
    i_13_207_781_0, i_13_207_1024_0, i_13_207_1085_0, i_13_207_1087_0,
    i_13_207_1088_0, i_13_207_1411_0, i_13_207_1429_0, i_13_207_1430_0,
    i_13_207_1443_0, i_13_207_1475_0, i_13_207_1484_0, i_13_207_1573_0,
    i_13_207_1574_0, i_13_207_1623_0, i_13_207_1624_0, i_13_207_1625_0,
    i_13_207_1634_0, i_13_207_1651_0, i_13_207_1659_0, i_13_207_1736_0,
    i_13_207_1786_0, i_13_207_1816_0, i_13_207_1817_0, i_13_207_1844_0,
    i_13_207_1915_0, i_13_207_1939_0, i_13_207_2005_0, i_13_207_2123_0,
    i_13_207_2137_0, i_13_207_2276_0, i_13_207_2347_0, i_13_207_2348_0,
    i_13_207_2437_0, i_13_207_2455_0, i_13_207_2489_0, i_13_207_2501_0,
    i_13_207_2543_0, i_13_207_2555_0, i_13_207_2712_0, i_13_207_2715_0,
    i_13_207_2716_0, i_13_207_2717_0, i_13_207_2725_0, i_13_207_2726_0,
    i_13_207_2788_0, i_13_207_2858_0, i_13_207_2876_0, i_13_207_3047_0,
    i_13_207_3068_0, i_13_207_3148_0, i_13_207_3149_0, i_13_207_3166_0,
    i_13_207_3221_0, i_13_207_3238_0, i_13_207_3274_0, i_13_207_3328_0,
    i_13_207_3419_0, i_13_207_3454_0, i_13_207_3455_0, i_13_207_3525_0,
    i_13_207_3527_0, i_13_207_3554_0, i_13_207_3685_0, i_13_207_3688_0,
    i_13_207_3689_0, i_13_207_3724_0, i_13_207_3922_0, i_13_207_3932_0,
    i_13_207_3939_0, i_13_207_4036_0, i_13_207_4057_0, i_13_207_4094_0,
    i_13_207_4184_0, i_13_207_4274_0, i_13_207_4328_0, i_13_207_4400_0,
    i_13_207_4408_0, i_13_207_4522_0, i_13_207_4525_0, i_13_207_4544_0,
    o_13_207_0_0  );
  input  i_13_207_112_0, i_13_207_143_0, i_13_207_205_0, i_13_207_210_0,
    i_13_207_223_0, i_13_207_251_0, i_13_207_277_0, i_13_207_278_0,
    i_13_207_287_0, i_13_207_322_0, i_13_207_340_0, i_13_207_341_0,
    i_13_207_386_0, i_13_207_447_0, i_13_207_457_0, i_13_207_512_0,
    i_13_207_562_0, i_13_207_563_0, i_13_207_619_0, i_13_207_746_0,
    i_13_207_781_0, i_13_207_1024_0, i_13_207_1085_0, i_13_207_1087_0,
    i_13_207_1088_0, i_13_207_1411_0, i_13_207_1429_0, i_13_207_1430_0,
    i_13_207_1443_0, i_13_207_1475_0, i_13_207_1484_0, i_13_207_1573_0,
    i_13_207_1574_0, i_13_207_1623_0, i_13_207_1624_0, i_13_207_1625_0,
    i_13_207_1634_0, i_13_207_1651_0, i_13_207_1659_0, i_13_207_1736_0,
    i_13_207_1786_0, i_13_207_1816_0, i_13_207_1817_0, i_13_207_1844_0,
    i_13_207_1915_0, i_13_207_1939_0, i_13_207_2005_0, i_13_207_2123_0,
    i_13_207_2137_0, i_13_207_2276_0, i_13_207_2347_0, i_13_207_2348_0,
    i_13_207_2437_0, i_13_207_2455_0, i_13_207_2489_0, i_13_207_2501_0,
    i_13_207_2543_0, i_13_207_2555_0, i_13_207_2712_0, i_13_207_2715_0,
    i_13_207_2716_0, i_13_207_2717_0, i_13_207_2725_0, i_13_207_2726_0,
    i_13_207_2788_0, i_13_207_2858_0, i_13_207_2876_0, i_13_207_3047_0,
    i_13_207_3068_0, i_13_207_3148_0, i_13_207_3149_0, i_13_207_3166_0,
    i_13_207_3221_0, i_13_207_3238_0, i_13_207_3274_0, i_13_207_3328_0,
    i_13_207_3419_0, i_13_207_3454_0, i_13_207_3455_0, i_13_207_3525_0,
    i_13_207_3527_0, i_13_207_3554_0, i_13_207_3685_0, i_13_207_3688_0,
    i_13_207_3689_0, i_13_207_3724_0, i_13_207_3922_0, i_13_207_3932_0,
    i_13_207_3939_0, i_13_207_4036_0, i_13_207_4057_0, i_13_207_4094_0,
    i_13_207_4184_0, i_13_207_4274_0, i_13_207_4328_0, i_13_207_4400_0,
    i_13_207_4408_0, i_13_207_4522_0, i_13_207_4525_0, i_13_207_4544_0;
  output o_13_207_0_0;
  assign o_13_207_0_0 = ~((~i_13_207_3688_0 & ~i_13_207_4328_0) | (~i_13_207_1429_0 & ~i_13_207_1475_0 & ~i_13_207_1573_0 & ~i_13_207_3689_0) | (~i_13_207_277_0 & ~i_13_207_2717_0 & ~i_13_207_2788_0 & ~i_13_207_3685_0));
endmodule



// Benchmark "kernel_13_208" written by ABC on Sun Jul 19 10:48:19 2020

module kernel_13_208 ( 
    i_13_208_32_0, i_13_208_49_0, i_13_208_104_0, i_13_208_106_0,
    i_13_208_117_0, i_13_208_175_0, i_13_208_185_0, i_13_208_189_0,
    i_13_208_193_0, i_13_208_196_0, i_13_208_216_0, i_13_208_337_0,
    i_13_208_526_0, i_13_208_569_0, i_13_208_575_0, i_13_208_602_0,
    i_13_208_616_0, i_13_208_625_0, i_13_208_626_0, i_13_208_643_0,
    i_13_208_711_0, i_13_208_742_0, i_13_208_746_0, i_13_208_757_0,
    i_13_208_780_0, i_13_208_839_0, i_13_208_845_0, i_13_208_895_0,
    i_13_208_897_0, i_13_208_1018_0, i_13_208_1093_0, i_13_208_1099_0,
    i_13_208_1226_0, i_13_208_1251_0, i_13_208_1310_0, i_13_208_1360_0,
    i_13_208_1381_0, i_13_208_1405_0, i_13_208_1464_0, i_13_208_1478_0,
    i_13_208_1480_0, i_13_208_1481_0, i_13_208_1499_0, i_13_208_1507_0,
    i_13_208_1643_0, i_13_208_1667_0, i_13_208_1678_0, i_13_208_1714_0,
    i_13_208_1720_0, i_13_208_1748_0, i_13_208_1750_0, i_13_208_1754_0,
    i_13_208_1760_0, i_13_208_1805_0, i_13_208_1808_0, i_13_208_1858_0,
    i_13_208_1930_0, i_13_208_2002_0, i_13_208_2119_0, i_13_208_2120_0,
    i_13_208_2138_0, i_13_208_2274_0, i_13_208_2309_0, i_13_208_2395_0,
    i_13_208_2408_0, i_13_208_2447_0, i_13_208_2458_0, i_13_208_2470_0,
    i_13_208_2506_0, i_13_208_2542_0, i_13_208_2621_0, i_13_208_2747_0,
    i_13_208_2751_0, i_13_208_2825_0, i_13_208_2848_0, i_13_208_2876_0,
    i_13_208_2999_0, i_13_208_3173_0, i_13_208_3220_0, i_13_208_3221_0,
    i_13_208_3260_0, i_13_208_3379_0, i_13_208_3380_0, i_13_208_3466_0,
    i_13_208_3721_0, i_13_208_3782_0, i_13_208_3790_0, i_13_208_3791_0,
    i_13_208_3937_0, i_13_208_3942_0, i_13_208_3989_0, i_13_208_4046_0,
    i_13_208_4101_0, i_13_208_4121_0, i_13_208_4238_0, i_13_208_4295_0,
    i_13_208_4315_0, i_13_208_4519_0, i_13_208_4523_0, i_13_208_4525_0,
    o_13_208_0_0  );
  input  i_13_208_32_0, i_13_208_49_0, i_13_208_104_0, i_13_208_106_0,
    i_13_208_117_0, i_13_208_175_0, i_13_208_185_0, i_13_208_189_0,
    i_13_208_193_0, i_13_208_196_0, i_13_208_216_0, i_13_208_337_0,
    i_13_208_526_0, i_13_208_569_0, i_13_208_575_0, i_13_208_602_0,
    i_13_208_616_0, i_13_208_625_0, i_13_208_626_0, i_13_208_643_0,
    i_13_208_711_0, i_13_208_742_0, i_13_208_746_0, i_13_208_757_0,
    i_13_208_780_0, i_13_208_839_0, i_13_208_845_0, i_13_208_895_0,
    i_13_208_897_0, i_13_208_1018_0, i_13_208_1093_0, i_13_208_1099_0,
    i_13_208_1226_0, i_13_208_1251_0, i_13_208_1310_0, i_13_208_1360_0,
    i_13_208_1381_0, i_13_208_1405_0, i_13_208_1464_0, i_13_208_1478_0,
    i_13_208_1480_0, i_13_208_1481_0, i_13_208_1499_0, i_13_208_1507_0,
    i_13_208_1643_0, i_13_208_1667_0, i_13_208_1678_0, i_13_208_1714_0,
    i_13_208_1720_0, i_13_208_1748_0, i_13_208_1750_0, i_13_208_1754_0,
    i_13_208_1760_0, i_13_208_1805_0, i_13_208_1808_0, i_13_208_1858_0,
    i_13_208_1930_0, i_13_208_2002_0, i_13_208_2119_0, i_13_208_2120_0,
    i_13_208_2138_0, i_13_208_2274_0, i_13_208_2309_0, i_13_208_2395_0,
    i_13_208_2408_0, i_13_208_2447_0, i_13_208_2458_0, i_13_208_2470_0,
    i_13_208_2506_0, i_13_208_2542_0, i_13_208_2621_0, i_13_208_2747_0,
    i_13_208_2751_0, i_13_208_2825_0, i_13_208_2848_0, i_13_208_2876_0,
    i_13_208_2999_0, i_13_208_3173_0, i_13_208_3220_0, i_13_208_3221_0,
    i_13_208_3260_0, i_13_208_3379_0, i_13_208_3380_0, i_13_208_3466_0,
    i_13_208_3721_0, i_13_208_3782_0, i_13_208_3790_0, i_13_208_3791_0,
    i_13_208_3937_0, i_13_208_3942_0, i_13_208_3989_0, i_13_208_4046_0,
    i_13_208_4101_0, i_13_208_4121_0, i_13_208_4238_0, i_13_208_4295_0,
    i_13_208_4315_0, i_13_208_4519_0, i_13_208_4523_0, i_13_208_4525_0;
  output o_13_208_0_0;
  assign o_13_208_0_0 = ~((~i_13_208_1481_0 & ((i_13_208_175_0 & ((~i_13_208_189_0 & ~i_13_208_616_0 & ~i_13_208_897_0 & i_13_208_1678_0 & ~i_13_208_2408_0) | (~i_13_208_569_0 & ~i_13_208_1251_0 & ~i_13_208_1480_0 & i_13_208_2002_0 & ~i_13_208_4315_0))) | (~i_13_208_189_0 & ~i_13_208_895_0 & ~i_13_208_897_0 & ~i_13_208_1714_0 & ~i_13_208_1754_0 & ~i_13_208_2274_0 & ~i_13_208_2848_0))) | (i_13_208_526_0 & ((~i_13_208_104_0 & ~i_13_208_1750_0 & ~i_13_208_2458_0) | (~i_13_208_117_0 & ~i_13_208_575_0 & ~i_13_208_897_0 & ~i_13_208_1405_0 & ~i_13_208_2848_0))) | (~i_13_208_3782_0 & ((i_13_208_104_0 & i_13_208_1310_0 & i_13_208_2876_0) | (~i_13_208_895_0 & i_13_208_2002_0 & ~i_13_208_2848_0 & ~i_13_208_3220_0))) | (~i_13_208_189_0 & ~i_13_208_1405_0 & ~i_13_208_1480_0 & ~i_13_208_1750_0 & ~i_13_208_2876_0));
endmodule



// Benchmark "kernel_13_209" written by ABC on Sun Jul 19 10:48:20 2020

module kernel_13_209 ( 
    i_13_209_19_0, i_13_209_69_0, i_13_209_77_0, i_13_209_107_0,
    i_13_209_109_0, i_13_209_112_0, i_13_209_113_0, i_13_209_124_0,
    i_13_209_125_0, i_13_209_130_0, i_13_209_132_0, i_13_209_211_0,
    i_13_209_368_0, i_13_209_463_0, i_13_209_525_0, i_13_209_589_0,
    i_13_209_680_0, i_13_209_949_0, i_13_209_950_0, i_13_209_1061_0,
    i_13_209_1085_0, i_13_209_1087_0, i_13_209_1284_0, i_13_209_1311_0,
    i_13_209_1327_0, i_13_209_1428_0, i_13_209_1489_0, i_13_209_1490_0,
    i_13_209_1519_0, i_13_209_1525_0, i_13_209_1571_0, i_13_209_1574_0,
    i_13_209_1633_0, i_13_209_1634_0, i_13_209_1637_0, i_13_209_1643_0,
    i_13_209_1815_0, i_13_209_1840_0, i_13_209_1841_0, i_13_209_2045_0,
    i_13_209_2128_0, i_13_209_2137_0, i_13_209_2173_0, i_13_209_2266_0,
    i_13_209_2337_0, i_13_209_2380_0, i_13_209_2407_0, i_13_209_2435_0,
    i_13_209_2438_0, i_13_209_2501_0, i_13_209_2512_0, i_13_209_2542_0,
    i_13_209_2543_0, i_13_209_2713_0, i_13_209_2716_0, i_13_209_2717_0,
    i_13_209_2785_0, i_13_209_2923_0, i_13_209_3100_0, i_13_209_3144_0,
    i_13_209_3146_0, i_13_209_3148_0, i_13_209_3149_0, i_13_209_3166_0,
    i_13_209_3167_0, i_13_209_3227_0, i_13_209_3370_0, i_13_209_3371_0,
    i_13_209_3406_0, i_13_209_3418_0, i_13_209_3419_0, i_13_209_3455_0,
    i_13_209_3506_0, i_13_209_3530_0, i_13_209_3553_0, i_13_209_3623_0,
    i_13_209_3686_0, i_13_209_3688_0, i_13_209_3734_0, i_13_209_3770_0,
    i_13_209_3878_0, i_13_209_3892_0, i_13_209_3912_0, i_13_209_3919_0,
    i_13_209_4021_0, i_13_209_4048_0, i_13_209_4120_0, i_13_209_4174_0,
    i_13_209_4256_0, i_13_209_4355_0, i_13_209_4409_0, i_13_209_4417_0,
    i_13_209_4418_0, i_13_209_4513_0, i_13_209_4522_0, i_13_209_4523_0,
    i_13_209_4525_0, i_13_209_4544_0, i_13_209_4555_0, i_13_209_4561_0,
    o_13_209_0_0  );
  input  i_13_209_19_0, i_13_209_69_0, i_13_209_77_0, i_13_209_107_0,
    i_13_209_109_0, i_13_209_112_0, i_13_209_113_0, i_13_209_124_0,
    i_13_209_125_0, i_13_209_130_0, i_13_209_132_0, i_13_209_211_0,
    i_13_209_368_0, i_13_209_463_0, i_13_209_525_0, i_13_209_589_0,
    i_13_209_680_0, i_13_209_949_0, i_13_209_950_0, i_13_209_1061_0,
    i_13_209_1085_0, i_13_209_1087_0, i_13_209_1284_0, i_13_209_1311_0,
    i_13_209_1327_0, i_13_209_1428_0, i_13_209_1489_0, i_13_209_1490_0,
    i_13_209_1519_0, i_13_209_1525_0, i_13_209_1571_0, i_13_209_1574_0,
    i_13_209_1633_0, i_13_209_1634_0, i_13_209_1637_0, i_13_209_1643_0,
    i_13_209_1815_0, i_13_209_1840_0, i_13_209_1841_0, i_13_209_2045_0,
    i_13_209_2128_0, i_13_209_2137_0, i_13_209_2173_0, i_13_209_2266_0,
    i_13_209_2337_0, i_13_209_2380_0, i_13_209_2407_0, i_13_209_2435_0,
    i_13_209_2438_0, i_13_209_2501_0, i_13_209_2512_0, i_13_209_2542_0,
    i_13_209_2543_0, i_13_209_2713_0, i_13_209_2716_0, i_13_209_2717_0,
    i_13_209_2785_0, i_13_209_2923_0, i_13_209_3100_0, i_13_209_3144_0,
    i_13_209_3146_0, i_13_209_3148_0, i_13_209_3149_0, i_13_209_3166_0,
    i_13_209_3167_0, i_13_209_3227_0, i_13_209_3370_0, i_13_209_3371_0,
    i_13_209_3406_0, i_13_209_3418_0, i_13_209_3419_0, i_13_209_3455_0,
    i_13_209_3506_0, i_13_209_3530_0, i_13_209_3553_0, i_13_209_3623_0,
    i_13_209_3686_0, i_13_209_3688_0, i_13_209_3734_0, i_13_209_3770_0,
    i_13_209_3878_0, i_13_209_3892_0, i_13_209_3912_0, i_13_209_3919_0,
    i_13_209_4021_0, i_13_209_4048_0, i_13_209_4120_0, i_13_209_4174_0,
    i_13_209_4256_0, i_13_209_4355_0, i_13_209_4409_0, i_13_209_4417_0,
    i_13_209_4418_0, i_13_209_4513_0, i_13_209_4522_0, i_13_209_4523_0,
    i_13_209_4525_0, i_13_209_4544_0, i_13_209_4555_0, i_13_209_4561_0;
  output o_13_209_0_0;
  assign o_13_209_0_0 = ~((~i_13_209_680_0 & ((~i_13_209_949_0 & ~i_13_209_1085_0) | (~i_13_209_2923_0 & ~i_13_209_3146_0))) | (~i_13_209_4355_0 & (i_13_209_4513_0 | (~i_13_209_3892_0 & ~i_13_209_4048_0))) | (~i_13_209_4418_0 & (i_13_209_2380_0 | (i_13_209_2713_0 & ~i_13_209_4561_0))) | (~i_13_209_69_0 & ~i_13_209_2543_0 & ~i_13_209_3149_0 & ~i_13_209_4561_0) | (i_13_209_2137_0 & ~i_13_209_3878_0));
endmodule



// Benchmark "kernel_13_210" written by ABC on Sun Jul 19 10:48:20 2020

module kernel_13_210 ( 
    i_13_210_35_0, i_13_210_77_0, i_13_210_103_0, i_13_210_107_0,
    i_13_210_121_0, i_13_210_140_0, i_13_210_161_0, i_13_210_358_0,
    i_13_210_368_0, i_13_210_382_0, i_13_210_383_0, i_13_210_386_0,
    i_13_210_458_0, i_13_210_584_0, i_13_210_592_0, i_13_210_737_0,
    i_13_210_745_0, i_13_210_746_0, i_13_210_934_0, i_13_210_950_0,
    i_13_210_953_0, i_13_210_1066_0, i_13_210_1087_0, i_13_210_1132_0,
    i_13_210_1214_0, i_13_210_1220_0, i_13_210_1304_0, i_13_210_1348_0,
    i_13_210_1349_0, i_13_210_1411_0, i_13_210_1438_0, i_13_210_1462_0,
    i_13_210_1474_0, i_13_210_1624_0, i_13_210_1724_0, i_13_210_1726_0,
    i_13_210_1768_0, i_13_210_1772_0, i_13_210_1840_0, i_13_210_1934_0,
    i_13_210_1942_0, i_13_210_2059_0, i_13_210_2060_0, i_13_210_2284_0,
    i_13_210_2285_0, i_13_210_2348_0, i_13_210_2408_0, i_13_210_2515_0,
    i_13_210_2518_0, i_13_210_2555_0, i_13_210_2617_0, i_13_210_2716_0,
    i_13_210_2717_0, i_13_210_2860_0, i_13_210_2861_0, i_13_210_2884_0,
    i_13_210_3130_0, i_13_210_3139_0, i_13_210_3148_0, i_13_210_3325_0,
    i_13_210_3326_0, i_13_210_3388_0, i_13_210_3391_0, i_13_210_3392_0,
    i_13_210_3526_0, i_13_210_3551_0, i_13_210_3562_0, i_13_210_3598_0,
    i_13_210_3599_0, i_13_210_3622_0, i_13_210_3623_0, i_13_210_3634_0,
    i_13_210_3635_0, i_13_210_3686_0, i_13_210_3734_0, i_13_210_3742_0,
    i_13_210_3743_0, i_13_210_3847_0, i_13_210_3923_0, i_13_210_4055_0,
    i_13_210_4085_0, i_13_210_4093_0, i_13_210_4100_0, i_13_210_4103_0,
    i_13_210_4121_0, i_13_210_4165_0, i_13_210_4166_0, i_13_210_4237_0,
    i_13_210_4255_0, i_13_210_4333_0, i_13_210_4345_0, i_13_210_4346_0,
    i_13_210_4388_0, i_13_210_4399_0, i_13_210_4400_0, i_13_210_4418_0,
    i_13_210_4454_0, i_13_210_4514_0, i_13_210_4525_0, i_13_210_4568_0,
    o_13_210_0_0  );
  input  i_13_210_35_0, i_13_210_77_0, i_13_210_103_0, i_13_210_107_0,
    i_13_210_121_0, i_13_210_140_0, i_13_210_161_0, i_13_210_358_0,
    i_13_210_368_0, i_13_210_382_0, i_13_210_383_0, i_13_210_386_0,
    i_13_210_458_0, i_13_210_584_0, i_13_210_592_0, i_13_210_737_0,
    i_13_210_745_0, i_13_210_746_0, i_13_210_934_0, i_13_210_950_0,
    i_13_210_953_0, i_13_210_1066_0, i_13_210_1087_0, i_13_210_1132_0,
    i_13_210_1214_0, i_13_210_1220_0, i_13_210_1304_0, i_13_210_1348_0,
    i_13_210_1349_0, i_13_210_1411_0, i_13_210_1438_0, i_13_210_1462_0,
    i_13_210_1474_0, i_13_210_1624_0, i_13_210_1724_0, i_13_210_1726_0,
    i_13_210_1768_0, i_13_210_1772_0, i_13_210_1840_0, i_13_210_1934_0,
    i_13_210_1942_0, i_13_210_2059_0, i_13_210_2060_0, i_13_210_2284_0,
    i_13_210_2285_0, i_13_210_2348_0, i_13_210_2408_0, i_13_210_2515_0,
    i_13_210_2518_0, i_13_210_2555_0, i_13_210_2617_0, i_13_210_2716_0,
    i_13_210_2717_0, i_13_210_2860_0, i_13_210_2861_0, i_13_210_2884_0,
    i_13_210_3130_0, i_13_210_3139_0, i_13_210_3148_0, i_13_210_3325_0,
    i_13_210_3326_0, i_13_210_3388_0, i_13_210_3391_0, i_13_210_3392_0,
    i_13_210_3526_0, i_13_210_3551_0, i_13_210_3562_0, i_13_210_3598_0,
    i_13_210_3599_0, i_13_210_3622_0, i_13_210_3623_0, i_13_210_3634_0,
    i_13_210_3635_0, i_13_210_3686_0, i_13_210_3734_0, i_13_210_3742_0,
    i_13_210_3743_0, i_13_210_3847_0, i_13_210_3923_0, i_13_210_4055_0,
    i_13_210_4085_0, i_13_210_4093_0, i_13_210_4100_0, i_13_210_4103_0,
    i_13_210_4121_0, i_13_210_4165_0, i_13_210_4166_0, i_13_210_4237_0,
    i_13_210_4255_0, i_13_210_4333_0, i_13_210_4345_0, i_13_210_4346_0,
    i_13_210_4388_0, i_13_210_4399_0, i_13_210_4400_0, i_13_210_4418_0,
    i_13_210_4454_0, i_13_210_4514_0, i_13_210_4525_0, i_13_210_4568_0;
  output o_13_210_0_0;
  assign o_13_210_0_0 = ~((~i_13_210_2861_0 & ~i_13_210_4454_0) | (~i_13_210_1348_0 & i_13_210_2617_0));
endmodule



// Benchmark "kernel_13_211" written by ABC on Sun Jul 19 10:48:21 2020

module kernel_13_211 ( 
    i_13_211_14_0, i_13_211_38_0, i_13_211_112_0, i_13_211_120_0,
    i_13_211_127_0, i_13_211_128_0, i_13_211_180_0, i_13_211_236_0,
    i_13_211_248_0, i_13_211_260_0, i_13_211_319_0, i_13_211_320_0,
    i_13_211_418_0, i_13_211_527_0, i_13_211_531_0, i_13_211_533_0,
    i_13_211_576_0, i_13_211_577_0, i_13_211_596_0, i_13_211_607_0,
    i_13_211_615_0, i_13_211_671_0, i_13_211_695_0, i_13_211_769_0,
    i_13_211_892_0, i_13_211_928_0, i_13_211_945_0, i_13_211_977_0,
    i_13_211_1022_0, i_13_211_1089_0, i_13_211_1117_0, i_13_211_1121_0,
    i_13_211_1301_0, i_13_211_1318_0, i_13_211_1396_0, i_13_211_1397_0,
    i_13_211_1462_0, i_13_211_1480_0, i_13_211_1674_0, i_13_211_1706_0,
    i_13_211_1714_0, i_13_211_1757_0, i_13_211_1760_0, i_13_211_1777_0,
    i_13_211_1805_0, i_13_211_1814_0, i_13_211_1904_0, i_13_211_1918_0,
    i_13_211_2137_0, i_13_211_2138_0, i_13_211_2141_0, i_13_211_2147_0,
    i_13_211_2165_0, i_13_211_2173_0, i_13_211_2181_0, i_13_211_2225_0,
    i_13_211_2300_0, i_13_211_2443_0, i_13_211_2444_0, i_13_211_2458_0,
    i_13_211_2459_0, i_13_211_2630_0, i_13_211_2748_0, i_13_211_2749_0,
    i_13_211_2755_0, i_13_211_2785_0, i_13_211_2786_0, i_13_211_2821_0,
    i_13_211_2822_0, i_13_211_2921_0, i_13_211_2935_0, i_13_211_3105_0,
    i_13_211_3128_0, i_13_211_3206_0, i_13_211_3218_0, i_13_211_3254_0,
    i_13_211_3371_0, i_13_211_3560_0, i_13_211_3593_0, i_13_211_3619_0,
    i_13_211_3620_0, i_13_211_3631_0, i_13_211_3721_0, i_13_211_3791_0,
    i_13_211_3911_0, i_13_211_3928_0, i_13_211_3929_0, i_13_211_3988_0,
    i_13_211_3989_0, i_13_211_4015_0, i_13_211_4082_0, i_13_211_4207_0,
    i_13_211_4312_0, i_13_211_4369_0, i_13_211_4379_0, i_13_211_4391_0,
    i_13_211_4519_0, i_13_211_4522_0, i_13_211_4525_0, i_13_211_4566_0,
    o_13_211_0_0  );
  input  i_13_211_14_0, i_13_211_38_0, i_13_211_112_0, i_13_211_120_0,
    i_13_211_127_0, i_13_211_128_0, i_13_211_180_0, i_13_211_236_0,
    i_13_211_248_0, i_13_211_260_0, i_13_211_319_0, i_13_211_320_0,
    i_13_211_418_0, i_13_211_527_0, i_13_211_531_0, i_13_211_533_0,
    i_13_211_576_0, i_13_211_577_0, i_13_211_596_0, i_13_211_607_0,
    i_13_211_615_0, i_13_211_671_0, i_13_211_695_0, i_13_211_769_0,
    i_13_211_892_0, i_13_211_928_0, i_13_211_945_0, i_13_211_977_0,
    i_13_211_1022_0, i_13_211_1089_0, i_13_211_1117_0, i_13_211_1121_0,
    i_13_211_1301_0, i_13_211_1318_0, i_13_211_1396_0, i_13_211_1397_0,
    i_13_211_1462_0, i_13_211_1480_0, i_13_211_1674_0, i_13_211_1706_0,
    i_13_211_1714_0, i_13_211_1757_0, i_13_211_1760_0, i_13_211_1777_0,
    i_13_211_1805_0, i_13_211_1814_0, i_13_211_1904_0, i_13_211_1918_0,
    i_13_211_2137_0, i_13_211_2138_0, i_13_211_2141_0, i_13_211_2147_0,
    i_13_211_2165_0, i_13_211_2173_0, i_13_211_2181_0, i_13_211_2225_0,
    i_13_211_2300_0, i_13_211_2443_0, i_13_211_2444_0, i_13_211_2458_0,
    i_13_211_2459_0, i_13_211_2630_0, i_13_211_2748_0, i_13_211_2749_0,
    i_13_211_2755_0, i_13_211_2785_0, i_13_211_2786_0, i_13_211_2821_0,
    i_13_211_2822_0, i_13_211_2921_0, i_13_211_2935_0, i_13_211_3105_0,
    i_13_211_3128_0, i_13_211_3206_0, i_13_211_3218_0, i_13_211_3254_0,
    i_13_211_3371_0, i_13_211_3560_0, i_13_211_3593_0, i_13_211_3619_0,
    i_13_211_3620_0, i_13_211_3631_0, i_13_211_3721_0, i_13_211_3791_0,
    i_13_211_3911_0, i_13_211_3928_0, i_13_211_3929_0, i_13_211_3988_0,
    i_13_211_3989_0, i_13_211_4015_0, i_13_211_4082_0, i_13_211_4207_0,
    i_13_211_4312_0, i_13_211_4369_0, i_13_211_4379_0, i_13_211_4391_0,
    i_13_211_4519_0, i_13_211_4522_0, i_13_211_4525_0, i_13_211_4566_0;
  output o_13_211_0_0;
  assign o_13_211_0_0 = ~((~i_13_211_928_0 & (~i_13_211_1397_0 | ~i_13_211_4379_0)) | (~i_13_211_1318_0 & ~i_13_211_2443_0) | (~i_13_211_3911_0 & ~i_13_211_3989_0));
endmodule



// Benchmark "kernel_13_212" written by ABC on Sun Jul 19 10:48:22 2020

module kernel_13_212 ( 
    i_13_212_94_0, i_13_212_95_0, i_13_212_139_0, i_13_212_140_0,
    i_13_212_175_0, i_13_212_177_0, i_13_212_178_0, i_13_212_187_0,
    i_13_212_310_0, i_13_212_319_0, i_13_212_321_0, i_13_212_415_0,
    i_13_212_457_0, i_13_212_510_0, i_13_212_553_0, i_13_212_555_0,
    i_13_212_571_0, i_13_212_574_0, i_13_212_580_0, i_13_212_607_0,
    i_13_212_609_0, i_13_212_610_0, i_13_212_646_0, i_13_212_660_0,
    i_13_212_668_0, i_13_212_714_0, i_13_212_771_0, i_13_212_796_0,
    i_13_212_850_0, i_13_212_853_0, i_13_212_952_0, i_13_212_987_0,
    i_13_212_988_0, i_13_212_1080_0, i_13_212_1123_0, i_13_212_1184_0,
    i_13_212_1203_0, i_13_212_1226_0, i_13_212_1264_0, i_13_212_1282_0,
    i_13_212_1300_0, i_13_212_1302_0, i_13_212_1432_0, i_13_212_1457_0,
    i_13_212_1650_0, i_13_212_1818_0, i_13_212_1828_0, i_13_212_1831_0,
    i_13_212_1861_0, i_13_212_2092_0, i_13_212_2100_0, i_13_212_2140_0,
    i_13_212_2172_0, i_13_212_2175_0, i_13_212_2176_0, i_13_212_2177_0,
    i_13_212_2346_0, i_13_212_2425_0, i_13_212_2427_0, i_13_212_2446_0,
    i_13_212_2470_0, i_13_212_2624_0, i_13_212_2676_0, i_13_212_2695_0,
    i_13_212_2860_0, i_13_212_2887_0, i_13_212_2901_0, i_13_212_3014_0,
    i_13_212_3108_0, i_13_212_3109_0, i_13_212_3112_0, i_13_212_3208_0,
    i_13_212_3217_0, i_13_212_3271_0, i_13_212_3415_0, i_13_212_3418_0,
    i_13_212_3423_0, i_13_212_3426_0, i_13_212_3488_0, i_13_212_3615_0,
    i_13_212_3616_0, i_13_212_3641_0, i_13_212_3685_0, i_13_212_3819_0,
    i_13_212_3820_0, i_13_212_3874_0, i_13_212_3994_0, i_13_212_4054_0,
    i_13_212_4080_0, i_13_212_4084_0, i_13_212_4251_0, i_13_212_4359_0,
    i_13_212_4436_0, i_13_212_4522_0, i_13_212_4523_0, i_13_212_4566_0,
    i_13_212_4567_0, i_13_212_4569_0, i_13_212_4570_0, i_13_212_4593_0,
    o_13_212_0_0  );
  input  i_13_212_94_0, i_13_212_95_0, i_13_212_139_0, i_13_212_140_0,
    i_13_212_175_0, i_13_212_177_0, i_13_212_178_0, i_13_212_187_0,
    i_13_212_310_0, i_13_212_319_0, i_13_212_321_0, i_13_212_415_0,
    i_13_212_457_0, i_13_212_510_0, i_13_212_553_0, i_13_212_555_0,
    i_13_212_571_0, i_13_212_574_0, i_13_212_580_0, i_13_212_607_0,
    i_13_212_609_0, i_13_212_610_0, i_13_212_646_0, i_13_212_660_0,
    i_13_212_668_0, i_13_212_714_0, i_13_212_771_0, i_13_212_796_0,
    i_13_212_850_0, i_13_212_853_0, i_13_212_952_0, i_13_212_987_0,
    i_13_212_988_0, i_13_212_1080_0, i_13_212_1123_0, i_13_212_1184_0,
    i_13_212_1203_0, i_13_212_1226_0, i_13_212_1264_0, i_13_212_1282_0,
    i_13_212_1300_0, i_13_212_1302_0, i_13_212_1432_0, i_13_212_1457_0,
    i_13_212_1650_0, i_13_212_1818_0, i_13_212_1828_0, i_13_212_1831_0,
    i_13_212_1861_0, i_13_212_2092_0, i_13_212_2100_0, i_13_212_2140_0,
    i_13_212_2172_0, i_13_212_2175_0, i_13_212_2176_0, i_13_212_2177_0,
    i_13_212_2346_0, i_13_212_2425_0, i_13_212_2427_0, i_13_212_2446_0,
    i_13_212_2470_0, i_13_212_2624_0, i_13_212_2676_0, i_13_212_2695_0,
    i_13_212_2860_0, i_13_212_2887_0, i_13_212_2901_0, i_13_212_3014_0,
    i_13_212_3108_0, i_13_212_3109_0, i_13_212_3112_0, i_13_212_3208_0,
    i_13_212_3217_0, i_13_212_3271_0, i_13_212_3415_0, i_13_212_3418_0,
    i_13_212_3423_0, i_13_212_3426_0, i_13_212_3488_0, i_13_212_3615_0,
    i_13_212_3616_0, i_13_212_3641_0, i_13_212_3685_0, i_13_212_3819_0,
    i_13_212_3820_0, i_13_212_3874_0, i_13_212_3994_0, i_13_212_4054_0,
    i_13_212_4080_0, i_13_212_4084_0, i_13_212_4251_0, i_13_212_4359_0,
    i_13_212_4436_0, i_13_212_4522_0, i_13_212_4523_0, i_13_212_4566_0,
    i_13_212_4567_0, i_13_212_4569_0, i_13_212_4570_0, i_13_212_4593_0;
  output o_13_212_0_0;
  assign o_13_212_0_0 = ~((~i_13_212_4570_0 & ((~i_13_212_319_0 & ~i_13_212_574_0 & ~i_13_212_987_0 & ~i_13_212_2695_0) | (~i_13_212_177_0 & ~i_13_212_4436_0 & ~i_13_212_4566_0))) | (~i_13_212_94_0 & ~i_13_212_178_0 & ~i_13_212_2427_0 & ~i_13_212_3819_0) | (~i_13_212_571_0 & ~i_13_212_2175_0 & ~i_13_212_3208_0 & ~i_13_212_3820_0) | (~i_13_212_988_0 & ~i_13_212_3108_0 & ~i_13_212_4080_0) | (i_13_212_139_0 & i_13_212_4359_0 & ~i_13_212_4567_0));
endmodule



// Benchmark "kernel_13_213" written by ABC on Sun Jul 19 10:48:23 2020

module kernel_13_213 ( 
    i_13_213_70_0, i_13_213_71_0, i_13_213_78_0, i_13_213_79_0,
    i_13_213_176_0, i_13_213_223_0, i_13_213_313_0, i_13_213_338_0,
    i_13_213_448_0, i_13_213_601_0, i_13_213_608_0, i_13_213_610_0,
    i_13_213_611_0, i_13_213_661_0, i_13_213_662_0, i_13_213_664_0,
    i_13_213_682_0, i_13_213_689_0, i_13_213_760_0, i_13_213_764_0,
    i_13_213_823_0, i_13_213_953_0, i_13_213_985_0, i_13_213_1103_0,
    i_13_213_1105_0, i_13_213_1123_0, i_13_213_1151_0, i_13_213_1232_0,
    i_13_213_1275_0, i_13_213_1276_0, i_13_213_1313_0, i_13_213_1318_0,
    i_13_213_1399_0, i_13_213_1511_0, i_13_213_1542_0, i_13_213_1601_0,
    i_13_213_1627_0, i_13_213_1645_0, i_13_213_1733_0, i_13_213_1736_0,
    i_13_213_1764_0, i_13_213_1768_0, i_13_213_1797_0, i_13_213_1798_0,
    i_13_213_1799_0, i_13_213_1843_0, i_13_213_1888_0, i_13_213_1947_0,
    i_13_213_1948_0, i_13_213_1996_0, i_13_213_2023_0, i_13_213_2024_0,
    i_13_213_2177_0, i_13_213_2426_0, i_13_213_2437_0, i_13_213_2507_0,
    i_13_213_2679_0, i_13_213_2680_0, i_13_213_2681_0, i_13_213_2697_0,
    i_13_213_2788_0, i_13_213_2851_0, i_13_213_2929_0, i_13_213_2930_0,
    i_13_213_3001_0, i_13_213_3130_0, i_13_213_3146_0, i_13_213_3220_0,
    i_13_213_3274_0, i_13_213_3370_0, i_13_213_3418_0, i_13_213_3652_0,
    i_13_213_3656_0, i_13_213_3761_0, i_13_213_3822_0, i_13_213_3823_0,
    i_13_213_3847_0, i_13_213_3895_0, i_13_213_3931_0, i_13_213_3941_0,
    i_13_213_3970_0, i_13_213_3994_0, i_13_213_4019_0, i_13_213_4040_0,
    i_13_213_4063_0, i_13_213_4084_0, i_13_213_4175_0, i_13_213_4189_0,
    i_13_213_4252_0, i_13_213_4297_0, i_13_213_4325_0, i_13_213_4450_0,
    i_13_213_4453_0, i_13_213_4517_0, i_13_213_4522_0, i_13_213_4597_0,
    i_13_213_4598_0, i_13_213_4602_0, i_13_213_4606_0, i_13_213_4607_0,
    o_13_213_0_0  );
  input  i_13_213_70_0, i_13_213_71_0, i_13_213_78_0, i_13_213_79_0,
    i_13_213_176_0, i_13_213_223_0, i_13_213_313_0, i_13_213_338_0,
    i_13_213_448_0, i_13_213_601_0, i_13_213_608_0, i_13_213_610_0,
    i_13_213_611_0, i_13_213_661_0, i_13_213_662_0, i_13_213_664_0,
    i_13_213_682_0, i_13_213_689_0, i_13_213_760_0, i_13_213_764_0,
    i_13_213_823_0, i_13_213_953_0, i_13_213_985_0, i_13_213_1103_0,
    i_13_213_1105_0, i_13_213_1123_0, i_13_213_1151_0, i_13_213_1232_0,
    i_13_213_1275_0, i_13_213_1276_0, i_13_213_1313_0, i_13_213_1318_0,
    i_13_213_1399_0, i_13_213_1511_0, i_13_213_1542_0, i_13_213_1601_0,
    i_13_213_1627_0, i_13_213_1645_0, i_13_213_1733_0, i_13_213_1736_0,
    i_13_213_1764_0, i_13_213_1768_0, i_13_213_1797_0, i_13_213_1798_0,
    i_13_213_1799_0, i_13_213_1843_0, i_13_213_1888_0, i_13_213_1947_0,
    i_13_213_1948_0, i_13_213_1996_0, i_13_213_2023_0, i_13_213_2024_0,
    i_13_213_2177_0, i_13_213_2426_0, i_13_213_2437_0, i_13_213_2507_0,
    i_13_213_2679_0, i_13_213_2680_0, i_13_213_2681_0, i_13_213_2697_0,
    i_13_213_2788_0, i_13_213_2851_0, i_13_213_2929_0, i_13_213_2930_0,
    i_13_213_3001_0, i_13_213_3130_0, i_13_213_3146_0, i_13_213_3220_0,
    i_13_213_3274_0, i_13_213_3370_0, i_13_213_3418_0, i_13_213_3652_0,
    i_13_213_3656_0, i_13_213_3761_0, i_13_213_3822_0, i_13_213_3823_0,
    i_13_213_3847_0, i_13_213_3895_0, i_13_213_3931_0, i_13_213_3941_0,
    i_13_213_3970_0, i_13_213_3994_0, i_13_213_4019_0, i_13_213_4040_0,
    i_13_213_4063_0, i_13_213_4084_0, i_13_213_4175_0, i_13_213_4189_0,
    i_13_213_4252_0, i_13_213_4297_0, i_13_213_4325_0, i_13_213_4450_0,
    i_13_213_4453_0, i_13_213_4517_0, i_13_213_4522_0, i_13_213_4597_0,
    i_13_213_4598_0, i_13_213_4602_0, i_13_213_4606_0, i_13_213_4607_0;
  output o_13_213_0_0;
  assign o_13_213_0_0 = ~(~i_13_213_1511_0 | ~i_13_213_1799_0);
endmodule



// Benchmark "kernel_13_214" written by ABC on Sun Jul 19 10:48:24 2020

module kernel_13_214 ( 
    i_13_214_4_0, i_13_214_70_0, i_13_214_111_0, i_13_214_139_0,
    i_13_214_193_0, i_13_214_229_0, i_13_214_382_0, i_13_214_480_0,
    i_13_214_519_0, i_13_214_607_0, i_13_214_610_0, i_13_214_628_0,
    i_13_214_655_0, i_13_214_661_0, i_13_214_663_0, i_13_214_682_0,
    i_13_214_683_0, i_13_214_886_0, i_13_214_934_0, i_13_214_939_0,
    i_13_214_940_0, i_13_214_988_0, i_13_214_1065_0, i_13_214_1086_0,
    i_13_214_1087_0, i_13_214_1132_0, i_13_214_1147_0, i_13_214_1156_0,
    i_13_214_1321_0, i_13_214_1330_0, i_13_214_1335_0, i_13_214_1519_0,
    i_13_214_1573_0, i_13_214_1660_0, i_13_214_1678_0, i_13_214_1735_0,
    i_13_214_1744_0, i_13_214_1745_0, i_13_214_1798_0, i_13_214_1994_0,
    i_13_214_2020_0, i_13_214_2022_0, i_13_214_2023_0, i_13_214_2024_0,
    i_13_214_2027_0, i_13_214_2198_0, i_13_214_2274_0, i_13_214_2338_0,
    i_13_214_2345_0, i_13_214_2455_0, i_13_214_2471_0, i_13_214_2482_0,
    i_13_214_2501_0, i_13_214_2507_0, i_13_214_2573_0, i_13_214_2715_0,
    i_13_214_2743_0, i_13_214_2765_0, i_13_214_2939_0, i_13_214_3031_0,
    i_13_214_3075_0, i_13_214_3076_0, i_13_214_3094_0, i_13_214_3234_0,
    i_13_214_3244_0, i_13_214_3265_0, i_13_214_3355_0, i_13_214_3452_0,
    i_13_214_3453_0, i_13_214_3454_0, i_13_214_3455_0, i_13_214_3549_0,
    i_13_214_3616_0, i_13_214_3635_0, i_13_214_3643_0, i_13_214_3647_0,
    i_13_214_3649_0, i_13_214_3670_0, i_13_214_3742_0, i_13_214_3822_0,
    i_13_214_3823_0, i_13_214_3939_0, i_13_214_4063_0, i_13_214_4126_0,
    i_13_214_4164_0, i_13_214_4165_0, i_13_214_4166_0, i_13_214_4171_0,
    i_13_214_4175_0, i_13_214_4189_0, i_13_214_4192_0, i_13_214_4201_0,
    i_13_214_4209_0, i_13_214_4324_0, i_13_214_4370_0, i_13_214_4596_0,
    i_13_214_4597_0, i_13_214_4603_0, i_13_214_4606_0, i_13_214_4607_0,
    o_13_214_0_0  );
  input  i_13_214_4_0, i_13_214_70_0, i_13_214_111_0, i_13_214_139_0,
    i_13_214_193_0, i_13_214_229_0, i_13_214_382_0, i_13_214_480_0,
    i_13_214_519_0, i_13_214_607_0, i_13_214_610_0, i_13_214_628_0,
    i_13_214_655_0, i_13_214_661_0, i_13_214_663_0, i_13_214_682_0,
    i_13_214_683_0, i_13_214_886_0, i_13_214_934_0, i_13_214_939_0,
    i_13_214_940_0, i_13_214_988_0, i_13_214_1065_0, i_13_214_1086_0,
    i_13_214_1087_0, i_13_214_1132_0, i_13_214_1147_0, i_13_214_1156_0,
    i_13_214_1321_0, i_13_214_1330_0, i_13_214_1335_0, i_13_214_1519_0,
    i_13_214_1573_0, i_13_214_1660_0, i_13_214_1678_0, i_13_214_1735_0,
    i_13_214_1744_0, i_13_214_1745_0, i_13_214_1798_0, i_13_214_1994_0,
    i_13_214_2020_0, i_13_214_2022_0, i_13_214_2023_0, i_13_214_2024_0,
    i_13_214_2027_0, i_13_214_2198_0, i_13_214_2274_0, i_13_214_2338_0,
    i_13_214_2345_0, i_13_214_2455_0, i_13_214_2471_0, i_13_214_2482_0,
    i_13_214_2501_0, i_13_214_2507_0, i_13_214_2573_0, i_13_214_2715_0,
    i_13_214_2743_0, i_13_214_2765_0, i_13_214_2939_0, i_13_214_3031_0,
    i_13_214_3075_0, i_13_214_3076_0, i_13_214_3094_0, i_13_214_3234_0,
    i_13_214_3244_0, i_13_214_3265_0, i_13_214_3355_0, i_13_214_3452_0,
    i_13_214_3453_0, i_13_214_3454_0, i_13_214_3455_0, i_13_214_3549_0,
    i_13_214_3616_0, i_13_214_3635_0, i_13_214_3643_0, i_13_214_3647_0,
    i_13_214_3649_0, i_13_214_3670_0, i_13_214_3742_0, i_13_214_3822_0,
    i_13_214_3823_0, i_13_214_3939_0, i_13_214_4063_0, i_13_214_4126_0,
    i_13_214_4164_0, i_13_214_4165_0, i_13_214_4166_0, i_13_214_4171_0,
    i_13_214_4175_0, i_13_214_4189_0, i_13_214_4192_0, i_13_214_4201_0,
    i_13_214_4209_0, i_13_214_4324_0, i_13_214_4370_0, i_13_214_4596_0,
    i_13_214_4597_0, i_13_214_4603_0, i_13_214_4606_0, i_13_214_4607_0;
  output o_13_214_0_0;
  assign o_13_214_0_0 = ~((~i_13_214_2023_0 & ((~i_13_214_70_0 & i_13_214_229_0 & ~i_13_214_988_0 & ~i_13_214_2743_0) | (~i_13_214_682_0 & ~i_13_214_939_0 & ~i_13_214_2939_0 & ~i_13_214_3455_0))) | (~i_13_214_1660_0 & i_13_214_1678_0 & ~i_13_214_3616_0) | (~i_13_214_886_0 & ~i_13_214_2274_0 & ~i_13_214_4166_0 & ~i_13_214_4192_0) | (~i_13_214_683_0 & ~i_13_214_2024_0 & ~i_13_214_3742_0 & ~i_13_214_4324_0));
endmodule



// Benchmark "kernel_13_215" written by ABC on Sun Jul 19 10:48:25 2020

module kernel_13_215 ( 
    i_13_215_40_0, i_13_215_136_0, i_13_215_193_0, i_13_215_228_0,
    i_13_215_229_0, i_13_215_265_0, i_13_215_378_0, i_13_215_445_0,
    i_13_215_586_0, i_13_215_639_0, i_13_215_643_0, i_13_215_680_0,
    i_13_215_692_0, i_13_215_711_0, i_13_215_738_0, i_13_215_768_0,
    i_13_215_975_0, i_13_215_1117_0, i_13_215_1124_0, i_13_215_1246_0,
    i_13_215_1269_0, i_13_215_1270_0, i_13_215_1314_0, i_13_215_1341_0,
    i_13_215_1342_0, i_13_215_1387_0, i_13_215_1388_0, i_13_215_1390_0,
    i_13_215_1440_0, i_13_215_1467_0, i_13_215_1468_0, i_13_215_1512_0,
    i_13_215_1513_0, i_13_215_1520_0, i_13_215_1567_0, i_13_215_1587_0,
    i_13_215_1633_0, i_13_215_1638_0, i_13_215_1722_0, i_13_215_1723_0,
    i_13_215_1726_0, i_13_215_1740_0, i_13_215_1767_0, i_13_215_1792_0,
    i_13_215_1793_0, i_13_215_1801_0, i_13_215_1903_0, i_13_215_1926_0,
    i_13_215_1944_0, i_13_215_1945_0, i_13_215_2029_0, i_13_215_2056_0,
    i_13_215_2134_0, i_13_215_2277_0, i_13_215_2278_0, i_13_215_2377_0,
    i_13_215_2411_0, i_13_215_2458_0, i_13_215_2461_0, i_13_215_2646_0,
    i_13_215_2721_0, i_13_215_2745_0, i_13_215_2746_0, i_13_215_2847_0,
    i_13_215_2874_0, i_13_215_3123_0, i_13_215_3135_0, i_13_215_3221_0,
    i_13_215_3340_0, i_13_215_3343_0, i_13_215_3366_0, i_13_215_3367_0,
    i_13_215_3384_0, i_13_215_3385_0, i_13_215_3439_0, i_13_215_3443_0,
    i_13_215_3636_0, i_13_215_3730_0, i_13_215_3784_0, i_13_215_3790_0,
    i_13_215_3793_0, i_13_215_3927_0, i_13_215_3928_0, i_13_215_4017_0,
    i_13_215_4018_0, i_13_215_4041_0, i_13_215_4042_0, i_13_215_4186_0,
    i_13_215_4216_0, i_13_215_4230_0, i_13_215_4231_0, i_13_215_4266_0,
    i_13_215_4293_0, i_13_215_4294_0, i_13_215_4338_0, i_13_215_4375_0,
    i_13_215_4410_0, i_13_215_4411_0, i_13_215_4447_0, i_13_215_4538_0,
    o_13_215_0_0  );
  input  i_13_215_40_0, i_13_215_136_0, i_13_215_193_0, i_13_215_228_0,
    i_13_215_229_0, i_13_215_265_0, i_13_215_378_0, i_13_215_445_0,
    i_13_215_586_0, i_13_215_639_0, i_13_215_643_0, i_13_215_680_0,
    i_13_215_692_0, i_13_215_711_0, i_13_215_738_0, i_13_215_768_0,
    i_13_215_975_0, i_13_215_1117_0, i_13_215_1124_0, i_13_215_1246_0,
    i_13_215_1269_0, i_13_215_1270_0, i_13_215_1314_0, i_13_215_1341_0,
    i_13_215_1342_0, i_13_215_1387_0, i_13_215_1388_0, i_13_215_1390_0,
    i_13_215_1440_0, i_13_215_1467_0, i_13_215_1468_0, i_13_215_1512_0,
    i_13_215_1513_0, i_13_215_1520_0, i_13_215_1567_0, i_13_215_1587_0,
    i_13_215_1633_0, i_13_215_1638_0, i_13_215_1722_0, i_13_215_1723_0,
    i_13_215_1726_0, i_13_215_1740_0, i_13_215_1767_0, i_13_215_1792_0,
    i_13_215_1793_0, i_13_215_1801_0, i_13_215_1903_0, i_13_215_1926_0,
    i_13_215_1944_0, i_13_215_1945_0, i_13_215_2029_0, i_13_215_2056_0,
    i_13_215_2134_0, i_13_215_2277_0, i_13_215_2278_0, i_13_215_2377_0,
    i_13_215_2411_0, i_13_215_2458_0, i_13_215_2461_0, i_13_215_2646_0,
    i_13_215_2721_0, i_13_215_2745_0, i_13_215_2746_0, i_13_215_2847_0,
    i_13_215_2874_0, i_13_215_3123_0, i_13_215_3135_0, i_13_215_3221_0,
    i_13_215_3340_0, i_13_215_3343_0, i_13_215_3366_0, i_13_215_3367_0,
    i_13_215_3384_0, i_13_215_3385_0, i_13_215_3439_0, i_13_215_3443_0,
    i_13_215_3636_0, i_13_215_3730_0, i_13_215_3784_0, i_13_215_3790_0,
    i_13_215_3793_0, i_13_215_3927_0, i_13_215_3928_0, i_13_215_4017_0,
    i_13_215_4018_0, i_13_215_4041_0, i_13_215_4042_0, i_13_215_4186_0,
    i_13_215_4216_0, i_13_215_4230_0, i_13_215_4231_0, i_13_215_4266_0,
    i_13_215_4293_0, i_13_215_4294_0, i_13_215_4338_0, i_13_215_4375_0,
    i_13_215_4410_0, i_13_215_4411_0, i_13_215_4447_0, i_13_215_4538_0;
  output o_13_215_0_0;
  assign o_13_215_0_0 = ~((~i_13_215_4230_0 & (~i_13_215_1270_0 | (~i_13_215_2134_0 & ~i_13_215_3439_0) | (~i_13_215_3384_0 & ~i_13_215_4411_0))) | (~i_13_215_1567_0 & ~i_13_215_3927_0 & ~i_13_215_4410_0));
endmodule



// Benchmark "kernel_13_216" written by ABC on Sun Jul 19 10:48:25 2020

module kernel_13_216 ( 
    i_13_216_75_0, i_13_216_132_0, i_13_216_240_0, i_13_216_250_0,
    i_13_216_258_0, i_13_216_274_0, i_13_216_277_0, i_13_216_321_0,
    i_13_216_339_0, i_13_216_357_0, i_13_216_456_0, i_13_216_561_0,
    i_13_216_588_0, i_13_216_618_0, i_13_216_642_0, i_13_216_699_0,
    i_13_216_844_0, i_13_216_850_0, i_13_216_858_0, i_13_216_943_0,
    i_13_216_1077_0, i_13_216_1084_0, i_13_216_1105_0, i_13_216_1326_0,
    i_13_216_1363_0, i_13_216_1399_0, i_13_216_1431_0, i_13_216_1437_0,
    i_13_216_1470_0, i_13_216_1488_0, i_13_216_1489_0, i_13_216_1507_0,
    i_13_216_1527_0, i_13_216_1528_0, i_13_216_1552_0, i_13_216_1570_0,
    i_13_216_1591_0, i_13_216_1608_0, i_13_216_1693_0, i_13_216_1807_0,
    i_13_216_1908_0, i_13_216_1917_0, i_13_216_1920_0, i_13_216_2002_0,
    i_13_216_2004_0, i_13_216_2016_0, i_13_216_2032_0, i_13_216_2110_0,
    i_13_216_2302_0, i_13_216_2437_0, i_13_216_2502_0, i_13_216_2535_0,
    i_13_216_2544_0, i_13_216_2545_0, i_13_216_2589_0, i_13_216_2751_0,
    i_13_216_2766_0, i_13_216_2769_0, i_13_216_2787_0, i_13_216_2937_0,
    i_13_216_3024_0, i_13_216_3025_0, i_13_216_3064_0, i_13_216_3070_0,
    i_13_216_3129_0, i_13_216_3130_0, i_13_216_3220_0, i_13_216_3315_0,
    i_13_216_3372_0, i_13_216_3417_0, i_13_216_3418_0, i_13_216_3448_0,
    i_13_216_3471_0, i_13_216_3489_0, i_13_216_3552_0, i_13_216_3598_0,
    i_13_216_3613_0, i_13_216_3643_0, i_13_216_3646_0, i_13_216_3687_0,
    i_13_216_3705_0, i_13_216_3711_0, i_13_216_3714_0, i_13_216_3856_0,
    i_13_216_3876_0, i_13_216_3903_0, i_13_216_3904_0, i_13_216_4083_0,
    i_13_216_4084_0, i_13_216_4090_0, i_13_216_4117_0, i_13_216_4160_0,
    i_13_216_4189_0, i_13_216_4360_0, i_13_216_4362_0, i_13_216_4378_0,
    i_13_216_4452_0, i_13_216_4540_0, i_13_216_4543_0, i_13_216_4588_0,
    o_13_216_0_0  );
  input  i_13_216_75_0, i_13_216_132_0, i_13_216_240_0, i_13_216_250_0,
    i_13_216_258_0, i_13_216_274_0, i_13_216_277_0, i_13_216_321_0,
    i_13_216_339_0, i_13_216_357_0, i_13_216_456_0, i_13_216_561_0,
    i_13_216_588_0, i_13_216_618_0, i_13_216_642_0, i_13_216_699_0,
    i_13_216_844_0, i_13_216_850_0, i_13_216_858_0, i_13_216_943_0,
    i_13_216_1077_0, i_13_216_1084_0, i_13_216_1105_0, i_13_216_1326_0,
    i_13_216_1363_0, i_13_216_1399_0, i_13_216_1431_0, i_13_216_1437_0,
    i_13_216_1470_0, i_13_216_1488_0, i_13_216_1489_0, i_13_216_1507_0,
    i_13_216_1527_0, i_13_216_1528_0, i_13_216_1552_0, i_13_216_1570_0,
    i_13_216_1591_0, i_13_216_1608_0, i_13_216_1693_0, i_13_216_1807_0,
    i_13_216_1908_0, i_13_216_1917_0, i_13_216_1920_0, i_13_216_2002_0,
    i_13_216_2004_0, i_13_216_2016_0, i_13_216_2032_0, i_13_216_2110_0,
    i_13_216_2302_0, i_13_216_2437_0, i_13_216_2502_0, i_13_216_2535_0,
    i_13_216_2544_0, i_13_216_2545_0, i_13_216_2589_0, i_13_216_2751_0,
    i_13_216_2766_0, i_13_216_2769_0, i_13_216_2787_0, i_13_216_2937_0,
    i_13_216_3024_0, i_13_216_3025_0, i_13_216_3064_0, i_13_216_3070_0,
    i_13_216_3129_0, i_13_216_3130_0, i_13_216_3220_0, i_13_216_3315_0,
    i_13_216_3372_0, i_13_216_3417_0, i_13_216_3418_0, i_13_216_3448_0,
    i_13_216_3471_0, i_13_216_3489_0, i_13_216_3552_0, i_13_216_3598_0,
    i_13_216_3613_0, i_13_216_3643_0, i_13_216_3646_0, i_13_216_3687_0,
    i_13_216_3705_0, i_13_216_3711_0, i_13_216_3714_0, i_13_216_3856_0,
    i_13_216_3876_0, i_13_216_3903_0, i_13_216_3904_0, i_13_216_4083_0,
    i_13_216_4084_0, i_13_216_4090_0, i_13_216_4117_0, i_13_216_4160_0,
    i_13_216_4189_0, i_13_216_4360_0, i_13_216_4362_0, i_13_216_4378_0,
    i_13_216_4452_0, i_13_216_4540_0, i_13_216_4543_0, i_13_216_4588_0;
  output o_13_216_0_0;
  assign o_13_216_0_0 = ~((~i_13_216_2787_0 & ((~i_13_216_3064_0 & ~i_13_216_3315_0) | (~i_13_216_3903_0 & ~i_13_216_4452_0))) | (~i_13_216_3315_0 & ~i_13_216_4452_0) | (i_13_216_2437_0 & ~i_13_216_4090_0) | (~i_13_216_699_0 & i_13_216_4189_0));
endmodule



// Benchmark "kernel_13_217" written by ABC on Sun Jul 19 10:48:26 2020

module kernel_13_217 ( 
    i_13_217_97_0, i_13_217_116_0, i_13_217_117_0, i_13_217_121_0,
    i_13_217_122_0, i_13_217_124_0, i_13_217_125_0, i_13_217_171_0,
    i_13_217_229_0, i_13_217_279_0, i_13_217_340_0, i_13_217_427_0,
    i_13_217_575_0, i_13_217_589_0, i_13_217_602_0, i_13_217_657_0,
    i_13_217_728_0, i_13_217_741_0, i_13_217_800_0, i_13_217_823_0,
    i_13_217_931_0, i_13_217_949_0, i_13_217_951_0, i_13_217_985_0,
    i_13_217_1024_0, i_13_217_1096_0, i_13_217_1123_0, i_13_217_1224_0,
    i_13_217_1282_0, i_13_217_1283_0, i_13_217_1304_0, i_13_217_1489_0,
    i_13_217_1490_0, i_13_217_1597_0, i_13_217_1600_0, i_13_217_1713_0,
    i_13_217_1787_0, i_13_217_1817_0, i_13_217_1844_0, i_13_217_1848_0,
    i_13_217_2056_0, i_13_217_2090_0, i_13_217_2118_0, i_13_217_2205_0,
    i_13_217_2209_0, i_13_217_2404_0, i_13_217_2429_0, i_13_217_2458_0,
    i_13_217_2461_0, i_13_217_2465_0, i_13_217_2614_0, i_13_217_2615_0,
    i_13_217_2639_0, i_13_217_2698_0, i_13_217_2785_0, i_13_217_2884_0,
    i_13_217_2980_0, i_13_217_3023_0, i_13_217_3047_0, i_13_217_3105_0,
    i_13_217_3146_0, i_13_217_3166_0, i_13_217_3167_0, i_13_217_3176_0,
    i_13_217_3208_0, i_13_217_3214_0, i_13_217_3220_0, i_13_217_3221_0,
    i_13_217_3267_0, i_13_217_3418_0, i_13_217_3420_0, i_13_217_3421_0,
    i_13_217_3425_0, i_13_217_3506_0, i_13_217_3532_0, i_13_217_3535_0,
    i_13_217_3553_0, i_13_217_3688_0, i_13_217_3699_0, i_13_217_3700_0,
    i_13_217_3788_0, i_13_217_3875_0, i_13_217_3877_0, i_13_217_3878_0,
    i_13_217_3928_0, i_13_217_3981_0, i_13_217_3985_0, i_13_217_4008_0,
    i_13_217_4013_0, i_13_217_4018_0, i_13_217_4036_0, i_13_217_4261_0,
    i_13_217_4328_0, i_13_217_4522_0, i_13_217_4523_0, i_13_217_4543_0,
    i_13_217_4544_0, i_13_217_4554_0, i_13_217_4561_0, i_13_217_4597_0,
    o_13_217_0_0  );
  input  i_13_217_97_0, i_13_217_116_0, i_13_217_117_0, i_13_217_121_0,
    i_13_217_122_0, i_13_217_124_0, i_13_217_125_0, i_13_217_171_0,
    i_13_217_229_0, i_13_217_279_0, i_13_217_340_0, i_13_217_427_0,
    i_13_217_575_0, i_13_217_589_0, i_13_217_602_0, i_13_217_657_0,
    i_13_217_728_0, i_13_217_741_0, i_13_217_800_0, i_13_217_823_0,
    i_13_217_931_0, i_13_217_949_0, i_13_217_951_0, i_13_217_985_0,
    i_13_217_1024_0, i_13_217_1096_0, i_13_217_1123_0, i_13_217_1224_0,
    i_13_217_1282_0, i_13_217_1283_0, i_13_217_1304_0, i_13_217_1489_0,
    i_13_217_1490_0, i_13_217_1597_0, i_13_217_1600_0, i_13_217_1713_0,
    i_13_217_1787_0, i_13_217_1817_0, i_13_217_1844_0, i_13_217_1848_0,
    i_13_217_2056_0, i_13_217_2090_0, i_13_217_2118_0, i_13_217_2205_0,
    i_13_217_2209_0, i_13_217_2404_0, i_13_217_2429_0, i_13_217_2458_0,
    i_13_217_2461_0, i_13_217_2465_0, i_13_217_2614_0, i_13_217_2615_0,
    i_13_217_2639_0, i_13_217_2698_0, i_13_217_2785_0, i_13_217_2884_0,
    i_13_217_2980_0, i_13_217_3023_0, i_13_217_3047_0, i_13_217_3105_0,
    i_13_217_3146_0, i_13_217_3166_0, i_13_217_3167_0, i_13_217_3176_0,
    i_13_217_3208_0, i_13_217_3214_0, i_13_217_3220_0, i_13_217_3221_0,
    i_13_217_3267_0, i_13_217_3418_0, i_13_217_3420_0, i_13_217_3421_0,
    i_13_217_3425_0, i_13_217_3506_0, i_13_217_3532_0, i_13_217_3535_0,
    i_13_217_3553_0, i_13_217_3688_0, i_13_217_3699_0, i_13_217_3700_0,
    i_13_217_3788_0, i_13_217_3875_0, i_13_217_3877_0, i_13_217_3878_0,
    i_13_217_3928_0, i_13_217_3981_0, i_13_217_3985_0, i_13_217_4008_0,
    i_13_217_4013_0, i_13_217_4018_0, i_13_217_4036_0, i_13_217_4261_0,
    i_13_217_4328_0, i_13_217_4522_0, i_13_217_4523_0, i_13_217_4543_0,
    i_13_217_4544_0, i_13_217_4554_0, i_13_217_4561_0, i_13_217_4597_0;
  output o_13_217_0_0;
  assign o_13_217_0_0 = ~((~i_13_217_3167_0 & ((i_13_217_589_0 & (i_13_217_1597_0 | i_13_217_1600_0)) | (~i_13_217_340_0 & ~i_13_217_2465_0 & ~i_13_217_3421_0 & ~i_13_217_4008_0))) | (~i_13_217_1597_0 & i_13_217_3421_0) | (~i_13_217_116_0 & ~i_13_217_3875_0 & ~i_13_217_3877_0 & ~i_13_217_4013_0) | (i_13_217_2884_0 & ~i_13_217_4328_0));
endmodule



// Benchmark "kernel_13_218" written by ABC on Sun Jul 19 10:48:27 2020

module kernel_13_218 ( 
    i_13_218_58_0, i_13_218_121_0, i_13_218_183_0, i_13_218_185_0,
    i_13_218_192_0, i_13_218_199_0, i_13_218_225_0, i_13_218_324_0,
    i_13_218_325_0, i_13_218_378_0, i_13_218_380_0, i_13_218_396_0,
    i_13_218_441_0, i_13_218_486_0, i_13_218_526_0, i_13_218_570_0,
    i_13_218_576_0, i_13_218_588_0, i_13_218_589_0, i_13_218_640_0,
    i_13_218_660_0, i_13_218_669_0, i_13_218_697_0, i_13_218_714_0,
    i_13_218_715_0, i_13_218_741_0, i_13_218_756_0, i_13_218_828_0,
    i_13_218_829_0, i_13_218_858_0, i_13_218_859_0, i_13_218_893_0,
    i_13_218_927_0, i_13_218_929_0, i_13_218_948_0, i_13_218_1084_0,
    i_13_218_1102_0, i_13_218_1118_0, i_13_218_1210_0, i_13_218_1219_0,
    i_13_218_1224_0, i_13_218_1225_0, i_13_218_1227_0, i_13_218_1254_0,
    i_13_218_1296_0, i_13_218_1369_0, i_13_218_1408_0, i_13_218_1413_0,
    i_13_218_1434_0, i_13_218_1488_0, i_13_218_1489_0, i_13_218_1507_0,
    i_13_218_1629_0, i_13_218_1719_0, i_13_218_1720_0, i_13_218_1782_0,
    i_13_218_1800_0, i_13_218_1818_0, i_13_218_1819_0, i_13_218_1882_0,
    i_13_218_1990_0, i_13_218_2011_0, i_13_218_2055_0, i_13_218_2128_0,
    i_13_218_2210_0, i_13_218_2224_0, i_13_218_2262_0, i_13_218_2343_0,
    i_13_218_2358_0, i_13_218_2503_0, i_13_218_2532_0, i_13_218_2722_0,
    i_13_218_2757_0, i_13_218_2766_0, i_13_218_2980_0, i_13_218_2981_0,
    i_13_218_3024_0, i_13_218_3114_0, i_13_218_3171_0, i_13_218_3259_0,
    i_13_218_3285_0, i_13_218_3286_0, i_13_218_3287_0, i_13_218_3420_0,
    i_13_218_3421_0, i_13_218_3423_0, i_13_218_3424_0, i_13_218_3451_0,
    i_13_218_3577_0, i_13_218_3649_0, i_13_218_3873_0, i_13_218_4008_0,
    i_13_218_4009_0, i_13_218_4050_0, i_13_218_4077_0, i_13_218_4087_0,
    i_13_218_4167_0, i_13_218_4232_0, i_13_218_4557_0, i_13_218_4582_0,
    o_13_218_0_0  );
  input  i_13_218_58_0, i_13_218_121_0, i_13_218_183_0, i_13_218_185_0,
    i_13_218_192_0, i_13_218_199_0, i_13_218_225_0, i_13_218_324_0,
    i_13_218_325_0, i_13_218_378_0, i_13_218_380_0, i_13_218_396_0,
    i_13_218_441_0, i_13_218_486_0, i_13_218_526_0, i_13_218_570_0,
    i_13_218_576_0, i_13_218_588_0, i_13_218_589_0, i_13_218_640_0,
    i_13_218_660_0, i_13_218_669_0, i_13_218_697_0, i_13_218_714_0,
    i_13_218_715_0, i_13_218_741_0, i_13_218_756_0, i_13_218_828_0,
    i_13_218_829_0, i_13_218_858_0, i_13_218_859_0, i_13_218_893_0,
    i_13_218_927_0, i_13_218_929_0, i_13_218_948_0, i_13_218_1084_0,
    i_13_218_1102_0, i_13_218_1118_0, i_13_218_1210_0, i_13_218_1219_0,
    i_13_218_1224_0, i_13_218_1225_0, i_13_218_1227_0, i_13_218_1254_0,
    i_13_218_1296_0, i_13_218_1369_0, i_13_218_1408_0, i_13_218_1413_0,
    i_13_218_1434_0, i_13_218_1488_0, i_13_218_1489_0, i_13_218_1507_0,
    i_13_218_1629_0, i_13_218_1719_0, i_13_218_1720_0, i_13_218_1782_0,
    i_13_218_1800_0, i_13_218_1818_0, i_13_218_1819_0, i_13_218_1882_0,
    i_13_218_1990_0, i_13_218_2011_0, i_13_218_2055_0, i_13_218_2128_0,
    i_13_218_2210_0, i_13_218_2224_0, i_13_218_2262_0, i_13_218_2343_0,
    i_13_218_2358_0, i_13_218_2503_0, i_13_218_2532_0, i_13_218_2722_0,
    i_13_218_2757_0, i_13_218_2766_0, i_13_218_2980_0, i_13_218_2981_0,
    i_13_218_3024_0, i_13_218_3114_0, i_13_218_3171_0, i_13_218_3259_0,
    i_13_218_3285_0, i_13_218_3286_0, i_13_218_3287_0, i_13_218_3420_0,
    i_13_218_3421_0, i_13_218_3423_0, i_13_218_3424_0, i_13_218_3451_0,
    i_13_218_3577_0, i_13_218_3649_0, i_13_218_3873_0, i_13_218_4008_0,
    i_13_218_4009_0, i_13_218_4050_0, i_13_218_4077_0, i_13_218_4087_0,
    i_13_218_4167_0, i_13_218_4232_0, i_13_218_4557_0, i_13_218_4582_0;
  output o_13_218_0_0;
  assign o_13_218_0_0 = ~(~i_13_218_927_0 | ~i_13_218_3424_0);
endmodule



// Benchmark "kernel_13_219" written by ABC on Sun Jul 19 10:48:28 2020

module kernel_13_219 ( 
    i_13_219_49_0, i_13_219_101_0, i_13_219_109_0, i_13_219_112_0,
    i_13_219_141_0, i_13_219_175_0, i_13_219_210_0, i_13_219_220_0,
    i_13_219_279_0, i_13_219_281_0, i_13_219_284_0, i_13_219_287_0,
    i_13_219_317_0, i_13_219_337_0, i_13_219_382_0, i_13_219_425_0,
    i_13_219_445_0, i_13_219_534_0, i_13_219_550_0, i_13_219_551_0,
    i_13_219_554_0, i_13_219_613_0, i_13_219_652_0, i_13_219_653_0,
    i_13_219_654_0, i_13_219_655_0, i_13_219_658_0, i_13_219_668_0,
    i_13_219_676_0, i_13_219_677_0, i_13_219_679_0, i_13_219_688_0,
    i_13_219_844_0, i_13_219_852_0, i_13_219_853_0, i_13_219_1018_0,
    i_13_219_1144_0, i_13_219_1216_0, i_13_219_1300_0, i_13_219_1400_0,
    i_13_219_1423_0, i_13_219_1424_0, i_13_219_1516_0, i_13_219_1624_0,
    i_13_219_1643_0, i_13_219_1658_0, i_13_219_1668_0, i_13_219_1671_0,
    i_13_219_1748_0, i_13_219_1774_0, i_13_219_1801_0, i_13_219_1804_0,
    i_13_219_1840_0, i_13_219_1842_0, i_13_219_1921_0, i_13_219_1945_0,
    i_13_219_2000_0, i_13_219_2101_0, i_13_219_2146_0, i_13_219_2170_0,
    i_13_219_2331_0, i_13_219_2380_0, i_13_219_2433_0, i_13_219_2472_0,
    i_13_219_2473_0, i_13_219_2611_0, i_13_219_2674_0, i_13_219_2693_0,
    i_13_219_2697_0, i_13_219_2722_0, i_13_219_2767_0, i_13_219_2847_0,
    i_13_219_2850_0, i_13_219_2938_0, i_13_219_2956_0, i_13_219_2999_0,
    i_13_219_3054_0, i_13_219_3108_0, i_13_219_3368_0, i_13_219_3502_0,
    i_13_219_3523_0, i_13_219_3524_0, i_13_219_3637_0, i_13_219_3640_0,
    i_13_219_3767_0, i_13_219_3863_0, i_13_219_3889_0, i_13_219_3890_0,
    i_13_219_4034_0, i_13_219_4045_0, i_13_219_4117_0, i_13_219_4121_0,
    i_13_219_4270_0, i_13_219_4314_0, i_13_219_4377_0, i_13_219_4413_0,
    i_13_219_4556_0, i_13_219_4558_0, i_13_219_4600_0, i_13_219_4601_0,
    o_13_219_0_0  );
  input  i_13_219_49_0, i_13_219_101_0, i_13_219_109_0, i_13_219_112_0,
    i_13_219_141_0, i_13_219_175_0, i_13_219_210_0, i_13_219_220_0,
    i_13_219_279_0, i_13_219_281_0, i_13_219_284_0, i_13_219_287_0,
    i_13_219_317_0, i_13_219_337_0, i_13_219_382_0, i_13_219_425_0,
    i_13_219_445_0, i_13_219_534_0, i_13_219_550_0, i_13_219_551_0,
    i_13_219_554_0, i_13_219_613_0, i_13_219_652_0, i_13_219_653_0,
    i_13_219_654_0, i_13_219_655_0, i_13_219_658_0, i_13_219_668_0,
    i_13_219_676_0, i_13_219_677_0, i_13_219_679_0, i_13_219_688_0,
    i_13_219_844_0, i_13_219_852_0, i_13_219_853_0, i_13_219_1018_0,
    i_13_219_1144_0, i_13_219_1216_0, i_13_219_1300_0, i_13_219_1400_0,
    i_13_219_1423_0, i_13_219_1424_0, i_13_219_1516_0, i_13_219_1624_0,
    i_13_219_1643_0, i_13_219_1658_0, i_13_219_1668_0, i_13_219_1671_0,
    i_13_219_1748_0, i_13_219_1774_0, i_13_219_1801_0, i_13_219_1804_0,
    i_13_219_1840_0, i_13_219_1842_0, i_13_219_1921_0, i_13_219_1945_0,
    i_13_219_2000_0, i_13_219_2101_0, i_13_219_2146_0, i_13_219_2170_0,
    i_13_219_2331_0, i_13_219_2380_0, i_13_219_2433_0, i_13_219_2472_0,
    i_13_219_2473_0, i_13_219_2611_0, i_13_219_2674_0, i_13_219_2693_0,
    i_13_219_2697_0, i_13_219_2722_0, i_13_219_2767_0, i_13_219_2847_0,
    i_13_219_2850_0, i_13_219_2938_0, i_13_219_2956_0, i_13_219_2999_0,
    i_13_219_3054_0, i_13_219_3108_0, i_13_219_3368_0, i_13_219_3502_0,
    i_13_219_3523_0, i_13_219_3524_0, i_13_219_3637_0, i_13_219_3640_0,
    i_13_219_3767_0, i_13_219_3863_0, i_13_219_3889_0, i_13_219_3890_0,
    i_13_219_4034_0, i_13_219_4045_0, i_13_219_4117_0, i_13_219_4121_0,
    i_13_219_4270_0, i_13_219_4314_0, i_13_219_4377_0, i_13_219_4413_0,
    i_13_219_4556_0, i_13_219_4558_0, i_13_219_4600_0, i_13_219_4601_0;
  output o_13_219_0_0;
  assign o_13_219_0_0 = ~((~i_13_219_3890_0 & ((~i_13_219_668_0 & ~i_13_219_676_0) | (~i_13_219_281_0 & ~i_13_219_1018_0 & ~i_13_219_2433_0))) | (~i_13_219_317_0 & ~i_13_219_1144_0 & i_13_219_2938_0));
endmodule



// Benchmark "kernel_13_220" written by ABC on Sun Jul 19 10:48:29 2020

module kernel_13_220 ( 
    i_13_220_48_0, i_13_220_134_0, i_13_220_184_0, i_13_220_234_0,
    i_13_220_238_0, i_13_220_322_0, i_13_220_351_0, i_13_220_354_0,
    i_13_220_357_0, i_13_220_358_0, i_13_220_374_0, i_13_220_455_0,
    i_13_220_480_0, i_13_220_525_0, i_13_220_529_0, i_13_220_530_0,
    i_13_220_558_0, i_13_220_1024_0, i_13_220_1053_0, i_13_220_1079_0,
    i_13_220_1080_0, i_13_220_1085_0, i_13_220_1210_0, i_13_220_1371_0,
    i_13_220_1396_0, i_13_220_1399_0, i_13_220_1422_0, i_13_220_1426_0,
    i_13_220_1430_0, i_13_220_1458_0, i_13_220_1497_0, i_13_220_1498_0,
    i_13_220_1501_0, i_13_220_1502_0, i_13_220_1504_0, i_13_220_1555_0,
    i_13_220_1556_0, i_13_220_1620_0, i_13_220_1629_0, i_13_220_1637_0,
    i_13_220_1917_0, i_13_220_1921_0, i_13_220_1950_0, i_13_220_2006_0,
    i_13_220_2031_0, i_13_220_2033_0, i_13_220_2109_0, i_13_220_2203_0,
    i_13_220_2300_0, i_13_220_2368_0, i_13_220_2510_0, i_13_220_2511_0,
    i_13_220_2542_0, i_13_220_2691_0, i_13_220_2723_0, i_13_220_2767_0,
    i_13_220_2768_0, i_13_220_2788_0, i_13_220_2924_0, i_13_220_2934_0,
    i_13_220_2939_0, i_13_220_2955_0, i_13_220_2959_0, i_13_220_3014_0,
    i_13_220_3065_0, i_13_220_3069_0, i_13_220_3110_0, i_13_220_3123_0,
    i_13_220_3221_0, i_13_220_3235_0, i_13_220_3316_0, i_13_220_3373_0,
    i_13_220_3374_0, i_13_220_3403_0, i_13_220_3405_0, i_13_220_3432_0,
    i_13_220_3439_0, i_13_220_3464_0, i_13_220_3491_0, i_13_220_3576_0,
    i_13_220_3581_0, i_13_220_3594_0, i_13_220_3598_0, i_13_220_3599_0,
    i_13_220_3618_0, i_13_220_3646_0, i_13_220_3733_0, i_13_220_3781_0,
    i_13_220_3860_0, i_13_220_3904_0, i_13_220_3987_0, i_13_220_4067_0,
    i_13_220_4108_0, i_13_220_4212_0, i_13_220_4249_0, i_13_220_4271_0,
    i_13_220_4329_0, i_13_220_4453_0, i_13_220_4454_0, i_13_220_4561_0,
    o_13_220_0_0  );
  input  i_13_220_48_0, i_13_220_134_0, i_13_220_184_0, i_13_220_234_0,
    i_13_220_238_0, i_13_220_322_0, i_13_220_351_0, i_13_220_354_0,
    i_13_220_357_0, i_13_220_358_0, i_13_220_374_0, i_13_220_455_0,
    i_13_220_480_0, i_13_220_525_0, i_13_220_529_0, i_13_220_530_0,
    i_13_220_558_0, i_13_220_1024_0, i_13_220_1053_0, i_13_220_1079_0,
    i_13_220_1080_0, i_13_220_1085_0, i_13_220_1210_0, i_13_220_1371_0,
    i_13_220_1396_0, i_13_220_1399_0, i_13_220_1422_0, i_13_220_1426_0,
    i_13_220_1430_0, i_13_220_1458_0, i_13_220_1497_0, i_13_220_1498_0,
    i_13_220_1501_0, i_13_220_1502_0, i_13_220_1504_0, i_13_220_1555_0,
    i_13_220_1556_0, i_13_220_1620_0, i_13_220_1629_0, i_13_220_1637_0,
    i_13_220_1917_0, i_13_220_1921_0, i_13_220_1950_0, i_13_220_2006_0,
    i_13_220_2031_0, i_13_220_2033_0, i_13_220_2109_0, i_13_220_2203_0,
    i_13_220_2300_0, i_13_220_2368_0, i_13_220_2510_0, i_13_220_2511_0,
    i_13_220_2542_0, i_13_220_2691_0, i_13_220_2723_0, i_13_220_2767_0,
    i_13_220_2768_0, i_13_220_2788_0, i_13_220_2924_0, i_13_220_2934_0,
    i_13_220_2939_0, i_13_220_2955_0, i_13_220_2959_0, i_13_220_3014_0,
    i_13_220_3065_0, i_13_220_3069_0, i_13_220_3110_0, i_13_220_3123_0,
    i_13_220_3221_0, i_13_220_3235_0, i_13_220_3316_0, i_13_220_3373_0,
    i_13_220_3374_0, i_13_220_3403_0, i_13_220_3405_0, i_13_220_3432_0,
    i_13_220_3439_0, i_13_220_3464_0, i_13_220_3491_0, i_13_220_3576_0,
    i_13_220_3581_0, i_13_220_3594_0, i_13_220_3598_0, i_13_220_3599_0,
    i_13_220_3618_0, i_13_220_3646_0, i_13_220_3733_0, i_13_220_3781_0,
    i_13_220_3860_0, i_13_220_3904_0, i_13_220_3987_0, i_13_220_4067_0,
    i_13_220_4108_0, i_13_220_4212_0, i_13_220_4249_0, i_13_220_4271_0,
    i_13_220_4329_0, i_13_220_4453_0, i_13_220_4454_0, i_13_220_4561_0;
  output o_13_220_0_0;
  assign o_13_220_0_0 = ~((~i_13_220_3904_0 & (~i_13_220_2300_0 | ~i_13_220_3581_0)) | (~i_13_220_1430_0 & ~i_13_220_2924_0) | (~i_13_220_3014_0 & ~i_13_220_3464_0 & ~i_13_220_3599_0));
endmodule



// Benchmark "kernel_13_221" written by ABC on Sun Jul 19 10:48:30 2020

module kernel_13_221 ( 
    i_13_221_37_0, i_13_221_73_0, i_13_221_74_0, i_13_221_109_0,
    i_13_221_110_0, i_13_221_113_0, i_13_221_116_0, i_13_221_122_0,
    i_13_221_157_0, i_13_221_262_0, i_13_221_365_0, i_13_221_366_0,
    i_13_221_551_0, i_13_221_559_0, i_13_221_562_0, i_13_221_604_0,
    i_13_221_605_0, i_13_221_613_0, i_13_221_639_0, i_13_221_676_0,
    i_13_221_677_0, i_13_221_814_0, i_13_221_821_0, i_13_221_947_0,
    i_13_221_992_0, i_13_221_1081_0, i_13_221_1084_0, i_13_221_1085_0,
    i_13_221_1120_0, i_13_221_1144_0, i_13_221_1217_0, i_13_221_1220_0,
    i_13_221_1283_0, i_13_221_1408_0, i_13_221_1424_0, i_13_221_1521_0,
    i_13_221_1541_0, i_13_221_1567_0, i_13_221_1621_0, i_13_221_1631_0,
    i_13_221_1720_0, i_13_221_1721_0, i_13_221_1775_0, i_13_221_1837_0,
    i_13_221_1838_0, i_13_221_1840_0, i_13_221_1841_0, i_13_221_1898_0,
    i_13_221_1945_0, i_13_221_1957_0, i_13_221_2021_0, i_13_221_2054_0,
    i_13_221_2134_0, i_13_221_2170_0, i_13_221_2171_0, i_13_221_2341_0,
    i_13_221_2345_0, i_13_221_2404_0, i_13_221_2432_0, i_13_221_2498_0,
    i_13_221_2611_0, i_13_221_2702_0, i_13_221_2746_0, i_13_221_2767_0,
    i_13_221_2818_0, i_13_221_2845_0, i_13_221_2846_0, i_13_221_2956_0,
    i_13_221_2958_0, i_13_221_3044_0, i_13_221_3098_0, i_13_221_3099_0,
    i_13_221_3100_0, i_13_221_3110_0, i_13_221_3125_0, i_13_221_3142_0,
    i_13_221_3146_0, i_13_221_3148_0, i_13_221_3152_0, i_13_221_3376_0,
    i_13_221_3377_0, i_13_221_3404_0, i_13_221_3452_0, i_13_221_3503_0,
    i_13_221_3524_0, i_13_221_3552_0, i_13_221_3686_0, i_13_221_3731_0,
    i_13_221_3736_0, i_13_221_3737_0, i_13_221_3802_0, i_13_221_3836_0,
    i_13_221_3910_0, i_13_221_3917_0, i_13_221_4051_0, i_13_221_4118_0,
    i_13_221_4160_0, i_13_221_4339_0, i_13_221_4541_0, i_13_221_4542_0,
    o_13_221_0_0  );
  input  i_13_221_37_0, i_13_221_73_0, i_13_221_74_0, i_13_221_109_0,
    i_13_221_110_0, i_13_221_113_0, i_13_221_116_0, i_13_221_122_0,
    i_13_221_157_0, i_13_221_262_0, i_13_221_365_0, i_13_221_366_0,
    i_13_221_551_0, i_13_221_559_0, i_13_221_562_0, i_13_221_604_0,
    i_13_221_605_0, i_13_221_613_0, i_13_221_639_0, i_13_221_676_0,
    i_13_221_677_0, i_13_221_814_0, i_13_221_821_0, i_13_221_947_0,
    i_13_221_992_0, i_13_221_1081_0, i_13_221_1084_0, i_13_221_1085_0,
    i_13_221_1120_0, i_13_221_1144_0, i_13_221_1217_0, i_13_221_1220_0,
    i_13_221_1283_0, i_13_221_1408_0, i_13_221_1424_0, i_13_221_1521_0,
    i_13_221_1541_0, i_13_221_1567_0, i_13_221_1621_0, i_13_221_1631_0,
    i_13_221_1720_0, i_13_221_1721_0, i_13_221_1775_0, i_13_221_1837_0,
    i_13_221_1838_0, i_13_221_1840_0, i_13_221_1841_0, i_13_221_1898_0,
    i_13_221_1945_0, i_13_221_1957_0, i_13_221_2021_0, i_13_221_2054_0,
    i_13_221_2134_0, i_13_221_2170_0, i_13_221_2171_0, i_13_221_2341_0,
    i_13_221_2345_0, i_13_221_2404_0, i_13_221_2432_0, i_13_221_2498_0,
    i_13_221_2611_0, i_13_221_2702_0, i_13_221_2746_0, i_13_221_2767_0,
    i_13_221_2818_0, i_13_221_2845_0, i_13_221_2846_0, i_13_221_2956_0,
    i_13_221_2958_0, i_13_221_3044_0, i_13_221_3098_0, i_13_221_3099_0,
    i_13_221_3100_0, i_13_221_3110_0, i_13_221_3125_0, i_13_221_3142_0,
    i_13_221_3146_0, i_13_221_3148_0, i_13_221_3152_0, i_13_221_3376_0,
    i_13_221_3377_0, i_13_221_3404_0, i_13_221_3452_0, i_13_221_3503_0,
    i_13_221_3524_0, i_13_221_3552_0, i_13_221_3686_0, i_13_221_3731_0,
    i_13_221_3736_0, i_13_221_3737_0, i_13_221_3802_0, i_13_221_3836_0,
    i_13_221_3910_0, i_13_221_3917_0, i_13_221_4051_0, i_13_221_4118_0,
    i_13_221_4160_0, i_13_221_4339_0, i_13_221_4541_0, i_13_221_4542_0;
  output o_13_221_0_0;
  assign o_13_221_0_0 = ~((~i_13_221_2171_0 & (i_13_221_613_0 | i_13_221_3917_0)) | (~i_13_221_1217_0 & ~i_13_221_2845_0 & ~i_13_221_3098_0) | (~i_13_221_2170_0 & ~i_13_221_3142_0) | (i_13_221_2767_0 & i_13_221_3736_0) | (~i_13_221_73_0 & ~i_13_221_110_0 & ~i_13_221_1775_0 & ~i_13_221_3737_0));
endmodule



// Benchmark "kernel_13_222" written by ABC on Sun Jul 19 10:48:31 2020

module kernel_13_222 ( 
    i_13_222_40_0, i_13_222_100_0, i_13_222_106_0, i_13_222_115_0,
    i_13_222_116_0, i_13_222_125_0, i_13_222_184_0, i_13_222_197_0,
    i_13_222_269_0, i_13_222_278_0, i_13_222_602_0, i_13_222_610_0,
    i_13_222_611_0, i_13_222_664_0, i_13_222_665_0, i_13_222_700_0,
    i_13_222_701_0, i_13_222_763_0, i_13_222_772_0, i_13_222_832_0,
    i_13_222_862_0, i_13_222_863_0, i_13_222_872_0, i_13_222_932_0,
    i_13_222_943_0, i_13_222_944_0, i_13_222_950_0, i_13_222_953_0,
    i_13_222_1075_0, i_13_222_1085_0, i_13_222_1262_0, i_13_222_1277_0,
    i_13_222_1286_0, i_13_222_1298_0, i_13_222_1411_0, i_13_222_1438_0,
    i_13_222_1481_0, i_13_222_1501_0, i_13_222_1539_0, i_13_222_1625_0,
    i_13_222_1636_0, i_13_222_1637_0, i_13_222_1660_0, i_13_222_1661_0,
    i_13_222_1682_0, i_13_222_1734_0, i_13_222_1843_0, i_13_222_1844_0,
    i_13_222_1931_0, i_13_222_1961_0, i_13_222_1996_0, i_13_222_2003_0,
    i_13_222_2006_0, i_13_222_2140_0, i_13_222_2303_0, i_13_222_2320_0,
    i_13_222_2438_0, i_13_222_2456_0, i_13_222_2536_0, i_13_222_2544_0,
    i_13_222_2545_0, i_13_222_2546_0, i_13_222_2616_0, i_13_222_2617_0,
    i_13_222_2618_0, i_13_222_2663_0, i_13_222_2798_0, i_13_222_2887_0,
    i_13_222_2888_0, i_13_222_2959_0, i_13_222_3004_0, i_13_222_3050_0,
    i_13_222_3113_0, i_13_222_3262_0, i_13_222_3316_0, i_13_222_3464_0,
    i_13_222_3490_0, i_13_222_3535_0, i_13_222_3571_0, i_13_222_3604_0,
    i_13_222_3731_0, i_13_222_3733_0, i_13_222_3769_0, i_13_222_3770_0,
    i_13_222_3878_0, i_13_222_3904_0, i_13_222_3905_0, i_13_222_3910_0,
    i_13_222_4090_0, i_13_222_4091_0, i_13_222_4166_0, i_13_222_4211_0,
    i_13_222_4343_0, i_13_222_4358_0, i_13_222_4372_0, i_13_222_4373_0,
    i_13_222_4391_0, i_13_222_4433_0, i_13_222_4517_0, i_13_222_4586_0,
    o_13_222_0_0  );
  input  i_13_222_40_0, i_13_222_100_0, i_13_222_106_0, i_13_222_115_0,
    i_13_222_116_0, i_13_222_125_0, i_13_222_184_0, i_13_222_197_0,
    i_13_222_269_0, i_13_222_278_0, i_13_222_602_0, i_13_222_610_0,
    i_13_222_611_0, i_13_222_664_0, i_13_222_665_0, i_13_222_700_0,
    i_13_222_701_0, i_13_222_763_0, i_13_222_772_0, i_13_222_832_0,
    i_13_222_862_0, i_13_222_863_0, i_13_222_872_0, i_13_222_932_0,
    i_13_222_943_0, i_13_222_944_0, i_13_222_950_0, i_13_222_953_0,
    i_13_222_1075_0, i_13_222_1085_0, i_13_222_1262_0, i_13_222_1277_0,
    i_13_222_1286_0, i_13_222_1298_0, i_13_222_1411_0, i_13_222_1438_0,
    i_13_222_1481_0, i_13_222_1501_0, i_13_222_1539_0, i_13_222_1625_0,
    i_13_222_1636_0, i_13_222_1637_0, i_13_222_1660_0, i_13_222_1661_0,
    i_13_222_1682_0, i_13_222_1734_0, i_13_222_1843_0, i_13_222_1844_0,
    i_13_222_1931_0, i_13_222_1961_0, i_13_222_1996_0, i_13_222_2003_0,
    i_13_222_2006_0, i_13_222_2140_0, i_13_222_2303_0, i_13_222_2320_0,
    i_13_222_2438_0, i_13_222_2456_0, i_13_222_2536_0, i_13_222_2544_0,
    i_13_222_2545_0, i_13_222_2546_0, i_13_222_2616_0, i_13_222_2617_0,
    i_13_222_2618_0, i_13_222_2663_0, i_13_222_2798_0, i_13_222_2887_0,
    i_13_222_2888_0, i_13_222_2959_0, i_13_222_3004_0, i_13_222_3050_0,
    i_13_222_3113_0, i_13_222_3262_0, i_13_222_3316_0, i_13_222_3464_0,
    i_13_222_3490_0, i_13_222_3535_0, i_13_222_3571_0, i_13_222_3604_0,
    i_13_222_3731_0, i_13_222_3733_0, i_13_222_3769_0, i_13_222_3770_0,
    i_13_222_3878_0, i_13_222_3904_0, i_13_222_3905_0, i_13_222_3910_0,
    i_13_222_4090_0, i_13_222_4091_0, i_13_222_4166_0, i_13_222_4211_0,
    i_13_222_4343_0, i_13_222_4358_0, i_13_222_4372_0, i_13_222_4373_0,
    i_13_222_4391_0, i_13_222_4433_0, i_13_222_4517_0, i_13_222_4586_0;
  output o_13_222_0_0;
  assign o_13_222_0_0 = ~(i_13_222_2544_0 | (~i_13_222_700_0 & ~i_13_222_3113_0) | (i_13_222_1996_0 & ~i_13_222_2303_0 & ~i_13_222_4166_0) | (~i_13_222_943_0 & ~i_13_222_950_0 & ~i_13_222_4091_0 & ~i_13_222_4373_0));
endmodule



// Benchmark "kernel_13_223" written by ABC on Sun Jul 19 10:48:32 2020

module kernel_13_223 ( 
    i_13_223_76_0, i_13_223_118_0, i_13_223_156_0, i_13_223_162_0,
    i_13_223_163_0, i_13_223_244_0, i_13_223_310_0, i_13_223_319_0,
    i_13_223_336_0, i_13_223_337_0, i_13_223_381_0, i_13_223_453_0,
    i_13_223_561_0, i_13_223_567_0, i_13_223_615_0, i_13_223_633_0,
    i_13_223_654_0, i_13_223_757_0, i_13_223_841_0, i_13_223_855_0,
    i_13_223_960_0, i_13_223_1063_0, i_13_223_1120_0, i_13_223_1218_0,
    i_13_223_1219_0, i_13_223_1300_0, i_13_223_1344_0, i_13_223_1434_0,
    i_13_223_1458_0, i_13_223_1522_0, i_13_223_1566_0, i_13_223_1593_0,
    i_13_223_1620_0, i_13_223_1693_0, i_13_223_1734_0, i_13_223_1783_0,
    i_13_223_1785_0, i_13_223_1786_0, i_13_223_1803_0, i_13_223_1813_0,
    i_13_223_1815_0, i_13_223_1816_0, i_13_223_1854_0, i_13_223_1992_0,
    i_13_223_2115_0, i_13_223_2116_0, i_13_223_2133_0, i_13_223_2205_0,
    i_13_223_2208_0, i_13_223_2212_0, i_13_223_2213_0, i_13_223_2403_0,
    i_13_223_2404_0, i_13_223_2421_0, i_13_223_2556_0, i_13_223_2584_0,
    i_13_223_2712_0, i_13_223_2935_0, i_13_223_2937_0, i_13_223_2938_0,
    i_13_223_3015_0, i_13_223_3034_0, i_13_223_3036_0, i_13_223_3060_0,
    i_13_223_3106_0, i_13_223_3145_0, i_13_223_3160_0, i_13_223_3213_0,
    i_13_223_3214_0, i_13_223_3216_0, i_13_223_3217_0, i_13_223_3220_0,
    i_13_223_3234_0, i_13_223_3268_0, i_13_223_3325_0, i_13_223_3438_0,
    i_13_223_3717_0, i_13_223_3741_0, i_13_223_3745_0, i_13_223_3816_0,
    i_13_223_3817_0, i_13_223_3843_0, i_13_223_3870_0, i_13_223_3884_0,
    i_13_223_3891_0, i_13_223_3982_0, i_13_223_4006_0, i_13_223_4041_0,
    i_13_223_4053_0, i_13_223_4207_0, i_13_223_4261_0, i_13_223_4302_0,
    i_13_223_4314_0, i_13_223_4321_0, i_13_223_4522_0, i_13_223_4530_0,
    i_13_223_4533_0, i_13_223_4582_0, i_13_223_4591_0, i_13_223_4600_0,
    o_13_223_0_0  );
  input  i_13_223_76_0, i_13_223_118_0, i_13_223_156_0, i_13_223_162_0,
    i_13_223_163_0, i_13_223_244_0, i_13_223_310_0, i_13_223_319_0,
    i_13_223_336_0, i_13_223_337_0, i_13_223_381_0, i_13_223_453_0,
    i_13_223_561_0, i_13_223_567_0, i_13_223_615_0, i_13_223_633_0,
    i_13_223_654_0, i_13_223_757_0, i_13_223_841_0, i_13_223_855_0,
    i_13_223_960_0, i_13_223_1063_0, i_13_223_1120_0, i_13_223_1218_0,
    i_13_223_1219_0, i_13_223_1300_0, i_13_223_1344_0, i_13_223_1434_0,
    i_13_223_1458_0, i_13_223_1522_0, i_13_223_1566_0, i_13_223_1593_0,
    i_13_223_1620_0, i_13_223_1693_0, i_13_223_1734_0, i_13_223_1783_0,
    i_13_223_1785_0, i_13_223_1786_0, i_13_223_1803_0, i_13_223_1813_0,
    i_13_223_1815_0, i_13_223_1816_0, i_13_223_1854_0, i_13_223_1992_0,
    i_13_223_2115_0, i_13_223_2116_0, i_13_223_2133_0, i_13_223_2205_0,
    i_13_223_2208_0, i_13_223_2212_0, i_13_223_2213_0, i_13_223_2403_0,
    i_13_223_2404_0, i_13_223_2421_0, i_13_223_2556_0, i_13_223_2584_0,
    i_13_223_2712_0, i_13_223_2935_0, i_13_223_2937_0, i_13_223_2938_0,
    i_13_223_3015_0, i_13_223_3034_0, i_13_223_3036_0, i_13_223_3060_0,
    i_13_223_3106_0, i_13_223_3145_0, i_13_223_3160_0, i_13_223_3213_0,
    i_13_223_3214_0, i_13_223_3216_0, i_13_223_3217_0, i_13_223_3220_0,
    i_13_223_3234_0, i_13_223_3268_0, i_13_223_3325_0, i_13_223_3438_0,
    i_13_223_3717_0, i_13_223_3741_0, i_13_223_3745_0, i_13_223_3816_0,
    i_13_223_3817_0, i_13_223_3843_0, i_13_223_3870_0, i_13_223_3884_0,
    i_13_223_3891_0, i_13_223_3982_0, i_13_223_4006_0, i_13_223_4041_0,
    i_13_223_4053_0, i_13_223_4207_0, i_13_223_4261_0, i_13_223_4302_0,
    i_13_223_4314_0, i_13_223_4321_0, i_13_223_4522_0, i_13_223_4530_0,
    i_13_223_4533_0, i_13_223_4582_0, i_13_223_4591_0, i_13_223_4600_0;
  output o_13_223_0_0;
  assign o_13_223_0_0 = ~((~i_13_223_3216_0 & (i_13_223_1120_0 | ~i_13_223_3214_0)) | (~i_13_223_4053_0 & (i_13_223_76_0 | ~i_13_223_3982_0)) | (~i_13_223_4041_0 & ((~i_13_223_337_0 & ~i_13_223_1522_0 & ~i_13_223_1815_0) | (~i_13_223_118_0 & ~i_13_223_1344_0 & ~i_13_223_1816_0) | (~i_13_223_1300_0 & ~i_13_223_3160_0))) | (i_13_223_319_0 & ~i_13_223_561_0 & ~i_13_223_3036_0) | (~i_13_223_2937_0 & i_13_223_3106_0 & i_13_223_3145_0) | (~i_13_223_2205_0 & ~i_13_223_3217_0));
endmodule



// Benchmark "kernel_13_224" written by ABC on Sun Jul 19 10:48:33 2020

module kernel_13_224 ( 
    i_13_224_41_0, i_13_224_74_0, i_13_224_76_0, i_13_224_103_0,
    i_13_224_112_0, i_13_224_113_0, i_13_224_184_0, i_13_224_185_0,
    i_13_224_193_0, i_13_224_208_0, i_13_224_316_0, i_13_224_317_0,
    i_13_224_374_0, i_13_224_571_0, i_13_224_572_0, i_13_224_575_0,
    i_13_224_643_0, i_13_224_644_0, i_13_224_685_0, i_13_224_689_0,
    i_13_224_715_0, i_13_224_778_0, i_13_224_811_0, i_13_224_814_0,
    i_13_224_895_0, i_13_224_982_0, i_13_224_983_0, i_13_224_1064_0,
    i_13_224_1067_0, i_13_224_1096_0, i_13_224_1102_0, i_13_224_1120_0,
    i_13_224_1121_0, i_13_224_1282_0, i_13_224_1507_0, i_13_224_1525_0,
    i_13_224_1678_0, i_13_224_1747_0, i_13_224_1750_0, i_13_224_1751_0,
    i_13_224_1804_0, i_13_224_1805_0, i_13_224_1829_0, i_13_224_1832_0,
    i_13_224_1834_0, i_13_224_1858_0, i_13_224_1907_0, i_13_224_1912_0,
    i_13_224_1921_0, i_13_224_2002_0, i_13_224_2044_0, i_13_224_2116_0,
    i_13_224_2120_0, i_13_224_2135_0, i_13_224_2137_0, i_13_224_2180_0,
    i_13_224_2264_0, i_13_224_2273_0, i_13_224_2404_0, i_13_224_2408_0,
    i_13_224_2434_0, i_13_224_2470_0, i_13_224_2542_0, i_13_224_2567_0,
    i_13_224_2651_0, i_13_224_2677_0, i_13_224_2692_0, i_13_224_2693_0,
    i_13_224_2696_0, i_13_224_2713_0, i_13_224_2737_0, i_13_224_2746_0,
    i_13_224_2747_0, i_13_224_2798_0, i_13_224_2920_0, i_13_224_2936_0,
    i_13_224_3206_0, i_13_224_3208_0, i_13_224_3209_0, i_13_224_3272_0,
    i_13_224_3406_0, i_13_224_3407_0, i_13_224_3427_0, i_13_224_3478_0,
    i_13_224_3607_0, i_13_224_3650_0, i_13_224_3686_0, i_13_224_3719_0,
    i_13_224_3817_0, i_13_224_3818_0, i_13_224_3854_0, i_13_224_3892_0,
    i_13_224_3989_0, i_13_224_4033_0, i_13_224_4036_0, i_13_224_4042_0,
    i_13_224_4141_0, i_13_224_4396_0, i_13_224_4421_0, i_13_224_4567_0,
    o_13_224_0_0  );
  input  i_13_224_41_0, i_13_224_74_0, i_13_224_76_0, i_13_224_103_0,
    i_13_224_112_0, i_13_224_113_0, i_13_224_184_0, i_13_224_185_0,
    i_13_224_193_0, i_13_224_208_0, i_13_224_316_0, i_13_224_317_0,
    i_13_224_374_0, i_13_224_571_0, i_13_224_572_0, i_13_224_575_0,
    i_13_224_643_0, i_13_224_644_0, i_13_224_685_0, i_13_224_689_0,
    i_13_224_715_0, i_13_224_778_0, i_13_224_811_0, i_13_224_814_0,
    i_13_224_895_0, i_13_224_982_0, i_13_224_983_0, i_13_224_1064_0,
    i_13_224_1067_0, i_13_224_1096_0, i_13_224_1102_0, i_13_224_1120_0,
    i_13_224_1121_0, i_13_224_1282_0, i_13_224_1507_0, i_13_224_1525_0,
    i_13_224_1678_0, i_13_224_1747_0, i_13_224_1750_0, i_13_224_1751_0,
    i_13_224_1804_0, i_13_224_1805_0, i_13_224_1829_0, i_13_224_1832_0,
    i_13_224_1834_0, i_13_224_1858_0, i_13_224_1907_0, i_13_224_1912_0,
    i_13_224_1921_0, i_13_224_2002_0, i_13_224_2044_0, i_13_224_2116_0,
    i_13_224_2120_0, i_13_224_2135_0, i_13_224_2137_0, i_13_224_2180_0,
    i_13_224_2264_0, i_13_224_2273_0, i_13_224_2404_0, i_13_224_2408_0,
    i_13_224_2434_0, i_13_224_2470_0, i_13_224_2542_0, i_13_224_2567_0,
    i_13_224_2651_0, i_13_224_2677_0, i_13_224_2692_0, i_13_224_2693_0,
    i_13_224_2696_0, i_13_224_2713_0, i_13_224_2737_0, i_13_224_2746_0,
    i_13_224_2747_0, i_13_224_2798_0, i_13_224_2920_0, i_13_224_2936_0,
    i_13_224_3206_0, i_13_224_3208_0, i_13_224_3209_0, i_13_224_3272_0,
    i_13_224_3406_0, i_13_224_3407_0, i_13_224_3427_0, i_13_224_3478_0,
    i_13_224_3607_0, i_13_224_3650_0, i_13_224_3686_0, i_13_224_3719_0,
    i_13_224_3817_0, i_13_224_3818_0, i_13_224_3854_0, i_13_224_3892_0,
    i_13_224_3989_0, i_13_224_4033_0, i_13_224_4036_0, i_13_224_4042_0,
    i_13_224_4141_0, i_13_224_4396_0, i_13_224_4421_0, i_13_224_4567_0;
  output o_13_224_0_0;
  assign o_13_224_0_0 = ~((~i_13_224_571_0 & (~i_13_224_1805_0 | ~i_13_224_1858_0)) | (~i_13_224_572_0 & ~i_13_224_811_0 & ~i_13_224_1747_0) | (~i_13_224_814_0 & i_13_224_1834_0) | (~i_13_224_1805_0 & ~i_13_224_2137_0) | (~i_13_224_2180_0 & ~i_13_224_2677_0) | (~i_13_224_1832_0 & i_13_224_3686_0 & i_13_224_3989_0) | (~i_13_224_1751_0 & ~i_13_224_3989_0));
endmodule



// Benchmark "kernel_13_225" written by ABC on Sun Jul 19 10:48:33 2020

module kernel_13_225 ( 
    i_13_225_51_0, i_13_225_69_0, i_13_225_153_0, i_13_225_169_0,
    i_13_225_186_0, i_13_225_283_0, i_13_225_285_0, i_13_225_286_0,
    i_13_225_310_0, i_13_225_318_0, i_13_225_319_0, i_13_225_328_0,
    i_13_225_364_0, i_13_225_384_0, i_13_225_385_0, i_13_225_448_0,
    i_13_225_569_0, i_13_225_625_0, i_13_225_642_0, i_13_225_646_0,
    i_13_225_673_0, i_13_225_681_0, i_13_225_688_0, i_13_225_690_0,
    i_13_225_697_0, i_13_225_759_0, i_13_225_816_0, i_13_225_817_0,
    i_13_225_844_0, i_13_225_1122_0, i_13_225_1254_0, i_13_225_1255_0,
    i_13_225_1303_0, i_13_225_1438_0, i_13_225_1542_0, i_13_225_1572_0,
    i_13_225_1599_0, i_13_225_1644_0, i_13_225_1677_0, i_13_225_1723_0,
    i_13_225_1777_0, i_13_225_1851_0, i_13_225_1852_0, i_13_225_1933_0,
    i_13_225_1954_0, i_13_225_2001_0, i_13_225_2055_0, i_13_225_2058_0,
    i_13_225_2119_0, i_13_225_2184_0, i_13_225_2280_0, i_13_225_2319_0,
    i_13_225_2407_0, i_13_225_2409_0, i_13_225_2410_0, i_13_225_2578_0,
    i_13_225_2614_0, i_13_225_2626_0, i_13_225_2679_0, i_13_225_2697_0,
    i_13_225_2698_0, i_13_225_2923_0, i_13_225_2940_0, i_13_225_2941_0,
    i_13_225_3112_0, i_13_225_3117_0, i_13_225_3129_0, i_13_225_3145_0,
    i_13_225_3210_0, i_13_225_3291_0, i_13_225_3399_0, i_13_225_3400_0,
    i_13_225_3417_0, i_13_225_3460_0, i_13_225_3541_0, i_13_225_3613_0,
    i_13_225_3705_0, i_13_225_3768_0, i_13_225_3820_0, i_13_225_3858_0,
    i_13_225_3993_0, i_13_225_3994_0, i_13_225_4021_0, i_13_225_4038_0,
    i_13_225_4056_0, i_13_225_4065_0, i_13_225_4066_0, i_13_225_4162_0,
    i_13_225_4308_0, i_13_225_4309_0, i_13_225_4317_0, i_13_225_4318_0,
    i_13_225_4341_0, i_13_225_4344_0, i_13_225_4378_0, i_13_225_4381_0,
    i_13_225_4440_0, i_13_225_4461_0, i_13_225_4594_0, i_13_225_4597_0,
    o_13_225_0_0  );
  input  i_13_225_51_0, i_13_225_69_0, i_13_225_153_0, i_13_225_169_0,
    i_13_225_186_0, i_13_225_283_0, i_13_225_285_0, i_13_225_286_0,
    i_13_225_310_0, i_13_225_318_0, i_13_225_319_0, i_13_225_328_0,
    i_13_225_364_0, i_13_225_384_0, i_13_225_385_0, i_13_225_448_0,
    i_13_225_569_0, i_13_225_625_0, i_13_225_642_0, i_13_225_646_0,
    i_13_225_673_0, i_13_225_681_0, i_13_225_688_0, i_13_225_690_0,
    i_13_225_697_0, i_13_225_759_0, i_13_225_816_0, i_13_225_817_0,
    i_13_225_844_0, i_13_225_1122_0, i_13_225_1254_0, i_13_225_1255_0,
    i_13_225_1303_0, i_13_225_1438_0, i_13_225_1542_0, i_13_225_1572_0,
    i_13_225_1599_0, i_13_225_1644_0, i_13_225_1677_0, i_13_225_1723_0,
    i_13_225_1777_0, i_13_225_1851_0, i_13_225_1852_0, i_13_225_1933_0,
    i_13_225_1954_0, i_13_225_2001_0, i_13_225_2055_0, i_13_225_2058_0,
    i_13_225_2119_0, i_13_225_2184_0, i_13_225_2280_0, i_13_225_2319_0,
    i_13_225_2407_0, i_13_225_2409_0, i_13_225_2410_0, i_13_225_2578_0,
    i_13_225_2614_0, i_13_225_2626_0, i_13_225_2679_0, i_13_225_2697_0,
    i_13_225_2698_0, i_13_225_2923_0, i_13_225_2940_0, i_13_225_2941_0,
    i_13_225_3112_0, i_13_225_3117_0, i_13_225_3129_0, i_13_225_3145_0,
    i_13_225_3210_0, i_13_225_3291_0, i_13_225_3399_0, i_13_225_3400_0,
    i_13_225_3417_0, i_13_225_3460_0, i_13_225_3541_0, i_13_225_3613_0,
    i_13_225_3705_0, i_13_225_3768_0, i_13_225_3820_0, i_13_225_3858_0,
    i_13_225_3993_0, i_13_225_3994_0, i_13_225_4021_0, i_13_225_4038_0,
    i_13_225_4056_0, i_13_225_4065_0, i_13_225_4066_0, i_13_225_4162_0,
    i_13_225_4308_0, i_13_225_4309_0, i_13_225_4317_0, i_13_225_4318_0,
    i_13_225_4341_0, i_13_225_4344_0, i_13_225_4378_0, i_13_225_4381_0,
    i_13_225_4440_0, i_13_225_4461_0, i_13_225_4594_0, i_13_225_4597_0;
  output o_13_225_0_0;
  assign o_13_225_0_0 = ~((~i_13_225_4317_0 & ((~i_13_225_384_0 & ~i_13_225_1851_0 & ~i_13_225_1852_0) | (~i_13_225_2280_0 & ~i_13_225_2410_0 & ~i_13_225_3768_0))) | (~i_13_225_3994_0 & ~i_13_225_4065_0 & ~i_13_225_4309_0));
endmodule



// Benchmark "kernel_13_226" written by ABC on Sun Jul 19 10:48:34 2020

module kernel_13_226 ( 
    i_13_226_91_0, i_13_226_94_0, i_13_226_114_0, i_13_226_118_0,
    i_13_226_121_0, i_13_226_123_0, i_13_226_136_0, i_13_226_190_0,
    i_13_226_231_0, i_13_226_276_0, i_13_226_376_0, i_13_226_396_0,
    i_13_226_474_0, i_13_226_517_0, i_13_226_597_0, i_13_226_609_0,
    i_13_226_732_0, i_13_226_793_0, i_13_226_832_0, i_13_226_840_0,
    i_13_226_841_0, i_13_226_861_0, i_13_226_862_0, i_13_226_879_0,
    i_13_226_913_0, i_13_226_950_0, i_13_226_1257_0, i_13_226_1272_0,
    i_13_226_1309_0, i_13_226_1491_0, i_13_226_1532_0, i_13_226_1599_0,
    i_13_226_1626_0, i_13_226_1736_0, i_13_226_1748_0, i_13_226_1786_0,
    i_13_226_1831_0, i_13_226_1839_0, i_13_226_1840_0, i_13_226_1842_0,
    i_13_226_1843_0, i_13_226_1930_0, i_13_226_1993_0, i_13_226_2117_0,
    i_13_226_2175_0, i_13_226_2206_0, i_13_226_2208_0, i_13_226_2211_0,
    i_13_226_2306_0, i_13_226_2361_0, i_13_226_2424_0, i_13_226_2426_0,
    i_13_226_2431_0, i_13_226_2436_0, i_13_226_2437_0, i_13_226_2459_0,
    i_13_226_2461_0, i_13_226_2463_0, i_13_226_2470_0, i_13_226_2541_0,
    i_13_226_2544_0, i_13_226_2616_0, i_13_226_2727_0, i_13_226_2744_0,
    i_13_226_3037_0, i_13_226_3163_0, i_13_226_3206_0, i_13_226_3369_0,
    i_13_226_3377_0, i_13_226_3422_0, i_13_226_3423_0, i_13_226_3426_0,
    i_13_226_3455_0, i_13_226_3530_0, i_13_226_3534_0, i_13_226_3651_0,
    i_13_226_3702_0, i_13_226_3849_0, i_13_226_3870_0, i_13_226_3871_0,
    i_13_226_3873_0, i_13_226_3874_0, i_13_226_3876_0, i_13_226_3877_0,
    i_13_226_3912_0, i_13_226_3991_0, i_13_226_4036_0, i_13_226_4086_0,
    i_13_226_4115_0, i_13_226_4180_0, i_13_226_4192_0, i_13_226_4206_0,
    i_13_226_4258_0, i_13_226_4271_0, i_13_226_4325_0, i_13_226_4349_0,
    i_13_226_4350_0, i_13_226_4351_0, i_13_226_4415_0, i_13_226_4582_0,
    o_13_226_0_0  );
  input  i_13_226_91_0, i_13_226_94_0, i_13_226_114_0, i_13_226_118_0,
    i_13_226_121_0, i_13_226_123_0, i_13_226_136_0, i_13_226_190_0,
    i_13_226_231_0, i_13_226_276_0, i_13_226_376_0, i_13_226_396_0,
    i_13_226_474_0, i_13_226_517_0, i_13_226_597_0, i_13_226_609_0,
    i_13_226_732_0, i_13_226_793_0, i_13_226_832_0, i_13_226_840_0,
    i_13_226_841_0, i_13_226_861_0, i_13_226_862_0, i_13_226_879_0,
    i_13_226_913_0, i_13_226_950_0, i_13_226_1257_0, i_13_226_1272_0,
    i_13_226_1309_0, i_13_226_1491_0, i_13_226_1532_0, i_13_226_1599_0,
    i_13_226_1626_0, i_13_226_1736_0, i_13_226_1748_0, i_13_226_1786_0,
    i_13_226_1831_0, i_13_226_1839_0, i_13_226_1840_0, i_13_226_1842_0,
    i_13_226_1843_0, i_13_226_1930_0, i_13_226_1993_0, i_13_226_2117_0,
    i_13_226_2175_0, i_13_226_2206_0, i_13_226_2208_0, i_13_226_2211_0,
    i_13_226_2306_0, i_13_226_2361_0, i_13_226_2424_0, i_13_226_2426_0,
    i_13_226_2431_0, i_13_226_2436_0, i_13_226_2437_0, i_13_226_2459_0,
    i_13_226_2461_0, i_13_226_2463_0, i_13_226_2470_0, i_13_226_2541_0,
    i_13_226_2544_0, i_13_226_2616_0, i_13_226_2727_0, i_13_226_2744_0,
    i_13_226_3037_0, i_13_226_3163_0, i_13_226_3206_0, i_13_226_3369_0,
    i_13_226_3377_0, i_13_226_3422_0, i_13_226_3423_0, i_13_226_3426_0,
    i_13_226_3455_0, i_13_226_3530_0, i_13_226_3534_0, i_13_226_3651_0,
    i_13_226_3702_0, i_13_226_3849_0, i_13_226_3870_0, i_13_226_3871_0,
    i_13_226_3873_0, i_13_226_3874_0, i_13_226_3876_0, i_13_226_3877_0,
    i_13_226_3912_0, i_13_226_3991_0, i_13_226_4036_0, i_13_226_4086_0,
    i_13_226_4115_0, i_13_226_4180_0, i_13_226_4192_0, i_13_226_4206_0,
    i_13_226_4258_0, i_13_226_4271_0, i_13_226_4325_0, i_13_226_4349_0,
    i_13_226_4350_0, i_13_226_4351_0, i_13_226_4415_0, i_13_226_4582_0;
  output o_13_226_0_0;
  assign o_13_226_0_0 = ~((~i_13_226_3534_0 & ((~i_13_226_2206_0 & ~i_13_226_2424_0) | (~i_13_226_1839_0 & ~i_13_226_3874_0 & i_13_226_4036_0))) | i_13_226_3206_0 | (i_13_226_841_0 & ~i_13_226_1626_0 & i_13_226_4036_0) | i_13_226_4258_0 | (i_13_226_840_0 & ~i_13_226_3423_0 & i_13_226_3870_0));
endmodule



// Benchmark "kernel_13_227" written by ABC on Sun Jul 19 10:48:35 2020

module kernel_13_227 ( 
    i_13_227_31_0, i_13_227_45_0, i_13_227_174_0, i_13_227_262_0,
    i_13_227_352_0, i_13_227_373_0, i_13_227_489_0, i_13_227_507_0,
    i_13_227_553_0, i_13_227_567_0, i_13_227_606_0, i_13_227_607_0,
    i_13_227_625_0, i_13_227_627_0, i_13_227_657_0, i_13_227_658_0,
    i_13_227_679_0, i_13_227_697_0, i_13_227_819_0, i_13_227_823_0,
    i_13_227_850_0, i_13_227_931_0, i_13_227_936_0, i_13_227_960_0,
    i_13_227_981_0, i_13_227_1021_0, i_13_227_1129_0, i_13_227_1224_0,
    i_13_227_1225_0, i_13_227_1228_0, i_13_227_1327_0, i_13_227_1359_0,
    i_13_227_1515_0, i_13_227_1522_0, i_13_227_1609_0, i_13_227_1677_0,
    i_13_227_1729_0, i_13_227_1732_0, i_13_227_1764_0, i_13_227_1767_0,
    i_13_227_1768_0, i_13_227_1771_0, i_13_227_1794_0, i_13_227_1795_0,
    i_13_227_1831_0, i_13_227_1832_0, i_13_227_2019_0, i_13_227_2020_0,
    i_13_227_2113_0, i_13_227_2120_0, i_13_227_2146_0, i_13_227_2237_0,
    i_13_227_2469_0, i_13_227_2470_0, i_13_227_2473_0, i_13_227_2541_0,
    i_13_227_2562_0, i_13_227_2566_0, i_13_227_2592_0, i_13_227_2767_0,
    i_13_227_2835_0, i_13_227_2848_0, i_13_227_2901_0, i_13_227_2908_0,
    i_13_227_2983_0, i_13_227_3028_0, i_13_227_3087_0, i_13_227_3123_0,
    i_13_227_3132_0, i_13_227_3208_0, i_13_227_3220_0, i_13_227_3234_0,
    i_13_227_3261_0, i_13_227_3262_0, i_13_227_3264_0, i_13_227_3270_0,
    i_13_227_3381_0, i_13_227_3417_0, i_13_227_3418_0, i_13_227_3483_0,
    i_13_227_3546_0, i_13_227_3613_0, i_13_227_3651_0, i_13_227_3720_0,
    i_13_227_3729_0, i_13_227_3730_0, i_13_227_3819_0, i_13_227_3820_0,
    i_13_227_3897_0, i_13_227_3901_0, i_13_227_3978_0, i_13_227_4035_0,
    i_13_227_4161_0, i_13_227_4162_0, i_13_227_4164_0, i_13_227_4321_0,
    i_13_227_4344_0, i_13_227_4350_0, i_13_227_4476_0, i_13_227_4603_0,
    o_13_227_0_0  );
  input  i_13_227_31_0, i_13_227_45_0, i_13_227_174_0, i_13_227_262_0,
    i_13_227_352_0, i_13_227_373_0, i_13_227_489_0, i_13_227_507_0,
    i_13_227_553_0, i_13_227_567_0, i_13_227_606_0, i_13_227_607_0,
    i_13_227_625_0, i_13_227_627_0, i_13_227_657_0, i_13_227_658_0,
    i_13_227_679_0, i_13_227_697_0, i_13_227_819_0, i_13_227_823_0,
    i_13_227_850_0, i_13_227_931_0, i_13_227_936_0, i_13_227_960_0,
    i_13_227_981_0, i_13_227_1021_0, i_13_227_1129_0, i_13_227_1224_0,
    i_13_227_1225_0, i_13_227_1228_0, i_13_227_1327_0, i_13_227_1359_0,
    i_13_227_1515_0, i_13_227_1522_0, i_13_227_1609_0, i_13_227_1677_0,
    i_13_227_1729_0, i_13_227_1732_0, i_13_227_1764_0, i_13_227_1767_0,
    i_13_227_1768_0, i_13_227_1771_0, i_13_227_1794_0, i_13_227_1795_0,
    i_13_227_1831_0, i_13_227_1832_0, i_13_227_2019_0, i_13_227_2020_0,
    i_13_227_2113_0, i_13_227_2120_0, i_13_227_2146_0, i_13_227_2237_0,
    i_13_227_2469_0, i_13_227_2470_0, i_13_227_2473_0, i_13_227_2541_0,
    i_13_227_2562_0, i_13_227_2566_0, i_13_227_2592_0, i_13_227_2767_0,
    i_13_227_2835_0, i_13_227_2848_0, i_13_227_2901_0, i_13_227_2908_0,
    i_13_227_2983_0, i_13_227_3028_0, i_13_227_3087_0, i_13_227_3123_0,
    i_13_227_3132_0, i_13_227_3208_0, i_13_227_3220_0, i_13_227_3234_0,
    i_13_227_3261_0, i_13_227_3262_0, i_13_227_3264_0, i_13_227_3270_0,
    i_13_227_3381_0, i_13_227_3417_0, i_13_227_3418_0, i_13_227_3483_0,
    i_13_227_3546_0, i_13_227_3613_0, i_13_227_3651_0, i_13_227_3720_0,
    i_13_227_3729_0, i_13_227_3730_0, i_13_227_3819_0, i_13_227_3820_0,
    i_13_227_3897_0, i_13_227_3901_0, i_13_227_3978_0, i_13_227_4035_0,
    i_13_227_4161_0, i_13_227_4162_0, i_13_227_4164_0, i_13_227_4321_0,
    i_13_227_4344_0, i_13_227_4350_0, i_13_227_4476_0, i_13_227_4603_0;
  output o_13_227_0_0;
  assign o_13_227_0_0 = ~((~i_13_227_4321_0 & ((~i_13_227_1677_0 & ~i_13_227_2237_0 & ~i_13_227_3483_0 & ~i_13_227_3819_0) | (i_13_227_697_0 & i_13_227_1732_0 & ~i_13_227_3978_0 & ~i_13_227_4161_0))) | (~i_13_227_3978_0 & ((~i_13_227_2020_0 & ~i_13_227_3261_0) | (~i_13_227_31_0 & ~i_13_227_1522_0 & ~i_13_227_3264_0 & ~i_13_227_3546_0 & ~i_13_227_3730_0 & ~i_13_227_4035_0))) | (~i_13_227_4161_0 & ((~i_13_227_489_0 & ~i_13_227_1729_0 & ~i_13_227_1795_0) | (~i_13_227_1327_0 & ~i_13_227_1764_0 & ~i_13_227_2019_0 & ~i_13_227_3234_0) | (~i_13_227_174_0 & i_13_227_4164_0))) | (i_13_227_2237_0 & ~i_13_227_2848_0 & ~i_13_227_3220_0));
endmodule



// Benchmark "kernel_13_228" written by ABC on Sun Jul 19 10:48:36 2020

module kernel_13_228 ( 
    i_13_228_73_0, i_13_228_94_0, i_13_228_96_0, i_13_228_120_0,
    i_13_228_192_0, i_13_228_199_0, i_13_228_228_0, i_13_228_323_0,
    i_13_228_373_0, i_13_228_380_0, i_13_228_441_0, i_13_228_485_0,
    i_13_228_492_0, i_13_228_526_0, i_13_228_570_0, i_13_228_588_0,
    i_13_228_593_0, i_13_228_647_0, i_13_228_661_0, i_13_228_712_0,
    i_13_228_714_0, i_13_228_735_0, i_13_228_819_0, i_13_228_841_0,
    i_13_228_858_0, i_13_228_899_0, i_13_228_917_0, i_13_228_948_0,
    i_13_228_950_0, i_13_228_1066_0, i_13_228_1080_0, i_13_228_1298_0,
    i_13_228_1327_0, i_13_228_1394_0, i_13_228_1400_0, i_13_228_1407_0,
    i_13_228_1443_0, i_13_228_1569_0, i_13_228_1570_0, i_13_228_1627_0,
    i_13_228_1639_0, i_13_228_1673_0, i_13_228_1691_0, i_13_228_1722_0,
    i_13_228_1800_0, i_13_228_1831_0, i_13_228_1956_0, i_13_228_2011_0,
    i_13_228_2141_0, i_13_228_2210_0, i_13_228_2238_0, i_13_228_2239_0,
    i_13_228_2281_0, i_13_228_2407_0, i_13_228_2424_0, i_13_228_2425_0,
    i_13_228_2474_0, i_13_228_2532_0, i_13_228_2589_0, i_13_228_2636_0,
    i_13_228_2705_0, i_13_228_2739_0, i_13_228_2874_0, i_13_228_2935_0,
    i_13_228_2955_0, i_13_228_2986_0, i_13_228_3024_0, i_13_228_3026_0,
    i_13_228_3240_0, i_13_228_3241_0, i_13_228_3258_0, i_13_228_3370_0,
    i_13_228_3395_0, i_13_228_3421_0, i_13_228_3424_0, i_13_228_3426_0,
    i_13_228_3450_0, i_13_228_3463_0, i_13_228_3521_0, i_13_228_3595_0,
    i_13_228_3666_0, i_13_228_3753_0, i_13_228_3791_0, i_13_228_3797_0,
    i_13_228_3842_0, i_13_228_3846_0, i_13_228_3873_0, i_13_228_3893_0,
    i_13_228_3918_0, i_13_228_3919_0, i_13_228_3932_0, i_13_228_3981_0,
    i_13_228_4008_0, i_13_228_4009_0, i_13_228_4043_0, i_13_228_4077_0,
    i_13_228_4090_0, i_13_228_4193_0, i_13_228_4353_0, i_13_228_4584_0,
    o_13_228_0_0  );
  input  i_13_228_73_0, i_13_228_94_0, i_13_228_96_0, i_13_228_120_0,
    i_13_228_192_0, i_13_228_199_0, i_13_228_228_0, i_13_228_323_0,
    i_13_228_373_0, i_13_228_380_0, i_13_228_441_0, i_13_228_485_0,
    i_13_228_492_0, i_13_228_526_0, i_13_228_570_0, i_13_228_588_0,
    i_13_228_593_0, i_13_228_647_0, i_13_228_661_0, i_13_228_712_0,
    i_13_228_714_0, i_13_228_735_0, i_13_228_819_0, i_13_228_841_0,
    i_13_228_858_0, i_13_228_899_0, i_13_228_917_0, i_13_228_948_0,
    i_13_228_950_0, i_13_228_1066_0, i_13_228_1080_0, i_13_228_1298_0,
    i_13_228_1327_0, i_13_228_1394_0, i_13_228_1400_0, i_13_228_1407_0,
    i_13_228_1443_0, i_13_228_1569_0, i_13_228_1570_0, i_13_228_1627_0,
    i_13_228_1639_0, i_13_228_1673_0, i_13_228_1691_0, i_13_228_1722_0,
    i_13_228_1800_0, i_13_228_1831_0, i_13_228_1956_0, i_13_228_2011_0,
    i_13_228_2141_0, i_13_228_2210_0, i_13_228_2238_0, i_13_228_2239_0,
    i_13_228_2281_0, i_13_228_2407_0, i_13_228_2424_0, i_13_228_2425_0,
    i_13_228_2474_0, i_13_228_2532_0, i_13_228_2589_0, i_13_228_2636_0,
    i_13_228_2705_0, i_13_228_2739_0, i_13_228_2874_0, i_13_228_2935_0,
    i_13_228_2955_0, i_13_228_2986_0, i_13_228_3024_0, i_13_228_3026_0,
    i_13_228_3240_0, i_13_228_3241_0, i_13_228_3258_0, i_13_228_3370_0,
    i_13_228_3395_0, i_13_228_3421_0, i_13_228_3424_0, i_13_228_3426_0,
    i_13_228_3450_0, i_13_228_3463_0, i_13_228_3521_0, i_13_228_3595_0,
    i_13_228_3666_0, i_13_228_3753_0, i_13_228_3791_0, i_13_228_3797_0,
    i_13_228_3842_0, i_13_228_3846_0, i_13_228_3873_0, i_13_228_3893_0,
    i_13_228_3918_0, i_13_228_3919_0, i_13_228_3932_0, i_13_228_3981_0,
    i_13_228_4008_0, i_13_228_4009_0, i_13_228_4043_0, i_13_228_4077_0,
    i_13_228_4090_0, i_13_228_4193_0, i_13_228_4353_0, i_13_228_4584_0;
  output o_13_228_0_0;
  assign o_13_228_0_0 = ~((i_13_228_3919_0 & ((~i_13_228_2874_0 & ~i_13_228_4009_0) | (~i_13_228_858_0 & ~i_13_228_4353_0))) | (~i_13_228_4009_0 & ((i_13_228_1570_0 & ~i_13_228_1627_0 & i_13_228_2407_0) | (~i_13_228_2532_0 & i_13_228_3595_0 & ~i_13_228_3753_0))) | (~i_13_228_2532_0 & ((~i_13_228_735_0 & ~i_13_228_1800_0 & ~i_13_228_3426_0 & ~i_13_228_3873_0) | (i_13_228_1956_0 & i_13_228_3918_0 & ~i_13_228_4077_0))) | (i_13_228_96_0 & ~i_13_228_570_0 & ~i_13_228_3424_0) | (i_13_228_841_0 & ~i_13_228_1407_0 & ~i_13_228_3918_0));
endmodule



// Benchmark "kernel_13_229" written by ABC on Sun Jul 19 10:48:37 2020

module kernel_13_229 ( 
    i_13_229_48_0, i_13_229_66_0, i_13_229_67_0, i_13_229_105_0,
    i_13_229_136_0, i_13_229_447_0, i_13_229_469_0, i_13_229_529_0,
    i_13_229_568_0, i_13_229_609_0, i_13_229_615_0, i_13_229_619_0,
    i_13_229_627_0, i_13_229_628_0, i_13_229_645_0, i_13_229_646_0,
    i_13_229_669_0, i_13_229_760_0, i_13_229_763_0, i_13_229_781_0,
    i_13_229_933_0, i_13_229_994_0, i_13_229_1074_0, i_13_229_1084_0,
    i_13_229_1086_0, i_13_229_1095_0, i_13_229_1122_0, i_13_229_1131_0,
    i_13_229_1132_0, i_13_229_1167_0, i_13_229_1317_0, i_13_229_1482_0,
    i_13_229_1483_0, i_13_229_1501_0, i_13_229_1525_0, i_13_229_1634_0,
    i_13_229_1645_0, i_13_229_1716_0, i_13_229_1752_0, i_13_229_1770_0,
    i_13_229_1788_0, i_13_229_1798_0, i_13_229_1806_0, i_13_229_1807_0,
    i_13_229_1857_0, i_13_229_1914_0, i_13_229_1995_0, i_13_229_2022_0,
    i_13_229_2023_0, i_13_229_2091_0, i_13_229_2122_0, i_13_229_2134_0,
    i_13_229_2291_0, i_13_229_2364_0, i_13_229_2462_0, i_13_229_2472_0,
    i_13_229_2473_0, i_13_229_2488_0, i_13_229_2515_0, i_13_229_2569_0,
    i_13_229_2581_0, i_13_229_2676_0, i_13_229_2722_0, i_13_229_2857_0,
    i_13_229_2909_0, i_13_229_2912_0, i_13_229_2940_0, i_13_229_2981_0,
    i_13_229_3030_0, i_13_229_3031_0, i_13_229_3076_0, i_13_229_3211_0,
    i_13_229_3264_0, i_13_229_3435_0, i_13_229_3459_0, i_13_229_3479_0,
    i_13_229_3487_0, i_13_229_3505_0, i_13_229_3669_0, i_13_229_3759_0,
    i_13_229_3783_0, i_13_229_3822_0, i_13_229_3856_0, i_13_229_3900_0,
    i_13_229_3901_0, i_13_229_3907_0, i_13_229_4017_0, i_13_229_4063_0,
    i_13_229_4101_0, i_13_229_4161_0, i_13_229_4164_0, i_13_229_4165_0,
    i_13_229_4270_0, i_13_229_4272_0, i_13_229_4296_0, i_13_229_4324_0,
    i_13_229_4416_0, i_13_229_4521_0, i_13_229_4523_0, i_13_229_4606_0,
    o_13_229_0_0  );
  input  i_13_229_48_0, i_13_229_66_0, i_13_229_67_0, i_13_229_105_0,
    i_13_229_136_0, i_13_229_447_0, i_13_229_469_0, i_13_229_529_0,
    i_13_229_568_0, i_13_229_609_0, i_13_229_615_0, i_13_229_619_0,
    i_13_229_627_0, i_13_229_628_0, i_13_229_645_0, i_13_229_646_0,
    i_13_229_669_0, i_13_229_760_0, i_13_229_763_0, i_13_229_781_0,
    i_13_229_933_0, i_13_229_994_0, i_13_229_1074_0, i_13_229_1084_0,
    i_13_229_1086_0, i_13_229_1095_0, i_13_229_1122_0, i_13_229_1131_0,
    i_13_229_1132_0, i_13_229_1167_0, i_13_229_1317_0, i_13_229_1482_0,
    i_13_229_1483_0, i_13_229_1501_0, i_13_229_1525_0, i_13_229_1634_0,
    i_13_229_1645_0, i_13_229_1716_0, i_13_229_1752_0, i_13_229_1770_0,
    i_13_229_1788_0, i_13_229_1798_0, i_13_229_1806_0, i_13_229_1807_0,
    i_13_229_1857_0, i_13_229_1914_0, i_13_229_1995_0, i_13_229_2022_0,
    i_13_229_2023_0, i_13_229_2091_0, i_13_229_2122_0, i_13_229_2134_0,
    i_13_229_2291_0, i_13_229_2364_0, i_13_229_2462_0, i_13_229_2472_0,
    i_13_229_2473_0, i_13_229_2488_0, i_13_229_2515_0, i_13_229_2569_0,
    i_13_229_2581_0, i_13_229_2676_0, i_13_229_2722_0, i_13_229_2857_0,
    i_13_229_2909_0, i_13_229_2912_0, i_13_229_2940_0, i_13_229_2981_0,
    i_13_229_3030_0, i_13_229_3031_0, i_13_229_3076_0, i_13_229_3211_0,
    i_13_229_3264_0, i_13_229_3435_0, i_13_229_3459_0, i_13_229_3479_0,
    i_13_229_3487_0, i_13_229_3505_0, i_13_229_3669_0, i_13_229_3759_0,
    i_13_229_3783_0, i_13_229_3822_0, i_13_229_3856_0, i_13_229_3900_0,
    i_13_229_3901_0, i_13_229_3907_0, i_13_229_4017_0, i_13_229_4063_0,
    i_13_229_4101_0, i_13_229_4161_0, i_13_229_4164_0, i_13_229_4165_0,
    i_13_229_4270_0, i_13_229_4272_0, i_13_229_4296_0, i_13_229_4324_0,
    i_13_229_4416_0, i_13_229_4521_0, i_13_229_4523_0, i_13_229_4606_0;
  output o_13_229_0_0;
  assign o_13_229_0_0 = ~((~i_13_229_1716_0 & ((~i_13_229_615_0 & ~i_13_229_2022_0) | (i_13_229_1084_0 & ~i_13_229_4164_0))) | ~i_13_229_3264_0 | (~i_13_229_619_0 & ~i_13_229_2023_0));
endmodule



// Benchmark "kernel_13_230" written by ABC on Sun Jul 19 10:48:38 2020

module kernel_13_230 ( 
    i_13_230_26_0, i_13_230_38_0, i_13_230_40_0, i_13_230_79_0,
    i_13_230_103_0, i_13_230_105_0, i_13_230_266_0, i_13_230_431_0,
    i_13_230_599_0, i_13_230_607_0, i_13_230_677_0, i_13_230_679_0,
    i_13_230_685_0, i_13_230_686_0, i_13_230_717_0, i_13_230_761_0,
    i_13_230_778_0, i_13_230_815_0, i_13_230_816_0, i_13_230_839_0,
    i_13_230_895_0, i_13_230_924_0, i_13_230_983_0, i_13_230_1088_0,
    i_13_230_1150_0, i_13_230_1187_0, i_13_230_1270_0, i_13_230_1271_0,
    i_13_230_1437_0, i_13_230_1456_0, i_13_230_1462_0, i_13_230_1490_0,
    i_13_230_1518_0, i_13_230_1571_0, i_13_230_1594_0, i_13_230_1655_0,
    i_13_230_1747_0, i_13_230_1748_0, i_13_230_1750_0, i_13_230_1751_0,
    i_13_230_1805_0, i_13_230_1806_0, i_13_230_1815_0, i_13_230_1841_0,
    i_13_230_1856_0, i_13_230_1858_0, i_13_230_1909_0, i_13_230_1914_0,
    i_13_230_2047_0, i_13_230_2049_0, i_13_230_2112_0, i_13_230_2137_0,
    i_13_230_2138_0, i_13_230_2139_0, i_13_230_2140_0, i_13_230_2141_0,
    i_13_230_2224_0, i_13_230_2354_0, i_13_230_2357_0, i_13_230_2407_0,
    i_13_230_2408_0, i_13_230_2557_0, i_13_230_2562_0, i_13_230_2579_0,
    i_13_230_2650_0, i_13_230_2651_0, i_13_230_2652_0, i_13_230_2692_0,
    i_13_230_2722_0, i_13_230_2749_0, i_13_230_2750_0, i_13_230_2751_0,
    i_13_230_2752_0, i_13_230_2822_0, i_13_230_2823_0, i_13_230_2939_0,
    i_13_230_2999_0, i_13_230_3206_0, i_13_230_3208_0, i_13_230_3273_0,
    i_13_230_3290_0, i_13_230_3374_0, i_13_230_3430_0, i_13_230_3449_0,
    i_13_230_3533_0, i_13_230_3534_0, i_13_230_3556_0, i_13_230_3876_0,
    i_13_230_3911_0, i_13_230_3912_0, i_13_230_3943_0, i_13_230_3989_0,
    i_13_230_3991_0, i_13_230_4048_0, i_13_230_4161_0, i_13_230_4187_0,
    i_13_230_4309_0, i_13_230_4369_0, i_13_230_4381_0, i_13_230_4426_0,
    o_13_230_0_0  );
  input  i_13_230_26_0, i_13_230_38_0, i_13_230_40_0, i_13_230_79_0,
    i_13_230_103_0, i_13_230_105_0, i_13_230_266_0, i_13_230_431_0,
    i_13_230_599_0, i_13_230_607_0, i_13_230_677_0, i_13_230_679_0,
    i_13_230_685_0, i_13_230_686_0, i_13_230_717_0, i_13_230_761_0,
    i_13_230_778_0, i_13_230_815_0, i_13_230_816_0, i_13_230_839_0,
    i_13_230_895_0, i_13_230_924_0, i_13_230_983_0, i_13_230_1088_0,
    i_13_230_1150_0, i_13_230_1187_0, i_13_230_1270_0, i_13_230_1271_0,
    i_13_230_1437_0, i_13_230_1456_0, i_13_230_1462_0, i_13_230_1490_0,
    i_13_230_1518_0, i_13_230_1571_0, i_13_230_1594_0, i_13_230_1655_0,
    i_13_230_1747_0, i_13_230_1748_0, i_13_230_1750_0, i_13_230_1751_0,
    i_13_230_1805_0, i_13_230_1806_0, i_13_230_1815_0, i_13_230_1841_0,
    i_13_230_1856_0, i_13_230_1858_0, i_13_230_1909_0, i_13_230_1914_0,
    i_13_230_2047_0, i_13_230_2049_0, i_13_230_2112_0, i_13_230_2137_0,
    i_13_230_2138_0, i_13_230_2139_0, i_13_230_2140_0, i_13_230_2141_0,
    i_13_230_2224_0, i_13_230_2354_0, i_13_230_2357_0, i_13_230_2407_0,
    i_13_230_2408_0, i_13_230_2557_0, i_13_230_2562_0, i_13_230_2579_0,
    i_13_230_2650_0, i_13_230_2651_0, i_13_230_2652_0, i_13_230_2692_0,
    i_13_230_2722_0, i_13_230_2749_0, i_13_230_2750_0, i_13_230_2751_0,
    i_13_230_2752_0, i_13_230_2822_0, i_13_230_2823_0, i_13_230_2939_0,
    i_13_230_2999_0, i_13_230_3206_0, i_13_230_3208_0, i_13_230_3273_0,
    i_13_230_3290_0, i_13_230_3374_0, i_13_230_3430_0, i_13_230_3449_0,
    i_13_230_3533_0, i_13_230_3534_0, i_13_230_3556_0, i_13_230_3876_0,
    i_13_230_3911_0, i_13_230_3912_0, i_13_230_3943_0, i_13_230_3989_0,
    i_13_230_3991_0, i_13_230_4048_0, i_13_230_4161_0, i_13_230_4187_0,
    i_13_230_4309_0, i_13_230_4369_0, i_13_230_4381_0, i_13_230_4426_0;
  output o_13_230_0_0;
  assign o_13_230_0_0 = ~(~i_13_230_2939_0 | ~i_13_230_3989_0);
endmodule



// Benchmark "kernel_13_231" written by ABC on Sun Jul 19 10:48:38 2020

module kernel_13_231 ( 
    i_13_231_76_0, i_13_231_106_0, i_13_231_107_0, i_13_231_139_0,
    i_13_231_170_0, i_13_231_229_0, i_13_231_232_0, i_13_231_269_0,
    i_13_231_313_0, i_13_231_340_0, i_13_231_357_0, i_13_231_395_0,
    i_13_231_510_0, i_13_231_515_0, i_13_231_524_0, i_13_231_667_0,
    i_13_231_691_0, i_13_231_695_0, i_13_231_817_0, i_13_231_818_0,
    i_13_231_820_0, i_13_231_911_0, i_13_231_980_0, i_13_231_1069_0,
    i_13_231_1070_0, i_13_231_1208_0, i_13_231_1217_0, i_13_231_1222_0,
    i_13_231_1307_0, i_13_231_1316_0, i_13_231_1329_0, i_13_231_1330_0,
    i_13_231_1489_0, i_13_231_1573_0, i_13_231_1750_0, i_13_231_1807_0,
    i_13_231_1808_0, i_13_231_1815_0, i_13_231_1852_0, i_13_231_1882_0,
    i_13_231_1912_0, i_13_231_1999_0, i_13_231_2000_0, i_13_231_2059_0,
    i_13_231_2125_0, i_13_231_2126_0, i_13_231_2135_0, i_13_231_2139_0,
    i_13_231_2140_0, i_13_231_2185_0, i_13_231_2188_0, i_13_231_2225_0,
    i_13_231_2380_0, i_13_231_2409_0, i_13_231_2410_0, i_13_231_2411_0,
    i_13_231_2536_0, i_13_231_2586_0, i_13_231_2614_0, i_13_231_2656_0,
    i_13_231_2698_0, i_13_231_2722_0, i_13_231_2744_0, i_13_231_2751_0,
    i_13_231_2752_0, i_13_231_2797_0, i_13_231_2941_0, i_13_231_3003_0,
    i_13_231_3208_0, i_13_231_3220_0, i_13_231_3237_0, i_13_231_3238_0,
    i_13_231_3269_0, i_13_231_3273_0, i_13_231_3291_0, i_13_231_3292_0,
    i_13_231_3346_0, i_13_231_3372_0, i_13_231_3373_0, i_13_231_3505_0,
    i_13_231_3532_0, i_13_231_3538_0, i_13_231_3539_0, i_13_231_3727_0,
    i_13_231_3728_0, i_13_231_3853_0, i_13_231_3877_0, i_13_231_3895_0,
    i_13_231_3910_0, i_13_231_4021_0, i_13_231_4048_0, i_13_231_4063_0,
    i_13_231_4065_0, i_13_231_4066_0, i_13_231_4088_0, i_13_231_4252_0,
    i_13_231_4274_0, i_13_231_4318_0, i_13_231_4319_0, i_13_231_4448_0,
    o_13_231_0_0  );
  input  i_13_231_76_0, i_13_231_106_0, i_13_231_107_0, i_13_231_139_0,
    i_13_231_170_0, i_13_231_229_0, i_13_231_232_0, i_13_231_269_0,
    i_13_231_313_0, i_13_231_340_0, i_13_231_357_0, i_13_231_395_0,
    i_13_231_510_0, i_13_231_515_0, i_13_231_524_0, i_13_231_667_0,
    i_13_231_691_0, i_13_231_695_0, i_13_231_817_0, i_13_231_818_0,
    i_13_231_820_0, i_13_231_911_0, i_13_231_980_0, i_13_231_1069_0,
    i_13_231_1070_0, i_13_231_1208_0, i_13_231_1217_0, i_13_231_1222_0,
    i_13_231_1307_0, i_13_231_1316_0, i_13_231_1329_0, i_13_231_1330_0,
    i_13_231_1489_0, i_13_231_1573_0, i_13_231_1750_0, i_13_231_1807_0,
    i_13_231_1808_0, i_13_231_1815_0, i_13_231_1852_0, i_13_231_1882_0,
    i_13_231_1912_0, i_13_231_1999_0, i_13_231_2000_0, i_13_231_2059_0,
    i_13_231_2125_0, i_13_231_2126_0, i_13_231_2135_0, i_13_231_2139_0,
    i_13_231_2140_0, i_13_231_2185_0, i_13_231_2188_0, i_13_231_2225_0,
    i_13_231_2380_0, i_13_231_2409_0, i_13_231_2410_0, i_13_231_2411_0,
    i_13_231_2536_0, i_13_231_2586_0, i_13_231_2614_0, i_13_231_2656_0,
    i_13_231_2698_0, i_13_231_2722_0, i_13_231_2744_0, i_13_231_2751_0,
    i_13_231_2752_0, i_13_231_2797_0, i_13_231_2941_0, i_13_231_3003_0,
    i_13_231_3208_0, i_13_231_3220_0, i_13_231_3237_0, i_13_231_3238_0,
    i_13_231_3269_0, i_13_231_3273_0, i_13_231_3291_0, i_13_231_3292_0,
    i_13_231_3346_0, i_13_231_3372_0, i_13_231_3373_0, i_13_231_3505_0,
    i_13_231_3532_0, i_13_231_3538_0, i_13_231_3539_0, i_13_231_3727_0,
    i_13_231_3728_0, i_13_231_3853_0, i_13_231_3877_0, i_13_231_3895_0,
    i_13_231_3910_0, i_13_231_4021_0, i_13_231_4048_0, i_13_231_4063_0,
    i_13_231_4065_0, i_13_231_4066_0, i_13_231_4088_0, i_13_231_4252_0,
    i_13_231_4274_0, i_13_231_4318_0, i_13_231_4319_0, i_13_231_4448_0;
  output o_13_231_0_0;
  assign o_13_231_0_0 = ~(~i_13_231_2410_0);
endmodule



// Benchmark "kernel_13_232" written by ABC on Sun Jul 19 10:48:39 2020

module kernel_13_232 ( 
    i_13_232_39_0, i_13_232_40_0, i_13_232_43_0, i_13_232_105_0,
    i_13_232_114_0, i_13_232_186_0, i_13_232_187_0, i_13_232_373_0,
    i_13_232_445_0, i_13_232_529_0, i_13_232_533_0, i_13_232_547_0,
    i_13_232_556_0, i_13_232_573_0, i_13_232_600_0, i_13_232_607_0,
    i_13_232_629_0, i_13_232_682_0, i_13_232_717_0, i_13_232_732_0,
    i_13_232_780_0, i_13_232_817_0, i_13_232_897_0, i_13_232_940_0,
    i_13_232_1069_0, i_13_232_1084_0, i_13_232_1123_0, i_13_232_1159_0,
    i_13_232_1210_0, i_13_232_1266_0, i_13_232_1276_0, i_13_232_1464_0,
    i_13_232_1465_0, i_13_232_1482_0, i_13_232_1483_0, i_13_232_1501_0,
    i_13_232_1502_0, i_13_232_1645_0, i_13_232_1677_0, i_13_232_1690_0,
    i_13_232_1732_0, i_13_232_1749_0, i_13_232_1750_0, i_13_232_1752_0,
    i_13_232_1753_0, i_13_232_1770_0, i_13_232_1776_0, i_13_232_1788_0,
    i_13_232_1806_0, i_13_232_1807_0, i_13_232_1826_0, i_13_232_1862_0,
    i_13_232_1914_0, i_13_232_2051_0, i_13_232_2122_0, i_13_232_2139_0,
    i_13_232_2140_0, i_13_232_2149_0, i_13_232_2266_0, i_13_232_2310_0,
    i_13_232_2365_0, i_13_232_2582_0, i_13_232_2653_0, i_13_232_2722_0,
    i_13_232_2751_0, i_13_232_2752_0, i_13_232_2823_0, i_13_232_2824_0,
    i_13_232_2874_0, i_13_232_2883_0, i_13_232_2940_0, i_13_232_2941_0,
    i_13_232_2983_0, i_13_232_3030_0, i_13_232_3032_0, i_13_232_3119_0,
    i_13_232_3121_0, i_13_232_3122_0, i_13_232_3293_0, i_13_232_3345_0,
    i_13_232_3373_0, i_13_232_3400_0, i_13_232_3417_0, i_13_232_3418_0,
    i_13_232_3471_0, i_13_232_3525_0, i_13_232_3526_0, i_13_232_3562_0,
    i_13_232_3864_0, i_13_232_3895_0, i_13_232_3994_0, i_13_232_4047_0,
    i_13_232_4049_0, i_13_232_4080_0, i_13_232_4101_0, i_13_232_4156_0,
    i_13_232_4272_0, i_13_232_4318_0, i_13_232_4381_0, i_13_232_4443_0,
    o_13_232_0_0  );
  input  i_13_232_39_0, i_13_232_40_0, i_13_232_43_0, i_13_232_105_0,
    i_13_232_114_0, i_13_232_186_0, i_13_232_187_0, i_13_232_373_0,
    i_13_232_445_0, i_13_232_529_0, i_13_232_533_0, i_13_232_547_0,
    i_13_232_556_0, i_13_232_573_0, i_13_232_600_0, i_13_232_607_0,
    i_13_232_629_0, i_13_232_682_0, i_13_232_717_0, i_13_232_732_0,
    i_13_232_780_0, i_13_232_817_0, i_13_232_897_0, i_13_232_940_0,
    i_13_232_1069_0, i_13_232_1084_0, i_13_232_1123_0, i_13_232_1159_0,
    i_13_232_1210_0, i_13_232_1266_0, i_13_232_1276_0, i_13_232_1464_0,
    i_13_232_1465_0, i_13_232_1482_0, i_13_232_1483_0, i_13_232_1501_0,
    i_13_232_1502_0, i_13_232_1645_0, i_13_232_1677_0, i_13_232_1690_0,
    i_13_232_1732_0, i_13_232_1749_0, i_13_232_1750_0, i_13_232_1752_0,
    i_13_232_1753_0, i_13_232_1770_0, i_13_232_1776_0, i_13_232_1788_0,
    i_13_232_1806_0, i_13_232_1807_0, i_13_232_1826_0, i_13_232_1862_0,
    i_13_232_1914_0, i_13_232_2051_0, i_13_232_2122_0, i_13_232_2139_0,
    i_13_232_2140_0, i_13_232_2149_0, i_13_232_2266_0, i_13_232_2310_0,
    i_13_232_2365_0, i_13_232_2582_0, i_13_232_2653_0, i_13_232_2722_0,
    i_13_232_2751_0, i_13_232_2752_0, i_13_232_2823_0, i_13_232_2824_0,
    i_13_232_2874_0, i_13_232_2883_0, i_13_232_2940_0, i_13_232_2941_0,
    i_13_232_2983_0, i_13_232_3030_0, i_13_232_3032_0, i_13_232_3119_0,
    i_13_232_3121_0, i_13_232_3122_0, i_13_232_3293_0, i_13_232_3345_0,
    i_13_232_3373_0, i_13_232_3400_0, i_13_232_3417_0, i_13_232_3418_0,
    i_13_232_3471_0, i_13_232_3525_0, i_13_232_3526_0, i_13_232_3562_0,
    i_13_232_3864_0, i_13_232_3895_0, i_13_232_3994_0, i_13_232_4047_0,
    i_13_232_4049_0, i_13_232_4080_0, i_13_232_4101_0, i_13_232_4156_0,
    i_13_232_4272_0, i_13_232_4318_0, i_13_232_4381_0, i_13_232_4443_0;
  output o_13_232_0_0;
  assign o_13_232_0_0 = ~((~i_13_232_3345_0 & ((~i_13_232_2140_0 & ~i_13_232_2149_0) | (~i_13_232_2941_0 & ~i_13_232_3994_0))) | (~i_13_232_186_0 & ~i_13_232_940_0 & ~i_13_232_1862_0));
endmodule



// Benchmark "kernel_13_233" written by ABC on Sun Jul 19 10:48:40 2020

module kernel_13_233 ( 
    i_13_233_48_0, i_13_233_165_0, i_13_233_211_0, i_13_233_217_0,
    i_13_233_441_0, i_13_233_531_0, i_13_233_532_0, i_13_233_558_0,
    i_13_233_570_0, i_13_233_640_0, i_13_233_676_0, i_13_233_679_0,
    i_13_233_837_0, i_13_233_928_0, i_13_233_931_0, i_13_233_945_0,
    i_13_233_1098_0, i_13_233_1117_0, i_13_233_1270_0, i_13_233_1380_0,
    i_13_233_1381_0, i_13_233_1396_0, i_13_233_1399_0, i_13_233_1434_0,
    i_13_233_1471_0, i_13_233_1530_0, i_13_233_1593_0, i_13_233_1657_0,
    i_13_233_1674_0, i_13_233_1719_0, i_13_233_1746_0, i_13_233_1777_0,
    i_13_233_1791_0, i_13_233_1792_0, i_13_233_1795_0, i_13_233_1908_0,
    i_13_233_1917_0, i_13_233_1930_0, i_13_233_2011_0, i_13_233_2016_0,
    i_13_233_2046_0, i_13_233_2115_0, i_13_233_2191_0, i_13_233_2259_0,
    i_13_233_2397_0, i_13_233_2466_0, i_13_233_2505_0, i_13_233_2673_0,
    i_13_233_2722_0, i_13_233_2748_0, i_13_233_2749_0, i_13_233_2818_0,
    i_13_233_2844_0, i_13_233_2857_0, i_13_233_2901_0, i_13_233_2911_0,
    i_13_233_2916_0, i_13_233_3024_0, i_13_233_3025_0, i_13_233_3060_0,
    i_13_233_3069_0, i_13_233_3090_0, i_13_233_3258_0, i_13_233_3348_0,
    i_13_233_3349_0, i_13_233_3375_0, i_13_233_3414_0, i_13_233_3415_0,
    i_13_233_3421_0, i_13_233_3532_0, i_13_233_3573_0, i_13_233_3685_0,
    i_13_233_3735_0, i_13_233_3765_0, i_13_233_3766_0, i_13_233_3783_0,
    i_13_233_3784_0, i_13_233_3846_0, i_13_233_3855_0, i_13_233_3862_0,
    i_13_233_3888_0, i_13_233_3924_0, i_13_233_3925_0, i_13_233_3987_0,
    i_13_233_3988_0, i_13_233_4054_0, i_13_233_4077_0, i_13_233_4086_0,
    i_13_233_4122_0, i_13_233_4123_0, i_13_233_4203_0, i_13_233_4204_0,
    i_13_233_4212_0, i_13_233_4447_0, i_13_233_4590_0, i_13_233_4591_0,
    i_13_233_4594_0, i_13_233_4599_0, i_13_233_4600_0, i_13_233_4604_0,
    o_13_233_0_0  );
  input  i_13_233_48_0, i_13_233_165_0, i_13_233_211_0, i_13_233_217_0,
    i_13_233_441_0, i_13_233_531_0, i_13_233_532_0, i_13_233_558_0,
    i_13_233_570_0, i_13_233_640_0, i_13_233_676_0, i_13_233_679_0,
    i_13_233_837_0, i_13_233_928_0, i_13_233_931_0, i_13_233_945_0,
    i_13_233_1098_0, i_13_233_1117_0, i_13_233_1270_0, i_13_233_1380_0,
    i_13_233_1381_0, i_13_233_1396_0, i_13_233_1399_0, i_13_233_1434_0,
    i_13_233_1471_0, i_13_233_1530_0, i_13_233_1593_0, i_13_233_1657_0,
    i_13_233_1674_0, i_13_233_1719_0, i_13_233_1746_0, i_13_233_1777_0,
    i_13_233_1791_0, i_13_233_1792_0, i_13_233_1795_0, i_13_233_1908_0,
    i_13_233_1917_0, i_13_233_1930_0, i_13_233_2011_0, i_13_233_2016_0,
    i_13_233_2046_0, i_13_233_2115_0, i_13_233_2191_0, i_13_233_2259_0,
    i_13_233_2397_0, i_13_233_2466_0, i_13_233_2505_0, i_13_233_2673_0,
    i_13_233_2722_0, i_13_233_2748_0, i_13_233_2749_0, i_13_233_2818_0,
    i_13_233_2844_0, i_13_233_2857_0, i_13_233_2901_0, i_13_233_2911_0,
    i_13_233_2916_0, i_13_233_3024_0, i_13_233_3025_0, i_13_233_3060_0,
    i_13_233_3069_0, i_13_233_3090_0, i_13_233_3258_0, i_13_233_3348_0,
    i_13_233_3349_0, i_13_233_3375_0, i_13_233_3414_0, i_13_233_3415_0,
    i_13_233_3421_0, i_13_233_3532_0, i_13_233_3573_0, i_13_233_3685_0,
    i_13_233_3735_0, i_13_233_3765_0, i_13_233_3766_0, i_13_233_3783_0,
    i_13_233_3784_0, i_13_233_3846_0, i_13_233_3855_0, i_13_233_3862_0,
    i_13_233_3888_0, i_13_233_3924_0, i_13_233_3925_0, i_13_233_3987_0,
    i_13_233_3988_0, i_13_233_4054_0, i_13_233_4077_0, i_13_233_4086_0,
    i_13_233_4122_0, i_13_233_4123_0, i_13_233_4203_0, i_13_233_4204_0,
    i_13_233_4212_0, i_13_233_4447_0, i_13_233_4590_0, i_13_233_4591_0,
    i_13_233_4594_0, i_13_233_4599_0, i_13_233_4600_0, i_13_233_4604_0;
  output o_13_233_0_0;
  assign o_13_233_0_0 = ~((~i_13_233_3924_0 & (~i_13_233_532_0 | ~i_13_233_1792_0)) | (~i_13_233_676_0 & ~i_13_233_1746_0 & ~i_13_233_3987_0 & ~i_13_233_4086_0));
endmodule



// Benchmark "kernel_13_234" written by ABC on Sun Jul 19 10:48:41 2020

module kernel_13_234 ( 
    i_13_234_81_0, i_13_234_137_0, i_13_234_140_0, i_13_234_142_0,
    i_13_234_143_0, i_13_234_166_0, i_13_234_232_0, i_13_234_279_0,
    i_13_234_280_0, i_13_234_355_0, i_13_234_454_0, i_13_234_534_0,
    i_13_234_539_0, i_13_234_582_0, i_13_234_595_0, i_13_234_603_0,
    i_13_234_611_0, i_13_234_620_0, i_13_234_691_0, i_13_234_700_0,
    i_13_234_725_0, i_13_234_726_0, i_13_234_780_0, i_13_234_824_0,
    i_13_234_894_0, i_13_234_1215_0, i_13_234_1222_0, i_13_234_1276_0,
    i_13_234_1277_0, i_13_234_1486_0, i_13_234_1498_0, i_13_234_1552_0,
    i_13_234_1678_0, i_13_234_1710_0, i_13_234_1711_0, i_13_234_1714_0,
    i_13_234_1715_0, i_13_234_1722_0, i_13_234_1725_0, i_13_234_1726_0,
    i_13_234_1727_0, i_13_234_1731_0, i_13_234_1761_0, i_13_234_1780_0,
    i_13_234_1781_0, i_13_234_1846_0, i_13_234_1881_0, i_13_234_1884_0,
    i_13_234_1885_0, i_13_234_1886_0, i_13_234_1888_0, i_13_234_1889_0,
    i_13_234_1999_0, i_13_234_2009_0, i_13_234_2158_0, i_13_234_2380_0,
    i_13_234_2461_0, i_13_234_2462_0, i_13_234_2470_0, i_13_234_2629_0,
    i_13_234_2647_0, i_13_234_2650_0, i_13_234_2651_0, i_13_234_2714_0,
    i_13_234_2848_0, i_13_234_2849_0, i_13_234_2875_0, i_13_234_2878_0,
    i_13_234_2887_0, i_13_234_2916_0, i_13_234_2917_0, i_13_234_3004_0,
    i_13_234_3040_0, i_13_234_3041_0, i_13_234_3109_0, i_13_234_3145_0,
    i_13_234_3146_0, i_13_234_3293_0, i_13_234_3406_0, i_13_234_3429_0,
    i_13_234_3689_0, i_13_234_3707_0, i_13_234_3781_0, i_13_234_3794_0,
    i_13_234_3964_0, i_13_234_4083_0, i_13_234_4095_0, i_13_234_4096_0,
    i_13_234_4100_0, i_13_234_4153_0, i_13_234_4190_0, i_13_234_4253_0,
    i_13_234_4390_0, i_13_234_4414_0, i_13_234_4426_0, i_13_234_4437_0,
    i_13_234_4440_0, i_13_234_4513_0, i_13_234_4519_0, i_13_234_4526_0,
    o_13_234_0_0  );
  input  i_13_234_81_0, i_13_234_137_0, i_13_234_140_0, i_13_234_142_0,
    i_13_234_143_0, i_13_234_166_0, i_13_234_232_0, i_13_234_279_0,
    i_13_234_280_0, i_13_234_355_0, i_13_234_454_0, i_13_234_534_0,
    i_13_234_539_0, i_13_234_582_0, i_13_234_595_0, i_13_234_603_0,
    i_13_234_611_0, i_13_234_620_0, i_13_234_691_0, i_13_234_700_0,
    i_13_234_725_0, i_13_234_726_0, i_13_234_780_0, i_13_234_824_0,
    i_13_234_894_0, i_13_234_1215_0, i_13_234_1222_0, i_13_234_1276_0,
    i_13_234_1277_0, i_13_234_1486_0, i_13_234_1498_0, i_13_234_1552_0,
    i_13_234_1678_0, i_13_234_1710_0, i_13_234_1711_0, i_13_234_1714_0,
    i_13_234_1715_0, i_13_234_1722_0, i_13_234_1725_0, i_13_234_1726_0,
    i_13_234_1727_0, i_13_234_1731_0, i_13_234_1761_0, i_13_234_1780_0,
    i_13_234_1781_0, i_13_234_1846_0, i_13_234_1881_0, i_13_234_1884_0,
    i_13_234_1885_0, i_13_234_1886_0, i_13_234_1888_0, i_13_234_1889_0,
    i_13_234_1999_0, i_13_234_2009_0, i_13_234_2158_0, i_13_234_2380_0,
    i_13_234_2461_0, i_13_234_2462_0, i_13_234_2470_0, i_13_234_2629_0,
    i_13_234_2647_0, i_13_234_2650_0, i_13_234_2651_0, i_13_234_2714_0,
    i_13_234_2848_0, i_13_234_2849_0, i_13_234_2875_0, i_13_234_2878_0,
    i_13_234_2887_0, i_13_234_2916_0, i_13_234_2917_0, i_13_234_3004_0,
    i_13_234_3040_0, i_13_234_3041_0, i_13_234_3109_0, i_13_234_3145_0,
    i_13_234_3146_0, i_13_234_3293_0, i_13_234_3406_0, i_13_234_3429_0,
    i_13_234_3689_0, i_13_234_3707_0, i_13_234_3781_0, i_13_234_3794_0,
    i_13_234_3964_0, i_13_234_4083_0, i_13_234_4095_0, i_13_234_4096_0,
    i_13_234_4100_0, i_13_234_4153_0, i_13_234_4190_0, i_13_234_4253_0,
    i_13_234_4390_0, i_13_234_4414_0, i_13_234_4426_0, i_13_234_4437_0,
    i_13_234_4440_0, i_13_234_4513_0, i_13_234_4519_0, i_13_234_4526_0;
  output o_13_234_0_0;
  assign o_13_234_0_0 = ~((i_13_234_1498_0 & ((~i_13_234_1780_0 & ~i_13_234_1781_0 & ~i_13_234_2875_0 & ~i_13_234_2878_0) | (i_13_234_2887_0 & ~i_13_234_4253_0))) | (~i_13_234_1714_0 & ((~i_13_234_143_0 & ~i_13_234_280_0 & ~i_13_234_1222_0) | (~i_13_234_1277_0 & ~i_13_234_2849_0 & ~i_13_234_3145_0))) | (~i_13_234_1780_0 & ((~i_13_234_2461_0 & ~i_13_234_2848_0 & ~i_13_234_2849_0) | (~i_13_234_1999_0 & ~i_13_234_2714_0 & ~i_13_234_4253_0))) | (~i_13_234_2849_0 & ((~i_13_234_539_0 & ~i_13_234_620_0 & ~i_13_234_1715_0 & ~i_13_234_2878_0) | (~i_13_234_3040_0 & ~i_13_234_4190_0))) | (~i_13_234_3689_0 & ~i_13_234_4190_0 & i_13_234_4253_0));
endmodule



// Benchmark "kernel_13_235" written by ABC on Sun Jul 19 10:48:42 2020

module kernel_13_235 ( 
    i_13_235_67_0, i_13_235_68_0, i_13_235_70_0, i_13_235_97_0,
    i_13_235_173_0, i_13_235_233_0, i_13_235_234_0, i_13_235_311_0,
    i_13_235_319_0, i_13_235_349_0, i_13_235_389_0, i_13_235_412_0,
    i_13_235_444_0, i_13_235_534_0, i_13_235_538_0, i_13_235_539_0,
    i_13_235_643_0, i_13_235_644_0, i_13_235_646_0, i_13_235_682_0,
    i_13_235_797_0, i_13_235_841_0, i_13_235_898_0, i_13_235_930_0,
    i_13_235_932_0, i_13_235_938_0, i_13_235_1105_0, i_13_235_1120_0,
    i_13_235_1121_0, i_13_235_1222_0, i_13_235_1259_0, i_13_235_1274_0,
    i_13_235_1281_0, i_13_235_1390_0, i_13_235_1391_0, i_13_235_1400_0,
    i_13_235_1428_0, i_13_235_1461_0, i_13_235_1491_0, i_13_235_1511_0,
    i_13_235_1512_0, i_13_235_1552_0, i_13_235_1642_0, i_13_235_1733_0,
    i_13_235_1765_0, i_13_235_1795_0, i_13_235_1796_0, i_13_235_1798_0,
    i_13_235_1804_0, i_13_235_1867_0, i_13_235_1881_0, i_13_235_1886_0,
    i_13_235_1924_0, i_13_235_1945_0, i_13_235_1946_0, i_13_235_2017_0,
    i_13_235_2021_0, i_13_235_2032_0, i_13_235_2056_0, i_13_235_2142_0,
    i_13_235_2315_0, i_13_235_2461_0, i_13_235_2542_0, i_13_235_2594_0,
    i_13_235_2678_0, i_13_235_2847_0, i_13_235_2848_0, i_13_235_2849_0,
    i_13_235_2878_0, i_13_235_2884_0, i_13_235_2966_0, i_13_235_3040_0,
    i_13_235_3075_0, i_13_235_3101_0, i_13_235_3172_0, i_13_235_3176_0,
    i_13_235_3367_0, i_13_235_3523_0, i_13_235_3730_0, i_13_235_3736_0,
    i_13_235_3740_0, i_13_235_3757_0, i_13_235_3784_0, i_13_235_3889_0,
    i_13_235_3910_0, i_13_235_3928_0, i_13_235_3930_0, i_13_235_3931_0,
    i_13_235_4038_0, i_13_235_4186_0, i_13_235_4187_0, i_13_235_4189_0,
    i_13_235_4294_0, i_13_235_4297_0, i_13_235_4303_0, i_13_235_4351_0,
    i_13_235_4453_0, i_13_235_4595_0, i_13_235_4597_0, i_13_235_4606_0,
    o_13_235_0_0  );
  input  i_13_235_67_0, i_13_235_68_0, i_13_235_70_0, i_13_235_97_0,
    i_13_235_173_0, i_13_235_233_0, i_13_235_234_0, i_13_235_311_0,
    i_13_235_319_0, i_13_235_349_0, i_13_235_389_0, i_13_235_412_0,
    i_13_235_444_0, i_13_235_534_0, i_13_235_538_0, i_13_235_539_0,
    i_13_235_643_0, i_13_235_644_0, i_13_235_646_0, i_13_235_682_0,
    i_13_235_797_0, i_13_235_841_0, i_13_235_898_0, i_13_235_930_0,
    i_13_235_932_0, i_13_235_938_0, i_13_235_1105_0, i_13_235_1120_0,
    i_13_235_1121_0, i_13_235_1222_0, i_13_235_1259_0, i_13_235_1274_0,
    i_13_235_1281_0, i_13_235_1390_0, i_13_235_1391_0, i_13_235_1400_0,
    i_13_235_1428_0, i_13_235_1461_0, i_13_235_1491_0, i_13_235_1511_0,
    i_13_235_1512_0, i_13_235_1552_0, i_13_235_1642_0, i_13_235_1733_0,
    i_13_235_1765_0, i_13_235_1795_0, i_13_235_1796_0, i_13_235_1798_0,
    i_13_235_1804_0, i_13_235_1867_0, i_13_235_1881_0, i_13_235_1886_0,
    i_13_235_1924_0, i_13_235_1945_0, i_13_235_1946_0, i_13_235_2017_0,
    i_13_235_2021_0, i_13_235_2032_0, i_13_235_2056_0, i_13_235_2142_0,
    i_13_235_2315_0, i_13_235_2461_0, i_13_235_2542_0, i_13_235_2594_0,
    i_13_235_2678_0, i_13_235_2847_0, i_13_235_2848_0, i_13_235_2849_0,
    i_13_235_2878_0, i_13_235_2884_0, i_13_235_2966_0, i_13_235_3040_0,
    i_13_235_3075_0, i_13_235_3101_0, i_13_235_3172_0, i_13_235_3176_0,
    i_13_235_3367_0, i_13_235_3523_0, i_13_235_3730_0, i_13_235_3736_0,
    i_13_235_3740_0, i_13_235_3757_0, i_13_235_3784_0, i_13_235_3889_0,
    i_13_235_3910_0, i_13_235_3928_0, i_13_235_3930_0, i_13_235_3931_0,
    i_13_235_4038_0, i_13_235_4186_0, i_13_235_4187_0, i_13_235_4189_0,
    i_13_235_4294_0, i_13_235_4297_0, i_13_235_4303_0, i_13_235_4351_0,
    i_13_235_4453_0, i_13_235_4595_0, i_13_235_4597_0, i_13_235_4606_0;
  output o_13_235_0_0;
  assign o_13_235_0_0 = ~((~i_13_235_173_0 & (i_13_235_3736_0 | (~i_13_235_1222_0 & ~i_13_235_1796_0 & ~i_13_235_4186_0))) | (i_13_235_3784_0 & ((~i_13_235_2056_0 & ~i_13_235_3757_0) | (~i_13_235_319_0 & ~i_13_235_3176_0 & ~i_13_235_4303_0))) | (~i_13_235_1642_0 & ~i_13_235_1795_0) | (~i_13_235_1121_0 & ~i_13_235_1765_0 & i_13_235_1804_0) | (~i_13_235_444_0 & ~i_13_235_3523_0 & ~i_13_235_3740_0) | (~i_13_235_234_0 & ~i_13_235_898_0 & ~i_13_235_932_0 & ~i_13_235_2849_0 & ~i_13_235_3930_0 & ~i_13_235_4187_0));
endmodule



// Benchmark "kernel_13_236" written by ABC on Sun Jul 19 10:48:42 2020

module kernel_13_236 ( 
    i_13_236_76_0, i_13_236_77_0, i_13_236_79_0, i_13_236_94_0,
    i_13_236_116_0, i_13_236_251_0, i_13_236_329_0, i_13_236_431_0,
    i_13_236_450_0, i_13_236_494_0, i_13_236_518_0, i_13_236_571_0,
    i_13_236_604_0, i_13_236_605_0, i_13_236_619_0, i_13_236_658_0,
    i_13_236_670_0, i_13_236_697_0, i_13_236_698_0, i_13_236_700_0,
    i_13_236_845_0, i_13_236_928_0, i_13_236_940_0, i_13_236_1024_0,
    i_13_236_1078_0, i_13_236_1079_0, i_13_236_1081_0, i_13_236_1082_0,
    i_13_236_1213_0, i_13_236_1276_0, i_13_236_1277_0, i_13_236_1317_0,
    i_13_236_1318_0, i_13_236_1341_0, i_13_236_1408_0, i_13_236_1427_0,
    i_13_236_1429_0, i_13_236_1430_0, i_13_236_1444_0, i_13_236_1573_0,
    i_13_236_1629_0, i_13_236_1637_0, i_13_236_1711_0, i_13_236_1731_0,
    i_13_236_1736_0, i_13_236_1781_0, i_13_236_1888_0, i_13_236_2027_0,
    i_13_236_2029_0, i_13_236_2060_0, i_13_236_2104_0, i_13_236_2198_0,
    i_13_236_2209_0, i_13_236_2236_0, i_13_236_2448_0, i_13_236_2453_0,
    i_13_236_2455_0, i_13_236_2511_0, i_13_236_2617_0, i_13_236_2632_0,
    i_13_236_2710_0, i_13_236_2726_0, i_13_236_2764_0, i_13_236_2809_0,
    i_13_236_2821_0, i_13_236_2854_0, i_13_236_2887_0, i_13_236_2888_0,
    i_13_236_2959_0, i_13_236_2986_0, i_13_236_3061_0, i_13_236_3208_0,
    i_13_236_3343_0, i_13_236_3392_0, i_13_236_3419_0, i_13_236_3452_0,
    i_13_236_3454_0, i_13_236_3460_0, i_13_236_3464_0, i_13_236_3490_0,
    i_13_236_3536_0, i_13_236_3571_0, i_13_236_3572_0, i_13_236_3593_0,
    i_13_236_3601_0, i_13_236_3662_0, i_13_236_3688_0, i_13_236_3717_0,
    i_13_236_3847_0, i_13_236_3850_0, i_13_236_4009_0, i_13_236_4063_0,
    i_13_236_4087_0, i_13_236_4094_0, i_13_236_4252_0, i_13_236_4264_0,
    i_13_236_4267_0, i_13_236_4330_0, i_13_236_4365_0, i_13_236_4562_0,
    o_13_236_0_0  );
  input  i_13_236_76_0, i_13_236_77_0, i_13_236_79_0, i_13_236_94_0,
    i_13_236_116_0, i_13_236_251_0, i_13_236_329_0, i_13_236_431_0,
    i_13_236_450_0, i_13_236_494_0, i_13_236_518_0, i_13_236_571_0,
    i_13_236_604_0, i_13_236_605_0, i_13_236_619_0, i_13_236_658_0,
    i_13_236_670_0, i_13_236_697_0, i_13_236_698_0, i_13_236_700_0,
    i_13_236_845_0, i_13_236_928_0, i_13_236_940_0, i_13_236_1024_0,
    i_13_236_1078_0, i_13_236_1079_0, i_13_236_1081_0, i_13_236_1082_0,
    i_13_236_1213_0, i_13_236_1276_0, i_13_236_1277_0, i_13_236_1317_0,
    i_13_236_1318_0, i_13_236_1341_0, i_13_236_1408_0, i_13_236_1427_0,
    i_13_236_1429_0, i_13_236_1430_0, i_13_236_1444_0, i_13_236_1573_0,
    i_13_236_1629_0, i_13_236_1637_0, i_13_236_1711_0, i_13_236_1731_0,
    i_13_236_1736_0, i_13_236_1781_0, i_13_236_1888_0, i_13_236_2027_0,
    i_13_236_2029_0, i_13_236_2060_0, i_13_236_2104_0, i_13_236_2198_0,
    i_13_236_2209_0, i_13_236_2236_0, i_13_236_2448_0, i_13_236_2453_0,
    i_13_236_2455_0, i_13_236_2511_0, i_13_236_2617_0, i_13_236_2632_0,
    i_13_236_2710_0, i_13_236_2726_0, i_13_236_2764_0, i_13_236_2809_0,
    i_13_236_2821_0, i_13_236_2854_0, i_13_236_2887_0, i_13_236_2888_0,
    i_13_236_2959_0, i_13_236_2986_0, i_13_236_3061_0, i_13_236_3208_0,
    i_13_236_3343_0, i_13_236_3392_0, i_13_236_3419_0, i_13_236_3452_0,
    i_13_236_3454_0, i_13_236_3460_0, i_13_236_3464_0, i_13_236_3490_0,
    i_13_236_3536_0, i_13_236_3571_0, i_13_236_3572_0, i_13_236_3593_0,
    i_13_236_3601_0, i_13_236_3662_0, i_13_236_3688_0, i_13_236_3717_0,
    i_13_236_3847_0, i_13_236_3850_0, i_13_236_4009_0, i_13_236_4063_0,
    i_13_236_4087_0, i_13_236_4094_0, i_13_236_4252_0, i_13_236_4264_0,
    i_13_236_4267_0, i_13_236_4330_0, i_13_236_4365_0, i_13_236_4562_0;
  output o_13_236_0_0;
  assign o_13_236_0_0 = ~((~i_13_236_2453_0 & (~i_13_236_1078_0 | (~i_13_236_1024_0 & i_13_236_3847_0))) | (~i_13_236_2726_0 & (i_13_236_1408_0 | (~i_13_236_1888_0 & ~i_13_236_4009_0))) | (~i_13_236_700_0 & ~i_13_236_3464_0) | (~i_13_236_1430_0 & i_13_236_3343_0 & ~i_13_236_3572_0) | (~i_13_236_2887_0 & i_13_236_4009_0));
endmodule



// Benchmark "kernel_13_237" written by ABC on Sun Jul 19 10:48:43 2020

module kernel_13_237 ( 
    i_13_237_97_0, i_13_237_106_0, i_13_237_125_0, i_13_237_134_0,
    i_13_237_233_0, i_13_237_358_0, i_13_237_376_0, i_13_237_409_0,
    i_13_237_512_0, i_13_237_529_0, i_13_237_530_0, i_13_237_573_0,
    i_13_237_574_0, i_13_237_575_0, i_13_237_607_0, i_13_237_718_0,
    i_13_237_799_0, i_13_237_800_0, i_13_237_845_0, i_13_237_1101_0,
    i_13_237_1304_0, i_13_237_1322_0, i_13_237_1410_0, i_13_237_1447_0,
    i_13_237_1492_0, i_13_237_1493_0, i_13_237_1501_0, i_13_237_1502_0,
    i_13_237_1511_0, i_13_237_1538_0, i_13_237_1543_0, i_13_237_1555_0,
    i_13_237_1556_0, i_13_237_1642_0, i_13_237_1643_0, i_13_237_1711_0,
    i_13_237_1744_0, i_13_237_1760_0, i_13_237_1796_0, i_13_237_1840_0,
    i_13_237_1933_0, i_13_237_1951_0, i_13_237_1990_0, i_13_237_1991_0,
    i_13_237_2015_0, i_13_237_2104_0, i_13_237_2239_0, i_13_237_2240_0,
    i_13_237_2246_0, i_13_237_2266_0, i_13_237_2318_0, i_13_237_2362_0,
    i_13_237_2428_0, i_13_237_2429_0, i_13_237_2458_0, i_13_237_2483_0,
    i_13_237_2536_0, i_13_237_2825_0, i_13_237_2906_0, i_13_237_2935_0,
    i_13_237_2936_0, i_13_237_2938_0, i_13_237_2947_0, i_13_237_2971_0,
    i_13_237_2983_0, i_13_237_3028_0, i_13_237_3065_0, i_13_237_3100_0,
    i_13_237_3117_0, i_13_237_3127_0, i_13_237_3207_0, i_13_237_3208_0,
    i_13_237_3244_0, i_13_237_3245_0, i_13_237_3425_0, i_13_237_3427_0,
    i_13_237_3428_0, i_13_237_3455_0, i_13_237_3478_0, i_13_237_3544_0,
    i_13_237_3722_0, i_13_237_3788_0, i_13_237_3794_0, i_13_237_3806_0,
    i_13_237_3859_0, i_13_237_3860_0, i_13_237_3914_0, i_13_237_3968_0,
    i_13_237_3985_0, i_13_237_4012_0, i_13_237_4013_0, i_13_237_4120_0,
    i_13_237_4219_0, i_13_237_4308_0, i_13_237_4313_0, i_13_237_4433_0,
    i_13_237_4444_0, i_13_237_4541_0, i_13_237_4567_0, i_13_237_4588_0,
    o_13_237_0_0  );
  input  i_13_237_97_0, i_13_237_106_0, i_13_237_125_0, i_13_237_134_0,
    i_13_237_233_0, i_13_237_358_0, i_13_237_376_0, i_13_237_409_0,
    i_13_237_512_0, i_13_237_529_0, i_13_237_530_0, i_13_237_573_0,
    i_13_237_574_0, i_13_237_575_0, i_13_237_607_0, i_13_237_718_0,
    i_13_237_799_0, i_13_237_800_0, i_13_237_845_0, i_13_237_1101_0,
    i_13_237_1304_0, i_13_237_1322_0, i_13_237_1410_0, i_13_237_1447_0,
    i_13_237_1492_0, i_13_237_1493_0, i_13_237_1501_0, i_13_237_1502_0,
    i_13_237_1511_0, i_13_237_1538_0, i_13_237_1543_0, i_13_237_1555_0,
    i_13_237_1556_0, i_13_237_1642_0, i_13_237_1643_0, i_13_237_1711_0,
    i_13_237_1744_0, i_13_237_1760_0, i_13_237_1796_0, i_13_237_1840_0,
    i_13_237_1933_0, i_13_237_1951_0, i_13_237_1990_0, i_13_237_1991_0,
    i_13_237_2015_0, i_13_237_2104_0, i_13_237_2239_0, i_13_237_2240_0,
    i_13_237_2246_0, i_13_237_2266_0, i_13_237_2318_0, i_13_237_2362_0,
    i_13_237_2428_0, i_13_237_2429_0, i_13_237_2458_0, i_13_237_2483_0,
    i_13_237_2536_0, i_13_237_2825_0, i_13_237_2906_0, i_13_237_2935_0,
    i_13_237_2936_0, i_13_237_2938_0, i_13_237_2947_0, i_13_237_2971_0,
    i_13_237_2983_0, i_13_237_3028_0, i_13_237_3065_0, i_13_237_3100_0,
    i_13_237_3117_0, i_13_237_3127_0, i_13_237_3207_0, i_13_237_3208_0,
    i_13_237_3244_0, i_13_237_3245_0, i_13_237_3425_0, i_13_237_3427_0,
    i_13_237_3428_0, i_13_237_3455_0, i_13_237_3478_0, i_13_237_3544_0,
    i_13_237_3722_0, i_13_237_3788_0, i_13_237_3794_0, i_13_237_3806_0,
    i_13_237_3859_0, i_13_237_3860_0, i_13_237_3914_0, i_13_237_3968_0,
    i_13_237_3985_0, i_13_237_4012_0, i_13_237_4013_0, i_13_237_4120_0,
    i_13_237_4219_0, i_13_237_4308_0, i_13_237_4313_0, i_13_237_4433_0,
    i_13_237_4444_0, i_13_237_4541_0, i_13_237_4567_0, i_13_237_4588_0;
  output o_13_237_0_0;
  assign o_13_237_0_0 = ~((~i_13_237_97_0 & i_13_237_4567_0) | (~i_13_237_575_0 & ~i_13_237_4433_0 & ~i_13_237_4567_0) | (~i_13_237_1556_0 & ~i_13_237_2536_0 & ~i_13_237_4013_0));
endmodule



// Benchmark "kernel_13_238" written by ABC on Sun Jul 19 10:48:44 2020

module kernel_13_238 ( 
    i_13_238_49_0, i_13_238_93_0, i_13_238_117_0, i_13_238_180_0,
    i_13_238_181_0, i_13_238_183_0, i_13_238_184_0, i_13_238_190_0,
    i_13_238_193_0, i_13_238_381_0, i_13_238_382_0, i_13_238_489_0,
    i_13_238_527_0, i_13_238_531_0, i_13_238_567_0, i_13_238_589_0,
    i_13_238_621_0, i_13_238_624_0, i_13_238_689_0, i_13_238_712_0,
    i_13_238_713_0, i_13_238_715_0, i_13_238_858_0, i_13_238_948_0,
    i_13_238_1099_0, i_13_238_1116_0, i_13_238_1117_0, i_13_238_1146_0,
    i_13_238_1219_0, i_13_238_1225_0, i_13_238_1251_0, i_13_238_1254_0,
    i_13_238_1255_0, i_13_238_1280_0, i_13_238_1387_0, i_13_238_1404_0,
    i_13_238_1407_0, i_13_238_1408_0, i_13_238_1488_0, i_13_238_1489_0,
    i_13_238_1512_0, i_13_238_1513_0, i_13_238_1677_0, i_13_238_1680_0,
    i_13_238_1760_0, i_13_238_1765_0, i_13_238_1786_0, i_13_238_1792_0,
    i_13_238_1801_0, i_13_238_1857_0, i_13_238_1862_0, i_13_238_1991_0,
    i_13_238_2002_0, i_13_238_2123_0, i_13_238_2242_0, i_13_238_2263_0,
    i_13_238_2281_0, i_13_238_2314_0, i_13_238_2533_0, i_13_238_2690_0,
    i_13_238_2836_0, i_13_238_2848_0, i_13_238_2856_0, i_13_238_2857_0,
    i_13_238_2908_0, i_13_238_2967_0, i_13_238_3025_0, i_13_238_3064_0,
    i_13_238_3126_0, i_13_238_3148_0, i_13_238_3153_0, i_13_238_3260_0,
    i_13_238_3262_0, i_13_238_3348_0, i_13_238_3352_0, i_13_238_3427_0,
    i_13_238_3456_0, i_13_238_3466_0, i_13_238_3478_0, i_13_238_3486_0,
    i_13_238_3489_0, i_13_238_3612_0, i_13_238_3638_0, i_13_238_3685_0,
    i_13_238_3699_0, i_13_238_3753_0, i_13_238_3754_0, i_13_238_3756_0,
    i_13_238_3757_0, i_13_238_3762_0, i_13_238_3874_0, i_13_238_3890_0,
    i_13_238_3978_0, i_13_238_4045_0, i_13_238_4261_0, i_13_238_4404_0,
    i_13_238_4509_0, i_13_238_4510_0, i_13_238_4538_0, i_13_238_4563_0,
    o_13_238_0_0  );
  input  i_13_238_49_0, i_13_238_93_0, i_13_238_117_0, i_13_238_180_0,
    i_13_238_181_0, i_13_238_183_0, i_13_238_184_0, i_13_238_190_0,
    i_13_238_193_0, i_13_238_381_0, i_13_238_382_0, i_13_238_489_0,
    i_13_238_527_0, i_13_238_531_0, i_13_238_567_0, i_13_238_589_0,
    i_13_238_621_0, i_13_238_624_0, i_13_238_689_0, i_13_238_712_0,
    i_13_238_713_0, i_13_238_715_0, i_13_238_858_0, i_13_238_948_0,
    i_13_238_1099_0, i_13_238_1116_0, i_13_238_1117_0, i_13_238_1146_0,
    i_13_238_1219_0, i_13_238_1225_0, i_13_238_1251_0, i_13_238_1254_0,
    i_13_238_1255_0, i_13_238_1280_0, i_13_238_1387_0, i_13_238_1404_0,
    i_13_238_1407_0, i_13_238_1408_0, i_13_238_1488_0, i_13_238_1489_0,
    i_13_238_1512_0, i_13_238_1513_0, i_13_238_1677_0, i_13_238_1680_0,
    i_13_238_1760_0, i_13_238_1765_0, i_13_238_1786_0, i_13_238_1792_0,
    i_13_238_1801_0, i_13_238_1857_0, i_13_238_1862_0, i_13_238_1991_0,
    i_13_238_2002_0, i_13_238_2123_0, i_13_238_2242_0, i_13_238_2263_0,
    i_13_238_2281_0, i_13_238_2314_0, i_13_238_2533_0, i_13_238_2690_0,
    i_13_238_2836_0, i_13_238_2848_0, i_13_238_2856_0, i_13_238_2857_0,
    i_13_238_2908_0, i_13_238_2967_0, i_13_238_3025_0, i_13_238_3064_0,
    i_13_238_3126_0, i_13_238_3148_0, i_13_238_3153_0, i_13_238_3260_0,
    i_13_238_3262_0, i_13_238_3348_0, i_13_238_3352_0, i_13_238_3427_0,
    i_13_238_3456_0, i_13_238_3466_0, i_13_238_3478_0, i_13_238_3486_0,
    i_13_238_3489_0, i_13_238_3612_0, i_13_238_3638_0, i_13_238_3685_0,
    i_13_238_3699_0, i_13_238_3753_0, i_13_238_3754_0, i_13_238_3756_0,
    i_13_238_3757_0, i_13_238_3762_0, i_13_238_3874_0, i_13_238_3890_0,
    i_13_238_3978_0, i_13_238_4045_0, i_13_238_4261_0, i_13_238_4404_0,
    i_13_238_4509_0, i_13_238_4510_0, i_13_238_4538_0, i_13_238_4563_0;
  output o_13_238_0_0;
  assign o_13_238_0_0 = ~((~i_13_238_1792_0 & ((~i_13_238_1857_0 & ~i_13_238_2242_0 & ~i_13_238_3753_0) | (~i_13_238_1488_0 & ~i_13_238_1765_0 & ~i_13_238_3762_0))) | (~i_13_238_1677_0 & ~i_13_238_1801_0) | (~i_13_238_3612_0 & ~i_13_238_3874_0) | (~i_13_238_1404_0 & ~i_13_238_1408_0 & ~i_13_238_3978_0) | (i_13_238_93_0 & ~i_13_238_190_0 & ~i_13_238_4509_0));
endmodule



// Benchmark "kernel_13_239" written by ABC on Sun Jul 19 10:48:45 2020

module kernel_13_239 ( 
    i_13_239_24_0, i_13_239_44_0, i_13_239_66_0, i_13_239_112_0,
    i_13_239_115_0, i_13_239_183_0, i_13_239_210_0, i_13_239_268_0,
    i_13_239_357_0, i_13_239_391_0, i_13_239_465_0, i_13_239_466_0,
    i_13_239_527_0, i_13_239_529_0, i_13_239_552_0, i_13_239_591_0,
    i_13_239_744_0, i_13_239_762_0, i_13_239_795_0, i_13_239_831_0,
    i_13_239_859_0, i_13_239_1083_0, i_13_239_1084_0, i_13_239_1131_0,
    i_13_239_1302_0, i_13_239_1303_0, i_13_239_1321_0, i_13_239_1419_0,
    i_13_239_1434_0, i_13_239_1474_0, i_13_239_1565_0, i_13_239_1597_0,
    i_13_239_1605_0, i_13_239_1607_0, i_13_239_1627_0, i_13_239_1677_0,
    i_13_239_1753_0, i_13_239_1806_0, i_13_239_1842_0, i_13_239_1843_0,
    i_13_239_1849_0, i_13_239_1914_0, i_13_239_1960_0, i_13_239_2029_0,
    i_13_239_2139_0, i_13_239_2145_0, i_13_239_2202_0, i_13_239_2203_0,
    i_13_239_2239_0, i_13_239_2284_0, i_13_239_2397_0, i_13_239_2401_0,
    i_13_239_2472_0, i_13_239_2506_0, i_13_239_2544_0, i_13_239_2545_0,
    i_13_239_2553_0, i_13_239_2578_0, i_13_239_2699_0, i_13_239_2704_0,
    i_13_239_2759_0, i_13_239_2762_0, i_13_239_2824_0, i_13_239_3003_0,
    i_13_239_3075_0, i_13_239_3092_0, i_13_239_3166_0, i_13_239_3243_0,
    i_13_239_3326_0, i_13_239_3345_0, i_13_239_3346_0, i_13_239_3373_0,
    i_13_239_3391_0, i_13_239_3477_0, i_13_239_3481_0, i_13_239_3579_0,
    i_13_239_3597_0, i_13_239_3633_0, i_13_239_3669_0, i_13_239_3724_0,
    i_13_239_3768_0, i_13_239_3805_0, i_13_239_3823_0, i_13_239_3859_0,
    i_13_239_3860_0, i_13_239_3894_0, i_13_239_3939_0, i_13_239_4038_0,
    i_13_239_4099_0, i_13_239_4164_0, i_13_239_4254_0, i_13_239_4264_0,
    i_13_239_4265_0, i_13_239_4272_0, i_13_239_4309_0, i_13_239_4315_0,
    i_13_239_4380_0, i_13_239_4381_0, i_13_239_4452_0, i_13_239_4453_0,
    o_13_239_0_0  );
  input  i_13_239_24_0, i_13_239_44_0, i_13_239_66_0, i_13_239_112_0,
    i_13_239_115_0, i_13_239_183_0, i_13_239_210_0, i_13_239_268_0,
    i_13_239_357_0, i_13_239_391_0, i_13_239_465_0, i_13_239_466_0,
    i_13_239_527_0, i_13_239_529_0, i_13_239_552_0, i_13_239_591_0,
    i_13_239_744_0, i_13_239_762_0, i_13_239_795_0, i_13_239_831_0,
    i_13_239_859_0, i_13_239_1083_0, i_13_239_1084_0, i_13_239_1131_0,
    i_13_239_1302_0, i_13_239_1303_0, i_13_239_1321_0, i_13_239_1419_0,
    i_13_239_1434_0, i_13_239_1474_0, i_13_239_1565_0, i_13_239_1597_0,
    i_13_239_1605_0, i_13_239_1607_0, i_13_239_1627_0, i_13_239_1677_0,
    i_13_239_1753_0, i_13_239_1806_0, i_13_239_1842_0, i_13_239_1843_0,
    i_13_239_1849_0, i_13_239_1914_0, i_13_239_1960_0, i_13_239_2029_0,
    i_13_239_2139_0, i_13_239_2145_0, i_13_239_2202_0, i_13_239_2203_0,
    i_13_239_2239_0, i_13_239_2284_0, i_13_239_2397_0, i_13_239_2401_0,
    i_13_239_2472_0, i_13_239_2506_0, i_13_239_2544_0, i_13_239_2545_0,
    i_13_239_2553_0, i_13_239_2578_0, i_13_239_2699_0, i_13_239_2704_0,
    i_13_239_2759_0, i_13_239_2762_0, i_13_239_2824_0, i_13_239_3003_0,
    i_13_239_3075_0, i_13_239_3092_0, i_13_239_3166_0, i_13_239_3243_0,
    i_13_239_3326_0, i_13_239_3345_0, i_13_239_3346_0, i_13_239_3373_0,
    i_13_239_3391_0, i_13_239_3477_0, i_13_239_3481_0, i_13_239_3579_0,
    i_13_239_3597_0, i_13_239_3633_0, i_13_239_3669_0, i_13_239_3724_0,
    i_13_239_3768_0, i_13_239_3805_0, i_13_239_3823_0, i_13_239_3859_0,
    i_13_239_3860_0, i_13_239_3894_0, i_13_239_3939_0, i_13_239_4038_0,
    i_13_239_4099_0, i_13_239_4164_0, i_13_239_4254_0, i_13_239_4264_0,
    i_13_239_4265_0, i_13_239_4272_0, i_13_239_4309_0, i_13_239_4315_0,
    i_13_239_4380_0, i_13_239_4381_0, i_13_239_4452_0, i_13_239_4453_0;
  output o_13_239_0_0;
  assign o_13_239_0_0 = ~((~i_13_239_1605_0 & ((~i_13_239_1753_0 & i_13_239_4164_0) | (~i_13_239_2139_0 & ~i_13_239_3859_0 & ~i_13_239_4453_0))) | (i_13_239_2762_0 & ~i_13_239_3346_0) | (~i_13_239_762_0 & ~i_13_239_2139_0 & ~i_13_239_3391_0) | (i_13_239_3166_0 & ~i_13_239_4038_0 & ~i_13_239_4309_0 & ~i_13_239_4380_0));
endmodule



// Benchmark "kernel_13_240" written by ABC on Sun Jul 19 10:48:45 2020

module kernel_13_240 ( 
    i_13_240_65_0, i_13_240_131_0, i_13_240_163_0, i_13_240_252_0,
    i_13_240_256_0, i_13_240_266_0, i_13_240_269_0, i_13_240_272_0,
    i_13_240_308_0, i_13_240_340_0, i_13_240_354_0, i_13_240_379_0,
    i_13_240_380_0, i_13_240_458_0, i_13_240_463_0, i_13_240_466_0,
    i_13_240_467_0, i_13_240_475_0, i_13_240_535_0, i_13_240_592_0,
    i_13_240_684_0, i_13_240_821_0, i_13_240_829_0, i_13_240_895_0,
    i_13_240_1116_0, i_13_240_1120_0, i_13_240_1121_0, i_13_240_1307_0,
    i_13_240_1397_0, i_13_240_1444_0, i_13_240_1448_0, i_13_240_1467_0,
    i_13_240_1480_0, i_13_240_1496_0, i_13_240_1553_0, i_13_240_1594_0,
    i_13_240_1595_0, i_13_240_1697_0, i_13_240_1710_0, i_13_240_1723_0,
    i_13_240_1802_0, i_13_240_1844_0, i_13_240_1846_0, i_13_240_1847_0,
    i_13_240_1885_0, i_13_240_1908_0, i_13_240_1927_0, i_13_240_1928_0,
    i_13_240_1958_0, i_13_240_1989_0, i_13_240_1991_0, i_13_240_2101_0,
    i_13_240_2108_0, i_13_240_2261_0, i_13_240_2297_0, i_13_240_2366_0,
    i_13_240_2650_0, i_13_240_2677_0, i_13_240_2848_0, i_13_240_2849_0,
    i_13_240_2871_0, i_13_240_2935_0, i_13_240_2936_0, i_13_240_3035_0,
    i_13_240_3050_0, i_13_240_3167_0, i_13_240_3232_0, i_13_240_3241_0,
    i_13_240_3242_0, i_13_240_3415_0, i_13_240_3447_0, i_13_240_3519_0,
    i_13_240_3523_0, i_13_240_3569_0, i_13_240_3597_0, i_13_240_3598_0,
    i_13_240_3667_0, i_13_240_3730_0, i_13_240_3818_0, i_13_240_3857_0,
    i_13_240_3859_0, i_13_240_4017_0, i_13_240_4052_0, i_13_240_4060_0,
    i_13_240_4061_0, i_13_240_4063_0, i_13_240_4088_0, i_13_240_4165_0,
    i_13_240_4187_0, i_13_240_4189_0, i_13_240_4204_0, i_13_240_4205_0,
    i_13_240_4214_0, i_13_240_4267_0, i_13_240_4268_0, i_13_240_4313_0,
    i_13_240_4413_0, i_13_240_4430_0, i_13_240_4530_0, i_13_240_4562_0,
    o_13_240_0_0  );
  input  i_13_240_65_0, i_13_240_131_0, i_13_240_163_0, i_13_240_252_0,
    i_13_240_256_0, i_13_240_266_0, i_13_240_269_0, i_13_240_272_0,
    i_13_240_308_0, i_13_240_340_0, i_13_240_354_0, i_13_240_379_0,
    i_13_240_380_0, i_13_240_458_0, i_13_240_463_0, i_13_240_466_0,
    i_13_240_467_0, i_13_240_475_0, i_13_240_535_0, i_13_240_592_0,
    i_13_240_684_0, i_13_240_821_0, i_13_240_829_0, i_13_240_895_0,
    i_13_240_1116_0, i_13_240_1120_0, i_13_240_1121_0, i_13_240_1307_0,
    i_13_240_1397_0, i_13_240_1444_0, i_13_240_1448_0, i_13_240_1467_0,
    i_13_240_1480_0, i_13_240_1496_0, i_13_240_1553_0, i_13_240_1594_0,
    i_13_240_1595_0, i_13_240_1697_0, i_13_240_1710_0, i_13_240_1723_0,
    i_13_240_1802_0, i_13_240_1844_0, i_13_240_1846_0, i_13_240_1847_0,
    i_13_240_1885_0, i_13_240_1908_0, i_13_240_1927_0, i_13_240_1928_0,
    i_13_240_1958_0, i_13_240_1989_0, i_13_240_1991_0, i_13_240_2101_0,
    i_13_240_2108_0, i_13_240_2261_0, i_13_240_2297_0, i_13_240_2366_0,
    i_13_240_2650_0, i_13_240_2677_0, i_13_240_2848_0, i_13_240_2849_0,
    i_13_240_2871_0, i_13_240_2935_0, i_13_240_2936_0, i_13_240_3035_0,
    i_13_240_3050_0, i_13_240_3167_0, i_13_240_3232_0, i_13_240_3241_0,
    i_13_240_3242_0, i_13_240_3415_0, i_13_240_3447_0, i_13_240_3519_0,
    i_13_240_3523_0, i_13_240_3569_0, i_13_240_3597_0, i_13_240_3598_0,
    i_13_240_3667_0, i_13_240_3730_0, i_13_240_3818_0, i_13_240_3857_0,
    i_13_240_3859_0, i_13_240_4017_0, i_13_240_4052_0, i_13_240_4060_0,
    i_13_240_4061_0, i_13_240_4063_0, i_13_240_4088_0, i_13_240_4165_0,
    i_13_240_4187_0, i_13_240_4189_0, i_13_240_4204_0, i_13_240_4205_0,
    i_13_240_4214_0, i_13_240_4267_0, i_13_240_4268_0, i_13_240_4313_0,
    i_13_240_4413_0, i_13_240_4430_0, i_13_240_4530_0, i_13_240_4562_0;
  output o_13_240_0_0;
  assign o_13_240_0_0 = ~((~i_13_240_829_0 & ~i_13_240_4088_0) | (~i_13_240_3730_0 & ~i_13_240_4061_0) | (~i_13_240_1595_0 & ~i_13_240_1802_0 & ~i_13_240_4063_0));
endmodule



// Benchmark "kernel_13_241" written by ABC on Sun Jul 19 10:48:46 2020

module kernel_13_241 ( 
    i_13_241_69_0, i_13_241_101_0, i_13_241_230_0, i_13_241_326_0,
    i_13_241_336_0, i_13_241_379_0, i_13_241_505_0, i_13_241_573_0,
    i_13_241_578_0, i_13_241_623_0, i_13_241_641_0, i_13_241_690_0,
    i_13_241_717_0, i_13_241_780_0, i_13_241_1063_0, i_13_241_1064_0,
    i_13_241_1297_0, i_13_241_1298_0, i_13_241_1342_0, i_13_241_1410_0,
    i_13_241_1499_0, i_13_241_1529_0, i_13_241_1609_0, i_13_241_1627_0,
    i_13_241_1635_0, i_13_241_1712_0, i_13_241_1723_0, i_13_241_1777_0,
    i_13_241_1778_0, i_13_241_1801_0, i_13_241_1802_0, i_13_241_1810_0,
    i_13_241_1900_0, i_13_241_1906_0, i_13_241_1939_0, i_13_241_1990_0,
    i_13_241_1991_0, i_13_241_1993_0, i_13_241_2003_0, i_13_241_2012_0,
    i_13_241_2107_0, i_13_241_2134_0, i_13_241_2135_0, i_13_241_2209_0,
    i_13_241_2260_0, i_13_241_2261_0, i_13_241_2302_0, i_13_241_2309_0,
    i_13_241_2341_0, i_13_241_2359_0, i_13_241_2396_0, i_13_241_2404_0,
    i_13_241_2512_0, i_13_241_2522_0, i_13_241_2576_0, i_13_241_2614_0,
    i_13_241_2648_0, i_13_241_2746_0, i_13_241_2859_0, i_13_241_2935_0,
    i_13_241_2936_0, i_13_241_2939_0, i_13_241_2980_0, i_13_241_3012_0,
    i_13_241_3037_0, i_13_241_3143_0, i_13_241_3213_0, i_13_241_3286_0,
    i_13_241_3287_0, i_13_241_3340_0, i_13_241_3385_0, i_13_241_3386_0,
    i_13_241_3416_0, i_13_241_3421_0, i_13_241_3466_0, i_13_241_3476_0,
    i_13_241_3532_0, i_13_241_3642_0, i_13_241_3665_0, i_13_241_3729_0,
    i_13_241_3739_0, i_13_241_3747_0, i_13_241_3791_0, i_13_241_3876_0,
    i_13_241_4009_0, i_13_241_4011_0, i_13_241_4012_0, i_13_241_4015_0,
    i_13_241_4043_0, i_13_241_4055_0, i_13_241_4209_0, i_13_241_4230_0,
    i_13_241_4231_0, i_13_241_4232_0, i_13_241_4393_0, i_13_241_4398_0,
    i_13_241_4412_0, i_13_241_4531_0, i_13_241_4533_0, i_13_241_4587_0,
    o_13_241_0_0  );
  input  i_13_241_69_0, i_13_241_101_0, i_13_241_230_0, i_13_241_326_0,
    i_13_241_336_0, i_13_241_379_0, i_13_241_505_0, i_13_241_573_0,
    i_13_241_578_0, i_13_241_623_0, i_13_241_641_0, i_13_241_690_0,
    i_13_241_717_0, i_13_241_780_0, i_13_241_1063_0, i_13_241_1064_0,
    i_13_241_1297_0, i_13_241_1298_0, i_13_241_1342_0, i_13_241_1410_0,
    i_13_241_1499_0, i_13_241_1529_0, i_13_241_1609_0, i_13_241_1627_0,
    i_13_241_1635_0, i_13_241_1712_0, i_13_241_1723_0, i_13_241_1777_0,
    i_13_241_1778_0, i_13_241_1801_0, i_13_241_1802_0, i_13_241_1810_0,
    i_13_241_1900_0, i_13_241_1906_0, i_13_241_1939_0, i_13_241_1990_0,
    i_13_241_1991_0, i_13_241_1993_0, i_13_241_2003_0, i_13_241_2012_0,
    i_13_241_2107_0, i_13_241_2134_0, i_13_241_2135_0, i_13_241_2209_0,
    i_13_241_2260_0, i_13_241_2261_0, i_13_241_2302_0, i_13_241_2309_0,
    i_13_241_2341_0, i_13_241_2359_0, i_13_241_2396_0, i_13_241_2404_0,
    i_13_241_2512_0, i_13_241_2522_0, i_13_241_2576_0, i_13_241_2614_0,
    i_13_241_2648_0, i_13_241_2746_0, i_13_241_2859_0, i_13_241_2935_0,
    i_13_241_2936_0, i_13_241_2939_0, i_13_241_2980_0, i_13_241_3012_0,
    i_13_241_3037_0, i_13_241_3143_0, i_13_241_3213_0, i_13_241_3286_0,
    i_13_241_3287_0, i_13_241_3340_0, i_13_241_3385_0, i_13_241_3386_0,
    i_13_241_3416_0, i_13_241_3421_0, i_13_241_3466_0, i_13_241_3476_0,
    i_13_241_3532_0, i_13_241_3642_0, i_13_241_3665_0, i_13_241_3729_0,
    i_13_241_3739_0, i_13_241_3747_0, i_13_241_3791_0, i_13_241_3876_0,
    i_13_241_4009_0, i_13_241_4011_0, i_13_241_4012_0, i_13_241_4015_0,
    i_13_241_4043_0, i_13_241_4055_0, i_13_241_4209_0, i_13_241_4230_0,
    i_13_241_4231_0, i_13_241_4232_0, i_13_241_4393_0, i_13_241_4398_0,
    i_13_241_4412_0, i_13_241_4531_0, i_13_241_4533_0, i_13_241_4587_0;
  output o_13_241_0_0;
  assign o_13_241_0_0 = ~((~i_13_241_1298_0 & ~i_13_241_3037_0) | (~i_13_241_1063_0 & ~i_13_241_2135_0 & ~i_13_241_3386_0 & ~i_13_241_4412_0));
endmodule



// Benchmark "kernel_13_242" written by ABC on Sun Jul 19 10:48:47 2020

module kernel_13_242 ( 
    i_13_242_94_0, i_13_242_121_0, i_13_242_229_0, i_13_242_230_0,
    i_13_242_232_0, i_13_242_518_0, i_13_242_520_0, i_13_242_521_0,
    i_13_242_535_0, i_13_242_645_0, i_13_242_661_0, i_13_242_739_0,
    i_13_242_756_0, i_13_242_820_0, i_13_242_850_0, i_13_242_851_0,
    i_13_242_870_0, i_13_242_938_0, i_13_242_1072_0, i_13_242_1073_0,
    i_13_242_1075_0, i_13_242_1201_0, i_13_242_1219_0, i_13_242_1262_0,
    i_13_242_1423_0, i_13_242_1424_0, i_13_242_1549_0, i_13_242_1550_0,
    i_13_242_1624_0, i_13_242_1630_0, i_13_242_1723_0, i_13_242_1758_0,
    i_13_242_1774_0, i_13_242_1787_0, i_13_242_1858_0, i_13_242_1939_0,
    i_13_242_1970_0, i_13_242_2027_0, i_13_242_2029_0, i_13_242_2033_0,
    i_13_242_2201_0, i_13_242_2209_0, i_13_242_2425_0, i_13_242_2451_0,
    i_13_242_2452_0, i_13_242_2454_0, i_13_242_2455_0, i_13_242_2558_0,
    i_13_242_2567_0, i_13_242_2612_0, i_13_242_2693_0, i_13_242_2764_0,
    i_13_242_2848_0, i_13_242_2850_0, i_13_242_3010_0, i_13_242_3011_0,
    i_13_242_3014_0, i_13_242_3037_0, i_13_242_3040_0, i_13_242_3143_0,
    i_13_242_3163_0, i_13_242_3217_0, i_13_242_3251_0, i_13_242_3272_0,
    i_13_242_3424_0, i_13_242_3442_0, i_13_242_3467_0, i_13_242_3472_0,
    i_13_242_3473_0, i_13_242_3485_0, i_13_242_3487_0, i_13_242_3488_0,
    i_13_242_3539_0, i_13_242_3541_0, i_13_242_3575_0, i_13_242_3731_0,
    i_13_242_3784_0, i_13_242_3853_0, i_13_242_3856_0, i_13_242_3863_0,
    i_13_242_3866_0, i_13_242_3893_0, i_13_242_3991_0, i_13_242_4038_0,
    i_13_242_4210_0, i_13_242_4216_0, i_13_242_4252_0, i_13_242_4253_0,
    i_13_242_4261_0, i_13_242_4262_0, i_13_242_4264_0, i_13_242_4265_0,
    i_13_242_4355_0, i_13_242_4370_0, i_13_242_4372_0, i_13_242_4379_0,
    i_13_242_4380_0, i_13_242_4511_0, i_13_242_4540_0, i_13_242_4558_0,
    o_13_242_0_0  );
  input  i_13_242_94_0, i_13_242_121_0, i_13_242_229_0, i_13_242_230_0,
    i_13_242_232_0, i_13_242_518_0, i_13_242_520_0, i_13_242_521_0,
    i_13_242_535_0, i_13_242_645_0, i_13_242_661_0, i_13_242_739_0,
    i_13_242_756_0, i_13_242_820_0, i_13_242_850_0, i_13_242_851_0,
    i_13_242_870_0, i_13_242_938_0, i_13_242_1072_0, i_13_242_1073_0,
    i_13_242_1075_0, i_13_242_1201_0, i_13_242_1219_0, i_13_242_1262_0,
    i_13_242_1423_0, i_13_242_1424_0, i_13_242_1549_0, i_13_242_1550_0,
    i_13_242_1624_0, i_13_242_1630_0, i_13_242_1723_0, i_13_242_1758_0,
    i_13_242_1774_0, i_13_242_1787_0, i_13_242_1858_0, i_13_242_1939_0,
    i_13_242_1970_0, i_13_242_2027_0, i_13_242_2029_0, i_13_242_2033_0,
    i_13_242_2201_0, i_13_242_2209_0, i_13_242_2425_0, i_13_242_2451_0,
    i_13_242_2452_0, i_13_242_2454_0, i_13_242_2455_0, i_13_242_2558_0,
    i_13_242_2567_0, i_13_242_2612_0, i_13_242_2693_0, i_13_242_2764_0,
    i_13_242_2848_0, i_13_242_2850_0, i_13_242_3010_0, i_13_242_3011_0,
    i_13_242_3014_0, i_13_242_3037_0, i_13_242_3040_0, i_13_242_3143_0,
    i_13_242_3163_0, i_13_242_3217_0, i_13_242_3251_0, i_13_242_3272_0,
    i_13_242_3424_0, i_13_242_3442_0, i_13_242_3467_0, i_13_242_3472_0,
    i_13_242_3473_0, i_13_242_3485_0, i_13_242_3487_0, i_13_242_3488_0,
    i_13_242_3539_0, i_13_242_3541_0, i_13_242_3575_0, i_13_242_3731_0,
    i_13_242_3784_0, i_13_242_3853_0, i_13_242_3856_0, i_13_242_3863_0,
    i_13_242_3866_0, i_13_242_3893_0, i_13_242_3991_0, i_13_242_4038_0,
    i_13_242_4210_0, i_13_242_4216_0, i_13_242_4252_0, i_13_242_4253_0,
    i_13_242_4261_0, i_13_242_4262_0, i_13_242_4264_0, i_13_242_4265_0,
    i_13_242_4355_0, i_13_242_4370_0, i_13_242_4372_0, i_13_242_4379_0,
    i_13_242_4380_0, i_13_242_4511_0, i_13_242_4540_0, i_13_242_4558_0;
  output o_13_242_0_0;
  assign o_13_242_0_0 = ~((~i_13_242_518_0 & ((~i_13_242_521_0 & i_13_242_2209_0 & ~i_13_242_2455_0) | (~i_13_242_3014_0 & i_13_242_3893_0 & i_13_242_4355_0))) | (~i_13_242_1423_0 & ((~i_13_242_2029_0 & i_13_242_3784_0 & ~i_13_242_3856_0) | (i_13_242_121_0 & i_13_242_3217_0 & ~i_13_242_4262_0 & i_13_242_4558_0))) | (~i_13_242_3488_0 & ((i_13_242_1423_0 & ~i_13_242_3541_0 & ~i_13_242_3784_0) | (i_13_242_1624_0 & ~i_13_242_4370_0))) | (~i_13_242_4370_0 & ((i_13_242_229_0 & ~i_13_242_2454_0 & ~i_13_242_3011_0 & ~i_13_242_3853_0) | (~i_13_242_1424_0 & ~i_13_242_1549_0 & ~i_13_242_2029_0 & ~i_13_242_3575_0 & ~i_13_242_4265_0 & ~i_13_242_4379_0))) | (~i_13_242_230_0 & ~i_13_242_3010_0 & ~i_13_242_3040_0 & i_13_242_3217_0 & ~i_13_242_4262_0) | (~i_13_242_521_0 & ~i_13_242_2451_0 & ~i_13_242_4253_0 & ~i_13_242_4261_0 & ~i_13_242_4355_0));
endmodule



// Benchmark "kernel_13_243" written by ABC on Sun Jul 19 10:48:48 2020

module kernel_13_243 ( 
    i_13_243_37_0, i_13_243_77_0, i_13_243_104_0, i_13_243_112_0,
    i_13_243_117_0, i_13_243_337_0, i_13_243_379_0, i_13_243_451_0,
    i_13_243_452_0, i_13_243_461_0, i_13_243_561_0, i_13_243_583_0,
    i_13_243_586_0, i_13_243_589_0, i_13_243_643_0, i_13_243_676_0,
    i_13_243_724_0, i_13_243_769_0, i_13_243_914_0, i_13_243_949_0,
    i_13_243_950_0, i_13_243_1062_0, i_13_243_1064_0, i_13_243_1208_0,
    i_13_243_1243_0, i_13_243_1270_0, i_13_243_1297_0, i_13_243_1341_0,
    i_13_243_1342_0, i_13_243_1423_0, i_13_243_1427_0, i_13_243_1441_0,
    i_13_243_1495_0, i_13_243_1516_0, i_13_243_1594_0, i_13_243_1633_0,
    i_13_243_1693_0, i_13_243_1764_0, i_13_243_1811_0, i_13_243_1893_0,
    i_13_243_1945_0, i_13_243_2003_0, i_13_243_2099_0, i_13_243_2107_0,
    i_13_243_2108_0, i_13_243_2147_0, i_13_243_2197_0, i_13_243_2233_0,
    i_13_243_2234_0, i_13_243_2278_0, i_13_243_2542_0, i_13_243_2615_0,
    i_13_243_2650_0, i_13_243_2705_0, i_13_243_2710_0, i_13_243_2765_0,
    i_13_243_2782_0, i_13_243_2854_0, i_13_243_2898_0, i_13_243_2917_0,
    i_13_243_2918_0, i_13_243_2921_0, i_13_243_2926_0, i_13_243_3016_0,
    i_13_243_3017_0, i_13_243_3037_0, i_13_243_3064_0, i_13_243_3092_0,
    i_13_243_3136_0, i_13_243_3154_0, i_13_243_3199_0, i_13_243_3215_0,
    i_13_243_3218_0, i_13_243_3232_0, i_13_243_3289_0, i_13_243_3367_0,
    i_13_243_3415_0, i_13_243_3416_0, i_13_243_3532_0, i_13_243_3593_0,
    i_13_243_3739_0, i_13_243_3818_0, i_13_243_3874_0, i_13_243_3925_0,
    i_13_243_4019_0, i_13_243_4051_0, i_13_243_4087_0, i_13_243_4088_0,
    i_13_243_4106_0, i_13_243_4231_0, i_13_243_4232_0, i_13_243_4234_0,
    i_13_243_4250_0, i_13_243_4258_0, i_13_243_4267_0, i_13_243_4268_0,
    i_13_243_4393_0, i_13_243_4394_0, i_13_243_4448_0, i_13_243_4591_0,
    o_13_243_0_0  );
  input  i_13_243_37_0, i_13_243_77_0, i_13_243_104_0, i_13_243_112_0,
    i_13_243_117_0, i_13_243_337_0, i_13_243_379_0, i_13_243_451_0,
    i_13_243_452_0, i_13_243_461_0, i_13_243_561_0, i_13_243_583_0,
    i_13_243_586_0, i_13_243_589_0, i_13_243_643_0, i_13_243_676_0,
    i_13_243_724_0, i_13_243_769_0, i_13_243_914_0, i_13_243_949_0,
    i_13_243_950_0, i_13_243_1062_0, i_13_243_1064_0, i_13_243_1208_0,
    i_13_243_1243_0, i_13_243_1270_0, i_13_243_1297_0, i_13_243_1341_0,
    i_13_243_1342_0, i_13_243_1423_0, i_13_243_1427_0, i_13_243_1441_0,
    i_13_243_1495_0, i_13_243_1516_0, i_13_243_1594_0, i_13_243_1633_0,
    i_13_243_1693_0, i_13_243_1764_0, i_13_243_1811_0, i_13_243_1893_0,
    i_13_243_1945_0, i_13_243_2003_0, i_13_243_2099_0, i_13_243_2107_0,
    i_13_243_2108_0, i_13_243_2147_0, i_13_243_2197_0, i_13_243_2233_0,
    i_13_243_2234_0, i_13_243_2278_0, i_13_243_2542_0, i_13_243_2615_0,
    i_13_243_2650_0, i_13_243_2705_0, i_13_243_2710_0, i_13_243_2765_0,
    i_13_243_2782_0, i_13_243_2854_0, i_13_243_2898_0, i_13_243_2917_0,
    i_13_243_2918_0, i_13_243_2921_0, i_13_243_2926_0, i_13_243_3016_0,
    i_13_243_3017_0, i_13_243_3037_0, i_13_243_3064_0, i_13_243_3092_0,
    i_13_243_3136_0, i_13_243_3154_0, i_13_243_3199_0, i_13_243_3215_0,
    i_13_243_3218_0, i_13_243_3232_0, i_13_243_3289_0, i_13_243_3367_0,
    i_13_243_3415_0, i_13_243_3416_0, i_13_243_3532_0, i_13_243_3593_0,
    i_13_243_3739_0, i_13_243_3818_0, i_13_243_3874_0, i_13_243_3925_0,
    i_13_243_4019_0, i_13_243_4051_0, i_13_243_4087_0, i_13_243_4088_0,
    i_13_243_4106_0, i_13_243_4231_0, i_13_243_4232_0, i_13_243_4234_0,
    i_13_243_4250_0, i_13_243_4258_0, i_13_243_4267_0, i_13_243_4268_0,
    i_13_243_4393_0, i_13_243_4394_0, i_13_243_4448_0, i_13_243_4591_0;
  output o_13_243_0_0;
  assign o_13_243_0_0 = ~((~i_13_243_4088_0 & ~i_13_243_4267_0) | (~i_13_243_379_0 & ~i_13_243_4051_0) | (~i_13_243_1945_0 & ~i_13_243_2234_0) | (~i_13_243_112_0 & ~i_13_243_1811_0));
endmodule



// Benchmark "kernel_13_244" written by ABC on Sun Jul 19 10:48:49 2020

module kernel_13_244 ( 
    i_13_244_37_0, i_13_244_53_0, i_13_244_61_0, i_13_244_180_0,
    i_13_244_227_0, i_13_244_279_0, i_13_244_280_0, i_13_244_325_0,
    i_13_244_414_0, i_13_244_558_0, i_13_244_595_0, i_13_244_598_0,
    i_13_244_642_0, i_13_244_670_0, i_13_244_690_0, i_13_244_777_0,
    i_13_244_794_0, i_13_244_846_0, i_13_244_847_0, i_13_244_848_0,
    i_13_244_855_0, i_13_244_1073_0, i_13_244_1225_0, i_13_244_1252_0,
    i_13_244_1302_0, i_13_244_1314_0, i_13_244_1322_0, i_13_244_1404_0,
    i_13_244_1405_0, i_13_244_1444_0, i_13_244_1465_0, i_13_244_1479_0,
    i_13_244_1481_0, i_13_244_1483_0, i_13_244_1486_0, i_13_244_1548_0,
    i_13_244_1549_0, i_13_244_1574_0, i_13_244_1660_0, i_13_244_1746_0,
    i_13_244_1749_0, i_13_244_1776_0, i_13_244_1807_0, i_13_244_1854_0,
    i_13_244_1855_0, i_13_244_1856_0, i_13_244_1857_0, i_13_244_1858_0,
    i_13_244_1954_0, i_13_244_2022_0, i_13_244_2113_0, i_13_244_2134_0,
    i_13_244_2278_0, i_13_244_2281_0, i_13_244_2304_0, i_13_244_2307_0,
    i_13_244_2310_0, i_13_244_2311_0, i_13_244_2457_0, i_13_244_2458_0,
    i_13_244_2459_0, i_13_244_2553_0, i_13_244_2610_0, i_13_244_2629_0,
    i_13_244_2630_0, i_13_244_2636_0, i_13_244_2710_0, i_13_244_2877_0,
    i_13_244_2926_0, i_13_244_2937_0, i_13_244_3007_0, i_13_244_3019_0,
    i_13_244_3097_0, i_13_244_3129_0, i_13_244_3169_0, i_13_244_3170_0,
    i_13_244_3429_0, i_13_244_3448_0, i_13_244_3539_0, i_13_244_3579_0,
    i_13_244_3633_0, i_13_244_3741_0, i_13_244_3781_0, i_13_244_3791_0,
    i_13_244_3853_0, i_13_244_3907_0, i_13_244_3908_0, i_13_244_3910_0,
    i_13_244_3915_0, i_13_244_3987_0, i_13_244_4036_0, i_13_244_4059_0,
    i_13_244_4237_0, i_13_244_4267_0, i_13_244_4374_0, i_13_244_4375_0,
    i_13_244_4378_0, i_13_244_4381_0, i_13_244_4413_0, i_13_244_4518_0,
    o_13_244_0_0  );
  input  i_13_244_37_0, i_13_244_53_0, i_13_244_61_0, i_13_244_180_0,
    i_13_244_227_0, i_13_244_279_0, i_13_244_280_0, i_13_244_325_0,
    i_13_244_414_0, i_13_244_558_0, i_13_244_595_0, i_13_244_598_0,
    i_13_244_642_0, i_13_244_670_0, i_13_244_690_0, i_13_244_777_0,
    i_13_244_794_0, i_13_244_846_0, i_13_244_847_0, i_13_244_848_0,
    i_13_244_855_0, i_13_244_1073_0, i_13_244_1225_0, i_13_244_1252_0,
    i_13_244_1302_0, i_13_244_1314_0, i_13_244_1322_0, i_13_244_1404_0,
    i_13_244_1405_0, i_13_244_1444_0, i_13_244_1465_0, i_13_244_1479_0,
    i_13_244_1481_0, i_13_244_1483_0, i_13_244_1486_0, i_13_244_1548_0,
    i_13_244_1549_0, i_13_244_1574_0, i_13_244_1660_0, i_13_244_1746_0,
    i_13_244_1749_0, i_13_244_1776_0, i_13_244_1807_0, i_13_244_1854_0,
    i_13_244_1855_0, i_13_244_1856_0, i_13_244_1857_0, i_13_244_1858_0,
    i_13_244_1954_0, i_13_244_2022_0, i_13_244_2113_0, i_13_244_2134_0,
    i_13_244_2278_0, i_13_244_2281_0, i_13_244_2304_0, i_13_244_2307_0,
    i_13_244_2310_0, i_13_244_2311_0, i_13_244_2457_0, i_13_244_2458_0,
    i_13_244_2459_0, i_13_244_2553_0, i_13_244_2610_0, i_13_244_2629_0,
    i_13_244_2630_0, i_13_244_2636_0, i_13_244_2710_0, i_13_244_2877_0,
    i_13_244_2926_0, i_13_244_2937_0, i_13_244_3007_0, i_13_244_3019_0,
    i_13_244_3097_0, i_13_244_3129_0, i_13_244_3169_0, i_13_244_3170_0,
    i_13_244_3429_0, i_13_244_3448_0, i_13_244_3539_0, i_13_244_3579_0,
    i_13_244_3633_0, i_13_244_3741_0, i_13_244_3781_0, i_13_244_3791_0,
    i_13_244_3853_0, i_13_244_3907_0, i_13_244_3908_0, i_13_244_3910_0,
    i_13_244_3915_0, i_13_244_3987_0, i_13_244_4036_0, i_13_244_4059_0,
    i_13_244_4237_0, i_13_244_4267_0, i_13_244_4374_0, i_13_244_4375_0,
    i_13_244_4378_0, i_13_244_4381_0, i_13_244_4413_0, i_13_244_4518_0;
  output o_13_244_0_0;
  assign o_13_244_0_0 = ~((i_13_244_2281_0 & i_13_244_3097_0) | (~i_13_244_1405_0 & ~i_13_244_1776_0 & i_13_244_2710_0) | (~i_13_244_414_0 & ~i_13_244_1855_0 & ~i_13_244_2457_0) | (~i_13_244_1854_0 & ~i_13_244_2459_0 & ~i_13_244_3169_0 & ~i_13_244_4374_0) | (~i_13_244_1858_0 & ~i_13_244_2710_0 & ~i_13_244_3097_0 & i_13_244_3169_0) | (~i_13_244_279_0 & ~i_13_244_1252_0 & ~i_13_244_1954_0 & ~i_13_244_3781_0 & ~i_13_244_4375_0));
endmodule



// Benchmark "kernel_13_245" written by ABC on Sun Jul 19 10:48:49 2020

module kernel_13_245 ( 
    i_13_245_41_0, i_13_245_45_0, i_13_245_46_0, i_13_245_59_0,
    i_13_245_163_0, i_13_245_213_0, i_13_245_234_0, i_13_245_236_0,
    i_13_245_241_0, i_13_245_274_0, i_13_245_333_0, i_13_245_355_0,
    i_13_245_370_0, i_13_245_384_0, i_13_245_450_0, i_13_245_453_0,
    i_13_245_457_0, i_13_245_535_0, i_13_245_586_0, i_13_245_612_0,
    i_13_245_810_0, i_13_245_816_0, i_13_245_832_0, i_13_245_894_0,
    i_13_245_954_0, i_13_245_956_0, i_13_245_1219_0, i_13_245_1342_0,
    i_13_245_1459_0, i_13_245_1509_0, i_13_245_1521_0, i_13_245_1522_0,
    i_13_245_1524_0, i_13_245_1551_0, i_13_245_1552_0, i_13_245_1568_0,
    i_13_245_1696_0, i_13_245_1750_0, i_13_245_1765_0, i_13_245_1767_0,
    i_13_245_1891_0, i_13_245_1903_0, i_13_245_1927_0, i_13_245_2121_0,
    i_13_245_2142_0, i_13_245_2143_0, i_13_245_2144_0, i_13_245_2296_0,
    i_13_245_2394_0, i_13_245_2461_0, i_13_245_2560_0, i_13_245_2565_0,
    i_13_245_2568_0, i_13_245_2613_0, i_13_245_2691_0, i_13_245_2715_0,
    i_13_245_2716_0, i_13_245_2764_0, i_13_245_2766_0, i_13_245_2781_0,
    i_13_245_2782_0, i_13_245_2845_0, i_13_245_2881_0, i_13_245_2935_0,
    i_13_245_3028_0, i_13_245_3108_0, i_13_245_3142_0, i_13_245_3145_0,
    i_13_245_3146_0, i_13_245_3207_0, i_13_245_3231_0, i_13_245_3238_0,
    i_13_245_3274_0, i_13_245_3342_0, i_13_245_3366_0, i_13_245_3382_0,
    i_13_245_3546_0, i_13_245_3636_0, i_13_245_3754_0, i_13_245_3836_0,
    i_13_245_3856_0, i_13_245_3889_0, i_13_245_3900_0, i_13_245_3902_0,
    i_13_245_3916_0, i_13_245_3921_0, i_13_245_3982_0, i_13_245_4017_0,
    i_13_245_4052_0, i_13_245_4081_0, i_13_245_4086_0, i_13_245_4249_0,
    i_13_245_4269_0, i_13_245_4270_0, i_13_245_4311_0, i_13_245_4312_0,
    i_13_245_4428_0, i_13_245_4509_0, i_13_245_4510_0, i_13_245_4533_0,
    o_13_245_0_0  );
  input  i_13_245_41_0, i_13_245_45_0, i_13_245_46_0, i_13_245_59_0,
    i_13_245_163_0, i_13_245_213_0, i_13_245_234_0, i_13_245_236_0,
    i_13_245_241_0, i_13_245_274_0, i_13_245_333_0, i_13_245_355_0,
    i_13_245_370_0, i_13_245_384_0, i_13_245_450_0, i_13_245_453_0,
    i_13_245_457_0, i_13_245_535_0, i_13_245_586_0, i_13_245_612_0,
    i_13_245_810_0, i_13_245_816_0, i_13_245_832_0, i_13_245_894_0,
    i_13_245_954_0, i_13_245_956_0, i_13_245_1219_0, i_13_245_1342_0,
    i_13_245_1459_0, i_13_245_1509_0, i_13_245_1521_0, i_13_245_1522_0,
    i_13_245_1524_0, i_13_245_1551_0, i_13_245_1552_0, i_13_245_1568_0,
    i_13_245_1696_0, i_13_245_1750_0, i_13_245_1765_0, i_13_245_1767_0,
    i_13_245_1891_0, i_13_245_1903_0, i_13_245_1927_0, i_13_245_2121_0,
    i_13_245_2142_0, i_13_245_2143_0, i_13_245_2144_0, i_13_245_2296_0,
    i_13_245_2394_0, i_13_245_2461_0, i_13_245_2560_0, i_13_245_2565_0,
    i_13_245_2568_0, i_13_245_2613_0, i_13_245_2691_0, i_13_245_2715_0,
    i_13_245_2716_0, i_13_245_2764_0, i_13_245_2766_0, i_13_245_2781_0,
    i_13_245_2782_0, i_13_245_2845_0, i_13_245_2881_0, i_13_245_2935_0,
    i_13_245_3028_0, i_13_245_3108_0, i_13_245_3142_0, i_13_245_3145_0,
    i_13_245_3146_0, i_13_245_3207_0, i_13_245_3231_0, i_13_245_3238_0,
    i_13_245_3274_0, i_13_245_3342_0, i_13_245_3366_0, i_13_245_3382_0,
    i_13_245_3546_0, i_13_245_3636_0, i_13_245_3754_0, i_13_245_3836_0,
    i_13_245_3856_0, i_13_245_3889_0, i_13_245_3900_0, i_13_245_3902_0,
    i_13_245_3916_0, i_13_245_3921_0, i_13_245_3982_0, i_13_245_4017_0,
    i_13_245_4052_0, i_13_245_4081_0, i_13_245_4086_0, i_13_245_4249_0,
    i_13_245_4269_0, i_13_245_4270_0, i_13_245_4311_0, i_13_245_4312_0,
    i_13_245_4428_0, i_13_245_4509_0, i_13_245_4510_0, i_13_245_4533_0;
  output o_13_245_0_0;
  assign o_13_245_0_0 = ~((~i_13_245_4311_0 & ((~i_13_245_832_0 & ~i_13_245_2144_0 & ~i_13_245_3231_0) | (~i_13_245_2782_0 & ~i_13_245_4052_0 & ~i_13_245_4081_0))) | (~i_13_245_1552_0 & ~i_13_245_1568_0 & ~i_13_245_4269_0 & ~i_13_245_4312_0) | (~i_13_245_234_0 & ~i_13_245_1522_0 & ~i_13_245_2143_0 & ~i_13_245_4428_0));
endmodule



// Benchmark "kernel_13_246" written by ABC on Sun Jul 19 10:48:50 2020

module kernel_13_246 ( 
    i_13_246_53_0, i_13_246_76_0, i_13_246_77_0, i_13_246_116_0,
    i_13_246_166_0, i_13_246_184_0, i_13_246_193_0, i_13_246_203_0,
    i_13_246_446_0, i_13_246_530_0, i_13_246_554_0, i_13_246_561_0,
    i_13_246_571_0, i_13_246_592_0, i_13_246_655_0, i_13_246_656_0,
    i_13_246_671_0, i_13_246_697_0, i_13_246_698_0, i_13_246_700_0,
    i_13_246_826_0, i_13_246_944_0, i_13_246_1084_0, i_13_246_1085_0,
    i_13_246_1147_0, i_13_246_1148_0, i_13_246_1211_0, i_13_246_1223_0,
    i_13_246_1267_0, i_13_246_1285_0, i_13_246_1430_0, i_13_246_1502_0,
    i_13_246_1508_0, i_13_246_1517_0, i_13_246_1525_0, i_13_246_1552_0,
    i_13_246_1636_0, i_13_246_1637_0, i_13_246_1660_0, i_13_246_1661_0,
    i_13_246_1664_0, i_13_246_1741_0, i_13_246_1831_0, i_13_246_1840_0,
    i_13_246_1843_0, i_13_246_1844_0, i_13_246_1885_0, i_13_246_1886_0,
    i_13_246_2033_0, i_13_246_2172_0, i_13_246_2245_0, i_13_246_2314_0,
    i_13_246_2321_0, i_13_246_2354_0, i_13_246_2398_0, i_13_246_2438_0,
    i_13_246_2455_0, i_13_246_2456_0, i_13_246_2510_0, i_13_246_2762_0,
    i_13_246_2848_0, i_13_246_2849_0, i_13_246_2887_0, i_13_246_2924_0,
    i_13_246_2959_0, i_13_246_2983_0, i_13_246_3001_0, i_13_246_3002_0,
    i_13_246_3004_0, i_13_246_3050_0, i_13_246_3130_0, i_13_246_3383_0,
    i_13_246_3436_0, i_13_246_3467_0, i_13_246_3476_0, i_13_246_3505_0,
    i_13_246_3571_0, i_13_246_3572_0, i_13_246_3599_0, i_13_246_3602_0,
    i_13_246_3649_0, i_13_246_3650_0, i_13_246_3689_0, i_13_246_3740_0,
    i_13_246_3742_0, i_13_246_3866_0, i_13_246_3875_0, i_13_246_4021_0,
    i_13_246_4045_0, i_13_246_4063_0, i_13_246_4190_0, i_13_246_4264_0,
    i_13_246_4279_0, i_13_246_4301_0, i_13_246_4333_0, i_13_246_4378_0,
    i_13_246_4417_0, i_13_246_4594_0, i_13_246_4603_0, i_13_246_4604_0,
    o_13_246_0_0  );
  input  i_13_246_53_0, i_13_246_76_0, i_13_246_77_0, i_13_246_116_0,
    i_13_246_166_0, i_13_246_184_0, i_13_246_193_0, i_13_246_203_0,
    i_13_246_446_0, i_13_246_530_0, i_13_246_554_0, i_13_246_561_0,
    i_13_246_571_0, i_13_246_592_0, i_13_246_655_0, i_13_246_656_0,
    i_13_246_671_0, i_13_246_697_0, i_13_246_698_0, i_13_246_700_0,
    i_13_246_826_0, i_13_246_944_0, i_13_246_1084_0, i_13_246_1085_0,
    i_13_246_1147_0, i_13_246_1148_0, i_13_246_1211_0, i_13_246_1223_0,
    i_13_246_1267_0, i_13_246_1285_0, i_13_246_1430_0, i_13_246_1502_0,
    i_13_246_1508_0, i_13_246_1517_0, i_13_246_1525_0, i_13_246_1552_0,
    i_13_246_1636_0, i_13_246_1637_0, i_13_246_1660_0, i_13_246_1661_0,
    i_13_246_1664_0, i_13_246_1741_0, i_13_246_1831_0, i_13_246_1840_0,
    i_13_246_1843_0, i_13_246_1844_0, i_13_246_1885_0, i_13_246_1886_0,
    i_13_246_2033_0, i_13_246_2172_0, i_13_246_2245_0, i_13_246_2314_0,
    i_13_246_2321_0, i_13_246_2354_0, i_13_246_2398_0, i_13_246_2438_0,
    i_13_246_2455_0, i_13_246_2456_0, i_13_246_2510_0, i_13_246_2762_0,
    i_13_246_2848_0, i_13_246_2849_0, i_13_246_2887_0, i_13_246_2924_0,
    i_13_246_2959_0, i_13_246_2983_0, i_13_246_3001_0, i_13_246_3002_0,
    i_13_246_3004_0, i_13_246_3050_0, i_13_246_3130_0, i_13_246_3383_0,
    i_13_246_3436_0, i_13_246_3467_0, i_13_246_3476_0, i_13_246_3505_0,
    i_13_246_3571_0, i_13_246_3572_0, i_13_246_3599_0, i_13_246_3602_0,
    i_13_246_3649_0, i_13_246_3650_0, i_13_246_3689_0, i_13_246_3740_0,
    i_13_246_3742_0, i_13_246_3866_0, i_13_246_3875_0, i_13_246_4021_0,
    i_13_246_4045_0, i_13_246_4063_0, i_13_246_4190_0, i_13_246_4264_0,
    i_13_246_4279_0, i_13_246_4301_0, i_13_246_4333_0, i_13_246_4378_0,
    i_13_246_4417_0, i_13_246_4594_0, i_13_246_4603_0, i_13_246_4604_0;
  output o_13_246_0_0;
  assign o_13_246_0_0 = 0;
endmodule



// Benchmark "kernel_13_247" written by ABC on Sun Jul 19 10:48:51 2020

module kernel_13_247 ( 
    i_13_247_74_0, i_13_247_91_0, i_13_247_94_0, i_13_247_103_0,
    i_13_247_104_0, i_13_247_109_0, i_13_247_112_0, i_13_247_118_0,
    i_13_247_166_0, i_13_247_201_0, i_13_247_263_0, i_13_247_364_0,
    i_13_247_607_0, i_13_247_643_0, i_13_247_730_0, i_13_247_733_0,
    i_13_247_768_0, i_13_247_793_0, i_13_247_794_0, i_13_247_856_0,
    i_13_247_946_0, i_13_247_1084_0, i_13_247_1086_0, i_13_247_1102_0,
    i_13_247_1144_0, i_13_247_1217_0, i_13_247_1273_0, i_13_247_1486_0,
    i_13_247_1487_0, i_13_247_1552_0, i_13_247_1621_0, i_13_247_1630_0,
    i_13_247_1692_0, i_13_247_1774_0, i_13_247_1775_0, i_13_247_1836_0,
    i_13_247_1837_0, i_13_247_1839_0, i_13_247_1846_0, i_13_247_2000_0,
    i_13_247_2009_0, i_13_247_2137_0, i_13_247_2170_0, i_13_247_2172_0,
    i_13_247_2173_0, i_13_247_2201_0, i_13_247_2381_0, i_13_247_2407_0,
    i_13_247_2422_0, i_13_247_2430_0, i_13_247_2431_0, i_13_247_2434_0,
    i_13_247_2497_0, i_13_247_2498_0, i_13_247_2539_0, i_13_247_2542_0,
    i_13_247_2569_0, i_13_247_2579_0, i_13_247_2611_0, i_13_247_2875_0,
    i_13_247_2943_0, i_13_247_2958_0, i_13_247_3024_0, i_13_247_3054_0,
    i_13_247_3100_0, i_13_247_3143_0, i_13_247_3145_0, i_13_247_3146_0,
    i_13_247_3370_0, i_13_247_3375_0, i_13_247_3452_0, i_13_247_3525_0,
    i_13_247_3529_0, i_13_247_3530_0, i_13_247_3646_0, i_13_247_3696_0,
    i_13_247_3739_0, i_13_247_3864_0, i_13_247_3871_0, i_13_247_3872_0,
    i_13_247_3891_0, i_13_247_4036_0, i_13_247_4063_0, i_13_247_4091_0,
    i_13_247_4106_0, i_13_247_4118_0, i_13_247_4119_0, i_13_247_4122_0,
    i_13_247_4234_0, i_13_247_4252_0, i_13_247_4263_0, i_13_247_4339_0,
    i_13_247_4351_0, i_13_247_4367_0, i_13_247_4413_0, i_13_247_4417_0,
    i_13_247_4431_0, i_13_247_4542_0, i_13_247_4559_0, i_13_247_4560_0,
    o_13_247_0_0  );
  input  i_13_247_74_0, i_13_247_91_0, i_13_247_94_0, i_13_247_103_0,
    i_13_247_104_0, i_13_247_109_0, i_13_247_112_0, i_13_247_118_0,
    i_13_247_166_0, i_13_247_201_0, i_13_247_263_0, i_13_247_364_0,
    i_13_247_607_0, i_13_247_643_0, i_13_247_730_0, i_13_247_733_0,
    i_13_247_768_0, i_13_247_793_0, i_13_247_794_0, i_13_247_856_0,
    i_13_247_946_0, i_13_247_1084_0, i_13_247_1086_0, i_13_247_1102_0,
    i_13_247_1144_0, i_13_247_1217_0, i_13_247_1273_0, i_13_247_1486_0,
    i_13_247_1487_0, i_13_247_1552_0, i_13_247_1621_0, i_13_247_1630_0,
    i_13_247_1692_0, i_13_247_1774_0, i_13_247_1775_0, i_13_247_1836_0,
    i_13_247_1837_0, i_13_247_1839_0, i_13_247_1846_0, i_13_247_2000_0,
    i_13_247_2009_0, i_13_247_2137_0, i_13_247_2170_0, i_13_247_2172_0,
    i_13_247_2173_0, i_13_247_2201_0, i_13_247_2381_0, i_13_247_2407_0,
    i_13_247_2422_0, i_13_247_2430_0, i_13_247_2431_0, i_13_247_2434_0,
    i_13_247_2497_0, i_13_247_2498_0, i_13_247_2539_0, i_13_247_2542_0,
    i_13_247_2569_0, i_13_247_2579_0, i_13_247_2611_0, i_13_247_2875_0,
    i_13_247_2943_0, i_13_247_2958_0, i_13_247_3024_0, i_13_247_3054_0,
    i_13_247_3100_0, i_13_247_3143_0, i_13_247_3145_0, i_13_247_3146_0,
    i_13_247_3370_0, i_13_247_3375_0, i_13_247_3452_0, i_13_247_3525_0,
    i_13_247_3529_0, i_13_247_3530_0, i_13_247_3646_0, i_13_247_3696_0,
    i_13_247_3739_0, i_13_247_3864_0, i_13_247_3871_0, i_13_247_3872_0,
    i_13_247_3891_0, i_13_247_4036_0, i_13_247_4063_0, i_13_247_4091_0,
    i_13_247_4106_0, i_13_247_4118_0, i_13_247_4119_0, i_13_247_4122_0,
    i_13_247_4234_0, i_13_247_4252_0, i_13_247_4263_0, i_13_247_4339_0,
    i_13_247_4351_0, i_13_247_4367_0, i_13_247_4413_0, i_13_247_4417_0,
    i_13_247_4431_0, i_13_247_4542_0, i_13_247_4559_0, i_13_247_4560_0;
  output o_13_247_0_0;
  assign o_13_247_0_0 = ~(~i_13_247_3529_0 | ~i_13_247_109_0 | (~i_13_247_1775_0 & ~i_13_247_3143_0));
endmodule



// Benchmark "kernel_13_248" written by ABC on Sun Jul 19 10:48:52 2020

module kernel_13_248 ( 
    i_13_248_97_0, i_13_248_154_0, i_13_248_164_0, i_13_248_217_0,
    i_13_248_251_0, i_13_248_272_0, i_13_248_319_0, i_13_248_355_0,
    i_13_248_451_0, i_13_248_559_0, i_13_248_688_0, i_13_248_895_0,
    i_13_248_928_0, i_13_248_929_0, i_13_248_966_0, i_13_248_974_0,
    i_13_248_1081_0, i_13_248_1099_0, i_13_248_1120_0, i_13_248_1252_0,
    i_13_248_1262_0, i_13_248_1283_0, i_13_248_1298_0, i_13_248_1340_0,
    i_13_248_1372_0, i_13_248_1396_0, i_13_248_1397_0, i_13_248_1468_0,
    i_13_248_1502_0, i_13_248_1505_0, i_13_248_1568_0, i_13_248_1606_0,
    i_13_248_1628_0, i_13_248_1633_0, i_13_248_1786_0, i_13_248_1811_0,
    i_13_248_1855_0, i_13_248_1858_0, i_13_248_1891_0, i_13_248_1910_0,
    i_13_248_1928_0, i_13_248_1990_0, i_13_248_2003_0, i_13_248_2108_0,
    i_13_248_2117_0, i_13_248_2180_0, i_13_248_2234_0, i_13_248_2314_0,
    i_13_248_2333_0, i_13_248_2430_0, i_13_248_2467_0, i_13_248_2483_0,
    i_13_248_2542_0, i_13_248_2543_0, i_13_248_2696_0, i_13_248_2711_0,
    i_13_248_2755_0, i_13_248_2764_0, i_13_248_2765_0, i_13_248_2785_0,
    i_13_248_2786_0, i_13_248_2935_0, i_13_248_2936_0, i_13_248_2958_0,
    i_13_248_3016_0, i_13_248_3017_0, i_13_248_3061_0, i_13_248_3062_0,
    i_13_248_3206_0, i_13_248_3218_0, i_13_248_3231_0, i_13_248_3234_0,
    i_13_248_3239_0, i_13_248_3242_0, i_13_248_3271_0, i_13_248_3312_0,
    i_13_248_3313_0, i_13_248_3340_0, i_13_248_3341_0, i_13_248_3532_0,
    i_13_248_3601_0, i_13_248_3683_0, i_13_248_3709_0, i_13_248_3723_0,
    i_13_248_3851_0, i_13_248_3920_0, i_13_248_4081_0, i_13_248_4082_0,
    i_13_248_4087_0, i_13_248_4160_0, i_13_248_4214_0, i_13_248_4266_0,
    i_13_248_4268_0, i_13_248_4313_0, i_13_248_4361_0, i_13_248_4430_0,
    i_13_248_4453_0, i_13_248_4462_0, i_13_248_4466_0, i_13_248_4595_0,
    o_13_248_0_0  );
  input  i_13_248_97_0, i_13_248_154_0, i_13_248_164_0, i_13_248_217_0,
    i_13_248_251_0, i_13_248_272_0, i_13_248_319_0, i_13_248_355_0,
    i_13_248_451_0, i_13_248_559_0, i_13_248_688_0, i_13_248_895_0,
    i_13_248_928_0, i_13_248_929_0, i_13_248_966_0, i_13_248_974_0,
    i_13_248_1081_0, i_13_248_1099_0, i_13_248_1120_0, i_13_248_1252_0,
    i_13_248_1262_0, i_13_248_1283_0, i_13_248_1298_0, i_13_248_1340_0,
    i_13_248_1372_0, i_13_248_1396_0, i_13_248_1397_0, i_13_248_1468_0,
    i_13_248_1502_0, i_13_248_1505_0, i_13_248_1568_0, i_13_248_1606_0,
    i_13_248_1628_0, i_13_248_1633_0, i_13_248_1786_0, i_13_248_1811_0,
    i_13_248_1855_0, i_13_248_1858_0, i_13_248_1891_0, i_13_248_1910_0,
    i_13_248_1928_0, i_13_248_1990_0, i_13_248_2003_0, i_13_248_2108_0,
    i_13_248_2117_0, i_13_248_2180_0, i_13_248_2234_0, i_13_248_2314_0,
    i_13_248_2333_0, i_13_248_2430_0, i_13_248_2467_0, i_13_248_2483_0,
    i_13_248_2542_0, i_13_248_2543_0, i_13_248_2696_0, i_13_248_2711_0,
    i_13_248_2755_0, i_13_248_2764_0, i_13_248_2765_0, i_13_248_2785_0,
    i_13_248_2786_0, i_13_248_2935_0, i_13_248_2936_0, i_13_248_2958_0,
    i_13_248_3016_0, i_13_248_3017_0, i_13_248_3061_0, i_13_248_3062_0,
    i_13_248_3206_0, i_13_248_3218_0, i_13_248_3231_0, i_13_248_3234_0,
    i_13_248_3239_0, i_13_248_3242_0, i_13_248_3271_0, i_13_248_3312_0,
    i_13_248_3313_0, i_13_248_3340_0, i_13_248_3341_0, i_13_248_3532_0,
    i_13_248_3601_0, i_13_248_3683_0, i_13_248_3709_0, i_13_248_3723_0,
    i_13_248_3851_0, i_13_248_3920_0, i_13_248_4081_0, i_13_248_4082_0,
    i_13_248_4087_0, i_13_248_4160_0, i_13_248_4214_0, i_13_248_4266_0,
    i_13_248_4268_0, i_13_248_4313_0, i_13_248_4361_0, i_13_248_4430_0,
    i_13_248_4453_0, i_13_248_4462_0, i_13_248_4466_0, i_13_248_4595_0;
  output o_13_248_0_0;
  assign o_13_248_0_0 = ~((~i_13_248_2542_0 & ~i_13_248_4430_0) | (~i_13_248_2935_0 & ~i_13_248_3313_0) | (~i_13_248_1396_0 & ~i_13_248_1397_0 & ~i_13_248_4268_0) | (i_13_248_2785_0 & ~i_13_248_3061_0 & ~i_13_248_3601_0 & ~i_13_248_4214_0) | (~i_13_248_1468_0 & ~i_13_248_2711_0 & ~i_13_248_2936_0 & ~i_13_248_3234_0));
endmodule



// Benchmark "kernel_13_249" written by ABC on Sun Jul 19 10:48:53 2020

module kernel_13_249 ( 
    i_13_249_34_0, i_13_249_47_0, i_13_249_139_0, i_13_249_143_0,
    i_13_249_184_0, i_13_249_233_0, i_13_249_380_0, i_13_249_383_0,
    i_13_249_385_0, i_13_249_386_0, i_13_249_529_0, i_13_249_649_0,
    i_13_249_666_0, i_13_249_675_0, i_13_249_701_0, i_13_249_763_0,
    i_13_249_824_0, i_13_249_871_0, i_13_249_883_0, i_13_249_985_0,
    i_13_249_1082_0, i_13_249_1206_0, i_13_249_1220_0, i_13_249_1281_0,
    i_13_249_1326_0, i_13_249_1403_0, i_13_249_1442_0, i_13_249_1445_0,
    i_13_249_1502_0, i_13_249_1511_0, i_13_249_1516_0, i_13_249_1600_0,
    i_13_249_1664_0, i_13_249_1678_0, i_13_249_1684_0, i_13_249_1750_0,
    i_13_249_1780_0, i_13_249_1787_0, i_13_249_1817_0, i_13_249_1861_0,
    i_13_249_1912_0, i_13_249_1930_0, i_13_249_2002_0, i_13_249_2003_0,
    i_13_249_2005_0, i_13_249_2006_0, i_13_249_2054_0, i_13_249_2177_0,
    i_13_249_2189_0, i_13_249_2196_0, i_13_249_2210_0, i_13_249_2246_0,
    i_13_249_2259_0, i_13_249_2266_0, i_13_249_2279_0, i_13_249_2351_0,
    i_13_249_2537_0, i_13_249_2543_0, i_13_249_2677_0, i_13_249_2708_0,
    i_13_249_2719_0, i_13_249_2722_0, i_13_249_2723_0, i_13_249_2725_0,
    i_13_249_2726_0, i_13_249_2854_0, i_13_249_2855_0, i_13_249_2858_0,
    i_13_249_2861_0, i_13_249_2969_0, i_13_249_3218_0, i_13_249_3347_0,
    i_13_249_3379_0, i_13_249_3392_0, i_13_249_3418_0, i_13_249_3419_0,
    i_13_249_3442_0, i_13_249_3577_0, i_13_249_3593_0, i_13_249_3614_0,
    i_13_249_3653_0, i_13_249_3686_0, i_13_249_3730_0, i_13_249_3844_0,
    i_13_249_3865_0, i_13_249_3873_0, i_13_249_3892_0, i_13_249_3917_0,
    i_13_249_4052_0, i_13_249_4057_0, i_13_249_4058_0, i_13_249_4171_0,
    i_13_249_4268_0, i_13_249_4273_0, i_13_249_4282_0, i_13_249_4345_0,
    i_13_249_4394_0, i_13_249_4400_0, i_13_249_4568_0, i_13_249_4583_0,
    o_13_249_0_0  );
  input  i_13_249_34_0, i_13_249_47_0, i_13_249_139_0, i_13_249_143_0,
    i_13_249_184_0, i_13_249_233_0, i_13_249_380_0, i_13_249_383_0,
    i_13_249_385_0, i_13_249_386_0, i_13_249_529_0, i_13_249_649_0,
    i_13_249_666_0, i_13_249_675_0, i_13_249_701_0, i_13_249_763_0,
    i_13_249_824_0, i_13_249_871_0, i_13_249_883_0, i_13_249_985_0,
    i_13_249_1082_0, i_13_249_1206_0, i_13_249_1220_0, i_13_249_1281_0,
    i_13_249_1326_0, i_13_249_1403_0, i_13_249_1442_0, i_13_249_1445_0,
    i_13_249_1502_0, i_13_249_1511_0, i_13_249_1516_0, i_13_249_1600_0,
    i_13_249_1664_0, i_13_249_1678_0, i_13_249_1684_0, i_13_249_1750_0,
    i_13_249_1780_0, i_13_249_1787_0, i_13_249_1817_0, i_13_249_1861_0,
    i_13_249_1912_0, i_13_249_1930_0, i_13_249_2002_0, i_13_249_2003_0,
    i_13_249_2005_0, i_13_249_2006_0, i_13_249_2054_0, i_13_249_2177_0,
    i_13_249_2189_0, i_13_249_2196_0, i_13_249_2210_0, i_13_249_2246_0,
    i_13_249_2259_0, i_13_249_2266_0, i_13_249_2279_0, i_13_249_2351_0,
    i_13_249_2537_0, i_13_249_2543_0, i_13_249_2677_0, i_13_249_2708_0,
    i_13_249_2719_0, i_13_249_2722_0, i_13_249_2723_0, i_13_249_2725_0,
    i_13_249_2726_0, i_13_249_2854_0, i_13_249_2855_0, i_13_249_2858_0,
    i_13_249_2861_0, i_13_249_2969_0, i_13_249_3218_0, i_13_249_3347_0,
    i_13_249_3379_0, i_13_249_3392_0, i_13_249_3418_0, i_13_249_3419_0,
    i_13_249_3442_0, i_13_249_3577_0, i_13_249_3593_0, i_13_249_3614_0,
    i_13_249_3653_0, i_13_249_3686_0, i_13_249_3730_0, i_13_249_3844_0,
    i_13_249_3865_0, i_13_249_3873_0, i_13_249_3892_0, i_13_249_3917_0,
    i_13_249_4052_0, i_13_249_4057_0, i_13_249_4058_0, i_13_249_4171_0,
    i_13_249_4268_0, i_13_249_4273_0, i_13_249_4282_0, i_13_249_4345_0,
    i_13_249_4394_0, i_13_249_4400_0, i_13_249_4568_0, i_13_249_4583_0;
  output o_13_249_0_0;
  assign o_13_249_0_0 = ~((i_13_249_985_0 & ~i_13_249_3442_0) | (~i_13_249_383_0 & ~i_13_249_2861_0) | (~i_13_249_386_0 & ~i_13_249_701_0));
endmodule



// Benchmark "kernel_13_250" written by ABC on Sun Jul 19 10:48:54 2020

module kernel_13_250 ( 
    i_13_250_47_0, i_13_250_65_0, i_13_250_169_0, i_13_250_170_0,
    i_13_250_319_0, i_13_250_438_0, i_13_250_463_0, i_13_250_524_0,
    i_13_250_538_0, i_13_250_623_0, i_13_250_659_0, i_13_250_667_0,
    i_13_250_848_0, i_13_250_937_0, i_13_250_938_0, i_13_250_1018_0,
    i_13_250_1019_0, i_13_250_1072_0, i_13_250_1073_0, i_13_250_1086_0,
    i_13_250_1095_0, i_13_250_1096_0, i_13_250_1100_0, i_13_250_1252_0,
    i_13_250_1253_0, i_13_250_1315_0, i_13_250_1365_0, i_13_250_1400_0,
    i_13_250_1428_0, i_13_250_1488_0, i_13_250_1550_0, i_13_250_1596_0,
    i_13_250_1662_0, i_13_250_1694_0, i_13_250_1778_0, i_13_250_1792_0,
    i_13_250_1825_0, i_13_250_1913_0, i_13_250_1947_0, i_13_250_2026_0,
    i_13_250_2027_0, i_13_250_2056_0, i_13_250_2103_0, i_13_250_2122_0,
    i_13_250_2197_0, i_13_250_2227_0, i_13_250_2360_0, i_13_250_2364_0,
    i_13_250_2373_0, i_13_250_2770_0, i_13_250_2910_0, i_13_250_2915_0,
    i_13_250_2918_0, i_13_250_2975_0, i_13_250_3001_0, i_13_250_3008_0,
    i_13_250_3010_0, i_13_250_3103_0, i_13_250_3120_0, i_13_250_3166_0,
    i_13_250_3265_0, i_13_250_3352_0, i_13_250_3353_0, i_13_250_3382_0,
    i_13_250_3432_0, i_13_250_3452_0, i_13_250_3454_0, i_13_250_3459_0,
    i_13_250_3484_0, i_13_250_3534_0, i_13_250_3538_0, i_13_250_3539_0,
    i_13_250_3574_0, i_13_250_3575_0, i_13_250_3727_0, i_13_250_3741_0,
    i_13_250_3781_0, i_13_250_3782_0, i_13_250_3783_0, i_13_250_3820_0,
    i_13_250_3840_0, i_13_250_3847_0, i_13_250_3853_0, i_13_250_3859_0,
    i_13_250_3893_0, i_13_250_3908_0, i_13_250_3918_0, i_13_250_4063_0,
    i_13_250_4108_0, i_13_250_4150_0, i_13_250_4250_0, i_13_250_4253_0,
    i_13_250_4259_0, i_13_250_4335_0, i_13_250_4336_0, i_13_250_4344_0,
    i_13_250_4448_0, i_13_250_4583_0, i_13_250_4604_0, i_13_250_4605_0,
    o_13_250_0_0  );
  input  i_13_250_47_0, i_13_250_65_0, i_13_250_169_0, i_13_250_170_0,
    i_13_250_319_0, i_13_250_438_0, i_13_250_463_0, i_13_250_524_0,
    i_13_250_538_0, i_13_250_623_0, i_13_250_659_0, i_13_250_667_0,
    i_13_250_848_0, i_13_250_937_0, i_13_250_938_0, i_13_250_1018_0,
    i_13_250_1019_0, i_13_250_1072_0, i_13_250_1073_0, i_13_250_1086_0,
    i_13_250_1095_0, i_13_250_1096_0, i_13_250_1100_0, i_13_250_1252_0,
    i_13_250_1253_0, i_13_250_1315_0, i_13_250_1365_0, i_13_250_1400_0,
    i_13_250_1428_0, i_13_250_1488_0, i_13_250_1550_0, i_13_250_1596_0,
    i_13_250_1662_0, i_13_250_1694_0, i_13_250_1778_0, i_13_250_1792_0,
    i_13_250_1825_0, i_13_250_1913_0, i_13_250_1947_0, i_13_250_2026_0,
    i_13_250_2027_0, i_13_250_2056_0, i_13_250_2103_0, i_13_250_2122_0,
    i_13_250_2197_0, i_13_250_2227_0, i_13_250_2360_0, i_13_250_2364_0,
    i_13_250_2373_0, i_13_250_2770_0, i_13_250_2910_0, i_13_250_2915_0,
    i_13_250_2918_0, i_13_250_2975_0, i_13_250_3001_0, i_13_250_3008_0,
    i_13_250_3010_0, i_13_250_3103_0, i_13_250_3120_0, i_13_250_3166_0,
    i_13_250_3265_0, i_13_250_3352_0, i_13_250_3353_0, i_13_250_3382_0,
    i_13_250_3432_0, i_13_250_3452_0, i_13_250_3454_0, i_13_250_3459_0,
    i_13_250_3484_0, i_13_250_3534_0, i_13_250_3538_0, i_13_250_3539_0,
    i_13_250_3574_0, i_13_250_3575_0, i_13_250_3727_0, i_13_250_3741_0,
    i_13_250_3781_0, i_13_250_3782_0, i_13_250_3783_0, i_13_250_3820_0,
    i_13_250_3840_0, i_13_250_3847_0, i_13_250_3853_0, i_13_250_3859_0,
    i_13_250_3893_0, i_13_250_3908_0, i_13_250_3918_0, i_13_250_4063_0,
    i_13_250_4108_0, i_13_250_4150_0, i_13_250_4250_0, i_13_250_4253_0,
    i_13_250_4259_0, i_13_250_4335_0, i_13_250_4336_0, i_13_250_4344_0,
    i_13_250_4448_0, i_13_250_4583_0, i_13_250_4604_0, i_13_250_4605_0;
  output o_13_250_0_0;
  assign o_13_250_0_0 = ~(~i_13_250_3574_0 | (~i_13_250_3575_0 & (~i_13_250_1315_0 | ~i_13_250_2918_0)));
endmodule



// Benchmark "kernel_13_251" written by ABC on Sun Jul 19 10:48:55 2020

module kernel_13_251 ( 
    i_13_251_37_0, i_13_251_38_0, i_13_251_51_0, i_13_251_75_0,
    i_13_251_76_0, i_13_251_103_0, i_13_251_112_0, i_13_251_165_0,
    i_13_251_173_0, i_13_251_181_0, i_13_251_184_0, i_13_251_240_0,
    i_13_251_252_0, i_13_251_280_0, i_13_251_281_0, i_13_251_324_0,
    i_13_251_325_0, i_13_251_339_0, i_13_251_571_0, i_13_251_577_0,
    i_13_251_596_0, i_13_251_597_0, i_13_251_598_0, i_13_251_618_0,
    i_13_251_640_0, i_13_251_643_0, i_13_251_685_0, i_13_251_715_0,
    i_13_251_744_0, i_13_251_778_0, i_13_251_814_0, i_13_251_840_0,
    i_13_251_891_0, i_13_251_892_0, i_13_251_894_0, i_13_251_896_0,
    i_13_251_1031_0, i_13_251_1093_0, i_13_251_1248_0, i_13_251_1249_0,
    i_13_251_1462_0, i_13_251_1480_0, i_13_251_1541_0, i_13_251_1711_0,
    i_13_251_1746_0, i_13_251_1747_0, i_13_251_1786_0, i_13_251_1804_0,
    i_13_251_1805_0, i_13_251_1806_0, i_13_251_1854_0, i_13_251_1855_0,
    i_13_251_1856_0, i_13_251_1858_0, i_13_251_2119_0, i_13_251_2121_0,
    i_13_251_2137_0, i_13_251_2138_0, i_13_251_2165_0, i_13_251_2344_0,
    i_13_251_2360_0, i_13_251_2403_0, i_13_251_2452_0, i_13_251_2557_0,
    i_13_251_2559_0, i_13_251_2630_0, i_13_251_2647_0, i_13_251_2650_0,
    i_13_251_2719_0, i_13_251_2722_0, i_13_251_2749_0, i_13_251_2751_0,
    i_13_251_2821_0, i_13_251_2881_0, i_13_251_2896_0, i_13_251_2938_0,
    i_13_251_3019_0, i_13_251_3064_0, i_13_251_3205_0, i_13_251_3290_0,
    i_13_251_3325_0, i_13_251_3372_0, i_13_251_3430_0, i_13_251_3439_0,
    i_13_251_3520_0, i_13_251_3524_0, i_13_251_3525_0, i_13_251_3910_0,
    i_13_251_3919_0, i_13_251_3925_0, i_13_251_3926_0, i_13_251_3974_0,
    i_13_251_3987_0, i_13_251_3992_0, i_13_251_4032_0, i_13_251_4078_0,
    i_13_251_4183_0, i_13_251_4270_0, i_13_251_4294_0, i_13_251_4369_0,
    o_13_251_0_0  );
  input  i_13_251_37_0, i_13_251_38_0, i_13_251_51_0, i_13_251_75_0,
    i_13_251_76_0, i_13_251_103_0, i_13_251_112_0, i_13_251_165_0,
    i_13_251_173_0, i_13_251_181_0, i_13_251_184_0, i_13_251_240_0,
    i_13_251_252_0, i_13_251_280_0, i_13_251_281_0, i_13_251_324_0,
    i_13_251_325_0, i_13_251_339_0, i_13_251_571_0, i_13_251_577_0,
    i_13_251_596_0, i_13_251_597_0, i_13_251_598_0, i_13_251_618_0,
    i_13_251_640_0, i_13_251_643_0, i_13_251_685_0, i_13_251_715_0,
    i_13_251_744_0, i_13_251_778_0, i_13_251_814_0, i_13_251_840_0,
    i_13_251_891_0, i_13_251_892_0, i_13_251_894_0, i_13_251_896_0,
    i_13_251_1031_0, i_13_251_1093_0, i_13_251_1248_0, i_13_251_1249_0,
    i_13_251_1462_0, i_13_251_1480_0, i_13_251_1541_0, i_13_251_1711_0,
    i_13_251_1746_0, i_13_251_1747_0, i_13_251_1786_0, i_13_251_1804_0,
    i_13_251_1805_0, i_13_251_1806_0, i_13_251_1854_0, i_13_251_1855_0,
    i_13_251_1856_0, i_13_251_1858_0, i_13_251_2119_0, i_13_251_2121_0,
    i_13_251_2137_0, i_13_251_2138_0, i_13_251_2165_0, i_13_251_2344_0,
    i_13_251_2360_0, i_13_251_2403_0, i_13_251_2452_0, i_13_251_2557_0,
    i_13_251_2559_0, i_13_251_2630_0, i_13_251_2647_0, i_13_251_2650_0,
    i_13_251_2719_0, i_13_251_2722_0, i_13_251_2749_0, i_13_251_2751_0,
    i_13_251_2821_0, i_13_251_2881_0, i_13_251_2896_0, i_13_251_2938_0,
    i_13_251_3019_0, i_13_251_3064_0, i_13_251_3205_0, i_13_251_3290_0,
    i_13_251_3325_0, i_13_251_3372_0, i_13_251_3430_0, i_13_251_3439_0,
    i_13_251_3520_0, i_13_251_3524_0, i_13_251_3525_0, i_13_251_3910_0,
    i_13_251_3919_0, i_13_251_3925_0, i_13_251_3926_0, i_13_251_3974_0,
    i_13_251_3987_0, i_13_251_3992_0, i_13_251_4032_0, i_13_251_4078_0,
    i_13_251_4183_0, i_13_251_4270_0, i_13_251_4294_0, i_13_251_4369_0;
  output o_13_251_0_0;
  assign o_13_251_0_0 = ~((~i_13_251_618_0 & ((~i_13_251_184_0 & ~i_13_251_892_0) | (~i_13_251_894_0 & ~i_13_251_1747_0 & ~i_13_251_2138_0))) | (~i_13_251_3205_0 & ((~i_13_251_1806_0 & ~i_13_251_3064_0 & ~i_13_251_3524_0) | (i_13_251_3524_0 & ~i_13_251_3992_0))) | (i_13_251_618_0 & ~i_13_251_2137_0) | (~i_13_251_3910_0 & ~i_13_251_4032_0) | (~i_13_251_51_0 & ~i_13_251_2938_0 & ~i_13_251_4078_0) | (~i_13_251_571_0 & ~i_13_251_840_0 & ~i_13_251_4270_0));
endmodule



// Benchmark "kernel_13_252" written by ABC on Sun Jul 19 10:48:55 2020

module kernel_13_252 ( 
    i_13_252_37_0, i_13_252_49_0, i_13_252_100_0, i_13_252_127_0,
    i_13_252_136_0, i_13_252_154_0, i_13_252_166_0, i_13_252_167_0,
    i_13_252_269_0, i_13_252_271_0, i_13_252_280_0, i_13_252_283_0,
    i_13_252_316_0, i_13_252_379_0, i_13_252_385_0, i_13_252_386_0,
    i_13_252_415_0, i_13_252_450_0, i_13_252_451_0, i_13_252_558_0,
    i_13_252_571_0, i_13_252_639_0, i_13_252_640_0, i_13_252_658_0,
    i_13_252_676_0, i_13_252_677_0, i_13_252_720_0, i_13_252_758_0,
    i_13_252_869_0, i_13_252_940_0, i_13_252_982_0, i_13_252_1062_0,
    i_13_252_1063_0, i_13_252_1082_0, i_13_252_1093_0, i_13_252_1210_0,
    i_13_252_1300_0, i_13_252_1324_0, i_13_252_1390_0, i_13_252_1423_0,
    i_13_252_1436_0, i_13_252_1494_0, i_13_252_1525_0, i_13_252_1567_0,
    i_13_252_1633_0, i_13_252_1714_0, i_13_252_1807_0, i_13_252_1850_0,
    i_13_252_1909_0, i_13_252_1991_0, i_13_252_2054_0, i_13_252_2107_0,
    i_13_252_2108_0, i_13_252_2116_0, i_13_252_2233_0, i_13_252_2234_0,
    i_13_252_2297_0, i_13_252_2313_0, i_13_252_2361_0, i_13_252_2398_0,
    i_13_252_2467_0, i_13_252_2507_0, i_13_252_2542_0, i_13_252_2547_0,
    i_13_252_2663_0, i_13_252_2692_0, i_13_252_2766_0, i_13_252_2848_0,
    i_13_252_2872_0, i_13_252_3016_0, i_13_252_3106_0, i_13_252_3107_0,
    i_13_252_3109_0, i_13_252_3110_0, i_13_252_3307_0, i_13_252_3406_0,
    i_13_252_3433_0, i_13_252_3522_0, i_13_252_3528_0, i_13_252_3646_0,
    i_13_252_3708_0, i_13_252_3763_0, i_13_252_3766_0, i_13_252_3768_0,
    i_13_252_3817_0, i_13_252_3818_0, i_13_252_3901_0, i_13_252_4015_0,
    i_13_252_4078_0, i_13_252_4087_0, i_13_252_4117_0, i_13_252_4207_0,
    i_13_252_4230_0, i_13_252_4259_0, i_13_252_4266_0, i_13_252_4267_0,
    i_13_252_4302_0, i_13_252_4510_0, i_13_252_4555_0, i_13_252_4564_0,
    o_13_252_0_0  );
  input  i_13_252_37_0, i_13_252_49_0, i_13_252_100_0, i_13_252_127_0,
    i_13_252_136_0, i_13_252_154_0, i_13_252_166_0, i_13_252_167_0,
    i_13_252_269_0, i_13_252_271_0, i_13_252_280_0, i_13_252_283_0,
    i_13_252_316_0, i_13_252_379_0, i_13_252_385_0, i_13_252_386_0,
    i_13_252_415_0, i_13_252_450_0, i_13_252_451_0, i_13_252_558_0,
    i_13_252_571_0, i_13_252_639_0, i_13_252_640_0, i_13_252_658_0,
    i_13_252_676_0, i_13_252_677_0, i_13_252_720_0, i_13_252_758_0,
    i_13_252_869_0, i_13_252_940_0, i_13_252_982_0, i_13_252_1062_0,
    i_13_252_1063_0, i_13_252_1082_0, i_13_252_1093_0, i_13_252_1210_0,
    i_13_252_1300_0, i_13_252_1324_0, i_13_252_1390_0, i_13_252_1423_0,
    i_13_252_1436_0, i_13_252_1494_0, i_13_252_1525_0, i_13_252_1567_0,
    i_13_252_1633_0, i_13_252_1714_0, i_13_252_1807_0, i_13_252_1850_0,
    i_13_252_1909_0, i_13_252_1991_0, i_13_252_2054_0, i_13_252_2107_0,
    i_13_252_2108_0, i_13_252_2116_0, i_13_252_2233_0, i_13_252_2234_0,
    i_13_252_2297_0, i_13_252_2313_0, i_13_252_2361_0, i_13_252_2398_0,
    i_13_252_2467_0, i_13_252_2507_0, i_13_252_2542_0, i_13_252_2547_0,
    i_13_252_2663_0, i_13_252_2692_0, i_13_252_2766_0, i_13_252_2848_0,
    i_13_252_2872_0, i_13_252_3016_0, i_13_252_3106_0, i_13_252_3107_0,
    i_13_252_3109_0, i_13_252_3110_0, i_13_252_3307_0, i_13_252_3406_0,
    i_13_252_3433_0, i_13_252_3522_0, i_13_252_3528_0, i_13_252_3646_0,
    i_13_252_3708_0, i_13_252_3763_0, i_13_252_3766_0, i_13_252_3768_0,
    i_13_252_3817_0, i_13_252_3818_0, i_13_252_3901_0, i_13_252_4015_0,
    i_13_252_4078_0, i_13_252_4087_0, i_13_252_4117_0, i_13_252_4207_0,
    i_13_252_4230_0, i_13_252_4259_0, i_13_252_4266_0, i_13_252_4267_0,
    i_13_252_4302_0, i_13_252_4510_0, i_13_252_4555_0, i_13_252_4564_0;
  output o_13_252_0_0;
  assign o_13_252_0_0 = ~(~i_13_252_1324_0 | (i_13_252_2872_0 & ~i_13_252_4510_0) | (~i_13_252_2107_0 & i_13_252_3522_0) | (~i_13_252_100_0 & i_13_252_415_0 & ~i_13_252_4555_0) | (~i_13_252_3646_0 & ~i_13_252_3817_0 & ~i_13_252_3818_0));
endmodule



// Benchmark "kernel_13_253" written by ABC on Sun Jul 19 10:48:56 2020

module kernel_13_253 ( 
    i_13_253_93_0, i_13_253_94_0, i_13_253_112_0, i_13_253_121_0,
    i_13_253_165_0, i_13_253_192_0, i_13_253_193_0, i_13_253_199_0,
    i_13_253_225_0, i_13_253_504_0, i_13_253_531_0, i_13_253_570_0,
    i_13_253_571_0, i_13_253_588_0, i_13_253_639_0, i_13_253_714_0,
    i_13_253_715_0, i_13_253_729_0, i_13_253_814_0, i_13_253_891_0,
    i_13_253_927_0, i_13_253_948_0, i_13_253_999_0, i_13_253_1053_0,
    i_13_253_1200_0, i_13_253_1209_0, i_13_253_1210_0, i_13_253_1227_0,
    i_13_253_1317_0, i_13_253_1386_0, i_13_253_1407_0, i_13_253_1426_0,
    i_13_253_1467_0, i_13_253_1488_0, i_13_253_1512_0, i_13_253_1720_0,
    i_13_253_1764_0, i_13_253_1767_0, i_13_253_1782_0, i_13_253_1783_0,
    i_13_253_1785_0, i_13_253_1800_0, i_13_253_1801_0, i_13_253_1908_0,
    i_13_253_1990_0, i_13_253_1992_0, i_13_253_2011_0, i_13_253_2056_0,
    i_13_253_2109_0, i_13_253_2116_0, i_13_253_2128_0, i_13_253_2164_0,
    i_13_253_2206_0, i_13_253_2209_0, i_13_253_2225_0, i_13_253_2235_0,
    i_13_253_2452_0, i_13_253_2505_0, i_13_253_2532_0, i_13_253_2568_0,
    i_13_253_2623_0, i_13_253_2722_0, i_13_253_2875_0, i_13_253_2889_0,
    i_13_253_2934_0, i_13_253_3024_0, i_13_253_3046_0, i_13_253_3087_0,
    i_13_253_3154_0, i_13_253_3162_0, i_13_253_3163_0, i_13_253_3214_0,
    i_13_253_3286_0, i_13_253_3304_0, i_13_253_3375_0, i_13_253_3420_0,
    i_13_253_3421_0, i_13_253_3423_0, i_13_253_3451_0, i_13_253_3522_0,
    i_13_253_3753_0, i_13_253_3790_0, i_13_253_3873_0, i_13_253_3883_0,
    i_13_253_3918_0, i_13_253_3924_0, i_13_253_3981_0, i_13_253_4008_0,
    i_13_253_4009_0, i_13_253_4077_0, i_13_253_4167_0, i_13_253_4194_0,
    i_13_253_4212_0, i_13_253_4305_0, i_13_253_4320_0, i_13_253_4497_0,
    i_13_253_4530_0, i_13_253_4539_0, i_13_253_4584_0, i_13_253_4594_0,
    o_13_253_0_0  );
  input  i_13_253_93_0, i_13_253_94_0, i_13_253_112_0, i_13_253_121_0,
    i_13_253_165_0, i_13_253_192_0, i_13_253_193_0, i_13_253_199_0,
    i_13_253_225_0, i_13_253_504_0, i_13_253_531_0, i_13_253_570_0,
    i_13_253_571_0, i_13_253_588_0, i_13_253_639_0, i_13_253_714_0,
    i_13_253_715_0, i_13_253_729_0, i_13_253_814_0, i_13_253_891_0,
    i_13_253_927_0, i_13_253_948_0, i_13_253_999_0, i_13_253_1053_0,
    i_13_253_1200_0, i_13_253_1209_0, i_13_253_1210_0, i_13_253_1227_0,
    i_13_253_1317_0, i_13_253_1386_0, i_13_253_1407_0, i_13_253_1426_0,
    i_13_253_1467_0, i_13_253_1488_0, i_13_253_1512_0, i_13_253_1720_0,
    i_13_253_1764_0, i_13_253_1767_0, i_13_253_1782_0, i_13_253_1783_0,
    i_13_253_1785_0, i_13_253_1800_0, i_13_253_1801_0, i_13_253_1908_0,
    i_13_253_1990_0, i_13_253_1992_0, i_13_253_2011_0, i_13_253_2056_0,
    i_13_253_2109_0, i_13_253_2116_0, i_13_253_2128_0, i_13_253_2164_0,
    i_13_253_2206_0, i_13_253_2209_0, i_13_253_2225_0, i_13_253_2235_0,
    i_13_253_2452_0, i_13_253_2505_0, i_13_253_2532_0, i_13_253_2568_0,
    i_13_253_2623_0, i_13_253_2722_0, i_13_253_2875_0, i_13_253_2889_0,
    i_13_253_2934_0, i_13_253_3024_0, i_13_253_3046_0, i_13_253_3087_0,
    i_13_253_3154_0, i_13_253_3162_0, i_13_253_3163_0, i_13_253_3214_0,
    i_13_253_3286_0, i_13_253_3304_0, i_13_253_3375_0, i_13_253_3420_0,
    i_13_253_3421_0, i_13_253_3423_0, i_13_253_3451_0, i_13_253_3522_0,
    i_13_253_3753_0, i_13_253_3790_0, i_13_253_3873_0, i_13_253_3883_0,
    i_13_253_3918_0, i_13_253_3924_0, i_13_253_3981_0, i_13_253_4008_0,
    i_13_253_4009_0, i_13_253_4077_0, i_13_253_4167_0, i_13_253_4194_0,
    i_13_253_4212_0, i_13_253_4305_0, i_13_253_4320_0, i_13_253_4497_0,
    i_13_253_4530_0, i_13_253_4539_0, i_13_253_4584_0, i_13_253_4594_0;
  output o_13_253_0_0;
  assign o_13_253_0_0 = ~(i_13_253_1210_0 | (~i_13_253_1767_0 & ~i_13_253_4212_0 & i_13_253_4305_0) | (~i_13_253_927_0 & ~i_13_253_3420_0 & ~i_13_253_4008_0));
endmodule



// Benchmark "kernel_13_254" written by ABC on Sun Jul 19 10:48:57 2020

module kernel_13_254 ( 
    i_13_254_0_0, i_13_254_46_0, i_13_254_55_0, i_13_254_121_0,
    i_13_254_164_0, i_13_254_172_0, i_13_254_208_0, i_13_254_243_0,
    i_13_254_346_0, i_13_254_416_0, i_13_254_482_0, i_13_254_490_0,
    i_13_254_606_0, i_13_254_625_0, i_13_254_644_0, i_13_254_676_0,
    i_13_254_695_0, i_13_254_712_0, i_13_254_764_0, i_13_254_782_0,
    i_13_254_841_0, i_13_254_850_0, i_13_254_882_0, i_13_254_884_0,
    i_13_254_936_0, i_13_254_982_0, i_13_254_983_0, i_13_254_1242_0,
    i_13_254_1252_0, i_13_254_1263_0, i_13_254_1307_0, i_13_254_1484_0,
    i_13_254_1489_0, i_13_254_1507_0, i_13_254_1521_0, i_13_254_1525_0,
    i_13_254_1564_0, i_13_254_1570_0, i_13_254_1611_0, i_13_254_1643_0,
    i_13_254_1750_0, i_13_254_1751_0, i_13_254_1757_0, i_13_254_1841_0,
    i_13_254_1940_0, i_13_254_1943_0, i_13_254_1953_0, i_13_254_2024_0,
    i_13_254_2047_0, i_13_254_2097_0, i_13_254_2389_0, i_13_254_2443_0,
    i_13_254_2515_0, i_13_254_2539_0, i_13_254_2542_0, i_13_254_2605_0,
    i_13_254_2614_0, i_13_254_2692_0, i_13_254_2763_0, i_13_254_2782_0,
    i_13_254_2880_0, i_13_254_2963_0, i_13_254_3073_0, i_13_254_3077_0,
    i_13_254_3091_0, i_13_254_3106_0, i_13_254_3172_0, i_13_254_3261_0,
    i_13_254_3320_0, i_13_254_3352_0, i_13_254_3412_0, i_13_254_3566_0,
    i_13_254_3638_0, i_13_254_3657_0, i_13_254_3753_0, i_13_254_3781_0,
    i_13_254_3838_0, i_13_254_3845_0, i_13_254_3852_0, i_13_254_3865_0,
    i_13_254_3898_0, i_13_254_3983_0, i_13_254_3988_0, i_13_254_3991_0,
    i_13_254_3996_0, i_13_254_4036_0, i_13_254_4187_0, i_13_254_4214_0,
    i_13_254_4242_0, i_13_254_4270_0, i_13_254_4272_0, i_13_254_4295_0,
    i_13_254_4297_0, i_13_254_4307_0, i_13_254_4311_0, i_13_254_4375_0,
    i_13_254_4378_0, i_13_254_4511_0, i_13_254_4513_0, i_13_254_4603_0,
    o_13_254_0_0  );
  input  i_13_254_0_0, i_13_254_46_0, i_13_254_55_0, i_13_254_121_0,
    i_13_254_164_0, i_13_254_172_0, i_13_254_208_0, i_13_254_243_0,
    i_13_254_346_0, i_13_254_416_0, i_13_254_482_0, i_13_254_490_0,
    i_13_254_606_0, i_13_254_625_0, i_13_254_644_0, i_13_254_676_0,
    i_13_254_695_0, i_13_254_712_0, i_13_254_764_0, i_13_254_782_0,
    i_13_254_841_0, i_13_254_850_0, i_13_254_882_0, i_13_254_884_0,
    i_13_254_936_0, i_13_254_982_0, i_13_254_983_0, i_13_254_1242_0,
    i_13_254_1252_0, i_13_254_1263_0, i_13_254_1307_0, i_13_254_1484_0,
    i_13_254_1489_0, i_13_254_1507_0, i_13_254_1521_0, i_13_254_1525_0,
    i_13_254_1564_0, i_13_254_1570_0, i_13_254_1611_0, i_13_254_1643_0,
    i_13_254_1750_0, i_13_254_1751_0, i_13_254_1757_0, i_13_254_1841_0,
    i_13_254_1940_0, i_13_254_1943_0, i_13_254_1953_0, i_13_254_2024_0,
    i_13_254_2047_0, i_13_254_2097_0, i_13_254_2389_0, i_13_254_2443_0,
    i_13_254_2515_0, i_13_254_2539_0, i_13_254_2542_0, i_13_254_2605_0,
    i_13_254_2614_0, i_13_254_2692_0, i_13_254_2763_0, i_13_254_2782_0,
    i_13_254_2880_0, i_13_254_2963_0, i_13_254_3073_0, i_13_254_3077_0,
    i_13_254_3091_0, i_13_254_3106_0, i_13_254_3172_0, i_13_254_3261_0,
    i_13_254_3320_0, i_13_254_3352_0, i_13_254_3412_0, i_13_254_3566_0,
    i_13_254_3638_0, i_13_254_3657_0, i_13_254_3753_0, i_13_254_3781_0,
    i_13_254_3838_0, i_13_254_3845_0, i_13_254_3852_0, i_13_254_3865_0,
    i_13_254_3898_0, i_13_254_3983_0, i_13_254_3988_0, i_13_254_3991_0,
    i_13_254_3996_0, i_13_254_4036_0, i_13_254_4187_0, i_13_254_4214_0,
    i_13_254_4242_0, i_13_254_4270_0, i_13_254_4272_0, i_13_254_4295_0,
    i_13_254_4297_0, i_13_254_4307_0, i_13_254_4311_0, i_13_254_4375_0,
    i_13_254_4378_0, i_13_254_4511_0, i_13_254_4513_0, i_13_254_4603_0;
  output o_13_254_0_0;
  assign o_13_254_0_0 = 0;
endmodule



// Benchmark "kernel_13_255" written by ABC on Sun Jul 19 10:48:58 2020

module kernel_13_255 ( 
    i_13_255_0_0, i_13_255_1_0, i_13_255_136_0, i_13_255_298_0,
    i_13_255_326_0, i_13_255_364_0, i_13_255_544_0, i_13_255_550_0,
    i_13_255_568_0, i_13_255_625_0, i_13_255_626_0, i_13_255_712_0,
    i_13_255_730_0, i_13_255_847_0, i_13_255_850_0, i_13_255_901_0,
    i_13_255_941_0, i_13_255_1044_0, i_13_255_1125_0, i_13_255_1129_0,
    i_13_255_1225_0, i_13_255_1226_0, i_13_255_1252_0, i_13_255_1270_0,
    i_13_255_1279_0, i_13_255_1310_0, i_13_255_1480_0, i_13_255_1486_0,
    i_13_255_1522_0, i_13_255_1552_0, i_13_255_1584_0, i_13_255_1585_0,
    i_13_255_1604_0, i_13_255_1749_0, i_13_255_1765_0, i_13_255_1810_0,
    i_13_255_1828_0, i_13_255_1854_0, i_13_255_1891_0, i_13_255_2020_0,
    i_13_255_2098_0, i_13_255_2116_0, i_13_255_2119_0, i_13_255_2214_0,
    i_13_255_2395_0, i_13_255_2422_0, i_13_255_2566_0, i_13_255_2593_0,
    i_13_255_2642_0, i_13_255_2647_0, i_13_255_2740_0, i_13_255_2755_0,
    i_13_255_2803_0, i_13_255_2875_0, i_13_255_2876_0, i_13_255_2917_0,
    i_13_255_2971_0, i_13_255_2972_0, i_13_255_2974_0, i_13_255_3019_0,
    i_13_255_3044_0, i_13_255_3091_0, i_13_255_3100_0, i_13_255_3101_0,
    i_13_255_3115_0, i_13_255_3127_0, i_13_255_3133_0, i_13_255_3145_0,
    i_13_255_3190_0, i_13_255_3213_0, i_13_255_3214_0, i_13_255_3262_0,
    i_13_255_3304_0, i_13_255_3331_0, i_13_255_3380_0, i_13_255_3416_0,
    i_13_255_3460_0, i_13_255_3485_0, i_13_255_3573_0, i_13_255_3822_0,
    i_13_255_3853_0, i_13_255_3899_0, i_13_255_3916_0, i_13_255_3944_0,
    i_13_255_3964_0, i_13_255_3979_0, i_13_255_3981_0, i_13_255_4033_0,
    i_13_255_4078_0, i_13_255_4091_0, i_13_255_4160_0, i_13_255_4266_0,
    i_13_255_4270_0, i_13_255_4303_0, i_13_255_4320_0, i_13_255_4325_0,
    i_13_255_4460_0, i_13_255_4475_0, i_13_255_4504_0, i_13_255_4529_0,
    o_13_255_0_0  );
  input  i_13_255_0_0, i_13_255_1_0, i_13_255_136_0, i_13_255_298_0,
    i_13_255_326_0, i_13_255_364_0, i_13_255_544_0, i_13_255_550_0,
    i_13_255_568_0, i_13_255_625_0, i_13_255_626_0, i_13_255_712_0,
    i_13_255_730_0, i_13_255_847_0, i_13_255_850_0, i_13_255_901_0,
    i_13_255_941_0, i_13_255_1044_0, i_13_255_1125_0, i_13_255_1129_0,
    i_13_255_1225_0, i_13_255_1226_0, i_13_255_1252_0, i_13_255_1270_0,
    i_13_255_1279_0, i_13_255_1310_0, i_13_255_1480_0, i_13_255_1486_0,
    i_13_255_1522_0, i_13_255_1552_0, i_13_255_1584_0, i_13_255_1585_0,
    i_13_255_1604_0, i_13_255_1749_0, i_13_255_1765_0, i_13_255_1810_0,
    i_13_255_1828_0, i_13_255_1854_0, i_13_255_1891_0, i_13_255_2020_0,
    i_13_255_2098_0, i_13_255_2116_0, i_13_255_2119_0, i_13_255_2214_0,
    i_13_255_2395_0, i_13_255_2422_0, i_13_255_2566_0, i_13_255_2593_0,
    i_13_255_2642_0, i_13_255_2647_0, i_13_255_2740_0, i_13_255_2755_0,
    i_13_255_2803_0, i_13_255_2875_0, i_13_255_2876_0, i_13_255_2917_0,
    i_13_255_2971_0, i_13_255_2972_0, i_13_255_2974_0, i_13_255_3019_0,
    i_13_255_3044_0, i_13_255_3091_0, i_13_255_3100_0, i_13_255_3101_0,
    i_13_255_3115_0, i_13_255_3127_0, i_13_255_3133_0, i_13_255_3145_0,
    i_13_255_3190_0, i_13_255_3213_0, i_13_255_3214_0, i_13_255_3262_0,
    i_13_255_3304_0, i_13_255_3331_0, i_13_255_3380_0, i_13_255_3416_0,
    i_13_255_3460_0, i_13_255_3485_0, i_13_255_3573_0, i_13_255_3822_0,
    i_13_255_3853_0, i_13_255_3899_0, i_13_255_3916_0, i_13_255_3944_0,
    i_13_255_3964_0, i_13_255_3979_0, i_13_255_3981_0, i_13_255_4033_0,
    i_13_255_4078_0, i_13_255_4091_0, i_13_255_4160_0, i_13_255_4266_0,
    i_13_255_4270_0, i_13_255_4303_0, i_13_255_4320_0, i_13_255_4325_0,
    i_13_255_4460_0, i_13_255_4475_0, i_13_255_4504_0, i_13_255_4529_0;
  output o_13_255_0_0;
  assign o_13_255_0_0 = 0;
endmodule



// Benchmark "kernel_13_256" written by ABC on Sun Jul 19 10:48:59 2020

module kernel_13_256 ( 
    i_13_256_27_0, i_13_256_30_0, i_13_256_63_0, i_13_256_64_0,
    i_13_256_130_0, i_13_256_135_0, i_13_256_136_0, i_13_256_156_0,
    i_13_256_202_0, i_13_256_207_0, i_13_256_208_0, i_13_256_225_0,
    i_13_256_354_0, i_13_256_355_0, i_13_256_378_0, i_13_256_453_0,
    i_13_256_454_0, i_13_256_468_0, i_13_256_469_0, i_13_256_489_0,
    i_13_256_549_0, i_13_256_612_0, i_13_256_643_0, i_13_256_675_0,
    i_13_256_730_0, i_13_256_732_0, i_13_256_793_0, i_13_256_796_0,
    i_13_256_810_0, i_13_256_831_0, i_13_256_840_0, i_13_256_946_0,
    i_13_256_954_0, i_13_256_1021_0, i_13_256_1063_0, i_13_256_1120_0,
    i_13_256_1128_0, i_13_256_1273_0, i_13_256_1300_0, i_13_256_1344_0,
    i_13_256_1486_0, i_13_256_1522_0, i_13_256_1525_0, i_13_256_1620_0,
    i_13_256_1621_0, i_13_256_1677_0, i_13_256_1692_0, i_13_256_1696_0,
    i_13_256_1719_0, i_13_256_1720_0, i_13_256_1836_0, i_13_256_1846_0,
    i_13_256_2002_0, i_13_256_2100_0, i_13_256_2173_0, i_13_256_2296_0,
    i_13_256_2316_0, i_13_256_2340_0, i_13_256_2341_0, i_13_256_2421_0,
    i_13_256_2431_0, i_13_256_2538_0, i_13_256_2550_0, i_13_256_2676_0,
    i_13_256_2677_0, i_13_256_2694_0, i_13_256_2718_0, i_13_256_2719_0,
    i_13_256_2748_0, i_13_256_2880_0, i_13_256_2946_0, i_13_256_3033_0,
    i_13_256_3072_0, i_13_256_3109_0, i_13_256_3231_0, i_13_256_3241_0,
    i_13_256_3421_0, i_13_256_3466_0, i_13_256_3528_0, i_13_256_3594_0,
    i_13_256_3610_0, i_13_256_3618_0, i_13_256_3619_0, i_13_256_3636_0,
    i_13_256_3637_0, i_13_256_3666_0, i_13_256_3681_0, i_13_256_3726_0,
    i_13_256_3843_0, i_13_256_3982_0, i_13_256_4233_0, i_13_256_4261_0,
    i_13_256_4269_0, i_13_256_4279_0, i_13_256_4315_0, i_13_256_4329_0,
    i_13_256_4396_0, i_13_256_4509_0, i_13_256_4519_0, i_13_256_4537_0,
    o_13_256_0_0  );
  input  i_13_256_27_0, i_13_256_30_0, i_13_256_63_0, i_13_256_64_0,
    i_13_256_130_0, i_13_256_135_0, i_13_256_136_0, i_13_256_156_0,
    i_13_256_202_0, i_13_256_207_0, i_13_256_208_0, i_13_256_225_0,
    i_13_256_354_0, i_13_256_355_0, i_13_256_378_0, i_13_256_453_0,
    i_13_256_454_0, i_13_256_468_0, i_13_256_469_0, i_13_256_489_0,
    i_13_256_549_0, i_13_256_612_0, i_13_256_643_0, i_13_256_675_0,
    i_13_256_730_0, i_13_256_732_0, i_13_256_793_0, i_13_256_796_0,
    i_13_256_810_0, i_13_256_831_0, i_13_256_840_0, i_13_256_946_0,
    i_13_256_954_0, i_13_256_1021_0, i_13_256_1063_0, i_13_256_1120_0,
    i_13_256_1128_0, i_13_256_1273_0, i_13_256_1300_0, i_13_256_1344_0,
    i_13_256_1486_0, i_13_256_1522_0, i_13_256_1525_0, i_13_256_1620_0,
    i_13_256_1621_0, i_13_256_1677_0, i_13_256_1692_0, i_13_256_1696_0,
    i_13_256_1719_0, i_13_256_1720_0, i_13_256_1836_0, i_13_256_1846_0,
    i_13_256_2002_0, i_13_256_2100_0, i_13_256_2173_0, i_13_256_2296_0,
    i_13_256_2316_0, i_13_256_2340_0, i_13_256_2341_0, i_13_256_2421_0,
    i_13_256_2431_0, i_13_256_2538_0, i_13_256_2550_0, i_13_256_2676_0,
    i_13_256_2677_0, i_13_256_2694_0, i_13_256_2718_0, i_13_256_2719_0,
    i_13_256_2748_0, i_13_256_2880_0, i_13_256_2946_0, i_13_256_3033_0,
    i_13_256_3072_0, i_13_256_3109_0, i_13_256_3231_0, i_13_256_3241_0,
    i_13_256_3421_0, i_13_256_3466_0, i_13_256_3528_0, i_13_256_3594_0,
    i_13_256_3610_0, i_13_256_3618_0, i_13_256_3619_0, i_13_256_3636_0,
    i_13_256_3637_0, i_13_256_3666_0, i_13_256_3681_0, i_13_256_3726_0,
    i_13_256_3843_0, i_13_256_3982_0, i_13_256_4233_0, i_13_256_4261_0,
    i_13_256_4269_0, i_13_256_4279_0, i_13_256_4315_0, i_13_256_4329_0,
    i_13_256_4396_0, i_13_256_4509_0, i_13_256_4519_0, i_13_256_4537_0;
  output o_13_256_0_0;
  assign o_13_256_0_0 = ~(~i_13_256_468_0 & ~i_13_256_1836_0);
endmodule



// Benchmark "kernel_13_257" written by ABC on Sun Jul 19 10:49:00 2020

module kernel_13_257 ( 
    i_13_257_171_0, i_13_257_172_0, i_13_257_174_0, i_13_257_175_0,
    i_13_257_279_0, i_13_257_280_0, i_13_257_283_0, i_13_257_465_0,
    i_13_257_472_0, i_13_257_523_0, i_13_257_525_0, i_13_257_562_0,
    i_13_257_612_0, i_13_257_657_0, i_13_257_661_0, i_13_257_793_0,
    i_13_257_820_0, i_13_257_822_0, i_13_257_823_0, i_13_257_847_0,
    i_13_257_849_0, i_13_257_1017_0, i_13_257_1071_0, i_13_257_1072_0,
    i_13_257_1224_0, i_13_257_1225_0, i_13_257_1227_0, i_13_257_1308_0,
    i_13_257_1309_0, i_13_257_1363_0, i_13_257_1422_0, i_13_257_1425_0,
    i_13_257_1485_0, i_13_257_1489_0, i_13_257_1494_0, i_13_257_1495_0,
    i_13_257_1549_0, i_13_257_1629_0, i_13_257_1641_0, i_13_257_1855_0,
    i_13_257_1858_0, i_13_257_1881_0, i_13_257_1999_0, i_13_257_2070_0,
    i_13_257_2190_0, i_13_257_2206_0, i_13_257_2314_0, i_13_257_2347_0,
    i_13_257_2422_0, i_13_257_2448_0, i_13_257_2449_0, i_13_257_2539_0,
    i_13_257_2658_0, i_13_257_2673_0, i_13_257_2676_0, i_13_257_2692_0,
    i_13_257_2746_0, i_13_257_3007_0, i_13_257_3009_0, i_13_257_3096_0,
    i_13_257_3133_0, i_13_257_3216_0, i_13_257_3235_0, i_13_257_3267_0,
    i_13_257_3268_0, i_13_257_3270_0, i_13_257_3271_0, i_13_257_3414_0,
    i_13_257_3420_0, i_13_257_3421_0, i_13_257_3423_0, i_13_257_3523_0,
    i_13_257_3537_0, i_13_257_3538_0, i_13_257_3540_0, i_13_257_3643_0,
    i_13_257_3730_0, i_13_257_3741_0, i_13_257_3781_0, i_13_257_3798_0,
    i_13_257_3834_0, i_13_257_4015_0, i_13_257_4080_0, i_13_257_4195_0,
    i_13_257_4248_0, i_13_257_4249_0, i_13_257_4251_0, i_13_257_4252_0,
    i_13_257_4257_0, i_13_257_4258_0, i_13_257_4260_0, i_13_257_4275_0,
    i_13_257_4293_0, i_13_257_4338_0, i_13_257_4351_0, i_13_257_4375_0,
    i_13_257_4381_0, i_13_257_4414_0, i_13_257_4494_0, i_13_257_4555_0,
    o_13_257_0_0  );
  input  i_13_257_171_0, i_13_257_172_0, i_13_257_174_0, i_13_257_175_0,
    i_13_257_279_0, i_13_257_280_0, i_13_257_283_0, i_13_257_465_0,
    i_13_257_472_0, i_13_257_523_0, i_13_257_525_0, i_13_257_562_0,
    i_13_257_612_0, i_13_257_657_0, i_13_257_661_0, i_13_257_793_0,
    i_13_257_820_0, i_13_257_822_0, i_13_257_823_0, i_13_257_847_0,
    i_13_257_849_0, i_13_257_1017_0, i_13_257_1071_0, i_13_257_1072_0,
    i_13_257_1224_0, i_13_257_1225_0, i_13_257_1227_0, i_13_257_1308_0,
    i_13_257_1309_0, i_13_257_1363_0, i_13_257_1422_0, i_13_257_1425_0,
    i_13_257_1485_0, i_13_257_1489_0, i_13_257_1494_0, i_13_257_1495_0,
    i_13_257_1549_0, i_13_257_1629_0, i_13_257_1641_0, i_13_257_1855_0,
    i_13_257_1858_0, i_13_257_1881_0, i_13_257_1999_0, i_13_257_2070_0,
    i_13_257_2190_0, i_13_257_2206_0, i_13_257_2314_0, i_13_257_2347_0,
    i_13_257_2422_0, i_13_257_2448_0, i_13_257_2449_0, i_13_257_2539_0,
    i_13_257_2658_0, i_13_257_2673_0, i_13_257_2676_0, i_13_257_2692_0,
    i_13_257_2746_0, i_13_257_3007_0, i_13_257_3009_0, i_13_257_3096_0,
    i_13_257_3133_0, i_13_257_3216_0, i_13_257_3235_0, i_13_257_3267_0,
    i_13_257_3268_0, i_13_257_3270_0, i_13_257_3271_0, i_13_257_3414_0,
    i_13_257_3420_0, i_13_257_3421_0, i_13_257_3423_0, i_13_257_3523_0,
    i_13_257_3537_0, i_13_257_3538_0, i_13_257_3540_0, i_13_257_3643_0,
    i_13_257_3730_0, i_13_257_3741_0, i_13_257_3781_0, i_13_257_3798_0,
    i_13_257_3834_0, i_13_257_4015_0, i_13_257_4080_0, i_13_257_4195_0,
    i_13_257_4248_0, i_13_257_4249_0, i_13_257_4251_0, i_13_257_4252_0,
    i_13_257_4257_0, i_13_257_4258_0, i_13_257_4260_0, i_13_257_4275_0,
    i_13_257_4293_0, i_13_257_4338_0, i_13_257_4351_0, i_13_257_4375_0,
    i_13_257_4381_0, i_13_257_4414_0, i_13_257_4494_0, i_13_257_4555_0;
  output o_13_257_0_0;
  assign o_13_257_0_0 = ~(~i_13_257_1549_0 | (~i_13_257_2206_0 & ~i_13_257_4252_0) | (~i_13_257_2449_0 & ~i_13_257_3423_0) | (~i_13_257_2448_0 & ~i_13_257_4251_0 & ~i_13_257_4414_0) | (~i_13_257_1858_0 & ~i_13_257_3540_0 & ~i_13_257_4257_0));
endmodule



// Benchmark "kernel_13_258" written by ABC on Sun Jul 19 10:49:00 2020

module kernel_13_258 ( 
    i_13_258_105_0, i_13_258_106_0, i_13_258_213_0, i_13_258_420_0,
    i_13_258_600_0, i_13_258_609_0, i_13_258_619_0, i_13_258_742_0,
    i_13_258_745_0, i_13_258_858_0, i_13_258_1024_0, i_13_258_1068_0,
    i_13_258_1069_0, i_13_258_1086_0, i_13_258_1087_0, i_13_258_1095_0,
    i_13_258_1347_0, i_13_258_1488_0, i_13_258_1500_0, i_13_258_1507_0,
    i_13_258_1518_0, i_13_258_1519_0, i_13_258_1536_0, i_13_258_1561_0,
    i_13_258_1570_0, i_13_258_1572_0, i_13_258_1795_0, i_13_258_1813_0,
    i_13_258_1860_0, i_13_258_1930_0, i_13_258_2058_0, i_13_258_2059_0,
    i_13_258_2095_0, i_13_258_2149_0, i_13_258_2265_0, i_13_258_2280_0,
    i_13_258_2380_0, i_13_258_2400_0, i_13_258_2496_0, i_13_258_2500_0,
    i_13_258_2541_0, i_13_258_2551_0, i_13_258_2598_0, i_13_258_2599_0,
    i_13_258_2617_0, i_13_258_2679_0, i_13_258_2707_0, i_13_258_2715_0,
    i_13_258_2751_0, i_13_258_2851_0, i_13_258_2938_0, i_13_258_2985_0,
    i_13_258_2986_0, i_13_258_3012_0, i_13_258_3019_0, i_13_258_3031_0,
    i_13_258_3067_0, i_13_258_3073_0, i_13_258_3147_0, i_13_258_3148_0,
    i_13_258_3210_0, i_13_258_3211_0, i_13_258_3217_0, i_13_258_3328_0,
    i_13_258_3343_0, i_13_258_3346_0, i_13_258_3388_0, i_13_258_3400_0,
    i_13_258_3417_0, i_13_258_3418_0, i_13_258_3453_0, i_13_258_3454_0,
    i_13_258_3478_0, i_13_258_3525_0, i_13_258_3526_0, i_13_258_3531_0,
    i_13_258_3532_0, i_13_258_3732_0, i_13_258_3769_0, i_13_258_3891_0,
    i_13_258_4020_0, i_13_258_4039_0, i_13_258_4047_0, i_13_258_4048_0,
    i_13_258_4093_0, i_13_258_4119_0, i_13_258_4120_0, i_13_258_4234_0,
    i_13_258_4236_0, i_13_258_4254_0, i_13_258_4270_0, i_13_258_4317_0,
    i_13_258_4327_0, i_13_258_4353_0, i_13_258_4396_0, i_13_258_4416_0,
    i_13_258_4417_0, i_13_258_4476_0, i_13_258_4543_0, i_13_258_4557_0,
    o_13_258_0_0  );
  input  i_13_258_105_0, i_13_258_106_0, i_13_258_213_0, i_13_258_420_0,
    i_13_258_600_0, i_13_258_609_0, i_13_258_619_0, i_13_258_742_0,
    i_13_258_745_0, i_13_258_858_0, i_13_258_1024_0, i_13_258_1068_0,
    i_13_258_1069_0, i_13_258_1086_0, i_13_258_1087_0, i_13_258_1095_0,
    i_13_258_1347_0, i_13_258_1488_0, i_13_258_1500_0, i_13_258_1507_0,
    i_13_258_1518_0, i_13_258_1519_0, i_13_258_1536_0, i_13_258_1561_0,
    i_13_258_1570_0, i_13_258_1572_0, i_13_258_1795_0, i_13_258_1813_0,
    i_13_258_1860_0, i_13_258_1930_0, i_13_258_2058_0, i_13_258_2059_0,
    i_13_258_2095_0, i_13_258_2149_0, i_13_258_2265_0, i_13_258_2280_0,
    i_13_258_2380_0, i_13_258_2400_0, i_13_258_2496_0, i_13_258_2500_0,
    i_13_258_2541_0, i_13_258_2551_0, i_13_258_2598_0, i_13_258_2599_0,
    i_13_258_2617_0, i_13_258_2679_0, i_13_258_2707_0, i_13_258_2715_0,
    i_13_258_2751_0, i_13_258_2851_0, i_13_258_2938_0, i_13_258_2985_0,
    i_13_258_2986_0, i_13_258_3012_0, i_13_258_3019_0, i_13_258_3031_0,
    i_13_258_3067_0, i_13_258_3073_0, i_13_258_3147_0, i_13_258_3148_0,
    i_13_258_3210_0, i_13_258_3211_0, i_13_258_3217_0, i_13_258_3328_0,
    i_13_258_3343_0, i_13_258_3346_0, i_13_258_3388_0, i_13_258_3400_0,
    i_13_258_3417_0, i_13_258_3418_0, i_13_258_3453_0, i_13_258_3454_0,
    i_13_258_3478_0, i_13_258_3525_0, i_13_258_3526_0, i_13_258_3531_0,
    i_13_258_3532_0, i_13_258_3732_0, i_13_258_3769_0, i_13_258_3891_0,
    i_13_258_4020_0, i_13_258_4039_0, i_13_258_4047_0, i_13_258_4048_0,
    i_13_258_4093_0, i_13_258_4119_0, i_13_258_4120_0, i_13_258_4234_0,
    i_13_258_4236_0, i_13_258_4254_0, i_13_258_4270_0, i_13_258_4317_0,
    i_13_258_4327_0, i_13_258_4353_0, i_13_258_4396_0, i_13_258_4416_0,
    i_13_258_4417_0, i_13_258_4476_0, i_13_258_4543_0, i_13_258_4557_0;
  output o_13_258_0_0;
  assign o_13_258_0_0 = ~((~i_13_258_1087_0 & ((~i_13_258_1068_0 & i_13_258_2851_0 & ~i_13_258_3453_0) | (~i_13_258_1860_0 & ~i_13_258_2715_0 & ~i_13_258_2986_0 & ~i_13_258_4236_0))) | (i_13_258_3343_0 & (~i_13_258_4417_0 | (i_13_258_2149_0 & ~i_13_258_4236_0))) | (~i_13_258_4236_0 & ((~i_13_258_2986_0 & ~i_13_258_3400_0) | (~i_13_258_1488_0 & ~i_13_258_3067_0 & ~i_13_258_3769_0))) | (~i_13_258_1069_0 & ~i_13_258_2851_0 & ~i_13_258_3147_0) | (~i_13_258_858_0 & i_13_258_4234_0) | (i_13_258_3388_0 & ~i_13_258_4416_0));
endmodule



// Benchmark "kernel_13_259" written by ABC on Sun Jul 19 10:49:01 2020

module kernel_13_259 ( 
    i_13_259_49_0, i_13_259_64_0, i_13_259_118_0, i_13_259_166_0,
    i_13_259_233_0, i_13_259_238_0, i_13_259_308_0, i_13_259_311_0,
    i_13_259_317_0, i_13_259_328_0, i_13_259_569_0, i_13_259_586_0,
    i_13_259_587_0, i_13_259_640_0, i_13_259_641_0, i_13_259_712_0,
    i_13_259_739_0, i_13_259_740_0, i_13_259_757_0, i_13_259_838_0,
    i_13_259_839_0, i_13_259_856_0, i_13_259_929_0, i_13_259_1017_0,
    i_13_259_1082_0, i_13_259_1201_0, i_13_259_1253_0, i_13_259_1324_0,
    i_13_259_1325_0, i_13_259_1350_0, i_13_259_1442_0, i_13_259_1468_0,
    i_13_259_1486_0, i_13_259_1505_0, i_13_259_1526_0, i_13_259_1550_0,
    i_13_259_1568_0, i_13_259_1830_0, i_13_259_1832_0, i_13_259_1908_0,
    i_13_259_1990_0, i_13_259_2002_0, i_13_259_2045_0, i_13_259_2053_0,
    i_13_259_2054_0, i_13_259_2056_0, i_13_259_2108_0, i_13_259_2117_0,
    i_13_259_2234_0, i_13_259_2245_0, i_13_259_2259_0, i_13_259_2260_0,
    i_13_259_2261_0, i_13_259_2263_0, i_13_259_2264_0, i_13_259_2277_0,
    i_13_259_2278_0, i_13_259_2279_0, i_13_259_2407_0, i_13_259_2709_0,
    i_13_259_2711_0, i_13_259_2722_0, i_13_259_2750_0, i_13_259_2855_0,
    i_13_259_2945_0, i_13_259_3037_0, i_13_259_3061_0, i_13_259_3064_0,
    i_13_259_3065_0, i_13_259_3109_0, i_13_259_3110_0, i_13_259_3288_0,
    i_13_259_3388_0, i_13_259_3438_0, i_13_259_3439_0, i_13_259_3476_0,
    i_13_259_3483_0, i_13_259_3611_0, i_13_259_3614_0, i_13_259_3688_0,
    i_13_259_3703_0, i_13_259_3757_0, i_13_259_3766_0, i_13_259_3817_0,
    i_13_259_3818_0, i_13_259_3901_0, i_13_259_3928_0, i_13_259_3993_0,
    i_13_259_4007_0, i_13_259_4033_0, i_13_259_4186_0, i_13_259_4187_0,
    i_13_259_4276_0, i_13_259_4303_0, i_13_259_4304_0, i_13_259_4306_0,
    i_13_259_4315_0, i_13_259_4339_0, i_13_259_4394_0, i_13_259_4601_0,
    o_13_259_0_0  );
  input  i_13_259_49_0, i_13_259_64_0, i_13_259_118_0, i_13_259_166_0,
    i_13_259_233_0, i_13_259_238_0, i_13_259_308_0, i_13_259_311_0,
    i_13_259_317_0, i_13_259_328_0, i_13_259_569_0, i_13_259_586_0,
    i_13_259_587_0, i_13_259_640_0, i_13_259_641_0, i_13_259_712_0,
    i_13_259_739_0, i_13_259_740_0, i_13_259_757_0, i_13_259_838_0,
    i_13_259_839_0, i_13_259_856_0, i_13_259_929_0, i_13_259_1017_0,
    i_13_259_1082_0, i_13_259_1201_0, i_13_259_1253_0, i_13_259_1324_0,
    i_13_259_1325_0, i_13_259_1350_0, i_13_259_1442_0, i_13_259_1468_0,
    i_13_259_1486_0, i_13_259_1505_0, i_13_259_1526_0, i_13_259_1550_0,
    i_13_259_1568_0, i_13_259_1830_0, i_13_259_1832_0, i_13_259_1908_0,
    i_13_259_1990_0, i_13_259_2002_0, i_13_259_2045_0, i_13_259_2053_0,
    i_13_259_2054_0, i_13_259_2056_0, i_13_259_2108_0, i_13_259_2117_0,
    i_13_259_2234_0, i_13_259_2245_0, i_13_259_2259_0, i_13_259_2260_0,
    i_13_259_2261_0, i_13_259_2263_0, i_13_259_2264_0, i_13_259_2277_0,
    i_13_259_2278_0, i_13_259_2279_0, i_13_259_2407_0, i_13_259_2709_0,
    i_13_259_2711_0, i_13_259_2722_0, i_13_259_2750_0, i_13_259_2855_0,
    i_13_259_2945_0, i_13_259_3037_0, i_13_259_3061_0, i_13_259_3064_0,
    i_13_259_3065_0, i_13_259_3109_0, i_13_259_3110_0, i_13_259_3288_0,
    i_13_259_3388_0, i_13_259_3438_0, i_13_259_3439_0, i_13_259_3476_0,
    i_13_259_3483_0, i_13_259_3611_0, i_13_259_3614_0, i_13_259_3688_0,
    i_13_259_3703_0, i_13_259_3757_0, i_13_259_3766_0, i_13_259_3817_0,
    i_13_259_3818_0, i_13_259_3901_0, i_13_259_3928_0, i_13_259_3993_0,
    i_13_259_4007_0, i_13_259_4033_0, i_13_259_4186_0, i_13_259_4187_0,
    i_13_259_4276_0, i_13_259_4303_0, i_13_259_4304_0, i_13_259_4306_0,
    i_13_259_4315_0, i_13_259_4339_0, i_13_259_4394_0, i_13_259_4601_0;
  output o_13_259_0_0;
  assign o_13_259_0_0 = ~((~i_13_259_2054_0 & ((i_13_259_2234_0 & ~i_13_259_2711_0) | (~i_13_259_2855_0 & ~i_13_259_3928_0 & i_13_259_4033_0 & ~i_13_259_4187_0))) | (~i_13_259_4394_0 & ((~i_13_259_757_0 & ~i_13_259_3064_0) | (~i_13_259_3061_0 & ~i_13_259_3818_0))) | (~i_13_259_3064_0 & ~i_13_259_3818_0 & (i_13_259_118_0 | ~i_13_259_2002_0)) | (~i_13_259_49_0 & ~i_13_259_2278_0 & ~i_13_259_2279_0) | (~i_13_259_2056_0 & ~i_13_259_3614_0 & ~i_13_259_3817_0));
endmodule



// Benchmark "kernel_13_260" written by ABC on Sun Jul 19 10:49:02 2020

module kernel_13_260 ( 
    i_13_260_20_0, i_13_260_39_0, i_13_260_64_0, i_13_260_65_0,
    i_13_260_73_0, i_13_260_173_0, i_13_260_356_0, i_13_260_357_0,
    i_13_260_379_0, i_13_260_406_0, i_13_260_443_0, i_13_260_469_0,
    i_13_260_526_0, i_13_260_527_0, i_13_260_530_0, i_13_260_667_0,
    i_13_260_668_0, i_13_260_676_0, i_13_260_677_0, i_13_260_695_0,
    i_13_260_700_0, i_13_260_758_0, i_13_260_829_0, i_13_260_830_0,
    i_13_260_838_0, i_13_260_839_0, i_13_260_853_0, i_13_260_854_0,
    i_13_260_947_0, i_13_260_949_0, i_13_260_950_0, i_13_260_1024_0,
    i_13_260_1099_0, i_13_260_1118_0, i_13_260_1397_0, i_13_260_1438_0,
    i_13_260_1487_0, i_13_260_1499_0, i_13_260_1505_0, i_13_260_1594_0,
    i_13_260_1658_0, i_13_260_1720_0, i_13_260_1742_0, i_13_260_1744_0,
    i_13_260_1751_0, i_13_260_1792_0, i_13_260_1883_0, i_13_260_1913_0,
    i_13_260_1928_0, i_13_260_1950_0, i_13_260_2030_0, i_13_260_2032_0,
    i_13_260_2224_0, i_13_260_2242_0, i_13_260_2341_0, i_13_260_2454_0,
    i_13_260_2467_0, i_13_260_2468_0, i_13_260_2512_0, i_13_260_2514_0,
    i_13_260_2692_0, i_13_260_2693_0, i_13_260_2720_0, i_13_260_2750_0,
    i_13_260_2764_0, i_13_260_2912_0, i_13_260_3010_0, i_13_260_3026_0,
    i_13_260_3044_0, i_13_260_3061_0, i_13_260_3062_0, i_13_260_3128_0,
    i_13_260_3134_0, i_13_260_3146_0, i_13_260_3370_0, i_13_260_3371_0,
    i_13_260_3373_0, i_13_260_3382_0, i_13_260_3533_0, i_13_260_3596_0,
    i_13_260_3597_0, i_13_260_3598_0, i_13_260_3620_0, i_13_260_3632_0,
    i_13_260_3633_0, i_13_260_3638_0, i_13_260_3733_0, i_13_260_3783_0,
    i_13_260_3860_0, i_13_260_3925_0, i_13_260_3926_0, i_13_260_3988_0,
    i_13_260_4264_0, i_13_260_4312_0, i_13_260_4330_0, i_13_260_4331_0,
    i_13_260_4332_0, i_13_260_4414_0, i_13_260_4430_0, i_13_260_4451_0,
    o_13_260_0_0  );
  input  i_13_260_20_0, i_13_260_39_0, i_13_260_64_0, i_13_260_65_0,
    i_13_260_73_0, i_13_260_173_0, i_13_260_356_0, i_13_260_357_0,
    i_13_260_379_0, i_13_260_406_0, i_13_260_443_0, i_13_260_469_0,
    i_13_260_526_0, i_13_260_527_0, i_13_260_530_0, i_13_260_667_0,
    i_13_260_668_0, i_13_260_676_0, i_13_260_677_0, i_13_260_695_0,
    i_13_260_700_0, i_13_260_758_0, i_13_260_829_0, i_13_260_830_0,
    i_13_260_838_0, i_13_260_839_0, i_13_260_853_0, i_13_260_854_0,
    i_13_260_947_0, i_13_260_949_0, i_13_260_950_0, i_13_260_1024_0,
    i_13_260_1099_0, i_13_260_1118_0, i_13_260_1397_0, i_13_260_1438_0,
    i_13_260_1487_0, i_13_260_1499_0, i_13_260_1505_0, i_13_260_1594_0,
    i_13_260_1658_0, i_13_260_1720_0, i_13_260_1742_0, i_13_260_1744_0,
    i_13_260_1751_0, i_13_260_1792_0, i_13_260_1883_0, i_13_260_1913_0,
    i_13_260_1928_0, i_13_260_1950_0, i_13_260_2030_0, i_13_260_2032_0,
    i_13_260_2224_0, i_13_260_2242_0, i_13_260_2341_0, i_13_260_2454_0,
    i_13_260_2467_0, i_13_260_2468_0, i_13_260_2512_0, i_13_260_2514_0,
    i_13_260_2692_0, i_13_260_2693_0, i_13_260_2720_0, i_13_260_2750_0,
    i_13_260_2764_0, i_13_260_2912_0, i_13_260_3010_0, i_13_260_3026_0,
    i_13_260_3044_0, i_13_260_3061_0, i_13_260_3062_0, i_13_260_3128_0,
    i_13_260_3134_0, i_13_260_3146_0, i_13_260_3370_0, i_13_260_3371_0,
    i_13_260_3373_0, i_13_260_3382_0, i_13_260_3533_0, i_13_260_3596_0,
    i_13_260_3597_0, i_13_260_3598_0, i_13_260_3620_0, i_13_260_3632_0,
    i_13_260_3633_0, i_13_260_3638_0, i_13_260_3733_0, i_13_260_3783_0,
    i_13_260_3860_0, i_13_260_3925_0, i_13_260_3926_0, i_13_260_3988_0,
    i_13_260_4264_0, i_13_260_4312_0, i_13_260_4330_0, i_13_260_4331_0,
    i_13_260_4332_0, i_13_260_4414_0, i_13_260_4430_0, i_13_260_4451_0;
  output o_13_260_0_0;
  assign o_13_260_0_0 = ~(~i_13_260_4430_0 | (~i_13_260_65_0 & ~i_13_260_1397_0));
endmodule



// Benchmark "kernel_13_261" written by ABC on Sun Jul 19 10:49:03 2020

module kernel_13_261 ( 
    i_13_261_31_0, i_13_261_116_0, i_13_261_197_0, i_13_261_219_0,
    i_13_261_226_0, i_13_261_359_0, i_13_261_370_0, i_13_261_382_0,
    i_13_261_396_0, i_13_261_405_0, i_13_261_441_0, i_13_261_450_0,
    i_13_261_473_0, i_13_261_553_0, i_13_261_558_0, i_13_261_607_0,
    i_13_261_651_0, i_13_261_666_0, i_13_261_667_0, i_13_261_671_0,
    i_13_261_675_0, i_13_261_676_0, i_13_261_823_0, i_13_261_828_0,
    i_13_261_829_0, i_13_261_833_0, i_13_261_1062_0, i_13_261_1098_0,
    i_13_261_1116_0, i_13_261_1147_0, i_13_261_1148_0, i_13_261_1454_0,
    i_13_261_1492_0, i_13_261_1507_0, i_13_261_1530_0, i_13_261_1624_0,
    i_13_261_1642_0, i_13_261_1729_0, i_13_261_1754_0, i_13_261_1777_0,
    i_13_261_1795_0, i_13_261_1837_0, i_13_261_1840_0, i_13_261_1858_0,
    i_13_261_1908_0, i_13_261_1993_0, i_13_261_2020_0, i_13_261_2024_0,
    i_13_261_2045_0, i_13_261_2186_0, i_13_261_2280_0, i_13_261_2281_0,
    i_13_261_2307_0, i_13_261_2413_0, i_13_261_2431_0, i_13_261_2438_0,
    i_13_261_2456_0, i_13_261_2461_0, i_13_261_2466_0, i_13_261_2471_0,
    i_13_261_2709_0, i_13_261_2938_0, i_13_261_3097_0, i_13_261_3098_0,
    i_13_261_3104_0, i_13_261_3267_0, i_13_261_3388_0, i_13_261_3490_0,
    i_13_261_3505_0, i_13_261_3541_0, i_13_261_3599_0, i_13_261_3670_0,
    i_13_261_3725_0, i_13_261_3740_0, i_13_261_3753_0, i_13_261_3766_0,
    i_13_261_3769_0, i_13_261_3819_0, i_13_261_3910_0, i_13_261_3925_0,
    i_13_261_3987_0, i_13_261_4086_0, i_13_261_4096_0, i_13_261_4126_0,
    i_13_261_4158_0, i_13_261_4162_0, i_13_261_4165_0, i_13_261_4212_0,
    i_13_261_4213_0, i_13_261_4343_0, i_13_261_4354_0, i_13_261_4355_0,
    i_13_261_4394_0, i_13_261_4429_0, i_13_261_4433_0, i_13_261_4514_0,
    i_13_261_4540_0, i_13_261_4571_0, i_13_261_4590_0, i_13_261_4600_0,
    o_13_261_0_0  );
  input  i_13_261_31_0, i_13_261_116_0, i_13_261_197_0, i_13_261_219_0,
    i_13_261_226_0, i_13_261_359_0, i_13_261_370_0, i_13_261_382_0,
    i_13_261_396_0, i_13_261_405_0, i_13_261_441_0, i_13_261_450_0,
    i_13_261_473_0, i_13_261_553_0, i_13_261_558_0, i_13_261_607_0,
    i_13_261_651_0, i_13_261_666_0, i_13_261_667_0, i_13_261_671_0,
    i_13_261_675_0, i_13_261_676_0, i_13_261_823_0, i_13_261_828_0,
    i_13_261_829_0, i_13_261_833_0, i_13_261_1062_0, i_13_261_1098_0,
    i_13_261_1116_0, i_13_261_1147_0, i_13_261_1148_0, i_13_261_1454_0,
    i_13_261_1492_0, i_13_261_1507_0, i_13_261_1530_0, i_13_261_1624_0,
    i_13_261_1642_0, i_13_261_1729_0, i_13_261_1754_0, i_13_261_1777_0,
    i_13_261_1795_0, i_13_261_1837_0, i_13_261_1840_0, i_13_261_1858_0,
    i_13_261_1908_0, i_13_261_1993_0, i_13_261_2020_0, i_13_261_2024_0,
    i_13_261_2045_0, i_13_261_2186_0, i_13_261_2280_0, i_13_261_2281_0,
    i_13_261_2307_0, i_13_261_2413_0, i_13_261_2431_0, i_13_261_2438_0,
    i_13_261_2456_0, i_13_261_2461_0, i_13_261_2466_0, i_13_261_2471_0,
    i_13_261_2709_0, i_13_261_2938_0, i_13_261_3097_0, i_13_261_3098_0,
    i_13_261_3104_0, i_13_261_3267_0, i_13_261_3388_0, i_13_261_3490_0,
    i_13_261_3505_0, i_13_261_3541_0, i_13_261_3599_0, i_13_261_3670_0,
    i_13_261_3725_0, i_13_261_3740_0, i_13_261_3753_0, i_13_261_3766_0,
    i_13_261_3769_0, i_13_261_3819_0, i_13_261_3910_0, i_13_261_3925_0,
    i_13_261_3987_0, i_13_261_4086_0, i_13_261_4096_0, i_13_261_4126_0,
    i_13_261_4158_0, i_13_261_4162_0, i_13_261_4165_0, i_13_261_4212_0,
    i_13_261_4213_0, i_13_261_4343_0, i_13_261_4354_0, i_13_261_4355_0,
    i_13_261_4394_0, i_13_261_4429_0, i_13_261_4433_0, i_13_261_4514_0,
    i_13_261_4540_0, i_13_261_4571_0, i_13_261_4590_0, i_13_261_4600_0;
  output o_13_261_0_0;
  assign o_13_261_0_0 = ~((i_13_261_3910_0 & ~i_13_261_4162_0) | (i_13_261_382_0 & ~i_13_261_3766_0) | (~i_13_261_441_0 & ~i_13_261_3098_0) | (~i_13_261_558_0 & i_13_261_1993_0) | (~i_13_261_1116_0 & ~i_13_261_1837_0));
endmodule



// Benchmark "kernel_13_262" written by ABC on Sun Jul 19 10:49:03 2020

module kernel_13_262 ( 
    i_13_262_58_0, i_13_262_61_0, i_13_262_136_0, i_13_262_220_0,
    i_13_262_283_0, i_13_262_310_0, i_13_262_493_0, i_13_262_554_0,
    i_13_262_577_0, i_13_262_628_0, i_13_262_684_0, i_13_262_698_0,
    i_13_262_891_0, i_13_262_897_0, i_13_262_917_0, i_13_262_1071_0,
    i_13_262_1096_0, i_13_262_1111_0, i_13_262_1129_0, i_13_262_1142_0,
    i_13_262_1263_0, i_13_262_1271_0, i_13_262_1282_0, i_13_262_1299_0,
    i_13_262_1302_0, i_13_262_1304_0, i_13_262_1317_0, i_13_262_1321_0,
    i_13_262_1322_0, i_13_262_1380_0, i_13_262_1441_0, i_13_262_1462_0,
    i_13_262_1464_0, i_13_262_1480_0, i_13_262_1484_0, i_13_262_1498_0,
    i_13_262_1633_0, i_13_262_1673_0, i_13_262_1742_0, i_13_262_1756_0,
    i_13_262_1770_0, i_13_262_1774_0, i_13_262_1781_0, i_13_262_1796_0,
    i_13_262_1806_0, i_13_262_1840_0, i_13_262_1849_0, i_13_262_2002_0,
    i_13_262_2380_0, i_13_262_2382_0, i_13_262_2407_0, i_13_262_2409_0,
    i_13_262_2425_0, i_13_262_2442_0, i_13_262_2443_0, i_13_262_2446_0,
    i_13_262_2447_0, i_13_262_2498_0, i_13_262_2650_0, i_13_262_2749_0,
    i_13_262_2785_0, i_13_262_2820_0, i_13_262_2835_0, i_13_262_2871_0,
    i_13_262_2872_0, i_13_262_3035_0, i_13_262_3056_0, i_13_262_3093_0,
    i_13_262_3094_0, i_13_262_3113_0, i_13_262_3118_0, i_13_262_3145_0,
    i_13_262_3253_0, i_13_262_3311_0, i_13_262_3312_0, i_13_262_3356_0,
    i_13_262_3390_0, i_13_262_3418_0, i_13_262_3419_0, i_13_262_3516_0,
    i_13_262_3542_0, i_13_262_3766_0, i_13_262_3817_0, i_13_262_3855_0,
    i_13_262_3869_0, i_13_262_3887_0, i_13_262_3960_0, i_13_262_3963_0,
    i_13_262_3981_0, i_13_262_4018_0, i_13_262_4019_0, i_13_262_4026_0,
    i_13_262_4238_0, i_13_262_4336_0, i_13_262_4349_0, i_13_262_4377_0,
    i_13_262_4382_0, i_13_262_4407_0, i_13_262_4519_0, i_13_262_4567_0,
    o_13_262_0_0  );
  input  i_13_262_58_0, i_13_262_61_0, i_13_262_136_0, i_13_262_220_0,
    i_13_262_283_0, i_13_262_310_0, i_13_262_493_0, i_13_262_554_0,
    i_13_262_577_0, i_13_262_628_0, i_13_262_684_0, i_13_262_698_0,
    i_13_262_891_0, i_13_262_897_0, i_13_262_917_0, i_13_262_1071_0,
    i_13_262_1096_0, i_13_262_1111_0, i_13_262_1129_0, i_13_262_1142_0,
    i_13_262_1263_0, i_13_262_1271_0, i_13_262_1282_0, i_13_262_1299_0,
    i_13_262_1302_0, i_13_262_1304_0, i_13_262_1317_0, i_13_262_1321_0,
    i_13_262_1322_0, i_13_262_1380_0, i_13_262_1441_0, i_13_262_1462_0,
    i_13_262_1464_0, i_13_262_1480_0, i_13_262_1484_0, i_13_262_1498_0,
    i_13_262_1633_0, i_13_262_1673_0, i_13_262_1742_0, i_13_262_1756_0,
    i_13_262_1770_0, i_13_262_1774_0, i_13_262_1781_0, i_13_262_1796_0,
    i_13_262_1806_0, i_13_262_1840_0, i_13_262_1849_0, i_13_262_2002_0,
    i_13_262_2380_0, i_13_262_2382_0, i_13_262_2407_0, i_13_262_2409_0,
    i_13_262_2425_0, i_13_262_2442_0, i_13_262_2443_0, i_13_262_2446_0,
    i_13_262_2447_0, i_13_262_2498_0, i_13_262_2650_0, i_13_262_2749_0,
    i_13_262_2785_0, i_13_262_2820_0, i_13_262_2835_0, i_13_262_2871_0,
    i_13_262_2872_0, i_13_262_3035_0, i_13_262_3056_0, i_13_262_3093_0,
    i_13_262_3094_0, i_13_262_3113_0, i_13_262_3118_0, i_13_262_3145_0,
    i_13_262_3253_0, i_13_262_3311_0, i_13_262_3312_0, i_13_262_3356_0,
    i_13_262_3390_0, i_13_262_3418_0, i_13_262_3419_0, i_13_262_3516_0,
    i_13_262_3542_0, i_13_262_3766_0, i_13_262_3817_0, i_13_262_3855_0,
    i_13_262_3869_0, i_13_262_3887_0, i_13_262_3960_0, i_13_262_3963_0,
    i_13_262_3981_0, i_13_262_4018_0, i_13_262_4019_0, i_13_262_4026_0,
    i_13_262_4238_0, i_13_262_4336_0, i_13_262_4349_0, i_13_262_4377_0,
    i_13_262_4382_0, i_13_262_4407_0, i_13_262_4519_0, i_13_262_4567_0;
  output o_13_262_0_0;
  assign o_13_262_0_0 = ~((~i_13_262_2447_0 & ((~i_13_262_1271_0 & ((~i_13_262_58_0 & ~i_13_262_1849_0 & i_13_262_2002_0) | (~i_13_262_136_0 & ~i_13_262_1302_0 & ~i_13_262_1484_0 & ~i_13_262_2382_0 & ~i_13_262_2872_0 & ~i_13_262_3312_0))) | (~i_13_262_1480_0 & i_13_262_3766_0 & ~i_13_262_4377_0))) | (~i_13_262_58_0 & ((~i_13_262_1142_0 & ~i_13_262_1796_0 & ~i_13_262_3035_0 & ~i_13_262_3094_0) | (~i_13_262_493_0 & i_13_262_3145_0) | (~i_13_262_1480_0 & ~i_13_262_3542_0))) | (i_13_262_283_0 & i_13_262_1271_0) | (i_13_262_310_0 & i_13_262_2407_0 & ~i_13_262_2785_0 & ~i_13_262_3855_0 & ~i_13_262_4382_0));
endmodule



// Benchmark "kernel_13_263" written by ABC on Sun Jul 19 10:49:04 2020

module kernel_13_263 ( 
    i_13_263_104_0, i_13_263_124_0, i_13_263_169_0, i_13_263_197_0,
    i_13_263_203_0, i_13_263_217_0, i_13_263_382_0, i_13_263_383_0,
    i_13_263_590_0, i_13_263_607_0, i_13_263_619_0, i_13_263_626_0,
    i_13_263_718_0, i_13_263_719_0, i_13_263_838_0, i_13_263_862_0,
    i_13_263_863_0, i_13_263_932_0, i_13_263_952_0, i_13_263_1024_0,
    i_13_263_1025_0, i_13_263_1033_0, i_13_263_1147_0, i_13_263_1232_0,
    i_13_263_1243_0, i_13_263_1259_0, i_13_263_1301_0, i_13_263_1411_0,
    i_13_263_1412_0, i_13_263_1493_0, i_13_263_1529_0, i_13_263_1628_0,
    i_13_263_1711_0, i_13_263_1780_0, i_13_263_1786_0, i_13_263_1789_0,
    i_13_263_1814_0, i_13_263_1961_0, i_13_263_1990_0, i_13_263_1994_0,
    i_13_263_2006_0, i_13_263_2015_0, i_13_263_2021_0, i_13_263_2104_0,
    i_13_263_2126_0, i_13_263_2212_0, i_13_263_2213_0, i_13_263_2237_0,
    i_13_263_2246_0, i_13_263_2264_0, i_13_263_2434_0, i_13_263_2464_0,
    i_13_263_2465_0, i_13_263_2507_0, i_13_263_2536_0, i_13_263_2537_0,
    i_13_263_2545_0, i_13_263_2617_0, i_13_263_2618_0, i_13_263_2714_0,
    i_13_263_2923_0, i_13_263_2934_0, i_13_263_2938_0, i_13_263_2939_0,
    i_13_263_3040_0, i_13_263_3041_0, i_13_263_3176_0, i_13_263_3218_0,
    i_13_263_3220_0, i_13_263_3286_0, i_13_263_3290_0, i_13_263_3344_0,
    i_13_263_3388_0, i_13_263_3395_0, i_13_263_3424_0, i_13_263_3425_0,
    i_13_263_3467_0, i_13_263_3536_0, i_13_263_3613_0, i_13_263_3643_0,
    i_13_263_3644_0, i_13_263_3790_0, i_13_263_3796_0, i_13_263_3806_0,
    i_13_263_3865_0, i_13_263_3877_0, i_13_263_3878_0, i_13_263_4008_0,
    i_13_263_4012_0, i_13_263_4013_0, i_13_263_4022_0, i_13_263_4078_0,
    i_13_263_4091_0, i_13_263_4162_0, i_13_263_4333_0, i_13_263_4369_0,
    i_13_263_4410_0, i_13_263_4414_0, i_13_263_4534_0, i_13_263_4600_0,
    o_13_263_0_0  );
  input  i_13_263_104_0, i_13_263_124_0, i_13_263_169_0, i_13_263_197_0,
    i_13_263_203_0, i_13_263_217_0, i_13_263_382_0, i_13_263_383_0,
    i_13_263_590_0, i_13_263_607_0, i_13_263_619_0, i_13_263_626_0,
    i_13_263_718_0, i_13_263_719_0, i_13_263_838_0, i_13_263_862_0,
    i_13_263_863_0, i_13_263_932_0, i_13_263_952_0, i_13_263_1024_0,
    i_13_263_1025_0, i_13_263_1033_0, i_13_263_1147_0, i_13_263_1232_0,
    i_13_263_1243_0, i_13_263_1259_0, i_13_263_1301_0, i_13_263_1411_0,
    i_13_263_1412_0, i_13_263_1493_0, i_13_263_1529_0, i_13_263_1628_0,
    i_13_263_1711_0, i_13_263_1780_0, i_13_263_1786_0, i_13_263_1789_0,
    i_13_263_1814_0, i_13_263_1961_0, i_13_263_1990_0, i_13_263_1994_0,
    i_13_263_2006_0, i_13_263_2015_0, i_13_263_2021_0, i_13_263_2104_0,
    i_13_263_2126_0, i_13_263_2212_0, i_13_263_2213_0, i_13_263_2237_0,
    i_13_263_2246_0, i_13_263_2264_0, i_13_263_2434_0, i_13_263_2464_0,
    i_13_263_2465_0, i_13_263_2507_0, i_13_263_2536_0, i_13_263_2537_0,
    i_13_263_2545_0, i_13_263_2617_0, i_13_263_2618_0, i_13_263_2714_0,
    i_13_263_2923_0, i_13_263_2934_0, i_13_263_2938_0, i_13_263_2939_0,
    i_13_263_3040_0, i_13_263_3041_0, i_13_263_3176_0, i_13_263_3218_0,
    i_13_263_3220_0, i_13_263_3286_0, i_13_263_3290_0, i_13_263_3344_0,
    i_13_263_3388_0, i_13_263_3395_0, i_13_263_3424_0, i_13_263_3425_0,
    i_13_263_3467_0, i_13_263_3536_0, i_13_263_3613_0, i_13_263_3643_0,
    i_13_263_3644_0, i_13_263_3790_0, i_13_263_3796_0, i_13_263_3806_0,
    i_13_263_3865_0, i_13_263_3877_0, i_13_263_3878_0, i_13_263_4008_0,
    i_13_263_4012_0, i_13_263_4013_0, i_13_263_4022_0, i_13_263_4078_0,
    i_13_263_4091_0, i_13_263_4162_0, i_13_263_4333_0, i_13_263_4369_0,
    i_13_263_4410_0, i_13_263_4414_0, i_13_263_4534_0, i_13_263_4600_0;
  output o_13_263_0_0;
  assign o_13_263_0_0 = ~(~i_13_263_2939_0 | (~i_13_263_1025_0 & i_13_263_3865_0) | (~i_13_263_1628_0 & ~i_13_263_2212_0));
endmodule



// Benchmark "kernel_13_264" written by ABC on Sun Jul 19 10:49:05 2020

module kernel_13_264 ( 
    i_13_264_76_0, i_13_264_118_0, i_13_264_119_0, i_13_264_122_0,
    i_13_264_181_0, i_13_264_182_0, i_13_264_184_0, i_13_264_202_0,
    i_13_264_226_0, i_13_264_227_0, i_13_264_229_0, i_13_264_380_0,
    i_13_264_418_0, i_13_264_491_0, i_13_264_518_0, i_13_264_524_0,
    i_13_264_532_0, i_13_264_533_0, i_13_264_562_0, i_13_264_572_0,
    i_13_264_715_0, i_13_264_725_0, i_13_264_831_0, i_13_264_833_0,
    i_13_264_841_0, i_13_264_911_0, i_13_264_946_0, i_13_264_1046_0,
    i_13_264_1109_0, i_13_264_1112_0, i_13_264_1128_0, i_13_264_1226_0,
    i_13_264_1406_0, i_13_264_1523_0, i_13_264_1540_0, i_13_264_1690_0,
    i_13_264_1720_0, i_13_264_1721_0, i_13_264_1723_0, i_13_264_1757_0,
    i_13_264_1783_0, i_13_264_1784_0, i_13_264_1786_0, i_13_264_1787_0,
    i_13_264_1837_0, i_13_264_1838_0, i_13_264_1921_0, i_13_264_1940_0,
    i_13_264_1967_0, i_13_264_2054_0, i_13_264_2056_0, i_13_264_2110_0,
    i_13_264_2116_0, i_13_264_2120_0, i_13_264_2165_0, i_13_264_2206_0,
    i_13_264_2207_0, i_13_264_2210_0, i_13_264_2213_0, i_13_264_2225_0,
    i_13_264_2236_0, i_13_264_2295_0, i_13_264_2426_0, i_13_264_2563_0,
    i_13_264_2579_0, i_13_264_2630_0, i_13_264_2639_0, i_13_264_2786_0,
    i_13_264_3010_0, i_13_264_3020_0, i_13_264_3037_0, i_13_264_3044_0,
    i_13_264_3163_0, i_13_264_3164_0, i_13_264_3214_0, i_13_264_3260_0,
    i_13_264_3278_0, i_13_264_3422_0, i_13_264_3425_0, i_13_264_3524_0,
    i_13_264_3533_0, i_13_264_3700_0, i_13_264_3791_0, i_13_264_3836_0,
    i_13_264_3871_0, i_13_264_3872_0, i_13_264_3874_0, i_13_264_3884_0,
    i_13_264_3919_0, i_13_264_3983_0, i_13_264_4010_0, i_13_264_4087_0,
    i_13_264_4111_0, i_13_264_4258_0, i_13_264_4276_0, i_13_264_4448_0,
    i_13_264_4519_0, i_13_264_4531_0, i_13_264_4537_0, i_13_264_4583_0,
    o_13_264_0_0  );
  input  i_13_264_76_0, i_13_264_118_0, i_13_264_119_0, i_13_264_122_0,
    i_13_264_181_0, i_13_264_182_0, i_13_264_184_0, i_13_264_202_0,
    i_13_264_226_0, i_13_264_227_0, i_13_264_229_0, i_13_264_380_0,
    i_13_264_418_0, i_13_264_491_0, i_13_264_518_0, i_13_264_524_0,
    i_13_264_532_0, i_13_264_533_0, i_13_264_562_0, i_13_264_572_0,
    i_13_264_715_0, i_13_264_725_0, i_13_264_831_0, i_13_264_833_0,
    i_13_264_841_0, i_13_264_911_0, i_13_264_946_0, i_13_264_1046_0,
    i_13_264_1109_0, i_13_264_1112_0, i_13_264_1128_0, i_13_264_1226_0,
    i_13_264_1406_0, i_13_264_1523_0, i_13_264_1540_0, i_13_264_1690_0,
    i_13_264_1720_0, i_13_264_1721_0, i_13_264_1723_0, i_13_264_1757_0,
    i_13_264_1783_0, i_13_264_1784_0, i_13_264_1786_0, i_13_264_1787_0,
    i_13_264_1837_0, i_13_264_1838_0, i_13_264_1921_0, i_13_264_1940_0,
    i_13_264_1967_0, i_13_264_2054_0, i_13_264_2056_0, i_13_264_2110_0,
    i_13_264_2116_0, i_13_264_2120_0, i_13_264_2165_0, i_13_264_2206_0,
    i_13_264_2207_0, i_13_264_2210_0, i_13_264_2213_0, i_13_264_2225_0,
    i_13_264_2236_0, i_13_264_2295_0, i_13_264_2426_0, i_13_264_2563_0,
    i_13_264_2579_0, i_13_264_2630_0, i_13_264_2639_0, i_13_264_2786_0,
    i_13_264_3010_0, i_13_264_3020_0, i_13_264_3037_0, i_13_264_3044_0,
    i_13_264_3163_0, i_13_264_3164_0, i_13_264_3214_0, i_13_264_3260_0,
    i_13_264_3278_0, i_13_264_3422_0, i_13_264_3425_0, i_13_264_3524_0,
    i_13_264_3533_0, i_13_264_3700_0, i_13_264_3791_0, i_13_264_3836_0,
    i_13_264_3871_0, i_13_264_3872_0, i_13_264_3874_0, i_13_264_3884_0,
    i_13_264_3919_0, i_13_264_3983_0, i_13_264_4010_0, i_13_264_4087_0,
    i_13_264_4111_0, i_13_264_4258_0, i_13_264_4276_0, i_13_264_4448_0,
    i_13_264_4519_0, i_13_264_4531_0, i_13_264_4537_0, i_13_264_4583_0;
  output o_13_264_0_0;
  assign o_13_264_0_0 = ~(~i_13_264_3164_0 | (~i_13_264_118_0 & ~i_13_264_2207_0));
endmodule



// Benchmark "kernel_13_265" written by ABC on Sun Jul 19 10:49:06 2020

module kernel_13_265 ( 
    i_13_265_64_0, i_13_265_94_0, i_13_265_183_0, i_13_265_184_0,
    i_13_265_279_0, i_13_265_280_0, i_13_265_306_0, i_13_265_307_0,
    i_13_265_315_0, i_13_265_316_0, i_13_265_324_0, i_13_265_372_0,
    i_13_265_517_0, i_13_265_531_0, i_13_265_554_0, i_13_265_570_0,
    i_13_265_571_0, i_13_265_573_0, i_13_265_639_0, i_13_265_640_0,
    i_13_265_642_0, i_13_265_643_0, i_13_265_684_0, i_13_265_685_0,
    i_13_265_688_0, i_13_265_697_0, i_13_265_714_0, i_13_265_741_0,
    i_13_265_819_0, i_13_265_825_0, i_13_265_978_0, i_13_265_1089_0,
    i_13_265_1120_0, i_13_265_1206_0, i_13_265_1246_0, i_13_265_1269_0,
    i_13_265_1270_0, i_13_265_1380_0, i_13_265_1387_0, i_13_265_1426_0,
    i_13_265_1438_0, i_13_265_1503_0, i_13_265_1593_0, i_13_265_1594_0,
    i_13_265_1638_0, i_13_265_1639_0, i_13_265_1677_0, i_13_265_1693_0,
    i_13_265_1710_0, i_13_265_1720_0, i_13_265_1752_0, i_13_265_1804_0,
    i_13_265_1857_0, i_13_265_1858_0, i_13_265_1873_0, i_13_265_1914_0,
    i_13_265_1915_0, i_13_265_1959_0, i_13_265_2022_0, i_13_265_2023_0,
    i_13_265_2133_0, i_13_265_2134_0, i_13_265_2259_0, i_13_265_2260_0,
    i_13_265_2268_0, i_13_265_2272_0, i_13_265_2452_0, i_13_265_2472_0,
    i_13_265_2550_0, i_13_265_2646_0, i_13_265_2650_0, i_13_265_2673_0,
    i_13_265_2674_0, i_13_265_2845_0, i_13_265_2916_0, i_13_265_3024_0,
    i_13_265_3198_0, i_13_265_3205_0, i_13_265_3208_0, i_13_265_3267_0,
    i_13_265_3270_0, i_13_265_3384_0, i_13_265_3423_0, i_13_265_3735_0,
    i_13_265_3760_0, i_13_265_3817_0, i_13_265_3924_0, i_13_265_4032_0,
    i_13_265_4077_0, i_13_265_4078_0, i_13_265_4252_0, i_13_265_4344_0,
    i_13_265_4357_0, i_13_265_4369_0, i_13_265_4411_0, i_13_265_4566_0,
    i_13_265_4587_0, i_13_265_4590_0, i_13_265_4591_0, i_13_265_4592_0,
    o_13_265_0_0  );
  input  i_13_265_64_0, i_13_265_94_0, i_13_265_183_0, i_13_265_184_0,
    i_13_265_279_0, i_13_265_280_0, i_13_265_306_0, i_13_265_307_0,
    i_13_265_315_0, i_13_265_316_0, i_13_265_324_0, i_13_265_372_0,
    i_13_265_517_0, i_13_265_531_0, i_13_265_554_0, i_13_265_570_0,
    i_13_265_571_0, i_13_265_573_0, i_13_265_639_0, i_13_265_640_0,
    i_13_265_642_0, i_13_265_643_0, i_13_265_684_0, i_13_265_685_0,
    i_13_265_688_0, i_13_265_697_0, i_13_265_714_0, i_13_265_741_0,
    i_13_265_819_0, i_13_265_825_0, i_13_265_978_0, i_13_265_1089_0,
    i_13_265_1120_0, i_13_265_1206_0, i_13_265_1246_0, i_13_265_1269_0,
    i_13_265_1270_0, i_13_265_1380_0, i_13_265_1387_0, i_13_265_1426_0,
    i_13_265_1438_0, i_13_265_1503_0, i_13_265_1593_0, i_13_265_1594_0,
    i_13_265_1638_0, i_13_265_1639_0, i_13_265_1677_0, i_13_265_1693_0,
    i_13_265_1710_0, i_13_265_1720_0, i_13_265_1752_0, i_13_265_1804_0,
    i_13_265_1857_0, i_13_265_1858_0, i_13_265_1873_0, i_13_265_1914_0,
    i_13_265_1915_0, i_13_265_1959_0, i_13_265_2022_0, i_13_265_2023_0,
    i_13_265_2133_0, i_13_265_2134_0, i_13_265_2259_0, i_13_265_2260_0,
    i_13_265_2268_0, i_13_265_2272_0, i_13_265_2452_0, i_13_265_2472_0,
    i_13_265_2550_0, i_13_265_2646_0, i_13_265_2650_0, i_13_265_2673_0,
    i_13_265_2674_0, i_13_265_2845_0, i_13_265_2916_0, i_13_265_3024_0,
    i_13_265_3198_0, i_13_265_3205_0, i_13_265_3208_0, i_13_265_3267_0,
    i_13_265_3270_0, i_13_265_3384_0, i_13_265_3423_0, i_13_265_3735_0,
    i_13_265_3760_0, i_13_265_3817_0, i_13_265_3924_0, i_13_265_4032_0,
    i_13_265_4077_0, i_13_265_4078_0, i_13_265_4252_0, i_13_265_4344_0,
    i_13_265_4357_0, i_13_265_4369_0, i_13_265_4411_0, i_13_265_4566_0,
    i_13_265_4587_0, i_13_265_4590_0, i_13_265_4591_0, i_13_265_4592_0;
  output o_13_265_0_0;
  assign o_13_265_0_0 = ~((i_13_265_2272_0 & ((~i_13_265_372_0 & ~i_13_265_1270_0) | (~i_13_265_316_0 & ~i_13_265_2268_0 & ~i_13_265_2845_0))) | (~i_13_265_4077_0 & (i_13_265_697_0 | (~i_13_265_184_0 & ~i_13_265_570_0 & ~i_13_265_2650_0))) | (~i_13_265_307_0 & ~i_13_265_1639_0 & ~i_13_265_2646_0) | (~i_13_265_685_0 & ~i_13_265_3924_0));
endmodule



// Benchmark "kernel_13_266" written by ABC on Sun Jul 19 10:49:07 2020

module kernel_13_266 ( 
    i_13_266_40_0, i_13_266_48_0, i_13_266_49_0, i_13_266_51_0,
    i_13_266_101_0, i_13_266_112_0, i_13_266_139_0, i_13_266_165_0,
    i_13_266_166_0, i_13_266_216_0, i_13_266_229_0, i_13_266_265_0,
    i_13_266_282_0, i_13_266_328_0, i_13_266_365_0, i_13_266_452_0,
    i_13_266_488_0, i_13_266_500_0, i_13_266_570_0, i_13_266_676_0,
    i_13_266_737_0, i_13_266_813_0, i_13_266_814_0, i_13_266_815_0,
    i_13_266_823_0, i_13_266_840_0, i_13_266_869_0, i_13_266_960_0,
    i_13_266_1063_0, i_13_266_1166_0, i_13_266_1226_0, i_13_266_1242_0,
    i_13_266_1524_0, i_13_266_1525_0, i_13_266_1570_0, i_13_266_1624_0,
    i_13_266_1741_0, i_13_266_1753_0, i_13_266_1776_0, i_13_266_1811_0,
    i_13_266_1831_0, i_13_266_1848_0, i_13_266_1849_0, i_13_266_1882_0,
    i_13_266_1885_0, i_13_266_1943_0, i_13_266_1997_0, i_13_266_2029_0,
    i_13_266_2056_0, i_13_266_2136_0, i_13_266_2184_0, i_13_266_2201_0,
    i_13_266_2380_0, i_13_266_2403_0, i_13_266_2404_0, i_13_266_2407_0,
    i_13_266_2408_0, i_13_266_2465_0, i_13_266_2551_0, i_13_266_2693_0,
    i_13_266_2695_0, i_13_266_2756_0, i_13_266_2760_0, i_13_266_2848_0,
    i_13_266_2938_0, i_13_266_3003_0, i_13_266_3010_0, i_13_266_3092_0,
    i_13_266_3108_0, i_13_266_3109_0, i_13_266_3274_0, i_13_266_3352_0,
    i_13_266_3370_0, i_13_266_3440_0, i_13_266_3502_0, i_13_266_3505_0,
    i_13_266_3506_0, i_13_266_3640_0, i_13_266_3738_0, i_13_266_3739_0,
    i_13_266_3817_0, i_13_266_3838_0, i_13_266_3889_0, i_13_266_3892_0,
    i_13_266_3980_0, i_13_266_4017_0, i_13_266_4018_0, i_13_266_4063_0,
    i_13_266_4064_0, i_13_266_4085_0, i_13_266_4297_0, i_13_266_4315_0,
    i_13_266_4316_0, i_13_266_4318_0, i_13_266_4319_0, i_13_266_4378_0,
    i_13_266_4418_0, i_13_266_4425_0, i_13_266_4432_0, i_13_266_4544_0,
    o_13_266_0_0  );
  input  i_13_266_40_0, i_13_266_48_0, i_13_266_49_0, i_13_266_51_0,
    i_13_266_101_0, i_13_266_112_0, i_13_266_139_0, i_13_266_165_0,
    i_13_266_166_0, i_13_266_216_0, i_13_266_229_0, i_13_266_265_0,
    i_13_266_282_0, i_13_266_328_0, i_13_266_365_0, i_13_266_452_0,
    i_13_266_488_0, i_13_266_500_0, i_13_266_570_0, i_13_266_676_0,
    i_13_266_737_0, i_13_266_813_0, i_13_266_814_0, i_13_266_815_0,
    i_13_266_823_0, i_13_266_840_0, i_13_266_869_0, i_13_266_960_0,
    i_13_266_1063_0, i_13_266_1166_0, i_13_266_1226_0, i_13_266_1242_0,
    i_13_266_1524_0, i_13_266_1525_0, i_13_266_1570_0, i_13_266_1624_0,
    i_13_266_1741_0, i_13_266_1753_0, i_13_266_1776_0, i_13_266_1811_0,
    i_13_266_1831_0, i_13_266_1848_0, i_13_266_1849_0, i_13_266_1882_0,
    i_13_266_1885_0, i_13_266_1943_0, i_13_266_1997_0, i_13_266_2029_0,
    i_13_266_2056_0, i_13_266_2136_0, i_13_266_2184_0, i_13_266_2201_0,
    i_13_266_2380_0, i_13_266_2403_0, i_13_266_2404_0, i_13_266_2407_0,
    i_13_266_2408_0, i_13_266_2465_0, i_13_266_2551_0, i_13_266_2693_0,
    i_13_266_2695_0, i_13_266_2756_0, i_13_266_2760_0, i_13_266_2848_0,
    i_13_266_2938_0, i_13_266_3003_0, i_13_266_3010_0, i_13_266_3092_0,
    i_13_266_3108_0, i_13_266_3109_0, i_13_266_3274_0, i_13_266_3352_0,
    i_13_266_3370_0, i_13_266_3440_0, i_13_266_3502_0, i_13_266_3505_0,
    i_13_266_3506_0, i_13_266_3640_0, i_13_266_3738_0, i_13_266_3739_0,
    i_13_266_3817_0, i_13_266_3838_0, i_13_266_3889_0, i_13_266_3892_0,
    i_13_266_3980_0, i_13_266_4017_0, i_13_266_4018_0, i_13_266_4063_0,
    i_13_266_4064_0, i_13_266_4085_0, i_13_266_4297_0, i_13_266_4315_0,
    i_13_266_4316_0, i_13_266_4318_0, i_13_266_4319_0, i_13_266_4378_0,
    i_13_266_4418_0, i_13_266_4425_0, i_13_266_4432_0, i_13_266_4544_0;
  output o_13_266_0_0;
  assign o_13_266_0_0 = ~((~i_13_266_1524_0 & ((~i_13_266_2184_0 & ~i_13_266_4315_0) | (~i_13_266_1525_0 & i_13_266_3505_0 & i_13_266_4432_0))) | (~i_13_266_1525_0 & ((i_13_266_2380_0 & ~i_13_266_3108_0 & ~i_13_266_3889_0) | (~i_13_266_2136_0 & i_13_266_4432_0))) | (~i_13_266_1848_0 & (i_13_266_282_0 | (~i_13_266_737_0 & ~i_13_266_3108_0 & ~i_13_266_3817_0))) | (~i_13_266_3817_0 & (~i_13_266_3109_0 | (~i_13_266_813_0 & ~i_13_266_1753_0 & ~i_13_266_4085_0 & ~i_13_266_4319_0))) | (~i_13_266_1831_0 & ~i_13_266_1849_0 & ~i_13_266_4319_0) | (i_13_266_139_0 & i_13_266_3505_0) | (i_13_266_229_0 & i_13_266_1753_0 & i_13_266_4316_0) | (i_13_266_112_0 & ~i_13_266_4316_0));
endmodule



// Benchmark "kernel_13_267" written by ABC on Sun Jul 19 10:49:07 2020

module kernel_13_267 ( 
    i_13_267_28_0, i_13_267_31_0, i_13_267_63_0, i_13_267_64_0,
    i_13_267_90_0, i_13_267_91_0, i_13_267_94_0, i_13_267_95_0,
    i_13_267_225_0, i_13_267_226_0, i_13_267_287_0, i_13_267_306_0,
    i_13_267_307_0, i_13_267_355_0, i_13_267_367_0, i_13_267_369_0,
    i_13_267_380_0, i_13_267_468_0, i_13_267_538_0, i_13_267_606_0,
    i_13_267_607_0, i_13_267_616_0, i_13_267_649_0, i_13_267_667_0,
    i_13_267_729_0, i_13_267_756_0, i_13_267_757_0, i_13_267_814_0,
    i_13_267_829_0, i_13_267_945_0, i_13_267_946_0, i_13_267_953_0,
    i_13_267_1075_0, i_13_267_1076_0, i_13_267_1099_0, i_13_267_1215_0,
    i_13_267_1218_0, i_13_267_1219_0, i_13_267_1228_0, i_13_267_1306_0,
    i_13_267_1318_0, i_13_267_1444_0, i_13_267_1462_0, i_13_267_1594_0,
    i_13_267_1678_0, i_13_267_1719_0, i_13_267_1720_0, i_13_267_1777_0,
    i_13_267_1790_0, i_13_267_1840_0, i_13_267_1843_0, i_13_267_1844_0,
    i_13_267_1858_0, i_13_267_1926_0, i_13_267_1999_0, i_13_267_2001_0,
    i_13_267_2172_0, i_13_267_2176_0, i_13_267_2407_0, i_13_267_2421_0,
    i_13_267_2478_0, i_13_267_2534_0, i_13_267_2676_0, i_13_267_2718_0,
    i_13_267_2719_0, i_13_267_2749_0, i_13_267_2785_0, i_13_267_2821_0,
    i_13_267_2881_0, i_13_267_3028_0, i_13_267_3060_0, i_13_267_3063_0,
    i_13_267_3109_0, i_13_267_3116_0, i_13_267_3119_0, i_13_267_3149_0,
    i_13_267_3241_0, i_13_267_3316_0, i_13_267_3416_0, i_13_267_3460_0,
    i_13_267_3464_0, i_13_267_3636_0, i_13_267_3712_0, i_13_267_3738_0,
    i_13_267_3760_0, i_13_267_3797_0, i_13_267_3875_0, i_13_267_3910_0,
    i_13_267_3925_0, i_13_267_3929_0, i_13_267_3932_0, i_13_267_3979_0,
    i_13_267_4060_0, i_13_267_4093_0, i_13_267_4120_0, i_13_267_4212_0,
    i_13_267_4213_0, i_13_267_4351_0, i_13_267_4354_0, i_13_267_4544_0,
    o_13_267_0_0  );
  input  i_13_267_28_0, i_13_267_31_0, i_13_267_63_0, i_13_267_64_0,
    i_13_267_90_0, i_13_267_91_0, i_13_267_94_0, i_13_267_95_0,
    i_13_267_225_0, i_13_267_226_0, i_13_267_287_0, i_13_267_306_0,
    i_13_267_307_0, i_13_267_355_0, i_13_267_367_0, i_13_267_369_0,
    i_13_267_380_0, i_13_267_468_0, i_13_267_538_0, i_13_267_606_0,
    i_13_267_607_0, i_13_267_616_0, i_13_267_649_0, i_13_267_667_0,
    i_13_267_729_0, i_13_267_756_0, i_13_267_757_0, i_13_267_814_0,
    i_13_267_829_0, i_13_267_945_0, i_13_267_946_0, i_13_267_953_0,
    i_13_267_1075_0, i_13_267_1076_0, i_13_267_1099_0, i_13_267_1215_0,
    i_13_267_1218_0, i_13_267_1219_0, i_13_267_1228_0, i_13_267_1306_0,
    i_13_267_1318_0, i_13_267_1444_0, i_13_267_1462_0, i_13_267_1594_0,
    i_13_267_1678_0, i_13_267_1719_0, i_13_267_1720_0, i_13_267_1777_0,
    i_13_267_1790_0, i_13_267_1840_0, i_13_267_1843_0, i_13_267_1844_0,
    i_13_267_1858_0, i_13_267_1926_0, i_13_267_1999_0, i_13_267_2001_0,
    i_13_267_2172_0, i_13_267_2176_0, i_13_267_2407_0, i_13_267_2421_0,
    i_13_267_2478_0, i_13_267_2534_0, i_13_267_2676_0, i_13_267_2718_0,
    i_13_267_2719_0, i_13_267_2749_0, i_13_267_2785_0, i_13_267_2821_0,
    i_13_267_2881_0, i_13_267_3028_0, i_13_267_3060_0, i_13_267_3063_0,
    i_13_267_3109_0, i_13_267_3116_0, i_13_267_3119_0, i_13_267_3149_0,
    i_13_267_3241_0, i_13_267_3316_0, i_13_267_3416_0, i_13_267_3460_0,
    i_13_267_3464_0, i_13_267_3636_0, i_13_267_3712_0, i_13_267_3738_0,
    i_13_267_3760_0, i_13_267_3797_0, i_13_267_3875_0, i_13_267_3910_0,
    i_13_267_3925_0, i_13_267_3929_0, i_13_267_3932_0, i_13_267_3979_0,
    i_13_267_4060_0, i_13_267_4093_0, i_13_267_4120_0, i_13_267_4212_0,
    i_13_267_4213_0, i_13_267_4351_0, i_13_267_4354_0, i_13_267_4544_0;
  output o_13_267_0_0;
  assign o_13_267_0_0 = ~(~i_13_267_226_0 | (~i_13_267_1306_0 & i_13_267_3875_0) | (~i_13_267_95_0 & ~i_13_267_945_0 & ~i_13_267_1215_0) | (~i_13_267_64_0 & ~i_13_267_1218_0 & ~i_13_267_1219_0 & ~i_13_267_2421_0) | (~i_13_267_306_0 & ~i_13_267_380_0 & ~i_13_267_468_0 & ~i_13_267_3063_0 & ~i_13_267_3241_0));
endmodule



// Benchmark "kernel_13_268" written by ABC on Sun Jul 19 10:49:08 2020

module kernel_13_268 ( 
    i_13_268_103_0, i_13_268_133_0, i_13_268_134_0, i_13_268_139_0,
    i_13_268_237_0, i_13_268_252_0, i_13_268_280_0, i_13_268_319_0,
    i_13_268_326_0, i_13_268_429_0, i_13_268_469_0, i_13_268_524_0,
    i_13_268_588_0, i_13_268_608_0, i_13_268_668_0, i_13_268_821_0,
    i_13_268_852_0, i_13_268_951_0, i_13_268_1021_0, i_13_268_1066_0,
    i_13_268_1076_0, i_13_268_1122_0, i_13_268_1230_0, i_13_268_1275_0,
    i_13_268_1311_0, i_13_268_1343_0, i_13_268_1401_0, i_13_268_1426_0,
    i_13_268_1428_0, i_13_268_1468_0, i_13_268_1499_0, i_13_268_1509_0,
    i_13_268_1599_0, i_13_268_1634_0, i_13_268_1644_0, i_13_268_1651_0,
    i_13_268_1680_0, i_13_268_1691_0, i_13_268_1696_0, i_13_268_1712_0,
    i_13_268_1777_0, i_13_268_1778_0, i_13_268_1794_0, i_13_268_1797_0,
    i_13_268_1811_0, i_13_268_1882_0, i_13_268_1883_0, i_13_268_1914_0,
    i_13_268_1929_0, i_13_268_1990_0, i_13_268_1991_0, i_13_268_1999_0,
    i_13_268_2000_0, i_13_268_2002_0, i_13_268_2003_0, i_13_268_2115_0,
    i_13_268_2134_0, i_13_268_2198_0, i_13_268_2237_0, i_13_268_2265_0,
    i_13_268_2377_0, i_13_268_2461_0, i_13_268_2470_0, i_13_268_2647_0,
    i_13_268_2711_0, i_13_268_2763_0, i_13_268_2845_0, i_13_268_2854_0,
    i_13_268_2935_0, i_13_268_2983_0, i_13_268_3142_0, i_13_268_3143_0,
    i_13_268_3172_0, i_13_268_3273_0, i_13_268_3448_0, i_13_268_3461_0,
    i_13_268_3503_0, i_13_268_3727_0, i_13_268_3728_0, i_13_268_3731_0,
    i_13_268_3783_0, i_13_268_3816_0, i_13_268_3838_0, i_13_268_3874_0,
    i_13_268_4015_0, i_13_268_4016_0, i_13_268_4038_0, i_13_268_4083_0,
    i_13_268_4097_0, i_13_268_4162_0, i_13_268_4259_0, i_13_268_4268_0,
    i_13_268_4270_0, i_13_268_4314_0, i_13_268_4393_0, i_13_268_4411_0,
    i_13_268_4554_0, i_13_268_4558_0, i_13_268_4567_0, i_13_268_4568_0,
    o_13_268_0_0  );
  input  i_13_268_103_0, i_13_268_133_0, i_13_268_134_0, i_13_268_139_0,
    i_13_268_237_0, i_13_268_252_0, i_13_268_280_0, i_13_268_319_0,
    i_13_268_326_0, i_13_268_429_0, i_13_268_469_0, i_13_268_524_0,
    i_13_268_588_0, i_13_268_608_0, i_13_268_668_0, i_13_268_821_0,
    i_13_268_852_0, i_13_268_951_0, i_13_268_1021_0, i_13_268_1066_0,
    i_13_268_1076_0, i_13_268_1122_0, i_13_268_1230_0, i_13_268_1275_0,
    i_13_268_1311_0, i_13_268_1343_0, i_13_268_1401_0, i_13_268_1426_0,
    i_13_268_1428_0, i_13_268_1468_0, i_13_268_1499_0, i_13_268_1509_0,
    i_13_268_1599_0, i_13_268_1634_0, i_13_268_1644_0, i_13_268_1651_0,
    i_13_268_1680_0, i_13_268_1691_0, i_13_268_1696_0, i_13_268_1712_0,
    i_13_268_1777_0, i_13_268_1778_0, i_13_268_1794_0, i_13_268_1797_0,
    i_13_268_1811_0, i_13_268_1882_0, i_13_268_1883_0, i_13_268_1914_0,
    i_13_268_1929_0, i_13_268_1990_0, i_13_268_1991_0, i_13_268_1999_0,
    i_13_268_2000_0, i_13_268_2002_0, i_13_268_2003_0, i_13_268_2115_0,
    i_13_268_2134_0, i_13_268_2198_0, i_13_268_2237_0, i_13_268_2265_0,
    i_13_268_2377_0, i_13_268_2461_0, i_13_268_2470_0, i_13_268_2647_0,
    i_13_268_2711_0, i_13_268_2763_0, i_13_268_2845_0, i_13_268_2854_0,
    i_13_268_2935_0, i_13_268_2983_0, i_13_268_3142_0, i_13_268_3143_0,
    i_13_268_3172_0, i_13_268_3273_0, i_13_268_3448_0, i_13_268_3461_0,
    i_13_268_3503_0, i_13_268_3727_0, i_13_268_3728_0, i_13_268_3731_0,
    i_13_268_3783_0, i_13_268_3816_0, i_13_268_3838_0, i_13_268_3874_0,
    i_13_268_4015_0, i_13_268_4016_0, i_13_268_4038_0, i_13_268_4083_0,
    i_13_268_4097_0, i_13_268_4162_0, i_13_268_4259_0, i_13_268_4268_0,
    i_13_268_4270_0, i_13_268_4314_0, i_13_268_4393_0, i_13_268_4411_0,
    i_13_268_4554_0, i_13_268_4558_0, i_13_268_4567_0, i_13_268_4568_0;
  output o_13_268_0_0;
  assign o_13_268_0_0 = ~((~i_13_268_1778_0 & ~i_13_268_4411_0) | (i_13_268_1066_0 & ~i_13_268_4162_0) | (~i_13_268_2845_0 & ~i_13_268_3461_0 & ~i_13_268_3731_0) | (~i_13_268_1883_0 & ~i_13_268_2647_0 & ~i_13_268_3728_0));
endmodule



// Benchmark "kernel_13_269" written by ABC on Sun Jul 19 10:49:09 2020

module kernel_13_269 ( 
    i_13_269_30_0, i_13_269_75_0, i_13_269_111_0, i_13_269_114_0,
    i_13_269_115_0, i_13_269_123_0, i_13_269_124_0, i_13_269_247_0,
    i_13_269_265_0, i_13_269_276_0, i_13_269_363_0, i_13_269_366_0,
    i_13_269_418_0, i_13_269_444_0, i_13_269_561_0, i_13_269_564_0,
    i_13_269_606_0, i_13_269_607_0, i_13_269_609_0, i_13_269_654_0,
    i_13_269_663_0, i_13_269_670_0, i_13_269_672_0, i_13_269_688_0,
    i_13_269_814_0, i_13_269_817_0, i_13_269_939_0, i_13_269_949_0,
    i_13_269_1083_0, i_13_269_1084_0, i_13_269_1086_0, i_13_269_1114_0,
    i_13_269_1408_0, i_13_269_1434_0, i_13_269_1446_0, i_13_269_1470_0,
    i_13_269_1626_0, i_13_269_1653_0, i_13_269_1750_0, i_13_269_1776_0,
    i_13_269_1804_0, i_13_269_1839_0, i_13_269_1840_0, i_13_269_1842_0,
    i_13_269_1843_0, i_13_269_2056_0, i_13_269_2130_0, i_13_269_2136_0,
    i_13_269_2157_0, i_13_269_2172_0, i_13_269_2173_0, i_13_269_2175_0,
    i_13_269_2247_0, i_13_269_2299_0, i_13_269_2347_0, i_13_269_2407_0,
    i_13_269_2425_0, i_13_269_2434_0, i_13_269_2436_0, i_13_269_2437_0,
    i_13_269_2452_0, i_13_269_2497_0, i_13_269_2581_0, i_13_269_2704_0,
    i_13_269_2748_0, i_13_269_2938_0, i_13_269_3031_0, i_13_269_3049_0,
    i_13_269_3099_0, i_13_269_3100_0, i_13_269_3103_0, i_13_269_3147_0,
    i_13_269_3148_0, i_13_269_3156_0, i_13_269_3165_0, i_13_269_3261_0,
    i_13_269_3504_0, i_13_269_3505_0, i_13_269_3541_0, i_13_269_3615_0,
    i_13_269_3688_0, i_13_269_3741_0, i_13_269_3760_0, i_13_269_3769_0,
    i_13_269_3784_0, i_13_269_3877_0, i_13_269_3891_0, i_13_269_3909_0,
    i_13_269_3910_0, i_13_269_4044_0, i_13_269_4084_0, i_13_269_4119_0,
    i_13_269_4120_0, i_13_269_4162_0, i_13_269_4327_0, i_13_269_4353_0,
    i_13_269_4354_0, i_13_269_4449_0, i_13_269_4528_0, i_13_269_4543_0,
    o_13_269_0_0  );
  input  i_13_269_30_0, i_13_269_75_0, i_13_269_111_0, i_13_269_114_0,
    i_13_269_115_0, i_13_269_123_0, i_13_269_124_0, i_13_269_247_0,
    i_13_269_265_0, i_13_269_276_0, i_13_269_363_0, i_13_269_366_0,
    i_13_269_418_0, i_13_269_444_0, i_13_269_561_0, i_13_269_564_0,
    i_13_269_606_0, i_13_269_607_0, i_13_269_609_0, i_13_269_654_0,
    i_13_269_663_0, i_13_269_670_0, i_13_269_672_0, i_13_269_688_0,
    i_13_269_814_0, i_13_269_817_0, i_13_269_939_0, i_13_269_949_0,
    i_13_269_1083_0, i_13_269_1084_0, i_13_269_1086_0, i_13_269_1114_0,
    i_13_269_1408_0, i_13_269_1434_0, i_13_269_1446_0, i_13_269_1470_0,
    i_13_269_1626_0, i_13_269_1653_0, i_13_269_1750_0, i_13_269_1776_0,
    i_13_269_1804_0, i_13_269_1839_0, i_13_269_1840_0, i_13_269_1842_0,
    i_13_269_1843_0, i_13_269_2056_0, i_13_269_2130_0, i_13_269_2136_0,
    i_13_269_2157_0, i_13_269_2172_0, i_13_269_2173_0, i_13_269_2175_0,
    i_13_269_2247_0, i_13_269_2299_0, i_13_269_2347_0, i_13_269_2407_0,
    i_13_269_2425_0, i_13_269_2434_0, i_13_269_2436_0, i_13_269_2437_0,
    i_13_269_2452_0, i_13_269_2497_0, i_13_269_2581_0, i_13_269_2704_0,
    i_13_269_2748_0, i_13_269_2938_0, i_13_269_3031_0, i_13_269_3049_0,
    i_13_269_3099_0, i_13_269_3100_0, i_13_269_3103_0, i_13_269_3147_0,
    i_13_269_3148_0, i_13_269_3156_0, i_13_269_3165_0, i_13_269_3261_0,
    i_13_269_3504_0, i_13_269_3505_0, i_13_269_3541_0, i_13_269_3615_0,
    i_13_269_3688_0, i_13_269_3741_0, i_13_269_3760_0, i_13_269_3769_0,
    i_13_269_3784_0, i_13_269_3877_0, i_13_269_3891_0, i_13_269_3909_0,
    i_13_269_3910_0, i_13_269_4044_0, i_13_269_4084_0, i_13_269_4119_0,
    i_13_269_4120_0, i_13_269_4162_0, i_13_269_4327_0, i_13_269_4353_0,
    i_13_269_4354_0, i_13_269_4449_0, i_13_269_4528_0, i_13_269_4543_0;
  output o_13_269_0_0;
  assign o_13_269_0_0 = ~(~i_13_269_1843_0 | (~i_13_269_1626_0 & ~i_13_269_4354_0) | (~i_13_269_3099_0 & ~i_13_269_4353_0));
endmodule



// Benchmark "kernel_13_270" written by ABC on Sun Jul 19 10:49:10 2020

module kernel_13_270 ( 
    i_13_270_25_0, i_13_270_61_0, i_13_270_76_0, i_13_270_119_0,
    i_13_270_163_0, i_13_270_164_0, i_13_270_177_0, i_13_270_182_0,
    i_13_270_184_0, i_13_270_185_0, i_13_270_186_0, i_13_270_187_0,
    i_13_270_192_0, i_13_270_193_0, i_13_270_194_0, i_13_270_196_0,
    i_13_270_347_0, i_13_270_382_0, i_13_270_419_0, i_13_270_518_0,
    i_13_270_571_0, i_13_270_573_0, i_13_270_574_0, i_13_270_625_0,
    i_13_270_628_0, i_13_270_661_0, i_13_270_697_0, i_13_270_715_0,
    i_13_270_717_0, i_13_270_811_0, i_13_270_837_0, i_13_270_841_0,
    i_13_270_850_0, i_13_270_853_0, i_13_270_1151_0, i_13_270_1210_0,
    i_13_270_1211_0, i_13_270_1285_0, i_13_270_1406_0, i_13_270_1407_0,
    i_13_270_1408_0, i_13_270_1409_0, i_13_270_1411_0, i_13_270_1416_0,
    i_13_270_1426_0, i_13_270_1471_0, i_13_270_1516_0, i_13_270_1525_0,
    i_13_270_1681_0, i_13_270_1770_0, i_13_270_1771_0, i_13_270_1805_0,
    i_13_270_1831_0, i_13_270_1832_0, i_13_270_1834_0, i_13_270_1908_0,
    i_13_270_1912_0, i_13_270_1959_0, i_13_270_1960_0, i_13_270_2002_0,
    i_13_270_2146_0, i_13_270_2178_0, i_13_270_2403_0, i_13_270_2452_0,
    i_13_270_2504_0, i_13_270_2563_0, i_13_270_2572_0, i_13_270_2612_0,
    i_13_270_2723_0, i_13_270_2736_0, i_13_270_2857_0, i_13_270_2983_0,
    i_13_270_3049_0, i_13_270_3064_0, i_13_270_3065_0, i_13_270_3108_0,
    i_13_270_3145_0, i_13_270_3164_0, i_13_270_3165_0, i_13_270_3166_0,
    i_13_270_3208_0, i_13_270_3209_0, i_13_270_3212_0, i_13_270_3215_0,
    i_13_270_3261_0, i_13_270_3446_0, i_13_270_3602_0, i_13_270_3604_0,
    i_13_270_3616_0, i_13_270_3685_0, i_13_270_3730_0, i_13_270_3733_0,
    i_13_270_3901_0, i_13_270_3979_0, i_13_270_4073_0, i_13_270_4162_0,
    i_13_270_4261_0, i_13_270_4396_0, i_13_270_4421_0, i_13_270_4569_0,
    o_13_270_0_0  );
  input  i_13_270_25_0, i_13_270_61_0, i_13_270_76_0, i_13_270_119_0,
    i_13_270_163_0, i_13_270_164_0, i_13_270_177_0, i_13_270_182_0,
    i_13_270_184_0, i_13_270_185_0, i_13_270_186_0, i_13_270_187_0,
    i_13_270_192_0, i_13_270_193_0, i_13_270_194_0, i_13_270_196_0,
    i_13_270_347_0, i_13_270_382_0, i_13_270_419_0, i_13_270_518_0,
    i_13_270_571_0, i_13_270_573_0, i_13_270_574_0, i_13_270_625_0,
    i_13_270_628_0, i_13_270_661_0, i_13_270_697_0, i_13_270_715_0,
    i_13_270_717_0, i_13_270_811_0, i_13_270_837_0, i_13_270_841_0,
    i_13_270_850_0, i_13_270_853_0, i_13_270_1151_0, i_13_270_1210_0,
    i_13_270_1211_0, i_13_270_1285_0, i_13_270_1406_0, i_13_270_1407_0,
    i_13_270_1408_0, i_13_270_1409_0, i_13_270_1411_0, i_13_270_1416_0,
    i_13_270_1426_0, i_13_270_1471_0, i_13_270_1516_0, i_13_270_1525_0,
    i_13_270_1681_0, i_13_270_1770_0, i_13_270_1771_0, i_13_270_1805_0,
    i_13_270_1831_0, i_13_270_1832_0, i_13_270_1834_0, i_13_270_1908_0,
    i_13_270_1912_0, i_13_270_1959_0, i_13_270_1960_0, i_13_270_2002_0,
    i_13_270_2146_0, i_13_270_2178_0, i_13_270_2403_0, i_13_270_2452_0,
    i_13_270_2504_0, i_13_270_2563_0, i_13_270_2572_0, i_13_270_2612_0,
    i_13_270_2723_0, i_13_270_2736_0, i_13_270_2857_0, i_13_270_2983_0,
    i_13_270_3049_0, i_13_270_3064_0, i_13_270_3065_0, i_13_270_3108_0,
    i_13_270_3145_0, i_13_270_3164_0, i_13_270_3165_0, i_13_270_3166_0,
    i_13_270_3208_0, i_13_270_3209_0, i_13_270_3212_0, i_13_270_3215_0,
    i_13_270_3261_0, i_13_270_3446_0, i_13_270_3602_0, i_13_270_3604_0,
    i_13_270_3616_0, i_13_270_3685_0, i_13_270_3730_0, i_13_270_3733_0,
    i_13_270_3901_0, i_13_270_3979_0, i_13_270_4073_0, i_13_270_4162_0,
    i_13_270_4261_0, i_13_270_4396_0, i_13_270_4421_0, i_13_270_4569_0;
  output o_13_270_0_0;
  assign o_13_270_0_0 = ~((~i_13_270_185_0 & ~i_13_270_1407_0 & ((~i_13_270_194_0 & ~i_13_270_1408_0 & ~i_13_270_1681_0 & ~i_13_270_3108_0) | (~i_13_270_182_0 & ~i_13_270_187_0 & ~i_13_270_811_0 & ~i_13_270_4569_0))) | (i_13_270_2002_0 & ((~i_13_270_2146_0 & i_13_270_2403_0) | (~i_13_270_61_0 & ~i_13_270_1409_0 & ~i_13_270_3212_0 & ~i_13_270_3261_0 & ~i_13_270_4569_0))) | (i_13_270_2452_0 & i_13_270_3145_0 & ~i_13_270_3166_0 & i_13_270_3209_0) | (i_13_270_1210_0 & ~i_13_270_1408_0 & ~i_13_270_1960_0 & ~i_13_270_3215_0) | (~i_13_270_3208_0 & i_13_270_3730_0 & ~i_13_270_4569_0));
endmodule



// Benchmark "kernel_13_271" written by ABC on Sun Jul 19 10:49:10 2020

module kernel_13_271 ( 
    i_13_271_46_0, i_13_271_48_0, i_13_271_117_0, i_13_271_118_0,
    i_13_271_127_0, i_13_271_164_0, i_13_271_189_0, i_13_271_323_0,
    i_13_271_409_0, i_13_271_504_0, i_13_271_532_0, i_13_271_572_0,
    i_13_271_604_0, i_13_271_616_0, i_13_271_711_0, i_13_271_712_0,
    i_13_271_832_0, i_13_271_909_0, i_13_271_918_0, i_13_271_935_0,
    i_13_271_1081_0, i_13_271_1147_0, i_13_271_1226_0, i_13_271_1252_0,
    i_13_271_1378_0, i_13_271_1404_0, i_13_271_1426_0, i_13_271_1435_0,
    i_13_271_1440_0, i_13_271_1495_0, i_13_271_1503_0, i_13_271_1513_0,
    i_13_271_1514_0, i_13_271_1534_0, i_13_271_1548_0, i_13_271_1549_0,
    i_13_271_1595_0, i_13_271_1664_0, i_13_271_1695_0, i_13_271_1711_0,
    i_13_271_1728_0, i_13_271_1764_0, i_13_271_1766_0, i_13_271_1768_0,
    i_13_271_1795_0, i_13_271_1906_0, i_13_271_1916_0, i_13_271_2025_0,
    i_13_271_2056_0, i_13_271_2097_0, i_13_271_2143_0, i_13_271_2149_0,
    i_13_271_2172_0, i_13_271_2286_0, i_13_271_2296_0, i_13_271_2360_0,
    i_13_271_2379_0, i_13_271_2430_0, i_13_271_2529_0, i_13_271_2744_0,
    i_13_271_2901_0, i_13_271_2978_0, i_13_271_3106_0, i_13_271_3113_0,
    i_13_271_3123_0, i_13_271_3132_0, i_13_271_3214_0, i_13_271_3261_0,
    i_13_271_3367_0, i_13_271_3547_0, i_13_271_3565_0, i_13_271_3574_0,
    i_13_271_3637_0, i_13_271_3645_0, i_13_271_3782_0, i_13_271_3843_0,
    i_13_271_3844_0, i_13_271_3888_0, i_13_271_3897_0, i_13_271_3898_0,
    i_13_271_3908_0, i_13_271_3910_0, i_13_271_3913_0, i_13_271_3916_0,
    i_13_271_3979_0, i_13_271_3982_0, i_13_271_4019_0, i_13_271_4042_0,
    i_13_271_4097_0, i_13_271_4159_0, i_13_271_4230_0, i_13_271_4266_0,
    i_13_271_4293_0, i_13_271_4321_0, i_13_271_4331_0, i_13_271_4401_0,
    i_13_271_4509_0, i_13_271_4510_0, i_13_271_4536_0, i_13_271_4606_0,
    o_13_271_0_0  );
  input  i_13_271_46_0, i_13_271_48_0, i_13_271_117_0, i_13_271_118_0,
    i_13_271_127_0, i_13_271_164_0, i_13_271_189_0, i_13_271_323_0,
    i_13_271_409_0, i_13_271_504_0, i_13_271_532_0, i_13_271_572_0,
    i_13_271_604_0, i_13_271_616_0, i_13_271_711_0, i_13_271_712_0,
    i_13_271_832_0, i_13_271_909_0, i_13_271_918_0, i_13_271_935_0,
    i_13_271_1081_0, i_13_271_1147_0, i_13_271_1226_0, i_13_271_1252_0,
    i_13_271_1378_0, i_13_271_1404_0, i_13_271_1426_0, i_13_271_1435_0,
    i_13_271_1440_0, i_13_271_1495_0, i_13_271_1503_0, i_13_271_1513_0,
    i_13_271_1514_0, i_13_271_1534_0, i_13_271_1548_0, i_13_271_1549_0,
    i_13_271_1595_0, i_13_271_1664_0, i_13_271_1695_0, i_13_271_1711_0,
    i_13_271_1728_0, i_13_271_1764_0, i_13_271_1766_0, i_13_271_1768_0,
    i_13_271_1795_0, i_13_271_1906_0, i_13_271_1916_0, i_13_271_2025_0,
    i_13_271_2056_0, i_13_271_2097_0, i_13_271_2143_0, i_13_271_2149_0,
    i_13_271_2172_0, i_13_271_2286_0, i_13_271_2296_0, i_13_271_2360_0,
    i_13_271_2379_0, i_13_271_2430_0, i_13_271_2529_0, i_13_271_2744_0,
    i_13_271_2901_0, i_13_271_2978_0, i_13_271_3106_0, i_13_271_3113_0,
    i_13_271_3123_0, i_13_271_3132_0, i_13_271_3214_0, i_13_271_3261_0,
    i_13_271_3367_0, i_13_271_3547_0, i_13_271_3565_0, i_13_271_3574_0,
    i_13_271_3637_0, i_13_271_3645_0, i_13_271_3782_0, i_13_271_3843_0,
    i_13_271_3844_0, i_13_271_3888_0, i_13_271_3897_0, i_13_271_3898_0,
    i_13_271_3908_0, i_13_271_3910_0, i_13_271_3913_0, i_13_271_3916_0,
    i_13_271_3979_0, i_13_271_3982_0, i_13_271_4019_0, i_13_271_4042_0,
    i_13_271_4097_0, i_13_271_4159_0, i_13_271_4230_0, i_13_271_4266_0,
    i_13_271_4293_0, i_13_271_4321_0, i_13_271_4331_0, i_13_271_4401_0,
    i_13_271_4509_0, i_13_271_4510_0, i_13_271_4536_0, i_13_271_4606_0;
  output o_13_271_0_0;
  assign o_13_271_0_0 = ~((~i_13_271_118_0 & (~i_13_271_3547_0 | (~i_13_271_3261_0 & ~i_13_271_4266_0))) | (~i_13_271_1226_0 & ~i_13_271_1549_0 & ~i_13_271_2529_0 & ~i_13_271_4266_0) | (~i_13_271_832_0 & ~i_13_271_1503_0 & i_13_271_3910_0) | (~i_13_271_3106_0 & ~i_13_271_3214_0 & ~i_13_271_3910_0) | (~i_13_271_1404_0 & ~i_13_271_3979_0 & ~i_13_271_4331_0 & ~i_13_271_4509_0));
endmodule



// Benchmark "kernel_13_272" written by ABC on Sun Jul 19 10:49:11 2020

module kernel_13_272 ( 
    i_13_272_29_0, i_13_272_47_0, i_13_272_71_0, i_13_272_155_0,
    i_13_272_209_0, i_13_272_231_0, i_13_272_269_0, i_13_272_300_0,
    i_13_272_314_0, i_13_272_352_0, i_13_272_416_0, i_13_272_445_0,
    i_13_272_583_0, i_13_272_610_0, i_13_272_628_0, i_13_272_646_0,
    i_13_272_647_0, i_13_272_689_0, i_13_272_713_0, i_13_272_764_0,
    i_13_272_854_0, i_13_272_953_0, i_13_272_985_0, i_13_272_986_0,
    i_13_272_1086_0, i_13_272_1106_0, i_13_272_1132_0, i_13_272_1136_0,
    i_13_272_1226_0, i_13_272_1303_0, i_13_272_1408_0, i_13_272_1495_0,
    i_13_272_1511_0, i_13_272_1525_0, i_13_272_1551_0, i_13_272_1606_0,
    i_13_272_1644_0, i_13_272_1717_0, i_13_272_1753_0, i_13_272_1754_0,
    i_13_272_1799_0, i_13_272_1802_0, i_13_272_1808_0, i_13_272_1918_0,
    i_13_272_1945_0, i_13_272_1996_0, i_13_272_2122_0, i_13_272_2123_0,
    i_13_272_2193_0, i_13_272_2195_0, i_13_272_2240_0, i_13_272_2294_0,
    i_13_272_2373_0, i_13_272_2390_0, i_13_272_2473_0, i_13_272_2515_0,
    i_13_272_2518_0, i_13_272_2545_0, i_13_272_2567_0, i_13_272_2680_0,
    i_13_272_2695_0, i_13_272_2698_0, i_13_272_2699_0, i_13_272_2715_0,
    i_13_272_2786_0, i_13_272_2816_0, i_13_272_2911_0, i_13_272_2941_0,
    i_13_272_3014_0, i_13_272_3021_0, i_13_272_3031_0, i_13_272_3032_0,
    i_13_272_3128_0, i_13_272_3133_0, i_13_272_3134_0, i_13_272_3212_0,
    i_13_272_3232_0, i_13_272_3262_0, i_13_272_3264_0, i_13_272_3347_0,
    i_13_272_3355_0, i_13_272_3399_0, i_13_272_3453_0, i_13_272_3589_0,
    i_13_272_3700_0, i_13_272_3760_0, i_13_272_3782_0, i_13_272_3853_0,
    i_13_272_3916_0, i_13_272_4038_0, i_13_272_4046_0, i_13_272_4085_0,
    i_13_272_4254_0, i_13_272_4273_0, i_13_272_4326_0, i_13_272_4396_0,
    i_13_272_4398_0, i_13_272_4557_0, i_13_272_4597_0, i_13_272_4607_0,
    o_13_272_0_0  );
  input  i_13_272_29_0, i_13_272_47_0, i_13_272_71_0, i_13_272_155_0,
    i_13_272_209_0, i_13_272_231_0, i_13_272_269_0, i_13_272_300_0,
    i_13_272_314_0, i_13_272_352_0, i_13_272_416_0, i_13_272_445_0,
    i_13_272_583_0, i_13_272_610_0, i_13_272_628_0, i_13_272_646_0,
    i_13_272_647_0, i_13_272_689_0, i_13_272_713_0, i_13_272_764_0,
    i_13_272_854_0, i_13_272_953_0, i_13_272_985_0, i_13_272_986_0,
    i_13_272_1086_0, i_13_272_1106_0, i_13_272_1132_0, i_13_272_1136_0,
    i_13_272_1226_0, i_13_272_1303_0, i_13_272_1408_0, i_13_272_1495_0,
    i_13_272_1511_0, i_13_272_1525_0, i_13_272_1551_0, i_13_272_1606_0,
    i_13_272_1644_0, i_13_272_1717_0, i_13_272_1753_0, i_13_272_1754_0,
    i_13_272_1799_0, i_13_272_1802_0, i_13_272_1808_0, i_13_272_1918_0,
    i_13_272_1945_0, i_13_272_1996_0, i_13_272_2122_0, i_13_272_2123_0,
    i_13_272_2193_0, i_13_272_2195_0, i_13_272_2240_0, i_13_272_2294_0,
    i_13_272_2373_0, i_13_272_2390_0, i_13_272_2473_0, i_13_272_2515_0,
    i_13_272_2518_0, i_13_272_2545_0, i_13_272_2567_0, i_13_272_2680_0,
    i_13_272_2695_0, i_13_272_2698_0, i_13_272_2699_0, i_13_272_2715_0,
    i_13_272_2786_0, i_13_272_2816_0, i_13_272_2911_0, i_13_272_2941_0,
    i_13_272_3014_0, i_13_272_3021_0, i_13_272_3031_0, i_13_272_3032_0,
    i_13_272_3128_0, i_13_272_3133_0, i_13_272_3134_0, i_13_272_3212_0,
    i_13_272_3232_0, i_13_272_3262_0, i_13_272_3264_0, i_13_272_3347_0,
    i_13_272_3355_0, i_13_272_3399_0, i_13_272_3453_0, i_13_272_3589_0,
    i_13_272_3700_0, i_13_272_3760_0, i_13_272_3782_0, i_13_272_3853_0,
    i_13_272_3916_0, i_13_272_4038_0, i_13_272_4046_0, i_13_272_4085_0,
    i_13_272_4254_0, i_13_272_4273_0, i_13_272_4326_0, i_13_272_4396_0,
    i_13_272_4398_0, i_13_272_4557_0, i_13_272_4597_0, i_13_272_4607_0;
  output o_13_272_0_0;
  assign o_13_272_0_0 = 0;
endmodule



// Benchmark "kernel_13_273" written by ABC on Sun Jul 19 10:49:12 2020

module kernel_13_273 ( 
    i_13_273_106_0, i_13_273_107_0, i_13_273_124_0, i_13_273_142_0,
    i_13_273_170_0, i_13_273_184_0, i_13_273_269_0, i_13_273_320_0,
    i_13_273_340_0, i_13_273_341_0, i_13_273_380_0, i_13_273_449_0,
    i_13_273_458_0, i_13_273_511_0, i_13_273_618_0, i_13_273_746_0,
    i_13_273_781_0, i_13_273_817_0, i_13_273_818_0, i_13_273_836_0,
    i_13_273_934_0, i_13_273_980_0, i_13_273_1055_0, i_13_273_1220_0,
    i_13_273_1222_0, i_13_273_1303_0, i_13_273_1304_0, i_13_273_1309_0,
    i_13_273_1349_0, i_13_273_1465_0, i_13_273_1573_0, i_13_273_1574_0,
    i_13_273_1723_0, i_13_273_1789_0, i_13_273_1808_0, i_13_273_1817_0,
    i_13_273_1825_0, i_13_273_1996_0, i_13_273_1997_0, i_13_273_2053_0,
    i_13_273_2060_0, i_13_273_2122_0, i_13_273_2123_0, i_13_273_2140_0,
    i_13_273_2141_0, i_13_273_2411_0, i_13_273_2438_0, i_13_273_2461_0,
    i_13_273_2506_0, i_13_273_2573_0, i_13_273_2582_0, i_13_273_2728_0,
    i_13_273_2729_0, i_13_273_2752_0, i_13_273_2861_0, i_13_273_2940_0,
    i_13_273_2941_0, i_13_273_2942_0, i_13_273_3001_0, i_13_273_3022_0,
    i_13_273_3023_0, i_13_273_3030_0, i_13_273_3220_0, i_13_273_3221_0,
    i_13_273_3238_0, i_13_273_3272_0, i_13_273_3292_0, i_13_273_3293_0,
    i_13_273_3346_0, i_13_273_3347_0, i_13_273_3386_0, i_13_273_3391_0,
    i_13_273_3392_0, i_13_273_3400_0, i_13_273_3401_0, i_13_273_3418_0,
    i_13_273_3419_0, i_13_273_3437_0, i_13_273_3505_0, i_13_273_3526_0,
    i_13_273_3527_0, i_13_273_3560_0, i_13_273_3670_0, i_13_273_3824_0,
    i_13_273_3881_0, i_13_273_3911_0, i_13_273_3926_0, i_13_273_4049_0,
    i_13_273_4058_0, i_13_273_4067_0, i_13_273_4166_0, i_13_273_4273_0,
    i_13_273_4318_0, i_13_273_4319_0, i_13_273_4332_0, i_13_273_4372_0,
    i_13_273_4396_0, i_13_273_4400_0, i_13_273_4416_0, i_13_273_4594_0,
    o_13_273_0_0  );
  input  i_13_273_106_0, i_13_273_107_0, i_13_273_124_0, i_13_273_142_0,
    i_13_273_170_0, i_13_273_184_0, i_13_273_269_0, i_13_273_320_0,
    i_13_273_340_0, i_13_273_341_0, i_13_273_380_0, i_13_273_449_0,
    i_13_273_458_0, i_13_273_511_0, i_13_273_618_0, i_13_273_746_0,
    i_13_273_781_0, i_13_273_817_0, i_13_273_818_0, i_13_273_836_0,
    i_13_273_934_0, i_13_273_980_0, i_13_273_1055_0, i_13_273_1220_0,
    i_13_273_1222_0, i_13_273_1303_0, i_13_273_1304_0, i_13_273_1309_0,
    i_13_273_1349_0, i_13_273_1465_0, i_13_273_1573_0, i_13_273_1574_0,
    i_13_273_1723_0, i_13_273_1789_0, i_13_273_1808_0, i_13_273_1817_0,
    i_13_273_1825_0, i_13_273_1996_0, i_13_273_1997_0, i_13_273_2053_0,
    i_13_273_2060_0, i_13_273_2122_0, i_13_273_2123_0, i_13_273_2140_0,
    i_13_273_2141_0, i_13_273_2411_0, i_13_273_2438_0, i_13_273_2461_0,
    i_13_273_2506_0, i_13_273_2573_0, i_13_273_2582_0, i_13_273_2728_0,
    i_13_273_2729_0, i_13_273_2752_0, i_13_273_2861_0, i_13_273_2940_0,
    i_13_273_2941_0, i_13_273_2942_0, i_13_273_3001_0, i_13_273_3022_0,
    i_13_273_3023_0, i_13_273_3030_0, i_13_273_3220_0, i_13_273_3221_0,
    i_13_273_3238_0, i_13_273_3272_0, i_13_273_3292_0, i_13_273_3293_0,
    i_13_273_3346_0, i_13_273_3347_0, i_13_273_3386_0, i_13_273_3391_0,
    i_13_273_3392_0, i_13_273_3400_0, i_13_273_3401_0, i_13_273_3418_0,
    i_13_273_3419_0, i_13_273_3437_0, i_13_273_3505_0, i_13_273_3526_0,
    i_13_273_3527_0, i_13_273_3560_0, i_13_273_3670_0, i_13_273_3824_0,
    i_13_273_3881_0, i_13_273_3911_0, i_13_273_3926_0, i_13_273_4049_0,
    i_13_273_4058_0, i_13_273_4067_0, i_13_273_4166_0, i_13_273_4273_0,
    i_13_273_4318_0, i_13_273_4319_0, i_13_273_4332_0, i_13_273_4372_0,
    i_13_273_4396_0, i_13_273_4400_0, i_13_273_4416_0, i_13_273_4594_0;
  output o_13_273_0_0;
  assign o_13_273_0_0 = ~((i_13_273_4332_0 & ((~i_13_273_3526_0 & (~i_13_273_2140_0 | (~i_13_273_340_0 & ~i_13_273_3220_0))) | ~i_13_273_4273_0 | (i_13_273_1222_0 & ~i_13_273_4416_0))) | (~i_13_273_1303_0 & ~i_13_273_1573_0 & ~i_13_273_3346_0 & ~i_13_273_3527_0));
endmodule



// Benchmark "kernel_13_274" written by ABC on Sun Jul 19 10:49:13 2020

module kernel_13_274 ( 
    i_13_274_177_0, i_13_274_274_0, i_13_274_281_0, i_13_274_310_0,
    i_13_274_312_0, i_13_274_313_0, i_13_274_314_0, i_13_274_315_0,
    i_13_274_318_0, i_13_274_320_0, i_13_274_554_0, i_13_274_587_0,
    i_13_274_642_0, i_13_274_643_0, i_13_274_645_0, i_13_274_647_0,
    i_13_274_688_0, i_13_274_689_0, i_13_274_691_0, i_13_274_692_0,
    i_13_274_820_0, i_13_274_840_0, i_13_274_854_0, i_13_274_871_0,
    i_13_274_1106_0, i_13_274_1119_0, i_13_274_1123_0, i_13_274_1124_0,
    i_13_274_1211_0, i_13_274_1223_0, i_13_274_1276_0, i_13_274_1277_0,
    i_13_274_1283_0, i_13_274_1308_0, i_13_274_1311_0, i_13_274_1343_0,
    i_13_274_1391_0, i_13_274_1394_0, i_13_274_1399_0, i_13_274_1442_0,
    i_13_274_1511_0, i_13_274_1593_0, i_13_274_1597_0, i_13_274_1600_0,
    i_13_274_1633_0, i_13_274_1642_0, i_13_274_1649_0, i_13_274_1791_0,
    i_13_274_1798_0, i_13_274_1799_0, i_13_274_1853_0, i_13_274_1997_0,
    i_13_274_2000_0, i_13_274_2001_0, i_13_274_2003_0, i_13_274_2004_0,
    i_13_274_2055_0, i_13_274_2057_0, i_13_274_2194_0, i_13_274_2262_0,
    i_13_274_2270_0, i_13_274_2272_0, i_13_274_2303_0, i_13_274_2434_0,
    i_13_274_2555_0, i_13_274_2588_0, i_13_274_2651_0, i_13_274_2680_0,
    i_13_274_2681_0, i_13_274_2711_0, i_13_274_3011_0, i_13_274_3037_0,
    i_13_274_3246_0, i_13_274_3272_0, i_13_274_3368_0, i_13_274_3415_0,
    i_13_274_3419_0, i_13_274_3653_0, i_13_274_3666_0, i_13_274_3736_0,
    i_13_274_3743_0, i_13_274_3782_0, i_13_274_3868_0, i_13_274_3931_0,
    i_13_274_3990_0, i_13_274_3995_0, i_13_274_4043_0, i_13_274_4081_0,
    i_13_274_4085_0, i_13_274_4090_0, i_13_274_4190_0, i_13_274_4193_0,
    i_13_274_4207_0, i_13_274_4232_0, i_13_274_4297_0, i_13_274_4531_0,
    i_13_274_4594_0, i_13_274_4595_0, i_13_274_4598_0, i_13_274_4604_0,
    o_13_274_0_0  );
  input  i_13_274_177_0, i_13_274_274_0, i_13_274_281_0, i_13_274_310_0,
    i_13_274_312_0, i_13_274_313_0, i_13_274_314_0, i_13_274_315_0,
    i_13_274_318_0, i_13_274_320_0, i_13_274_554_0, i_13_274_587_0,
    i_13_274_642_0, i_13_274_643_0, i_13_274_645_0, i_13_274_647_0,
    i_13_274_688_0, i_13_274_689_0, i_13_274_691_0, i_13_274_692_0,
    i_13_274_820_0, i_13_274_840_0, i_13_274_854_0, i_13_274_871_0,
    i_13_274_1106_0, i_13_274_1119_0, i_13_274_1123_0, i_13_274_1124_0,
    i_13_274_1211_0, i_13_274_1223_0, i_13_274_1276_0, i_13_274_1277_0,
    i_13_274_1283_0, i_13_274_1308_0, i_13_274_1311_0, i_13_274_1343_0,
    i_13_274_1391_0, i_13_274_1394_0, i_13_274_1399_0, i_13_274_1442_0,
    i_13_274_1511_0, i_13_274_1593_0, i_13_274_1597_0, i_13_274_1600_0,
    i_13_274_1633_0, i_13_274_1642_0, i_13_274_1649_0, i_13_274_1791_0,
    i_13_274_1798_0, i_13_274_1799_0, i_13_274_1853_0, i_13_274_1997_0,
    i_13_274_2000_0, i_13_274_2001_0, i_13_274_2003_0, i_13_274_2004_0,
    i_13_274_2055_0, i_13_274_2057_0, i_13_274_2194_0, i_13_274_2262_0,
    i_13_274_2270_0, i_13_274_2272_0, i_13_274_2303_0, i_13_274_2434_0,
    i_13_274_2555_0, i_13_274_2588_0, i_13_274_2651_0, i_13_274_2680_0,
    i_13_274_2681_0, i_13_274_2711_0, i_13_274_3011_0, i_13_274_3037_0,
    i_13_274_3246_0, i_13_274_3272_0, i_13_274_3368_0, i_13_274_3415_0,
    i_13_274_3419_0, i_13_274_3653_0, i_13_274_3666_0, i_13_274_3736_0,
    i_13_274_3743_0, i_13_274_3782_0, i_13_274_3868_0, i_13_274_3931_0,
    i_13_274_3990_0, i_13_274_3995_0, i_13_274_4043_0, i_13_274_4081_0,
    i_13_274_4085_0, i_13_274_4090_0, i_13_274_4190_0, i_13_274_4193_0,
    i_13_274_4207_0, i_13_274_4232_0, i_13_274_4297_0, i_13_274_4531_0,
    i_13_274_4594_0, i_13_274_4595_0, i_13_274_4598_0, i_13_274_4604_0;
  output o_13_274_0_0;
  assign o_13_274_0_0 = ~((i_13_274_2434_0 & ~i_13_274_3931_0) | (~i_13_274_1600_0 & i_13_274_2272_0) | (~i_13_274_1798_0 & i_13_274_2001_0) | (~i_13_274_692_0 & ~i_13_274_1123_0 & ~i_13_274_1799_0));
endmodule



// Benchmark "kernel_13_275" written by ABC on Sun Jul 19 10:49:13 2020

module kernel_13_275 ( 
    i_13_275_63_0, i_13_275_64_0, i_13_275_75_0, i_13_275_103_0,
    i_13_275_174_0, i_13_275_184_0, i_13_275_211_0, i_13_275_379_0,
    i_13_275_453_0, i_13_275_523_0, i_13_275_558_0, i_13_275_567_0,
    i_13_275_585_0, i_13_275_696_0, i_13_275_707_0, i_13_275_738_0,
    i_13_275_741_0, i_13_275_759_0, i_13_275_840_0, i_13_275_855_0,
    i_13_275_1092_0, i_13_275_1093_0, i_13_275_1137_0, i_13_275_1180_0,
    i_13_275_1192_0, i_13_275_1200_0, i_13_275_1206_0, i_13_275_1207_0,
    i_13_275_1209_0, i_13_275_1341_0, i_13_275_1342_0, i_13_275_1425_0,
    i_13_275_1441_0, i_13_275_1467_0, i_13_275_1468_0, i_13_275_1569_0,
    i_13_275_1604_0, i_13_275_1649_0, i_13_275_1755_0, i_13_275_1810_0,
    i_13_275_1855_0, i_13_275_1857_0, i_13_275_1858_0, i_13_275_1920_0,
    i_13_275_1927_0, i_13_275_1944_0, i_13_275_1946_0, i_13_275_2001_0,
    i_13_275_2052_0, i_13_275_2053_0, i_13_275_2055_0, i_13_275_2187_0,
    i_13_275_2262_0, i_13_275_2277_0, i_13_275_2278_0, i_13_275_2341_0,
    i_13_275_2350_0, i_13_275_2376_0, i_13_275_2563_0, i_13_275_2596_0,
    i_13_275_2676_0, i_13_275_2709_0, i_13_275_2719_0, i_13_275_2722_0,
    i_13_275_2766_0, i_13_275_2767_0, i_13_275_2856_0, i_13_275_2857_0,
    i_13_275_2934_0, i_13_275_3060_0, i_13_275_3061_0, i_13_275_3063_0,
    i_13_275_3098_0, i_13_275_3126_0, i_13_275_3366_0, i_13_275_3369_0,
    i_13_275_3414_0, i_13_275_3415_0, i_13_275_3438_0, i_13_275_3439_0,
    i_13_275_3592_0, i_13_275_3627_0, i_13_275_3681_0, i_13_275_3684_0,
    i_13_275_3726_0, i_13_275_3910_0, i_13_275_4015_0, i_13_275_4033_0,
    i_13_275_4152_0, i_13_275_4203_0, i_13_275_4230_0, i_13_275_4302_0,
    i_13_275_4305_0, i_13_275_4306_0, i_13_275_4348_0, i_13_275_4393_0,
    i_13_275_4395_0, i_13_275_4410_0, i_13_275_4441_0, i_13_275_4554_0,
    o_13_275_0_0  );
  input  i_13_275_63_0, i_13_275_64_0, i_13_275_75_0, i_13_275_103_0,
    i_13_275_174_0, i_13_275_184_0, i_13_275_211_0, i_13_275_379_0,
    i_13_275_453_0, i_13_275_523_0, i_13_275_558_0, i_13_275_567_0,
    i_13_275_585_0, i_13_275_696_0, i_13_275_707_0, i_13_275_738_0,
    i_13_275_741_0, i_13_275_759_0, i_13_275_840_0, i_13_275_855_0,
    i_13_275_1092_0, i_13_275_1093_0, i_13_275_1137_0, i_13_275_1180_0,
    i_13_275_1192_0, i_13_275_1200_0, i_13_275_1206_0, i_13_275_1207_0,
    i_13_275_1209_0, i_13_275_1341_0, i_13_275_1342_0, i_13_275_1425_0,
    i_13_275_1441_0, i_13_275_1467_0, i_13_275_1468_0, i_13_275_1569_0,
    i_13_275_1604_0, i_13_275_1649_0, i_13_275_1755_0, i_13_275_1810_0,
    i_13_275_1855_0, i_13_275_1857_0, i_13_275_1858_0, i_13_275_1920_0,
    i_13_275_1927_0, i_13_275_1944_0, i_13_275_1946_0, i_13_275_2001_0,
    i_13_275_2052_0, i_13_275_2053_0, i_13_275_2055_0, i_13_275_2187_0,
    i_13_275_2262_0, i_13_275_2277_0, i_13_275_2278_0, i_13_275_2341_0,
    i_13_275_2350_0, i_13_275_2376_0, i_13_275_2563_0, i_13_275_2596_0,
    i_13_275_2676_0, i_13_275_2709_0, i_13_275_2719_0, i_13_275_2722_0,
    i_13_275_2766_0, i_13_275_2767_0, i_13_275_2856_0, i_13_275_2857_0,
    i_13_275_2934_0, i_13_275_3060_0, i_13_275_3061_0, i_13_275_3063_0,
    i_13_275_3098_0, i_13_275_3126_0, i_13_275_3366_0, i_13_275_3369_0,
    i_13_275_3414_0, i_13_275_3415_0, i_13_275_3438_0, i_13_275_3439_0,
    i_13_275_3592_0, i_13_275_3627_0, i_13_275_3681_0, i_13_275_3684_0,
    i_13_275_3726_0, i_13_275_3910_0, i_13_275_4015_0, i_13_275_4033_0,
    i_13_275_4152_0, i_13_275_4203_0, i_13_275_4230_0, i_13_275_4302_0,
    i_13_275_4305_0, i_13_275_4306_0, i_13_275_4348_0, i_13_275_4393_0,
    i_13_275_4395_0, i_13_275_4410_0, i_13_275_4441_0, i_13_275_4554_0;
  output o_13_275_0_0;
  assign o_13_275_0_0 = ~((~i_13_275_2052_0 & ~i_13_275_3438_0) | (~i_13_275_1341_0 & ~i_13_275_2277_0 & ~i_13_275_3061_0));
endmodule



// Benchmark "kernel_13_276" written by ABC on Sun Jul 19 10:49:14 2020

module kernel_13_276 ( 
    i_13_276_37_0, i_13_276_61_0, i_13_276_117_0, i_13_276_189_0,
    i_13_276_190_0, i_13_276_222_0, i_13_276_223_0, i_13_276_226_0,
    i_13_276_273_0, i_13_276_333_0, i_13_276_387_0, i_13_276_396_0,
    i_13_276_408_0, i_13_276_561_0, i_13_276_567_0, i_13_276_585_0,
    i_13_276_603_0, i_13_276_604_0, i_13_276_607_0, i_13_276_608_0,
    i_13_276_629_0, i_13_276_657_0, i_13_276_669_0, i_13_276_742_0,
    i_13_276_855_0, i_13_276_945_0, i_13_276_1083_0, i_13_276_1112_0,
    i_13_276_1368_0, i_13_276_1404_0, i_13_276_1440_0, i_13_276_1486_0,
    i_13_276_1516_0, i_13_276_1620_0, i_13_276_1623_0, i_13_276_1729_0,
    i_13_276_1745_0, i_13_276_1785_0, i_13_276_1813_0, i_13_276_1836_0,
    i_13_276_1837_0, i_13_276_1840_0, i_13_276_1844_0, i_13_276_1924_0,
    i_13_276_2019_0, i_13_276_2020_0, i_13_276_2023_0, i_13_276_2137_0,
    i_13_276_2214_0, i_13_276_2359_0, i_13_276_2422_0, i_13_276_2431_0,
    i_13_276_2497_0, i_13_276_2529_0, i_13_276_2622_0, i_13_276_2650_0,
    i_13_276_2907_0, i_13_276_3043_0, i_13_276_3099_0, i_13_276_3101_0,
    i_13_276_3114_0, i_13_276_3126_0, i_13_276_3160_0, i_13_276_3163_0,
    i_13_276_3261_0, i_13_276_3274_0, i_13_276_3307_0, i_13_276_3322_0,
    i_13_276_3465_0, i_13_276_3475_0, i_13_276_3523_0, i_13_276_3565_0,
    i_13_276_3567_0, i_13_276_3598_0, i_13_276_3600_0, i_13_276_3648_0,
    i_13_276_3730_0, i_13_276_3738_0, i_13_276_3762_0, i_13_276_3763_0,
    i_13_276_3784_0, i_13_276_3819_0, i_13_276_3843_0, i_13_276_3897_0,
    i_13_276_3978_0, i_13_276_4005_0, i_13_276_4116_0, i_13_276_4117_0,
    i_13_276_4158_0, i_13_276_4159_0, i_13_276_4161_0, i_13_276_4162_0,
    i_13_276_4260_0, i_13_276_4315_0, i_13_276_4324_0, i_13_276_4355_0,
    i_13_276_4366_0, i_13_276_4467_0, i_13_276_4507_0, i_13_276_4537_0,
    o_13_276_0_0  );
  input  i_13_276_37_0, i_13_276_61_0, i_13_276_117_0, i_13_276_189_0,
    i_13_276_190_0, i_13_276_222_0, i_13_276_223_0, i_13_276_226_0,
    i_13_276_273_0, i_13_276_333_0, i_13_276_387_0, i_13_276_396_0,
    i_13_276_408_0, i_13_276_561_0, i_13_276_567_0, i_13_276_585_0,
    i_13_276_603_0, i_13_276_604_0, i_13_276_607_0, i_13_276_608_0,
    i_13_276_629_0, i_13_276_657_0, i_13_276_669_0, i_13_276_742_0,
    i_13_276_855_0, i_13_276_945_0, i_13_276_1083_0, i_13_276_1112_0,
    i_13_276_1368_0, i_13_276_1404_0, i_13_276_1440_0, i_13_276_1486_0,
    i_13_276_1516_0, i_13_276_1620_0, i_13_276_1623_0, i_13_276_1729_0,
    i_13_276_1745_0, i_13_276_1785_0, i_13_276_1813_0, i_13_276_1836_0,
    i_13_276_1837_0, i_13_276_1840_0, i_13_276_1844_0, i_13_276_1924_0,
    i_13_276_2019_0, i_13_276_2020_0, i_13_276_2023_0, i_13_276_2137_0,
    i_13_276_2214_0, i_13_276_2359_0, i_13_276_2422_0, i_13_276_2431_0,
    i_13_276_2497_0, i_13_276_2529_0, i_13_276_2622_0, i_13_276_2650_0,
    i_13_276_2907_0, i_13_276_3043_0, i_13_276_3099_0, i_13_276_3101_0,
    i_13_276_3114_0, i_13_276_3126_0, i_13_276_3160_0, i_13_276_3163_0,
    i_13_276_3261_0, i_13_276_3274_0, i_13_276_3307_0, i_13_276_3322_0,
    i_13_276_3465_0, i_13_276_3475_0, i_13_276_3523_0, i_13_276_3565_0,
    i_13_276_3567_0, i_13_276_3598_0, i_13_276_3600_0, i_13_276_3648_0,
    i_13_276_3730_0, i_13_276_3738_0, i_13_276_3762_0, i_13_276_3763_0,
    i_13_276_3784_0, i_13_276_3819_0, i_13_276_3843_0, i_13_276_3897_0,
    i_13_276_3978_0, i_13_276_4005_0, i_13_276_4116_0, i_13_276_4117_0,
    i_13_276_4158_0, i_13_276_4159_0, i_13_276_4161_0, i_13_276_4162_0,
    i_13_276_4260_0, i_13_276_4315_0, i_13_276_4324_0, i_13_276_4355_0,
    i_13_276_4366_0, i_13_276_4467_0, i_13_276_4507_0, i_13_276_4537_0;
  output o_13_276_0_0;
  assign o_13_276_0_0 = ~(~i_13_276_3763_0 | (~i_13_276_1083_0 & ~i_13_276_1836_0 & ~i_13_276_3819_0));
endmodule



// Benchmark "kernel_13_277" written by ABC on Sun Jul 19 10:49:15 2020

module kernel_13_277 ( 
    i_13_277_130_0, i_13_277_170_0, i_13_277_286_0, i_13_277_352_0,
    i_13_277_383_0, i_13_277_422_0, i_13_277_461_0, i_13_277_466_0,
    i_13_277_467_0, i_13_277_512_0, i_13_277_526_0, i_13_277_527_0,
    i_13_277_529_0, i_13_277_530_0, i_13_277_535_0, i_13_277_547_0,
    i_13_277_625_0, i_13_277_800_0, i_13_277_817_0, i_13_277_881_0,
    i_13_277_1025_0, i_13_277_1148_0, i_13_277_1273_0, i_13_277_1313_0,
    i_13_277_1516_0, i_13_277_1553_0, i_13_277_1556_0, i_13_277_1600_0,
    i_13_277_1634_0, i_13_277_1636_0, i_13_277_1678_0, i_13_277_1849_0,
    i_13_277_1940_0, i_13_277_2005_0, i_13_277_2006_0, i_13_277_2033_0,
    i_13_277_2105_0, i_13_277_2131_0, i_13_277_2137_0, i_13_277_2200_0,
    i_13_277_2203_0, i_13_277_2204_0, i_13_277_2267_0, i_13_277_2278_0,
    i_13_277_2363_0, i_13_277_2408_0, i_13_277_2462_0, i_13_277_2465_0,
    i_13_277_2474_0, i_13_277_2510_0, i_13_277_2545_0, i_13_277_2546_0,
    i_13_277_2557_0, i_13_277_2618_0, i_13_277_2690_0, i_13_277_2711_0,
    i_13_277_2747_0, i_13_277_2806_0, i_13_277_2852_0, i_13_277_2939_0,
    i_13_277_3100_0, i_13_277_3118_0, i_13_277_3125_0, i_13_277_3235_0,
    i_13_277_3265_0, i_13_277_3346_0, i_13_277_3368_0, i_13_277_3461_0,
    i_13_277_3541_0, i_13_277_3598_0, i_13_277_3644_0, i_13_277_3667_0,
    i_13_277_3670_0, i_13_277_3730_0, i_13_277_3731_0, i_13_277_3733_0,
    i_13_277_3734_0, i_13_277_3742_0, i_13_277_3787_0, i_13_277_3860_0,
    i_13_277_3910_0, i_13_277_3913_0, i_13_277_3914_0, i_13_277_3920_0,
    i_13_277_4018_0, i_13_277_4019_0, i_13_277_4063_0, i_13_277_4064_0,
    i_13_277_4210_0, i_13_277_4255_0, i_13_277_4256_0, i_13_277_4265_0,
    i_13_277_4298_0, i_13_277_4316_0, i_13_277_4342_0, i_13_277_4393_0,
    i_13_277_4423_0, i_13_277_4543_0, i_13_277_4561_0, i_13_277_4603_0,
    o_13_277_0_0  );
  input  i_13_277_130_0, i_13_277_170_0, i_13_277_286_0, i_13_277_352_0,
    i_13_277_383_0, i_13_277_422_0, i_13_277_461_0, i_13_277_466_0,
    i_13_277_467_0, i_13_277_512_0, i_13_277_526_0, i_13_277_527_0,
    i_13_277_529_0, i_13_277_530_0, i_13_277_535_0, i_13_277_547_0,
    i_13_277_625_0, i_13_277_800_0, i_13_277_817_0, i_13_277_881_0,
    i_13_277_1025_0, i_13_277_1148_0, i_13_277_1273_0, i_13_277_1313_0,
    i_13_277_1516_0, i_13_277_1553_0, i_13_277_1556_0, i_13_277_1600_0,
    i_13_277_1634_0, i_13_277_1636_0, i_13_277_1678_0, i_13_277_1849_0,
    i_13_277_1940_0, i_13_277_2005_0, i_13_277_2006_0, i_13_277_2033_0,
    i_13_277_2105_0, i_13_277_2131_0, i_13_277_2137_0, i_13_277_2200_0,
    i_13_277_2203_0, i_13_277_2204_0, i_13_277_2267_0, i_13_277_2278_0,
    i_13_277_2363_0, i_13_277_2408_0, i_13_277_2462_0, i_13_277_2465_0,
    i_13_277_2474_0, i_13_277_2510_0, i_13_277_2545_0, i_13_277_2546_0,
    i_13_277_2557_0, i_13_277_2618_0, i_13_277_2690_0, i_13_277_2711_0,
    i_13_277_2747_0, i_13_277_2806_0, i_13_277_2852_0, i_13_277_2939_0,
    i_13_277_3100_0, i_13_277_3118_0, i_13_277_3125_0, i_13_277_3235_0,
    i_13_277_3265_0, i_13_277_3346_0, i_13_277_3368_0, i_13_277_3461_0,
    i_13_277_3541_0, i_13_277_3598_0, i_13_277_3644_0, i_13_277_3667_0,
    i_13_277_3670_0, i_13_277_3730_0, i_13_277_3731_0, i_13_277_3733_0,
    i_13_277_3734_0, i_13_277_3742_0, i_13_277_3787_0, i_13_277_3860_0,
    i_13_277_3910_0, i_13_277_3913_0, i_13_277_3914_0, i_13_277_3920_0,
    i_13_277_4018_0, i_13_277_4019_0, i_13_277_4063_0, i_13_277_4064_0,
    i_13_277_4210_0, i_13_277_4255_0, i_13_277_4256_0, i_13_277_4265_0,
    i_13_277_4298_0, i_13_277_4316_0, i_13_277_4342_0, i_13_277_4393_0,
    i_13_277_4423_0, i_13_277_4543_0, i_13_277_4561_0, i_13_277_4603_0;
  output o_13_277_0_0;
  assign o_13_277_0_0 = ~((~i_13_277_2939_0 & ~i_13_277_4561_0) | (~i_13_277_3541_0 & ~i_13_277_3920_0) | (~i_13_277_422_0 & ~i_13_277_2203_0));
endmodule



// Benchmark "kernel_13_278" written by ABC on Sun Jul 19 10:49:16 2020

module kernel_13_278 ( 
    i_13_278_0_0, i_13_278_14_0, i_13_278_22_0, i_13_278_64_0,
    i_13_278_76_0, i_13_278_168_0, i_13_278_182_0, i_13_278_199_0,
    i_13_278_225_0, i_13_278_228_0, i_13_278_247_0, i_13_278_280_0,
    i_13_278_336_0, i_13_278_339_0, i_13_278_378_0, i_13_278_381_0,
    i_13_278_531_0, i_13_278_536_0, i_13_278_573_0, i_13_278_585_0,
    i_13_278_586_0, i_13_278_639_0, i_13_278_640_0, i_13_278_717_0,
    i_13_278_781_0, i_13_278_927_0, i_13_278_1004_0, i_13_278_1064_0,
    i_13_278_1081_0, i_13_278_1116_0, i_13_278_1117_0, i_13_278_1141_0,
    i_13_278_1142_0, i_13_278_1181_0, i_13_278_1296_0, i_13_278_1467_0,
    i_13_278_1468_0, i_13_278_1470_0, i_13_278_1497_0, i_13_278_1503_0,
    i_13_278_1647_0, i_13_278_1648_0, i_13_278_1710_0, i_13_278_1711_0,
    i_13_278_1719_0, i_13_278_1731_0, i_13_278_1782_0, i_13_278_1786_0,
    i_13_278_1791_0, i_13_278_1792_0, i_13_278_1800_0, i_13_278_1802_0,
    i_13_278_1851_0, i_13_278_1989_0, i_13_278_1990_0, i_13_278_1993_0,
    i_13_278_2115_0, i_13_278_2116_0, i_13_278_2259_0, i_13_278_2265_0,
    i_13_278_2290_0, i_13_278_2358_0, i_13_278_2377_0, i_13_278_2379_0,
    i_13_278_2536_0, i_13_278_2667_0, i_13_278_2672_0, i_13_278_2673_0,
    i_13_278_2709_0, i_13_278_2844_0, i_13_278_2845_0, i_13_278_2934_0,
    i_13_278_3036_0, i_13_278_3040_0, i_13_278_3061_0, i_13_278_3123_0,
    i_13_278_3153_0, i_13_278_3215_0, i_13_278_3285_0, i_13_278_3286_0,
    i_13_278_3468_0, i_13_278_3475_0, i_13_278_3550_0, i_13_278_3554_0,
    i_13_278_3581_0, i_13_278_3610_0, i_13_278_3639_0, i_13_278_3818_0,
    i_13_278_3924_0, i_13_278_4008_0, i_13_278_4011_0, i_13_278_4042_0,
    i_13_278_4230_0, i_13_278_4232_0, i_13_278_4302_0, i_13_278_4303_0,
    i_13_278_4390_0, i_13_278_4391_0, i_13_278_4410_0, i_13_278_4411_0,
    o_13_278_0_0  );
  input  i_13_278_0_0, i_13_278_14_0, i_13_278_22_0, i_13_278_64_0,
    i_13_278_76_0, i_13_278_168_0, i_13_278_182_0, i_13_278_199_0,
    i_13_278_225_0, i_13_278_228_0, i_13_278_247_0, i_13_278_280_0,
    i_13_278_336_0, i_13_278_339_0, i_13_278_378_0, i_13_278_381_0,
    i_13_278_531_0, i_13_278_536_0, i_13_278_573_0, i_13_278_585_0,
    i_13_278_586_0, i_13_278_639_0, i_13_278_640_0, i_13_278_717_0,
    i_13_278_781_0, i_13_278_927_0, i_13_278_1004_0, i_13_278_1064_0,
    i_13_278_1081_0, i_13_278_1116_0, i_13_278_1117_0, i_13_278_1141_0,
    i_13_278_1142_0, i_13_278_1181_0, i_13_278_1296_0, i_13_278_1467_0,
    i_13_278_1468_0, i_13_278_1470_0, i_13_278_1497_0, i_13_278_1503_0,
    i_13_278_1647_0, i_13_278_1648_0, i_13_278_1710_0, i_13_278_1711_0,
    i_13_278_1719_0, i_13_278_1731_0, i_13_278_1782_0, i_13_278_1786_0,
    i_13_278_1791_0, i_13_278_1792_0, i_13_278_1800_0, i_13_278_1802_0,
    i_13_278_1851_0, i_13_278_1989_0, i_13_278_1990_0, i_13_278_1993_0,
    i_13_278_2115_0, i_13_278_2116_0, i_13_278_2259_0, i_13_278_2265_0,
    i_13_278_2290_0, i_13_278_2358_0, i_13_278_2377_0, i_13_278_2379_0,
    i_13_278_2536_0, i_13_278_2667_0, i_13_278_2672_0, i_13_278_2673_0,
    i_13_278_2709_0, i_13_278_2844_0, i_13_278_2845_0, i_13_278_2934_0,
    i_13_278_3036_0, i_13_278_3040_0, i_13_278_3061_0, i_13_278_3123_0,
    i_13_278_3153_0, i_13_278_3215_0, i_13_278_3285_0, i_13_278_3286_0,
    i_13_278_3468_0, i_13_278_3475_0, i_13_278_3550_0, i_13_278_3554_0,
    i_13_278_3581_0, i_13_278_3610_0, i_13_278_3639_0, i_13_278_3818_0,
    i_13_278_3924_0, i_13_278_4008_0, i_13_278_4011_0, i_13_278_4042_0,
    i_13_278_4230_0, i_13_278_4232_0, i_13_278_4302_0, i_13_278_4303_0,
    i_13_278_4390_0, i_13_278_4391_0, i_13_278_4410_0, i_13_278_4411_0;
  output o_13_278_0_0;
  assign o_13_278_0_0 = ~(~i_13_278_1710_0 & ~i_13_278_3285_0);
endmodule



// Benchmark "kernel_13_279" written by ABC on Sun Jul 19 10:49:17 2020

module kernel_13_279 ( 
    i_13_279_46_0, i_13_279_53_0, i_13_279_80_0, i_13_279_91_0,
    i_13_279_114_0, i_13_279_140_0, i_13_279_161_0, i_13_279_171_0,
    i_13_279_178_0, i_13_279_216_0, i_13_279_228_0, i_13_279_237_0,
    i_13_279_251_0, i_13_279_273_0, i_13_279_278_0, i_13_279_441_0,
    i_13_279_455_0, i_13_279_518_0, i_13_279_544_0, i_13_279_562_0,
    i_13_279_576_0, i_13_279_619_0, i_13_279_700_0, i_13_279_723_0,
    i_13_279_885_0, i_13_279_888_0, i_13_279_936_0, i_13_279_944_0,
    i_13_279_945_0, i_13_279_1071_0, i_13_279_1131_0, i_13_279_1262_0,
    i_13_279_1265_0, i_13_279_1329_0, i_13_279_1483_0, i_13_279_1515_0,
    i_13_279_1517_0, i_13_279_1569_0, i_13_279_1626_0, i_13_279_1642_0,
    i_13_279_1643_0, i_13_279_1742_0, i_13_279_1757_0, i_13_279_1777_0,
    i_13_279_1921_0, i_13_279_1948_0, i_13_279_1953_0, i_13_279_2020_0,
    i_13_279_2024_0, i_13_279_2087_0, i_13_279_2185_0, i_13_279_2294_0,
    i_13_279_2302_0, i_13_279_2321_0, i_13_279_2370_0, i_13_279_2424_0,
    i_13_279_2442_0, i_13_279_2446_0, i_13_279_2447_0, i_13_279_2455_0,
    i_13_279_2466_0, i_13_279_2716_0, i_13_279_2742_0, i_13_279_2743_0,
    i_13_279_2744_0, i_13_279_2955_0, i_13_279_2959_0, i_13_279_3042_0,
    i_13_279_3043_0, i_13_279_3208_0, i_13_279_3316_0, i_13_279_3374_0,
    i_13_279_3490_0, i_13_279_3541_0, i_13_279_3546_0, i_13_279_3599_0,
    i_13_279_3604_0, i_13_279_3683_0, i_13_279_3767_0, i_13_279_3769_0,
    i_13_279_3870_0, i_13_279_3904_0, i_13_279_4110_0, i_13_279_4158_0,
    i_13_279_4159_0, i_13_279_4161_0, i_13_279_4166_0, i_13_279_4249_0,
    i_13_279_4321_0, i_13_279_4364_0, i_13_279_4365_0, i_13_279_4432_0,
    i_13_279_4451_0, i_13_279_4454_0, i_13_279_4495_0, i_13_279_4516_0,
    i_13_279_4518_0, i_13_279_4536_0, i_13_279_4542_0, i_13_279_4575_0,
    o_13_279_0_0  );
  input  i_13_279_46_0, i_13_279_53_0, i_13_279_80_0, i_13_279_91_0,
    i_13_279_114_0, i_13_279_140_0, i_13_279_161_0, i_13_279_171_0,
    i_13_279_178_0, i_13_279_216_0, i_13_279_228_0, i_13_279_237_0,
    i_13_279_251_0, i_13_279_273_0, i_13_279_278_0, i_13_279_441_0,
    i_13_279_455_0, i_13_279_518_0, i_13_279_544_0, i_13_279_562_0,
    i_13_279_576_0, i_13_279_619_0, i_13_279_700_0, i_13_279_723_0,
    i_13_279_885_0, i_13_279_888_0, i_13_279_936_0, i_13_279_944_0,
    i_13_279_945_0, i_13_279_1071_0, i_13_279_1131_0, i_13_279_1262_0,
    i_13_279_1265_0, i_13_279_1329_0, i_13_279_1483_0, i_13_279_1515_0,
    i_13_279_1517_0, i_13_279_1569_0, i_13_279_1626_0, i_13_279_1642_0,
    i_13_279_1643_0, i_13_279_1742_0, i_13_279_1757_0, i_13_279_1777_0,
    i_13_279_1921_0, i_13_279_1948_0, i_13_279_1953_0, i_13_279_2020_0,
    i_13_279_2024_0, i_13_279_2087_0, i_13_279_2185_0, i_13_279_2294_0,
    i_13_279_2302_0, i_13_279_2321_0, i_13_279_2370_0, i_13_279_2424_0,
    i_13_279_2442_0, i_13_279_2446_0, i_13_279_2447_0, i_13_279_2455_0,
    i_13_279_2466_0, i_13_279_2716_0, i_13_279_2742_0, i_13_279_2743_0,
    i_13_279_2744_0, i_13_279_2955_0, i_13_279_2959_0, i_13_279_3042_0,
    i_13_279_3043_0, i_13_279_3208_0, i_13_279_3316_0, i_13_279_3374_0,
    i_13_279_3490_0, i_13_279_3541_0, i_13_279_3546_0, i_13_279_3599_0,
    i_13_279_3604_0, i_13_279_3683_0, i_13_279_3767_0, i_13_279_3769_0,
    i_13_279_3870_0, i_13_279_3904_0, i_13_279_4110_0, i_13_279_4158_0,
    i_13_279_4159_0, i_13_279_4161_0, i_13_279_4166_0, i_13_279_4249_0,
    i_13_279_4321_0, i_13_279_4364_0, i_13_279_4365_0, i_13_279_4432_0,
    i_13_279_4451_0, i_13_279_4454_0, i_13_279_4495_0, i_13_279_4516_0,
    i_13_279_4518_0, i_13_279_4536_0, i_13_279_4542_0, i_13_279_4575_0;
  output o_13_279_0_0;
  assign o_13_279_0_0 = ~(~i_13_279_3604_0 & ((~i_13_279_237_0 & ~i_13_279_3316_0) | (~i_13_279_278_0 & ~i_13_279_2743_0 & ~i_13_279_4161_0)));
endmodule



// Benchmark "kernel_13_280" written by ABC on Sun Jul 19 10:49:17 2020

module kernel_13_280 ( 
    i_13_280_32_0, i_13_280_52_0, i_13_280_70_0, i_13_280_71_0,
    i_13_280_79_0, i_13_280_80_0, i_13_280_140_0, i_13_280_176_0,
    i_13_280_230_0, i_13_280_314_0, i_13_280_322_0, i_13_280_323_0,
    i_13_280_377_0, i_13_280_526_0, i_13_280_527_0, i_13_280_557_0,
    i_13_280_589_0, i_13_280_608_0, i_13_280_610_0, i_13_280_647_0,
    i_13_280_674_0, i_13_280_683_0, i_13_280_734_0, i_13_280_853_0,
    i_13_280_986_0, i_13_280_1105_0, i_13_280_1202_0, i_13_280_1222_0,
    i_13_280_1228_0, i_13_280_1229_0, i_13_280_1231_0, i_13_280_1277_0,
    i_13_280_1283_0, i_13_280_1312_0, i_13_280_1313_0, i_13_280_1336_0,
    i_13_280_1394_0, i_13_280_1426_0, i_13_280_1430_0, i_13_280_1510_0,
    i_13_280_1511_0, i_13_280_1664_0, i_13_280_1724_0, i_13_280_1736_0,
    i_13_280_1750_0, i_13_280_1751_0, i_13_280_1781_0, i_13_280_1799_0,
    i_13_280_1843_0, i_13_280_1844_0, i_13_280_1858_0, i_13_280_1886_0,
    i_13_280_1912_0, i_13_280_1931_0, i_13_280_1934_0, i_13_280_1948_0,
    i_13_280_2119_0, i_13_280_2194_0, i_13_280_2195_0, i_13_280_2287_0,
    i_13_280_2426_0, i_13_280_2462_0, i_13_280_2509_0, i_13_280_2552_0,
    i_13_280_2600_0, i_13_280_2722_0, i_13_280_2851_0, i_13_280_2852_0,
    i_13_280_3095_0, i_13_280_3104_0, i_13_280_3118_0, i_13_280_3146_0,
    i_13_280_3271_0, i_13_280_3272_0, i_13_280_3398_0, i_13_280_3418_0,
    i_13_280_3419_0, i_13_280_3433_0, i_13_280_3439_0, i_13_280_3479_0,
    i_13_280_3548_0, i_13_280_3614_0, i_13_280_3743_0, i_13_280_3761_0,
    i_13_280_3769_0, i_13_280_3869_0, i_13_280_3896_0, i_13_280_3932_0,
    i_13_280_3994_0, i_13_280_4040_0, i_13_280_4063_0, i_13_280_4085_0,
    i_13_280_4190_0, i_13_280_4252_0, i_13_280_4297_0, i_13_280_4298_0,
    i_13_280_4382_0, i_13_280_4534_0, i_13_280_4597_0, i_13_280_4598_0,
    o_13_280_0_0  );
  input  i_13_280_32_0, i_13_280_52_0, i_13_280_70_0, i_13_280_71_0,
    i_13_280_79_0, i_13_280_80_0, i_13_280_140_0, i_13_280_176_0,
    i_13_280_230_0, i_13_280_314_0, i_13_280_322_0, i_13_280_323_0,
    i_13_280_377_0, i_13_280_526_0, i_13_280_527_0, i_13_280_557_0,
    i_13_280_589_0, i_13_280_608_0, i_13_280_610_0, i_13_280_647_0,
    i_13_280_674_0, i_13_280_683_0, i_13_280_734_0, i_13_280_853_0,
    i_13_280_986_0, i_13_280_1105_0, i_13_280_1202_0, i_13_280_1222_0,
    i_13_280_1228_0, i_13_280_1229_0, i_13_280_1231_0, i_13_280_1277_0,
    i_13_280_1283_0, i_13_280_1312_0, i_13_280_1313_0, i_13_280_1336_0,
    i_13_280_1394_0, i_13_280_1426_0, i_13_280_1430_0, i_13_280_1510_0,
    i_13_280_1511_0, i_13_280_1664_0, i_13_280_1724_0, i_13_280_1736_0,
    i_13_280_1750_0, i_13_280_1751_0, i_13_280_1781_0, i_13_280_1799_0,
    i_13_280_1843_0, i_13_280_1844_0, i_13_280_1858_0, i_13_280_1886_0,
    i_13_280_1912_0, i_13_280_1931_0, i_13_280_1934_0, i_13_280_1948_0,
    i_13_280_2119_0, i_13_280_2194_0, i_13_280_2195_0, i_13_280_2287_0,
    i_13_280_2426_0, i_13_280_2462_0, i_13_280_2509_0, i_13_280_2552_0,
    i_13_280_2600_0, i_13_280_2722_0, i_13_280_2851_0, i_13_280_2852_0,
    i_13_280_3095_0, i_13_280_3104_0, i_13_280_3118_0, i_13_280_3146_0,
    i_13_280_3271_0, i_13_280_3272_0, i_13_280_3398_0, i_13_280_3418_0,
    i_13_280_3419_0, i_13_280_3433_0, i_13_280_3439_0, i_13_280_3479_0,
    i_13_280_3548_0, i_13_280_3614_0, i_13_280_3743_0, i_13_280_3761_0,
    i_13_280_3769_0, i_13_280_3869_0, i_13_280_3896_0, i_13_280_3932_0,
    i_13_280_3994_0, i_13_280_4040_0, i_13_280_4063_0, i_13_280_4085_0,
    i_13_280_4190_0, i_13_280_4252_0, i_13_280_4297_0, i_13_280_4298_0,
    i_13_280_4382_0, i_13_280_4534_0, i_13_280_4597_0, i_13_280_4598_0;
  output o_13_280_0_0;
  assign o_13_280_0_0 = ~(~i_13_280_674_0 | (~i_13_280_683_0 & ~i_13_280_3104_0) | (~i_13_280_323_0 & ~i_13_280_1510_0 & ~i_13_280_2852_0));
endmodule



// Benchmark "kernel_13_281" written by ABC on Sun Jul 19 10:49:18 2020

module kernel_13_281 ( 
    i_13_281_31_0, i_13_281_58_0, i_13_281_94_0, i_13_281_184_0,
    i_13_281_192_0, i_13_281_310_0, i_13_281_324_0, i_13_281_463_0,
    i_13_281_570_0, i_13_281_575_0, i_13_281_628_0, i_13_281_660_0,
    i_13_281_661_0, i_13_281_714_0, i_13_281_760_0, i_13_281_796_0,
    i_13_281_840_0, i_13_281_858_0, i_13_281_859_0, i_13_281_861_0,
    i_13_281_927_0, i_13_281_1224_0, i_13_281_1225_0, i_13_281_1227_0,
    i_13_281_1228_0, i_13_281_1230_0, i_13_281_1231_0, i_13_281_1254_0,
    i_13_281_1255_0, i_13_281_1345_0, i_13_281_1407_0, i_13_281_1408_0,
    i_13_281_1452_0, i_13_281_1470_0, i_13_281_1488_0, i_13_281_1489_0,
    i_13_281_1507_0, i_13_281_1596_0, i_13_281_1597_0, i_13_281_1632_0,
    i_13_281_1686_0, i_13_281_1687_0, i_13_281_1714_0, i_13_281_1740_0,
    i_13_281_1758_0, i_13_281_1769_0, i_13_281_1854_0, i_13_281_1857_0,
    i_13_281_1858_0, i_13_281_1917_0, i_13_281_1918_0, i_13_281_1930_0,
    i_13_281_1957_0, i_13_281_2011_0, i_13_281_2055_0, i_13_281_2056_0,
    i_13_281_2226_0, i_13_281_2312_0, i_13_281_2425_0, i_13_281_2458_0,
    i_13_281_2568_0, i_13_281_2618_0, i_13_281_2629_0, i_13_281_2676_0,
    i_13_281_2695_0, i_13_281_2856_0, i_13_281_2857_0, i_13_281_2946_0,
    i_13_281_3031_0, i_13_281_3063_0, i_13_281_3064_0, i_13_281_3100_0,
    i_13_281_3114_0, i_13_281_3171_0, i_13_281_3172_0, i_13_281_3204_0,
    i_13_281_3414_0, i_13_281_3421_0, i_13_281_3459_0, i_13_281_3460_0,
    i_13_281_3487_0, i_13_281_3531_0, i_13_281_3532_0, i_13_281_3718_0,
    i_13_281_3802_0, i_13_281_3854_0, i_13_281_3855_0, i_13_281_3856_0,
    i_13_281_3873_0, i_13_281_3874_0, i_13_281_3982_0, i_13_281_4050_0,
    i_13_281_4216_0, i_13_281_4306_0, i_13_281_4341_0, i_13_281_4363_0,
    i_13_281_4396_0, i_13_281_4423_0, i_13_281_4446_0, i_13_281_4507_0,
    o_13_281_0_0  );
  input  i_13_281_31_0, i_13_281_58_0, i_13_281_94_0, i_13_281_184_0,
    i_13_281_192_0, i_13_281_310_0, i_13_281_324_0, i_13_281_463_0,
    i_13_281_570_0, i_13_281_575_0, i_13_281_628_0, i_13_281_660_0,
    i_13_281_661_0, i_13_281_714_0, i_13_281_760_0, i_13_281_796_0,
    i_13_281_840_0, i_13_281_858_0, i_13_281_859_0, i_13_281_861_0,
    i_13_281_927_0, i_13_281_1224_0, i_13_281_1225_0, i_13_281_1227_0,
    i_13_281_1228_0, i_13_281_1230_0, i_13_281_1231_0, i_13_281_1254_0,
    i_13_281_1255_0, i_13_281_1345_0, i_13_281_1407_0, i_13_281_1408_0,
    i_13_281_1452_0, i_13_281_1470_0, i_13_281_1488_0, i_13_281_1489_0,
    i_13_281_1507_0, i_13_281_1596_0, i_13_281_1597_0, i_13_281_1632_0,
    i_13_281_1686_0, i_13_281_1687_0, i_13_281_1714_0, i_13_281_1740_0,
    i_13_281_1758_0, i_13_281_1769_0, i_13_281_1854_0, i_13_281_1857_0,
    i_13_281_1858_0, i_13_281_1917_0, i_13_281_1918_0, i_13_281_1930_0,
    i_13_281_1957_0, i_13_281_2011_0, i_13_281_2055_0, i_13_281_2056_0,
    i_13_281_2226_0, i_13_281_2312_0, i_13_281_2425_0, i_13_281_2458_0,
    i_13_281_2568_0, i_13_281_2618_0, i_13_281_2629_0, i_13_281_2676_0,
    i_13_281_2695_0, i_13_281_2856_0, i_13_281_2857_0, i_13_281_2946_0,
    i_13_281_3031_0, i_13_281_3063_0, i_13_281_3064_0, i_13_281_3100_0,
    i_13_281_3114_0, i_13_281_3171_0, i_13_281_3172_0, i_13_281_3204_0,
    i_13_281_3414_0, i_13_281_3421_0, i_13_281_3459_0, i_13_281_3460_0,
    i_13_281_3487_0, i_13_281_3531_0, i_13_281_3532_0, i_13_281_3718_0,
    i_13_281_3802_0, i_13_281_3854_0, i_13_281_3855_0, i_13_281_3856_0,
    i_13_281_3873_0, i_13_281_3874_0, i_13_281_3982_0, i_13_281_4050_0,
    i_13_281_4216_0, i_13_281_4306_0, i_13_281_4341_0, i_13_281_4363_0,
    i_13_281_4396_0, i_13_281_4423_0, i_13_281_4446_0, i_13_281_4507_0;
  output o_13_281_0_0;
  assign o_13_281_0_0 = ~((~i_13_281_1489_0 & ((~i_13_281_1488_0 & ~i_13_281_3459_0) | (~i_13_281_1452_0 & ~i_13_281_4446_0))) | (~i_13_281_1488_0 & (~i_13_281_1408_0 | ~i_13_281_1858_0)) | (~i_13_281_3855_0 & ((~i_13_281_1407_0 & ~i_13_281_1769_0) | (~i_13_281_2425_0 & i_13_281_4306_0))) | (~i_13_281_3856_0 & (~i_13_281_3171_0 | ~i_13_281_3982_0)) | (~i_13_281_1255_0 & i_13_281_1596_0) | (i_13_281_1597_0 & ~i_13_281_2458_0) | i_13_281_2857_0 | (~i_13_281_1857_0 & ~i_13_281_3459_0 & ~i_13_281_3874_0));
endmodule



// Benchmark "kernel_13_282" written by ABC on Sun Jul 19 10:49:19 2020

module kernel_13_282 ( 
    i_13_282_92_0, i_13_282_96_0, i_13_282_97_0, i_13_282_105_0,
    i_13_282_112_0, i_13_282_175_0, i_13_282_237_0, i_13_282_310_0,
    i_13_282_319_0, i_13_282_519_0, i_13_282_578_0, i_13_282_604_0,
    i_13_282_618_0, i_13_282_643_0, i_13_282_652_0, i_13_282_653_0,
    i_13_282_740_0, i_13_282_771_0, i_13_282_816_0, i_13_282_884_0,
    i_13_282_913_0, i_13_282_921_0, i_13_282_929_0, i_13_282_940_0,
    i_13_282_979_0, i_13_282_1077_0, i_13_282_1084_0, i_13_282_1109_0,
    i_13_282_1280_0, i_13_282_1329_0, i_13_282_1337_0, i_13_282_1441_0,
    i_13_282_1464_0, i_13_282_1480_0, i_13_282_1535_0, i_13_282_1597_0,
    i_13_282_1607_0, i_13_282_1609_0, i_13_282_1667_0, i_13_282_1776_0,
    i_13_282_1786_0, i_13_282_1816_0, i_13_282_1841_0, i_13_282_1894_0,
    i_13_282_1924_0, i_13_282_1948_0, i_13_282_2020_0, i_13_282_2029_0,
    i_13_282_2144_0, i_13_282_2156_0, i_13_282_2173_0, i_13_282_2317_0,
    i_13_282_2425_0, i_13_282_2444_0, i_13_282_2468_0, i_13_282_2498_0,
    i_13_282_2667_0, i_13_282_2749_0, i_13_282_2750_0, i_13_282_2813_0,
    i_13_282_2838_0, i_13_282_2884_0, i_13_282_2940_0, i_13_282_3110_0,
    i_13_282_3155_0, i_13_282_3218_0, i_13_282_3230_0, i_13_282_3268_0,
    i_13_282_3315_0, i_13_282_3350_0, i_13_282_3380_0, i_13_282_3460_0,
    i_13_282_3491_0, i_13_282_3504_0, i_13_282_3522_0, i_13_282_3620_0,
    i_13_282_3649_0, i_13_282_3746_0, i_13_282_3757_0, i_13_282_3824_0,
    i_13_282_3874_0, i_13_282_3910_0, i_13_282_3913_0, i_13_282_4036_0,
    i_13_282_4089_0, i_13_282_4091_0, i_13_282_4124_0, i_13_282_4126_0,
    i_13_282_4187_0, i_13_282_4360_0, i_13_282_4361_0, i_13_282_4366_0,
    i_13_282_4372_0, i_13_282_4396_0, i_13_282_4412_0, i_13_282_4416_0,
    i_13_282_4465_0, i_13_282_4492_0, i_13_282_4519_0, i_13_282_4523_0,
    o_13_282_0_0  );
  input  i_13_282_92_0, i_13_282_96_0, i_13_282_97_0, i_13_282_105_0,
    i_13_282_112_0, i_13_282_175_0, i_13_282_237_0, i_13_282_310_0,
    i_13_282_319_0, i_13_282_519_0, i_13_282_578_0, i_13_282_604_0,
    i_13_282_618_0, i_13_282_643_0, i_13_282_652_0, i_13_282_653_0,
    i_13_282_740_0, i_13_282_771_0, i_13_282_816_0, i_13_282_884_0,
    i_13_282_913_0, i_13_282_921_0, i_13_282_929_0, i_13_282_940_0,
    i_13_282_979_0, i_13_282_1077_0, i_13_282_1084_0, i_13_282_1109_0,
    i_13_282_1280_0, i_13_282_1329_0, i_13_282_1337_0, i_13_282_1441_0,
    i_13_282_1464_0, i_13_282_1480_0, i_13_282_1535_0, i_13_282_1597_0,
    i_13_282_1607_0, i_13_282_1609_0, i_13_282_1667_0, i_13_282_1776_0,
    i_13_282_1786_0, i_13_282_1816_0, i_13_282_1841_0, i_13_282_1894_0,
    i_13_282_1924_0, i_13_282_1948_0, i_13_282_2020_0, i_13_282_2029_0,
    i_13_282_2144_0, i_13_282_2156_0, i_13_282_2173_0, i_13_282_2317_0,
    i_13_282_2425_0, i_13_282_2444_0, i_13_282_2468_0, i_13_282_2498_0,
    i_13_282_2667_0, i_13_282_2749_0, i_13_282_2750_0, i_13_282_2813_0,
    i_13_282_2838_0, i_13_282_2884_0, i_13_282_2940_0, i_13_282_3110_0,
    i_13_282_3155_0, i_13_282_3218_0, i_13_282_3230_0, i_13_282_3268_0,
    i_13_282_3315_0, i_13_282_3350_0, i_13_282_3380_0, i_13_282_3460_0,
    i_13_282_3491_0, i_13_282_3504_0, i_13_282_3522_0, i_13_282_3620_0,
    i_13_282_3649_0, i_13_282_3746_0, i_13_282_3757_0, i_13_282_3824_0,
    i_13_282_3874_0, i_13_282_3910_0, i_13_282_3913_0, i_13_282_4036_0,
    i_13_282_4089_0, i_13_282_4091_0, i_13_282_4124_0, i_13_282_4126_0,
    i_13_282_4187_0, i_13_282_4360_0, i_13_282_4361_0, i_13_282_4366_0,
    i_13_282_4372_0, i_13_282_4396_0, i_13_282_4412_0, i_13_282_4416_0,
    i_13_282_4465_0, i_13_282_4492_0, i_13_282_4519_0, i_13_282_4523_0;
  output o_13_282_0_0;
  assign o_13_282_0_0 = 0;
endmodule



// Benchmark "kernel_13_283" written by ABC on Sun Jul 19 10:49:20 2020

module kernel_13_283 ( 
    i_13_283_27_0, i_13_283_28_0, i_13_283_102_0, i_13_283_103_0,
    i_13_283_126_0, i_13_283_153_0, i_13_283_154_0, i_13_283_190_0,
    i_13_283_282_0, i_13_283_585_0, i_13_283_586_0, i_13_283_669_0,
    i_13_283_846_0, i_13_283_856_0, i_13_283_914_0, i_13_283_949_0,
    i_13_283_1080_0, i_13_283_1081_0, i_13_283_1206_0, i_13_283_1305_0,
    i_13_283_1341_0, i_13_283_1342_0, i_13_283_1422_0, i_13_283_1434_0,
    i_13_283_1441_0, i_13_283_1443_0, i_13_283_1467_0, i_13_283_1504_0,
    i_13_283_1540_0, i_13_283_1632_0, i_13_283_1678_0, i_13_283_1750_0,
    i_13_283_1782_0, i_13_283_1803_0, i_13_283_1810_0, i_13_283_1839_0,
    i_13_283_1840_0, i_13_283_1926_0, i_13_283_1927_0, i_13_283_1999_0,
    i_13_283_2001_0, i_13_283_2052_0, i_13_283_2053_0, i_13_283_2054_0,
    i_13_283_2109_0, i_13_283_2119_0, i_13_283_2197_0, i_13_283_2259_0,
    i_13_283_2277_0, i_13_283_2278_0, i_13_283_2341_0, i_13_283_2407_0,
    i_13_283_2433_0, i_13_283_2443_0, i_13_283_2512_0, i_13_283_2541_0,
    i_13_283_2542_0, i_13_283_2550_0, i_13_283_2614_0, i_13_283_2619_0,
    i_13_283_2629_0, i_13_283_2686_0, i_13_283_2709_0, i_13_283_2710_0,
    i_13_283_2853_0, i_13_283_2854_0, i_13_283_2858_0, i_13_283_2917_0,
    i_13_283_2946_0, i_13_283_3061_0, i_13_283_3150_0, i_13_283_3205_0,
    i_13_283_3307_0, i_13_283_3315_0, i_13_283_3415_0, i_13_283_3432_0,
    i_13_283_3528_0, i_13_283_3532_0, i_13_283_3610_0, i_13_283_3627_0,
    i_13_283_3730_0, i_13_283_3862_0, i_13_283_3979_0, i_13_283_4014_0,
    i_13_283_4050_0, i_13_283_4059_0, i_13_283_4087_0, i_13_283_4114_0,
    i_13_283_4230_0, i_13_283_4231_0, i_13_283_4248_0, i_13_283_4257_0,
    i_13_283_4268_0, i_13_283_4270_0, i_13_283_4338_0, i_13_283_4342_0,
    i_13_283_4392_0, i_13_283_4393_0, i_13_283_4394_0, i_13_283_4536_0,
    o_13_283_0_0  );
  input  i_13_283_27_0, i_13_283_28_0, i_13_283_102_0, i_13_283_103_0,
    i_13_283_126_0, i_13_283_153_0, i_13_283_154_0, i_13_283_190_0,
    i_13_283_282_0, i_13_283_585_0, i_13_283_586_0, i_13_283_669_0,
    i_13_283_846_0, i_13_283_856_0, i_13_283_914_0, i_13_283_949_0,
    i_13_283_1080_0, i_13_283_1081_0, i_13_283_1206_0, i_13_283_1305_0,
    i_13_283_1341_0, i_13_283_1342_0, i_13_283_1422_0, i_13_283_1434_0,
    i_13_283_1441_0, i_13_283_1443_0, i_13_283_1467_0, i_13_283_1504_0,
    i_13_283_1540_0, i_13_283_1632_0, i_13_283_1678_0, i_13_283_1750_0,
    i_13_283_1782_0, i_13_283_1803_0, i_13_283_1810_0, i_13_283_1839_0,
    i_13_283_1840_0, i_13_283_1926_0, i_13_283_1927_0, i_13_283_1999_0,
    i_13_283_2001_0, i_13_283_2052_0, i_13_283_2053_0, i_13_283_2054_0,
    i_13_283_2109_0, i_13_283_2119_0, i_13_283_2197_0, i_13_283_2259_0,
    i_13_283_2277_0, i_13_283_2278_0, i_13_283_2341_0, i_13_283_2407_0,
    i_13_283_2433_0, i_13_283_2443_0, i_13_283_2512_0, i_13_283_2541_0,
    i_13_283_2542_0, i_13_283_2550_0, i_13_283_2614_0, i_13_283_2619_0,
    i_13_283_2629_0, i_13_283_2686_0, i_13_283_2709_0, i_13_283_2710_0,
    i_13_283_2853_0, i_13_283_2854_0, i_13_283_2858_0, i_13_283_2917_0,
    i_13_283_2946_0, i_13_283_3061_0, i_13_283_3150_0, i_13_283_3205_0,
    i_13_283_3307_0, i_13_283_3315_0, i_13_283_3415_0, i_13_283_3432_0,
    i_13_283_3528_0, i_13_283_3532_0, i_13_283_3610_0, i_13_283_3627_0,
    i_13_283_3730_0, i_13_283_3862_0, i_13_283_3979_0, i_13_283_4014_0,
    i_13_283_4050_0, i_13_283_4059_0, i_13_283_4087_0, i_13_283_4114_0,
    i_13_283_4230_0, i_13_283_4231_0, i_13_283_4248_0, i_13_283_4257_0,
    i_13_283_4268_0, i_13_283_4270_0, i_13_283_4338_0, i_13_283_4342_0,
    i_13_283_4392_0, i_13_283_4393_0, i_13_283_4394_0, i_13_283_4536_0;
  output o_13_283_0_0;
  assign o_13_283_0_0 = ~(~i_13_283_2710_0 | (~i_13_283_1342_0 & ~i_13_283_4230_0) | (~i_13_283_1504_0 & ~i_13_283_2854_0 & ~i_13_283_4392_0));
endmodule



// Benchmark "kernel_13_284" written by ABC on Sun Jul 19 10:49:20 2020

module kernel_13_284 ( 
    i_13_284_39_0, i_13_284_40_0, i_13_284_66_0, i_13_284_125_0,
    i_13_284_178_0, i_13_284_268_0, i_13_284_308_0, i_13_284_310_0,
    i_13_284_318_0, i_13_284_319_0, i_13_284_463_0, i_13_284_466_0,
    i_13_284_489_0, i_13_284_536_0, i_13_284_589_0, i_13_284_591_0,
    i_13_284_592_0, i_13_284_625_0, i_13_284_640_0, i_13_284_645_0,
    i_13_284_646_0, i_13_284_690_0, i_13_284_691_0, i_13_284_763_0,
    i_13_284_817_0, i_13_284_841_0, i_13_284_933_0, i_13_284_1122_0,
    i_13_284_1228_0, i_13_284_1284_0, i_13_284_1347_0, i_13_284_1348_0,
    i_13_284_1411_0, i_13_284_1437_0, i_13_284_1542_0, i_13_284_1596_0,
    i_13_284_1597_0, i_13_284_1599_0, i_13_284_1671_0, i_13_284_1754_0,
    i_13_284_1852_0, i_13_284_1941_0, i_13_284_1959_0, i_13_284_2001_0,
    i_13_284_2002_0, i_13_284_2058_0, i_13_284_2059_0, i_13_284_2139_0,
    i_13_284_2181_0, i_13_284_2182_0, i_13_284_2193_0, i_13_284_2265_0,
    i_13_284_2275_0, i_13_284_2283_0, i_13_284_2284_0, i_13_284_2410_0,
    i_13_284_2554_0, i_13_284_2614_0, i_13_284_2617_0, i_13_284_2652_0,
    i_13_284_2653_0, i_13_284_2673_0, i_13_284_2679_0, i_13_284_2697_0,
    i_13_284_2698_0, i_13_284_2760_0, i_13_284_2823_0, i_13_284_2856_0,
    i_13_284_2859_0, i_13_284_2860_0, i_13_284_2997_0, i_13_284_3004_0,
    i_13_284_3212_0, i_13_284_3275_0, i_13_284_3372_0, i_13_284_3390_0,
    i_13_284_3391_0, i_13_284_3392_0, i_13_284_3415_0, i_13_284_3487_0,
    i_13_284_3532_0, i_13_284_3535_0, i_13_284_3616_0, i_13_284_3721_0,
    i_13_284_3877_0, i_13_284_3930_0, i_13_284_4034_0, i_13_284_4035_0,
    i_13_284_4207_0, i_13_284_4218_0, i_13_284_4308_0, i_13_284_4309_0,
    i_13_284_4341_0, i_13_284_4363_0, i_13_284_4372_0, i_13_284_4399_0,
    i_13_284_4540_0, i_13_284_4543_0, i_13_284_4585_0, i_13_284_4597_0,
    o_13_284_0_0  );
  input  i_13_284_39_0, i_13_284_40_0, i_13_284_66_0, i_13_284_125_0,
    i_13_284_178_0, i_13_284_268_0, i_13_284_308_0, i_13_284_310_0,
    i_13_284_318_0, i_13_284_319_0, i_13_284_463_0, i_13_284_466_0,
    i_13_284_489_0, i_13_284_536_0, i_13_284_589_0, i_13_284_591_0,
    i_13_284_592_0, i_13_284_625_0, i_13_284_640_0, i_13_284_645_0,
    i_13_284_646_0, i_13_284_690_0, i_13_284_691_0, i_13_284_763_0,
    i_13_284_817_0, i_13_284_841_0, i_13_284_933_0, i_13_284_1122_0,
    i_13_284_1228_0, i_13_284_1284_0, i_13_284_1347_0, i_13_284_1348_0,
    i_13_284_1411_0, i_13_284_1437_0, i_13_284_1542_0, i_13_284_1596_0,
    i_13_284_1597_0, i_13_284_1599_0, i_13_284_1671_0, i_13_284_1754_0,
    i_13_284_1852_0, i_13_284_1941_0, i_13_284_1959_0, i_13_284_2001_0,
    i_13_284_2002_0, i_13_284_2058_0, i_13_284_2059_0, i_13_284_2139_0,
    i_13_284_2181_0, i_13_284_2182_0, i_13_284_2193_0, i_13_284_2265_0,
    i_13_284_2275_0, i_13_284_2283_0, i_13_284_2284_0, i_13_284_2410_0,
    i_13_284_2554_0, i_13_284_2614_0, i_13_284_2617_0, i_13_284_2652_0,
    i_13_284_2653_0, i_13_284_2673_0, i_13_284_2679_0, i_13_284_2697_0,
    i_13_284_2698_0, i_13_284_2760_0, i_13_284_2823_0, i_13_284_2856_0,
    i_13_284_2859_0, i_13_284_2860_0, i_13_284_2997_0, i_13_284_3004_0,
    i_13_284_3212_0, i_13_284_3275_0, i_13_284_3372_0, i_13_284_3390_0,
    i_13_284_3391_0, i_13_284_3392_0, i_13_284_3415_0, i_13_284_3487_0,
    i_13_284_3532_0, i_13_284_3535_0, i_13_284_3616_0, i_13_284_3721_0,
    i_13_284_3877_0, i_13_284_3930_0, i_13_284_4034_0, i_13_284_4035_0,
    i_13_284_4207_0, i_13_284_4218_0, i_13_284_4308_0, i_13_284_4309_0,
    i_13_284_4341_0, i_13_284_4363_0, i_13_284_4372_0, i_13_284_4399_0,
    i_13_284_4540_0, i_13_284_4543_0, i_13_284_4585_0, i_13_284_4597_0;
  output o_13_284_0_0;
  assign o_13_284_0_0 = ~((i_13_284_2614_0 & ((i_13_284_763_0 & ~i_13_284_3390_0) | (~i_13_284_2139_0 & ~i_13_284_3212_0 & ~i_13_284_4309_0))) | (~i_13_284_1596_0 & (i_13_284_489_0 | ~i_13_284_2059_0 | (~i_13_284_2856_0 & i_13_284_3535_0))) | (~i_13_284_2760_0 & ~i_13_284_3391_0) | (~i_13_284_2284_0 & ~i_13_284_2698_0 & ~i_13_284_3930_0));
endmodule



// Benchmark "kernel_13_285" written by ABC on Sun Jul 19 10:49:21 2020

module kernel_13_285 ( 
    i_13_285_25_0, i_13_285_40_0, i_13_285_67_0, i_13_285_70_0,
    i_13_285_87_0, i_13_285_276_0, i_13_285_310_0, i_13_285_319_0,
    i_13_285_382_0, i_13_285_411_0, i_13_285_492_0, i_13_285_520_0,
    i_13_285_609_0, i_13_285_628_0, i_13_285_660_0, i_13_285_663_0,
    i_13_285_744_0, i_13_285_746_0, i_13_285_805_0, i_13_285_835_0,
    i_13_285_912_0, i_13_285_934_0, i_13_285_939_0, i_13_285_1020_0,
    i_13_285_1021_0, i_13_285_1074_0, i_13_285_1086_0, i_13_285_1087_0,
    i_13_285_1095_0, i_13_285_1096_0, i_13_285_1111_0, i_13_285_1147_0,
    i_13_285_1156_0, i_13_285_1330_0, i_13_285_1403_0, i_13_285_1470_0,
    i_13_285_1474_0, i_13_285_1597_0, i_13_285_1716_0, i_13_285_1735_0,
    i_13_285_1744_0, i_13_285_1750_0, i_13_285_1767_0, i_13_285_1795_0,
    i_13_285_1798_0, i_13_285_1857_0, i_13_285_1965_0, i_13_285_2022_0,
    i_13_285_2023_0, i_13_285_2028_0, i_13_285_2059_0, i_13_285_2060_0,
    i_13_285_2199_0, i_13_285_2235_0, i_13_285_2454_0, i_13_285_2472_0,
    i_13_285_2473_0, i_13_285_2500_0, i_13_285_2617_0, i_13_285_2676_0,
    i_13_285_2715_0, i_13_285_2733_0, i_13_285_2743_0, i_13_285_2769_0,
    i_13_285_2884_0, i_13_285_3030_0, i_13_285_3031_0, i_13_285_3076_0,
    i_13_285_3093_0, i_13_285_3121_0, i_13_285_3144_0, i_13_285_3264_0,
    i_13_285_3265_0, i_13_285_3306_0, i_13_285_3355_0, i_13_285_3435_0,
    i_13_285_3453_0, i_13_285_3454_0, i_13_285_3486_0, i_13_285_3527_0,
    i_13_285_3549_0, i_13_285_3576_0, i_13_285_3613_0, i_13_285_3741_0,
    i_13_285_3742_0, i_13_285_3822_0, i_13_285_3823_0, i_13_285_3927_0,
    i_13_285_3981_0, i_13_285_4092_0, i_13_285_4093_0, i_13_285_4119_0,
    i_13_285_4161_0, i_13_285_4164_0, i_13_285_4165_0, i_13_285_4254_0,
    i_13_285_4417_0, i_13_285_4461_0, i_13_285_4596_0, i_13_285_4606_0,
    o_13_285_0_0  );
  input  i_13_285_25_0, i_13_285_40_0, i_13_285_67_0, i_13_285_70_0,
    i_13_285_87_0, i_13_285_276_0, i_13_285_310_0, i_13_285_319_0,
    i_13_285_382_0, i_13_285_411_0, i_13_285_492_0, i_13_285_520_0,
    i_13_285_609_0, i_13_285_628_0, i_13_285_660_0, i_13_285_663_0,
    i_13_285_744_0, i_13_285_746_0, i_13_285_805_0, i_13_285_835_0,
    i_13_285_912_0, i_13_285_934_0, i_13_285_939_0, i_13_285_1020_0,
    i_13_285_1021_0, i_13_285_1074_0, i_13_285_1086_0, i_13_285_1087_0,
    i_13_285_1095_0, i_13_285_1096_0, i_13_285_1111_0, i_13_285_1147_0,
    i_13_285_1156_0, i_13_285_1330_0, i_13_285_1403_0, i_13_285_1470_0,
    i_13_285_1474_0, i_13_285_1597_0, i_13_285_1716_0, i_13_285_1735_0,
    i_13_285_1744_0, i_13_285_1750_0, i_13_285_1767_0, i_13_285_1795_0,
    i_13_285_1798_0, i_13_285_1857_0, i_13_285_1965_0, i_13_285_2022_0,
    i_13_285_2023_0, i_13_285_2028_0, i_13_285_2059_0, i_13_285_2060_0,
    i_13_285_2199_0, i_13_285_2235_0, i_13_285_2454_0, i_13_285_2472_0,
    i_13_285_2473_0, i_13_285_2500_0, i_13_285_2617_0, i_13_285_2676_0,
    i_13_285_2715_0, i_13_285_2733_0, i_13_285_2743_0, i_13_285_2769_0,
    i_13_285_2884_0, i_13_285_3030_0, i_13_285_3031_0, i_13_285_3076_0,
    i_13_285_3093_0, i_13_285_3121_0, i_13_285_3144_0, i_13_285_3264_0,
    i_13_285_3265_0, i_13_285_3306_0, i_13_285_3355_0, i_13_285_3435_0,
    i_13_285_3453_0, i_13_285_3454_0, i_13_285_3486_0, i_13_285_3527_0,
    i_13_285_3549_0, i_13_285_3576_0, i_13_285_3613_0, i_13_285_3741_0,
    i_13_285_3742_0, i_13_285_3822_0, i_13_285_3823_0, i_13_285_3927_0,
    i_13_285_3981_0, i_13_285_4092_0, i_13_285_4093_0, i_13_285_4119_0,
    i_13_285_4161_0, i_13_285_4164_0, i_13_285_4165_0, i_13_285_4254_0,
    i_13_285_4417_0, i_13_285_4461_0, i_13_285_4596_0, i_13_285_4606_0;
  output o_13_285_0_0;
  assign o_13_285_0_0 = ~(~i_13_285_3741_0 | ~i_13_285_3454_0 | (~i_13_285_934_0 & ~i_13_285_4165_0));
endmodule



// Benchmark "kernel_13_286" written by ABC on Sun Jul 19 10:49:22 2020

module kernel_13_286 ( 
    i_13_286_24_0, i_13_286_87_0, i_13_286_133_0, i_13_286_165_0,
    i_13_286_168_0, i_13_286_183_0, i_13_286_192_0, i_13_286_318_0,
    i_13_286_319_0, i_13_286_334_0, i_13_286_336_0, i_13_286_447_0,
    i_13_286_468_0, i_13_286_469_0, i_13_286_492_0, i_13_286_516_0,
    i_13_286_594_0, i_13_286_615_0, i_13_286_619_0, i_13_286_627_0,
    i_13_286_628_0, i_13_286_648_0, i_13_286_762_0, i_13_286_945_0,
    i_13_286_946_0, i_13_286_951_0, i_13_286_999_0, i_13_286_1018_0,
    i_13_286_1095_0, i_13_286_1227_0, i_13_286_1257_0, i_13_286_1314_0,
    i_13_286_1482_0, i_13_286_1483_0, i_13_286_1495_0, i_13_286_1525_0,
    i_13_286_1537_0, i_13_286_1542_0, i_13_286_1548_0, i_13_286_1620_0,
    i_13_286_1626_0, i_13_286_1627_0, i_13_286_1633_0, i_13_286_1723_0,
    i_13_286_1725_0, i_13_286_1734_0, i_13_286_1770_0, i_13_286_1806_0,
    i_13_286_1924_0, i_13_286_1941_0, i_13_286_1959_0, i_13_286_2002_0,
    i_13_286_2052_0, i_13_286_2103_0, i_13_286_2142_0, i_13_286_2238_0,
    i_13_286_2258_0, i_13_286_2364_0, i_13_286_2382_0, i_13_286_2445_0,
    i_13_286_2538_0, i_13_286_2727_0, i_13_286_2730_0, i_13_286_2850_0,
    i_13_286_2940_0, i_13_286_2985_0, i_13_286_2998_0, i_13_286_3021_0,
    i_13_286_3075_0, i_13_286_3220_0, i_13_286_3240_0, i_13_286_3241_0,
    i_13_286_3246_0, i_13_286_3264_0, i_13_286_3265_0, i_13_286_3282_0,
    i_13_286_3310_0, i_13_286_3345_0, i_13_286_3355_0, i_13_286_3528_0,
    i_13_286_3534_0, i_13_286_3535_0, i_13_286_3639_0, i_13_286_3702_0,
    i_13_286_3733_0, i_13_286_3759_0, i_13_286_3877_0, i_13_286_3889_0,
    i_13_286_3891_0, i_13_286_3892_0, i_13_286_3984_0, i_13_286_3985_0,
    i_13_286_4018_0, i_13_286_4044_0, i_13_286_4137_0, i_13_286_4185_0,
    i_13_286_4272_0, i_13_286_4294_0, i_13_286_4296_0, i_13_286_4425_0,
    o_13_286_0_0  );
  input  i_13_286_24_0, i_13_286_87_0, i_13_286_133_0, i_13_286_165_0,
    i_13_286_168_0, i_13_286_183_0, i_13_286_192_0, i_13_286_318_0,
    i_13_286_319_0, i_13_286_334_0, i_13_286_336_0, i_13_286_447_0,
    i_13_286_468_0, i_13_286_469_0, i_13_286_492_0, i_13_286_516_0,
    i_13_286_594_0, i_13_286_615_0, i_13_286_619_0, i_13_286_627_0,
    i_13_286_628_0, i_13_286_648_0, i_13_286_762_0, i_13_286_945_0,
    i_13_286_946_0, i_13_286_951_0, i_13_286_999_0, i_13_286_1018_0,
    i_13_286_1095_0, i_13_286_1227_0, i_13_286_1257_0, i_13_286_1314_0,
    i_13_286_1482_0, i_13_286_1483_0, i_13_286_1495_0, i_13_286_1525_0,
    i_13_286_1537_0, i_13_286_1542_0, i_13_286_1548_0, i_13_286_1620_0,
    i_13_286_1626_0, i_13_286_1627_0, i_13_286_1633_0, i_13_286_1723_0,
    i_13_286_1725_0, i_13_286_1734_0, i_13_286_1770_0, i_13_286_1806_0,
    i_13_286_1924_0, i_13_286_1941_0, i_13_286_1959_0, i_13_286_2002_0,
    i_13_286_2052_0, i_13_286_2103_0, i_13_286_2142_0, i_13_286_2238_0,
    i_13_286_2258_0, i_13_286_2364_0, i_13_286_2382_0, i_13_286_2445_0,
    i_13_286_2538_0, i_13_286_2727_0, i_13_286_2730_0, i_13_286_2850_0,
    i_13_286_2940_0, i_13_286_2985_0, i_13_286_2998_0, i_13_286_3021_0,
    i_13_286_3075_0, i_13_286_3220_0, i_13_286_3240_0, i_13_286_3241_0,
    i_13_286_3246_0, i_13_286_3264_0, i_13_286_3265_0, i_13_286_3282_0,
    i_13_286_3310_0, i_13_286_3345_0, i_13_286_3355_0, i_13_286_3528_0,
    i_13_286_3534_0, i_13_286_3535_0, i_13_286_3639_0, i_13_286_3702_0,
    i_13_286_3733_0, i_13_286_3759_0, i_13_286_3877_0, i_13_286_3889_0,
    i_13_286_3891_0, i_13_286_3892_0, i_13_286_3984_0, i_13_286_3985_0,
    i_13_286_4018_0, i_13_286_4044_0, i_13_286_4137_0, i_13_286_4185_0,
    i_13_286_4272_0, i_13_286_4294_0, i_13_286_4296_0, i_13_286_4425_0;
  output o_13_286_0_0;
  assign o_13_286_0_0 = ~((~i_13_286_3984_0 & ((~i_13_286_615_0 & ~i_13_286_1482_0 & ~i_13_286_1806_0) | (~i_13_286_2445_0 & ~i_13_286_3534_0 & ~i_13_286_3877_0))) | (~i_13_286_492_0 & i_13_286_2002_0) | (~i_13_286_447_0 & ~i_13_286_1627_0 & ~i_13_286_2850_0));
endmodule



// Benchmark "kernel_13_287" written by ABC on Sun Jul 19 10:49:23 2020

module kernel_13_287 ( 
    i_13_287_40_0, i_13_287_53_0, i_13_287_95_0, i_13_287_96_0,
    i_13_287_143_0, i_13_287_274_0, i_13_287_287_0, i_13_287_341_0,
    i_13_287_476_0, i_13_287_521_0, i_13_287_529_0, i_13_287_565_0,
    i_13_287_592_0, i_13_287_644_0, i_13_287_646_0, i_13_287_647_0,
    i_13_287_688_0, i_13_287_689_0, i_13_287_691_0, i_13_287_692_0,
    i_13_287_797_0, i_13_287_980_0, i_13_287_1025_0, i_13_287_1101_0,
    i_13_287_1121_0, i_13_287_1123_0, i_13_287_1124_0, i_13_287_1204_0,
    i_13_287_1256_0, i_13_287_1273_0, i_13_287_1277_0, i_13_287_1384_0,
    i_13_287_1391_0, i_13_287_1444_0, i_13_287_1445_0, i_13_287_1465_0,
    i_13_287_1484_0, i_13_287_1489_0, i_13_287_1502_0, i_13_287_1627_0,
    i_13_287_1643_0, i_13_287_1714_0, i_13_287_1715_0, i_13_287_1885_0,
    i_13_287_1886_0, i_13_287_1888_0, i_13_287_1991_0, i_13_287_2059_0,
    i_13_287_2140_0, i_13_287_2267_0, i_13_287_2285_0, i_13_287_2354_0,
    i_13_287_2428_0, i_13_287_2447_0, i_13_287_2464_0, i_13_287_2497_0,
    i_13_287_2506_0, i_13_287_2509_0, i_13_287_2510_0, i_13_287_2511_0,
    i_13_287_2533_0, i_13_287_2542_0, i_13_287_2569_0, i_13_287_2648_0,
    i_13_287_2650_0, i_13_287_2651_0, i_13_287_2653_0, i_13_287_2654_0,
    i_13_287_2677_0, i_13_287_2752_0, i_13_287_2753_0, i_13_287_2825_0,
    i_13_287_2848_0, i_13_287_2849_0, i_13_287_2920_0, i_13_287_3004_0,
    i_13_287_3126_0, i_13_287_3146_0, i_13_287_3217_0, i_13_287_3391_0,
    i_13_287_3392_0, i_13_287_3424_0, i_13_287_3445_0, i_13_287_3550_0,
    i_13_287_3794_0, i_13_287_3874_0, i_13_287_3914_0, i_13_287_3982_0,
    i_13_287_3991_0, i_13_287_3992_0, i_13_287_3995_0, i_13_287_4057_0,
    i_13_287_4081_0, i_13_287_4085_0, i_13_287_4153_0, i_13_287_4162_0,
    i_13_287_4318_0, i_13_287_4372_0, i_13_287_4381_0, i_13_287_4444_0,
    o_13_287_0_0  );
  input  i_13_287_40_0, i_13_287_53_0, i_13_287_95_0, i_13_287_96_0,
    i_13_287_143_0, i_13_287_274_0, i_13_287_287_0, i_13_287_341_0,
    i_13_287_476_0, i_13_287_521_0, i_13_287_529_0, i_13_287_565_0,
    i_13_287_592_0, i_13_287_644_0, i_13_287_646_0, i_13_287_647_0,
    i_13_287_688_0, i_13_287_689_0, i_13_287_691_0, i_13_287_692_0,
    i_13_287_797_0, i_13_287_980_0, i_13_287_1025_0, i_13_287_1101_0,
    i_13_287_1121_0, i_13_287_1123_0, i_13_287_1124_0, i_13_287_1204_0,
    i_13_287_1256_0, i_13_287_1273_0, i_13_287_1277_0, i_13_287_1384_0,
    i_13_287_1391_0, i_13_287_1444_0, i_13_287_1445_0, i_13_287_1465_0,
    i_13_287_1484_0, i_13_287_1489_0, i_13_287_1502_0, i_13_287_1627_0,
    i_13_287_1643_0, i_13_287_1714_0, i_13_287_1715_0, i_13_287_1885_0,
    i_13_287_1886_0, i_13_287_1888_0, i_13_287_1991_0, i_13_287_2059_0,
    i_13_287_2140_0, i_13_287_2267_0, i_13_287_2285_0, i_13_287_2354_0,
    i_13_287_2428_0, i_13_287_2447_0, i_13_287_2464_0, i_13_287_2497_0,
    i_13_287_2506_0, i_13_287_2509_0, i_13_287_2510_0, i_13_287_2511_0,
    i_13_287_2533_0, i_13_287_2542_0, i_13_287_2569_0, i_13_287_2648_0,
    i_13_287_2650_0, i_13_287_2651_0, i_13_287_2653_0, i_13_287_2654_0,
    i_13_287_2677_0, i_13_287_2752_0, i_13_287_2753_0, i_13_287_2825_0,
    i_13_287_2848_0, i_13_287_2849_0, i_13_287_2920_0, i_13_287_3004_0,
    i_13_287_3126_0, i_13_287_3146_0, i_13_287_3217_0, i_13_287_3391_0,
    i_13_287_3392_0, i_13_287_3424_0, i_13_287_3445_0, i_13_287_3550_0,
    i_13_287_3794_0, i_13_287_3874_0, i_13_287_3914_0, i_13_287_3982_0,
    i_13_287_3991_0, i_13_287_3992_0, i_13_287_3995_0, i_13_287_4057_0,
    i_13_287_4081_0, i_13_287_4085_0, i_13_287_4153_0, i_13_287_4162_0,
    i_13_287_4318_0, i_13_287_4372_0, i_13_287_4381_0, i_13_287_4444_0;
  output o_13_287_0_0;
  assign o_13_287_0_0 = ~((~i_13_287_2140_0 & i_13_287_3550_0) | (~i_13_287_688_0 & ~i_13_287_2848_0) | (~i_13_287_1121_0 & ~i_13_287_1124_0) | (~i_13_287_287_0 & ~i_13_287_1888_0 & ~i_13_287_4381_0));
endmodule



// Benchmark "kernel_13_288" written by ABC on Sun Jul 19 10:49:23 2020

module kernel_13_288 ( 
    i_13_288_49_0, i_13_288_167_0, i_13_288_173_0, i_13_288_190_0,
    i_13_288_211_0, i_13_288_255_0, i_13_288_280_0, i_13_288_283_0,
    i_13_288_314_0, i_13_288_379_0, i_13_288_380_0, i_13_288_472_0,
    i_13_288_526_0, i_13_288_530_0, i_13_288_571_0, i_13_288_640_0,
    i_13_288_641_0, i_13_288_659_0, i_13_288_661_0, i_13_288_662_0,
    i_13_288_668_0, i_13_288_676_0, i_13_288_677_0, i_13_288_810_0,
    i_13_288_928_0, i_13_288_941_0, i_13_288_992_0, i_13_288_1063_0,
    i_13_288_1081_0, i_13_288_1082_0, i_13_288_1306_0, i_13_288_1307_0,
    i_13_288_1411_0, i_13_288_1444_0, i_13_288_1498_0, i_13_288_1499_0,
    i_13_288_1504_0, i_13_288_1505_0, i_13_288_1633_0, i_13_288_1636_0,
    i_13_288_1730_0, i_13_288_1783_0, i_13_288_1801_0, i_13_288_1838_0,
    i_13_288_1846_0, i_13_288_1880_0, i_13_288_1927_0, i_13_288_1942_0,
    i_13_288_2054_0, i_13_288_2170_0, i_13_288_2315_0, i_13_288_2425_0,
    i_13_288_2431_0, i_13_288_2432_0, i_13_288_2674_0, i_13_288_2923_0,
    i_13_288_3107_0, i_13_288_3142_0, i_13_288_3143_0, i_13_288_3242_0,
    i_13_288_3267_0, i_13_288_3269_0, i_13_288_3271_0, i_13_288_3371_0,
    i_13_288_3420_0, i_13_288_3421_0, i_13_288_3422_0, i_13_288_3424_0,
    i_13_288_3425_0, i_13_288_3545_0, i_13_288_3646_0, i_13_288_3730_0,
    i_13_288_3731_0, i_13_288_3767_0, i_13_288_3817_0, i_13_288_3818_0,
    i_13_288_3925_0, i_13_288_3971_0, i_13_288_3989_0, i_13_288_4015_0,
    i_13_288_4016_0, i_13_288_4018_0, i_13_288_4019_0, i_13_288_4044_0,
    i_13_288_4060_0, i_13_288_4061_0, i_13_288_4078_0, i_13_288_4214_0,
    i_13_288_4249_0, i_13_288_4250_0, i_13_288_4253_0, i_13_288_4261_0,
    i_13_288_4313_0, i_13_288_4340_0, i_13_288_4351_0, i_13_288_4430_0,
    i_13_288_4556_0, i_13_288_4558_0, i_13_288_4567_0, i_13_288_4591_0,
    o_13_288_0_0  );
  input  i_13_288_49_0, i_13_288_167_0, i_13_288_173_0, i_13_288_190_0,
    i_13_288_211_0, i_13_288_255_0, i_13_288_280_0, i_13_288_283_0,
    i_13_288_314_0, i_13_288_379_0, i_13_288_380_0, i_13_288_472_0,
    i_13_288_526_0, i_13_288_530_0, i_13_288_571_0, i_13_288_640_0,
    i_13_288_641_0, i_13_288_659_0, i_13_288_661_0, i_13_288_662_0,
    i_13_288_668_0, i_13_288_676_0, i_13_288_677_0, i_13_288_810_0,
    i_13_288_928_0, i_13_288_941_0, i_13_288_992_0, i_13_288_1063_0,
    i_13_288_1081_0, i_13_288_1082_0, i_13_288_1306_0, i_13_288_1307_0,
    i_13_288_1411_0, i_13_288_1444_0, i_13_288_1498_0, i_13_288_1499_0,
    i_13_288_1504_0, i_13_288_1505_0, i_13_288_1633_0, i_13_288_1636_0,
    i_13_288_1730_0, i_13_288_1783_0, i_13_288_1801_0, i_13_288_1838_0,
    i_13_288_1846_0, i_13_288_1880_0, i_13_288_1927_0, i_13_288_1942_0,
    i_13_288_2054_0, i_13_288_2170_0, i_13_288_2315_0, i_13_288_2425_0,
    i_13_288_2431_0, i_13_288_2432_0, i_13_288_2674_0, i_13_288_2923_0,
    i_13_288_3107_0, i_13_288_3142_0, i_13_288_3143_0, i_13_288_3242_0,
    i_13_288_3267_0, i_13_288_3269_0, i_13_288_3271_0, i_13_288_3371_0,
    i_13_288_3420_0, i_13_288_3421_0, i_13_288_3422_0, i_13_288_3424_0,
    i_13_288_3425_0, i_13_288_3545_0, i_13_288_3646_0, i_13_288_3730_0,
    i_13_288_3731_0, i_13_288_3767_0, i_13_288_3817_0, i_13_288_3818_0,
    i_13_288_3925_0, i_13_288_3971_0, i_13_288_3989_0, i_13_288_4015_0,
    i_13_288_4016_0, i_13_288_4018_0, i_13_288_4019_0, i_13_288_4044_0,
    i_13_288_4060_0, i_13_288_4061_0, i_13_288_4078_0, i_13_288_4214_0,
    i_13_288_4249_0, i_13_288_4250_0, i_13_288_4253_0, i_13_288_4261_0,
    i_13_288_4313_0, i_13_288_4340_0, i_13_288_4351_0, i_13_288_4430_0,
    i_13_288_4556_0, i_13_288_4558_0, i_13_288_4567_0, i_13_288_4591_0;
  output o_13_288_0_0;
  assign o_13_288_0_0 = ~((~i_13_288_1499_0 & ~i_13_288_4060_0) | (~i_13_288_1730_0 & ~i_13_288_1838_0 & ~i_13_288_3818_0));
endmodule



// Benchmark "kernel_13_289" written by ABC on Sun Jul 19 10:49:24 2020

module kernel_13_289 ( 
    i_13_289_120_0, i_13_289_139_0, i_13_289_140_0, i_13_289_142_0,
    i_13_289_175_0, i_13_289_177_0, i_13_289_227_0, i_13_289_228_0,
    i_13_289_281_0, i_13_289_310_0, i_13_289_338_0, i_13_289_371_0,
    i_13_289_418_0, i_13_289_532_0, i_13_289_538_0, i_13_289_617_0,
    i_13_289_654_0, i_13_289_700_0, i_13_289_769_0, i_13_289_817_0,
    i_13_289_821_0, i_13_289_892_0, i_13_289_897_0, i_13_289_918_0,
    i_13_289_982_0, i_13_289_985_0, i_13_289_1114_0, i_13_289_1219_0,
    i_13_289_1220_0, i_13_289_1228_0, i_13_289_1327_0, i_13_289_1424_0,
    i_13_289_1473_0, i_13_289_1525_0, i_13_289_1599_0, i_13_289_1627_0,
    i_13_289_1711_0, i_13_289_1714_0, i_13_289_1720_0, i_13_289_1723_0,
    i_13_289_1724_0, i_13_289_1831_0, i_13_289_1841_0, i_13_289_1844_0,
    i_13_289_1849_0, i_13_289_1882_0, i_13_289_1883_0, i_13_289_1885_0,
    i_13_289_1888_0, i_13_289_2104_0, i_13_289_2110_0, i_13_289_2206_0,
    i_13_289_2407_0, i_13_289_2410_0, i_13_289_2424_0, i_13_289_2463_0,
    i_13_289_2499_0, i_13_289_2663_0, i_13_289_2678_0, i_13_289_2695_0,
    i_13_289_2845_0, i_13_289_2846_0, i_13_289_2857_0, i_13_289_2875_0,
    i_13_289_2983_0, i_13_289_3005_0, i_13_289_3010_0, i_13_289_3109_0,
    i_13_289_3142_0, i_13_289_3143_0, i_13_289_3165_0, i_13_289_3444_0,
    i_13_289_3450_0, i_13_289_3451_0, i_13_289_3482_0, i_13_289_3503_0,
    i_13_289_3505_0, i_13_289_3506_0, i_13_289_3524_0, i_13_289_3571_0,
    i_13_289_3685_0, i_13_289_3686_0, i_13_289_3688_0, i_13_289_3736_0,
    i_13_289_3737_0, i_13_289_3740_0, i_13_289_3820_0, i_13_289_3836_0,
    i_13_289_3900_0, i_13_289_3928_0, i_13_289_4015_0, i_13_289_4066_0,
    i_13_289_4082_0, i_13_289_4204_0, i_13_289_4315_0, i_13_289_4388_0,
    i_13_289_4412_0, i_13_289_4459_0, i_13_289_4520_0, i_13_289_4567_0,
    o_13_289_0_0  );
  input  i_13_289_120_0, i_13_289_139_0, i_13_289_140_0, i_13_289_142_0,
    i_13_289_175_0, i_13_289_177_0, i_13_289_227_0, i_13_289_228_0,
    i_13_289_281_0, i_13_289_310_0, i_13_289_338_0, i_13_289_371_0,
    i_13_289_418_0, i_13_289_532_0, i_13_289_538_0, i_13_289_617_0,
    i_13_289_654_0, i_13_289_700_0, i_13_289_769_0, i_13_289_817_0,
    i_13_289_821_0, i_13_289_892_0, i_13_289_897_0, i_13_289_918_0,
    i_13_289_982_0, i_13_289_985_0, i_13_289_1114_0, i_13_289_1219_0,
    i_13_289_1220_0, i_13_289_1228_0, i_13_289_1327_0, i_13_289_1424_0,
    i_13_289_1473_0, i_13_289_1525_0, i_13_289_1599_0, i_13_289_1627_0,
    i_13_289_1711_0, i_13_289_1714_0, i_13_289_1720_0, i_13_289_1723_0,
    i_13_289_1724_0, i_13_289_1831_0, i_13_289_1841_0, i_13_289_1844_0,
    i_13_289_1849_0, i_13_289_1882_0, i_13_289_1883_0, i_13_289_1885_0,
    i_13_289_1888_0, i_13_289_2104_0, i_13_289_2110_0, i_13_289_2206_0,
    i_13_289_2407_0, i_13_289_2410_0, i_13_289_2424_0, i_13_289_2463_0,
    i_13_289_2499_0, i_13_289_2663_0, i_13_289_2678_0, i_13_289_2695_0,
    i_13_289_2845_0, i_13_289_2846_0, i_13_289_2857_0, i_13_289_2875_0,
    i_13_289_2983_0, i_13_289_3005_0, i_13_289_3010_0, i_13_289_3109_0,
    i_13_289_3142_0, i_13_289_3143_0, i_13_289_3165_0, i_13_289_3444_0,
    i_13_289_3450_0, i_13_289_3451_0, i_13_289_3482_0, i_13_289_3503_0,
    i_13_289_3505_0, i_13_289_3506_0, i_13_289_3524_0, i_13_289_3571_0,
    i_13_289_3685_0, i_13_289_3686_0, i_13_289_3688_0, i_13_289_3736_0,
    i_13_289_3737_0, i_13_289_3740_0, i_13_289_3820_0, i_13_289_3836_0,
    i_13_289_3900_0, i_13_289_3928_0, i_13_289_4015_0, i_13_289_4066_0,
    i_13_289_4082_0, i_13_289_4204_0, i_13_289_4315_0, i_13_289_4388_0,
    i_13_289_4412_0, i_13_289_4459_0, i_13_289_4520_0, i_13_289_4567_0;
  output o_13_289_0_0;
  assign o_13_289_0_0 = ~((i_13_289_1831_0 & ((~i_13_289_1220_0 & ~i_13_289_1711_0 & ~i_13_289_3688_0 & ~i_13_289_3737_0) | (~i_13_289_1219_0 & ~i_13_289_3736_0 & ~i_13_289_4412_0))) | (~i_13_289_2845_0 & ((~i_13_289_1841_0 & ~i_13_289_2424_0 & ~i_13_289_2857_0 & ~i_13_289_3450_0 & ~i_13_289_3524_0 & ~i_13_289_3571_0) | (~i_13_289_140_0 & ~i_13_289_310_0 & ~i_13_289_3444_0 & ~i_13_289_3685_0))) | (i_13_289_3571_0 & (i_13_289_3109_0 | ~i_13_289_3451_0)) | (~i_13_289_617_0 & ~i_13_289_2678_0 & i_13_289_2695_0) | (i_13_289_2983_0 & ~i_13_289_3506_0) | (i_13_289_1599_0 & ~i_13_289_1627_0 & i_13_289_2407_0 & ~i_13_289_3685_0) | (i_13_289_1327_0 & ~i_13_289_3737_0 & ~i_13_289_4082_0) | (~i_13_289_3505_0 & i_13_289_4315_0));
endmodule



// Benchmark "kernel_13_290" written by ABC on Sun Jul 19 10:49:25 2020

module kernel_13_290 ( 
    i_13_290_127_0, i_13_290_130_0, i_13_290_131_0, i_13_290_272_0,
    i_13_290_280_0, i_13_290_329_0, i_13_290_354_0, i_13_290_355_0,
    i_13_290_364_0, i_13_290_442_0, i_13_290_469_0, i_13_290_490_0,
    i_13_290_667_0, i_13_290_668_0, i_13_290_694_0, i_13_290_820_0,
    i_13_290_828_0, i_13_290_829_0, i_13_290_830_0, i_13_290_939_0,
    i_13_290_946_0, i_13_290_1022_0, i_13_290_1081_0, i_13_290_1100_0,
    i_13_290_1256_0, i_13_290_1271_0, i_13_290_1306_0, i_13_290_1307_0,
    i_13_290_1397_0, i_13_290_1435_0, i_13_290_1499_0, i_13_290_1504_0,
    i_13_290_1620_0, i_13_290_1639_0, i_13_290_1640_0, i_13_290_1657_0,
    i_13_290_1696_0, i_13_290_1697_0, i_13_290_1721_0, i_13_290_1777_0,
    i_13_290_1792_0, i_13_290_1793_0, i_13_290_1846_0, i_13_290_2029_0,
    i_13_290_2142_0, i_13_290_2143_0, i_13_290_2191_0, i_13_290_2296_0,
    i_13_290_2297_0, i_13_290_2317_0, i_13_290_2431_0, i_13_290_2432_0,
    i_13_290_2444_0, i_13_290_2468_0, i_13_290_2511_0, i_13_290_2512_0,
    i_13_290_2549_0, i_13_290_2552_0, i_13_290_2692_0, i_13_290_2719_0,
    i_13_290_2720_0, i_13_290_2880_0, i_13_290_2881_0, i_13_290_2882_0,
    i_13_290_2921_0, i_13_290_2935_0, i_13_290_3097_0, i_13_290_3136_0,
    i_13_290_3241_0, i_13_290_3242_0, i_13_290_3416_0, i_13_290_3421_0,
    i_13_290_3523_0, i_13_290_3595_0, i_13_290_3619_0, i_13_290_3620_0,
    i_13_290_3631_0, i_13_290_3632_0, i_13_290_3731_0, i_13_290_3754_0,
    i_13_290_3780_0, i_13_290_3802_0, i_13_290_3925_0, i_13_290_3935_0,
    i_13_290_3989_0, i_13_290_3991_0, i_13_290_3992_0, i_13_290_4198_0,
    i_13_290_4212_0, i_13_290_4214_0, i_13_290_4311_0, i_13_290_4313_0,
    i_13_290_4329_0, i_13_290_4330_0, i_13_290_4331_0, i_13_290_4339_0,
    i_13_290_4429_0, i_13_290_4430_0, i_13_290_4450_0, i_13_290_4510_0,
    o_13_290_0_0  );
  input  i_13_290_127_0, i_13_290_130_0, i_13_290_131_0, i_13_290_272_0,
    i_13_290_280_0, i_13_290_329_0, i_13_290_354_0, i_13_290_355_0,
    i_13_290_364_0, i_13_290_442_0, i_13_290_469_0, i_13_290_490_0,
    i_13_290_667_0, i_13_290_668_0, i_13_290_694_0, i_13_290_820_0,
    i_13_290_828_0, i_13_290_829_0, i_13_290_830_0, i_13_290_939_0,
    i_13_290_946_0, i_13_290_1022_0, i_13_290_1081_0, i_13_290_1100_0,
    i_13_290_1256_0, i_13_290_1271_0, i_13_290_1306_0, i_13_290_1307_0,
    i_13_290_1397_0, i_13_290_1435_0, i_13_290_1499_0, i_13_290_1504_0,
    i_13_290_1620_0, i_13_290_1639_0, i_13_290_1640_0, i_13_290_1657_0,
    i_13_290_1696_0, i_13_290_1697_0, i_13_290_1721_0, i_13_290_1777_0,
    i_13_290_1792_0, i_13_290_1793_0, i_13_290_1846_0, i_13_290_2029_0,
    i_13_290_2142_0, i_13_290_2143_0, i_13_290_2191_0, i_13_290_2296_0,
    i_13_290_2297_0, i_13_290_2317_0, i_13_290_2431_0, i_13_290_2432_0,
    i_13_290_2444_0, i_13_290_2468_0, i_13_290_2511_0, i_13_290_2512_0,
    i_13_290_2549_0, i_13_290_2552_0, i_13_290_2692_0, i_13_290_2719_0,
    i_13_290_2720_0, i_13_290_2880_0, i_13_290_2881_0, i_13_290_2882_0,
    i_13_290_2921_0, i_13_290_2935_0, i_13_290_3097_0, i_13_290_3136_0,
    i_13_290_3241_0, i_13_290_3242_0, i_13_290_3416_0, i_13_290_3421_0,
    i_13_290_3523_0, i_13_290_3595_0, i_13_290_3619_0, i_13_290_3620_0,
    i_13_290_3631_0, i_13_290_3632_0, i_13_290_3731_0, i_13_290_3754_0,
    i_13_290_3780_0, i_13_290_3802_0, i_13_290_3925_0, i_13_290_3935_0,
    i_13_290_3989_0, i_13_290_3991_0, i_13_290_3992_0, i_13_290_4198_0,
    i_13_290_4212_0, i_13_290_4214_0, i_13_290_4311_0, i_13_290_4313_0,
    i_13_290_4329_0, i_13_290_4330_0, i_13_290_4331_0, i_13_290_4339_0,
    i_13_290_4429_0, i_13_290_4430_0, i_13_290_4450_0, i_13_290_4510_0;
  output o_13_290_0_0;
  assign o_13_290_0_0 = ~((~i_13_290_694_0 & ~i_13_290_1639_0 & ~i_13_290_3241_0) | (~i_13_290_1081_0 & ~i_13_290_3242_0 & ~i_13_290_4429_0 & ~i_13_290_4510_0) | (~i_13_290_355_0 & ~i_13_290_830_0 & ~i_13_290_1504_0 & ~i_13_290_2432_0));
endmodule



// Benchmark "kernel_13_291" written by ABC on Sun Jul 19 10:49:26 2020

module kernel_13_291 ( 
    i_13_291_31_0, i_13_291_48_0, i_13_291_49_0, i_13_291_51_0,
    i_13_291_94_0, i_13_291_121_0, i_13_291_137_0, i_13_291_166_0,
    i_13_291_229_0, i_13_291_316_0, i_13_291_514_0, i_13_291_550_0,
    i_13_291_558_0, i_13_291_640_0, i_13_291_652_0, i_13_291_657_0,
    i_13_291_676_0, i_13_291_677_0, i_13_291_678_0, i_13_291_756_0,
    i_13_291_757_0, i_13_291_838_0, i_13_291_839_0, i_13_291_855_0,
    i_13_291_928_0, i_13_291_939_0, i_13_291_940_0, i_13_291_981_0,
    i_13_291_982_0, i_13_291_1063_0, i_13_291_1072_0, i_13_291_1080_0,
    i_13_291_1098_0, i_13_291_1323_0, i_13_291_1324_0, i_13_291_1327_0,
    i_13_291_1486_0, i_13_291_1570_0, i_13_291_1647_0, i_13_291_1747_0,
    i_13_291_1809_0, i_13_291_1831_0, i_13_291_1908_0, i_13_291_1911_0,
    i_13_291_2016_0, i_13_291_2017_0, i_13_291_2052_0, i_13_291_2055_0,
    i_13_291_2107_0, i_13_291_2116_0, i_13_291_2260_0, i_13_291_2380_0,
    i_13_291_2407_0, i_13_291_2433_0, i_13_291_2448_0, i_13_291_2449_0,
    i_13_291_2467_0, i_13_291_2505_0, i_13_291_2506_0, i_13_291_2592_0,
    i_13_291_2674_0, i_13_291_2702_0, i_13_291_2710_0, i_13_291_2749_0,
    i_13_291_2817_0, i_13_291_2908_0, i_13_291_2939_0, i_13_291_2979_0,
    i_13_291_2980_0, i_13_291_3025_0, i_13_291_3096_0, i_13_291_3109_0,
    i_13_291_3110_0, i_13_291_3142_0, i_13_291_3291_0, i_13_291_3519_0,
    i_13_291_3532_0, i_13_291_3541_0, i_13_291_3549_0, i_13_291_3550_0,
    i_13_291_3646_0, i_13_291_3737_0, i_13_291_3765_0, i_13_291_3766_0,
    i_13_291_3817_0, i_13_291_3818_0, i_13_291_3862_0, i_13_291_3889_0,
    i_13_291_3987_0, i_13_291_3988_0, i_13_291_4063_0, i_13_291_4087_0,
    i_13_291_4122_0, i_13_291_4158_0, i_13_291_4185_0, i_13_291_4279_0,
    i_13_291_4320_0, i_13_291_4393_0, i_13_291_4591_0, i_13_291_4600_0,
    o_13_291_0_0  );
  input  i_13_291_31_0, i_13_291_48_0, i_13_291_49_0, i_13_291_51_0,
    i_13_291_94_0, i_13_291_121_0, i_13_291_137_0, i_13_291_166_0,
    i_13_291_229_0, i_13_291_316_0, i_13_291_514_0, i_13_291_550_0,
    i_13_291_558_0, i_13_291_640_0, i_13_291_652_0, i_13_291_657_0,
    i_13_291_676_0, i_13_291_677_0, i_13_291_678_0, i_13_291_756_0,
    i_13_291_757_0, i_13_291_838_0, i_13_291_839_0, i_13_291_855_0,
    i_13_291_928_0, i_13_291_939_0, i_13_291_940_0, i_13_291_981_0,
    i_13_291_982_0, i_13_291_1063_0, i_13_291_1072_0, i_13_291_1080_0,
    i_13_291_1098_0, i_13_291_1323_0, i_13_291_1324_0, i_13_291_1327_0,
    i_13_291_1486_0, i_13_291_1570_0, i_13_291_1647_0, i_13_291_1747_0,
    i_13_291_1809_0, i_13_291_1831_0, i_13_291_1908_0, i_13_291_1911_0,
    i_13_291_2016_0, i_13_291_2017_0, i_13_291_2052_0, i_13_291_2055_0,
    i_13_291_2107_0, i_13_291_2116_0, i_13_291_2260_0, i_13_291_2380_0,
    i_13_291_2407_0, i_13_291_2433_0, i_13_291_2448_0, i_13_291_2449_0,
    i_13_291_2467_0, i_13_291_2505_0, i_13_291_2506_0, i_13_291_2592_0,
    i_13_291_2674_0, i_13_291_2702_0, i_13_291_2710_0, i_13_291_2749_0,
    i_13_291_2817_0, i_13_291_2908_0, i_13_291_2939_0, i_13_291_2979_0,
    i_13_291_2980_0, i_13_291_3025_0, i_13_291_3096_0, i_13_291_3109_0,
    i_13_291_3110_0, i_13_291_3142_0, i_13_291_3291_0, i_13_291_3519_0,
    i_13_291_3532_0, i_13_291_3541_0, i_13_291_3549_0, i_13_291_3550_0,
    i_13_291_3646_0, i_13_291_3737_0, i_13_291_3765_0, i_13_291_3766_0,
    i_13_291_3817_0, i_13_291_3818_0, i_13_291_3862_0, i_13_291_3889_0,
    i_13_291_3987_0, i_13_291_3988_0, i_13_291_4063_0, i_13_291_4087_0,
    i_13_291_4122_0, i_13_291_4158_0, i_13_291_4185_0, i_13_291_4279_0,
    i_13_291_4320_0, i_13_291_4393_0, i_13_291_4591_0, i_13_291_4600_0;
  output o_13_291_0_0;
  assign o_13_291_0_0 = ~((i_13_291_3818_0 & ((~i_13_291_3142_0 & i_13_291_4393_0) | (~i_13_291_1327_0 & ~i_13_291_4393_0))) | i_13_291_3737_0 | (~i_13_291_316_0 & ~i_13_291_3519_0) | (~i_13_291_839_0 & ~i_13_291_2448_0 & ~i_13_291_3765_0) | (~i_13_291_3109_0 & ~i_13_291_3988_0 & ~i_13_291_4087_0) | (~i_13_291_756_0 & ~i_13_291_3817_0 & ~i_13_291_4158_0));
endmodule



// Benchmark "kernel_13_292" written by ABC on Sun Jul 19 10:49:26 2020

module kernel_13_292 ( 
    i_13_292_49_0, i_13_292_70_0, i_13_292_71_0, i_13_292_78_0,
    i_13_292_79_0, i_13_292_80_0, i_13_292_105_0, i_13_292_232_0,
    i_13_292_312_0, i_13_292_313_0, i_13_292_314_0, i_13_292_319_0,
    i_13_292_320_0, i_13_292_358_0, i_13_292_448_0, i_13_292_457_0,
    i_13_292_525_0, i_13_292_553_0, i_13_292_624_0, i_13_292_644_0,
    i_13_292_646_0, i_13_292_673_0, i_13_292_682_0, i_13_292_688_0,
    i_13_292_689_0, i_13_292_692_0, i_13_292_844_0, i_13_292_935_0,
    i_13_292_969_0, i_13_292_1050_0, i_13_292_1104_0, i_13_292_1105_0,
    i_13_292_1110_0, i_13_292_1123_0, i_13_292_1274_0, i_13_292_1311_0,
    i_13_292_1312_0, i_13_292_1330_0, i_13_292_1402_0, i_13_292_1403_0,
    i_13_292_1429_0, i_13_292_1508_0, i_13_292_1510_0, i_13_292_1541_0,
    i_13_292_1645_0, i_13_292_1646_0, i_13_292_1798_0, i_13_292_1799_0,
    i_13_292_1843_0, i_13_292_1853_0, i_13_292_1887_0, i_13_292_1912_0,
    i_13_292_1945_0, i_13_292_1946_0, i_13_292_1948_0, i_13_292_2027_0,
    i_13_292_2104_0, i_13_292_2203_0, i_13_292_2229_0, i_13_292_2245_0,
    i_13_292_2291_0, i_13_292_2415_0, i_13_292_2680_0, i_13_292_2697_0,
    i_13_292_2698_0, i_13_292_2699_0, i_13_292_2852_0, i_13_292_2853_0,
    i_13_292_2858_0, i_13_292_2923_0, i_13_292_3031_0, i_13_292_3054_0,
    i_13_292_3067_0, i_13_292_3130_0, i_13_292_3138_0, i_13_292_3245_0,
    i_13_292_3370_0, i_13_292_3373_0, i_13_292_3418_0, i_13_292_3561_0,
    i_13_292_3595_0, i_13_292_3622_0, i_13_292_3623_0, i_13_292_3652_0,
    i_13_292_3787_0, i_13_292_3895_0, i_13_292_3931_0, i_13_292_3940_0,
    i_13_292_3994_0, i_13_292_3995_0, i_13_292_4068_0, i_13_292_4084_0,
    i_13_292_4111_0, i_13_292_4156_0, i_13_292_4435_0, i_13_292_4454_0,
    i_13_292_4595_0, i_13_292_4596_0, i_13_292_4597_0, i_13_292_4598_0,
    o_13_292_0_0  );
  input  i_13_292_49_0, i_13_292_70_0, i_13_292_71_0, i_13_292_78_0,
    i_13_292_79_0, i_13_292_80_0, i_13_292_105_0, i_13_292_232_0,
    i_13_292_312_0, i_13_292_313_0, i_13_292_314_0, i_13_292_319_0,
    i_13_292_320_0, i_13_292_358_0, i_13_292_448_0, i_13_292_457_0,
    i_13_292_525_0, i_13_292_553_0, i_13_292_624_0, i_13_292_644_0,
    i_13_292_646_0, i_13_292_673_0, i_13_292_682_0, i_13_292_688_0,
    i_13_292_689_0, i_13_292_692_0, i_13_292_844_0, i_13_292_935_0,
    i_13_292_969_0, i_13_292_1050_0, i_13_292_1104_0, i_13_292_1105_0,
    i_13_292_1110_0, i_13_292_1123_0, i_13_292_1274_0, i_13_292_1311_0,
    i_13_292_1312_0, i_13_292_1330_0, i_13_292_1402_0, i_13_292_1403_0,
    i_13_292_1429_0, i_13_292_1508_0, i_13_292_1510_0, i_13_292_1541_0,
    i_13_292_1645_0, i_13_292_1646_0, i_13_292_1798_0, i_13_292_1799_0,
    i_13_292_1843_0, i_13_292_1853_0, i_13_292_1887_0, i_13_292_1912_0,
    i_13_292_1945_0, i_13_292_1946_0, i_13_292_1948_0, i_13_292_2027_0,
    i_13_292_2104_0, i_13_292_2203_0, i_13_292_2229_0, i_13_292_2245_0,
    i_13_292_2291_0, i_13_292_2415_0, i_13_292_2680_0, i_13_292_2697_0,
    i_13_292_2698_0, i_13_292_2699_0, i_13_292_2852_0, i_13_292_2853_0,
    i_13_292_2858_0, i_13_292_2923_0, i_13_292_3031_0, i_13_292_3054_0,
    i_13_292_3067_0, i_13_292_3130_0, i_13_292_3138_0, i_13_292_3245_0,
    i_13_292_3370_0, i_13_292_3373_0, i_13_292_3418_0, i_13_292_3561_0,
    i_13_292_3595_0, i_13_292_3622_0, i_13_292_3623_0, i_13_292_3652_0,
    i_13_292_3787_0, i_13_292_3895_0, i_13_292_3931_0, i_13_292_3940_0,
    i_13_292_3994_0, i_13_292_3995_0, i_13_292_4068_0, i_13_292_4084_0,
    i_13_292_4111_0, i_13_292_4156_0, i_13_292_4435_0, i_13_292_4454_0,
    i_13_292_4595_0, i_13_292_4596_0, i_13_292_4597_0, i_13_292_4598_0;
  output o_13_292_0_0;
  assign o_13_292_0_0 = 0;
endmodule



// Benchmark "kernel_13_293" written by ABC on Sun Jul 19 10:49:27 2020

module kernel_13_293 ( 
    i_13_293_49_0, i_13_293_74_0, i_13_293_77_0, i_13_293_113_0,
    i_13_293_166_0, i_13_293_172_0, i_13_293_175_0, i_13_293_176_0,
    i_13_293_200_0, i_13_293_326_0, i_13_293_337_0, i_13_293_523_0,
    i_13_293_544_0, i_13_293_658_0, i_13_293_661_0, i_13_293_662_0,
    i_13_293_694_0, i_13_293_824_0, i_13_293_839_0, i_13_293_841_0,
    i_13_293_848_0, i_13_293_853_0, i_13_293_859_0, i_13_293_1018_0,
    i_13_293_1019_0, i_13_293_1072_0, i_13_293_1073_0, i_13_293_1148_0,
    i_13_293_1225_0, i_13_293_1226_0, i_13_293_1229_0, i_13_293_1231_0,
    i_13_293_1253_0, i_13_293_1310_0, i_13_293_1315_0, i_13_293_1316_0,
    i_13_293_1324_0, i_13_293_1378_0, i_13_293_1424_0, i_13_293_1427_0,
    i_13_293_1441_0, i_13_293_1486_0, i_13_293_1487_0, i_13_293_1549_0,
    i_13_293_1550_0, i_13_293_1630_0, i_13_293_1778_0, i_13_293_1849_0,
    i_13_293_1883_0, i_13_293_1885_0, i_13_293_1886_0, i_13_293_1909_0,
    i_13_293_2021_0, i_13_293_2137_0, i_13_293_2173_0, i_13_293_2371_0,
    i_13_293_2452_0, i_13_293_2453_0, i_13_293_2462_0, i_13_293_2539_0,
    i_13_293_2540_0, i_13_293_2561_0, i_13_293_2611_0, i_13_293_2749_0,
    i_13_293_2917_0, i_13_293_2984_0, i_13_293_3269_0, i_13_293_3367_0,
    i_13_293_3370_0, i_13_293_3395_0, i_13_293_3484_0, i_13_293_3485_0,
    i_13_293_3488_0, i_13_293_3502_0, i_13_293_3503_0, i_13_293_3530_0,
    i_13_293_3538_0, i_13_293_3539_0, i_13_293_3541_0, i_13_293_3542_0,
    i_13_293_3548_0, i_13_293_3574_0, i_13_293_3575_0, i_13_293_3703_0,
    i_13_293_3740_0, i_13_293_3812_0, i_13_293_3854_0, i_13_293_3866_0,
    i_13_293_3892_0, i_13_293_3916_0, i_13_293_4063_0, i_13_293_4064_0,
    i_13_293_4249_0, i_13_293_4250_0, i_13_293_4252_0, i_13_293_4253_0,
    i_13_293_4366_0, i_13_293_4369_0, i_13_293_4376_0, i_13_293_4448_0,
    o_13_293_0_0  );
  input  i_13_293_49_0, i_13_293_74_0, i_13_293_77_0, i_13_293_113_0,
    i_13_293_166_0, i_13_293_172_0, i_13_293_175_0, i_13_293_176_0,
    i_13_293_200_0, i_13_293_326_0, i_13_293_337_0, i_13_293_523_0,
    i_13_293_544_0, i_13_293_658_0, i_13_293_661_0, i_13_293_662_0,
    i_13_293_694_0, i_13_293_824_0, i_13_293_839_0, i_13_293_841_0,
    i_13_293_848_0, i_13_293_853_0, i_13_293_859_0, i_13_293_1018_0,
    i_13_293_1019_0, i_13_293_1072_0, i_13_293_1073_0, i_13_293_1148_0,
    i_13_293_1225_0, i_13_293_1226_0, i_13_293_1229_0, i_13_293_1231_0,
    i_13_293_1253_0, i_13_293_1310_0, i_13_293_1315_0, i_13_293_1316_0,
    i_13_293_1324_0, i_13_293_1378_0, i_13_293_1424_0, i_13_293_1427_0,
    i_13_293_1441_0, i_13_293_1486_0, i_13_293_1487_0, i_13_293_1549_0,
    i_13_293_1550_0, i_13_293_1630_0, i_13_293_1778_0, i_13_293_1849_0,
    i_13_293_1883_0, i_13_293_1885_0, i_13_293_1886_0, i_13_293_1909_0,
    i_13_293_2021_0, i_13_293_2137_0, i_13_293_2173_0, i_13_293_2371_0,
    i_13_293_2452_0, i_13_293_2453_0, i_13_293_2462_0, i_13_293_2539_0,
    i_13_293_2540_0, i_13_293_2561_0, i_13_293_2611_0, i_13_293_2749_0,
    i_13_293_2917_0, i_13_293_2984_0, i_13_293_3269_0, i_13_293_3367_0,
    i_13_293_3370_0, i_13_293_3395_0, i_13_293_3484_0, i_13_293_3485_0,
    i_13_293_3488_0, i_13_293_3502_0, i_13_293_3503_0, i_13_293_3530_0,
    i_13_293_3538_0, i_13_293_3539_0, i_13_293_3541_0, i_13_293_3542_0,
    i_13_293_3548_0, i_13_293_3574_0, i_13_293_3575_0, i_13_293_3703_0,
    i_13_293_3740_0, i_13_293_3812_0, i_13_293_3854_0, i_13_293_3866_0,
    i_13_293_3892_0, i_13_293_3916_0, i_13_293_4063_0, i_13_293_4064_0,
    i_13_293_4249_0, i_13_293_4250_0, i_13_293_4252_0, i_13_293_4253_0,
    i_13_293_4366_0, i_13_293_4369_0, i_13_293_4376_0, i_13_293_4448_0;
  output o_13_293_0_0;
  assign o_13_293_0_0 = ~(~i_13_293_4252_0 | (~i_13_293_1427_0 & ~i_13_293_4366_0) | (~i_13_293_3740_0 & ~i_13_293_4250_0) | (~i_13_293_824_0 & ~i_13_293_3530_0) | (~i_13_293_74_0 & ~i_13_293_3548_0 & ~i_13_293_3575_0) | (i_13_293_1324_0 & ~i_13_293_3854_0 & ~i_13_293_3892_0 & ~i_13_293_4369_0));
endmodule



// Benchmark "kernel_13_294" written by ABC on Sun Jul 19 10:49:28 2020

module kernel_13_294 ( 
    i_13_294_28_0, i_13_294_29_0, i_13_294_52_0, i_13_294_65_0,
    i_13_294_103_0, i_13_294_124_0, i_13_294_140_0, i_13_294_175_0,
    i_13_294_211_0, i_13_294_257_0, i_13_294_266_0, i_13_294_308_0,
    i_13_294_316_0, i_13_294_340_0, i_13_294_358_0, i_13_294_359_0,
    i_13_294_371_0, i_13_294_418_0, i_13_294_419_0, i_13_294_584_0,
    i_13_294_587_0, i_13_294_604_0, i_13_294_640_0, i_13_294_641_0,
    i_13_294_668_0, i_13_294_679_0, i_13_294_757_0, i_13_294_758_0,
    i_13_294_856_0, i_13_294_928_0, i_13_294_1081_0, i_13_294_1082_0,
    i_13_294_1117_0, i_13_294_1300_0, i_13_294_1342_0, i_13_294_1343_0,
    i_13_294_1345_0, i_13_294_1501_0, i_13_294_1502_0, i_13_294_1567_0,
    i_13_294_1637_0, i_13_294_1793_0, i_13_294_1804_0, i_13_294_1813_0,
    i_13_294_1840_0, i_13_294_1841_0, i_13_294_1928_0, i_13_294_1991_0,
    i_13_294_2002_0, i_13_294_2032_0, i_13_294_2033_0, i_13_294_2054_0,
    i_13_294_2119_0, i_13_294_2137_0, i_13_294_2260_0, i_13_294_2432_0,
    i_13_294_2549_0, i_13_294_2554_0, i_13_294_2674_0, i_13_294_2675_0,
    i_13_294_2710_0, i_13_294_2719_0, i_13_294_2846_0, i_13_294_2848_0,
    i_13_294_2924_0, i_13_294_2938_0, i_13_294_2960_0, i_13_294_3061_0,
    i_13_294_3073_0, i_13_294_3088_0, i_13_294_3217_0, i_13_294_3289_0,
    i_13_294_3343_0, i_13_294_3386_0, i_13_294_3415_0, i_13_294_3416_0,
    i_13_294_3440_0, i_13_294_3485_0, i_13_294_3501_0, i_13_294_3502_0,
    i_13_294_3503_0, i_13_294_3634_0, i_13_294_3737_0, i_13_294_3788_0,
    i_13_294_3800_0, i_13_294_3806_0, i_13_294_3851_0, i_13_294_3893_0,
    i_13_294_4018_0, i_13_294_4034_0, i_13_294_4078_0, i_13_294_4234_0,
    i_13_294_4267_0, i_13_294_4268_0, i_13_294_4270_0, i_13_294_4274_0,
    i_13_294_4411_0, i_13_294_4454_0, i_13_294_4591_0, i_13_294_4592_0,
    o_13_294_0_0  );
  input  i_13_294_28_0, i_13_294_29_0, i_13_294_52_0, i_13_294_65_0,
    i_13_294_103_0, i_13_294_124_0, i_13_294_140_0, i_13_294_175_0,
    i_13_294_211_0, i_13_294_257_0, i_13_294_266_0, i_13_294_308_0,
    i_13_294_316_0, i_13_294_340_0, i_13_294_358_0, i_13_294_359_0,
    i_13_294_371_0, i_13_294_418_0, i_13_294_419_0, i_13_294_584_0,
    i_13_294_587_0, i_13_294_604_0, i_13_294_640_0, i_13_294_641_0,
    i_13_294_668_0, i_13_294_679_0, i_13_294_757_0, i_13_294_758_0,
    i_13_294_856_0, i_13_294_928_0, i_13_294_1081_0, i_13_294_1082_0,
    i_13_294_1117_0, i_13_294_1300_0, i_13_294_1342_0, i_13_294_1343_0,
    i_13_294_1345_0, i_13_294_1501_0, i_13_294_1502_0, i_13_294_1567_0,
    i_13_294_1637_0, i_13_294_1793_0, i_13_294_1804_0, i_13_294_1813_0,
    i_13_294_1840_0, i_13_294_1841_0, i_13_294_1928_0, i_13_294_1991_0,
    i_13_294_2002_0, i_13_294_2032_0, i_13_294_2033_0, i_13_294_2054_0,
    i_13_294_2119_0, i_13_294_2137_0, i_13_294_2260_0, i_13_294_2432_0,
    i_13_294_2549_0, i_13_294_2554_0, i_13_294_2674_0, i_13_294_2675_0,
    i_13_294_2710_0, i_13_294_2719_0, i_13_294_2846_0, i_13_294_2848_0,
    i_13_294_2924_0, i_13_294_2938_0, i_13_294_2960_0, i_13_294_3061_0,
    i_13_294_3073_0, i_13_294_3088_0, i_13_294_3217_0, i_13_294_3289_0,
    i_13_294_3343_0, i_13_294_3386_0, i_13_294_3415_0, i_13_294_3416_0,
    i_13_294_3440_0, i_13_294_3485_0, i_13_294_3501_0, i_13_294_3502_0,
    i_13_294_3503_0, i_13_294_3634_0, i_13_294_3737_0, i_13_294_3788_0,
    i_13_294_3800_0, i_13_294_3806_0, i_13_294_3851_0, i_13_294_3893_0,
    i_13_294_4018_0, i_13_294_4034_0, i_13_294_4078_0, i_13_294_4234_0,
    i_13_294_4267_0, i_13_294_4268_0, i_13_294_4270_0, i_13_294_4274_0,
    i_13_294_4411_0, i_13_294_4454_0, i_13_294_4591_0, i_13_294_4592_0;
  output o_13_294_0_0;
  assign o_13_294_0_0 = ~(~i_13_294_1082_0 | (~i_13_294_3737_0 & i_13_294_4234_0) | (~i_13_294_29_0 & ~i_13_294_316_0));
endmodule



// Benchmark "kernel_13_295" written by ABC on Sun Jul 19 10:49:29 2020

module kernel_13_295 ( 
    i_13_295_39_0, i_13_295_94_0, i_13_295_95_0, i_13_295_97_0,
    i_13_295_102_0, i_13_295_176_0, i_13_295_178_0, i_13_295_179_0,
    i_13_295_241_0, i_13_295_310_0, i_13_295_311_0, i_13_295_313_0,
    i_13_295_314_0, i_13_295_318_0, i_13_295_319_0, i_13_295_320_0,
    i_13_295_337_0, i_13_295_418_0, i_13_295_510_0, i_13_295_527_0,
    i_13_295_574_0, i_13_295_575_0, i_13_295_580_0, i_13_295_643_0,
    i_13_295_646_0, i_13_295_647_0, i_13_295_674_0, i_13_295_689_0,
    i_13_295_872_0, i_13_295_931_0, i_13_295_985_0, i_13_295_988_0,
    i_13_295_989_0, i_13_295_1123_0, i_13_295_1124_0, i_13_295_1186_0,
    i_13_295_1444_0, i_13_295_1516_0, i_13_295_1526_0, i_13_295_1598_0,
    i_13_295_1641_0, i_13_295_1642_0, i_13_295_1813_0, i_13_295_1850_0,
    i_13_295_1934_0, i_13_295_2137_0, i_13_295_2176_0, i_13_295_2177_0,
    i_13_295_2264_0, i_13_295_2314_0, i_13_295_2408_0, i_13_295_2567_0,
    i_13_295_2614_0, i_13_295_2678_0, i_13_295_2680_0, i_13_295_2681_0,
    i_13_295_2698_0, i_13_295_2699_0, i_13_295_2788_0, i_13_295_2887_0,
    i_13_295_2923_0, i_13_295_2983_0, i_13_295_3010_0, i_13_295_3113_0,
    i_13_295_3127_0, i_13_295_3128_0, i_13_295_3212_0, i_13_295_3217_0,
    i_13_295_3274_0, i_13_295_3370_0, i_13_295_3379_0, i_13_295_3408_0,
    i_13_295_3409_0, i_13_295_3410_0, i_13_295_3415_0, i_13_295_3426_0,
    i_13_295_3469_0, i_13_295_3554_0, i_13_295_3688_0, i_13_295_3821_0,
    i_13_295_3901_0, i_13_295_3931_0, i_13_295_3932_0, i_13_295_4034_0,
    i_13_295_4036_0, i_13_295_4037_0, i_13_295_4084_0, i_13_295_4208_0,
    i_13_295_4261_0, i_13_295_4327_0, i_13_295_4342_0, i_13_295_4354_0,
    i_13_295_4522_0, i_13_295_4523_0, i_13_295_4568_0, i_13_295_4569_0,
    i_13_295_4570_0, i_13_295_4571_0, i_13_295_4595_0, i_13_295_4598_0,
    o_13_295_0_0  );
  input  i_13_295_39_0, i_13_295_94_0, i_13_295_95_0, i_13_295_97_0,
    i_13_295_102_0, i_13_295_176_0, i_13_295_178_0, i_13_295_179_0,
    i_13_295_241_0, i_13_295_310_0, i_13_295_311_0, i_13_295_313_0,
    i_13_295_314_0, i_13_295_318_0, i_13_295_319_0, i_13_295_320_0,
    i_13_295_337_0, i_13_295_418_0, i_13_295_510_0, i_13_295_527_0,
    i_13_295_574_0, i_13_295_575_0, i_13_295_580_0, i_13_295_643_0,
    i_13_295_646_0, i_13_295_647_0, i_13_295_674_0, i_13_295_689_0,
    i_13_295_872_0, i_13_295_931_0, i_13_295_985_0, i_13_295_988_0,
    i_13_295_989_0, i_13_295_1123_0, i_13_295_1124_0, i_13_295_1186_0,
    i_13_295_1444_0, i_13_295_1516_0, i_13_295_1526_0, i_13_295_1598_0,
    i_13_295_1641_0, i_13_295_1642_0, i_13_295_1813_0, i_13_295_1850_0,
    i_13_295_1934_0, i_13_295_2137_0, i_13_295_2176_0, i_13_295_2177_0,
    i_13_295_2264_0, i_13_295_2314_0, i_13_295_2408_0, i_13_295_2567_0,
    i_13_295_2614_0, i_13_295_2678_0, i_13_295_2680_0, i_13_295_2681_0,
    i_13_295_2698_0, i_13_295_2699_0, i_13_295_2788_0, i_13_295_2887_0,
    i_13_295_2923_0, i_13_295_2983_0, i_13_295_3010_0, i_13_295_3113_0,
    i_13_295_3127_0, i_13_295_3128_0, i_13_295_3212_0, i_13_295_3217_0,
    i_13_295_3274_0, i_13_295_3370_0, i_13_295_3379_0, i_13_295_3408_0,
    i_13_295_3409_0, i_13_295_3410_0, i_13_295_3415_0, i_13_295_3426_0,
    i_13_295_3469_0, i_13_295_3554_0, i_13_295_3688_0, i_13_295_3821_0,
    i_13_295_3901_0, i_13_295_3931_0, i_13_295_3932_0, i_13_295_4034_0,
    i_13_295_4036_0, i_13_295_4037_0, i_13_295_4084_0, i_13_295_4208_0,
    i_13_295_4261_0, i_13_295_4327_0, i_13_295_4342_0, i_13_295_4354_0,
    i_13_295_4522_0, i_13_295_4523_0, i_13_295_4568_0, i_13_295_4569_0,
    i_13_295_4570_0, i_13_295_4571_0, i_13_295_4595_0, i_13_295_4598_0;
  output o_13_295_0_0;
  assign o_13_295_0_0 = ~(i_13_295_3426_0 | (~i_13_295_3931_0 & ~i_13_295_4571_0) | (~i_13_295_1934_0 & ~i_13_295_4354_0) | (~i_13_295_527_0 & ~i_13_295_1123_0 & ~i_13_295_3212_0));
endmodule



// Benchmark "kernel_13_296" written by ABC on Sun Jul 19 10:49:29 2020

module kernel_13_296 ( 
    i_13_296_106_0, i_13_296_116_0, i_13_296_139_0, i_13_296_213_0,
    i_13_296_229_0, i_13_296_241_0, i_13_296_319_0, i_13_296_326_0,
    i_13_296_359_0, i_13_296_492_0, i_13_296_744_0, i_13_296_745_0,
    i_13_296_826_0, i_13_296_948_0, i_13_296_1066_0, i_13_296_1071_0,
    i_13_296_1087_0, i_13_296_1095_0, i_13_296_1096_0, i_13_296_1097_0,
    i_13_296_1131_0, i_13_296_1239_0, i_13_296_1267_0, i_13_296_1274_0,
    i_13_296_1302_0, i_13_296_1303_0, i_13_296_1347_0, i_13_296_1348_0,
    i_13_296_1349_0, i_13_296_1402_0, i_13_296_1435_0, i_13_296_1438_0,
    i_13_296_1446_0, i_13_296_1464_0, i_13_296_1529_0, i_13_296_1721_0,
    i_13_296_1722_0, i_13_296_1723_0, i_13_296_1755_0, i_13_296_1803_0,
    i_13_296_1815_0, i_13_296_1816_0, i_13_296_1817_0, i_13_296_1916_0,
    i_13_296_2023_0, i_13_296_2111_0, i_13_296_2123_0, i_13_296_2199_0,
    i_13_296_2238_0, i_13_296_2239_0, i_13_296_2273_0, i_13_296_2347_0,
    i_13_296_2348_0, i_13_296_2447_0, i_13_296_2500_0, i_13_296_2550_0,
    i_13_296_2715_0, i_13_296_2716_0, i_13_296_2717_0, i_13_296_2760_0,
    i_13_296_2789_0, i_13_296_2814_0, i_13_296_2822_0, i_13_296_2825_0,
    i_13_296_2853_0, i_13_296_2875_0, i_13_296_3023_0, i_13_296_3028_0,
    i_13_296_3036_0, i_13_296_3112_0, i_13_296_3328_0, i_13_296_3391_0,
    i_13_296_3422_0, i_13_296_3443_0, i_13_296_3446_0, i_13_296_3479_0,
    i_13_296_3482_0, i_13_296_3532_0, i_13_296_3594_0, i_13_296_3595_0,
    i_13_296_3622_0, i_13_296_3742_0, i_13_296_3817_0, i_13_296_3820_0,
    i_13_296_3830_0, i_13_296_3893_0, i_13_296_3921_0, i_13_296_3984_0,
    i_13_296_3985_0, i_13_296_4093_0, i_13_296_4120_0, i_13_296_4237_0,
    i_13_296_4252_0, i_13_296_4261_0, i_13_296_4272_0, i_13_296_4327_0,
    i_13_296_4328_0, i_13_296_4396_0, i_13_296_4399_0, i_13_296_4417_0,
    o_13_296_0_0  );
  input  i_13_296_106_0, i_13_296_116_0, i_13_296_139_0, i_13_296_213_0,
    i_13_296_229_0, i_13_296_241_0, i_13_296_319_0, i_13_296_326_0,
    i_13_296_359_0, i_13_296_492_0, i_13_296_744_0, i_13_296_745_0,
    i_13_296_826_0, i_13_296_948_0, i_13_296_1066_0, i_13_296_1071_0,
    i_13_296_1087_0, i_13_296_1095_0, i_13_296_1096_0, i_13_296_1097_0,
    i_13_296_1131_0, i_13_296_1239_0, i_13_296_1267_0, i_13_296_1274_0,
    i_13_296_1302_0, i_13_296_1303_0, i_13_296_1347_0, i_13_296_1348_0,
    i_13_296_1349_0, i_13_296_1402_0, i_13_296_1435_0, i_13_296_1438_0,
    i_13_296_1446_0, i_13_296_1464_0, i_13_296_1529_0, i_13_296_1721_0,
    i_13_296_1722_0, i_13_296_1723_0, i_13_296_1755_0, i_13_296_1803_0,
    i_13_296_1815_0, i_13_296_1816_0, i_13_296_1817_0, i_13_296_1916_0,
    i_13_296_2023_0, i_13_296_2111_0, i_13_296_2123_0, i_13_296_2199_0,
    i_13_296_2238_0, i_13_296_2239_0, i_13_296_2273_0, i_13_296_2347_0,
    i_13_296_2348_0, i_13_296_2447_0, i_13_296_2500_0, i_13_296_2550_0,
    i_13_296_2715_0, i_13_296_2716_0, i_13_296_2717_0, i_13_296_2760_0,
    i_13_296_2789_0, i_13_296_2814_0, i_13_296_2822_0, i_13_296_2825_0,
    i_13_296_2853_0, i_13_296_2875_0, i_13_296_3023_0, i_13_296_3028_0,
    i_13_296_3036_0, i_13_296_3112_0, i_13_296_3328_0, i_13_296_3391_0,
    i_13_296_3422_0, i_13_296_3443_0, i_13_296_3446_0, i_13_296_3479_0,
    i_13_296_3482_0, i_13_296_3532_0, i_13_296_3594_0, i_13_296_3595_0,
    i_13_296_3622_0, i_13_296_3742_0, i_13_296_3817_0, i_13_296_3820_0,
    i_13_296_3830_0, i_13_296_3893_0, i_13_296_3921_0, i_13_296_3984_0,
    i_13_296_3985_0, i_13_296_4093_0, i_13_296_4120_0, i_13_296_4237_0,
    i_13_296_4252_0, i_13_296_4261_0, i_13_296_4272_0, i_13_296_4327_0,
    i_13_296_4328_0, i_13_296_4396_0, i_13_296_4399_0, i_13_296_4417_0;
  output o_13_296_0_0;
  assign o_13_296_0_0 = ~((~i_13_296_2239_0 & ~i_13_296_3532_0 & ~i_13_296_4327_0) | (~i_13_296_1347_0 & ~i_13_296_2789_0 & ~i_13_296_3984_0 & ~i_13_296_4237_0));
endmodule



// Benchmark "kernel_13_297" written by ABC on Sun Jul 19 10:49:31 2020

module kernel_13_297 ( 
    i_13_297_69_0, i_13_297_124_0, i_13_297_154_0, i_13_297_166_0,
    i_13_297_178_0, i_13_297_195_0, i_13_297_210_0, i_13_297_211_0,
    i_13_297_228_0, i_13_297_231_0, i_13_297_232_0, i_13_297_247_0,
    i_13_297_376_0, i_13_297_528_0, i_13_297_534_0, i_13_297_640_0,
    i_13_297_642_0, i_13_297_646_0, i_13_297_714_0, i_13_297_717_0,
    i_13_297_771_0, i_13_297_826_0, i_13_297_861_0, i_13_297_862_0,
    i_13_297_895_0, i_13_297_951_0, i_13_297_952_0, i_13_297_1066_0,
    i_13_297_1075_0, i_13_297_1221_0, i_13_297_1222_0, i_13_297_1275_0,
    i_13_297_1293_0, i_13_297_1390_0, i_13_297_1410_0, i_13_297_1432_0,
    i_13_297_1491_0, i_13_297_1492_0, i_13_297_1627_0, i_13_297_1635_0,
    i_13_297_1641_0, i_13_297_1713_0, i_13_297_1726_0, i_13_297_1795_0,
    i_13_297_1842_0, i_13_297_1843_0, i_13_297_1884_0, i_13_297_1885_0,
    i_13_297_1929_0, i_13_297_1989_0, i_13_297_1993_0, i_13_297_2014_0,
    i_13_297_2028_0, i_13_297_2110_0, i_13_297_2175_0, i_13_297_2262_0,
    i_13_297_2410_0, i_13_297_2425_0, i_13_297_2463_0, i_13_297_2506_0,
    i_13_297_2535_0, i_13_297_2536_0, i_13_297_2616_0, i_13_297_2760_0,
    i_13_297_2847_0, i_13_297_2850_0, i_13_297_2851_0, i_13_297_3097_0,
    i_13_297_3345_0, i_13_297_3384_0, i_13_297_3387_0, i_13_297_3418_0,
    i_13_297_3426_0, i_13_297_3504_0, i_13_297_3505_0, i_13_297_3594_0,
    i_13_297_3669_0, i_13_297_3706_0, i_13_297_3766_0, i_13_297_3838_0,
    i_13_297_3876_0, i_13_297_3895_0, i_13_297_3931_0, i_13_297_4003_0,
    i_13_297_4011_0, i_13_297_4048_0, i_13_297_4080_0, i_13_297_4081_0,
    i_13_297_4086_0, i_13_297_4087_0, i_13_297_4114_0, i_13_297_4189_0,
    i_13_297_4210_0, i_13_297_4218_0, i_13_297_4273_0, i_13_297_4296_0,
    i_13_297_4297_0, i_13_297_4315_0, i_13_297_4543_0, i_13_297_4557_0,
    o_13_297_0_0  );
  input  i_13_297_69_0, i_13_297_124_0, i_13_297_154_0, i_13_297_166_0,
    i_13_297_178_0, i_13_297_195_0, i_13_297_210_0, i_13_297_211_0,
    i_13_297_228_0, i_13_297_231_0, i_13_297_232_0, i_13_297_247_0,
    i_13_297_376_0, i_13_297_528_0, i_13_297_534_0, i_13_297_640_0,
    i_13_297_642_0, i_13_297_646_0, i_13_297_714_0, i_13_297_717_0,
    i_13_297_771_0, i_13_297_826_0, i_13_297_861_0, i_13_297_862_0,
    i_13_297_895_0, i_13_297_951_0, i_13_297_952_0, i_13_297_1066_0,
    i_13_297_1075_0, i_13_297_1221_0, i_13_297_1222_0, i_13_297_1275_0,
    i_13_297_1293_0, i_13_297_1390_0, i_13_297_1410_0, i_13_297_1432_0,
    i_13_297_1491_0, i_13_297_1492_0, i_13_297_1627_0, i_13_297_1635_0,
    i_13_297_1641_0, i_13_297_1713_0, i_13_297_1726_0, i_13_297_1795_0,
    i_13_297_1842_0, i_13_297_1843_0, i_13_297_1884_0, i_13_297_1885_0,
    i_13_297_1929_0, i_13_297_1989_0, i_13_297_1993_0, i_13_297_2014_0,
    i_13_297_2028_0, i_13_297_2110_0, i_13_297_2175_0, i_13_297_2262_0,
    i_13_297_2410_0, i_13_297_2425_0, i_13_297_2463_0, i_13_297_2506_0,
    i_13_297_2535_0, i_13_297_2536_0, i_13_297_2616_0, i_13_297_2760_0,
    i_13_297_2847_0, i_13_297_2850_0, i_13_297_2851_0, i_13_297_3097_0,
    i_13_297_3345_0, i_13_297_3384_0, i_13_297_3387_0, i_13_297_3418_0,
    i_13_297_3426_0, i_13_297_3504_0, i_13_297_3505_0, i_13_297_3594_0,
    i_13_297_3669_0, i_13_297_3706_0, i_13_297_3766_0, i_13_297_3838_0,
    i_13_297_3876_0, i_13_297_3895_0, i_13_297_3931_0, i_13_297_4003_0,
    i_13_297_4011_0, i_13_297_4048_0, i_13_297_4080_0, i_13_297_4081_0,
    i_13_297_4086_0, i_13_297_4087_0, i_13_297_4114_0, i_13_297_4189_0,
    i_13_297_4210_0, i_13_297_4218_0, i_13_297_4273_0, i_13_297_4296_0,
    i_13_297_4297_0, i_13_297_4315_0, i_13_297_4543_0, i_13_297_4557_0;
  output o_13_297_0_0;
  assign o_13_297_0_0 = ~((~i_13_297_2851_0 & ((~i_13_297_3876_0 & ~i_13_297_4080_0) | (i_13_297_69_0 & ~i_13_297_4218_0))) | (~i_13_297_1221_0 & ~i_13_297_3876_0) | (~i_13_297_3426_0 & ~i_13_297_3931_0) | (i_13_297_1075_0 & ~i_13_297_1275_0 & ~i_13_297_4011_0));
endmodule



// Benchmark "kernel_13_298" written by ABC on Sun Jul 19 10:49:32 2020

module kernel_13_298 ( 
    i_13_298_31_0, i_13_298_39_0, i_13_298_63_0, i_13_298_64_0,
    i_13_298_98_0, i_13_298_128_0, i_13_298_137_0, i_13_298_175_0,
    i_13_298_184_0, i_13_298_214_0, i_13_298_229_0, i_13_298_269_0,
    i_13_298_279_0, i_13_298_280_0, i_13_298_306_0, i_13_298_323_0,
    i_13_298_337_0, i_13_298_352_0, i_13_298_379_0, i_13_298_525_0,
    i_13_298_605_0, i_13_298_616_0, i_13_298_683_0, i_13_298_768_0,
    i_13_298_824_0, i_13_298_1066_0, i_13_298_1070_0, i_13_298_1142_0,
    i_13_298_1150_0, i_13_298_1216_0, i_13_298_1218_0, i_13_298_1306_0,
    i_13_298_1309_0, i_13_298_1326_0, i_13_298_1553_0, i_13_298_1561_0,
    i_13_298_1570_0, i_13_298_1593_0, i_13_298_1594_0, i_13_298_1604_0,
    i_13_298_1638_0, i_13_298_1720_0, i_13_298_1748_0, i_13_298_1792_0,
    i_13_298_1804_0, i_13_298_1831_0, i_13_298_1835_0, i_13_298_1847_0,
    i_13_298_1882_0, i_13_298_1930_0, i_13_298_1998_0, i_13_298_1999_0,
    i_13_298_2233_0, i_13_298_2267_0, i_13_298_2407_0, i_13_298_2426_0,
    i_13_298_2429_0, i_13_298_2505_0, i_13_298_2657_0, i_13_298_2673_0,
    i_13_298_2677_0, i_13_298_2718_0, i_13_298_2739_0, i_13_298_2740_0,
    i_13_298_2853_0, i_13_298_2856_0, i_13_298_2872_0, i_13_298_2986_0,
    i_13_298_3028_0, i_13_298_3073_0, i_13_298_3141_0, i_13_298_3149_0,
    i_13_298_3211_0, i_13_298_3446_0, i_13_298_3488_0, i_13_298_3501_0,
    i_13_298_3502_0, i_13_298_3523_0, i_13_298_3538_0, i_13_298_3539_0,
    i_13_298_3541_0, i_13_298_3609_0, i_13_298_3638_0, i_13_298_3641_0,
    i_13_298_3727_0, i_13_298_3728_0, i_13_298_3857_0, i_13_298_3860_0,
    i_13_298_3934_0, i_13_298_4022_0, i_13_298_4063_0, i_13_298_4085_0,
    i_13_298_4121_0, i_13_298_4126_0, i_13_298_4162_0, i_13_298_4315_0,
    i_13_298_4318_0, i_13_298_4355_0, i_13_298_4395_0, i_13_298_4570_0,
    o_13_298_0_0  );
  input  i_13_298_31_0, i_13_298_39_0, i_13_298_63_0, i_13_298_64_0,
    i_13_298_98_0, i_13_298_128_0, i_13_298_137_0, i_13_298_175_0,
    i_13_298_184_0, i_13_298_214_0, i_13_298_229_0, i_13_298_269_0,
    i_13_298_279_0, i_13_298_280_0, i_13_298_306_0, i_13_298_323_0,
    i_13_298_337_0, i_13_298_352_0, i_13_298_379_0, i_13_298_525_0,
    i_13_298_605_0, i_13_298_616_0, i_13_298_683_0, i_13_298_768_0,
    i_13_298_824_0, i_13_298_1066_0, i_13_298_1070_0, i_13_298_1142_0,
    i_13_298_1150_0, i_13_298_1216_0, i_13_298_1218_0, i_13_298_1306_0,
    i_13_298_1309_0, i_13_298_1326_0, i_13_298_1553_0, i_13_298_1561_0,
    i_13_298_1570_0, i_13_298_1593_0, i_13_298_1594_0, i_13_298_1604_0,
    i_13_298_1638_0, i_13_298_1720_0, i_13_298_1748_0, i_13_298_1792_0,
    i_13_298_1804_0, i_13_298_1831_0, i_13_298_1835_0, i_13_298_1847_0,
    i_13_298_1882_0, i_13_298_1930_0, i_13_298_1998_0, i_13_298_1999_0,
    i_13_298_2233_0, i_13_298_2267_0, i_13_298_2407_0, i_13_298_2426_0,
    i_13_298_2429_0, i_13_298_2505_0, i_13_298_2657_0, i_13_298_2673_0,
    i_13_298_2677_0, i_13_298_2718_0, i_13_298_2739_0, i_13_298_2740_0,
    i_13_298_2853_0, i_13_298_2856_0, i_13_298_2872_0, i_13_298_2986_0,
    i_13_298_3028_0, i_13_298_3073_0, i_13_298_3141_0, i_13_298_3149_0,
    i_13_298_3211_0, i_13_298_3446_0, i_13_298_3488_0, i_13_298_3501_0,
    i_13_298_3502_0, i_13_298_3523_0, i_13_298_3538_0, i_13_298_3539_0,
    i_13_298_3541_0, i_13_298_3609_0, i_13_298_3638_0, i_13_298_3641_0,
    i_13_298_3727_0, i_13_298_3728_0, i_13_298_3857_0, i_13_298_3860_0,
    i_13_298_3934_0, i_13_298_4022_0, i_13_298_4063_0, i_13_298_4085_0,
    i_13_298_4121_0, i_13_298_4126_0, i_13_298_4162_0, i_13_298_4315_0,
    i_13_298_4318_0, i_13_298_4355_0, i_13_298_4395_0, i_13_298_4570_0;
  output o_13_298_0_0;
  assign o_13_298_0_0 = ~((~i_13_298_525_0 & ~i_13_298_3538_0 & ((i_13_298_337_0 & i_13_298_616_0 & ~i_13_298_1594_0 & ~i_13_298_1999_0) | (~i_13_298_64_0 & ~i_13_298_1070_0 & ~i_13_298_1150_0 & ~i_13_298_2673_0))) | (~i_13_298_683_0 & ((~i_13_298_63_0 & ~i_13_298_137_0 & ~i_13_298_3149_0 & ~i_13_298_3501_0 & ~i_13_298_3502_0) | (i_13_298_616_0 & i_13_298_4355_0))) | (~i_13_298_1309_0 & ((i_13_298_1831_0 & i_13_298_4162_0) | (~i_13_298_2429_0 & ~i_13_298_2673_0 & ~i_13_298_4395_0))) | (i_13_298_3523_0 & (i_13_298_4085_0 | (~i_13_298_184_0 & ~i_13_298_1847_0 & i_13_298_4162_0))) | (~i_13_298_1593_0 & i_13_298_1804_0 & ~i_13_298_1999_0 & ~i_13_298_2426_0));
endmodule



// Benchmark "kernel_13_299" written by ABC on Sun Jul 19 10:49:32 2020

module kernel_13_299 ( 
    i_13_299_31_0, i_13_299_58_0, i_13_299_64_0, i_13_299_103_0,
    i_13_299_104_0, i_13_299_130_0, i_13_299_162_0, i_13_299_184_0,
    i_13_299_237_0, i_13_299_307_0, i_13_299_553_0, i_13_299_556_0,
    i_13_299_586_0, i_13_299_598_0, i_13_299_612_0, i_13_299_684_0,
    i_13_299_693_0, i_13_299_814_0, i_13_299_822_0, i_13_299_828_0,
    i_13_299_837_0, i_13_299_1065_0, i_13_299_1066_0, i_13_299_1117_0,
    i_13_299_1120_0, i_13_299_1206_0, i_13_299_1213_0, i_13_299_1305_0,
    i_13_299_1306_0, i_13_299_1309_0, i_13_299_1387_0, i_13_299_1390_0,
    i_13_299_1425_0, i_13_299_1507_0, i_13_299_1624_0, i_13_299_1639_0,
    i_13_299_1644_0, i_13_299_1648_0, i_13_299_1669_0, i_13_299_1741_0,
    i_13_299_1846_0, i_13_299_1926_0, i_13_299_1927_0, i_13_299_1957_0,
    i_13_299_2008_0, i_13_299_2100_0, i_13_299_2142_0, i_13_299_2143_0,
    i_13_299_2188_0, i_13_299_2199_0, i_13_299_2377_0, i_13_299_2380_0,
    i_13_299_2407_0, i_13_299_2461_0, i_13_299_2462_0, i_13_299_2676_0,
    i_13_299_2692_0, i_13_299_2718_0, i_13_299_2754_0, i_13_299_2848_0,
    i_13_299_2858_0, i_13_299_2881_0, i_13_299_2935_0, i_13_299_2938_0,
    i_13_299_3009_0, i_13_299_3047_0, i_13_299_3205_0, i_13_299_3208_0,
    i_13_299_3486_0, i_13_299_3537_0, i_13_299_3637_0, i_13_299_3719_0,
    i_13_299_3738_0, i_13_299_3753_0, i_13_299_3754_0, i_13_299_3853_0,
    i_13_299_3907_0, i_13_299_3910_0, i_13_299_3924_0, i_13_299_3927_0,
    i_13_299_3928_0, i_13_299_3936_0, i_13_299_4032_0, i_13_299_4033_0,
    i_13_299_4034_0, i_13_299_4035_0, i_13_299_4063_0, i_13_299_4214_0,
    i_13_299_4216_0, i_13_299_4294_0, i_13_299_4311_0, i_13_299_4315_0,
    i_13_299_4318_0, i_13_299_4325_0, i_13_299_4330_0, i_13_299_4341_0,
    i_13_299_4509_0, i_13_299_4522_0, i_13_299_4591_0, i_13_299_4593_0,
    o_13_299_0_0  );
  input  i_13_299_31_0, i_13_299_58_0, i_13_299_64_0, i_13_299_103_0,
    i_13_299_104_0, i_13_299_130_0, i_13_299_162_0, i_13_299_184_0,
    i_13_299_237_0, i_13_299_307_0, i_13_299_553_0, i_13_299_556_0,
    i_13_299_586_0, i_13_299_598_0, i_13_299_612_0, i_13_299_684_0,
    i_13_299_693_0, i_13_299_814_0, i_13_299_822_0, i_13_299_828_0,
    i_13_299_837_0, i_13_299_1065_0, i_13_299_1066_0, i_13_299_1117_0,
    i_13_299_1120_0, i_13_299_1206_0, i_13_299_1213_0, i_13_299_1305_0,
    i_13_299_1306_0, i_13_299_1309_0, i_13_299_1387_0, i_13_299_1390_0,
    i_13_299_1425_0, i_13_299_1507_0, i_13_299_1624_0, i_13_299_1639_0,
    i_13_299_1644_0, i_13_299_1648_0, i_13_299_1669_0, i_13_299_1741_0,
    i_13_299_1846_0, i_13_299_1926_0, i_13_299_1927_0, i_13_299_1957_0,
    i_13_299_2008_0, i_13_299_2100_0, i_13_299_2142_0, i_13_299_2143_0,
    i_13_299_2188_0, i_13_299_2199_0, i_13_299_2377_0, i_13_299_2380_0,
    i_13_299_2407_0, i_13_299_2461_0, i_13_299_2462_0, i_13_299_2676_0,
    i_13_299_2692_0, i_13_299_2718_0, i_13_299_2754_0, i_13_299_2848_0,
    i_13_299_2858_0, i_13_299_2881_0, i_13_299_2935_0, i_13_299_2938_0,
    i_13_299_3009_0, i_13_299_3047_0, i_13_299_3205_0, i_13_299_3208_0,
    i_13_299_3486_0, i_13_299_3537_0, i_13_299_3637_0, i_13_299_3719_0,
    i_13_299_3738_0, i_13_299_3753_0, i_13_299_3754_0, i_13_299_3853_0,
    i_13_299_3907_0, i_13_299_3910_0, i_13_299_3924_0, i_13_299_3927_0,
    i_13_299_3928_0, i_13_299_3936_0, i_13_299_4032_0, i_13_299_4033_0,
    i_13_299_4034_0, i_13_299_4035_0, i_13_299_4063_0, i_13_299_4214_0,
    i_13_299_4216_0, i_13_299_4294_0, i_13_299_4311_0, i_13_299_4315_0,
    i_13_299_4318_0, i_13_299_4325_0, i_13_299_4330_0, i_13_299_4341_0,
    i_13_299_4509_0, i_13_299_4522_0, i_13_299_4591_0, i_13_299_4593_0;
  output o_13_299_0_0;
  assign o_13_299_0_0 = ~((~i_13_299_1507_0 & ((~i_13_299_64_0 & ~i_13_299_822_0 & ~i_13_299_3009_0) | (~i_13_299_3754_0 & ~i_13_299_4311_0 & ~i_13_299_4330_0))) | (~i_13_299_693_0 & ~i_13_299_2377_0 & ~i_13_299_3754_0) | (~i_13_299_837_0 & ~i_13_299_1306_0 & i_13_299_3205_0) | (i_13_299_1624_0 & ~i_13_299_4035_0 & ~i_13_299_4214_0) | (~i_13_299_58_0 & ~i_13_299_2881_0 & i_13_299_4325_0));
endmodule



// Benchmark "kernel_13_300" written by ABC on Sun Jul 19 10:49:33 2020

module kernel_13_300 ( 
    i_13_300_91_0, i_13_300_93_0, i_13_300_94_0, i_13_300_95_0,
    i_13_300_121_0, i_13_300_125_0, i_13_300_165_0, i_13_300_184_0,
    i_13_300_238_0, i_13_300_309_0, i_13_300_367_0, i_13_300_564_0,
    i_13_300_571_0, i_13_300_572_0, i_13_300_697_0, i_13_300_730_0,
    i_13_300_733_0, i_13_300_793_0, i_13_300_797_0, i_13_300_859_0,
    i_13_300_1120_0, i_13_300_1179_0, i_13_300_1180_0, i_13_300_1188_0,
    i_13_300_1210_0, i_13_300_1218_0, i_13_300_1273_0, i_13_300_1390_0,
    i_13_300_1408_0, i_13_300_1441_0, i_13_300_1489_0, i_13_300_1624_0,
    i_13_300_1632_0, i_13_300_1660_0, i_13_300_1683_0, i_13_300_1786_0,
    i_13_300_1832_0, i_13_300_1843_0, i_13_300_1844_0, i_13_300_1921_0,
    i_13_300_2088_0, i_13_300_2127_0, i_13_300_2128_0, i_13_300_2169_0,
    i_13_300_2173_0, i_13_300_2175_0, i_13_300_2176_0, i_13_300_2208_0,
    i_13_300_2209_0, i_13_300_2237_0, i_13_300_2380_0, i_13_300_2424_0,
    i_13_300_2425_0, i_13_300_2426_0, i_13_300_2427_0, i_13_300_2428_0,
    i_13_300_2446_0, i_13_300_2533_0, i_13_300_2541_0, i_13_300_2542_0,
    i_13_300_2551_0, i_13_300_2567_0, i_13_300_2614_0, i_13_300_2652_0,
    i_13_300_2722_0, i_13_300_2848_0, i_13_300_2884_0, i_13_300_2985_0,
    i_13_300_3109_0, i_13_300_3112_0, i_13_300_3147_0, i_13_300_3163_0,
    i_13_300_3165_0, i_13_300_3211_0, i_13_300_3216_0, i_13_300_3348_0,
    i_13_300_3373_0, i_13_300_3388_0, i_13_300_3390_0, i_13_300_3424_0,
    i_13_300_3425_0, i_13_300_3532_0, i_13_300_3732_0, i_13_300_3767_0,
    i_13_300_3846_0, i_13_300_3870_0, i_13_300_3872_0, i_13_300_3874_0,
    i_13_300_3875_0, i_13_300_4006_0, i_13_300_4008_0, i_13_300_4121_0,
    i_13_300_4189_0, i_13_300_4346_0, i_13_300_4351_0, i_13_300_4353_0,
    i_13_300_4354_0, i_13_300_4355_0, i_13_300_4570_0, i_13_300_4579_0,
    o_13_300_0_0  );
  input  i_13_300_91_0, i_13_300_93_0, i_13_300_94_0, i_13_300_95_0,
    i_13_300_121_0, i_13_300_125_0, i_13_300_165_0, i_13_300_184_0,
    i_13_300_238_0, i_13_300_309_0, i_13_300_367_0, i_13_300_564_0,
    i_13_300_571_0, i_13_300_572_0, i_13_300_697_0, i_13_300_730_0,
    i_13_300_733_0, i_13_300_793_0, i_13_300_797_0, i_13_300_859_0,
    i_13_300_1120_0, i_13_300_1179_0, i_13_300_1180_0, i_13_300_1188_0,
    i_13_300_1210_0, i_13_300_1218_0, i_13_300_1273_0, i_13_300_1390_0,
    i_13_300_1408_0, i_13_300_1441_0, i_13_300_1489_0, i_13_300_1624_0,
    i_13_300_1632_0, i_13_300_1660_0, i_13_300_1683_0, i_13_300_1786_0,
    i_13_300_1832_0, i_13_300_1843_0, i_13_300_1844_0, i_13_300_1921_0,
    i_13_300_2088_0, i_13_300_2127_0, i_13_300_2128_0, i_13_300_2169_0,
    i_13_300_2173_0, i_13_300_2175_0, i_13_300_2176_0, i_13_300_2208_0,
    i_13_300_2209_0, i_13_300_2237_0, i_13_300_2380_0, i_13_300_2424_0,
    i_13_300_2425_0, i_13_300_2426_0, i_13_300_2427_0, i_13_300_2428_0,
    i_13_300_2446_0, i_13_300_2533_0, i_13_300_2541_0, i_13_300_2542_0,
    i_13_300_2551_0, i_13_300_2567_0, i_13_300_2614_0, i_13_300_2652_0,
    i_13_300_2722_0, i_13_300_2848_0, i_13_300_2884_0, i_13_300_2985_0,
    i_13_300_3109_0, i_13_300_3112_0, i_13_300_3147_0, i_13_300_3163_0,
    i_13_300_3165_0, i_13_300_3211_0, i_13_300_3216_0, i_13_300_3348_0,
    i_13_300_3373_0, i_13_300_3388_0, i_13_300_3390_0, i_13_300_3424_0,
    i_13_300_3425_0, i_13_300_3532_0, i_13_300_3732_0, i_13_300_3767_0,
    i_13_300_3846_0, i_13_300_3870_0, i_13_300_3872_0, i_13_300_3874_0,
    i_13_300_3875_0, i_13_300_4006_0, i_13_300_4008_0, i_13_300_4121_0,
    i_13_300_4189_0, i_13_300_4346_0, i_13_300_4351_0, i_13_300_4353_0,
    i_13_300_4354_0, i_13_300_4355_0, i_13_300_4570_0, i_13_300_4579_0;
  output o_13_300_0_0;
  assign o_13_300_0_0 = ~((~i_13_300_4353_0 & (i_13_300_2884_0 | ~i_13_300_3211_0)) | (i_13_300_4355_0 & (~i_13_300_1408_0 | ~i_13_300_2428_0)) | i_13_300_1273_0 | (~i_13_300_1844_0 & ~i_13_300_2541_0) | (~i_13_300_184_0 & ~i_13_300_4008_0));
endmodule



// Benchmark "kernel_13_301" written by ABC on Sun Jul 19 10:49:34 2020

module kernel_13_301 ( 
    i_13_301_124_0, i_13_301_143_0, i_13_301_187_0, i_13_301_188_0,
    i_13_301_229_0, i_13_301_283_0, i_13_301_287_0, i_13_301_340_0,
    i_13_301_374_0, i_13_301_446_0, i_13_301_508_0, i_13_301_535_0,
    i_13_301_536_0, i_13_301_543_0, i_13_301_548_0, i_13_301_571_0,
    i_13_301_574_0, i_13_301_580_0, i_13_301_594_0, i_13_301_599_0,
    i_13_301_616_0, i_13_301_644_0, i_13_301_718_0, i_13_301_728_0,
    i_13_301_777_0, i_13_301_781_0, i_13_301_845_0, i_13_301_895_0,
    i_13_301_914_0, i_13_301_941_0, i_13_301_1069_0, i_13_301_1231_0,
    i_13_301_1249_0, i_13_301_1435_0, i_13_301_1439_0, i_13_301_1444_0,
    i_13_301_1465_0, i_13_301_1484_0, i_13_301_1499_0, i_13_301_1502_0,
    i_13_301_1543_0, i_13_301_1634_0, i_13_301_1636_0, i_13_301_1643_0,
    i_13_301_1694_0, i_13_301_1724_0, i_13_301_1742_0, i_13_301_1750_0,
    i_13_301_1762_0, i_13_301_1771_0, i_13_301_1772_0, i_13_301_1796_0,
    i_13_301_1804_0, i_13_301_1827_0, i_13_301_1853_0, i_13_301_1912_0,
    i_13_301_1930_0, i_13_301_2150_0, i_13_301_2168_0, i_13_301_2183_0,
    i_13_301_2200_0, i_13_301_2201_0, i_13_301_2228_0, i_13_301_2264_0,
    i_13_301_2311_0, i_13_301_2425_0, i_13_301_2510_0, i_13_301_2542_0,
    i_13_301_2554_0, i_13_301_2579_0, i_13_301_2633_0, i_13_301_2650_0,
    i_13_301_2660_0, i_13_301_2695_0, i_13_301_2848_0, i_13_301_2917_0,
    i_13_301_2920_0, i_13_301_3131_0, i_13_301_3169_0, i_13_301_3220_0,
    i_13_301_3221_0, i_13_301_3433_0, i_13_301_3523_0, i_13_301_3536_0,
    i_13_301_3636_0, i_13_301_3722_0, i_13_301_3794_0, i_13_301_3839_0,
    i_13_301_3901_0, i_13_301_4012_0, i_13_301_4013_0, i_13_301_4193_0,
    i_13_301_4238_0, i_13_301_4271_0, i_13_301_4408_0, i_13_301_4444_0,
    i_13_301_4526_0, i_13_301_4544_0, i_13_301_4586_0, i_13_301_4588_0,
    o_13_301_0_0  );
  input  i_13_301_124_0, i_13_301_143_0, i_13_301_187_0, i_13_301_188_0,
    i_13_301_229_0, i_13_301_283_0, i_13_301_287_0, i_13_301_340_0,
    i_13_301_374_0, i_13_301_446_0, i_13_301_508_0, i_13_301_535_0,
    i_13_301_536_0, i_13_301_543_0, i_13_301_548_0, i_13_301_571_0,
    i_13_301_574_0, i_13_301_580_0, i_13_301_594_0, i_13_301_599_0,
    i_13_301_616_0, i_13_301_644_0, i_13_301_718_0, i_13_301_728_0,
    i_13_301_777_0, i_13_301_781_0, i_13_301_845_0, i_13_301_895_0,
    i_13_301_914_0, i_13_301_941_0, i_13_301_1069_0, i_13_301_1231_0,
    i_13_301_1249_0, i_13_301_1435_0, i_13_301_1439_0, i_13_301_1444_0,
    i_13_301_1465_0, i_13_301_1484_0, i_13_301_1499_0, i_13_301_1502_0,
    i_13_301_1543_0, i_13_301_1634_0, i_13_301_1636_0, i_13_301_1643_0,
    i_13_301_1694_0, i_13_301_1724_0, i_13_301_1742_0, i_13_301_1750_0,
    i_13_301_1762_0, i_13_301_1771_0, i_13_301_1772_0, i_13_301_1796_0,
    i_13_301_1804_0, i_13_301_1827_0, i_13_301_1853_0, i_13_301_1912_0,
    i_13_301_1930_0, i_13_301_2150_0, i_13_301_2168_0, i_13_301_2183_0,
    i_13_301_2200_0, i_13_301_2201_0, i_13_301_2228_0, i_13_301_2264_0,
    i_13_301_2311_0, i_13_301_2425_0, i_13_301_2510_0, i_13_301_2542_0,
    i_13_301_2554_0, i_13_301_2579_0, i_13_301_2633_0, i_13_301_2650_0,
    i_13_301_2660_0, i_13_301_2695_0, i_13_301_2848_0, i_13_301_2917_0,
    i_13_301_2920_0, i_13_301_3131_0, i_13_301_3169_0, i_13_301_3220_0,
    i_13_301_3221_0, i_13_301_3433_0, i_13_301_3523_0, i_13_301_3536_0,
    i_13_301_3636_0, i_13_301_3722_0, i_13_301_3794_0, i_13_301_3839_0,
    i_13_301_3901_0, i_13_301_4012_0, i_13_301_4013_0, i_13_301_4193_0,
    i_13_301_4238_0, i_13_301_4271_0, i_13_301_4408_0, i_13_301_4444_0,
    i_13_301_4526_0, i_13_301_4544_0, i_13_301_4586_0, i_13_301_4588_0;
  output o_13_301_0_0;
  assign o_13_301_0_0 = 0;
endmodule



// Benchmark "kernel_13_302" written by ABC on Sun Jul 19 10:49:35 2020

module kernel_13_302 ( 
    i_13_302_29_0, i_13_302_48_0, i_13_302_69_0, i_13_302_70_0,
    i_13_302_124_0, i_13_302_140_0, i_13_302_160_0, i_13_302_231_0,
    i_13_302_240_0, i_13_302_245_0, i_13_302_313_0, i_13_302_380_0,
    i_13_302_385_0, i_13_302_447_0, i_13_302_610_0, i_13_302_645_0,
    i_13_302_688_0, i_13_302_742_0, i_13_302_762_0, i_13_302_870_0,
    i_13_302_1020_0, i_13_302_1069_0, i_13_302_1084_0, i_13_302_1086_0,
    i_13_302_1104_0, i_13_302_1123_0, i_13_302_1132_0, i_13_302_1218_0,
    i_13_302_1221_0, i_13_302_1257_0, i_13_302_1276_0, i_13_302_1312_0,
    i_13_302_1441_0, i_13_302_1444_0, i_13_302_1507_0, i_13_302_1510_0,
    i_13_302_1522_0, i_13_302_1529_0, i_13_302_1598_0, i_13_302_1609_0,
    i_13_302_1626_0, i_13_302_1716_0, i_13_302_1726_0, i_13_302_1798_0,
    i_13_302_1803_0, i_13_302_1887_0, i_13_302_1932_0, i_13_302_1933_0,
    i_13_302_1939_0, i_13_302_1947_0, i_13_302_1995_0, i_13_302_2001_0,
    i_13_302_2032_0, i_13_302_2122_0, i_13_302_2175_0, i_13_302_2193_0,
    i_13_302_2194_0, i_13_302_2235_0, i_13_302_2236_0, i_13_302_2266_0,
    i_13_302_2459_0, i_13_302_2472_0, i_13_302_2679_0, i_13_302_2680_0,
    i_13_302_2697_0, i_13_302_2724_0, i_13_302_2748_0, i_13_302_2757_0,
    i_13_302_2810_0, i_13_302_2855_0, i_13_302_2929_0, i_13_302_3003_0,
    i_13_302_3031_0, i_13_302_3044_0, i_13_302_3147_0, i_13_302_3211_0,
    i_13_302_3290_0, i_13_302_3370_0, i_13_302_3417_0, i_13_302_3418_0,
    i_13_302_3553_0, i_13_302_3616_0, i_13_302_3637_0, i_13_302_3640_0,
    i_13_302_3796_0, i_13_302_3822_0, i_13_302_3823_0, i_13_302_3891_0,
    i_13_302_3892_0, i_13_302_3930_0, i_13_302_4038_0, i_13_302_4039_0,
    i_13_302_4056_0, i_13_302_4083_0, i_13_302_4084_0, i_13_302_4308_0,
    i_13_302_4312_0, i_13_302_4596_0, i_13_302_4597_0, i_13_302_4606_0,
    o_13_302_0_0  );
  input  i_13_302_29_0, i_13_302_48_0, i_13_302_69_0, i_13_302_70_0,
    i_13_302_124_0, i_13_302_140_0, i_13_302_160_0, i_13_302_231_0,
    i_13_302_240_0, i_13_302_245_0, i_13_302_313_0, i_13_302_380_0,
    i_13_302_385_0, i_13_302_447_0, i_13_302_610_0, i_13_302_645_0,
    i_13_302_688_0, i_13_302_742_0, i_13_302_762_0, i_13_302_870_0,
    i_13_302_1020_0, i_13_302_1069_0, i_13_302_1084_0, i_13_302_1086_0,
    i_13_302_1104_0, i_13_302_1123_0, i_13_302_1132_0, i_13_302_1218_0,
    i_13_302_1221_0, i_13_302_1257_0, i_13_302_1276_0, i_13_302_1312_0,
    i_13_302_1441_0, i_13_302_1444_0, i_13_302_1507_0, i_13_302_1510_0,
    i_13_302_1522_0, i_13_302_1529_0, i_13_302_1598_0, i_13_302_1609_0,
    i_13_302_1626_0, i_13_302_1716_0, i_13_302_1726_0, i_13_302_1798_0,
    i_13_302_1803_0, i_13_302_1887_0, i_13_302_1932_0, i_13_302_1933_0,
    i_13_302_1939_0, i_13_302_1947_0, i_13_302_1995_0, i_13_302_2001_0,
    i_13_302_2032_0, i_13_302_2122_0, i_13_302_2175_0, i_13_302_2193_0,
    i_13_302_2194_0, i_13_302_2235_0, i_13_302_2236_0, i_13_302_2266_0,
    i_13_302_2459_0, i_13_302_2472_0, i_13_302_2679_0, i_13_302_2680_0,
    i_13_302_2697_0, i_13_302_2724_0, i_13_302_2748_0, i_13_302_2757_0,
    i_13_302_2810_0, i_13_302_2855_0, i_13_302_2929_0, i_13_302_3003_0,
    i_13_302_3031_0, i_13_302_3044_0, i_13_302_3147_0, i_13_302_3211_0,
    i_13_302_3290_0, i_13_302_3370_0, i_13_302_3417_0, i_13_302_3418_0,
    i_13_302_3553_0, i_13_302_3616_0, i_13_302_3637_0, i_13_302_3640_0,
    i_13_302_3796_0, i_13_302_3822_0, i_13_302_3823_0, i_13_302_3891_0,
    i_13_302_3892_0, i_13_302_3930_0, i_13_302_4038_0, i_13_302_4039_0,
    i_13_302_4056_0, i_13_302_4083_0, i_13_302_4084_0, i_13_302_4308_0,
    i_13_302_4312_0, i_13_302_4596_0, i_13_302_4597_0, i_13_302_4606_0;
  output o_13_302_0_0;
  assign o_13_302_0_0 = ~((~i_13_302_4083_0 & ((~i_13_302_1123_0 & ~i_13_302_1510_0) | (~i_13_302_70_0 & ~i_13_302_1803_0))) | i_13_302_1529_0 | (i_13_302_1598_0 & ~i_13_302_3553_0) | (i_13_302_124_0 & ~i_13_302_3290_0 & ~i_13_302_4038_0 & ~i_13_302_4308_0));
endmodule



// Benchmark "kernel_13_303" written by ABC on Sun Jul 19 10:49:36 2020

module kernel_13_303 ( 
    i_13_303_103_0, i_13_303_105_0, i_13_303_106_0, i_13_303_159_0,
    i_13_303_160_0, i_13_303_175_0, i_13_303_227_0, i_13_303_339_0,
    i_13_303_357_0, i_13_303_372_0, i_13_303_421_0, i_13_303_456_0,
    i_13_303_457_0, i_13_303_471_0, i_13_303_486_0, i_13_303_492_0,
    i_13_303_696_0, i_13_303_697_0, i_13_303_735_0, i_13_303_797_0,
    i_13_303_825_0, i_13_303_949_0, i_13_303_1086_0, i_13_303_1131_0,
    i_13_303_1213_0, i_13_303_1299_0, i_13_303_1302_0, i_13_303_1303_0,
    i_13_303_1346_0, i_13_303_1347_0, i_13_303_1348_0, i_13_303_1437_0,
    i_13_303_1446_0, i_13_303_1463_0, i_13_303_1464_0, i_13_303_1473_0,
    i_13_303_1474_0, i_13_303_1528_0, i_13_303_1609_0, i_13_303_1721_0,
    i_13_303_1722_0, i_13_303_1743_0, i_13_303_1771_0, i_13_303_1815_0,
    i_13_303_1816_0, i_13_303_1883_0, i_13_303_1951_0, i_13_303_2031_0,
    i_13_303_2045_0, i_13_303_2056_0, i_13_303_2103_0, i_13_303_2110_0,
    i_13_303_2223_0, i_13_303_2238_0, i_13_303_2239_0, i_13_303_2378_0,
    i_13_303_2404_0, i_13_303_2407_0, i_13_303_2422_0, i_13_303_2445_0,
    i_13_303_2446_0, i_13_303_2553_0, i_13_303_2697_0, i_13_303_2715_0,
    i_13_303_2716_0, i_13_303_2823_0, i_13_303_2824_0, i_13_303_2846_0,
    i_13_303_2911_0, i_13_303_2922_0, i_13_303_3009_0, i_13_303_3058_0,
    i_13_303_3112_0, i_13_303_3219_0, i_13_303_3220_0, i_13_303_3255_0,
    i_13_303_3390_0, i_13_303_3391_0, i_13_303_3418_0, i_13_303_3420_0,
    i_13_303_3531_0, i_13_303_3595_0, i_13_303_3612_0, i_13_303_3621_0,
    i_13_303_3622_0, i_13_303_3706_0, i_13_303_3741_0, i_13_303_3985_0,
    i_13_303_3999_0, i_13_303_4042_0, i_13_303_4083_0, i_13_303_4092_0,
    i_13_303_4236_0, i_13_303_4237_0, i_13_303_4326_0, i_13_303_4327_0,
    i_13_303_4398_0, i_13_303_4512_0, i_13_303_4521_0, i_13_303_4567_0,
    o_13_303_0_0  );
  input  i_13_303_103_0, i_13_303_105_0, i_13_303_106_0, i_13_303_159_0,
    i_13_303_160_0, i_13_303_175_0, i_13_303_227_0, i_13_303_339_0,
    i_13_303_357_0, i_13_303_372_0, i_13_303_421_0, i_13_303_456_0,
    i_13_303_457_0, i_13_303_471_0, i_13_303_486_0, i_13_303_492_0,
    i_13_303_696_0, i_13_303_697_0, i_13_303_735_0, i_13_303_797_0,
    i_13_303_825_0, i_13_303_949_0, i_13_303_1086_0, i_13_303_1131_0,
    i_13_303_1213_0, i_13_303_1299_0, i_13_303_1302_0, i_13_303_1303_0,
    i_13_303_1346_0, i_13_303_1347_0, i_13_303_1348_0, i_13_303_1437_0,
    i_13_303_1446_0, i_13_303_1463_0, i_13_303_1464_0, i_13_303_1473_0,
    i_13_303_1474_0, i_13_303_1528_0, i_13_303_1609_0, i_13_303_1721_0,
    i_13_303_1722_0, i_13_303_1743_0, i_13_303_1771_0, i_13_303_1815_0,
    i_13_303_1816_0, i_13_303_1883_0, i_13_303_1951_0, i_13_303_2031_0,
    i_13_303_2045_0, i_13_303_2056_0, i_13_303_2103_0, i_13_303_2110_0,
    i_13_303_2223_0, i_13_303_2238_0, i_13_303_2239_0, i_13_303_2378_0,
    i_13_303_2404_0, i_13_303_2407_0, i_13_303_2422_0, i_13_303_2445_0,
    i_13_303_2446_0, i_13_303_2553_0, i_13_303_2697_0, i_13_303_2715_0,
    i_13_303_2716_0, i_13_303_2823_0, i_13_303_2824_0, i_13_303_2846_0,
    i_13_303_2911_0, i_13_303_2922_0, i_13_303_3009_0, i_13_303_3058_0,
    i_13_303_3112_0, i_13_303_3219_0, i_13_303_3220_0, i_13_303_3255_0,
    i_13_303_3390_0, i_13_303_3391_0, i_13_303_3418_0, i_13_303_3420_0,
    i_13_303_3531_0, i_13_303_3595_0, i_13_303_3612_0, i_13_303_3621_0,
    i_13_303_3622_0, i_13_303_3706_0, i_13_303_3741_0, i_13_303_3985_0,
    i_13_303_3999_0, i_13_303_4042_0, i_13_303_4083_0, i_13_303_4092_0,
    i_13_303_4236_0, i_13_303_4237_0, i_13_303_4326_0, i_13_303_4327_0,
    i_13_303_4398_0, i_13_303_4512_0, i_13_303_4521_0, i_13_303_4567_0;
  output o_13_303_0_0;
  assign o_13_303_0_0 = ~((~i_13_303_105_0 & ~i_13_303_1348_0) | (~i_13_303_357_0 & ~i_13_303_2922_0 & ~i_13_303_3531_0) | (~i_13_303_106_0 & i_13_303_175_0 & ~i_13_303_3391_0));
endmodule



// Benchmark "kernel_13_304" written by ABC on Sun Jul 19 10:49:37 2020

module kernel_13_304 ( 
    i_13_304_59_0, i_13_304_70_0, i_13_304_112_0, i_13_304_119_0,
    i_13_304_157_0, i_13_304_171_0, i_13_304_172_0, i_13_304_175_0,
    i_13_304_184_0, i_13_304_280_0, i_13_304_282_0, i_13_304_283_0,
    i_13_304_313_0, i_13_304_319_0, i_13_304_370_0, i_13_304_489_0,
    i_13_304_523_0, i_13_304_532_0, i_13_304_598_0, i_13_304_607_0,
    i_13_304_657_0, i_13_304_658_0, i_13_304_660_0, i_13_304_675_0,
    i_13_304_694_0, i_13_304_695_0, i_13_304_939_0, i_13_304_1018_0,
    i_13_304_1020_0, i_13_304_1066_0, i_13_304_1072_0, i_13_304_1074_0,
    i_13_304_1075_0, i_13_304_1206_0, i_13_304_1224_0, i_13_304_1225_0,
    i_13_304_1300_0, i_13_304_1305_0, i_13_304_1422_0, i_13_304_1423_0,
    i_13_304_1444_0, i_13_304_1494_0, i_13_304_1630_0, i_13_304_1631_0,
    i_13_304_1632_0, i_13_304_1633_0, i_13_304_1639_0, i_13_304_1657_0,
    i_13_304_1720_0, i_13_304_1729_0, i_13_304_1732_0, i_13_304_1779_0,
    i_13_304_1838_0, i_13_304_1936_0, i_13_304_1954_0, i_13_304_2196_0,
    i_13_304_2235_0, i_13_304_2377_0, i_13_304_2448_0, i_13_304_2449_0,
    i_13_304_2451_0, i_13_304_2452_0, i_13_304_3141_0, i_13_304_3142_0,
    i_13_304_3217_0, i_13_304_3244_0, i_13_304_3264_0, i_13_304_3388_0,
    i_13_304_3447_0, i_13_304_3483_0, i_13_304_3484_0, i_13_304_3538_0,
    i_13_304_3568_0, i_13_304_3574_0, i_13_304_3612_0, i_13_304_3726_0,
    i_13_304_3880_0, i_13_304_3888_0, i_13_304_3889_0, i_13_304_3994_0,
    i_13_304_4017_0, i_13_304_4086_0, i_13_304_4087_0, i_13_304_4186_0,
    i_13_304_4248_0, i_13_304_4249_0, i_13_304_4251_0, i_13_304_4252_0,
    i_13_304_4254_0, i_13_304_4258_0, i_13_304_4260_0, i_13_304_4261_0,
    i_13_304_4393_0, i_13_304_4415_0, i_13_304_4455_0, i_13_304_4521_0,
    i_13_304_4541_0, i_13_304_4554_0, i_13_304_4558_0, i_13_304_4591_0,
    o_13_304_0_0  );
  input  i_13_304_59_0, i_13_304_70_0, i_13_304_112_0, i_13_304_119_0,
    i_13_304_157_0, i_13_304_171_0, i_13_304_172_0, i_13_304_175_0,
    i_13_304_184_0, i_13_304_280_0, i_13_304_282_0, i_13_304_283_0,
    i_13_304_313_0, i_13_304_319_0, i_13_304_370_0, i_13_304_489_0,
    i_13_304_523_0, i_13_304_532_0, i_13_304_598_0, i_13_304_607_0,
    i_13_304_657_0, i_13_304_658_0, i_13_304_660_0, i_13_304_675_0,
    i_13_304_694_0, i_13_304_695_0, i_13_304_939_0, i_13_304_1018_0,
    i_13_304_1020_0, i_13_304_1066_0, i_13_304_1072_0, i_13_304_1074_0,
    i_13_304_1075_0, i_13_304_1206_0, i_13_304_1224_0, i_13_304_1225_0,
    i_13_304_1300_0, i_13_304_1305_0, i_13_304_1422_0, i_13_304_1423_0,
    i_13_304_1444_0, i_13_304_1494_0, i_13_304_1630_0, i_13_304_1631_0,
    i_13_304_1632_0, i_13_304_1633_0, i_13_304_1639_0, i_13_304_1657_0,
    i_13_304_1720_0, i_13_304_1729_0, i_13_304_1732_0, i_13_304_1779_0,
    i_13_304_1838_0, i_13_304_1936_0, i_13_304_1954_0, i_13_304_2196_0,
    i_13_304_2235_0, i_13_304_2377_0, i_13_304_2448_0, i_13_304_2449_0,
    i_13_304_2451_0, i_13_304_2452_0, i_13_304_3141_0, i_13_304_3142_0,
    i_13_304_3217_0, i_13_304_3244_0, i_13_304_3264_0, i_13_304_3388_0,
    i_13_304_3447_0, i_13_304_3483_0, i_13_304_3484_0, i_13_304_3538_0,
    i_13_304_3568_0, i_13_304_3574_0, i_13_304_3612_0, i_13_304_3726_0,
    i_13_304_3880_0, i_13_304_3888_0, i_13_304_3889_0, i_13_304_3994_0,
    i_13_304_4017_0, i_13_304_4086_0, i_13_304_4087_0, i_13_304_4186_0,
    i_13_304_4248_0, i_13_304_4249_0, i_13_304_4251_0, i_13_304_4252_0,
    i_13_304_4254_0, i_13_304_4258_0, i_13_304_4260_0, i_13_304_4261_0,
    i_13_304_4393_0, i_13_304_4415_0, i_13_304_4455_0, i_13_304_4521_0,
    i_13_304_4541_0, i_13_304_4554_0, i_13_304_4558_0, i_13_304_4591_0;
  output o_13_304_0_0;
  assign o_13_304_0_0 = ~((~i_13_304_1018_0 & ~i_13_304_3888_0) | (~i_13_304_2448_0 & ~i_13_304_2451_0) | (i_13_304_1300_0 & ~i_13_304_2196_0));
endmodule



// Benchmark "kernel_13_305" written by ABC on Sun Jul 19 10:49:38 2020

module kernel_13_305 ( 
    i_13_305_70_0, i_13_305_98_0, i_13_305_229_0, i_13_305_268_0,
    i_13_305_359_0, i_13_305_562_0, i_13_305_607_0, i_13_305_608_0,
    i_13_305_610_0, i_13_305_611_0, i_13_305_646_0, i_13_305_655_0,
    i_13_305_661_0, i_13_305_662_0, i_13_305_671_0, i_13_305_673_0,
    i_13_305_701_0, i_13_305_814_0, i_13_305_825_0, i_13_305_950_0,
    i_13_305_1024_0, i_13_305_1085_0, i_13_305_1102_0, i_13_305_1120_0,
    i_13_305_1123_0, i_13_305_1148_0, i_13_305_1167_0, i_13_305_1220_0,
    i_13_305_1430_0, i_13_305_1660_0, i_13_305_1661_0, i_13_305_1672_0,
    i_13_305_1727_0, i_13_305_1733_0, i_13_305_1735_0, i_13_305_1736_0,
    i_13_305_1745_0, i_13_305_1840_0, i_13_305_1841_0, i_13_305_1843_0,
    i_13_305_1844_0, i_13_305_1858_0, i_13_305_2020_0, i_13_305_2021_0,
    i_13_305_2024_0, i_13_305_2099_0, i_13_305_2137_0, i_13_305_2173_0,
    i_13_305_2348_0, i_13_305_2435_0, i_13_305_2471_0, i_13_305_2716_0,
    i_13_305_2787_0, i_13_305_2885_0, i_13_305_2902_0, i_13_305_2959_0,
    i_13_305_3029_0, i_13_305_3047_0, i_13_305_3050_0, i_13_305_3092_0,
    i_13_305_3100_0, i_13_305_3101_0, i_13_305_3145_0, i_13_305_3262_0,
    i_13_305_3352_0, i_13_305_3417_0, i_13_305_3479_0, i_13_305_3527_0,
    i_13_305_3613_0, i_13_305_3649_0, i_13_305_3662_0, i_13_305_3667_0,
    i_13_305_3730_0, i_13_305_3743_0, i_13_305_3751_0, i_13_305_3866_0,
    i_13_305_3896_0, i_13_305_3910_0, i_13_305_3911_0, i_13_305_3931_0,
    i_13_305_4063_0, i_13_305_4162_0, i_13_305_4163_0, i_13_305_4166_0,
    i_13_305_4189_0, i_13_305_4190_0, i_13_305_4192_0, i_13_305_4193_0,
    i_13_305_4294_0, i_13_305_4296_0, i_13_305_4297_0, i_13_305_4328_0,
    i_13_305_4343_0, i_13_305_4364_0, i_13_305_4530_0, i_13_305_4594_0,
    i_13_305_4597_0, i_13_305_4603_0, i_13_305_4604_0, i_13_305_4607_0,
    o_13_305_0_0  );
  input  i_13_305_70_0, i_13_305_98_0, i_13_305_229_0, i_13_305_268_0,
    i_13_305_359_0, i_13_305_562_0, i_13_305_607_0, i_13_305_608_0,
    i_13_305_610_0, i_13_305_611_0, i_13_305_646_0, i_13_305_655_0,
    i_13_305_661_0, i_13_305_662_0, i_13_305_671_0, i_13_305_673_0,
    i_13_305_701_0, i_13_305_814_0, i_13_305_825_0, i_13_305_950_0,
    i_13_305_1024_0, i_13_305_1085_0, i_13_305_1102_0, i_13_305_1120_0,
    i_13_305_1123_0, i_13_305_1148_0, i_13_305_1167_0, i_13_305_1220_0,
    i_13_305_1430_0, i_13_305_1660_0, i_13_305_1661_0, i_13_305_1672_0,
    i_13_305_1727_0, i_13_305_1733_0, i_13_305_1735_0, i_13_305_1736_0,
    i_13_305_1745_0, i_13_305_1840_0, i_13_305_1841_0, i_13_305_1843_0,
    i_13_305_1844_0, i_13_305_1858_0, i_13_305_2020_0, i_13_305_2021_0,
    i_13_305_2024_0, i_13_305_2099_0, i_13_305_2137_0, i_13_305_2173_0,
    i_13_305_2348_0, i_13_305_2435_0, i_13_305_2471_0, i_13_305_2716_0,
    i_13_305_2787_0, i_13_305_2885_0, i_13_305_2902_0, i_13_305_2959_0,
    i_13_305_3029_0, i_13_305_3047_0, i_13_305_3050_0, i_13_305_3092_0,
    i_13_305_3100_0, i_13_305_3101_0, i_13_305_3145_0, i_13_305_3262_0,
    i_13_305_3352_0, i_13_305_3417_0, i_13_305_3479_0, i_13_305_3527_0,
    i_13_305_3613_0, i_13_305_3649_0, i_13_305_3662_0, i_13_305_3667_0,
    i_13_305_3730_0, i_13_305_3743_0, i_13_305_3751_0, i_13_305_3866_0,
    i_13_305_3896_0, i_13_305_3910_0, i_13_305_3911_0, i_13_305_3931_0,
    i_13_305_4063_0, i_13_305_4162_0, i_13_305_4163_0, i_13_305_4166_0,
    i_13_305_4189_0, i_13_305_4190_0, i_13_305_4192_0, i_13_305_4193_0,
    i_13_305_4294_0, i_13_305_4296_0, i_13_305_4297_0, i_13_305_4328_0,
    i_13_305_4343_0, i_13_305_4364_0, i_13_305_4530_0, i_13_305_4594_0,
    i_13_305_4597_0, i_13_305_4603_0, i_13_305_4604_0, i_13_305_4607_0;
  output o_13_305_0_0;
  assign o_13_305_0_0 = ~((~i_13_305_359_0 & ((~i_13_305_1736_0 & ~i_13_305_2021_0) | (~i_13_305_1024_0 & i_13_305_1733_0 & ~i_13_305_3649_0 & i_13_305_4163_0))) | (~i_13_305_1085_0 & (~i_13_305_4193_0 | (~i_13_305_1660_0 & i_13_305_4190_0))) | (~i_13_305_1661_0 & ~i_13_305_1844_0) | (~i_13_305_950_0 & ~i_13_305_3751_0) | (~i_13_305_2021_0 & ~i_13_305_4328_0));
endmodule



// Benchmark "kernel_13_306" written by ABC on Sun Jul 19 10:49:38 2020

module kernel_13_306 ( 
    i_13_306_53_0, i_13_306_71_0, i_13_306_108_0, i_13_306_173_0,
    i_13_306_193_0, i_13_306_241_0, i_13_306_311_0, i_13_306_314_0,
    i_13_306_466_0, i_13_306_538_0, i_13_306_557_0, i_13_306_620_0,
    i_13_306_628_0, i_13_306_629_0, i_13_306_644_0, i_13_306_646_0,
    i_13_306_647_0, i_13_306_683_0, i_13_306_686_0, i_13_306_689_0,
    i_13_306_698_0, i_13_306_758_0, i_13_306_827_0, i_13_306_859_0,
    i_13_306_985_0, i_13_306_1066_0, i_13_306_1124_0, i_13_306_1133_0,
    i_13_306_1151_0, i_13_306_1228_0, i_13_306_1274_0, i_13_306_1277_0,
    i_13_306_1378_0, i_13_306_1394_0, i_13_306_1459_0, i_13_306_1484_0,
    i_13_306_1511_0, i_13_306_1549_0, i_13_306_1624_0, i_13_306_1645_0,
    i_13_306_1646_0, i_13_306_1660_0, i_13_306_1670_0, i_13_306_1673_0,
    i_13_306_1727_0, i_13_306_1745_0, i_13_306_1796_0, i_13_306_1798_0,
    i_13_306_1799_0, i_13_306_1889_0, i_13_306_1912_0, i_13_306_2119_0,
    i_13_306_2134_0, i_13_306_2384_0, i_13_306_2651_0, i_13_306_2654_0,
    i_13_306_2690_0, i_13_306_2851_0, i_13_306_2852_0, i_13_306_2876_0,
    i_13_306_2878_0, i_13_306_2906_0, i_13_306_2983_0, i_13_306_3095_0,
    i_13_306_3097_0, i_13_306_3131_0, i_13_306_3157_0, i_13_306_3265_0,
    i_13_306_3274_0, i_13_306_3343_0, i_13_306_3356_0, i_13_306_3397_0,
    i_13_306_3479_0, i_13_306_3575_0, i_13_306_3663_0, i_13_306_3742_0,
    i_13_306_3743_0, i_13_306_3785_0, i_13_306_3797_0, i_13_306_3842_0,
    i_13_306_3869_0, i_13_306_3896_0, i_13_306_3931_0, i_13_306_3941_0,
    i_13_306_3995_0, i_13_306_4033_0, i_13_306_4055_0, i_13_306_4059_0,
    i_13_306_4084_0, i_13_306_4085_0, i_13_306_4190_0, i_13_306_4297_0,
    i_13_306_4298_0, i_13_306_4301_0, i_13_306_4436_0, i_13_306_4448_0,
    i_13_306_4463_0, i_13_306_4530_0, i_13_306_4598_0, i_13_306_4607_0,
    o_13_306_0_0  );
  input  i_13_306_53_0, i_13_306_71_0, i_13_306_108_0, i_13_306_173_0,
    i_13_306_193_0, i_13_306_241_0, i_13_306_311_0, i_13_306_314_0,
    i_13_306_466_0, i_13_306_538_0, i_13_306_557_0, i_13_306_620_0,
    i_13_306_628_0, i_13_306_629_0, i_13_306_644_0, i_13_306_646_0,
    i_13_306_647_0, i_13_306_683_0, i_13_306_686_0, i_13_306_689_0,
    i_13_306_698_0, i_13_306_758_0, i_13_306_827_0, i_13_306_859_0,
    i_13_306_985_0, i_13_306_1066_0, i_13_306_1124_0, i_13_306_1133_0,
    i_13_306_1151_0, i_13_306_1228_0, i_13_306_1274_0, i_13_306_1277_0,
    i_13_306_1378_0, i_13_306_1394_0, i_13_306_1459_0, i_13_306_1484_0,
    i_13_306_1511_0, i_13_306_1549_0, i_13_306_1624_0, i_13_306_1645_0,
    i_13_306_1646_0, i_13_306_1660_0, i_13_306_1670_0, i_13_306_1673_0,
    i_13_306_1727_0, i_13_306_1745_0, i_13_306_1796_0, i_13_306_1798_0,
    i_13_306_1799_0, i_13_306_1889_0, i_13_306_1912_0, i_13_306_2119_0,
    i_13_306_2134_0, i_13_306_2384_0, i_13_306_2651_0, i_13_306_2654_0,
    i_13_306_2690_0, i_13_306_2851_0, i_13_306_2852_0, i_13_306_2876_0,
    i_13_306_2878_0, i_13_306_2906_0, i_13_306_2983_0, i_13_306_3095_0,
    i_13_306_3097_0, i_13_306_3131_0, i_13_306_3157_0, i_13_306_3265_0,
    i_13_306_3274_0, i_13_306_3343_0, i_13_306_3356_0, i_13_306_3397_0,
    i_13_306_3479_0, i_13_306_3575_0, i_13_306_3663_0, i_13_306_3742_0,
    i_13_306_3743_0, i_13_306_3785_0, i_13_306_3797_0, i_13_306_3842_0,
    i_13_306_3869_0, i_13_306_3896_0, i_13_306_3931_0, i_13_306_3941_0,
    i_13_306_3995_0, i_13_306_4033_0, i_13_306_4055_0, i_13_306_4059_0,
    i_13_306_4084_0, i_13_306_4085_0, i_13_306_4190_0, i_13_306_4297_0,
    i_13_306_4298_0, i_13_306_4301_0, i_13_306_4436_0, i_13_306_4448_0,
    i_13_306_4463_0, i_13_306_4530_0, i_13_306_4598_0, i_13_306_4607_0;
  output o_13_306_0_0;
  assign o_13_306_0_0 = ~(~i_13_306_1645_0 | ~i_13_306_2852_0);
endmodule



// Benchmark "kernel_13_307" written by ABC on Sun Jul 19 10:49:39 2020

module kernel_13_307 ( 
    i_13_307_31_0, i_13_307_32_0, i_13_307_64_0, i_13_307_121_0,
    i_13_307_207_0, i_13_307_208_0, i_13_307_307_0, i_13_307_374_0,
    i_13_307_399_0, i_13_307_412_0, i_13_307_489_0, i_13_307_524_0,
    i_13_307_586_0, i_13_307_598_0, i_13_307_612_0, i_13_307_613_0,
    i_13_307_671_0, i_13_307_715_0, i_13_307_738_0, i_13_307_759_0,
    i_13_307_760_0, i_13_307_796_0, i_13_307_829_0, i_13_307_1066_0,
    i_13_307_1121_0, i_13_307_1128_0, i_13_307_1129_0, i_13_307_1207_0,
    i_13_307_1223_0, i_13_307_1281_0, i_13_307_1286_0, i_13_307_1306_0,
    i_13_307_1372_0, i_13_307_1423_0, i_13_307_1441_0, i_13_307_1507_0,
    i_13_307_1523_0, i_13_307_1559_0, i_13_307_1562_0, i_13_307_1639_0,
    i_13_307_1696_0, i_13_307_1697_0, i_13_307_1720_0, i_13_307_1792_0,
    i_13_307_1795_0, i_13_307_1927_0, i_13_307_1928_0, i_13_307_1945_0,
    i_13_307_1964_0, i_13_307_2101_0, i_13_307_2126_0, i_13_307_2172_0,
    i_13_307_2200_0, i_13_307_2237_0, i_13_307_2351_0, i_13_307_2365_0,
    i_13_307_2377_0, i_13_307_2438_0, i_13_307_2542_0, i_13_307_2552_0,
    i_13_307_2593_0, i_13_307_2677_0, i_13_307_2719_0, i_13_307_2749_0,
    i_13_307_2759_0, i_13_307_2771_0, i_13_307_2857_0, i_13_307_2881_0,
    i_13_307_2882_0, i_13_307_3127_0, i_13_307_3172_0, i_13_307_3242_0,
    i_13_307_3269_0, i_13_307_3367_0, i_13_307_3438_0, i_13_307_3446_0,
    i_13_307_3572_0, i_13_307_3591_0, i_13_307_3605_0, i_13_307_3637_0,
    i_13_307_3638_0, i_13_307_3889_0, i_13_307_3910_0, i_13_307_3916_0,
    i_13_307_3925_0, i_13_307_3928_0, i_13_307_3934_0, i_13_307_4033_0,
    i_13_307_4034_0, i_13_307_4036_0, i_13_307_4042_0, i_13_307_4045_0,
    i_13_307_4052_0, i_13_307_4166_0, i_13_307_4313_0, i_13_307_4337_0,
    i_13_307_4494_0, i_13_307_4510_0, i_13_307_4522_0, i_13_307_4591_0,
    o_13_307_0_0  );
  input  i_13_307_31_0, i_13_307_32_0, i_13_307_64_0, i_13_307_121_0,
    i_13_307_207_0, i_13_307_208_0, i_13_307_307_0, i_13_307_374_0,
    i_13_307_399_0, i_13_307_412_0, i_13_307_489_0, i_13_307_524_0,
    i_13_307_586_0, i_13_307_598_0, i_13_307_612_0, i_13_307_613_0,
    i_13_307_671_0, i_13_307_715_0, i_13_307_738_0, i_13_307_759_0,
    i_13_307_760_0, i_13_307_796_0, i_13_307_829_0, i_13_307_1066_0,
    i_13_307_1121_0, i_13_307_1128_0, i_13_307_1129_0, i_13_307_1207_0,
    i_13_307_1223_0, i_13_307_1281_0, i_13_307_1286_0, i_13_307_1306_0,
    i_13_307_1372_0, i_13_307_1423_0, i_13_307_1441_0, i_13_307_1507_0,
    i_13_307_1523_0, i_13_307_1559_0, i_13_307_1562_0, i_13_307_1639_0,
    i_13_307_1696_0, i_13_307_1697_0, i_13_307_1720_0, i_13_307_1792_0,
    i_13_307_1795_0, i_13_307_1927_0, i_13_307_1928_0, i_13_307_1945_0,
    i_13_307_1964_0, i_13_307_2101_0, i_13_307_2126_0, i_13_307_2172_0,
    i_13_307_2200_0, i_13_307_2237_0, i_13_307_2351_0, i_13_307_2365_0,
    i_13_307_2377_0, i_13_307_2438_0, i_13_307_2542_0, i_13_307_2552_0,
    i_13_307_2593_0, i_13_307_2677_0, i_13_307_2719_0, i_13_307_2749_0,
    i_13_307_2759_0, i_13_307_2771_0, i_13_307_2857_0, i_13_307_2881_0,
    i_13_307_2882_0, i_13_307_3127_0, i_13_307_3172_0, i_13_307_3242_0,
    i_13_307_3269_0, i_13_307_3367_0, i_13_307_3438_0, i_13_307_3446_0,
    i_13_307_3572_0, i_13_307_3591_0, i_13_307_3605_0, i_13_307_3637_0,
    i_13_307_3638_0, i_13_307_3889_0, i_13_307_3910_0, i_13_307_3916_0,
    i_13_307_3925_0, i_13_307_3928_0, i_13_307_3934_0, i_13_307_4033_0,
    i_13_307_4034_0, i_13_307_4036_0, i_13_307_4042_0, i_13_307_4045_0,
    i_13_307_4052_0, i_13_307_4166_0, i_13_307_4313_0, i_13_307_4337_0,
    i_13_307_4494_0, i_13_307_4510_0, i_13_307_4522_0, i_13_307_4591_0;
  output o_13_307_0_0;
  assign o_13_307_0_0 = ~((~i_13_307_524_0 & ~i_13_307_3925_0 & ~i_13_307_4042_0) | (~i_13_307_1306_0 & ~i_13_307_2882_0 & ~i_13_307_3928_0 & ~i_13_307_4510_0) | (~i_13_307_64_0 & ~i_13_307_2881_0 & ~i_13_307_3438_0 & ~i_13_307_4313_0) | (~i_13_307_32_0 & ~i_13_307_613_0 & ~i_13_307_2200_0 & ~i_13_307_3242_0 & ~i_13_307_3591_0));
endmodule



// Benchmark "kernel_13_308" written by ABC on Sun Jul 19 10:49:40 2020

module kernel_13_308 ( 
    i_13_308_64_0, i_13_308_65_0, i_13_308_118_0, i_13_308_188_0,
    i_13_308_190_0, i_13_308_226_0, i_13_308_274_0, i_13_308_308_0,
    i_13_308_320_0, i_13_308_357_0, i_13_308_359_0, i_13_308_373_0,
    i_13_308_464_0, i_13_308_544_0, i_13_308_589_0, i_13_308_601_0,
    i_13_308_695_0, i_13_308_712_0, i_13_308_758_0, i_13_308_839_0,
    i_13_308_890_0, i_13_308_949_0, i_13_308_1100_0, i_13_308_1190_0,
    i_13_308_1207_0, i_13_308_1208_0, i_13_308_1271_0, i_13_308_1306_0,
    i_13_308_1307_0, i_13_308_1319_0, i_13_308_1345_0, i_13_308_1346_0,
    i_13_308_1436_0, i_13_308_1486_0, i_13_308_1504_0, i_13_308_1505_0,
    i_13_308_1594_0, i_13_308_1595_0, i_13_308_1639_0, i_13_308_1640_0,
    i_13_308_1688_0, i_13_308_1768_0, i_13_308_1792_0, i_13_308_1831_0,
    i_13_308_1913_0, i_13_308_1928_0, i_13_308_1948_0, i_13_308_2003_0,
    i_13_308_2030_0, i_13_308_2053_0, i_13_308_2054_0, i_13_308_2056_0,
    i_13_308_2099_0, i_13_308_2101_0, i_13_308_2189_0, i_13_308_2281_0,
    i_13_308_2282_0, i_13_308_2345_0, i_13_308_2398_0, i_13_308_2494_0,
    i_13_308_2552_0, i_13_308_2674_0, i_13_308_2675_0, i_13_308_2720_0,
    i_13_308_2846_0, i_13_308_2854_0, i_13_308_2861_0, i_13_308_2900_0,
    i_13_308_2917_0, i_13_308_2918_0, i_13_308_2983_0, i_13_308_3062_0,
    i_13_308_3089_0, i_13_308_3136_0, i_13_308_3169_0, i_13_308_3377_0,
    i_13_308_3380_0, i_13_308_3389_0, i_13_308_3479_0, i_13_308_3595_0,
    i_13_308_3596_0, i_13_308_3631_0, i_13_308_3730_0, i_13_308_3781_0,
    i_13_308_3916_0, i_13_308_3935_0, i_13_308_3979_0, i_13_308_3989_0,
    i_13_308_4034_0, i_13_308_4052_0, i_13_308_4097_0, i_13_308_4127_0,
    i_13_308_4204_0, i_13_308_4262_0, i_13_308_4394_0, i_13_308_4447_0,
    i_13_308_4555_0, i_13_308_4586_0, i_13_308_4591_0, i_13_308_4592_0,
    o_13_308_0_0  );
  input  i_13_308_64_0, i_13_308_65_0, i_13_308_118_0, i_13_308_188_0,
    i_13_308_190_0, i_13_308_226_0, i_13_308_274_0, i_13_308_308_0,
    i_13_308_320_0, i_13_308_357_0, i_13_308_359_0, i_13_308_373_0,
    i_13_308_464_0, i_13_308_544_0, i_13_308_589_0, i_13_308_601_0,
    i_13_308_695_0, i_13_308_712_0, i_13_308_758_0, i_13_308_839_0,
    i_13_308_890_0, i_13_308_949_0, i_13_308_1100_0, i_13_308_1190_0,
    i_13_308_1207_0, i_13_308_1208_0, i_13_308_1271_0, i_13_308_1306_0,
    i_13_308_1307_0, i_13_308_1319_0, i_13_308_1345_0, i_13_308_1346_0,
    i_13_308_1436_0, i_13_308_1486_0, i_13_308_1504_0, i_13_308_1505_0,
    i_13_308_1594_0, i_13_308_1595_0, i_13_308_1639_0, i_13_308_1640_0,
    i_13_308_1688_0, i_13_308_1768_0, i_13_308_1792_0, i_13_308_1831_0,
    i_13_308_1913_0, i_13_308_1928_0, i_13_308_1948_0, i_13_308_2003_0,
    i_13_308_2030_0, i_13_308_2053_0, i_13_308_2054_0, i_13_308_2056_0,
    i_13_308_2099_0, i_13_308_2101_0, i_13_308_2189_0, i_13_308_2281_0,
    i_13_308_2282_0, i_13_308_2345_0, i_13_308_2398_0, i_13_308_2494_0,
    i_13_308_2552_0, i_13_308_2674_0, i_13_308_2675_0, i_13_308_2720_0,
    i_13_308_2846_0, i_13_308_2854_0, i_13_308_2861_0, i_13_308_2900_0,
    i_13_308_2917_0, i_13_308_2918_0, i_13_308_2983_0, i_13_308_3062_0,
    i_13_308_3089_0, i_13_308_3136_0, i_13_308_3169_0, i_13_308_3377_0,
    i_13_308_3380_0, i_13_308_3389_0, i_13_308_3479_0, i_13_308_3595_0,
    i_13_308_3596_0, i_13_308_3631_0, i_13_308_3730_0, i_13_308_3781_0,
    i_13_308_3916_0, i_13_308_3935_0, i_13_308_3979_0, i_13_308_3989_0,
    i_13_308_4034_0, i_13_308_4052_0, i_13_308_4097_0, i_13_308_4127_0,
    i_13_308_4204_0, i_13_308_4262_0, i_13_308_4394_0, i_13_308_4447_0,
    i_13_308_4555_0, i_13_308_4586_0, i_13_308_4591_0, i_13_308_4592_0;
  output o_13_308_0_0;
  assign o_13_308_0_0 = ~((~i_13_308_1307_0 & (~i_13_308_2054_0 | ~i_13_308_3389_0)) | ~i_13_308_2674_0 | (~i_13_308_1208_0 & ~i_13_308_1319_0 & ~i_13_308_3916_0));
endmodule



// Benchmark "kernel_13_309" written by ABC on Sun Jul 19 10:49:41 2020

module kernel_13_309 ( 
    i_13_309_72_0, i_13_309_121_0, i_13_309_156_0, i_13_309_175_0,
    i_13_309_192_0, i_13_309_207_0, i_13_309_244_0, i_13_309_264_0,
    i_13_309_265_0, i_13_309_336_0, i_13_309_354_0, i_13_309_367_0,
    i_13_309_372_0, i_13_309_381_0, i_13_309_462_0, i_13_309_463_0,
    i_13_309_516_0, i_13_309_588_0, i_13_309_607_0, i_13_309_660_0,
    i_13_309_670_0, i_13_309_768_0, i_13_309_811_0, i_13_309_813_0,
    i_13_309_831_0, i_13_309_1072_0, i_13_309_1116_0, i_13_309_1200_0,
    i_13_309_1203_0, i_13_309_1227_0, i_13_309_1228_0, i_13_309_1252_0,
    i_13_309_1306_0, i_13_309_1344_0, i_13_309_1345_0, i_13_309_1407_0,
    i_13_309_1488_0, i_13_309_1593_0, i_13_309_1602_0, i_13_309_1633_0,
    i_13_309_1723_0, i_13_309_1813_0, i_13_309_1839_0, i_13_309_1840_0,
    i_13_309_1845_0, i_13_309_1846_0, i_13_309_1996_0, i_13_309_2029_0,
    i_13_309_2055_0, i_13_309_2124_0, i_13_309_2133_0, i_13_309_2136_0,
    i_13_309_2142_0, i_13_309_2190_0, i_13_309_2199_0, i_13_309_2200_0,
    i_13_309_2208_0, i_13_309_2280_0, i_13_309_2281_0, i_13_309_2395_0,
    i_13_309_2469_0, i_13_309_2506_0, i_13_309_2538_0, i_13_309_2613_0,
    i_13_309_2820_0, i_13_309_2934_0, i_13_309_3136_0, i_13_309_3241_0,
    i_13_309_3342_0, i_13_309_3343_0, i_13_309_3370_0, i_13_309_3387_0,
    i_13_309_3486_0, i_13_309_3502_0, i_13_309_3532_0, i_13_309_3549_0,
    i_13_309_3550_0, i_13_309_3567_0, i_13_309_3594_0, i_13_309_3595_0,
    i_13_309_3618_0, i_13_309_3619_0, i_13_309_3630_0, i_13_309_3663_0,
    i_13_309_3666_0, i_13_309_3667_0, i_13_309_3670_0, i_13_309_3691_0,
    i_13_309_3934_0, i_13_309_3988_0, i_13_309_4059_0, i_13_309_4060_0,
    i_13_309_4162_0, i_13_309_4233_0, i_13_309_4311_0, i_13_309_4312_0,
    i_13_309_4408_0, i_13_309_4449_0, i_13_309_4545_0, i_13_309_4599_0,
    o_13_309_0_0  );
  input  i_13_309_72_0, i_13_309_121_0, i_13_309_156_0, i_13_309_175_0,
    i_13_309_192_0, i_13_309_207_0, i_13_309_244_0, i_13_309_264_0,
    i_13_309_265_0, i_13_309_336_0, i_13_309_354_0, i_13_309_367_0,
    i_13_309_372_0, i_13_309_381_0, i_13_309_462_0, i_13_309_463_0,
    i_13_309_516_0, i_13_309_588_0, i_13_309_607_0, i_13_309_660_0,
    i_13_309_670_0, i_13_309_768_0, i_13_309_811_0, i_13_309_813_0,
    i_13_309_831_0, i_13_309_1072_0, i_13_309_1116_0, i_13_309_1200_0,
    i_13_309_1203_0, i_13_309_1227_0, i_13_309_1228_0, i_13_309_1252_0,
    i_13_309_1306_0, i_13_309_1344_0, i_13_309_1345_0, i_13_309_1407_0,
    i_13_309_1488_0, i_13_309_1593_0, i_13_309_1602_0, i_13_309_1633_0,
    i_13_309_1723_0, i_13_309_1813_0, i_13_309_1839_0, i_13_309_1840_0,
    i_13_309_1845_0, i_13_309_1846_0, i_13_309_1996_0, i_13_309_2029_0,
    i_13_309_2055_0, i_13_309_2124_0, i_13_309_2133_0, i_13_309_2136_0,
    i_13_309_2142_0, i_13_309_2190_0, i_13_309_2199_0, i_13_309_2200_0,
    i_13_309_2208_0, i_13_309_2280_0, i_13_309_2281_0, i_13_309_2395_0,
    i_13_309_2469_0, i_13_309_2506_0, i_13_309_2538_0, i_13_309_2613_0,
    i_13_309_2820_0, i_13_309_2934_0, i_13_309_3136_0, i_13_309_3241_0,
    i_13_309_3342_0, i_13_309_3343_0, i_13_309_3370_0, i_13_309_3387_0,
    i_13_309_3486_0, i_13_309_3502_0, i_13_309_3532_0, i_13_309_3549_0,
    i_13_309_3550_0, i_13_309_3567_0, i_13_309_3594_0, i_13_309_3595_0,
    i_13_309_3618_0, i_13_309_3619_0, i_13_309_3630_0, i_13_309_3663_0,
    i_13_309_3666_0, i_13_309_3667_0, i_13_309_3670_0, i_13_309_3691_0,
    i_13_309_3934_0, i_13_309_3988_0, i_13_309_4059_0, i_13_309_4060_0,
    i_13_309_4162_0, i_13_309_4233_0, i_13_309_4311_0, i_13_309_4312_0,
    i_13_309_4408_0, i_13_309_4449_0, i_13_309_4545_0, i_13_309_4599_0;
  output o_13_309_0_0;
  assign o_13_309_0_0 = ~(~i_13_309_2281_0 | ~i_13_309_462_0 | i_13_309_2208_0);
endmodule



// Benchmark "kernel_13_310" written by ABC on Sun Jul 19 10:49:42 2020

module kernel_13_310 ( 
    i_13_310_71_0, i_13_310_79_0, i_13_310_125_0, i_13_310_139_0,
    i_13_310_172_0, i_13_310_175_0, i_13_310_179_0, i_13_310_205_0,
    i_13_310_279_0, i_13_310_285_0, i_13_310_310_0, i_13_310_313_0,
    i_13_310_358_0, i_13_310_373_0, i_13_310_448_0, i_13_310_522_0,
    i_13_310_538_0, i_13_310_604_0, i_13_310_607_0, i_13_310_646_0,
    i_13_310_657_0, i_13_310_672_0, i_13_310_682_0, i_13_310_683_0,
    i_13_310_685_0, i_13_310_688_0, i_13_310_691_0, i_13_310_820_0,
    i_13_310_844_0, i_13_310_1123_0, i_13_310_1124_0, i_13_310_1215_0,
    i_13_310_1224_0, i_13_310_1275_0, i_13_310_1276_0, i_13_310_1277_0,
    i_13_310_1286_0, i_13_310_1305_0, i_13_310_1311_0, i_13_310_1501_0,
    i_13_310_1511_0, i_13_310_1599_0, i_13_310_1645_0, i_13_310_1672_0,
    i_13_310_1732_0, i_13_310_1771_0, i_13_310_1799_0, i_13_310_1881_0,
    i_13_310_1886_0, i_13_310_1934_0, i_13_310_2175_0, i_13_310_2481_0,
    i_13_310_2646_0, i_13_310_2650_0, i_13_310_2677_0, i_13_310_2680_0,
    i_13_310_2698_0, i_13_310_2851_0, i_13_310_2878_0, i_13_310_2916_0,
    i_13_310_2938_0, i_13_310_3014_0, i_13_310_3204_0, i_13_310_3217_0,
    i_13_310_3235_0, i_13_310_3270_0, i_13_310_3271_0, i_13_310_3275_0,
    i_13_310_3356_0, i_13_310_3392_0, i_13_310_3418_0, i_13_310_3421_0,
    i_13_310_3574_0, i_13_310_3652_0, i_13_310_3742_0, i_13_310_3761_0,
    i_13_310_3895_0, i_13_310_3994_0, i_13_310_4083_0, i_13_310_4084_0,
    i_13_310_4186_0, i_13_310_4248_0, i_13_310_4251_0, i_13_310_4252_0,
    i_13_310_4260_0, i_13_310_4293_0, i_13_310_4296_0, i_13_310_4306_0,
    i_13_310_4307_0, i_13_310_4309_0, i_13_310_4400_0, i_13_310_4435_0,
    i_13_310_4446_0, i_13_310_4447_0, i_13_310_4557_0, i_13_310_4590_0,
    i_13_310_4593_0, i_13_310_4594_0, i_13_310_4597_0, i_13_310_4598_0,
    o_13_310_0_0  );
  input  i_13_310_71_0, i_13_310_79_0, i_13_310_125_0, i_13_310_139_0,
    i_13_310_172_0, i_13_310_175_0, i_13_310_179_0, i_13_310_205_0,
    i_13_310_279_0, i_13_310_285_0, i_13_310_310_0, i_13_310_313_0,
    i_13_310_358_0, i_13_310_373_0, i_13_310_448_0, i_13_310_522_0,
    i_13_310_538_0, i_13_310_604_0, i_13_310_607_0, i_13_310_646_0,
    i_13_310_657_0, i_13_310_672_0, i_13_310_682_0, i_13_310_683_0,
    i_13_310_685_0, i_13_310_688_0, i_13_310_691_0, i_13_310_820_0,
    i_13_310_844_0, i_13_310_1123_0, i_13_310_1124_0, i_13_310_1215_0,
    i_13_310_1224_0, i_13_310_1275_0, i_13_310_1276_0, i_13_310_1277_0,
    i_13_310_1286_0, i_13_310_1305_0, i_13_310_1311_0, i_13_310_1501_0,
    i_13_310_1511_0, i_13_310_1599_0, i_13_310_1645_0, i_13_310_1672_0,
    i_13_310_1732_0, i_13_310_1771_0, i_13_310_1799_0, i_13_310_1881_0,
    i_13_310_1886_0, i_13_310_1934_0, i_13_310_2175_0, i_13_310_2481_0,
    i_13_310_2646_0, i_13_310_2650_0, i_13_310_2677_0, i_13_310_2680_0,
    i_13_310_2698_0, i_13_310_2851_0, i_13_310_2878_0, i_13_310_2916_0,
    i_13_310_2938_0, i_13_310_3014_0, i_13_310_3204_0, i_13_310_3217_0,
    i_13_310_3235_0, i_13_310_3270_0, i_13_310_3271_0, i_13_310_3275_0,
    i_13_310_3356_0, i_13_310_3392_0, i_13_310_3418_0, i_13_310_3421_0,
    i_13_310_3574_0, i_13_310_3652_0, i_13_310_3742_0, i_13_310_3761_0,
    i_13_310_3895_0, i_13_310_3994_0, i_13_310_4083_0, i_13_310_4084_0,
    i_13_310_4186_0, i_13_310_4248_0, i_13_310_4251_0, i_13_310_4252_0,
    i_13_310_4260_0, i_13_310_4293_0, i_13_310_4296_0, i_13_310_4306_0,
    i_13_310_4307_0, i_13_310_4309_0, i_13_310_4400_0, i_13_310_4435_0,
    i_13_310_4446_0, i_13_310_4447_0, i_13_310_4557_0, i_13_310_4590_0,
    i_13_310_4593_0, i_13_310_4594_0, i_13_310_4597_0, i_13_310_4598_0;
  output o_13_310_0_0;
  assign o_13_310_0_0 = ~((~i_13_310_4083_0 & (~i_13_310_1123_0 | (~i_13_310_1277_0 & i_13_310_4309_0))) | (~i_13_310_1276_0 & ~i_13_310_3014_0 & ~i_13_310_4260_0) | (~i_13_310_313_0 & ~i_13_310_4435_0));
endmodule



// Benchmark "kernel_13_311" written by ABC on Sun Jul 19 10:49:42 2020

module kernel_13_311 ( 
    i_13_311_75_0, i_13_311_76_0, i_13_311_79_0, i_13_311_94_0,
    i_13_311_95_0, i_13_311_122_0, i_13_311_143_0, i_13_311_166_0,
    i_13_311_193_0, i_13_311_322_0, i_13_311_406_0, i_13_311_518_0,
    i_13_311_586_0, i_13_311_698_0, i_13_311_700_0, i_13_311_701_0,
    i_13_311_827_0, i_13_311_841_0, i_13_311_932_0, i_13_311_943_0,
    i_13_311_979_0, i_13_311_1025_0, i_13_311_1078_0, i_13_311_1079_0,
    i_13_311_1084_0, i_13_311_1115_0, i_13_311_1209_0, i_13_311_1276_0,
    i_13_311_1330_0, i_13_311_1408_0, i_13_311_1429_0, i_13_311_1430_0,
    i_13_311_1439_0, i_13_311_1546_0, i_13_311_1596_0, i_13_311_1610_0,
    i_13_311_1632_0, i_13_311_1636_0, i_13_311_1675_0, i_13_311_1777_0,
    i_13_311_1778_0, i_13_311_1831_0, i_13_311_1888_0, i_13_311_1908_0,
    i_13_311_1947_0, i_13_311_2028_0, i_13_311_2119_0, i_13_311_2343_0,
    i_13_311_2450_0, i_13_311_2455_0, i_13_311_2610_0, i_13_311_2618_0,
    i_13_311_2709_0, i_13_311_2788_0, i_13_311_2858_0, i_13_311_2880_0,
    i_13_311_2887_0, i_13_311_2888_0, i_13_311_2919_0, i_13_311_2955_0,
    i_13_311_2959_0, i_13_311_2983_0, i_13_311_3141_0, i_13_311_3208_0,
    i_13_311_3211_0, i_13_311_3244_0, i_13_311_3437_0, i_13_311_3448_0,
    i_13_311_3451_0, i_13_311_3454_0, i_13_311_3455_0, i_13_311_3464_0,
    i_13_311_3482_0, i_13_311_3486_0, i_13_311_3526_0, i_13_311_3528_0,
    i_13_311_3532_0, i_13_311_3571_0, i_13_311_3572_0, i_13_311_3576_0,
    i_13_311_3618_0, i_13_311_3640_0, i_13_311_3649_0, i_13_311_3688_0,
    i_13_311_3767_0, i_13_311_3783_0, i_13_311_3799_0, i_13_311_3837_0,
    i_13_311_3846_0, i_13_311_3888_0, i_13_311_3967_0, i_13_311_4009_0,
    i_13_311_4086_0, i_13_311_4170_0, i_13_311_4190_0, i_13_311_4248_0,
    i_13_311_4252_0, i_13_311_4265_0, i_13_311_4301_0, i_13_311_4451_0,
    o_13_311_0_0  );
  input  i_13_311_75_0, i_13_311_76_0, i_13_311_79_0, i_13_311_94_0,
    i_13_311_95_0, i_13_311_122_0, i_13_311_143_0, i_13_311_166_0,
    i_13_311_193_0, i_13_311_322_0, i_13_311_406_0, i_13_311_518_0,
    i_13_311_586_0, i_13_311_698_0, i_13_311_700_0, i_13_311_701_0,
    i_13_311_827_0, i_13_311_841_0, i_13_311_932_0, i_13_311_943_0,
    i_13_311_979_0, i_13_311_1025_0, i_13_311_1078_0, i_13_311_1079_0,
    i_13_311_1084_0, i_13_311_1115_0, i_13_311_1209_0, i_13_311_1276_0,
    i_13_311_1330_0, i_13_311_1408_0, i_13_311_1429_0, i_13_311_1430_0,
    i_13_311_1439_0, i_13_311_1546_0, i_13_311_1596_0, i_13_311_1610_0,
    i_13_311_1632_0, i_13_311_1636_0, i_13_311_1675_0, i_13_311_1777_0,
    i_13_311_1778_0, i_13_311_1831_0, i_13_311_1888_0, i_13_311_1908_0,
    i_13_311_1947_0, i_13_311_2028_0, i_13_311_2119_0, i_13_311_2343_0,
    i_13_311_2450_0, i_13_311_2455_0, i_13_311_2610_0, i_13_311_2618_0,
    i_13_311_2709_0, i_13_311_2788_0, i_13_311_2858_0, i_13_311_2880_0,
    i_13_311_2887_0, i_13_311_2888_0, i_13_311_2919_0, i_13_311_2955_0,
    i_13_311_2959_0, i_13_311_2983_0, i_13_311_3141_0, i_13_311_3208_0,
    i_13_311_3211_0, i_13_311_3244_0, i_13_311_3437_0, i_13_311_3448_0,
    i_13_311_3451_0, i_13_311_3454_0, i_13_311_3455_0, i_13_311_3464_0,
    i_13_311_3482_0, i_13_311_3486_0, i_13_311_3526_0, i_13_311_3528_0,
    i_13_311_3532_0, i_13_311_3571_0, i_13_311_3572_0, i_13_311_3576_0,
    i_13_311_3618_0, i_13_311_3640_0, i_13_311_3649_0, i_13_311_3688_0,
    i_13_311_3767_0, i_13_311_3783_0, i_13_311_3799_0, i_13_311_3837_0,
    i_13_311_3846_0, i_13_311_3888_0, i_13_311_3967_0, i_13_311_4009_0,
    i_13_311_4086_0, i_13_311_4170_0, i_13_311_4190_0, i_13_311_4248_0,
    i_13_311_4252_0, i_13_311_4265_0, i_13_311_4301_0, i_13_311_4451_0;
  output o_13_311_0_0;
  assign o_13_311_0_0 = ~((i_13_311_2983_0 & ((~i_13_311_943_0 & i_13_311_3783_0) | (~i_13_311_1276_0 & ~i_13_311_4451_0))) | (~i_13_311_3572_0 & ((~i_13_311_701_0 & ~i_13_311_3576_0 & ~i_13_311_3649_0) | (~i_13_311_2888_0 & ~i_13_311_3688_0))) | (i_13_311_94_0 & i_13_311_193_0 & ~i_13_311_3464_0) | (~i_13_311_2788_0 & i_13_311_3688_0) | i_13_311_3846_0 | (i_13_311_3783_0 & ~i_13_311_4252_0));
endmodule



// Benchmark "kernel_13_312" written by ABC on Sun Jul 19 10:49:43 2020

module kernel_13_312 ( 
    i_13_312_25_0, i_13_312_30_0, i_13_312_48_0, i_13_312_69_0,
    i_13_312_70_0, i_13_312_177_0, i_13_312_186_0, i_13_312_193_0,
    i_13_312_321_0, i_13_312_381_0, i_13_312_411_0, i_13_312_417_0,
    i_13_312_492_0, i_13_312_498_0, i_13_312_570_0, i_13_312_609_0,
    i_13_312_645_0, i_13_312_678_0, i_13_312_699_0, i_13_312_759_0,
    i_13_312_760_0, i_13_312_762_0, i_13_312_763_0, i_13_312_870_0,
    i_13_312_933_0, i_13_312_994_0, i_13_312_1021_0, i_13_312_1083_0,
    i_13_312_1084_0, i_13_312_1086_0, i_13_312_1095_0, i_13_312_1104_0,
    i_13_312_1131_0, i_13_312_1132_0, i_13_312_1224_0, i_13_312_1302_0,
    i_13_312_1303_0, i_13_312_1308_0, i_13_312_1347_0, i_13_312_1407_0,
    i_13_312_1525_0, i_13_312_1528_0, i_13_312_1551_0, i_13_312_1605_0,
    i_13_312_1632_0, i_13_312_1644_0, i_13_312_1714_0, i_13_312_1716_0,
    i_13_312_1789_0, i_13_312_1797_0, i_13_312_1798_0, i_13_312_1806_0,
    i_13_312_1807_0, i_13_312_1843_0, i_13_312_1942_0, i_13_312_1992_0,
    i_13_312_1995_0, i_13_312_2023_0, i_13_312_2055_0, i_13_312_2122_0,
    i_13_312_2224_0, i_13_312_2472_0, i_13_312_2473_0, i_13_312_2505_0,
    i_13_312_2536_0, i_13_312_2541_0, i_13_312_2542_0, i_13_312_2722_0,
    i_13_312_2757_0, i_13_312_2955_0, i_13_312_3022_0, i_13_312_3030_0,
    i_13_312_3031_0, i_13_312_3118_0, i_13_312_3121_0, i_13_312_3198_0,
    i_13_312_3264_0, i_13_312_3346_0, i_13_312_3375_0, i_13_312_3399_0,
    i_13_312_3453_0, i_13_312_3702_0, i_13_312_3739_0, i_13_312_3804_0,
    i_13_312_3822_0, i_13_312_4038_0, i_13_312_4081_0, i_13_312_4090_0,
    i_13_312_4093_0, i_13_312_4117_0, i_13_312_4189_0, i_13_312_4233_0,
    i_13_312_4255_0, i_13_312_4272_0, i_13_312_4273_0, i_13_312_4308_0,
    i_13_312_4336_0, i_13_312_4596_0, i_13_312_4605_0, i_13_312_4606_0,
    o_13_312_0_0  );
  input  i_13_312_25_0, i_13_312_30_0, i_13_312_48_0, i_13_312_69_0,
    i_13_312_70_0, i_13_312_177_0, i_13_312_186_0, i_13_312_193_0,
    i_13_312_321_0, i_13_312_381_0, i_13_312_411_0, i_13_312_417_0,
    i_13_312_492_0, i_13_312_498_0, i_13_312_570_0, i_13_312_609_0,
    i_13_312_645_0, i_13_312_678_0, i_13_312_699_0, i_13_312_759_0,
    i_13_312_760_0, i_13_312_762_0, i_13_312_763_0, i_13_312_870_0,
    i_13_312_933_0, i_13_312_994_0, i_13_312_1021_0, i_13_312_1083_0,
    i_13_312_1084_0, i_13_312_1086_0, i_13_312_1095_0, i_13_312_1104_0,
    i_13_312_1131_0, i_13_312_1132_0, i_13_312_1224_0, i_13_312_1302_0,
    i_13_312_1303_0, i_13_312_1308_0, i_13_312_1347_0, i_13_312_1407_0,
    i_13_312_1525_0, i_13_312_1528_0, i_13_312_1551_0, i_13_312_1605_0,
    i_13_312_1632_0, i_13_312_1644_0, i_13_312_1714_0, i_13_312_1716_0,
    i_13_312_1789_0, i_13_312_1797_0, i_13_312_1798_0, i_13_312_1806_0,
    i_13_312_1807_0, i_13_312_1843_0, i_13_312_1942_0, i_13_312_1992_0,
    i_13_312_1995_0, i_13_312_2023_0, i_13_312_2055_0, i_13_312_2122_0,
    i_13_312_2224_0, i_13_312_2472_0, i_13_312_2473_0, i_13_312_2505_0,
    i_13_312_2536_0, i_13_312_2541_0, i_13_312_2542_0, i_13_312_2722_0,
    i_13_312_2757_0, i_13_312_2955_0, i_13_312_3022_0, i_13_312_3030_0,
    i_13_312_3031_0, i_13_312_3118_0, i_13_312_3121_0, i_13_312_3198_0,
    i_13_312_3264_0, i_13_312_3346_0, i_13_312_3375_0, i_13_312_3399_0,
    i_13_312_3453_0, i_13_312_3702_0, i_13_312_3739_0, i_13_312_3804_0,
    i_13_312_3822_0, i_13_312_4038_0, i_13_312_4081_0, i_13_312_4090_0,
    i_13_312_4093_0, i_13_312_4117_0, i_13_312_4189_0, i_13_312_4233_0,
    i_13_312_4255_0, i_13_312_4272_0, i_13_312_4273_0, i_13_312_4308_0,
    i_13_312_4336_0, i_13_312_4596_0, i_13_312_4605_0, i_13_312_4606_0;
  output o_13_312_0_0;
  assign o_13_312_0_0 = ~((~i_13_312_1605_0 & i_13_312_3739_0) | (~i_13_312_763_0 & i_13_312_4081_0 & ~i_13_312_4273_0) | (~i_13_312_1302_0 & ~i_13_312_1347_0 & ~i_13_312_3822_0));
endmodule



// Benchmark "kernel_13_313" written by ABC on Sun Jul 19 10:49:44 2020

module kernel_13_313 ( 
    i_13_313_136_0, i_13_313_137_0, i_13_313_139_0, i_13_313_140_0,
    i_13_313_175_0, i_13_313_226_0, i_13_313_227_0, i_13_313_230_0,
    i_13_313_268_0, i_13_313_362_0, i_13_313_419_0, i_13_313_533_0,
    i_13_313_536_0, i_13_313_641_0, i_13_313_695_0, i_13_313_824_0,
    i_13_313_850_0, i_13_313_892_0, i_13_313_976_0, i_13_313_982_0,
    i_13_313_985_0, i_13_313_1201_0, i_13_313_1217_0, i_13_313_1219_0,
    i_13_313_1220_0, i_13_313_1274_0, i_13_313_1283_0, i_13_313_1343_0,
    i_13_313_1467_0, i_13_313_1607_0, i_13_313_1711_0, i_13_313_1712_0,
    i_13_313_1722_0, i_13_313_1723_0, i_13_313_1778_0, i_13_313_1882_0,
    i_13_313_1883_0, i_13_313_1885_0, i_13_313_1886_0, i_13_313_1958_0,
    i_13_313_2003_0, i_13_313_2098_0, i_13_313_2189_0, i_13_313_2210_0,
    i_13_313_2297_0, i_13_313_2426_0, i_13_313_2549_0, i_13_313_2647_0,
    i_13_313_2648_0, i_13_313_2708_0, i_13_313_2747_0, i_13_313_2846_0,
    i_13_313_2848_0, i_13_313_2855_0, i_13_313_2858_0, i_13_313_2872_0,
    i_13_313_2885_0, i_13_313_2909_0, i_13_313_2935_0, i_13_313_2956_0,
    i_13_313_2983_0, i_13_313_3001_0, i_13_313_3004_0, i_13_313_3005_0,
    i_13_313_3010_0, i_13_313_3037_0, i_13_313_3038_0, i_13_313_3056_0,
    i_13_313_3109_0, i_13_313_3143_0, i_13_313_3322_0, i_13_313_3370_0,
    i_13_313_3382_0, i_13_313_3385_0, i_13_313_3386_0, i_13_313_3425_0,
    i_13_313_3439_0, i_13_313_3449_0, i_13_313_3487_0, i_13_313_3503_0,
    i_13_313_3542_0, i_13_313_3743_0, i_13_313_3820_0, i_13_313_3836_0,
    i_13_313_3839_0, i_13_313_3865_0, i_13_313_4016_0, i_13_313_4054_0,
    i_13_313_4060_0, i_13_313_4063_0, i_13_313_4181_0, i_13_313_4190_0,
    i_13_313_4211_0, i_13_313_4342_0, i_13_313_4388_0, i_13_313_4394_0,
    i_13_313_4411_0, i_13_313_4414_0, i_13_313_4522_0, i_13_313_4531_0,
    o_13_313_0_0  );
  input  i_13_313_136_0, i_13_313_137_0, i_13_313_139_0, i_13_313_140_0,
    i_13_313_175_0, i_13_313_226_0, i_13_313_227_0, i_13_313_230_0,
    i_13_313_268_0, i_13_313_362_0, i_13_313_419_0, i_13_313_533_0,
    i_13_313_536_0, i_13_313_641_0, i_13_313_695_0, i_13_313_824_0,
    i_13_313_850_0, i_13_313_892_0, i_13_313_976_0, i_13_313_982_0,
    i_13_313_985_0, i_13_313_1201_0, i_13_313_1217_0, i_13_313_1219_0,
    i_13_313_1220_0, i_13_313_1274_0, i_13_313_1283_0, i_13_313_1343_0,
    i_13_313_1467_0, i_13_313_1607_0, i_13_313_1711_0, i_13_313_1712_0,
    i_13_313_1722_0, i_13_313_1723_0, i_13_313_1778_0, i_13_313_1882_0,
    i_13_313_1883_0, i_13_313_1885_0, i_13_313_1886_0, i_13_313_1958_0,
    i_13_313_2003_0, i_13_313_2098_0, i_13_313_2189_0, i_13_313_2210_0,
    i_13_313_2297_0, i_13_313_2426_0, i_13_313_2549_0, i_13_313_2647_0,
    i_13_313_2648_0, i_13_313_2708_0, i_13_313_2747_0, i_13_313_2846_0,
    i_13_313_2848_0, i_13_313_2855_0, i_13_313_2858_0, i_13_313_2872_0,
    i_13_313_2885_0, i_13_313_2909_0, i_13_313_2935_0, i_13_313_2956_0,
    i_13_313_2983_0, i_13_313_3001_0, i_13_313_3004_0, i_13_313_3005_0,
    i_13_313_3010_0, i_13_313_3037_0, i_13_313_3038_0, i_13_313_3056_0,
    i_13_313_3109_0, i_13_313_3143_0, i_13_313_3322_0, i_13_313_3370_0,
    i_13_313_3382_0, i_13_313_3385_0, i_13_313_3386_0, i_13_313_3425_0,
    i_13_313_3439_0, i_13_313_3449_0, i_13_313_3487_0, i_13_313_3503_0,
    i_13_313_3542_0, i_13_313_3743_0, i_13_313_3820_0, i_13_313_3836_0,
    i_13_313_3839_0, i_13_313_3865_0, i_13_313_4016_0, i_13_313_4054_0,
    i_13_313_4060_0, i_13_313_4063_0, i_13_313_4181_0, i_13_313_4190_0,
    i_13_313_4211_0, i_13_313_4342_0, i_13_313_4388_0, i_13_313_4394_0,
    i_13_313_4411_0, i_13_313_4414_0, i_13_313_4522_0, i_13_313_4531_0;
  output o_13_313_0_0;
  assign o_13_313_0_0 = ~((~i_13_313_1220_0 & ~i_13_313_2872_0 & (i_13_313_175_0 | i_13_313_1958_0)) | (i_13_313_3010_0 & (i_13_313_1467_0 | (~i_13_313_1343_0 & ~i_13_313_1711_0))) | (~i_13_313_1607_0 & ~i_13_313_2858_0 & ~i_13_313_2935_0 & ~i_13_313_3385_0 & ~i_13_313_3425_0) | (i_13_313_3542_0 & i_13_313_3743_0) | (~i_13_313_136_0 & ~i_13_313_1886_0 & ~i_13_313_2426_0 & ~i_13_313_4394_0));
endmodule



// Benchmark "kernel_13_314" written by ABC on Sun Jul 19 10:49:45 2020

module kernel_13_314 ( 
    i_13_314_45_0, i_13_314_99_0, i_13_314_102_0, i_13_314_157_0,
    i_13_314_192_0, i_13_314_193_0, i_13_314_195_0, i_13_314_333_0,
    i_13_314_442_0, i_13_314_450_0, i_13_314_451_0, i_13_314_577_0,
    i_13_314_612_0, i_13_314_624_0, i_13_314_640_0, i_13_314_657_0,
    i_13_314_714_0, i_13_314_721_0, i_13_314_858_0, i_13_314_946_0,
    i_13_314_948_0, i_13_314_955_0, i_13_314_982_0, i_13_314_1062_0,
    i_13_314_1116_0, i_13_314_1147_0, i_13_314_1224_0, i_13_314_1225_0,
    i_13_314_1227_0, i_13_314_1231_0, i_13_314_1282_0, i_13_314_1297_0,
    i_13_314_1314_0, i_13_314_1345_0, i_13_314_1407_0, i_13_314_1435_0,
    i_13_314_1443_0, i_13_314_1458_0, i_13_314_1468_0, i_13_314_1488_0,
    i_13_314_1494_0, i_13_314_1566_0, i_13_314_1567_0, i_13_314_1764_0,
    i_13_314_1776_0, i_13_314_1800_0, i_13_314_1801_0, i_13_314_1803_0,
    i_13_314_1891_0, i_13_314_1926_0, i_13_314_1990_0, i_13_314_1999_0,
    i_13_314_2056_0, i_13_314_2107_0, i_13_314_2137_0, i_13_314_2145_0,
    i_13_314_2205_0, i_13_314_2209_0, i_13_314_2296_0, i_13_314_2425_0,
    i_13_314_2532_0, i_13_314_2568_0, i_13_314_2613_0, i_13_314_2614_0,
    i_13_314_2691_0, i_13_314_2745_0, i_13_314_2820_0, i_13_314_3006_0,
    i_13_314_3024_0, i_13_314_3052_0, i_13_314_3055_0, i_13_314_3144_0,
    i_13_314_3214_0, i_13_314_3267_0, i_13_314_3286_0, i_13_314_3339_0,
    i_13_314_3342_0, i_13_314_3420_0, i_13_314_3421_0, i_13_314_3474_0,
    i_13_314_3486_0, i_13_314_3753_0, i_13_314_3873_0, i_13_314_3978_0,
    i_13_314_4017_0, i_13_314_4086_0, i_13_314_4087_0, i_13_314_4230_0,
    i_13_314_4231_0, i_13_314_4233_0, i_13_314_4266_0, i_13_314_4267_0,
    i_13_314_4302_0, i_13_314_4339_0, i_13_314_4341_0, i_13_314_4404_0,
    i_13_314_4431_0, i_13_314_4468_0, i_13_314_4509_0, i_13_314_4513_0,
    o_13_314_0_0  );
  input  i_13_314_45_0, i_13_314_99_0, i_13_314_102_0, i_13_314_157_0,
    i_13_314_192_0, i_13_314_193_0, i_13_314_195_0, i_13_314_333_0,
    i_13_314_442_0, i_13_314_450_0, i_13_314_451_0, i_13_314_577_0,
    i_13_314_612_0, i_13_314_624_0, i_13_314_640_0, i_13_314_657_0,
    i_13_314_714_0, i_13_314_721_0, i_13_314_858_0, i_13_314_946_0,
    i_13_314_948_0, i_13_314_955_0, i_13_314_982_0, i_13_314_1062_0,
    i_13_314_1116_0, i_13_314_1147_0, i_13_314_1224_0, i_13_314_1225_0,
    i_13_314_1227_0, i_13_314_1231_0, i_13_314_1282_0, i_13_314_1297_0,
    i_13_314_1314_0, i_13_314_1345_0, i_13_314_1407_0, i_13_314_1435_0,
    i_13_314_1443_0, i_13_314_1458_0, i_13_314_1468_0, i_13_314_1488_0,
    i_13_314_1494_0, i_13_314_1566_0, i_13_314_1567_0, i_13_314_1764_0,
    i_13_314_1776_0, i_13_314_1800_0, i_13_314_1801_0, i_13_314_1803_0,
    i_13_314_1891_0, i_13_314_1926_0, i_13_314_1990_0, i_13_314_1999_0,
    i_13_314_2056_0, i_13_314_2107_0, i_13_314_2137_0, i_13_314_2145_0,
    i_13_314_2205_0, i_13_314_2209_0, i_13_314_2296_0, i_13_314_2425_0,
    i_13_314_2532_0, i_13_314_2568_0, i_13_314_2613_0, i_13_314_2614_0,
    i_13_314_2691_0, i_13_314_2745_0, i_13_314_2820_0, i_13_314_3006_0,
    i_13_314_3024_0, i_13_314_3052_0, i_13_314_3055_0, i_13_314_3144_0,
    i_13_314_3214_0, i_13_314_3267_0, i_13_314_3286_0, i_13_314_3339_0,
    i_13_314_3342_0, i_13_314_3420_0, i_13_314_3421_0, i_13_314_3474_0,
    i_13_314_3486_0, i_13_314_3753_0, i_13_314_3873_0, i_13_314_3978_0,
    i_13_314_4017_0, i_13_314_4086_0, i_13_314_4087_0, i_13_314_4230_0,
    i_13_314_4231_0, i_13_314_4233_0, i_13_314_4266_0, i_13_314_4267_0,
    i_13_314_4302_0, i_13_314_4339_0, i_13_314_4341_0, i_13_314_4404_0,
    i_13_314_4431_0, i_13_314_4468_0, i_13_314_4509_0, i_13_314_4513_0;
  output o_13_314_0_0;
  assign o_13_314_0_0 = ~((~i_13_314_3339_0 & ~i_13_314_4302_0) | (~i_13_314_192_0 & ~i_13_314_1566_0));
endmodule



// Benchmark "kernel_13_315" written by ABC on Sun Jul 19 10:49:46 2020

module kernel_13_315 ( 
    i_13_315_26_0, i_13_315_69_0, i_13_315_93_0, i_13_315_96_0,
    i_13_315_97_0, i_13_315_106_0, i_13_315_107_0, i_13_315_117_0,
    i_13_315_121_0, i_13_315_159_0, i_13_315_180_0, i_13_315_183_0,
    i_13_315_352_0, i_13_315_386_0, i_13_315_409_0, i_13_315_410_0,
    i_13_315_415_0, i_13_315_457_0, i_13_315_529_0, i_13_315_565_0,
    i_13_315_654_0, i_13_315_697_0, i_13_315_746_0, i_13_315_760_0,
    i_13_315_800_0, i_13_315_832_0, i_13_315_933_0, i_13_315_944_0,
    i_13_315_1086_0, i_13_315_1087_0, i_13_315_1088_0, i_13_315_1097_0,
    i_13_315_1303_0, i_13_315_1491_0, i_13_315_1507_0, i_13_315_1529_0,
    i_13_315_1725_0, i_13_315_1789_0, i_13_315_1790_0, i_13_315_1797_0,
    i_13_315_1807_0, i_13_315_1815_0, i_13_315_1995_0, i_13_315_1996_0,
    i_13_315_2122_0, i_13_315_2177_0, i_13_315_2211_0, i_13_315_2212_0,
    i_13_315_2239_0, i_13_315_2240_0, i_13_315_2303_0, i_13_315_2429_0,
    i_13_315_2614_0, i_13_315_2713_0, i_13_315_2716_0, i_13_315_2760_0,
    i_13_315_2848_0, i_13_315_2942_0, i_13_315_3022_0, i_13_315_3030_0,
    i_13_315_3066_0, i_13_315_3103_0, i_13_315_3147_0, i_13_315_3153_0,
    i_13_315_3237_0, i_13_315_3326_0, i_13_315_3345_0, i_13_315_3391_0,
    i_13_315_3399_0, i_13_315_3400_0, i_13_315_3525_0, i_13_315_3527_0,
    i_13_315_3580_0, i_13_315_3607_0, i_13_315_3686_0, i_13_315_3702_0,
    i_13_315_3739_0, i_13_315_3797_0, i_13_315_3846_0, i_13_315_3985_0,
    i_13_315_3986_0, i_13_315_4006_0, i_13_315_4008_0, i_13_315_4009_0,
    i_13_315_4046_0, i_13_315_4047_0, i_13_315_4094_0, i_13_315_4193_0,
    i_13_315_4235_0, i_13_315_4238_0, i_13_315_4261_0, i_13_315_4264_0,
    i_13_315_4273_0, i_13_315_4310_0, i_13_315_4327_0, i_13_315_4343_0,
    i_13_315_4399_0, i_13_315_4416_0, i_13_315_4417_0, i_13_315_4463_0,
    o_13_315_0_0  );
  input  i_13_315_26_0, i_13_315_69_0, i_13_315_93_0, i_13_315_96_0,
    i_13_315_97_0, i_13_315_106_0, i_13_315_107_0, i_13_315_117_0,
    i_13_315_121_0, i_13_315_159_0, i_13_315_180_0, i_13_315_183_0,
    i_13_315_352_0, i_13_315_386_0, i_13_315_409_0, i_13_315_410_0,
    i_13_315_415_0, i_13_315_457_0, i_13_315_529_0, i_13_315_565_0,
    i_13_315_654_0, i_13_315_697_0, i_13_315_746_0, i_13_315_760_0,
    i_13_315_800_0, i_13_315_832_0, i_13_315_933_0, i_13_315_944_0,
    i_13_315_1086_0, i_13_315_1087_0, i_13_315_1088_0, i_13_315_1097_0,
    i_13_315_1303_0, i_13_315_1491_0, i_13_315_1507_0, i_13_315_1529_0,
    i_13_315_1725_0, i_13_315_1789_0, i_13_315_1790_0, i_13_315_1797_0,
    i_13_315_1807_0, i_13_315_1815_0, i_13_315_1995_0, i_13_315_1996_0,
    i_13_315_2122_0, i_13_315_2177_0, i_13_315_2211_0, i_13_315_2212_0,
    i_13_315_2239_0, i_13_315_2240_0, i_13_315_2303_0, i_13_315_2429_0,
    i_13_315_2614_0, i_13_315_2713_0, i_13_315_2716_0, i_13_315_2760_0,
    i_13_315_2848_0, i_13_315_2942_0, i_13_315_3022_0, i_13_315_3030_0,
    i_13_315_3066_0, i_13_315_3103_0, i_13_315_3147_0, i_13_315_3153_0,
    i_13_315_3237_0, i_13_315_3326_0, i_13_315_3345_0, i_13_315_3391_0,
    i_13_315_3399_0, i_13_315_3400_0, i_13_315_3525_0, i_13_315_3527_0,
    i_13_315_3580_0, i_13_315_3607_0, i_13_315_3686_0, i_13_315_3702_0,
    i_13_315_3739_0, i_13_315_3797_0, i_13_315_3846_0, i_13_315_3985_0,
    i_13_315_3986_0, i_13_315_4006_0, i_13_315_4008_0, i_13_315_4009_0,
    i_13_315_4046_0, i_13_315_4047_0, i_13_315_4094_0, i_13_315_4193_0,
    i_13_315_4235_0, i_13_315_4238_0, i_13_315_4261_0, i_13_315_4264_0,
    i_13_315_4273_0, i_13_315_4310_0, i_13_315_4327_0, i_13_315_4343_0,
    i_13_315_4399_0, i_13_315_4416_0, i_13_315_4417_0, i_13_315_4463_0;
  output o_13_315_0_0;
  assign o_13_315_0_0 = ~((~i_13_315_3345_0 & ((~i_13_315_386_0 & ~i_13_315_1996_0) | (~i_13_315_3400_0 & i_13_315_3739_0))) | (i_13_315_2848_0 & ~i_13_315_3391_0 & ~i_13_315_3400_0 & ~i_13_315_3739_0) | (~i_13_315_1995_0 & ~i_13_315_2716_0 & ~i_13_315_4047_0 & ~i_13_315_4310_0 & ~i_13_315_4327_0) | (~i_13_315_97_0 & ~i_13_315_933_0 & ~i_13_315_2429_0 & ~i_13_315_4416_0) | (i_13_315_4235_0 & ~i_13_315_4417_0));
endmodule



// Benchmark "kernel_13_316" written by ABC on Sun Jul 19 10:49:47 2020

module kernel_13_316 ( 
    i_13_316_40_0, i_13_316_58_0, i_13_316_259_0, i_13_316_276_0,
    i_13_316_369_0, i_13_316_450_0, i_13_316_513_0, i_13_316_526_0,
    i_13_316_552_0, i_13_316_604_0, i_13_316_606_0, i_13_316_607_0,
    i_13_316_610_0, i_13_316_657_0, i_13_316_658_0, i_13_316_660_0,
    i_13_316_661_0, i_13_316_663_0, i_13_316_670_0, i_13_316_678_0,
    i_13_316_829_0, i_13_316_840_0, i_13_316_931_0, i_13_316_936_0,
    i_13_316_939_0, i_13_316_1056_0, i_13_316_1059_0, i_13_316_1060_0,
    i_13_316_1072_0, i_13_316_1102_0, i_13_316_1119_0, i_13_316_1147_0,
    i_13_316_1516_0, i_13_316_1534_0, i_13_316_1606_0, i_13_316_1659_0,
    i_13_316_1660_0, i_13_316_1663_0, i_13_316_1729_0, i_13_316_1731_0,
    i_13_316_1732_0, i_13_316_1764_0, i_13_316_1767_0, i_13_316_1891_0,
    i_13_316_1897_0, i_13_316_1911_0, i_13_316_1998_0, i_13_316_1999_0,
    i_13_316_2001_0, i_13_316_2019_0, i_13_316_2020_0, i_13_316_2148_0,
    i_13_316_2425_0, i_13_316_2437_0, i_13_316_2448_0, i_13_316_2467_0,
    i_13_316_2469_0, i_13_316_2514_0, i_13_316_2515_0, i_13_316_2626_0,
    i_13_316_2740_0, i_13_316_2910_0, i_13_316_2955_0, i_13_316_2958_0,
    i_13_316_3027_0, i_13_316_3046_0, i_13_316_3072_0, i_13_316_3073_0,
    i_13_316_3108_0, i_13_316_3127_0, i_13_316_3261_0, i_13_316_3262_0,
    i_13_316_3486_0, i_13_316_3549_0, i_13_316_3550_0, i_13_316_3565_0,
    i_13_316_3567_0, i_13_316_3573_0, i_13_316_3648_0, i_13_316_3819_0,
    i_13_316_3891_0, i_13_316_3897_0, i_13_316_3909_0, i_13_316_3910_0,
    i_13_316_3990_0, i_13_316_4158_0, i_13_316_4159_0, i_13_316_4161_0,
    i_13_316_4162_0, i_13_316_4251_0, i_13_316_4293_0, i_13_316_4333_0,
    i_13_316_4336_0, i_13_316_4365_0, i_13_316_4368_0, i_13_316_4369_0,
    i_13_316_4434_0, i_13_316_4510_0, i_13_316_4602_0, i_13_316_4603_0,
    o_13_316_0_0  );
  input  i_13_316_40_0, i_13_316_58_0, i_13_316_259_0, i_13_316_276_0,
    i_13_316_369_0, i_13_316_450_0, i_13_316_513_0, i_13_316_526_0,
    i_13_316_552_0, i_13_316_604_0, i_13_316_606_0, i_13_316_607_0,
    i_13_316_610_0, i_13_316_657_0, i_13_316_658_0, i_13_316_660_0,
    i_13_316_661_0, i_13_316_663_0, i_13_316_670_0, i_13_316_678_0,
    i_13_316_829_0, i_13_316_840_0, i_13_316_931_0, i_13_316_936_0,
    i_13_316_939_0, i_13_316_1056_0, i_13_316_1059_0, i_13_316_1060_0,
    i_13_316_1072_0, i_13_316_1102_0, i_13_316_1119_0, i_13_316_1147_0,
    i_13_316_1516_0, i_13_316_1534_0, i_13_316_1606_0, i_13_316_1659_0,
    i_13_316_1660_0, i_13_316_1663_0, i_13_316_1729_0, i_13_316_1731_0,
    i_13_316_1732_0, i_13_316_1764_0, i_13_316_1767_0, i_13_316_1891_0,
    i_13_316_1897_0, i_13_316_1911_0, i_13_316_1998_0, i_13_316_1999_0,
    i_13_316_2001_0, i_13_316_2019_0, i_13_316_2020_0, i_13_316_2148_0,
    i_13_316_2425_0, i_13_316_2437_0, i_13_316_2448_0, i_13_316_2467_0,
    i_13_316_2469_0, i_13_316_2514_0, i_13_316_2515_0, i_13_316_2626_0,
    i_13_316_2740_0, i_13_316_2910_0, i_13_316_2955_0, i_13_316_2958_0,
    i_13_316_3027_0, i_13_316_3046_0, i_13_316_3072_0, i_13_316_3073_0,
    i_13_316_3108_0, i_13_316_3127_0, i_13_316_3261_0, i_13_316_3262_0,
    i_13_316_3486_0, i_13_316_3549_0, i_13_316_3550_0, i_13_316_3565_0,
    i_13_316_3567_0, i_13_316_3573_0, i_13_316_3648_0, i_13_316_3819_0,
    i_13_316_3891_0, i_13_316_3897_0, i_13_316_3909_0, i_13_316_3910_0,
    i_13_316_3990_0, i_13_316_4158_0, i_13_316_4159_0, i_13_316_4161_0,
    i_13_316_4162_0, i_13_316_4251_0, i_13_316_4293_0, i_13_316_4333_0,
    i_13_316_4336_0, i_13_316_4365_0, i_13_316_4368_0, i_13_316_4369_0,
    i_13_316_4434_0, i_13_316_4510_0, i_13_316_4602_0, i_13_316_4603_0;
  output o_13_316_0_0;
  assign o_13_316_0_0 = ~(~i_13_316_4369_0 | (~i_13_316_936_0 & ~i_13_316_3648_0) | (~i_13_316_1767_0 & ~i_13_316_3486_0 & ~i_13_316_3549_0));
endmodule



// Benchmark "kernel_13_317" written by ABC on Sun Jul 19 10:49:47 2020

module kernel_13_317 ( 
    i_13_317_32_0, i_13_317_69_0, i_13_317_93_0, i_13_317_94_0,
    i_13_317_120_0, i_13_317_121_0, i_13_317_157_0, i_13_317_229_0,
    i_13_317_276_0, i_13_317_382_0, i_13_317_446_0, i_13_317_447_0,
    i_13_317_508_0, i_13_317_542_0, i_13_317_564_0, i_13_317_672_0,
    i_13_317_697_0, i_13_317_732_0, i_13_317_733_0, i_13_317_886_0,
    i_13_317_951_0, i_13_317_952_0, i_13_317_1185_0, i_13_317_1226_0,
    i_13_317_1231_0, i_13_317_1303_0, i_13_317_1318_0, i_13_317_1443_0,
    i_13_317_1444_0, i_13_317_1446_0, i_13_317_1498_0, i_13_317_1602_0,
    i_13_317_1626_0, i_13_317_1632_0, i_13_317_1758_0, i_13_317_1786_0,
    i_13_317_1813_0, i_13_317_2012_0, i_13_317_2173_0, i_13_317_2175_0,
    i_13_317_2176_0, i_13_317_2189_0, i_13_317_2208_0, i_13_317_2209_0,
    i_13_317_2262_0, i_13_317_2424_0, i_13_317_2425_0, i_13_317_2427_0,
    i_13_317_2436_0, i_13_317_2463_0, i_13_317_2541_0, i_13_317_2565_0,
    i_13_317_2581_0, i_13_317_2698_0, i_13_317_2749_0, i_13_317_2857_0,
    i_13_317_2939_0, i_13_317_3000_0, i_13_317_3004_0, i_13_317_3019_0,
    i_13_317_3020_0, i_13_317_3037_0, i_13_317_3063_0, i_13_317_3066_0,
    i_13_317_3067_0, i_13_317_3102_0, i_13_317_3129_0, i_13_317_3130_0,
    i_13_317_3147_0, i_13_317_3160_0, i_13_317_3165_0, i_13_317_3274_0,
    i_13_317_3287_0, i_13_317_3307_0, i_13_317_3399_0, i_13_317_3417_0,
    i_13_317_3418_0, i_13_317_3424_0, i_13_317_3426_0, i_13_317_3427_0,
    i_13_317_3441_0, i_13_317_3534_0, i_13_317_3541_0, i_13_317_3702_0,
    i_13_317_3739_0, i_13_317_3801_0, i_13_317_3843_0, i_13_317_3844_0,
    i_13_317_3980_0, i_13_317_3990_0, i_13_317_4008_0, i_13_317_4009_0,
    i_13_317_4021_0, i_13_317_4054_0, i_13_317_4251_0, i_13_317_4341_0,
    i_13_317_4353_0, i_13_317_4380_0, i_13_317_4560_0, i_13_317_4561_0,
    o_13_317_0_0  );
  input  i_13_317_32_0, i_13_317_69_0, i_13_317_93_0, i_13_317_94_0,
    i_13_317_120_0, i_13_317_121_0, i_13_317_157_0, i_13_317_229_0,
    i_13_317_276_0, i_13_317_382_0, i_13_317_446_0, i_13_317_447_0,
    i_13_317_508_0, i_13_317_542_0, i_13_317_564_0, i_13_317_672_0,
    i_13_317_697_0, i_13_317_732_0, i_13_317_733_0, i_13_317_886_0,
    i_13_317_951_0, i_13_317_952_0, i_13_317_1185_0, i_13_317_1226_0,
    i_13_317_1231_0, i_13_317_1303_0, i_13_317_1318_0, i_13_317_1443_0,
    i_13_317_1444_0, i_13_317_1446_0, i_13_317_1498_0, i_13_317_1602_0,
    i_13_317_1626_0, i_13_317_1632_0, i_13_317_1758_0, i_13_317_1786_0,
    i_13_317_1813_0, i_13_317_2012_0, i_13_317_2173_0, i_13_317_2175_0,
    i_13_317_2176_0, i_13_317_2189_0, i_13_317_2208_0, i_13_317_2209_0,
    i_13_317_2262_0, i_13_317_2424_0, i_13_317_2425_0, i_13_317_2427_0,
    i_13_317_2436_0, i_13_317_2463_0, i_13_317_2541_0, i_13_317_2565_0,
    i_13_317_2581_0, i_13_317_2698_0, i_13_317_2749_0, i_13_317_2857_0,
    i_13_317_2939_0, i_13_317_3000_0, i_13_317_3004_0, i_13_317_3019_0,
    i_13_317_3020_0, i_13_317_3037_0, i_13_317_3063_0, i_13_317_3066_0,
    i_13_317_3067_0, i_13_317_3102_0, i_13_317_3129_0, i_13_317_3130_0,
    i_13_317_3147_0, i_13_317_3160_0, i_13_317_3165_0, i_13_317_3274_0,
    i_13_317_3287_0, i_13_317_3307_0, i_13_317_3399_0, i_13_317_3417_0,
    i_13_317_3418_0, i_13_317_3424_0, i_13_317_3426_0, i_13_317_3427_0,
    i_13_317_3441_0, i_13_317_3534_0, i_13_317_3541_0, i_13_317_3702_0,
    i_13_317_3739_0, i_13_317_3801_0, i_13_317_3843_0, i_13_317_3844_0,
    i_13_317_3980_0, i_13_317_3990_0, i_13_317_4008_0, i_13_317_4009_0,
    i_13_317_4021_0, i_13_317_4054_0, i_13_317_4251_0, i_13_317_4341_0,
    i_13_317_4353_0, i_13_317_4380_0, i_13_317_4560_0, i_13_317_4561_0;
  output o_13_317_0_0;
  assign o_13_317_0_0 = ~((~i_13_317_2436_0 & (~i_13_317_951_0 | (~i_13_317_3441_0 & ~i_13_317_4009_0))) | (~i_13_317_447_0 & ~i_13_317_3427_0) | (~i_13_317_1813_0 & ~i_13_317_3102_0 & ~i_13_317_3147_0 & ~i_13_317_4008_0));
endmodule



// Benchmark "kernel_13_318" written by ABC on Sun Jul 19 10:49:48 2020

module kernel_13_318 ( 
    i_13_318_73_0, i_13_318_74_0, i_13_318_121_0, i_13_318_139_0,
    i_13_318_182_0, i_13_318_184_0, i_13_318_185_0, i_13_318_193_0,
    i_13_318_229_0, i_13_318_235_0, i_13_318_253_0, i_13_318_355_0,
    i_13_318_415_0, i_13_318_469_0, i_13_318_470_0, i_13_318_590_0,
    i_13_318_668_0, i_13_318_694_0, i_13_318_695_0, i_13_318_743_0,
    i_13_318_829_0, i_13_318_947_0, i_13_318_1072_0, i_13_318_1073_0,
    i_13_318_1118_0, i_13_318_1145_0, i_13_318_1208_0, i_13_318_1247_0,
    i_13_318_1307_0, i_13_318_1408_0, i_13_318_1424_0, i_13_318_1522_0,
    i_13_318_1523_0, i_13_318_1536_0, i_13_318_1549_0, i_13_318_1658_0,
    i_13_318_1667_0, i_13_318_1723_0, i_13_318_1742_0, i_13_318_1774_0,
    i_13_318_1849_0, i_13_318_1919_0, i_13_318_1998_0, i_13_318_2000_0,
    i_13_318_2017_0, i_13_318_2021_0, i_13_318_2056_0, i_13_318_2057_0,
    i_13_318_2126_0, i_13_318_2143_0, i_13_318_2144_0, i_13_318_2308_0,
    i_13_318_2425_0, i_13_318_2444_0, i_13_318_2449_0, i_13_318_2450_0,
    i_13_318_2512_0, i_13_318_2513_0, i_13_318_2539_0, i_13_318_2660_0,
    i_13_318_2692_0, i_13_318_2855_0, i_13_318_2881_0, i_13_318_2882_0,
    i_13_318_2907_0, i_13_318_3010_0, i_13_318_3025_0, i_13_318_3037_0,
    i_13_318_3128_0, i_13_318_3254_0, i_13_318_3269_0, i_13_318_3415_0,
    i_13_318_3416_0, i_13_318_3610_0, i_13_318_3620_0, i_13_318_3683_0,
    i_13_318_3863_0, i_13_318_3865_0, i_13_318_3874_0, i_13_318_3916_0,
    i_13_318_3919_0, i_13_318_3921_0, i_13_318_3988_0, i_13_318_4009_0,
    i_13_318_4118_0, i_13_318_4180_0, i_13_318_4253_0, i_13_318_4262_0,
    i_13_318_4271_0, i_13_318_4330_0, i_13_318_4331_0, i_13_318_4366_0,
    i_13_318_4430_0, i_13_318_4529_0, i_13_318_4538_0, i_13_318_4583_0,
    i_13_318_4591_0, i_13_318_4592_0, i_13_318_4601_0, i_13_318_4604_0,
    o_13_318_0_0  );
  input  i_13_318_73_0, i_13_318_74_0, i_13_318_121_0, i_13_318_139_0,
    i_13_318_182_0, i_13_318_184_0, i_13_318_185_0, i_13_318_193_0,
    i_13_318_229_0, i_13_318_235_0, i_13_318_253_0, i_13_318_355_0,
    i_13_318_415_0, i_13_318_469_0, i_13_318_470_0, i_13_318_590_0,
    i_13_318_668_0, i_13_318_694_0, i_13_318_695_0, i_13_318_743_0,
    i_13_318_829_0, i_13_318_947_0, i_13_318_1072_0, i_13_318_1073_0,
    i_13_318_1118_0, i_13_318_1145_0, i_13_318_1208_0, i_13_318_1247_0,
    i_13_318_1307_0, i_13_318_1408_0, i_13_318_1424_0, i_13_318_1522_0,
    i_13_318_1523_0, i_13_318_1536_0, i_13_318_1549_0, i_13_318_1658_0,
    i_13_318_1667_0, i_13_318_1723_0, i_13_318_1742_0, i_13_318_1774_0,
    i_13_318_1849_0, i_13_318_1919_0, i_13_318_1998_0, i_13_318_2000_0,
    i_13_318_2017_0, i_13_318_2021_0, i_13_318_2056_0, i_13_318_2057_0,
    i_13_318_2126_0, i_13_318_2143_0, i_13_318_2144_0, i_13_318_2308_0,
    i_13_318_2425_0, i_13_318_2444_0, i_13_318_2449_0, i_13_318_2450_0,
    i_13_318_2512_0, i_13_318_2513_0, i_13_318_2539_0, i_13_318_2660_0,
    i_13_318_2692_0, i_13_318_2855_0, i_13_318_2881_0, i_13_318_2882_0,
    i_13_318_2907_0, i_13_318_3010_0, i_13_318_3025_0, i_13_318_3037_0,
    i_13_318_3128_0, i_13_318_3254_0, i_13_318_3269_0, i_13_318_3415_0,
    i_13_318_3416_0, i_13_318_3610_0, i_13_318_3620_0, i_13_318_3683_0,
    i_13_318_3863_0, i_13_318_3865_0, i_13_318_3874_0, i_13_318_3916_0,
    i_13_318_3919_0, i_13_318_3921_0, i_13_318_3988_0, i_13_318_4009_0,
    i_13_318_4118_0, i_13_318_4180_0, i_13_318_4253_0, i_13_318_4262_0,
    i_13_318_4271_0, i_13_318_4330_0, i_13_318_4331_0, i_13_318_4366_0,
    i_13_318_4430_0, i_13_318_4529_0, i_13_318_4538_0, i_13_318_4583_0,
    i_13_318_4591_0, i_13_318_4592_0, i_13_318_4601_0, i_13_318_4604_0;
  output o_13_318_0_0;
  assign o_13_318_0_0 = ~((~i_13_318_2021_0 & ~i_13_318_4331_0) | (~i_13_318_1424_0 & ~i_13_318_2126_0 & ~i_13_318_4330_0));
endmodule



// Benchmark "kernel_13_319" written by ABC on Sun Jul 19 10:49:49 2020

module kernel_13_319 ( 
    i_13_319_95_0, i_13_319_136_0, i_13_319_137_0, i_13_319_139_0,
    i_13_319_140_0, i_13_319_202_0, i_13_319_226_0, i_13_319_230_0,
    i_13_319_262_0, i_13_319_383_0, i_13_319_384_0, i_13_319_418_0,
    i_13_319_607_0, i_13_319_618_0, i_13_319_686_0, i_13_319_688_0,
    i_13_319_725_0, i_13_319_779_0, i_13_319_824_0, i_13_319_985_0,
    i_13_319_1094_0, i_13_319_1217_0, i_13_319_1265_0, i_13_319_1270_0,
    i_13_319_1274_0, i_13_319_1282_0, i_13_319_1442_0, i_13_319_1462_0,
    i_13_319_1499_0, i_13_319_1552_0, i_13_319_1712_0, i_13_319_1723_0,
    i_13_319_1778_0, i_13_319_1802_0, i_13_319_1832_0, i_13_319_1837_0,
    i_13_319_1882_0, i_13_319_1883_0, i_13_319_1885_0, i_13_319_1886_0,
    i_13_319_1993_0, i_13_319_1994_0, i_13_319_1999_0, i_13_319_2000_0,
    i_13_319_2018_0, i_13_319_2054_0, i_13_319_2120_0, i_13_319_2170_0,
    i_13_319_2192_0, i_13_319_2207_0, i_13_319_2224_0, i_13_319_2314_0,
    i_13_319_2426_0, i_13_319_2593_0, i_13_319_2647_0, i_13_319_2648_0,
    i_13_319_2651_0, i_13_319_2845_0, i_13_319_2848_0, i_13_319_2849_0,
    i_13_319_2857_0, i_13_319_2875_0, i_13_319_2885_0, i_13_319_3044_0,
    i_13_319_3065_0, i_13_319_3091_0, i_13_319_3143_0, i_13_319_3154_0,
    i_13_319_3164_0, i_13_319_3322_0, i_13_319_3368_0, i_13_319_3389_0,
    i_13_319_3424_0, i_13_319_3425_0, i_13_319_3444_0, i_13_319_3478_0,
    i_13_319_3487_0, i_13_319_3488_0, i_13_319_3556_0, i_13_319_3686_0,
    i_13_319_3791_0, i_13_319_3794_0, i_13_319_3799_0, i_13_319_3836_0,
    i_13_319_3841_0, i_13_319_3992_0, i_13_319_4025_0, i_13_319_4051_0,
    i_13_319_4097_0, i_13_319_4124_0, i_13_319_4186_0, i_13_319_4187_0,
    i_13_319_4235_0, i_13_319_4295_0, i_13_319_4301_0, i_13_319_4369_0,
    i_13_319_4394_0, i_13_319_4397_0, i_13_319_4501_0, i_13_319_4568_0,
    o_13_319_0_0  );
  input  i_13_319_95_0, i_13_319_136_0, i_13_319_137_0, i_13_319_139_0,
    i_13_319_140_0, i_13_319_202_0, i_13_319_226_0, i_13_319_230_0,
    i_13_319_262_0, i_13_319_383_0, i_13_319_384_0, i_13_319_418_0,
    i_13_319_607_0, i_13_319_618_0, i_13_319_686_0, i_13_319_688_0,
    i_13_319_725_0, i_13_319_779_0, i_13_319_824_0, i_13_319_985_0,
    i_13_319_1094_0, i_13_319_1217_0, i_13_319_1265_0, i_13_319_1270_0,
    i_13_319_1274_0, i_13_319_1282_0, i_13_319_1442_0, i_13_319_1462_0,
    i_13_319_1499_0, i_13_319_1552_0, i_13_319_1712_0, i_13_319_1723_0,
    i_13_319_1778_0, i_13_319_1802_0, i_13_319_1832_0, i_13_319_1837_0,
    i_13_319_1882_0, i_13_319_1883_0, i_13_319_1885_0, i_13_319_1886_0,
    i_13_319_1993_0, i_13_319_1994_0, i_13_319_1999_0, i_13_319_2000_0,
    i_13_319_2018_0, i_13_319_2054_0, i_13_319_2120_0, i_13_319_2170_0,
    i_13_319_2192_0, i_13_319_2207_0, i_13_319_2224_0, i_13_319_2314_0,
    i_13_319_2426_0, i_13_319_2593_0, i_13_319_2647_0, i_13_319_2648_0,
    i_13_319_2651_0, i_13_319_2845_0, i_13_319_2848_0, i_13_319_2849_0,
    i_13_319_2857_0, i_13_319_2875_0, i_13_319_2885_0, i_13_319_3044_0,
    i_13_319_3065_0, i_13_319_3091_0, i_13_319_3143_0, i_13_319_3154_0,
    i_13_319_3164_0, i_13_319_3322_0, i_13_319_3368_0, i_13_319_3389_0,
    i_13_319_3424_0, i_13_319_3425_0, i_13_319_3444_0, i_13_319_3478_0,
    i_13_319_3487_0, i_13_319_3488_0, i_13_319_3556_0, i_13_319_3686_0,
    i_13_319_3791_0, i_13_319_3794_0, i_13_319_3799_0, i_13_319_3836_0,
    i_13_319_3841_0, i_13_319_3992_0, i_13_319_4025_0, i_13_319_4051_0,
    i_13_319_4097_0, i_13_319_4124_0, i_13_319_4186_0, i_13_319_4187_0,
    i_13_319_4235_0, i_13_319_4295_0, i_13_319_4301_0, i_13_319_4369_0,
    i_13_319_4394_0, i_13_319_4397_0, i_13_319_4501_0, i_13_319_4568_0;
  output o_13_319_0_0;
  assign o_13_319_0_0 = ~(~i_13_319_1886_0 | (~i_13_319_1712_0 & ~i_13_319_2207_0));
endmodule



// Benchmark "kernel_13_320" written by ABC on Sun Jul 19 10:49:50 2020

module kernel_13_320 ( 
    i_13_320_61_0, i_13_320_65_0, i_13_320_76_0, i_13_320_111_0,
    i_13_320_112_0, i_13_320_186_0, i_13_320_187_0, i_13_320_283_0,
    i_13_320_309_0, i_13_320_382_0, i_13_320_406_0, i_13_320_473_0,
    i_13_320_532_0, i_13_320_571_0, i_13_320_573_0, i_13_320_574_0,
    i_13_320_623_0, i_13_320_643_0, i_13_320_646_0, i_13_320_717_0,
    i_13_320_780_0, i_13_320_814_0, i_13_320_889_0, i_13_320_1073_0,
    i_13_320_1201_0, i_13_320_1210_0, i_13_320_1271_0, i_13_320_1388_0,
    i_13_320_1390_0, i_13_320_1426_0, i_13_320_1492_0, i_13_320_1525_0,
    i_13_320_1528_0, i_13_320_1542_0, i_13_320_1633_0, i_13_320_1640_0,
    i_13_320_1641_0, i_13_320_1642_0, i_13_320_1677_0, i_13_320_1680_0,
    i_13_320_1721_0, i_13_320_1749_0, i_13_320_1793_0, i_13_320_1803_0,
    i_13_320_1804_0, i_13_320_1870_0, i_13_320_1993_0, i_13_320_2014_0,
    i_13_320_2103_0, i_13_320_2197_0, i_13_320_2211_0, i_13_320_2212_0,
    i_13_320_2262_0, i_13_320_2272_0, i_13_320_2407_0, i_13_320_2428_0,
    i_13_320_2452_0, i_13_320_2535_0, i_13_320_2616_0, i_13_320_2649_0,
    i_13_320_2653_0, i_13_320_2679_0, i_13_320_2846_0, i_13_320_3027_0,
    i_13_320_3028_0, i_13_320_3089_0, i_13_320_3166_0, i_13_320_3207_0,
    i_13_320_3208_0, i_13_320_3292_0, i_13_320_3378_0, i_13_320_3387_0,
    i_13_320_3424_0, i_13_320_3426_0, i_13_320_3476_0, i_13_320_3480_0,
    i_13_320_3561_0, i_13_320_3610_0, i_13_320_3649_0, i_13_320_3755_0,
    i_13_320_3836_0, i_13_320_3859_0, i_13_320_3904_0, i_13_320_3991_0,
    i_13_320_3994_0, i_13_320_4011_0, i_13_320_4012_0, i_13_320_4021_0,
    i_13_320_4073_0, i_13_320_4079_0, i_13_320_4080_0, i_13_320_4083_0,
    i_13_320_4183_0, i_13_320_4188_0, i_13_320_4264_0, i_13_320_4295_0,
    i_13_320_4411_0, i_13_320_4558_0, i_13_320_4587_0, i_13_320_4596_0,
    o_13_320_0_0  );
  input  i_13_320_61_0, i_13_320_65_0, i_13_320_76_0, i_13_320_111_0,
    i_13_320_112_0, i_13_320_186_0, i_13_320_187_0, i_13_320_283_0,
    i_13_320_309_0, i_13_320_382_0, i_13_320_406_0, i_13_320_473_0,
    i_13_320_532_0, i_13_320_571_0, i_13_320_573_0, i_13_320_574_0,
    i_13_320_623_0, i_13_320_643_0, i_13_320_646_0, i_13_320_717_0,
    i_13_320_780_0, i_13_320_814_0, i_13_320_889_0, i_13_320_1073_0,
    i_13_320_1201_0, i_13_320_1210_0, i_13_320_1271_0, i_13_320_1388_0,
    i_13_320_1390_0, i_13_320_1426_0, i_13_320_1492_0, i_13_320_1525_0,
    i_13_320_1528_0, i_13_320_1542_0, i_13_320_1633_0, i_13_320_1640_0,
    i_13_320_1641_0, i_13_320_1642_0, i_13_320_1677_0, i_13_320_1680_0,
    i_13_320_1721_0, i_13_320_1749_0, i_13_320_1793_0, i_13_320_1803_0,
    i_13_320_1804_0, i_13_320_1870_0, i_13_320_1993_0, i_13_320_2014_0,
    i_13_320_2103_0, i_13_320_2197_0, i_13_320_2211_0, i_13_320_2212_0,
    i_13_320_2262_0, i_13_320_2272_0, i_13_320_2407_0, i_13_320_2428_0,
    i_13_320_2452_0, i_13_320_2535_0, i_13_320_2616_0, i_13_320_2649_0,
    i_13_320_2653_0, i_13_320_2679_0, i_13_320_2846_0, i_13_320_3027_0,
    i_13_320_3028_0, i_13_320_3089_0, i_13_320_3166_0, i_13_320_3207_0,
    i_13_320_3208_0, i_13_320_3292_0, i_13_320_3378_0, i_13_320_3387_0,
    i_13_320_3424_0, i_13_320_3426_0, i_13_320_3476_0, i_13_320_3480_0,
    i_13_320_3561_0, i_13_320_3610_0, i_13_320_3649_0, i_13_320_3755_0,
    i_13_320_3836_0, i_13_320_3859_0, i_13_320_3904_0, i_13_320_3991_0,
    i_13_320_3994_0, i_13_320_4011_0, i_13_320_4012_0, i_13_320_4021_0,
    i_13_320_4073_0, i_13_320_4079_0, i_13_320_4080_0, i_13_320_4083_0,
    i_13_320_4183_0, i_13_320_4188_0, i_13_320_4264_0, i_13_320_4295_0,
    i_13_320_4411_0, i_13_320_4558_0, i_13_320_4587_0, i_13_320_4596_0;
  output o_13_320_0_0;
  assign o_13_320_0_0 = ~((~i_13_320_3166_0 & ((~i_13_320_1642_0 & ~i_13_320_2212_0) | (i_13_320_2452_0 & ~i_13_320_3426_0))) | (~i_13_320_1749_0 & ~i_13_320_1803_0) | (~i_13_320_382_0 & ~i_13_320_2407_0 & ~i_13_320_4012_0) | (~i_13_320_1993_0 & ~i_13_320_4083_0) | (~i_13_320_1641_0 & i_13_320_4188_0) | (~i_13_320_309_0 & ~i_13_320_4188_0));
endmodule



// Benchmark "kernel_13_321" written by ABC on Sun Jul 19 10:49:50 2020

module kernel_13_321 ( 
    i_13_321_36_0, i_13_321_39_0, i_13_321_40_0, i_13_321_42_0,
    i_13_321_49_0, i_13_321_70_0, i_13_321_137_0, i_13_321_306_0,
    i_13_321_454_0, i_13_321_492_0, i_13_321_585_0, i_13_321_643_0,
    i_13_321_688_0, i_13_321_689_0, i_13_321_690_0, i_13_321_697_0,
    i_13_321_726_0, i_13_321_823_0, i_13_321_826_0, i_13_321_1084_0,
    i_13_321_1271_0, i_13_321_1272_0, i_13_321_1278_0, i_13_321_1279_0,
    i_13_321_1299_0, i_13_321_1303_0, i_13_321_1347_0, i_13_321_1391_0,
    i_13_321_1465_0, i_13_321_1593_0, i_13_321_1600_0, i_13_321_1638_0,
    i_13_321_1642_0, i_13_321_1669_0, i_13_321_1672_0, i_13_321_1759_0,
    i_13_321_1792_0, i_13_321_1831_0, i_13_321_1837_0, i_13_321_1845_0,
    i_13_321_1884_0, i_13_321_1885_0, i_13_321_2059_0, i_13_321_2082_0,
    i_13_321_2104_0, i_13_321_2140_0, i_13_321_2161_0, i_13_321_2199_0,
    i_13_321_2239_0, i_13_321_2378_0, i_13_321_2380_0, i_13_321_2434_0,
    i_13_321_2554_0, i_13_321_2589_0, i_13_321_2650_0, i_13_321_2652_0,
    i_13_321_2653_0, i_13_321_2694_0, i_13_321_2761_0, i_13_321_2823_0,
    i_13_321_2824_0, i_13_321_2848_0, i_13_321_2871_0, i_13_321_3001_0,
    i_13_321_3006_0, i_13_321_3114_0, i_13_321_3130_0, i_13_321_3151_0,
    i_13_321_3156_0, i_13_321_3387_0, i_13_321_3388_0, i_13_321_3390_0,
    i_13_321_3391_0, i_13_321_3394_0, i_13_321_3538_0, i_13_321_3541_0,
    i_13_321_3597_0, i_13_321_3633_0, i_13_321_3766_0, i_13_321_3816_0,
    i_13_321_3874_0, i_13_321_3877_0, i_13_321_3895_0, i_13_321_3912_0,
    i_13_321_3925_0, i_13_321_4014_0, i_13_321_4039_0, i_13_321_4162_0,
    i_13_321_4187_0, i_13_321_4197_0, i_13_321_4203_0, i_13_321_4297_0,
    i_13_321_4341_0, i_13_321_4351_0, i_13_321_4356_0, i_13_321_4368_0,
    i_13_321_4369_0, i_13_321_4381_0, i_13_321_4429_0, i_13_321_4554_0,
    o_13_321_0_0  );
  input  i_13_321_36_0, i_13_321_39_0, i_13_321_40_0, i_13_321_42_0,
    i_13_321_49_0, i_13_321_70_0, i_13_321_137_0, i_13_321_306_0,
    i_13_321_454_0, i_13_321_492_0, i_13_321_585_0, i_13_321_643_0,
    i_13_321_688_0, i_13_321_689_0, i_13_321_690_0, i_13_321_697_0,
    i_13_321_726_0, i_13_321_823_0, i_13_321_826_0, i_13_321_1084_0,
    i_13_321_1271_0, i_13_321_1272_0, i_13_321_1278_0, i_13_321_1279_0,
    i_13_321_1299_0, i_13_321_1303_0, i_13_321_1347_0, i_13_321_1391_0,
    i_13_321_1465_0, i_13_321_1593_0, i_13_321_1600_0, i_13_321_1638_0,
    i_13_321_1642_0, i_13_321_1669_0, i_13_321_1672_0, i_13_321_1759_0,
    i_13_321_1792_0, i_13_321_1831_0, i_13_321_1837_0, i_13_321_1845_0,
    i_13_321_1884_0, i_13_321_1885_0, i_13_321_2059_0, i_13_321_2082_0,
    i_13_321_2104_0, i_13_321_2140_0, i_13_321_2161_0, i_13_321_2199_0,
    i_13_321_2239_0, i_13_321_2378_0, i_13_321_2380_0, i_13_321_2434_0,
    i_13_321_2554_0, i_13_321_2589_0, i_13_321_2650_0, i_13_321_2652_0,
    i_13_321_2653_0, i_13_321_2694_0, i_13_321_2761_0, i_13_321_2823_0,
    i_13_321_2824_0, i_13_321_2848_0, i_13_321_2871_0, i_13_321_3001_0,
    i_13_321_3006_0, i_13_321_3114_0, i_13_321_3130_0, i_13_321_3151_0,
    i_13_321_3156_0, i_13_321_3387_0, i_13_321_3388_0, i_13_321_3390_0,
    i_13_321_3391_0, i_13_321_3394_0, i_13_321_3538_0, i_13_321_3541_0,
    i_13_321_3597_0, i_13_321_3633_0, i_13_321_3766_0, i_13_321_3816_0,
    i_13_321_3874_0, i_13_321_3877_0, i_13_321_3895_0, i_13_321_3912_0,
    i_13_321_3925_0, i_13_321_4014_0, i_13_321_4039_0, i_13_321_4162_0,
    i_13_321_4187_0, i_13_321_4197_0, i_13_321_4203_0, i_13_321_4297_0,
    i_13_321_4341_0, i_13_321_4351_0, i_13_321_4356_0, i_13_321_4368_0,
    i_13_321_4369_0, i_13_321_4381_0, i_13_321_4429_0, i_13_321_4554_0;
  output o_13_321_0_0;
  assign o_13_321_0_0 = ~((i_13_321_1831_0 & ~i_13_321_4381_0 & (i_13_321_2434_0 | (~i_13_321_697_0 & ~i_13_321_3538_0 & ~i_13_321_3912_0))) | (~i_13_321_2650_0 & (~i_13_321_1642_0 | (~i_13_321_3541_0 & i_13_321_3766_0))) | (~i_13_321_1885_0 & ~i_13_321_3391_0 & ~i_13_321_3597_0) | (~i_13_321_2140_0 & ~i_13_321_3387_0 & ~i_13_321_3633_0 & ~i_13_321_3912_0));
endmodule



// Benchmark "kernel_13_322" written by ABC on Sun Jul 19 10:49:51 2020

module kernel_13_322 ( 
    i_13_322_45_0, i_13_322_103_0, i_13_322_120_0, i_13_322_139_0,
    i_13_322_172_0, i_13_322_189_0, i_13_322_202_0, i_13_322_229_0,
    i_13_322_408_0, i_13_322_414_0, i_13_322_549_0, i_13_322_568_0,
    i_13_322_604_0, i_13_322_606_0, i_13_322_625_0, i_13_322_642_0,
    i_13_322_643_0, i_13_322_648_0, i_13_322_657_0, i_13_322_684_0,
    i_13_322_685_0, i_13_322_796_0, i_13_322_936_0, i_13_322_982_0,
    i_13_322_1071_0, i_13_322_1191_0, i_13_322_1225_0, i_13_322_1228_0,
    i_13_322_1272_0, i_13_322_1282_0, i_13_322_1300_0, i_13_322_1404_0,
    i_13_322_1432_0, i_13_322_1498_0, i_13_322_1521_0, i_13_322_1548_0,
    i_13_322_1560_0, i_13_322_1629_0, i_13_322_1674_0, i_13_322_1677_0,
    i_13_322_1729_0, i_13_322_1750_0, i_13_322_1767_0, i_13_322_1768_0,
    i_13_322_1795_0, i_13_322_1803_0, i_13_322_1804_0, i_13_322_1808_0,
    i_13_322_1854_0, i_13_322_1896_0, i_13_322_1911_0, i_13_322_2001_0,
    i_13_322_2019_0, i_13_322_2020_0, i_13_322_2047_0, i_13_322_2119_0,
    i_13_322_2286_0, i_13_322_2314_0, i_13_322_2361_0, i_13_322_2469_0,
    i_13_322_2470_0, i_13_322_2542_0, i_13_322_2578_0, i_13_322_2691_0,
    i_13_322_2979_0, i_13_322_3000_0, i_13_322_3006_0, i_13_322_3009_0,
    i_13_322_3027_0, i_13_322_3028_0, i_13_322_3105_0, i_13_322_3204_0,
    i_13_322_3205_0, i_13_322_3208_0, i_13_322_3261_0, i_13_322_3396_0,
    i_13_322_3420_0, i_13_322_3475_0, i_13_322_3483_0, i_13_322_3522_0,
    i_13_322_3546_0, i_13_322_3573_0, i_13_322_3657_0, i_13_322_3811_0,
    i_13_322_3819_0, i_13_322_3820_0, i_13_322_3897_0, i_13_322_3898_0,
    i_13_322_3907_0, i_13_322_3978_0, i_13_322_3990_0, i_13_322_4248_0,
    i_13_322_4251_0, i_13_322_4269_0, i_13_322_4332_0, i_13_322_4392_0,
    i_13_322_4404_0, i_13_322_4582_0, i_13_322_4594_0, i_13_322_4603_0,
    o_13_322_0_0  );
  input  i_13_322_45_0, i_13_322_103_0, i_13_322_120_0, i_13_322_139_0,
    i_13_322_172_0, i_13_322_189_0, i_13_322_202_0, i_13_322_229_0,
    i_13_322_408_0, i_13_322_414_0, i_13_322_549_0, i_13_322_568_0,
    i_13_322_604_0, i_13_322_606_0, i_13_322_625_0, i_13_322_642_0,
    i_13_322_643_0, i_13_322_648_0, i_13_322_657_0, i_13_322_684_0,
    i_13_322_685_0, i_13_322_796_0, i_13_322_936_0, i_13_322_982_0,
    i_13_322_1071_0, i_13_322_1191_0, i_13_322_1225_0, i_13_322_1228_0,
    i_13_322_1272_0, i_13_322_1282_0, i_13_322_1300_0, i_13_322_1404_0,
    i_13_322_1432_0, i_13_322_1498_0, i_13_322_1521_0, i_13_322_1548_0,
    i_13_322_1560_0, i_13_322_1629_0, i_13_322_1674_0, i_13_322_1677_0,
    i_13_322_1729_0, i_13_322_1750_0, i_13_322_1767_0, i_13_322_1768_0,
    i_13_322_1795_0, i_13_322_1803_0, i_13_322_1804_0, i_13_322_1808_0,
    i_13_322_1854_0, i_13_322_1896_0, i_13_322_1911_0, i_13_322_2001_0,
    i_13_322_2019_0, i_13_322_2020_0, i_13_322_2047_0, i_13_322_2119_0,
    i_13_322_2286_0, i_13_322_2314_0, i_13_322_2361_0, i_13_322_2469_0,
    i_13_322_2470_0, i_13_322_2542_0, i_13_322_2578_0, i_13_322_2691_0,
    i_13_322_2979_0, i_13_322_3000_0, i_13_322_3006_0, i_13_322_3009_0,
    i_13_322_3027_0, i_13_322_3028_0, i_13_322_3105_0, i_13_322_3204_0,
    i_13_322_3205_0, i_13_322_3208_0, i_13_322_3261_0, i_13_322_3396_0,
    i_13_322_3420_0, i_13_322_3475_0, i_13_322_3483_0, i_13_322_3522_0,
    i_13_322_3546_0, i_13_322_3573_0, i_13_322_3657_0, i_13_322_3811_0,
    i_13_322_3819_0, i_13_322_3820_0, i_13_322_3897_0, i_13_322_3898_0,
    i_13_322_3907_0, i_13_322_3978_0, i_13_322_3990_0, i_13_322_4248_0,
    i_13_322_4251_0, i_13_322_4269_0, i_13_322_4332_0, i_13_322_4392_0,
    i_13_322_4404_0, i_13_322_4582_0, i_13_322_4594_0, i_13_322_4603_0;
  output o_13_322_0_0;
  assign o_13_322_0_0 = ~((~i_13_322_172_0 & ~i_13_322_3396_0) | (~i_13_322_1404_0 & ~i_13_322_2020_0) | (~i_13_322_45_0 & ~i_13_322_1803_0) | (~i_13_322_414_0 & ~i_13_322_648_0 & ~i_13_322_1071_0));
endmodule



// Benchmark "kernel_13_323" written by ABC on Sun Jul 19 10:49:52 2020

module kernel_13_323 ( 
    i_13_323_112_0, i_13_323_142_0, i_13_323_143_0, i_13_323_188_0,
    i_13_323_203_0, i_13_323_229_0, i_13_323_232_0, i_13_323_233_0,
    i_13_323_283_0, i_13_323_341_0, i_13_323_428_0, i_13_323_607_0,
    i_13_323_619_0, i_13_323_643_0, i_13_323_644_0, i_13_323_647_0,
    i_13_323_689_0, i_13_323_692_0, i_13_323_827_0, i_13_323_859_0,
    i_13_323_887_0, i_13_323_931_0, i_13_323_941_0, i_13_323_1079_0,
    i_13_323_1120_0, i_13_323_1121_0, i_13_323_1124_0, i_13_323_1147_0,
    i_13_323_1204_0, i_13_323_1276_0, i_13_323_1277_0, i_13_323_1283_0,
    i_13_323_1346_0, i_13_323_1411_0, i_13_323_1426_0, i_13_323_1448_0,
    i_13_323_1502_0, i_13_323_1520_0, i_13_323_1637_0, i_13_323_1714_0,
    i_13_323_1715_0, i_13_323_1726_0, i_13_323_1786_0, i_13_323_1790_0,
    i_13_323_1796_0, i_13_323_1885_0, i_13_323_1994_0, i_13_323_2005_0,
    i_13_323_2056_0, i_13_323_2137_0, i_13_323_2138_0, i_13_323_2186_0,
    i_13_323_2212_0, i_13_323_2213_0, i_13_323_2263_0, i_13_323_2408_0,
    i_13_323_2428_0, i_13_323_2429_0, i_13_323_2464_0, i_13_323_2542_0,
    i_13_323_2597_0, i_13_323_2614_0, i_13_323_2617_0, i_13_323_2650_0,
    i_13_323_2651_0, i_13_323_2654_0, i_13_323_2848_0, i_13_323_2857_0,
    i_13_323_3040_0, i_13_323_3041_0, i_13_323_3257_0, i_13_323_3308_0,
    i_13_323_3389_0, i_13_323_3392_0, i_13_323_3425_0, i_13_323_3427_0,
    i_13_323_3428_0, i_13_323_3482_0, i_13_323_3541_0, i_13_323_3661_0,
    i_13_323_3724_0, i_13_323_3725_0, i_13_323_3733_0, i_13_323_3856_0,
    i_13_323_3865_0, i_13_323_4012_0, i_13_323_4013_0, i_13_323_4018_0,
    i_13_323_4019_0, i_13_323_4057_0, i_13_323_4081_0, i_13_323_4235_0,
    i_13_323_4307_0, i_13_323_4333_0, i_13_323_4334_0, i_13_323_4369_0,
    i_13_323_4370_0, i_13_323_4415_0, i_13_323_4534_0, i_13_323_4595_0,
    o_13_323_0_0  );
  input  i_13_323_112_0, i_13_323_142_0, i_13_323_143_0, i_13_323_188_0,
    i_13_323_203_0, i_13_323_229_0, i_13_323_232_0, i_13_323_233_0,
    i_13_323_283_0, i_13_323_341_0, i_13_323_428_0, i_13_323_607_0,
    i_13_323_619_0, i_13_323_643_0, i_13_323_644_0, i_13_323_647_0,
    i_13_323_689_0, i_13_323_692_0, i_13_323_827_0, i_13_323_859_0,
    i_13_323_887_0, i_13_323_931_0, i_13_323_941_0, i_13_323_1079_0,
    i_13_323_1120_0, i_13_323_1121_0, i_13_323_1124_0, i_13_323_1147_0,
    i_13_323_1204_0, i_13_323_1276_0, i_13_323_1277_0, i_13_323_1283_0,
    i_13_323_1346_0, i_13_323_1411_0, i_13_323_1426_0, i_13_323_1448_0,
    i_13_323_1502_0, i_13_323_1520_0, i_13_323_1637_0, i_13_323_1714_0,
    i_13_323_1715_0, i_13_323_1726_0, i_13_323_1786_0, i_13_323_1790_0,
    i_13_323_1796_0, i_13_323_1885_0, i_13_323_1994_0, i_13_323_2005_0,
    i_13_323_2056_0, i_13_323_2137_0, i_13_323_2138_0, i_13_323_2186_0,
    i_13_323_2212_0, i_13_323_2213_0, i_13_323_2263_0, i_13_323_2408_0,
    i_13_323_2428_0, i_13_323_2429_0, i_13_323_2464_0, i_13_323_2542_0,
    i_13_323_2597_0, i_13_323_2614_0, i_13_323_2617_0, i_13_323_2650_0,
    i_13_323_2651_0, i_13_323_2654_0, i_13_323_2848_0, i_13_323_2857_0,
    i_13_323_3040_0, i_13_323_3041_0, i_13_323_3257_0, i_13_323_3308_0,
    i_13_323_3389_0, i_13_323_3392_0, i_13_323_3425_0, i_13_323_3427_0,
    i_13_323_3428_0, i_13_323_3482_0, i_13_323_3541_0, i_13_323_3661_0,
    i_13_323_3724_0, i_13_323_3725_0, i_13_323_3733_0, i_13_323_3856_0,
    i_13_323_3865_0, i_13_323_4012_0, i_13_323_4013_0, i_13_323_4018_0,
    i_13_323_4019_0, i_13_323_4057_0, i_13_323_4081_0, i_13_323_4235_0,
    i_13_323_4307_0, i_13_323_4333_0, i_13_323_4334_0, i_13_323_4369_0,
    i_13_323_4370_0, i_13_323_4415_0, i_13_323_4534_0, i_13_323_4595_0;
  output o_13_323_0_0;
  assign o_13_323_0_0 = ~((i_13_323_3541_0 & ~i_13_323_4307_0) | (~i_13_323_2005_0 & ~i_13_323_3428_0) | (~i_13_323_2213_0 & ~i_13_323_2650_0) | (~i_13_323_2138_0 & ~i_13_323_2428_0) | (~i_13_323_1079_0 & ~i_13_323_1714_0 & ~i_13_323_2857_0));
endmodule



// Benchmark "kernel_13_324" written by ABC on Sun Jul 19 10:49:53 2020

module kernel_13_324 ( 
    i_13_324_37_0, i_13_324_64_0, i_13_324_121_0, i_13_324_274_0,
    i_13_324_280_0, i_13_324_331_0, i_13_324_338_0, i_13_324_401_0,
    i_13_324_463_0, i_13_324_526_0, i_13_324_561_0, i_13_324_562_0,
    i_13_324_589_0, i_13_324_608_0, i_13_324_662_0, i_13_324_694_0,
    i_13_324_724_0, i_13_324_823_0, i_13_324_914_0, i_13_324_1066_0,
    i_13_324_1256_0, i_13_324_1309_0, i_13_324_1310_0, i_13_324_1327_0,
    i_13_324_1483_0, i_13_324_1499_0, i_13_324_1561_0, i_13_324_1594_0,
    i_13_324_1595_0, i_13_324_1624_0, i_13_324_1639_0, i_13_324_1661_0,
    i_13_324_1684_0, i_13_324_1729_0, i_13_324_1732_0, i_13_324_1775_0,
    i_13_324_1778_0, i_13_324_1793_0, i_13_324_1795_0, i_13_324_1882_0,
    i_13_324_1883_0, i_13_324_1885_0, i_13_324_1925_0, i_13_324_1927_0,
    i_13_324_1942_0, i_13_324_1943_0, i_13_324_1999_0, i_13_324_2233_0,
    i_13_324_2380_0, i_13_324_2443_0, i_13_324_2558_0, i_13_324_2585_0,
    i_13_324_2650_0, i_13_324_2651_0, i_13_324_2821_0, i_13_324_2872_0,
    i_13_324_2900_0, i_13_324_2914_0, i_13_324_2983_0, i_13_324_3109_0,
    i_13_324_3142_0, i_13_324_3163_0, i_13_324_3215_0, i_13_324_3235_0,
    i_13_324_3271_0, i_13_324_3289_0, i_13_324_3388_0, i_13_324_3389_0,
    i_13_324_3395_0, i_13_324_3523_0, i_13_324_3538_0, i_13_324_3539_0,
    i_13_324_3542_0, i_13_324_3662_0, i_13_324_3667_0, i_13_324_3668_0,
    i_13_324_3728_0, i_13_324_3730_0, i_13_324_3731_0, i_13_324_3739_0,
    i_13_324_3740_0, i_13_324_3766_0, i_13_324_3792_0, i_13_324_3803_0,
    i_13_324_3901_0, i_13_324_3904_0, i_13_324_3916_0, i_13_324_3935_0,
    i_13_324_3989_0, i_13_324_4099_0, i_13_324_4162_0, i_13_324_4324_0,
    i_13_324_4351_0, i_13_324_4364_0, i_13_324_4369_0, i_13_324_4379_0,
    i_13_324_4396_0, i_13_324_4443_0, i_13_324_4540_0, i_13_324_4567_0,
    o_13_324_0_0  );
  input  i_13_324_37_0, i_13_324_64_0, i_13_324_121_0, i_13_324_274_0,
    i_13_324_280_0, i_13_324_331_0, i_13_324_338_0, i_13_324_401_0,
    i_13_324_463_0, i_13_324_526_0, i_13_324_561_0, i_13_324_562_0,
    i_13_324_589_0, i_13_324_608_0, i_13_324_662_0, i_13_324_694_0,
    i_13_324_724_0, i_13_324_823_0, i_13_324_914_0, i_13_324_1066_0,
    i_13_324_1256_0, i_13_324_1309_0, i_13_324_1310_0, i_13_324_1327_0,
    i_13_324_1483_0, i_13_324_1499_0, i_13_324_1561_0, i_13_324_1594_0,
    i_13_324_1595_0, i_13_324_1624_0, i_13_324_1639_0, i_13_324_1661_0,
    i_13_324_1684_0, i_13_324_1729_0, i_13_324_1732_0, i_13_324_1775_0,
    i_13_324_1778_0, i_13_324_1793_0, i_13_324_1795_0, i_13_324_1882_0,
    i_13_324_1883_0, i_13_324_1885_0, i_13_324_1925_0, i_13_324_1927_0,
    i_13_324_1942_0, i_13_324_1943_0, i_13_324_1999_0, i_13_324_2233_0,
    i_13_324_2380_0, i_13_324_2443_0, i_13_324_2558_0, i_13_324_2585_0,
    i_13_324_2650_0, i_13_324_2651_0, i_13_324_2821_0, i_13_324_2872_0,
    i_13_324_2900_0, i_13_324_2914_0, i_13_324_2983_0, i_13_324_3109_0,
    i_13_324_3142_0, i_13_324_3163_0, i_13_324_3215_0, i_13_324_3235_0,
    i_13_324_3271_0, i_13_324_3289_0, i_13_324_3388_0, i_13_324_3389_0,
    i_13_324_3395_0, i_13_324_3523_0, i_13_324_3538_0, i_13_324_3539_0,
    i_13_324_3542_0, i_13_324_3662_0, i_13_324_3667_0, i_13_324_3668_0,
    i_13_324_3728_0, i_13_324_3730_0, i_13_324_3731_0, i_13_324_3739_0,
    i_13_324_3740_0, i_13_324_3766_0, i_13_324_3792_0, i_13_324_3803_0,
    i_13_324_3901_0, i_13_324_3904_0, i_13_324_3916_0, i_13_324_3935_0,
    i_13_324_3989_0, i_13_324_4099_0, i_13_324_4162_0, i_13_324_4324_0,
    i_13_324_4351_0, i_13_324_4364_0, i_13_324_4369_0, i_13_324_4379_0,
    i_13_324_4396_0, i_13_324_4443_0, i_13_324_4540_0, i_13_324_4567_0;
  output o_13_324_0_0;
  assign o_13_324_0_0 = ~((~i_13_324_694_0 & (~i_13_324_2900_0 | (~i_13_324_280_0 & ~i_13_324_3539_0))) | (~i_13_324_1661_0 & ((~i_13_324_2651_0 & i_13_324_3523_0 & ~i_13_324_3539_0) | (~i_13_324_64_0 & ~i_13_324_1793_0 & ~i_13_324_3728_0 & ~i_13_324_3731_0))) | (~i_13_324_2900_0 & (i_13_324_1624_0 | ~i_13_324_4396_0)) | i_13_324_561_0 | (~i_13_324_1885_0 & ~i_13_324_2872_0 & ~i_13_324_3731_0) | (~i_13_324_1883_0 & ~i_13_324_3389_0 & i_13_324_4162_0));
endmodule



// Benchmark "kernel_13_325" written by ABC on Sun Jul 19 10:49:54 2020

module kernel_13_325 ( 
    i_13_325_61_0, i_13_325_62_0, i_13_325_76_0, i_13_325_106_0,
    i_13_325_112_0, i_13_325_166_0, i_13_325_169_0, i_13_325_193_0,
    i_13_325_220_0, i_13_325_382_0, i_13_325_484_0, i_13_325_535_0,
    i_13_325_544_0, i_13_325_573_0, i_13_325_574_0, i_13_325_575_0,
    i_13_325_601_0, i_13_325_728_0, i_13_325_815_0, i_13_325_895_0,
    i_13_325_914_0, i_13_325_1040_0, i_13_325_1093_0, i_13_325_1120_0,
    i_13_325_1124_0, i_13_325_1258_0, i_13_325_1277_0, i_13_325_1393_0,
    i_13_325_1394_0, i_13_325_1411_0, i_13_325_1466_0, i_13_325_1483_0,
    i_13_325_1484_0, i_13_325_1537_0, i_13_325_1561_0, i_13_325_1628_0,
    i_13_325_1643_0, i_13_325_1660_0, i_13_325_1691_0, i_13_325_1723_0,
    i_13_325_1726_0, i_13_325_1727_0, i_13_325_1750_0, i_13_325_1760_0,
    i_13_325_1771_0, i_13_325_1781_0, i_13_325_1786_0, i_13_325_1789_0,
    i_13_325_1796_0, i_13_325_1804_0, i_13_325_1834_0, i_13_325_1858_0,
    i_13_325_1894_0, i_13_325_1907_0, i_13_325_2002_0, i_13_325_2005_0,
    i_13_325_2041_0, i_13_325_2049_0, i_13_325_2150_0, i_13_325_2168_0,
    i_13_325_2212_0, i_13_325_2213_0, i_13_325_2263_0, i_13_325_2408_0,
    i_13_325_2446_0, i_13_325_2542_0, i_13_325_2618_0, i_13_325_2633_0,
    i_13_325_2642_0, i_13_325_2650_0, i_13_325_2654_0, i_13_325_2687_0,
    i_13_325_2750_0, i_13_325_2767_0, i_13_325_2785_0, i_13_325_3001_0,
    i_13_325_3027_0, i_13_325_3041_0, i_13_325_3157_0, i_13_325_3158_0,
    i_13_325_3200_0, i_13_325_3238_0, i_13_325_3308_0, i_13_325_3427_0,
    i_13_325_3433_0, i_13_325_3469_0, i_13_325_3472_0, i_13_325_3522_0,
    i_13_325_3527_0, i_13_325_3562_0, i_13_325_3730_0, i_13_325_3794_0,
    i_13_325_3884_0, i_13_325_3887_0, i_13_325_3976_0, i_13_325_4012_0,
    i_13_325_4081_0, i_13_325_4156_0, i_13_325_4157_0, i_13_325_4325_0,
    o_13_325_0_0  );
  input  i_13_325_61_0, i_13_325_62_0, i_13_325_76_0, i_13_325_106_0,
    i_13_325_112_0, i_13_325_166_0, i_13_325_169_0, i_13_325_193_0,
    i_13_325_220_0, i_13_325_382_0, i_13_325_484_0, i_13_325_535_0,
    i_13_325_544_0, i_13_325_573_0, i_13_325_574_0, i_13_325_575_0,
    i_13_325_601_0, i_13_325_728_0, i_13_325_815_0, i_13_325_895_0,
    i_13_325_914_0, i_13_325_1040_0, i_13_325_1093_0, i_13_325_1120_0,
    i_13_325_1124_0, i_13_325_1258_0, i_13_325_1277_0, i_13_325_1393_0,
    i_13_325_1394_0, i_13_325_1411_0, i_13_325_1466_0, i_13_325_1483_0,
    i_13_325_1484_0, i_13_325_1537_0, i_13_325_1561_0, i_13_325_1628_0,
    i_13_325_1643_0, i_13_325_1660_0, i_13_325_1691_0, i_13_325_1723_0,
    i_13_325_1726_0, i_13_325_1727_0, i_13_325_1750_0, i_13_325_1760_0,
    i_13_325_1771_0, i_13_325_1781_0, i_13_325_1786_0, i_13_325_1789_0,
    i_13_325_1796_0, i_13_325_1804_0, i_13_325_1834_0, i_13_325_1858_0,
    i_13_325_1894_0, i_13_325_1907_0, i_13_325_2002_0, i_13_325_2005_0,
    i_13_325_2041_0, i_13_325_2049_0, i_13_325_2150_0, i_13_325_2168_0,
    i_13_325_2212_0, i_13_325_2213_0, i_13_325_2263_0, i_13_325_2408_0,
    i_13_325_2446_0, i_13_325_2542_0, i_13_325_2618_0, i_13_325_2633_0,
    i_13_325_2642_0, i_13_325_2650_0, i_13_325_2654_0, i_13_325_2687_0,
    i_13_325_2750_0, i_13_325_2767_0, i_13_325_2785_0, i_13_325_3001_0,
    i_13_325_3027_0, i_13_325_3041_0, i_13_325_3157_0, i_13_325_3158_0,
    i_13_325_3200_0, i_13_325_3238_0, i_13_325_3308_0, i_13_325_3427_0,
    i_13_325_3433_0, i_13_325_3469_0, i_13_325_3472_0, i_13_325_3522_0,
    i_13_325_3527_0, i_13_325_3562_0, i_13_325_3730_0, i_13_325_3794_0,
    i_13_325_3884_0, i_13_325_3887_0, i_13_325_3976_0, i_13_325_4012_0,
    i_13_325_4081_0, i_13_325_4156_0, i_13_325_4157_0, i_13_325_4325_0;
  output o_13_325_0_0;
  assign o_13_325_0_0 = ~((~i_13_325_4012_0 & ((~i_13_325_573_0 & ~i_13_325_1277_0) | (~i_13_325_575_0 & ~i_13_325_2446_0))) | (~i_13_325_4325_0 & (~i_13_325_193_0 | (~i_13_325_1643_0 & ~i_13_325_2213_0 & ~i_13_325_3427_0))) | (i_13_325_2005_0 & ~i_13_325_2650_0 & ~i_13_325_4157_0));
endmodule



// Benchmark "kernel_13_326" written by ABC on Sun Jul 19 10:49:54 2020

module kernel_13_326 ( 
    i_13_326_48_0, i_13_326_72_0, i_13_326_73_0, i_13_326_77_0,
    i_13_326_162_0, i_13_326_217_0, i_13_326_226_0, i_13_326_286_0,
    i_13_326_370_0, i_13_326_406_0, i_13_326_463_0, i_13_326_480_0,
    i_13_326_558_0, i_13_326_582_0, i_13_326_583_0, i_13_326_651_0,
    i_13_326_652_0, i_13_326_659_0, i_13_326_675_0, i_13_326_676_0,
    i_13_326_696_0, i_13_326_811_0, i_13_326_939_0, i_13_326_1071_0,
    i_13_326_1074_0, i_13_326_1116_0, i_13_326_1141_0, i_13_326_1143_0,
    i_13_326_1144_0, i_13_326_1145_0, i_13_326_1200_0, i_13_326_1281_0,
    i_13_326_1362_0, i_13_326_1437_0, i_13_326_1549_0, i_13_326_1632_0,
    i_13_326_1656_0, i_13_326_1657_0, i_13_326_1658_0, i_13_326_1720_0,
    i_13_326_1837_0, i_13_326_1839_0, i_13_326_1841_0, i_13_326_2017_0,
    i_13_326_2047_0, i_13_326_2241_0, i_13_326_2317_0, i_13_326_2394_0,
    i_13_326_2404_0, i_13_326_2451_0, i_13_326_2452_0, i_13_326_2468_0,
    i_13_326_2511_0, i_13_326_2550_0, i_13_326_2745_0, i_13_326_2754_0,
    i_13_326_2791_0, i_13_326_2844_0, i_13_326_2845_0, i_13_326_2854_0,
    i_13_326_2883_0, i_13_326_2925_0, i_13_326_2944_0, i_13_326_2955_0,
    i_13_326_2959_0, i_13_326_2986_0, i_13_326_2997_0, i_13_326_2998_0,
    i_13_326_3096_0, i_13_326_3100_0, i_13_326_3105_0, i_13_326_3204_0,
    i_13_326_3447_0, i_13_326_3448_0, i_13_326_3501_0, i_13_326_3522_0,
    i_13_326_3549_0, i_13_326_3567_0, i_13_326_3568_0, i_13_326_3577_0,
    i_13_326_3645_0, i_13_326_3646_0, i_13_326_3663_0, i_13_326_3735_0,
    i_13_326_3847_0, i_13_326_3891_0, i_13_326_3907_0, i_13_326_3933_0,
    i_13_326_4017_0, i_13_326_4095_0, i_13_326_4160_0, i_13_326_4186_0,
    i_13_326_4258_0, i_13_326_4311_0, i_13_326_4329_0, i_13_326_4590_0,
    i_13_326_4591_0, i_13_326_4599_0, i_13_326_4600_0, i_13_326_4601_0,
    o_13_326_0_0  );
  input  i_13_326_48_0, i_13_326_72_0, i_13_326_73_0, i_13_326_77_0,
    i_13_326_162_0, i_13_326_217_0, i_13_326_226_0, i_13_326_286_0,
    i_13_326_370_0, i_13_326_406_0, i_13_326_463_0, i_13_326_480_0,
    i_13_326_558_0, i_13_326_582_0, i_13_326_583_0, i_13_326_651_0,
    i_13_326_652_0, i_13_326_659_0, i_13_326_675_0, i_13_326_676_0,
    i_13_326_696_0, i_13_326_811_0, i_13_326_939_0, i_13_326_1071_0,
    i_13_326_1074_0, i_13_326_1116_0, i_13_326_1141_0, i_13_326_1143_0,
    i_13_326_1144_0, i_13_326_1145_0, i_13_326_1200_0, i_13_326_1281_0,
    i_13_326_1362_0, i_13_326_1437_0, i_13_326_1549_0, i_13_326_1632_0,
    i_13_326_1656_0, i_13_326_1657_0, i_13_326_1658_0, i_13_326_1720_0,
    i_13_326_1837_0, i_13_326_1839_0, i_13_326_1841_0, i_13_326_2017_0,
    i_13_326_2047_0, i_13_326_2241_0, i_13_326_2317_0, i_13_326_2394_0,
    i_13_326_2404_0, i_13_326_2451_0, i_13_326_2452_0, i_13_326_2468_0,
    i_13_326_2511_0, i_13_326_2550_0, i_13_326_2745_0, i_13_326_2754_0,
    i_13_326_2791_0, i_13_326_2844_0, i_13_326_2845_0, i_13_326_2854_0,
    i_13_326_2883_0, i_13_326_2925_0, i_13_326_2944_0, i_13_326_2955_0,
    i_13_326_2959_0, i_13_326_2986_0, i_13_326_2997_0, i_13_326_2998_0,
    i_13_326_3096_0, i_13_326_3100_0, i_13_326_3105_0, i_13_326_3204_0,
    i_13_326_3447_0, i_13_326_3448_0, i_13_326_3501_0, i_13_326_3522_0,
    i_13_326_3549_0, i_13_326_3567_0, i_13_326_3568_0, i_13_326_3577_0,
    i_13_326_3645_0, i_13_326_3646_0, i_13_326_3663_0, i_13_326_3735_0,
    i_13_326_3847_0, i_13_326_3891_0, i_13_326_3907_0, i_13_326_3933_0,
    i_13_326_4017_0, i_13_326_4095_0, i_13_326_4160_0, i_13_326_4186_0,
    i_13_326_4258_0, i_13_326_4311_0, i_13_326_4329_0, i_13_326_4590_0,
    i_13_326_4591_0, i_13_326_4599_0, i_13_326_4600_0, i_13_326_4601_0;
  output o_13_326_0_0;
  assign o_13_326_0_0 = ~(i_13_326_2404_0 | ~i_13_326_1657_0 | (~i_13_326_651_0 & ~i_13_326_3646_0));
endmodule



// Benchmark "kernel_13_327" written by ABC on Sun Jul 19 10:49:55 2020

module kernel_13_327 ( 
    i_13_327_48_0, i_13_327_67_0, i_13_327_69_0, i_13_327_186_0,
    i_13_327_229_0, i_13_327_258_0, i_13_327_285_0, i_13_327_310_0,
    i_13_327_411_0, i_13_327_438_0, i_13_327_520_0, i_13_327_610_0,
    i_13_327_616_0, i_13_327_627_0, i_13_327_628_0, i_13_327_760_0,
    i_13_327_762_0, i_13_327_853_0, i_13_327_934_0, i_13_327_939_0,
    i_13_327_1023_0, i_13_327_1105_0, i_13_327_1132_0, i_13_327_1149_0,
    i_13_327_1150_0, i_13_327_1191_0, i_13_327_1227_0, i_13_327_1317_0,
    i_13_327_1381_0, i_13_327_1402_0, i_13_327_1429_0, i_13_327_1482_0,
    i_13_327_1509_0, i_13_327_1537_0, i_13_327_1563_0, i_13_327_1596_0,
    i_13_327_1597_0, i_13_327_1610_0, i_13_327_1644_0, i_13_327_1651_0,
    i_13_327_1744_0, i_13_327_1753_0, i_13_327_1770_0, i_13_327_1794_0,
    i_13_327_1798_0, i_13_327_1829_0, i_13_327_1838_0, i_13_327_1884_0,
    i_13_327_1922_0, i_13_327_1923_0, i_13_327_1947_0, i_13_327_2022_0,
    i_13_327_2122_0, i_13_327_2199_0, i_13_327_2311_0, i_13_327_2427_0,
    i_13_327_2428_0, i_13_327_2454_0, i_13_327_2472_0, i_13_327_2473_0,
    i_13_327_2506_0, i_13_327_2517_0, i_13_327_2742_0, i_13_327_2743_0,
    i_13_327_2770_0, i_13_327_2940_0, i_13_327_2968_0, i_13_327_3009_0,
    i_13_327_3012_0, i_13_327_3030_0, i_13_327_3031_0, i_13_327_3075_0,
    i_13_327_3076_0, i_13_327_3091_0, i_13_327_3093_0, i_13_327_3211_0,
    i_13_327_3264_0, i_13_327_3273_0, i_13_327_3292_0, i_13_327_3345_0,
    i_13_327_3354_0, i_13_327_3381_0, i_13_327_3382_0, i_13_327_3418_0,
    i_13_327_3435_0, i_13_327_3540_0, i_13_327_3576_0, i_13_327_3759_0,
    i_13_327_3822_0, i_13_327_3900_0, i_13_327_3929_0, i_13_327_4036_0,
    i_13_327_4083_0, i_13_327_4164_0, i_13_327_4272_0, i_13_327_4362_0,
    i_13_327_4450_0, i_13_327_4497_0, i_13_327_4605_0, i_13_327_4606_0,
    o_13_327_0_0  );
  input  i_13_327_48_0, i_13_327_67_0, i_13_327_69_0, i_13_327_186_0,
    i_13_327_229_0, i_13_327_258_0, i_13_327_285_0, i_13_327_310_0,
    i_13_327_411_0, i_13_327_438_0, i_13_327_520_0, i_13_327_610_0,
    i_13_327_616_0, i_13_327_627_0, i_13_327_628_0, i_13_327_760_0,
    i_13_327_762_0, i_13_327_853_0, i_13_327_934_0, i_13_327_939_0,
    i_13_327_1023_0, i_13_327_1105_0, i_13_327_1132_0, i_13_327_1149_0,
    i_13_327_1150_0, i_13_327_1191_0, i_13_327_1227_0, i_13_327_1317_0,
    i_13_327_1381_0, i_13_327_1402_0, i_13_327_1429_0, i_13_327_1482_0,
    i_13_327_1509_0, i_13_327_1537_0, i_13_327_1563_0, i_13_327_1596_0,
    i_13_327_1597_0, i_13_327_1610_0, i_13_327_1644_0, i_13_327_1651_0,
    i_13_327_1744_0, i_13_327_1753_0, i_13_327_1770_0, i_13_327_1794_0,
    i_13_327_1798_0, i_13_327_1829_0, i_13_327_1838_0, i_13_327_1884_0,
    i_13_327_1922_0, i_13_327_1923_0, i_13_327_1947_0, i_13_327_2022_0,
    i_13_327_2122_0, i_13_327_2199_0, i_13_327_2311_0, i_13_327_2427_0,
    i_13_327_2428_0, i_13_327_2454_0, i_13_327_2472_0, i_13_327_2473_0,
    i_13_327_2506_0, i_13_327_2517_0, i_13_327_2742_0, i_13_327_2743_0,
    i_13_327_2770_0, i_13_327_2940_0, i_13_327_2968_0, i_13_327_3009_0,
    i_13_327_3012_0, i_13_327_3030_0, i_13_327_3031_0, i_13_327_3075_0,
    i_13_327_3076_0, i_13_327_3091_0, i_13_327_3093_0, i_13_327_3211_0,
    i_13_327_3264_0, i_13_327_3273_0, i_13_327_3292_0, i_13_327_3345_0,
    i_13_327_3354_0, i_13_327_3381_0, i_13_327_3382_0, i_13_327_3418_0,
    i_13_327_3435_0, i_13_327_3540_0, i_13_327_3576_0, i_13_327_3759_0,
    i_13_327_3822_0, i_13_327_3900_0, i_13_327_3929_0, i_13_327_4036_0,
    i_13_327_4083_0, i_13_327_4164_0, i_13_327_4272_0, i_13_327_4362_0,
    i_13_327_4450_0, i_13_327_4497_0, i_13_327_4605_0, i_13_327_4606_0;
  output o_13_327_0_0;
  assign o_13_327_0_0 = ~((~i_13_327_1150_0 & ((~i_13_327_48_0 & ~i_13_327_1923_0) | (i_13_327_1596_0 & i_13_327_2427_0))) | (~i_13_327_1798_0 & ((~i_13_327_285_0 & ~i_13_327_1402_0 & ~i_13_327_1770_0 & ~i_13_327_1947_0) | (~i_13_327_2022_0 & ~i_13_327_2454_0 & ~i_13_327_3576_0 & i_13_327_4036_0))) | (~i_13_327_4036_0 & (i_13_327_1794_0 | (~i_13_327_2743_0 & i_13_327_4272_0))) | (i_13_327_1922_0 & ~i_13_327_4450_0));
endmodule



// Benchmark "kernel_13_328" written by ABC on Sun Jul 19 10:49:56 2020

module kernel_13_328 ( 
    i_13_328_18_0, i_13_328_58_0, i_13_328_102_0, i_13_328_130_0,
    i_13_328_131_0, i_13_328_132_0, i_13_328_223_0, i_13_328_355_0,
    i_13_328_371_0, i_13_328_374_0, i_13_328_415_0, i_13_328_489_0,
    i_13_328_614_0, i_13_328_736_0, i_13_328_955_0, i_13_328_956_0,
    i_13_328_1084_0, i_13_328_1100_0, i_13_328_1128_0, i_13_328_1227_0,
    i_13_328_1256_0, i_13_328_1300_0, i_13_328_1302_0, i_13_328_1305_0,
    i_13_328_1306_0, i_13_328_1322_0, i_13_328_1409_0, i_13_328_1445_0,
    i_13_328_1451_0, i_13_328_1472_0, i_13_328_1494_0, i_13_328_1503_0,
    i_13_328_1517_0, i_13_328_1522_0, i_13_328_1551_0, i_13_328_1552_0,
    i_13_328_1553_0, i_13_328_1554_0, i_13_328_1638_0, i_13_328_1639_0,
    i_13_328_1736_0, i_13_328_1778_0, i_13_328_1801_0, i_13_328_1802_0,
    i_13_328_1814_0, i_13_328_1846_0, i_13_328_1957_0, i_13_328_2090_0,
    i_13_328_2093_0, i_13_328_2100_0, i_13_328_2101_0, i_13_328_2142_0,
    i_13_328_2199_0, i_13_328_2235_0, i_13_328_2236_0, i_13_328_2296_0,
    i_13_328_2297_0, i_13_328_2522_0, i_13_328_2744_0, i_13_328_2789_0,
    i_13_328_2821_0, i_13_328_2822_0, i_13_328_2935_0, i_13_328_2936_0,
    i_13_328_2997_0, i_13_328_3024_0, i_13_328_3064_0, i_13_328_3100_0,
    i_13_328_3119_0, i_13_328_3145_0, i_13_328_3206_0, i_13_328_3241_0,
    i_13_328_3242_0, i_13_328_3308_0, i_13_328_3383_0, i_13_328_3388_0,
    i_13_328_3420_0, i_13_328_3433_0, i_13_328_3451_0, i_13_328_3477_0,
    i_13_328_3523_0, i_13_328_3537_0, i_13_328_3539_0, i_13_328_3617_0,
    i_13_328_3638_0, i_13_328_3685_0, i_13_328_3686_0, i_13_328_3754_0,
    i_13_328_3855_0, i_13_328_3856_0, i_13_328_3857_0, i_13_328_3916_0,
    i_13_328_4018_0, i_13_328_4060_0, i_13_328_4311_0, i_13_328_4312_0,
    i_13_328_4378_0, i_13_328_4382_0, i_13_328_4509_0, i_13_328_4592_0,
    o_13_328_0_0  );
  input  i_13_328_18_0, i_13_328_58_0, i_13_328_102_0, i_13_328_130_0,
    i_13_328_131_0, i_13_328_132_0, i_13_328_223_0, i_13_328_355_0,
    i_13_328_371_0, i_13_328_374_0, i_13_328_415_0, i_13_328_489_0,
    i_13_328_614_0, i_13_328_736_0, i_13_328_955_0, i_13_328_956_0,
    i_13_328_1084_0, i_13_328_1100_0, i_13_328_1128_0, i_13_328_1227_0,
    i_13_328_1256_0, i_13_328_1300_0, i_13_328_1302_0, i_13_328_1305_0,
    i_13_328_1306_0, i_13_328_1322_0, i_13_328_1409_0, i_13_328_1445_0,
    i_13_328_1451_0, i_13_328_1472_0, i_13_328_1494_0, i_13_328_1503_0,
    i_13_328_1517_0, i_13_328_1522_0, i_13_328_1551_0, i_13_328_1552_0,
    i_13_328_1553_0, i_13_328_1554_0, i_13_328_1638_0, i_13_328_1639_0,
    i_13_328_1736_0, i_13_328_1778_0, i_13_328_1801_0, i_13_328_1802_0,
    i_13_328_1814_0, i_13_328_1846_0, i_13_328_1957_0, i_13_328_2090_0,
    i_13_328_2093_0, i_13_328_2100_0, i_13_328_2101_0, i_13_328_2142_0,
    i_13_328_2199_0, i_13_328_2235_0, i_13_328_2236_0, i_13_328_2296_0,
    i_13_328_2297_0, i_13_328_2522_0, i_13_328_2744_0, i_13_328_2789_0,
    i_13_328_2821_0, i_13_328_2822_0, i_13_328_2935_0, i_13_328_2936_0,
    i_13_328_2997_0, i_13_328_3024_0, i_13_328_3064_0, i_13_328_3100_0,
    i_13_328_3119_0, i_13_328_3145_0, i_13_328_3206_0, i_13_328_3241_0,
    i_13_328_3242_0, i_13_328_3308_0, i_13_328_3383_0, i_13_328_3388_0,
    i_13_328_3420_0, i_13_328_3433_0, i_13_328_3451_0, i_13_328_3477_0,
    i_13_328_3523_0, i_13_328_3537_0, i_13_328_3539_0, i_13_328_3617_0,
    i_13_328_3638_0, i_13_328_3685_0, i_13_328_3686_0, i_13_328_3754_0,
    i_13_328_3855_0, i_13_328_3856_0, i_13_328_3857_0, i_13_328_3916_0,
    i_13_328_4018_0, i_13_328_4060_0, i_13_328_4311_0, i_13_328_4312_0,
    i_13_328_4378_0, i_13_328_4382_0, i_13_328_4509_0, i_13_328_4592_0;
  output o_13_328_0_0;
  assign o_13_328_0_0 = ~((~i_13_328_1639_0 & ((~i_13_328_1472_0 & ~i_13_328_3451_0) | (i_13_328_3145_0 & ~i_13_328_4312_0))) | (~i_13_328_1409_0 & i_13_328_3617_0) | (~i_13_328_1451_0 & ~i_13_328_1846_0 & ~i_13_328_3206_0 & i_13_328_3685_0) | (~i_13_328_1256_0 & ~i_13_328_1553_0 & ~i_13_328_3539_0 & ~i_13_328_3855_0 & ~i_13_328_4311_0) | (i_13_328_736_0 & ~i_13_328_4378_0) | (~i_13_328_1778_0 & ~i_13_328_3523_0 & ~i_13_328_3916_0 & ~i_13_328_4382_0) | (~i_13_328_1552_0 & ~i_13_328_3754_0 & ~i_13_328_3856_0 & ~i_13_328_4509_0));
endmodule



// Benchmark "kernel_13_329" written by ABC on Sun Jul 19 10:49:57 2020

module kernel_13_329 ( 
    i_13_329_45_0, i_13_329_46_0, i_13_329_169_0, i_13_329_175_0,
    i_13_329_179_0, i_13_329_187_0, i_13_329_283_0, i_13_329_310_0,
    i_13_329_343_0, i_13_329_444_0, i_13_329_515_0, i_13_329_532_0,
    i_13_329_554_0, i_13_329_567_0, i_13_329_568_0, i_13_329_574_0,
    i_13_329_649_0, i_13_329_719_0, i_13_329_730_0, i_13_329_847_0,
    i_13_329_854_0, i_13_329_886_0, i_13_329_986_0, i_13_329_1037_0,
    i_13_329_1072_0, i_13_329_1105_0, i_13_329_1228_0, i_13_329_1232_0,
    i_13_329_1309_0, i_13_329_1316_0, i_13_329_1550_0, i_13_329_1729_0,
    i_13_329_1741_0, i_13_329_1765_0, i_13_329_1804_0, i_13_329_1805_0,
    i_13_329_1822_0, i_13_329_1832_0, i_13_329_1846_0, i_13_329_1850_0,
    i_13_329_1852_0, i_13_329_1895_0, i_13_329_1992_0, i_13_329_1996_0,
    i_13_329_2020_0, i_13_329_2288_0, i_13_329_2314_0, i_13_329_2365_0,
    i_13_329_2372_0, i_13_329_2408_0, i_13_329_2422_0, i_13_329_2434_0,
    i_13_329_2443_0, i_13_329_2449_0, i_13_329_2450_0, i_13_329_2470_0,
    i_13_329_2473_0, i_13_329_2479_0, i_13_329_2680_0, i_13_329_2681_0,
    i_13_329_2897_0, i_13_329_3010_0, i_13_329_3011_0, i_13_329_3032_0,
    i_13_329_3110_0, i_13_329_3168_0, i_13_329_3207_0, i_13_329_3208_0,
    i_13_329_3212_0, i_13_329_3272_0, i_13_329_3400_0, i_13_329_3420_0,
    i_13_329_3421_0, i_13_329_3483_0, i_13_329_3502_0, i_13_329_3578_0,
    i_13_329_3637_0, i_13_329_3748_0, i_13_329_3871_0, i_13_329_3872_0,
    i_13_329_3907_0, i_13_329_3914_0, i_13_329_3955_0, i_13_329_4015_0,
    i_13_329_4036_0, i_13_329_4041_0, i_13_329_4042_0, i_13_329_4095_0,
    i_13_329_4190_0, i_13_329_4248_0, i_13_329_4252_0, i_13_329_4253_0,
    i_13_329_4270_0, i_13_329_4368_0, i_13_329_4369_0, i_13_329_4374_0,
    i_13_329_4379_0, i_13_329_4441_0, i_13_329_4514_0, i_13_329_4607_0,
    o_13_329_0_0  );
  input  i_13_329_45_0, i_13_329_46_0, i_13_329_169_0, i_13_329_175_0,
    i_13_329_179_0, i_13_329_187_0, i_13_329_283_0, i_13_329_310_0,
    i_13_329_343_0, i_13_329_444_0, i_13_329_515_0, i_13_329_532_0,
    i_13_329_554_0, i_13_329_567_0, i_13_329_568_0, i_13_329_574_0,
    i_13_329_649_0, i_13_329_719_0, i_13_329_730_0, i_13_329_847_0,
    i_13_329_854_0, i_13_329_886_0, i_13_329_986_0, i_13_329_1037_0,
    i_13_329_1072_0, i_13_329_1105_0, i_13_329_1228_0, i_13_329_1232_0,
    i_13_329_1309_0, i_13_329_1316_0, i_13_329_1550_0, i_13_329_1729_0,
    i_13_329_1741_0, i_13_329_1765_0, i_13_329_1804_0, i_13_329_1805_0,
    i_13_329_1822_0, i_13_329_1832_0, i_13_329_1846_0, i_13_329_1850_0,
    i_13_329_1852_0, i_13_329_1895_0, i_13_329_1992_0, i_13_329_1996_0,
    i_13_329_2020_0, i_13_329_2288_0, i_13_329_2314_0, i_13_329_2365_0,
    i_13_329_2372_0, i_13_329_2408_0, i_13_329_2422_0, i_13_329_2434_0,
    i_13_329_2443_0, i_13_329_2449_0, i_13_329_2450_0, i_13_329_2470_0,
    i_13_329_2473_0, i_13_329_2479_0, i_13_329_2680_0, i_13_329_2681_0,
    i_13_329_2897_0, i_13_329_3010_0, i_13_329_3011_0, i_13_329_3032_0,
    i_13_329_3110_0, i_13_329_3168_0, i_13_329_3207_0, i_13_329_3208_0,
    i_13_329_3212_0, i_13_329_3272_0, i_13_329_3400_0, i_13_329_3420_0,
    i_13_329_3421_0, i_13_329_3483_0, i_13_329_3502_0, i_13_329_3578_0,
    i_13_329_3637_0, i_13_329_3748_0, i_13_329_3871_0, i_13_329_3872_0,
    i_13_329_3907_0, i_13_329_3914_0, i_13_329_3955_0, i_13_329_4015_0,
    i_13_329_4036_0, i_13_329_4041_0, i_13_329_4042_0, i_13_329_4095_0,
    i_13_329_4190_0, i_13_329_4248_0, i_13_329_4252_0, i_13_329_4253_0,
    i_13_329_4270_0, i_13_329_4368_0, i_13_329_4369_0, i_13_329_4374_0,
    i_13_329_4379_0, i_13_329_4441_0, i_13_329_4514_0, i_13_329_4607_0;
  output o_13_329_0_0;
  assign o_13_329_0_0 = 0;
endmodule



// Benchmark "kernel_13_330" written by ABC on Sun Jul 19 10:49:58 2020

module kernel_13_330 ( 
    i_13_330_50_0, i_13_330_80_0, i_13_330_201_0, i_13_330_203_0,
    i_13_330_229_0, i_13_330_286_0, i_13_330_421_0, i_13_330_535_0,
    i_13_330_626_0, i_13_330_661_0, i_13_330_792_0, i_13_330_823_0,
    i_13_330_847_0, i_13_330_850_0, i_13_330_851_0, i_13_330_867_0,
    i_13_330_869_0, i_13_330_941_0, i_13_330_1018_0, i_13_330_1021_0,
    i_13_330_1022_0, i_13_330_1060_0, i_13_330_1075_0, i_13_330_1076_0,
    i_13_330_1232_0, i_13_330_1318_0, i_13_330_1427_0, i_13_330_1530_0,
    i_13_330_1541_0, i_13_330_1549_0, i_13_330_1550_0, i_13_330_1551_0,
    i_13_330_1598_0, i_13_330_1679_0, i_13_330_1774_0, i_13_330_1780_0,
    i_13_330_1855_0, i_13_330_1858_0, i_13_330_2030_0, i_13_330_2197_0,
    i_13_330_2199_0, i_13_330_2200_0, i_13_330_2202_0, i_13_330_2452_0,
    i_13_330_2539_0, i_13_330_2543_0, i_13_330_2617_0, i_13_330_2703_0,
    i_13_330_2913_0, i_13_330_2920_0, i_13_330_2999_0, i_13_330_3007_0,
    i_13_330_3010_0, i_13_330_3011_0, i_13_330_3013_0, i_13_330_3064_0,
    i_13_330_3087_0, i_13_330_3104_0, i_13_330_3169_0, i_13_330_3172_0,
    i_13_330_3399_0, i_13_330_3453_0, i_13_330_3454_0, i_13_330_3461_0,
    i_13_330_3484_0, i_13_330_3486_0, i_13_330_3487_0, i_13_330_3488_0,
    i_13_330_3535_0, i_13_330_3539_0, i_13_330_3541_0, i_13_330_3542_0,
    i_13_330_3576_0, i_13_330_3577_0, i_13_330_3578_0, i_13_330_3616_0,
    i_13_330_3703_0, i_13_330_3730_0, i_13_330_3764_0, i_13_330_3781_0,
    i_13_330_3782_0, i_13_330_3784_0, i_13_330_3785_0, i_13_330_3854_0,
    i_13_330_3865_0, i_13_330_3866_0, i_13_330_3868_0, i_13_330_3885_0,
    i_13_330_3889_0, i_13_330_3892_0, i_13_330_3906_0, i_13_330_4176_0,
    i_13_330_4179_0, i_13_330_4249_0, i_13_330_4252_0, i_13_330_4256_0,
    i_13_330_4262_0, i_13_330_4378_0, i_13_330_4379_0, i_13_330_4561_0,
    o_13_330_0_0  );
  input  i_13_330_50_0, i_13_330_80_0, i_13_330_201_0, i_13_330_203_0,
    i_13_330_229_0, i_13_330_286_0, i_13_330_421_0, i_13_330_535_0,
    i_13_330_626_0, i_13_330_661_0, i_13_330_792_0, i_13_330_823_0,
    i_13_330_847_0, i_13_330_850_0, i_13_330_851_0, i_13_330_867_0,
    i_13_330_869_0, i_13_330_941_0, i_13_330_1018_0, i_13_330_1021_0,
    i_13_330_1022_0, i_13_330_1060_0, i_13_330_1075_0, i_13_330_1076_0,
    i_13_330_1232_0, i_13_330_1318_0, i_13_330_1427_0, i_13_330_1530_0,
    i_13_330_1541_0, i_13_330_1549_0, i_13_330_1550_0, i_13_330_1551_0,
    i_13_330_1598_0, i_13_330_1679_0, i_13_330_1774_0, i_13_330_1780_0,
    i_13_330_1855_0, i_13_330_1858_0, i_13_330_2030_0, i_13_330_2197_0,
    i_13_330_2199_0, i_13_330_2200_0, i_13_330_2202_0, i_13_330_2452_0,
    i_13_330_2539_0, i_13_330_2543_0, i_13_330_2617_0, i_13_330_2703_0,
    i_13_330_2913_0, i_13_330_2920_0, i_13_330_2999_0, i_13_330_3007_0,
    i_13_330_3010_0, i_13_330_3011_0, i_13_330_3013_0, i_13_330_3064_0,
    i_13_330_3087_0, i_13_330_3104_0, i_13_330_3169_0, i_13_330_3172_0,
    i_13_330_3399_0, i_13_330_3453_0, i_13_330_3454_0, i_13_330_3461_0,
    i_13_330_3484_0, i_13_330_3486_0, i_13_330_3487_0, i_13_330_3488_0,
    i_13_330_3535_0, i_13_330_3539_0, i_13_330_3541_0, i_13_330_3542_0,
    i_13_330_3576_0, i_13_330_3577_0, i_13_330_3578_0, i_13_330_3616_0,
    i_13_330_3703_0, i_13_330_3730_0, i_13_330_3764_0, i_13_330_3781_0,
    i_13_330_3782_0, i_13_330_3784_0, i_13_330_3785_0, i_13_330_3854_0,
    i_13_330_3865_0, i_13_330_3866_0, i_13_330_3868_0, i_13_330_3885_0,
    i_13_330_3889_0, i_13_330_3892_0, i_13_330_3906_0, i_13_330_4176_0,
    i_13_330_4179_0, i_13_330_4249_0, i_13_330_4252_0, i_13_330_4256_0,
    i_13_330_4262_0, i_13_330_4378_0, i_13_330_4379_0, i_13_330_4561_0;
  output o_13_330_0_0;
  assign o_13_330_0_0 = ~((~i_13_330_4561_0 & ((~i_13_330_1318_0 & ~i_13_330_3487_0) | (~i_13_330_3011_0 & ~i_13_330_3488_0 & ~i_13_330_4252_0))) | (~i_13_330_2617_0 & i_13_330_3453_0) | (~i_13_330_1021_0 & i_13_330_3865_0 & i_13_330_3906_0) | (~i_13_330_1858_0 & ~i_13_330_3007_0 & ~i_13_330_3782_0 & ~i_13_330_3868_0 & ~i_13_330_3892_0 & ~i_13_330_4262_0) | (i_13_330_535_0 & ~i_13_330_3781_0 & i_13_330_4378_0) | (~i_13_330_3461_0 & ~i_13_330_3539_0 & ~i_13_330_3577_0 & ~i_13_330_4379_0));
endmodule



// Benchmark "kernel_13_331" written by ABC on Sun Jul 19 10:49:59 2020

module kernel_13_331 ( 
    i_13_331_28_0, i_13_331_29_0, i_13_331_31_0, i_13_331_32_0,
    i_13_331_64_0, i_13_331_65_0, i_13_331_91_0, i_13_331_136_0,
    i_13_331_137_0, i_13_331_184_0, i_13_331_226_0, i_13_331_227_0,
    i_13_331_228_0, i_13_331_307_0, i_13_331_308_0, i_13_331_309_0,
    i_13_331_316_0, i_13_331_317_0, i_13_331_380_0, i_13_331_418_0,
    i_13_331_419_0, i_13_331_459_0, i_13_331_535_0, i_13_331_553_0,
    i_13_331_639_0, i_13_331_718_0, i_13_331_873_0, i_13_331_950_0,
    i_13_331_1075_0, i_13_331_1143_0, i_13_331_1208_0, i_13_331_1216_0,
    i_13_331_1217_0, i_13_331_1308_0, i_13_331_1318_0, i_13_331_1341_0,
    i_13_331_1408_0, i_13_331_1422_0, i_13_331_1435_0, i_13_331_1445_0,
    i_13_331_1526_0, i_13_331_1594_0, i_13_331_1596_0, i_13_331_1678_0,
    i_13_331_1720_0, i_13_331_1785_0, i_13_331_1841_0, i_13_331_1848_0,
    i_13_331_1858_0, i_13_331_1922_0, i_13_331_1999_0, i_13_331_2000_0,
    i_13_331_2002_0, i_13_331_2003_0, i_13_331_2052_0, i_13_331_2055_0,
    i_13_331_2142_0, i_13_331_2146_0, i_13_331_2174_0, i_13_331_2189_0,
    i_13_331_2259_0, i_13_331_2280_0, i_13_331_2345_0, i_13_331_2403_0,
    i_13_331_2422_0, i_13_331_2423_0, i_13_331_2547_0, i_13_331_2552_0,
    i_13_331_2674_0, i_13_331_2694_0, i_13_331_2710_0, i_13_331_2719_0,
    i_13_331_2720_0, i_13_331_2740_0, i_13_331_2854_0, i_13_331_2855_0,
    i_13_331_2857_0, i_13_331_2884_0, i_13_331_2937_0, i_13_331_3034_0,
    i_13_331_3036_0, i_13_331_3127_0, i_13_331_3204_0, i_13_331_3207_0,
    i_13_331_3366_0, i_13_331_3487_0, i_13_331_3523_0, i_13_331_3529_0,
    i_13_331_3663_0, i_13_331_3727_0, i_13_331_3764_0, i_13_331_3902_0,
    i_13_331_3990_0, i_13_331_4034_0, i_13_331_4036_0, i_13_331_4082_0,
    i_13_331_4349_0, i_13_331_4351_0, i_13_331_4397_0, i_13_331_4514_0,
    o_13_331_0_0  );
  input  i_13_331_28_0, i_13_331_29_0, i_13_331_31_0, i_13_331_32_0,
    i_13_331_64_0, i_13_331_65_0, i_13_331_91_0, i_13_331_136_0,
    i_13_331_137_0, i_13_331_184_0, i_13_331_226_0, i_13_331_227_0,
    i_13_331_228_0, i_13_331_307_0, i_13_331_308_0, i_13_331_309_0,
    i_13_331_316_0, i_13_331_317_0, i_13_331_380_0, i_13_331_418_0,
    i_13_331_419_0, i_13_331_459_0, i_13_331_535_0, i_13_331_553_0,
    i_13_331_639_0, i_13_331_718_0, i_13_331_873_0, i_13_331_950_0,
    i_13_331_1075_0, i_13_331_1143_0, i_13_331_1208_0, i_13_331_1216_0,
    i_13_331_1217_0, i_13_331_1308_0, i_13_331_1318_0, i_13_331_1341_0,
    i_13_331_1408_0, i_13_331_1422_0, i_13_331_1435_0, i_13_331_1445_0,
    i_13_331_1526_0, i_13_331_1594_0, i_13_331_1596_0, i_13_331_1678_0,
    i_13_331_1720_0, i_13_331_1785_0, i_13_331_1841_0, i_13_331_1848_0,
    i_13_331_1858_0, i_13_331_1922_0, i_13_331_1999_0, i_13_331_2000_0,
    i_13_331_2002_0, i_13_331_2003_0, i_13_331_2052_0, i_13_331_2055_0,
    i_13_331_2142_0, i_13_331_2146_0, i_13_331_2174_0, i_13_331_2189_0,
    i_13_331_2259_0, i_13_331_2280_0, i_13_331_2345_0, i_13_331_2403_0,
    i_13_331_2422_0, i_13_331_2423_0, i_13_331_2547_0, i_13_331_2552_0,
    i_13_331_2674_0, i_13_331_2694_0, i_13_331_2710_0, i_13_331_2719_0,
    i_13_331_2720_0, i_13_331_2740_0, i_13_331_2854_0, i_13_331_2855_0,
    i_13_331_2857_0, i_13_331_2884_0, i_13_331_2937_0, i_13_331_3034_0,
    i_13_331_3036_0, i_13_331_3127_0, i_13_331_3204_0, i_13_331_3207_0,
    i_13_331_3366_0, i_13_331_3487_0, i_13_331_3523_0, i_13_331_3529_0,
    i_13_331_3663_0, i_13_331_3727_0, i_13_331_3764_0, i_13_331_3902_0,
    i_13_331_3990_0, i_13_331_4034_0, i_13_331_4036_0, i_13_331_4082_0,
    i_13_331_4349_0, i_13_331_4351_0, i_13_331_4397_0, i_13_331_4514_0;
  output o_13_331_0_0;
  assign o_13_331_0_0 = ~((~i_13_331_316_0 & i_13_331_3036_0) | (~i_13_331_65_0 & ~i_13_331_1216_0) | (~i_13_331_32_0 & ~i_13_331_380_0 & ~i_13_331_1848_0 & i_13_331_2710_0));
endmodule



// Benchmark "kernel_13_332" written by ABC on Sun Jul 19 10:49:59 2020

module kernel_13_332 ( 
    i_13_332_16_0, i_13_332_40_0, i_13_332_119_0, i_13_332_138_0,
    i_13_332_139_0, i_13_332_141_0, i_13_332_225_0, i_13_332_231_0,
    i_13_332_273_0, i_13_332_369_0, i_13_332_431_0, i_13_332_447_0,
    i_13_332_469_0, i_13_332_537_0, i_13_332_613_0, i_13_332_646_0,
    i_13_332_690_0, i_13_332_691_0, i_13_332_717_0, i_13_332_727_0,
    i_13_332_760_0, i_13_332_780_0, i_13_332_811_0, i_13_332_894_0,
    i_13_332_940_0, i_13_332_984_0, i_13_332_1092_0, i_13_332_1203_0,
    i_13_332_1221_0, i_13_332_1249_0, i_13_332_1251_0, i_13_332_1260_0,
    i_13_332_1276_0, i_13_332_1299_0, i_13_332_1383_0, i_13_332_1386_0,
    i_13_332_1393_0, i_13_332_1464_0, i_13_332_1470_0, i_13_332_1567_0,
    i_13_332_1642_0, i_13_332_1671_0, i_13_332_1672_0, i_13_332_1713_0,
    i_13_332_1725_0, i_13_332_1726_0, i_13_332_1731_0, i_13_332_1884_0,
    i_13_332_1885_0, i_13_332_1887_0, i_13_332_1906_0, i_13_332_1990_0,
    i_13_332_1996_0, i_13_332_2136_0, i_13_332_2139_0, i_13_332_2167_0,
    i_13_332_2187_0, i_13_332_2464_0, i_13_332_2470_0, i_13_332_2577_0,
    i_13_332_2632_0, i_13_332_2649_0, i_13_332_2650_0, i_13_332_2652_0,
    i_13_332_2653_0, i_13_332_2680_0, i_13_332_2709_0, i_13_332_2755_0,
    i_13_332_2847_0, i_13_332_2877_0, i_13_332_2884_0, i_13_332_2914_0,
    i_13_332_3009_0, i_13_332_3108_0, i_13_332_3174_0, i_13_332_3219_0,
    i_13_332_3273_0, i_13_332_3279_0, i_13_332_3387_0, i_13_332_3391_0,
    i_13_332_3432_0, i_13_332_3474_0, i_13_332_3487_0, i_13_332_3528_0,
    i_13_332_3532_0, i_13_332_3682_0, i_13_332_3766_0, i_13_332_3793_0,
    i_13_332_3801_0, i_13_332_3838_0, i_13_332_3874_0, i_13_332_3906_0,
    i_13_332_4126_0, i_13_332_4156_0, i_13_332_4162_0, i_13_332_4308_0,
    i_13_332_4371_0, i_13_332_4443_0, i_13_332_4521_0, i_13_332_4533_0,
    o_13_332_0_0  );
  input  i_13_332_16_0, i_13_332_40_0, i_13_332_119_0, i_13_332_138_0,
    i_13_332_139_0, i_13_332_141_0, i_13_332_225_0, i_13_332_231_0,
    i_13_332_273_0, i_13_332_369_0, i_13_332_431_0, i_13_332_447_0,
    i_13_332_469_0, i_13_332_537_0, i_13_332_613_0, i_13_332_646_0,
    i_13_332_690_0, i_13_332_691_0, i_13_332_717_0, i_13_332_727_0,
    i_13_332_760_0, i_13_332_780_0, i_13_332_811_0, i_13_332_894_0,
    i_13_332_940_0, i_13_332_984_0, i_13_332_1092_0, i_13_332_1203_0,
    i_13_332_1221_0, i_13_332_1249_0, i_13_332_1251_0, i_13_332_1260_0,
    i_13_332_1276_0, i_13_332_1299_0, i_13_332_1383_0, i_13_332_1386_0,
    i_13_332_1393_0, i_13_332_1464_0, i_13_332_1470_0, i_13_332_1567_0,
    i_13_332_1642_0, i_13_332_1671_0, i_13_332_1672_0, i_13_332_1713_0,
    i_13_332_1725_0, i_13_332_1726_0, i_13_332_1731_0, i_13_332_1884_0,
    i_13_332_1885_0, i_13_332_1887_0, i_13_332_1906_0, i_13_332_1990_0,
    i_13_332_1996_0, i_13_332_2136_0, i_13_332_2139_0, i_13_332_2167_0,
    i_13_332_2187_0, i_13_332_2464_0, i_13_332_2470_0, i_13_332_2577_0,
    i_13_332_2632_0, i_13_332_2649_0, i_13_332_2650_0, i_13_332_2652_0,
    i_13_332_2653_0, i_13_332_2680_0, i_13_332_2709_0, i_13_332_2755_0,
    i_13_332_2847_0, i_13_332_2877_0, i_13_332_2884_0, i_13_332_2914_0,
    i_13_332_3009_0, i_13_332_3108_0, i_13_332_3174_0, i_13_332_3219_0,
    i_13_332_3273_0, i_13_332_3279_0, i_13_332_3387_0, i_13_332_3391_0,
    i_13_332_3432_0, i_13_332_3474_0, i_13_332_3487_0, i_13_332_3528_0,
    i_13_332_3532_0, i_13_332_3682_0, i_13_332_3766_0, i_13_332_3793_0,
    i_13_332_3801_0, i_13_332_3838_0, i_13_332_3874_0, i_13_332_3906_0,
    i_13_332_4126_0, i_13_332_4156_0, i_13_332_4162_0, i_13_332_4308_0,
    i_13_332_4371_0, i_13_332_4443_0, i_13_332_4521_0, i_13_332_4533_0;
  output o_13_332_0_0;
  assign o_13_332_0_0 = ~((~i_13_332_1713_0 & (~i_13_332_894_0 | (~i_13_332_3219_0 & ~i_13_332_3874_0))) | (~i_13_332_2650_0 & i_13_332_3528_0 & ~i_13_332_3682_0));
endmodule



// Benchmark "kernel_13_333" written by ABC on Sun Jul 19 10:50:00 2020

module kernel_13_333 ( 
    i_13_333_34_0, i_13_333_35_0, i_13_333_74_0, i_13_333_104_0,
    i_13_333_117_0, i_13_333_118_0, i_13_333_122_0, i_13_333_137_0,
    i_13_333_139_0, i_13_333_175_0, i_13_333_190_0, i_13_333_226_0,
    i_13_333_227_0, i_13_333_374_0, i_13_333_377_0, i_13_333_460_0,
    i_13_333_463_0, i_13_333_490_0, i_13_333_526_0, i_13_333_527_0,
    i_13_333_533_0, i_13_333_535_0, i_13_333_536_0, i_13_333_617_0,
    i_13_333_667_0, i_13_333_715_0, i_13_333_895_0, i_13_333_946_0,
    i_13_333_1084_0, i_13_333_1093_0, i_13_333_1094_0, i_13_333_1313_0,
    i_13_333_1444_0, i_13_333_1471_0, i_13_333_1597_0, i_13_333_1621_0,
    i_13_333_1684_0, i_13_333_1720_0, i_13_333_1721_0, i_13_333_1724_0,
    i_13_333_1784_0, i_13_333_1786_0, i_13_333_1787_0, i_13_333_1838_0,
    i_13_333_1841_0, i_13_333_1844_0, i_13_333_1849_0, i_13_333_1931_0,
    i_13_333_2056_0, i_13_333_2120_0, i_13_333_2177_0, i_13_333_2197_0,
    i_13_333_2263_0, i_13_333_2345_0, i_13_333_2459_0, i_13_333_2501_0,
    i_13_333_2611_0, i_13_333_2705_0, i_13_333_2714_0, i_13_333_2872_0,
    i_13_333_3010_0, i_13_333_3034_0, i_13_333_3037_0, i_13_333_3044_0,
    i_13_333_3047_0, i_13_333_3101_0, i_13_333_3159_0, i_13_333_3161_0,
    i_13_333_3162_0, i_13_333_3163_0, i_13_333_3164_0, i_13_333_3275_0,
    i_13_333_3326_0, i_13_333_3353_0, i_13_333_3376_0, i_13_333_3407_0,
    i_13_333_3449_0, i_13_333_3524_0, i_13_333_3539_0, i_13_333_3653_0,
    i_13_333_3685_0, i_13_333_3731_0, i_13_333_3737_0, i_13_333_3740_0,
    i_13_333_3857_0, i_13_333_3917_0, i_13_333_3919_0, i_13_333_3982_0,
    i_13_333_4106_0, i_13_333_4234_0, i_13_333_4235_0, i_13_333_4258_0,
    i_13_333_4316_0, i_13_333_4325_0, i_13_333_4414_0, i_13_333_4415_0,
    i_13_333_4492_0, i_13_333_4519_0, i_13_333_4540_0, i_13_333_4541_0,
    o_13_333_0_0  );
  input  i_13_333_34_0, i_13_333_35_0, i_13_333_74_0, i_13_333_104_0,
    i_13_333_117_0, i_13_333_118_0, i_13_333_122_0, i_13_333_137_0,
    i_13_333_139_0, i_13_333_175_0, i_13_333_190_0, i_13_333_226_0,
    i_13_333_227_0, i_13_333_374_0, i_13_333_377_0, i_13_333_460_0,
    i_13_333_463_0, i_13_333_490_0, i_13_333_526_0, i_13_333_527_0,
    i_13_333_533_0, i_13_333_535_0, i_13_333_536_0, i_13_333_617_0,
    i_13_333_667_0, i_13_333_715_0, i_13_333_895_0, i_13_333_946_0,
    i_13_333_1084_0, i_13_333_1093_0, i_13_333_1094_0, i_13_333_1313_0,
    i_13_333_1444_0, i_13_333_1471_0, i_13_333_1597_0, i_13_333_1621_0,
    i_13_333_1684_0, i_13_333_1720_0, i_13_333_1721_0, i_13_333_1724_0,
    i_13_333_1784_0, i_13_333_1786_0, i_13_333_1787_0, i_13_333_1838_0,
    i_13_333_1841_0, i_13_333_1844_0, i_13_333_1849_0, i_13_333_1931_0,
    i_13_333_2056_0, i_13_333_2120_0, i_13_333_2177_0, i_13_333_2197_0,
    i_13_333_2263_0, i_13_333_2345_0, i_13_333_2459_0, i_13_333_2501_0,
    i_13_333_2611_0, i_13_333_2705_0, i_13_333_2714_0, i_13_333_2872_0,
    i_13_333_3010_0, i_13_333_3034_0, i_13_333_3037_0, i_13_333_3044_0,
    i_13_333_3047_0, i_13_333_3101_0, i_13_333_3159_0, i_13_333_3161_0,
    i_13_333_3162_0, i_13_333_3163_0, i_13_333_3164_0, i_13_333_3275_0,
    i_13_333_3326_0, i_13_333_3353_0, i_13_333_3376_0, i_13_333_3407_0,
    i_13_333_3449_0, i_13_333_3524_0, i_13_333_3539_0, i_13_333_3653_0,
    i_13_333_3685_0, i_13_333_3731_0, i_13_333_3737_0, i_13_333_3740_0,
    i_13_333_3857_0, i_13_333_3917_0, i_13_333_3919_0, i_13_333_3982_0,
    i_13_333_4106_0, i_13_333_4234_0, i_13_333_4235_0, i_13_333_4258_0,
    i_13_333_4316_0, i_13_333_4325_0, i_13_333_4414_0, i_13_333_4415_0,
    i_13_333_4492_0, i_13_333_4519_0, i_13_333_4540_0, i_13_333_4541_0;
  output o_13_333_0_0;
  assign o_13_333_0_0 = ~((~i_13_333_139_0 & (~i_13_333_490_0 | (i_13_333_526_0 & ~i_13_333_1621_0 & ~i_13_333_4325_0))) | (~i_13_333_4415_0 & ((~i_13_333_1621_0 & ~i_13_333_1844_0 & ~i_13_333_3163_0) | (~i_13_333_3164_0 & i_13_333_3524_0))) | (i_13_333_463_0 & ~i_13_333_2056_0 & ~i_13_333_2714_0) | (~i_13_333_117_0 & ~i_13_333_227_0 & i_13_333_526_0 & ~i_13_333_3161_0) | (~i_13_333_226_0 & ~i_13_333_895_0 & ~i_13_333_3524_0) | (~i_13_333_1084_0 & i_13_333_3162_0 & ~i_13_333_3982_0));
endmodule



// Benchmark "kernel_13_334" written by ABC on Sun Jul 19 10:50:01 2020

module kernel_13_334 ( 
    i_13_334_41_0, i_13_334_274_0, i_13_334_283_0, i_13_334_284_0,
    i_13_334_383_0, i_13_334_422_0, i_13_334_454_0, i_13_334_529_0,
    i_13_334_553_0, i_13_334_554_0, i_13_334_558_0, i_13_334_565_0,
    i_13_334_599_0, i_13_334_607_0, i_13_334_666_0, i_13_334_820_0,
    i_13_334_821_0, i_13_334_896_0, i_13_334_1024_0, i_13_334_1099_0,
    i_13_334_1120_0, i_13_334_1147_0, i_13_334_1270_0, i_13_334_1314_0,
    i_13_334_1387_0, i_13_334_1433_0, i_13_334_1609_0, i_13_334_1635_0,
    i_13_334_1636_0, i_13_334_1637_0, i_13_334_1665_0, i_13_334_1687_0,
    i_13_334_1715_0, i_13_334_1716_0, i_13_334_1720_0, i_13_334_1732_0,
    i_13_334_1737_0, i_13_334_1774_0, i_13_334_1775_0, i_13_334_1788_0,
    i_13_334_1840_0, i_13_334_1859_0, i_13_334_1886_0, i_13_334_1960_0,
    i_13_334_1994_0, i_13_334_2005_0, i_13_334_2015_0, i_13_334_2121_0,
    i_13_334_2137_0, i_13_334_2302_0, i_13_334_2381_0, i_13_334_2459_0,
    i_13_334_2461_0, i_13_334_2462_0, i_13_334_2464_0, i_13_334_2493_0,
    i_13_334_2593_0, i_13_334_2630_0, i_13_334_2677_0, i_13_334_2678_0,
    i_13_334_2722_0, i_13_334_2839_0, i_13_334_2884_0, i_13_334_2983_0,
    i_13_334_3100_0, i_13_334_3172_0, i_13_334_3173_0, i_13_334_3175_0,
    i_13_334_3367_0, i_13_334_3448_0, i_13_334_3464_0, i_13_334_3545_0,
    i_13_334_3667_0, i_13_334_3730_0, i_13_334_3731_0, i_13_334_3733_0,
    i_13_334_3734_0, i_13_334_3787_0, i_13_334_3909_0, i_13_334_3910_0,
    i_13_334_3911_0, i_13_334_3913_0, i_13_334_3914_0, i_13_334_3931_0,
    i_13_334_4018_0, i_13_334_4091_0, i_13_334_4097_0, i_13_334_4162_0,
    i_13_334_4216_0, i_13_334_4255_0, i_13_334_4315_0, i_13_334_4351_0,
    i_13_334_4369_0, i_13_334_4372_0, i_13_334_4432_0, i_13_334_4514_0,
    i_13_334_4561_0, i_13_334_4568_0, i_13_334_4594_0, i_13_334_4603_0,
    o_13_334_0_0  );
  input  i_13_334_41_0, i_13_334_274_0, i_13_334_283_0, i_13_334_284_0,
    i_13_334_383_0, i_13_334_422_0, i_13_334_454_0, i_13_334_529_0,
    i_13_334_553_0, i_13_334_554_0, i_13_334_558_0, i_13_334_565_0,
    i_13_334_599_0, i_13_334_607_0, i_13_334_666_0, i_13_334_820_0,
    i_13_334_821_0, i_13_334_896_0, i_13_334_1024_0, i_13_334_1099_0,
    i_13_334_1120_0, i_13_334_1147_0, i_13_334_1270_0, i_13_334_1314_0,
    i_13_334_1387_0, i_13_334_1433_0, i_13_334_1609_0, i_13_334_1635_0,
    i_13_334_1636_0, i_13_334_1637_0, i_13_334_1665_0, i_13_334_1687_0,
    i_13_334_1715_0, i_13_334_1716_0, i_13_334_1720_0, i_13_334_1732_0,
    i_13_334_1737_0, i_13_334_1774_0, i_13_334_1775_0, i_13_334_1788_0,
    i_13_334_1840_0, i_13_334_1859_0, i_13_334_1886_0, i_13_334_1960_0,
    i_13_334_1994_0, i_13_334_2005_0, i_13_334_2015_0, i_13_334_2121_0,
    i_13_334_2137_0, i_13_334_2302_0, i_13_334_2381_0, i_13_334_2459_0,
    i_13_334_2461_0, i_13_334_2462_0, i_13_334_2464_0, i_13_334_2493_0,
    i_13_334_2593_0, i_13_334_2630_0, i_13_334_2677_0, i_13_334_2678_0,
    i_13_334_2722_0, i_13_334_2839_0, i_13_334_2884_0, i_13_334_2983_0,
    i_13_334_3100_0, i_13_334_3172_0, i_13_334_3173_0, i_13_334_3175_0,
    i_13_334_3367_0, i_13_334_3448_0, i_13_334_3464_0, i_13_334_3545_0,
    i_13_334_3667_0, i_13_334_3730_0, i_13_334_3731_0, i_13_334_3733_0,
    i_13_334_3734_0, i_13_334_3787_0, i_13_334_3909_0, i_13_334_3910_0,
    i_13_334_3911_0, i_13_334_3913_0, i_13_334_3914_0, i_13_334_3931_0,
    i_13_334_4018_0, i_13_334_4091_0, i_13_334_4097_0, i_13_334_4162_0,
    i_13_334_4216_0, i_13_334_4255_0, i_13_334_4315_0, i_13_334_4351_0,
    i_13_334_4369_0, i_13_334_4372_0, i_13_334_4432_0, i_13_334_4514_0,
    i_13_334_4561_0, i_13_334_4568_0, i_13_334_4594_0, i_13_334_4603_0;
  output o_13_334_0_0;
  assign o_13_334_0_0 = ~((~i_13_334_3175_0 & ((~i_13_334_821_0 & ~i_13_334_2464_0) | (~i_13_334_1775_0 & ~i_13_334_3914_0 & ~i_13_334_4091_0))) | (~i_13_334_565_0 & ~i_13_334_1609_0 & i_13_334_2983_0) | (~i_13_334_3911_0 & ~i_13_334_4315_0) | (i_13_334_1147_0 & i_13_334_4369_0) | (~i_13_334_3914_0 & ~i_13_334_4091_0 & ~i_13_334_4369_0 & ~i_13_334_4561_0));
endmodule



// Benchmark "kernel_13_335" written by ABC on Sun Jul 19 10:50:02 2020

module kernel_13_335 ( 
    i_13_335_77_0, i_13_335_92_0, i_13_335_203_0, i_13_335_259_0,
    i_13_335_265_0, i_13_335_266_0, i_13_335_353_0, i_13_335_374_0,
    i_13_335_382_0, i_13_335_413_0, i_13_335_451_0, i_13_335_520_0,
    i_13_335_569_0, i_13_335_605_0, i_13_335_607_0, i_13_335_608_0,
    i_13_335_658_0, i_13_335_661_0, i_13_335_670_0, i_13_335_671_0,
    i_13_335_680_0, i_13_335_929_0, i_13_335_940_0, i_13_335_943_0,
    i_13_335_950_0, i_13_335_1081_0, i_13_335_1082_0, i_13_335_1145_0,
    i_13_335_1148_0, i_13_335_1229_0, i_13_335_1300_0, i_13_335_1307_0,
    i_13_335_1385_0, i_13_335_1444_0, i_13_335_1454_0, i_13_335_1486_0,
    i_13_335_1663_0, i_13_335_1730_0, i_13_335_1733_0, i_13_335_1765_0,
    i_13_335_1766_0, i_13_335_1841_0, i_13_335_1865_0, i_13_335_1885_0,
    i_13_335_1892_0, i_13_335_1927_0, i_13_335_2020_0, i_13_335_2054_0,
    i_13_335_2137_0, i_13_335_2281_0, i_13_335_2300_0, i_13_335_2365_0,
    i_13_335_2423_0, i_13_335_2435_0, i_13_335_2468_0, i_13_335_2546_0,
    i_13_335_2570_0, i_13_335_2614_0, i_13_335_2615_0, i_13_335_2650_0,
    i_13_335_2858_0, i_13_335_2887_0, i_13_335_2980_0, i_13_335_3017_0,
    i_13_335_3047_0, i_13_335_3077_0, i_13_335_3142_0, i_13_335_3259_0,
    i_13_335_3269_0, i_13_335_3343_0, i_13_335_3359_0, i_13_335_3445_0,
    i_13_335_3449_0, i_13_335_3476_0, i_13_335_3484_0, i_13_335_3485_0,
    i_13_335_3646_0, i_13_335_3731_0, i_13_335_3764_0, i_13_335_3781_0,
    i_13_335_3872_0, i_13_335_3875_0, i_13_335_3979_0, i_13_335_4018_0,
    i_13_335_4054_0, i_13_335_4079_0, i_13_335_4160_0, i_13_335_4162_0,
    i_13_335_4163_0, i_13_335_4166_0, i_13_335_4199_0, i_13_335_4369_0,
    i_13_335_4370_0, i_13_335_4372_0, i_13_335_4394_0, i_13_335_4430_0,
    i_13_335_4441_0, i_13_335_4477_0, i_13_335_4555_0, i_13_335_4568_0,
    o_13_335_0_0  );
  input  i_13_335_77_0, i_13_335_92_0, i_13_335_203_0, i_13_335_259_0,
    i_13_335_265_0, i_13_335_266_0, i_13_335_353_0, i_13_335_374_0,
    i_13_335_382_0, i_13_335_413_0, i_13_335_451_0, i_13_335_520_0,
    i_13_335_569_0, i_13_335_605_0, i_13_335_607_0, i_13_335_608_0,
    i_13_335_658_0, i_13_335_661_0, i_13_335_670_0, i_13_335_671_0,
    i_13_335_680_0, i_13_335_929_0, i_13_335_940_0, i_13_335_943_0,
    i_13_335_950_0, i_13_335_1081_0, i_13_335_1082_0, i_13_335_1145_0,
    i_13_335_1148_0, i_13_335_1229_0, i_13_335_1300_0, i_13_335_1307_0,
    i_13_335_1385_0, i_13_335_1444_0, i_13_335_1454_0, i_13_335_1486_0,
    i_13_335_1663_0, i_13_335_1730_0, i_13_335_1733_0, i_13_335_1765_0,
    i_13_335_1766_0, i_13_335_1841_0, i_13_335_1865_0, i_13_335_1885_0,
    i_13_335_1892_0, i_13_335_1927_0, i_13_335_2020_0, i_13_335_2054_0,
    i_13_335_2137_0, i_13_335_2281_0, i_13_335_2300_0, i_13_335_2365_0,
    i_13_335_2423_0, i_13_335_2435_0, i_13_335_2468_0, i_13_335_2546_0,
    i_13_335_2570_0, i_13_335_2614_0, i_13_335_2615_0, i_13_335_2650_0,
    i_13_335_2858_0, i_13_335_2887_0, i_13_335_2980_0, i_13_335_3017_0,
    i_13_335_3047_0, i_13_335_3077_0, i_13_335_3142_0, i_13_335_3259_0,
    i_13_335_3269_0, i_13_335_3343_0, i_13_335_3359_0, i_13_335_3445_0,
    i_13_335_3449_0, i_13_335_3476_0, i_13_335_3484_0, i_13_335_3485_0,
    i_13_335_3646_0, i_13_335_3731_0, i_13_335_3764_0, i_13_335_3781_0,
    i_13_335_3872_0, i_13_335_3875_0, i_13_335_3979_0, i_13_335_4018_0,
    i_13_335_4054_0, i_13_335_4079_0, i_13_335_4160_0, i_13_335_4162_0,
    i_13_335_4163_0, i_13_335_4166_0, i_13_335_4199_0, i_13_335_4369_0,
    i_13_335_4370_0, i_13_335_4372_0, i_13_335_4394_0, i_13_335_4430_0,
    i_13_335_4441_0, i_13_335_4477_0, i_13_335_4555_0, i_13_335_4568_0;
  output o_13_335_0_0;
  assign o_13_335_0_0 = ~((~i_13_335_940_0 & ((~i_13_335_943_0 & ~i_13_335_1082_0 & ~i_13_335_1766_0 & ~i_13_335_3485_0) | (i_13_335_382_0 & ~i_13_335_1454_0 & ~i_13_335_4163_0))) | (~i_13_335_1307_0 & ((~i_13_335_671_0 & i_13_335_2435_0 & ~i_13_335_3872_0 & i_13_335_4370_0) | (~i_13_335_92_0 & ~i_13_335_1730_0 & i_13_335_3142_0 & ~i_13_335_3484_0 & ~i_13_335_4163_0 & ~i_13_335_4555_0))) | (~i_13_335_1765_0 & ((i_13_335_2137_0 & ~i_13_335_4079_0) | (~i_13_335_77_0 & ~i_13_335_353_0 & ~i_13_335_3781_0 & ~i_13_335_4370_0))) | (~i_13_335_1081_0 & ~i_13_335_1841_0 & ~i_13_335_2650_0 & ~i_13_335_4370_0) | (~i_13_335_929_0 & ~i_13_335_943_0 & ~i_13_335_2137_0 & ~i_13_335_2858_0 & ~i_13_335_3646_0 & ~i_13_335_3875_0 & ~i_13_335_3979_0 & ~i_13_335_4160_0) | (i_13_335_1486_0 & ~i_13_335_2435_0 & ~i_13_335_4162_0));
endmodule



// Benchmark "kernel_13_336" written by ABC on Sun Jul 19 10:50:03 2020

module kernel_13_336 ( 
    i_13_336_39_0, i_13_336_76_0, i_13_336_137_0, i_13_336_156_0,
    i_13_336_157_0, i_13_336_193_0, i_13_336_238_0, i_13_336_279_0,
    i_13_336_280_0, i_13_336_310_0, i_13_336_313_0, i_13_336_316_0,
    i_13_336_337_0, i_13_336_360_0, i_13_336_373_0, i_13_336_428_0,
    i_13_336_454_0, i_13_336_490_0, i_13_336_550_0, i_13_336_562_0,
    i_13_336_641_0, i_13_336_643_0, i_13_336_685_0, i_13_336_686_0,
    i_13_336_688_0, i_13_336_756_0, i_13_336_757_0, i_13_336_770_0,
    i_13_336_819_0, i_13_336_895_0, i_13_336_949_0, i_13_336_1057_0,
    i_13_336_1118_0, i_13_336_1120_0, i_13_336_1121_0, i_13_336_1122_0,
    i_13_336_1272_0, i_13_336_1273_0, i_13_336_1364_0, i_13_336_1371_0,
    i_13_336_1498_0, i_13_336_1552_0, i_13_336_1669_0, i_13_336_1722_0,
    i_13_336_1750_0, i_13_336_1813_0, i_13_336_1858_0, i_13_336_1884_0,
    i_13_336_1943_0, i_13_336_2053_0, i_13_336_2101_0, i_13_336_2153_0,
    i_13_336_2190_0, i_13_336_2200_0, i_13_336_2296_0, i_13_336_2548_0,
    i_13_336_2592_0, i_13_336_2614_0, i_13_336_2647_0, i_13_336_2650_0,
    i_13_336_2677_0, i_13_336_2695_0, i_13_336_2722_0, i_13_336_2767_0,
    i_13_336_2857_0, i_13_336_3002_0, i_13_336_3088_0, i_13_336_3127_0,
    i_13_336_3217_0, i_13_336_3235_0, i_13_336_3262_0, i_13_336_3303_0,
    i_13_336_3384_0, i_13_336_3403_0, i_13_336_3478_0, i_13_336_3847_0,
    i_13_336_3889_0, i_13_336_3928_0, i_13_336_3982_0, i_13_336_3990_0,
    i_13_336_3991_0, i_13_336_3992_0, i_13_336_4032_0, i_13_336_4033_0,
    i_13_336_4045_0, i_13_336_4075_0, i_13_336_4078_0, i_13_336_4081_0,
    i_13_336_4082_0, i_13_336_4153_0, i_13_336_4186_0, i_13_336_4187_0,
    i_13_336_4258_0, i_13_336_4270_0, i_13_336_4540_0, i_13_336_4560_0,
    i_13_336_4592_0, i_13_336_4594_0, i_13_336_4595_0, i_13_336_4600_0,
    o_13_336_0_0  );
  input  i_13_336_39_0, i_13_336_76_0, i_13_336_137_0, i_13_336_156_0,
    i_13_336_157_0, i_13_336_193_0, i_13_336_238_0, i_13_336_279_0,
    i_13_336_280_0, i_13_336_310_0, i_13_336_313_0, i_13_336_316_0,
    i_13_336_337_0, i_13_336_360_0, i_13_336_373_0, i_13_336_428_0,
    i_13_336_454_0, i_13_336_490_0, i_13_336_550_0, i_13_336_562_0,
    i_13_336_641_0, i_13_336_643_0, i_13_336_685_0, i_13_336_686_0,
    i_13_336_688_0, i_13_336_756_0, i_13_336_757_0, i_13_336_770_0,
    i_13_336_819_0, i_13_336_895_0, i_13_336_949_0, i_13_336_1057_0,
    i_13_336_1118_0, i_13_336_1120_0, i_13_336_1121_0, i_13_336_1122_0,
    i_13_336_1272_0, i_13_336_1273_0, i_13_336_1364_0, i_13_336_1371_0,
    i_13_336_1498_0, i_13_336_1552_0, i_13_336_1669_0, i_13_336_1722_0,
    i_13_336_1750_0, i_13_336_1813_0, i_13_336_1858_0, i_13_336_1884_0,
    i_13_336_1943_0, i_13_336_2053_0, i_13_336_2101_0, i_13_336_2153_0,
    i_13_336_2190_0, i_13_336_2200_0, i_13_336_2296_0, i_13_336_2548_0,
    i_13_336_2592_0, i_13_336_2614_0, i_13_336_2647_0, i_13_336_2650_0,
    i_13_336_2677_0, i_13_336_2695_0, i_13_336_2722_0, i_13_336_2767_0,
    i_13_336_2857_0, i_13_336_3002_0, i_13_336_3088_0, i_13_336_3127_0,
    i_13_336_3217_0, i_13_336_3235_0, i_13_336_3262_0, i_13_336_3303_0,
    i_13_336_3384_0, i_13_336_3403_0, i_13_336_3478_0, i_13_336_3847_0,
    i_13_336_3889_0, i_13_336_3928_0, i_13_336_3982_0, i_13_336_3990_0,
    i_13_336_3991_0, i_13_336_3992_0, i_13_336_4032_0, i_13_336_4033_0,
    i_13_336_4045_0, i_13_336_4075_0, i_13_336_4078_0, i_13_336_4081_0,
    i_13_336_4082_0, i_13_336_4153_0, i_13_336_4186_0, i_13_336_4187_0,
    i_13_336_4258_0, i_13_336_4270_0, i_13_336_4540_0, i_13_336_4560_0,
    i_13_336_4592_0, i_13_336_4594_0, i_13_336_4595_0, i_13_336_4600_0;
  output o_13_336_0_0;
  assign o_13_336_0_0 = ~((i_13_336_3217_0 & ((~i_13_336_1122_0 & ~i_13_336_4186_0) | (~i_13_336_279_0 & i_13_336_949_0 & ~i_13_336_4187_0))) | (~i_13_336_4033_0 & (~i_13_336_1750_0 | (~i_13_336_4187_0 & i_13_336_4270_0))) | (~i_13_336_819_0 & i_13_336_1498_0 & i_13_336_4270_0) | (~i_13_336_1273_0 & i_13_336_4045_0 & ~i_13_336_4078_0) | (~i_13_336_685_0 & ~i_13_336_1272_0 & ~i_13_336_4082_0) | (i_13_336_1552_0 & ~i_13_336_2650_0 & ~i_13_336_4258_0));
endmodule



// Benchmark "kernel_13_337" written by ABC on Sun Jul 19 10:50:03 2020

module kernel_13_337 ( 
    i_13_337_102_0, i_13_337_103_0, i_13_337_276_0, i_13_337_307_0,
    i_13_337_448_0, i_13_337_450_0, i_13_337_460_0, i_13_337_585_0,
    i_13_337_586_0, i_13_337_598_0, i_13_337_610_0, i_13_337_704_0,
    i_13_337_828_0, i_13_337_843_0, i_13_337_844_0, i_13_337_940_0,
    i_13_337_1063_0, i_13_337_1081_0, i_13_337_1093_0, i_13_337_1095_0,
    i_13_337_1206_0, i_13_337_1305_0, i_13_337_1309_0, i_13_337_1341_0,
    i_13_337_1342_0, i_13_337_1380_0, i_13_337_1399_0, i_13_337_1402_0,
    i_13_337_1440_0, i_13_337_1441_0, i_13_337_1442_0, i_13_337_1473_0,
    i_13_337_1495_0, i_13_337_1529_0, i_13_337_1531_0, i_13_337_1652_0,
    i_13_337_1671_0, i_13_337_1698_0, i_13_337_1744_0, i_13_337_1765_0,
    i_13_337_1795_0, i_13_337_1810_0, i_13_337_1845_0, i_13_337_1927_0,
    i_13_337_1944_0, i_13_337_1990_0, i_13_337_1993_0, i_13_337_2001_0,
    i_13_337_2023_0, i_13_337_2197_0, i_13_337_2236_0, i_13_337_2260_0,
    i_13_337_2277_0, i_13_337_2278_0, i_13_337_2382_0, i_13_337_2448_0,
    i_13_337_2500_0, i_13_337_2547_0, i_13_337_2614_0, i_13_337_2650_0,
    i_13_337_2709_0, i_13_337_2718_0, i_13_337_2719_0, i_13_337_2722_0,
    i_13_337_2742_0, i_13_337_2766_0, i_13_337_2821_0, i_13_337_2919_0,
    i_13_337_2935_0, i_13_337_2949_0, i_13_337_2950_0, i_13_337_3016_0,
    i_13_337_3019_0, i_13_337_3061_0, i_13_337_3122_0, i_13_337_3345_0,
    i_13_337_3366_0, i_13_337_3367_0, i_13_337_3368_0, i_13_337_3390_0,
    i_13_337_3420_0, i_13_337_3454_0, i_13_337_3525_0, i_13_337_3592_0,
    i_13_337_3689_0, i_13_337_3730_0, i_13_337_3741_0, i_13_337_3754_0,
    i_13_337_3856_0, i_13_337_4051_0, i_13_337_4086_0, i_13_337_4165_0,
    i_13_337_4231_0, i_13_337_4257_0, i_13_337_4266_0, i_13_337_4267_0,
    i_13_337_4294_0, i_13_337_4302_0, i_13_337_4393_0, i_13_337_4448_0,
    o_13_337_0_0  );
  input  i_13_337_102_0, i_13_337_103_0, i_13_337_276_0, i_13_337_307_0,
    i_13_337_448_0, i_13_337_450_0, i_13_337_460_0, i_13_337_585_0,
    i_13_337_586_0, i_13_337_598_0, i_13_337_610_0, i_13_337_704_0,
    i_13_337_828_0, i_13_337_843_0, i_13_337_844_0, i_13_337_940_0,
    i_13_337_1063_0, i_13_337_1081_0, i_13_337_1093_0, i_13_337_1095_0,
    i_13_337_1206_0, i_13_337_1305_0, i_13_337_1309_0, i_13_337_1341_0,
    i_13_337_1342_0, i_13_337_1380_0, i_13_337_1399_0, i_13_337_1402_0,
    i_13_337_1440_0, i_13_337_1441_0, i_13_337_1442_0, i_13_337_1473_0,
    i_13_337_1495_0, i_13_337_1529_0, i_13_337_1531_0, i_13_337_1652_0,
    i_13_337_1671_0, i_13_337_1698_0, i_13_337_1744_0, i_13_337_1765_0,
    i_13_337_1795_0, i_13_337_1810_0, i_13_337_1845_0, i_13_337_1927_0,
    i_13_337_1944_0, i_13_337_1990_0, i_13_337_1993_0, i_13_337_2001_0,
    i_13_337_2023_0, i_13_337_2197_0, i_13_337_2236_0, i_13_337_2260_0,
    i_13_337_2277_0, i_13_337_2278_0, i_13_337_2382_0, i_13_337_2448_0,
    i_13_337_2500_0, i_13_337_2547_0, i_13_337_2614_0, i_13_337_2650_0,
    i_13_337_2709_0, i_13_337_2718_0, i_13_337_2719_0, i_13_337_2722_0,
    i_13_337_2742_0, i_13_337_2766_0, i_13_337_2821_0, i_13_337_2919_0,
    i_13_337_2935_0, i_13_337_2949_0, i_13_337_2950_0, i_13_337_3016_0,
    i_13_337_3019_0, i_13_337_3061_0, i_13_337_3122_0, i_13_337_3345_0,
    i_13_337_3366_0, i_13_337_3367_0, i_13_337_3368_0, i_13_337_3390_0,
    i_13_337_3420_0, i_13_337_3454_0, i_13_337_3525_0, i_13_337_3592_0,
    i_13_337_3689_0, i_13_337_3730_0, i_13_337_3741_0, i_13_337_3754_0,
    i_13_337_3856_0, i_13_337_4051_0, i_13_337_4086_0, i_13_337_4165_0,
    i_13_337_4231_0, i_13_337_4257_0, i_13_337_4266_0, i_13_337_4267_0,
    i_13_337_4294_0, i_13_337_4302_0, i_13_337_4393_0, i_13_337_4448_0;
  output o_13_337_0_0;
  assign o_13_337_0_0 = ~((~i_13_337_828_0 & ~i_13_337_1342_0) | (~i_13_337_1206_0 & ~i_13_337_1495_0 & ~i_13_337_4302_0) | (i_13_337_103_0 & ~i_13_337_4266_0 & ~i_13_337_4267_0));
endmodule



// Benchmark "kernel_13_338" written by ABC on Sun Jul 19 10:50:04 2020

module kernel_13_338 ( 
    i_13_338_76_0, i_13_338_118_0, i_13_338_121_0, i_13_338_158_0,
    i_13_338_184_0, i_13_338_186_0, i_13_338_376_0, i_13_338_508_0,
    i_13_338_517_0, i_13_338_526_0, i_13_338_535_0, i_13_338_557_0,
    i_13_338_600_0, i_13_338_616_0, i_13_338_617_0, i_13_338_661_0,
    i_13_338_670_0, i_13_338_737_0, i_13_338_778_0, i_13_338_850_0,
    i_13_338_931_0, i_13_338_945_0, i_13_338_946_0, i_13_338_1067_0,
    i_13_338_1069_0, i_13_338_1084_0, i_13_338_1191_0, i_13_338_1210_0,
    i_13_338_1276_0, i_13_338_1406_0, i_13_338_1424_0, i_13_338_1444_0,
    i_13_338_1545_0, i_13_338_1552_0, i_13_338_1558_0, i_13_338_1624_0,
    i_13_338_1631_0, i_13_338_1723_0, i_13_338_1725_0, i_13_338_1786_0,
    i_13_338_1814_0, i_13_338_1841_0, i_13_338_1938_0, i_13_338_1940_0,
    i_13_338_2120_0, i_13_338_2200_0, i_13_338_2209_0, i_13_338_2211_0,
    i_13_338_2212_0, i_13_338_2365_0, i_13_338_2427_0, i_13_338_2434_0,
    i_13_338_2459_0, i_13_338_2461_0, i_13_338_2713_0, i_13_338_2938_0,
    i_13_338_2939_0, i_13_338_3019_0, i_13_338_3020_0, i_13_338_3028_0,
    i_13_338_3029_0, i_13_338_3037_0, i_13_338_3039_0, i_13_338_3040_0,
    i_13_338_3044_0, i_13_338_3139_0, i_13_338_3160_0, i_13_338_3162_0,
    i_13_338_3163_0, i_13_338_3164_0, i_13_338_3165_0, i_13_338_3205_0,
    i_13_338_3209_0, i_13_338_3217_0, i_13_338_3218_0, i_13_338_3250_0,
    i_13_338_3289_0, i_13_338_3292_0, i_13_338_3413_0, i_13_338_3421_0,
    i_13_338_3424_0, i_13_338_3541_0, i_13_338_3545_0, i_13_338_3595_0,
    i_13_338_3874_0, i_13_338_3899_0, i_13_338_4009_0, i_13_338_4194_0,
    i_13_338_4233_0, i_13_338_4234_0, i_13_338_4271_0, i_13_338_4312_0,
    i_13_338_4333_0, i_13_338_4352_0, i_13_338_4360_0, i_13_338_4361_0,
    i_13_338_4414_0, i_13_338_4498_0, i_13_338_4526_0, i_13_338_4544_0,
    o_13_338_0_0  );
  input  i_13_338_76_0, i_13_338_118_0, i_13_338_121_0, i_13_338_158_0,
    i_13_338_184_0, i_13_338_186_0, i_13_338_376_0, i_13_338_508_0,
    i_13_338_517_0, i_13_338_526_0, i_13_338_535_0, i_13_338_557_0,
    i_13_338_600_0, i_13_338_616_0, i_13_338_617_0, i_13_338_661_0,
    i_13_338_670_0, i_13_338_737_0, i_13_338_778_0, i_13_338_850_0,
    i_13_338_931_0, i_13_338_945_0, i_13_338_946_0, i_13_338_1067_0,
    i_13_338_1069_0, i_13_338_1084_0, i_13_338_1191_0, i_13_338_1210_0,
    i_13_338_1276_0, i_13_338_1406_0, i_13_338_1424_0, i_13_338_1444_0,
    i_13_338_1545_0, i_13_338_1552_0, i_13_338_1558_0, i_13_338_1624_0,
    i_13_338_1631_0, i_13_338_1723_0, i_13_338_1725_0, i_13_338_1786_0,
    i_13_338_1814_0, i_13_338_1841_0, i_13_338_1938_0, i_13_338_1940_0,
    i_13_338_2120_0, i_13_338_2200_0, i_13_338_2209_0, i_13_338_2211_0,
    i_13_338_2212_0, i_13_338_2365_0, i_13_338_2427_0, i_13_338_2434_0,
    i_13_338_2459_0, i_13_338_2461_0, i_13_338_2713_0, i_13_338_2938_0,
    i_13_338_2939_0, i_13_338_3019_0, i_13_338_3020_0, i_13_338_3028_0,
    i_13_338_3029_0, i_13_338_3037_0, i_13_338_3039_0, i_13_338_3040_0,
    i_13_338_3044_0, i_13_338_3139_0, i_13_338_3160_0, i_13_338_3162_0,
    i_13_338_3163_0, i_13_338_3164_0, i_13_338_3165_0, i_13_338_3205_0,
    i_13_338_3209_0, i_13_338_3217_0, i_13_338_3218_0, i_13_338_3250_0,
    i_13_338_3289_0, i_13_338_3292_0, i_13_338_3413_0, i_13_338_3421_0,
    i_13_338_3424_0, i_13_338_3541_0, i_13_338_3545_0, i_13_338_3595_0,
    i_13_338_3874_0, i_13_338_3899_0, i_13_338_4009_0, i_13_338_4194_0,
    i_13_338_4233_0, i_13_338_4234_0, i_13_338_4271_0, i_13_338_4312_0,
    i_13_338_4333_0, i_13_338_4352_0, i_13_338_4360_0, i_13_338_4361_0,
    i_13_338_4414_0, i_13_338_4498_0, i_13_338_4526_0, i_13_338_4544_0;
  output o_13_338_0_0;
  assign o_13_338_0_0 = ~((i_13_338_1210_0 & (i_13_338_517_0 | i_13_338_3541_0)) | (~i_13_338_2212_0 & ((~i_13_338_3205_0 & ~i_13_338_3292_0 & ~i_13_338_3421_0 & ~i_13_338_3899_0) | (i_13_338_3595_0 & ~i_13_338_4352_0))) | (i_13_338_3541_0 & ((~i_13_338_931_0 & ~i_13_338_3205_0) | (~i_13_338_3218_0 & ~i_13_338_4414_0))) | (~i_13_338_3218_0 & ((i_13_338_670_0 & ~i_13_338_945_0 & ~i_13_338_946_0 & ~i_13_338_3040_0) | (~i_13_338_186_0 & ~i_13_338_616_0 & ~i_13_338_1084_0 & ~i_13_338_2713_0 & ~i_13_338_3164_0 & ~i_13_338_4233_0 & ~i_13_338_4312_0))) | (~i_13_338_737_0 & ~i_13_338_1067_0 & ~i_13_338_2209_0 & ~i_13_338_3162_0) | (i_13_338_3162_0 & ~i_13_338_3217_0 & ~i_13_338_4414_0));
endmodule



// Benchmark "kernel_13_339" written by ABC on Sun Jul 19 10:50:05 2020

module kernel_13_339 ( 
    i_13_339_110_0, i_13_339_184_0, i_13_339_186_0, i_13_339_192_0,
    i_13_339_193_0, i_13_339_194_0, i_13_339_195_0, i_13_339_328_0,
    i_13_339_333_0, i_13_339_572_0, i_13_339_573_0, i_13_339_618_0,
    i_13_339_625_0, i_13_339_641_0, i_13_339_658_0, i_13_339_715_0,
    i_13_339_716_0, i_13_339_858_0, i_13_339_859_0, i_13_339_867_0,
    i_13_339_868_0, i_13_339_928_0, i_13_339_955_0, i_13_339_1116_0,
    i_13_339_1117_0, i_13_339_1148_0, i_13_339_1149_0, i_13_339_1210_0,
    i_13_339_1225_0, i_13_339_1226_0, i_13_339_1228_0, i_13_339_1229_0,
    i_13_339_1256_0, i_13_339_1258_0, i_13_339_1259_0, i_13_339_1329_0,
    i_13_339_1404_0, i_13_339_1405_0, i_13_339_1408_0, i_13_339_1411_0,
    i_13_339_1507_0, i_13_339_1513_0, i_13_339_1570_0, i_13_339_1597_0,
    i_13_339_1678_0, i_13_339_1680_0, i_13_339_1729_0, i_13_339_1734_0,
    i_13_339_1765_0, i_13_339_1768_0, i_13_339_1801_0, i_13_339_1802_0,
    i_13_339_1829_0, i_13_339_1956_0, i_13_339_1991_0, i_13_339_2002_0,
    i_13_339_2056_0, i_13_339_2059_0, i_13_339_2225_0, i_13_339_2281_0,
    i_13_339_2302_0, i_13_339_2341_0, i_13_339_2532_0, i_13_339_2614_0,
    i_13_339_2619_0, i_13_339_2648_0, i_13_339_2705_0, i_13_339_2746_0,
    i_13_339_2857_0, i_13_339_2981_0, i_13_339_3034_0, i_13_339_3064_0,
    i_13_339_3118_0, i_13_339_3145_0, i_13_339_3214_0, i_13_339_3258_0,
    i_13_339_3268_0, i_13_339_3269_0, i_13_339_3287_0, i_13_339_3291_0,
    i_13_339_3310_0, i_13_339_3386_0, i_13_339_3421_0, i_13_339_3424_0,
    i_13_339_3546_0, i_13_339_3562_0, i_13_339_3606_0, i_13_339_3755_0,
    i_13_339_3763_0, i_13_339_3764_0, i_13_339_3979_0, i_13_339_4018_0,
    i_13_339_4078_0, i_13_339_4201_0, i_13_339_4202_0, i_13_339_4213_0,
    i_13_339_4267_0, i_13_339_4297_0, i_13_339_4362_0, i_13_339_4515_0,
    o_13_339_0_0  );
  input  i_13_339_110_0, i_13_339_184_0, i_13_339_186_0, i_13_339_192_0,
    i_13_339_193_0, i_13_339_194_0, i_13_339_195_0, i_13_339_328_0,
    i_13_339_333_0, i_13_339_572_0, i_13_339_573_0, i_13_339_618_0,
    i_13_339_625_0, i_13_339_641_0, i_13_339_658_0, i_13_339_715_0,
    i_13_339_716_0, i_13_339_858_0, i_13_339_859_0, i_13_339_867_0,
    i_13_339_868_0, i_13_339_928_0, i_13_339_955_0, i_13_339_1116_0,
    i_13_339_1117_0, i_13_339_1148_0, i_13_339_1149_0, i_13_339_1210_0,
    i_13_339_1225_0, i_13_339_1226_0, i_13_339_1228_0, i_13_339_1229_0,
    i_13_339_1256_0, i_13_339_1258_0, i_13_339_1259_0, i_13_339_1329_0,
    i_13_339_1404_0, i_13_339_1405_0, i_13_339_1408_0, i_13_339_1411_0,
    i_13_339_1507_0, i_13_339_1513_0, i_13_339_1570_0, i_13_339_1597_0,
    i_13_339_1678_0, i_13_339_1680_0, i_13_339_1729_0, i_13_339_1734_0,
    i_13_339_1765_0, i_13_339_1768_0, i_13_339_1801_0, i_13_339_1802_0,
    i_13_339_1829_0, i_13_339_1956_0, i_13_339_1991_0, i_13_339_2002_0,
    i_13_339_2056_0, i_13_339_2059_0, i_13_339_2225_0, i_13_339_2281_0,
    i_13_339_2302_0, i_13_339_2341_0, i_13_339_2532_0, i_13_339_2614_0,
    i_13_339_2619_0, i_13_339_2648_0, i_13_339_2705_0, i_13_339_2746_0,
    i_13_339_2857_0, i_13_339_2981_0, i_13_339_3034_0, i_13_339_3064_0,
    i_13_339_3118_0, i_13_339_3145_0, i_13_339_3214_0, i_13_339_3258_0,
    i_13_339_3268_0, i_13_339_3269_0, i_13_339_3287_0, i_13_339_3291_0,
    i_13_339_3310_0, i_13_339_3386_0, i_13_339_3421_0, i_13_339_3424_0,
    i_13_339_3546_0, i_13_339_3562_0, i_13_339_3606_0, i_13_339_3755_0,
    i_13_339_3763_0, i_13_339_3764_0, i_13_339_3979_0, i_13_339_4018_0,
    i_13_339_4078_0, i_13_339_4201_0, i_13_339_4202_0, i_13_339_4213_0,
    i_13_339_4267_0, i_13_339_4297_0, i_13_339_4362_0, i_13_339_4515_0;
  output o_13_339_0_0;
  assign o_13_339_0_0 = ~((i_13_339_2532_0 & ~i_13_339_3763_0) | (~i_13_339_1678_0 & ~i_13_339_1802_0) | (~i_13_339_194_0 & ~i_13_339_1408_0) | (~i_13_339_333_0 & ~i_13_339_2648_0 & ~i_13_339_3755_0));
endmodule



// Benchmark "kernel_13_340" written by ABC on Sun Jul 19 10:50:06 2020

module kernel_13_340 ( 
    i_13_340_45_0, i_13_340_46_0, i_13_340_55_0, i_13_340_103_0,
    i_13_340_138_0, i_13_340_154_0, i_13_340_186_0, i_13_340_255_0,
    i_13_340_258_0, i_13_340_259_0, i_13_340_307_0, i_13_340_309_0,
    i_13_340_352_0, i_13_340_408_0, i_13_340_450_0, i_13_340_505_0,
    i_13_340_644_0, i_13_340_660_0, i_13_340_667_0, i_13_340_848_0,
    i_13_340_894_0, i_13_340_930_0, i_13_340_936_0, i_13_340_937_0,
    i_13_340_1108_0, i_13_340_1227_0, i_13_340_1228_0, i_13_340_1243_0,
    i_13_340_1326_0, i_13_340_1328_0, i_13_340_1399_0, i_13_340_1479_0,
    i_13_340_1513_0, i_13_340_1623_0, i_13_340_1660_0, i_13_340_1677_0,
    i_13_340_1723_0, i_13_340_1764_0, i_13_340_1767_0, i_13_340_1801_0,
    i_13_340_1803_0, i_13_340_1804_0, i_13_340_1944_0, i_13_340_1945_0,
    i_13_340_1948_0, i_13_340_2025_0, i_13_340_2026_0, i_13_340_2053_0,
    i_13_340_2134_0, i_13_340_2145_0, i_13_340_2197_0, i_13_340_2206_0,
    i_13_340_2277_0, i_13_340_2297_0, i_13_340_2403_0, i_13_340_2404_0,
    i_13_340_2430_0, i_13_340_2471_0, i_13_340_2578_0, i_13_340_2611_0,
    i_13_340_2613_0, i_13_340_2622_0, i_13_340_2745_0, i_13_340_2793_0,
    i_13_340_2848_0, i_13_340_2916_0, i_13_340_2980_0, i_13_340_3001_0,
    i_13_340_3027_0, i_13_340_3028_0, i_13_340_3073_0, i_13_340_3133_0,
    i_13_340_3213_0, i_13_340_3352_0, i_13_340_3367_0, i_13_340_3378_0,
    i_13_340_3439_0, i_13_340_3591_0, i_13_340_3592_0, i_13_340_3703_0,
    i_13_340_3763_0, i_13_340_3780_0, i_13_340_3820_0, i_13_340_3898_0,
    i_13_340_3978_0, i_13_340_3979_0, i_13_340_4017_0, i_13_340_4158_0,
    i_13_340_4231_0, i_13_340_4249_0, i_13_340_4302_0, i_13_340_4332_0,
    i_13_340_4351_0, i_13_340_4360_0, i_13_340_4367_0, i_13_340_4387_0,
    i_13_340_4438_0, i_13_340_4446_0, i_13_340_4563_0, i_13_340_4602_0,
    o_13_340_0_0  );
  input  i_13_340_45_0, i_13_340_46_0, i_13_340_55_0, i_13_340_103_0,
    i_13_340_138_0, i_13_340_154_0, i_13_340_186_0, i_13_340_255_0,
    i_13_340_258_0, i_13_340_259_0, i_13_340_307_0, i_13_340_309_0,
    i_13_340_352_0, i_13_340_408_0, i_13_340_450_0, i_13_340_505_0,
    i_13_340_644_0, i_13_340_660_0, i_13_340_667_0, i_13_340_848_0,
    i_13_340_894_0, i_13_340_930_0, i_13_340_936_0, i_13_340_937_0,
    i_13_340_1108_0, i_13_340_1227_0, i_13_340_1228_0, i_13_340_1243_0,
    i_13_340_1326_0, i_13_340_1328_0, i_13_340_1399_0, i_13_340_1479_0,
    i_13_340_1513_0, i_13_340_1623_0, i_13_340_1660_0, i_13_340_1677_0,
    i_13_340_1723_0, i_13_340_1764_0, i_13_340_1767_0, i_13_340_1801_0,
    i_13_340_1803_0, i_13_340_1804_0, i_13_340_1944_0, i_13_340_1945_0,
    i_13_340_1948_0, i_13_340_2025_0, i_13_340_2026_0, i_13_340_2053_0,
    i_13_340_2134_0, i_13_340_2145_0, i_13_340_2197_0, i_13_340_2206_0,
    i_13_340_2277_0, i_13_340_2297_0, i_13_340_2403_0, i_13_340_2404_0,
    i_13_340_2430_0, i_13_340_2471_0, i_13_340_2578_0, i_13_340_2611_0,
    i_13_340_2613_0, i_13_340_2622_0, i_13_340_2745_0, i_13_340_2793_0,
    i_13_340_2848_0, i_13_340_2916_0, i_13_340_2980_0, i_13_340_3001_0,
    i_13_340_3027_0, i_13_340_3028_0, i_13_340_3073_0, i_13_340_3133_0,
    i_13_340_3213_0, i_13_340_3352_0, i_13_340_3367_0, i_13_340_3378_0,
    i_13_340_3439_0, i_13_340_3591_0, i_13_340_3592_0, i_13_340_3703_0,
    i_13_340_3763_0, i_13_340_3780_0, i_13_340_3820_0, i_13_340_3898_0,
    i_13_340_3978_0, i_13_340_3979_0, i_13_340_4017_0, i_13_340_4158_0,
    i_13_340_4231_0, i_13_340_4249_0, i_13_340_4302_0, i_13_340_4332_0,
    i_13_340_4351_0, i_13_340_4360_0, i_13_340_4367_0, i_13_340_4387_0,
    i_13_340_4438_0, i_13_340_4446_0, i_13_340_4563_0, i_13_340_4602_0;
  output o_13_340_0_0;
  assign o_13_340_0_0 = ~((~i_13_340_2025_0 & (~i_13_340_2980_0 | (~i_13_340_930_0 & ~i_13_340_1764_0 & ~i_13_340_2916_0 & ~i_13_340_3898_0))) | (~i_13_340_936_0 & ~i_13_340_2404_0 & ~i_13_340_4563_0));
endmodule



// Benchmark "kernel_13_341" written by ABC on Sun Jul 19 10:50:07 2020

module kernel_13_341 ( 
    i_13_341_97_0, i_13_341_107_0, i_13_341_119_0, i_13_341_121_0,
    i_13_341_122_0, i_13_341_181_0, i_13_341_285_0, i_13_341_286_0,
    i_13_341_311_0, i_13_341_320_0, i_13_341_430_0, i_13_341_535_0,
    i_13_341_538_0, i_13_341_569_0, i_13_341_599_0, i_13_341_697_0,
    i_13_341_712_0, i_13_341_746_0, i_13_341_781_0, i_13_341_850_0,
    i_13_341_934_0, i_13_341_976_0, i_13_341_985_0, i_13_341_1034_0,
    i_13_341_1093_0, i_13_341_1094_0, i_13_341_1216_0, i_13_341_1279_0,
    i_13_341_1283_0, i_13_341_1284_0, i_13_341_1300_0, i_13_341_1471_0,
    i_13_341_1526_0, i_13_341_1552_0, i_13_341_1714_0, i_13_341_1721_0,
    i_13_341_1726_0, i_13_341_1757_0, i_13_341_1760_0, i_13_341_1783_0,
    i_13_341_1786_0, i_13_341_1787_0, i_13_341_1789_0, i_13_341_1817_0,
    i_13_341_2072_0, i_13_341_2120_0, i_13_341_2123_0, i_13_341_2209_0,
    i_13_341_2308_0, i_13_341_2312_0, i_13_341_2365_0, i_13_341_2458_0,
    i_13_341_2459_0, i_13_341_2465_0, i_13_341_2551_0, i_13_341_2630_0,
    i_13_341_2633_0, i_13_341_2663_0, i_13_341_2939_0, i_13_341_3040_0,
    i_13_341_3148_0, i_13_341_3161_0, i_13_341_3163_0, i_13_341_3167_0,
    i_13_341_3211_0, i_13_341_3212_0, i_13_341_3218_0, i_13_341_3265_0,
    i_13_341_3271_0, i_13_341_3347_0, i_13_341_3424_0, i_13_341_3482_0,
    i_13_341_3483_0, i_13_341_3506_0, i_13_341_3523_0, i_13_341_3527_0,
    i_13_341_3688_0, i_13_341_3689_0, i_13_341_3700_0, i_13_341_3746_0,
    i_13_341_3844_0, i_13_341_3871_0, i_13_341_3878_0, i_13_341_3935_0,
    i_13_341_3962_0, i_13_341_4009_0, i_13_341_4012_0, i_13_341_4048_0,
    i_13_341_4093_0, i_13_341_4105_0, i_13_341_4106_0, i_13_341_4235_0,
    i_13_341_4237_0, i_13_341_4238_0, i_13_341_4261_0, i_13_341_4273_0,
    i_13_341_4414_0, i_13_341_4417_0, i_13_341_4450_0, i_13_341_4519_0,
    o_13_341_0_0  );
  input  i_13_341_97_0, i_13_341_107_0, i_13_341_119_0, i_13_341_121_0,
    i_13_341_122_0, i_13_341_181_0, i_13_341_285_0, i_13_341_286_0,
    i_13_341_311_0, i_13_341_320_0, i_13_341_430_0, i_13_341_535_0,
    i_13_341_538_0, i_13_341_569_0, i_13_341_599_0, i_13_341_697_0,
    i_13_341_712_0, i_13_341_746_0, i_13_341_781_0, i_13_341_850_0,
    i_13_341_934_0, i_13_341_976_0, i_13_341_985_0, i_13_341_1034_0,
    i_13_341_1093_0, i_13_341_1094_0, i_13_341_1216_0, i_13_341_1279_0,
    i_13_341_1283_0, i_13_341_1284_0, i_13_341_1300_0, i_13_341_1471_0,
    i_13_341_1526_0, i_13_341_1552_0, i_13_341_1714_0, i_13_341_1721_0,
    i_13_341_1726_0, i_13_341_1757_0, i_13_341_1760_0, i_13_341_1783_0,
    i_13_341_1786_0, i_13_341_1787_0, i_13_341_1789_0, i_13_341_1817_0,
    i_13_341_2072_0, i_13_341_2120_0, i_13_341_2123_0, i_13_341_2209_0,
    i_13_341_2308_0, i_13_341_2312_0, i_13_341_2365_0, i_13_341_2458_0,
    i_13_341_2459_0, i_13_341_2465_0, i_13_341_2551_0, i_13_341_2630_0,
    i_13_341_2633_0, i_13_341_2663_0, i_13_341_2939_0, i_13_341_3040_0,
    i_13_341_3148_0, i_13_341_3161_0, i_13_341_3163_0, i_13_341_3167_0,
    i_13_341_3211_0, i_13_341_3212_0, i_13_341_3218_0, i_13_341_3265_0,
    i_13_341_3271_0, i_13_341_3347_0, i_13_341_3424_0, i_13_341_3482_0,
    i_13_341_3483_0, i_13_341_3506_0, i_13_341_3523_0, i_13_341_3527_0,
    i_13_341_3688_0, i_13_341_3689_0, i_13_341_3700_0, i_13_341_3746_0,
    i_13_341_3844_0, i_13_341_3871_0, i_13_341_3878_0, i_13_341_3935_0,
    i_13_341_3962_0, i_13_341_4009_0, i_13_341_4012_0, i_13_341_4048_0,
    i_13_341_4093_0, i_13_341_4105_0, i_13_341_4106_0, i_13_341_4235_0,
    i_13_341_4237_0, i_13_341_4238_0, i_13_341_4261_0, i_13_341_4273_0,
    i_13_341_4414_0, i_13_341_4417_0, i_13_341_4450_0, i_13_341_4519_0;
  output o_13_341_0_0;
  assign o_13_341_0_0 = ~((~i_13_341_2209_0 & ((~i_13_341_538_0 & i_13_341_985_0 & ~i_13_341_3689_0 & ~i_13_341_4238_0) | (~i_13_341_121_0 & ~i_13_341_4417_0))) | (~i_13_341_4009_0 & ((~i_13_341_122_0 & i_13_341_286_0) | (~i_13_341_1471_0 & i_13_341_4012_0))) | (~i_13_341_4235_0 & ((i_13_341_1471_0 & ~i_13_341_1714_0 & ~i_13_341_4273_0) | (~i_13_341_1817_0 & ~i_13_341_3040_0 & ~i_13_341_4417_0))) | (~i_13_341_535_0 & ~i_13_341_3218_0 & i_13_341_4414_0) | (~i_13_341_3347_0 & ~i_13_341_3689_0 & ~i_13_341_4012_0 & i_13_341_4450_0));
endmodule



// Benchmark "kernel_13_342" written by ABC on Sun Jul 19 10:50:07 2020

module kernel_13_342 ( 
    i_13_342_31_0, i_13_342_93_0, i_13_342_94_0, i_13_342_97_0,
    i_13_342_114_0, i_13_342_121_0, i_13_342_123_0, i_13_342_159_0,
    i_13_342_184_0, i_13_342_328_0, i_13_342_435_0, i_13_342_517_0,
    i_13_342_564_0, i_13_342_570_0, i_13_342_571_0, i_13_342_574_0,
    i_13_342_614_0, i_13_342_696_0, i_13_342_697_0, i_13_342_732_0,
    i_13_342_733_0, i_13_342_742_0, i_13_342_796_0, i_13_342_799_0,
    i_13_342_822_0, i_13_342_1210_0, i_13_342_1254_0, i_13_342_1390_0,
    i_13_342_1408_0, i_13_342_1446_0, i_13_342_1447_0, i_13_342_1456_0,
    i_13_342_1473_0, i_13_342_1489_0, i_13_342_1551_0, i_13_342_1552_0,
    i_13_342_1569_0, i_13_342_1642_0, i_13_342_1761_0, i_13_342_1786_0,
    i_13_342_1789_0, i_13_342_1860_0, i_13_342_1910_0, i_13_342_2018_0,
    i_13_342_2056_0, i_13_342_2103_0, i_13_342_2175_0, i_13_342_2176_0,
    i_13_342_2202_0, i_13_342_2208_0, i_13_342_2235_0, i_13_342_2238_0,
    i_13_342_2269_0, i_13_342_2427_0, i_13_342_2434_0, i_13_342_2541_0,
    i_13_342_2680_0, i_13_342_2767_0, i_13_342_2914_0, i_13_342_2985_0,
    i_13_342_3009_0, i_13_342_3022_0, i_13_342_3028_0, i_13_342_3053_0,
    i_13_342_3091_0, i_13_342_3163_0, i_13_342_3207_0, i_13_342_3243_0,
    i_13_342_3244_0, i_13_342_3415_0, i_13_342_3422_0, i_13_342_3423_0,
    i_13_342_3424_0, i_13_342_3426_0, i_13_342_3427_0, i_13_342_3432_0,
    i_13_342_3451_0, i_13_342_3521_0, i_13_342_3571_0, i_13_342_3649_0,
    i_13_342_3665_0, i_13_342_3702_0, i_13_342_3739_0, i_13_342_3846_0,
    i_13_342_3847_0, i_13_342_3850_0, i_13_342_3873_0, i_13_342_3874_0,
    i_13_342_3876_0, i_13_342_3967_0, i_13_342_4009_0, i_13_342_4038_0,
    i_13_342_4119_0, i_13_342_4188_0, i_13_342_4189_0, i_13_342_4195_0,
    i_13_342_4236_0, i_13_342_4351_0, i_13_342_4353_0, i_13_342_4569_0,
    o_13_342_0_0  );
  input  i_13_342_31_0, i_13_342_93_0, i_13_342_94_0, i_13_342_97_0,
    i_13_342_114_0, i_13_342_121_0, i_13_342_123_0, i_13_342_159_0,
    i_13_342_184_0, i_13_342_328_0, i_13_342_435_0, i_13_342_517_0,
    i_13_342_564_0, i_13_342_570_0, i_13_342_571_0, i_13_342_574_0,
    i_13_342_614_0, i_13_342_696_0, i_13_342_697_0, i_13_342_732_0,
    i_13_342_733_0, i_13_342_742_0, i_13_342_796_0, i_13_342_799_0,
    i_13_342_822_0, i_13_342_1210_0, i_13_342_1254_0, i_13_342_1390_0,
    i_13_342_1408_0, i_13_342_1446_0, i_13_342_1447_0, i_13_342_1456_0,
    i_13_342_1473_0, i_13_342_1489_0, i_13_342_1551_0, i_13_342_1552_0,
    i_13_342_1569_0, i_13_342_1642_0, i_13_342_1761_0, i_13_342_1786_0,
    i_13_342_1789_0, i_13_342_1860_0, i_13_342_1910_0, i_13_342_2018_0,
    i_13_342_2056_0, i_13_342_2103_0, i_13_342_2175_0, i_13_342_2176_0,
    i_13_342_2202_0, i_13_342_2208_0, i_13_342_2235_0, i_13_342_2238_0,
    i_13_342_2269_0, i_13_342_2427_0, i_13_342_2434_0, i_13_342_2541_0,
    i_13_342_2680_0, i_13_342_2767_0, i_13_342_2914_0, i_13_342_2985_0,
    i_13_342_3009_0, i_13_342_3022_0, i_13_342_3028_0, i_13_342_3053_0,
    i_13_342_3091_0, i_13_342_3163_0, i_13_342_3207_0, i_13_342_3243_0,
    i_13_342_3244_0, i_13_342_3415_0, i_13_342_3422_0, i_13_342_3423_0,
    i_13_342_3424_0, i_13_342_3426_0, i_13_342_3427_0, i_13_342_3432_0,
    i_13_342_3451_0, i_13_342_3521_0, i_13_342_3571_0, i_13_342_3649_0,
    i_13_342_3665_0, i_13_342_3702_0, i_13_342_3739_0, i_13_342_3846_0,
    i_13_342_3847_0, i_13_342_3850_0, i_13_342_3873_0, i_13_342_3874_0,
    i_13_342_3876_0, i_13_342_3967_0, i_13_342_4009_0, i_13_342_4038_0,
    i_13_342_4119_0, i_13_342_4188_0, i_13_342_4189_0, i_13_342_4195_0,
    i_13_342_4236_0, i_13_342_4351_0, i_13_342_4353_0, i_13_342_4569_0;
  output o_13_342_0_0;
  assign o_13_342_0_0 = ~((~i_13_342_3244_0 & ((~i_13_342_3423_0 & ~i_13_342_3424_0 & ~i_13_342_3426_0) | (~i_13_342_3009_0 & ~i_13_342_3846_0 & ~i_13_342_3873_0 & ~i_13_342_3874_0))) | (~i_13_342_3874_0 & ((~i_13_342_2176_0 & ~i_13_342_3873_0 & ~i_13_342_4009_0 & ~i_13_342_4353_0) | (i_13_342_1552_0 & ~i_13_342_2175_0 & ~i_13_342_4569_0))) | (i_13_342_697_0 & ~i_13_342_1489_0) | (~i_13_342_570_0 & ~i_13_342_1456_0 & ~i_13_342_2541_0 & i_13_342_3091_0) | (~i_13_342_3091_0 & ~i_13_342_4009_0));
endmodule



// Benchmark "kernel_13_343" written by ABC on Sun Jul 19 10:50:08 2020

module kernel_13_343 ( 
    i_13_343_39_0, i_13_343_48_0, i_13_343_139_0, i_13_343_163_0,
    i_13_343_174_0, i_13_343_274_0, i_13_343_279_0, i_13_343_280_0,
    i_13_343_307_0, i_13_343_310_0, i_13_343_315_0, i_13_343_316_0,
    i_13_343_514_0, i_13_343_549_0, i_13_343_550_0, i_13_343_639_0,
    i_13_343_640_0, i_13_343_646_0, i_13_343_667_0, i_13_343_670_0,
    i_13_343_675_0, i_13_343_676_0, i_13_343_684_0, i_13_343_685_0,
    i_13_343_687_0, i_13_343_688_0, i_13_343_691_0, i_13_343_757_0,
    i_13_343_875_0, i_13_343_981_0, i_13_343_1055_0, i_13_343_1099_0,
    i_13_343_1116_0, i_13_343_1270_0, i_13_343_1363_0, i_13_343_1438_0,
    i_13_343_1445_0, i_13_343_1449_0, i_13_343_1593_0, i_13_343_1594_0,
    i_13_343_1597_0, i_13_343_1632_0, i_13_343_1803_0, i_13_343_1813_0,
    i_13_343_1847_0, i_13_343_2053_0, i_13_343_2236_0, i_13_343_2274_0,
    i_13_343_2313_0, i_13_343_2396_0, i_13_343_2397_0, i_13_343_2422_0,
    i_13_343_2507_0, i_13_343_2614_0, i_13_343_2648_0, i_13_343_2649_0,
    i_13_343_2650_0, i_13_343_2673_0, i_13_343_2674_0, i_13_343_2693_0,
    i_13_343_2694_0, i_13_343_2695_0, i_13_343_2698_0, i_13_343_2929_0,
    i_13_343_3011_0, i_13_343_3034_0, i_13_343_3142_0, i_13_343_3145_0,
    i_13_343_3217_0, i_13_343_3385_0, i_13_343_3415_0, i_13_343_3532_0,
    i_13_343_3610_0, i_13_343_3685_0, i_13_343_3730_0, i_13_343_3736_0,
    i_13_343_3739_0, i_13_343_3816_0, i_13_343_3817_0, i_13_343_3888_0,
    i_13_343_3889_0, i_13_343_3987_0, i_13_343_3991_0, i_13_343_4017_0,
    i_13_343_4032_0, i_13_343_4033_0, i_13_343_4034_0, i_13_343_4077_0,
    i_13_343_4086_0, i_13_343_4187_0, i_13_343_4278_0, i_13_343_4306_0,
    i_13_343_4338_0, i_13_343_4458_0, i_13_343_4531_0, i_13_343_4540_0,
    i_13_343_4590_0, i_13_343_4591_0, i_13_343_4594_0, i_13_343_4600_0,
    o_13_343_0_0  );
  input  i_13_343_39_0, i_13_343_48_0, i_13_343_139_0, i_13_343_163_0,
    i_13_343_174_0, i_13_343_274_0, i_13_343_279_0, i_13_343_280_0,
    i_13_343_307_0, i_13_343_310_0, i_13_343_315_0, i_13_343_316_0,
    i_13_343_514_0, i_13_343_549_0, i_13_343_550_0, i_13_343_639_0,
    i_13_343_640_0, i_13_343_646_0, i_13_343_667_0, i_13_343_670_0,
    i_13_343_675_0, i_13_343_676_0, i_13_343_684_0, i_13_343_685_0,
    i_13_343_687_0, i_13_343_688_0, i_13_343_691_0, i_13_343_757_0,
    i_13_343_875_0, i_13_343_981_0, i_13_343_1055_0, i_13_343_1099_0,
    i_13_343_1116_0, i_13_343_1270_0, i_13_343_1363_0, i_13_343_1438_0,
    i_13_343_1445_0, i_13_343_1449_0, i_13_343_1593_0, i_13_343_1594_0,
    i_13_343_1597_0, i_13_343_1632_0, i_13_343_1803_0, i_13_343_1813_0,
    i_13_343_1847_0, i_13_343_2053_0, i_13_343_2236_0, i_13_343_2274_0,
    i_13_343_2313_0, i_13_343_2396_0, i_13_343_2397_0, i_13_343_2422_0,
    i_13_343_2507_0, i_13_343_2614_0, i_13_343_2648_0, i_13_343_2649_0,
    i_13_343_2650_0, i_13_343_2673_0, i_13_343_2674_0, i_13_343_2693_0,
    i_13_343_2694_0, i_13_343_2695_0, i_13_343_2698_0, i_13_343_2929_0,
    i_13_343_3011_0, i_13_343_3034_0, i_13_343_3142_0, i_13_343_3145_0,
    i_13_343_3217_0, i_13_343_3385_0, i_13_343_3415_0, i_13_343_3532_0,
    i_13_343_3610_0, i_13_343_3685_0, i_13_343_3730_0, i_13_343_3736_0,
    i_13_343_3739_0, i_13_343_3816_0, i_13_343_3817_0, i_13_343_3888_0,
    i_13_343_3889_0, i_13_343_3987_0, i_13_343_3991_0, i_13_343_4017_0,
    i_13_343_4032_0, i_13_343_4033_0, i_13_343_4034_0, i_13_343_4077_0,
    i_13_343_4086_0, i_13_343_4187_0, i_13_343_4278_0, i_13_343_4306_0,
    i_13_343_4338_0, i_13_343_4458_0, i_13_343_4531_0, i_13_343_4540_0,
    i_13_343_4590_0, i_13_343_4591_0, i_13_343_4594_0, i_13_343_4600_0;
  output o_13_343_0_0;
  assign o_13_343_0_0 = ~((i_13_343_4187_0 & (~i_13_343_280_0 | (~i_13_343_1270_0 & ~i_13_343_2053_0) | (~i_13_343_3736_0 & ~i_13_343_3817_0))) | (~i_13_343_307_0 & ~i_13_343_316_0) | (~i_13_343_675_0 & ~i_13_343_3991_0) | (~i_13_343_3730_0 & ~i_13_343_4032_0 & ~i_13_343_4187_0));
endmodule



// Benchmark "kernel_13_344" written by ABC on Sun Jul 19 10:50:09 2020

module kernel_13_344 ( 
    i_13_344_112_0, i_13_344_121_0, i_13_344_122_0, i_13_344_139_0,
    i_13_344_193_0, i_13_344_230_0, i_13_344_267_0, i_13_344_274_0,
    i_13_344_275_0, i_13_344_320_0, i_13_344_382_0, i_13_344_409_0,
    i_13_344_410_0, i_13_344_418_0, i_13_344_454_0, i_13_344_466_0,
    i_13_344_528_0, i_13_344_562_0, i_13_344_589_0, i_13_344_590_0,
    i_13_344_591_0, i_13_344_597_0, i_13_344_625_0, i_13_344_646_0,
    i_13_344_688_0, i_13_344_718_0, i_13_344_760_0, i_13_344_761_0,
    i_13_344_824_0, i_13_344_839_0, i_13_344_843_0, i_13_344_915_0,
    i_13_344_949_0, i_13_344_1208_0, i_13_344_1211_0, i_13_344_1274_0,
    i_13_344_1307_0, i_13_344_1310_0, i_13_344_1348_0, i_13_344_1391_0,
    i_13_344_1531_0, i_13_344_1597_0, i_13_344_1598_0, i_13_344_1624_0,
    i_13_344_1640_0, i_13_344_1643_0, i_13_344_1646_0, i_13_344_1670_0,
    i_13_344_1886_0, i_13_344_1938_0, i_13_344_2138_0, i_13_344_2140_0,
    i_13_344_2192_0, i_13_344_2209_0, i_13_344_2248_0, i_13_344_2363_0,
    i_13_344_2434_0, i_13_344_2542_0, i_13_344_2550_0, i_13_344_2551_0,
    i_13_344_2552_0, i_13_344_2623_0, i_13_344_2651_0, i_13_344_2678_0,
    i_13_344_2821_0, i_13_344_2822_0, i_13_344_2857_0, i_13_344_2998_0,
    i_13_344_3108_0, i_13_344_3109_0, i_13_344_3110_0, i_13_344_3116_0,
    i_13_344_3163_0, i_13_344_3235_0, i_13_344_3269_0, i_13_344_3323_0,
    i_13_344_3361_0, i_13_344_3370_0, i_13_344_3388_0, i_13_344_3389_0,
    i_13_344_3391_0, i_13_344_3491_0, i_13_344_3595_0, i_13_344_3633_0,
    i_13_344_3668_0, i_13_344_3685_0, i_13_344_3767_0, i_13_344_3882_0,
    i_13_344_4036_0, i_13_344_4037_0, i_13_344_4055_0, i_13_344_4162_0,
    i_13_344_4262_0, i_13_344_4351_0, i_13_344_4372_0, i_13_344_4397_0,
    i_13_344_4451_0, i_13_344_4559_0, i_13_344_4567_0, i_13_344_4596_0,
    o_13_344_0_0  );
  input  i_13_344_112_0, i_13_344_121_0, i_13_344_122_0, i_13_344_139_0,
    i_13_344_193_0, i_13_344_230_0, i_13_344_267_0, i_13_344_274_0,
    i_13_344_275_0, i_13_344_320_0, i_13_344_382_0, i_13_344_409_0,
    i_13_344_410_0, i_13_344_418_0, i_13_344_454_0, i_13_344_466_0,
    i_13_344_528_0, i_13_344_562_0, i_13_344_589_0, i_13_344_590_0,
    i_13_344_591_0, i_13_344_597_0, i_13_344_625_0, i_13_344_646_0,
    i_13_344_688_0, i_13_344_718_0, i_13_344_760_0, i_13_344_761_0,
    i_13_344_824_0, i_13_344_839_0, i_13_344_843_0, i_13_344_915_0,
    i_13_344_949_0, i_13_344_1208_0, i_13_344_1211_0, i_13_344_1274_0,
    i_13_344_1307_0, i_13_344_1310_0, i_13_344_1348_0, i_13_344_1391_0,
    i_13_344_1531_0, i_13_344_1597_0, i_13_344_1598_0, i_13_344_1624_0,
    i_13_344_1640_0, i_13_344_1643_0, i_13_344_1646_0, i_13_344_1670_0,
    i_13_344_1886_0, i_13_344_1938_0, i_13_344_2138_0, i_13_344_2140_0,
    i_13_344_2192_0, i_13_344_2209_0, i_13_344_2248_0, i_13_344_2363_0,
    i_13_344_2434_0, i_13_344_2542_0, i_13_344_2550_0, i_13_344_2551_0,
    i_13_344_2552_0, i_13_344_2623_0, i_13_344_2651_0, i_13_344_2678_0,
    i_13_344_2821_0, i_13_344_2822_0, i_13_344_2857_0, i_13_344_2998_0,
    i_13_344_3108_0, i_13_344_3109_0, i_13_344_3110_0, i_13_344_3116_0,
    i_13_344_3163_0, i_13_344_3235_0, i_13_344_3269_0, i_13_344_3323_0,
    i_13_344_3361_0, i_13_344_3370_0, i_13_344_3388_0, i_13_344_3389_0,
    i_13_344_3391_0, i_13_344_3491_0, i_13_344_3595_0, i_13_344_3633_0,
    i_13_344_3668_0, i_13_344_3685_0, i_13_344_3767_0, i_13_344_3882_0,
    i_13_344_4036_0, i_13_344_4037_0, i_13_344_4055_0, i_13_344_4162_0,
    i_13_344_4262_0, i_13_344_4351_0, i_13_344_4372_0, i_13_344_4397_0,
    i_13_344_4451_0, i_13_344_4559_0, i_13_344_4567_0, i_13_344_4596_0;
  output o_13_344_0_0;
  assign o_13_344_0_0 = ~((i_13_344_949_0 & (i_13_344_3235_0 | (i_13_344_1598_0 & ~i_13_344_2857_0 & ~i_13_344_3163_0))) | i_13_344_3767_0 | ~i_13_344_4037_0 | (~i_13_344_1208_0 & ~i_13_344_4262_0 & ~i_13_344_4397_0) | (~i_13_344_1640_0 & i_13_344_4262_0 & i_13_344_4559_0));
endmodule



// Benchmark "kernel_13_345" written by ABC on Sun Jul 19 10:50:12 2020

module kernel_13_345 ( 
    i_13_345_48_0, i_13_345_61_0, i_13_345_93_0, i_13_345_106_0,
    i_13_345_136_0, i_13_345_259_0, i_13_345_492_0, i_13_345_619_0,
    i_13_345_624_0, i_13_345_625_0, i_13_345_627_0, i_13_345_673_0,
    i_13_345_697_0, i_13_345_707_0, i_13_345_823_0, i_13_345_825_0,
    i_13_345_826_0, i_13_345_948_0, i_13_345_978_0, i_13_345_979_0,
    i_13_345_1024_0, i_13_345_1072_0, i_13_345_1095_0, i_13_345_1102_0,
    i_13_345_1200_0, i_13_345_1279_0, i_13_345_1303_0, i_13_345_1320_0,
    i_13_345_1321_0, i_13_345_1428_0, i_13_345_1434_0, i_13_345_1444_0,
    i_13_345_1464_0, i_13_345_1465_0, i_13_345_1480_0, i_13_345_1483_0,
    i_13_345_1547_0, i_13_345_1572_0, i_13_345_1752_0, i_13_345_1757_0,
    i_13_345_1786_0, i_13_345_1807_0, i_13_345_1911_0, i_13_345_1960_0,
    i_13_345_2010_0, i_13_345_2103_0, i_13_345_2238_0, i_13_345_2244_0,
    i_13_345_2245_0, i_13_345_2263_0, i_13_345_2343_0, i_13_345_2424_0,
    i_13_345_2442_0, i_13_345_2443_0, i_13_345_2445_0, i_13_345_2446_0,
    i_13_345_2454_0, i_13_345_2554_0, i_13_345_2743_0, i_13_345_2752_0,
    i_13_345_2823_0, i_13_345_2824_0, i_13_345_2857_0, i_13_345_2883_0,
    i_13_345_3073_0, i_13_345_3135_0, i_13_345_3153_0, i_13_345_3310_0,
    i_13_345_3345_0, i_13_345_3381_0, i_13_345_3418_0, i_13_345_3432_0,
    i_13_345_3437_0, i_13_345_3475_0, i_13_345_3489_0, i_13_345_3594_0,
    i_13_345_3618_0, i_13_345_3622_0, i_13_345_3766_0, i_13_345_3786_0,
    i_13_345_3874_0, i_13_345_3936_0, i_13_345_3937_0, i_13_345_4018_0,
    i_13_345_4209_0, i_13_345_4210_0, i_13_345_4237_0, i_13_345_4330_0,
    i_13_345_4332_0, i_13_345_4333_0, i_13_345_4341_0, i_13_345_4344_0,
    i_13_345_4351_0, i_13_345_4381_0, i_13_345_4396_0, i_13_345_4452_0,
    i_13_345_4453_0, i_13_345_4509_0, i_13_345_4567_0, i_13_345_4587_0,
    o_13_345_0_0  );
  input  i_13_345_48_0, i_13_345_61_0, i_13_345_93_0, i_13_345_106_0,
    i_13_345_136_0, i_13_345_259_0, i_13_345_492_0, i_13_345_619_0,
    i_13_345_624_0, i_13_345_625_0, i_13_345_627_0, i_13_345_673_0,
    i_13_345_697_0, i_13_345_707_0, i_13_345_823_0, i_13_345_825_0,
    i_13_345_826_0, i_13_345_948_0, i_13_345_978_0, i_13_345_979_0,
    i_13_345_1024_0, i_13_345_1072_0, i_13_345_1095_0, i_13_345_1102_0,
    i_13_345_1200_0, i_13_345_1279_0, i_13_345_1303_0, i_13_345_1320_0,
    i_13_345_1321_0, i_13_345_1428_0, i_13_345_1434_0, i_13_345_1444_0,
    i_13_345_1464_0, i_13_345_1465_0, i_13_345_1480_0, i_13_345_1483_0,
    i_13_345_1547_0, i_13_345_1572_0, i_13_345_1752_0, i_13_345_1757_0,
    i_13_345_1786_0, i_13_345_1807_0, i_13_345_1911_0, i_13_345_1960_0,
    i_13_345_2010_0, i_13_345_2103_0, i_13_345_2238_0, i_13_345_2244_0,
    i_13_345_2245_0, i_13_345_2263_0, i_13_345_2343_0, i_13_345_2424_0,
    i_13_345_2442_0, i_13_345_2443_0, i_13_345_2445_0, i_13_345_2446_0,
    i_13_345_2454_0, i_13_345_2554_0, i_13_345_2743_0, i_13_345_2752_0,
    i_13_345_2823_0, i_13_345_2824_0, i_13_345_2857_0, i_13_345_2883_0,
    i_13_345_3073_0, i_13_345_3135_0, i_13_345_3153_0, i_13_345_3310_0,
    i_13_345_3345_0, i_13_345_3381_0, i_13_345_3418_0, i_13_345_3432_0,
    i_13_345_3437_0, i_13_345_3475_0, i_13_345_3489_0, i_13_345_3594_0,
    i_13_345_3618_0, i_13_345_3622_0, i_13_345_3766_0, i_13_345_3786_0,
    i_13_345_3874_0, i_13_345_3936_0, i_13_345_3937_0, i_13_345_4018_0,
    i_13_345_4209_0, i_13_345_4210_0, i_13_345_4237_0, i_13_345_4330_0,
    i_13_345_4332_0, i_13_345_4333_0, i_13_345_4341_0, i_13_345_4344_0,
    i_13_345_4351_0, i_13_345_4381_0, i_13_345_4396_0, i_13_345_4452_0,
    i_13_345_4453_0, i_13_345_4509_0, i_13_345_4567_0, i_13_345_4587_0;
  output o_13_345_0_0;
  assign o_13_345_0_0 = ~((~i_13_345_2446_0 & ((~i_13_345_61_0 & ~i_13_345_2445_0) | (~i_13_345_3489_0 & ~i_13_345_3622_0))) | (~i_13_345_106_0 & ~i_13_345_2244_0 & ~i_13_345_2245_0 & ~i_13_345_4333_0) | (i_13_345_259_0 & ~i_13_345_1483_0 & ~i_13_345_4452_0));
endmodule



// Benchmark "kernel_13_346" written by ABC on Sun Jul 19 10:50:13 2020

module kernel_13_346 ( 
    i_13_346_40_0, i_13_346_117_0, i_13_346_121_0, i_13_346_162_0,
    i_13_346_166_0, i_13_346_183_0, i_13_346_189_0, i_13_346_192_0,
    i_13_346_283_0, i_13_346_315_0, i_13_346_333_0, i_13_346_454_0,
    i_13_346_517_0, i_13_346_532_0, i_13_346_576_0, i_13_346_661_0,
    i_13_346_714_0, i_13_346_760_0, i_13_346_862_0, i_13_346_927_0,
    i_13_346_948_0, i_13_346_1098_0, i_13_346_1135_0, i_13_346_1227_0,
    i_13_346_1254_0, i_13_346_1259_0, i_13_346_1261_0, i_13_346_1279_0,
    i_13_346_1407_0, i_13_346_1430_0, i_13_346_1458_0, i_13_346_1468_0,
    i_13_346_1479_0, i_13_346_1488_0, i_13_346_1507_0, i_13_346_1522_0,
    i_13_346_1570_0, i_13_346_1597_0, i_13_346_1624_0, i_13_346_1647_0,
    i_13_346_1685_0, i_13_346_1710_0, i_13_346_1723_0, i_13_346_1767_0,
    i_13_346_1771_0, i_13_346_1782_0, i_13_346_1786_0, i_13_346_1800_0,
    i_13_346_1939_0, i_13_346_2011_0, i_13_346_2056_0, i_13_346_2100_0,
    i_13_346_2115_0, i_13_346_2208_0, i_13_346_2209_0, i_13_346_2223_0,
    i_13_346_2224_0, i_13_346_2235_0, i_13_346_2236_0, i_13_346_2358_0,
    i_13_346_2394_0, i_13_346_2407_0, i_13_346_2438_0, i_13_346_2457_0,
    i_13_346_2532_0, i_13_346_2565_0, i_13_346_2595_0, i_13_346_2835_0,
    i_13_346_2902_0, i_13_346_3036_0, i_13_346_3136_0, i_13_346_3216_0,
    i_13_346_3217_0, i_13_346_3221_0, i_13_346_3286_0, i_13_346_3339_0,
    i_13_346_3369_0, i_13_346_3414_0, i_13_346_3424_0, i_13_346_3429_0,
    i_13_346_3468_0, i_13_346_3549_0, i_13_346_3613_0, i_13_346_3699_0,
    i_13_346_3855_0, i_13_346_3873_0, i_13_346_3877_0, i_13_346_3883_0,
    i_13_346_3982_0, i_13_346_4008_0, i_13_346_4009_0, i_13_346_4260_0,
    i_13_346_4261_0, i_13_346_4297_0, i_13_346_4360_0, i_13_346_4518_0,
    i_13_346_4527_0, i_13_346_4530_0, i_13_346_4540_0, i_13_346_4594_0,
    o_13_346_0_0  );
  input  i_13_346_40_0, i_13_346_117_0, i_13_346_121_0, i_13_346_162_0,
    i_13_346_166_0, i_13_346_183_0, i_13_346_189_0, i_13_346_192_0,
    i_13_346_283_0, i_13_346_315_0, i_13_346_333_0, i_13_346_454_0,
    i_13_346_517_0, i_13_346_532_0, i_13_346_576_0, i_13_346_661_0,
    i_13_346_714_0, i_13_346_760_0, i_13_346_862_0, i_13_346_927_0,
    i_13_346_948_0, i_13_346_1098_0, i_13_346_1135_0, i_13_346_1227_0,
    i_13_346_1254_0, i_13_346_1259_0, i_13_346_1261_0, i_13_346_1279_0,
    i_13_346_1407_0, i_13_346_1430_0, i_13_346_1458_0, i_13_346_1468_0,
    i_13_346_1479_0, i_13_346_1488_0, i_13_346_1507_0, i_13_346_1522_0,
    i_13_346_1570_0, i_13_346_1597_0, i_13_346_1624_0, i_13_346_1647_0,
    i_13_346_1685_0, i_13_346_1710_0, i_13_346_1723_0, i_13_346_1767_0,
    i_13_346_1771_0, i_13_346_1782_0, i_13_346_1786_0, i_13_346_1800_0,
    i_13_346_1939_0, i_13_346_2011_0, i_13_346_2056_0, i_13_346_2100_0,
    i_13_346_2115_0, i_13_346_2208_0, i_13_346_2209_0, i_13_346_2223_0,
    i_13_346_2224_0, i_13_346_2235_0, i_13_346_2236_0, i_13_346_2358_0,
    i_13_346_2394_0, i_13_346_2407_0, i_13_346_2438_0, i_13_346_2457_0,
    i_13_346_2532_0, i_13_346_2565_0, i_13_346_2595_0, i_13_346_2835_0,
    i_13_346_2902_0, i_13_346_3036_0, i_13_346_3136_0, i_13_346_3216_0,
    i_13_346_3217_0, i_13_346_3221_0, i_13_346_3286_0, i_13_346_3339_0,
    i_13_346_3369_0, i_13_346_3414_0, i_13_346_3424_0, i_13_346_3429_0,
    i_13_346_3468_0, i_13_346_3549_0, i_13_346_3613_0, i_13_346_3699_0,
    i_13_346_3855_0, i_13_346_3873_0, i_13_346_3877_0, i_13_346_3883_0,
    i_13_346_3982_0, i_13_346_4008_0, i_13_346_4009_0, i_13_346_4260_0,
    i_13_346_4261_0, i_13_346_4297_0, i_13_346_4360_0, i_13_346_4518_0,
    i_13_346_4527_0, i_13_346_4530_0, i_13_346_4540_0, i_13_346_4594_0;
  output o_13_346_0_0;
  assign o_13_346_0_0 = ~(~i_13_346_2208_0 | ~i_13_346_3982_0 | (i_13_346_1597_0 & ~i_13_346_3549_0) | (~i_13_346_2236_0 & i_13_346_3549_0) | (~i_13_346_1488_0 & ~i_13_346_1710_0));
endmodule



// Benchmark "kernel_13_347" written by ABC on Sun Jul 19 10:50:14 2020

module kernel_13_347 ( 
    i_13_347_161_0, i_13_347_232_0, i_13_347_242_0, i_13_347_285_0,
    i_13_347_359_0, i_13_347_412_0, i_13_347_469_0, i_13_347_503_0,
    i_13_347_526_0, i_13_347_528_0, i_13_347_529_0, i_13_347_535_0,
    i_13_347_706_0, i_13_347_843_0, i_13_347_853_0, i_13_347_882_0,
    i_13_347_895_0, i_13_347_897_0, i_13_347_1024_0, i_13_347_1203_0,
    i_13_347_1309_0, i_13_347_1310_0, i_13_347_1312_0, i_13_347_1390_0,
    i_13_347_1426_0, i_13_347_1428_0, i_13_347_1438_0, i_13_347_1496_0,
    i_13_347_1500_0, i_13_347_1501_0, i_13_347_1550_0, i_13_347_1552_0,
    i_13_347_1574_0, i_13_347_1631_0, i_13_347_1723_0, i_13_347_1726_0,
    i_13_347_1786_0, i_13_347_1834_0, i_13_347_1917_0, i_13_347_1950_0,
    i_13_347_2004_0, i_13_347_2033_0, i_13_347_2114_0, i_13_347_2200_0,
    i_13_347_2201_0, i_13_347_2202_0, i_13_347_2263_0, i_13_347_2407_0,
    i_13_347_2449_0, i_13_347_2452_0, i_13_347_2454_0, i_13_347_2455_0,
    i_13_347_2721_0, i_13_347_2764_0, i_13_347_2767_0, i_13_347_2924_0,
    i_13_347_3012_0, i_13_347_3163_0, i_13_347_3217_0, i_13_347_3323_0,
    i_13_347_3373_0, i_13_347_3460_0, i_13_347_3464_0, i_13_347_3533_0,
    i_13_347_3539_0, i_13_347_3545_0, i_13_347_3579_0, i_13_347_3581_0,
    i_13_347_3597_0, i_13_347_3623_0, i_13_347_3635_0, i_13_347_3646_0,
    i_13_347_3666_0, i_13_347_3669_0, i_13_347_3730_0, i_13_347_3731_0,
    i_13_347_3733_0, i_13_347_3734_0, i_13_347_3786_0, i_13_347_3787_0,
    i_13_347_3856_0, i_13_347_3865_0, i_13_347_3892_0, i_13_347_3931_0,
    i_13_347_4016_0, i_13_347_4081_0, i_13_347_4234_0, i_13_347_4252_0,
    i_13_347_4253_0, i_13_347_4261_0, i_13_347_4263_0, i_13_347_4264_0,
    i_13_347_4279_0, i_13_347_4369_0, i_13_347_4380_0, i_13_347_4435_0,
    i_13_347_4452_0, i_13_347_4554_0, i_13_347_4555_0, i_13_347_4558_0,
    o_13_347_0_0  );
  input  i_13_347_161_0, i_13_347_232_0, i_13_347_242_0, i_13_347_285_0,
    i_13_347_359_0, i_13_347_412_0, i_13_347_469_0, i_13_347_503_0,
    i_13_347_526_0, i_13_347_528_0, i_13_347_529_0, i_13_347_535_0,
    i_13_347_706_0, i_13_347_843_0, i_13_347_853_0, i_13_347_882_0,
    i_13_347_895_0, i_13_347_897_0, i_13_347_1024_0, i_13_347_1203_0,
    i_13_347_1309_0, i_13_347_1310_0, i_13_347_1312_0, i_13_347_1390_0,
    i_13_347_1426_0, i_13_347_1428_0, i_13_347_1438_0, i_13_347_1496_0,
    i_13_347_1500_0, i_13_347_1501_0, i_13_347_1550_0, i_13_347_1552_0,
    i_13_347_1574_0, i_13_347_1631_0, i_13_347_1723_0, i_13_347_1726_0,
    i_13_347_1786_0, i_13_347_1834_0, i_13_347_1917_0, i_13_347_1950_0,
    i_13_347_2004_0, i_13_347_2033_0, i_13_347_2114_0, i_13_347_2200_0,
    i_13_347_2201_0, i_13_347_2202_0, i_13_347_2263_0, i_13_347_2407_0,
    i_13_347_2449_0, i_13_347_2452_0, i_13_347_2454_0, i_13_347_2455_0,
    i_13_347_2721_0, i_13_347_2764_0, i_13_347_2767_0, i_13_347_2924_0,
    i_13_347_3012_0, i_13_347_3163_0, i_13_347_3217_0, i_13_347_3323_0,
    i_13_347_3373_0, i_13_347_3460_0, i_13_347_3464_0, i_13_347_3533_0,
    i_13_347_3539_0, i_13_347_3545_0, i_13_347_3579_0, i_13_347_3581_0,
    i_13_347_3597_0, i_13_347_3623_0, i_13_347_3635_0, i_13_347_3646_0,
    i_13_347_3666_0, i_13_347_3669_0, i_13_347_3730_0, i_13_347_3731_0,
    i_13_347_3733_0, i_13_347_3734_0, i_13_347_3786_0, i_13_347_3787_0,
    i_13_347_3856_0, i_13_347_3865_0, i_13_347_3892_0, i_13_347_3931_0,
    i_13_347_4016_0, i_13_347_4081_0, i_13_347_4234_0, i_13_347_4252_0,
    i_13_347_4253_0, i_13_347_4261_0, i_13_347_4263_0, i_13_347_4264_0,
    i_13_347_4279_0, i_13_347_4369_0, i_13_347_4380_0, i_13_347_4435_0,
    i_13_347_4452_0, i_13_347_4554_0, i_13_347_4555_0, i_13_347_4558_0;
  output o_13_347_0_0;
  assign o_13_347_0_0 = ~(~i_13_347_3579_0 | ~i_13_347_2767_0 | (~i_13_347_2454_0 & ~i_13_347_3892_0 & ~i_13_347_4264_0));
endmodule



// Benchmark "kernel_13_348" written by ABC on Sun Jul 19 10:50:14 2020

module kernel_13_348 ( 
    i_13_348_49_0, i_13_348_76_0, i_13_348_77_0, i_13_348_100_0,
    i_13_348_329_0, i_13_348_353_0, i_13_348_356_0, i_13_348_409_0,
    i_13_348_410_0, i_13_348_419_0, i_13_348_529_0, i_13_348_530_0,
    i_13_348_562_0, i_13_348_611_0, i_13_348_698_0, i_13_348_742_0,
    i_13_348_827_0, i_13_348_853_0, i_13_348_854_0, i_13_348_953_0,
    i_13_348_1025_0, i_13_348_1076_0, i_13_348_1109_0, i_13_348_1142_0,
    i_13_348_1232_0, i_13_348_1305_0, i_13_348_1309_0, i_13_348_1310_0,
    i_13_348_1313_0, i_13_348_1321_0, i_13_348_1322_0, i_13_348_1330_0,
    i_13_348_1430_0, i_13_348_1444_0, i_13_348_1462_0, i_13_348_1493_0,
    i_13_348_1552_0, i_13_348_1553_0, i_13_348_1694_0, i_13_348_1723_0,
    i_13_348_1741_0, i_13_348_1771_0, i_13_348_1777_0, i_13_348_1846_0,
    i_13_348_1889_0, i_13_348_1948_0, i_13_348_1951_0, i_13_348_1961_0,
    i_13_348_2011_0, i_13_348_2033_0, i_13_348_2141_0, i_13_348_2203_0,
    i_13_348_2236_0, i_13_348_2237_0, i_13_348_2282_0, i_13_348_2354_0,
    i_13_348_2402_0, i_13_348_2428_0, i_13_348_2546_0, i_13_348_2596_0,
    i_13_348_2654_0, i_13_348_2923_0, i_13_348_2924_0, i_13_348_3013_0,
    i_13_348_3014_0, i_13_348_3016_0, i_13_348_3034_0, i_13_348_3071_0,
    i_13_348_3197_0, i_13_348_3274_0, i_13_348_3419_0, i_13_348_3427_0,
    i_13_348_3442_0, i_13_348_3542_0, i_13_348_3544_0, i_13_348_3580_0,
    i_13_348_3595_0, i_13_348_3726_0, i_13_348_3730_0, i_13_348_3734_0,
    i_13_348_3787_0, i_13_348_3788_0, i_13_348_3806_0, i_13_348_3896_0,
    i_13_348_3913_0, i_13_348_3914_0, i_13_348_3929_0, i_13_348_3938_0,
    i_13_348_4060_0, i_13_348_4238_0, i_13_348_4256_0, i_13_348_4264_0,
    i_13_348_4265_0, i_13_348_4334_0, i_13_348_4381_0, i_13_348_4382_0,
    i_13_348_4450_0, i_13_348_4454_0, i_13_348_4478_0, i_13_348_4600_0,
    o_13_348_0_0  );
  input  i_13_348_49_0, i_13_348_76_0, i_13_348_77_0, i_13_348_100_0,
    i_13_348_329_0, i_13_348_353_0, i_13_348_356_0, i_13_348_409_0,
    i_13_348_410_0, i_13_348_419_0, i_13_348_529_0, i_13_348_530_0,
    i_13_348_562_0, i_13_348_611_0, i_13_348_698_0, i_13_348_742_0,
    i_13_348_827_0, i_13_348_853_0, i_13_348_854_0, i_13_348_953_0,
    i_13_348_1025_0, i_13_348_1076_0, i_13_348_1109_0, i_13_348_1142_0,
    i_13_348_1232_0, i_13_348_1305_0, i_13_348_1309_0, i_13_348_1310_0,
    i_13_348_1313_0, i_13_348_1321_0, i_13_348_1322_0, i_13_348_1330_0,
    i_13_348_1430_0, i_13_348_1444_0, i_13_348_1462_0, i_13_348_1493_0,
    i_13_348_1552_0, i_13_348_1553_0, i_13_348_1694_0, i_13_348_1723_0,
    i_13_348_1741_0, i_13_348_1771_0, i_13_348_1777_0, i_13_348_1846_0,
    i_13_348_1889_0, i_13_348_1948_0, i_13_348_1951_0, i_13_348_1961_0,
    i_13_348_2011_0, i_13_348_2033_0, i_13_348_2141_0, i_13_348_2203_0,
    i_13_348_2236_0, i_13_348_2237_0, i_13_348_2282_0, i_13_348_2354_0,
    i_13_348_2402_0, i_13_348_2428_0, i_13_348_2546_0, i_13_348_2596_0,
    i_13_348_2654_0, i_13_348_2923_0, i_13_348_2924_0, i_13_348_3013_0,
    i_13_348_3014_0, i_13_348_3016_0, i_13_348_3034_0, i_13_348_3071_0,
    i_13_348_3197_0, i_13_348_3274_0, i_13_348_3419_0, i_13_348_3427_0,
    i_13_348_3442_0, i_13_348_3542_0, i_13_348_3544_0, i_13_348_3580_0,
    i_13_348_3595_0, i_13_348_3726_0, i_13_348_3730_0, i_13_348_3734_0,
    i_13_348_3787_0, i_13_348_3788_0, i_13_348_3806_0, i_13_348_3896_0,
    i_13_348_3913_0, i_13_348_3914_0, i_13_348_3929_0, i_13_348_3938_0,
    i_13_348_4060_0, i_13_348_4238_0, i_13_348_4256_0, i_13_348_4264_0,
    i_13_348_4265_0, i_13_348_4334_0, i_13_348_4381_0, i_13_348_4382_0,
    i_13_348_4450_0, i_13_348_4454_0, i_13_348_4478_0, i_13_348_4600_0;
  output o_13_348_0_0;
  assign o_13_348_0_0 = ~((~i_13_348_3914_0 & ~i_13_348_4238_0 & ~i_13_348_4454_0) | (~i_13_348_2033_0 & ~i_13_348_3896_0 & ~i_13_348_4381_0));
endmodule



// Benchmark "kernel_13_349" written by ABC on Sun Jul 19 10:50:15 2020

module kernel_13_349 ( 
    i_13_349_205_0, i_13_349_210_0, i_13_349_285_0, i_13_349_363_0,
    i_13_349_417_0, i_13_349_465_0, i_13_349_520_0, i_13_349_525_0,
    i_13_349_528_0, i_13_349_529_0, i_13_349_537_0, i_13_349_690_0,
    i_13_349_736_0, i_13_349_825_0, i_13_349_852_0, i_13_349_853_0,
    i_13_349_1020_0, i_13_349_1023_0, i_13_349_1024_0, i_13_349_1075_0,
    i_13_349_1120_0, i_13_349_1131_0, i_13_349_1212_0, i_13_349_1311_0,
    i_13_349_1312_0, i_13_349_1317_0, i_13_349_1320_0, i_13_349_1461_0,
    i_13_349_1498_0, i_13_349_1551_0, i_13_349_1552_0, i_13_349_1554_0,
    i_13_349_1555_0, i_13_349_1605_0, i_13_349_1699_0, i_13_349_1749_0,
    i_13_349_1906_0, i_13_349_1920_0, i_13_349_1932_0, i_13_349_1941_0,
    i_13_349_1959_0, i_13_349_1960_0, i_13_349_2032_0, i_13_349_2127_0,
    i_13_349_2136_0, i_13_349_2139_0, i_13_349_2199_0, i_13_349_2202_0,
    i_13_349_2454_0, i_13_349_2491_0, i_13_349_2506_0, i_13_349_2572_0,
    i_13_349_2677_0, i_13_349_3012_0, i_13_349_3013_0, i_13_349_3103_0,
    i_13_349_3118_0, i_13_349_3156_0, i_13_349_3172_0, i_13_349_3271_0,
    i_13_349_3378_0, i_13_349_3432_0, i_13_349_3453_0, i_13_349_3460_0,
    i_13_349_3478_0, i_13_349_3505_0, i_13_349_3540_0, i_13_349_3541_0,
    i_13_349_3543_0, i_13_349_3571_0, i_13_349_3579_0, i_13_349_3580_0,
    i_13_349_3597_0, i_13_349_3633_0, i_13_349_3669_0, i_13_349_3670_0,
    i_13_349_3729_0, i_13_349_3732_0, i_13_349_3733_0, i_13_349_3786_0,
    i_13_349_3787_0, i_13_349_3805_0, i_13_349_3858_0, i_13_349_3912_0,
    i_13_349_3918_0, i_13_349_3919_0, i_13_349_3985_0, i_13_349_4039_0,
    i_13_349_4120_0, i_13_349_4164_0, i_13_349_4254_0, i_13_349_4255_0,
    i_13_349_4260_0, i_13_349_4341_0, i_13_349_4351_0, i_13_349_4354_0,
    i_13_349_4378_0, i_13_349_4380_0, i_13_349_4381_0, i_13_349_4578_0,
    o_13_349_0_0  );
  input  i_13_349_205_0, i_13_349_210_0, i_13_349_285_0, i_13_349_363_0,
    i_13_349_417_0, i_13_349_465_0, i_13_349_520_0, i_13_349_525_0,
    i_13_349_528_0, i_13_349_529_0, i_13_349_537_0, i_13_349_690_0,
    i_13_349_736_0, i_13_349_825_0, i_13_349_852_0, i_13_349_853_0,
    i_13_349_1020_0, i_13_349_1023_0, i_13_349_1024_0, i_13_349_1075_0,
    i_13_349_1120_0, i_13_349_1131_0, i_13_349_1212_0, i_13_349_1311_0,
    i_13_349_1312_0, i_13_349_1317_0, i_13_349_1320_0, i_13_349_1461_0,
    i_13_349_1498_0, i_13_349_1551_0, i_13_349_1552_0, i_13_349_1554_0,
    i_13_349_1555_0, i_13_349_1605_0, i_13_349_1699_0, i_13_349_1749_0,
    i_13_349_1906_0, i_13_349_1920_0, i_13_349_1932_0, i_13_349_1941_0,
    i_13_349_1959_0, i_13_349_1960_0, i_13_349_2032_0, i_13_349_2127_0,
    i_13_349_2136_0, i_13_349_2139_0, i_13_349_2199_0, i_13_349_2202_0,
    i_13_349_2454_0, i_13_349_2491_0, i_13_349_2506_0, i_13_349_2572_0,
    i_13_349_2677_0, i_13_349_3012_0, i_13_349_3013_0, i_13_349_3103_0,
    i_13_349_3118_0, i_13_349_3156_0, i_13_349_3172_0, i_13_349_3271_0,
    i_13_349_3378_0, i_13_349_3432_0, i_13_349_3453_0, i_13_349_3460_0,
    i_13_349_3478_0, i_13_349_3505_0, i_13_349_3540_0, i_13_349_3541_0,
    i_13_349_3543_0, i_13_349_3571_0, i_13_349_3579_0, i_13_349_3580_0,
    i_13_349_3597_0, i_13_349_3633_0, i_13_349_3669_0, i_13_349_3670_0,
    i_13_349_3729_0, i_13_349_3732_0, i_13_349_3733_0, i_13_349_3786_0,
    i_13_349_3787_0, i_13_349_3805_0, i_13_349_3858_0, i_13_349_3912_0,
    i_13_349_3918_0, i_13_349_3919_0, i_13_349_3985_0, i_13_349_4039_0,
    i_13_349_4120_0, i_13_349_4164_0, i_13_349_4254_0, i_13_349_4255_0,
    i_13_349_4260_0, i_13_349_4341_0, i_13_349_4351_0, i_13_349_4354_0,
    i_13_349_4378_0, i_13_349_4380_0, i_13_349_4381_0, i_13_349_4578_0;
  output o_13_349_0_0;
  assign o_13_349_0_0 = ~((~i_13_349_3543_0 & ((~i_13_349_1212_0 & ~i_13_349_3579_0) | (i_13_349_528_0 & ~i_13_349_3633_0))) | ~i_13_349_1555_0 | (~i_13_349_3579_0 & ~i_13_349_3858_0) | (i_13_349_3103_0 & ~i_13_349_3786_0 & ~i_13_349_4380_0 & ~i_13_349_4381_0));
endmodule



// Benchmark "kernel_13_350" written by ABC on Sun Jul 19 10:50:16 2020

module kernel_13_350 ( 
    i_13_350_31_0, i_13_350_46_0, i_13_350_47_0, i_13_350_163_0,
    i_13_350_164_0, i_13_350_173_0, i_13_350_174_0, i_13_350_245_0,
    i_13_350_273_0, i_13_350_299_0, i_13_350_326_0, i_13_350_415_0,
    i_13_350_416_0, i_13_350_518_0, i_13_350_533_0, i_13_350_568_0,
    i_13_350_626_0, i_13_350_658_0, i_13_350_659_0, i_13_350_688_0,
    i_13_350_721_0, i_13_350_757_0, i_13_350_758_0, i_13_350_761_0,
    i_13_350_848_0, i_13_350_856_0, i_13_350_937_0, i_13_350_938_0,
    i_13_350_1023_0, i_13_350_1072_0, i_13_350_1073_0, i_13_350_1129_0,
    i_13_350_1130_0, i_13_350_1201_0, i_13_350_1219_0, i_13_350_1252_0,
    i_13_350_1253_0, i_13_350_1280_0, i_13_350_1445_0, i_13_350_1495_0,
    i_13_350_1522_0, i_13_350_1523_0, i_13_350_1535_0, i_13_350_1549_0,
    i_13_350_1550_0, i_13_350_1603_0, i_13_350_1604_0, i_13_350_1725_0,
    i_13_350_1751_0, i_13_350_1946_0, i_13_350_1991_0, i_13_350_2026_0,
    i_13_350_2027_0, i_13_350_2116_0, i_13_350_2297_0, i_13_350_2425_0,
    i_13_350_2443_0, i_13_350_2471_0, i_13_350_2472_0, i_13_350_2539_0,
    i_13_350_2540_0, i_13_350_2722_0, i_13_350_2724_0, i_13_350_2801_0,
    i_13_350_2920_0, i_13_350_2981_0, i_13_350_3000_0, i_13_350_3001_0,
    i_13_350_3003_0, i_13_350_3007_0, i_13_350_3029_0, i_13_350_3124_0,
    i_13_350_3215_0, i_13_350_3218_0, i_13_350_3262_0, i_13_350_3457_0,
    i_13_350_3458_0, i_13_350_3485_0, i_13_350_3538_0, i_13_350_3539_0,
    i_13_350_3547_0, i_13_350_3575_0, i_13_350_3638_0, i_13_350_3818_0,
    i_13_350_3822_0, i_13_350_3844_0, i_13_350_3894_0, i_13_350_3898_0,
    i_13_350_3899_0, i_13_350_3908_0, i_13_350_4018_0, i_13_350_4053_0,
    i_13_350_4061_0, i_13_350_4102_0, i_13_350_4322_0, i_13_350_4331_0,
    i_13_350_4339_0, i_13_350_4511_0, i_13_350_4604_0, i_13_350_4605_0,
    o_13_350_0_0  );
  input  i_13_350_31_0, i_13_350_46_0, i_13_350_47_0, i_13_350_163_0,
    i_13_350_164_0, i_13_350_173_0, i_13_350_174_0, i_13_350_245_0,
    i_13_350_273_0, i_13_350_299_0, i_13_350_326_0, i_13_350_415_0,
    i_13_350_416_0, i_13_350_518_0, i_13_350_533_0, i_13_350_568_0,
    i_13_350_626_0, i_13_350_658_0, i_13_350_659_0, i_13_350_688_0,
    i_13_350_721_0, i_13_350_757_0, i_13_350_758_0, i_13_350_761_0,
    i_13_350_848_0, i_13_350_856_0, i_13_350_937_0, i_13_350_938_0,
    i_13_350_1023_0, i_13_350_1072_0, i_13_350_1073_0, i_13_350_1129_0,
    i_13_350_1130_0, i_13_350_1201_0, i_13_350_1219_0, i_13_350_1252_0,
    i_13_350_1253_0, i_13_350_1280_0, i_13_350_1445_0, i_13_350_1495_0,
    i_13_350_1522_0, i_13_350_1523_0, i_13_350_1535_0, i_13_350_1549_0,
    i_13_350_1550_0, i_13_350_1603_0, i_13_350_1604_0, i_13_350_1725_0,
    i_13_350_1751_0, i_13_350_1946_0, i_13_350_1991_0, i_13_350_2026_0,
    i_13_350_2027_0, i_13_350_2116_0, i_13_350_2297_0, i_13_350_2425_0,
    i_13_350_2443_0, i_13_350_2471_0, i_13_350_2472_0, i_13_350_2539_0,
    i_13_350_2540_0, i_13_350_2722_0, i_13_350_2724_0, i_13_350_2801_0,
    i_13_350_2920_0, i_13_350_2981_0, i_13_350_3000_0, i_13_350_3001_0,
    i_13_350_3003_0, i_13_350_3007_0, i_13_350_3029_0, i_13_350_3124_0,
    i_13_350_3215_0, i_13_350_3218_0, i_13_350_3262_0, i_13_350_3457_0,
    i_13_350_3458_0, i_13_350_3485_0, i_13_350_3538_0, i_13_350_3539_0,
    i_13_350_3547_0, i_13_350_3575_0, i_13_350_3638_0, i_13_350_3818_0,
    i_13_350_3822_0, i_13_350_3844_0, i_13_350_3894_0, i_13_350_3898_0,
    i_13_350_3899_0, i_13_350_3908_0, i_13_350_4018_0, i_13_350_4053_0,
    i_13_350_4061_0, i_13_350_4102_0, i_13_350_4322_0, i_13_350_4331_0,
    i_13_350_4339_0, i_13_350_4511_0, i_13_350_4604_0, i_13_350_4605_0;
  output o_13_350_0_0;
  assign o_13_350_0_0 = ~((~i_13_350_173_0 & ~i_13_350_3457_0 & (~i_13_350_856_0 | ~i_13_350_1751_0)) | ~i_13_350_518_0 | (~i_13_350_326_0 & ~i_13_350_3262_0) | (~i_13_350_568_0 & ~i_13_350_2026_0 & ~i_13_350_4061_0));
endmodule



// Benchmark "kernel_13_351" written by ABC on Sun Jul 19 10:50:17 2020

module kernel_13_351 ( 
    i_13_351_33_0, i_13_351_46_0, i_13_351_160_0, i_13_351_167_0,
    i_13_351_175_0, i_13_351_200_0, i_13_351_238_0, i_13_351_248_0,
    i_13_351_274_0, i_13_351_275_0, i_13_351_277_0, i_13_351_278_0,
    i_13_351_283_0, i_13_351_284_0, i_13_351_315_0, i_13_351_340_0,
    i_13_351_376_0, i_13_351_454_0, i_13_351_457_0, i_13_351_492_0,
    i_13_351_494_0, i_13_351_521_0, i_13_351_565_0, i_13_351_566_0,
    i_13_351_575_0, i_13_351_584_0, i_13_351_615_0, i_13_351_644_0,
    i_13_351_688_0, i_13_351_713_0, i_13_351_741_0, i_13_351_742_0,
    i_13_351_745_0, i_13_351_823_0, i_13_351_824_0, i_13_351_960_0,
    i_13_351_1092_0, i_13_351_1201_0, i_13_351_1221_0, i_13_351_1349_0,
    i_13_351_1400_0, i_13_351_1494_0, i_13_351_1499_0, i_13_351_1715_0,
    i_13_351_1722_0, i_13_351_1770_0, i_13_351_1817_0, i_13_351_1858_0,
    i_13_351_1861_0, i_13_351_1890_0, i_13_351_1920_0, i_13_351_2147_0,
    i_13_351_2300_0, i_13_351_2524_0, i_13_351_2540_0, i_13_351_2651_0,
    i_13_351_2676_0, i_13_351_2721_0, i_13_351_2723_0, i_13_351_2725_0,
    i_13_351_2726_0, i_13_351_2771_0, i_13_351_2785_0, i_13_351_3036_0,
    i_13_351_3076_0, i_13_351_3214_0, i_13_351_3216_0, i_13_351_3218_0,
    i_13_351_3234_0, i_13_351_3235_0, i_13_351_3366_0, i_13_351_3423_0,
    i_13_351_3426_0, i_13_351_3432_0, i_13_351_3461_0, i_13_351_3477_0,
    i_13_351_3549_0, i_13_351_3639_0, i_13_351_3689_0, i_13_351_3723_0,
    i_13_351_3730_0, i_13_351_3858_0, i_13_351_3892_0, i_13_351_3897_0,
    i_13_351_3901_0, i_13_351_3904_0, i_13_351_3923_0, i_13_351_3981_0,
    i_13_351_3986_0, i_13_351_4011_0, i_13_351_4089_0, i_13_351_4163_0,
    i_13_351_4218_0, i_13_351_4261_0, i_13_351_4273_0, i_13_351_4363_0,
    i_13_351_4472_0, i_13_351_4512_0, i_13_351_4569_0, i_13_351_4598_0,
    o_13_351_0_0  );
  input  i_13_351_33_0, i_13_351_46_0, i_13_351_160_0, i_13_351_167_0,
    i_13_351_175_0, i_13_351_200_0, i_13_351_238_0, i_13_351_248_0,
    i_13_351_274_0, i_13_351_275_0, i_13_351_277_0, i_13_351_278_0,
    i_13_351_283_0, i_13_351_284_0, i_13_351_315_0, i_13_351_340_0,
    i_13_351_376_0, i_13_351_454_0, i_13_351_457_0, i_13_351_492_0,
    i_13_351_494_0, i_13_351_521_0, i_13_351_565_0, i_13_351_566_0,
    i_13_351_575_0, i_13_351_584_0, i_13_351_615_0, i_13_351_644_0,
    i_13_351_688_0, i_13_351_713_0, i_13_351_741_0, i_13_351_742_0,
    i_13_351_745_0, i_13_351_823_0, i_13_351_824_0, i_13_351_960_0,
    i_13_351_1092_0, i_13_351_1201_0, i_13_351_1221_0, i_13_351_1349_0,
    i_13_351_1400_0, i_13_351_1494_0, i_13_351_1499_0, i_13_351_1715_0,
    i_13_351_1722_0, i_13_351_1770_0, i_13_351_1817_0, i_13_351_1858_0,
    i_13_351_1861_0, i_13_351_1890_0, i_13_351_1920_0, i_13_351_2147_0,
    i_13_351_2300_0, i_13_351_2524_0, i_13_351_2540_0, i_13_351_2651_0,
    i_13_351_2676_0, i_13_351_2721_0, i_13_351_2723_0, i_13_351_2725_0,
    i_13_351_2726_0, i_13_351_2771_0, i_13_351_2785_0, i_13_351_3036_0,
    i_13_351_3076_0, i_13_351_3214_0, i_13_351_3216_0, i_13_351_3218_0,
    i_13_351_3234_0, i_13_351_3235_0, i_13_351_3366_0, i_13_351_3423_0,
    i_13_351_3426_0, i_13_351_3432_0, i_13_351_3461_0, i_13_351_3477_0,
    i_13_351_3549_0, i_13_351_3639_0, i_13_351_3689_0, i_13_351_3723_0,
    i_13_351_3730_0, i_13_351_3858_0, i_13_351_3892_0, i_13_351_3897_0,
    i_13_351_3901_0, i_13_351_3904_0, i_13_351_3923_0, i_13_351_3981_0,
    i_13_351_3986_0, i_13_351_4011_0, i_13_351_4089_0, i_13_351_4163_0,
    i_13_351_4218_0, i_13_351_4261_0, i_13_351_4273_0, i_13_351_4363_0,
    i_13_351_4472_0, i_13_351_4512_0, i_13_351_4569_0, i_13_351_4598_0;
  output o_13_351_0_0;
  assign o_13_351_0_0 = ~((~i_13_351_238_0 & ((~i_13_351_274_0 & ~i_13_351_1349_0) | (~i_13_351_3218_0 & ~i_13_351_3892_0 & ~i_13_351_3986_0 & ~i_13_351_4569_0))) | (i_13_351_688_0 & ((i_13_351_824_0 & ~i_13_351_2147_0) | (~i_13_351_3218_0 & ~i_13_351_3986_0))) | (~i_13_351_3214_0 & ((~i_13_351_1817_0 & ~i_13_351_2785_0 & ~i_13_351_3036_0 & ~i_13_351_3923_0) | (~i_13_351_2726_0 & ~i_13_351_3461_0 & ~i_13_351_4089_0))) | (~i_13_351_3923_0 & (~i_13_351_3235_0 | (~i_13_351_1499_0 & ~i_13_351_4273_0))) | (i_13_351_283_0 & ~i_13_351_565_0 & i_13_351_4089_0));
endmodule



// Benchmark "kernel_13_352" written by ABC on Sun Jul 19 10:50:18 2020

module kernel_13_352 ( 
    i_13_352_74_0, i_13_352_77_0, i_13_352_137_0, i_13_352_170_0,
    i_13_352_265_0, i_13_352_266_0, i_13_352_283_0, i_13_352_319_0,
    i_13_352_337_0, i_13_352_492_0, i_13_352_518_0, i_13_352_571_0,
    i_13_352_582_0, i_13_352_662_0, i_13_352_688_0, i_13_352_697_0,
    i_13_352_814_0, i_13_352_886_0, i_13_352_888_0, i_13_352_935_0,
    i_13_352_939_0, i_13_352_1066_0, i_13_352_1112_0, i_13_352_1145_0,
    i_13_352_1148_0, i_13_352_1208_0, i_13_352_1210_0, i_13_352_1217_0,
    i_13_352_1226_0, i_13_352_1253_0, i_13_352_1266_0, i_13_352_1426_0,
    i_13_352_1530_0, i_13_352_1633_0, i_13_352_1660_0, i_13_352_1662_0,
    i_13_352_1730_0, i_13_352_1731_0, i_13_352_1733_0, i_13_352_1734_0,
    i_13_352_1849_0, i_13_352_1886_0, i_13_352_2020_0, i_13_352_2021_0,
    i_13_352_2031_0, i_13_352_2117_0, i_13_352_2137_0, i_13_352_2209_0,
    i_13_352_2263_0, i_13_352_2297_0, i_13_352_2407_0, i_13_352_2408_0,
    i_13_352_2432_0, i_13_352_2445_0, i_13_352_2498_0, i_13_352_2501_0,
    i_13_352_2517_0, i_13_352_2725_0, i_13_352_2812_0, i_13_352_2884_0,
    i_13_352_2938_0, i_13_352_3047_0, i_13_352_3076_0, i_13_352_3089_0,
    i_13_352_3115_0, i_13_352_3208_0, i_13_352_3209_0, i_13_352_3424_0,
    i_13_352_3476_0, i_13_352_3505_0, i_13_352_3565_0, i_13_352_3569_0,
    i_13_352_3597_0, i_13_352_3611_0, i_13_352_3614_0, i_13_352_3730_0,
    i_13_352_3739_0, i_13_352_3740_0, i_13_352_3741_0, i_13_352_3747_0,
    i_13_352_4036_0, i_13_352_4063_0, i_13_352_4064_0, i_13_352_4160_0,
    i_13_352_4163_0, i_13_352_4164_0, i_13_352_4202_0, i_13_352_4316_0,
    i_13_352_4327_0, i_13_352_4330_0, i_13_352_4331_0, i_13_352_4340_0,
    i_13_352_4367_0, i_13_352_4369_0, i_13_352_4370_0, i_13_352_4372_0,
    i_13_352_4517_0, i_13_352_4600_0, i_13_352_4604_0, i_13_352_4606_0,
    o_13_352_0_0  );
  input  i_13_352_74_0, i_13_352_77_0, i_13_352_137_0, i_13_352_170_0,
    i_13_352_265_0, i_13_352_266_0, i_13_352_283_0, i_13_352_319_0,
    i_13_352_337_0, i_13_352_492_0, i_13_352_518_0, i_13_352_571_0,
    i_13_352_582_0, i_13_352_662_0, i_13_352_688_0, i_13_352_697_0,
    i_13_352_814_0, i_13_352_886_0, i_13_352_888_0, i_13_352_935_0,
    i_13_352_939_0, i_13_352_1066_0, i_13_352_1112_0, i_13_352_1145_0,
    i_13_352_1148_0, i_13_352_1208_0, i_13_352_1210_0, i_13_352_1217_0,
    i_13_352_1226_0, i_13_352_1253_0, i_13_352_1266_0, i_13_352_1426_0,
    i_13_352_1530_0, i_13_352_1633_0, i_13_352_1660_0, i_13_352_1662_0,
    i_13_352_1730_0, i_13_352_1731_0, i_13_352_1733_0, i_13_352_1734_0,
    i_13_352_1849_0, i_13_352_1886_0, i_13_352_2020_0, i_13_352_2021_0,
    i_13_352_2031_0, i_13_352_2117_0, i_13_352_2137_0, i_13_352_2209_0,
    i_13_352_2263_0, i_13_352_2297_0, i_13_352_2407_0, i_13_352_2408_0,
    i_13_352_2432_0, i_13_352_2445_0, i_13_352_2498_0, i_13_352_2501_0,
    i_13_352_2517_0, i_13_352_2725_0, i_13_352_2812_0, i_13_352_2884_0,
    i_13_352_2938_0, i_13_352_3047_0, i_13_352_3076_0, i_13_352_3089_0,
    i_13_352_3115_0, i_13_352_3208_0, i_13_352_3209_0, i_13_352_3424_0,
    i_13_352_3476_0, i_13_352_3505_0, i_13_352_3565_0, i_13_352_3569_0,
    i_13_352_3597_0, i_13_352_3611_0, i_13_352_3614_0, i_13_352_3730_0,
    i_13_352_3739_0, i_13_352_3740_0, i_13_352_3741_0, i_13_352_3747_0,
    i_13_352_4036_0, i_13_352_4063_0, i_13_352_4064_0, i_13_352_4160_0,
    i_13_352_4163_0, i_13_352_4164_0, i_13_352_4202_0, i_13_352_4316_0,
    i_13_352_4327_0, i_13_352_4330_0, i_13_352_4331_0, i_13_352_4340_0,
    i_13_352_4367_0, i_13_352_4369_0, i_13_352_4370_0, i_13_352_4372_0,
    i_13_352_4517_0, i_13_352_4600_0, i_13_352_4604_0, i_13_352_4606_0;
  output o_13_352_0_0;
  assign o_13_352_0_0 = ~((~i_13_352_4517_0 & (i_13_352_814_0 | (i_13_352_337_0 & ((~i_13_352_697_0 & ~i_13_352_1145_0 & ~i_13_352_1208_0) | (~i_13_352_1660_0 & ~i_13_352_3424_0 & ~i_13_352_3565_0))))) | (~i_13_352_1208_0 & ((~i_13_352_2020_0 & ~i_13_352_2432_0 & ~i_13_352_3569_0) | (~i_13_352_1253_0 & i_13_352_3424_0 & ~i_13_352_4164_0 & ~i_13_352_4330_0 & ~i_13_352_4370_0))) | (~i_13_352_697_0 & i_13_352_2407_0) | (~i_13_352_77_0 & ~i_13_352_935_0 & ~i_13_352_2297_0 & ~i_13_352_3565_0 & ~i_13_352_3740_0 & ~i_13_352_4164_0) | (i_13_352_283_0 & ~i_13_352_688_0 & i_13_352_3747_0) | (~i_13_352_137_0 & ~i_13_352_1660_0 & i_13_352_4064_0) | (~i_13_352_1210_0 & ~i_13_352_1253_0 & ~i_13_352_4160_0) | (~i_13_352_1145_0 & ~i_13_352_1426_0 & ~i_13_352_3209_0 & ~i_13_352_4331_0 & ~i_13_352_4372_0));
endmodule



// Benchmark "kernel_13_353" written by ABC on Sun Jul 19 10:50:19 2020

module kernel_13_353 ( 
    i_13_353_52_0, i_13_353_111_0, i_13_353_124_0, i_13_353_140_0,
    i_13_353_169_0, i_13_353_170_0, i_13_353_269_0, i_13_353_273_0,
    i_13_353_283_0, i_13_353_287_0, i_13_353_371_0, i_13_353_373_0,
    i_13_353_417_0, i_13_353_463_0, i_13_353_509_0, i_13_353_692_0,
    i_13_353_817_0, i_13_353_818_0, i_13_353_849_0, i_13_353_851_0,
    i_13_353_853_0, i_13_353_886_0, i_13_353_887_0, i_13_353_916_0,
    i_13_353_939_0, i_13_353_943_0, i_13_353_985_0, i_13_353_1053_0,
    i_13_353_1067_0, i_13_353_1110_0, i_13_353_1121_0, i_13_353_1122_0,
    i_13_353_1328_0, i_13_353_1329_0, i_13_353_1492_0, i_13_353_1573_0,
    i_13_353_1623_0, i_13_353_1808_0, i_13_353_1830_0, i_13_353_1840_0,
    i_13_353_1852_0, i_13_353_1853_0, i_13_353_1857_0, i_13_353_1924_0,
    i_13_353_2006_0, i_13_353_2051_0, i_13_353_2123_0, i_13_353_2136_0,
    i_13_353_2140_0, i_13_353_2141_0, i_13_353_2173_0, i_13_353_2237_0,
    i_13_353_2407_0, i_13_353_2408_0, i_13_353_2410_0, i_13_353_2411_0,
    i_13_353_2460_0, i_13_353_2552_0, i_13_353_2696_0, i_13_353_2823_0,
    i_13_353_2848_0, i_13_353_2875_0, i_13_353_2941_0, i_13_353_2942_0,
    i_13_353_3011_0, i_13_353_3031_0, i_13_353_3037_0, i_13_353_3050_0,
    i_13_353_3108_0, i_13_353_3346_0, i_13_353_3400_0, i_13_353_3424_0,
    i_13_353_3453_0, i_13_353_3478_0, i_13_353_3479_0, i_13_353_3505_0,
    i_13_353_3525_0, i_13_353_3526_0, i_13_353_3567_0, i_13_353_3741_0,
    i_13_353_3742_0, i_13_353_3765_0, i_13_353_3821_0, i_13_353_3867_0,
    i_13_353_3911_0, i_13_353_3928_0, i_13_353_3984_0, i_13_353_4022_0,
    i_13_353_4063_0, i_13_353_4064_0, i_13_353_4066_0, i_13_353_4067_0,
    i_13_353_4164_0, i_13_353_4209_0, i_13_353_4309_0, i_13_353_4318_0,
    i_13_353_4319_0, i_13_353_4434_0, i_13_353_4441_0, i_13_353_4451_0,
    o_13_353_0_0  );
  input  i_13_353_52_0, i_13_353_111_0, i_13_353_124_0, i_13_353_140_0,
    i_13_353_169_0, i_13_353_170_0, i_13_353_269_0, i_13_353_273_0,
    i_13_353_283_0, i_13_353_287_0, i_13_353_371_0, i_13_353_373_0,
    i_13_353_417_0, i_13_353_463_0, i_13_353_509_0, i_13_353_692_0,
    i_13_353_817_0, i_13_353_818_0, i_13_353_849_0, i_13_353_851_0,
    i_13_353_853_0, i_13_353_886_0, i_13_353_887_0, i_13_353_916_0,
    i_13_353_939_0, i_13_353_943_0, i_13_353_985_0, i_13_353_1053_0,
    i_13_353_1067_0, i_13_353_1110_0, i_13_353_1121_0, i_13_353_1122_0,
    i_13_353_1328_0, i_13_353_1329_0, i_13_353_1492_0, i_13_353_1573_0,
    i_13_353_1623_0, i_13_353_1808_0, i_13_353_1830_0, i_13_353_1840_0,
    i_13_353_1852_0, i_13_353_1853_0, i_13_353_1857_0, i_13_353_1924_0,
    i_13_353_2006_0, i_13_353_2051_0, i_13_353_2123_0, i_13_353_2136_0,
    i_13_353_2140_0, i_13_353_2141_0, i_13_353_2173_0, i_13_353_2237_0,
    i_13_353_2407_0, i_13_353_2408_0, i_13_353_2410_0, i_13_353_2411_0,
    i_13_353_2460_0, i_13_353_2552_0, i_13_353_2696_0, i_13_353_2823_0,
    i_13_353_2848_0, i_13_353_2875_0, i_13_353_2941_0, i_13_353_2942_0,
    i_13_353_3011_0, i_13_353_3031_0, i_13_353_3037_0, i_13_353_3050_0,
    i_13_353_3108_0, i_13_353_3346_0, i_13_353_3400_0, i_13_353_3424_0,
    i_13_353_3453_0, i_13_353_3478_0, i_13_353_3479_0, i_13_353_3505_0,
    i_13_353_3525_0, i_13_353_3526_0, i_13_353_3567_0, i_13_353_3741_0,
    i_13_353_3742_0, i_13_353_3765_0, i_13_353_3821_0, i_13_353_3867_0,
    i_13_353_3911_0, i_13_353_3928_0, i_13_353_3984_0, i_13_353_4022_0,
    i_13_353_4063_0, i_13_353_4064_0, i_13_353_4066_0, i_13_353_4067_0,
    i_13_353_4164_0, i_13_353_4209_0, i_13_353_4309_0, i_13_353_4318_0,
    i_13_353_4319_0, i_13_353_4434_0, i_13_353_4441_0, i_13_353_4451_0;
  output o_13_353_0_0;
  assign o_13_353_0_0 = ~((~i_13_353_4066_0 & (~i_13_353_287_0 | ~i_13_353_2141_0)) | i_13_353_3741_0 | (~i_13_353_817_0 & ~i_13_353_2411_0 & ~i_13_353_4064_0) | (i_13_353_1121_0 & ~i_13_353_4067_0));
endmodule



// Benchmark "kernel_13_354" written by ABC on Sun Jul 19 10:50:19 2020

module kernel_13_354 ( 
    i_13_354_73_0, i_13_354_74_0, i_13_354_123_0, i_13_354_186_0,
    i_13_354_235_0, i_13_354_280_0, i_13_354_284_0, i_13_354_442_0,
    i_13_354_523_0, i_13_354_532_0, i_13_354_533_0, i_13_354_640_0,
    i_13_354_668_0, i_13_354_676_0, i_13_354_677_0, i_13_354_680_0,
    i_13_354_717_0, i_13_354_832_0, i_13_354_839_0, i_13_354_958_0,
    i_13_354_982_0, i_13_354_1084_0, i_13_354_1099_0, i_13_354_1145_0,
    i_13_354_1256_0, i_13_354_1270_0, i_13_354_1271_0, i_13_354_1302_0,
    i_13_354_1400_0, i_13_354_1464_0, i_13_354_1504_0, i_13_354_1505_0,
    i_13_354_1594_0, i_13_354_1658_0, i_13_354_1720_0, i_13_354_1723_0,
    i_13_354_1744_0, i_13_354_1775_0, i_13_354_1792_0, i_13_354_1796_0,
    i_13_354_1881_0, i_13_354_1915_0, i_13_354_1989_0, i_13_354_2017_0,
    i_13_354_2026_0, i_13_354_2116_0, i_13_354_2223_0, i_13_354_2446_0,
    i_13_354_2511_0, i_13_354_2512_0, i_13_354_2539_0, i_13_354_2575_0,
    i_13_354_2576_0, i_13_354_2611_0, i_13_354_2750_0, i_13_354_2844_0,
    i_13_354_2845_0, i_13_354_2854_0, i_13_354_2921_0, i_13_354_2922_0,
    i_13_354_2935_0, i_13_354_3001_0, i_13_354_3135_0, i_13_354_3259_0,
    i_13_354_3260_0, i_13_354_3287_0, i_13_354_3289_0, i_13_354_3321_0,
    i_13_354_3350_0, i_13_354_3371_0, i_13_354_3396_0, i_13_354_3449_0,
    i_13_354_3452_0, i_13_354_3477_0, i_13_354_3578_0, i_13_354_3593_0,
    i_13_354_3647_0, i_13_354_3784_0, i_13_354_3865_0, i_13_354_3889_0,
    i_13_354_3907_0, i_13_354_3924_0, i_13_354_3925_0, i_13_354_3926_0,
    i_13_354_3984_0, i_13_354_3988_0, i_13_354_3989_0, i_13_354_4078_0,
    i_13_354_4079_0, i_13_354_4099_0, i_13_354_4106_0, i_13_354_4163_0,
    i_13_354_4186_0, i_13_354_4187_0, i_13_354_4331_0, i_13_354_4340_0,
    i_13_354_4430_0, i_13_354_4452_0, i_13_354_4543_0, i_13_354_4592_0,
    o_13_354_0_0  );
  input  i_13_354_73_0, i_13_354_74_0, i_13_354_123_0, i_13_354_186_0,
    i_13_354_235_0, i_13_354_280_0, i_13_354_284_0, i_13_354_442_0,
    i_13_354_523_0, i_13_354_532_0, i_13_354_533_0, i_13_354_640_0,
    i_13_354_668_0, i_13_354_676_0, i_13_354_677_0, i_13_354_680_0,
    i_13_354_717_0, i_13_354_832_0, i_13_354_839_0, i_13_354_958_0,
    i_13_354_982_0, i_13_354_1084_0, i_13_354_1099_0, i_13_354_1145_0,
    i_13_354_1256_0, i_13_354_1270_0, i_13_354_1271_0, i_13_354_1302_0,
    i_13_354_1400_0, i_13_354_1464_0, i_13_354_1504_0, i_13_354_1505_0,
    i_13_354_1594_0, i_13_354_1658_0, i_13_354_1720_0, i_13_354_1723_0,
    i_13_354_1744_0, i_13_354_1775_0, i_13_354_1792_0, i_13_354_1796_0,
    i_13_354_1881_0, i_13_354_1915_0, i_13_354_1989_0, i_13_354_2017_0,
    i_13_354_2026_0, i_13_354_2116_0, i_13_354_2223_0, i_13_354_2446_0,
    i_13_354_2511_0, i_13_354_2512_0, i_13_354_2539_0, i_13_354_2575_0,
    i_13_354_2576_0, i_13_354_2611_0, i_13_354_2750_0, i_13_354_2844_0,
    i_13_354_2845_0, i_13_354_2854_0, i_13_354_2921_0, i_13_354_2922_0,
    i_13_354_2935_0, i_13_354_3001_0, i_13_354_3135_0, i_13_354_3259_0,
    i_13_354_3260_0, i_13_354_3287_0, i_13_354_3289_0, i_13_354_3321_0,
    i_13_354_3350_0, i_13_354_3371_0, i_13_354_3396_0, i_13_354_3449_0,
    i_13_354_3452_0, i_13_354_3477_0, i_13_354_3578_0, i_13_354_3593_0,
    i_13_354_3647_0, i_13_354_3784_0, i_13_354_3865_0, i_13_354_3889_0,
    i_13_354_3907_0, i_13_354_3924_0, i_13_354_3925_0, i_13_354_3926_0,
    i_13_354_3984_0, i_13_354_3988_0, i_13_354_3989_0, i_13_354_4078_0,
    i_13_354_4079_0, i_13_354_4099_0, i_13_354_4106_0, i_13_354_4163_0,
    i_13_354_4186_0, i_13_354_4187_0, i_13_354_4331_0, i_13_354_4340_0,
    i_13_354_4430_0, i_13_354_4452_0, i_13_354_4543_0, i_13_354_4592_0;
  output o_13_354_0_0;
  assign o_13_354_0_0 = ~((~i_13_354_3988_0 & ~i_13_354_4078_0) | (~i_13_354_280_0 & ~i_13_354_533_0 & ~i_13_354_1504_0) | (i_13_354_523_0 & ~i_13_354_676_0 & i_13_354_2026_0 & ~i_13_354_2844_0 & ~i_13_354_3989_0 & ~i_13_354_4187_0));
endmodule



// Benchmark "kernel_13_355" written by ABC on Sun Jul 19 10:50:20 2020

module kernel_13_355 ( 
    i_13_355_45_0, i_13_355_172_0, i_13_355_175_0, i_13_355_178_0,
    i_13_355_179_0, i_13_355_229_0, i_13_355_280_0, i_13_355_283_0,
    i_13_355_284_0, i_13_355_286_0, i_13_355_287_0, i_13_355_335_0,
    i_13_355_360_0, i_13_355_454_0, i_13_355_562_0, i_13_355_574_0,
    i_13_355_589_0, i_13_355_645_0, i_13_355_687_0, i_13_355_688_0,
    i_13_355_691_0, i_13_355_742_0, i_13_355_760_0, i_13_355_823_0,
    i_13_355_832_0, i_13_355_867_0, i_13_355_871_0, i_13_355_872_0,
    i_13_355_1078_0, i_13_355_1085_0, i_13_355_1122_0, i_13_355_1228_0,
    i_13_355_1229_0, i_13_355_1469_0, i_13_355_1573_0, i_13_355_1636_0,
    i_13_355_1710_0, i_13_355_1712_0, i_13_355_1716_0, i_13_355_1732_0,
    i_13_355_1747_0, i_13_355_1750_0, i_13_355_1751_0, i_13_355_1855_0,
    i_13_355_1858_0, i_13_355_1859_0, i_13_355_1861_0, i_13_355_1864_0,
    i_13_355_1933_0, i_13_355_2239_0, i_13_355_2341_0, i_13_355_2428_0,
    i_13_355_2624_0, i_13_355_2652_0, i_13_355_2653_0, i_13_355_2654_0,
    i_13_355_2708_0, i_13_355_2722_0, i_13_355_2731_0, i_13_355_2752_0,
    i_13_355_2785_0, i_13_355_2851_0, i_13_355_3092_0, i_13_355_3100_0,
    i_13_355_3113_0, i_13_355_3172_0, i_13_355_3174_0, i_13_355_3235_0,
    i_13_355_3267_0, i_13_355_3268_0, i_13_355_3271_0, i_13_355_3274_0,
    i_13_355_3293_0, i_13_355_3371_0, i_13_355_3400_0, i_13_355_3424_0,
    i_13_355_3426_0, i_13_355_3427_0, i_13_355_3428_0, i_13_355_3646_0,
    i_13_355_3686_0, i_13_355_3783_0, i_13_355_3890_0, i_13_355_3910_0,
    i_13_355_3911_0, i_13_355_3913_0, i_13_355_3914_0, i_13_355_3995_0,
    i_13_355_4017_0, i_13_355_4018_0, i_13_355_4019_0, i_13_355_4021_0,
    i_13_355_4090_0, i_13_355_4097_0, i_13_355_4295_0, i_13_355_4322_0,
    i_13_355_4556_0, i_13_355_4559_0, i_13_355_4561_0, i_13_355_4573_0,
    o_13_355_0_0  );
  input  i_13_355_45_0, i_13_355_172_0, i_13_355_175_0, i_13_355_178_0,
    i_13_355_179_0, i_13_355_229_0, i_13_355_280_0, i_13_355_283_0,
    i_13_355_284_0, i_13_355_286_0, i_13_355_287_0, i_13_355_335_0,
    i_13_355_360_0, i_13_355_454_0, i_13_355_562_0, i_13_355_574_0,
    i_13_355_589_0, i_13_355_645_0, i_13_355_687_0, i_13_355_688_0,
    i_13_355_691_0, i_13_355_742_0, i_13_355_760_0, i_13_355_823_0,
    i_13_355_832_0, i_13_355_867_0, i_13_355_871_0, i_13_355_872_0,
    i_13_355_1078_0, i_13_355_1085_0, i_13_355_1122_0, i_13_355_1228_0,
    i_13_355_1229_0, i_13_355_1469_0, i_13_355_1573_0, i_13_355_1636_0,
    i_13_355_1710_0, i_13_355_1712_0, i_13_355_1716_0, i_13_355_1732_0,
    i_13_355_1747_0, i_13_355_1750_0, i_13_355_1751_0, i_13_355_1855_0,
    i_13_355_1858_0, i_13_355_1859_0, i_13_355_1861_0, i_13_355_1864_0,
    i_13_355_1933_0, i_13_355_2239_0, i_13_355_2341_0, i_13_355_2428_0,
    i_13_355_2624_0, i_13_355_2652_0, i_13_355_2653_0, i_13_355_2654_0,
    i_13_355_2708_0, i_13_355_2722_0, i_13_355_2731_0, i_13_355_2752_0,
    i_13_355_2785_0, i_13_355_2851_0, i_13_355_3092_0, i_13_355_3100_0,
    i_13_355_3113_0, i_13_355_3172_0, i_13_355_3174_0, i_13_355_3235_0,
    i_13_355_3267_0, i_13_355_3268_0, i_13_355_3271_0, i_13_355_3274_0,
    i_13_355_3293_0, i_13_355_3371_0, i_13_355_3400_0, i_13_355_3424_0,
    i_13_355_3426_0, i_13_355_3427_0, i_13_355_3428_0, i_13_355_3646_0,
    i_13_355_3686_0, i_13_355_3783_0, i_13_355_3890_0, i_13_355_3910_0,
    i_13_355_3911_0, i_13_355_3913_0, i_13_355_3914_0, i_13_355_3995_0,
    i_13_355_4017_0, i_13_355_4018_0, i_13_355_4019_0, i_13_355_4021_0,
    i_13_355_4090_0, i_13_355_4097_0, i_13_355_4295_0, i_13_355_4322_0,
    i_13_355_4556_0, i_13_355_4559_0, i_13_355_4561_0, i_13_355_4573_0;
  output o_13_355_0_0;
  assign o_13_355_0_0 = ~((~i_13_355_1861_0 & (~i_13_355_3424_0 | (~i_13_355_1469_0 & ~i_13_355_3293_0 & ~i_13_355_4559_0))) | (~i_13_355_1858_0 & ((~i_13_355_691_0 & ~i_13_355_1750_0) | ~i_13_355_4559_0 | (~i_13_355_1859_0 & ~i_13_355_2851_0))) | (i_13_355_3235_0 & ~i_13_355_3913_0) | (~i_13_355_283_0 & ~i_13_355_1078_0 & ~i_13_355_2653_0 & ~i_13_355_3995_0));
endmodule



// Benchmark "kernel_13_356" written by ABC on Sun Jul 19 10:50:21 2020

module kernel_13_356 ( 
    i_13_356_44_0, i_13_356_79_0, i_13_356_80_0, i_13_356_168_0,
    i_13_356_276_0, i_13_356_537_0, i_13_356_539_0, i_13_356_554_0,
    i_13_356_591_0, i_13_356_608_0, i_13_356_611_0, i_13_356_645_0,
    i_13_356_647_0, i_13_356_672_0, i_13_356_673_0, i_13_356_674_0,
    i_13_356_682_0, i_13_356_683_0, i_13_356_691_0, i_13_356_692_0,
    i_13_356_701_0, i_13_356_718_0, i_13_356_823_0, i_13_356_844_0,
    i_13_356_978_0, i_13_356_1065_0, i_13_356_1104_0, i_13_356_1123_0,
    i_13_356_1124_0, i_13_356_1218_0, i_13_356_1223_0, i_13_356_1283_0,
    i_13_356_1410_0, i_13_356_1423_0, i_13_356_1426_0, i_13_356_1429_0,
    i_13_356_1470_0, i_13_356_1659_0, i_13_356_1660_0, i_13_356_1663_0,
    i_13_356_1689_0, i_13_356_1727_0, i_13_356_1734_0, i_13_356_1736_0,
    i_13_356_1799_0, i_13_356_1803_0, i_13_356_1842_0, i_13_356_1849_0,
    i_13_356_1992_0, i_13_356_2022_0, i_13_356_2024_0, i_13_356_2058_0,
    i_13_356_2104_0, i_13_356_2450_0, i_13_356_2496_0, i_13_356_2570_0,
    i_13_356_2698_0, i_13_356_2715_0, i_13_356_2887_0, i_13_356_2938_0,
    i_13_356_2982_0, i_13_356_3027_0, i_13_356_3067_0, i_13_356_3068_0,
    i_13_356_3088_0, i_13_356_3089_0, i_13_356_3102_0, i_13_356_3104_0,
    i_13_356_3244_0, i_13_356_3289_0, i_13_356_3454_0, i_13_356_3525_0,
    i_13_356_3572_0, i_13_356_3653_0, i_13_356_3682_0, i_13_356_3739_0,
    i_13_356_3742_0, i_13_356_3743_0, i_13_356_3787_0, i_13_356_3797_0,
    i_13_356_3858_0, i_13_356_3930_0, i_13_356_3931_0, i_13_356_3932_0,
    i_13_356_3994_0, i_13_356_3995_0, i_13_356_4063_0, i_13_356_4084_0,
    i_13_356_4189_0, i_13_356_4190_0, i_13_356_4191_0, i_13_356_4193_0,
    i_13_356_4249_0, i_13_356_4368_0, i_13_356_4515_0, i_13_356_4533_0,
    i_13_356_4595_0, i_13_356_4596_0, i_13_356_4597_0, i_13_356_4598_0,
    o_13_356_0_0  );
  input  i_13_356_44_0, i_13_356_79_0, i_13_356_80_0, i_13_356_168_0,
    i_13_356_276_0, i_13_356_537_0, i_13_356_539_0, i_13_356_554_0,
    i_13_356_591_0, i_13_356_608_0, i_13_356_611_0, i_13_356_645_0,
    i_13_356_647_0, i_13_356_672_0, i_13_356_673_0, i_13_356_674_0,
    i_13_356_682_0, i_13_356_683_0, i_13_356_691_0, i_13_356_692_0,
    i_13_356_701_0, i_13_356_718_0, i_13_356_823_0, i_13_356_844_0,
    i_13_356_978_0, i_13_356_1065_0, i_13_356_1104_0, i_13_356_1123_0,
    i_13_356_1124_0, i_13_356_1218_0, i_13_356_1223_0, i_13_356_1283_0,
    i_13_356_1410_0, i_13_356_1423_0, i_13_356_1426_0, i_13_356_1429_0,
    i_13_356_1470_0, i_13_356_1659_0, i_13_356_1660_0, i_13_356_1663_0,
    i_13_356_1689_0, i_13_356_1727_0, i_13_356_1734_0, i_13_356_1736_0,
    i_13_356_1799_0, i_13_356_1803_0, i_13_356_1842_0, i_13_356_1849_0,
    i_13_356_1992_0, i_13_356_2022_0, i_13_356_2024_0, i_13_356_2058_0,
    i_13_356_2104_0, i_13_356_2450_0, i_13_356_2496_0, i_13_356_2570_0,
    i_13_356_2698_0, i_13_356_2715_0, i_13_356_2887_0, i_13_356_2938_0,
    i_13_356_2982_0, i_13_356_3027_0, i_13_356_3067_0, i_13_356_3068_0,
    i_13_356_3088_0, i_13_356_3089_0, i_13_356_3102_0, i_13_356_3104_0,
    i_13_356_3244_0, i_13_356_3289_0, i_13_356_3454_0, i_13_356_3525_0,
    i_13_356_3572_0, i_13_356_3653_0, i_13_356_3682_0, i_13_356_3739_0,
    i_13_356_3742_0, i_13_356_3743_0, i_13_356_3787_0, i_13_356_3797_0,
    i_13_356_3858_0, i_13_356_3930_0, i_13_356_3931_0, i_13_356_3932_0,
    i_13_356_3994_0, i_13_356_3995_0, i_13_356_4063_0, i_13_356_4084_0,
    i_13_356_4189_0, i_13_356_4190_0, i_13_356_4191_0, i_13_356_4193_0,
    i_13_356_4249_0, i_13_356_4368_0, i_13_356_4515_0, i_13_356_4533_0,
    i_13_356_4595_0, i_13_356_4596_0, i_13_356_4597_0, i_13_356_4598_0;
  output o_13_356_0_0;
  assign o_13_356_0_0 = ~((~i_13_356_1124_0 & ((~i_13_356_80_0 & ~i_13_356_1429_0 & ~i_13_356_3931_0) | (~i_13_356_674_0 & ~i_13_356_701_0 & ~i_13_356_3994_0 & ~i_13_356_4191_0))) | (~i_13_356_4193_0 & ((~i_13_356_79_0 & ~i_13_356_1223_0) | (~i_13_356_539_0 & ~i_13_356_1123_0 & ~i_13_356_3244_0))) | (i_13_356_4063_0 & (~i_13_356_823_0 | i_13_356_3787_0 | ~i_13_356_4190_0)));
endmodule



// Benchmark "kernel_13_357" written by ABC on Sun Jul 19 10:50:22 2020

module kernel_13_357 ( 
    i_13_357_27_0, i_13_357_28_0, i_13_357_35_0, i_13_357_37_0,
    i_13_357_54_0, i_13_357_63_0, i_13_357_64_0, i_13_357_80_0,
    i_13_357_135_0, i_13_357_172_0, i_13_357_178_0, i_13_357_306_0,
    i_13_357_307_0, i_13_357_316_0, i_13_357_325_0, i_13_357_379_0,
    i_13_357_383_0, i_13_357_588_0, i_13_357_612_0, i_13_357_639_0,
    i_13_357_642_0, i_13_357_647_0, i_13_357_694_0, i_13_357_772_0,
    i_13_357_944_0, i_13_357_1121_0, i_13_357_1131_0, i_13_357_1198_0,
    i_13_357_1206_0, i_13_357_1227_0, i_13_357_1269_0, i_13_357_1270_0,
    i_13_357_1272_0, i_13_357_1305_0, i_13_357_1309_0, i_13_357_1342_0,
    i_13_357_1351_0, i_13_357_1390_0, i_13_357_1396_0, i_13_357_1489_0,
    i_13_357_1504_0, i_13_357_1593_0, i_13_357_1594_0, i_13_357_1638_0,
    i_13_357_1639_0, i_13_357_1792_0, i_13_357_1828_0, i_13_357_1881_0,
    i_13_357_1882_0, i_13_357_1909_0, i_13_357_1918_0, i_13_357_1926_0,
    i_13_357_1927_0, i_13_357_1931_0, i_13_357_2008_0, i_13_357_2011_0,
    i_13_357_2126_0, i_13_357_2537_0, i_13_357_2596_0, i_13_357_2673_0,
    i_13_357_2674_0, i_13_357_2719_0, i_13_357_2848_0, i_13_357_2849_0,
    i_13_357_2875_0, i_13_357_2880_0, i_13_357_2881_0, i_13_357_2934_0,
    i_13_357_3040_0, i_13_357_3060_0, i_13_357_3061_0, i_13_357_3204_0,
    i_13_357_3208_0, i_13_357_3218_0, i_13_357_3241_0, i_13_357_3387_0,
    i_13_357_3397_0, i_13_357_3505_0, i_13_357_3636_0, i_13_357_3738_0,
    i_13_357_3853_0, i_13_357_3916_0, i_13_357_3925_0, i_13_357_3932_0,
    i_13_357_3934_0, i_13_357_3973_0, i_13_357_4033_0, i_13_357_4064_0,
    i_13_357_4091_0, i_13_357_4185_0, i_13_357_4213_0, i_13_357_4215_0,
    i_13_357_4260_0, i_13_357_4294_0, i_13_357_4302_0, i_13_357_4308_0,
    i_13_357_4315_0, i_13_357_4393_0, i_13_357_4396_0, i_13_357_4593_0,
    o_13_357_0_0  );
  input  i_13_357_27_0, i_13_357_28_0, i_13_357_35_0, i_13_357_37_0,
    i_13_357_54_0, i_13_357_63_0, i_13_357_64_0, i_13_357_80_0,
    i_13_357_135_0, i_13_357_172_0, i_13_357_178_0, i_13_357_306_0,
    i_13_357_307_0, i_13_357_316_0, i_13_357_325_0, i_13_357_379_0,
    i_13_357_383_0, i_13_357_588_0, i_13_357_612_0, i_13_357_639_0,
    i_13_357_642_0, i_13_357_647_0, i_13_357_694_0, i_13_357_772_0,
    i_13_357_944_0, i_13_357_1121_0, i_13_357_1131_0, i_13_357_1198_0,
    i_13_357_1206_0, i_13_357_1227_0, i_13_357_1269_0, i_13_357_1270_0,
    i_13_357_1272_0, i_13_357_1305_0, i_13_357_1309_0, i_13_357_1342_0,
    i_13_357_1351_0, i_13_357_1390_0, i_13_357_1396_0, i_13_357_1489_0,
    i_13_357_1504_0, i_13_357_1593_0, i_13_357_1594_0, i_13_357_1638_0,
    i_13_357_1639_0, i_13_357_1792_0, i_13_357_1828_0, i_13_357_1881_0,
    i_13_357_1882_0, i_13_357_1909_0, i_13_357_1918_0, i_13_357_1926_0,
    i_13_357_1927_0, i_13_357_1931_0, i_13_357_2008_0, i_13_357_2011_0,
    i_13_357_2126_0, i_13_357_2537_0, i_13_357_2596_0, i_13_357_2673_0,
    i_13_357_2674_0, i_13_357_2719_0, i_13_357_2848_0, i_13_357_2849_0,
    i_13_357_2875_0, i_13_357_2880_0, i_13_357_2881_0, i_13_357_2934_0,
    i_13_357_3040_0, i_13_357_3060_0, i_13_357_3061_0, i_13_357_3204_0,
    i_13_357_3208_0, i_13_357_3218_0, i_13_357_3241_0, i_13_357_3387_0,
    i_13_357_3397_0, i_13_357_3505_0, i_13_357_3636_0, i_13_357_3738_0,
    i_13_357_3853_0, i_13_357_3916_0, i_13_357_3925_0, i_13_357_3932_0,
    i_13_357_3934_0, i_13_357_3973_0, i_13_357_4033_0, i_13_357_4064_0,
    i_13_357_4091_0, i_13_357_4185_0, i_13_357_4213_0, i_13_357_4215_0,
    i_13_357_4260_0, i_13_357_4294_0, i_13_357_4302_0, i_13_357_4308_0,
    i_13_357_4315_0, i_13_357_4393_0, i_13_357_4396_0, i_13_357_4593_0;
  output o_13_357_0_0;
  assign o_13_357_0_0 = ~((~i_13_357_54_0 & ((~i_13_357_63_0 & ~i_13_357_612_0 & ~i_13_357_1121_0 & ~i_13_357_1792_0 & ~i_13_357_2881_0) | (~i_13_357_316_0 & ~i_13_357_1593_0 & ~i_13_357_4393_0 & ~i_13_357_4396_0))) | (~i_13_357_2673_0 & ((~i_13_357_694_0 & ~i_13_357_2881_0) | (i_13_357_1828_0 & i_13_357_4396_0))) | (~i_13_357_306_0 & ~i_13_357_379_0 & ~i_13_357_2934_0 & ~i_13_357_3060_0));
endmodule



// Benchmark "kernel_13_358" written by ABC on Sun Jul 19 10:50:22 2020

module kernel_13_358 ( 
    i_13_358_67_0, i_13_358_105_0, i_13_358_106_0, i_13_358_165_0,
    i_13_358_241_0, i_13_358_258_0, i_13_358_339_0, i_13_358_527_0,
    i_13_358_662_0, i_13_358_697_0, i_13_358_771_0, i_13_358_793_0,
    i_13_358_817_0, i_13_358_831_0, i_13_358_832_0, i_13_358_851_0,
    i_13_358_855_0, i_13_358_856_0, i_13_358_897_0, i_13_358_1068_0,
    i_13_358_1069_0, i_13_358_1076_0, i_13_358_1099_0, i_13_358_1279_0,
    i_13_358_1309_0, i_13_358_1464_0, i_13_358_1470_0, i_13_358_1485_0,
    i_13_358_1497_0, i_13_358_1572_0, i_13_358_1573_0, i_13_358_1597_0,
    i_13_358_1642_0, i_13_358_1679_0, i_13_358_1735_0, i_13_358_1788_0,
    i_13_358_1852_0, i_13_358_1914_0, i_13_358_1935_0, i_13_358_1996_0,
    i_13_358_2120_0, i_13_358_2122_0, i_13_358_2123_0, i_13_358_2139_0,
    i_13_358_2140_0, i_13_358_2184_0, i_13_358_2209_0, i_13_358_2280_0,
    i_13_358_2409_0, i_13_358_2453_0, i_13_358_2460_0, i_13_358_2461_0,
    i_13_358_2464_0, i_13_358_2536_0, i_13_358_2640_0, i_13_358_2722_0,
    i_13_358_2751_0, i_13_358_2757_0, i_13_358_2760_0, i_13_358_2940_0,
    i_13_358_2941_0, i_13_358_2942_0, i_13_358_2982_0, i_13_358_3014_0,
    i_13_358_3030_0, i_13_358_3031_0, i_13_358_3040_0, i_13_358_3106_0,
    i_13_358_3148_0, i_13_358_3244_0, i_13_358_3291_0, i_13_358_3292_0,
    i_13_358_3322_0, i_13_358_3346_0, i_13_358_3399_0, i_13_358_3400_0,
    i_13_358_3402_0, i_13_358_3417_0, i_13_358_3418_0, i_13_358_3423_0,
    i_13_358_3525_0, i_13_358_3526_0, i_13_358_3732_0, i_13_358_3785_0,
    i_13_358_3866_0, i_13_358_3909_0, i_13_358_3911_0, i_13_358_4047_0,
    i_13_358_4056_0, i_13_358_4066_0, i_13_358_4120_0, i_13_358_4216_0,
    i_13_358_4317_0, i_13_358_4318_0, i_13_358_4357_0, i_13_358_4366_0,
    i_13_358_4391_0, i_13_358_4524_0, i_13_358_4559_0, i_13_358_4562_0,
    o_13_358_0_0  );
  input  i_13_358_67_0, i_13_358_105_0, i_13_358_106_0, i_13_358_165_0,
    i_13_358_241_0, i_13_358_258_0, i_13_358_339_0, i_13_358_527_0,
    i_13_358_662_0, i_13_358_697_0, i_13_358_771_0, i_13_358_793_0,
    i_13_358_817_0, i_13_358_831_0, i_13_358_832_0, i_13_358_851_0,
    i_13_358_855_0, i_13_358_856_0, i_13_358_897_0, i_13_358_1068_0,
    i_13_358_1069_0, i_13_358_1076_0, i_13_358_1099_0, i_13_358_1279_0,
    i_13_358_1309_0, i_13_358_1464_0, i_13_358_1470_0, i_13_358_1485_0,
    i_13_358_1497_0, i_13_358_1572_0, i_13_358_1573_0, i_13_358_1597_0,
    i_13_358_1642_0, i_13_358_1679_0, i_13_358_1735_0, i_13_358_1788_0,
    i_13_358_1852_0, i_13_358_1914_0, i_13_358_1935_0, i_13_358_1996_0,
    i_13_358_2120_0, i_13_358_2122_0, i_13_358_2123_0, i_13_358_2139_0,
    i_13_358_2140_0, i_13_358_2184_0, i_13_358_2209_0, i_13_358_2280_0,
    i_13_358_2409_0, i_13_358_2453_0, i_13_358_2460_0, i_13_358_2461_0,
    i_13_358_2464_0, i_13_358_2536_0, i_13_358_2640_0, i_13_358_2722_0,
    i_13_358_2751_0, i_13_358_2757_0, i_13_358_2760_0, i_13_358_2940_0,
    i_13_358_2941_0, i_13_358_2942_0, i_13_358_2982_0, i_13_358_3014_0,
    i_13_358_3030_0, i_13_358_3031_0, i_13_358_3040_0, i_13_358_3106_0,
    i_13_358_3148_0, i_13_358_3244_0, i_13_358_3291_0, i_13_358_3292_0,
    i_13_358_3322_0, i_13_358_3346_0, i_13_358_3399_0, i_13_358_3400_0,
    i_13_358_3402_0, i_13_358_3417_0, i_13_358_3418_0, i_13_358_3423_0,
    i_13_358_3525_0, i_13_358_3526_0, i_13_358_3732_0, i_13_358_3785_0,
    i_13_358_3866_0, i_13_358_3909_0, i_13_358_3911_0, i_13_358_4047_0,
    i_13_358_4056_0, i_13_358_4066_0, i_13_358_4120_0, i_13_358_4216_0,
    i_13_358_4317_0, i_13_358_4318_0, i_13_358_4357_0, i_13_358_4366_0,
    i_13_358_4391_0, i_13_358_4524_0, i_13_358_4559_0, i_13_358_4562_0;
  output o_13_358_0_0;
  assign o_13_358_0_0 = ~(i_13_358_1076_0 | (i_13_358_1642_0 & i_13_358_3785_0) | (~i_13_358_1069_0 & ~i_13_358_2941_0 & i_13_358_4216_0) | (~i_13_358_1068_0 & ~i_13_358_1573_0 & ~i_13_358_3291_0 & ~i_13_358_4317_0));
endmodule



// Benchmark "kernel_13_359" written by ABC on Sun Jul 19 10:50:23 2020

module kernel_13_359 ( 
    i_13_359_40_0, i_13_359_48_0, i_13_359_64_0, i_13_359_72_0,
    i_13_359_139_0, i_13_359_163_0, i_13_359_174_0, i_13_359_237_0,
    i_13_359_241_0, i_13_359_273_0, i_13_359_274_0, i_13_359_336_0,
    i_13_359_378_0, i_13_359_379_0, i_13_359_450_0, i_13_359_453_0,
    i_13_359_513_0, i_13_359_558_0, i_13_359_559_0, i_13_359_561_0,
    i_13_359_586_0, i_13_359_817_0, i_13_359_840_0, i_13_359_849_0,
    i_13_359_850_0, i_13_359_889_0, i_13_359_927_0, i_13_359_928_0,
    i_13_359_1078_0, i_13_359_1080_0, i_13_359_1081_0, i_13_359_1200_0,
    i_13_359_1261_0, i_13_359_1327_0, i_13_359_1359_0, i_13_359_1371_0,
    i_13_359_1396_0, i_13_359_1494_0, i_13_359_1620_0, i_13_359_1623_0,
    i_13_359_1657_0, i_13_359_1731_0, i_13_359_1732_0, i_13_359_1750_0,
    i_13_359_1785_0, i_13_359_1809_0, i_13_359_1810_0, i_13_359_1917_0,
    i_13_359_1935_0, i_13_359_1936_0, i_13_359_2055_0, i_13_359_2091_0,
    i_13_359_2229_0, i_13_359_2388_0, i_13_359_2430_0, i_13_359_2506_0,
    i_13_359_2512_0, i_13_359_2560_0, i_13_359_2565_0, i_13_359_2650_0,
    i_13_359_2709_0, i_13_359_2938_0, i_13_359_2955_0, i_13_359_3016_0,
    i_13_359_3043_0, i_13_359_3060_0, i_13_359_3096_0, i_13_359_3097_0,
    i_13_359_3141_0, i_13_359_3150_0, i_13_359_3162_0, i_13_359_3204_0,
    i_13_359_3205_0, i_13_359_3213_0, i_13_359_3216_0, i_13_359_3217_0,
    i_13_359_3231_0, i_13_359_3234_0, i_13_359_3312_0, i_13_359_3519_0,
    i_13_359_3549_0, i_13_359_3600_0, i_13_359_3681_0, i_13_359_3684_0,
    i_13_359_3720_0, i_13_359_3853_0, i_13_359_3873_0, i_13_359_3900_0,
    i_13_359_4087_0, i_13_359_4159_0, i_13_359_4162_0, i_13_359_4170_0,
    i_13_359_4207_0, i_13_359_4339_0, i_13_359_4359_0, i_13_359_4410_0,
    i_13_359_4530_0, i_13_359_4554_0, i_13_359_4594_0, i_13_359_4603_0,
    o_13_359_0_0  );
  input  i_13_359_40_0, i_13_359_48_0, i_13_359_64_0, i_13_359_72_0,
    i_13_359_139_0, i_13_359_163_0, i_13_359_174_0, i_13_359_237_0,
    i_13_359_241_0, i_13_359_273_0, i_13_359_274_0, i_13_359_336_0,
    i_13_359_378_0, i_13_359_379_0, i_13_359_450_0, i_13_359_453_0,
    i_13_359_513_0, i_13_359_558_0, i_13_359_559_0, i_13_359_561_0,
    i_13_359_586_0, i_13_359_817_0, i_13_359_840_0, i_13_359_849_0,
    i_13_359_850_0, i_13_359_889_0, i_13_359_927_0, i_13_359_928_0,
    i_13_359_1078_0, i_13_359_1080_0, i_13_359_1081_0, i_13_359_1200_0,
    i_13_359_1261_0, i_13_359_1327_0, i_13_359_1359_0, i_13_359_1371_0,
    i_13_359_1396_0, i_13_359_1494_0, i_13_359_1620_0, i_13_359_1623_0,
    i_13_359_1657_0, i_13_359_1731_0, i_13_359_1732_0, i_13_359_1750_0,
    i_13_359_1785_0, i_13_359_1809_0, i_13_359_1810_0, i_13_359_1917_0,
    i_13_359_1935_0, i_13_359_1936_0, i_13_359_2055_0, i_13_359_2091_0,
    i_13_359_2229_0, i_13_359_2388_0, i_13_359_2430_0, i_13_359_2506_0,
    i_13_359_2512_0, i_13_359_2560_0, i_13_359_2565_0, i_13_359_2650_0,
    i_13_359_2709_0, i_13_359_2938_0, i_13_359_2955_0, i_13_359_3016_0,
    i_13_359_3043_0, i_13_359_3060_0, i_13_359_3096_0, i_13_359_3097_0,
    i_13_359_3141_0, i_13_359_3150_0, i_13_359_3162_0, i_13_359_3204_0,
    i_13_359_3205_0, i_13_359_3213_0, i_13_359_3216_0, i_13_359_3217_0,
    i_13_359_3231_0, i_13_359_3234_0, i_13_359_3312_0, i_13_359_3519_0,
    i_13_359_3549_0, i_13_359_3600_0, i_13_359_3681_0, i_13_359_3684_0,
    i_13_359_3720_0, i_13_359_3853_0, i_13_359_3873_0, i_13_359_3900_0,
    i_13_359_4087_0, i_13_359_4159_0, i_13_359_4162_0, i_13_359_4170_0,
    i_13_359_4207_0, i_13_359_4339_0, i_13_359_4359_0, i_13_359_4410_0,
    i_13_359_4530_0, i_13_359_4554_0, i_13_359_4594_0, i_13_359_4603_0;
  output o_13_359_0_0;
  assign o_13_359_0_0 = ~(~i_13_359_2430_0 | (~i_13_359_1080_0 & ~i_13_359_3681_0) | (~i_13_359_558_0 & ~i_13_359_3097_0));
endmodule



// Benchmark "kernel_13_360" written by ABC on Sun Jul 19 10:50:24 2020

module kernel_13_360 ( 
    i_13_360_66_0, i_13_360_108_0, i_13_360_121_0, i_13_360_124_0,
    i_13_360_125_0, i_13_360_140_0, i_13_360_229_0, i_13_360_230_0,
    i_13_360_232_0, i_13_360_268_0, i_13_360_282_0, i_13_360_341_0,
    i_13_360_353_0, i_13_360_381_0, i_13_360_387_0, i_13_360_418_0,
    i_13_360_449_0, i_13_360_517_0, i_13_360_532_0, i_13_360_535_0,
    i_13_360_538_0, i_13_360_539_0, i_13_360_575_0, i_13_360_637_0,
    i_13_360_729_0, i_13_360_734_0, i_13_360_792_0, i_13_360_855_0,
    i_13_360_949_0, i_13_360_985_0, i_13_360_1049_0, i_13_360_1215_0,
    i_13_360_1301_0, i_13_360_1318_0, i_13_360_1367_0, i_13_360_1376_0,
    i_13_360_1394_0, i_13_360_1448_0, i_13_360_1465_0, i_13_360_1485_0,
    i_13_360_1512_0, i_13_360_1723_0, i_13_360_1724_0, i_13_360_1783_0,
    i_13_360_1786_0, i_13_360_1787_0, i_13_360_1789_0, i_13_360_1790_0,
    i_13_360_1827_0, i_13_360_1840_0, i_13_360_1841_0, i_13_360_1843_0,
    i_13_360_1844_0, i_13_360_2128_0, i_13_360_2169_0, i_13_360_2224_0,
    i_13_360_2240_0, i_13_360_2429_0, i_13_360_2430_0, i_13_360_2435_0,
    i_13_360_2849_0, i_13_360_2861_0, i_13_360_2873_0, i_13_360_3023_0,
    i_13_360_3038_0, i_13_360_3047_0, i_13_360_3159_0, i_13_360_3166_0,
    i_13_360_3167_0, i_13_360_3220_0, i_13_360_3236_0, i_13_360_3266_0,
    i_13_360_3410_0, i_13_360_3420_0, i_13_360_3425_0, i_13_360_3428_0,
    i_13_360_3431_0, i_13_360_3487_0, i_13_360_3541_0, i_13_360_3616_0,
    i_13_360_3725_0, i_13_360_3794_0, i_13_360_3839_0, i_13_360_3878_0,
    i_13_360_3906_0, i_13_360_3978_0, i_13_360_3985_0, i_13_360_4005_0,
    i_13_360_4009_0, i_13_360_4011_0, i_13_360_4012_0, i_13_360_4013_0,
    i_13_360_4185_0, i_13_360_4237_0, i_13_360_4238_0, i_13_360_4328_0,
    i_13_360_4370_0, i_13_360_4418_0, i_13_360_4498_0, i_13_360_4536_0,
    o_13_360_0_0  );
  input  i_13_360_66_0, i_13_360_108_0, i_13_360_121_0, i_13_360_124_0,
    i_13_360_125_0, i_13_360_140_0, i_13_360_229_0, i_13_360_230_0,
    i_13_360_232_0, i_13_360_268_0, i_13_360_282_0, i_13_360_341_0,
    i_13_360_353_0, i_13_360_381_0, i_13_360_387_0, i_13_360_418_0,
    i_13_360_449_0, i_13_360_517_0, i_13_360_532_0, i_13_360_535_0,
    i_13_360_538_0, i_13_360_539_0, i_13_360_575_0, i_13_360_637_0,
    i_13_360_729_0, i_13_360_734_0, i_13_360_792_0, i_13_360_855_0,
    i_13_360_949_0, i_13_360_985_0, i_13_360_1049_0, i_13_360_1215_0,
    i_13_360_1301_0, i_13_360_1318_0, i_13_360_1367_0, i_13_360_1376_0,
    i_13_360_1394_0, i_13_360_1448_0, i_13_360_1465_0, i_13_360_1485_0,
    i_13_360_1512_0, i_13_360_1723_0, i_13_360_1724_0, i_13_360_1783_0,
    i_13_360_1786_0, i_13_360_1787_0, i_13_360_1789_0, i_13_360_1790_0,
    i_13_360_1827_0, i_13_360_1840_0, i_13_360_1841_0, i_13_360_1843_0,
    i_13_360_1844_0, i_13_360_2128_0, i_13_360_2169_0, i_13_360_2224_0,
    i_13_360_2240_0, i_13_360_2429_0, i_13_360_2430_0, i_13_360_2435_0,
    i_13_360_2849_0, i_13_360_2861_0, i_13_360_2873_0, i_13_360_3023_0,
    i_13_360_3038_0, i_13_360_3047_0, i_13_360_3159_0, i_13_360_3166_0,
    i_13_360_3167_0, i_13_360_3220_0, i_13_360_3236_0, i_13_360_3266_0,
    i_13_360_3410_0, i_13_360_3420_0, i_13_360_3425_0, i_13_360_3428_0,
    i_13_360_3431_0, i_13_360_3487_0, i_13_360_3541_0, i_13_360_3616_0,
    i_13_360_3725_0, i_13_360_3794_0, i_13_360_3839_0, i_13_360_3878_0,
    i_13_360_3906_0, i_13_360_3978_0, i_13_360_3985_0, i_13_360_4005_0,
    i_13_360_4009_0, i_13_360_4011_0, i_13_360_4012_0, i_13_360_4013_0,
    i_13_360_4185_0, i_13_360_4237_0, i_13_360_4238_0, i_13_360_4328_0,
    i_13_360_4370_0, i_13_360_4418_0, i_13_360_4498_0, i_13_360_4536_0;
  output o_13_360_0_0;
  assign o_13_360_0_0 = ~((~i_13_360_341_0 & ~i_13_360_2429_0) | (~i_13_360_2849_0 & ~i_13_360_4009_0 & ~i_13_360_4012_0) | (~i_13_360_535_0 & ~i_13_360_539_0 & ~i_13_360_3878_0));
endmodule



// Benchmark "kernel_13_361" written by ABC on Sun Jul 19 10:50:25 2020

module kernel_13_361 ( 
    i_13_361_49_0, i_13_361_50_0, i_13_361_52_0, i_13_361_71_0,
    i_13_361_94_0, i_13_361_97_0, i_13_361_98_0, i_13_361_248_0,
    i_13_361_251_0, i_13_361_259_0, i_13_361_278_0, i_13_361_310_0,
    i_13_361_319_0, i_13_361_364_0, i_13_361_521_0, i_13_361_575_0,
    i_13_361_619_0, i_13_361_620_0, i_13_361_700_0, i_13_361_800_0,
    i_13_361_889_0, i_13_361_979_0, i_13_361_980_0, i_13_361_1025_0,
    i_13_361_1079_0, i_13_361_1087_0, i_13_361_1265_0, i_13_361_1331_0,
    i_13_361_1403_0, i_13_361_1427_0, i_13_361_1429_0, i_13_361_1430_0,
    i_13_361_1435_0, i_13_361_1436_0, i_13_361_1573_0, i_13_361_1637_0,
    i_13_361_1652_0, i_13_361_1661_0, i_13_361_1664_0, i_13_361_1735_0,
    i_13_361_1736_0, i_13_361_1777_0, i_13_361_1808_0, i_13_361_1817_0,
    i_13_361_1921_0, i_13_361_1933_0, i_13_361_2023_0, i_13_361_2024_0,
    i_13_361_2030_0, i_13_361_2051_0, i_13_361_2059_0, i_13_361_2230_0,
    i_13_361_2344_0, i_13_361_2455_0, i_13_361_2456_0, i_13_361_2588_0,
    i_13_361_2716_0, i_13_361_2726_0, i_13_361_2743_0, i_13_361_2744_0,
    i_13_361_2788_0, i_13_361_2789_0, i_13_361_2959_0, i_13_361_3002_0,
    i_13_361_3032_0, i_13_361_3058_0, i_13_361_3076_0, i_13_361_3077_0,
    i_13_361_3119_0, i_13_361_3128_0, i_13_361_3272_0, i_13_361_3292_0,
    i_13_361_3316_0, i_13_361_3370_0, i_13_361_3380_0, i_13_361_3419_0,
    i_13_361_3452_0, i_13_361_3454_0, i_13_361_3464_0, i_13_361_3472_0,
    i_13_361_3481_0, i_13_361_3514_0, i_13_361_3653_0, i_13_361_3685_0,
    i_13_361_3689_0, i_13_361_3707_0, i_13_361_3802_0, i_13_361_3905_0,
    i_13_361_3923_0, i_13_361_4022_0, i_13_361_4031_0, i_13_361_4256_0,
    i_13_361_4265_0, i_13_361_4274_0, i_13_361_4336_0, i_13_361_4342_0,
    i_13_361_4391_0, i_13_361_4450_0, i_13_361_4451_0, i_13_361_4558_0,
    o_13_361_0_0  );
  input  i_13_361_49_0, i_13_361_50_0, i_13_361_52_0, i_13_361_71_0,
    i_13_361_94_0, i_13_361_97_0, i_13_361_98_0, i_13_361_248_0,
    i_13_361_251_0, i_13_361_259_0, i_13_361_278_0, i_13_361_310_0,
    i_13_361_319_0, i_13_361_364_0, i_13_361_521_0, i_13_361_575_0,
    i_13_361_619_0, i_13_361_620_0, i_13_361_700_0, i_13_361_800_0,
    i_13_361_889_0, i_13_361_979_0, i_13_361_980_0, i_13_361_1025_0,
    i_13_361_1079_0, i_13_361_1087_0, i_13_361_1265_0, i_13_361_1331_0,
    i_13_361_1403_0, i_13_361_1427_0, i_13_361_1429_0, i_13_361_1430_0,
    i_13_361_1435_0, i_13_361_1436_0, i_13_361_1573_0, i_13_361_1637_0,
    i_13_361_1652_0, i_13_361_1661_0, i_13_361_1664_0, i_13_361_1735_0,
    i_13_361_1736_0, i_13_361_1777_0, i_13_361_1808_0, i_13_361_1817_0,
    i_13_361_1921_0, i_13_361_1933_0, i_13_361_2023_0, i_13_361_2024_0,
    i_13_361_2030_0, i_13_361_2051_0, i_13_361_2059_0, i_13_361_2230_0,
    i_13_361_2344_0, i_13_361_2455_0, i_13_361_2456_0, i_13_361_2588_0,
    i_13_361_2716_0, i_13_361_2726_0, i_13_361_2743_0, i_13_361_2744_0,
    i_13_361_2788_0, i_13_361_2789_0, i_13_361_2959_0, i_13_361_3002_0,
    i_13_361_3032_0, i_13_361_3058_0, i_13_361_3076_0, i_13_361_3077_0,
    i_13_361_3119_0, i_13_361_3128_0, i_13_361_3272_0, i_13_361_3292_0,
    i_13_361_3316_0, i_13_361_3370_0, i_13_361_3380_0, i_13_361_3419_0,
    i_13_361_3452_0, i_13_361_3454_0, i_13_361_3464_0, i_13_361_3472_0,
    i_13_361_3481_0, i_13_361_3514_0, i_13_361_3653_0, i_13_361_3685_0,
    i_13_361_3689_0, i_13_361_3707_0, i_13_361_3802_0, i_13_361_3905_0,
    i_13_361_3923_0, i_13_361_4022_0, i_13_361_4031_0, i_13_361_4256_0,
    i_13_361_4265_0, i_13_361_4274_0, i_13_361_4336_0, i_13_361_4342_0,
    i_13_361_4391_0, i_13_361_4450_0, i_13_361_4451_0, i_13_361_4558_0;
  output o_13_361_0_0;
  assign o_13_361_0_0 = ~((~i_13_361_3464_0 & (~i_13_361_1430_0 | ~i_13_361_2024_0)) | (~i_13_361_521_0 & ~i_13_361_3316_0) | (~i_13_361_700_0 & ~i_13_361_4274_0) | (i_13_361_94_0 & ~i_13_361_4336_0 & ~i_13_361_4450_0));
endmodule



// Benchmark "kernel_13_362" written by ABC on Sun Jul 19 10:50:25 2020

module kernel_13_362 ( 
    i_13_362_38_0, i_13_362_40_0, i_13_362_72_0, i_13_362_73_0,
    i_13_362_108_0, i_13_362_173_0, i_13_362_226_0, i_13_362_252_0,
    i_13_362_271_0, i_13_362_355_0, i_13_362_363_0, i_13_362_364_0,
    i_13_362_441_0, i_13_362_442_0, i_13_362_453_0, i_13_362_468_0,
    i_13_362_469_0, i_13_362_558_0, i_13_362_559_0, i_13_362_643_0,
    i_13_362_666_0, i_13_362_667_0, i_13_362_732_0, i_13_362_796_0,
    i_13_362_839_0, i_13_362_945_0, i_13_362_946_0, i_13_362_947_0,
    i_13_362_1081_0, i_13_362_1099_0, i_13_362_1100_0, i_13_362_1143_0,
    i_13_362_1144_0, i_13_362_1307_0, i_13_362_1344_0, i_13_362_1407_0,
    i_13_362_1443_0, i_13_362_1620_0, i_13_362_1621_0, i_13_362_1719_0,
    i_13_362_1720_0, i_13_362_1729_0, i_13_362_1773_0, i_13_362_1802_0,
    i_13_362_1836_0, i_13_362_1837_0, i_13_362_2016_0, i_13_362_2169_0,
    i_13_362_2210_0, i_13_362_2281_0, i_13_362_2299_0, i_13_362_2358_0,
    i_13_362_2430_0, i_13_362_2431_0, i_13_362_2433_0, i_13_362_2448_0,
    i_13_362_2468_0, i_13_362_2511_0, i_13_362_2610_0, i_13_362_2611_0,
    i_13_362_2712_0, i_13_362_2719_0, i_13_362_2757_0, i_13_362_2784_0,
    i_13_362_2874_0, i_13_362_2880_0, i_13_362_2920_0, i_13_362_2955_0,
    i_13_362_3026_0, i_13_362_3033_0, i_13_362_3048_0, i_13_362_3060_0,
    i_13_362_3097_0, i_13_362_3107_0, i_13_362_3127_0, i_13_362_3162_0,
    i_13_362_3216_0, i_13_362_3231_0, i_13_362_3369_0, i_13_362_3421_0,
    i_13_362_3467_0, i_13_362_3481_0, i_13_362_3521_0, i_13_362_3528_0,
    i_13_362_3550_0, i_13_362_3592_0, i_13_362_3595_0, i_13_362_3619_0,
    i_13_362_3720_0, i_13_362_3727_0, i_13_362_3908_0, i_13_362_4126_0,
    i_13_362_4215_0, i_13_362_4258_0, i_13_362_4329_0, i_13_362_4340_0,
    i_13_362_4350_0, i_13_362_4351_0, i_13_362_4446_0, i_13_362_4540_0,
    o_13_362_0_0  );
  input  i_13_362_38_0, i_13_362_40_0, i_13_362_72_0, i_13_362_73_0,
    i_13_362_108_0, i_13_362_173_0, i_13_362_226_0, i_13_362_252_0,
    i_13_362_271_0, i_13_362_355_0, i_13_362_363_0, i_13_362_364_0,
    i_13_362_441_0, i_13_362_442_0, i_13_362_453_0, i_13_362_468_0,
    i_13_362_469_0, i_13_362_558_0, i_13_362_559_0, i_13_362_643_0,
    i_13_362_666_0, i_13_362_667_0, i_13_362_732_0, i_13_362_796_0,
    i_13_362_839_0, i_13_362_945_0, i_13_362_946_0, i_13_362_947_0,
    i_13_362_1081_0, i_13_362_1099_0, i_13_362_1100_0, i_13_362_1143_0,
    i_13_362_1144_0, i_13_362_1307_0, i_13_362_1344_0, i_13_362_1407_0,
    i_13_362_1443_0, i_13_362_1620_0, i_13_362_1621_0, i_13_362_1719_0,
    i_13_362_1720_0, i_13_362_1729_0, i_13_362_1773_0, i_13_362_1802_0,
    i_13_362_1836_0, i_13_362_1837_0, i_13_362_2016_0, i_13_362_2169_0,
    i_13_362_2210_0, i_13_362_2281_0, i_13_362_2299_0, i_13_362_2358_0,
    i_13_362_2430_0, i_13_362_2431_0, i_13_362_2433_0, i_13_362_2448_0,
    i_13_362_2468_0, i_13_362_2511_0, i_13_362_2610_0, i_13_362_2611_0,
    i_13_362_2712_0, i_13_362_2719_0, i_13_362_2757_0, i_13_362_2784_0,
    i_13_362_2874_0, i_13_362_2880_0, i_13_362_2920_0, i_13_362_2955_0,
    i_13_362_3026_0, i_13_362_3033_0, i_13_362_3048_0, i_13_362_3060_0,
    i_13_362_3097_0, i_13_362_3107_0, i_13_362_3127_0, i_13_362_3162_0,
    i_13_362_3216_0, i_13_362_3231_0, i_13_362_3369_0, i_13_362_3421_0,
    i_13_362_3467_0, i_13_362_3481_0, i_13_362_3521_0, i_13_362_3528_0,
    i_13_362_3550_0, i_13_362_3592_0, i_13_362_3595_0, i_13_362_3619_0,
    i_13_362_3720_0, i_13_362_3727_0, i_13_362_3908_0, i_13_362_4126_0,
    i_13_362_4215_0, i_13_362_4258_0, i_13_362_4329_0, i_13_362_4340_0,
    i_13_362_4350_0, i_13_362_4351_0, i_13_362_4446_0, i_13_362_4540_0;
  output o_13_362_0_0;
  assign o_13_362_0_0 = ~((~i_13_362_2757_0 & ~i_13_362_4351_0) | (~i_13_362_73_0 & ~i_13_362_945_0) | (~i_13_362_469_0 & ~i_13_362_1620_0 & ~i_13_362_1836_0));
endmodule



// Benchmark "kernel_13_363" written by ABC on Sun Jul 19 10:50:26 2020

module kernel_13_363 ( 
    i_13_363_77_0, i_13_363_94_0, i_13_363_230_0, i_13_363_259_0,
    i_13_363_518_0, i_13_363_536_0, i_13_363_554_0, i_13_363_611_0,
    i_13_363_616_0, i_13_363_627_0, i_13_363_647_0, i_13_363_655_0,
    i_13_363_664_0, i_13_363_689_0, i_13_363_692_0, i_13_363_697_0,
    i_13_363_698_0, i_13_363_700_0, i_13_363_862_0, i_13_363_943_0,
    i_13_363_980_0, i_13_363_1025_0, i_13_363_1076_0, i_13_363_1079_0,
    i_13_363_1121_0, i_13_363_1124_0, i_13_363_1183_0, i_13_363_1214_0,
    i_13_363_1304_0, i_13_363_1330_0, i_13_363_1331_0, i_13_363_1483_0,
    i_13_363_1517_0, i_13_363_1519_0, i_13_363_1678_0, i_13_363_1682_0,
    i_13_363_1735_0, i_13_363_1745_0, i_13_363_1778_0, i_13_363_1795_0,
    i_13_363_1889_0, i_13_363_1922_0, i_13_363_2024_0, i_13_363_2113_0,
    i_13_363_2209_0, i_13_363_2212_0, i_13_363_2321_0, i_13_363_2447_0,
    i_13_363_2455_0, i_13_363_2651_0, i_13_363_2654_0, i_13_363_2696_0,
    i_13_363_2851_0, i_13_363_2887_0, i_13_363_2888_0, i_13_363_2894_0,
    i_13_363_2959_0, i_13_363_3030_0, i_13_363_3037_0, i_13_363_3073_0,
    i_13_363_3091_0, i_13_363_3157_0, i_13_363_3203_0, i_13_363_3208_0,
    i_13_363_3217_0, i_13_363_3238_0, i_13_363_3265_0, i_13_363_3310_0,
    i_13_363_3418_0, i_13_363_3482_0, i_13_363_3526_0, i_13_363_3527_0,
    i_13_363_3571_0, i_13_363_3572_0, i_13_363_3695_0, i_13_363_3742_0,
    i_13_363_3743_0, i_13_363_3847_0, i_13_363_3866_0, i_13_363_3874_0,
    i_13_363_3887_0, i_13_363_3930_0, i_13_363_4045_0, i_13_363_4064_0,
    i_13_363_4081_0, i_13_363_4091_0, i_13_363_4130_0, i_13_363_4162_0,
    i_13_363_4190_0, i_13_363_4192_0, i_13_363_4193_0, i_13_363_4256_0,
    i_13_363_4270_0, i_13_363_4336_0, i_13_363_4372_0, i_13_363_4382_0,
    i_13_363_4460_0, i_13_363_4598_0, i_13_363_4603_0, i_13_363_4604_0,
    o_13_363_0_0  );
  input  i_13_363_77_0, i_13_363_94_0, i_13_363_230_0, i_13_363_259_0,
    i_13_363_518_0, i_13_363_536_0, i_13_363_554_0, i_13_363_611_0,
    i_13_363_616_0, i_13_363_627_0, i_13_363_647_0, i_13_363_655_0,
    i_13_363_664_0, i_13_363_689_0, i_13_363_692_0, i_13_363_697_0,
    i_13_363_698_0, i_13_363_700_0, i_13_363_862_0, i_13_363_943_0,
    i_13_363_980_0, i_13_363_1025_0, i_13_363_1076_0, i_13_363_1079_0,
    i_13_363_1121_0, i_13_363_1124_0, i_13_363_1183_0, i_13_363_1214_0,
    i_13_363_1304_0, i_13_363_1330_0, i_13_363_1331_0, i_13_363_1483_0,
    i_13_363_1517_0, i_13_363_1519_0, i_13_363_1678_0, i_13_363_1682_0,
    i_13_363_1735_0, i_13_363_1745_0, i_13_363_1778_0, i_13_363_1795_0,
    i_13_363_1889_0, i_13_363_1922_0, i_13_363_2024_0, i_13_363_2113_0,
    i_13_363_2209_0, i_13_363_2212_0, i_13_363_2321_0, i_13_363_2447_0,
    i_13_363_2455_0, i_13_363_2651_0, i_13_363_2654_0, i_13_363_2696_0,
    i_13_363_2851_0, i_13_363_2887_0, i_13_363_2888_0, i_13_363_2894_0,
    i_13_363_2959_0, i_13_363_3030_0, i_13_363_3037_0, i_13_363_3073_0,
    i_13_363_3091_0, i_13_363_3157_0, i_13_363_3203_0, i_13_363_3208_0,
    i_13_363_3217_0, i_13_363_3238_0, i_13_363_3265_0, i_13_363_3310_0,
    i_13_363_3418_0, i_13_363_3482_0, i_13_363_3526_0, i_13_363_3527_0,
    i_13_363_3571_0, i_13_363_3572_0, i_13_363_3695_0, i_13_363_3742_0,
    i_13_363_3743_0, i_13_363_3847_0, i_13_363_3866_0, i_13_363_3874_0,
    i_13_363_3887_0, i_13_363_3930_0, i_13_363_4045_0, i_13_363_4064_0,
    i_13_363_4081_0, i_13_363_4091_0, i_13_363_4130_0, i_13_363_4162_0,
    i_13_363_4190_0, i_13_363_4192_0, i_13_363_4193_0, i_13_363_4256_0,
    i_13_363_4270_0, i_13_363_4336_0, i_13_363_4372_0, i_13_363_4382_0,
    i_13_363_4460_0, i_13_363_4598_0, i_13_363_4603_0, i_13_363_4604_0;
  output o_13_363_0_0;
  assign o_13_363_0_0 = ~(~i_13_363_1121_0 | (i_13_363_94_0 & ~i_13_363_3526_0) | (~i_13_363_1124_0 & ~i_13_363_2887_0) | (~i_13_363_697_0 & ~i_13_363_2696_0) | (~i_13_363_536_0 & ~i_13_363_1079_0 & ~i_13_363_4064_0 & ~i_13_363_4256_0));
endmodule



// Benchmark "kernel_13_364" written by ABC on Sun Jul 19 10:50:27 2020

module kernel_13_364 ( 
    i_13_364_34_0, i_13_364_51_0, i_13_364_52_0, i_13_364_75_0,
    i_13_364_93_0, i_13_364_129_0, i_13_364_130_0, i_13_364_141_0,
    i_13_364_240_0, i_13_364_250_0, i_13_364_258_0, i_13_364_340_0,
    i_13_364_561_0, i_13_364_570_0, i_13_364_585_0, i_13_364_618_0,
    i_13_364_619_0, i_13_364_642_0, i_13_364_699_0, i_13_364_700_0,
    i_13_364_714_0, i_13_364_763_0, i_13_364_840_0, i_13_364_843_0,
    i_13_364_844_0, i_13_364_931_0, i_13_364_1077_0, i_13_364_1078_0,
    i_13_364_1342_0, i_13_364_1399_0, i_13_364_1401_0, i_13_364_1408_0,
    i_13_364_1471_0, i_13_364_1482_0, i_13_364_1527_0, i_13_364_1552_0,
    i_13_364_1572_0, i_13_364_1608_0, i_13_364_1635_0, i_13_364_1636_0,
    i_13_364_1660_0, i_13_364_1710_0, i_13_364_1734_0, i_13_364_1912_0,
    i_13_364_1920_0, i_13_364_1921_0, i_13_364_1992_0, i_13_364_2019_0,
    i_13_364_2032_0, i_13_364_2055_0, i_13_364_2277_0, i_13_364_2280_0,
    i_13_364_2311_0, i_13_364_2454_0, i_13_364_2505_0, i_13_364_2551_0,
    i_13_364_2569_0, i_13_364_2670_0, i_13_364_2724_0, i_13_364_2787_0,
    i_13_364_2847_0, i_13_364_2854_0, i_13_364_2857_0, i_13_364_2886_0,
    i_13_364_2887_0, i_13_364_2958_0, i_13_364_2959_0, i_13_364_3063_0,
    i_13_364_3145_0, i_13_364_3244_0, i_13_364_3315_0, i_13_364_3322_0,
    i_13_364_3372_0, i_13_364_3379_0, i_13_364_3382_0, i_13_364_3451_0,
    i_13_364_3463_0, i_13_364_3525_0, i_13_364_3540_0, i_13_364_3552_0,
    i_13_364_3553_0, i_13_364_3613_0, i_13_364_3630_0, i_13_364_3643_0,
    i_13_364_3646_0, i_13_364_3649_0, i_13_364_3667_0, i_13_364_3687_0,
    i_13_364_3688_0, i_13_364_3694_0, i_13_364_3724_0, i_13_364_3739_0,
    i_13_364_4104_0, i_13_364_4162_0, i_13_364_4209_0, i_13_364_4254_0,
    i_13_364_4390_0, i_13_364_4392_0, i_13_364_4393_0, i_13_364_4395_0,
    o_13_364_0_0  );
  input  i_13_364_34_0, i_13_364_51_0, i_13_364_52_0, i_13_364_75_0,
    i_13_364_93_0, i_13_364_129_0, i_13_364_130_0, i_13_364_141_0,
    i_13_364_240_0, i_13_364_250_0, i_13_364_258_0, i_13_364_340_0,
    i_13_364_561_0, i_13_364_570_0, i_13_364_585_0, i_13_364_618_0,
    i_13_364_619_0, i_13_364_642_0, i_13_364_699_0, i_13_364_700_0,
    i_13_364_714_0, i_13_364_763_0, i_13_364_840_0, i_13_364_843_0,
    i_13_364_844_0, i_13_364_931_0, i_13_364_1077_0, i_13_364_1078_0,
    i_13_364_1342_0, i_13_364_1399_0, i_13_364_1401_0, i_13_364_1408_0,
    i_13_364_1471_0, i_13_364_1482_0, i_13_364_1527_0, i_13_364_1552_0,
    i_13_364_1572_0, i_13_364_1608_0, i_13_364_1635_0, i_13_364_1636_0,
    i_13_364_1660_0, i_13_364_1710_0, i_13_364_1734_0, i_13_364_1912_0,
    i_13_364_1920_0, i_13_364_1921_0, i_13_364_1992_0, i_13_364_2019_0,
    i_13_364_2032_0, i_13_364_2055_0, i_13_364_2277_0, i_13_364_2280_0,
    i_13_364_2311_0, i_13_364_2454_0, i_13_364_2505_0, i_13_364_2551_0,
    i_13_364_2569_0, i_13_364_2670_0, i_13_364_2724_0, i_13_364_2787_0,
    i_13_364_2847_0, i_13_364_2854_0, i_13_364_2857_0, i_13_364_2886_0,
    i_13_364_2887_0, i_13_364_2958_0, i_13_364_2959_0, i_13_364_3063_0,
    i_13_364_3145_0, i_13_364_3244_0, i_13_364_3315_0, i_13_364_3322_0,
    i_13_364_3372_0, i_13_364_3379_0, i_13_364_3382_0, i_13_364_3451_0,
    i_13_364_3463_0, i_13_364_3525_0, i_13_364_3540_0, i_13_364_3552_0,
    i_13_364_3553_0, i_13_364_3613_0, i_13_364_3630_0, i_13_364_3643_0,
    i_13_364_3646_0, i_13_364_3649_0, i_13_364_3667_0, i_13_364_3687_0,
    i_13_364_3688_0, i_13_364_3694_0, i_13_364_3724_0, i_13_364_3739_0,
    i_13_364_4104_0, i_13_364_4162_0, i_13_364_4209_0, i_13_364_4254_0,
    i_13_364_4390_0, i_13_364_4392_0, i_13_364_4393_0, i_13_364_4395_0;
  output o_13_364_0_0;
  assign o_13_364_0_0 = ~((~i_13_364_2886_0 & ~i_13_364_3451_0) | (i_13_364_34_0 & ~i_13_364_1401_0) | (~i_13_364_141_0 & ~i_13_364_618_0));
endmodule



// Benchmark "kernel_13_365" written by ABC on Sun Jul 19 10:50:28 2020

module kernel_13_365 ( 
    i_13_365_39_0, i_13_365_66_0, i_13_365_75_0, i_13_365_96_0,
    i_13_365_106_0, i_13_365_168_0, i_13_365_268_0, i_13_365_284_0,
    i_13_365_357_0, i_13_365_410_0, i_13_365_411_0, i_13_365_465_0,
    i_13_365_466_0, i_13_365_515_0, i_13_365_529_0, i_13_365_569_0,
    i_13_365_591_0, i_13_365_592_0, i_13_365_654_0, i_13_365_794_0,
    i_13_365_824_0, i_13_365_914_0, i_13_365_1019_0, i_13_365_1021_0,
    i_13_365_1118_0, i_13_365_1212_0, i_13_365_1229_0, i_13_365_1347_0,
    i_13_365_1348_0, i_13_365_1391_0, i_13_365_1409_0, i_13_365_1443_0,
    i_13_365_1446_0, i_13_365_1490_0, i_13_365_1492_0, i_13_365_1501_0,
    i_13_365_1596_0, i_13_365_1713_0, i_13_365_1776_0, i_13_365_1777_0,
    i_13_365_1802_0, i_13_365_1884_0, i_13_365_1931_0, i_13_365_1950_0,
    i_13_365_1960_0, i_13_365_2032_0, i_13_365_2058_0, i_13_365_2059_0,
    i_13_365_2103_0, i_13_365_2110_0, i_13_365_2202_0, i_13_365_2283_0,
    i_13_365_2284_0, i_13_365_2347_0, i_13_365_2409_0, i_13_365_2410_0,
    i_13_365_2444_0, i_13_365_2446_0, i_13_365_2465_0, i_13_365_2514_0,
    i_13_365_2553_0, i_13_365_2554_0, i_13_365_3173_0, i_13_365_3215_0,
    i_13_365_3263_0, i_13_365_3353_0, i_13_365_3372_0, i_13_365_3373_0,
    i_13_365_3390_0, i_13_365_3391_0, i_13_365_3418_0, i_13_365_3425_0,
    i_13_365_3530_0, i_13_365_3535_0, i_13_365_3579_0, i_13_365_3597_0,
    i_13_365_3598_0, i_13_365_3621_0, i_13_365_3633_0, i_13_365_3638_0,
    i_13_365_3755_0, i_13_365_3783_0, i_13_365_3784_0, i_13_365_3785_0,
    i_13_365_3786_0, i_13_365_3787_0, i_13_365_3800_0, i_13_365_3874_0,
    i_13_365_3983_0, i_13_365_3990_0, i_13_365_4236_0, i_13_365_4250_0,
    i_13_365_4263_0, i_13_365_4264_0, i_13_365_4332_0, i_13_365_4367_0,
    i_13_365_4432_0, i_13_365_4452_0, i_13_365_4453_0, i_13_365_4543_0,
    o_13_365_0_0  );
  input  i_13_365_39_0, i_13_365_66_0, i_13_365_75_0, i_13_365_96_0,
    i_13_365_106_0, i_13_365_168_0, i_13_365_268_0, i_13_365_284_0,
    i_13_365_357_0, i_13_365_410_0, i_13_365_411_0, i_13_365_465_0,
    i_13_365_466_0, i_13_365_515_0, i_13_365_529_0, i_13_365_569_0,
    i_13_365_591_0, i_13_365_592_0, i_13_365_654_0, i_13_365_794_0,
    i_13_365_824_0, i_13_365_914_0, i_13_365_1019_0, i_13_365_1021_0,
    i_13_365_1118_0, i_13_365_1212_0, i_13_365_1229_0, i_13_365_1347_0,
    i_13_365_1348_0, i_13_365_1391_0, i_13_365_1409_0, i_13_365_1443_0,
    i_13_365_1446_0, i_13_365_1490_0, i_13_365_1492_0, i_13_365_1501_0,
    i_13_365_1596_0, i_13_365_1713_0, i_13_365_1776_0, i_13_365_1777_0,
    i_13_365_1802_0, i_13_365_1884_0, i_13_365_1931_0, i_13_365_1950_0,
    i_13_365_1960_0, i_13_365_2032_0, i_13_365_2058_0, i_13_365_2059_0,
    i_13_365_2103_0, i_13_365_2110_0, i_13_365_2202_0, i_13_365_2283_0,
    i_13_365_2284_0, i_13_365_2347_0, i_13_365_2409_0, i_13_365_2410_0,
    i_13_365_2444_0, i_13_365_2446_0, i_13_365_2465_0, i_13_365_2514_0,
    i_13_365_2553_0, i_13_365_2554_0, i_13_365_3173_0, i_13_365_3215_0,
    i_13_365_3263_0, i_13_365_3353_0, i_13_365_3372_0, i_13_365_3373_0,
    i_13_365_3390_0, i_13_365_3391_0, i_13_365_3418_0, i_13_365_3425_0,
    i_13_365_3530_0, i_13_365_3535_0, i_13_365_3579_0, i_13_365_3597_0,
    i_13_365_3598_0, i_13_365_3621_0, i_13_365_3633_0, i_13_365_3638_0,
    i_13_365_3755_0, i_13_365_3783_0, i_13_365_3784_0, i_13_365_3785_0,
    i_13_365_3786_0, i_13_365_3787_0, i_13_365_3800_0, i_13_365_3874_0,
    i_13_365_3983_0, i_13_365_3990_0, i_13_365_4236_0, i_13_365_4250_0,
    i_13_365_4263_0, i_13_365_4264_0, i_13_365_4332_0, i_13_365_4367_0,
    i_13_365_4432_0, i_13_365_4452_0, i_13_365_4453_0, i_13_365_4543_0;
  output o_13_365_0_0;
  assign o_13_365_0_0 = ~(~i_13_365_1950_0 | ~i_13_365_3391_0);
endmodule



// Benchmark "kernel_13_366" written by ABC on Sun Jul 19 10:50:29 2020

module kernel_13_366 ( 
    i_13_366_46_0, i_13_366_119_0, i_13_366_154_0, i_13_366_157_0,
    i_13_366_164_0, i_13_366_167_0, i_13_366_214_0, i_13_366_259_0,
    i_13_366_269_0, i_13_366_275_0, i_13_366_278_0, i_13_366_334_0,
    i_13_366_352_0, i_13_366_353_0, i_13_366_451_0, i_13_366_455_0,
    i_13_366_506_0, i_13_366_518_0, i_13_366_617_0, i_13_366_667_0,
    i_13_366_814_0, i_13_366_815_0, i_13_366_841_0, i_13_366_845_0,
    i_13_366_932_0, i_13_366_961_0, i_13_366_977_0, i_13_366_1066_0,
    i_13_366_1103_0, i_13_366_1244_0, i_13_366_1327_0, i_13_366_1342_0,
    i_13_366_1400_0, i_13_366_1402_0, i_13_366_1445_0, i_13_366_1480_0,
    i_13_366_1508_0, i_13_366_1543_0, i_13_366_1570_0, i_13_366_1573_0,
    i_13_366_1594_0, i_13_366_1604_0, i_13_366_1649_0, i_13_366_1766_0,
    i_13_366_1801_0, i_13_366_1805_0, i_13_366_1807_0, i_13_366_1850_0,
    i_13_366_1852_0, i_13_366_1931_0, i_13_366_1946_0, i_13_366_2026_0,
    i_13_366_2146_0, i_13_366_2149_0, i_13_366_2201_0, i_13_366_2237_0,
    i_13_366_2278_0, i_13_366_2303_0, i_13_366_2408_0, i_13_366_2569_0,
    i_13_366_2585_0, i_13_366_2591_0, i_13_366_2600_0, i_13_366_2621_0,
    i_13_366_2768_0, i_13_366_2899_0, i_13_366_2965_0, i_13_366_2972_0,
    i_13_366_3106_0, i_13_366_3112_0, i_13_366_3127_0, i_13_366_3128_0,
    i_13_366_3215_0, i_13_366_3274_0, i_13_366_3313_0, i_13_366_3379_0,
    i_13_366_3397_0, i_13_366_3398_0, i_13_366_3400_0, i_13_366_3439_0,
    i_13_366_3521_0, i_13_366_3592_0, i_13_366_3628_0, i_13_366_3664_0,
    i_13_366_3739_0, i_13_366_3821_0, i_13_366_3889_0, i_13_366_3899_0,
    i_13_366_4042_0, i_13_366_4043_0, i_13_366_4061_0, i_13_366_4063_0,
    i_13_366_4231_0, i_13_366_4253_0, i_13_366_4318_0, i_13_366_4319_0,
    i_13_366_4348_0, i_13_366_4375_0, i_13_366_4534_0, i_13_366_4556_0,
    o_13_366_0_0  );
  input  i_13_366_46_0, i_13_366_119_0, i_13_366_154_0, i_13_366_157_0,
    i_13_366_164_0, i_13_366_167_0, i_13_366_214_0, i_13_366_259_0,
    i_13_366_269_0, i_13_366_275_0, i_13_366_278_0, i_13_366_334_0,
    i_13_366_352_0, i_13_366_353_0, i_13_366_451_0, i_13_366_455_0,
    i_13_366_506_0, i_13_366_518_0, i_13_366_617_0, i_13_366_667_0,
    i_13_366_814_0, i_13_366_815_0, i_13_366_841_0, i_13_366_845_0,
    i_13_366_932_0, i_13_366_961_0, i_13_366_977_0, i_13_366_1066_0,
    i_13_366_1103_0, i_13_366_1244_0, i_13_366_1327_0, i_13_366_1342_0,
    i_13_366_1400_0, i_13_366_1402_0, i_13_366_1445_0, i_13_366_1480_0,
    i_13_366_1508_0, i_13_366_1543_0, i_13_366_1570_0, i_13_366_1573_0,
    i_13_366_1594_0, i_13_366_1604_0, i_13_366_1649_0, i_13_366_1766_0,
    i_13_366_1801_0, i_13_366_1805_0, i_13_366_1807_0, i_13_366_1850_0,
    i_13_366_1852_0, i_13_366_1931_0, i_13_366_1946_0, i_13_366_2026_0,
    i_13_366_2146_0, i_13_366_2149_0, i_13_366_2201_0, i_13_366_2237_0,
    i_13_366_2278_0, i_13_366_2303_0, i_13_366_2408_0, i_13_366_2569_0,
    i_13_366_2585_0, i_13_366_2591_0, i_13_366_2600_0, i_13_366_2621_0,
    i_13_366_2768_0, i_13_366_2899_0, i_13_366_2965_0, i_13_366_2972_0,
    i_13_366_3106_0, i_13_366_3112_0, i_13_366_3127_0, i_13_366_3128_0,
    i_13_366_3215_0, i_13_366_3274_0, i_13_366_3313_0, i_13_366_3379_0,
    i_13_366_3397_0, i_13_366_3398_0, i_13_366_3400_0, i_13_366_3439_0,
    i_13_366_3521_0, i_13_366_3592_0, i_13_366_3628_0, i_13_366_3664_0,
    i_13_366_3739_0, i_13_366_3821_0, i_13_366_3889_0, i_13_366_3899_0,
    i_13_366_4042_0, i_13_366_4043_0, i_13_366_4061_0, i_13_366_4063_0,
    i_13_366_4231_0, i_13_366_4253_0, i_13_366_4318_0, i_13_366_4319_0,
    i_13_366_4348_0, i_13_366_4375_0, i_13_366_4534_0, i_13_366_4556_0;
  output o_13_366_0_0;
  assign o_13_366_0_0 = ~((~i_13_366_334_0 & i_13_366_4375_0) | (~i_13_366_1400_0 & ~i_13_366_3313_0) | (~i_13_366_352_0 & ~i_13_366_1852_0) | (~i_13_366_46_0 & ~i_13_366_1805_0) | (~i_13_366_814_0 & ~i_13_366_1931_0 & ~i_13_366_4375_0) | (~i_13_366_3398_0 & ~i_13_366_3439_0 & ~i_13_366_4348_0) | (~i_13_366_1508_0 & ~i_13_366_3592_0 & ~i_13_366_4253_0));
endmodule



// Benchmark "kernel_13_367" written by ABC on Sun Jul 19 10:50:30 2020

module kernel_13_367 ( 
    i_13_367_139_0, i_13_367_357_0, i_13_367_382_0, i_13_367_399_0,
    i_13_367_409_0, i_13_367_441_0, i_13_367_456_0, i_13_367_468_0,
    i_13_367_472_0, i_13_367_478_0, i_13_367_572_0, i_13_367_594_0,
    i_13_367_605_0, i_13_367_622_0, i_13_367_652_0, i_13_367_654_0,
    i_13_367_657_0, i_13_367_660_0, i_13_367_661_0, i_13_367_663_0,
    i_13_367_885_0, i_13_367_889_0, i_13_367_939_0, i_13_367_943_0,
    i_13_367_1076_0, i_13_367_1114_0, i_13_367_1119_0, i_13_367_1143_0,
    i_13_367_1144_0, i_13_367_1147_0, i_13_367_1270_0, i_13_367_1515_0,
    i_13_367_1656_0, i_13_367_1657_0, i_13_367_1660_0, i_13_367_1723_0,
    i_13_367_1734_0, i_13_367_1741_0, i_13_367_1768_0, i_13_367_1791_0,
    i_13_367_1792_0, i_13_367_1832_0, i_13_367_1922_0, i_13_367_2002_0,
    i_13_367_2016_0, i_13_367_2017_0, i_13_367_2019_0, i_13_367_2020_0,
    i_13_367_2023_0, i_13_367_2057_0, i_13_367_2131_0, i_13_367_2295_0,
    i_13_367_2320_0, i_13_367_2407_0, i_13_367_2461_0, i_13_367_2469_0,
    i_13_367_2470_0, i_13_367_2512_0, i_13_367_2534_0, i_13_367_2819_0,
    i_13_367_2847_0, i_13_367_2955_0, i_13_367_2958_0, i_13_367_3057_0,
    i_13_367_3075_0, i_13_367_3115_0, i_13_367_3259_0, i_13_367_3352_0,
    i_13_367_3418_0, i_13_367_3486_0, i_13_367_3489_0, i_13_367_3658_0,
    i_13_367_3666_0, i_13_367_3729_0, i_13_367_3730_0, i_13_367_3739_0,
    i_13_367_3742_0, i_13_367_3756_0, i_13_367_3865_0, i_13_367_3901_0,
    i_13_367_3903_0, i_13_367_3909_0, i_13_367_3910_0, i_13_367_3924_0,
    i_13_367_4161_0, i_13_367_4162_0, i_13_367_4165_0, i_13_367_4186_0,
    i_13_367_4217_0, i_13_367_4315_0, i_13_367_4330_0, i_13_367_4332_0,
    i_13_367_4363_0, i_13_367_4429_0, i_13_367_4432_0, i_13_367_4516_0,
    i_13_367_4591_0, i_13_367_4599_0, i_13_367_4600_0, i_13_367_4602_0,
    o_13_367_0_0  );
  input  i_13_367_139_0, i_13_367_357_0, i_13_367_382_0, i_13_367_399_0,
    i_13_367_409_0, i_13_367_441_0, i_13_367_456_0, i_13_367_468_0,
    i_13_367_472_0, i_13_367_478_0, i_13_367_572_0, i_13_367_594_0,
    i_13_367_605_0, i_13_367_622_0, i_13_367_652_0, i_13_367_654_0,
    i_13_367_657_0, i_13_367_660_0, i_13_367_661_0, i_13_367_663_0,
    i_13_367_885_0, i_13_367_889_0, i_13_367_939_0, i_13_367_943_0,
    i_13_367_1076_0, i_13_367_1114_0, i_13_367_1119_0, i_13_367_1143_0,
    i_13_367_1144_0, i_13_367_1147_0, i_13_367_1270_0, i_13_367_1515_0,
    i_13_367_1656_0, i_13_367_1657_0, i_13_367_1660_0, i_13_367_1723_0,
    i_13_367_1734_0, i_13_367_1741_0, i_13_367_1768_0, i_13_367_1791_0,
    i_13_367_1792_0, i_13_367_1832_0, i_13_367_1922_0, i_13_367_2002_0,
    i_13_367_2016_0, i_13_367_2017_0, i_13_367_2019_0, i_13_367_2020_0,
    i_13_367_2023_0, i_13_367_2057_0, i_13_367_2131_0, i_13_367_2295_0,
    i_13_367_2320_0, i_13_367_2407_0, i_13_367_2461_0, i_13_367_2469_0,
    i_13_367_2470_0, i_13_367_2512_0, i_13_367_2534_0, i_13_367_2819_0,
    i_13_367_2847_0, i_13_367_2955_0, i_13_367_2958_0, i_13_367_3057_0,
    i_13_367_3075_0, i_13_367_3115_0, i_13_367_3259_0, i_13_367_3352_0,
    i_13_367_3418_0, i_13_367_3486_0, i_13_367_3489_0, i_13_367_3658_0,
    i_13_367_3666_0, i_13_367_3729_0, i_13_367_3730_0, i_13_367_3739_0,
    i_13_367_3742_0, i_13_367_3756_0, i_13_367_3865_0, i_13_367_3901_0,
    i_13_367_3903_0, i_13_367_3909_0, i_13_367_3910_0, i_13_367_3924_0,
    i_13_367_4161_0, i_13_367_4162_0, i_13_367_4165_0, i_13_367_4186_0,
    i_13_367_4217_0, i_13_367_4315_0, i_13_367_4330_0, i_13_367_4332_0,
    i_13_367_4363_0, i_13_367_4429_0, i_13_367_4432_0, i_13_367_4516_0,
    i_13_367_4591_0, i_13_367_4599_0, i_13_367_4600_0, i_13_367_4602_0;
  output o_13_367_0_0;
  assign o_13_367_0_0 = ~((~i_13_367_4432_0 & ((~i_13_367_1791_0 & ((~i_13_367_2016_0 & ~i_13_367_4162_0) | (i_13_367_2002_0 & ~i_13_367_4161_0 & ~i_13_367_4429_0))) | (~i_13_367_441_0 & ~i_13_367_2017_0 & ~i_13_367_3865_0) | (~i_13_367_1660_0 & i_13_367_4315_0))) | (i_13_367_382_0 & ~i_13_367_885_0 & ~i_13_367_4162_0) | (~i_13_367_1792_0 & ~i_13_367_3756_0 & ~i_13_367_3865_0) | (~i_13_367_1144_0 & ~i_13_367_2016_0 & ~i_13_367_2847_0 & ~i_13_367_3901_0 & ~i_13_367_3903_0 & ~i_13_367_4363_0));
endmodule



// Benchmark "kernel_13_368" written by ABC on Sun Jul 19 10:50:31 2020

module kernel_13_368 ( 
    i_13_368_25_0, i_13_368_28_0, i_13_368_64_0, i_13_368_65_0,
    i_13_368_131_0, i_13_368_156_0, i_13_368_212_0, i_13_368_253_0,
    i_13_368_308_0, i_13_368_356_0, i_13_368_373_0, i_13_368_376_0,
    i_13_368_397_0, i_13_368_469_0, i_13_368_524_0, i_13_368_535_0,
    i_13_368_667_0, i_13_368_668_0, i_13_368_712_0, i_13_368_725_0,
    i_13_368_758_0, i_13_368_829_0, i_13_368_830_0, i_13_368_850_0,
    i_13_368_896_0, i_13_368_929_0, i_13_368_947_0, i_13_368_1081_0,
    i_13_368_1082_0, i_13_368_1099_0, i_13_368_1246_0, i_13_368_1273_0,
    i_13_368_1274_0, i_13_368_1306_0, i_13_368_1307_0, i_13_368_1397_0,
    i_13_368_1443_0, i_13_368_1504_0, i_13_368_1505_0, i_13_368_1550_0,
    i_13_368_1639_0, i_13_368_1714_0, i_13_368_1721_0, i_13_368_1723_0,
    i_13_368_1774_0, i_13_368_1786_0, i_13_368_1838_0, i_13_368_1847_0,
    i_13_368_1918_0, i_13_368_1927_0, i_13_368_1999_0, i_13_368_2000_0,
    i_13_368_2030_0, i_13_368_2101_0, i_13_368_2297_0, i_13_368_2378_0,
    i_13_368_2395_0, i_13_368_2468_0, i_13_368_2507_0, i_13_368_2512_0,
    i_13_368_2693_0, i_13_368_2764_0, i_13_368_2875_0, i_13_368_2881_0,
    i_13_368_2935_0, i_13_368_2936_0, i_13_368_2938_0, i_13_368_3001_0,
    i_13_368_3037_0, i_13_368_3241_0, i_13_368_3242_0, i_13_368_3251_0,
    i_13_368_3259_0, i_13_368_3290_0, i_13_368_3376_0, i_13_368_3377_0,
    i_13_368_3397_0, i_13_368_3415_0, i_13_368_3529_0, i_13_368_3596_0,
    i_13_368_3620_0, i_13_368_3728_0, i_13_368_3730_0, i_13_368_3754_0,
    i_13_368_3755_0, i_13_368_3857_0, i_13_368_3935_0, i_13_368_3988_0,
    i_13_368_4060_0, i_13_368_4213_0, i_13_368_4262_0, i_13_368_4313_0,
    i_13_368_4330_0, i_13_368_4340_0, i_13_368_4341_0, i_13_368_4429_0,
    i_13_368_4430_0, i_13_368_4448_0, i_13_368_4511_0, i_13_368_4592_0,
    o_13_368_0_0  );
  input  i_13_368_25_0, i_13_368_28_0, i_13_368_64_0, i_13_368_65_0,
    i_13_368_131_0, i_13_368_156_0, i_13_368_212_0, i_13_368_253_0,
    i_13_368_308_0, i_13_368_356_0, i_13_368_373_0, i_13_368_376_0,
    i_13_368_397_0, i_13_368_469_0, i_13_368_524_0, i_13_368_535_0,
    i_13_368_667_0, i_13_368_668_0, i_13_368_712_0, i_13_368_725_0,
    i_13_368_758_0, i_13_368_829_0, i_13_368_830_0, i_13_368_850_0,
    i_13_368_896_0, i_13_368_929_0, i_13_368_947_0, i_13_368_1081_0,
    i_13_368_1082_0, i_13_368_1099_0, i_13_368_1246_0, i_13_368_1273_0,
    i_13_368_1274_0, i_13_368_1306_0, i_13_368_1307_0, i_13_368_1397_0,
    i_13_368_1443_0, i_13_368_1504_0, i_13_368_1505_0, i_13_368_1550_0,
    i_13_368_1639_0, i_13_368_1714_0, i_13_368_1721_0, i_13_368_1723_0,
    i_13_368_1774_0, i_13_368_1786_0, i_13_368_1838_0, i_13_368_1847_0,
    i_13_368_1918_0, i_13_368_1927_0, i_13_368_1999_0, i_13_368_2000_0,
    i_13_368_2030_0, i_13_368_2101_0, i_13_368_2297_0, i_13_368_2378_0,
    i_13_368_2395_0, i_13_368_2468_0, i_13_368_2507_0, i_13_368_2512_0,
    i_13_368_2693_0, i_13_368_2764_0, i_13_368_2875_0, i_13_368_2881_0,
    i_13_368_2935_0, i_13_368_2936_0, i_13_368_2938_0, i_13_368_3001_0,
    i_13_368_3037_0, i_13_368_3241_0, i_13_368_3242_0, i_13_368_3251_0,
    i_13_368_3259_0, i_13_368_3290_0, i_13_368_3376_0, i_13_368_3377_0,
    i_13_368_3397_0, i_13_368_3415_0, i_13_368_3529_0, i_13_368_3596_0,
    i_13_368_3620_0, i_13_368_3728_0, i_13_368_3730_0, i_13_368_3754_0,
    i_13_368_3755_0, i_13_368_3857_0, i_13_368_3935_0, i_13_368_3988_0,
    i_13_368_4060_0, i_13_368_4213_0, i_13_368_4262_0, i_13_368_4313_0,
    i_13_368_4330_0, i_13_368_4340_0, i_13_368_4341_0, i_13_368_4429_0,
    i_13_368_4430_0, i_13_368_4448_0, i_13_368_4511_0, i_13_368_4592_0;
  output o_13_368_0_0;
  assign o_13_368_0_0 = ~((~i_13_368_3730_0 & (~i_13_368_469_0 | (~i_13_368_2881_0 & ~i_13_368_3857_0))) | (~i_13_368_830_0 & ~i_13_368_1504_0) | (~i_13_368_667_0 & ~i_13_368_3529_0 & ~i_13_368_3728_0));
endmodule



// Benchmark "kernel_13_369" written by ABC on Sun Jul 19 10:50:32 2020

module kernel_13_369 ( 
    i_13_369_48_0, i_13_369_126_0, i_13_369_127_0, i_13_369_159_0,
    i_13_369_162_0, i_13_369_188_0, i_13_369_210_0, i_13_369_275_0,
    i_13_369_318_0, i_13_369_431_0, i_13_369_456_0, i_13_369_465_0,
    i_13_369_519_0, i_13_369_520_0, i_13_369_535_0, i_13_369_665_0,
    i_13_369_679_0, i_13_369_744_0, i_13_369_762_0, i_13_369_763_0,
    i_13_369_823_0, i_13_369_939_0, i_13_369_944_0, i_13_369_1103_0,
    i_13_369_1131_0, i_13_369_1132_0, i_13_369_1230_0, i_13_369_1303_0,
    i_13_369_1320_0, i_13_369_1392_0, i_13_369_1524_0, i_13_369_1525_0,
    i_13_369_1551_0, i_13_369_1555_0, i_13_369_1556_0, i_13_369_1602_0,
    i_13_369_1605_0, i_13_369_1606_0, i_13_369_1698_0, i_13_369_1699_0,
    i_13_369_1753_0, i_13_369_1803_0, i_13_369_1806_0, i_13_369_1903_0,
    i_13_369_1961_0, i_13_369_1998_0, i_13_369_2025_0, i_13_369_2106_0,
    i_13_369_2145_0, i_13_369_2239_0, i_13_369_2277_0, i_13_369_2299_0,
    i_13_369_2400_0, i_13_369_2472_0, i_13_369_2473_0, i_13_369_2508_0,
    i_13_369_2709_0, i_13_369_2724_0, i_13_369_2787_0, i_13_369_3075_0,
    i_13_369_3076_0, i_13_369_3144_0, i_13_369_3198_0, i_13_369_3234_0,
    i_13_369_3263_0, i_13_369_3264_0, i_13_369_3345_0, i_13_369_3366_0,
    i_13_369_3368_0, i_13_369_3399_0, i_13_369_3402_0, i_13_369_3460_0,
    i_13_369_3553_0, i_13_369_3581_0, i_13_369_3639_0, i_13_369_3640_0,
    i_13_369_3744_0, i_13_369_3780_0, i_13_369_3788_0, i_13_369_3822_0,
    i_13_369_3823_0, i_13_369_3867_0, i_13_369_3891_0, i_13_369_3900_0,
    i_13_369_3914_0, i_13_369_3922_0, i_13_369_3933_0, i_13_369_4038_0,
    i_13_369_4062_0, i_13_369_4206_0, i_13_369_4252_0, i_13_369_4256_0,
    i_13_369_4272_0, i_13_369_4341_0, i_13_369_4342_0, i_13_369_4448_0,
    i_13_369_4514_0, i_13_369_4517_0, i_13_369_4576_0, i_13_369_4596_0,
    o_13_369_0_0  );
  input  i_13_369_48_0, i_13_369_126_0, i_13_369_127_0, i_13_369_159_0,
    i_13_369_162_0, i_13_369_188_0, i_13_369_210_0, i_13_369_275_0,
    i_13_369_318_0, i_13_369_431_0, i_13_369_456_0, i_13_369_465_0,
    i_13_369_519_0, i_13_369_520_0, i_13_369_535_0, i_13_369_665_0,
    i_13_369_679_0, i_13_369_744_0, i_13_369_762_0, i_13_369_763_0,
    i_13_369_823_0, i_13_369_939_0, i_13_369_944_0, i_13_369_1103_0,
    i_13_369_1131_0, i_13_369_1132_0, i_13_369_1230_0, i_13_369_1303_0,
    i_13_369_1320_0, i_13_369_1392_0, i_13_369_1524_0, i_13_369_1525_0,
    i_13_369_1551_0, i_13_369_1555_0, i_13_369_1556_0, i_13_369_1602_0,
    i_13_369_1605_0, i_13_369_1606_0, i_13_369_1698_0, i_13_369_1699_0,
    i_13_369_1753_0, i_13_369_1803_0, i_13_369_1806_0, i_13_369_1903_0,
    i_13_369_1961_0, i_13_369_1998_0, i_13_369_2025_0, i_13_369_2106_0,
    i_13_369_2145_0, i_13_369_2239_0, i_13_369_2277_0, i_13_369_2299_0,
    i_13_369_2400_0, i_13_369_2472_0, i_13_369_2473_0, i_13_369_2508_0,
    i_13_369_2709_0, i_13_369_2724_0, i_13_369_2787_0, i_13_369_3075_0,
    i_13_369_3076_0, i_13_369_3144_0, i_13_369_3198_0, i_13_369_3234_0,
    i_13_369_3263_0, i_13_369_3264_0, i_13_369_3345_0, i_13_369_3366_0,
    i_13_369_3368_0, i_13_369_3399_0, i_13_369_3402_0, i_13_369_3460_0,
    i_13_369_3553_0, i_13_369_3581_0, i_13_369_3639_0, i_13_369_3640_0,
    i_13_369_3744_0, i_13_369_3780_0, i_13_369_3788_0, i_13_369_3822_0,
    i_13_369_3823_0, i_13_369_3867_0, i_13_369_3891_0, i_13_369_3900_0,
    i_13_369_3914_0, i_13_369_3922_0, i_13_369_3933_0, i_13_369_4038_0,
    i_13_369_4062_0, i_13_369_4206_0, i_13_369_4252_0, i_13_369_4256_0,
    i_13_369_4272_0, i_13_369_4341_0, i_13_369_4342_0, i_13_369_4448_0,
    i_13_369_4514_0, i_13_369_4517_0, i_13_369_4576_0, i_13_369_4596_0;
  output o_13_369_0_0;
  assign o_13_369_0_0 = ~((~i_13_369_4038_0 & ~i_13_369_4514_0) | (~i_13_369_1606_0 & ~i_13_369_4252_0) | (~i_13_369_1524_0 & ~i_13_369_3234_0 & ~i_13_369_3914_0) | (~i_13_369_1753_0 & ~i_13_369_3345_0 & ~i_13_369_3900_0) | (~i_13_369_465_0 & ~i_13_369_520_0 & ~i_13_369_3399_0));
endmodule



// Benchmark "kernel_13_370" written by ABC on Sun Jul 19 10:50:32 2020

module kernel_13_370 ( 
    i_13_370_69_0, i_13_370_282_0, i_13_370_285_0, i_13_370_321_0,
    i_13_370_327_0, i_13_370_328_0, i_13_370_411_0, i_13_370_448_0,
    i_13_370_457_0, i_13_370_528_0, i_13_370_529_0, i_13_370_573_0,
    i_13_370_579_0, i_13_370_598_0, i_13_370_601_0, i_13_370_640_0,
    i_13_370_676_0, i_13_370_717_0, i_13_370_745_0, i_13_370_762_0,
    i_13_370_780_0, i_13_370_825_0, i_13_370_826_0, i_13_370_861_0,
    i_13_370_862_0, i_13_370_894_0, i_13_370_913_0, i_13_370_1023_0,
    i_13_370_1024_0, i_13_370_1095_0, i_13_370_1134_0, i_13_370_1182_0,
    i_13_370_1230_0, i_13_370_1258_0, i_13_370_1320_0, i_13_370_1326_0,
    i_13_370_1347_0, i_13_370_1410_0, i_13_370_1464_0, i_13_370_1635_0,
    i_13_370_1636_0, i_13_370_1690_0, i_13_370_1713_0, i_13_370_1732_0,
    i_13_370_1749_0, i_13_370_1816_0, i_13_370_1858_0, i_13_370_1861_0,
    i_13_370_1884_0, i_13_370_1923_0, i_13_370_2005_0, i_13_370_2110_0,
    i_13_370_2139_0, i_13_370_2310_0, i_13_370_2454_0, i_13_370_2461_0,
    i_13_370_2464_0, i_13_370_2502_0, i_13_370_2544_0, i_13_370_2545_0,
    i_13_370_2559_0, i_13_370_2616_0, i_13_370_2632_0, i_13_370_2652_0,
    i_13_370_2653_0, i_13_370_2770_0, i_13_370_2874_0, i_13_370_3001_0,
    i_13_370_3088_0, i_13_370_3174_0, i_13_370_3175_0, i_13_370_3219_0,
    i_13_370_3321_0, i_13_370_3370_0, i_13_370_3399_0, i_13_370_3432_0,
    i_13_370_3562_0, i_13_370_3565_0, i_13_370_3630_0, i_13_370_3640_0,
    i_13_370_3721_0, i_13_370_3732_0, i_13_370_3793_0, i_13_370_3858_0,
    i_13_370_3876_0, i_13_370_3912_0, i_13_370_3913_0, i_13_370_3922_0,
    i_13_370_3924_0, i_13_370_4015_0, i_13_370_4078_0, i_13_370_4237_0,
    i_13_370_4254_0, i_13_370_4255_0, i_13_370_4263_0, i_13_370_4350_0,
    i_13_370_4380_0, i_13_370_4381_0, i_13_370_4443_0, i_13_370_4567_0,
    o_13_370_0_0  );
  input  i_13_370_69_0, i_13_370_282_0, i_13_370_285_0, i_13_370_321_0,
    i_13_370_327_0, i_13_370_328_0, i_13_370_411_0, i_13_370_448_0,
    i_13_370_457_0, i_13_370_528_0, i_13_370_529_0, i_13_370_573_0,
    i_13_370_579_0, i_13_370_598_0, i_13_370_601_0, i_13_370_640_0,
    i_13_370_676_0, i_13_370_717_0, i_13_370_745_0, i_13_370_762_0,
    i_13_370_780_0, i_13_370_825_0, i_13_370_826_0, i_13_370_861_0,
    i_13_370_862_0, i_13_370_894_0, i_13_370_913_0, i_13_370_1023_0,
    i_13_370_1024_0, i_13_370_1095_0, i_13_370_1134_0, i_13_370_1182_0,
    i_13_370_1230_0, i_13_370_1258_0, i_13_370_1320_0, i_13_370_1326_0,
    i_13_370_1347_0, i_13_370_1410_0, i_13_370_1464_0, i_13_370_1635_0,
    i_13_370_1636_0, i_13_370_1690_0, i_13_370_1713_0, i_13_370_1732_0,
    i_13_370_1749_0, i_13_370_1816_0, i_13_370_1858_0, i_13_370_1861_0,
    i_13_370_1884_0, i_13_370_1923_0, i_13_370_2005_0, i_13_370_2110_0,
    i_13_370_2139_0, i_13_370_2310_0, i_13_370_2454_0, i_13_370_2461_0,
    i_13_370_2464_0, i_13_370_2502_0, i_13_370_2544_0, i_13_370_2545_0,
    i_13_370_2559_0, i_13_370_2616_0, i_13_370_2632_0, i_13_370_2652_0,
    i_13_370_2653_0, i_13_370_2770_0, i_13_370_2874_0, i_13_370_3001_0,
    i_13_370_3088_0, i_13_370_3174_0, i_13_370_3175_0, i_13_370_3219_0,
    i_13_370_3321_0, i_13_370_3370_0, i_13_370_3399_0, i_13_370_3432_0,
    i_13_370_3562_0, i_13_370_3565_0, i_13_370_3630_0, i_13_370_3640_0,
    i_13_370_3721_0, i_13_370_3732_0, i_13_370_3793_0, i_13_370_3858_0,
    i_13_370_3876_0, i_13_370_3912_0, i_13_370_3913_0, i_13_370_3922_0,
    i_13_370_3924_0, i_13_370_4015_0, i_13_370_4078_0, i_13_370_4237_0,
    i_13_370_4254_0, i_13_370_4255_0, i_13_370_4263_0, i_13_370_4350_0,
    i_13_370_4380_0, i_13_370_4381_0, i_13_370_4443_0, i_13_370_4567_0;
  output o_13_370_0_0;
  assign o_13_370_0_0 = ~(~i_13_370_327_0 | ~i_13_370_3175_0);
endmodule



// Benchmark "kernel_13_371" written by ABC on Sun Jul 19 10:50:33 2020

module kernel_13_371 ( 
    i_13_371_69_0, i_13_371_70_0, i_13_371_94_0, i_13_371_258_0,
    i_13_371_372_0, i_13_371_373_0, i_13_371_645_0, i_13_371_673_0,
    i_13_371_686_0, i_13_371_797_0, i_13_371_820_0, i_13_371_921_0,
    i_13_371_1065_0, i_13_371_1103_0, i_13_371_1104_0, i_13_371_1148_0,
    i_13_371_1274_0, i_13_371_1275_0, i_13_371_1276_0, i_13_371_1297_0,
    i_13_371_1317_0, i_13_371_1401_0, i_13_371_1402_0, i_13_371_1428_0,
    i_13_371_1456_0, i_13_371_1469_0, i_13_371_1599_0, i_13_371_1600_0,
    i_13_371_1644_0, i_13_371_1649_0, i_13_371_1720_0, i_13_371_1722_0,
    i_13_371_1726_0, i_13_371_1777_0, i_13_371_1780_0, i_13_371_1807_0,
    i_13_371_1914_0, i_13_371_1923_0, i_13_371_1939_0, i_13_371_1945_0,
    i_13_371_1946_0, i_13_371_1947_0, i_13_371_1995_0, i_13_371_2026_0,
    i_13_371_2054_0, i_13_371_2107_0, i_13_371_2193_0, i_13_371_2197_0,
    i_13_371_2265_0, i_13_371_2279_0, i_13_371_2302_0, i_13_371_2406_0,
    i_13_371_2472_0, i_13_371_2548_0, i_13_371_2549_0, i_13_371_2568_0,
    i_13_371_2697_0, i_13_371_2742_0, i_13_371_2747_0, i_13_371_2755_0,
    i_13_371_2786_0, i_13_371_2884_0, i_13_371_2886_0, i_13_371_2887_0,
    i_13_371_2899_0, i_13_371_2901_0, i_13_371_2919_0, i_13_371_2940_0,
    i_13_371_2954_0, i_13_371_3030_0, i_13_371_3130_0, i_13_371_3291_0,
    i_13_371_3292_0, i_13_371_3367_0, i_13_371_3368_0, i_13_371_3399_0,
    i_13_371_3459_0, i_13_371_3525_0, i_13_371_3534_0, i_13_371_3570_0,
    i_13_371_3592_0, i_13_371_3593_0, i_13_371_3594_0, i_13_371_3595_0,
    i_13_371_3759_0, i_13_371_3785_0, i_13_371_3787_0, i_13_371_3822_0,
    i_13_371_3908_0, i_13_371_3927_0, i_13_371_3992_0, i_13_371_4037_0,
    i_13_371_4231_0, i_13_371_4305_0, i_13_371_4308_0, i_13_371_4317_0,
    i_13_371_4434_0, i_13_371_4448_0, i_13_371_4449_0, i_13_371_4450_0,
    o_13_371_0_0  );
  input  i_13_371_69_0, i_13_371_70_0, i_13_371_94_0, i_13_371_258_0,
    i_13_371_372_0, i_13_371_373_0, i_13_371_645_0, i_13_371_673_0,
    i_13_371_686_0, i_13_371_797_0, i_13_371_820_0, i_13_371_921_0,
    i_13_371_1065_0, i_13_371_1103_0, i_13_371_1104_0, i_13_371_1148_0,
    i_13_371_1274_0, i_13_371_1275_0, i_13_371_1276_0, i_13_371_1297_0,
    i_13_371_1317_0, i_13_371_1401_0, i_13_371_1402_0, i_13_371_1428_0,
    i_13_371_1456_0, i_13_371_1469_0, i_13_371_1599_0, i_13_371_1600_0,
    i_13_371_1644_0, i_13_371_1649_0, i_13_371_1720_0, i_13_371_1722_0,
    i_13_371_1726_0, i_13_371_1777_0, i_13_371_1780_0, i_13_371_1807_0,
    i_13_371_1914_0, i_13_371_1923_0, i_13_371_1939_0, i_13_371_1945_0,
    i_13_371_1946_0, i_13_371_1947_0, i_13_371_1995_0, i_13_371_2026_0,
    i_13_371_2054_0, i_13_371_2107_0, i_13_371_2193_0, i_13_371_2197_0,
    i_13_371_2265_0, i_13_371_2279_0, i_13_371_2302_0, i_13_371_2406_0,
    i_13_371_2472_0, i_13_371_2548_0, i_13_371_2549_0, i_13_371_2568_0,
    i_13_371_2697_0, i_13_371_2742_0, i_13_371_2747_0, i_13_371_2755_0,
    i_13_371_2786_0, i_13_371_2884_0, i_13_371_2886_0, i_13_371_2887_0,
    i_13_371_2899_0, i_13_371_2901_0, i_13_371_2919_0, i_13_371_2940_0,
    i_13_371_2954_0, i_13_371_3030_0, i_13_371_3130_0, i_13_371_3291_0,
    i_13_371_3292_0, i_13_371_3367_0, i_13_371_3368_0, i_13_371_3399_0,
    i_13_371_3459_0, i_13_371_3525_0, i_13_371_3534_0, i_13_371_3570_0,
    i_13_371_3592_0, i_13_371_3593_0, i_13_371_3594_0, i_13_371_3595_0,
    i_13_371_3759_0, i_13_371_3785_0, i_13_371_3787_0, i_13_371_3822_0,
    i_13_371_3908_0, i_13_371_3927_0, i_13_371_3992_0, i_13_371_4037_0,
    i_13_371_4231_0, i_13_371_4305_0, i_13_371_4308_0, i_13_371_4317_0,
    i_13_371_4434_0, i_13_371_4448_0, i_13_371_4449_0, i_13_371_4450_0;
  output o_13_371_0_0;
  assign o_13_371_0_0 = ~(~i_13_371_1780_0 | (~i_13_371_3822_0 & ~i_13_371_4450_0) | (~i_13_371_1644_0 & ~i_13_371_2742_0));
endmodule



// Benchmark "kernel_13_372" written by ABC on Sun Jul 19 10:50:34 2020

module kernel_13_372 ( 
    i_13_372_118_0, i_13_372_125_0, i_13_372_179_0, i_13_372_191_0,
    i_13_372_195_0, i_13_372_196_0, i_13_372_197_0, i_13_372_303_0,
    i_13_372_575_0, i_13_372_614_0, i_13_372_664_0, i_13_372_712_0,
    i_13_372_719_0, i_13_372_772_0, i_13_372_800_0, i_13_372_862_0,
    i_13_372_863_0, i_13_372_932_0, i_13_372_943_0, i_13_372_952_0,
    i_13_372_953_0, i_13_372_1073_0, i_13_372_1079_0, i_13_372_1226_0,
    i_13_372_1228_0, i_13_372_1231_0, i_13_372_1232_0, i_13_372_1252_0,
    i_13_372_1253_0, i_13_372_1259_0, i_13_372_1285_0, i_13_372_1315_0,
    i_13_372_1318_0, i_13_372_1321_0, i_13_372_1322_0, i_13_372_1410_0,
    i_13_372_1411_0, i_13_372_1491_0, i_13_372_1492_0, i_13_372_1493_0,
    i_13_372_1502_0, i_13_372_1538_0, i_13_372_1550_0, i_13_372_1556_0,
    i_13_372_1573_0, i_13_372_1739_0, i_13_372_1741_0, i_13_372_1781_0,
    i_13_372_1919_0, i_13_372_1960_0, i_13_372_1961_0, i_13_372_2002_0,
    i_13_372_2015_0, i_13_372_2059_0, i_13_372_2195_0, i_13_372_2207_0,
    i_13_372_2242_0, i_13_372_2265_0, i_13_372_2300_0, i_13_372_2314_0,
    i_13_372_2359_0, i_13_372_2423_0, i_13_372_2536_0, i_13_372_2545_0,
    i_13_372_2573_0, i_13_372_2617_0, i_13_372_2618_0, i_13_372_2712_0,
    i_13_372_2918_0, i_13_372_3049_0, i_13_372_3050_0, i_13_372_3117_0,
    i_13_372_3170_0, i_13_372_3212_0, i_13_372_3220_0, i_13_372_3221_0,
    i_13_372_3290_0, i_13_372_3346_0, i_13_372_3391_0, i_13_372_3471_0,
    i_13_372_3475_0, i_13_372_3491_0, i_13_372_3535_0, i_13_372_3536_0,
    i_13_372_3560_0, i_13_372_3565_0, i_13_372_3575_0, i_13_372_3781_0,
    i_13_372_3782_0, i_13_372_3859_0, i_13_372_3878_0, i_13_372_4012_0,
    i_13_372_4013_0, i_13_372_4091_0, i_13_372_4094_0, i_13_372_4252_0,
    i_13_372_4372_0, i_13_372_4381_0, i_13_372_4520_0, i_13_372_4559_0,
    o_13_372_0_0  );
  input  i_13_372_118_0, i_13_372_125_0, i_13_372_179_0, i_13_372_191_0,
    i_13_372_195_0, i_13_372_196_0, i_13_372_197_0, i_13_372_303_0,
    i_13_372_575_0, i_13_372_614_0, i_13_372_664_0, i_13_372_712_0,
    i_13_372_719_0, i_13_372_772_0, i_13_372_800_0, i_13_372_862_0,
    i_13_372_863_0, i_13_372_932_0, i_13_372_943_0, i_13_372_952_0,
    i_13_372_953_0, i_13_372_1073_0, i_13_372_1079_0, i_13_372_1226_0,
    i_13_372_1228_0, i_13_372_1231_0, i_13_372_1232_0, i_13_372_1252_0,
    i_13_372_1253_0, i_13_372_1259_0, i_13_372_1285_0, i_13_372_1315_0,
    i_13_372_1318_0, i_13_372_1321_0, i_13_372_1322_0, i_13_372_1410_0,
    i_13_372_1411_0, i_13_372_1491_0, i_13_372_1492_0, i_13_372_1493_0,
    i_13_372_1502_0, i_13_372_1538_0, i_13_372_1550_0, i_13_372_1556_0,
    i_13_372_1573_0, i_13_372_1739_0, i_13_372_1741_0, i_13_372_1781_0,
    i_13_372_1919_0, i_13_372_1960_0, i_13_372_1961_0, i_13_372_2002_0,
    i_13_372_2015_0, i_13_372_2059_0, i_13_372_2195_0, i_13_372_2207_0,
    i_13_372_2242_0, i_13_372_2265_0, i_13_372_2300_0, i_13_372_2314_0,
    i_13_372_2359_0, i_13_372_2423_0, i_13_372_2536_0, i_13_372_2545_0,
    i_13_372_2573_0, i_13_372_2617_0, i_13_372_2618_0, i_13_372_2712_0,
    i_13_372_2918_0, i_13_372_3049_0, i_13_372_3050_0, i_13_372_3117_0,
    i_13_372_3170_0, i_13_372_3212_0, i_13_372_3220_0, i_13_372_3221_0,
    i_13_372_3290_0, i_13_372_3346_0, i_13_372_3391_0, i_13_372_3471_0,
    i_13_372_3475_0, i_13_372_3491_0, i_13_372_3535_0, i_13_372_3536_0,
    i_13_372_3560_0, i_13_372_3565_0, i_13_372_3575_0, i_13_372_3781_0,
    i_13_372_3782_0, i_13_372_3859_0, i_13_372_3878_0, i_13_372_4012_0,
    i_13_372_4013_0, i_13_372_4091_0, i_13_372_4094_0, i_13_372_4252_0,
    i_13_372_4372_0, i_13_372_4381_0, i_13_372_4520_0, i_13_372_4559_0;
  output o_13_372_0_0;
  assign o_13_372_0_0 = ~((~i_13_372_2618_0 & ~i_13_372_4012_0) | (i_13_372_3220_0 & ~i_13_372_3290_0) | (i_13_372_2002_0 & i_13_372_2712_0) | (~i_13_372_863_0 & ~i_13_372_1493_0 & ~i_13_372_4372_0) | (i_13_372_3346_0 & ~i_13_372_3535_0 & ~i_13_372_3859_0));
endmodule



// Benchmark "kernel_13_373" written by ABC on Sun Jul 19 10:50:35 2020

module kernel_13_373 ( 
    i_13_373_40_0, i_13_373_43_0, i_13_373_112_0, i_13_373_113_0,
    i_13_373_141_0, i_13_373_142_0, i_13_373_193_0, i_13_373_241_0,
    i_13_373_251_0, i_13_373_380_0, i_13_373_389_0, i_13_373_562_0,
    i_13_373_581_0, i_13_373_583_0, i_13_373_619_0, i_13_373_776_0,
    i_13_373_819_0, i_13_373_843_0, i_13_373_1083_0, i_13_373_1084_0,
    i_13_373_1087_0, i_13_373_1098_0, i_13_373_1212_0, i_13_373_1219_0,
    i_13_373_1273_0, i_13_373_1318_0, i_13_373_1427_0, i_13_373_1429_0,
    i_13_373_1444_0, i_13_373_1473_0, i_13_373_1474_0, i_13_373_1552_0,
    i_13_373_1572_0, i_13_373_1602_0, i_13_373_1624_0, i_13_373_1636_0,
    i_13_373_1681_0, i_13_373_1750_0, i_13_373_1800_0, i_13_373_1804_0,
    i_13_373_1817_0, i_13_373_1840_0, i_13_373_1924_0, i_13_373_1933_0,
    i_13_373_1943_0, i_13_373_1960_0, i_13_373_1996_0, i_13_373_2005_0,
    i_13_373_2006_0, i_13_373_2124_0, i_13_373_2187_0, i_13_373_2196_0,
    i_13_373_2276_0, i_13_373_2428_0, i_13_373_2434_0, i_13_373_2437_0,
    i_13_373_2455_0, i_13_373_2646_0, i_13_373_2713_0, i_13_373_2716_0,
    i_13_373_2717_0, i_13_373_2726_0, i_13_373_2858_0, i_13_373_2958_0,
    i_13_373_3010_0, i_13_373_3038_0, i_13_373_3064_0, i_13_373_3066_0,
    i_13_373_3067_0, i_13_373_3146_0, i_13_373_3227_0, i_13_373_3258_0,
    i_13_373_3326_0, i_13_373_3373_0, i_13_373_3374_0, i_13_373_3440_0,
    i_13_373_3442_0, i_13_373_3526_0, i_13_373_3537_0, i_13_373_3541_0,
    i_13_373_3559_0, i_13_373_3564_0, i_13_373_3573_0, i_13_373_3649_0,
    i_13_373_3653_0, i_13_373_3685_0, i_13_373_3686_0, i_13_373_3687_0,
    i_13_373_3688_0, i_13_373_3689_0, i_13_373_3726_0, i_13_373_3780_0,
    i_13_373_3852_0, i_13_373_3856_0, i_13_373_4021_0, i_13_373_4057_0,
    i_13_373_4093_0, i_13_373_4230_0, i_13_373_4257_0, i_13_373_4400_0,
    o_13_373_0_0  );
  input  i_13_373_40_0, i_13_373_43_0, i_13_373_112_0, i_13_373_113_0,
    i_13_373_141_0, i_13_373_142_0, i_13_373_193_0, i_13_373_241_0,
    i_13_373_251_0, i_13_373_380_0, i_13_373_389_0, i_13_373_562_0,
    i_13_373_581_0, i_13_373_583_0, i_13_373_619_0, i_13_373_776_0,
    i_13_373_819_0, i_13_373_843_0, i_13_373_1083_0, i_13_373_1084_0,
    i_13_373_1087_0, i_13_373_1098_0, i_13_373_1212_0, i_13_373_1219_0,
    i_13_373_1273_0, i_13_373_1318_0, i_13_373_1427_0, i_13_373_1429_0,
    i_13_373_1444_0, i_13_373_1473_0, i_13_373_1474_0, i_13_373_1552_0,
    i_13_373_1572_0, i_13_373_1602_0, i_13_373_1624_0, i_13_373_1636_0,
    i_13_373_1681_0, i_13_373_1750_0, i_13_373_1800_0, i_13_373_1804_0,
    i_13_373_1817_0, i_13_373_1840_0, i_13_373_1924_0, i_13_373_1933_0,
    i_13_373_1943_0, i_13_373_1960_0, i_13_373_1996_0, i_13_373_2005_0,
    i_13_373_2006_0, i_13_373_2124_0, i_13_373_2187_0, i_13_373_2196_0,
    i_13_373_2276_0, i_13_373_2428_0, i_13_373_2434_0, i_13_373_2437_0,
    i_13_373_2455_0, i_13_373_2646_0, i_13_373_2713_0, i_13_373_2716_0,
    i_13_373_2717_0, i_13_373_2726_0, i_13_373_2858_0, i_13_373_2958_0,
    i_13_373_3010_0, i_13_373_3038_0, i_13_373_3064_0, i_13_373_3066_0,
    i_13_373_3067_0, i_13_373_3146_0, i_13_373_3227_0, i_13_373_3258_0,
    i_13_373_3326_0, i_13_373_3373_0, i_13_373_3374_0, i_13_373_3440_0,
    i_13_373_3442_0, i_13_373_3526_0, i_13_373_3537_0, i_13_373_3541_0,
    i_13_373_3559_0, i_13_373_3564_0, i_13_373_3573_0, i_13_373_3649_0,
    i_13_373_3653_0, i_13_373_3685_0, i_13_373_3686_0, i_13_373_3687_0,
    i_13_373_3688_0, i_13_373_3689_0, i_13_373_3726_0, i_13_373_3780_0,
    i_13_373_3852_0, i_13_373_3856_0, i_13_373_4021_0, i_13_373_4057_0,
    i_13_373_4093_0, i_13_373_4230_0, i_13_373_4257_0, i_13_373_4400_0;
  output o_13_373_0_0;
  assign o_13_373_0_0 = ~((~i_13_373_2716_0 & (~i_13_373_1084_0 | (~i_13_373_562_0 & ~i_13_373_1083_0 & ~i_13_373_3653_0))) | (~i_13_373_241_0 & ~i_13_373_1572_0 & ~i_13_373_3067_0) | (~i_13_373_3685_0 & ~i_13_373_4093_0 & ~i_13_373_4400_0));
endmodule



// Benchmark "kernel_13_374" written by ABC on Sun Jul 19 10:50:36 2020

module kernel_13_374 ( 
    i_13_374_30_0, i_13_374_63_0, i_13_374_64_0, i_13_374_79_0,
    i_13_374_99_0, i_13_374_112_0, i_13_374_162_0, i_13_374_199_0,
    i_13_374_225_0, i_13_374_272_0, i_13_374_357_0, i_13_374_370_0,
    i_13_374_396_0, i_13_374_405_0, i_13_374_428_0, i_13_374_445_0,
    i_13_374_468_0, i_13_374_470_0, i_13_374_489_0, i_13_374_568_0,
    i_13_374_622_0, i_13_374_684_0, i_13_374_695_0, i_13_374_810_0,
    i_13_374_956_0, i_13_374_1017_0, i_13_374_1098_0, i_13_374_1263_0,
    i_13_374_1269_0, i_13_374_1296_0, i_13_374_1363_0, i_13_374_1424_0,
    i_13_374_1432_0, i_13_374_1478_0, i_13_374_1503_0, i_13_374_1504_0,
    i_13_374_1593_0, i_13_374_1638_0, i_13_374_1642_0, i_13_374_1643_0,
    i_13_374_1688_0, i_13_374_1719_0, i_13_374_1720_0, i_13_374_1791_0,
    i_13_374_1792_0, i_13_374_1828_0, i_13_374_1881_0, i_13_374_1927_0,
    i_13_374_2015_0, i_13_374_2100_0, i_13_374_2103_0, i_13_374_2111_0,
    i_13_374_2179_0, i_13_374_2235_0, i_13_374_2238_0, i_13_374_2246_0,
    i_13_374_2376_0, i_13_374_2377_0, i_13_374_2378_0, i_13_374_2444_0,
    i_13_374_2558_0, i_13_374_2720_0, i_13_374_2749_0, i_13_374_2917_0,
    i_13_374_2934_0, i_13_374_2935_0, i_13_374_3171_0, i_13_374_3241_0,
    i_13_374_3262_0, i_13_374_3305_0, i_13_374_3396_0, i_13_374_3450_0,
    i_13_374_3451_0, i_13_374_3479_0, i_13_374_3566_0, i_13_374_3648_0,
    i_13_374_3762_0, i_13_374_3763_0, i_13_374_3790_0, i_13_374_3859_0,
    i_13_374_3865_0, i_13_374_3893_0, i_13_374_3987_0, i_13_374_3988_0,
    i_13_374_4050_0, i_13_374_4051_0, i_13_374_4078_0, i_13_374_4159_0,
    i_13_374_4212_0, i_13_374_4215_0, i_13_374_4234_0, i_13_374_4303_0,
    i_13_374_4312_0, i_13_374_4369_0, i_13_374_4375_0, i_13_374_4379_0,
    i_13_374_4410_0, i_13_374_4432_0, i_13_374_4512_0, i_13_374_4582_0,
    o_13_374_0_0  );
  input  i_13_374_30_0, i_13_374_63_0, i_13_374_64_0, i_13_374_79_0,
    i_13_374_99_0, i_13_374_112_0, i_13_374_162_0, i_13_374_199_0,
    i_13_374_225_0, i_13_374_272_0, i_13_374_357_0, i_13_374_370_0,
    i_13_374_396_0, i_13_374_405_0, i_13_374_428_0, i_13_374_445_0,
    i_13_374_468_0, i_13_374_470_0, i_13_374_489_0, i_13_374_568_0,
    i_13_374_622_0, i_13_374_684_0, i_13_374_695_0, i_13_374_810_0,
    i_13_374_956_0, i_13_374_1017_0, i_13_374_1098_0, i_13_374_1263_0,
    i_13_374_1269_0, i_13_374_1296_0, i_13_374_1363_0, i_13_374_1424_0,
    i_13_374_1432_0, i_13_374_1478_0, i_13_374_1503_0, i_13_374_1504_0,
    i_13_374_1593_0, i_13_374_1638_0, i_13_374_1642_0, i_13_374_1643_0,
    i_13_374_1688_0, i_13_374_1719_0, i_13_374_1720_0, i_13_374_1791_0,
    i_13_374_1792_0, i_13_374_1828_0, i_13_374_1881_0, i_13_374_1927_0,
    i_13_374_2015_0, i_13_374_2100_0, i_13_374_2103_0, i_13_374_2111_0,
    i_13_374_2179_0, i_13_374_2235_0, i_13_374_2238_0, i_13_374_2246_0,
    i_13_374_2376_0, i_13_374_2377_0, i_13_374_2378_0, i_13_374_2444_0,
    i_13_374_2558_0, i_13_374_2720_0, i_13_374_2749_0, i_13_374_2917_0,
    i_13_374_2934_0, i_13_374_2935_0, i_13_374_3171_0, i_13_374_3241_0,
    i_13_374_3262_0, i_13_374_3305_0, i_13_374_3396_0, i_13_374_3450_0,
    i_13_374_3451_0, i_13_374_3479_0, i_13_374_3566_0, i_13_374_3648_0,
    i_13_374_3762_0, i_13_374_3763_0, i_13_374_3790_0, i_13_374_3859_0,
    i_13_374_3865_0, i_13_374_3893_0, i_13_374_3987_0, i_13_374_3988_0,
    i_13_374_4050_0, i_13_374_4051_0, i_13_374_4078_0, i_13_374_4159_0,
    i_13_374_4212_0, i_13_374_4215_0, i_13_374_4234_0, i_13_374_4303_0,
    i_13_374_4312_0, i_13_374_4369_0, i_13_374_4375_0, i_13_374_4379_0,
    i_13_374_4410_0, i_13_374_4432_0, i_13_374_4512_0, i_13_374_4582_0;
  output o_13_374_0_0;
  assign o_13_374_0_0 = ~((i_13_374_3865_0 & i_13_374_4379_0) | (~i_13_374_64_0 & ~i_13_374_1791_0 & ~i_13_374_1881_0) | (~i_13_374_1424_0 & ~i_13_374_1593_0 & ~i_13_374_2246_0 & ~i_13_374_4050_0));
endmodule



// Benchmark "kernel_13_375" written by ABC on Sun Jul 19 10:50:37 2020

module kernel_13_375 ( 
    i_13_375_46_0, i_13_375_49_0, i_13_375_71_0, i_13_375_136_0,
    i_13_375_190_0, i_13_375_316_0, i_13_375_338_0, i_13_375_362_0,
    i_13_375_373_0, i_13_375_412_0, i_13_375_415_0, i_13_375_550_0,
    i_13_375_568_0, i_13_375_626_0, i_13_375_651_0, i_13_375_662_0,
    i_13_375_811_0, i_13_375_836_0, i_13_375_851_0, i_13_375_934_0,
    i_13_375_937_0, i_13_375_939_0, i_13_375_940_0, i_13_375_1018_0,
    i_13_375_1022_0, i_13_375_1072_0, i_13_375_1101_0, i_13_375_1102_0,
    i_13_375_1104_0, i_13_375_1105_0, i_13_375_1119_0, i_13_375_1120_0,
    i_13_375_1230_0, i_13_375_1391_0, i_13_375_1407_0, i_13_375_1508_0,
    i_13_375_1544_0, i_13_375_1549_0, i_13_375_1603_0, i_13_375_1661_0,
    i_13_375_1668_0, i_13_375_1736_0, i_13_375_1768_0, i_13_375_1796_0,
    i_13_375_1798_0, i_13_375_1799_0, i_13_375_1858_0, i_13_375_2020_0,
    i_13_375_2021_0, i_13_375_2145_0, i_13_375_2301_0, i_13_375_2381_0,
    i_13_375_2461_0, i_13_375_2469_0, i_13_375_2470_0, i_13_375_2471_0,
    i_13_375_2473_0, i_13_375_2474_0, i_13_375_2677_0, i_13_375_2857_0,
    i_13_375_2858_0, i_13_375_2907_0, i_13_375_2966_0, i_13_375_2969_0,
    i_13_375_2986_0, i_13_375_3029_0, i_13_375_3031_0, i_13_375_3032_0,
    i_13_375_3077_0, i_13_375_3117_0, i_13_375_3128_0, i_13_375_3204_0,
    i_13_375_3210_0, i_13_375_3261_0, i_13_375_3265_0, i_13_375_3272_0,
    i_13_375_3380_0, i_13_375_3404_0, i_13_375_3457_0, i_13_375_3476_0,
    i_13_375_3482_0, i_13_375_3484_0, i_13_375_3505_0, i_13_375_3548_0,
    i_13_375_3568_0, i_13_375_3666_0, i_13_375_3823_0, i_13_375_3898_0,
    i_13_375_3899_0, i_13_375_3901_0, i_13_375_3964_0, i_13_375_4018_0,
    i_13_375_4069_0, i_13_375_4090_0, i_13_375_4116_0, i_13_375_4204_0,
    i_13_375_4298_0, i_13_375_4505_0, i_13_375_4604_0, i_13_375_4607_0,
    o_13_375_0_0  );
  input  i_13_375_46_0, i_13_375_49_0, i_13_375_71_0, i_13_375_136_0,
    i_13_375_190_0, i_13_375_316_0, i_13_375_338_0, i_13_375_362_0,
    i_13_375_373_0, i_13_375_412_0, i_13_375_415_0, i_13_375_550_0,
    i_13_375_568_0, i_13_375_626_0, i_13_375_651_0, i_13_375_662_0,
    i_13_375_811_0, i_13_375_836_0, i_13_375_851_0, i_13_375_934_0,
    i_13_375_937_0, i_13_375_939_0, i_13_375_940_0, i_13_375_1018_0,
    i_13_375_1022_0, i_13_375_1072_0, i_13_375_1101_0, i_13_375_1102_0,
    i_13_375_1104_0, i_13_375_1105_0, i_13_375_1119_0, i_13_375_1120_0,
    i_13_375_1230_0, i_13_375_1391_0, i_13_375_1407_0, i_13_375_1508_0,
    i_13_375_1544_0, i_13_375_1549_0, i_13_375_1603_0, i_13_375_1661_0,
    i_13_375_1668_0, i_13_375_1736_0, i_13_375_1768_0, i_13_375_1796_0,
    i_13_375_1798_0, i_13_375_1799_0, i_13_375_1858_0, i_13_375_2020_0,
    i_13_375_2021_0, i_13_375_2145_0, i_13_375_2301_0, i_13_375_2381_0,
    i_13_375_2461_0, i_13_375_2469_0, i_13_375_2470_0, i_13_375_2471_0,
    i_13_375_2473_0, i_13_375_2474_0, i_13_375_2677_0, i_13_375_2857_0,
    i_13_375_2858_0, i_13_375_2907_0, i_13_375_2966_0, i_13_375_2969_0,
    i_13_375_2986_0, i_13_375_3029_0, i_13_375_3031_0, i_13_375_3032_0,
    i_13_375_3077_0, i_13_375_3117_0, i_13_375_3128_0, i_13_375_3204_0,
    i_13_375_3210_0, i_13_375_3261_0, i_13_375_3265_0, i_13_375_3272_0,
    i_13_375_3380_0, i_13_375_3404_0, i_13_375_3457_0, i_13_375_3476_0,
    i_13_375_3482_0, i_13_375_3484_0, i_13_375_3505_0, i_13_375_3548_0,
    i_13_375_3568_0, i_13_375_3666_0, i_13_375_3823_0, i_13_375_3898_0,
    i_13_375_3899_0, i_13_375_3901_0, i_13_375_3964_0, i_13_375_4018_0,
    i_13_375_4069_0, i_13_375_4090_0, i_13_375_4116_0, i_13_375_4204_0,
    i_13_375_4298_0, i_13_375_4505_0, i_13_375_4604_0, i_13_375_4607_0;
  output o_13_375_0_0;
  assign o_13_375_0_0 = 0;
endmodule



// Benchmark "kernel_13_376" written by ABC on Sun Jul 19 10:50:37 2020

module kernel_13_376 ( 
    i_13_376_49_0, i_13_376_67_0, i_13_376_70_0, i_13_376_178_0,
    i_13_376_259_0, i_13_376_276_0, i_13_376_277_0, i_13_376_310_0,
    i_13_376_355_0, i_13_376_476_0, i_13_376_520_0, i_13_376_535_0,
    i_13_376_619_0, i_13_376_642_0, i_13_376_651_0, i_13_376_673_0,
    i_13_376_745_0, i_13_376_922_0, i_13_376_934_0, i_13_376_1024_0,
    i_13_376_1104_0, i_13_376_1105_0, i_13_376_1132_0, i_13_376_1276_0,
    i_13_376_1330_0, i_13_376_1401_0, i_13_376_1402_0, i_13_376_1481_0,
    i_13_376_1510_0, i_13_376_1564_0, i_13_376_1573_0, i_13_376_1574_0,
    i_13_376_1597_0, i_13_376_1641_0, i_13_376_1653_0, i_13_376_1659_0,
    i_13_376_1723_0, i_13_376_1735_0, i_13_376_1779_0, i_13_376_1835_0,
    i_13_376_1914_0, i_13_376_1923_0, i_13_376_1924_0, i_13_376_1932_0,
    i_13_376_1947_0, i_13_376_2019_0, i_13_376_2022_0, i_13_376_2028_0,
    i_13_376_2029_0, i_13_376_2185_0, i_13_376_2196_0, i_13_376_2199_0,
    i_13_376_2302_0, i_13_376_2436_0, i_13_376_2454_0, i_13_376_2469_0,
    i_13_376_2473_0, i_13_376_2518_0, i_13_376_2677_0, i_13_376_2697_0,
    i_13_376_2742_0, i_13_376_2743_0, i_13_376_2769_0, i_13_376_2770_0,
    i_13_376_2850_0, i_13_376_2923_0, i_13_376_2940_0, i_13_376_2968_0,
    i_13_376_3030_0, i_13_376_3031_0, i_13_376_3077_0, i_13_376_3110_0,
    i_13_376_3121_0, i_13_376_3130_0, i_13_376_3246_0, i_13_376_3291_0,
    i_13_376_3315_0, i_13_376_3381_0, i_13_376_3418_0, i_13_376_3453_0,
    i_13_376_3525_0, i_13_376_3577_0, i_13_376_3595_0, i_13_376_3625_0,
    i_13_376_3785_0, i_13_376_3786_0, i_13_376_3787_0, i_13_376_3819_0,
    i_13_376_3822_0, i_13_376_3901_0, i_13_376_3930_0, i_13_376_4029_0,
    i_13_376_4093_0, i_13_376_4323_0, i_13_376_4324_0, i_13_376_4325_0,
    i_13_376_4390_0, i_13_376_4434_0, i_13_376_4516_0, i_13_376_4606_0,
    o_13_376_0_0  );
  input  i_13_376_49_0, i_13_376_67_0, i_13_376_70_0, i_13_376_178_0,
    i_13_376_259_0, i_13_376_276_0, i_13_376_277_0, i_13_376_310_0,
    i_13_376_355_0, i_13_376_476_0, i_13_376_520_0, i_13_376_535_0,
    i_13_376_619_0, i_13_376_642_0, i_13_376_651_0, i_13_376_673_0,
    i_13_376_745_0, i_13_376_922_0, i_13_376_934_0, i_13_376_1024_0,
    i_13_376_1104_0, i_13_376_1105_0, i_13_376_1132_0, i_13_376_1276_0,
    i_13_376_1330_0, i_13_376_1401_0, i_13_376_1402_0, i_13_376_1481_0,
    i_13_376_1510_0, i_13_376_1564_0, i_13_376_1573_0, i_13_376_1574_0,
    i_13_376_1597_0, i_13_376_1641_0, i_13_376_1653_0, i_13_376_1659_0,
    i_13_376_1723_0, i_13_376_1735_0, i_13_376_1779_0, i_13_376_1835_0,
    i_13_376_1914_0, i_13_376_1923_0, i_13_376_1924_0, i_13_376_1932_0,
    i_13_376_1947_0, i_13_376_2019_0, i_13_376_2022_0, i_13_376_2028_0,
    i_13_376_2029_0, i_13_376_2185_0, i_13_376_2196_0, i_13_376_2199_0,
    i_13_376_2302_0, i_13_376_2436_0, i_13_376_2454_0, i_13_376_2469_0,
    i_13_376_2473_0, i_13_376_2518_0, i_13_376_2677_0, i_13_376_2697_0,
    i_13_376_2742_0, i_13_376_2743_0, i_13_376_2769_0, i_13_376_2770_0,
    i_13_376_2850_0, i_13_376_2923_0, i_13_376_2940_0, i_13_376_2968_0,
    i_13_376_3030_0, i_13_376_3031_0, i_13_376_3077_0, i_13_376_3110_0,
    i_13_376_3121_0, i_13_376_3130_0, i_13_376_3246_0, i_13_376_3291_0,
    i_13_376_3315_0, i_13_376_3381_0, i_13_376_3418_0, i_13_376_3453_0,
    i_13_376_3525_0, i_13_376_3577_0, i_13_376_3595_0, i_13_376_3625_0,
    i_13_376_3785_0, i_13_376_3786_0, i_13_376_3787_0, i_13_376_3819_0,
    i_13_376_3822_0, i_13_376_3901_0, i_13_376_3930_0, i_13_376_4029_0,
    i_13_376_4093_0, i_13_376_4323_0, i_13_376_4324_0, i_13_376_4325_0,
    i_13_376_4390_0, i_13_376_4434_0, i_13_376_4516_0, i_13_376_4606_0;
  output o_13_376_0_0;
  assign o_13_376_0_0 = ~((~i_13_376_4434_0 & ((~i_13_376_520_0 & ~i_13_376_1401_0 & ~i_13_376_2185_0 & ~i_13_376_2742_0) | (~i_13_376_1779_0 & i_13_376_2850_0))) | (~i_13_376_49_0 & ~i_13_376_2022_0 & ~i_13_376_3453_0) | (~i_13_376_1573_0 & ~i_13_376_2850_0 & ~i_13_376_3246_0 & ~i_13_376_4324_0));
endmodule



// Benchmark "kernel_13_377" written by ABC on Sun Jul 19 10:50:38 2020

module kernel_13_377 ( 
    i_13_377_98_0, i_13_377_107_0, i_13_377_113_0, i_13_377_140_0,
    i_13_377_251_0, i_13_377_262_0, i_13_377_368_0, i_13_377_370_0,
    i_13_377_538_0, i_13_377_554_0, i_13_377_562_0, i_13_377_608_0,
    i_13_377_620_0, i_13_377_647_0, i_13_377_655_0, i_13_377_661_0,
    i_13_377_671_0, i_13_377_680_0, i_13_377_845_0, i_13_377_949_0,
    i_13_377_1070_0, i_13_377_1087_0, i_13_377_1145_0, i_13_377_1148_0,
    i_13_377_1219_0, i_13_377_1220_0, i_13_377_1264_0, i_13_377_1318_0,
    i_13_377_1348_0, i_13_377_1474_0, i_13_377_1519_0, i_13_377_1520_0,
    i_13_377_1574_0, i_13_377_1624_0, i_13_377_1727_0, i_13_377_1742_0,
    i_13_377_1745_0, i_13_377_1789_0, i_13_377_1840_0, i_13_377_1841_0,
    i_13_377_2024_0, i_13_377_2137_0, i_13_377_2173_0, i_13_377_2284_0,
    i_13_377_2285_0, i_13_377_2348_0, i_13_377_2380_0, i_13_377_2417_0,
    i_13_377_2435_0, i_13_377_2437_0, i_13_377_2438_0, i_13_377_2501_0,
    i_13_377_2510_0, i_13_377_2599_0, i_13_377_2680_0, i_13_377_2716_0,
    i_13_377_2717_0, i_13_377_2749_0, i_13_377_2879_0, i_13_377_2906_0,
    i_13_377_2987_0, i_13_377_3047_0, i_13_377_3053_0, i_13_377_3059_0,
    i_13_377_3067_0, i_13_377_3100_0, i_13_377_3130_0, i_13_377_3131_0,
    i_13_377_3148_0, i_13_377_3149_0, i_13_377_3166_0, i_13_377_3167_0,
    i_13_377_3329_0, i_13_377_3343_0, i_13_377_3347_0, i_13_377_3373_0,
    i_13_377_3455_0, i_13_377_3464_0, i_13_377_3478_0, i_13_377_3527_0,
    i_13_377_3623_0, i_13_377_3632_0, i_13_377_4021_0, i_13_377_4049_0,
    i_13_377_4100_0, i_13_377_4120_0, i_13_377_4121_0, i_13_377_4192_0,
    i_13_377_4262_0, i_13_377_4264_0, i_13_377_4321_0, i_13_377_4328_0,
    i_13_377_4343_0, i_13_377_4354_0, i_13_377_4418_0, i_13_377_4460_0,
    i_13_377_4463_0, i_13_377_4543_0, i_13_377_4544_0, i_13_377_4604_0,
    o_13_377_0_0  );
  input  i_13_377_98_0, i_13_377_107_0, i_13_377_113_0, i_13_377_140_0,
    i_13_377_251_0, i_13_377_262_0, i_13_377_368_0, i_13_377_370_0,
    i_13_377_538_0, i_13_377_554_0, i_13_377_562_0, i_13_377_608_0,
    i_13_377_620_0, i_13_377_647_0, i_13_377_655_0, i_13_377_661_0,
    i_13_377_671_0, i_13_377_680_0, i_13_377_845_0, i_13_377_949_0,
    i_13_377_1070_0, i_13_377_1087_0, i_13_377_1145_0, i_13_377_1148_0,
    i_13_377_1219_0, i_13_377_1220_0, i_13_377_1264_0, i_13_377_1318_0,
    i_13_377_1348_0, i_13_377_1474_0, i_13_377_1519_0, i_13_377_1520_0,
    i_13_377_1574_0, i_13_377_1624_0, i_13_377_1727_0, i_13_377_1742_0,
    i_13_377_1745_0, i_13_377_1789_0, i_13_377_1840_0, i_13_377_1841_0,
    i_13_377_2024_0, i_13_377_2137_0, i_13_377_2173_0, i_13_377_2284_0,
    i_13_377_2285_0, i_13_377_2348_0, i_13_377_2380_0, i_13_377_2417_0,
    i_13_377_2435_0, i_13_377_2437_0, i_13_377_2438_0, i_13_377_2501_0,
    i_13_377_2510_0, i_13_377_2599_0, i_13_377_2680_0, i_13_377_2716_0,
    i_13_377_2717_0, i_13_377_2749_0, i_13_377_2879_0, i_13_377_2906_0,
    i_13_377_2987_0, i_13_377_3047_0, i_13_377_3053_0, i_13_377_3059_0,
    i_13_377_3067_0, i_13_377_3100_0, i_13_377_3130_0, i_13_377_3131_0,
    i_13_377_3148_0, i_13_377_3149_0, i_13_377_3166_0, i_13_377_3167_0,
    i_13_377_3329_0, i_13_377_3343_0, i_13_377_3347_0, i_13_377_3373_0,
    i_13_377_3455_0, i_13_377_3464_0, i_13_377_3478_0, i_13_377_3527_0,
    i_13_377_3623_0, i_13_377_3632_0, i_13_377_4021_0, i_13_377_4049_0,
    i_13_377_4100_0, i_13_377_4120_0, i_13_377_4121_0, i_13_377_4192_0,
    i_13_377_4262_0, i_13_377_4264_0, i_13_377_4321_0, i_13_377_4328_0,
    i_13_377_4343_0, i_13_377_4354_0, i_13_377_4418_0, i_13_377_4460_0,
    i_13_377_4463_0, i_13_377_4543_0, i_13_377_4544_0, i_13_377_4604_0;
  output o_13_377_0_0;
  assign o_13_377_0_0 = ~(~i_13_377_3149_0 | (~i_13_377_1624_0 & ~i_13_377_1841_0));
endmodule



// Benchmark "kernel_13_378" written by ABC on Sun Jul 19 10:50:39 2020

module kernel_13_378 ( 
    i_13_378_31_0, i_13_378_99_0, i_13_378_139_0, i_13_378_155_0,
    i_13_378_210_0, i_13_378_228_0, i_13_378_229_0, i_13_378_237_0,
    i_13_378_247_0, i_13_378_372_0, i_13_378_513_0, i_13_378_514_0,
    i_13_378_517_0, i_13_378_535_0, i_13_378_569_0, i_13_378_606_0,
    i_13_378_652_0, i_13_378_823_0, i_13_378_840_0, i_13_378_983_0,
    i_13_378_984_0, i_13_378_985_0, i_13_378_1025_0, i_13_378_1063_0,
    i_13_378_1075_0, i_13_378_1112_0, i_13_378_1192_0, i_13_378_1219_0,
    i_13_378_1300_0, i_13_378_1324_0, i_13_378_1326_0, i_13_378_1327_0,
    i_13_378_1447_0, i_13_378_1476_0, i_13_378_1489_0, i_13_378_1525_0,
    i_13_378_1549_0, i_13_378_1569_0, i_13_378_1570_0, i_13_378_1584_0,
    i_13_378_1670_0, i_13_378_1714_0, i_13_378_1723_0, i_13_378_1746_0,
    i_13_378_1831_0, i_13_378_1848_0, i_13_378_1936_0, i_13_378_2002_0,
    i_13_378_2025_0, i_13_378_2029_0, i_13_378_2107_0, i_13_378_2108_0,
    i_13_378_2116_0, i_13_378_2182_0, i_13_378_2233_0, i_13_378_2259_0,
    i_13_378_2377_0, i_13_378_2406_0, i_13_378_2489_0, i_13_378_2557_0,
    i_13_378_2673_0, i_13_378_2677_0, i_13_378_2736_0, i_13_378_2848_0,
    i_13_378_2966_0, i_13_378_3006_0, i_13_378_3007_0, i_13_378_3108_0,
    i_13_378_3109_0, i_13_378_3150_0, i_13_378_3151_0, i_13_378_3209_0,
    i_13_378_3226_0, i_13_378_3313_0, i_13_378_3376_0, i_13_378_3388_0,
    i_13_378_3406_0, i_13_378_3439_0, i_13_378_3460_0, i_13_378_3485_0,
    i_13_378_3546_0, i_13_378_3554_0, i_13_378_3730_0, i_13_378_3763_0,
    i_13_378_3766_0, i_13_378_3817_0, i_13_378_3861_0, i_13_378_3900_0,
    i_13_378_3977_0, i_13_378_4063_0, i_13_378_4123_0, i_13_378_4158_0,
    i_13_378_4452_0, i_13_378_4455_0, i_13_378_4513_0, i_13_378_4554_0,
    i_13_378_4556_0, i_13_378_4564_0, i_13_378_4568_0, i_13_378_4600_0,
    o_13_378_0_0  );
  input  i_13_378_31_0, i_13_378_99_0, i_13_378_139_0, i_13_378_155_0,
    i_13_378_210_0, i_13_378_228_0, i_13_378_229_0, i_13_378_237_0,
    i_13_378_247_0, i_13_378_372_0, i_13_378_513_0, i_13_378_514_0,
    i_13_378_517_0, i_13_378_535_0, i_13_378_569_0, i_13_378_606_0,
    i_13_378_652_0, i_13_378_823_0, i_13_378_840_0, i_13_378_983_0,
    i_13_378_984_0, i_13_378_985_0, i_13_378_1025_0, i_13_378_1063_0,
    i_13_378_1075_0, i_13_378_1112_0, i_13_378_1192_0, i_13_378_1219_0,
    i_13_378_1300_0, i_13_378_1324_0, i_13_378_1326_0, i_13_378_1327_0,
    i_13_378_1447_0, i_13_378_1476_0, i_13_378_1489_0, i_13_378_1525_0,
    i_13_378_1549_0, i_13_378_1569_0, i_13_378_1570_0, i_13_378_1584_0,
    i_13_378_1670_0, i_13_378_1714_0, i_13_378_1723_0, i_13_378_1746_0,
    i_13_378_1831_0, i_13_378_1848_0, i_13_378_1936_0, i_13_378_2002_0,
    i_13_378_2025_0, i_13_378_2029_0, i_13_378_2107_0, i_13_378_2108_0,
    i_13_378_2116_0, i_13_378_2182_0, i_13_378_2233_0, i_13_378_2259_0,
    i_13_378_2377_0, i_13_378_2406_0, i_13_378_2489_0, i_13_378_2557_0,
    i_13_378_2673_0, i_13_378_2677_0, i_13_378_2736_0, i_13_378_2848_0,
    i_13_378_2966_0, i_13_378_3006_0, i_13_378_3007_0, i_13_378_3108_0,
    i_13_378_3109_0, i_13_378_3150_0, i_13_378_3151_0, i_13_378_3209_0,
    i_13_378_3226_0, i_13_378_3313_0, i_13_378_3376_0, i_13_378_3388_0,
    i_13_378_3406_0, i_13_378_3439_0, i_13_378_3460_0, i_13_378_3485_0,
    i_13_378_3546_0, i_13_378_3554_0, i_13_378_3730_0, i_13_378_3763_0,
    i_13_378_3766_0, i_13_378_3817_0, i_13_378_3861_0, i_13_378_3900_0,
    i_13_378_3977_0, i_13_378_4063_0, i_13_378_4123_0, i_13_378_4158_0,
    i_13_378_4452_0, i_13_378_4455_0, i_13_378_4513_0, i_13_378_4554_0,
    i_13_378_4556_0, i_13_378_4564_0, i_13_378_4568_0, i_13_378_4600_0;
  output o_13_378_0_0;
  assign o_13_378_0_0 = ~((~i_13_378_985_0 & (~i_13_378_1831_0 | i_13_378_4452_0)) | (~i_13_378_1326_0 & ((~i_13_378_983_0 & ~i_13_378_2182_0 & ~i_13_378_2673_0) | (~i_13_378_3439_0 & ~i_13_378_3900_0 & ~i_13_378_4554_0 & ~i_13_378_4568_0))) | (~i_13_378_1570_0 & ~i_13_378_3900_0 & ((~i_13_378_1525_0 & ~i_13_378_3006_0 & ~i_13_378_3485_0) | (~i_13_378_1848_0 & ~i_13_378_3763_0))) | (~i_13_378_1525_0 & ((i_13_378_4063_0 & i_13_378_4513_0) | (~i_13_378_1327_0 & ~i_13_378_4513_0))) | (~i_13_378_517_0 & ~i_13_378_652_0 & i_13_378_2406_0 & ~i_13_378_3108_0) | (~i_13_378_1848_0 & i_13_378_2002_0 & i_13_378_3108_0 & i_13_378_3730_0) | (i_13_378_31_0 & ~i_13_378_2406_0 & ~i_13_378_3817_0 & ~i_13_378_3861_0 & ~i_13_378_4452_0) | (~i_13_378_237_0 & i_13_378_535_0 & ~i_13_378_4564_0) | (i_13_378_1219_0 & i_13_378_4568_0));
endmodule



// Benchmark "kernel_13_379" written by ABC on Sun Jul 19 10:50:40 2020

module kernel_13_379 ( 
    i_13_379_28_0, i_13_379_100_0, i_13_379_109_0, i_13_379_163_0,
    i_13_379_184_0, i_13_379_298_0, i_13_379_317_0, i_13_379_382_0,
    i_13_379_415_0, i_13_379_416_0, i_13_379_470_0, i_13_379_568_0,
    i_13_379_640_0, i_13_379_686_0, i_13_379_743_0, i_13_379_794_0,
    i_13_379_797_0, i_13_379_856_0, i_13_379_886_0, i_13_379_947_0,
    i_13_379_1072_0, i_13_379_1073_0, i_13_379_1093_0, i_13_379_1129_0,
    i_13_379_1225_0, i_13_379_1252_0, i_13_379_1253_0, i_13_379_1268_0,
    i_13_379_1280_0, i_13_379_1301_0, i_13_379_1361_0, i_13_379_1424_0,
    i_13_379_1484_0, i_13_379_1486_0, i_13_379_1499_0, i_13_379_1526_0,
    i_13_379_1550_0, i_13_379_1603_0, i_13_379_1621_0, i_13_379_1631_0,
    i_13_379_1690_0, i_13_379_1691_0, i_13_379_1720_0, i_13_379_1814_0,
    i_13_379_2000_0, i_13_379_2237_0, i_13_379_2260_0, i_13_379_2444_0,
    i_13_379_2458_0, i_13_379_2459_0, i_13_379_2498_0, i_13_379_2503_0,
    i_13_379_2506_0, i_13_379_2530_0, i_13_379_2535_0, i_13_379_2539_0,
    i_13_379_2560_0, i_13_379_2567_0, i_13_379_2576_0, i_13_379_2600_0,
    i_13_379_2611_0, i_13_379_2612_0, i_13_379_2675_0, i_13_379_2882_0,
    i_13_379_2948_0, i_13_379_3136_0, i_13_379_3344_0, i_13_379_3349_0,
    i_13_379_3388_0, i_13_379_3457_0, i_13_379_3458_0, i_13_379_3476_0,
    i_13_379_3529_0, i_13_379_3539_0, i_13_379_3544_0, i_13_379_3566_0,
    i_13_379_3619_0, i_13_379_3620_0, i_13_379_3638_0, i_13_379_3683_0,
    i_13_379_3718_0, i_13_379_3739_0, i_13_379_3766_0, i_13_379_3818_0,
    i_13_379_3844_0, i_13_379_3845_0, i_13_379_3908_0, i_13_379_3920_0,
    i_13_379_3983_0, i_13_379_4007_0, i_13_379_4186_0, i_13_379_4204_0,
    i_13_379_4315_0, i_13_379_4330_0, i_13_379_4339_0, i_13_379_4340_0,
    i_13_379_4342_0, i_13_379_4519_0, i_13_379_4582_0, i_13_379_4595_0,
    o_13_379_0_0  );
  input  i_13_379_28_0, i_13_379_100_0, i_13_379_109_0, i_13_379_163_0,
    i_13_379_184_0, i_13_379_298_0, i_13_379_317_0, i_13_379_382_0,
    i_13_379_415_0, i_13_379_416_0, i_13_379_470_0, i_13_379_568_0,
    i_13_379_640_0, i_13_379_686_0, i_13_379_743_0, i_13_379_794_0,
    i_13_379_797_0, i_13_379_856_0, i_13_379_886_0, i_13_379_947_0,
    i_13_379_1072_0, i_13_379_1073_0, i_13_379_1093_0, i_13_379_1129_0,
    i_13_379_1225_0, i_13_379_1252_0, i_13_379_1253_0, i_13_379_1268_0,
    i_13_379_1280_0, i_13_379_1301_0, i_13_379_1361_0, i_13_379_1424_0,
    i_13_379_1484_0, i_13_379_1486_0, i_13_379_1499_0, i_13_379_1526_0,
    i_13_379_1550_0, i_13_379_1603_0, i_13_379_1621_0, i_13_379_1631_0,
    i_13_379_1690_0, i_13_379_1691_0, i_13_379_1720_0, i_13_379_1814_0,
    i_13_379_2000_0, i_13_379_2237_0, i_13_379_2260_0, i_13_379_2444_0,
    i_13_379_2458_0, i_13_379_2459_0, i_13_379_2498_0, i_13_379_2503_0,
    i_13_379_2506_0, i_13_379_2530_0, i_13_379_2535_0, i_13_379_2539_0,
    i_13_379_2560_0, i_13_379_2567_0, i_13_379_2576_0, i_13_379_2600_0,
    i_13_379_2611_0, i_13_379_2612_0, i_13_379_2675_0, i_13_379_2882_0,
    i_13_379_2948_0, i_13_379_3136_0, i_13_379_3344_0, i_13_379_3349_0,
    i_13_379_3388_0, i_13_379_3457_0, i_13_379_3458_0, i_13_379_3476_0,
    i_13_379_3529_0, i_13_379_3539_0, i_13_379_3544_0, i_13_379_3566_0,
    i_13_379_3619_0, i_13_379_3620_0, i_13_379_3638_0, i_13_379_3683_0,
    i_13_379_3718_0, i_13_379_3739_0, i_13_379_3766_0, i_13_379_3818_0,
    i_13_379_3844_0, i_13_379_3845_0, i_13_379_3908_0, i_13_379_3920_0,
    i_13_379_3983_0, i_13_379_4007_0, i_13_379_4186_0, i_13_379_4204_0,
    i_13_379_4315_0, i_13_379_4330_0, i_13_379_4339_0, i_13_379_4340_0,
    i_13_379_4342_0, i_13_379_4519_0, i_13_379_4582_0, i_13_379_4595_0;
  output o_13_379_0_0;
  assign o_13_379_0_0 = ~((~i_13_379_2530_0 & ((~i_13_379_28_0 & ~i_13_379_416_0 & ~i_13_379_947_0) | (~i_13_379_1072_0 & ~i_13_379_3458_0))) | (~i_13_379_2948_0 & (~i_13_379_1486_0 | ~i_13_379_2539_0 | ~i_13_379_3844_0)) | (~i_13_379_415_0 & ~i_13_379_2612_0 & i_13_379_3766_0) | (~i_13_379_1603_0 & ~i_13_379_3766_0) | (~i_13_379_3529_0 & ~i_13_379_3983_0 & ~i_13_379_4330_0));
endmodule



// Benchmark "kernel_13_380" written by ABC on Sun Jul 19 10:50:41 2020

module kernel_13_380 ( 
    i_13_380_48_0, i_13_380_78_0, i_13_380_102_0, i_13_380_121_0,
    i_13_380_157_0, i_13_380_169_0, i_13_380_188_0, i_13_380_197_0,
    i_13_380_259_0, i_13_380_274_0, i_13_380_275_0, i_13_380_283_0,
    i_13_380_337_0, i_13_380_338_0, i_13_380_431_0, i_13_380_454_0,
    i_13_380_556_0, i_13_380_588_0, i_13_380_612_0, i_13_380_616_0,
    i_13_380_620_0, i_13_380_664_0, i_13_380_669_0, i_13_380_709_0,
    i_13_380_850_0, i_13_380_926_0, i_13_380_953_0, i_13_380_1191_0,
    i_13_380_1301_0, i_13_380_1329_0, i_13_380_1346_0, i_13_380_1377_0,
    i_13_380_1399_0, i_13_380_1400_0, i_13_380_1469_0, i_13_380_1529_0,
    i_13_380_1571_0, i_13_380_1643_0, i_13_380_1678_0, i_13_380_1724_0,
    i_13_380_1727_0, i_13_380_1735_0, i_13_380_1736_0, i_13_380_1750_0,
    i_13_380_1852_0, i_13_380_1921_0, i_13_380_1993_0, i_13_380_2002_0,
    i_13_380_2081_0, i_13_380_2118_0, i_13_380_2137_0, i_13_380_2138_0,
    i_13_380_2148_0, i_13_380_2191_0, i_13_380_2210_0, i_13_380_2363_0,
    i_13_380_2408_0, i_13_380_2425_0, i_13_380_2542_0, i_13_380_2617_0,
    i_13_380_2618_0, i_13_380_2699_0, i_13_380_2708_0, i_13_380_2786_0,
    i_13_380_2885_0, i_13_380_2888_0, i_13_380_3027_0, i_13_380_3038_0,
    i_13_380_3039_0, i_13_380_3040_0, i_13_380_3041_0, i_13_380_3050_0,
    i_13_380_3145_0, i_13_380_3217_0, i_13_380_3386_0, i_13_380_3491_0,
    i_13_380_3536_0, i_13_380_3640_0, i_13_380_3641_0, i_13_380_3644_0,
    i_13_380_3702_0, i_13_380_3705_0, i_13_380_3730_0, i_13_380_3758_0,
    i_13_380_3787_0, i_13_380_3892_0, i_13_380_4089_0, i_13_380_4136_0,
    i_13_380_4230_0, i_13_380_4232_0, i_13_380_4234_0, i_13_380_4235_0,
    i_13_380_4261_0, i_13_380_4262_0, i_13_380_4305_0, i_13_380_4360_0,
    i_13_380_4436_0, i_13_380_4449_0, i_13_380_4513_0, i_13_380_4531_0,
    o_13_380_0_0  );
  input  i_13_380_48_0, i_13_380_78_0, i_13_380_102_0, i_13_380_121_0,
    i_13_380_157_0, i_13_380_169_0, i_13_380_188_0, i_13_380_197_0,
    i_13_380_259_0, i_13_380_274_0, i_13_380_275_0, i_13_380_283_0,
    i_13_380_337_0, i_13_380_338_0, i_13_380_431_0, i_13_380_454_0,
    i_13_380_556_0, i_13_380_588_0, i_13_380_612_0, i_13_380_616_0,
    i_13_380_620_0, i_13_380_664_0, i_13_380_669_0, i_13_380_709_0,
    i_13_380_850_0, i_13_380_926_0, i_13_380_953_0, i_13_380_1191_0,
    i_13_380_1301_0, i_13_380_1329_0, i_13_380_1346_0, i_13_380_1377_0,
    i_13_380_1399_0, i_13_380_1400_0, i_13_380_1469_0, i_13_380_1529_0,
    i_13_380_1571_0, i_13_380_1643_0, i_13_380_1678_0, i_13_380_1724_0,
    i_13_380_1727_0, i_13_380_1735_0, i_13_380_1736_0, i_13_380_1750_0,
    i_13_380_1852_0, i_13_380_1921_0, i_13_380_1993_0, i_13_380_2002_0,
    i_13_380_2081_0, i_13_380_2118_0, i_13_380_2137_0, i_13_380_2138_0,
    i_13_380_2148_0, i_13_380_2191_0, i_13_380_2210_0, i_13_380_2363_0,
    i_13_380_2408_0, i_13_380_2425_0, i_13_380_2542_0, i_13_380_2617_0,
    i_13_380_2618_0, i_13_380_2699_0, i_13_380_2708_0, i_13_380_2786_0,
    i_13_380_2885_0, i_13_380_2888_0, i_13_380_3027_0, i_13_380_3038_0,
    i_13_380_3039_0, i_13_380_3040_0, i_13_380_3041_0, i_13_380_3050_0,
    i_13_380_3145_0, i_13_380_3217_0, i_13_380_3386_0, i_13_380_3491_0,
    i_13_380_3536_0, i_13_380_3640_0, i_13_380_3641_0, i_13_380_3644_0,
    i_13_380_3702_0, i_13_380_3705_0, i_13_380_3730_0, i_13_380_3758_0,
    i_13_380_3787_0, i_13_380_3892_0, i_13_380_4089_0, i_13_380_4136_0,
    i_13_380_4230_0, i_13_380_4232_0, i_13_380_4234_0, i_13_380_4235_0,
    i_13_380_4261_0, i_13_380_4262_0, i_13_380_4305_0, i_13_380_4360_0,
    i_13_380_4436_0, i_13_380_4449_0, i_13_380_4513_0, i_13_380_4531_0;
  output o_13_380_0_0;
  assign o_13_380_0_0 = ~((~i_13_380_4436_0 & (~i_13_380_2617_0 | (~i_13_380_1329_0 & i_13_380_2542_0 & ~i_13_380_3758_0))) | (i_13_380_1750_0 & i_13_380_2425_0) | (~i_13_380_2888_0 & ~i_13_380_3039_0 & ~i_13_380_3536_0 & ~i_13_380_4305_0));
endmodule



// Benchmark "kernel_13_381" written by ABC on Sun Jul 19 10:50:42 2020

module kernel_13_381 ( 
    i_13_381_112_0, i_13_381_175_0, i_13_381_178_0, i_13_381_186_0,
    i_13_381_225_0, i_13_381_237_0, i_13_381_273_0, i_13_381_282_0,
    i_13_381_283_0, i_13_381_310_0, i_13_381_361_0, i_13_381_375_0,
    i_13_381_469_0, i_13_381_471_0, i_13_381_490_0, i_13_381_573_0,
    i_13_381_574_0, i_13_381_642_0, i_13_381_643_0, i_13_381_645_0,
    i_13_381_646_0, i_13_381_647_0, i_13_381_687_0, i_13_381_688_0,
    i_13_381_690_0, i_13_381_691_0, i_13_381_702_0, i_13_381_717_0,
    i_13_381_760_0, i_13_381_862_0, i_13_381_1123_0, i_13_381_1267_0,
    i_13_381_1308_0, i_13_381_1311_0, i_13_381_1313_0, i_13_381_1399_0,
    i_13_381_1597_0, i_13_381_1641_0, i_13_381_1642_0, i_13_381_1672_0,
    i_13_381_1804_0, i_13_381_1857_0, i_13_381_1860_0, i_13_381_1861_0,
    i_13_381_1884_0, i_13_381_1939_0, i_13_381_2002_0, i_13_381_2029_0,
    i_13_381_2055_0, i_13_381_2136_0, i_13_381_2137_0, i_13_381_2176_0,
    i_13_381_2193_0, i_13_381_2263_0, i_13_381_2310_0, i_13_381_2427_0,
    i_13_381_2586_0, i_13_381_2599_0, i_13_381_2649_0, i_13_381_2650_0,
    i_13_381_2652_0, i_13_381_2653_0, i_13_381_2654_0, i_13_381_2676_0,
    i_13_381_2677_0, i_13_381_2680_0, i_13_381_2770_0, i_13_381_2847_0,
    i_13_381_2851_0, i_13_381_2913_0, i_13_381_2964_0, i_13_381_3003_0,
    i_13_381_3270_0, i_13_381_3271_0, i_13_381_3273_0, i_13_381_3274_0,
    i_13_381_3315_0, i_13_381_3378_0, i_13_381_3387_0, i_13_381_3423_0,
    i_13_381_3424_0, i_13_381_3426_0, i_13_381_3427_0, i_13_381_3478_0,
    i_13_381_3535_0, i_13_381_3639_0, i_13_381_3732_0, i_13_381_3875_0,
    i_13_381_3913_0, i_13_381_4018_0, i_13_381_4020_0, i_13_381_4045_0,
    i_13_381_4077_0, i_13_381_4080_0, i_13_381_4084_0, i_13_381_4162_0,
    i_13_381_4174_0, i_13_381_4219_0, i_13_381_4426_0, i_13_381_4594_0,
    o_13_381_0_0  );
  input  i_13_381_112_0, i_13_381_175_0, i_13_381_178_0, i_13_381_186_0,
    i_13_381_225_0, i_13_381_237_0, i_13_381_273_0, i_13_381_282_0,
    i_13_381_283_0, i_13_381_310_0, i_13_381_361_0, i_13_381_375_0,
    i_13_381_469_0, i_13_381_471_0, i_13_381_490_0, i_13_381_573_0,
    i_13_381_574_0, i_13_381_642_0, i_13_381_643_0, i_13_381_645_0,
    i_13_381_646_0, i_13_381_647_0, i_13_381_687_0, i_13_381_688_0,
    i_13_381_690_0, i_13_381_691_0, i_13_381_702_0, i_13_381_717_0,
    i_13_381_760_0, i_13_381_862_0, i_13_381_1123_0, i_13_381_1267_0,
    i_13_381_1308_0, i_13_381_1311_0, i_13_381_1313_0, i_13_381_1399_0,
    i_13_381_1597_0, i_13_381_1641_0, i_13_381_1642_0, i_13_381_1672_0,
    i_13_381_1804_0, i_13_381_1857_0, i_13_381_1860_0, i_13_381_1861_0,
    i_13_381_1884_0, i_13_381_1939_0, i_13_381_2002_0, i_13_381_2029_0,
    i_13_381_2055_0, i_13_381_2136_0, i_13_381_2137_0, i_13_381_2176_0,
    i_13_381_2193_0, i_13_381_2263_0, i_13_381_2310_0, i_13_381_2427_0,
    i_13_381_2586_0, i_13_381_2599_0, i_13_381_2649_0, i_13_381_2650_0,
    i_13_381_2652_0, i_13_381_2653_0, i_13_381_2654_0, i_13_381_2676_0,
    i_13_381_2677_0, i_13_381_2680_0, i_13_381_2770_0, i_13_381_2847_0,
    i_13_381_2851_0, i_13_381_2913_0, i_13_381_2964_0, i_13_381_3003_0,
    i_13_381_3270_0, i_13_381_3271_0, i_13_381_3273_0, i_13_381_3274_0,
    i_13_381_3315_0, i_13_381_3378_0, i_13_381_3387_0, i_13_381_3423_0,
    i_13_381_3424_0, i_13_381_3426_0, i_13_381_3427_0, i_13_381_3478_0,
    i_13_381_3535_0, i_13_381_3639_0, i_13_381_3732_0, i_13_381_3875_0,
    i_13_381_3913_0, i_13_381_4018_0, i_13_381_4020_0, i_13_381_4045_0,
    i_13_381_4077_0, i_13_381_4080_0, i_13_381_4084_0, i_13_381_4162_0,
    i_13_381_4174_0, i_13_381_4219_0, i_13_381_4426_0, i_13_381_4594_0;
  output o_13_381_0_0;
  assign o_13_381_0_0 = ~(~i_13_381_4080_0 | (~i_13_381_690_0 & ~i_13_381_2652_0) | (~i_13_381_574_0 & ~i_13_381_2649_0));
endmodule



// Benchmark "kernel_13_382" written by ABC on Sun Jul 19 10:50:42 2020

module kernel_13_382 ( 
    i_13_382_51_0, i_13_382_52_0, i_13_382_105_0, i_13_382_106_0,
    i_13_382_312_0, i_13_382_313_0, i_13_382_337_0, i_13_382_381_0,
    i_13_382_409_0, i_13_382_420_0, i_13_382_427_0, i_13_382_484_0,
    i_13_382_507_0, i_13_382_526_0, i_13_382_553_0, i_13_382_609_0,
    i_13_382_654_0, i_13_382_678_0, i_13_382_679_0, i_13_382_691_0,
    i_13_382_735_0, i_13_382_843_0, i_13_382_844_0, i_13_382_961_0,
    i_13_382_1042_0, i_13_382_1303_0, i_13_382_1311_0, i_13_382_1329_0,
    i_13_382_1330_0, i_13_382_1345_0, i_13_382_1407_0, i_13_382_1462_0,
    i_13_382_1518_0, i_13_382_1519_0, i_13_382_1572_0, i_13_382_1573_0,
    i_13_382_1677_0, i_13_382_1686_0, i_13_382_1813_0, i_13_382_1861_0,
    i_13_382_1911_0, i_13_382_2004_0, i_13_382_2023_0, i_13_382_2031_0,
    i_13_382_2049_0, i_13_382_2094_0, i_13_382_2131_0, i_13_382_2191_0,
    i_13_382_2209_0, i_13_382_2281_0, i_13_382_2596_0, i_13_382_2640_0,
    i_13_382_2695_0, i_13_382_2698_0, i_13_382_2722_0, i_13_382_2856_0,
    i_13_382_2928_0, i_13_382_2938_0, i_13_382_2982_0, i_13_382_2985_0,
    i_13_382_3090_0, i_13_382_3127_0, i_13_382_3217_0, i_13_382_3291_0,
    i_13_382_3364_0, i_13_382_3370_0, i_13_382_3372_0, i_13_382_3400_0,
    i_13_382_3417_0, i_13_382_3439_0, i_13_382_3490_0, i_13_382_3525_0,
    i_13_382_3526_0, i_13_382_3535_0, i_13_382_3549_0, i_13_382_3561_0,
    i_13_382_3616_0, i_13_382_3618_0, i_13_382_3648_0, i_13_382_3768_0,
    i_13_382_3769_0, i_13_382_3822_0, i_13_382_3864_0, i_13_382_3865_0,
    i_13_382_3891_0, i_13_382_3993_0, i_13_382_4035_0, i_13_382_4047_0,
    i_13_382_4119_0, i_13_382_4120_0, i_13_382_4161_0, i_13_382_4162_0,
    i_13_382_4191_0, i_13_382_4270_0, i_13_382_4369_0, i_13_382_4567_0,
    i_13_382_4597_0, i_13_382_4599_0, i_13_382_4602_0, i_13_382_4603_0,
    o_13_382_0_0  );
  input  i_13_382_51_0, i_13_382_52_0, i_13_382_105_0, i_13_382_106_0,
    i_13_382_312_0, i_13_382_313_0, i_13_382_337_0, i_13_382_381_0,
    i_13_382_409_0, i_13_382_420_0, i_13_382_427_0, i_13_382_484_0,
    i_13_382_507_0, i_13_382_526_0, i_13_382_553_0, i_13_382_609_0,
    i_13_382_654_0, i_13_382_678_0, i_13_382_679_0, i_13_382_691_0,
    i_13_382_735_0, i_13_382_843_0, i_13_382_844_0, i_13_382_961_0,
    i_13_382_1042_0, i_13_382_1303_0, i_13_382_1311_0, i_13_382_1329_0,
    i_13_382_1330_0, i_13_382_1345_0, i_13_382_1407_0, i_13_382_1462_0,
    i_13_382_1518_0, i_13_382_1519_0, i_13_382_1572_0, i_13_382_1573_0,
    i_13_382_1677_0, i_13_382_1686_0, i_13_382_1813_0, i_13_382_1861_0,
    i_13_382_1911_0, i_13_382_2004_0, i_13_382_2023_0, i_13_382_2031_0,
    i_13_382_2049_0, i_13_382_2094_0, i_13_382_2131_0, i_13_382_2191_0,
    i_13_382_2209_0, i_13_382_2281_0, i_13_382_2596_0, i_13_382_2640_0,
    i_13_382_2695_0, i_13_382_2698_0, i_13_382_2722_0, i_13_382_2856_0,
    i_13_382_2928_0, i_13_382_2938_0, i_13_382_2982_0, i_13_382_2985_0,
    i_13_382_3090_0, i_13_382_3127_0, i_13_382_3217_0, i_13_382_3291_0,
    i_13_382_3364_0, i_13_382_3370_0, i_13_382_3372_0, i_13_382_3400_0,
    i_13_382_3417_0, i_13_382_3439_0, i_13_382_3490_0, i_13_382_3525_0,
    i_13_382_3526_0, i_13_382_3535_0, i_13_382_3549_0, i_13_382_3561_0,
    i_13_382_3616_0, i_13_382_3618_0, i_13_382_3648_0, i_13_382_3768_0,
    i_13_382_3769_0, i_13_382_3822_0, i_13_382_3864_0, i_13_382_3865_0,
    i_13_382_3891_0, i_13_382_3993_0, i_13_382_4035_0, i_13_382_4047_0,
    i_13_382_4119_0, i_13_382_4120_0, i_13_382_4161_0, i_13_382_4162_0,
    i_13_382_4191_0, i_13_382_4270_0, i_13_382_4369_0, i_13_382_4567_0,
    i_13_382_4597_0, i_13_382_4599_0, i_13_382_4602_0, i_13_382_4603_0;
  output o_13_382_0_0;
  assign o_13_382_0_0 = ~((~i_13_382_4047_0 & ~i_13_382_4369_0) | (~i_13_382_2698_0 & ~i_13_382_4191_0) | (i_13_382_3490_0 & ~i_13_382_4035_0) | (~i_13_382_691_0 & ~i_13_382_3822_0) | (~i_13_382_2131_0 & ~i_13_382_2985_0));
endmodule



// Benchmark "kernel_13_383" written by ABC on Sun Jul 19 10:50:43 2020

module kernel_13_383 ( 
    i_13_383_33_0, i_13_383_76_0, i_13_383_111_0, i_13_383_120_0,
    i_13_383_159_0, i_13_383_160_0, i_13_383_271_0, i_13_383_285_0,
    i_13_383_313_0, i_13_383_322_0, i_13_383_384_0, i_13_383_385_0,
    i_13_383_456_0, i_13_383_511_0, i_13_383_537_0, i_13_383_564_0,
    i_13_383_570_0, i_13_383_611_0, i_13_383_643_0, i_13_383_655_0,
    i_13_383_760_0, i_13_383_840_0, i_13_383_943_0, i_13_383_1086_0,
    i_13_383_1087_0, i_13_383_1218_0, i_13_383_1255_0, i_13_383_1302_0,
    i_13_383_1303_0, i_13_383_1443_0, i_13_383_1473_0, i_13_383_1477_0,
    i_13_383_1489_0, i_13_383_1509_0, i_13_383_1599_0, i_13_383_1635_0,
    i_13_383_1636_0, i_13_383_1650_0, i_13_383_1735_0, i_13_383_1789_0,
    i_13_383_1795_0, i_13_383_1995_0, i_13_383_2056_0, i_13_383_2112_0,
    i_13_383_2122_0, i_13_383_2173_0, i_13_383_2193_0, i_13_383_2208_0,
    i_13_383_2242_0, i_13_383_2400_0, i_13_383_2424_0, i_13_383_2436_0,
    i_13_383_2500_0, i_13_383_2532_0, i_13_383_2541_0, i_13_383_2715_0,
    i_13_383_2716_0, i_13_383_2847_0, i_13_383_2919_0, i_13_383_2941_0,
    i_13_383_3000_0, i_13_383_3004_0, i_13_383_3022_0, i_13_383_3028_0,
    i_13_383_3103_0, i_13_383_3129_0, i_13_383_3147_0, i_13_383_3163_0,
    i_13_383_3172_0, i_13_383_3261_0, i_13_383_3274_0, i_13_383_3321_0,
    i_13_383_3346_0, i_13_383_3382_0, i_13_383_3388_0, i_13_383_3580_0,
    i_13_383_3615_0, i_13_383_3616_0, i_13_383_3702_0, i_13_383_3720_0,
    i_13_383_3783_0, i_13_383_3796_0, i_13_383_3802_0, i_13_383_3846_0,
    i_13_383_3873_0, i_13_383_3874_0, i_13_383_3910_0, i_13_383_4008_0,
    i_13_383_4009_0, i_13_383_4036_0, i_13_383_4045_0, i_13_383_4083_0,
    i_13_383_4084_0, i_13_383_4093_0, i_13_383_4107_0, i_13_383_4120_0,
    i_13_383_4236_0, i_13_383_4282_0, i_13_383_4336_0, i_13_383_4417_0,
    o_13_383_0_0  );
  input  i_13_383_33_0, i_13_383_76_0, i_13_383_111_0, i_13_383_120_0,
    i_13_383_159_0, i_13_383_160_0, i_13_383_271_0, i_13_383_285_0,
    i_13_383_313_0, i_13_383_322_0, i_13_383_384_0, i_13_383_385_0,
    i_13_383_456_0, i_13_383_511_0, i_13_383_537_0, i_13_383_564_0,
    i_13_383_570_0, i_13_383_611_0, i_13_383_643_0, i_13_383_655_0,
    i_13_383_760_0, i_13_383_840_0, i_13_383_943_0, i_13_383_1086_0,
    i_13_383_1087_0, i_13_383_1218_0, i_13_383_1255_0, i_13_383_1302_0,
    i_13_383_1303_0, i_13_383_1443_0, i_13_383_1473_0, i_13_383_1477_0,
    i_13_383_1489_0, i_13_383_1509_0, i_13_383_1599_0, i_13_383_1635_0,
    i_13_383_1636_0, i_13_383_1650_0, i_13_383_1735_0, i_13_383_1789_0,
    i_13_383_1795_0, i_13_383_1995_0, i_13_383_2056_0, i_13_383_2112_0,
    i_13_383_2122_0, i_13_383_2173_0, i_13_383_2193_0, i_13_383_2208_0,
    i_13_383_2242_0, i_13_383_2400_0, i_13_383_2424_0, i_13_383_2436_0,
    i_13_383_2500_0, i_13_383_2532_0, i_13_383_2541_0, i_13_383_2715_0,
    i_13_383_2716_0, i_13_383_2847_0, i_13_383_2919_0, i_13_383_2941_0,
    i_13_383_3000_0, i_13_383_3004_0, i_13_383_3022_0, i_13_383_3028_0,
    i_13_383_3103_0, i_13_383_3129_0, i_13_383_3147_0, i_13_383_3163_0,
    i_13_383_3172_0, i_13_383_3261_0, i_13_383_3274_0, i_13_383_3321_0,
    i_13_383_3346_0, i_13_383_3382_0, i_13_383_3388_0, i_13_383_3580_0,
    i_13_383_3615_0, i_13_383_3616_0, i_13_383_3702_0, i_13_383_3720_0,
    i_13_383_3783_0, i_13_383_3796_0, i_13_383_3802_0, i_13_383_3846_0,
    i_13_383_3873_0, i_13_383_3874_0, i_13_383_3910_0, i_13_383_4008_0,
    i_13_383_4009_0, i_13_383_4036_0, i_13_383_4045_0, i_13_383_4083_0,
    i_13_383_4084_0, i_13_383_4093_0, i_13_383_4107_0, i_13_383_4120_0,
    i_13_383_4236_0, i_13_383_4282_0, i_13_383_4336_0, i_13_383_4417_0;
  output o_13_383_0_0;
  assign o_13_383_0_0 = ~((~i_13_383_2424_0 & ~i_13_383_2716_0) | (~i_13_383_537_0 & ~i_13_383_1509_0));
endmodule



// Benchmark "kernel_13_384" written by ABC on Sun Jul 19 10:50:44 2020

module kernel_13_384 ( 
    i_13_384_66_0, i_13_384_69_0, i_13_384_70_0, i_13_384_133_0,
    i_13_384_205_0, i_13_384_208_0, i_13_384_209_0, i_13_384_357_0,
    i_13_384_466_0, i_13_384_535_0, i_13_384_588_0, i_13_384_591_0,
    i_13_384_616_0, i_13_384_653_0, i_13_384_745_0, i_13_384_762_0,
    i_13_384_763_0, i_13_384_814_0, i_13_384_1073_0, i_13_384_1131_0,
    i_13_384_1132_0, i_13_384_1302_0, i_13_384_1303_0, i_13_384_1312_0,
    i_13_384_1347_0, i_13_384_1445_0, i_13_384_1453_0, i_13_384_1523_0,
    i_13_384_1524_0, i_13_384_1525_0, i_13_384_1605_0, i_13_384_1649_0,
    i_13_384_1650_0, i_13_384_1699_0, i_13_384_1717_0, i_13_384_1930_0,
    i_13_384_1932_0, i_13_384_1933_0, i_13_384_1995_0, i_13_384_2103_0,
    i_13_384_2125_0, i_13_384_2128_0, i_13_384_2135_0, i_13_384_2145_0,
    i_13_384_2193_0, i_13_384_2194_0, i_13_384_2195_0, i_13_384_2239_0,
    i_13_384_2380_0, i_13_384_2418_0, i_13_384_2435_0, i_13_384_2472_0,
    i_13_384_2553_0, i_13_384_2697_0, i_13_384_2698_0, i_13_384_2699_0,
    i_13_384_2721_0, i_13_384_2770_0, i_13_384_3129_0, i_13_384_3244_0,
    i_13_384_3272_0, i_13_384_3308_0, i_13_384_3344_0, i_13_384_3403_0,
    i_13_384_3541_0, i_13_384_3634_0, i_13_384_3637_0, i_13_384_3639_0,
    i_13_384_3640_0, i_13_384_3666_0, i_13_384_3718_0, i_13_384_3742_0,
    i_13_384_3757_0, i_13_384_3766_0, i_13_384_3844_0, i_13_384_3847_0,
    i_13_384_3871_0, i_13_384_3900_0, i_13_384_3918_0, i_13_384_3940_0,
    i_13_384_3973_0, i_13_384_3985_0, i_13_384_3994_0, i_13_384_4010_0,
    i_13_384_4035_0, i_13_384_4036_0, i_13_384_4038_0, i_13_384_4039_0,
    i_13_384_4060_0, i_13_384_4225_0, i_13_384_4236_0, i_13_384_4272_0,
    i_13_384_4273_0, i_13_384_4295_0, i_13_384_4309_0, i_13_384_4312_0,
    i_13_384_4398_0, i_13_384_4593_0, i_13_384_4596_0, i_13_384_4606_0,
    o_13_384_0_0  );
  input  i_13_384_66_0, i_13_384_69_0, i_13_384_70_0, i_13_384_133_0,
    i_13_384_205_0, i_13_384_208_0, i_13_384_209_0, i_13_384_357_0,
    i_13_384_466_0, i_13_384_535_0, i_13_384_588_0, i_13_384_591_0,
    i_13_384_616_0, i_13_384_653_0, i_13_384_745_0, i_13_384_762_0,
    i_13_384_763_0, i_13_384_814_0, i_13_384_1073_0, i_13_384_1131_0,
    i_13_384_1132_0, i_13_384_1302_0, i_13_384_1303_0, i_13_384_1312_0,
    i_13_384_1347_0, i_13_384_1445_0, i_13_384_1453_0, i_13_384_1523_0,
    i_13_384_1524_0, i_13_384_1525_0, i_13_384_1605_0, i_13_384_1649_0,
    i_13_384_1650_0, i_13_384_1699_0, i_13_384_1717_0, i_13_384_1930_0,
    i_13_384_1932_0, i_13_384_1933_0, i_13_384_1995_0, i_13_384_2103_0,
    i_13_384_2125_0, i_13_384_2128_0, i_13_384_2135_0, i_13_384_2145_0,
    i_13_384_2193_0, i_13_384_2194_0, i_13_384_2195_0, i_13_384_2239_0,
    i_13_384_2380_0, i_13_384_2418_0, i_13_384_2435_0, i_13_384_2472_0,
    i_13_384_2553_0, i_13_384_2697_0, i_13_384_2698_0, i_13_384_2699_0,
    i_13_384_2721_0, i_13_384_2770_0, i_13_384_3129_0, i_13_384_3244_0,
    i_13_384_3272_0, i_13_384_3308_0, i_13_384_3344_0, i_13_384_3403_0,
    i_13_384_3541_0, i_13_384_3634_0, i_13_384_3637_0, i_13_384_3639_0,
    i_13_384_3640_0, i_13_384_3666_0, i_13_384_3718_0, i_13_384_3742_0,
    i_13_384_3757_0, i_13_384_3766_0, i_13_384_3844_0, i_13_384_3847_0,
    i_13_384_3871_0, i_13_384_3900_0, i_13_384_3918_0, i_13_384_3940_0,
    i_13_384_3973_0, i_13_384_3985_0, i_13_384_3994_0, i_13_384_4010_0,
    i_13_384_4035_0, i_13_384_4036_0, i_13_384_4038_0, i_13_384_4039_0,
    i_13_384_4060_0, i_13_384_4225_0, i_13_384_4236_0, i_13_384_4272_0,
    i_13_384_4273_0, i_13_384_4295_0, i_13_384_4309_0, i_13_384_4312_0,
    i_13_384_4398_0, i_13_384_4593_0, i_13_384_4596_0, i_13_384_4606_0;
  output o_13_384_0_0;
  assign o_13_384_0_0 = ~(~i_13_384_762_0 | (~i_13_384_616_0 & i_13_384_3994_0));
endmodule



// Benchmark "kernel_13_385" written by ABC on Sun Jul 19 10:50:45 2020

module kernel_13_385 ( 
    i_13_385_76_0, i_13_385_79_0, i_13_385_115_0, i_13_385_285_0,
    i_13_385_409_0, i_13_385_471_0, i_13_385_520_0, i_13_385_525_0,
    i_13_385_597_0, i_13_385_609_0, i_13_385_660_0, i_13_385_663_0,
    i_13_385_664_0, i_13_385_700_0, i_13_385_798_0, i_13_385_825_0,
    i_13_385_831_0, i_13_385_841_0, i_13_385_852_0, i_13_385_940_0,
    i_13_385_942_0, i_13_385_1066_0, i_13_385_1104_0, i_13_385_1147_0,
    i_13_385_1150_0, i_13_385_1230_0, i_13_385_1231_0, i_13_385_1309_0,
    i_13_385_1311_0, i_13_385_1317_0, i_13_385_1492_0, i_13_385_1497_0,
    i_13_385_1524_0, i_13_385_1551_0, i_13_385_1599_0, i_13_385_1659_0,
    i_13_385_1660_0, i_13_385_1744_0, i_13_385_1794_0, i_13_385_1884_0,
    i_13_385_1921_0, i_13_385_1929_0, i_13_385_1959_0, i_13_385_1960_0,
    i_13_385_1965_0, i_13_385_2230_0, i_13_385_2299_0, i_13_385_2334_0,
    i_13_385_2356_0, i_13_385_2451_0, i_13_385_2454_0, i_13_385_2455_0,
    i_13_385_2469_0, i_13_385_2553_0, i_13_385_2724_0, i_13_385_2850_0,
    i_13_385_2883_0, i_13_385_2941_0, i_13_385_3012_0, i_13_385_3028_0,
    i_13_385_3049_0, i_13_385_3117_0, i_13_385_3135_0, i_13_385_3156_0,
    i_13_385_3388_0, i_13_385_3478_0, i_13_385_3486_0, i_13_385_3489_0,
    i_13_385_3490_0, i_13_385_3504_0, i_13_385_3541_0, i_13_385_3543_0,
    i_13_385_3544_0, i_13_385_3549_0, i_13_385_3579_0, i_13_385_3580_0,
    i_13_385_3648_0, i_13_385_3742_0, i_13_385_3894_0, i_13_385_4019_0,
    i_13_385_4054_0, i_13_385_4126_0, i_13_385_4164_0, i_13_385_4165_0,
    i_13_385_4201_0, i_13_385_4251_0, i_13_385_4254_0, i_13_385_4255_0,
    i_13_385_4263_0, i_13_385_4264_0, i_13_385_4269_0, i_13_385_4296_0,
    i_13_385_4318_0, i_13_385_4332_0, i_13_385_4333_0, i_13_385_4396_0,
    i_13_385_4431_0, i_13_385_4452_0, i_13_385_4461_0, i_13_385_4603_0,
    o_13_385_0_0  );
  input  i_13_385_76_0, i_13_385_79_0, i_13_385_115_0, i_13_385_285_0,
    i_13_385_409_0, i_13_385_471_0, i_13_385_520_0, i_13_385_525_0,
    i_13_385_597_0, i_13_385_609_0, i_13_385_660_0, i_13_385_663_0,
    i_13_385_664_0, i_13_385_700_0, i_13_385_798_0, i_13_385_825_0,
    i_13_385_831_0, i_13_385_841_0, i_13_385_852_0, i_13_385_940_0,
    i_13_385_942_0, i_13_385_1066_0, i_13_385_1104_0, i_13_385_1147_0,
    i_13_385_1150_0, i_13_385_1230_0, i_13_385_1231_0, i_13_385_1309_0,
    i_13_385_1311_0, i_13_385_1317_0, i_13_385_1492_0, i_13_385_1497_0,
    i_13_385_1524_0, i_13_385_1551_0, i_13_385_1599_0, i_13_385_1659_0,
    i_13_385_1660_0, i_13_385_1744_0, i_13_385_1794_0, i_13_385_1884_0,
    i_13_385_1921_0, i_13_385_1929_0, i_13_385_1959_0, i_13_385_1960_0,
    i_13_385_1965_0, i_13_385_2230_0, i_13_385_2299_0, i_13_385_2334_0,
    i_13_385_2356_0, i_13_385_2451_0, i_13_385_2454_0, i_13_385_2455_0,
    i_13_385_2469_0, i_13_385_2553_0, i_13_385_2724_0, i_13_385_2850_0,
    i_13_385_2883_0, i_13_385_2941_0, i_13_385_3012_0, i_13_385_3028_0,
    i_13_385_3049_0, i_13_385_3117_0, i_13_385_3135_0, i_13_385_3156_0,
    i_13_385_3388_0, i_13_385_3478_0, i_13_385_3486_0, i_13_385_3489_0,
    i_13_385_3490_0, i_13_385_3504_0, i_13_385_3541_0, i_13_385_3543_0,
    i_13_385_3544_0, i_13_385_3549_0, i_13_385_3579_0, i_13_385_3580_0,
    i_13_385_3648_0, i_13_385_3742_0, i_13_385_3894_0, i_13_385_4019_0,
    i_13_385_4054_0, i_13_385_4126_0, i_13_385_4164_0, i_13_385_4165_0,
    i_13_385_4201_0, i_13_385_4251_0, i_13_385_4254_0, i_13_385_4255_0,
    i_13_385_4263_0, i_13_385_4264_0, i_13_385_4269_0, i_13_385_4296_0,
    i_13_385_4318_0, i_13_385_4332_0, i_13_385_4333_0, i_13_385_4396_0,
    i_13_385_4431_0, i_13_385_4452_0, i_13_385_4461_0, i_13_385_4603_0;
  output o_13_385_0_0;
  assign o_13_385_0_0 = ~((~i_13_385_4251_0 & ~i_13_385_4452_0) | (~i_13_385_2883_0 & ~i_13_385_3012_0) | (~i_13_385_825_0 & ~i_13_385_1794_0 & ~i_13_385_3648_0) | (~i_13_385_115_0 & ~i_13_385_520_0 & ~i_13_385_2553_0));
endmodule



// Benchmark "kernel_13_386" written by ABC on Sun Jul 19 10:50:45 2020

module kernel_13_386 ( 
    i_13_386_36_0, i_13_386_37_0, i_13_386_72_0, i_13_386_130_0,
    i_13_386_136_0, i_13_386_163_0, i_13_386_182_0, i_13_386_186_0,
    i_13_386_216_0, i_13_386_225_0, i_13_386_279_0, i_13_386_280_0,
    i_13_386_324_0, i_13_386_375_0, i_13_386_382_0, i_13_386_407_0,
    i_13_386_532_0, i_13_386_544_0, i_13_386_595_0, i_13_386_641_0,
    i_13_386_670_0, i_13_386_680_0, i_13_386_694_0, i_13_386_714_0,
    i_13_386_724_0, i_13_386_777_0, i_13_386_823_0, i_13_386_828_0,
    i_13_386_831_0, i_13_386_848_0, i_13_386_850_0, i_13_386_891_0,
    i_13_386_976_0, i_13_386_1022_0, i_13_386_1065_0, i_13_386_1117_0,
    i_13_386_1217_0, i_13_386_1309_0, i_13_386_1332_0, i_13_386_1380_0,
    i_13_386_1390_0, i_13_386_1404_0, i_13_386_1461_0, i_13_386_1487_0,
    i_13_386_1667_0, i_13_386_1710_0, i_13_386_1711_0, i_13_386_1746_0,
    i_13_386_1828_0, i_13_386_1829_0, i_13_386_1831_0, i_13_386_1858_0,
    i_13_386_1881_0, i_13_386_1882_0, i_13_386_1884_0, i_13_386_1903_0,
    i_13_386_2093_0, i_13_386_2120_0, i_13_386_2296_0, i_13_386_2307_0,
    i_13_386_2342_0, i_13_386_2423_0, i_13_386_2435_0, i_13_386_2629_0,
    i_13_386_2646_0, i_13_386_2647_0, i_13_386_2649_0, i_13_386_2650_0,
    i_13_386_2700_0, i_13_386_2745_0, i_13_386_2844_0, i_13_386_2845_0,
    i_13_386_2871_0, i_13_386_2872_0, i_13_386_3029_0, i_13_386_3109_0,
    i_13_386_3142_0, i_13_386_3161_0, i_13_386_3171_0, i_13_386_3216_0,
    i_13_386_3241_0, i_13_386_3384_0, i_13_386_3429_0, i_13_386_3447_0,
    i_13_386_3559_0, i_13_386_3641_0, i_13_386_3784_0, i_13_386_3790_0,
    i_13_386_3817_0, i_13_386_3821_0, i_13_386_3854_0, i_13_386_3893_0,
    i_13_386_4077_0, i_13_386_4096_0, i_13_386_4162_0, i_13_386_4207_0,
    i_13_386_4348_0, i_13_386_4412_0, i_13_386_4440_0, i_13_386_4567_0,
    o_13_386_0_0  );
  input  i_13_386_36_0, i_13_386_37_0, i_13_386_72_0, i_13_386_130_0,
    i_13_386_136_0, i_13_386_163_0, i_13_386_182_0, i_13_386_186_0,
    i_13_386_216_0, i_13_386_225_0, i_13_386_279_0, i_13_386_280_0,
    i_13_386_324_0, i_13_386_375_0, i_13_386_382_0, i_13_386_407_0,
    i_13_386_532_0, i_13_386_544_0, i_13_386_595_0, i_13_386_641_0,
    i_13_386_670_0, i_13_386_680_0, i_13_386_694_0, i_13_386_714_0,
    i_13_386_724_0, i_13_386_777_0, i_13_386_823_0, i_13_386_828_0,
    i_13_386_831_0, i_13_386_848_0, i_13_386_850_0, i_13_386_891_0,
    i_13_386_976_0, i_13_386_1022_0, i_13_386_1065_0, i_13_386_1117_0,
    i_13_386_1217_0, i_13_386_1309_0, i_13_386_1332_0, i_13_386_1380_0,
    i_13_386_1390_0, i_13_386_1404_0, i_13_386_1461_0, i_13_386_1487_0,
    i_13_386_1667_0, i_13_386_1710_0, i_13_386_1711_0, i_13_386_1746_0,
    i_13_386_1828_0, i_13_386_1829_0, i_13_386_1831_0, i_13_386_1858_0,
    i_13_386_1881_0, i_13_386_1882_0, i_13_386_1884_0, i_13_386_1903_0,
    i_13_386_2093_0, i_13_386_2120_0, i_13_386_2296_0, i_13_386_2307_0,
    i_13_386_2342_0, i_13_386_2423_0, i_13_386_2435_0, i_13_386_2629_0,
    i_13_386_2646_0, i_13_386_2647_0, i_13_386_2649_0, i_13_386_2650_0,
    i_13_386_2700_0, i_13_386_2745_0, i_13_386_2844_0, i_13_386_2845_0,
    i_13_386_2871_0, i_13_386_2872_0, i_13_386_3029_0, i_13_386_3109_0,
    i_13_386_3142_0, i_13_386_3161_0, i_13_386_3171_0, i_13_386_3216_0,
    i_13_386_3241_0, i_13_386_3384_0, i_13_386_3429_0, i_13_386_3447_0,
    i_13_386_3559_0, i_13_386_3641_0, i_13_386_3784_0, i_13_386_3790_0,
    i_13_386_3817_0, i_13_386_3821_0, i_13_386_3854_0, i_13_386_3893_0,
    i_13_386_4077_0, i_13_386_4096_0, i_13_386_4162_0, i_13_386_4207_0,
    i_13_386_4348_0, i_13_386_4412_0, i_13_386_4440_0, i_13_386_4567_0;
  output o_13_386_0_0;
  assign o_13_386_0_0 = ~((~i_13_386_3142_0 & i_13_386_4412_0) | (i_13_386_182_0 & ~i_13_386_4162_0) | (~i_13_386_2650_0 & ~i_13_386_2871_0) | (~i_13_386_891_0 & ~i_13_386_2844_0 & ~i_13_386_4412_0) | (i_13_386_1831_0 & ~i_13_386_3384_0 & ~i_13_386_3447_0));
endmodule



// Benchmark "kernel_13_387" written by ABC on Sun Jul 19 10:50:46 2020

module kernel_13_387 ( 
    i_13_387_32_0, i_13_387_49_0, i_13_387_56_0, i_13_387_71_0,
    i_13_387_77_0, i_13_387_80_0, i_13_387_153_0, i_13_387_412_0,
    i_13_387_611_0, i_13_387_629_0, i_13_387_661_0, i_13_387_662_0,
    i_13_387_664_0, i_13_387_674_0, i_13_387_683_0, i_13_387_686_0,
    i_13_387_716_0, i_13_387_851_0, i_13_387_854_0, i_13_387_940_0,
    i_13_387_1060_0, i_13_387_1071_0, i_13_387_1076_0, i_13_387_1101_0,
    i_13_387_1105_0, i_13_387_1106_0, i_13_387_1133_0, i_13_387_1151_0,
    i_13_387_1188_0, i_13_387_1224_0, i_13_387_1228_0, i_13_387_1229_0,
    i_13_387_1232_0, i_13_387_1244_0, i_13_387_1256_0, i_13_387_1318_0,
    i_13_387_1345_0, i_13_387_1484_0, i_13_387_1733_0, i_13_387_1765_0,
    i_13_387_1766_0, i_13_387_1768_0, i_13_387_1787_0, i_13_387_1799_0,
    i_13_387_1892_0, i_13_387_1927_0, i_13_387_1962_0, i_13_387_2005_0,
    i_13_387_2023_0, i_13_387_2024_0, i_13_387_2026_0, i_13_387_2212_0,
    i_13_387_2284_0, i_13_387_2288_0, i_13_387_2434_0, i_13_387_2518_0,
    i_13_387_2582_0, i_13_387_2852_0, i_13_387_2903_0, i_13_387_2975_0,
    i_13_387_2987_0, i_13_387_3010_0, i_13_387_3013_0, i_13_387_3027_0,
    i_13_387_3032_0, i_13_387_3050_0, i_13_387_3064_0, i_13_387_3122_0,
    i_13_387_3261_0, i_13_387_3355_0, i_13_387_3356_0, i_13_387_3487_0,
    i_13_387_3539_0, i_13_387_3542_0, i_13_387_3573_0, i_13_387_3574_0,
    i_13_387_3731_0, i_13_387_3734_0, i_13_387_3755_0, i_13_387_3866_0,
    i_13_387_3869_0, i_13_387_3928_0, i_13_387_3978_0, i_13_387_4166_0,
    i_13_387_4212_0, i_13_387_4255_0, i_13_387_4256_0, i_13_387_4302_0,
    i_13_387_4322_0, i_13_387_4336_0, i_13_387_4343_0, i_13_387_4372_0,
    i_13_387_4373_0, i_13_387_4382_0, i_13_387_4450_0, i_13_387_4514_0,
    i_13_387_4516_0, i_13_387_4598_0, i_13_387_4606_0, i_13_387_4607_0,
    o_13_387_0_0  );
  input  i_13_387_32_0, i_13_387_49_0, i_13_387_56_0, i_13_387_71_0,
    i_13_387_77_0, i_13_387_80_0, i_13_387_153_0, i_13_387_412_0,
    i_13_387_611_0, i_13_387_629_0, i_13_387_661_0, i_13_387_662_0,
    i_13_387_664_0, i_13_387_674_0, i_13_387_683_0, i_13_387_686_0,
    i_13_387_716_0, i_13_387_851_0, i_13_387_854_0, i_13_387_940_0,
    i_13_387_1060_0, i_13_387_1071_0, i_13_387_1076_0, i_13_387_1101_0,
    i_13_387_1105_0, i_13_387_1106_0, i_13_387_1133_0, i_13_387_1151_0,
    i_13_387_1188_0, i_13_387_1224_0, i_13_387_1228_0, i_13_387_1229_0,
    i_13_387_1232_0, i_13_387_1244_0, i_13_387_1256_0, i_13_387_1318_0,
    i_13_387_1345_0, i_13_387_1484_0, i_13_387_1733_0, i_13_387_1765_0,
    i_13_387_1766_0, i_13_387_1768_0, i_13_387_1787_0, i_13_387_1799_0,
    i_13_387_1892_0, i_13_387_1927_0, i_13_387_1962_0, i_13_387_2005_0,
    i_13_387_2023_0, i_13_387_2024_0, i_13_387_2026_0, i_13_387_2212_0,
    i_13_387_2284_0, i_13_387_2288_0, i_13_387_2434_0, i_13_387_2518_0,
    i_13_387_2582_0, i_13_387_2852_0, i_13_387_2903_0, i_13_387_2975_0,
    i_13_387_2987_0, i_13_387_3010_0, i_13_387_3013_0, i_13_387_3027_0,
    i_13_387_3032_0, i_13_387_3050_0, i_13_387_3064_0, i_13_387_3122_0,
    i_13_387_3261_0, i_13_387_3355_0, i_13_387_3356_0, i_13_387_3487_0,
    i_13_387_3539_0, i_13_387_3542_0, i_13_387_3573_0, i_13_387_3574_0,
    i_13_387_3731_0, i_13_387_3734_0, i_13_387_3755_0, i_13_387_3866_0,
    i_13_387_3869_0, i_13_387_3928_0, i_13_387_3978_0, i_13_387_4166_0,
    i_13_387_4212_0, i_13_387_4255_0, i_13_387_4256_0, i_13_387_4302_0,
    i_13_387_4322_0, i_13_387_4336_0, i_13_387_4343_0, i_13_387_4372_0,
    i_13_387_4373_0, i_13_387_4382_0, i_13_387_4450_0, i_13_387_4514_0,
    i_13_387_4516_0, i_13_387_4598_0, i_13_387_4606_0, i_13_387_4607_0;
  output o_13_387_0_0;
  assign o_13_387_0_0 = ~(~i_13_387_940_0 | (~i_13_387_71_0 & ~i_13_387_2987_0));
endmodule



// Benchmark "kernel_13_388" written by ABC on Sun Jul 19 10:50:47 2020

module kernel_13_388 ( 
    i_13_388_31_0, i_13_388_53_0, i_13_388_103_0, i_13_388_125_0,
    i_13_388_142_0, i_13_388_143_0, i_13_388_241_0, i_13_388_251_0,
    i_13_388_278_0, i_13_388_322_0, i_13_388_340_0, i_13_388_449_0,
    i_13_388_508_0, i_13_388_575_0, i_13_388_619_0, i_13_388_620_0,
    i_13_388_728_0, i_13_388_781_0, i_13_388_850_0, i_13_388_980_0,
    i_13_388_1079_0, i_13_388_1084_0, i_13_388_1250_0, i_13_388_1265_0,
    i_13_388_1309_0, i_13_388_1364_0, i_13_388_1402_0, i_13_388_1436_0,
    i_13_388_1498_0, i_13_388_1502_0, i_13_388_1529_0, i_13_388_1566_0,
    i_13_388_1609_0, i_13_388_1636_0, i_13_388_1637_0, i_13_388_1726_0,
    i_13_388_1735_0, i_13_388_1796_0, i_13_388_1817_0, i_13_388_1907_0,
    i_13_388_1913_0, i_13_388_1921_0, i_13_388_1930_0, i_13_388_1989_0,
    i_13_388_2097_0, i_13_388_2120_0, i_13_388_2294_0, i_13_388_2358_0,
    i_13_388_2545_0, i_13_388_2564_0, i_13_388_2570_0, i_13_388_2596_0,
    i_13_388_2709_0, i_13_388_2768_0, i_13_388_2788_0, i_13_388_2789_0,
    i_13_388_2844_0, i_13_388_2848_0, i_13_388_2959_0, i_13_388_3004_0,
    i_13_388_3070_0, i_13_388_3130_0, i_13_388_3131_0, i_13_388_3167_0,
    i_13_388_3220_0, i_13_388_3221_0, i_13_388_3253_0, i_13_388_3374_0,
    i_13_388_3383_0, i_13_388_3411_0, i_13_388_3416_0, i_13_388_3418_0,
    i_13_388_3419_0, i_13_388_3447_0, i_13_388_3527_0, i_13_388_3554_0,
    i_13_388_3581_0, i_13_388_3641_0, i_13_388_3643_0, i_13_388_3662_0,
    i_13_388_3688_0, i_13_388_3740_0, i_13_388_3788_0, i_13_388_3847_0,
    i_13_388_3856_0, i_13_388_3874_0, i_13_388_3875_0, i_13_388_3914_0,
    i_13_388_4012_0, i_13_388_4057_0, i_13_388_4084_0, i_13_388_4090_0,
    i_13_388_4091_0, i_13_388_4108_0, i_13_388_4171_0, i_13_388_4271_0,
    i_13_388_4364_0, i_13_388_4391_0, i_13_388_4415_0, i_13_388_4526_0,
    o_13_388_0_0  );
  input  i_13_388_31_0, i_13_388_53_0, i_13_388_103_0, i_13_388_125_0,
    i_13_388_142_0, i_13_388_143_0, i_13_388_241_0, i_13_388_251_0,
    i_13_388_278_0, i_13_388_322_0, i_13_388_340_0, i_13_388_449_0,
    i_13_388_508_0, i_13_388_575_0, i_13_388_619_0, i_13_388_620_0,
    i_13_388_728_0, i_13_388_781_0, i_13_388_850_0, i_13_388_980_0,
    i_13_388_1079_0, i_13_388_1084_0, i_13_388_1250_0, i_13_388_1265_0,
    i_13_388_1309_0, i_13_388_1364_0, i_13_388_1402_0, i_13_388_1436_0,
    i_13_388_1498_0, i_13_388_1502_0, i_13_388_1529_0, i_13_388_1566_0,
    i_13_388_1609_0, i_13_388_1636_0, i_13_388_1637_0, i_13_388_1726_0,
    i_13_388_1735_0, i_13_388_1796_0, i_13_388_1817_0, i_13_388_1907_0,
    i_13_388_1913_0, i_13_388_1921_0, i_13_388_1930_0, i_13_388_1989_0,
    i_13_388_2097_0, i_13_388_2120_0, i_13_388_2294_0, i_13_388_2358_0,
    i_13_388_2545_0, i_13_388_2564_0, i_13_388_2570_0, i_13_388_2596_0,
    i_13_388_2709_0, i_13_388_2768_0, i_13_388_2788_0, i_13_388_2789_0,
    i_13_388_2844_0, i_13_388_2848_0, i_13_388_2959_0, i_13_388_3004_0,
    i_13_388_3070_0, i_13_388_3130_0, i_13_388_3131_0, i_13_388_3167_0,
    i_13_388_3220_0, i_13_388_3221_0, i_13_388_3253_0, i_13_388_3374_0,
    i_13_388_3383_0, i_13_388_3411_0, i_13_388_3416_0, i_13_388_3418_0,
    i_13_388_3419_0, i_13_388_3447_0, i_13_388_3527_0, i_13_388_3554_0,
    i_13_388_3581_0, i_13_388_3641_0, i_13_388_3643_0, i_13_388_3662_0,
    i_13_388_3688_0, i_13_388_3740_0, i_13_388_3788_0, i_13_388_3847_0,
    i_13_388_3856_0, i_13_388_3874_0, i_13_388_3875_0, i_13_388_3914_0,
    i_13_388_4012_0, i_13_388_4057_0, i_13_388_4084_0, i_13_388_4090_0,
    i_13_388_4091_0, i_13_388_4108_0, i_13_388_4171_0, i_13_388_4271_0,
    i_13_388_4364_0, i_13_388_4391_0, i_13_388_4415_0, i_13_388_4526_0;
  output o_13_388_0_0;
  assign o_13_388_0_0 = ~((i_13_388_31_0 & ~i_13_388_3554_0) | (~i_13_388_620_0 & ~i_13_388_3221_0));
endmodule



// Benchmark "kernel_13_389" written by ABC on Sun Jul 19 10:50:48 2020

module kernel_13_389 ( 
    i_13_389_28_0, i_13_389_37_0, i_13_389_48_0, i_13_389_63_0,
    i_13_389_64_0, i_13_389_65_0, i_13_389_198_0, i_13_389_352_0,
    i_13_389_354_0, i_13_389_361_0, i_13_389_378_0, i_13_389_462_0,
    i_13_389_588_0, i_13_389_668_0, i_13_389_685_0, i_13_389_694_0,
    i_13_389_712_0, i_13_389_756_0, i_13_389_823_0, i_13_389_828_0,
    i_13_389_838_0, i_13_389_859_0, i_13_389_909_0, i_13_389_1117_0,
    i_13_389_1137_0, i_13_389_1296_0, i_13_389_1304_0, i_13_389_1306_0,
    i_13_389_1309_0, i_13_389_1345_0, i_13_389_1372_0, i_13_389_1396_0,
    i_13_389_1405_0, i_13_389_1503_0, i_13_389_1504_0, i_13_389_1517_0,
    i_13_389_1543_0, i_13_389_1557_0, i_13_389_1593_0, i_13_389_1594_0,
    i_13_389_1638_0, i_13_389_1639_0, i_13_389_1669_0, i_13_389_1710_0,
    i_13_389_1732_0, i_13_389_1740_0, i_13_389_1858_0, i_13_389_1927_0,
    i_13_389_2056_0, i_13_389_2071_0, i_13_389_2124_0, i_13_389_2142_0,
    i_13_389_2189_0, i_13_389_2281_0, i_13_389_2317_0, i_13_389_2377_0,
    i_13_389_2395_0, i_13_389_2461_0, i_13_389_2478_0, i_13_389_2511_0,
    i_13_389_2539_0, i_13_389_2691_0, i_13_389_2718_0, i_13_389_2719_0,
    i_13_389_2720_0, i_13_389_2912_0, i_13_389_3052_0, i_13_389_3060_0,
    i_13_389_3109_0, i_13_389_3163_0, i_13_389_3172_0, i_13_389_3388_0,
    i_13_389_3414_0, i_13_389_3532_0, i_13_389_3594_0, i_13_389_3595_0,
    i_13_389_3609_0, i_13_389_3618_0, i_13_389_3637_0, i_13_389_3766_0,
    i_13_389_3863_0, i_13_389_3910_0, i_13_389_3916_0, i_13_389_3924_0,
    i_13_389_4032_0, i_13_389_4033_0, i_13_389_4036_0, i_13_389_4063_0,
    i_13_389_4213_0, i_13_389_4262_0, i_13_389_4302_0, i_13_389_4307_0,
    i_13_389_4312_0, i_13_389_4315_0, i_13_389_4330_0, i_13_389_4396_0,
    i_13_389_4429_0, i_13_389_4430_0, i_13_389_4477_0, i_13_389_4591_0,
    o_13_389_0_0  );
  input  i_13_389_28_0, i_13_389_37_0, i_13_389_48_0, i_13_389_63_0,
    i_13_389_64_0, i_13_389_65_0, i_13_389_198_0, i_13_389_352_0,
    i_13_389_354_0, i_13_389_361_0, i_13_389_378_0, i_13_389_462_0,
    i_13_389_588_0, i_13_389_668_0, i_13_389_685_0, i_13_389_694_0,
    i_13_389_712_0, i_13_389_756_0, i_13_389_823_0, i_13_389_828_0,
    i_13_389_838_0, i_13_389_859_0, i_13_389_909_0, i_13_389_1117_0,
    i_13_389_1137_0, i_13_389_1296_0, i_13_389_1304_0, i_13_389_1306_0,
    i_13_389_1309_0, i_13_389_1345_0, i_13_389_1372_0, i_13_389_1396_0,
    i_13_389_1405_0, i_13_389_1503_0, i_13_389_1504_0, i_13_389_1517_0,
    i_13_389_1543_0, i_13_389_1557_0, i_13_389_1593_0, i_13_389_1594_0,
    i_13_389_1638_0, i_13_389_1639_0, i_13_389_1669_0, i_13_389_1710_0,
    i_13_389_1732_0, i_13_389_1740_0, i_13_389_1858_0, i_13_389_1927_0,
    i_13_389_2056_0, i_13_389_2071_0, i_13_389_2124_0, i_13_389_2142_0,
    i_13_389_2189_0, i_13_389_2281_0, i_13_389_2317_0, i_13_389_2377_0,
    i_13_389_2395_0, i_13_389_2461_0, i_13_389_2478_0, i_13_389_2511_0,
    i_13_389_2539_0, i_13_389_2691_0, i_13_389_2718_0, i_13_389_2719_0,
    i_13_389_2720_0, i_13_389_2912_0, i_13_389_3052_0, i_13_389_3060_0,
    i_13_389_3109_0, i_13_389_3163_0, i_13_389_3172_0, i_13_389_3388_0,
    i_13_389_3414_0, i_13_389_3532_0, i_13_389_3594_0, i_13_389_3595_0,
    i_13_389_3609_0, i_13_389_3618_0, i_13_389_3637_0, i_13_389_3766_0,
    i_13_389_3863_0, i_13_389_3910_0, i_13_389_3916_0, i_13_389_3924_0,
    i_13_389_4032_0, i_13_389_4033_0, i_13_389_4036_0, i_13_389_4063_0,
    i_13_389_4213_0, i_13_389_4262_0, i_13_389_4302_0, i_13_389_4307_0,
    i_13_389_4312_0, i_13_389_4315_0, i_13_389_4330_0, i_13_389_4396_0,
    i_13_389_4429_0, i_13_389_4430_0, i_13_389_4477_0, i_13_389_4591_0;
  output o_13_389_0_0;
  assign o_13_389_0_0 = ~((~i_13_389_65_0 & ((~i_13_389_1309_0 & ~i_13_389_3618_0) | (~i_13_389_63_0 & ~i_13_389_828_0 & ~i_13_389_2056_0 & ~i_13_389_4330_0 & ~i_13_389_4429_0))) | (~i_13_389_4032_0 & ((i_13_389_859_0 & ~i_13_389_4312_0) | (~i_13_389_685_0 & ~i_13_389_4262_0 & ~i_13_389_4330_0))) | (~i_13_389_4429_0 & ((~i_13_389_4302_0 & (~i_13_389_1639_0 | ~i_13_389_4213_0)) | (i_13_389_3109_0 & i_13_389_4312_0))) | (~i_13_389_694_0 & ~i_13_389_1594_0 & ~i_13_389_2691_0));
endmodule



// Benchmark "kernel_13_390" written by ABC on Sun Jul 19 10:50:48 2020

module kernel_13_390 ( 
    i_13_390_72_0, i_13_390_121_0, i_13_390_139_0, i_13_390_165_0,
    i_13_390_173_0, i_13_390_175_0, i_13_390_311_0, i_13_390_523_0,
    i_13_390_526_0, i_13_390_532_0, i_13_390_535_0, i_13_390_796_0,
    i_13_390_798_0, i_13_390_811_0, i_13_390_814_0, i_13_390_848_0,
    i_13_390_850_0, i_13_390_851_0, i_13_390_958_0, i_13_390_985_0,
    i_13_390_1073_0, i_13_390_1079_0, i_13_390_1225_0, i_13_390_1228_0,
    i_13_390_1258_0, i_13_390_1411_0, i_13_390_1468_0, i_13_390_1471_0,
    i_13_390_1497_0, i_13_390_1549_0, i_13_390_1550_0, i_13_390_1552_0,
    i_13_390_1624_0, i_13_390_1750_0, i_13_390_1803_0, i_13_390_1831_0,
    i_13_390_1846_0, i_13_390_1858_0, i_13_390_1922_0, i_13_390_1925_0,
    i_13_390_1957_0, i_13_390_2124_0, i_13_390_2133_0, i_13_390_2203_0,
    i_13_390_2303_0, i_13_390_2408_0, i_13_390_2458_0, i_13_390_2570_0,
    i_13_390_2614_0, i_13_390_2785_0, i_13_390_2884_0, i_13_390_2918_0,
    i_13_390_3007_0, i_13_390_3010_0, i_13_390_3037_0, i_13_390_3061_0,
    i_13_390_3100_0, i_13_390_3108_0, i_13_390_3109_0, i_13_390_3268_0,
    i_13_390_3271_0, i_13_390_3274_0, i_13_390_3342_0, i_13_390_3396_0,
    i_13_390_3402_0, i_13_390_3409_0, i_13_390_3464_0, i_13_390_3469_0,
    i_13_390_3539_0, i_13_390_3541_0, i_13_390_3568_0, i_13_390_3604_0,
    i_13_390_3663_0, i_13_390_3666_0, i_13_390_3727_0, i_13_390_3728_0,
    i_13_390_3729_0, i_13_390_3838_0, i_13_390_3856_0, i_13_390_3869_0,
    i_13_390_3907_0, i_13_390_3909_0, i_13_390_3911_0, i_13_390_3928_0,
    i_13_390_4018_0, i_13_390_4054_0, i_13_390_4099_0, i_13_390_4249_0,
    i_13_390_4251_0, i_13_390_4252_0, i_13_390_4253_0, i_13_390_4255_0,
    i_13_390_4256_0, i_13_390_4258_0, i_13_390_4259_0, i_13_390_4277_0,
    i_13_390_4375_0, i_13_390_4376_0, i_13_390_4540_0, i_13_390_4557_0,
    o_13_390_0_0  );
  input  i_13_390_72_0, i_13_390_121_0, i_13_390_139_0, i_13_390_165_0,
    i_13_390_173_0, i_13_390_175_0, i_13_390_311_0, i_13_390_523_0,
    i_13_390_526_0, i_13_390_532_0, i_13_390_535_0, i_13_390_796_0,
    i_13_390_798_0, i_13_390_811_0, i_13_390_814_0, i_13_390_848_0,
    i_13_390_850_0, i_13_390_851_0, i_13_390_958_0, i_13_390_985_0,
    i_13_390_1073_0, i_13_390_1079_0, i_13_390_1225_0, i_13_390_1228_0,
    i_13_390_1258_0, i_13_390_1411_0, i_13_390_1468_0, i_13_390_1471_0,
    i_13_390_1497_0, i_13_390_1549_0, i_13_390_1550_0, i_13_390_1552_0,
    i_13_390_1624_0, i_13_390_1750_0, i_13_390_1803_0, i_13_390_1831_0,
    i_13_390_1846_0, i_13_390_1858_0, i_13_390_1922_0, i_13_390_1925_0,
    i_13_390_1957_0, i_13_390_2124_0, i_13_390_2133_0, i_13_390_2203_0,
    i_13_390_2303_0, i_13_390_2408_0, i_13_390_2458_0, i_13_390_2570_0,
    i_13_390_2614_0, i_13_390_2785_0, i_13_390_2884_0, i_13_390_2918_0,
    i_13_390_3007_0, i_13_390_3010_0, i_13_390_3037_0, i_13_390_3061_0,
    i_13_390_3100_0, i_13_390_3108_0, i_13_390_3109_0, i_13_390_3268_0,
    i_13_390_3271_0, i_13_390_3274_0, i_13_390_3342_0, i_13_390_3396_0,
    i_13_390_3402_0, i_13_390_3409_0, i_13_390_3464_0, i_13_390_3469_0,
    i_13_390_3539_0, i_13_390_3541_0, i_13_390_3568_0, i_13_390_3604_0,
    i_13_390_3663_0, i_13_390_3666_0, i_13_390_3727_0, i_13_390_3728_0,
    i_13_390_3729_0, i_13_390_3838_0, i_13_390_3856_0, i_13_390_3869_0,
    i_13_390_3907_0, i_13_390_3909_0, i_13_390_3911_0, i_13_390_3928_0,
    i_13_390_4018_0, i_13_390_4054_0, i_13_390_4099_0, i_13_390_4249_0,
    i_13_390_4251_0, i_13_390_4252_0, i_13_390_4253_0, i_13_390_4255_0,
    i_13_390_4256_0, i_13_390_4258_0, i_13_390_4259_0, i_13_390_4277_0,
    i_13_390_4375_0, i_13_390_4376_0, i_13_390_4540_0, i_13_390_4557_0;
  output o_13_390_0_0;
  assign o_13_390_0_0 = ~((i_13_390_1471_0 & ~i_13_390_3907_0 & ((~i_13_390_175_0 & i_13_390_1922_0 & ~i_13_390_3464_0) | (i_13_390_3037_0 & ~i_13_390_3342_0 & ~i_13_390_3911_0 & ~i_13_390_4253_0))) | (~i_13_390_1803_0 & ((~i_13_390_814_0 & ~i_13_390_3010_0 & ~i_13_390_3109_0 & ~i_13_390_3856_0 & i_13_390_3928_0 & ~i_13_390_4249_0) | (i_13_390_139_0 & ~i_13_390_811_0 & ~i_13_390_1079_0 & ~i_13_390_1552_0 & ~i_13_390_1957_0 & ~i_13_390_3108_0 & ~i_13_390_3727_0 & ~i_13_390_4258_0))) | (~i_13_390_173_0 & i_13_390_1624_0 & ~i_13_390_1846_0 & ~i_13_390_2408_0 & ~i_13_390_3010_0 & ~i_13_390_3396_0 & ~i_13_390_3541_0 & ~i_13_390_3909_0));
endmodule



// Benchmark "kernel_13_391" written by ABC on Sun Jul 19 10:50:49 2020

module kernel_13_391 ( 
    i_13_391_259_0, i_13_391_311_0, i_13_391_328_0, i_13_391_329_0,
    i_13_391_562_0, i_13_391_583_0, i_13_391_611_0, i_13_391_628_0,
    i_13_391_629_0, i_13_391_823_0, i_13_391_826_0, i_13_391_862_0,
    i_13_391_863_0, i_13_391_894_0, i_13_391_1024_0, i_13_391_1025_0,
    i_13_391_1033_0, i_13_391_1076_0, i_13_391_1096_0, i_13_391_1097_0,
    i_13_391_1228_0, i_13_391_1229_0, i_13_391_1232_0, i_13_391_1256_0,
    i_13_391_1258_0, i_13_391_1259_0, i_13_391_1320_0, i_13_391_1321_0,
    i_13_391_1327_0, i_13_391_1384_0, i_13_391_1439_0, i_13_391_1483_0,
    i_13_391_1484_0, i_13_391_1490_0, i_13_391_1492_0, i_13_391_1679_0,
    i_13_391_1691_0, i_13_391_1780_0, i_13_391_1781_0, i_13_391_1789_0,
    i_13_391_1858_0, i_13_391_1859_0, i_13_391_1861_0, i_13_391_1862_0,
    i_13_391_1886_0, i_13_391_1889_0, i_13_391_2030_0, i_13_391_2056_0,
    i_13_391_2123_0, i_13_391_2150_0, i_13_391_2230_0, i_13_391_2312_0,
    i_13_391_2461_0, i_13_391_2465_0, i_13_391_2509_0, i_13_391_2510_0,
    i_13_391_2570_0, i_13_391_2851_0, i_13_391_2852_0, i_13_391_2875_0,
    i_13_391_2876_0, i_13_391_2977_0, i_13_391_3001_0, i_13_391_3064_0,
    i_13_391_3094_0, i_13_391_3100_0, i_13_391_3101_0, i_13_391_3122_0,
    i_13_391_3157_0, i_13_391_3173_0, i_13_391_3176_0, i_13_391_3211_0,
    i_13_391_3432_0, i_13_391_3433_0, i_13_391_3460_0, i_13_391_3479_0,
    i_13_391_3488_0, i_13_391_3506_0, i_13_391_3524_0, i_13_391_3535_0,
    i_13_391_3536_0, i_13_391_3542_0, i_13_391_3545_0, i_13_391_3563_0,
    i_13_391_3707_0, i_13_391_3785_0, i_13_391_3835_0, i_13_391_3857_0,
    i_13_391_3895_0, i_13_391_3911_0, i_13_391_3914_0, i_13_391_4036_0,
    i_13_391_4207_0, i_13_391_4255_0, i_13_391_4342_0, i_13_391_4373_0,
    i_13_391_4378_0, i_13_391_4381_0, i_13_391_4382_0, i_13_391_4594_0,
    o_13_391_0_0  );
  input  i_13_391_259_0, i_13_391_311_0, i_13_391_328_0, i_13_391_329_0,
    i_13_391_562_0, i_13_391_583_0, i_13_391_611_0, i_13_391_628_0,
    i_13_391_629_0, i_13_391_823_0, i_13_391_826_0, i_13_391_862_0,
    i_13_391_863_0, i_13_391_894_0, i_13_391_1024_0, i_13_391_1025_0,
    i_13_391_1033_0, i_13_391_1076_0, i_13_391_1096_0, i_13_391_1097_0,
    i_13_391_1228_0, i_13_391_1229_0, i_13_391_1232_0, i_13_391_1256_0,
    i_13_391_1258_0, i_13_391_1259_0, i_13_391_1320_0, i_13_391_1321_0,
    i_13_391_1327_0, i_13_391_1384_0, i_13_391_1439_0, i_13_391_1483_0,
    i_13_391_1484_0, i_13_391_1490_0, i_13_391_1492_0, i_13_391_1679_0,
    i_13_391_1691_0, i_13_391_1780_0, i_13_391_1781_0, i_13_391_1789_0,
    i_13_391_1858_0, i_13_391_1859_0, i_13_391_1861_0, i_13_391_1862_0,
    i_13_391_1886_0, i_13_391_1889_0, i_13_391_2030_0, i_13_391_2056_0,
    i_13_391_2123_0, i_13_391_2150_0, i_13_391_2230_0, i_13_391_2312_0,
    i_13_391_2461_0, i_13_391_2465_0, i_13_391_2509_0, i_13_391_2510_0,
    i_13_391_2570_0, i_13_391_2851_0, i_13_391_2852_0, i_13_391_2875_0,
    i_13_391_2876_0, i_13_391_2977_0, i_13_391_3001_0, i_13_391_3064_0,
    i_13_391_3094_0, i_13_391_3100_0, i_13_391_3101_0, i_13_391_3122_0,
    i_13_391_3157_0, i_13_391_3173_0, i_13_391_3176_0, i_13_391_3211_0,
    i_13_391_3432_0, i_13_391_3433_0, i_13_391_3460_0, i_13_391_3479_0,
    i_13_391_3488_0, i_13_391_3506_0, i_13_391_3524_0, i_13_391_3535_0,
    i_13_391_3536_0, i_13_391_3542_0, i_13_391_3545_0, i_13_391_3563_0,
    i_13_391_3707_0, i_13_391_3785_0, i_13_391_3835_0, i_13_391_3857_0,
    i_13_391_3895_0, i_13_391_3911_0, i_13_391_3914_0, i_13_391_4036_0,
    i_13_391_4207_0, i_13_391_4255_0, i_13_391_4342_0, i_13_391_4373_0,
    i_13_391_4378_0, i_13_391_4381_0, i_13_391_4382_0, i_13_391_4594_0;
  output o_13_391_0_0;
  assign o_13_391_0_0 = ~((~i_13_391_329_0 & ((~i_13_391_1232_0 & ~i_13_391_2150_0 & ~i_13_391_3460_0) | (~i_13_391_3542_0 & ~i_13_391_4381_0))) | (~i_13_391_862_0 & i_13_391_3460_0 & ~i_13_391_4373_0));
endmodule



// Benchmark "kernel_13_392" written by ABC on Sun Jul 19 10:50:50 2020

module kernel_13_392 ( 
    i_13_392_30_0, i_13_392_67_0, i_13_392_72_0, i_13_392_73_0,
    i_13_392_103_0, i_13_392_108_0, i_13_392_255_0, i_13_392_282_0,
    i_13_392_297_0, i_13_392_354_0, i_13_392_355_0, i_13_392_358_0,
    i_13_392_360_0, i_13_392_369_0, i_13_392_373_0, i_13_392_396_0,
    i_13_392_468_0, i_13_392_523_0, i_13_392_588_0, i_13_392_603_0,
    i_13_392_639_0, i_13_392_666_0, i_13_392_667_0, i_13_392_741_0,
    i_13_392_742_0, i_13_392_759_0, i_13_392_828_0, i_13_392_838_0,
    i_13_392_945_0, i_13_392_946_0, i_13_392_975_0, i_13_392_1084_0,
    i_13_392_1209_0, i_13_392_1304_0, i_13_392_1344_0, i_13_392_1504_0,
    i_13_392_1620_0, i_13_392_1683_0, i_13_392_1693_0, i_13_392_1774_0,
    i_13_392_1777_0, i_13_392_1947_0, i_13_392_1999_0, i_13_392_2055_0,
    i_13_392_2056_0, i_13_392_2169_0, i_13_392_2181_0, i_13_392_2280_0,
    i_13_392_2281_0, i_13_392_2298_0, i_13_392_2348_0, i_13_392_2350_0,
    i_13_392_2430_0, i_13_392_2431_0, i_13_392_2469_0, i_13_392_2511_0,
    i_13_392_2512_0, i_13_392_2539_0, i_13_392_2613_0, i_13_392_2614_0,
    i_13_392_2691_0, i_13_392_2692_0, i_13_392_2721_0, i_13_392_2880_0,
    i_13_392_2881_0, i_13_392_2907_0, i_13_392_2916_0, i_13_392_3007_0,
    i_13_392_3385_0, i_13_392_3387_0, i_13_392_3528_0, i_13_392_3558_0,
    i_13_392_3594_0, i_13_392_3595_0, i_13_392_3599_0, i_13_392_3613_0,
    i_13_392_3618_0, i_13_392_3619_0, i_13_392_3631_0, i_13_392_3634_0,
    i_13_392_3636_0, i_13_392_3685_0, i_13_392_3726_0, i_13_392_3978_0,
    i_13_392_3987_0, i_13_392_4041_0, i_13_392_4117_0, i_13_392_4123_0,
    i_13_392_4188_0, i_13_392_4202_0, i_13_392_4233_0, i_13_392_4260_0,
    i_13_392_4329_0, i_13_392_4330_0, i_13_392_4365_0, i_13_392_4366_0,
    i_13_392_4410_0, i_13_392_4428_0, i_13_392_4429_0, i_13_392_4450_0,
    o_13_392_0_0  );
  input  i_13_392_30_0, i_13_392_67_0, i_13_392_72_0, i_13_392_73_0,
    i_13_392_103_0, i_13_392_108_0, i_13_392_255_0, i_13_392_282_0,
    i_13_392_297_0, i_13_392_354_0, i_13_392_355_0, i_13_392_358_0,
    i_13_392_360_0, i_13_392_369_0, i_13_392_373_0, i_13_392_396_0,
    i_13_392_468_0, i_13_392_523_0, i_13_392_588_0, i_13_392_603_0,
    i_13_392_639_0, i_13_392_666_0, i_13_392_667_0, i_13_392_741_0,
    i_13_392_742_0, i_13_392_759_0, i_13_392_828_0, i_13_392_838_0,
    i_13_392_945_0, i_13_392_946_0, i_13_392_975_0, i_13_392_1084_0,
    i_13_392_1209_0, i_13_392_1304_0, i_13_392_1344_0, i_13_392_1504_0,
    i_13_392_1620_0, i_13_392_1683_0, i_13_392_1693_0, i_13_392_1774_0,
    i_13_392_1777_0, i_13_392_1947_0, i_13_392_1999_0, i_13_392_2055_0,
    i_13_392_2056_0, i_13_392_2169_0, i_13_392_2181_0, i_13_392_2280_0,
    i_13_392_2281_0, i_13_392_2298_0, i_13_392_2348_0, i_13_392_2350_0,
    i_13_392_2430_0, i_13_392_2431_0, i_13_392_2469_0, i_13_392_2511_0,
    i_13_392_2512_0, i_13_392_2539_0, i_13_392_2613_0, i_13_392_2614_0,
    i_13_392_2691_0, i_13_392_2692_0, i_13_392_2721_0, i_13_392_2880_0,
    i_13_392_2881_0, i_13_392_2907_0, i_13_392_2916_0, i_13_392_3007_0,
    i_13_392_3385_0, i_13_392_3387_0, i_13_392_3528_0, i_13_392_3558_0,
    i_13_392_3594_0, i_13_392_3595_0, i_13_392_3599_0, i_13_392_3613_0,
    i_13_392_3618_0, i_13_392_3619_0, i_13_392_3631_0, i_13_392_3634_0,
    i_13_392_3636_0, i_13_392_3685_0, i_13_392_3726_0, i_13_392_3978_0,
    i_13_392_3987_0, i_13_392_4041_0, i_13_392_4117_0, i_13_392_4123_0,
    i_13_392_4188_0, i_13_392_4202_0, i_13_392_4233_0, i_13_392_4260_0,
    i_13_392_4329_0, i_13_392_4330_0, i_13_392_4365_0, i_13_392_4366_0,
    i_13_392_4410_0, i_13_392_4428_0, i_13_392_4429_0, i_13_392_4450_0;
  output o_13_392_0_0;
  assign o_13_392_0_0 = ~((~i_13_392_4429_0 & (~i_13_392_67_0 | (~i_13_392_103_0 & ~i_13_392_3685_0))) | (~i_13_392_1344_0 & ~i_13_392_3387_0) | (~i_13_392_468_0 & ~i_13_392_4260_0));
endmodule



// Benchmark "kernel_13_393" written by ABC on Sun Jul 19 10:50:51 2020

module kernel_13_393 ( 
    i_13_393_19_0, i_13_393_73_0, i_13_393_94_0, i_13_393_355_0,
    i_13_393_443_0, i_13_393_530_0, i_13_393_628_0, i_13_393_695_0,
    i_13_393_697_0, i_13_393_706_0, i_13_393_831_0, i_13_393_886_0,
    i_13_393_1022_0, i_13_393_1066_0, i_13_393_1072_0, i_13_393_1073_0,
    i_13_393_1100_0, i_13_393_1112_0, i_13_393_1208_0, i_13_393_1210_0,
    i_13_393_1217_0, i_13_393_1258_0, i_13_393_1286_0, i_13_393_1337_0,
    i_13_393_1399_0, i_13_393_1419_0, i_13_393_1424_0, i_13_393_1427_0,
    i_13_393_1491_0, i_13_393_1499_0, i_13_393_1522_0, i_13_393_1658_0,
    i_13_393_1732_0, i_13_393_1774_0, i_13_393_1775_0, i_13_393_1837_0,
    i_13_393_1960_0, i_13_393_1966_0, i_13_393_2006_0, i_13_393_2020_0,
    i_13_393_2021_0, i_13_393_2029_0, i_13_393_2045_0, i_13_393_2144_0,
    i_13_393_2209_0, i_13_393_2232_0, i_13_393_2281_0, i_13_393_2297_0,
    i_13_393_2347_0, i_13_393_2425_0, i_13_393_2443_0, i_13_393_2444_0,
    i_13_393_2446_0, i_13_393_2449_0, i_13_393_2453_0, i_13_393_2454_0,
    i_13_393_2512_0, i_13_393_2515_0, i_13_393_2555_0, i_13_393_2693_0,
    i_13_393_2719_0, i_13_393_2822_0, i_13_393_2884_0, i_13_393_2896_0,
    i_13_393_3037_0, i_13_393_3074_0, i_13_393_3307_0, i_13_393_3370_0,
    i_13_393_3416_0, i_13_393_3442_0, i_13_393_3547_0, i_13_393_3568_0,
    i_13_393_3578_0, i_13_393_3579_0, i_13_393_3598_0, i_13_393_3620_0,
    i_13_393_3634_0, i_13_393_3682_0, i_13_393_3740_0, i_13_393_3756_0,
    i_13_393_3806_0, i_13_393_3958_0, i_13_393_3967_0, i_13_393_3989_0,
    i_13_393_4018_0, i_13_393_4039_0, i_13_393_4208_0, i_13_393_4263_0,
    i_13_393_4272_0, i_13_393_4330_0, i_13_393_4332_0, i_13_393_4333_0,
    i_13_393_4379_0, i_13_393_4430_0, i_13_393_4453_0, i_13_393_4510_0,
    i_13_393_4513_0, i_13_393_4594_0, i_13_393_4596_0, i_13_393_4604_0,
    o_13_393_0_0  );
  input  i_13_393_19_0, i_13_393_73_0, i_13_393_94_0, i_13_393_355_0,
    i_13_393_443_0, i_13_393_530_0, i_13_393_628_0, i_13_393_695_0,
    i_13_393_697_0, i_13_393_706_0, i_13_393_831_0, i_13_393_886_0,
    i_13_393_1022_0, i_13_393_1066_0, i_13_393_1072_0, i_13_393_1073_0,
    i_13_393_1100_0, i_13_393_1112_0, i_13_393_1208_0, i_13_393_1210_0,
    i_13_393_1217_0, i_13_393_1258_0, i_13_393_1286_0, i_13_393_1337_0,
    i_13_393_1399_0, i_13_393_1419_0, i_13_393_1424_0, i_13_393_1427_0,
    i_13_393_1491_0, i_13_393_1499_0, i_13_393_1522_0, i_13_393_1658_0,
    i_13_393_1732_0, i_13_393_1774_0, i_13_393_1775_0, i_13_393_1837_0,
    i_13_393_1960_0, i_13_393_1966_0, i_13_393_2006_0, i_13_393_2020_0,
    i_13_393_2021_0, i_13_393_2029_0, i_13_393_2045_0, i_13_393_2144_0,
    i_13_393_2209_0, i_13_393_2232_0, i_13_393_2281_0, i_13_393_2297_0,
    i_13_393_2347_0, i_13_393_2425_0, i_13_393_2443_0, i_13_393_2444_0,
    i_13_393_2446_0, i_13_393_2449_0, i_13_393_2453_0, i_13_393_2454_0,
    i_13_393_2512_0, i_13_393_2515_0, i_13_393_2555_0, i_13_393_2693_0,
    i_13_393_2719_0, i_13_393_2822_0, i_13_393_2884_0, i_13_393_2896_0,
    i_13_393_3037_0, i_13_393_3074_0, i_13_393_3307_0, i_13_393_3370_0,
    i_13_393_3416_0, i_13_393_3442_0, i_13_393_3547_0, i_13_393_3568_0,
    i_13_393_3578_0, i_13_393_3579_0, i_13_393_3598_0, i_13_393_3620_0,
    i_13_393_3634_0, i_13_393_3682_0, i_13_393_3740_0, i_13_393_3756_0,
    i_13_393_3806_0, i_13_393_3958_0, i_13_393_3967_0, i_13_393_3989_0,
    i_13_393_4018_0, i_13_393_4039_0, i_13_393_4208_0, i_13_393_4263_0,
    i_13_393_4272_0, i_13_393_4330_0, i_13_393_4332_0, i_13_393_4333_0,
    i_13_393_4379_0, i_13_393_4430_0, i_13_393_4453_0, i_13_393_4510_0,
    i_13_393_4513_0, i_13_393_4594_0, i_13_393_4596_0, i_13_393_4604_0;
  output o_13_393_0_0;
  assign o_13_393_0_0 = 0;
endmodule



// Benchmark "kernel_13_394" written by ABC on Sun Jul 19 10:50:51 2020

module kernel_13_394 ( 
    i_13_394_58_0, i_13_394_59_0, i_13_394_140_0, i_13_394_190_0,
    i_13_394_256_0, i_13_394_259_0, i_13_394_334_0, i_13_394_428_0,
    i_13_394_484_0, i_13_394_485_0, i_13_394_612_0, i_13_394_625_0,
    i_13_394_626_0, i_13_394_628_0, i_13_394_629_0, i_13_394_657_0,
    i_13_394_685_0, i_13_394_779_0, i_13_394_781_0, i_13_394_913_0,
    i_13_394_914_0, i_13_394_977_0, i_13_394_980_0, i_13_394_1094_0,
    i_13_394_1115_0, i_13_394_1117_0, i_13_394_1228_0, i_13_394_1263_0,
    i_13_394_1274_0, i_13_394_1318_0, i_13_394_1343_0, i_13_394_1469_0,
    i_13_394_1480_0, i_13_394_1481_0, i_13_394_1484_0, i_13_394_1512_0,
    i_13_394_1561_0, i_13_394_1633_0, i_13_394_1639_0, i_13_394_1648_0,
    i_13_394_1649_0, i_13_394_1670_0, i_13_394_1673_0, i_13_394_1696_0,
    i_13_394_1733_0, i_13_394_1756_0, i_13_394_1778_0, i_13_394_1796_0,
    i_13_394_1801_0, i_13_394_1886_0, i_13_394_2180_0, i_13_394_2230_0,
    i_13_394_2307_0, i_13_394_2308_0, i_13_394_2366_0, i_13_394_2377_0,
    i_13_394_2380_0, i_13_394_2381_0, i_13_394_2425_0, i_13_394_2447_0,
    i_13_394_2461_0, i_13_394_2483_0, i_13_394_2647_0, i_13_394_2743_0,
    i_13_394_2781_0, i_13_394_2783_0, i_13_394_2849_0, i_13_394_2899_0,
    i_13_394_2950_0, i_13_394_2951_0, i_13_394_2953_0, i_13_394_3001_0,
    i_13_394_3005_0, i_13_394_3074_0, i_13_394_3091_0, i_13_394_3110_0,
    i_13_394_3135_0, i_13_394_3145_0, i_13_394_3153_0, i_13_394_3163_0,
    i_13_394_3308_0, i_13_394_3356_0, i_13_394_3433_0, i_13_394_3529_0,
    i_13_394_3637_0, i_13_394_3754_0, i_13_394_3766_0, i_13_394_3799_0,
    i_13_394_3842_0, i_13_394_3843_0, i_13_394_3874_0, i_13_394_4018_0,
    i_13_394_4187_0, i_13_394_4231_0, i_13_394_4294_0, i_13_394_4391_0,
    i_13_394_4448_0, i_13_394_4468_0, i_13_394_4481_0, i_13_394_4508_0,
    o_13_394_0_0  );
  input  i_13_394_58_0, i_13_394_59_0, i_13_394_140_0, i_13_394_190_0,
    i_13_394_256_0, i_13_394_259_0, i_13_394_334_0, i_13_394_428_0,
    i_13_394_484_0, i_13_394_485_0, i_13_394_612_0, i_13_394_625_0,
    i_13_394_626_0, i_13_394_628_0, i_13_394_629_0, i_13_394_657_0,
    i_13_394_685_0, i_13_394_779_0, i_13_394_781_0, i_13_394_913_0,
    i_13_394_914_0, i_13_394_977_0, i_13_394_980_0, i_13_394_1094_0,
    i_13_394_1115_0, i_13_394_1117_0, i_13_394_1228_0, i_13_394_1263_0,
    i_13_394_1274_0, i_13_394_1318_0, i_13_394_1343_0, i_13_394_1469_0,
    i_13_394_1480_0, i_13_394_1481_0, i_13_394_1484_0, i_13_394_1512_0,
    i_13_394_1561_0, i_13_394_1633_0, i_13_394_1639_0, i_13_394_1648_0,
    i_13_394_1649_0, i_13_394_1670_0, i_13_394_1673_0, i_13_394_1696_0,
    i_13_394_1733_0, i_13_394_1756_0, i_13_394_1778_0, i_13_394_1796_0,
    i_13_394_1801_0, i_13_394_1886_0, i_13_394_2180_0, i_13_394_2230_0,
    i_13_394_2307_0, i_13_394_2308_0, i_13_394_2366_0, i_13_394_2377_0,
    i_13_394_2380_0, i_13_394_2381_0, i_13_394_2425_0, i_13_394_2447_0,
    i_13_394_2461_0, i_13_394_2483_0, i_13_394_2647_0, i_13_394_2743_0,
    i_13_394_2781_0, i_13_394_2783_0, i_13_394_2849_0, i_13_394_2899_0,
    i_13_394_2950_0, i_13_394_2951_0, i_13_394_2953_0, i_13_394_3001_0,
    i_13_394_3005_0, i_13_394_3074_0, i_13_394_3091_0, i_13_394_3110_0,
    i_13_394_3135_0, i_13_394_3145_0, i_13_394_3153_0, i_13_394_3163_0,
    i_13_394_3308_0, i_13_394_3356_0, i_13_394_3433_0, i_13_394_3529_0,
    i_13_394_3637_0, i_13_394_3754_0, i_13_394_3766_0, i_13_394_3799_0,
    i_13_394_3842_0, i_13_394_3843_0, i_13_394_3874_0, i_13_394_4018_0,
    i_13_394_4187_0, i_13_394_4231_0, i_13_394_4294_0, i_13_394_4391_0,
    i_13_394_4448_0, i_13_394_4468_0, i_13_394_4481_0, i_13_394_4508_0;
  output o_13_394_0_0;
  assign o_13_394_0_0 = ~(~i_13_394_685_0 | ~i_13_394_2377_0 | (~i_13_394_2380_0 & i_13_394_3163_0) | (~i_13_394_58_0 & ~i_13_394_1778_0) | (~i_13_394_2781_0 & i_13_394_3145_0 & i_13_394_3529_0 & ~i_13_394_4187_0));
endmodule



// Benchmark "kernel_13_395" written by ABC on Sun Jul 19 10:50:52 2020

module kernel_13_395 ( 
    i_13_395_28_0, i_13_395_52_0, i_13_395_126_0, i_13_395_253_0,
    i_13_395_274_0, i_13_395_279_0, i_13_395_282_0, i_13_395_306_0,
    i_13_395_307_0, i_13_395_310_0, i_13_395_315_0, i_13_395_316_0,
    i_13_395_334_0, i_13_395_371_0, i_13_395_373_0, i_13_395_453_0,
    i_13_395_504_0, i_13_395_589_0, i_13_395_615_0, i_13_395_616_0,
    i_13_395_642_0, i_13_395_643_0, i_13_395_679_0, i_13_395_685_0,
    i_13_395_687_0, i_13_395_688_0, i_13_395_757_0, i_13_395_819_0,
    i_13_395_820_0, i_13_395_832_0, i_13_395_858_0, i_13_395_976_0,
    i_13_395_1075_0, i_13_395_1138_0, i_13_395_1222_0, i_13_395_1228_0,
    i_13_395_1284_0, i_13_395_1404_0, i_13_395_1422_0, i_13_395_1426_0,
    i_13_395_1518_0, i_13_395_1594_0, i_13_395_1597_0, i_13_395_1768_0,
    i_13_395_1813_0, i_13_395_1819_0, i_13_395_1827_0, i_13_395_1926_0,
    i_13_395_1999_0, i_13_395_2175_0, i_13_395_2200_0, i_13_395_2434_0,
    i_13_395_2436_0, i_13_395_2443_0, i_13_395_2497_0, i_13_395_2647_0,
    i_13_395_2673_0, i_13_395_2676_0, i_13_395_2695_0, i_13_395_2707_0,
    i_13_395_2713_0, i_13_395_2715_0, i_13_395_2740_0, i_13_395_2767_0,
    i_13_395_2845_0, i_13_395_2853_0, i_13_395_2883_0, i_13_395_2884_0,
    i_13_395_3087_0, i_13_395_3102_0, i_13_395_3106_0, i_13_395_3205_0,
    i_13_395_3207_0, i_13_395_3217_0, i_13_395_3415_0, i_13_395_3441_0,
    i_13_395_3457_0, i_13_395_3460_0, i_13_395_3486_0, i_13_395_3609_0,
    i_13_395_3688_0, i_13_395_3720_0, i_13_395_3726_0, i_13_395_3735_0,
    i_13_395_3736_0, i_13_395_3769_0, i_13_395_3888_0, i_13_395_3889_0,
    i_13_395_3919_0, i_13_395_4014_0, i_13_395_4015_0, i_13_395_4032_0,
    i_13_395_4033_0, i_13_395_4162_0, i_13_395_4269_0, i_13_395_4381_0,
    i_13_395_4392_0, i_13_395_4393_0, i_13_395_4513_0, i_13_395_4594_0,
    o_13_395_0_0  );
  input  i_13_395_28_0, i_13_395_52_0, i_13_395_126_0, i_13_395_253_0,
    i_13_395_274_0, i_13_395_279_0, i_13_395_282_0, i_13_395_306_0,
    i_13_395_307_0, i_13_395_310_0, i_13_395_315_0, i_13_395_316_0,
    i_13_395_334_0, i_13_395_371_0, i_13_395_373_0, i_13_395_453_0,
    i_13_395_504_0, i_13_395_589_0, i_13_395_615_0, i_13_395_616_0,
    i_13_395_642_0, i_13_395_643_0, i_13_395_679_0, i_13_395_685_0,
    i_13_395_687_0, i_13_395_688_0, i_13_395_757_0, i_13_395_819_0,
    i_13_395_820_0, i_13_395_832_0, i_13_395_858_0, i_13_395_976_0,
    i_13_395_1075_0, i_13_395_1138_0, i_13_395_1222_0, i_13_395_1228_0,
    i_13_395_1284_0, i_13_395_1404_0, i_13_395_1422_0, i_13_395_1426_0,
    i_13_395_1518_0, i_13_395_1594_0, i_13_395_1597_0, i_13_395_1768_0,
    i_13_395_1813_0, i_13_395_1819_0, i_13_395_1827_0, i_13_395_1926_0,
    i_13_395_1999_0, i_13_395_2175_0, i_13_395_2200_0, i_13_395_2434_0,
    i_13_395_2436_0, i_13_395_2443_0, i_13_395_2497_0, i_13_395_2647_0,
    i_13_395_2673_0, i_13_395_2676_0, i_13_395_2695_0, i_13_395_2707_0,
    i_13_395_2713_0, i_13_395_2715_0, i_13_395_2740_0, i_13_395_2767_0,
    i_13_395_2845_0, i_13_395_2853_0, i_13_395_2883_0, i_13_395_2884_0,
    i_13_395_3087_0, i_13_395_3102_0, i_13_395_3106_0, i_13_395_3205_0,
    i_13_395_3207_0, i_13_395_3217_0, i_13_395_3415_0, i_13_395_3441_0,
    i_13_395_3457_0, i_13_395_3460_0, i_13_395_3486_0, i_13_395_3609_0,
    i_13_395_3688_0, i_13_395_3720_0, i_13_395_3726_0, i_13_395_3735_0,
    i_13_395_3736_0, i_13_395_3769_0, i_13_395_3888_0, i_13_395_3889_0,
    i_13_395_3919_0, i_13_395_4014_0, i_13_395_4015_0, i_13_395_4032_0,
    i_13_395_4033_0, i_13_395_4162_0, i_13_395_4269_0, i_13_395_4381_0,
    i_13_395_4392_0, i_13_395_4393_0, i_13_395_4513_0, i_13_395_4594_0;
  output o_13_395_0_0;
  assign o_13_395_0_0 = ~((~i_13_395_3888_0 & (~i_13_395_1999_0 | (~i_13_395_315_0 & i_13_395_3609_0))) | (~i_13_395_1404_0 & ~i_13_395_2695_0) | (i_13_395_2767_0 & ~i_13_395_3609_0));
endmodule



// Benchmark "kernel_13_396" written by ABC on Sun Jul 19 10:50:53 2020

module kernel_13_396 ( 
    i_13_396_46_0, i_13_396_73_0, i_13_396_92_0, i_13_396_119_0,
    i_13_396_173_0, i_13_396_175_0, i_13_396_181_0, i_13_396_307_0,
    i_13_396_311_0, i_13_396_409_0, i_13_396_550_0, i_13_396_551_0,
    i_13_396_568_0, i_13_396_569_0, i_13_396_626_0, i_13_396_643_0,
    i_13_396_649_0, i_13_396_686_0, i_13_396_847_0, i_13_396_848_0,
    i_13_396_937_0, i_13_396_982_0, i_13_396_983_0, i_13_396_1120_0,
    i_13_396_1129_0, i_13_396_1130_0, i_13_396_1136_0, i_13_396_1253_0,
    i_13_396_1324_0, i_13_396_1328_0, i_13_396_1361_0, i_13_396_1372_0,
    i_13_396_1405_0, i_13_396_1406_0, i_13_396_1468_0, i_13_396_1523_0,
    i_13_396_1630_0, i_13_396_1750_0, i_13_396_1751_0, i_13_396_1778_0,
    i_13_396_1805_0, i_13_396_1936_0, i_13_396_2021_0, i_13_396_2098_0,
    i_13_396_2120_0, i_13_396_2264_0, i_13_396_2287_0, i_13_396_2384_0,
    i_13_396_2470_0, i_13_396_2507_0, i_13_396_2543_0, i_13_396_2567_0,
    i_13_396_2593_0, i_13_396_2692_0, i_13_396_2696_0, i_13_396_2851_0,
    i_13_396_2884_0, i_13_396_2900_0, i_13_396_2926_0, i_13_396_2980_0,
    i_13_396_2983_0, i_13_396_3002_0, i_13_396_3007_0, i_13_396_3029_0,
    i_13_396_3047_0, i_13_396_3106_0, i_13_396_3107_0, i_13_396_3172_0,
    i_13_396_3209_0, i_13_396_3262_0, i_13_396_3344_0, i_13_396_3403_0,
    i_13_396_3407_0, i_13_396_3485_0, i_13_396_3547_0, i_13_396_3568_0,
    i_13_396_3638_0, i_13_396_3640_0, i_13_396_3685_0, i_13_396_3754_0,
    i_13_396_3764_0, i_13_396_3802_0, i_13_396_3820_0, i_13_396_3821_0,
    i_13_396_3892_0, i_13_396_3898_0, i_13_396_3908_0, i_13_396_3992_0,
    i_13_396_4036_0, i_13_396_4081_0, i_13_396_4250_0, i_13_396_4262_0,
    i_13_396_4322_0, i_13_396_4399_0, i_13_396_4402_0, i_13_396_4495_0,
    i_13_396_4564_0, i_13_396_4565_0, i_13_396_4595_0, i_13_396_4604_0,
    o_13_396_0_0  );
  input  i_13_396_46_0, i_13_396_73_0, i_13_396_92_0, i_13_396_119_0,
    i_13_396_173_0, i_13_396_175_0, i_13_396_181_0, i_13_396_307_0,
    i_13_396_311_0, i_13_396_409_0, i_13_396_550_0, i_13_396_551_0,
    i_13_396_568_0, i_13_396_569_0, i_13_396_626_0, i_13_396_643_0,
    i_13_396_649_0, i_13_396_686_0, i_13_396_847_0, i_13_396_848_0,
    i_13_396_937_0, i_13_396_982_0, i_13_396_983_0, i_13_396_1120_0,
    i_13_396_1129_0, i_13_396_1130_0, i_13_396_1136_0, i_13_396_1253_0,
    i_13_396_1324_0, i_13_396_1328_0, i_13_396_1361_0, i_13_396_1372_0,
    i_13_396_1405_0, i_13_396_1406_0, i_13_396_1468_0, i_13_396_1523_0,
    i_13_396_1630_0, i_13_396_1750_0, i_13_396_1751_0, i_13_396_1778_0,
    i_13_396_1805_0, i_13_396_1936_0, i_13_396_2021_0, i_13_396_2098_0,
    i_13_396_2120_0, i_13_396_2264_0, i_13_396_2287_0, i_13_396_2384_0,
    i_13_396_2470_0, i_13_396_2507_0, i_13_396_2543_0, i_13_396_2567_0,
    i_13_396_2593_0, i_13_396_2692_0, i_13_396_2696_0, i_13_396_2851_0,
    i_13_396_2884_0, i_13_396_2900_0, i_13_396_2926_0, i_13_396_2980_0,
    i_13_396_2983_0, i_13_396_3002_0, i_13_396_3007_0, i_13_396_3029_0,
    i_13_396_3047_0, i_13_396_3106_0, i_13_396_3107_0, i_13_396_3172_0,
    i_13_396_3209_0, i_13_396_3262_0, i_13_396_3344_0, i_13_396_3403_0,
    i_13_396_3407_0, i_13_396_3485_0, i_13_396_3547_0, i_13_396_3568_0,
    i_13_396_3638_0, i_13_396_3640_0, i_13_396_3685_0, i_13_396_3754_0,
    i_13_396_3764_0, i_13_396_3802_0, i_13_396_3820_0, i_13_396_3821_0,
    i_13_396_3892_0, i_13_396_3898_0, i_13_396_3908_0, i_13_396_3992_0,
    i_13_396_4036_0, i_13_396_4081_0, i_13_396_4250_0, i_13_396_4262_0,
    i_13_396_4322_0, i_13_396_4399_0, i_13_396_4402_0, i_13_396_4495_0,
    i_13_396_4564_0, i_13_396_4565_0, i_13_396_4595_0, i_13_396_4604_0;
  output o_13_396_0_0;
  assign o_13_396_0_0 = ~(~i_13_396_569_0 | (~i_13_396_311_0 & ~i_13_396_3547_0 & ~i_13_396_4565_0));
endmodule



// Benchmark "kernel_13_397" written by ABC on Sun Jul 19 10:50:54 2020

module kernel_13_397 ( 
    i_13_397_30_0, i_13_397_31_0, i_13_397_58_0, i_13_397_90_0,
    i_13_397_91_0, i_13_397_108_0, i_13_397_228_0, i_13_397_459_0,
    i_13_397_534_0, i_13_397_660_0, i_13_397_685_0, i_13_397_732_0,
    i_13_397_742_0, i_13_397_757_0, i_13_397_793_0, i_13_397_811_0,
    i_13_397_850_0, i_13_397_855_0, i_13_397_957_0, i_13_397_958_0,
    i_13_397_1075_0, i_13_397_1083_0, i_13_397_1084_0, i_13_397_1117_0,
    i_13_397_1215_0, i_13_397_1228_0, i_13_397_1324_0, i_13_397_1462_0,
    i_13_397_1470_0, i_13_397_1485_0, i_13_397_1486_0, i_13_397_1677_0,
    i_13_397_1758_0, i_13_397_1813_0, i_13_397_1836_0, i_13_397_1899_0,
    i_13_397_1957_0, i_13_397_1998_0, i_13_397_1999_0, i_13_397_2043_0,
    i_13_397_2205_0, i_13_397_2227_0, i_13_397_2259_0, i_13_397_2286_0,
    i_13_397_2313_0, i_13_397_2421_0, i_13_397_2431_0, i_13_397_2497_0,
    i_13_397_2529_0, i_13_397_2538_0, i_13_397_2539_0, i_13_397_2563_0,
    i_13_397_2712_0, i_13_397_2731_0, i_13_397_2916_0, i_13_397_2917_0,
    i_13_397_2937_0, i_13_397_2979_0, i_13_397_3018_0, i_13_397_3019_0,
    i_13_397_3025_0, i_13_397_3043_0, i_13_397_3088_0, i_13_397_3099_0,
    i_13_397_3106_0, i_13_397_3126_0, i_13_397_3144_0, i_13_397_3145_0,
    i_13_397_3168_0, i_13_397_3325_0, i_13_397_3385_0, i_13_397_3457_0,
    i_13_397_3486_0, i_13_397_3487_0, i_13_397_3577_0, i_13_397_3609_0,
    i_13_397_3616_0, i_13_397_3622_0, i_13_397_3717_0, i_13_397_3802_0,
    i_13_397_3844_0, i_13_397_3846_0, i_13_397_3870_0, i_13_397_3871_0,
    i_13_397_3880_0, i_13_397_3906_0, i_13_397_3919_0, i_13_397_4006_0,
    i_13_397_4032_0, i_13_397_4054_0, i_13_397_4116_0, i_13_397_4121_0,
    i_13_397_4174_0, i_13_397_4186_0, i_13_397_4294_0, i_13_397_4347_0,
    i_13_397_4396_0, i_13_397_4521_0, i_13_397_4542_0, i_13_397_4557_0,
    o_13_397_0_0  );
  input  i_13_397_30_0, i_13_397_31_0, i_13_397_58_0, i_13_397_90_0,
    i_13_397_91_0, i_13_397_108_0, i_13_397_228_0, i_13_397_459_0,
    i_13_397_534_0, i_13_397_660_0, i_13_397_685_0, i_13_397_732_0,
    i_13_397_742_0, i_13_397_757_0, i_13_397_793_0, i_13_397_811_0,
    i_13_397_850_0, i_13_397_855_0, i_13_397_957_0, i_13_397_958_0,
    i_13_397_1075_0, i_13_397_1083_0, i_13_397_1084_0, i_13_397_1117_0,
    i_13_397_1215_0, i_13_397_1228_0, i_13_397_1324_0, i_13_397_1462_0,
    i_13_397_1470_0, i_13_397_1485_0, i_13_397_1486_0, i_13_397_1677_0,
    i_13_397_1758_0, i_13_397_1813_0, i_13_397_1836_0, i_13_397_1899_0,
    i_13_397_1957_0, i_13_397_1998_0, i_13_397_1999_0, i_13_397_2043_0,
    i_13_397_2205_0, i_13_397_2227_0, i_13_397_2259_0, i_13_397_2286_0,
    i_13_397_2313_0, i_13_397_2421_0, i_13_397_2431_0, i_13_397_2497_0,
    i_13_397_2529_0, i_13_397_2538_0, i_13_397_2539_0, i_13_397_2563_0,
    i_13_397_2712_0, i_13_397_2731_0, i_13_397_2916_0, i_13_397_2917_0,
    i_13_397_2937_0, i_13_397_2979_0, i_13_397_3018_0, i_13_397_3019_0,
    i_13_397_3025_0, i_13_397_3043_0, i_13_397_3088_0, i_13_397_3099_0,
    i_13_397_3106_0, i_13_397_3126_0, i_13_397_3144_0, i_13_397_3145_0,
    i_13_397_3168_0, i_13_397_3325_0, i_13_397_3385_0, i_13_397_3457_0,
    i_13_397_3486_0, i_13_397_3487_0, i_13_397_3577_0, i_13_397_3609_0,
    i_13_397_3616_0, i_13_397_3622_0, i_13_397_3717_0, i_13_397_3802_0,
    i_13_397_3844_0, i_13_397_3846_0, i_13_397_3870_0, i_13_397_3871_0,
    i_13_397_3880_0, i_13_397_3906_0, i_13_397_3919_0, i_13_397_4006_0,
    i_13_397_4032_0, i_13_397_4054_0, i_13_397_4116_0, i_13_397_4121_0,
    i_13_397_4174_0, i_13_397_4186_0, i_13_397_4294_0, i_13_397_4347_0,
    i_13_397_4396_0, i_13_397_4521_0, i_13_397_4542_0, i_13_397_4557_0;
  output o_13_397_0_0;
  assign o_13_397_0_0 = ~(~i_13_397_2529_0 | i_13_397_3487_0);
endmodule



// Benchmark "kernel_13_398" written by ABC on Sun Jul 19 10:50:55 2020

module kernel_13_398 ( 
    i_13_398_124_0, i_13_398_139_0, i_13_398_165_0, i_13_398_169_0,
    i_13_398_179_0, i_13_398_229_0, i_13_398_258_0, i_13_398_283_0,
    i_13_398_284_0, i_13_398_285_0, i_13_398_286_0, i_13_398_414_0,
    i_13_398_512_0, i_13_398_517_0, i_13_398_572_0, i_13_398_662_0,
    i_13_398_768_0, i_13_398_817_0, i_13_398_849_0, i_13_398_850_0,
    i_13_398_853_0, i_13_398_984_0, i_13_398_985_0, i_13_398_1019_0,
    i_13_398_1021_0, i_13_398_1022_0, i_13_398_1037_0, i_13_398_1226_0,
    i_13_398_1310_0, i_13_398_1313_0, i_13_398_1334_0, i_13_398_1344_0,
    i_13_398_1506_0, i_13_398_1549_0, i_13_398_1550_0, i_13_398_1714_0,
    i_13_398_1723_0, i_13_398_1749_0, i_13_398_1786_0, i_13_398_1858_0,
    i_13_398_1859_0, i_13_398_1860_0, i_13_398_1861_0, i_13_398_1921_0,
    i_13_398_2014_0, i_13_398_2142_0, i_13_398_2298_0, i_13_398_2407_0,
    i_13_398_2657_0, i_13_398_2680_0, i_13_398_2852_0, i_13_398_2857_0,
    i_13_398_2967_0, i_13_398_3010_0, i_13_398_3011_0, i_13_398_3014_0,
    i_13_398_3030_0, i_13_398_3037_0, i_13_398_3040_0, i_13_398_3108_0,
    i_13_398_3109_0, i_13_398_3112_0, i_13_398_3122_0, i_13_398_3163_0,
    i_13_398_3217_0, i_13_398_3218_0, i_13_398_3400_0, i_13_398_3542_0,
    i_13_398_3577_0, i_13_398_3636_0, i_13_398_3785_0, i_13_398_3838_0,
    i_13_398_3847_0, i_13_398_3856_0, i_13_398_3861_0, i_13_398_3865_0,
    i_13_398_3866_0, i_13_398_3868_0, i_13_398_3892_0, i_13_398_3910_0,
    i_13_398_3911_0, i_13_398_3913_0, i_13_398_3916_0, i_13_398_3936_0,
    i_13_398_3982_0, i_13_398_4047_0, i_13_398_4066_0, i_13_398_4162_0,
    i_13_398_4170_0, i_13_398_4204_0, i_13_398_4207_0, i_13_398_4250_0,
    i_13_398_4253_0, i_13_398_4258_0, i_13_398_4261_0, i_13_398_4304_0,
    i_13_398_4345_0, i_13_398_4351_0, i_13_398_4358_0, i_13_398_4379_0,
    o_13_398_0_0  );
  input  i_13_398_124_0, i_13_398_139_0, i_13_398_165_0, i_13_398_169_0,
    i_13_398_179_0, i_13_398_229_0, i_13_398_258_0, i_13_398_283_0,
    i_13_398_284_0, i_13_398_285_0, i_13_398_286_0, i_13_398_414_0,
    i_13_398_512_0, i_13_398_517_0, i_13_398_572_0, i_13_398_662_0,
    i_13_398_768_0, i_13_398_817_0, i_13_398_849_0, i_13_398_850_0,
    i_13_398_853_0, i_13_398_984_0, i_13_398_985_0, i_13_398_1019_0,
    i_13_398_1021_0, i_13_398_1022_0, i_13_398_1037_0, i_13_398_1226_0,
    i_13_398_1310_0, i_13_398_1313_0, i_13_398_1334_0, i_13_398_1344_0,
    i_13_398_1506_0, i_13_398_1549_0, i_13_398_1550_0, i_13_398_1714_0,
    i_13_398_1723_0, i_13_398_1749_0, i_13_398_1786_0, i_13_398_1858_0,
    i_13_398_1859_0, i_13_398_1860_0, i_13_398_1861_0, i_13_398_1921_0,
    i_13_398_2014_0, i_13_398_2142_0, i_13_398_2298_0, i_13_398_2407_0,
    i_13_398_2657_0, i_13_398_2680_0, i_13_398_2852_0, i_13_398_2857_0,
    i_13_398_2967_0, i_13_398_3010_0, i_13_398_3011_0, i_13_398_3014_0,
    i_13_398_3030_0, i_13_398_3037_0, i_13_398_3040_0, i_13_398_3108_0,
    i_13_398_3109_0, i_13_398_3112_0, i_13_398_3122_0, i_13_398_3163_0,
    i_13_398_3217_0, i_13_398_3218_0, i_13_398_3400_0, i_13_398_3542_0,
    i_13_398_3577_0, i_13_398_3636_0, i_13_398_3785_0, i_13_398_3838_0,
    i_13_398_3847_0, i_13_398_3856_0, i_13_398_3861_0, i_13_398_3865_0,
    i_13_398_3866_0, i_13_398_3868_0, i_13_398_3892_0, i_13_398_3910_0,
    i_13_398_3911_0, i_13_398_3913_0, i_13_398_3916_0, i_13_398_3936_0,
    i_13_398_3982_0, i_13_398_4047_0, i_13_398_4066_0, i_13_398_4162_0,
    i_13_398_4170_0, i_13_398_4204_0, i_13_398_4207_0, i_13_398_4250_0,
    i_13_398_4253_0, i_13_398_4258_0, i_13_398_4261_0, i_13_398_4304_0,
    i_13_398_4345_0, i_13_398_4351_0, i_13_398_4358_0, i_13_398_4379_0;
  output o_13_398_0_0;
  assign o_13_398_0_0 = ~(i_13_398_3037_0 | (i_13_398_3163_0 & ~i_13_398_4379_0) | (~i_13_398_3911_0 & ~i_13_398_3913_0) | (~i_13_398_2852_0 & ~i_13_398_3892_0 & ~i_13_398_4162_0));
endmodule



// Benchmark "kernel_13_399" written by ABC on Sun Jul 19 10:50:56 2020

module kernel_13_399 ( 
    i_13_399_29_0, i_13_399_91_0, i_13_399_95_0, i_13_399_104_0,
    i_13_399_118_0, i_13_399_119_0, i_13_399_158_0, i_13_399_164_0,
    i_13_399_181_0, i_13_399_182_0, i_13_399_224_0, i_13_399_383_0,
    i_13_399_395_0, i_13_399_454_0, i_13_399_515_0, i_13_399_523_0,
    i_13_399_568_0, i_13_399_572_0, i_13_399_697_0, i_13_399_824_0,
    i_13_399_856_0, i_13_399_868_0, i_13_399_913_0, i_13_399_946_0,
    i_13_399_1076_0, i_13_399_1085_0, i_13_399_1118_0, i_13_399_1190_0,
    i_13_399_1216_0, i_13_399_1301_0, i_13_399_1360_0, i_13_399_1361_0,
    i_13_399_1406_0, i_13_399_1606_0, i_13_399_1621_0, i_13_399_1694_0,
    i_13_399_1723_0, i_13_399_1786_0, i_13_399_1787_0, i_13_399_1805_0,
    i_13_399_1906_0, i_13_399_1907_0, i_13_399_1918_0, i_13_399_2000_0,
    i_13_399_2173_0, i_13_399_2174_0, i_13_399_2206_0, i_13_399_2209_0,
    i_13_399_2422_0, i_13_399_2431_0, i_13_399_2432_0, i_13_399_2434_0,
    i_13_399_2435_0, i_13_399_2552_0, i_13_399_2956_0, i_13_399_2984_0,
    i_13_399_3020_0, i_13_399_3101_0, i_13_399_3145_0, i_13_399_3146_0,
    i_13_399_3161_0, i_13_399_3163_0, i_13_399_3164_0, i_13_399_3205_0,
    i_13_399_3209_0, i_13_399_3235_0, i_13_399_3344_0, i_13_399_3380_0,
    i_13_399_3421_0, i_13_399_3461_0, i_13_399_3487_0, i_13_399_3488_0,
    i_13_399_3530_0, i_13_399_3533_0, i_13_399_3541_0, i_13_399_3542_0,
    i_13_399_3577_0, i_13_399_3700_0, i_13_399_3718_0, i_13_399_3728_0,
    i_13_399_3764_0, i_13_399_3784_0, i_13_399_3794_0, i_13_399_3844_0,
    i_13_399_3871_0, i_13_399_3872_0, i_13_399_3983_0, i_13_399_4006_0,
    i_13_399_4007_0, i_13_399_4118_0, i_13_399_4132_0, i_13_399_4204_0,
    i_13_399_4325_0, i_13_399_4348_0, i_13_399_4349_0, i_13_399_4351_0,
    i_13_399_4415_0, i_13_399_4583_0, i_13_399_4588_0, i_13_399_4589_0,
    o_13_399_0_0  );
  input  i_13_399_29_0, i_13_399_91_0, i_13_399_95_0, i_13_399_104_0,
    i_13_399_118_0, i_13_399_119_0, i_13_399_158_0, i_13_399_164_0,
    i_13_399_181_0, i_13_399_182_0, i_13_399_224_0, i_13_399_383_0,
    i_13_399_395_0, i_13_399_454_0, i_13_399_515_0, i_13_399_523_0,
    i_13_399_568_0, i_13_399_572_0, i_13_399_697_0, i_13_399_824_0,
    i_13_399_856_0, i_13_399_868_0, i_13_399_913_0, i_13_399_946_0,
    i_13_399_1076_0, i_13_399_1085_0, i_13_399_1118_0, i_13_399_1190_0,
    i_13_399_1216_0, i_13_399_1301_0, i_13_399_1360_0, i_13_399_1361_0,
    i_13_399_1406_0, i_13_399_1606_0, i_13_399_1621_0, i_13_399_1694_0,
    i_13_399_1723_0, i_13_399_1786_0, i_13_399_1787_0, i_13_399_1805_0,
    i_13_399_1906_0, i_13_399_1907_0, i_13_399_1918_0, i_13_399_2000_0,
    i_13_399_2173_0, i_13_399_2174_0, i_13_399_2206_0, i_13_399_2209_0,
    i_13_399_2422_0, i_13_399_2431_0, i_13_399_2432_0, i_13_399_2434_0,
    i_13_399_2435_0, i_13_399_2552_0, i_13_399_2956_0, i_13_399_2984_0,
    i_13_399_3020_0, i_13_399_3101_0, i_13_399_3145_0, i_13_399_3146_0,
    i_13_399_3161_0, i_13_399_3163_0, i_13_399_3164_0, i_13_399_3205_0,
    i_13_399_3209_0, i_13_399_3235_0, i_13_399_3344_0, i_13_399_3380_0,
    i_13_399_3421_0, i_13_399_3461_0, i_13_399_3487_0, i_13_399_3488_0,
    i_13_399_3530_0, i_13_399_3533_0, i_13_399_3541_0, i_13_399_3542_0,
    i_13_399_3577_0, i_13_399_3700_0, i_13_399_3718_0, i_13_399_3728_0,
    i_13_399_3764_0, i_13_399_3784_0, i_13_399_3794_0, i_13_399_3844_0,
    i_13_399_3871_0, i_13_399_3872_0, i_13_399_3983_0, i_13_399_4006_0,
    i_13_399_4007_0, i_13_399_4118_0, i_13_399_4132_0, i_13_399_4204_0,
    i_13_399_4325_0, i_13_399_4348_0, i_13_399_4349_0, i_13_399_4351_0,
    i_13_399_4415_0, i_13_399_4583_0, i_13_399_4588_0, i_13_399_4589_0;
  output o_13_399_0_0;
  assign o_13_399_0_0 = ~((~i_13_399_2435_0 & i_13_399_3487_0) | (~i_13_399_1406_0 & ~i_13_399_2422_0) | (~i_13_399_91_0 & ~i_13_399_1216_0));
endmodule



// Benchmark "kernel_13_400" written by ABC on Sun Jul 19 10:50:56 2020

module kernel_13_400 ( 
    i_13_400_71_0, i_13_400_74_0, i_13_400_76_0, i_13_400_79_0,
    i_13_400_80_0, i_13_400_139_0, i_13_400_176_0, i_13_400_309_0,
    i_13_400_323_0, i_13_400_358_0, i_13_400_376_0, i_13_400_610_0,
    i_13_400_647_0, i_13_400_672_0, i_13_400_673_0, i_13_400_674_0,
    i_13_400_683_0, i_13_400_772_0, i_13_400_814_0, i_13_400_821_0,
    i_13_400_841_0, i_13_400_952_0, i_13_400_1103_0, i_13_400_1106_0,
    i_13_400_1123_0, i_13_400_1151_0, i_13_400_1210_0, i_13_400_1276_0,
    i_13_400_1277_0, i_13_400_1282_0, i_13_400_1312_0, i_13_400_1403_0,
    i_13_400_1430_0, i_13_400_1468_0, i_13_400_1496_0, i_13_400_1509_0,
    i_13_400_1511_0, i_13_400_1600_0, i_13_400_1645_0, i_13_400_1687_0,
    i_13_400_1690_0, i_13_400_1726_0, i_13_400_1736_0, i_13_400_1750_0,
    i_13_400_1781_0, i_13_400_1798_0, i_13_400_1799_0, i_13_400_1857_0,
    i_13_400_1889_0, i_13_400_1912_0, i_13_400_1925_0, i_13_400_2002_0,
    i_13_400_2030_0, i_13_400_2032_0, i_13_400_2176_0, i_13_400_2177_0,
    i_13_400_2232_0, i_13_400_2240_0, i_13_400_2344_0, i_13_400_2407_0,
    i_13_400_2513_0, i_13_400_2654_0, i_13_400_2679_0, i_13_400_2680_0,
    i_13_400_2681_0, i_13_400_2698_0, i_13_400_2817_0, i_13_400_2818_0,
    i_13_400_2851_0, i_13_400_2852_0, i_13_400_2924_0, i_13_400_3028_0,
    i_13_400_3142_0, i_13_400_3221_0, i_13_400_3355_0, i_13_400_3386_0,
    i_13_400_3406_0, i_13_400_3607_0, i_13_400_3622_0, i_13_400_3739_0,
    i_13_400_3743_0, i_13_400_3784_0, i_13_400_3787_0, i_13_400_3797_0,
    i_13_400_3816_0, i_13_400_3860_0, i_13_400_3896_0, i_13_400_3930_0,
    i_13_400_3931_0, i_13_400_3932_0, i_13_400_3994_0, i_13_400_3995_0,
    i_13_400_4219_0, i_13_400_4372_0, i_13_400_4447_0, i_13_400_4453_0,
    i_13_400_4454_0, i_13_400_4596_0, i_13_400_4597_0, i_13_400_4598_0,
    o_13_400_0_0  );
  input  i_13_400_71_0, i_13_400_74_0, i_13_400_76_0, i_13_400_79_0,
    i_13_400_80_0, i_13_400_139_0, i_13_400_176_0, i_13_400_309_0,
    i_13_400_323_0, i_13_400_358_0, i_13_400_376_0, i_13_400_610_0,
    i_13_400_647_0, i_13_400_672_0, i_13_400_673_0, i_13_400_674_0,
    i_13_400_683_0, i_13_400_772_0, i_13_400_814_0, i_13_400_821_0,
    i_13_400_841_0, i_13_400_952_0, i_13_400_1103_0, i_13_400_1106_0,
    i_13_400_1123_0, i_13_400_1151_0, i_13_400_1210_0, i_13_400_1276_0,
    i_13_400_1277_0, i_13_400_1282_0, i_13_400_1312_0, i_13_400_1403_0,
    i_13_400_1430_0, i_13_400_1468_0, i_13_400_1496_0, i_13_400_1509_0,
    i_13_400_1511_0, i_13_400_1600_0, i_13_400_1645_0, i_13_400_1687_0,
    i_13_400_1690_0, i_13_400_1726_0, i_13_400_1736_0, i_13_400_1750_0,
    i_13_400_1781_0, i_13_400_1798_0, i_13_400_1799_0, i_13_400_1857_0,
    i_13_400_1889_0, i_13_400_1912_0, i_13_400_1925_0, i_13_400_2002_0,
    i_13_400_2030_0, i_13_400_2032_0, i_13_400_2176_0, i_13_400_2177_0,
    i_13_400_2232_0, i_13_400_2240_0, i_13_400_2344_0, i_13_400_2407_0,
    i_13_400_2513_0, i_13_400_2654_0, i_13_400_2679_0, i_13_400_2680_0,
    i_13_400_2681_0, i_13_400_2698_0, i_13_400_2817_0, i_13_400_2818_0,
    i_13_400_2851_0, i_13_400_2852_0, i_13_400_2924_0, i_13_400_3028_0,
    i_13_400_3142_0, i_13_400_3221_0, i_13_400_3355_0, i_13_400_3386_0,
    i_13_400_3406_0, i_13_400_3607_0, i_13_400_3622_0, i_13_400_3739_0,
    i_13_400_3743_0, i_13_400_3784_0, i_13_400_3787_0, i_13_400_3797_0,
    i_13_400_3816_0, i_13_400_3860_0, i_13_400_3896_0, i_13_400_3930_0,
    i_13_400_3931_0, i_13_400_3932_0, i_13_400_3994_0, i_13_400_3995_0,
    i_13_400_4219_0, i_13_400_4372_0, i_13_400_4447_0, i_13_400_4453_0,
    i_13_400_4454_0, i_13_400_4596_0, i_13_400_4597_0, i_13_400_4598_0;
  output o_13_400_0_0;
  assign o_13_400_0_0 = ~((~i_13_400_3932_0 & (~i_13_400_683_0 | i_13_400_2924_0)) | (~i_13_400_71_0 & ~i_13_400_1511_0 & ~i_13_400_2851_0));
endmodule



// Benchmark "kernel_13_401" written by ABC on Sun Jul 19 10:50:57 2020

module kernel_13_401 ( 
    i_13_401_112_0, i_13_401_171_0, i_13_401_189_0, i_13_401_316_0,
    i_13_401_325_0, i_13_401_414_0, i_13_401_415_0, i_13_401_416_0,
    i_13_401_558_0, i_13_401_562_0, i_13_401_625_0, i_13_401_778_0,
    i_13_401_826_0, i_13_401_841_0, i_13_401_847_0, i_13_401_849_0,
    i_13_401_850_0, i_13_401_891_0, i_13_401_918_0, i_13_401_984_0,
    i_13_401_1021_0, i_13_401_1072_0, i_13_401_1081_0, i_13_401_1092_0,
    i_13_401_1096_0, i_13_401_1200_0, i_13_401_1224_0, i_13_401_1225_0,
    i_13_401_1230_0, i_13_401_1255_0, i_13_401_1278_0, i_13_401_1302_0,
    i_13_401_1317_0, i_13_401_1318_0, i_13_401_1480_0, i_13_401_1486_0,
    i_13_401_1491_0, i_13_401_1548_0, i_13_401_1549_0, i_13_401_1674_0,
    i_13_401_1728_0, i_13_401_1740_0, i_13_401_1746_0, i_13_401_1749_0,
    i_13_401_1756_0, i_13_401_1777_0, i_13_401_1854_0, i_13_401_1855_0,
    i_13_401_1857_0, i_13_401_1858_0, i_13_401_1954_0, i_13_401_2307_0,
    i_13_401_2308_0, i_13_401_2353_0, i_13_401_2395_0, i_13_401_2434_0,
    i_13_401_2457_0, i_13_401_2505_0, i_13_401_2539_0, i_13_401_2556_0,
    i_13_401_2586_0, i_13_401_2629_0, i_13_401_2691_0, i_13_401_2722_0,
    i_13_401_2820_0, i_13_401_2821_0, i_13_401_2850_0, i_13_401_2875_0,
    i_13_401_3000_0, i_13_401_3008_0, i_13_401_3064_0, i_13_401_3092_0,
    i_13_401_3118_0, i_13_401_3153_0, i_13_401_3163_0, i_13_401_3168_0,
    i_13_401_3234_0, i_13_401_3244_0, i_13_401_3267_0, i_13_401_3304_0,
    i_13_401_3429_0, i_13_401_3432_0, i_13_401_3484_0, i_13_401_3519_0,
    i_13_401_3537_0, i_13_401_3538_0, i_13_401_3574_0, i_13_401_3575_0,
    i_13_401_3781_0, i_13_401_3852_0, i_13_401_3906_0, i_13_401_3907_0,
    i_13_401_3909_0, i_13_401_4018_0, i_13_401_4366_0, i_13_401_4374_0,
    i_13_401_4375_0, i_13_401_4378_0, i_13_401_4393_0, i_13_401_4519_0,
    o_13_401_0_0  );
  input  i_13_401_112_0, i_13_401_171_0, i_13_401_189_0, i_13_401_316_0,
    i_13_401_325_0, i_13_401_414_0, i_13_401_415_0, i_13_401_416_0,
    i_13_401_558_0, i_13_401_562_0, i_13_401_625_0, i_13_401_778_0,
    i_13_401_826_0, i_13_401_841_0, i_13_401_847_0, i_13_401_849_0,
    i_13_401_850_0, i_13_401_891_0, i_13_401_918_0, i_13_401_984_0,
    i_13_401_1021_0, i_13_401_1072_0, i_13_401_1081_0, i_13_401_1092_0,
    i_13_401_1096_0, i_13_401_1200_0, i_13_401_1224_0, i_13_401_1225_0,
    i_13_401_1230_0, i_13_401_1255_0, i_13_401_1278_0, i_13_401_1302_0,
    i_13_401_1317_0, i_13_401_1318_0, i_13_401_1480_0, i_13_401_1486_0,
    i_13_401_1491_0, i_13_401_1548_0, i_13_401_1549_0, i_13_401_1674_0,
    i_13_401_1728_0, i_13_401_1740_0, i_13_401_1746_0, i_13_401_1749_0,
    i_13_401_1756_0, i_13_401_1777_0, i_13_401_1854_0, i_13_401_1855_0,
    i_13_401_1857_0, i_13_401_1858_0, i_13_401_1954_0, i_13_401_2307_0,
    i_13_401_2308_0, i_13_401_2353_0, i_13_401_2395_0, i_13_401_2434_0,
    i_13_401_2457_0, i_13_401_2505_0, i_13_401_2539_0, i_13_401_2556_0,
    i_13_401_2586_0, i_13_401_2629_0, i_13_401_2691_0, i_13_401_2722_0,
    i_13_401_2820_0, i_13_401_2821_0, i_13_401_2850_0, i_13_401_2875_0,
    i_13_401_3000_0, i_13_401_3008_0, i_13_401_3064_0, i_13_401_3092_0,
    i_13_401_3118_0, i_13_401_3153_0, i_13_401_3163_0, i_13_401_3168_0,
    i_13_401_3234_0, i_13_401_3244_0, i_13_401_3267_0, i_13_401_3304_0,
    i_13_401_3429_0, i_13_401_3432_0, i_13_401_3484_0, i_13_401_3519_0,
    i_13_401_3537_0, i_13_401_3538_0, i_13_401_3574_0, i_13_401_3575_0,
    i_13_401_3781_0, i_13_401_3852_0, i_13_401_3906_0, i_13_401_3907_0,
    i_13_401_3909_0, i_13_401_4018_0, i_13_401_4366_0, i_13_401_4374_0,
    i_13_401_4375_0, i_13_401_4378_0, i_13_401_4393_0, i_13_401_4519_0;
  output o_13_401_0_0;
  assign o_13_401_0_0 = ~((i_13_401_4375_0 & i_13_401_4393_0) | (i_13_401_3092_0 & ~i_13_401_4366_0) | (i_13_401_2434_0 & i_13_401_3575_0) | (~i_13_401_414_0 & ~i_13_401_1857_0 & ~i_13_401_4378_0) | (~i_13_401_1021_0 & ~i_13_401_1749_0 & ~i_13_401_3906_0) | (~i_13_401_1486_0 & ~i_13_401_2457_0 & ~i_13_401_3537_0));
endmodule



// Benchmark "kernel_13_402" written by ABC on Sun Jul 19 10:50:58 2020

module kernel_13_402 ( 
    i_13_402_113_0, i_13_402_204_0, i_13_402_273_0, i_13_402_276_0,
    i_13_402_277_0, i_13_402_278_0, i_13_402_319_0, i_13_402_328_0,
    i_13_402_340_0, i_13_402_366_0, i_13_402_368_0, i_13_402_391_0,
    i_13_402_394_0, i_13_402_447_0, i_13_402_457_0, i_13_402_492_0,
    i_13_402_565_0, i_13_402_637_0, i_13_402_643_0, i_13_402_744_0,
    i_13_402_745_0, i_13_402_746_0, i_13_402_845_0, i_13_402_871_0,
    i_13_402_948_0, i_13_402_978_0, i_13_402_979_0, i_13_402_1023_0,
    i_13_402_1070_0, i_13_402_1086_0, i_13_402_1087_0, i_13_402_1088_0,
    i_13_402_1096_0, i_13_402_1141_0, i_13_402_1349_0, i_13_402_1465_0,
    i_13_402_1519_0, i_13_402_1623_0, i_13_402_1625_0, i_13_402_1815_0,
    i_13_402_1816_0, i_13_402_1943_0, i_13_402_1950_0, i_13_402_1951_0,
    i_13_402_2022_0, i_13_402_2060_0, i_13_402_2266_0, i_13_402_2347_0,
    i_13_402_2433_0, i_13_402_2437_0, i_13_402_2464_0, i_13_402_2480_0,
    i_13_402_2613_0, i_13_402_2677_0, i_13_402_2715_0, i_13_402_2716_0,
    i_13_402_2787_0, i_13_402_2788_0, i_13_402_2912_0, i_13_402_2921_0,
    i_13_402_2987_0, i_13_402_3003_0, i_13_402_3010_0, i_13_402_3068_0,
    i_13_402_3112_0, i_13_402_3127_0, i_13_402_3146_0, i_13_402_3166_0,
    i_13_402_3220_0, i_13_402_3229_0, i_13_402_3238_0, i_13_402_3417_0,
    i_13_402_3419_0, i_13_402_3451_0, i_13_402_3524_0, i_13_402_3568_0,
    i_13_402_3607_0, i_13_402_3658_0, i_13_402_3687_0, i_13_402_3688_0,
    i_13_402_3742_0, i_13_402_4001_0, i_13_402_4049_0, i_13_402_4093_0,
    i_13_402_4104_0, i_13_402_4120_0, i_13_402_4173_0, i_13_402_4237_0,
    i_13_402_4273_0, i_13_402_4297_0, i_13_402_4327_0, i_13_402_4333_0,
    i_13_402_4343_0, i_13_402_4399_0, i_13_402_4417_0, i_13_402_4495_0,
    i_13_402_4522_0, i_13_402_4533_0, i_13_402_4544_0, i_13_402_4578_0,
    o_13_402_0_0  );
  input  i_13_402_113_0, i_13_402_204_0, i_13_402_273_0, i_13_402_276_0,
    i_13_402_277_0, i_13_402_278_0, i_13_402_319_0, i_13_402_328_0,
    i_13_402_340_0, i_13_402_366_0, i_13_402_368_0, i_13_402_391_0,
    i_13_402_394_0, i_13_402_447_0, i_13_402_457_0, i_13_402_492_0,
    i_13_402_565_0, i_13_402_637_0, i_13_402_643_0, i_13_402_744_0,
    i_13_402_745_0, i_13_402_746_0, i_13_402_845_0, i_13_402_871_0,
    i_13_402_948_0, i_13_402_978_0, i_13_402_979_0, i_13_402_1023_0,
    i_13_402_1070_0, i_13_402_1086_0, i_13_402_1087_0, i_13_402_1088_0,
    i_13_402_1096_0, i_13_402_1141_0, i_13_402_1349_0, i_13_402_1465_0,
    i_13_402_1519_0, i_13_402_1623_0, i_13_402_1625_0, i_13_402_1815_0,
    i_13_402_1816_0, i_13_402_1943_0, i_13_402_1950_0, i_13_402_1951_0,
    i_13_402_2022_0, i_13_402_2060_0, i_13_402_2266_0, i_13_402_2347_0,
    i_13_402_2433_0, i_13_402_2437_0, i_13_402_2464_0, i_13_402_2480_0,
    i_13_402_2613_0, i_13_402_2677_0, i_13_402_2715_0, i_13_402_2716_0,
    i_13_402_2787_0, i_13_402_2788_0, i_13_402_2912_0, i_13_402_2921_0,
    i_13_402_2987_0, i_13_402_3003_0, i_13_402_3010_0, i_13_402_3068_0,
    i_13_402_3112_0, i_13_402_3127_0, i_13_402_3146_0, i_13_402_3166_0,
    i_13_402_3220_0, i_13_402_3229_0, i_13_402_3238_0, i_13_402_3417_0,
    i_13_402_3419_0, i_13_402_3451_0, i_13_402_3524_0, i_13_402_3568_0,
    i_13_402_3607_0, i_13_402_3658_0, i_13_402_3687_0, i_13_402_3688_0,
    i_13_402_3742_0, i_13_402_4001_0, i_13_402_4049_0, i_13_402_4093_0,
    i_13_402_4104_0, i_13_402_4120_0, i_13_402_4173_0, i_13_402_4237_0,
    i_13_402_4273_0, i_13_402_4297_0, i_13_402_4327_0, i_13_402_4333_0,
    i_13_402_4343_0, i_13_402_4399_0, i_13_402_4417_0, i_13_402_4495_0,
    i_13_402_4522_0, i_13_402_4533_0, i_13_402_4544_0, i_13_402_4578_0;
  output o_13_402_0_0;
  assign o_13_402_0_0 = ~((~i_13_402_1816_0 & ((~i_13_402_1086_0 & ~i_13_402_3688_0) | (~i_13_402_2716_0 & ~i_13_402_3742_0))) | (~i_13_402_3451_0 & ((~i_13_402_3238_0 & ~i_13_402_3742_0) | (~i_13_402_4093_0 & i_13_402_4333_0))) | (~i_13_402_2716_0 & ~i_13_402_3220_0) | (i_13_402_3524_0 & ~i_13_402_4273_0 & ~i_13_402_4327_0));
endmodule



// Benchmark "kernel_13_403" written by ABC on Sun Jul 19 10:50:59 2020

module kernel_13_403 ( 
    i_13_403_33_0, i_13_403_34_0, i_13_403_61_0, i_13_403_70_0,
    i_13_403_121_0, i_13_403_136_0, i_13_403_159_0, i_13_403_160_0,
    i_13_403_166_0, i_13_403_226_0, i_13_403_319_0, i_13_403_385_0,
    i_13_403_386_0, i_13_403_414_0, i_13_403_448_0, i_13_403_456_0,
    i_13_403_457_0, i_13_403_492_0, i_13_403_515_0, i_13_403_565_0,
    i_13_403_629_0, i_13_403_646_0, i_13_403_717_0, i_13_403_735_0,
    i_13_403_745_0, i_13_403_938_0, i_13_403_983_0, i_13_403_985_0,
    i_13_403_1023_0, i_13_403_1066_0, i_13_403_1096_0, i_13_403_1116_0,
    i_13_403_1132_0, i_13_403_1182_0, i_13_403_1208_0, i_13_403_1216_0,
    i_13_403_1217_0, i_13_403_1266_0, i_13_403_1275_0, i_13_403_1302_0,
    i_13_403_1304_0, i_13_403_1348_0, i_13_403_1380_0, i_13_403_1489_0,
    i_13_403_1521_0, i_13_403_1525_0, i_13_403_1605_0, i_13_403_1743_0,
    i_13_403_1774_0, i_13_403_1792_0, i_13_403_1793_0, i_13_403_1808_0,
    i_13_403_1816_0, i_13_403_1967_0, i_13_403_2056_0, i_13_403_2123_0,
    i_13_403_2209_0, i_13_403_2244_0, i_13_403_2248_0, i_13_403_2281_0,
    i_13_403_2364_0, i_13_403_2407_0, i_13_403_2705_0, i_13_403_2749_0,
    i_13_403_2851_0, i_13_403_2859_0, i_13_403_2876_0, i_13_403_3022_0,
    i_13_403_3034_0, i_13_403_3036_0, i_13_403_3094_0, i_13_403_3095_0,
    i_13_403_3101_0, i_13_403_3207_0, i_13_403_3265_0, i_13_403_3354_0,
    i_13_403_3391_0, i_13_403_3551_0, i_13_403_3564_0, i_13_403_3759_0,
    i_13_403_3768_0, i_13_403_3769_0, i_13_403_3820_0, i_13_403_3821_0,
    i_13_403_3847_0, i_13_403_3848_0, i_13_403_3859_0, i_13_403_3954_0,
    i_13_403_3985_0, i_13_403_3989_0, i_13_403_4076_0, i_13_403_4084_0,
    i_13_403_4090_0, i_13_403_4238_0, i_13_403_4273_0, i_13_403_4299_0,
    i_13_403_4328_0, i_13_403_4399_0, i_13_403_4400_0, i_13_403_4594_0,
    o_13_403_0_0  );
  input  i_13_403_33_0, i_13_403_34_0, i_13_403_61_0, i_13_403_70_0,
    i_13_403_121_0, i_13_403_136_0, i_13_403_159_0, i_13_403_160_0,
    i_13_403_166_0, i_13_403_226_0, i_13_403_319_0, i_13_403_385_0,
    i_13_403_386_0, i_13_403_414_0, i_13_403_448_0, i_13_403_456_0,
    i_13_403_457_0, i_13_403_492_0, i_13_403_515_0, i_13_403_565_0,
    i_13_403_629_0, i_13_403_646_0, i_13_403_717_0, i_13_403_735_0,
    i_13_403_745_0, i_13_403_938_0, i_13_403_983_0, i_13_403_985_0,
    i_13_403_1023_0, i_13_403_1066_0, i_13_403_1096_0, i_13_403_1116_0,
    i_13_403_1132_0, i_13_403_1182_0, i_13_403_1208_0, i_13_403_1216_0,
    i_13_403_1217_0, i_13_403_1266_0, i_13_403_1275_0, i_13_403_1302_0,
    i_13_403_1304_0, i_13_403_1348_0, i_13_403_1380_0, i_13_403_1489_0,
    i_13_403_1521_0, i_13_403_1525_0, i_13_403_1605_0, i_13_403_1743_0,
    i_13_403_1774_0, i_13_403_1792_0, i_13_403_1793_0, i_13_403_1808_0,
    i_13_403_1816_0, i_13_403_1967_0, i_13_403_2056_0, i_13_403_2123_0,
    i_13_403_2209_0, i_13_403_2244_0, i_13_403_2248_0, i_13_403_2281_0,
    i_13_403_2364_0, i_13_403_2407_0, i_13_403_2705_0, i_13_403_2749_0,
    i_13_403_2851_0, i_13_403_2859_0, i_13_403_2876_0, i_13_403_3022_0,
    i_13_403_3034_0, i_13_403_3036_0, i_13_403_3094_0, i_13_403_3095_0,
    i_13_403_3101_0, i_13_403_3207_0, i_13_403_3265_0, i_13_403_3354_0,
    i_13_403_3391_0, i_13_403_3551_0, i_13_403_3564_0, i_13_403_3759_0,
    i_13_403_3768_0, i_13_403_3769_0, i_13_403_3820_0, i_13_403_3821_0,
    i_13_403_3847_0, i_13_403_3848_0, i_13_403_3859_0, i_13_403_3954_0,
    i_13_403_3985_0, i_13_403_3989_0, i_13_403_4076_0, i_13_403_4084_0,
    i_13_403_4090_0, i_13_403_4238_0, i_13_403_4273_0, i_13_403_4299_0,
    i_13_403_4328_0, i_13_403_4399_0, i_13_403_4400_0, i_13_403_4594_0;
  output o_13_403_0_0;
  assign o_13_403_0_0 = ~((~i_13_403_1605_0 & (i_13_403_4090_0 | (~i_13_403_3036_0 & ~i_13_403_3095_0))) | (~i_13_403_2209_0 & ((~i_13_403_34_0 & ~i_13_403_3859_0) | (~i_13_403_3759_0 & ~i_13_403_3848_0 & ~i_13_403_4399_0))) | (~i_13_403_3859_0 & (~i_13_403_448_0 | (i_13_403_2407_0 & ~i_13_403_3391_0))) | (i_13_403_2407_0 & ((~i_13_403_1023_0 & ~i_13_403_3207_0 & ~i_13_403_4238_0) | (i_13_403_4238_0 & ~i_13_403_4273_0))) | (~i_13_403_3391_0 & ((i_13_403_3859_0 & ~i_13_403_4273_0) | (~i_13_403_2851_0 & ~i_13_403_4400_0))) | (~i_13_403_1816_0 & ~i_13_403_4273_0) | (i_13_403_319_0 & ~i_13_403_3551_0 & ~i_13_403_3768_0));
endmodule



// Benchmark "kernel_13_404" written by ABC on Sun Jul 19 10:50:59 2020

module kernel_13_404 ( 
    i_13_404_22_0, i_13_404_59_0, i_13_404_91_0, i_13_404_92_0,
    i_13_404_139_0, i_13_404_215_0, i_13_404_316_0, i_13_404_317_0,
    i_13_404_418_0, i_13_404_419_0, i_13_404_456_0, i_13_404_484_0,
    i_13_404_550_0, i_13_404_554_0, i_13_404_607_0, i_13_404_671_0,
    i_13_404_727_0, i_13_404_793_0, i_13_404_843_0, i_13_404_847_0,
    i_13_404_851_0, i_13_404_860_0, i_13_404_986_0, i_13_404_1018_0,
    i_13_404_1019_0, i_13_404_1083_0, i_13_404_1122_0, i_13_404_1129_0,
    i_13_404_1210_0, i_13_404_1226_0, i_13_404_1256_0, i_13_404_1300_0,
    i_13_404_1301_0, i_13_404_1306_0, i_13_404_1345_0, i_13_404_1361_0,
    i_13_404_1486_0, i_13_404_1487_0, i_13_404_1550_0, i_13_404_1599_0,
    i_13_404_1631_0, i_13_404_1644_0, i_13_404_1721_0, i_13_404_1733_0,
    i_13_404_1763_0, i_13_404_1769_0, i_13_404_1813_0, i_13_404_1855_0,
    i_13_404_1858_0, i_13_404_1859_0, i_13_404_1911_0, i_13_404_2016_0,
    i_13_404_2028_0, i_13_404_2173_0, i_13_404_2179_0, i_13_404_2207_0,
    i_13_404_2290_0, i_13_404_2296_0, i_13_404_2422_0, i_13_404_2450_0,
    i_13_404_2593_0, i_13_404_2615_0, i_13_404_2679_0, i_13_404_2697_0,
    i_13_404_2748_0, i_13_404_2857_0, i_13_404_2981_0, i_13_404_3007_0,
    i_13_404_3008_0, i_13_404_3010_0, i_13_404_3037_0, i_13_404_3110_0,
    i_13_404_3217_0, i_13_404_3389_0, i_13_404_3404_0, i_13_404_3428_0,
    i_13_404_3481_0, i_13_404_3530_0, i_13_404_3563_0, i_13_404_3570_0,
    i_13_404_3574_0, i_13_404_3767_0, i_13_404_3853_0, i_13_404_3854_0,
    i_13_404_3874_0, i_13_404_3889_0, i_13_404_3890_0, i_13_404_3893_0,
    i_13_404_3939_0, i_13_404_4016_0, i_13_404_4018_0, i_13_404_4055_0,
    i_13_404_4163_0, i_13_404_4232_0, i_13_404_4258_0, i_13_404_4369_0,
    i_13_404_4370_0, i_13_404_4376_0, i_13_404_4565_0, i_13_404_4568_0,
    o_13_404_0_0  );
  input  i_13_404_22_0, i_13_404_59_0, i_13_404_91_0, i_13_404_92_0,
    i_13_404_139_0, i_13_404_215_0, i_13_404_316_0, i_13_404_317_0,
    i_13_404_418_0, i_13_404_419_0, i_13_404_456_0, i_13_404_484_0,
    i_13_404_550_0, i_13_404_554_0, i_13_404_607_0, i_13_404_671_0,
    i_13_404_727_0, i_13_404_793_0, i_13_404_843_0, i_13_404_847_0,
    i_13_404_851_0, i_13_404_860_0, i_13_404_986_0, i_13_404_1018_0,
    i_13_404_1019_0, i_13_404_1083_0, i_13_404_1122_0, i_13_404_1129_0,
    i_13_404_1210_0, i_13_404_1226_0, i_13_404_1256_0, i_13_404_1300_0,
    i_13_404_1301_0, i_13_404_1306_0, i_13_404_1345_0, i_13_404_1361_0,
    i_13_404_1486_0, i_13_404_1487_0, i_13_404_1550_0, i_13_404_1599_0,
    i_13_404_1631_0, i_13_404_1644_0, i_13_404_1721_0, i_13_404_1733_0,
    i_13_404_1763_0, i_13_404_1769_0, i_13_404_1813_0, i_13_404_1855_0,
    i_13_404_1858_0, i_13_404_1859_0, i_13_404_1911_0, i_13_404_2016_0,
    i_13_404_2028_0, i_13_404_2173_0, i_13_404_2179_0, i_13_404_2207_0,
    i_13_404_2290_0, i_13_404_2296_0, i_13_404_2422_0, i_13_404_2450_0,
    i_13_404_2593_0, i_13_404_2615_0, i_13_404_2679_0, i_13_404_2697_0,
    i_13_404_2748_0, i_13_404_2857_0, i_13_404_2981_0, i_13_404_3007_0,
    i_13_404_3008_0, i_13_404_3010_0, i_13_404_3037_0, i_13_404_3110_0,
    i_13_404_3217_0, i_13_404_3389_0, i_13_404_3404_0, i_13_404_3428_0,
    i_13_404_3481_0, i_13_404_3530_0, i_13_404_3563_0, i_13_404_3570_0,
    i_13_404_3574_0, i_13_404_3767_0, i_13_404_3853_0, i_13_404_3854_0,
    i_13_404_3874_0, i_13_404_3889_0, i_13_404_3890_0, i_13_404_3893_0,
    i_13_404_3939_0, i_13_404_4016_0, i_13_404_4018_0, i_13_404_4055_0,
    i_13_404_4163_0, i_13_404_4232_0, i_13_404_4258_0, i_13_404_4369_0,
    i_13_404_4370_0, i_13_404_4376_0, i_13_404_4565_0, i_13_404_4568_0;
  output o_13_404_0_0;
  assign o_13_404_0_0 = ~(~i_13_404_3007_0 | (~i_13_404_92_0 & ~i_13_404_4232_0) | (~i_13_404_316_0 & ~i_13_404_2422_0 & ~i_13_404_3893_0) | (~i_13_404_1550_0 & i_13_404_2422_0 & ~i_13_404_3008_0));
endmodule



// Benchmark "kernel_13_405" written by ABC on Sun Jul 19 10:51:00 2020

module kernel_13_405 ( 
    i_13_405_52_0, i_13_405_78_0, i_13_405_94_0, i_13_405_118_0,
    i_13_405_124_0, i_13_405_142_0, i_13_405_159_0, i_13_405_241_0,
    i_13_405_251_0, i_13_405_259_0, i_13_405_327_0, i_13_405_485_0,
    i_13_405_526_0, i_13_405_552_0, i_13_405_553_0, i_13_405_555_0,
    i_13_405_584_0, i_13_405_591_0, i_13_405_619_0, i_13_405_620_0,
    i_13_405_680_0, i_13_405_713_0, i_13_405_732_0, i_13_405_742_0,
    i_13_405_796_0, i_13_405_943_0, i_13_405_944_0, i_13_405_961_0,
    i_13_405_980_0, i_13_405_1030_0, i_13_405_1078_0, i_13_405_1079_0,
    i_13_405_1249_0, i_13_405_1313_0, i_13_405_1366_0, i_13_405_1403_0,
    i_13_405_1472_0, i_13_405_1502_0, i_13_405_1552_0, i_13_405_1553_0,
    i_13_405_1636_0, i_13_405_1637_0, i_13_405_1661_0, i_13_405_1817_0,
    i_13_405_1951_0, i_13_405_1995_0, i_13_405_2118_0, i_13_405_2211_0,
    i_13_405_2238_0, i_13_405_2321_0, i_13_405_2402_0, i_13_405_2451_0,
    i_13_405_2455_0, i_13_405_2476_0, i_13_405_2555_0, i_13_405_2570_0,
    i_13_405_2596_0, i_13_405_2726_0, i_13_405_2788_0, i_13_405_2789_0,
    i_13_405_2861_0, i_13_405_2888_0, i_13_405_2959_0, i_13_405_3026_0,
    i_13_405_3037_0, i_13_405_3063_0, i_13_405_3207_0, i_13_405_3219_0,
    i_13_405_3373_0, i_13_405_3374_0, i_13_405_3452_0, i_13_405_3464_0,
    i_13_405_3554_0, i_13_405_3571_0, i_13_405_3572_0, i_13_405_3581_0,
    i_13_405_3650_0, i_13_405_3651_0, i_13_405_3689_0, i_13_405_3738_0,
    i_13_405_3894_0, i_13_405_3904_0, i_13_405_3905_0, i_13_405_3938_0,
    i_13_405_4057_0, i_13_405_4091_0, i_13_405_4118_0, i_13_405_4125_0,
    i_13_405_4254_0, i_13_405_4306_0, i_13_405_4318_0, i_13_405_4345_0,
    i_13_405_4364_0, i_13_405_4391_0, i_13_405_4414_0, i_13_405_4415_0,
    i_13_405_4526_0, i_13_405_4534_0, i_13_405_4556_0, i_13_405_4604_0,
    o_13_405_0_0  );
  input  i_13_405_52_0, i_13_405_78_0, i_13_405_94_0, i_13_405_118_0,
    i_13_405_124_0, i_13_405_142_0, i_13_405_159_0, i_13_405_241_0,
    i_13_405_251_0, i_13_405_259_0, i_13_405_327_0, i_13_405_485_0,
    i_13_405_526_0, i_13_405_552_0, i_13_405_553_0, i_13_405_555_0,
    i_13_405_584_0, i_13_405_591_0, i_13_405_619_0, i_13_405_620_0,
    i_13_405_680_0, i_13_405_713_0, i_13_405_732_0, i_13_405_742_0,
    i_13_405_796_0, i_13_405_943_0, i_13_405_944_0, i_13_405_961_0,
    i_13_405_980_0, i_13_405_1030_0, i_13_405_1078_0, i_13_405_1079_0,
    i_13_405_1249_0, i_13_405_1313_0, i_13_405_1366_0, i_13_405_1403_0,
    i_13_405_1472_0, i_13_405_1502_0, i_13_405_1552_0, i_13_405_1553_0,
    i_13_405_1636_0, i_13_405_1637_0, i_13_405_1661_0, i_13_405_1817_0,
    i_13_405_1951_0, i_13_405_1995_0, i_13_405_2118_0, i_13_405_2211_0,
    i_13_405_2238_0, i_13_405_2321_0, i_13_405_2402_0, i_13_405_2451_0,
    i_13_405_2455_0, i_13_405_2476_0, i_13_405_2555_0, i_13_405_2570_0,
    i_13_405_2596_0, i_13_405_2726_0, i_13_405_2788_0, i_13_405_2789_0,
    i_13_405_2861_0, i_13_405_2888_0, i_13_405_2959_0, i_13_405_3026_0,
    i_13_405_3037_0, i_13_405_3063_0, i_13_405_3207_0, i_13_405_3219_0,
    i_13_405_3373_0, i_13_405_3374_0, i_13_405_3452_0, i_13_405_3464_0,
    i_13_405_3554_0, i_13_405_3571_0, i_13_405_3572_0, i_13_405_3581_0,
    i_13_405_3650_0, i_13_405_3651_0, i_13_405_3689_0, i_13_405_3738_0,
    i_13_405_3894_0, i_13_405_3904_0, i_13_405_3905_0, i_13_405_3938_0,
    i_13_405_4057_0, i_13_405_4091_0, i_13_405_4118_0, i_13_405_4125_0,
    i_13_405_4254_0, i_13_405_4306_0, i_13_405_4318_0, i_13_405_4345_0,
    i_13_405_4364_0, i_13_405_4391_0, i_13_405_4414_0, i_13_405_4415_0,
    i_13_405_4526_0, i_13_405_4534_0, i_13_405_4556_0, i_13_405_4604_0;
  output o_13_405_0_0;
  assign o_13_405_0_0 = ~(~i_13_405_620_0);
endmodule



// Benchmark "kernel_13_406" written by ABC on Sun Jul 19 10:51:01 2020

module kernel_13_406 ( 
    i_13_406_76_0, i_13_406_111_0, i_13_406_129_0, i_13_406_179_0,
    i_13_406_266_0, i_13_406_277_0, i_13_406_282_0, i_13_406_283_0,
    i_13_406_302_0, i_13_406_358_0, i_13_406_366_0, i_13_406_471_0,
    i_13_406_472_0, i_13_406_509_0, i_13_406_510_0, i_13_406_545_0,
    i_13_406_591_0, i_13_406_598_0, i_13_406_664_0, i_13_406_726_0,
    i_13_406_799_0, i_13_406_832_0, i_13_406_854_0, i_13_406_862_0,
    i_13_406_894_0, i_13_406_1073_0, i_13_406_1203_0, i_13_406_1212_0,
    i_13_406_1213_0, i_13_406_1307_0, i_13_406_1308_0, i_13_406_1310_0,
    i_13_406_1390_0, i_13_406_1505_0, i_13_406_1623_0, i_13_406_1682_0,
    i_13_406_1698_0, i_13_406_1730_0, i_13_406_2020_0, i_13_406_2023_0,
    i_13_406_2024_0, i_13_406_2059_0, i_13_406_2285_0, i_13_406_2297_0,
    i_13_406_2299_0, i_13_406_2321_0, i_13_406_2445_0, i_13_406_2455_0,
    i_13_406_2456_0, i_13_406_2464_0, i_13_406_2554_0, i_13_406_2650_0,
    i_13_406_2715_0, i_13_406_2716_0, i_13_406_2722_0, i_13_406_2884_0,
    i_13_406_2897_0, i_13_406_2959_0, i_13_406_3046_0, i_13_406_3062_0,
    i_13_406_3076_0, i_13_406_3093_0, i_13_406_3145_0, i_13_406_3253_0,
    i_13_406_3327_0, i_13_406_3329_0, i_13_406_3374_0, i_13_406_3380_0,
    i_13_406_3388_0, i_13_406_3417_0, i_13_406_3418_0, i_13_406_3490_0,
    i_13_406_3550_0, i_13_406_3597_0, i_13_406_3599_0, i_13_406_3635_0,
    i_13_406_3659_0, i_13_406_3764_0, i_13_406_3846_0, i_13_406_3910_0,
    i_13_406_3923_0, i_13_406_3990_0, i_13_406_4119_0, i_13_406_4164_0,
    i_13_406_4192_0, i_13_406_4216_0, i_13_406_4255_0, i_13_406_4265_0,
    i_13_406_4332_0, i_13_406_4333_0, i_13_406_4334_0, i_13_406_4367_0,
    i_13_406_4369_0, i_13_406_4431_0, i_13_406_4433_0, i_13_406_4454_0,
    i_13_406_4461_0, i_13_406_4472_0, i_13_406_4510_0, i_13_406_4512_0,
    o_13_406_0_0  );
  input  i_13_406_76_0, i_13_406_111_0, i_13_406_129_0, i_13_406_179_0,
    i_13_406_266_0, i_13_406_277_0, i_13_406_282_0, i_13_406_283_0,
    i_13_406_302_0, i_13_406_358_0, i_13_406_366_0, i_13_406_471_0,
    i_13_406_472_0, i_13_406_509_0, i_13_406_510_0, i_13_406_545_0,
    i_13_406_591_0, i_13_406_598_0, i_13_406_664_0, i_13_406_726_0,
    i_13_406_799_0, i_13_406_832_0, i_13_406_854_0, i_13_406_862_0,
    i_13_406_894_0, i_13_406_1073_0, i_13_406_1203_0, i_13_406_1212_0,
    i_13_406_1213_0, i_13_406_1307_0, i_13_406_1308_0, i_13_406_1310_0,
    i_13_406_1390_0, i_13_406_1505_0, i_13_406_1623_0, i_13_406_1682_0,
    i_13_406_1698_0, i_13_406_1730_0, i_13_406_2020_0, i_13_406_2023_0,
    i_13_406_2024_0, i_13_406_2059_0, i_13_406_2285_0, i_13_406_2297_0,
    i_13_406_2299_0, i_13_406_2321_0, i_13_406_2445_0, i_13_406_2455_0,
    i_13_406_2456_0, i_13_406_2464_0, i_13_406_2554_0, i_13_406_2650_0,
    i_13_406_2715_0, i_13_406_2716_0, i_13_406_2722_0, i_13_406_2884_0,
    i_13_406_2897_0, i_13_406_2959_0, i_13_406_3046_0, i_13_406_3062_0,
    i_13_406_3076_0, i_13_406_3093_0, i_13_406_3145_0, i_13_406_3253_0,
    i_13_406_3327_0, i_13_406_3329_0, i_13_406_3374_0, i_13_406_3380_0,
    i_13_406_3388_0, i_13_406_3417_0, i_13_406_3418_0, i_13_406_3490_0,
    i_13_406_3550_0, i_13_406_3597_0, i_13_406_3599_0, i_13_406_3635_0,
    i_13_406_3659_0, i_13_406_3764_0, i_13_406_3846_0, i_13_406_3910_0,
    i_13_406_3923_0, i_13_406_3990_0, i_13_406_4119_0, i_13_406_4164_0,
    i_13_406_4192_0, i_13_406_4216_0, i_13_406_4255_0, i_13_406_4265_0,
    i_13_406_4332_0, i_13_406_4333_0, i_13_406_4334_0, i_13_406_4367_0,
    i_13_406_4369_0, i_13_406_4431_0, i_13_406_4433_0, i_13_406_4454_0,
    i_13_406_4461_0, i_13_406_4472_0, i_13_406_4510_0, i_13_406_4512_0;
  output o_13_406_0_0;
  assign o_13_406_0_0 = ~((~i_13_406_277_0 & ((i_13_406_1310_0 & ~i_13_406_4334_0 & ~i_13_406_4510_0) | (~i_13_406_832_0 & ~i_13_406_4333_0 & ~i_13_406_4512_0))) | (~i_13_406_472_0 & ((~i_13_406_894_0 & ~i_13_406_3062_0 & ~i_13_406_3846_0 & ~i_13_406_4255_0 & ~i_13_406_4334_0 & ~i_13_406_4433_0) | (~i_13_406_2884_0 & ~i_13_406_4510_0))) | (~i_13_406_4334_0 & ((~i_13_406_1203_0 & i_13_406_3910_0 & ~i_13_406_4255_0 & ~i_13_406_4431_0) | (i_13_406_3388_0 & ~i_13_406_4512_0))) | (~i_13_406_832_0 & ~i_13_406_3093_0 & ~i_13_406_3910_0));
endmodule



// Benchmark "kernel_13_407" written by ABC on Sun Jul 19 10:51:02 2020

module kernel_13_407 ( 
    i_13_407_19_0, i_13_407_64_0, i_13_407_111_0, i_13_407_165_0,
    i_13_407_166_0, i_13_407_237_0, i_13_407_325_0, i_13_407_336_0,
    i_13_407_450_0, i_13_407_495_0, i_13_407_585_0, i_13_407_615_0,
    i_13_407_639_0, i_13_407_756_0, i_13_407_811_0, i_13_407_813_0,
    i_13_407_855_0, i_13_407_882_0, i_13_407_984_0, i_13_407_1062_0,
    i_13_407_1063_0, i_13_407_1216_0, i_13_407_1219_0, i_13_407_1251_0,
    i_13_407_1395_0, i_13_407_1458_0, i_13_407_1503_0, i_13_407_1513_0,
    i_13_407_1524_0, i_13_407_1608_0, i_13_407_1714_0, i_13_407_1848_0,
    i_13_407_1927_0, i_13_407_1990_0, i_13_407_2052_0, i_13_407_2053_0,
    i_13_407_2107_0, i_13_407_2116_0, i_13_407_2124_0, i_13_407_2127_0,
    i_13_407_2133_0, i_13_407_2134_0, i_13_407_2136_0, i_13_407_2145_0,
    i_13_407_2172_0, i_13_407_2233_0, i_13_407_2259_0, i_13_407_2260_0,
    i_13_407_2277_0, i_13_407_2278_0, i_13_407_2340_0, i_13_407_2364_0,
    i_13_407_2403_0, i_13_407_2404_0, i_13_407_2520_0, i_13_407_2614_0,
    i_13_407_2709_0, i_13_407_2713_0, i_13_407_2745_0, i_13_407_2757_0,
    i_13_407_2781_0, i_13_407_2934_0, i_13_407_2937_0, i_13_407_2938_0,
    i_13_407_3010_0, i_13_407_3024_0, i_13_407_3127_0, i_13_407_3339_0,
    i_13_407_3376_0, i_13_407_3394_0, i_13_407_3612_0, i_13_407_3627_0,
    i_13_407_3628_0, i_13_407_3639_0, i_13_407_3663_0, i_13_407_3703_0,
    i_13_407_3708_0, i_13_407_3738_0, i_13_407_3739_0, i_13_407_3793_0,
    i_13_407_3817_0, i_13_407_3891_0, i_13_407_4017_0, i_13_407_4059_0,
    i_13_407_4060_0, i_13_407_4062_0, i_13_407_4086_0, i_13_407_4102_0,
    i_13_407_4267_0, i_13_407_4276_0, i_13_407_4303_0, i_13_407_4315_0,
    i_13_407_4329_0, i_13_407_4338_0, i_13_407_4377_0, i_13_407_4392_0,
    i_13_407_4446_0, i_13_407_4447_0, i_13_407_4530_0, i_13_407_4568_0,
    o_13_407_0_0  );
  input  i_13_407_19_0, i_13_407_64_0, i_13_407_111_0, i_13_407_165_0,
    i_13_407_166_0, i_13_407_237_0, i_13_407_325_0, i_13_407_336_0,
    i_13_407_450_0, i_13_407_495_0, i_13_407_585_0, i_13_407_615_0,
    i_13_407_639_0, i_13_407_756_0, i_13_407_811_0, i_13_407_813_0,
    i_13_407_855_0, i_13_407_882_0, i_13_407_984_0, i_13_407_1062_0,
    i_13_407_1063_0, i_13_407_1216_0, i_13_407_1219_0, i_13_407_1251_0,
    i_13_407_1395_0, i_13_407_1458_0, i_13_407_1503_0, i_13_407_1513_0,
    i_13_407_1524_0, i_13_407_1608_0, i_13_407_1714_0, i_13_407_1848_0,
    i_13_407_1927_0, i_13_407_1990_0, i_13_407_2052_0, i_13_407_2053_0,
    i_13_407_2107_0, i_13_407_2116_0, i_13_407_2124_0, i_13_407_2127_0,
    i_13_407_2133_0, i_13_407_2134_0, i_13_407_2136_0, i_13_407_2145_0,
    i_13_407_2172_0, i_13_407_2233_0, i_13_407_2259_0, i_13_407_2260_0,
    i_13_407_2277_0, i_13_407_2278_0, i_13_407_2340_0, i_13_407_2364_0,
    i_13_407_2403_0, i_13_407_2404_0, i_13_407_2520_0, i_13_407_2614_0,
    i_13_407_2709_0, i_13_407_2713_0, i_13_407_2745_0, i_13_407_2757_0,
    i_13_407_2781_0, i_13_407_2934_0, i_13_407_2937_0, i_13_407_2938_0,
    i_13_407_3010_0, i_13_407_3024_0, i_13_407_3127_0, i_13_407_3339_0,
    i_13_407_3376_0, i_13_407_3394_0, i_13_407_3612_0, i_13_407_3627_0,
    i_13_407_3628_0, i_13_407_3639_0, i_13_407_3663_0, i_13_407_3703_0,
    i_13_407_3708_0, i_13_407_3738_0, i_13_407_3739_0, i_13_407_3793_0,
    i_13_407_3817_0, i_13_407_3891_0, i_13_407_4017_0, i_13_407_4059_0,
    i_13_407_4060_0, i_13_407_4062_0, i_13_407_4086_0, i_13_407_4102_0,
    i_13_407_4267_0, i_13_407_4276_0, i_13_407_4303_0, i_13_407_4315_0,
    i_13_407_4329_0, i_13_407_4338_0, i_13_407_4377_0, i_13_407_4392_0,
    i_13_407_4446_0, i_13_407_4447_0, i_13_407_4530_0, i_13_407_4568_0;
  output o_13_407_0_0;
  assign o_13_407_0_0 = ~((~i_13_407_2403_0 & i_13_407_4329_0) | (~i_13_407_1062_0 & ~i_13_407_4059_0));
endmodule



// Benchmark "kernel_13_408" written by ABC on Sun Jul 19 10:51:03 2020

module kernel_13_408 ( 
    i_13_408_64_0, i_13_408_97_0, i_13_408_121_0, i_13_408_131_0,
    i_13_408_158_0, i_13_408_208_0, i_13_408_236_0, i_13_408_245_0,
    i_13_408_251_0, i_13_408_415_0, i_13_408_416_0, i_13_408_463_0,
    i_13_408_464_0, i_13_408_571_0, i_13_408_589_0, i_13_408_596_0,
    i_13_408_761_0, i_13_408_829_0, i_13_408_1073_0, i_13_408_1129_0,
    i_13_408_1207_0, i_13_408_1211_0, i_13_408_1318_0, i_13_408_1346_0,
    i_13_408_1361_0, i_13_408_1466_0, i_13_408_1510_0, i_13_408_1511_0,
    i_13_408_1522_0, i_13_408_1550_0, i_13_408_1570_0, i_13_408_1604_0,
    i_13_408_1640_0, i_13_408_1696_0, i_13_408_1697_0, i_13_408_1700_0,
    i_13_408_1751_0, i_13_408_1840_0, i_13_408_1847_0, i_13_408_1853_0,
    i_13_408_1874_0, i_13_408_1928_0, i_13_408_1958_0, i_13_408_1964_0,
    i_13_408_1994_0, i_13_408_2057_0, i_13_408_2101_0, i_13_408_2102_0,
    i_13_408_2143_0, i_13_408_2200_0, i_13_408_2201_0, i_13_408_2209_0,
    i_13_408_2297_0, i_13_408_2315_0, i_13_408_2434_0, i_13_408_2444_0,
    i_13_408_2551_0, i_13_408_2612_0, i_13_408_2798_0, i_13_408_2881_0,
    i_13_408_2936_0, i_13_408_2939_0, i_13_408_3056_0, i_13_408_3113_0,
    i_13_408_3143_0, i_13_408_3208_0, i_13_408_3242_0, i_13_408_3254_0,
    i_13_408_3347_0, i_13_408_3370_0, i_13_408_3388_0, i_13_408_3458_0,
    i_13_408_3551_0, i_13_408_3596_0, i_13_408_3610_0, i_13_408_3619_0,
    i_13_408_3632_0, i_13_408_3637_0, i_13_408_3638_0, i_13_408_3667_0,
    i_13_408_3704_0, i_13_408_3766_0, i_13_408_3844_0, i_13_408_3857_0,
    i_13_408_3916_0, i_13_408_3935_0, i_13_408_4009_0, i_13_408_4019_0,
    i_13_408_4037_0, i_13_408_4045_0, i_13_408_4105_0, i_13_408_4208_0,
    i_13_408_4214_0, i_13_408_4330_0, i_13_408_4378_0, i_13_408_4430_0,
    i_13_408_4451_0, i_13_408_4510_0, i_13_408_4559_0, i_13_408_4582_0,
    o_13_408_0_0  );
  input  i_13_408_64_0, i_13_408_97_0, i_13_408_121_0, i_13_408_131_0,
    i_13_408_158_0, i_13_408_208_0, i_13_408_236_0, i_13_408_245_0,
    i_13_408_251_0, i_13_408_415_0, i_13_408_416_0, i_13_408_463_0,
    i_13_408_464_0, i_13_408_571_0, i_13_408_589_0, i_13_408_596_0,
    i_13_408_761_0, i_13_408_829_0, i_13_408_1073_0, i_13_408_1129_0,
    i_13_408_1207_0, i_13_408_1211_0, i_13_408_1318_0, i_13_408_1346_0,
    i_13_408_1361_0, i_13_408_1466_0, i_13_408_1510_0, i_13_408_1511_0,
    i_13_408_1522_0, i_13_408_1550_0, i_13_408_1570_0, i_13_408_1604_0,
    i_13_408_1640_0, i_13_408_1696_0, i_13_408_1697_0, i_13_408_1700_0,
    i_13_408_1751_0, i_13_408_1840_0, i_13_408_1847_0, i_13_408_1853_0,
    i_13_408_1874_0, i_13_408_1928_0, i_13_408_1958_0, i_13_408_1964_0,
    i_13_408_1994_0, i_13_408_2057_0, i_13_408_2101_0, i_13_408_2102_0,
    i_13_408_2143_0, i_13_408_2200_0, i_13_408_2201_0, i_13_408_2209_0,
    i_13_408_2297_0, i_13_408_2315_0, i_13_408_2434_0, i_13_408_2444_0,
    i_13_408_2551_0, i_13_408_2612_0, i_13_408_2798_0, i_13_408_2881_0,
    i_13_408_2936_0, i_13_408_2939_0, i_13_408_3056_0, i_13_408_3113_0,
    i_13_408_3143_0, i_13_408_3208_0, i_13_408_3242_0, i_13_408_3254_0,
    i_13_408_3347_0, i_13_408_3370_0, i_13_408_3388_0, i_13_408_3458_0,
    i_13_408_3551_0, i_13_408_3596_0, i_13_408_3610_0, i_13_408_3619_0,
    i_13_408_3632_0, i_13_408_3637_0, i_13_408_3638_0, i_13_408_3667_0,
    i_13_408_3704_0, i_13_408_3766_0, i_13_408_3844_0, i_13_408_3857_0,
    i_13_408_3916_0, i_13_408_3935_0, i_13_408_4009_0, i_13_408_4019_0,
    i_13_408_4037_0, i_13_408_4045_0, i_13_408_4105_0, i_13_408_4208_0,
    i_13_408_4214_0, i_13_408_4330_0, i_13_408_4378_0, i_13_408_4430_0,
    i_13_408_4451_0, i_13_408_4510_0, i_13_408_4559_0, i_13_408_4582_0;
  output o_13_408_0_0;
  assign o_13_408_0_0 = ~(~i_13_408_1522_0 | (~i_13_408_1346_0 & ~i_13_408_1751_0));
endmodule



// Benchmark "kernel_13_409" written by ABC on Sun Jul 19 10:51:03 2020

module kernel_13_409 ( 
    i_13_409_20_0, i_13_409_91_0, i_13_409_92_0, i_13_409_100_0,
    i_13_409_155_0, i_13_409_166_0, i_13_409_169_0, i_13_409_174_0,
    i_13_409_203_0, i_13_409_280_0, i_13_409_284_0, i_13_409_316_0,
    i_13_409_381_0, i_13_409_490_0, i_13_409_517_0, i_13_409_571_0,
    i_13_409_607_0, i_13_409_697_0, i_13_409_931_0, i_13_409_1021_0,
    i_13_409_1063_0, i_13_409_1064_0, i_13_409_1066_0, i_13_409_1092_0,
    i_13_409_1093_0, i_13_409_1219_0, i_13_409_1268_0, i_13_409_1324_0,
    i_13_409_1364_0, i_13_409_1440_0, i_13_409_1496_0, i_13_409_1528_0,
    i_13_409_1570_0, i_13_409_1747_0, i_13_409_1810_0, i_13_409_1829_0,
    i_13_409_1848_0, i_13_409_1849_0, i_13_409_1870_0, i_13_409_1885_0,
    i_13_409_1909_0, i_13_409_2053_0, i_13_409_2107_0, i_13_409_2108_0,
    i_13_409_2116_0, i_13_409_2117_0, i_13_409_2233_0, i_13_409_2234_0,
    i_13_409_2260_0, i_13_409_2274_0, i_13_409_2332_0, i_13_409_2333_0,
    i_13_409_2396_0, i_13_409_2404_0, i_13_409_2406_0, i_13_409_2443_0,
    i_13_409_2597_0, i_13_409_2624_0, i_13_409_2701_0, i_13_409_2790_0,
    i_13_409_2793_0, i_13_409_2848_0, i_13_409_2853_0, i_13_409_2872_0,
    i_13_409_2935_0, i_13_409_2938_0, i_13_409_2980_0, i_13_409_3007_0,
    i_13_409_3089_0, i_13_409_3109_0, i_13_409_3143_0, i_13_409_3205_0,
    i_13_409_3339_0, i_13_409_3352_0, i_13_409_3397_0, i_13_409_3541_0,
    i_13_409_3603_0, i_13_409_3733_0, i_13_409_3739_0, i_13_409_3742_0,
    i_13_409_3764_0, i_13_409_3766_0, i_13_409_3816_0, i_13_409_3817_0,
    i_13_409_3818_0, i_13_409_3870_0, i_13_409_4012_0, i_13_409_4016_0,
    i_13_409_4018_0, i_13_409_4059_0, i_13_409_4060_0, i_13_409_4061_0,
    i_13_409_4062_0, i_13_409_4063_0, i_13_409_4143_0, i_13_409_4259_0,
    i_13_409_4267_0, i_13_409_4315_0, i_13_409_4352_0, i_13_409_4567_0,
    o_13_409_0_0  );
  input  i_13_409_20_0, i_13_409_91_0, i_13_409_92_0, i_13_409_100_0,
    i_13_409_155_0, i_13_409_166_0, i_13_409_169_0, i_13_409_174_0,
    i_13_409_203_0, i_13_409_280_0, i_13_409_284_0, i_13_409_316_0,
    i_13_409_381_0, i_13_409_490_0, i_13_409_517_0, i_13_409_571_0,
    i_13_409_607_0, i_13_409_697_0, i_13_409_931_0, i_13_409_1021_0,
    i_13_409_1063_0, i_13_409_1064_0, i_13_409_1066_0, i_13_409_1092_0,
    i_13_409_1093_0, i_13_409_1219_0, i_13_409_1268_0, i_13_409_1324_0,
    i_13_409_1364_0, i_13_409_1440_0, i_13_409_1496_0, i_13_409_1528_0,
    i_13_409_1570_0, i_13_409_1747_0, i_13_409_1810_0, i_13_409_1829_0,
    i_13_409_1848_0, i_13_409_1849_0, i_13_409_1870_0, i_13_409_1885_0,
    i_13_409_1909_0, i_13_409_2053_0, i_13_409_2107_0, i_13_409_2108_0,
    i_13_409_2116_0, i_13_409_2117_0, i_13_409_2233_0, i_13_409_2234_0,
    i_13_409_2260_0, i_13_409_2274_0, i_13_409_2332_0, i_13_409_2333_0,
    i_13_409_2396_0, i_13_409_2404_0, i_13_409_2406_0, i_13_409_2443_0,
    i_13_409_2597_0, i_13_409_2624_0, i_13_409_2701_0, i_13_409_2790_0,
    i_13_409_2793_0, i_13_409_2848_0, i_13_409_2853_0, i_13_409_2872_0,
    i_13_409_2935_0, i_13_409_2938_0, i_13_409_2980_0, i_13_409_3007_0,
    i_13_409_3089_0, i_13_409_3109_0, i_13_409_3143_0, i_13_409_3205_0,
    i_13_409_3339_0, i_13_409_3352_0, i_13_409_3397_0, i_13_409_3541_0,
    i_13_409_3603_0, i_13_409_3733_0, i_13_409_3739_0, i_13_409_3742_0,
    i_13_409_3764_0, i_13_409_3766_0, i_13_409_3816_0, i_13_409_3817_0,
    i_13_409_3818_0, i_13_409_3870_0, i_13_409_4012_0, i_13_409_4016_0,
    i_13_409_4018_0, i_13_409_4059_0, i_13_409_4060_0, i_13_409_4061_0,
    i_13_409_4062_0, i_13_409_4063_0, i_13_409_4143_0, i_13_409_4259_0,
    i_13_409_4267_0, i_13_409_4315_0, i_13_409_4352_0, i_13_409_4567_0;
  output o_13_409_0_0;
  assign o_13_409_0_0 = ~((i_13_409_3739_0 & ~i_13_409_4267_0) | (~i_13_409_1324_0 & ~i_13_409_3764_0) | (~i_13_409_1849_0 & ~i_13_409_2234_0 & ~i_13_409_3817_0));
endmodule



// Benchmark "kernel_13_410" written by ABC on Sun Jul 19 10:51:04 2020

module kernel_13_410 ( 
    i_13_410_18_0, i_13_410_34_0, i_13_410_45_0, i_13_410_67_0,
    i_13_410_70_0, i_13_410_94_0, i_13_410_128_0, i_13_410_129_0,
    i_13_410_156_0, i_13_410_157_0, i_13_410_160_0, i_13_410_218_0,
    i_13_410_222_0, i_13_410_275_0, i_13_410_333_0, i_13_410_385_0,
    i_13_410_409_0, i_13_410_473_0, i_13_410_490_0, i_13_410_493_0,
    i_13_410_615_0, i_13_410_643_0, i_13_410_644_0, i_13_410_737_0,
    i_13_410_738_0, i_13_410_741_0, i_13_410_742_0, i_13_410_745_0,
    i_13_410_829_0, i_13_410_841_0, i_13_410_934_0, i_13_410_950_0,
    i_13_410_956_0, i_13_410_1120_0, i_13_410_1211_0, i_13_410_1263_0,
    i_13_410_1300_0, i_13_410_1302_0, i_13_410_1395_0, i_13_410_1447_0,
    i_13_410_1522_0, i_13_410_1570_0, i_13_410_1605_0, i_13_410_1720_0,
    i_13_410_1760_0, i_13_410_1815_0, i_13_410_1847_0, i_13_410_1903_0,
    i_13_410_1939_0, i_13_410_2002_0, i_13_410_2007_0, i_13_410_2021_0,
    i_13_410_2101_0, i_13_410_2142_0, i_13_410_2154_0, i_13_410_2193_0,
    i_13_410_2235_0, i_13_410_2242_0, i_13_410_2297_0, i_13_410_2397_0,
    i_13_410_2584_0, i_13_410_2620_0, i_13_410_2676_0, i_13_410_2695_0,
    i_13_410_2781_0, i_13_410_2891_0, i_13_410_2998_0, i_13_410_3033_0,
    i_13_410_3213_0, i_13_410_3217_0, i_13_410_3240_0, i_13_410_3241_0,
    i_13_410_3242_0, i_13_410_3265_0, i_13_410_3531_0, i_13_410_3599_0,
    i_13_410_3618_0, i_13_410_3636_0, i_13_410_3637_0, i_13_410_3692_0,
    i_13_410_3702_0, i_13_410_3723_0, i_13_410_3766_0, i_13_410_3843_0,
    i_13_410_3846_0, i_13_410_3847_0, i_13_410_3876_0, i_13_410_3892_0,
    i_13_410_3915_0, i_13_410_3982_0, i_13_410_3985_0, i_13_410_4081_0,
    i_13_410_4117_0, i_13_410_4214_0, i_13_410_4273_0, i_13_410_4281_0,
    i_13_410_4327_0, i_13_410_4352_0, i_13_410_4461_0, i_13_410_4509_0,
    o_13_410_0_0  );
  input  i_13_410_18_0, i_13_410_34_0, i_13_410_45_0, i_13_410_67_0,
    i_13_410_70_0, i_13_410_94_0, i_13_410_128_0, i_13_410_129_0,
    i_13_410_156_0, i_13_410_157_0, i_13_410_160_0, i_13_410_218_0,
    i_13_410_222_0, i_13_410_275_0, i_13_410_333_0, i_13_410_385_0,
    i_13_410_409_0, i_13_410_473_0, i_13_410_490_0, i_13_410_493_0,
    i_13_410_615_0, i_13_410_643_0, i_13_410_644_0, i_13_410_737_0,
    i_13_410_738_0, i_13_410_741_0, i_13_410_742_0, i_13_410_745_0,
    i_13_410_829_0, i_13_410_841_0, i_13_410_934_0, i_13_410_950_0,
    i_13_410_956_0, i_13_410_1120_0, i_13_410_1211_0, i_13_410_1263_0,
    i_13_410_1300_0, i_13_410_1302_0, i_13_410_1395_0, i_13_410_1447_0,
    i_13_410_1522_0, i_13_410_1570_0, i_13_410_1605_0, i_13_410_1720_0,
    i_13_410_1760_0, i_13_410_1815_0, i_13_410_1847_0, i_13_410_1903_0,
    i_13_410_1939_0, i_13_410_2002_0, i_13_410_2007_0, i_13_410_2021_0,
    i_13_410_2101_0, i_13_410_2142_0, i_13_410_2154_0, i_13_410_2193_0,
    i_13_410_2235_0, i_13_410_2242_0, i_13_410_2297_0, i_13_410_2397_0,
    i_13_410_2584_0, i_13_410_2620_0, i_13_410_2676_0, i_13_410_2695_0,
    i_13_410_2781_0, i_13_410_2891_0, i_13_410_2998_0, i_13_410_3033_0,
    i_13_410_3213_0, i_13_410_3217_0, i_13_410_3240_0, i_13_410_3241_0,
    i_13_410_3242_0, i_13_410_3265_0, i_13_410_3531_0, i_13_410_3599_0,
    i_13_410_3618_0, i_13_410_3636_0, i_13_410_3637_0, i_13_410_3692_0,
    i_13_410_3702_0, i_13_410_3723_0, i_13_410_3766_0, i_13_410_3843_0,
    i_13_410_3846_0, i_13_410_3847_0, i_13_410_3876_0, i_13_410_3892_0,
    i_13_410_3915_0, i_13_410_3982_0, i_13_410_3985_0, i_13_410_4081_0,
    i_13_410_4117_0, i_13_410_4214_0, i_13_410_4273_0, i_13_410_4281_0,
    i_13_410_4327_0, i_13_410_4352_0, i_13_410_4461_0, i_13_410_4509_0;
  output o_13_410_0_0;
  assign o_13_410_0_0 = ~((~i_13_410_34_0 & ((i_13_410_841_0 & i_13_410_2695_0 & ~i_13_410_3240_0 & ~i_13_410_3876_0) | (~i_13_410_275_0 & ~i_13_410_1522_0 & ~i_13_410_3213_0 & ~i_13_410_3241_0 & ~i_13_410_3265_0 & ~i_13_410_3892_0 & i_13_410_4081_0))) | (~i_13_410_2002_0 & ((~i_13_410_1263_0 & ~i_13_410_3847_0 & ~i_13_410_3985_0) | (~i_13_410_3982_0 & ~i_13_410_4327_0))) | (~i_13_410_1263_0 & ~i_13_410_4081_0 & ((~i_13_410_1211_0 & i_13_410_1300_0 & ~i_13_410_2242_0) | (~i_13_410_950_0 & ~i_13_410_4214_0 & ~i_13_410_4273_0))) | (~i_13_410_3531_0 & ((~i_13_410_490_0 & ~i_13_410_934_0 & ~i_13_410_1815_0 & ~i_13_410_3846_0) | (i_13_410_841_0 & ~i_13_410_4273_0 & ~i_13_410_4509_0))) | (i_13_410_4352_0 & (~i_13_410_94_0 | (~i_13_410_3847_0 & ~i_13_410_4214_0))) | (~i_13_410_737_0 & ~i_13_410_1302_0 & ~i_13_410_1847_0 & ~i_13_410_3982_0) | (i_13_410_2695_0 & i_13_410_3985_0 & ~i_13_410_4273_0 & ~i_13_410_4327_0));
endmodule



// Benchmark "kernel_13_411" written by ABC on Sun Jul 19 10:51:05 2020

module kernel_13_411 ( 
    i_13_411_112_0, i_13_411_119_0, i_13_411_124_0, i_13_411_125_0,
    i_13_411_142_0, i_13_411_197_0, i_13_411_208_0, i_13_411_241_0,
    i_13_411_277_0, i_13_411_319_0, i_13_411_337_0, i_13_411_377_0,
    i_13_411_416_0, i_13_411_454_0, i_13_411_562_0, i_13_411_565_0,
    i_13_411_646_0, i_13_411_665_0, i_13_411_727_0, i_13_411_733_0,
    i_13_411_857_0, i_13_411_931_0, i_13_411_943_0, i_13_411_953_0,
    i_13_411_1019_0, i_13_411_1085_0, i_13_411_1225_0, i_13_411_1301_0,
    i_13_411_1302_0, i_13_411_1345_0, i_13_411_1375_0, i_13_411_1486_0,
    i_13_411_1487_0, i_13_411_1529_0, i_13_411_1627_0, i_13_411_1631_0,
    i_13_411_1726_0, i_13_411_1768_0, i_13_411_1787_0, i_13_411_1844_0,
    i_13_411_2015_0, i_13_411_2206_0, i_13_411_2212_0, i_13_411_2237_0,
    i_13_411_2438_0, i_13_411_2546_0, i_13_411_2618_0, i_13_411_2653_0,
    i_13_411_2680_0, i_13_411_2825_0, i_13_411_2917_0, i_13_411_2918_0,
    i_13_411_2920_0, i_13_411_3011_0, i_13_411_3020_0, i_13_411_3040_0,
    i_13_411_3113_0, i_13_411_3161_0, i_13_411_3167_0, i_13_411_3170_0,
    i_13_411_3212_0, i_13_411_3215_0, i_13_411_3217_0, i_13_411_3218_0,
    i_13_411_3238_0, i_13_411_3261_0, i_13_411_3328_0, i_13_411_3391_0,
    i_13_411_3421_0, i_13_411_3422_0, i_13_411_3463_0, i_13_411_3535_0,
    i_13_411_3536_0, i_13_411_3553_0, i_13_411_3644_0, i_13_411_3688_0,
    i_13_411_3689_0, i_13_411_3700_0, i_13_411_3781_0, i_13_411_3799_0,
    i_13_411_3821_0, i_13_411_3850_0, i_13_411_3872_0, i_13_411_3877_0,
    i_13_411_3878_0, i_13_411_3890_0, i_13_411_3898_0, i_13_411_3907_0,
    i_13_411_3983_0, i_13_411_3991_0, i_13_411_4012_0, i_13_411_4066_0,
    i_13_411_4067_0, i_13_411_4090_0, i_13_411_4270_0, i_13_411_4346_0,
    i_13_411_4534_0, i_13_411_4535_0, i_13_411_4543_0, i_13_411_4594_0,
    o_13_411_0_0  );
  input  i_13_411_112_0, i_13_411_119_0, i_13_411_124_0, i_13_411_125_0,
    i_13_411_142_0, i_13_411_197_0, i_13_411_208_0, i_13_411_241_0,
    i_13_411_277_0, i_13_411_319_0, i_13_411_337_0, i_13_411_377_0,
    i_13_411_416_0, i_13_411_454_0, i_13_411_562_0, i_13_411_565_0,
    i_13_411_646_0, i_13_411_665_0, i_13_411_727_0, i_13_411_733_0,
    i_13_411_857_0, i_13_411_931_0, i_13_411_943_0, i_13_411_953_0,
    i_13_411_1019_0, i_13_411_1085_0, i_13_411_1225_0, i_13_411_1301_0,
    i_13_411_1302_0, i_13_411_1345_0, i_13_411_1375_0, i_13_411_1486_0,
    i_13_411_1487_0, i_13_411_1529_0, i_13_411_1627_0, i_13_411_1631_0,
    i_13_411_1726_0, i_13_411_1768_0, i_13_411_1787_0, i_13_411_1844_0,
    i_13_411_2015_0, i_13_411_2206_0, i_13_411_2212_0, i_13_411_2237_0,
    i_13_411_2438_0, i_13_411_2546_0, i_13_411_2618_0, i_13_411_2653_0,
    i_13_411_2680_0, i_13_411_2825_0, i_13_411_2917_0, i_13_411_2918_0,
    i_13_411_2920_0, i_13_411_3011_0, i_13_411_3020_0, i_13_411_3040_0,
    i_13_411_3113_0, i_13_411_3161_0, i_13_411_3167_0, i_13_411_3170_0,
    i_13_411_3212_0, i_13_411_3215_0, i_13_411_3217_0, i_13_411_3218_0,
    i_13_411_3238_0, i_13_411_3261_0, i_13_411_3328_0, i_13_411_3391_0,
    i_13_411_3421_0, i_13_411_3422_0, i_13_411_3463_0, i_13_411_3535_0,
    i_13_411_3536_0, i_13_411_3553_0, i_13_411_3644_0, i_13_411_3688_0,
    i_13_411_3689_0, i_13_411_3700_0, i_13_411_3781_0, i_13_411_3799_0,
    i_13_411_3821_0, i_13_411_3850_0, i_13_411_3872_0, i_13_411_3877_0,
    i_13_411_3878_0, i_13_411_3890_0, i_13_411_3898_0, i_13_411_3907_0,
    i_13_411_3983_0, i_13_411_3991_0, i_13_411_4012_0, i_13_411_4066_0,
    i_13_411_4067_0, i_13_411_4090_0, i_13_411_4270_0, i_13_411_4346_0,
    i_13_411_4534_0, i_13_411_4535_0, i_13_411_4543_0, i_13_411_4594_0;
  output o_13_411_0_0;
  assign o_13_411_0_0 = ~((~i_13_411_3535_0 & ~i_13_411_3688_0) | (~i_13_411_277_0 & ~i_13_411_3218_0) | (~i_13_411_197_0 & ~i_13_411_2212_0 & ~i_13_411_3689_0) | (~i_13_411_1085_0 & ~i_13_411_1627_0 & i_13_411_1768_0) | (~i_13_411_112_0 & ~i_13_411_241_0 & ~i_13_411_953_0));
endmodule



// Benchmark "kernel_13_412" written by ABC on Sun Jul 19 10:51:06 2020

module kernel_13_412 ( 
    i_13_412_70_0, i_13_412_174_0, i_13_412_326_0, i_13_412_355_0,
    i_13_412_409_0, i_13_412_522_0, i_13_412_527_0, i_13_412_561_0,
    i_13_412_661_0, i_13_412_663_0, i_13_412_762_0, i_13_412_796_0,
    i_13_412_822_0, i_13_412_826_0, i_13_412_850_0, i_13_412_851_0,
    i_13_412_853_0, i_13_412_887_0, i_13_412_940_0, i_13_412_952_0,
    i_13_412_1020_0, i_13_412_1023_0, i_13_412_1075_0, i_13_412_1077_0,
    i_13_412_1186_0, i_13_412_1224_0, i_13_412_1227_0, i_13_412_1228_0,
    i_13_412_1230_0, i_13_412_1255_0, i_13_412_1275_0, i_13_412_1279_0,
    i_13_412_1303_0, i_13_412_1312_0, i_13_412_1317_0, i_13_412_1321_0,
    i_13_412_1345_0, i_13_412_1498_0, i_13_412_1551_0, i_13_412_1552_0,
    i_13_412_1570_0, i_13_412_1770_0, i_13_412_1780_0, i_13_412_1798_0,
    i_13_412_1854_0, i_13_412_1858_0, i_13_412_1860_0, i_13_412_1956_0,
    i_13_412_1957_0, i_13_412_2056_0, i_13_412_2110_0, i_13_412_2265_0,
    i_13_412_2281_0, i_13_412_2366_0, i_13_412_2452_0, i_13_412_2454_0,
    i_13_412_2460_0, i_13_412_2473_0, i_13_412_2505_0, i_13_412_2539_0,
    i_13_412_2541_0, i_13_412_2613_0, i_13_412_2622_0, i_13_412_2647_0,
    i_13_412_3031_0, i_13_412_3100_0, i_13_412_3120_0, i_13_412_3170_0,
    i_13_412_3172_0, i_13_412_3273_0, i_13_412_3381_0, i_13_412_3427_0,
    i_13_412_3429_0, i_13_412_3460_0, i_13_412_3468_0, i_13_412_3483_0,
    i_13_412_3503_0, i_13_412_3505_0, i_13_412_3541_0, i_13_412_3559_0,
    i_13_412_3570_0, i_13_412_3651_0, i_13_412_3729_0, i_13_412_3783_0,
    i_13_412_3822_0, i_13_412_3829_0, i_13_412_3856_0, i_13_412_3896_0,
    i_13_412_3910_0, i_13_412_3911_0, i_13_412_4252_0, i_13_412_4254_0,
    i_13_412_4256_0, i_13_412_4261_0, i_13_412_4377_0, i_13_412_4396_0,
    i_13_412_4415_0, i_13_412_4579_0, i_13_412_4597_0, i_13_412_4606_0,
    o_13_412_0_0  );
  input  i_13_412_70_0, i_13_412_174_0, i_13_412_326_0, i_13_412_355_0,
    i_13_412_409_0, i_13_412_522_0, i_13_412_527_0, i_13_412_561_0,
    i_13_412_661_0, i_13_412_663_0, i_13_412_762_0, i_13_412_796_0,
    i_13_412_822_0, i_13_412_826_0, i_13_412_850_0, i_13_412_851_0,
    i_13_412_853_0, i_13_412_887_0, i_13_412_940_0, i_13_412_952_0,
    i_13_412_1020_0, i_13_412_1023_0, i_13_412_1075_0, i_13_412_1077_0,
    i_13_412_1186_0, i_13_412_1224_0, i_13_412_1227_0, i_13_412_1228_0,
    i_13_412_1230_0, i_13_412_1255_0, i_13_412_1275_0, i_13_412_1279_0,
    i_13_412_1303_0, i_13_412_1312_0, i_13_412_1317_0, i_13_412_1321_0,
    i_13_412_1345_0, i_13_412_1498_0, i_13_412_1551_0, i_13_412_1552_0,
    i_13_412_1570_0, i_13_412_1770_0, i_13_412_1780_0, i_13_412_1798_0,
    i_13_412_1854_0, i_13_412_1858_0, i_13_412_1860_0, i_13_412_1956_0,
    i_13_412_1957_0, i_13_412_2056_0, i_13_412_2110_0, i_13_412_2265_0,
    i_13_412_2281_0, i_13_412_2366_0, i_13_412_2452_0, i_13_412_2454_0,
    i_13_412_2460_0, i_13_412_2473_0, i_13_412_2505_0, i_13_412_2539_0,
    i_13_412_2541_0, i_13_412_2613_0, i_13_412_2622_0, i_13_412_2647_0,
    i_13_412_3031_0, i_13_412_3100_0, i_13_412_3120_0, i_13_412_3170_0,
    i_13_412_3172_0, i_13_412_3273_0, i_13_412_3381_0, i_13_412_3427_0,
    i_13_412_3429_0, i_13_412_3460_0, i_13_412_3468_0, i_13_412_3483_0,
    i_13_412_3503_0, i_13_412_3505_0, i_13_412_3541_0, i_13_412_3559_0,
    i_13_412_3570_0, i_13_412_3651_0, i_13_412_3729_0, i_13_412_3783_0,
    i_13_412_3822_0, i_13_412_3829_0, i_13_412_3856_0, i_13_412_3896_0,
    i_13_412_3910_0, i_13_412_3911_0, i_13_412_4252_0, i_13_412_4254_0,
    i_13_412_4256_0, i_13_412_4261_0, i_13_412_4377_0, i_13_412_4396_0,
    i_13_412_4415_0, i_13_412_4579_0, i_13_412_4597_0, i_13_412_4606_0;
  output o_13_412_0_0;
  assign o_13_412_0_0 = ~((~i_13_412_1255_0 & (~i_13_412_4254_0 | (~i_13_412_3427_0 & ~i_13_412_3822_0))) | (~i_13_412_4254_0 & ((~i_13_412_2541_0 & ~i_13_412_3427_0) | (~i_13_412_1075_0 & i_13_412_3505_0))) | (~i_13_412_1023_0 & ~i_13_412_1956_0 & ~i_13_412_3822_0) | (i_13_412_1224_0 & i_13_412_1498_0 & ~i_13_412_4377_0));
endmodule



// Benchmark "kernel_13_413" written by ABC on Sun Jul 19 10:51:07 2020

module kernel_13_413 ( 
    i_13_413_78_0, i_13_413_79_0, i_13_413_103_0, i_13_413_157_0,
    i_13_413_158_0, i_13_413_185_0, i_13_413_219_0, i_13_413_374_0,
    i_13_413_379_0, i_13_413_515_0, i_13_413_533_0, i_13_413_536_0,
    i_13_413_550_0, i_13_413_551_0, i_13_413_644_0, i_13_413_648_0,
    i_13_413_652_0, i_13_413_653_0, i_13_413_676_0, i_13_413_685_0,
    i_13_413_689_0, i_13_413_823_0, i_13_413_833_0, i_13_413_839_0,
    i_13_413_842_0, i_13_413_1074_0, i_13_413_1104_0, i_13_413_1122_0,
    i_13_413_1145_0, i_13_413_1327_0, i_13_413_1514_0, i_13_413_1515_0,
    i_13_413_1516_0, i_13_413_1517_0, i_13_413_1632_0, i_13_413_1657_0,
    i_13_413_1675_0, i_13_413_1677_0, i_13_413_1678_0, i_13_413_1692_0,
    i_13_413_1739_0, i_13_413_1747_0, i_13_413_1752_0, i_13_413_1776_0,
    i_13_413_1792_0, i_13_413_1909_0, i_13_413_1912_0, i_13_413_1999_0,
    i_13_413_2002_0, i_13_413_2017_0, i_13_413_2025_0, i_13_413_2047_0,
    i_13_413_2101_0, i_13_413_2467_0, i_13_413_2468_0, i_13_413_2507_0,
    i_13_413_2512_0, i_13_413_2542_0, i_13_413_2547_0, i_13_413_2557_0,
    i_13_413_2570_0, i_13_413_2622_0, i_13_413_2722_0, i_13_413_2737_0,
    i_13_413_2740_0, i_13_413_2766_0, i_13_413_2850_0, i_13_413_2854_0,
    i_13_413_2898_0, i_13_413_2908_0, i_13_413_2917_0, i_13_413_2956_0,
    i_13_413_3052_0, i_13_413_3088_0, i_13_413_3235_0, i_13_413_3367_0,
    i_13_413_3377_0, i_13_413_3476_0, i_13_413_3486_0, i_13_413_3487_0,
    i_13_413_3523_0, i_13_413_3604_0, i_13_413_3727_0, i_13_413_3857_0,
    i_13_413_3862_0, i_13_413_3863_0, i_13_413_3925_0, i_13_413_3988_0,
    i_13_413_4123_0, i_13_413_4124_0, i_13_413_4160_0, i_13_413_4187_0,
    i_13_413_4188_0, i_13_413_4260_0, i_13_413_4512_0, i_13_413_4581_0,
    i_13_413_4591_0, i_13_413_4596_0, i_13_413_4600_0, i_13_413_4601_0,
    o_13_413_0_0  );
  input  i_13_413_78_0, i_13_413_79_0, i_13_413_103_0, i_13_413_157_0,
    i_13_413_158_0, i_13_413_185_0, i_13_413_219_0, i_13_413_374_0,
    i_13_413_379_0, i_13_413_515_0, i_13_413_533_0, i_13_413_536_0,
    i_13_413_550_0, i_13_413_551_0, i_13_413_644_0, i_13_413_648_0,
    i_13_413_652_0, i_13_413_653_0, i_13_413_676_0, i_13_413_685_0,
    i_13_413_689_0, i_13_413_823_0, i_13_413_833_0, i_13_413_839_0,
    i_13_413_842_0, i_13_413_1074_0, i_13_413_1104_0, i_13_413_1122_0,
    i_13_413_1145_0, i_13_413_1327_0, i_13_413_1514_0, i_13_413_1515_0,
    i_13_413_1516_0, i_13_413_1517_0, i_13_413_1632_0, i_13_413_1657_0,
    i_13_413_1675_0, i_13_413_1677_0, i_13_413_1678_0, i_13_413_1692_0,
    i_13_413_1739_0, i_13_413_1747_0, i_13_413_1752_0, i_13_413_1776_0,
    i_13_413_1792_0, i_13_413_1909_0, i_13_413_1912_0, i_13_413_1999_0,
    i_13_413_2002_0, i_13_413_2017_0, i_13_413_2025_0, i_13_413_2047_0,
    i_13_413_2101_0, i_13_413_2467_0, i_13_413_2468_0, i_13_413_2507_0,
    i_13_413_2512_0, i_13_413_2542_0, i_13_413_2547_0, i_13_413_2557_0,
    i_13_413_2570_0, i_13_413_2622_0, i_13_413_2722_0, i_13_413_2737_0,
    i_13_413_2740_0, i_13_413_2766_0, i_13_413_2850_0, i_13_413_2854_0,
    i_13_413_2898_0, i_13_413_2908_0, i_13_413_2917_0, i_13_413_2956_0,
    i_13_413_3052_0, i_13_413_3088_0, i_13_413_3235_0, i_13_413_3367_0,
    i_13_413_3377_0, i_13_413_3476_0, i_13_413_3486_0, i_13_413_3487_0,
    i_13_413_3523_0, i_13_413_3604_0, i_13_413_3727_0, i_13_413_3857_0,
    i_13_413_3862_0, i_13_413_3863_0, i_13_413_3925_0, i_13_413_3988_0,
    i_13_413_4123_0, i_13_413_4124_0, i_13_413_4160_0, i_13_413_4187_0,
    i_13_413_4188_0, i_13_413_4260_0, i_13_413_4512_0, i_13_413_4581_0,
    i_13_413_4591_0, i_13_413_4596_0, i_13_413_4600_0, i_13_413_4601_0;
  output o_13_413_0_0;
  assign o_13_413_0_0 = ~((~i_13_413_3862_0 & (i_13_413_1999_0 | i_13_413_2917_0)) | (i_13_413_379_0 & ~i_13_413_536_0 & i_13_413_3857_0) | (~i_13_413_648_0 & ~i_13_413_1657_0 & ~i_13_413_1747_0 & ~i_13_413_3863_0) | (~i_13_413_1074_0 & ~i_13_413_1327_0 & ~i_13_413_4187_0));
endmodule



// Benchmark "kernel_13_414" written by ABC on Sun Jul 19 10:51:08 2020

module kernel_13_414 ( 
    i_13_414_1_0, i_13_414_45_0, i_13_414_46_0, i_13_414_67_0,
    i_13_414_171_0, i_13_414_172_0, i_13_414_234_0, i_13_414_351_0,
    i_13_414_352_0, i_13_414_408_0, i_13_414_450_0, i_13_414_472_0,
    i_13_414_505_0, i_13_414_508_0, i_13_414_511_0, i_13_414_567_0,
    i_13_414_648_0, i_13_414_657_0, i_13_414_661_0, i_13_414_673_0,
    i_13_414_735_0, i_13_414_850_0, i_13_414_936_0, i_13_414_937_0,
    i_13_414_1071_0, i_13_414_1128_0, i_13_414_1129_0, i_13_414_1211_0,
    i_13_414_1243_0, i_13_414_1266_0, i_13_414_1272_0, i_13_414_1314_0,
    i_13_414_1326_0, i_13_414_1410_0, i_13_414_1422_0, i_13_414_1434_0,
    i_13_414_1480_0, i_13_414_1642_0, i_13_414_1663_0, i_13_414_1692_0,
    i_13_414_1729_0, i_13_414_1764_0, i_13_414_1786_0, i_13_414_1795_0,
    i_13_414_1915_0, i_13_414_1939_0, i_13_414_1944_0, i_13_414_1999_0,
    i_13_414_2019_0, i_13_414_2020_0, i_13_414_2026_0, i_13_414_2097_0,
    i_13_414_2176_0, i_13_414_2196_0, i_13_414_2299_0, i_13_414_2340_0,
    i_13_414_2448_0, i_13_414_2469_0, i_13_414_2470_0, i_13_414_2592_0,
    i_13_414_2637_0, i_13_414_2701_0, i_13_414_2704_0, i_13_414_3027_0,
    i_13_414_3028_0, i_13_414_3111_0, i_13_414_3112_0, i_13_414_3126_0,
    i_13_414_3127_0, i_13_414_3132_0, i_13_414_3261_0, i_13_414_3367_0,
    i_13_414_3418_0, i_13_414_3474_0, i_13_414_3478_0, i_13_414_3480_0,
    i_13_414_3481_0, i_13_414_3483_0, i_13_414_3484_0, i_13_414_3531_0,
    i_13_414_3546_0, i_13_414_3573_0, i_13_414_3574_0, i_13_414_3577_0,
    i_13_414_3726_0, i_13_414_3780_0, i_13_414_3781_0, i_13_414_3819_0,
    i_13_414_3897_0, i_13_414_3898_0, i_13_414_4015_0, i_13_414_4161_0,
    i_13_414_4230_0, i_13_414_4293_0, i_13_414_4321_0, i_13_414_4375_0,
    i_13_414_4521_0, i_13_414_4561_0, i_13_414_4563_0, i_13_414_4603_0,
    o_13_414_0_0  );
  input  i_13_414_1_0, i_13_414_45_0, i_13_414_46_0, i_13_414_67_0,
    i_13_414_171_0, i_13_414_172_0, i_13_414_234_0, i_13_414_351_0,
    i_13_414_352_0, i_13_414_408_0, i_13_414_450_0, i_13_414_472_0,
    i_13_414_505_0, i_13_414_508_0, i_13_414_511_0, i_13_414_567_0,
    i_13_414_648_0, i_13_414_657_0, i_13_414_661_0, i_13_414_673_0,
    i_13_414_735_0, i_13_414_850_0, i_13_414_936_0, i_13_414_937_0,
    i_13_414_1071_0, i_13_414_1128_0, i_13_414_1129_0, i_13_414_1211_0,
    i_13_414_1243_0, i_13_414_1266_0, i_13_414_1272_0, i_13_414_1314_0,
    i_13_414_1326_0, i_13_414_1410_0, i_13_414_1422_0, i_13_414_1434_0,
    i_13_414_1480_0, i_13_414_1642_0, i_13_414_1663_0, i_13_414_1692_0,
    i_13_414_1729_0, i_13_414_1764_0, i_13_414_1786_0, i_13_414_1795_0,
    i_13_414_1915_0, i_13_414_1939_0, i_13_414_1944_0, i_13_414_1999_0,
    i_13_414_2019_0, i_13_414_2020_0, i_13_414_2026_0, i_13_414_2097_0,
    i_13_414_2176_0, i_13_414_2196_0, i_13_414_2299_0, i_13_414_2340_0,
    i_13_414_2448_0, i_13_414_2469_0, i_13_414_2470_0, i_13_414_2592_0,
    i_13_414_2637_0, i_13_414_2701_0, i_13_414_2704_0, i_13_414_3027_0,
    i_13_414_3028_0, i_13_414_3111_0, i_13_414_3112_0, i_13_414_3126_0,
    i_13_414_3127_0, i_13_414_3132_0, i_13_414_3261_0, i_13_414_3367_0,
    i_13_414_3418_0, i_13_414_3474_0, i_13_414_3478_0, i_13_414_3480_0,
    i_13_414_3481_0, i_13_414_3483_0, i_13_414_3484_0, i_13_414_3531_0,
    i_13_414_3546_0, i_13_414_3573_0, i_13_414_3574_0, i_13_414_3577_0,
    i_13_414_3726_0, i_13_414_3780_0, i_13_414_3781_0, i_13_414_3819_0,
    i_13_414_3897_0, i_13_414_3898_0, i_13_414_4015_0, i_13_414_4161_0,
    i_13_414_4230_0, i_13_414_4293_0, i_13_414_4321_0, i_13_414_4375_0,
    i_13_414_4521_0, i_13_414_4561_0, i_13_414_4563_0, i_13_414_4603_0;
  output o_13_414_0_0;
  assign o_13_414_0_0 = ~((~i_13_414_4321_0 & (~i_13_414_1272_0 | ~i_13_414_1480_0 | ~i_13_414_3819_0)) | (~i_13_414_472_0 & ~i_13_414_3484_0 & ~i_13_414_3531_0) | (~i_13_414_1071_0 & ~i_13_414_1410_0 & ~i_13_414_1944_0 & ~i_13_414_4375_0));
endmodule



// Benchmark "kernel_13_415" written by ABC on Sun Jul 19 10:51:08 2020

module kernel_13_415 ( 
    i_13_415_162_0, i_13_415_174_0, i_13_415_201_0, i_13_415_363_0,
    i_13_415_412_0, i_13_415_468_0, i_13_415_604_0, i_13_415_657_0,
    i_13_415_658_0, i_13_415_660_0, i_13_415_661_0, i_13_415_667_0,
    i_13_415_694_0, i_13_415_822_0, i_13_415_828_0, i_13_415_829_0,
    i_13_415_831_0, i_13_415_853_0, i_13_415_946_0, i_13_415_954_0,
    i_13_415_955_0, i_13_415_984_0, i_13_415_1071_0, i_13_415_1075_0,
    i_13_415_1098_0, i_13_415_1224_0, i_13_415_1225_0, i_13_415_1269_0,
    i_13_415_1270_0, i_13_415_1305_0, i_13_415_1423_0, i_13_415_1435_0,
    i_13_415_1497_0, i_13_415_1503_0, i_13_415_1522_0, i_13_415_1534_0,
    i_13_415_1548_0, i_13_415_1620_0, i_13_415_1657_0, i_13_415_1722_0,
    i_13_415_1729_0, i_13_415_1764_0, i_13_415_1767_0, i_13_415_1791_0,
    i_13_415_1837_0, i_13_415_2019_0, i_13_415_2020_0, i_13_415_2142_0,
    i_13_415_2172_0, i_13_415_2296_0, i_13_415_2340_0, i_13_415_2365_0,
    i_13_415_2394_0, i_13_415_2430_0, i_13_415_2431_0, i_13_415_2448_0,
    i_13_415_2550_0, i_13_415_2647_0, i_13_415_2691_0, i_13_415_2721_0,
    i_13_415_2880_0, i_13_415_2881_0, i_13_415_2907_0, i_13_415_3000_0,
    i_13_415_3001_0, i_13_415_3060_0, i_13_415_3231_0, i_13_415_3324_0,
    i_13_415_3370_0, i_13_415_3456_0, i_13_415_3478_0, i_13_415_3483_0,
    i_13_415_3484_0, i_13_415_3486_0, i_13_415_3546_0, i_13_415_3547_0,
    i_13_415_3613_0, i_13_415_3619_0, i_13_415_3636_0, i_13_415_3637_0,
    i_13_415_3753_0, i_13_415_3843_0, i_13_415_3853_0, i_13_415_3910_0,
    i_13_415_3982_0, i_13_415_4063_0, i_13_415_4123_0, i_13_415_4161_0,
    i_13_415_4162_0, i_13_415_4251_0, i_13_415_4315_0, i_13_415_4329_0,
    i_13_415_4339_0, i_13_415_4378_0, i_13_415_4429_0, i_13_415_4449_0,
    i_13_415_4458_0, i_13_415_4509_0, i_13_415_4510_0, i_13_415_4600_0,
    o_13_415_0_0  );
  input  i_13_415_162_0, i_13_415_174_0, i_13_415_201_0, i_13_415_363_0,
    i_13_415_412_0, i_13_415_468_0, i_13_415_604_0, i_13_415_657_0,
    i_13_415_658_0, i_13_415_660_0, i_13_415_661_0, i_13_415_667_0,
    i_13_415_694_0, i_13_415_822_0, i_13_415_828_0, i_13_415_829_0,
    i_13_415_831_0, i_13_415_853_0, i_13_415_946_0, i_13_415_954_0,
    i_13_415_955_0, i_13_415_984_0, i_13_415_1071_0, i_13_415_1075_0,
    i_13_415_1098_0, i_13_415_1224_0, i_13_415_1225_0, i_13_415_1269_0,
    i_13_415_1270_0, i_13_415_1305_0, i_13_415_1423_0, i_13_415_1435_0,
    i_13_415_1497_0, i_13_415_1503_0, i_13_415_1522_0, i_13_415_1534_0,
    i_13_415_1548_0, i_13_415_1620_0, i_13_415_1657_0, i_13_415_1722_0,
    i_13_415_1729_0, i_13_415_1764_0, i_13_415_1767_0, i_13_415_1791_0,
    i_13_415_1837_0, i_13_415_2019_0, i_13_415_2020_0, i_13_415_2142_0,
    i_13_415_2172_0, i_13_415_2296_0, i_13_415_2340_0, i_13_415_2365_0,
    i_13_415_2394_0, i_13_415_2430_0, i_13_415_2431_0, i_13_415_2448_0,
    i_13_415_2550_0, i_13_415_2647_0, i_13_415_2691_0, i_13_415_2721_0,
    i_13_415_2880_0, i_13_415_2881_0, i_13_415_2907_0, i_13_415_3000_0,
    i_13_415_3001_0, i_13_415_3060_0, i_13_415_3231_0, i_13_415_3324_0,
    i_13_415_3370_0, i_13_415_3456_0, i_13_415_3478_0, i_13_415_3483_0,
    i_13_415_3484_0, i_13_415_3486_0, i_13_415_3546_0, i_13_415_3547_0,
    i_13_415_3613_0, i_13_415_3619_0, i_13_415_3636_0, i_13_415_3637_0,
    i_13_415_3753_0, i_13_415_3843_0, i_13_415_3853_0, i_13_415_3910_0,
    i_13_415_3982_0, i_13_415_4063_0, i_13_415_4123_0, i_13_415_4161_0,
    i_13_415_4162_0, i_13_415_4251_0, i_13_415_4315_0, i_13_415_4329_0,
    i_13_415_4339_0, i_13_415_4378_0, i_13_415_4429_0, i_13_415_4449_0,
    i_13_415_4458_0, i_13_415_4509_0, i_13_415_4510_0, i_13_415_4600_0;
  output o_13_415_0_0;
  assign o_13_415_0_0 = ~(~i_13_415_828_0);
endmodule



// Benchmark "kernel_13_416" written by ABC on Sun Jul 19 10:51:09 2020

module kernel_13_416 ( 
    i_13_416_33_0, i_13_416_40_0, i_13_416_93_0, i_13_416_96_0,
    i_13_416_105_0, i_13_416_106_0, i_13_416_159_0, i_13_416_185_0,
    i_13_416_268_0, i_13_416_286_0, i_13_416_318_0, i_13_416_321_0,
    i_13_416_338_0, i_13_416_372_0, i_13_416_569_0, i_13_416_699_0,
    i_13_416_700_0, i_13_416_744_0, i_13_416_816_0, i_13_416_817_0,
    i_13_416_843_0, i_13_416_931_0, i_13_416_984_0, i_13_416_985_0,
    i_13_416_1069_0, i_13_416_1122_0, i_13_416_1210_0, i_13_416_1308_0,
    i_13_416_1407_0, i_13_416_1429_0, i_13_416_1446_0, i_13_416_1481_0,
    i_13_416_1499_0, i_13_416_1518_0, i_13_416_1645_0, i_13_416_1652_0,
    i_13_416_1730_0, i_13_416_1733_0, i_13_416_1752_0, i_13_416_1753_0,
    i_13_416_1787_0, i_13_416_1813_0, i_13_416_1851_0, i_13_416_1933_0,
    i_13_416_1992_0, i_13_416_1995_0, i_13_416_2017_0, i_13_416_2058_0,
    i_13_416_2122_0, i_13_416_2139_0, i_13_416_2172_0, i_13_416_2266_0,
    i_13_416_2409_0, i_13_416_2410_0, i_13_416_2459_0, i_13_416_2472_0,
    i_13_416_2545_0, i_13_416_2617_0, i_13_416_2679_0, i_13_416_2680_0,
    i_13_416_2741_0, i_13_416_2787_0, i_13_416_2940_0, i_13_416_2981_0,
    i_13_416_2985_0, i_13_416_3022_0, i_13_416_3210_0, i_13_416_3211_0,
    i_13_416_3345_0, i_13_416_3371_0, i_13_416_3381_0, i_13_416_3390_0,
    i_13_416_3399_0, i_13_416_3400_0, i_13_416_3422_0, i_13_416_3449_0,
    i_13_416_3451_0, i_13_416_3488_0, i_13_416_3489_0, i_13_416_3521_0,
    i_13_416_3535_0, i_13_416_3702_0, i_13_416_3720_0, i_13_416_3764_0,
    i_13_416_3791_0, i_13_416_3911_0, i_13_416_3983_0, i_13_416_4047_0,
    i_13_416_4066_0, i_13_416_4083_0, i_13_416_4084_0, i_13_416_4191_0,
    i_13_416_4295_0, i_13_416_4350_0, i_13_416_4353_0, i_13_416_4395_0,
    i_13_416_4396_0, i_13_416_4416_0, i_13_416_4451_0, i_13_416_4538_0,
    o_13_416_0_0  );
  input  i_13_416_33_0, i_13_416_40_0, i_13_416_93_0, i_13_416_96_0,
    i_13_416_105_0, i_13_416_106_0, i_13_416_159_0, i_13_416_185_0,
    i_13_416_268_0, i_13_416_286_0, i_13_416_318_0, i_13_416_321_0,
    i_13_416_338_0, i_13_416_372_0, i_13_416_569_0, i_13_416_699_0,
    i_13_416_700_0, i_13_416_744_0, i_13_416_816_0, i_13_416_817_0,
    i_13_416_843_0, i_13_416_931_0, i_13_416_984_0, i_13_416_985_0,
    i_13_416_1069_0, i_13_416_1122_0, i_13_416_1210_0, i_13_416_1308_0,
    i_13_416_1407_0, i_13_416_1429_0, i_13_416_1446_0, i_13_416_1481_0,
    i_13_416_1499_0, i_13_416_1518_0, i_13_416_1645_0, i_13_416_1652_0,
    i_13_416_1730_0, i_13_416_1733_0, i_13_416_1752_0, i_13_416_1753_0,
    i_13_416_1787_0, i_13_416_1813_0, i_13_416_1851_0, i_13_416_1933_0,
    i_13_416_1992_0, i_13_416_1995_0, i_13_416_2017_0, i_13_416_2058_0,
    i_13_416_2122_0, i_13_416_2139_0, i_13_416_2172_0, i_13_416_2266_0,
    i_13_416_2409_0, i_13_416_2410_0, i_13_416_2459_0, i_13_416_2472_0,
    i_13_416_2545_0, i_13_416_2617_0, i_13_416_2679_0, i_13_416_2680_0,
    i_13_416_2741_0, i_13_416_2787_0, i_13_416_2940_0, i_13_416_2981_0,
    i_13_416_2985_0, i_13_416_3022_0, i_13_416_3210_0, i_13_416_3211_0,
    i_13_416_3345_0, i_13_416_3371_0, i_13_416_3381_0, i_13_416_3390_0,
    i_13_416_3399_0, i_13_416_3400_0, i_13_416_3422_0, i_13_416_3449_0,
    i_13_416_3451_0, i_13_416_3488_0, i_13_416_3489_0, i_13_416_3521_0,
    i_13_416_3535_0, i_13_416_3702_0, i_13_416_3720_0, i_13_416_3764_0,
    i_13_416_3791_0, i_13_416_3911_0, i_13_416_3983_0, i_13_416_4047_0,
    i_13_416_4066_0, i_13_416_4083_0, i_13_416_4084_0, i_13_416_4191_0,
    i_13_416_4295_0, i_13_416_4350_0, i_13_416_4353_0, i_13_416_4395_0,
    i_13_416_4396_0, i_13_416_4416_0, i_13_416_4451_0, i_13_416_4538_0;
  output o_13_416_0_0;
  assign o_13_416_0_0 = ~(~i_13_416_3400_0 | (~i_13_416_1122_0 & ~i_13_416_4083_0) | (i_13_416_843_0 & ~i_13_416_2172_0 & i_13_416_4083_0));
endmodule



// Benchmark "kernel_13_417" written by ABC on Sun Jul 19 10:51:10 2020

module kernel_13_417 ( 
    i_13_417_76_0, i_13_417_205_0, i_13_417_258_0, i_13_417_286_0,
    i_13_417_309_0, i_13_417_340_0, i_13_417_411_0, i_13_417_519_0,
    i_13_417_561_0, i_13_417_586_0, i_13_417_607_0, i_13_417_618_0,
    i_13_417_619_0, i_13_417_627_0, i_13_417_640_0, i_13_417_661_0,
    i_13_417_663_0, i_13_417_672_0, i_13_417_757_0, i_13_417_771_0,
    i_13_417_799_0, i_13_417_856_0, i_13_417_1021_0, i_13_417_1111_0,
    i_13_417_1147_0, i_13_417_1278_0, i_13_417_1279_0, i_13_417_1303_0,
    i_13_417_1329_0, i_13_417_1330_0, i_13_417_1429_0, i_13_417_1572_0,
    i_13_417_1596_0, i_13_417_1633_0, i_13_417_1659_0, i_13_417_1734_0,
    i_13_417_1735_0, i_13_417_1744_0, i_13_417_1767_0, i_13_417_1834_0,
    i_13_417_1843_0, i_13_417_1891_0, i_13_417_1932_0, i_13_417_1959_0,
    i_13_417_2019_0, i_13_417_2022_0, i_13_417_2023_0, i_13_417_2134_0,
    i_13_417_2211_0, i_13_417_2248_0, i_13_417_2260_0, i_13_417_2452_0,
    i_13_417_2454_0, i_13_417_2455_0, i_13_417_2469_0, i_13_417_2610_0,
    i_13_417_2707_0, i_13_417_2715_0, i_13_417_2742_0, i_13_417_2743_0,
    i_13_417_2746_0, i_13_417_2787_0, i_13_417_2886_0, i_13_417_2922_0,
    i_13_417_2958_0, i_13_417_3031_0, i_13_417_3075_0, i_13_417_3076_0,
    i_13_417_3102_0, i_13_417_3315_0, i_13_417_3448_0, i_13_417_3486_0,
    i_13_417_3489_0, i_13_417_3490_0, i_13_417_3519_0, i_13_417_3553_0,
    i_13_417_3570_0, i_13_417_3603_0, i_13_417_3822_0, i_13_417_3865_0,
    i_13_417_3901_0, i_13_417_4021_0, i_13_417_4119_0, i_13_417_4161_0,
    i_13_417_4164_0, i_13_417_4165_0, i_13_417_4179_0, i_13_417_4189_0,
    i_13_417_4191_0, i_13_417_4255_0, i_13_417_4293_0, i_13_417_4332_0,
    i_13_417_4333_0, i_13_417_4362_0, i_13_417_4374_0, i_13_417_4516_0,
    i_13_417_4600_0, i_13_417_4602_0, i_13_417_4605_0, i_13_417_4606_0,
    o_13_417_0_0  );
  input  i_13_417_76_0, i_13_417_205_0, i_13_417_258_0, i_13_417_286_0,
    i_13_417_309_0, i_13_417_340_0, i_13_417_411_0, i_13_417_519_0,
    i_13_417_561_0, i_13_417_586_0, i_13_417_607_0, i_13_417_618_0,
    i_13_417_619_0, i_13_417_627_0, i_13_417_640_0, i_13_417_661_0,
    i_13_417_663_0, i_13_417_672_0, i_13_417_757_0, i_13_417_771_0,
    i_13_417_799_0, i_13_417_856_0, i_13_417_1021_0, i_13_417_1111_0,
    i_13_417_1147_0, i_13_417_1278_0, i_13_417_1279_0, i_13_417_1303_0,
    i_13_417_1329_0, i_13_417_1330_0, i_13_417_1429_0, i_13_417_1572_0,
    i_13_417_1596_0, i_13_417_1633_0, i_13_417_1659_0, i_13_417_1734_0,
    i_13_417_1735_0, i_13_417_1744_0, i_13_417_1767_0, i_13_417_1834_0,
    i_13_417_1843_0, i_13_417_1891_0, i_13_417_1932_0, i_13_417_1959_0,
    i_13_417_2019_0, i_13_417_2022_0, i_13_417_2023_0, i_13_417_2134_0,
    i_13_417_2211_0, i_13_417_2248_0, i_13_417_2260_0, i_13_417_2452_0,
    i_13_417_2454_0, i_13_417_2455_0, i_13_417_2469_0, i_13_417_2610_0,
    i_13_417_2707_0, i_13_417_2715_0, i_13_417_2742_0, i_13_417_2743_0,
    i_13_417_2746_0, i_13_417_2787_0, i_13_417_2886_0, i_13_417_2922_0,
    i_13_417_2958_0, i_13_417_3031_0, i_13_417_3075_0, i_13_417_3076_0,
    i_13_417_3102_0, i_13_417_3315_0, i_13_417_3448_0, i_13_417_3486_0,
    i_13_417_3489_0, i_13_417_3490_0, i_13_417_3519_0, i_13_417_3553_0,
    i_13_417_3570_0, i_13_417_3603_0, i_13_417_3822_0, i_13_417_3865_0,
    i_13_417_3901_0, i_13_417_4021_0, i_13_417_4119_0, i_13_417_4161_0,
    i_13_417_4164_0, i_13_417_4165_0, i_13_417_4179_0, i_13_417_4189_0,
    i_13_417_4191_0, i_13_417_4255_0, i_13_417_4293_0, i_13_417_4332_0,
    i_13_417_4333_0, i_13_417_4362_0, i_13_417_4374_0, i_13_417_4516_0,
    i_13_417_4600_0, i_13_417_4602_0, i_13_417_4605_0, i_13_417_4606_0;
  output o_13_417_0_0;
  assign o_13_417_0_0 = ~((~i_13_417_619_0 & ~i_13_417_4161_0) | (~i_13_417_2022_0 & ~i_13_417_2454_0));
endmodule



// Benchmark "kernel_13_418" written by ABC on Sun Jul 19 10:51:11 2020

module kernel_13_418 ( 
    i_13_418_64_0, i_13_418_76_0, i_13_418_77_0, i_13_418_103_0,
    i_13_418_121_0, i_13_418_173_0, i_13_418_190_0, i_13_418_284_0,
    i_13_418_374_0, i_13_418_382_0, i_13_418_385_0, i_13_418_415_0,
    i_13_418_463_0, i_13_418_493_0, i_13_418_524_0, i_13_418_527_0,
    i_13_418_571_0, i_13_418_581_0, i_13_418_589_0, i_13_418_598_0,
    i_13_418_599_0, i_13_418_686_0, i_13_418_694_0, i_13_418_695_0,
    i_13_418_698_0, i_13_418_824_0, i_13_418_1207_0, i_13_418_1208_0,
    i_13_418_1211_0, i_13_418_1307_0, i_13_418_1309_0, i_13_418_1310_0,
    i_13_418_1343_0, i_13_418_1385_0, i_13_418_1403_0, i_13_418_1508_0,
    i_13_418_1516_0, i_13_418_1550_0, i_13_418_1594_0, i_13_418_1595_0,
    i_13_418_1597_0, i_13_418_1610_0, i_13_418_1685_0, i_13_418_1883_0,
    i_13_418_1886_0, i_13_418_1928_0, i_13_418_1931_0, i_13_418_1939_0,
    i_13_418_1945_0, i_13_418_2000_0, i_13_418_2002_0, i_13_418_2003_0,
    i_13_418_2125_0, i_13_418_2189_0, i_13_418_2201_0, i_13_418_2209_0,
    i_13_418_2239_0, i_13_418_2302_0, i_13_418_2449_0, i_13_418_2549_0,
    i_13_418_2657_0, i_13_418_2675_0, i_13_418_2719_0, i_13_418_2720_0,
    i_13_418_2824_0, i_13_418_2857_0, i_13_418_2858_0, i_13_418_2969_0,
    i_13_418_3010_0, i_13_418_3031_0, i_13_418_3062_0, i_13_418_3208_0,
    i_13_418_3217_0, i_13_418_3374_0, i_13_418_3400_0, i_13_418_3562_0,
    i_13_418_3563_0, i_13_418_3650_0, i_13_418_3667_0, i_13_418_3670_0,
    i_13_418_3727_0, i_13_418_3728_0, i_13_418_3731_0, i_13_418_3893_0,
    i_13_418_3916_0, i_13_418_3982_0, i_13_418_4015_0, i_13_418_4016_0,
    i_13_418_4019_0, i_13_418_4259_0, i_13_418_4261_0, i_13_418_4262_0,
    i_13_418_4303_0, i_13_418_4396_0, i_13_418_4397_0, i_13_418_4417_0,
    i_13_418_4447_0, i_13_418_4454_0, i_13_418_4540_0, i_13_418_4556_0,
    o_13_418_0_0  );
  input  i_13_418_64_0, i_13_418_76_0, i_13_418_77_0, i_13_418_103_0,
    i_13_418_121_0, i_13_418_173_0, i_13_418_190_0, i_13_418_284_0,
    i_13_418_374_0, i_13_418_382_0, i_13_418_385_0, i_13_418_415_0,
    i_13_418_463_0, i_13_418_493_0, i_13_418_524_0, i_13_418_527_0,
    i_13_418_571_0, i_13_418_581_0, i_13_418_589_0, i_13_418_598_0,
    i_13_418_599_0, i_13_418_686_0, i_13_418_694_0, i_13_418_695_0,
    i_13_418_698_0, i_13_418_824_0, i_13_418_1207_0, i_13_418_1208_0,
    i_13_418_1211_0, i_13_418_1307_0, i_13_418_1309_0, i_13_418_1310_0,
    i_13_418_1343_0, i_13_418_1385_0, i_13_418_1403_0, i_13_418_1508_0,
    i_13_418_1516_0, i_13_418_1550_0, i_13_418_1594_0, i_13_418_1595_0,
    i_13_418_1597_0, i_13_418_1610_0, i_13_418_1685_0, i_13_418_1883_0,
    i_13_418_1886_0, i_13_418_1928_0, i_13_418_1931_0, i_13_418_1939_0,
    i_13_418_1945_0, i_13_418_2000_0, i_13_418_2002_0, i_13_418_2003_0,
    i_13_418_2125_0, i_13_418_2189_0, i_13_418_2201_0, i_13_418_2209_0,
    i_13_418_2239_0, i_13_418_2302_0, i_13_418_2449_0, i_13_418_2549_0,
    i_13_418_2657_0, i_13_418_2675_0, i_13_418_2719_0, i_13_418_2720_0,
    i_13_418_2824_0, i_13_418_2857_0, i_13_418_2858_0, i_13_418_2969_0,
    i_13_418_3010_0, i_13_418_3031_0, i_13_418_3062_0, i_13_418_3208_0,
    i_13_418_3217_0, i_13_418_3374_0, i_13_418_3400_0, i_13_418_3562_0,
    i_13_418_3563_0, i_13_418_3650_0, i_13_418_3667_0, i_13_418_3670_0,
    i_13_418_3727_0, i_13_418_3728_0, i_13_418_3731_0, i_13_418_3893_0,
    i_13_418_3916_0, i_13_418_3982_0, i_13_418_4015_0, i_13_418_4016_0,
    i_13_418_4019_0, i_13_418_4259_0, i_13_418_4261_0, i_13_418_4262_0,
    i_13_418_4303_0, i_13_418_4396_0, i_13_418_4397_0, i_13_418_4417_0,
    i_13_418_4447_0, i_13_418_4454_0, i_13_418_4540_0, i_13_418_4556_0;
  output o_13_418_0_0;
  assign o_13_418_0_0 = ~((~i_13_418_2000_0 & (~i_13_418_589_0 | ~i_13_418_4556_0)) | (~i_13_418_2858_0 & ~i_13_418_3010_0 & ~i_13_418_3650_0) | (~i_13_418_2003_0 & ~i_13_418_3916_0) | (~i_13_418_3727_0 & ~i_13_418_4262_0 & ~i_13_418_4447_0));
endmodule



// Benchmark "kernel_13_419" written by ABC on Sun Jul 19 10:51:12 2020

module kernel_13_419 ( 
    i_13_419_121_0, i_13_419_171_0, i_13_419_175_0, i_13_419_202_0,
    i_13_419_324_0, i_13_419_325_0, i_13_419_414_0, i_13_419_415_0,
    i_13_419_432_0, i_13_419_558_0, i_13_419_566_0, i_13_419_568_0,
    i_13_419_822_0, i_13_419_823_0, i_13_419_868_0, i_13_419_891_0,
    i_13_419_1020_0, i_13_419_1071_0, i_13_419_1072_0, i_13_419_1092_0,
    i_13_419_1224_0, i_13_419_1225_0, i_13_419_1227_0, i_13_419_1251_0,
    i_13_419_1255_0, i_13_419_1278_0, i_13_419_1314_0, i_13_419_1317_0,
    i_13_419_1380_0, i_13_419_1414_0, i_13_419_1469_0, i_13_419_1511_0,
    i_13_419_1534_0, i_13_419_1540_0, i_13_419_1548_0, i_13_419_1549_0,
    i_13_419_1602_0, i_13_419_1668_0, i_13_419_1767_0, i_13_419_1775_0,
    i_13_419_1809_0, i_13_419_1854_0, i_13_419_1855_0, i_13_419_1881_0,
    i_13_419_1885_0, i_13_419_2171_0, i_13_419_2244_0, i_13_419_2405_0,
    i_13_419_2448_0, i_13_419_2457_0, i_13_419_2458_0, i_13_419_2539_0,
    i_13_419_2560_0, i_13_419_2566_0, i_13_419_2610_0, i_13_419_2629_0,
    i_13_419_2659_0, i_13_419_2883_0, i_13_419_2919_0, i_13_419_3007_0,
    i_13_419_3091_0, i_13_419_3168_0, i_13_419_3176_0, i_13_419_3236_0,
    i_13_419_3261_0, i_13_419_3307_0, i_13_419_3322_0, i_13_419_3415_0,
    i_13_419_3429_0, i_13_419_3456_0, i_13_419_3457_0, i_13_419_3459_0,
    i_13_419_3531_0, i_13_419_3537_0, i_13_419_3538_0, i_13_419_3540_0,
    i_13_419_3573_0, i_13_419_3726_0, i_13_419_3766_0, i_13_419_3784_0,
    i_13_419_3817_0, i_13_419_3855_0, i_13_419_3907_0, i_13_419_3909_0,
    i_13_419_3983_0, i_13_419_3988_0, i_13_419_4014_0, i_13_419_4015_0,
    i_13_419_4096_0, i_13_419_4248_0, i_13_419_4304_0, i_13_419_4338_0,
    i_13_419_4351_0, i_13_419_4374_0, i_13_419_4375_0, i_13_419_4378_0,
    i_13_419_4440_0, i_13_419_4447_0, i_13_419_4554_0, i_13_419_4557_0,
    o_13_419_0_0  );
  input  i_13_419_121_0, i_13_419_171_0, i_13_419_175_0, i_13_419_202_0,
    i_13_419_324_0, i_13_419_325_0, i_13_419_414_0, i_13_419_415_0,
    i_13_419_432_0, i_13_419_558_0, i_13_419_566_0, i_13_419_568_0,
    i_13_419_822_0, i_13_419_823_0, i_13_419_868_0, i_13_419_891_0,
    i_13_419_1020_0, i_13_419_1071_0, i_13_419_1072_0, i_13_419_1092_0,
    i_13_419_1224_0, i_13_419_1225_0, i_13_419_1227_0, i_13_419_1251_0,
    i_13_419_1255_0, i_13_419_1278_0, i_13_419_1314_0, i_13_419_1317_0,
    i_13_419_1380_0, i_13_419_1414_0, i_13_419_1469_0, i_13_419_1511_0,
    i_13_419_1534_0, i_13_419_1540_0, i_13_419_1548_0, i_13_419_1549_0,
    i_13_419_1602_0, i_13_419_1668_0, i_13_419_1767_0, i_13_419_1775_0,
    i_13_419_1809_0, i_13_419_1854_0, i_13_419_1855_0, i_13_419_1881_0,
    i_13_419_1885_0, i_13_419_2171_0, i_13_419_2244_0, i_13_419_2405_0,
    i_13_419_2448_0, i_13_419_2457_0, i_13_419_2458_0, i_13_419_2539_0,
    i_13_419_2560_0, i_13_419_2566_0, i_13_419_2610_0, i_13_419_2629_0,
    i_13_419_2659_0, i_13_419_2883_0, i_13_419_2919_0, i_13_419_3007_0,
    i_13_419_3091_0, i_13_419_3168_0, i_13_419_3176_0, i_13_419_3236_0,
    i_13_419_3261_0, i_13_419_3307_0, i_13_419_3322_0, i_13_419_3415_0,
    i_13_419_3429_0, i_13_419_3456_0, i_13_419_3457_0, i_13_419_3459_0,
    i_13_419_3531_0, i_13_419_3537_0, i_13_419_3538_0, i_13_419_3540_0,
    i_13_419_3573_0, i_13_419_3726_0, i_13_419_3766_0, i_13_419_3784_0,
    i_13_419_3817_0, i_13_419_3855_0, i_13_419_3907_0, i_13_419_3909_0,
    i_13_419_3983_0, i_13_419_3988_0, i_13_419_4014_0, i_13_419_4015_0,
    i_13_419_4096_0, i_13_419_4248_0, i_13_419_4304_0, i_13_419_4338_0,
    i_13_419_4351_0, i_13_419_4374_0, i_13_419_4375_0, i_13_419_4378_0,
    i_13_419_4440_0, i_13_419_4447_0, i_13_419_4554_0, i_13_419_4557_0;
  output o_13_419_0_0;
  assign o_13_419_0_0 = ~((~i_13_419_3538_0 & (~i_13_419_1225_0 | (~i_13_419_1071_0 & ~i_13_419_2919_0))) | (~i_13_419_2244_0 & ~i_13_419_3540_0));
endmodule



// Benchmark "kernel_13_420" written by ABC on Sun Jul 19 10:51:12 2020

module kernel_13_420 ( 
    i_13_420_0_0, i_13_420_45_0, i_13_420_46_0, i_13_420_63_0,
    i_13_420_64_0, i_13_420_66_0, i_13_420_121_0, i_13_420_183_0,
    i_13_420_234_0, i_13_420_255_0, i_13_420_256_0, i_13_420_310_0,
    i_13_420_414_0, i_13_420_415_0, i_13_420_444_0, i_13_420_468_0,
    i_13_420_469_0, i_13_420_489_0, i_13_420_490_0, i_13_420_586_0,
    i_13_420_603_0, i_13_420_612_0, i_13_420_613_0, i_13_420_666_0,
    i_13_420_685_0, i_13_420_694_0, i_13_420_695_0, i_13_420_760_0,
    i_13_420_839_0, i_13_420_928_0, i_13_420_945_0, i_13_420_1073_0,
    i_13_420_1101_0, i_13_420_1116_0, i_13_420_1129_0, i_13_420_1269_0,
    i_13_420_1270_0, i_13_420_1342_0, i_13_420_1422_0, i_13_420_1494_0,
    i_13_420_1506_0, i_13_420_1549_0, i_13_420_1596_0, i_13_420_1597_0,
    i_13_420_1603_0, i_13_420_1641_0, i_13_420_1669_0, i_13_420_1751_0,
    i_13_420_1777_0, i_13_420_1795_0, i_13_420_1926_0, i_13_420_1927_0,
    i_13_420_1930_0, i_13_420_1944_0, i_13_420_1998_0, i_13_420_1999_0,
    i_13_420_2070_0, i_13_420_2299_0, i_13_420_2377_0, i_13_420_2460_0,
    i_13_420_2505_0, i_13_420_2547_0, i_13_420_2676_0, i_13_420_2721_0,
    i_13_420_2722_0, i_13_420_2749_0, i_13_420_2880_0, i_13_420_2881_0,
    i_13_420_3091_0, i_13_420_3127_0, i_13_420_3261_0, i_13_420_3334_0,
    i_13_420_3366_0, i_13_420_3414_0, i_13_420_3415_0, i_13_420_3546_0,
    i_13_420_3547_0, i_13_420_3550_0, i_13_420_3610_0, i_13_420_3636_0,
    i_13_420_3637_0, i_13_420_3638_0, i_13_420_3699_0, i_13_420_3765_0,
    i_13_420_3766_0, i_13_420_3767_0, i_13_420_3781_0, i_13_420_3784_0,
    i_13_420_3793_0, i_13_420_3897_0, i_13_420_3937_0, i_13_420_3990_0,
    i_13_420_4036_0, i_13_420_4042_0, i_13_420_4080_0, i_13_420_4248_0,
    i_13_420_4257_0, i_13_420_4293_0, i_13_420_4294_0, i_13_420_4347_0,
    o_13_420_0_0  );
  input  i_13_420_0_0, i_13_420_45_0, i_13_420_46_0, i_13_420_63_0,
    i_13_420_64_0, i_13_420_66_0, i_13_420_121_0, i_13_420_183_0,
    i_13_420_234_0, i_13_420_255_0, i_13_420_256_0, i_13_420_310_0,
    i_13_420_414_0, i_13_420_415_0, i_13_420_444_0, i_13_420_468_0,
    i_13_420_469_0, i_13_420_489_0, i_13_420_490_0, i_13_420_586_0,
    i_13_420_603_0, i_13_420_612_0, i_13_420_613_0, i_13_420_666_0,
    i_13_420_685_0, i_13_420_694_0, i_13_420_695_0, i_13_420_760_0,
    i_13_420_839_0, i_13_420_928_0, i_13_420_945_0, i_13_420_1073_0,
    i_13_420_1101_0, i_13_420_1116_0, i_13_420_1129_0, i_13_420_1269_0,
    i_13_420_1270_0, i_13_420_1342_0, i_13_420_1422_0, i_13_420_1494_0,
    i_13_420_1506_0, i_13_420_1549_0, i_13_420_1596_0, i_13_420_1597_0,
    i_13_420_1603_0, i_13_420_1641_0, i_13_420_1669_0, i_13_420_1751_0,
    i_13_420_1777_0, i_13_420_1795_0, i_13_420_1926_0, i_13_420_1927_0,
    i_13_420_1930_0, i_13_420_1944_0, i_13_420_1998_0, i_13_420_1999_0,
    i_13_420_2070_0, i_13_420_2299_0, i_13_420_2377_0, i_13_420_2460_0,
    i_13_420_2505_0, i_13_420_2547_0, i_13_420_2676_0, i_13_420_2721_0,
    i_13_420_2722_0, i_13_420_2749_0, i_13_420_2880_0, i_13_420_2881_0,
    i_13_420_3091_0, i_13_420_3127_0, i_13_420_3261_0, i_13_420_3334_0,
    i_13_420_3366_0, i_13_420_3414_0, i_13_420_3415_0, i_13_420_3546_0,
    i_13_420_3547_0, i_13_420_3550_0, i_13_420_3610_0, i_13_420_3636_0,
    i_13_420_3637_0, i_13_420_3638_0, i_13_420_3699_0, i_13_420_3765_0,
    i_13_420_3766_0, i_13_420_3767_0, i_13_420_3781_0, i_13_420_3784_0,
    i_13_420_3793_0, i_13_420_3897_0, i_13_420_3937_0, i_13_420_3990_0,
    i_13_420_4036_0, i_13_420_4042_0, i_13_420_4080_0, i_13_420_4248_0,
    i_13_420_4257_0, i_13_420_4293_0, i_13_420_4294_0, i_13_420_4347_0;
  output o_13_420_0_0;
  assign o_13_420_0_0 = ~((~i_13_420_310_0 & ((~i_13_420_469_0 & ~i_13_420_2881_0 & i_13_420_4248_0) | (~i_13_420_234_0 & ~i_13_420_1603_0 & ~i_13_420_4248_0))) | (~i_13_420_2880_0 & ((~i_13_420_63_0 & ~i_13_420_468_0) | (~i_13_420_1506_0 & ~i_13_420_3990_0 & ~i_13_420_4042_0))) | (~i_13_420_613_0 & i_13_420_3766_0));
endmodule



// Benchmark "kernel_13_421" written by ABC on Sun Jul 19 10:51:13 2020

module kernel_13_421 ( 
    i_13_421_76_0, i_13_421_184_0, i_13_421_187_0, i_13_421_188_0,
    i_13_421_193_0, i_13_421_322_0, i_13_421_382_0, i_13_421_509_0,
    i_13_421_567_0, i_13_421_571_0, i_13_421_572_0, i_13_421_575_0,
    i_13_421_628_0, i_13_421_647_0, i_13_421_658_0, i_13_421_689_0,
    i_13_421_692_0, i_13_421_818_0, i_13_421_879_0, i_13_421_898_0,
    i_13_421_959_0, i_13_421_995_0, i_13_421_1020_0, i_13_421_1075_0,
    i_13_421_1098_0, i_13_421_1121_0, i_13_421_1123_0, i_13_421_1124_0,
    i_13_421_1143_0, i_13_421_1166_0, i_13_421_1224_0, i_13_421_1228_0,
    i_13_421_1232_0, i_13_421_1277_0, i_13_421_1346_0, i_13_421_1408_0,
    i_13_421_1411_0, i_13_421_1484_0, i_13_421_1516_0, i_13_421_1519_0,
    i_13_421_1645_0, i_13_421_1671_0, i_13_421_1678_0, i_13_421_1728_0,
    i_13_421_1729_0, i_13_421_1751_0, i_13_421_1754_0, i_13_421_1771_0,
    i_13_421_1804_0, i_13_421_1805_0, i_13_421_1807_0, i_13_421_1808_0,
    i_13_421_1858_0, i_13_421_1859_0, i_13_421_1862_0, i_13_421_2123_0,
    i_13_421_2136_0, i_13_421_2195_0, i_13_421_2267_0, i_13_421_2357_0,
    i_13_421_2473_0, i_13_421_2474_0, i_13_421_2624_0, i_13_421_2679_0,
    i_13_421_2681_0, i_13_421_2723_0, i_13_421_2823_0, i_13_421_2825_0,
    i_13_421_2857_0, i_13_421_2942_0, i_13_421_2983_0, i_13_421_2986_0,
    i_13_421_2987_0, i_13_421_3031_0, i_13_421_3032_0, i_13_421_3064_0,
    i_13_421_3074_0, i_13_421_3208_0, i_13_421_3209_0, i_13_421_3235_0,
    i_13_421_3265_0, i_13_421_3293_0, i_13_421_3347_0, i_13_421_3382_0,
    i_13_421_3401_0, i_13_421_3427_0, i_13_421_3506_0, i_13_421_3526_0,
    i_13_421_3681_0, i_13_421_3824_0, i_13_421_3861_0, i_13_421_3911_0,
    i_13_421_3913_0, i_13_421_4338_0, i_13_421_4396_0, i_13_421_4514_0,
    i_13_421_4540_0, i_13_421_4567_0, i_13_421_4598_0, i_13_421_4607_0,
    o_13_421_0_0  );
  input  i_13_421_76_0, i_13_421_184_0, i_13_421_187_0, i_13_421_188_0,
    i_13_421_193_0, i_13_421_322_0, i_13_421_382_0, i_13_421_509_0,
    i_13_421_567_0, i_13_421_571_0, i_13_421_572_0, i_13_421_575_0,
    i_13_421_628_0, i_13_421_647_0, i_13_421_658_0, i_13_421_689_0,
    i_13_421_692_0, i_13_421_818_0, i_13_421_879_0, i_13_421_898_0,
    i_13_421_959_0, i_13_421_995_0, i_13_421_1020_0, i_13_421_1075_0,
    i_13_421_1098_0, i_13_421_1121_0, i_13_421_1123_0, i_13_421_1124_0,
    i_13_421_1143_0, i_13_421_1166_0, i_13_421_1224_0, i_13_421_1228_0,
    i_13_421_1232_0, i_13_421_1277_0, i_13_421_1346_0, i_13_421_1408_0,
    i_13_421_1411_0, i_13_421_1484_0, i_13_421_1516_0, i_13_421_1519_0,
    i_13_421_1645_0, i_13_421_1671_0, i_13_421_1678_0, i_13_421_1728_0,
    i_13_421_1729_0, i_13_421_1751_0, i_13_421_1754_0, i_13_421_1771_0,
    i_13_421_1804_0, i_13_421_1805_0, i_13_421_1807_0, i_13_421_1808_0,
    i_13_421_1858_0, i_13_421_1859_0, i_13_421_1862_0, i_13_421_2123_0,
    i_13_421_2136_0, i_13_421_2195_0, i_13_421_2267_0, i_13_421_2357_0,
    i_13_421_2473_0, i_13_421_2474_0, i_13_421_2624_0, i_13_421_2679_0,
    i_13_421_2681_0, i_13_421_2723_0, i_13_421_2823_0, i_13_421_2825_0,
    i_13_421_2857_0, i_13_421_2942_0, i_13_421_2983_0, i_13_421_2986_0,
    i_13_421_2987_0, i_13_421_3031_0, i_13_421_3032_0, i_13_421_3064_0,
    i_13_421_3074_0, i_13_421_3208_0, i_13_421_3209_0, i_13_421_3235_0,
    i_13_421_3265_0, i_13_421_3293_0, i_13_421_3347_0, i_13_421_3382_0,
    i_13_421_3401_0, i_13_421_3427_0, i_13_421_3506_0, i_13_421_3526_0,
    i_13_421_3681_0, i_13_421_3824_0, i_13_421_3861_0, i_13_421_3911_0,
    i_13_421_3913_0, i_13_421_4338_0, i_13_421_4396_0, i_13_421_4514_0,
    i_13_421_4540_0, i_13_421_4567_0, i_13_421_4598_0, i_13_421_4607_0;
  output o_13_421_0_0;
  assign o_13_421_0_0 = ~((~i_13_421_1645_0 & (~i_13_421_2987_0 | (~i_13_421_188_0 & ~i_13_421_898_0))) | (~i_13_421_3911_0 & (~i_13_421_1804_0 | ~i_13_421_2983_0)) | (~i_13_421_1808_0 & ~i_13_421_1858_0) | (~i_13_421_1411_0 & ~i_13_421_3913_0 & ~i_13_421_4514_0) | (i_13_421_3235_0 & ~i_13_421_4567_0));
endmodule



// Benchmark "kernel_13_422" written by ABC on Sun Jul 19 10:51:14 2020

module kernel_13_422 ( 
    i_13_422_37_0, i_13_422_38_0, i_13_422_51_0, i_13_422_76_0,
    i_13_422_77_0, i_13_422_371_0, i_13_422_382_0, i_13_422_518_0,
    i_13_422_603_0, i_13_422_625_0, i_13_422_660_0, i_13_422_661_0,
    i_13_422_663_0, i_13_422_771_0, i_13_422_792_0, i_13_422_794_0,
    i_13_422_825_0, i_13_422_861_0, i_13_422_910_0, i_13_422_942_0,
    i_13_422_983_0, i_13_422_1018_0, i_13_422_1066_0, i_13_422_1077_0,
    i_13_422_1082_0, i_13_422_1120_0, i_13_422_1227_0, i_13_422_1284_0,
    i_13_422_1397_0, i_13_422_1425_0, i_13_422_1428_0, i_13_422_1429_0,
    i_13_422_1433_0, i_13_422_1571_0, i_13_422_1605_0, i_13_422_1631_0,
    i_13_422_1659_0, i_13_422_1681_0, i_13_422_1695_0, i_13_422_1744_0,
    i_13_422_1776_0, i_13_422_1777_0, i_13_422_1919_0, i_13_422_2027_0,
    i_13_422_2137_0, i_13_422_2189_0, i_13_422_2197_0, i_13_422_2209_0,
    i_13_422_2263_0, i_13_422_2297_0, i_13_422_2407_0, i_13_422_2451_0,
    i_13_422_2454_0, i_13_422_2553_0, i_13_422_2614_0, i_13_422_2662_0,
    i_13_422_2765_0, i_13_422_2821_0, i_13_422_3011_0, i_13_422_3037_0,
    i_13_422_3049_0, i_13_422_3135_0, i_13_422_3217_0, i_13_422_3322_0,
    i_13_422_3345_0, i_13_422_3377_0, i_13_422_3389_0, i_13_422_3397_0,
    i_13_422_3418_0, i_13_422_3461_0, i_13_422_3489_0, i_13_422_3490_0,
    i_13_422_3504_0, i_13_422_3505_0, i_13_422_3508_0, i_13_422_3567_0,
    i_13_422_3568_0, i_13_422_3570_0, i_13_422_3612_0, i_13_422_3618_0,
    i_13_422_3638_0, i_13_422_3651_0, i_13_422_3739_0, i_13_422_3740_0,
    i_13_422_3741_0, i_13_422_3742_0, i_13_422_3866_0, i_13_422_3891_0,
    i_13_422_3894_0, i_13_422_3895_0, i_13_422_4054_0, i_13_422_4088_0,
    i_13_422_4233_0, i_13_422_4254_0, i_13_422_4282_0, i_13_422_4356_0,
    i_13_422_4366_0, i_13_422_4368_0, i_13_422_4369_0, i_13_422_4603_0,
    o_13_422_0_0  );
  input  i_13_422_37_0, i_13_422_38_0, i_13_422_51_0, i_13_422_76_0,
    i_13_422_77_0, i_13_422_371_0, i_13_422_382_0, i_13_422_518_0,
    i_13_422_603_0, i_13_422_625_0, i_13_422_660_0, i_13_422_661_0,
    i_13_422_663_0, i_13_422_771_0, i_13_422_792_0, i_13_422_794_0,
    i_13_422_825_0, i_13_422_861_0, i_13_422_910_0, i_13_422_942_0,
    i_13_422_983_0, i_13_422_1018_0, i_13_422_1066_0, i_13_422_1077_0,
    i_13_422_1082_0, i_13_422_1120_0, i_13_422_1227_0, i_13_422_1284_0,
    i_13_422_1397_0, i_13_422_1425_0, i_13_422_1428_0, i_13_422_1429_0,
    i_13_422_1433_0, i_13_422_1571_0, i_13_422_1605_0, i_13_422_1631_0,
    i_13_422_1659_0, i_13_422_1681_0, i_13_422_1695_0, i_13_422_1744_0,
    i_13_422_1776_0, i_13_422_1777_0, i_13_422_1919_0, i_13_422_2027_0,
    i_13_422_2137_0, i_13_422_2189_0, i_13_422_2197_0, i_13_422_2209_0,
    i_13_422_2263_0, i_13_422_2297_0, i_13_422_2407_0, i_13_422_2451_0,
    i_13_422_2454_0, i_13_422_2553_0, i_13_422_2614_0, i_13_422_2662_0,
    i_13_422_2765_0, i_13_422_2821_0, i_13_422_3011_0, i_13_422_3037_0,
    i_13_422_3049_0, i_13_422_3135_0, i_13_422_3217_0, i_13_422_3322_0,
    i_13_422_3345_0, i_13_422_3377_0, i_13_422_3389_0, i_13_422_3397_0,
    i_13_422_3418_0, i_13_422_3461_0, i_13_422_3489_0, i_13_422_3490_0,
    i_13_422_3504_0, i_13_422_3505_0, i_13_422_3508_0, i_13_422_3567_0,
    i_13_422_3568_0, i_13_422_3570_0, i_13_422_3612_0, i_13_422_3618_0,
    i_13_422_3638_0, i_13_422_3651_0, i_13_422_3739_0, i_13_422_3740_0,
    i_13_422_3741_0, i_13_422_3742_0, i_13_422_3866_0, i_13_422_3891_0,
    i_13_422_3894_0, i_13_422_3895_0, i_13_422_4054_0, i_13_422_4088_0,
    i_13_422_4233_0, i_13_422_4254_0, i_13_422_4282_0, i_13_422_4356_0,
    i_13_422_4366_0, i_13_422_4368_0, i_13_422_4369_0, i_13_422_4603_0;
  output o_13_422_0_0;
  assign o_13_422_0_0 = ~((~i_13_422_3651_0 & ~i_13_422_4369_0) | (i_13_422_1066_0 & i_13_422_4054_0) | (~i_13_422_1425_0 & ~i_13_422_3742_0) | (~i_13_422_518_0 & i_13_422_2407_0 & ~i_13_422_4254_0) | (~i_13_422_1429_0 & ~i_13_422_2197_0 & ~i_13_422_3567_0 & ~i_13_422_4366_0) | (~i_13_422_1077_0 & ~i_13_422_1227_0 & ~i_13_422_3397_0 & ~i_13_422_3490_0));
endmodule



// Benchmark "kernel_13_423" written by ABC on Sun Jul 19 10:51:15 2020

module kernel_13_423 ( 
    i_13_423_38_0, i_13_423_193_0, i_13_423_209_0, i_13_423_274_0,
    i_13_423_284_0, i_13_423_287_0, i_13_423_310_0, i_13_423_317_0,
    i_13_423_382_0, i_13_423_525_0, i_13_423_528_0, i_13_423_529_0,
    i_13_423_561_0, i_13_423_679_0, i_13_423_682_0, i_13_423_826_0,
    i_13_423_852_0, i_13_423_863_0, i_13_423_914_0, i_13_423_979_0,
    i_13_423_1021_0, i_13_423_1022_0, i_13_423_1212_0, i_13_423_1227_0,
    i_13_423_1311_0, i_13_423_1312_0, i_13_423_1317_0, i_13_423_1327_0,
    i_13_423_1363_0, i_13_423_1429_0, i_13_423_1528_0, i_13_423_1565_0,
    i_13_423_1678_0, i_13_423_1726_0, i_13_423_1740_0, i_13_423_1780_0,
    i_13_423_1781_0, i_13_423_1871_0, i_13_423_1885_0, i_13_423_1886_0,
    i_13_423_1888_0, i_13_423_1960_0, i_13_423_2005_0, i_13_423_2108_0,
    i_13_423_2136_0, i_13_423_2146_0, i_13_423_2173_0, i_13_423_2261_0,
    i_13_423_2267_0, i_13_423_2302_0, i_13_423_2350_0, i_13_423_2394_0,
    i_13_423_2420_0, i_13_423_2462_0, i_13_423_2464_0, i_13_423_2470_0,
    i_13_423_2561_0, i_13_423_2653_0, i_13_423_2676_0, i_13_423_2740_0,
    i_13_423_2904_0, i_13_423_2962_0, i_13_423_3005_0, i_13_423_3012_0,
    i_13_423_3058_0, i_13_423_3100_0, i_13_423_3128_0, i_13_423_3130_0,
    i_13_423_3146_0, i_13_423_3197_0, i_13_423_3199_0, i_13_423_3262_0,
    i_13_423_3352_0, i_13_423_3509_0, i_13_423_3526_0, i_13_423_3541_0,
    i_13_423_3613_0, i_13_423_3614_0, i_13_423_3649_0, i_13_423_3709_0,
    i_13_423_3729_0, i_13_423_3730_0, i_13_423_3731_0, i_13_423_3733_0,
    i_13_423_3769_0, i_13_423_3854_0, i_13_423_3895_0, i_13_423_3913_0,
    i_13_423_4017_0, i_13_423_4057_0, i_13_423_4126_0, i_13_423_4255_0,
    i_13_423_4263_0, i_13_423_4264_0, i_13_423_4399_0, i_13_423_4432_0,
    i_13_423_4513_0, i_13_423_4557_0, i_13_423_4567_0, i_13_423_4597_0,
    o_13_423_0_0  );
  input  i_13_423_38_0, i_13_423_193_0, i_13_423_209_0, i_13_423_274_0,
    i_13_423_284_0, i_13_423_287_0, i_13_423_310_0, i_13_423_317_0,
    i_13_423_382_0, i_13_423_525_0, i_13_423_528_0, i_13_423_529_0,
    i_13_423_561_0, i_13_423_679_0, i_13_423_682_0, i_13_423_826_0,
    i_13_423_852_0, i_13_423_863_0, i_13_423_914_0, i_13_423_979_0,
    i_13_423_1021_0, i_13_423_1022_0, i_13_423_1212_0, i_13_423_1227_0,
    i_13_423_1311_0, i_13_423_1312_0, i_13_423_1317_0, i_13_423_1327_0,
    i_13_423_1363_0, i_13_423_1429_0, i_13_423_1528_0, i_13_423_1565_0,
    i_13_423_1678_0, i_13_423_1726_0, i_13_423_1740_0, i_13_423_1780_0,
    i_13_423_1781_0, i_13_423_1871_0, i_13_423_1885_0, i_13_423_1886_0,
    i_13_423_1888_0, i_13_423_1960_0, i_13_423_2005_0, i_13_423_2108_0,
    i_13_423_2136_0, i_13_423_2146_0, i_13_423_2173_0, i_13_423_2261_0,
    i_13_423_2267_0, i_13_423_2302_0, i_13_423_2350_0, i_13_423_2394_0,
    i_13_423_2420_0, i_13_423_2462_0, i_13_423_2464_0, i_13_423_2470_0,
    i_13_423_2561_0, i_13_423_2653_0, i_13_423_2676_0, i_13_423_2740_0,
    i_13_423_2904_0, i_13_423_2962_0, i_13_423_3005_0, i_13_423_3012_0,
    i_13_423_3058_0, i_13_423_3100_0, i_13_423_3128_0, i_13_423_3130_0,
    i_13_423_3146_0, i_13_423_3197_0, i_13_423_3199_0, i_13_423_3262_0,
    i_13_423_3352_0, i_13_423_3509_0, i_13_423_3526_0, i_13_423_3541_0,
    i_13_423_3613_0, i_13_423_3614_0, i_13_423_3649_0, i_13_423_3709_0,
    i_13_423_3729_0, i_13_423_3730_0, i_13_423_3731_0, i_13_423_3733_0,
    i_13_423_3769_0, i_13_423_3854_0, i_13_423_3895_0, i_13_423_3913_0,
    i_13_423_4017_0, i_13_423_4057_0, i_13_423_4126_0, i_13_423_4255_0,
    i_13_423_4263_0, i_13_423_4264_0, i_13_423_4399_0, i_13_423_4432_0,
    i_13_423_4513_0, i_13_423_4557_0, i_13_423_4567_0, i_13_423_4597_0;
  output o_13_423_0_0;
  assign o_13_423_0_0 = ~(~i_13_423_3541_0 | ~i_13_423_528_0 | (i_13_423_2464_0 & ~i_13_423_4264_0));
endmodule



// Benchmark "kernel_13_424" written by ABC on Sun Jul 19 10:51:16 2020

module kernel_13_424 ( 
    i_13_424_52_0, i_13_424_68_0, i_13_424_71_0, i_13_424_140_0,
    i_13_424_143_0, i_13_424_177_0, i_13_424_230_0, i_13_424_309_0,
    i_13_424_364_0, i_13_424_539_0, i_13_424_608_0, i_13_424_610_0,
    i_13_424_646_0, i_13_424_647_0, i_13_424_652_0, i_13_424_674_0,
    i_13_424_689_0, i_13_424_764_0, i_13_424_851_0, i_13_424_887_0,
    i_13_424_935_0, i_13_424_938_0, i_13_424_995_0, i_13_424_1117_0,
    i_13_424_1123_0, i_13_424_1124_0, i_13_424_1133_0, i_13_424_1145_0,
    i_13_424_1270_0, i_13_424_1277_0, i_13_424_1286_0, i_13_424_1342_0,
    i_13_424_1364_0, i_13_424_1403_0, i_13_424_1445_0, i_13_424_1472_0,
    i_13_424_1511_0, i_13_424_1660_0, i_13_424_1733_0, i_13_424_1735_0,
    i_13_424_1736_0, i_13_424_1768_0, i_13_424_1796_0, i_13_424_1798_0,
    i_13_424_1799_0, i_13_424_1809_0, i_13_424_1833_0, i_13_424_1920_0,
    i_13_424_1944_0, i_13_424_2052_0, i_13_424_2059_0, i_13_424_2115_0,
    i_13_424_2134_0, i_13_424_2265_0, i_13_424_2403_0, i_13_424_2406_0,
    i_13_424_2429_0, i_13_424_2462_0, i_13_424_2555_0, i_13_424_2679_0,
    i_13_424_2694_0, i_13_424_2725_0, i_13_424_2851_0, i_13_424_2852_0,
    i_13_424_2885_0, i_13_424_2983_0, i_13_424_3044_0, i_13_424_3050_0,
    i_13_424_3157_0, i_13_424_3208_0, i_13_424_3265_0, i_13_424_3339_0,
    i_13_424_3356_0, i_13_424_3371_0, i_13_424_3438_0, i_13_424_3451_0,
    i_13_424_3522_0, i_13_424_3532_0, i_13_424_3568_0, i_13_424_3569_0,
    i_13_424_3611_0, i_13_424_3653_0, i_13_424_3743_0, i_13_424_3787_0,
    i_13_424_3896_0, i_13_424_3913_0, i_13_424_3914_0, i_13_424_3927_0,
    i_13_424_3930_0, i_13_424_3931_0, i_13_424_3932_0, i_13_424_4040_0,
    i_13_424_4063_0, i_13_424_4190_0, i_13_424_4261_0, i_13_424_4279_0,
    i_13_424_4297_0, i_13_424_4298_0, i_13_424_4597_0, i_13_424_4598_0,
    o_13_424_0_0  );
  input  i_13_424_52_0, i_13_424_68_0, i_13_424_71_0, i_13_424_140_0,
    i_13_424_143_0, i_13_424_177_0, i_13_424_230_0, i_13_424_309_0,
    i_13_424_364_0, i_13_424_539_0, i_13_424_608_0, i_13_424_610_0,
    i_13_424_646_0, i_13_424_647_0, i_13_424_652_0, i_13_424_674_0,
    i_13_424_689_0, i_13_424_764_0, i_13_424_851_0, i_13_424_887_0,
    i_13_424_935_0, i_13_424_938_0, i_13_424_995_0, i_13_424_1117_0,
    i_13_424_1123_0, i_13_424_1124_0, i_13_424_1133_0, i_13_424_1145_0,
    i_13_424_1270_0, i_13_424_1277_0, i_13_424_1286_0, i_13_424_1342_0,
    i_13_424_1364_0, i_13_424_1403_0, i_13_424_1445_0, i_13_424_1472_0,
    i_13_424_1511_0, i_13_424_1660_0, i_13_424_1733_0, i_13_424_1735_0,
    i_13_424_1736_0, i_13_424_1768_0, i_13_424_1796_0, i_13_424_1798_0,
    i_13_424_1799_0, i_13_424_1809_0, i_13_424_1833_0, i_13_424_1920_0,
    i_13_424_1944_0, i_13_424_2052_0, i_13_424_2059_0, i_13_424_2115_0,
    i_13_424_2134_0, i_13_424_2265_0, i_13_424_2403_0, i_13_424_2406_0,
    i_13_424_2429_0, i_13_424_2462_0, i_13_424_2555_0, i_13_424_2679_0,
    i_13_424_2694_0, i_13_424_2725_0, i_13_424_2851_0, i_13_424_2852_0,
    i_13_424_2885_0, i_13_424_2983_0, i_13_424_3044_0, i_13_424_3050_0,
    i_13_424_3157_0, i_13_424_3208_0, i_13_424_3265_0, i_13_424_3339_0,
    i_13_424_3356_0, i_13_424_3371_0, i_13_424_3438_0, i_13_424_3451_0,
    i_13_424_3522_0, i_13_424_3532_0, i_13_424_3568_0, i_13_424_3569_0,
    i_13_424_3611_0, i_13_424_3653_0, i_13_424_3743_0, i_13_424_3787_0,
    i_13_424_3896_0, i_13_424_3913_0, i_13_424_3914_0, i_13_424_3927_0,
    i_13_424_3930_0, i_13_424_3931_0, i_13_424_3932_0, i_13_424_4040_0,
    i_13_424_4063_0, i_13_424_4190_0, i_13_424_4261_0, i_13_424_4279_0,
    i_13_424_4297_0, i_13_424_4298_0, i_13_424_4597_0, i_13_424_4598_0;
  output o_13_424_0_0;
  assign o_13_424_0_0 = ~((~i_13_424_935_0 & ((~i_13_424_1277_0 & ~i_13_424_1660_0) | (~i_13_424_1511_0 & ~i_13_424_3569_0))) | (~i_13_424_3932_0 & ((~i_13_424_1403_0 & ~i_13_424_2852_0 & i_13_424_3208_0) | (~i_13_424_2885_0 & ~i_13_424_3208_0))) | (i_13_424_689_0 & ~i_13_424_1123_0) | (~i_13_424_887_0 & ~i_13_424_1277_0 & i_13_424_4190_0));
endmodule



// Benchmark "kernel_13_425" written by ABC on Sun Jul 19 10:51:17 2020

module kernel_13_425 ( 
    i_13_425_28_0, i_13_425_31_0, i_13_425_67_0, i_13_425_136_0,
    i_13_425_157_0, i_13_425_184_0, i_13_425_193_0, i_13_425_206_0,
    i_13_425_266_0, i_13_425_316_0, i_13_425_335_0, i_13_425_338_0,
    i_13_425_373_0, i_13_425_381_0, i_13_425_383_0, i_13_425_459_0,
    i_13_425_543_0, i_13_425_581_0, i_13_425_590_0, i_13_425_715_0,
    i_13_425_742_0, i_13_425_746_0, i_13_425_795_0, i_13_425_813_0,
    i_13_425_870_0, i_13_425_1075_0, i_13_425_1120_0, i_13_425_1134_0,
    i_13_425_1216_0, i_13_425_1282_0, i_13_425_1300_0, i_13_425_1301_0,
    i_13_425_1327_0, i_13_425_1345_0, i_13_425_1400_0, i_13_425_1408_0,
    i_13_425_1444_0, i_13_425_1489_0, i_13_425_1495_0, i_13_425_1603_0,
    i_13_425_1633_0, i_13_425_1678_0, i_13_425_1717_0, i_13_425_1718_0,
    i_13_425_1811_0, i_13_425_1813_0, i_13_425_1831_0, i_13_425_1858_0,
    i_13_425_1993_0, i_13_425_1997_0, i_13_425_2056_0, i_13_425_2191_0,
    i_13_425_2208_0, i_13_425_2399_0, i_13_425_2480_0, i_13_425_2539_0,
    i_13_425_2540_0, i_13_425_2575_0, i_13_425_2632_0, i_13_425_2719_0,
    i_13_425_2721_0, i_13_425_2723_0, i_13_425_2857_0, i_13_425_2858_0,
    i_13_425_2860_0, i_13_425_2916_0, i_13_425_2970_0, i_13_425_2998_0,
    i_13_425_3016_0, i_13_425_3019_0, i_13_425_3061_0, i_13_425_3232_0,
    i_13_425_3235_0, i_13_425_3439_0, i_13_425_3441_0, i_13_425_3490_0,
    i_13_425_3615_0, i_13_425_3616_0, i_13_425_3619_0, i_13_425_3631_0,
    i_13_425_3666_0, i_13_425_3683_0, i_13_425_3685_0, i_13_425_3700_0,
    i_13_425_3727_0, i_13_425_3766_0, i_13_425_3844_0, i_13_425_3892_0,
    i_13_425_3921_0, i_13_425_3974_0, i_13_425_4055_0, i_13_425_4184_0,
    i_13_425_4186_0, i_13_425_4235_0, i_13_425_4369_0, i_13_425_4378_0,
    i_13_425_4395_0, i_13_425_4396_0, i_13_425_4397_0, i_13_425_4521_0,
    o_13_425_0_0  );
  input  i_13_425_28_0, i_13_425_31_0, i_13_425_67_0, i_13_425_136_0,
    i_13_425_157_0, i_13_425_184_0, i_13_425_193_0, i_13_425_206_0,
    i_13_425_266_0, i_13_425_316_0, i_13_425_335_0, i_13_425_338_0,
    i_13_425_373_0, i_13_425_381_0, i_13_425_383_0, i_13_425_459_0,
    i_13_425_543_0, i_13_425_581_0, i_13_425_590_0, i_13_425_715_0,
    i_13_425_742_0, i_13_425_746_0, i_13_425_795_0, i_13_425_813_0,
    i_13_425_870_0, i_13_425_1075_0, i_13_425_1120_0, i_13_425_1134_0,
    i_13_425_1216_0, i_13_425_1282_0, i_13_425_1300_0, i_13_425_1301_0,
    i_13_425_1327_0, i_13_425_1345_0, i_13_425_1400_0, i_13_425_1408_0,
    i_13_425_1444_0, i_13_425_1489_0, i_13_425_1495_0, i_13_425_1603_0,
    i_13_425_1633_0, i_13_425_1678_0, i_13_425_1717_0, i_13_425_1718_0,
    i_13_425_1811_0, i_13_425_1813_0, i_13_425_1831_0, i_13_425_1858_0,
    i_13_425_1993_0, i_13_425_1997_0, i_13_425_2056_0, i_13_425_2191_0,
    i_13_425_2208_0, i_13_425_2399_0, i_13_425_2480_0, i_13_425_2539_0,
    i_13_425_2540_0, i_13_425_2575_0, i_13_425_2632_0, i_13_425_2719_0,
    i_13_425_2721_0, i_13_425_2723_0, i_13_425_2857_0, i_13_425_2858_0,
    i_13_425_2860_0, i_13_425_2916_0, i_13_425_2970_0, i_13_425_2998_0,
    i_13_425_3016_0, i_13_425_3019_0, i_13_425_3061_0, i_13_425_3232_0,
    i_13_425_3235_0, i_13_425_3439_0, i_13_425_3441_0, i_13_425_3490_0,
    i_13_425_3615_0, i_13_425_3616_0, i_13_425_3619_0, i_13_425_3631_0,
    i_13_425_3666_0, i_13_425_3683_0, i_13_425_3685_0, i_13_425_3700_0,
    i_13_425_3727_0, i_13_425_3766_0, i_13_425_3844_0, i_13_425_3892_0,
    i_13_425_3921_0, i_13_425_3974_0, i_13_425_4055_0, i_13_425_4184_0,
    i_13_425_4186_0, i_13_425_4235_0, i_13_425_4369_0, i_13_425_4378_0,
    i_13_425_4395_0, i_13_425_4396_0, i_13_425_4397_0, i_13_425_4521_0;
  output o_13_425_0_0;
  assign o_13_425_0_0 = ~((~i_13_425_383_0 & (i_13_425_1678_0 | (~i_13_425_2056_0 & ~i_13_425_2916_0 & ~i_13_425_3727_0))) | (i_13_425_1831_0 & ((~i_13_425_2860_0 & i_13_425_3921_0) | (i_13_425_1327_0 & ~i_13_425_3683_0 & ~i_13_425_3844_0 & ~i_13_425_3921_0 & ~i_13_425_4378_0 & ~i_13_425_4397_0))) | (~i_13_425_4396_0 & (i_13_425_4369_0 | (~i_13_425_1301_0 & ~i_13_425_1831_0))) | (~i_13_425_1993_0 & ~i_13_425_3619_0) | (~i_13_425_2857_0 & ~i_13_425_3727_0 & ~i_13_425_3844_0 & i_13_425_4055_0) | (~i_13_425_381_0 & ~i_13_425_590_0 & ~i_13_425_1345_0 & ~i_13_425_2208_0 & ~i_13_425_4235_0));
endmodule



// Benchmark "kernel_13_426" written by ABC on Sun Jul 19 10:51:18 2020

module kernel_13_426 ( 
    i_13_426_32_0, i_13_426_36_0, i_13_426_179_0, i_13_426_184_0,
    i_13_426_279_0, i_13_426_286_0, i_13_426_315_0, i_13_426_319_0,
    i_13_426_320_0, i_13_426_337_0, i_13_426_454_0, i_13_426_553_0,
    i_13_426_592_0, i_13_426_645_0, i_13_426_646_0, i_13_426_647_0,
    i_13_426_655_0, i_13_426_670_0, i_13_426_679_0, i_13_426_680_0,
    i_13_426_684_0, i_13_426_691_0, i_13_426_692_0, i_13_426_835_0,
    i_13_426_844_0, i_13_426_898_0, i_13_426_952_0, i_13_426_1116_0,
    i_13_426_1121_0, i_13_426_1123_0, i_13_426_1124_0, i_13_426_1260_0,
    i_13_426_1262_0, i_13_426_1267_0, i_13_426_1274_0, i_13_426_1301_0,
    i_13_426_1519_0, i_13_426_1532_0, i_13_426_1553_0, i_13_426_1597_0,
    i_13_426_1643_0, i_13_426_1743_0, i_13_426_1813_0, i_13_426_1854_0,
    i_13_426_2058_0, i_13_426_2059_0, i_13_426_2104_0, i_13_426_2133_0,
    i_13_426_2210_0, i_13_426_2284_0, i_13_426_2466_0, i_13_426_2617_0,
    i_13_426_2677_0, i_13_426_2678_0, i_13_426_2708_0, i_13_426_2756_0,
    i_13_426_2781_0, i_13_426_2845_0, i_13_426_3012_0, i_13_426_3113_0,
    i_13_426_3145_0, i_13_426_3217_0, i_13_426_3218_0, i_13_426_3322_0,
    i_13_426_3379_0, i_13_426_3383_0, i_13_426_3401_0, i_13_426_3412_0,
    i_13_426_3418_0, i_13_426_3476_0, i_13_426_3533_0, i_13_426_3535_0,
    i_13_426_3538_0, i_13_426_3574_0, i_13_426_3598_0, i_13_426_3701_0,
    i_13_426_3724_0, i_13_426_3735_0, i_13_426_3739_0, i_13_426_3769_0,
    i_13_426_3770_0, i_13_426_3867_0, i_13_426_3892_0, i_13_426_3928_0,
    i_13_426_3935_0, i_13_426_3992_0, i_13_426_4021_0, i_13_426_4022_0,
    i_13_426_4032_0, i_13_426_4077_0, i_13_426_4081_0, i_13_426_4085_0,
    i_13_426_4090_0, i_13_426_4185_0, i_13_426_4270_0, i_13_426_4534_0,
    i_13_426_4586_0, i_13_426_4594_0, i_13_426_4595_0, i_13_426_4598_0,
    o_13_426_0_0  );
  input  i_13_426_32_0, i_13_426_36_0, i_13_426_179_0, i_13_426_184_0,
    i_13_426_279_0, i_13_426_286_0, i_13_426_315_0, i_13_426_319_0,
    i_13_426_320_0, i_13_426_337_0, i_13_426_454_0, i_13_426_553_0,
    i_13_426_592_0, i_13_426_645_0, i_13_426_646_0, i_13_426_647_0,
    i_13_426_655_0, i_13_426_670_0, i_13_426_679_0, i_13_426_680_0,
    i_13_426_684_0, i_13_426_691_0, i_13_426_692_0, i_13_426_835_0,
    i_13_426_844_0, i_13_426_898_0, i_13_426_952_0, i_13_426_1116_0,
    i_13_426_1121_0, i_13_426_1123_0, i_13_426_1124_0, i_13_426_1260_0,
    i_13_426_1262_0, i_13_426_1267_0, i_13_426_1274_0, i_13_426_1301_0,
    i_13_426_1519_0, i_13_426_1532_0, i_13_426_1553_0, i_13_426_1597_0,
    i_13_426_1643_0, i_13_426_1743_0, i_13_426_1813_0, i_13_426_1854_0,
    i_13_426_2058_0, i_13_426_2059_0, i_13_426_2104_0, i_13_426_2133_0,
    i_13_426_2210_0, i_13_426_2284_0, i_13_426_2466_0, i_13_426_2617_0,
    i_13_426_2677_0, i_13_426_2678_0, i_13_426_2708_0, i_13_426_2756_0,
    i_13_426_2781_0, i_13_426_2845_0, i_13_426_3012_0, i_13_426_3113_0,
    i_13_426_3145_0, i_13_426_3217_0, i_13_426_3218_0, i_13_426_3322_0,
    i_13_426_3379_0, i_13_426_3383_0, i_13_426_3401_0, i_13_426_3412_0,
    i_13_426_3418_0, i_13_426_3476_0, i_13_426_3533_0, i_13_426_3535_0,
    i_13_426_3538_0, i_13_426_3574_0, i_13_426_3598_0, i_13_426_3701_0,
    i_13_426_3724_0, i_13_426_3735_0, i_13_426_3739_0, i_13_426_3769_0,
    i_13_426_3770_0, i_13_426_3867_0, i_13_426_3892_0, i_13_426_3928_0,
    i_13_426_3935_0, i_13_426_3992_0, i_13_426_4021_0, i_13_426_4022_0,
    i_13_426_4032_0, i_13_426_4077_0, i_13_426_4081_0, i_13_426_4085_0,
    i_13_426_4090_0, i_13_426_4185_0, i_13_426_4270_0, i_13_426_4534_0,
    i_13_426_4586_0, i_13_426_4594_0, i_13_426_4595_0, i_13_426_4598_0;
  output o_13_426_0_0;
  assign o_13_426_0_0 = ~((~i_13_426_2058_0 & ((~i_13_426_898_0 & ~i_13_426_1116_0 & ~i_13_426_1124_0 & ~i_13_426_2284_0 & ~i_13_426_2845_0 & ~i_13_426_3574_0) | (~i_13_426_315_0 & ~i_13_426_320_0 & ~i_13_426_679_0 & ~i_13_426_3598_0))) | i_13_426_337_0 | (~i_13_426_179_0 & ~i_13_426_684_0 & ~i_13_426_844_0 & ~i_13_426_3892_0) | (~i_13_426_286_0 & ~i_13_426_670_0 & ~i_13_426_4085_0));
endmodule



// Benchmark "kernel_13_427" written by ABC on Sun Jul 19 10:51:18 2020

module kernel_13_427 ( 
    i_13_427_44_0, i_13_427_61_0, i_13_427_76_0, i_13_427_113_0,
    i_13_427_184_0, i_13_427_187_0, i_13_427_231_0, i_13_427_313_0,
    i_13_427_314_0, i_13_427_321_0, i_13_427_382_0, i_13_427_538_0,
    i_13_427_556_0, i_13_427_574_0, i_13_427_643_0, i_13_427_645_0,
    i_13_427_646_0, i_13_427_647_0, i_13_427_687_0, i_13_427_745_0,
    i_13_427_840_0, i_13_427_853_0, i_13_427_897_0, i_13_427_898_0,
    i_13_427_956_0, i_13_427_1021_0, i_13_427_1058_0, i_13_427_1112_0,
    i_13_427_1120_0, i_13_427_1121_0, i_13_427_1122_0, i_13_427_1123_0,
    i_13_427_1135_0, i_13_427_1275_0, i_13_427_1276_0, i_13_427_1426_0,
    i_13_427_1472_0, i_13_427_1516_0, i_13_427_1624_0, i_13_427_1633_0,
    i_13_427_1642_0, i_13_427_1643_0, i_13_427_1646_0, i_13_427_1678_0,
    i_13_427_1680_0, i_13_427_1716_0, i_13_427_1752_0, i_13_427_1789_0,
    i_13_427_1790_0, i_13_427_1800_0, i_13_427_1802_0, i_13_427_1804_0,
    i_13_427_1807_0, i_13_427_1816_0, i_13_427_1834_0, i_13_427_1853_0,
    i_13_427_1858_0, i_13_427_1861_0, i_13_427_1862_0, i_13_427_2002_0,
    i_13_427_2005_0, i_13_427_2057_0, i_13_427_2200_0, i_13_427_2213_0,
    i_13_427_2266_0, i_13_427_2267_0, i_13_427_2407_0, i_13_427_2408_0,
    i_13_427_2452_0, i_13_427_2528_0, i_13_427_2535_0, i_13_427_2542_0,
    i_13_427_2617_0, i_13_427_2697_0, i_13_427_2722_0, i_13_427_2850_0,
    i_13_427_2851_0, i_13_427_2903_0, i_13_427_2923_0, i_13_427_2965_0,
    i_13_427_2981_0, i_13_427_3028_0, i_13_427_3031_0, i_13_427_3065_0,
    i_13_427_3156_0, i_13_427_3292_0, i_13_427_3419_0, i_13_427_3703_0,
    i_13_427_3931_0, i_13_427_3993_0, i_13_427_3995_0, i_13_427_4044_0,
    i_13_427_4189_0, i_13_427_4190_0, i_13_427_4266_0, i_13_427_4297_0,
    i_13_427_4312_0, i_13_427_4356_0, i_13_427_4435_0, i_13_427_4598_0,
    o_13_427_0_0  );
  input  i_13_427_44_0, i_13_427_61_0, i_13_427_76_0, i_13_427_113_0,
    i_13_427_184_0, i_13_427_187_0, i_13_427_231_0, i_13_427_313_0,
    i_13_427_314_0, i_13_427_321_0, i_13_427_382_0, i_13_427_538_0,
    i_13_427_556_0, i_13_427_574_0, i_13_427_643_0, i_13_427_645_0,
    i_13_427_646_0, i_13_427_647_0, i_13_427_687_0, i_13_427_745_0,
    i_13_427_840_0, i_13_427_853_0, i_13_427_897_0, i_13_427_898_0,
    i_13_427_956_0, i_13_427_1021_0, i_13_427_1058_0, i_13_427_1112_0,
    i_13_427_1120_0, i_13_427_1121_0, i_13_427_1122_0, i_13_427_1123_0,
    i_13_427_1135_0, i_13_427_1275_0, i_13_427_1276_0, i_13_427_1426_0,
    i_13_427_1472_0, i_13_427_1516_0, i_13_427_1624_0, i_13_427_1633_0,
    i_13_427_1642_0, i_13_427_1643_0, i_13_427_1646_0, i_13_427_1678_0,
    i_13_427_1680_0, i_13_427_1716_0, i_13_427_1752_0, i_13_427_1789_0,
    i_13_427_1790_0, i_13_427_1800_0, i_13_427_1802_0, i_13_427_1804_0,
    i_13_427_1807_0, i_13_427_1816_0, i_13_427_1834_0, i_13_427_1853_0,
    i_13_427_1858_0, i_13_427_1861_0, i_13_427_1862_0, i_13_427_2002_0,
    i_13_427_2005_0, i_13_427_2057_0, i_13_427_2200_0, i_13_427_2213_0,
    i_13_427_2266_0, i_13_427_2267_0, i_13_427_2407_0, i_13_427_2408_0,
    i_13_427_2452_0, i_13_427_2528_0, i_13_427_2535_0, i_13_427_2542_0,
    i_13_427_2617_0, i_13_427_2697_0, i_13_427_2722_0, i_13_427_2850_0,
    i_13_427_2851_0, i_13_427_2903_0, i_13_427_2923_0, i_13_427_2965_0,
    i_13_427_2981_0, i_13_427_3028_0, i_13_427_3031_0, i_13_427_3065_0,
    i_13_427_3156_0, i_13_427_3292_0, i_13_427_3419_0, i_13_427_3703_0,
    i_13_427_3931_0, i_13_427_3993_0, i_13_427_3995_0, i_13_427_4044_0,
    i_13_427_4189_0, i_13_427_4190_0, i_13_427_4266_0, i_13_427_4297_0,
    i_13_427_4312_0, i_13_427_4356_0, i_13_427_4435_0, i_13_427_4598_0;
  output o_13_427_0_0;
  assign o_13_427_0_0 = ~((~i_13_427_1276_0 & ((i_13_427_61_0 & ~i_13_427_1472_0 & ~i_13_427_2535_0) | (~i_13_427_1646_0 & ~i_13_427_3993_0 & ~i_13_427_4435_0))) | (i_13_427_2923_0 & (i_13_427_2452_0 | (~i_13_427_61_0 & i_13_427_3065_0))) | (~i_13_427_313_0 & ~i_13_427_1678_0) | (~i_13_427_187_0 & ~i_13_427_1122_0 & ~i_13_427_4190_0));
endmodule



// Benchmark "kernel_13_428" written by ABC on Sun Jul 19 10:51:19 2020

module kernel_13_428 ( 
    i_13_428_41_0, i_13_428_67_0, i_13_428_135_0, i_13_428_136_0,
    i_13_428_137_0, i_13_428_138_0, i_13_428_139_0, i_13_428_166_0,
    i_13_428_181_0, i_13_428_283_0, i_13_428_373_0, i_13_428_489_0,
    i_13_428_493_0, i_13_428_535_0, i_13_428_539_0, i_13_428_621_0,
    i_13_428_625_0, i_13_428_694_0, i_13_428_695_0, i_13_428_696_0,
    i_13_428_814_0, i_13_428_856_0, i_13_428_864_0, i_13_428_884_0,
    i_13_428_1020_0, i_13_428_1021_0, i_13_428_1092_0, i_13_428_1129_0,
    i_13_428_1137_0, i_13_428_1218_0, i_13_428_1232_0, i_13_428_1306_0,
    i_13_428_1307_0, i_13_428_1404_0, i_13_428_1428_0, i_13_428_1431_0,
    i_13_428_1484_0, i_13_428_1516_0, i_13_428_1742_0, i_13_428_1759_0,
    i_13_428_1769_0, i_13_428_1795_0, i_13_428_1849_0, i_13_428_1882_0,
    i_13_428_1904_0, i_13_428_1947_0, i_13_428_1954_0, i_13_428_2119_0,
    i_13_428_2170_0, i_13_428_2200_0, i_13_428_2310_0, i_13_428_2354_0,
    i_13_428_2377_0, i_13_428_2407_0, i_13_428_2410_0, i_13_428_2445_0,
    i_13_428_2493_0, i_13_428_2505_0, i_13_428_2542_0, i_13_428_2720_0,
    i_13_428_2848_0, i_13_428_2849_0, i_13_428_2854_0, i_13_428_2872_0,
    i_13_428_2882_0, i_13_428_2997_0, i_13_428_2998_0, i_13_428_3021_0,
    i_13_428_3065_0, i_13_428_3109_0, i_13_428_3110_0, i_13_428_3130_0,
    i_13_428_3170_0, i_13_428_3371_0, i_13_428_3381_0, i_13_428_3481_0,
    i_13_428_3555_0, i_13_428_3684_0, i_13_428_3703_0, i_13_428_3723_0,
    i_13_428_3739_0, i_13_428_3740_0, i_13_428_3766_0, i_13_428_3818_0,
    i_13_428_3820_0, i_13_428_3836_0, i_13_428_3910_0, i_13_428_4006_0,
    i_13_428_4018_0, i_13_428_4063_0, i_13_428_4078_0, i_13_428_4152_0,
    i_13_428_4250_0, i_13_428_4294_0, i_13_428_4295_0, i_13_428_4316_0,
    i_13_428_4328_0, i_13_428_4341_0, i_13_428_4567_0, i_13_428_4581_0,
    o_13_428_0_0  );
  input  i_13_428_41_0, i_13_428_67_0, i_13_428_135_0, i_13_428_136_0,
    i_13_428_137_0, i_13_428_138_0, i_13_428_139_0, i_13_428_166_0,
    i_13_428_181_0, i_13_428_283_0, i_13_428_373_0, i_13_428_489_0,
    i_13_428_493_0, i_13_428_535_0, i_13_428_539_0, i_13_428_621_0,
    i_13_428_625_0, i_13_428_694_0, i_13_428_695_0, i_13_428_696_0,
    i_13_428_814_0, i_13_428_856_0, i_13_428_864_0, i_13_428_884_0,
    i_13_428_1020_0, i_13_428_1021_0, i_13_428_1092_0, i_13_428_1129_0,
    i_13_428_1137_0, i_13_428_1218_0, i_13_428_1232_0, i_13_428_1306_0,
    i_13_428_1307_0, i_13_428_1404_0, i_13_428_1428_0, i_13_428_1431_0,
    i_13_428_1484_0, i_13_428_1516_0, i_13_428_1742_0, i_13_428_1759_0,
    i_13_428_1769_0, i_13_428_1795_0, i_13_428_1849_0, i_13_428_1882_0,
    i_13_428_1904_0, i_13_428_1947_0, i_13_428_1954_0, i_13_428_2119_0,
    i_13_428_2170_0, i_13_428_2200_0, i_13_428_2310_0, i_13_428_2354_0,
    i_13_428_2377_0, i_13_428_2407_0, i_13_428_2410_0, i_13_428_2445_0,
    i_13_428_2493_0, i_13_428_2505_0, i_13_428_2542_0, i_13_428_2720_0,
    i_13_428_2848_0, i_13_428_2849_0, i_13_428_2854_0, i_13_428_2872_0,
    i_13_428_2882_0, i_13_428_2997_0, i_13_428_2998_0, i_13_428_3021_0,
    i_13_428_3065_0, i_13_428_3109_0, i_13_428_3110_0, i_13_428_3130_0,
    i_13_428_3170_0, i_13_428_3371_0, i_13_428_3381_0, i_13_428_3481_0,
    i_13_428_3555_0, i_13_428_3684_0, i_13_428_3703_0, i_13_428_3723_0,
    i_13_428_3739_0, i_13_428_3740_0, i_13_428_3766_0, i_13_428_3818_0,
    i_13_428_3820_0, i_13_428_3836_0, i_13_428_3910_0, i_13_428_4006_0,
    i_13_428_4018_0, i_13_428_4063_0, i_13_428_4078_0, i_13_428_4152_0,
    i_13_428_4250_0, i_13_428_4294_0, i_13_428_4295_0, i_13_428_4316_0,
    i_13_428_4328_0, i_13_428_4341_0, i_13_428_4567_0, i_13_428_4581_0;
  output o_13_428_0_0;
  assign o_13_428_0_0 = ~((~i_13_428_3739_0 & ((~i_13_428_2445_0 & ((i_13_428_283_0 & ~i_13_428_2377_0) | (~i_13_428_694_0 & ~i_13_428_2848_0 & ~i_13_428_3684_0 & ~i_13_428_3740_0))) | (~i_13_428_696_0 & i_13_428_814_0 & ~i_13_428_2848_0) | (~i_13_428_1428_0 & i_13_428_3684_0))) | (i_13_428_3109_0 & ((i_13_428_139_0 & ~i_13_428_1218_0 & i_13_428_3766_0 & ~i_13_428_4078_0) | (i_13_428_493_0 & i_13_428_4567_0) | (~i_13_428_535_0 & ~i_13_428_1795_0 & ~i_13_428_4567_0))) | (~i_13_428_489_0 & i_13_428_1428_0 & i_13_428_2542_0 & i_13_428_3910_0));
endmodule



// Benchmark "kernel_13_429" written by ABC on Sun Jul 19 10:51:20 2020

module kernel_13_429 ( 
    i_13_429_4_0, i_13_429_58_0, i_13_429_61_0, i_13_429_73_0,
    i_13_429_93_0, i_13_429_94_0, i_13_429_283_0, i_13_429_310_0,
    i_13_429_373_0, i_13_429_415_0, i_13_429_426_0, i_13_429_562_0,
    i_13_429_571_0, i_13_429_614_0, i_13_429_627_0, i_13_429_696_0,
    i_13_429_697_0, i_13_429_699_0, i_13_429_780_0, i_13_429_825_0,
    i_13_429_955_0, i_13_429_956_0, i_13_429_1006_0, i_13_429_1023_0,
    i_13_429_1071_0, i_13_429_1072_0, i_13_429_1098_0, i_13_429_1213_0,
    i_13_429_1225_0, i_13_429_1270_0, i_13_429_1301_0, i_13_429_1317_0,
    i_13_429_1318_0, i_13_429_1320_0, i_13_429_1380_0, i_13_429_1383_0,
    i_13_429_1428_0, i_13_429_1464_0, i_13_429_1479_0, i_13_429_1482_0,
    i_13_429_1483_0, i_13_429_1707_0, i_13_429_1721_0, i_13_429_1740_0,
    i_13_429_1759_0, i_13_429_1775_0, i_13_429_1795_0, i_13_429_1885_0,
    i_13_429_1888_0, i_13_429_1951_0, i_13_429_1957_0, i_13_429_2119_0,
    i_13_429_2244_0, i_13_429_2367_0, i_13_429_2407_0, i_13_429_2443_0,
    i_13_429_2444_0, i_13_429_2445_0, i_13_429_2446_0, i_13_429_2491_0,
    i_13_429_2512_0, i_13_429_2553_0, i_13_429_2554_0, i_13_429_2613_0,
    i_13_429_2676_0, i_13_429_2824_0, i_13_429_2857_0, i_13_429_2875_0,
    i_13_429_2964_0, i_13_429_2974_0, i_13_429_3093_0, i_13_429_3094_0,
    i_13_429_3119_0, i_13_429_3230_0, i_13_429_3235_0, i_13_429_3304_0,
    i_13_429_3307_0, i_13_429_3432_0, i_13_429_3479_0, i_13_429_3489_0,
    i_13_429_3540_0, i_13_429_3567_0, i_13_429_3580_0, i_13_429_3756_0,
    i_13_429_3820_0, i_13_429_3989_0, i_13_429_3991_0, i_13_429_4018_0,
    i_13_429_4205_0, i_13_429_4313_0, i_13_429_4315_0, i_13_429_4350_0,
    i_13_429_4353_0, i_13_429_4369_0, i_13_429_4378_0, i_13_429_4379_0,
    i_13_429_4380_0, i_13_429_4443_0, i_13_429_4498_0, i_13_429_4503_0,
    o_13_429_0_0  );
  input  i_13_429_4_0, i_13_429_58_0, i_13_429_61_0, i_13_429_73_0,
    i_13_429_93_0, i_13_429_94_0, i_13_429_283_0, i_13_429_310_0,
    i_13_429_373_0, i_13_429_415_0, i_13_429_426_0, i_13_429_562_0,
    i_13_429_571_0, i_13_429_614_0, i_13_429_627_0, i_13_429_696_0,
    i_13_429_697_0, i_13_429_699_0, i_13_429_780_0, i_13_429_825_0,
    i_13_429_955_0, i_13_429_956_0, i_13_429_1006_0, i_13_429_1023_0,
    i_13_429_1071_0, i_13_429_1072_0, i_13_429_1098_0, i_13_429_1213_0,
    i_13_429_1225_0, i_13_429_1270_0, i_13_429_1301_0, i_13_429_1317_0,
    i_13_429_1318_0, i_13_429_1320_0, i_13_429_1380_0, i_13_429_1383_0,
    i_13_429_1428_0, i_13_429_1464_0, i_13_429_1479_0, i_13_429_1482_0,
    i_13_429_1483_0, i_13_429_1707_0, i_13_429_1721_0, i_13_429_1740_0,
    i_13_429_1759_0, i_13_429_1775_0, i_13_429_1795_0, i_13_429_1885_0,
    i_13_429_1888_0, i_13_429_1951_0, i_13_429_1957_0, i_13_429_2119_0,
    i_13_429_2244_0, i_13_429_2367_0, i_13_429_2407_0, i_13_429_2443_0,
    i_13_429_2444_0, i_13_429_2445_0, i_13_429_2446_0, i_13_429_2491_0,
    i_13_429_2512_0, i_13_429_2553_0, i_13_429_2554_0, i_13_429_2613_0,
    i_13_429_2676_0, i_13_429_2824_0, i_13_429_2857_0, i_13_429_2875_0,
    i_13_429_2964_0, i_13_429_2974_0, i_13_429_3093_0, i_13_429_3094_0,
    i_13_429_3119_0, i_13_429_3230_0, i_13_429_3235_0, i_13_429_3304_0,
    i_13_429_3307_0, i_13_429_3432_0, i_13_429_3479_0, i_13_429_3489_0,
    i_13_429_3540_0, i_13_429_3567_0, i_13_429_3580_0, i_13_429_3756_0,
    i_13_429_3820_0, i_13_429_3989_0, i_13_429_3991_0, i_13_429_4018_0,
    i_13_429_4205_0, i_13_429_4313_0, i_13_429_4315_0, i_13_429_4350_0,
    i_13_429_4353_0, i_13_429_4369_0, i_13_429_4378_0, i_13_429_4379_0,
    i_13_429_4380_0, i_13_429_4443_0, i_13_429_4498_0, i_13_429_4503_0;
  output o_13_429_0_0;
  assign o_13_429_0_0 = ~((~i_13_429_697_0 & ((~i_13_429_696_0 & ~i_13_429_1320_0 & ~i_13_429_3567_0 & ~i_13_429_4369_0) | (i_13_429_4315_0 & i_13_429_4379_0))) | (~i_13_429_696_0 & ((i_13_429_571_0 & i_13_429_697_0 & ~i_13_429_3567_0 & ~i_13_429_3580_0 & ~i_13_429_4379_0) | (~i_13_429_1483_0 & ~i_13_429_2443_0 & ~i_13_429_4378_0 & ~i_13_429_4380_0))) | (~i_13_429_4353_0 & ((~i_13_429_571_0 & ~i_13_429_1885_0 & ~i_13_429_3540_0) | (~i_13_429_1225_0 & ~i_13_429_1301_0 & ~i_13_429_3093_0 & ~i_13_429_4315_0 & ~i_13_429_4379_0))) | (~i_13_429_4380_0 & ((~i_13_429_1023_0 & ~i_13_429_1071_0 & ~i_13_429_2875_0) | (~i_13_429_1795_0 & ~i_13_429_1957_0 & i_13_429_4315_0))) | (~i_13_429_426_0 & i_13_429_2407_0) | (i_13_429_94_0 & ~i_13_429_2244_0 & ~i_13_429_2613_0) | (~i_13_429_73_0 & i_13_429_283_0 & ~i_13_429_825_0 & ~i_13_429_1483_0 & ~i_13_429_3567_0));
endmodule



// Benchmark "kernel_13_430" written by ABC on Sun Jul 19 10:51:21 2020

module kernel_13_430 ( 
    i_13_430_33_0, i_13_430_114_0, i_13_430_159_0, i_13_430_183_0,
    i_13_430_384_0, i_13_430_385_0, i_13_430_406_0, i_13_430_537_0,
    i_13_430_570_0, i_13_430_571_0, i_13_430_589_0, i_13_430_591_0,
    i_13_430_681_0, i_13_430_724_0, i_13_430_760_0, i_13_430_762_0,
    i_13_430_795_0, i_13_430_816_0, i_13_430_913_0, i_13_430_931_0,
    i_13_430_942_0, i_13_430_1068_0, i_13_430_1084_0, i_13_430_1086_0,
    i_13_430_1266_0, i_13_430_1302_0, i_13_430_1303_0, i_13_430_1390_0,
    i_13_430_1408_0, i_13_430_1473_0, i_13_430_1509_0, i_13_430_1716_0,
    i_13_430_1788_0, i_13_430_1789_0, i_13_430_1803_0, i_13_430_1807_0,
    i_13_430_1815_0, i_13_430_1816_0, i_13_430_1951_0, i_13_430_1992_0,
    i_13_430_1995_0, i_13_430_1996_0, i_13_430_2001_0, i_13_430_2002_0,
    i_13_430_2122_0, i_13_430_2208_0, i_13_430_2226_0, i_13_430_2266_0,
    i_13_430_2424_0, i_13_430_2455_0, i_13_430_2472_0, i_13_430_2535_0,
    i_13_430_2541_0, i_13_430_2560_0, i_13_430_2577_0, i_13_430_2632_0,
    i_13_430_2790_0, i_13_430_2847_0, i_13_430_2919_0, i_13_430_2941_0,
    i_13_430_3003_0, i_13_430_3022_0, i_13_430_3031_0, i_13_430_3102_0,
    i_13_430_3126_0, i_13_430_3129_0, i_13_430_3147_0, i_13_430_3163_0,
    i_13_430_3265_0, i_13_430_3274_0, i_13_430_3328_0, i_13_430_3346_0,
    i_13_430_3381_0, i_13_430_3391_0, i_13_430_3399_0, i_13_430_3441_0,
    i_13_430_3453_0, i_13_430_3522_0, i_13_430_3535_0, i_13_430_3615_0,
    i_13_430_3624_0, i_13_430_3661_0, i_13_430_3702_0, i_13_430_3796_0,
    i_13_430_3846_0, i_13_430_3873_0, i_13_430_3928_0, i_13_430_3993_0,
    i_13_430_4057_0, i_13_430_4119_0, i_13_430_4165_0, i_13_430_4207_0,
    i_13_430_4236_0, i_13_430_4272_0, i_13_430_4273_0, i_13_430_4341_0,
    i_13_430_4399_0, i_13_430_4416_0, i_13_430_4417_0, i_13_430_4540_0,
    o_13_430_0_0  );
  input  i_13_430_33_0, i_13_430_114_0, i_13_430_159_0, i_13_430_183_0,
    i_13_430_384_0, i_13_430_385_0, i_13_430_406_0, i_13_430_537_0,
    i_13_430_570_0, i_13_430_571_0, i_13_430_589_0, i_13_430_591_0,
    i_13_430_681_0, i_13_430_724_0, i_13_430_760_0, i_13_430_762_0,
    i_13_430_795_0, i_13_430_816_0, i_13_430_913_0, i_13_430_931_0,
    i_13_430_942_0, i_13_430_1068_0, i_13_430_1084_0, i_13_430_1086_0,
    i_13_430_1266_0, i_13_430_1302_0, i_13_430_1303_0, i_13_430_1390_0,
    i_13_430_1408_0, i_13_430_1473_0, i_13_430_1509_0, i_13_430_1716_0,
    i_13_430_1788_0, i_13_430_1789_0, i_13_430_1803_0, i_13_430_1807_0,
    i_13_430_1815_0, i_13_430_1816_0, i_13_430_1951_0, i_13_430_1992_0,
    i_13_430_1995_0, i_13_430_1996_0, i_13_430_2001_0, i_13_430_2002_0,
    i_13_430_2122_0, i_13_430_2208_0, i_13_430_2226_0, i_13_430_2266_0,
    i_13_430_2424_0, i_13_430_2455_0, i_13_430_2472_0, i_13_430_2535_0,
    i_13_430_2541_0, i_13_430_2560_0, i_13_430_2577_0, i_13_430_2632_0,
    i_13_430_2790_0, i_13_430_2847_0, i_13_430_2919_0, i_13_430_2941_0,
    i_13_430_3003_0, i_13_430_3022_0, i_13_430_3031_0, i_13_430_3102_0,
    i_13_430_3126_0, i_13_430_3129_0, i_13_430_3147_0, i_13_430_3163_0,
    i_13_430_3265_0, i_13_430_3274_0, i_13_430_3328_0, i_13_430_3346_0,
    i_13_430_3381_0, i_13_430_3391_0, i_13_430_3399_0, i_13_430_3441_0,
    i_13_430_3453_0, i_13_430_3522_0, i_13_430_3535_0, i_13_430_3615_0,
    i_13_430_3624_0, i_13_430_3661_0, i_13_430_3702_0, i_13_430_3796_0,
    i_13_430_3846_0, i_13_430_3873_0, i_13_430_3928_0, i_13_430_3993_0,
    i_13_430_4057_0, i_13_430_4119_0, i_13_430_4165_0, i_13_430_4207_0,
    i_13_430_4236_0, i_13_430_4272_0, i_13_430_4273_0, i_13_430_4341_0,
    i_13_430_4399_0, i_13_430_4416_0, i_13_430_4417_0, i_13_430_4540_0;
  output o_13_430_0_0;
  assign o_13_430_0_0 = ~(~i_13_430_3346_0 | (~i_13_430_537_0 & i_13_430_4417_0) | (~i_13_430_1302_0 & ~i_13_430_1716_0) | (~i_13_430_1807_0 & ~i_13_430_3265_0 & ~i_13_430_3441_0 & i_13_430_4399_0));
endmodule



// Benchmark "kernel_13_431" written by ABC on Sun Jul 19 10:51:22 2020

module kernel_13_431 ( 
    i_13_431_37_0, i_13_431_93_0, i_13_431_102_0, i_13_431_138_0,
    i_13_431_139_0, i_13_431_174_0, i_13_431_229_0, i_13_431_267_0,
    i_13_431_373_0, i_13_431_505_0, i_13_431_549_0, i_13_431_550_0,
    i_13_431_603_0, i_13_431_604_0, i_13_431_657_0, i_13_431_660_0,
    i_13_431_661_0, i_13_431_663_0, i_13_431_669_0, i_13_431_675_0,
    i_13_431_676_0, i_13_431_855_0, i_13_431_1023_0, i_13_431_1072_0,
    i_13_431_1144_0, i_13_431_1219_0, i_13_431_1494_0, i_13_431_1515_0,
    i_13_431_1516_0, i_13_431_1521_0, i_13_431_1629_0, i_13_431_1630_0,
    i_13_431_1656_0, i_13_431_1711_0, i_13_431_1827_0, i_13_431_1828_0,
    i_13_431_1858_0, i_13_431_1881_0, i_13_431_1884_0, i_13_431_2001_0,
    i_13_431_2002_0, i_13_431_2016_0, i_13_431_2019_0, i_13_431_2020_0,
    i_13_431_2169_0, i_13_431_2340_0, i_13_431_2341_0, i_13_431_2362_0,
    i_13_431_2397_0, i_13_431_2398_0, i_13_431_2422_0, i_13_431_2448_0,
    i_13_431_2467_0, i_13_431_2497_0, i_13_431_2511_0, i_13_431_2611_0,
    i_13_431_2614_0, i_13_431_2718_0, i_13_431_2935_0, i_13_431_2982_0,
    i_13_431_3006_0, i_13_431_3009_0, i_13_431_3105_0, i_13_431_3108_0,
    i_13_431_3133_0, i_13_431_3159_0, i_13_431_3234_0, i_13_431_3385_0,
    i_13_431_3415_0, i_13_431_3475_0, i_13_431_3522_0, i_13_431_3639_0,
    i_13_431_3640_0, i_13_431_3738_0, i_13_431_3762_0, i_13_431_3763_0,
    i_13_431_3843_0, i_13_431_3861_0, i_13_431_3862_0, i_13_431_3889_0,
    i_13_431_3987_0, i_13_431_4077_0, i_13_431_4116_0, i_13_431_4159_0,
    i_13_431_4180_0, i_13_431_4186_0, i_13_431_4213_0, i_13_431_4248_0,
    i_13_431_4257_0, i_13_431_4320_0, i_13_431_4365_0, i_13_431_4366_0,
    i_13_431_4429_0, i_13_431_4521_0, i_13_431_4564_0, i_13_431_4566_0,
    i_13_431_4567_0, i_13_431_4590_0, i_13_431_4599_0, i_13_431_4600_0,
    o_13_431_0_0  );
  input  i_13_431_37_0, i_13_431_93_0, i_13_431_102_0, i_13_431_138_0,
    i_13_431_139_0, i_13_431_174_0, i_13_431_229_0, i_13_431_267_0,
    i_13_431_373_0, i_13_431_505_0, i_13_431_549_0, i_13_431_550_0,
    i_13_431_603_0, i_13_431_604_0, i_13_431_657_0, i_13_431_660_0,
    i_13_431_661_0, i_13_431_663_0, i_13_431_669_0, i_13_431_675_0,
    i_13_431_676_0, i_13_431_855_0, i_13_431_1023_0, i_13_431_1072_0,
    i_13_431_1144_0, i_13_431_1219_0, i_13_431_1494_0, i_13_431_1515_0,
    i_13_431_1516_0, i_13_431_1521_0, i_13_431_1629_0, i_13_431_1630_0,
    i_13_431_1656_0, i_13_431_1711_0, i_13_431_1827_0, i_13_431_1828_0,
    i_13_431_1858_0, i_13_431_1881_0, i_13_431_1884_0, i_13_431_2001_0,
    i_13_431_2002_0, i_13_431_2016_0, i_13_431_2019_0, i_13_431_2020_0,
    i_13_431_2169_0, i_13_431_2340_0, i_13_431_2341_0, i_13_431_2362_0,
    i_13_431_2397_0, i_13_431_2398_0, i_13_431_2422_0, i_13_431_2448_0,
    i_13_431_2467_0, i_13_431_2497_0, i_13_431_2511_0, i_13_431_2611_0,
    i_13_431_2614_0, i_13_431_2718_0, i_13_431_2935_0, i_13_431_2982_0,
    i_13_431_3006_0, i_13_431_3009_0, i_13_431_3105_0, i_13_431_3108_0,
    i_13_431_3133_0, i_13_431_3159_0, i_13_431_3234_0, i_13_431_3385_0,
    i_13_431_3415_0, i_13_431_3475_0, i_13_431_3522_0, i_13_431_3639_0,
    i_13_431_3640_0, i_13_431_3738_0, i_13_431_3762_0, i_13_431_3763_0,
    i_13_431_3843_0, i_13_431_3861_0, i_13_431_3862_0, i_13_431_3889_0,
    i_13_431_3987_0, i_13_431_4077_0, i_13_431_4116_0, i_13_431_4159_0,
    i_13_431_4180_0, i_13_431_4186_0, i_13_431_4213_0, i_13_431_4248_0,
    i_13_431_4257_0, i_13_431_4320_0, i_13_431_4365_0, i_13_431_4366_0,
    i_13_431_4429_0, i_13_431_4521_0, i_13_431_4564_0, i_13_431_4566_0,
    i_13_431_4567_0, i_13_431_4590_0, i_13_431_4599_0, i_13_431_4600_0;
  output o_13_431_0_0;
  assign o_13_431_0_0 = ~((i_13_431_139_0 & ((~i_13_431_1521_0 & ~i_13_431_3889_0) | (~i_13_431_4186_0 & ~i_13_431_4567_0))) | (~i_13_431_4365_0 & (i_13_431_1219_0 | (~i_13_431_675_0 & ~i_13_431_1144_0 & ~i_13_431_3762_0))) | (~i_13_431_2016_0 & ~i_13_431_2020_0 & ~i_13_431_3006_0) | (~i_13_431_3105_0 & ~i_13_431_4366_0) | (i_13_431_229_0 & ~i_13_431_3522_0 & ~i_13_431_4429_0));
endmodule



// Benchmark "kernel_13_432" written by ABC on Sun Jul 19 10:51:23 2020

module kernel_13_432 ( 
    i_13_432_49_0, i_13_432_75_0, i_13_432_76_0, i_13_432_94_0,
    i_13_432_133_0, i_13_432_139_0, i_13_432_183_0, i_13_432_187_0,
    i_13_432_192_0, i_13_432_193_0, i_13_432_195_0, i_13_432_207_0,
    i_13_432_321_0, i_13_432_526_0, i_13_432_542_0, i_13_432_570_0,
    i_13_432_574_0, i_13_432_612_0, i_13_432_663_0, i_13_432_668_0,
    i_13_432_697_0, i_13_432_714_0, i_13_432_798_0, i_13_432_831_0,
    i_13_432_847_0, i_13_432_853_0, i_13_432_854_0, i_13_432_985_0,
    i_13_432_988_0, i_13_432_1069_0, i_13_432_1149_0, i_13_432_1222_0,
    i_13_432_1230_0, i_13_432_1231_0, i_13_432_1321_0, i_13_432_1407_0,
    i_13_432_1408_0, i_13_432_1410_0, i_13_432_1521_0, i_13_432_1537_0,
    i_13_432_1548_0, i_13_432_1678_0, i_13_432_1732_0, i_13_432_1771_0,
    i_13_432_1804_0, i_13_432_1827_0, i_13_432_1834_0, i_13_432_1857_0,
    i_13_432_1860_0, i_13_432_1861_0, i_13_432_1885_0, i_13_432_2002_0,
    i_13_432_2100_0, i_13_432_2142_0, i_13_432_2145_0, i_13_432_2203_0,
    i_13_432_2299_0, i_13_432_2402_0, i_13_432_2422_0, i_13_432_2473_0,
    i_13_432_2680_0, i_13_432_2856_0, i_13_432_2857_0, i_13_432_2982_0,
    i_13_432_3000_0, i_13_432_3009_0, i_13_432_3064_0, i_13_432_3112_0,
    i_13_432_3159_0, i_13_432_3207_0, i_13_432_3208_0, i_13_432_3210_0,
    i_13_432_3212_0, i_13_432_3244_0, i_13_432_3409_0, i_13_432_3439_0,
    i_13_432_3442_0, i_13_432_3487_0, i_13_432_3531_0, i_13_432_3558_0,
    i_13_432_3667_0, i_13_432_3685_0, i_13_432_3730_0, i_13_432_3756_0,
    i_13_432_3763_0, i_13_432_3765_0, i_13_432_3979_0, i_13_432_3982_0,
    i_13_432_3984_0, i_13_432_4084_0, i_13_432_4357_0, i_13_432_4396_0,
    i_13_432_4432_0, i_13_432_4504_0, i_13_432_4512_0, i_13_432_4565_0,
    i_13_432_4566_0, i_13_432_4567_0, i_13_432_4569_0, i_13_432_4587_0,
    o_13_432_0_0  );
  input  i_13_432_49_0, i_13_432_75_0, i_13_432_76_0, i_13_432_94_0,
    i_13_432_133_0, i_13_432_139_0, i_13_432_183_0, i_13_432_187_0,
    i_13_432_192_0, i_13_432_193_0, i_13_432_195_0, i_13_432_207_0,
    i_13_432_321_0, i_13_432_526_0, i_13_432_542_0, i_13_432_570_0,
    i_13_432_574_0, i_13_432_612_0, i_13_432_663_0, i_13_432_668_0,
    i_13_432_697_0, i_13_432_714_0, i_13_432_798_0, i_13_432_831_0,
    i_13_432_847_0, i_13_432_853_0, i_13_432_854_0, i_13_432_985_0,
    i_13_432_988_0, i_13_432_1069_0, i_13_432_1149_0, i_13_432_1222_0,
    i_13_432_1230_0, i_13_432_1231_0, i_13_432_1321_0, i_13_432_1407_0,
    i_13_432_1408_0, i_13_432_1410_0, i_13_432_1521_0, i_13_432_1537_0,
    i_13_432_1548_0, i_13_432_1678_0, i_13_432_1732_0, i_13_432_1771_0,
    i_13_432_1804_0, i_13_432_1827_0, i_13_432_1834_0, i_13_432_1857_0,
    i_13_432_1860_0, i_13_432_1861_0, i_13_432_1885_0, i_13_432_2002_0,
    i_13_432_2100_0, i_13_432_2142_0, i_13_432_2145_0, i_13_432_2203_0,
    i_13_432_2299_0, i_13_432_2402_0, i_13_432_2422_0, i_13_432_2473_0,
    i_13_432_2680_0, i_13_432_2856_0, i_13_432_2857_0, i_13_432_2982_0,
    i_13_432_3000_0, i_13_432_3009_0, i_13_432_3064_0, i_13_432_3112_0,
    i_13_432_3159_0, i_13_432_3207_0, i_13_432_3208_0, i_13_432_3210_0,
    i_13_432_3212_0, i_13_432_3244_0, i_13_432_3409_0, i_13_432_3439_0,
    i_13_432_3442_0, i_13_432_3487_0, i_13_432_3531_0, i_13_432_3558_0,
    i_13_432_3667_0, i_13_432_3685_0, i_13_432_3730_0, i_13_432_3756_0,
    i_13_432_3763_0, i_13_432_3765_0, i_13_432_3979_0, i_13_432_3982_0,
    i_13_432_3984_0, i_13_432_4084_0, i_13_432_4357_0, i_13_432_4396_0,
    i_13_432_4432_0, i_13_432_4504_0, i_13_432_4512_0, i_13_432_4565_0,
    i_13_432_4566_0, i_13_432_4567_0, i_13_432_4569_0, i_13_432_4587_0;
  output o_13_432_0_0;
  assign o_13_432_0_0 = ~((~i_13_432_4569_0 & (~i_13_432_1408_0 | (i_13_432_2002_0 & ~i_13_432_3009_0))) | (i_13_432_2002_0 & (~i_13_432_2982_0 | (~i_13_432_2422_0 & ~i_13_432_3984_0))) | ~i_13_432_1407_0 | (~i_13_432_570_0 & ~i_13_432_1804_0) | (~i_13_432_2145_0 & i_13_432_3763_0) | (~i_13_432_3210_0 & ~i_13_432_3765_0) | (i_13_432_4432_0 & ~i_13_432_4512_0));
endmodule



// Benchmark "kernel_13_433" written by ABC on Sun Jul 19 10:51:24 2020

module kernel_13_433 ( 
    i_13_433_18_0, i_13_433_36_0, i_13_433_90_0, i_13_433_94_0,
    i_13_433_139_0, i_13_433_407_0, i_13_433_446_0, i_13_433_572_0,
    i_13_433_580_0, i_13_433_697_0, i_13_433_732_0, i_13_433_737_0,
    i_13_433_796_0, i_13_433_797_0, i_13_433_799_0, i_13_433_800_0,
    i_13_433_838_0, i_13_433_844_0, i_13_433_855_0, i_13_433_862_0,
    i_13_433_949_0, i_13_433_950_0, i_13_433_979_0, i_13_433_1030_0,
    i_13_433_1120_0, i_13_433_1196_0, i_13_433_1227_0, i_13_433_1303_0,
    i_13_433_1427_0, i_13_433_1445_0, i_13_433_1489_0, i_13_433_1492_0,
    i_13_433_1498_0, i_13_433_1499_0, i_13_433_1633_0, i_13_433_1732_0,
    i_13_433_1792_0, i_13_433_1854_0, i_13_433_1867_0, i_13_433_1996_0,
    i_13_433_2003_0, i_13_433_2005_0, i_13_433_2056_0, i_13_433_2208_0,
    i_13_433_2209_0, i_13_433_2272_0, i_13_433_2321_0, i_13_433_2357_0,
    i_13_433_2365_0, i_13_433_2425_0, i_13_433_2428_0, i_13_433_2434_0,
    i_13_433_2436_0, i_13_433_2437_0, i_13_433_2446_0, i_13_433_2461_0,
    i_13_433_2464_0, i_13_433_2465_0, i_13_433_2542_0, i_13_433_2544_0,
    i_13_433_2551_0, i_13_433_2614_0, i_13_433_2740_0, i_13_433_2749_0,
    i_13_433_2758_0, i_13_433_2919_0, i_13_433_2963_0, i_13_433_3001_0,
    i_13_433_3051_0, i_13_433_3059_0, i_13_433_3148_0, i_13_433_3163_0,
    i_13_433_3289_0, i_13_433_3424_0, i_13_433_3425_0, i_13_433_3476_0,
    i_13_433_3523_0, i_13_433_3531_0, i_13_433_3532_0, i_13_433_3535_0,
    i_13_433_3617_0, i_13_433_3726_0, i_13_433_3730_0, i_13_433_3733_0,
    i_13_433_3871_0, i_13_433_3873_0, i_13_433_3874_0, i_13_433_3877_0,
    i_13_433_3906_0, i_13_433_3910_0, i_13_433_4006_0, i_13_433_4036_0,
    i_13_433_4155_0, i_13_433_4189_0, i_13_433_4202_0, i_13_433_4236_0,
    i_13_433_4254_0, i_13_433_4450_0, i_13_433_4561_0, i_13_433_4603_0,
    o_13_433_0_0  );
  input  i_13_433_18_0, i_13_433_36_0, i_13_433_90_0, i_13_433_94_0,
    i_13_433_139_0, i_13_433_407_0, i_13_433_446_0, i_13_433_572_0,
    i_13_433_580_0, i_13_433_697_0, i_13_433_732_0, i_13_433_737_0,
    i_13_433_796_0, i_13_433_797_0, i_13_433_799_0, i_13_433_800_0,
    i_13_433_838_0, i_13_433_844_0, i_13_433_855_0, i_13_433_862_0,
    i_13_433_949_0, i_13_433_950_0, i_13_433_979_0, i_13_433_1030_0,
    i_13_433_1120_0, i_13_433_1196_0, i_13_433_1227_0, i_13_433_1303_0,
    i_13_433_1427_0, i_13_433_1445_0, i_13_433_1489_0, i_13_433_1492_0,
    i_13_433_1498_0, i_13_433_1499_0, i_13_433_1633_0, i_13_433_1732_0,
    i_13_433_1792_0, i_13_433_1854_0, i_13_433_1867_0, i_13_433_1996_0,
    i_13_433_2003_0, i_13_433_2005_0, i_13_433_2056_0, i_13_433_2208_0,
    i_13_433_2209_0, i_13_433_2272_0, i_13_433_2321_0, i_13_433_2357_0,
    i_13_433_2365_0, i_13_433_2425_0, i_13_433_2428_0, i_13_433_2434_0,
    i_13_433_2436_0, i_13_433_2437_0, i_13_433_2446_0, i_13_433_2461_0,
    i_13_433_2464_0, i_13_433_2465_0, i_13_433_2542_0, i_13_433_2544_0,
    i_13_433_2551_0, i_13_433_2614_0, i_13_433_2740_0, i_13_433_2749_0,
    i_13_433_2758_0, i_13_433_2919_0, i_13_433_2963_0, i_13_433_3001_0,
    i_13_433_3051_0, i_13_433_3059_0, i_13_433_3148_0, i_13_433_3163_0,
    i_13_433_3289_0, i_13_433_3424_0, i_13_433_3425_0, i_13_433_3476_0,
    i_13_433_3523_0, i_13_433_3531_0, i_13_433_3532_0, i_13_433_3535_0,
    i_13_433_3617_0, i_13_433_3726_0, i_13_433_3730_0, i_13_433_3733_0,
    i_13_433_3871_0, i_13_433_3873_0, i_13_433_3874_0, i_13_433_3877_0,
    i_13_433_3906_0, i_13_433_3910_0, i_13_433_4006_0, i_13_433_4036_0,
    i_13_433_4155_0, i_13_433_4189_0, i_13_433_4202_0, i_13_433_4236_0,
    i_13_433_4254_0, i_13_433_4450_0, i_13_433_4561_0, i_13_433_4603_0;
  output o_13_433_0_0;
  assign o_13_433_0_0 = ~((~i_13_433_3871_0 & ((~i_13_433_2437_0 & ((~i_13_433_1792_0 & ~i_13_433_3730_0) | (~i_13_433_732_0 & ~i_13_433_3535_0 & ~i_13_433_3906_0))) | (~i_13_433_90_0 & ~i_13_433_1498_0 & ~i_13_433_3874_0))) | (~i_13_433_2919_0 & ((i_13_433_2209_0 & ~i_13_433_3874_0) | (i_13_433_90_0 & i_13_433_3906_0))) | (~i_13_433_3531_0 & ((~i_13_433_2464_0 & ~i_13_433_2544_0 & ~i_13_433_3874_0) | (i_13_433_2056_0 & ~i_13_433_4155_0))) | (~i_13_433_2208_0 & ~i_13_433_2425_0 & ~i_13_433_2542_0) | (~i_13_433_1854_0 & ~i_13_433_1996_0 & ~i_13_433_3148_0 & ~i_13_433_3424_0) | (~i_13_433_3535_0 & i_13_433_4189_0));
endmodule



// Benchmark "kernel_13_434" written by ABC on Sun Jul 19 10:51:25 2020

module kernel_13_434 ( 
    i_13_434_94_0, i_13_434_141_0, i_13_434_142_0, i_13_434_168_0,
    i_13_434_240_0, i_13_434_258_0, i_13_434_264_0, i_13_434_310_0,
    i_13_434_322_0, i_13_434_339_0, i_13_434_340_0, i_13_434_373_0,
    i_13_434_430_0, i_13_434_526_0, i_13_434_553_0, i_13_434_582_0,
    i_13_434_598_0, i_13_434_607_0, i_13_434_618_0, i_13_434_619_0,
    i_13_434_717_0, i_13_434_727_0, i_13_434_780_0, i_13_434_799_0,
    i_13_434_979_0, i_13_434_1077_0, i_13_434_1078_0, i_13_434_1231_0,
    i_13_434_1276_0, i_13_434_1311_0, i_13_434_1402_0, i_13_434_1435_0,
    i_13_434_1470_0, i_13_434_1471_0, i_13_434_1483_0, i_13_434_1597_0,
    i_13_434_1626_0, i_13_434_1635_0, i_13_434_1650_0, i_13_434_1699_0,
    i_13_434_1725_0, i_13_434_1734_0, i_13_434_1776_0, i_13_434_1780_0,
    i_13_434_1783_0, i_13_434_1785_0, i_13_434_1816_0, i_13_434_1849_0,
    i_13_434_1960_0, i_13_434_1996_0, i_13_434_2059_0, i_13_434_2149_0,
    i_13_434_2293_0, i_13_434_2319_0, i_13_434_2347_0, i_13_434_2434_0,
    i_13_434_2649_0, i_13_434_2679_0, i_13_434_2742_0, i_13_434_2751_0,
    i_13_434_2787_0, i_13_434_2859_0, i_13_434_2886_0, i_13_434_2937_0,
    i_13_434_3013_0, i_13_434_3039_0, i_13_434_3291_0, i_13_434_3292_0,
    i_13_434_3414_0, i_13_434_3415_0, i_13_434_3444_0, i_13_434_3481_0,
    i_13_434_3525_0, i_13_434_3526_0, i_13_434_3532_0, i_13_434_3534_0,
    i_13_434_3541_0, i_13_434_3550_0, i_13_434_3642_0, i_13_434_3643_0,
    i_13_434_3687_0, i_13_434_3688_0, i_13_434_3706_0, i_13_434_3756_0,
    i_13_434_3757_0, i_13_434_4278_0, i_13_434_4318_0, i_13_434_4327_0,
    i_13_434_4335_0, i_13_434_4354_0, i_13_434_4360_0, i_13_434_4363_0,
    i_13_434_4389_0, i_13_434_4390_0, i_13_434_4395_0, i_13_434_4417_0,
    i_13_434_4432_0, i_13_434_4513_0, i_13_434_4525_0, i_13_434_4533_0,
    o_13_434_0_0  );
  input  i_13_434_94_0, i_13_434_141_0, i_13_434_142_0, i_13_434_168_0,
    i_13_434_240_0, i_13_434_258_0, i_13_434_264_0, i_13_434_310_0,
    i_13_434_322_0, i_13_434_339_0, i_13_434_340_0, i_13_434_373_0,
    i_13_434_430_0, i_13_434_526_0, i_13_434_553_0, i_13_434_582_0,
    i_13_434_598_0, i_13_434_607_0, i_13_434_618_0, i_13_434_619_0,
    i_13_434_717_0, i_13_434_727_0, i_13_434_780_0, i_13_434_799_0,
    i_13_434_979_0, i_13_434_1077_0, i_13_434_1078_0, i_13_434_1231_0,
    i_13_434_1276_0, i_13_434_1311_0, i_13_434_1402_0, i_13_434_1435_0,
    i_13_434_1470_0, i_13_434_1471_0, i_13_434_1483_0, i_13_434_1597_0,
    i_13_434_1626_0, i_13_434_1635_0, i_13_434_1650_0, i_13_434_1699_0,
    i_13_434_1725_0, i_13_434_1734_0, i_13_434_1776_0, i_13_434_1780_0,
    i_13_434_1783_0, i_13_434_1785_0, i_13_434_1816_0, i_13_434_1849_0,
    i_13_434_1960_0, i_13_434_1996_0, i_13_434_2059_0, i_13_434_2149_0,
    i_13_434_2293_0, i_13_434_2319_0, i_13_434_2347_0, i_13_434_2434_0,
    i_13_434_2649_0, i_13_434_2679_0, i_13_434_2742_0, i_13_434_2751_0,
    i_13_434_2787_0, i_13_434_2859_0, i_13_434_2886_0, i_13_434_2937_0,
    i_13_434_3013_0, i_13_434_3039_0, i_13_434_3291_0, i_13_434_3292_0,
    i_13_434_3414_0, i_13_434_3415_0, i_13_434_3444_0, i_13_434_3481_0,
    i_13_434_3525_0, i_13_434_3526_0, i_13_434_3532_0, i_13_434_3534_0,
    i_13_434_3541_0, i_13_434_3550_0, i_13_434_3642_0, i_13_434_3643_0,
    i_13_434_3687_0, i_13_434_3688_0, i_13_434_3706_0, i_13_434_3756_0,
    i_13_434_3757_0, i_13_434_4278_0, i_13_434_4318_0, i_13_434_4327_0,
    i_13_434_4335_0, i_13_434_4354_0, i_13_434_4360_0, i_13_434_4363_0,
    i_13_434_4389_0, i_13_434_4390_0, i_13_434_4395_0, i_13_434_4417_0,
    i_13_434_4432_0, i_13_434_4513_0, i_13_434_4525_0, i_13_434_4533_0;
  output o_13_434_0_0;
  assign o_13_434_0_0 = ~(~i_13_434_618_0 | ~i_13_434_1734_0);
endmodule



// Benchmark "kernel_13_435" written by ABC on Sun Jul 19 10:51:25 2020

module kernel_13_435 ( 
    i_13_435_34_0, i_13_435_67_0, i_13_435_71_0, i_13_435_95_0,
    i_13_435_136_0, i_13_435_137_0, i_13_435_185_0, i_13_435_200_0,
    i_13_435_448_0, i_13_435_449_0, i_13_435_517_0, i_13_435_535_0,
    i_13_435_536_0, i_13_435_538_0, i_13_435_605_0, i_13_435_613_0,
    i_13_435_614_0, i_13_435_644_0, i_13_435_682_0, i_13_435_686_0,
    i_13_435_703_0, i_13_435_934_0, i_13_435_1077_0, i_13_435_1087_0,
    i_13_435_1105_0, i_13_435_1123_0, i_13_435_1196_0, i_13_435_1215_0,
    i_13_435_1216_0, i_13_435_1218_0, i_13_435_1232_0, i_13_435_1274_0,
    i_13_435_1276_0, i_13_435_1283_0, i_13_435_1402_0, i_13_435_1403_0,
    i_13_435_1441_0, i_13_435_1598_0, i_13_435_1606_0, i_13_435_1643_0,
    i_13_435_1674_0, i_13_435_1736_0, i_13_435_1767_0, i_13_435_1796_0,
    i_13_435_1798_0, i_13_435_1799_0, i_13_435_1858_0, i_13_435_1889_0,
    i_13_435_1931_0, i_13_435_1934_0, i_13_435_1945_0, i_13_435_1998_0,
    i_13_435_2075_0, i_13_435_2123_0, i_13_435_2174_0, i_13_435_2176_0,
    i_13_435_2267_0, i_13_435_2421_0, i_13_435_2422_0, i_13_435_2425_0,
    i_13_435_2426_0, i_13_435_2567_0, i_13_435_2648_0, i_13_435_2917_0,
    i_13_435_3031_0, i_13_435_3032_0, i_13_435_3064_0, i_13_435_3103_0,
    i_13_435_3104_0, i_13_435_3128_0, i_13_435_3130_0, i_13_435_3212_0,
    i_13_435_3216_0, i_13_435_3239_0, i_13_435_3265_0, i_13_435_3367_0,
    i_13_435_3368_0, i_13_435_3406_0, i_13_435_3418_0, i_13_435_3419_0,
    i_13_435_3439_0, i_13_435_3456_0, i_13_435_3638_0, i_13_435_3699_0,
    i_13_435_3745_0, i_13_435_3787_0, i_13_435_3876_0, i_13_435_3899_0,
    i_13_435_3931_0, i_13_435_3932_0, i_13_435_3994_0, i_13_435_3995_0,
    i_13_435_4015_0, i_13_435_4042_0, i_13_435_4046_0, i_13_435_4066_0,
    i_13_435_4084_0, i_13_435_4085_0, i_13_435_4297_0, i_13_435_4606_0,
    o_13_435_0_0  );
  input  i_13_435_34_0, i_13_435_67_0, i_13_435_71_0, i_13_435_95_0,
    i_13_435_136_0, i_13_435_137_0, i_13_435_185_0, i_13_435_200_0,
    i_13_435_448_0, i_13_435_449_0, i_13_435_517_0, i_13_435_535_0,
    i_13_435_536_0, i_13_435_538_0, i_13_435_605_0, i_13_435_613_0,
    i_13_435_614_0, i_13_435_644_0, i_13_435_682_0, i_13_435_686_0,
    i_13_435_703_0, i_13_435_934_0, i_13_435_1077_0, i_13_435_1087_0,
    i_13_435_1105_0, i_13_435_1123_0, i_13_435_1196_0, i_13_435_1215_0,
    i_13_435_1216_0, i_13_435_1218_0, i_13_435_1232_0, i_13_435_1274_0,
    i_13_435_1276_0, i_13_435_1283_0, i_13_435_1402_0, i_13_435_1403_0,
    i_13_435_1441_0, i_13_435_1598_0, i_13_435_1606_0, i_13_435_1643_0,
    i_13_435_1674_0, i_13_435_1736_0, i_13_435_1767_0, i_13_435_1796_0,
    i_13_435_1798_0, i_13_435_1799_0, i_13_435_1858_0, i_13_435_1889_0,
    i_13_435_1931_0, i_13_435_1934_0, i_13_435_1945_0, i_13_435_1998_0,
    i_13_435_2075_0, i_13_435_2123_0, i_13_435_2174_0, i_13_435_2176_0,
    i_13_435_2267_0, i_13_435_2421_0, i_13_435_2422_0, i_13_435_2425_0,
    i_13_435_2426_0, i_13_435_2567_0, i_13_435_2648_0, i_13_435_2917_0,
    i_13_435_3031_0, i_13_435_3032_0, i_13_435_3064_0, i_13_435_3103_0,
    i_13_435_3104_0, i_13_435_3128_0, i_13_435_3130_0, i_13_435_3212_0,
    i_13_435_3216_0, i_13_435_3239_0, i_13_435_3265_0, i_13_435_3367_0,
    i_13_435_3368_0, i_13_435_3406_0, i_13_435_3418_0, i_13_435_3419_0,
    i_13_435_3439_0, i_13_435_3456_0, i_13_435_3638_0, i_13_435_3699_0,
    i_13_435_3745_0, i_13_435_3787_0, i_13_435_3876_0, i_13_435_3899_0,
    i_13_435_3931_0, i_13_435_3932_0, i_13_435_3994_0, i_13_435_3995_0,
    i_13_435_4015_0, i_13_435_4042_0, i_13_435_4046_0, i_13_435_4066_0,
    i_13_435_4084_0, i_13_435_4085_0, i_13_435_4297_0, i_13_435_4606_0;
  output o_13_435_0_0;
  assign o_13_435_0_0 = ~(~i_13_435_4085_0 | (~i_13_435_682_0 & (~i_13_435_1087_0 | ~i_13_435_3932_0)));
endmodule



// Benchmark "kernel_13_436" written by ABC on Sun Jul 19 10:51:26 2020

module kernel_13_436 ( 
    i_13_436_47_0, i_13_436_73_0, i_13_436_74_0, i_13_436_157_0,
    i_13_436_166_0, i_13_436_184_0, i_13_436_229_0, i_13_436_342_0,
    i_13_436_357_0, i_13_436_362_0, i_13_436_428_0, i_13_436_431_0,
    i_13_436_434_0, i_13_436_513_0, i_13_436_515_0, i_13_436_533_0,
    i_13_436_551_0, i_13_436_605_0, i_13_436_607_0, i_13_436_649_0,
    i_13_436_652_0, i_13_436_653_0, i_13_436_659_0, i_13_436_667_0,
    i_13_436_694_0, i_13_436_698_0, i_13_436_841_0, i_13_436_886_0,
    i_13_436_1110_0, i_13_436_1117_0, i_13_436_1144_0, i_13_436_1145_0,
    i_13_436_1207_0, i_13_436_1208_0, i_13_436_1658_0, i_13_436_1732_0,
    i_13_436_1742_0, i_13_436_1791_0, i_13_436_1792_0, i_13_436_1918_0,
    i_13_436_1920_0, i_13_436_1939_0, i_13_436_1950_0, i_13_436_1951_0,
    i_13_436_2017_0, i_13_436_2020_0, i_13_436_2030_0, i_13_436_2206_0,
    i_13_436_2209_0, i_13_436_2318_0, i_13_436_2377_0, i_13_436_2443_0,
    i_13_436_2452_0, i_13_436_2467_0, i_13_436_2514_0, i_13_436_2691_0,
    i_13_436_2785_0, i_13_436_2884_0, i_13_436_2906_0, i_13_436_2938_0,
    i_13_436_2939_0, i_13_436_2956_0, i_13_436_2958_0, i_13_436_3044_0,
    i_13_436_3101_0, i_13_436_3153_0, i_13_436_3241_0, i_13_436_3312_0,
    i_13_436_3313_0, i_13_436_3367_0, i_13_436_3476_0, i_13_436_3479_0,
    i_13_436_3488_0, i_13_436_3532_0, i_13_436_3550_0, i_13_436_3568_0,
    i_13_436_3569_0, i_13_436_3596_0, i_13_436_3598_0, i_13_436_3646_0,
    i_13_436_3739_0, i_13_436_3866_0, i_13_436_3910_0, i_13_436_4063_0,
    i_13_436_4158_0, i_13_436_4177_0, i_13_436_4186_0, i_13_436_4187_0,
    i_13_436_4190_0, i_13_436_4199_0, i_13_436_4257_0, i_13_436_4297_0,
    i_13_436_4306_0, i_13_436_4330_0, i_13_436_4331_0, i_13_436_4333_0,
    i_13_436_4448_0, i_13_436_4522_0, i_13_436_4540_0, i_13_436_4601_0,
    o_13_436_0_0  );
  input  i_13_436_47_0, i_13_436_73_0, i_13_436_74_0, i_13_436_157_0,
    i_13_436_166_0, i_13_436_184_0, i_13_436_229_0, i_13_436_342_0,
    i_13_436_357_0, i_13_436_362_0, i_13_436_428_0, i_13_436_431_0,
    i_13_436_434_0, i_13_436_513_0, i_13_436_515_0, i_13_436_533_0,
    i_13_436_551_0, i_13_436_605_0, i_13_436_607_0, i_13_436_649_0,
    i_13_436_652_0, i_13_436_653_0, i_13_436_659_0, i_13_436_667_0,
    i_13_436_694_0, i_13_436_698_0, i_13_436_841_0, i_13_436_886_0,
    i_13_436_1110_0, i_13_436_1117_0, i_13_436_1144_0, i_13_436_1145_0,
    i_13_436_1207_0, i_13_436_1208_0, i_13_436_1658_0, i_13_436_1732_0,
    i_13_436_1742_0, i_13_436_1791_0, i_13_436_1792_0, i_13_436_1918_0,
    i_13_436_1920_0, i_13_436_1939_0, i_13_436_1950_0, i_13_436_1951_0,
    i_13_436_2017_0, i_13_436_2020_0, i_13_436_2030_0, i_13_436_2206_0,
    i_13_436_2209_0, i_13_436_2318_0, i_13_436_2377_0, i_13_436_2443_0,
    i_13_436_2452_0, i_13_436_2467_0, i_13_436_2514_0, i_13_436_2691_0,
    i_13_436_2785_0, i_13_436_2884_0, i_13_436_2906_0, i_13_436_2938_0,
    i_13_436_2939_0, i_13_436_2956_0, i_13_436_2958_0, i_13_436_3044_0,
    i_13_436_3101_0, i_13_436_3153_0, i_13_436_3241_0, i_13_436_3312_0,
    i_13_436_3313_0, i_13_436_3367_0, i_13_436_3476_0, i_13_436_3479_0,
    i_13_436_3488_0, i_13_436_3532_0, i_13_436_3550_0, i_13_436_3568_0,
    i_13_436_3569_0, i_13_436_3596_0, i_13_436_3598_0, i_13_436_3646_0,
    i_13_436_3739_0, i_13_436_3866_0, i_13_436_3910_0, i_13_436_4063_0,
    i_13_436_4158_0, i_13_436_4177_0, i_13_436_4186_0, i_13_436_4187_0,
    i_13_436_4190_0, i_13_436_4199_0, i_13_436_4257_0, i_13_436_4297_0,
    i_13_436_4306_0, i_13_436_4330_0, i_13_436_4331_0, i_13_436_4333_0,
    i_13_436_4448_0, i_13_436_4522_0, i_13_436_4540_0, i_13_436_4601_0;
  output o_13_436_0_0;
  assign o_13_436_0_0 = ~((~i_13_436_2017_0 & (~i_13_436_4448_0 | (~i_13_436_694_0 & ~i_13_436_4333_0))) | ~i_13_436_2884_0 | (~i_13_436_1144_0 & i_13_436_3550_0) | (~i_13_436_47_0 & ~i_13_436_649_0 & ~i_13_436_4190_0 & ~i_13_436_4330_0));
endmodule



// Benchmark "kernel_13_437" written by ABC on Sun Jul 19 10:51:27 2020

module kernel_13_437 ( 
    i_13_437_47_0, i_13_437_65_0, i_13_437_109_0, i_13_437_110_0,
    i_13_437_111_0, i_13_437_112_0, i_13_437_206_0, i_13_437_276_0,
    i_13_437_382_0, i_13_437_411_0, i_13_437_520_0, i_13_437_605_0,
    i_13_437_626_0, i_13_437_659_0, i_13_437_680_0, i_13_437_816_0,
    i_13_437_856_0, i_13_437_927_0, i_13_437_932_0, i_13_437_937_0,
    i_13_437_938_0, i_13_437_1054_0, i_13_437_1072_0, i_13_437_1077_0,
    i_13_437_1086_0, i_13_437_1096_0, i_13_437_1212_0, i_13_437_1316_0,
    i_13_437_1424_0, i_13_437_1481_0, i_13_437_1495_0, i_13_437_1498_0,
    i_13_437_1519_0, i_13_437_1626_0, i_13_437_1653_0, i_13_437_1662_0,
    i_13_437_1735_0, i_13_437_1742_0, i_13_437_1746_0, i_13_437_1747_0,
    i_13_437_2020_0, i_13_437_2023_0, i_13_437_2136_0, i_13_437_2191_0,
    i_13_437_2248_0, i_13_437_2263_0, i_13_437_2320_0, i_13_437_2407_0,
    i_13_437_2481_0, i_13_437_2500_0, i_13_437_2529_0, i_13_437_2539_0,
    i_13_437_2562_0, i_13_437_2595_0, i_13_437_2677_0, i_13_437_2723_0,
    i_13_437_2884_0, i_13_437_2913_0, i_13_437_2935_0, i_13_437_3047_0,
    i_13_437_3089_0, i_13_437_3095_0, i_13_437_3100_0, i_13_437_3102_0,
    i_13_437_3103_0, i_13_437_3315_0, i_13_437_3326_0, i_13_437_3339_0,
    i_13_437_3355_0, i_13_437_3451_0, i_13_437_3452_0, i_13_437_3478_0,
    i_13_437_3550_0, i_13_437_3564_0, i_13_437_3570_0, i_13_437_3602_0,
    i_13_437_3606_0, i_13_437_3661_0, i_13_437_3685_0, i_13_437_3688_0,
    i_13_437_3730_0, i_13_437_3741_0, i_13_437_3859_0, i_13_437_4119_0,
    i_13_437_4159_0, i_13_437_4160_0, i_13_437_4162_0, i_13_437_4165_0,
    i_13_437_4173_0, i_13_437_4181_0, i_13_437_4184_0, i_13_437_4325_0,
    i_13_437_4332_0, i_13_437_4334_0, i_13_437_4335_0, i_13_437_4365_0,
    i_13_437_4366_0, i_13_437_4370_0, i_13_437_4372_0, i_13_437_4544_0,
    o_13_437_0_0  );
  input  i_13_437_47_0, i_13_437_65_0, i_13_437_109_0, i_13_437_110_0,
    i_13_437_111_0, i_13_437_112_0, i_13_437_206_0, i_13_437_276_0,
    i_13_437_382_0, i_13_437_411_0, i_13_437_520_0, i_13_437_605_0,
    i_13_437_626_0, i_13_437_659_0, i_13_437_680_0, i_13_437_816_0,
    i_13_437_856_0, i_13_437_927_0, i_13_437_932_0, i_13_437_937_0,
    i_13_437_938_0, i_13_437_1054_0, i_13_437_1072_0, i_13_437_1077_0,
    i_13_437_1086_0, i_13_437_1096_0, i_13_437_1212_0, i_13_437_1316_0,
    i_13_437_1424_0, i_13_437_1481_0, i_13_437_1495_0, i_13_437_1498_0,
    i_13_437_1519_0, i_13_437_1626_0, i_13_437_1653_0, i_13_437_1662_0,
    i_13_437_1735_0, i_13_437_1742_0, i_13_437_1746_0, i_13_437_1747_0,
    i_13_437_2020_0, i_13_437_2023_0, i_13_437_2136_0, i_13_437_2191_0,
    i_13_437_2248_0, i_13_437_2263_0, i_13_437_2320_0, i_13_437_2407_0,
    i_13_437_2481_0, i_13_437_2500_0, i_13_437_2529_0, i_13_437_2539_0,
    i_13_437_2562_0, i_13_437_2595_0, i_13_437_2677_0, i_13_437_2723_0,
    i_13_437_2884_0, i_13_437_2913_0, i_13_437_2935_0, i_13_437_3047_0,
    i_13_437_3089_0, i_13_437_3095_0, i_13_437_3100_0, i_13_437_3102_0,
    i_13_437_3103_0, i_13_437_3315_0, i_13_437_3326_0, i_13_437_3339_0,
    i_13_437_3355_0, i_13_437_3451_0, i_13_437_3452_0, i_13_437_3478_0,
    i_13_437_3550_0, i_13_437_3564_0, i_13_437_3570_0, i_13_437_3602_0,
    i_13_437_3606_0, i_13_437_3661_0, i_13_437_3685_0, i_13_437_3688_0,
    i_13_437_3730_0, i_13_437_3741_0, i_13_437_3859_0, i_13_437_4119_0,
    i_13_437_4159_0, i_13_437_4160_0, i_13_437_4162_0, i_13_437_4165_0,
    i_13_437_4173_0, i_13_437_4181_0, i_13_437_4184_0, i_13_437_4325_0,
    i_13_437_4332_0, i_13_437_4334_0, i_13_437_4335_0, i_13_437_4365_0,
    i_13_437_4366_0, i_13_437_4370_0, i_13_437_4372_0, i_13_437_4544_0;
  output o_13_437_0_0;
  assign o_13_437_0_0 = ~((~i_13_437_4160_0 & ((~i_13_437_927_0 & ~i_13_437_937_0 & ~i_13_437_1086_0 & ~i_13_437_1626_0 & ~i_13_437_2023_0) | (~i_13_437_3100_0 & ~i_13_437_3103_0 & ~i_13_437_4335_0))) | i_13_437_2935_0 | i_13_437_3339_0 | (~i_13_437_112_0 & ~i_13_437_3741_0 & i_13_437_3859_0) | (i_13_437_382_0 & ~i_13_437_2884_0 & ~i_13_437_4159_0) | (~i_13_437_110_0 & ~i_13_437_111_0 & ~i_13_437_4334_0 & ~i_13_437_4335_0));
endmodule



// Benchmark "kernel_13_438" written by ABC on Sun Jul 19 10:51:28 2020

module kernel_13_438 ( 
    i_13_438_29_0, i_13_438_45_0, i_13_438_107_0, i_13_438_271_0,
    i_13_438_300_0, i_13_438_352_0, i_13_438_374_0, i_13_438_422_0,
    i_13_438_451_0, i_13_438_559_0, i_13_438_561_0, i_13_438_562_0,
    i_13_438_569_0, i_13_438_604_0, i_13_438_605_0, i_13_438_607_0,
    i_13_438_608_0, i_13_438_610_0, i_13_438_658_0, i_13_438_659_0,
    i_13_438_661_0, i_13_438_662_0, i_13_438_670_0, i_13_438_680_0,
    i_13_438_829_0, i_13_438_832_0, i_13_438_833_0, i_13_438_882_0,
    i_13_438_885_0, i_13_438_886_0, i_13_438_946_0, i_13_438_1075_0,
    i_13_438_1084_0, i_13_438_1226_0, i_13_438_1281_0, i_13_438_1381_0,
    i_13_438_1404_0, i_13_438_1405_0, i_13_438_1467_0, i_13_438_1520_0,
    i_13_438_1522_0, i_13_438_1535_0, i_13_438_1660_0, i_13_438_1768_0,
    i_13_438_1787_0, i_13_438_1802_0, i_13_438_1838_0, i_13_438_1846_0,
    i_13_438_1885_0, i_13_438_1897_0, i_13_438_1927_0, i_13_438_2021_0,
    i_13_438_2137_0, i_13_438_2170_0, i_13_438_2297_0, i_13_438_2423_0,
    i_13_438_2431_0, i_13_438_2435_0, i_13_438_2647_0, i_13_438_2650_0,
    i_13_438_2749_0, i_13_438_2880_0, i_13_438_3047_0, i_13_438_3106_0,
    i_13_438_3117_0, i_13_438_3311_0, i_13_438_3457_0, i_13_438_3476_0,
    i_13_438_3547_0, i_13_438_3638_0, i_13_438_3664_0, i_13_438_3683_0,
    i_13_438_3740_0, i_13_438_3844_0, i_13_438_3871_0, i_13_438_3872_0,
    i_13_438_3889_0, i_13_438_3910_0, i_13_438_3932_0, i_13_438_3982_0,
    i_13_438_4006_0, i_13_438_4096_0, i_13_438_4115_0, i_13_438_4158_0,
    i_13_438_4160_0, i_13_438_4162_0, i_13_438_4163_0, i_13_438_4261_0,
    i_13_438_4313_0, i_13_438_4315_0, i_13_438_4324_0, i_13_438_4351_0,
    i_13_438_4369_0, i_13_438_4429_0, i_13_438_4441_0, i_13_438_4463_0,
    i_13_438_4510_0, i_13_438_4537_0, i_13_438_4540_0, i_13_438_4541_0,
    o_13_438_0_0  );
  input  i_13_438_29_0, i_13_438_45_0, i_13_438_107_0, i_13_438_271_0,
    i_13_438_300_0, i_13_438_352_0, i_13_438_374_0, i_13_438_422_0,
    i_13_438_451_0, i_13_438_559_0, i_13_438_561_0, i_13_438_562_0,
    i_13_438_569_0, i_13_438_604_0, i_13_438_605_0, i_13_438_607_0,
    i_13_438_608_0, i_13_438_610_0, i_13_438_658_0, i_13_438_659_0,
    i_13_438_661_0, i_13_438_662_0, i_13_438_670_0, i_13_438_680_0,
    i_13_438_829_0, i_13_438_832_0, i_13_438_833_0, i_13_438_882_0,
    i_13_438_885_0, i_13_438_886_0, i_13_438_946_0, i_13_438_1075_0,
    i_13_438_1084_0, i_13_438_1226_0, i_13_438_1281_0, i_13_438_1381_0,
    i_13_438_1404_0, i_13_438_1405_0, i_13_438_1467_0, i_13_438_1520_0,
    i_13_438_1522_0, i_13_438_1535_0, i_13_438_1660_0, i_13_438_1768_0,
    i_13_438_1787_0, i_13_438_1802_0, i_13_438_1838_0, i_13_438_1846_0,
    i_13_438_1885_0, i_13_438_1897_0, i_13_438_1927_0, i_13_438_2021_0,
    i_13_438_2137_0, i_13_438_2170_0, i_13_438_2297_0, i_13_438_2423_0,
    i_13_438_2431_0, i_13_438_2435_0, i_13_438_2647_0, i_13_438_2650_0,
    i_13_438_2749_0, i_13_438_2880_0, i_13_438_3047_0, i_13_438_3106_0,
    i_13_438_3117_0, i_13_438_3311_0, i_13_438_3457_0, i_13_438_3476_0,
    i_13_438_3547_0, i_13_438_3638_0, i_13_438_3664_0, i_13_438_3683_0,
    i_13_438_3740_0, i_13_438_3844_0, i_13_438_3871_0, i_13_438_3872_0,
    i_13_438_3889_0, i_13_438_3910_0, i_13_438_3932_0, i_13_438_3982_0,
    i_13_438_4006_0, i_13_438_4096_0, i_13_438_4115_0, i_13_438_4158_0,
    i_13_438_4160_0, i_13_438_4162_0, i_13_438_4163_0, i_13_438_4261_0,
    i_13_438_4313_0, i_13_438_4315_0, i_13_438_4324_0, i_13_438_4351_0,
    i_13_438_4369_0, i_13_438_4429_0, i_13_438_4441_0, i_13_438_4463_0,
    i_13_438_4510_0, i_13_438_4537_0, i_13_438_4540_0, i_13_438_4541_0;
  output o_13_438_0_0;
  assign o_13_438_0_0 = ~((~i_13_438_562_0 & ~i_13_438_4510_0) | (~i_13_438_1660_0 & i_13_438_1885_0 & ~i_13_438_2431_0) | (~i_13_438_1838_0 & ~i_13_438_3547_0 & ~i_13_438_4006_0 & ~i_13_438_4158_0));
endmodule



// Benchmark "kernel_13_439" written by ABC on Sun Jul 19 10:51:29 2020

module kernel_13_439 ( 
    i_13_439_108_0, i_13_439_112_0, i_13_439_171_0, i_13_439_282_0,
    i_13_439_336_0, i_13_439_594_0, i_13_439_639_0, i_13_439_739_0,
    i_13_439_793_0, i_13_439_819_0, i_13_439_820_0, i_13_439_847_0,
    i_13_439_855_0, i_13_439_856_0, i_13_439_868_0, i_13_439_894_0,
    i_13_439_1017_0, i_13_439_1120_0, i_13_439_1215_0, i_13_439_1224_0,
    i_13_439_1251_0, i_13_439_1252_0, i_13_439_1278_0, i_13_439_1279_0,
    i_13_439_1299_0, i_13_439_1309_0, i_13_439_1395_0, i_13_439_1422_0,
    i_13_439_1440_0, i_13_439_1467_0, i_13_439_1485_0, i_13_439_1486_0,
    i_13_439_1490_0, i_13_439_1494_0, i_13_439_1548_0, i_13_439_1549_0,
    i_13_439_1570_0, i_13_439_1629_0, i_13_439_1630_0, i_13_439_1693_0,
    i_13_439_1792_0, i_13_439_1827_0, i_13_439_1855_0, i_13_439_1857_0,
    i_13_439_1954_0, i_13_439_1998_0, i_13_439_1999_0, i_13_439_2044_0,
    i_13_439_2060_0, i_13_439_2172_0, i_13_439_2196_0, i_13_439_2377_0,
    i_13_439_2380_0, i_13_439_2394_0, i_13_439_2421_0, i_13_439_2422_0,
    i_13_439_2457_0, i_13_439_2494_0, i_13_439_2501_0, i_13_439_2529_0,
    i_13_439_2530_0, i_13_439_2538_0, i_13_439_2539_0, i_13_439_2542_0,
    i_13_439_2543_0, i_13_439_2592_0, i_13_439_2610_0, i_13_439_2712_0,
    i_13_439_2716_0, i_13_439_2728_0, i_13_439_2817_0, i_13_439_2902_0,
    i_13_439_2916_0, i_13_439_2917_0, i_13_439_2997_0, i_13_439_3025_0,
    i_13_439_3123_0, i_13_439_3144_0, i_13_439_3145_0, i_13_439_3168_0,
    i_13_439_3370_0, i_13_439_3420_0, i_13_439_3442_0, i_13_439_3465_0,
    i_13_439_3475_0, i_13_439_3483_0, i_13_439_3780_0, i_13_439_3870_0,
    i_13_439_3871_0, i_13_439_3991_0, i_13_439_4005_0, i_13_439_4006_0,
    i_13_439_4114_0, i_13_439_4185_0, i_13_439_4230_0, i_13_439_4248_0,
    i_13_439_4249_0, i_13_439_4251_0, i_13_439_4342_0, i_13_439_4374_0,
    o_13_439_0_0  );
  input  i_13_439_108_0, i_13_439_112_0, i_13_439_171_0, i_13_439_282_0,
    i_13_439_336_0, i_13_439_594_0, i_13_439_639_0, i_13_439_739_0,
    i_13_439_793_0, i_13_439_819_0, i_13_439_820_0, i_13_439_847_0,
    i_13_439_855_0, i_13_439_856_0, i_13_439_868_0, i_13_439_894_0,
    i_13_439_1017_0, i_13_439_1120_0, i_13_439_1215_0, i_13_439_1224_0,
    i_13_439_1251_0, i_13_439_1252_0, i_13_439_1278_0, i_13_439_1279_0,
    i_13_439_1299_0, i_13_439_1309_0, i_13_439_1395_0, i_13_439_1422_0,
    i_13_439_1440_0, i_13_439_1467_0, i_13_439_1485_0, i_13_439_1486_0,
    i_13_439_1490_0, i_13_439_1494_0, i_13_439_1548_0, i_13_439_1549_0,
    i_13_439_1570_0, i_13_439_1629_0, i_13_439_1630_0, i_13_439_1693_0,
    i_13_439_1792_0, i_13_439_1827_0, i_13_439_1855_0, i_13_439_1857_0,
    i_13_439_1954_0, i_13_439_1998_0, i_13_439_1999_0, i_13_439_2044_0,
    i_13_439_2060_0, i_13_439_2172_0, i_13_439_2196_0, i_13_439_2377_0,
    i_13_439_2380_0, i_13_439_2394_0, i_13_439_2421_0, i_13_439_2422_0,
    i_13_439_2457_0, i_13_439_2494_0, i_13_439_2501_0, i_13_439_2529_0,
    i_13_439_2530_0, i_13_439_2538_0, i_13_439_2539_0, i_13_439_2542_0,
    i_13_439_2543_0, i_13_439_2592_0, i_13_439_2610_0, i_13_439_2712_0,
    i_13_439_2716_0, i_13_439_2728_0, i_13_439_2817_0, i_13_439_2902_0,
    i_13_439_2916_0, i_13_439_2917_0, i_13_439_2997_0, i_13_439_3025_0,
    i_13_439_3123_0, i_13_439_3144_0, i_13_439_3145_0, i_13_439_3168_0,
    i_13_439_3370_0, i_13_439_3420_0, i_13_439_3442_0, i_13_439_3465_0,
    i_13_439_3475_0, i_13_439_3483_0, i_13_439_3780_0, i_13_439_3870_0,
    i_13_439_3871_0, i_13_439_3991_0, i_13_439_4005_0, i_13_439_4006_0,
    i_13_439_4114_0, i_13_439_4185_0, i_13_439_4230_0, i_13_439_4248_0,
    i_13_439_4249_0, i_13_439_4251_0, i_13_439_4342_0, i_13_439_4374_0;
  output o_13_439_0_0;
  assign o_13_439_0_0 = ~((~i_13_439_2172_0 & ~i_13_439_4249_0) | (~i_13_439_855_0 & ~i_13_439_1215_0 & i_13_439_2542_0) | (~i_13_439_1017_0 & ~i_13_439_1485_0 & ~i_13_439_3871_0 & ~i_13_439_4005_0));
endmodule



// Benchmark "kernel_13_440" written by ABC on Sun Jul 19 10:51:30 2020

module kernel_13_440 ( 
    i_13_440_52_0, i_13_440_71_0, i_13_440_76_0, i_13_440_112_0,
    i_13_440_113_0, i_13_440_241_0, i_13_440_251_0, i_13_440_273_0,
    i_13_440_278_0, i_13_440_284_0, i_13_440_341_0, i_13_440_594_0,
    i_13_440_619_0, i_13_440_855_0, i_13_440_878_0, i_13_440_1102_0,
    i_13_440_1120_0, i_13_440_1273_0, i_13_440_1309_0, i_13_440_1364_0,
    i_13_440_1426_0, i_13_440_1474_0, i_13_440_1525_0, i_13_440_1573_0,
    i_13_440_1597_0, i_13_440_1629_0, i_13_440_1633_0, i_13_440_1634_0,
    i_13_440_1642_0, i_13_440_1669_0, i_13_440_1741_0, i_13_440_1753_0,
    i_13_440_1795_0, i_13_440_1796_0, i_13_440_1816_0, i_13_440_1817_0,
    i_13_440_1939_0, i_13_440_2452_0, i_13_440_2455_0, i_13_440_2465_0,
    i_13_440_2497_0, i_13_440_2501_0, i_13_440_2561_0, i_13_440_2570_0,
    i_13_440_2712_0, i_13_440_2713_0, i_13_440_2715_0, i_13_440_2716_0,
    i_13_440_2761_0, i_13_440_2884_0, i_13_440_2920_0, i_13_440_2942_0,
    i_13_440_2983_0, i_13_440_3004_0, i_13_440_3010_0, i_13_440_3067_0,
    i_13_440_3101_0, i_13_440_3145_0, i_13_440_3148_0, i_13_440_3201_0,
    i_13_440_3238_0, i_13_440_3292_0, i_13_440_3310_0, i_13_440_3328_0,
    i_13_440_3329_0, i_13_440_3391_0, i_13_440_3406_0, i_13_440_3417_0,
    i_13_440_3451_0, i_13_440_3454_0, i_13_440_3455_0, i_13_440_3477_0,
    i_13_440_3527_0, i_13_440_3541_0, i_13_440_3599_0, i_13_440_3646_0,
    i_13_440_3660_0, i_13_440_3684_0, i_13_440_3687_0, i_13_440_3688_0,
    i_13_440_3689_0, i_13_440_3730_0, i_13_440_3832_0, i_13_440_3874_0,
    i_13_440_3922_0, i_13_440_3982_0, i_13_440_4021_0, i_13_440_4036_0,
    i_13_440_4057_0, i_13_440_4093_0, i_13_440_4157_0, i_13_440_4158_0,
    i_13_440_4274_0, i_13_440_4408_0, i_13_440_4409_0, i_13_440_4427_0,
    i_13_440_4522_0, i_13_440_4543_0, i_13_440_4558_0, i_13_440_4594_0,
    o_13_440_0_0  );
  input  i_13_440_52_0, i_13_440_71_0, i_13_440_76_0, i_13_440_112_0,
    i_13_440_113_0, i_13_440_241_0, i_13_440_251_0, i_13_440_273_0,
    i_13_440_278_0, i_13_440_284_0, i_13_440_341_0, i_13_440_594_0,
    i_13_440_619_0, i_13_440_855_0, i_13_440_878_0, i_13_440_1102_0,
    i_13_440_1120_0, i_13_440_1273_0, i_13_440_1309_0, i_13_440_1364_0,
    i_13_440_1426_0, i_13_440_1474_0, i_13_440_1525_0, i_13_440_1573_0,
    i_13_440_1597_0, i_13_440_1629_0, i_13_440_1633_0, i_13_440_1634_0,
    i_13_440_1642_0, i_13_440_1669_0, i_13_440_1741_0, i_13_440_1753_0,
    i_13_440_1795_0, i_13_440_1796_0, i_13_440_1816_0, i_13_440_1817_0,
    i_13_440_1939_0, i_13_440_2452_0, i_13_440_2455_0, i_13_440_2465_0,
    i_13_440_2497_0, i_13_440_2501_0, i_13_440_2561_0, i_13_440_2570_0,
    i_13_440_2712_0, i_13_440_2713_0, i_13_440_2715_0, i_13_440_2716_0,
    i_13_440_2761_0, i_13_440_2884_0, i_13_440_2920_0, i_13_440_2942_0,
    i_13_440_2983_0, i_13_440_3004_0, i_13_440_3010_0, i_13_440_3067_0,
    i_13_440_3101_0, i_13_440_3145_0, i_13_440_3148_0, i_13_440_3201_0,
    i_13_440_3238_0, i_13_440_3292_0, i_13_440_3310_0, i_13_440_3328_0,
    i_13_440_3329_0, i_13_440_3391_0, i_13_440_3406_0, i_13_440_3417_0,
    i_13_440_3451_0, i_13_440_3454_0, i_13_440_3455_0, i_13_440_3477_0,
    i_13_440_3527_0, i_13_440_3541_0, i_13_440_3599_0, i_13_440_3646_0,
    i_13_440_3660_0, i_13_440_3684_0, i_13_440_3687_0, i_13_440_3688_0,
    i_13_440_3689_0, i_13_440_3730_0, i_13_440_3832_0, i_13_440_3874_0,
    i_13_440_3922_0, i_13_440_3982_0, i_13_440_4021_0, i_13_440_4036_0,
    i_13_440_4057_0, i_13_440_4093_0, i_13_440_4157_0, i_13_440_4158_0,
    i_13_440_4274_0, i_13_440_4408_0, i_13_440_4409_0, i_13_440_4427_0,
    i_13_440_4522_0, i_13_440_4543_0, i_13_440_4558_0, i_13_440_4594_0;
  output o_13_440_0_0;
  assign o_13_440_0_0 = ~((~i_13_440_3455_0 & ((i_13_440_1597_0 & ~i_13_440_2455_0 & ~i_13_440_2920_0) | (~i_13_440_273_0 & ~i_13_440_2942_0 & ~i_13_440_3684_0))) | (~i_13_440_3688_0 & (~i_13_440_3148_0 | (i_13_440_4036_0 & ~i_13_440_4274_0))) | (~i_13_440_1573_0 & ~i_13_440_3689_0 & ~i_13_440_4558_0));
endmodule



// Benchmark "kernel_13_441" written by ABC on Sun Jul 19 10:51:31 2020

module kernel_13_441 ( 
    i_13_441_31_0, i_13_441_48_0, i_13_441_49_0, i_13_441_51_0,
    i_13_441_67_0, i_13_441_124_0, i_13_441_139_0, i_13_441_229_0,
    i_13_441_247_0, i_13_441_257_0, i_13_441_492_0, i_13_441_493_0,
    i_13_441_515_0, i_13_441_652_0, i_13_441_672_0, i_13_441_678_0,
    i_13_441_816_0, i_13_441_840_0, i_13_441_843_0, i_13_441_853_0,
    i_13_441_942_0, i_13_441_979_0, i_13_441_984_0, i_13_441_985_0,
    i_13_441_1191_0, i_13_441_1267_0, i_13_441_1326_0, i_13_441_1327_0,
    i_13_441_1329_0, i_13_441_1330_0, i_13_441_1509_0, i_13_441_1572_0,
    i_13_441_1681_0, i_13_441_1686_0, i_13_441_1723_0, i_13_441_1852_0,
    i_13_441_1908_0, i_13_441_2002_0, i_13_441_2022_0, i_13_441_2028_0,
    i_13_441_2148_0, i_13_441_2184_0, i_13_441_2229_0, i_13_441_2265_0,
    i_13_441_2277_0, i_13_441_2302_0, i_13_441_2318_0, i_13_441_2472_0,
    i_13_441_2506_0, i_13_441_2508_0, i_13_441_2509_0, i_13_441_2697_0,
    i_13_441_2698_0, i_13_441_2742_0, i_13_441_2743_0, i_13_441_2748_0,
    i_13_441_2751_0, i_13_441_2752_0, i_13_441_2874_0, i_13_441_2875_0,
    i_13_441_2958_0, i_13_441_2967_0, i_13_441_2973_0, i_13_441_3013_0,
    i_13_441_3058_0, i_13_441_3108_0, i_13_441_3115_0, i_13_441_3118_0,
    i_13_441_3144_0, i_13_441_3172_0, i_13_441_3210_0, i_13_441_3291_0,
    i_13_441_3315_0, i_13_441_3349_0, i_13_441_3372_0, i_13_441_3405_0,
    i_13_441_3418_0, i_13_441_3453_0, i_13_441_3463_0, i_13_441_3489_0,
    i_13_441_3490_0, i_13_441_3522_0, i_13_441_3525_0, i_13_441_3546_0,
    i_13_441_3552_0, i_13_441_3706_0, i_13_441_3765_0, i_13_441_3766_0,
    i_13_441_3769_0, i_13_441_3865_0, i_13_441_3876_0, i_13_441_3903_0,
    i_13_441_3994_0, i_13_441_4089_0, i_13_441_4161_0, i_13_441_4174_0,
    i_13_441_4318_0, i_13_441_4331_0, i_13_441_4495_0, i_13_441_4560_0,
    o_13_441_0_0  );
  input  i_13_441_31_0, i_13_441_48_0, i_13_441_49_0, i_13_441_51_0,
    i_13_441_67_0, i_13_441_124_0, i_13_441_139_0, i_13_441_229_0,
    i_13_441_247_0, i_13_441_257_0, i_13_441_492_0, i_13_441_493_0,
    i_13_441_515_0, i_13_441_652_0, i_13_441_672_0, i_13_441_678_0,
    i_13_441_816_0, i_13_441_840_0, i_13_441_843_0, i_13_441_853_0,
    i_13_441_942_0, i_13_441_979_0, i_13_441_984_0, i_13_441_985_0,
    i_13_441_1191_0, i_13_441_1267_0, i_13_441_1326_0, i_13_441_1327_0,
    i_13_441_1329_0, i_13_441_1330_0, i_13_441_1509_0, i_13_441_1572_0,
    i_13_441_1681_0, i_13_441_1686_0, i_13_441_1723_0, i_13_441_1852_0,
    i_13_441_1908_0, i_13_441_2002_0, i_13_441_2022_0, i_13_441_2028_0,
    i_13_441_2148_0, i_13_441_2184_0, i_13_441_2229_0, i_13_441_2265_0,
    i_13_441_2277_0, i_13_441_2302_0, i_13_441_2318_0, i_13_441_2472_0,
    i_13_441_2506_0, i_13_441_2508_0, i_13_441_2509_0, i_13_441_2697_0,
    i_13_441_2698_0, i_13_441_2742_0, i_13_441_2743_0, i_13_441_2748_0,
    i_13_441_2751_0, i_13_441_2752_0, i_13_441_2874_0, i_13_441_2875_0,
    i_13_441_2958_0, i_13_441_2967_0, i_13_441_2973_0, i_13_441_3013_0,
    i_13_441_3058_0, i_13_441_3108_0, i_13_441_3115_0, i_13_441_3118_0,
    i_13_441_3144_0, i_13_441_3172_0, i_13_441_3210_0, i_13_441_3291_0,
    i_13_441_3315_0, i_13_441_3349_0, i_13_441_3372_0, i_13_441_3405_0,
    i_13_441_3418_0, i_13_441_3453_0, i_13_441_3463_0, i_13_441_3489_0,
    i_13_441_3490_0, i_13_441_3522_0, i_13_441_3525_0, i_13_441_3546_0,
    i_13_441_3552_0, i_13_441_3706_0, i_13_441_3765_0, i_13_441_3766_0,
    i_13_441_3769_0, i_13_441_3865_0, i_13_441_3876_0, i_13_441_3903_0,
    i_13_441_3994_0, i_13_441_4089_0, i_13_441_4161_0, i_13_441_4174_0,
    i_13_441_4318_0, i_13_441_4331_0, i_13_441_4495_0, i_13_441_4560_0;
  output o_13_441_0_0;
  assign o_13_441_0_0 = ~((~i_13_441_984_0 & ~i_13_441_1326_0) | (~i_13_441_1330_0 & ~i_13_441_2697_0 & ~i_13_441_2742_0 & ~i_13_441_4318_0));
endmodule



// Benchmark "kernel_13_442" written by ABC on Sun Jul 19 10:51:31 2020

module kernel_13_442 ( 
    i_13_442_184_0, i_13_442_259_0, i_13_442_285_0, i_13_442_286_0,
    i_13_442_310_0, i_13_442_357_0, i_13_442_454_0, i_13_442_466_0,
    i_13_442_503_0, i_13_442_592_0, i_13_442_636_0, i_13_442_683_0,
    i_13_442_690_0, i_13_442_841_0, i_13_442_952_0, i_13_442_1111_0,
    i_13_442_1213_0, i_13_442_1218_0, i_13_442_1219_0, i_13_442_1261_0,
    i_13_442_1263_0, i_13_442_1313_0, i_13_442_1318_0, i_13_442_1347_0,
    i_13_442_1348_0, i_13_442_1364_0, i_13_442_1427_0, i_13_442_1447_0,
    i_13_442_1462_0, i_13_442_1525_0, i_13_442_1529_0, i_13_442_1561_0,
    i_13_442_1678_0, i_13_442_1868_0, i_13_442_1894_0, i_13_442_1933_0,
    i_13_442_1941_0, i_13_442_1993_0, i_13_442_2001_0, i_13_442_2002_0,
    i_13_442_2003_0, i_13_442_2005_0, i_13_442_2058_0, i_13_442_2059_0,
    i_13_442_2060_0, i_13_442_2146_0, i_13_442_2149_0, i_13_442_2236_0,
    i_13_442_2283_0, i_13_442_2284_0, i_13_442_2285_0, i_13_442_2299_0,
    i_13_442_2407_0, i_13_442_2425_0, i_13_442_2456_0, i_13_442_2554_0,
    i_13_442_2589_0, i_13_442_2590_0, i_13_442_2610_0, i_13_442_2653_0,
    i_13_442_2654_0, i_13_442_2658_0, i_13_442_2681_0, i_13_442_2743_0,
    i_13_442_2824_0, i_13_442_2856_0, i_13_442_2860_0, i_13_442_2906_0,
    i_13_442_2956_0, i_13_442_3146_0, i_13_442_3148_0, i_13_442_3220_0,
    i_13_442_3316_0, i_13_442_3345_0, i_13_442_3391_0, i_13_442_3392_0,
    i_13_442_3482_0, i_13_442_3553_0, i_13_442_3580_0, i_13_442_3598_0,
    i_13_442_3633_0, i_13_442_3729_0, i_13_442_3732_0, i_13_442_3734_0,
    i_13_442_3787_0, i_13_442_3994_0, i_13_442_4020_0, i_13_442_4114_0,
    i_13_442_4237_0, i_13_442_4263_0, i_13_442_4264_0, i_13_442_4310_0,
    i_13_442_4333_0, i_13_442_4363_0, i_13_442_4398_0, i_13_442_4399_0,
    i_13_442_4400_0, i_13_442_4534_0, i_13_442_4567_0, i_13_442_4598_0,
    o_13_442_0_0  );
  input  i_13_442_184_0, i_13_442_259_0, i_13_442_285_0, i_13_442_286_0,
    i_13_442_310_0, i_13_442_357_0, i_13_442_454_0, i_13_442_466_0,
    i_13_442_503_0, i_13_442_592_0, i_13_442_636_0, i_13_442_683_0,
    i_13_442_690_0, i_13_442_841_0, i_13_442_952_0, i_13_442_1111_0,
    i_13_442_1213_0, i_13_442_1218_0, i_13_442_1219_0, i_13_442_1261_0,
    i_13_442_1263_0, i_13_442_1313_0, i_13_442_1318_0, i_13_442_1347_0,
    i_13_442_1348_0, i_13_442_1364_0, i_13_442_1427_0, i_13_442_1447_0,
    i_13_442_1462_0, i_13_442_1525_0, i_13_442_1529_0, i_13_442_1561_0,
    i_13_442_1678_0, i_13_442_1868_0, i_13_442_1894_0, i_13_442_1933_0,
    i_13_442_1941_0, i_13_442_1993_0, i_13_442_2001_0, i_13_442_2002_0,
    i_13_442_2003_0, i_13_442_2005_0, i_13_442_2058_0, i_13_442_2059_0,
    i_13_442_2060_0, i_13_442_2146_0, i_13_442_2149_0, i_13_442_2236_0,
    i_13_442_2283_0, i_13_442_2284_0, i_13_442_2285_0, i_13_442_2299_0,
    i_13_442_2407_0, i_13_442_2425_0, i_13_442_2456_0, i_13_442_2554_0,
    i_13_442_2589_0, i_13_442_2590_0, i_13_442_2610_0, i_13_442_2653_0,
    i_13_442_2654_0, i_13_442_2658_0, i_13_442_2681_0, i_13_442_2743_0,
    i_13_442_2824_0, i_13_442_2856_0, i_13_442_2860_0, i_13_442_2906_0,
    i_13_442_2956_0, i_13_442_3146_0, i_13_442_3148_0, i_13_442_3220_0,
    i_13_442_3316_0, i_13_442_3345_0, i_13_442_3391_0, i_13_442_3392_0,
    i_13_442_3482_0, i_13_442_3553_0, i_13_442_3580_0, i_13_442_3598_0,
    i_13_442_3633_0, i_13_442_3729_0, i_13_442_3732_0, i_13_442_3734_0,
    i_13_442_3787_0, i_13_442_3994_0, i_13_442_4020_0, i_13_442_4114_0,
    i_13_442_4237_0, i_13_442_4263_0, i_13_442_4264_0, i_13_442_4310_0,
    i_13_442_4333_0, i_13_442_4363_0, i_13_442_4398_0, i_13_442_4399_0,
    i_13_442_4400_0, i_13_442_4534_0, i_13_442_4567_0, i_13_442_4598_0;
  output o_13_442_0_0;
  assign o_13_442_0_0 = ~((~i_13_442_2285_0 & ((~i_13_442_1348_0 & i_13_442_2149_0) | (~i_13_442_592_0 & ~i_13_442_3220_0 & ~i_13_442_3734_0 & ~i_13_442_4263_0))) | (i_13_442_1678_0 & ~i_13_442_2425_0 & ~i_13_442_4264_0 & ~i_13_442_4400_0));
endmodule



// Benchmark "kernel_13_443" written by ABC on Sun Jul 19 10:51:32 2020

module kernel_13_443 ( 
    i_13_443_62_0, i_13_443_117_0, i_13_443_134_0, i_13_443_136_0,
    i_13_443_174_0, i_13_443_283_0, i_13_443_333_0, i_13_443_351_0,
    i_13_443_489_0, i_13_443_493_0, i_13_443_599_0, i_13_443_612_0,
    i_13_443_617_0, i_13_443_624_0, i_13_443_828_0, i_13_443_889_0,
    i_13_443_1098_0, i_13_443_1099_0, i_13_443_1100_0, i_13_443_1116_0,
    i_13_443_1123_0, i_13_443_1128_0, i_13_443_1132_0, i_13_443_1208_0,
    i_13_443_1256_0, i_13_443_1394_0, i_13_443_1429_0, i_13_443_1442_0,
    i_13_443_1517_0, i_13_443_1521_0, i_13_443_1522_0, i_13_443_1639_0,
    i_13_443_1699_0, i_13_443_1745_0, i_13_443_1754_0, i_13_443_1811_0,
    i_13_443_1958_0, i_13_443_2111_0, i_13_443_2142_0, i_13_443_2143_0,
    i_13_443_2208_0, i_13_443_2295_0, i_13_443_2296_0, i_13_443_2300_0,
    i_13_443_2380_0, i_13_443_2402_0, i_13_443_2423_0, i_13_443_2438_0,
    i_13_443_2442_0, i_13_443_2464_0, i_13_443_2511_0, i_13_443_2781_0,
    i_13_443_2880_0, i_13_443_2986_0, i_13_443_3015_0, i_13_443_3065_0,
    i_13_443_3090_0, i_13_443_3094_0, i_13_443_3133_0, i_13_443_3171_0,
    i_13_443_3196_0, i_13_443_3241_0, i_13_443_3269_0, i_13_443_3307_0,
    i_13_443_3339_0, i_13_443_3366_0, i_13_443_3368_0, i_13_443_3429_0,
    i_13_443_3474_0, i_13_443_3537_0, i_13_443_3547_0, i_13_443_3636_0,
    i_13_443_3637_0, i_13_443_3685_0, i_13_443_3699_0, i_13_443_3753_0,
    i_13_443_3754_0, i_13_443_3765_0, i_13_443_3855_0, i_13_443_3889_0,
    i_13_443_3896_0, i_13_443_3910_0, i_13_443_3978_0, i_13_443_3985_0,
    i_13_443_4017_0, i_13_443_4018_0, i_13_443_4216_0, i_13_443_4297_0,
    i_13_443_4311_0, i_13_443_4312_0, i_13_443_4315_0, i_13_443_4321_0,
    i_13_443_4336_0, i_13_443_4394_0, i_13_443_4414_0, i_13_443_4509_0,
    i_13_443_4513_0, i_13_443_4514_0, i_13_443_4568_0, i_13_443_4598_0,
    o_13_443_0_0  );
  input  i_13_443_62_0, i_13_443_117_0, i_13_443_134_0, i_13_443_136_0,
    i_13_443_174_0, i_13_443_283_0, i_13_443_333_0, i_13_443_351_0,
    i_13_443_489_0, i_13_443_493_0, i_13_443_599_0, i_13_443_612_0,
    i_13_443_617_0, i_13_443_624_0, i_13_443_828_0, i_13_443_889_0,
    i_13_443_1098_0, i_13_443_1099_0, i_13_443_1100_0, i_13_443_1116_0,
    i_13_443_1123_0, i_13_443_1128_0, i_13_443_1132_0, i_13_443_1208_0,
    i_13_443_1256_0, i_13_443_1394_0, i_13_443_1429_0, i_13_443_1442_0,
    i_13_443_1517_0, i_13_443_1521_0, i_13_443_1522_0, i_13_443_1639_0,
    i_13_443_1699_0, i_13_443_1745_0, i_13_443_1754_0, i_13_443_1811_0,
    i_13_443_1958_0, i_13_443_2111_0, i_13_443_2142_0, i_13_443_2143_0,
    i_13_443_2208_0, i_13_443_2295_0, i_13_443_2296_0, i_13_443_2300_0,
    i_13_443_2380_0, i_13_443_2402_0, i_13_443_2423_0, i_13_443_2438_0,
    i_13_443_2442_0, i_13_443_2464_0, i_13_443_2511_0, i_13_443_2781_0,
    i_13_443_2880_0, i_13_443_2986_0, i_13_443_3015_0, i_13_443_3065_0,
    i_13_443_3090_0, i_13_443_3094_0, i_13_443_3133_0, i_13_443_3171_0,
    i_13_443_3196_0, i_13_443_3241_0, i_13_443_3269_0, i_13_443_3307_0,
    i_13_443_3339_0, i_13_443_3366_0, i_13_443_3368_0, i_13_443_3429_0,
    i_13_443_3474_0, i_13_443_3537_0, i_13_443_3547_0, i_13_443_3636_0,
    i_13_443_3637_0, i_13_443_3685_0, i_13_443_3699_0, i_13_443_3753_0,
    i_13_443_3754_0, i_13_443_3765_0, i_13_443_3855_0, i_13_443_3889_0,
    i_13_443_3896_0, i_13_443_3910_0, i_13_443_3978_0, i_13_443_3985_0,
    i_13_443_4017_0, i_13_443_4018_0, i_13_443_4216_0, i_13_443_4297_0,
    i_13_443_4311_0, i_13_443_4312_0, i_13_443_4315_0, i_13_443_4321_0,
    i_13_443_4336_0, i_13_443_4394_0, i_13_443_4414_0, i_13_443_4509_0,
    i_13_443_4513_0, i_13_443_4514_0, i_13_443_4568_0, i_13_443_4598_0;
  output o_13_443_0_0;
  assign o_13_443_0_0 = ~((~i_13_443_4509_0 & (i_13_443_3685_0 | (~i_13_443_1208_0 & ~i_13_443_3978_0) | (i_13_443_3910_0 & ~i_13_443_4216_0 & ~i_13_443_4311_0))) | (~i_13_443_2142_0 & ~i_13_443_3754_0 & ~i_13_443_4321_0) | (~i_13_443_4312_0 & i_13_443_4394_0));
endmodule



// Benchmark "kernel_13_444" written by ABC on Sun Jul 19 10:51:33 2020

module kernel_13_444 ( 
    i_13_444_48_0, i_13_444_49_0, i_13_444_70_0, i_13_444_107_0,
    i_13_444_178_0, i_13_444_411_0, i_13_444_448_0, i_13_444_535_0,
    i_13_444_570_0, i_13_444_610_0, i_13_444_616_0, i_13_444_645_0,
    i_13_444_760_0, i_13_444_762_0, i_13_444_797_0, i_13_444_933_0,
    i_13_444_934_0, i_13_444_939_0, i_13_444_1083_0, i_13_444_1101_0,
    i_13_444_1104_0, i_13_444_1131_0, i_13_444_1132_0, i_13_444_1137_0,
    i_13_444_1276_0, i_13_444_1285_0, i_13_444_1428_0, i_13_444_1482_0,
    i_13_444_1506_0, i_13_444_1509_0, i_13_444_1510_0, i_13_444_1515_0,
    i_13_444_1574_0, i_13_444_1626_0, i_13_444_1634_0, i_13_444_1644_0,
    i_13_444_1651_0, i_13_444_1716_0, i_13_444_1735_0, i_13_444_1767_0,
    i_13_444_1768_0, i_13_444_1770_0, i_13_444_1797_0, i_13_444_1798_0,
    i_13_444_1804_0, i_13_444_1841_0, i_13_444_1884_0, i_13_444_1945_0,
    i_13_444_1957_0, i_13_444_1995_0, i_13_444_2022_0, i_13_444_2023_0,
    i_13_444_2049_0, i_13_444_2122_0, i_13_444_2348_0, i_13_444_2454_0,
    i_13_444_2472_0, i_13_444_2473_0, i_13_444_2483_0, i_13_444_2501_0,
    i_13_444_2615_0, i_13_444_2679_0, i_13_444_2724_0, i_13_444_2913_0,
    i_13_444_2937_0, i_13_444_3031_0, i_13_444_3076_0, i_13_444_3120_0,
    i_13_444_3164_0, i_13_444_3263_0, i_13_444_3264_0, i_13_444_3274_0,
    i_13_444_3351_0, i_13_444_3389_0, i_13_444_3399_0, i_13_444_3417_0,
    i_13_444_3418_0, i_13_444_3455_0, i_13_444_3570_0, i_13_444_3613_0,
    i_13_444_3640_0, i_13_444_3651_0, i_13_444_3783_0, i_13_444_3813_0,
    i_13_444_3822_0, i_13_444_3823_0, i_13_444_3900_0, i_13_444_3940_0,
    i_13_444_3982_0, i_13_444_4084_0, i_13_444_4164_0, i_13_444_4193_0,
    i_13_444_4300_0, i_13_444_4308_0, i_13_444_4324_0, i_13_444_4400_0,
    i_13_444_4596_0, i_13_444_4597_0, i_13_444_4605_0, i_13_444_4606_0,
    o_13_444_0_0  );
  input  i_13_444_48_0, i_13_444_49_0, i_13_444_70_0, i_13_444_107_0,
    i_13_444_178_0, i_13_444_411_0, i_13_444_448_0, i_13_444_535_0,
    i_13_444_570_0, i_13_444_610_0, i_13_444_616_0, i_13_444_645_0,
    i_13_444_760_0, i_13_444_762_0, i_13_444_797_0, i_13_444_933_0,
    i_13_444_934_0, i_13_444_939_0, i_13_444_1083_0, i_13_444_1101_0,
    i_13_444_1104_0, i_13_444_1131_0, i_13_444_1132_0, i_13_444_1137_0,
    i_13_444_1276_0, i_13_444_1285_0, i_13_444_1428_0, i_13_444_1482_0,
    i_13_444_1506_0, i_13_444_1509_0, i_13_444_1510_0, i_13_444_1515_0,
    i_13_444_1574_0, i_13_444_1626_0, i_13_444_1634_0, i_13_444_1644_0,
    i_13_444_1651_0, i_13_444_1716_0, i_13_444_1735_0, i_13_444_1767_0,
    i_13_444_1768_0, i_13_444_1770_0, i_13_444_1797_0, i_13_444_1798_0,
    i_13_444_1804_0, i_13_444_1841_0, i_13_444_1884_0, i_13_444_1945_0,
    i_13_444_1957_0, i_13_444_1995_0, i_13_444_2022_0, i_13_444_2023_0,
    i_13_444_2049_0, i_13_444_2122_0, i_13_444_2348_0, i_13_444_2454_0,
    i_13_444_2472_0, i_13_444_2473_0, i_13_444_2483_0, i_13_444_2501_0,
    i_13_444_2615_0, i_13_444_2679_0, i_13_444_2724_0, i_13_444_2913_0,
    i_13_444_2937_0, i_13_444_3031_0, i_13_444_3076_0, i_13_444_3120_0,
    i_13_444_3164_0, i_13_444_3263_0, i_13_444_3264_0, i_13_444_3274_0,
    i_13_444_3351_0, i_13_444_3389_0, i_13_444_3399_0, i_13_444_3417_0,
    i_13_444_3418_0, i_13_444_3455_0, i_13_444_3570_0, i_13_444_3613_0,
    i_13_444_3640_0, i_13_444_3651_0, i_13_444_3783_0, i_13_444_3813_0,
    i_13_444_3822_0, i_13_444_3823_0, i_13_444_3900_0, i_13_444_3940_0,
    i_13_444_3982_0, i_13_444_4084_0, i_13_444_4164_0, i_13_444_4193_0,
    i_13_444_4300_0, i_13_444_4308_0, i_13_444_4324_0, i_13_444_4400_0,
    i_13_444_4596_0, i_13_444_4597_0, i_13_444_4605_0, i_13_444_4606_0;
  output o_13_444_0_0;
  assign o_13_444_0_0 = 0;
endmodule



// Benchmark "kernel_13_445" written by ABC on Sun Jul 19 10:51:34 2020

module kernel_13_445 ( 
    i_13_445_67_0, i_13_445_68_0, i_13_445_112_0, i_13_445_120_0,
    i_13_445_123_0, i_13_445_175_0, i_13_445_214_0, i_13_445_242_0,
    i_13_445_251_0, i_13_445_259_0, i_13_445_273_0, i_13_445_277_0,
    i_13_445_278_0, i_13_445_283_0, i_13_445_311_0, i_13_445_376_0,
    i_13_445_412_0, i_13_445_454_0, i_13_445_471_0, i_13_445_521_0,
    i_13_445_609_0, i_13_445_620_0, i_13_445_800_0, i_13_445_841_0,
    i_13_445_935_0, i_13_445_980_0, i_13_445_1070_0, i_13_445_1112_0,
    i_13_445_1330_0, i_13_445_1331_0, i_13_445_1389_0, i_13_445_1394_0,
    i_13_445_1398_0, i_13_445_1410_0, i_13_445_1455_0, i_13_445_1472_0,
    i_13_445_1483_0, i_13_445_1512_0, i_13_445_1520_0, i_13_445_1573_0,
    i_13_445_1597_0, i_13_445_1598_0, i_13_445_1642_0, i_13_445_1664_0,
    i_13_445_1674_0, i_13_445_1731_0, i_13_445_1807_0, i_13_445_1835_0,
    i_13_445_1836_0, i_13_445_1945_0, i_13_445_2023_0, i_13_445_2025_0,
    i_13_445_2029_0, i_13_445_2149_0, i_13_445_2186_0, i_13_445_2200_0,
    i_13_445_2303_0, i_13_445_2433_0, i_13_445_2456_0, i_13_445_2698_0,
    i_13_445_2743_0, i_13_445_2744_0, i_13_445_2789_0, i_13_445_2883_0,
    i_13_445_2888_0, i_13_445_2937_0, i_13_445_2942_0, i_13_445_2959_0,
    i_13_445_2969_0, i_13_445_3043_0, i_13_445_3050_0, i_13_445_3077_0,
    i_13_445_3212_0, i_13_445_3238_0, i_13_445_3292_0, i_13_445_3316_0,
    i_13_445_3329_0, i_13_445_3381_0, i_13_445_3419_0, i_13_445_3454_0,
    i_13_445_3526_0, i_13_445_3533_0, i_13_445_3553_0, i_13_445_3596_0,
    i_13_445_3613_0, i_13_445_3689_0, i_13_445_3730_0, i_13_445_3762_0,
    i_13_445_3928_0, i_13_445_4066_0, i_13_445_4173_0, i_13_445_4253_0,
    i_13_445_4274_0, i_13_445_4363_0, i_13_445_4446_0, i_13_445_4503_0,
    i_13_445_4506_0, i_13_445_4517_0, i_13_445_4526_0, i_13_445_4563_0,
    o_13_445_0_0  );
  input  i_13_445_67_0, i_13_445_68_0, i_13_445_112_0, i_13_445_120_0,
    i_13_445_123_0, i_13_445_175_0, i_13_445_214_0, i_13_445_242_0,
    i_13_445_251_0, i_13_445_259_0, i_13_445_273_0, i_13_445_277_0,
    i_13_445_278_0, i_13_445_283_0, i_13_445_311_0, i_13_445_376_0,
    i_13_445_412_0, i_13_445_454_0, i_13_445_471_0, i_13_445_521_0,
    i_13_445_609_0, i_13_445_620_0, i_13_445_800_0, i_13_445_841_0,
    i_13_445_935_0, i_13_445_980_0, i_13_445_1070_0, i_13_445_1112_0,
    i_13_445_1330_0, i_13_445_1331_0, i_13_445_1389_0, i_13_445_1394_0,
    i_13_445_1398_0, i_13_445_1410_0, i_13_445_1455_0, i_13_445_1472_0,
    i_13_445_1483_0, i_13_445_1512_0, i_13_445_1520_0, i_13_445_1573_0,
    i_13_445_1597_0, i_13_445_1598_0, i_13_445_1642_0, i_13_445_1664_0,
    i_13_445_1674_0, i_13_445_1731_0, i_13_445_1807_0, i_13_445_1835_0,
    i_13_445_1836_0, i_13_445_1945_0, i_13_445_2023_0, i_13_445_2025_0,
    i_13_445_2029_0, i_13_445_2149_0, i_13_445_2186_0, i_13_445_2200_0,
    i_13_445_2303_0, i_13_445_2433_0, i_13_445_2456_0, i_13_445_2698_0,
    i_13_445_2743_0, i_13_445_2744_0, i_13_445_2789_0, i_13_445_2883_0,
    i_13_445_2888_0, i_13_445_2937_0, i_13_445_2942_0, i_13_445_2959_0,
    i_13_445_2969_0, i_13_445_3043_0, i_13_445_3050_0, i_13_445_3077_0,
    i_13_445_3212_0, i_13_445_3238_0, i_13_445_3292_0, i_13_445_3316_0,
    i_13_445_3329_0, i_13_445_3381_0, i_13_445_3419_0, i_13_445_3454_0,
    i_13_445_3526_0, i_13_445_3533_0, i_13_445_3553_0, i_13_445_3596_0,
    i_13_445_3613_0, i_13_445_3689_0, i_13_445_3730_0, i_13_445_3762_0,
    i_13_445_3928_0, i_13_445_4066_0, i_13_445_4173_0, i_13_445_4253_0,
    i_13_445_4274_0, i_13_445_4363_0, i_13_445_4446_0, i_13_445_4503_0,
    i_13_445_4506_0, i_13_445_4517_0, i_13_445_4526_0, i_13_445_4563_0;
  output o_13_445_0_0;
  assign o_13_445_0_0 = ~((~i_13_445_3212_0 & ~i_13_445_4363_0) | (~i_13_445_2456_0 & ~i_13_445_2743_0) | (i_13_445_123_0 & i_13_445_175_0) | (~i_13_445_1483_0 & ~i_13_445_2149_0 & ~i_13_445_4517_0));
endmodule



// Benchmark "kernel_13_446" written by ABC on Sun Jul 19 10:51:35 2020

module kernel_13_446 ( 
    i_13_446_92_0, i_13_446_95_0, i_13_446_121_0, i_13_446_122_0,
    i_13_446_233_0, i_13_446_280_0, i_13_446_287_0, i_13_446_443_0,
    i_13_446_452_0, i_13_446_517_0, i_13_446_568_0, i_13_446_569_0,
    i_13_446_572_0, i_13_446_576_0, i_13_446_607_0, i_13_446_608_0,
    i_13_446_677_0, i_13_446_712_0, i_13_446_730_0, i_13_446_734_0,
    i_13_446_737_0, i_13_446_841_0, i_13_446_859_0, i_13_446_886_0,
    i_13_446_950_0, i_13_446_961_0, i_13_446_1058_0, i_13_446_1069_0,
    i_13_446_1225_0, i_13_446_1229_0, i_13_446_1327_0, i_13_446_1406_0,
    i_13_446_1448_0, i_13_446_1625_0, i_13_446_1720_0, i_13_446_1721_0,
    i_13_446_1783_0, i_13_446_1784_0, i_13_446_1787_0, i_13_446_1840_0,
    i_13_446_1855_0, i_13_446_1921_0, i_13_446_2056_0, i_13_446_2128_0,
    i_13_446_2129_0, i_13_446_2173_0, i_13_446_2206_0, i_13_446_2207_0,
    i_13_446_2359_0, i_13_446_2410_0, i_13_446_2422_0, i_13_446_2425_0,
    i_13_446_2426_0, i_13_446_2429_0, i_13_446_2458_0, i_13_446_2462_0,
    i_13_446_2465_0, i_13_446_2564_0, i_13_446_2654_0, i_13_446_2695_0,
    i_13_446_2741_0, i_13_446_2844_0, i_13_446_2941_0, i_13_446_2981_0,
    i_13_446_3015_0, i_13_446_3106_0, i_13_446_3142_0, i_13_446_3143_0,
    i_13_446_3161_0, i_13_446_3163_0, i_13_446_3164_0, i_13_446_3171_0,
    i_13_446_3214_0, i_13_446_3287_0, i_13_446_3421_0, i_13_446_3422_0,
    i_13_446_3424_0, i_13_446_3425_0, i_13_446_3428_0, i_13_446_3689_0,
    i_13_446_3769_0, i_13_446_3871_0, i_13_446_3874_0, i_13_446_3875_0,
    i_13_446_3878_0, i_13_446_3916_0, i_13_446_4006_0, i_13_446_4009_0,
    i_13_446_4010_0, i_13_446_4011_0, i_13_446_4015_0, i_13_446_4021_0,
    i_13_446_4048_0, i_13_446_4049_0, i_13_446_4066_0, i_13_446_4078_0,
    i_13_446_4318_0, i_13_446_4351_0, i_13_446_4357_0, i_13_446_4603_0,
    o_13_446_0_0  );
  input  i_13_446_92_0, i_13_446_95_0, i_13_446_121_0, i_13_446_122_0,
    i_13_446_233_0, i_13_446_280_0, i_13_446_287_0, i_13_446_443_0,
    i_13_446_452_0, i_13_446_517_0, i_13_446_568_0, i_13_446_569_0,
    i_13_446_572_0, i_13_446_576_0, i_13_446_607_0, i_13_446_608_0,
    i_13_446_677_0, i_13_446_712_0, i_13_446_730_0, i_13_446_734_0,
    i_13_446_737_0, i_13_446_841_0, i_13_446_859_0, i_13_446_886_0,
    i_13_446_950_0, i_13_446_961_0, i_13_446_1058_0, i_13_446_1069_0,
    i_13_446_1225_0, i_13_446_1229_0, i_13_446_1327_0, i_13_446_1406_0,
    i_13_446_1448_0, i_13_446_1625_0, i_13_446_1720_0, i_13_446_1721_0,
    i_13_446_1783_0, i_13_446_1784_0, i_13_446_1787_0, i_13_446_1840_0,
    i_13_446_1855_0, i_13_446_1921_0, i_13_446_2056_0, i_13_446_2128_0,
    i_13_446_2129_0, i_13_446_2173_0, i_13_446_2206_0, i_13_446_2207_0,
    i_13_446_2359_0, i_13_446_2410_0, i_13_446_2422_0, i_13_446_2425_0,
    i_13_446_2426_0, i_13_446_2429_0, i_13_446_2458_0, i_13_446_2462_0,
    i_13_446_2465_0, i_13_446_2564_0, i_13_446_2654_0, i_13_446_2695_0,
    i_13_446_2741_0, i_13_446_2844_0, i_13_446_2941_0, i_13_446_2981_0,
    i_13_446_3015_0, i_13_446_3106_0, i_13_446_3142_0, i_13_446_3143_0,
    i_13_446_3161_0, i_13_446_3163_0, i_13_446_3164_0, i_13_446_3171_0,
    i_13_446_3214_0, i_13_446_3287_0, i_13_446_3421_0, i_13_446_3422_0,
    i_13_446_3424_0, i_13_446_3425_0, i_13_446_3428_0, i_13_446_3689_0,
    i_13_446_3769_0, i_13_446_3871_0, i_13_446_3874_0, i_13_446_3875_0,
    i_13_446_3878_0, i_13_446_3916_0, i_13_446_4006_0, i_13_446_4009_0,
    i_13_446_4010_0, i_13_446_4011_0, i_13_446_4015_0, i_13_446_4021_0,
    i_13_446_4048_0, i_13_446_4049_0, i_13_446_4066_0, i_13_446_4078_0,
    i_13_446_4318_0, i_13_446_4351_0, i_13_446_4357_0, i_13_446_4603_0;
  output o_13_446_0_0;
  assign o_13_446_0_0 = ~((~i_13_446_4078_0 & (i_13_446_841_0 | (~i_13_446_3425_0 & ~i_13_446_3874_0))) | ~i_13_446_2207_0 | (~i_13_446_1625_0 & ~i_13_446_2426_0 & ~i_13_446_3875_0));
endmodule



// Benchmark "kernel_13_447" written by ABC on Sun Jul 19 10:51:35 2020

module kernel_13_447 ( 
    i_13_447_107_0, i_13_447_114_0, i_13_447_115_0, i_13_447_118_0,
    i_13_447_130_0, i_13_447_170_0, i_13_447_240_0, i_13_447_250_0,
    i_13_447_382_0, i_13_447_383_0, i_13_447_410_0, i_13_447_454_0,
    i_13_447_464_0, i_13_447_526_0, i_13_447_528_0, i_13_447_598_0,
    i_13_447_697_0, i_13_447_799_0, i_13_447_813_0, i_13_447_897_0,
    i_13_447_979_0, i_13_447_1066_0, i_13_447_1067_0, i_13_447_1085_0,
    i_13_447_1096_0, i_13_447_1300_0, i_13_447_1345_0, i_13_447_1444_0,
    i_13_447_1465_0, i_13_447_1500_0, i_13_447_1528_0, i_13_447_1544_0,
    i_13_447_1628_0, i_13_447_1636_0, i_13_447_1750_0, i_13_447_1813_0,
    i_13_447_1814_0, i_13_447_1851_0, i_13_447_1852_0, i_13_447_1867_0,
    i_13_447_1993_0, i_13_447_2005_0, i_13_447_2006_0, i_13_447_2045_0,
    i_13_447_2110_0, i_13_447_2200_0, i_13_447_2236_0, i_13_447_2435_0,
    i_13_447_2462_0, i_13_447_2464_0, i_13_447_2544_0, i_13_447_2545_0,
    i_13_447_2546_0, i_13_447_2572_0, i_13_447_2617_0, i_13_447_2618_0,
    i_13_447_2767_0, i_13_447_2825_0, i_13_447_2858_0, i_13_447_2938_0,
    i_13_447_2939_0, i_13_447_2985_0, i_13_447_3001_0, i_13_447_3014_0,
    i_13_447_3020_0, i_13_447_3112_0, i_13_447_3127_0, i_13_447_3140_0,
    i_13_447_3207_0, i_13_447_3234_0, i_13_447_3256_0, i_13_447_3262_0,
    i_13_447_3392_0, i_13_447_3418_0, i_13_447_3467_0, i_13_447_3526_0,
    i_13_447_3536_0, i_13_447_3643_0, i_13_447_3705_0, i_13_447_3722_0,
    i_13_447_3725_0, i_13_447_3733_0, i_13_447_3742_0, i_13_447_3850_0,
    i_13_447_3851_0, i_13_447_3865_0, i_13_447_3923_0, i_13_447_3963_0,
    i_13_447_4022_0, i_13_447_4063_0, i_13_447_4089_0, i_13_447_4090_0,
    i_13_447_4091_0, i_13_447_4234_0, i_13_447_4270_0, i_13_447_4271_0,
    i_13_447_4396_0, i_13_447_4533_0, i_13_447_4561_0, i_13_447_4579_0,
    o_13_447_0_0  );
  input  i_13_447_107_0, i_13_447_114_0, i_13_447_115_0, i_13_447_118_0,
    i_13_447_130_0, i_13_447_170_0, i_13_447_240_0, i_13_447_250_0,
    i_13_447_382_0, i_13_447_383_0, i_13_447_410_0, i_13_447_454_0,
    i_13_447_464_0, i_13_447_526_0, i_13_447_528_0, i_13_447_598_0,
    i_13_447_697_0, i_13_447_799_0, i_13_447_813_0, i_13_447_897_0,
    i_13_447_979_0, i_13_447_1066_0, i_13_447_1067_0, i_13_447_1085_0,
    i_13_447_1096_0, i_13_447_1300_0, i_13_447_1345_0, i_13_447_1444_0,
    i_13_447_1465_0, i_13_447_1500_0, i_13_447_1528_0, i_13_447_1544_0,
    i_13_447_1628_0, i_13_447_1636_0, i_13_447_1750_0, i_13_447_1813_0,
    i_13_447_1814_0, i_13_447_1851_0, i_13_447_1852_0, i_13_447_1867_0,
    i_13_447_1993_0, i_13_447_2005_0, i_13_447_2006_0, i_13_447_2045_0,
    i_13_447_2110_0, i_13_447_2200_0, i_13_447_2236_0, i_13_447_2435_0,
    i_13_447_2462_0, i_13_447_2464_0, i_13_447_2544_0, i_13_447_2545_0,
    i_13_447_2546_0, i_13_447_2572_0, i_13_447_2617_0, i_13_447_2618_0,
    i_13_447_2767_0, i_13_447_2825_0, i_13_447_2858_0, i_13_447_2938_0,
    i_13_447_2939_0, i_13_447_2985_0, i_13_447_3001_0, i_13_447_3014_0,
    i_13_447_3020_0, i_13_447_3112_0, i_13_447_3127_0, i_13_447_3140_0,
    i_13_447_3207_0, i_13_447_3234_0, i_13_447_3256_0, i_13_447_3262_0,
    i_13_447_3392_0, i_13_447_3418_0, i_13_447_3467_0, i_13_447_3526_0,
    i_13_447_3536_0, i_13_447_3643_0, i_13_447_3705_0, i_13_447_3722_0,
    i_13_447_3725_0, i_13_447_3733_0, i_13_447_3742_0, i_13_447_3850_0,
    i_13_447_3851_0, i_13_447_3865_0, i_13_447_3923_0, i_13_447_3963_0,
    i_13_447_4022_0, i_13_447_4063_0, i_13_447_4089_0, i_13_447_4090_0,
    i_13_447_4091_0, i_13_447_4234_0, i_13_447_4270_0, i_13_447_4271_0,
    i_13_447_4396_0, i_13_447_4533_0, i_13_447_4561_0, i_13_447_4579_0;
  output o_13_447_0_0;
  assign o_13_447_0_0 = ~((~i_13_447_2618_0 & ~i_13_447_4090_0) | (~i_13_447_115_0 & ~i_13_447_382_0) | (i_13_447_697_0 & ~i_13_447_1813_0 & ~i_13_447_4091_0) | (~i_13_447_1528_0 & ~i_13_447_1814_0 & ~i_13_447_2546_0 & ~i_13_447_3850_0) | (~i_13_447_1066_0 & ~i_13_447_1852_0 & ~i_13_447_2200_0 & ~i_13_447_2544_0));
endmodule



// Benchmark "kernel_13_448" written by ABC on Sun Jul 19 10:51:36 2020

module kernel_13_448 ( 
    i_13_448_93_0, i_13_448_106_0, i_13_448_121_0, i_13_448_183_0,
    i_13_448_184_0, i_13_448_285_0, i_13_448_322_0, i_13_448_410_0,
    i_13_448_445_0, i_13_448_466_0, i_13_448_490_0, i_13_448_537_0,
    i_13_448_571_0, i_13_448_588_0, i_13_448_645_0, i_13_448_646_0,
    i_13_448_691_0, i_13_448_697_0, i_13_448_832_0, i_13_448_845_0,
    i_13_448_898_0, i_13_448_1069_0, i_13_448_1088_0, i_13_448_1120_0,
    i_13_448_1210_0, i_13_448_1276_0, i_13_448_1303_0, i_13_448_1321_0,
    i_13_448_1329_0, i_13_448_1362_0, i_13_448_1473_0, i_13_448_1474_0,
    i_13_448_1492_0, i_13_448_1519_0, i_13_448_1520_0, i_13_448_1555_0,
    i_13_448_1789_0, i_13_448_1795_0, i_13_448_1807_0, i_13_448_1885_0,
    i_13_448_1921_0, i_13_448_1930_0, i_13_448_1933_0, i_13_448_1934_0,
    i_13_448_1960_0, i_13_448_2122_0, i_13_448_2244_0, i_13_448_2309_0,
    i_13_448_2365_0, i_13_448_2381_0, i_13_448_2473_0, i_13_448_2506_0,
    i_13_448_2695_0, i_13_448_2698_0, i_13_448_2941_0, i_13_448_2942_0,
    i_13_448_3002_0, i_13_448_3005_0, i_13_448_3022_0, i_13_448_3023_0,
    i_13_448_3064_0, i_13_448_3067_0, i_13_448_3103_0, i_13_448_3119_0,
    i_13_448_3122_0, i_13_448_3166_0, i_13_448_3210_0, i_13_448_3211_0,
    i_13_448_3346_0, i_13_448_3451_0, i_13_448_3490_0, i_13_448_3526_0,
    i_13_448_3527_0, i_13_448_3541_0, i_13_448_3544_0, i_13_448_3561_0,
    i_13_448_3631_0, i_13_448_3766_0, i_13_448_3796_0, i_13_448_3804_0,
    i_13_448_3806_0, i_13_448_3874_0, i_13_448_3910_0, i_13_448_4021_0,
    i_13_448_4048_0, i_13_448_4049_0, i_13_448_4057_0, i_13_448_4084_0,
    i_13_448_4090_0, i_13_448_4120_0, i_13_448_4273_0, i_13_448_4274_0,
    i_13_448_4353_0, i_13_448_4359_0, i_13_448_4381_0, i_13_448_4399_0,
    i_13_448_4417_0, i_13_448_4432_0, i_13_448_4593_0, i_13_448_4597_0,
    o_13_448_0_0  );
  input  i_13_448_93_0, i_13_448_106_0, i_13_448_121_0, i_13_448_183_0,
    i_13_448_184_0, i_13_448_285_0, i_13_448_322_0, i_13_448_410_0,
    i_13_448_445_0, i_13_448_466_0, i_13_448_490_0, i_13_448_537_0,
    i_13_448_571_0, i_13_448_588_0, i_13_448_645_0, i_13_448_646_0,
    i_13_448_691_0, i_13_448_697_0, i_13_448_832_0, i_13_448_845_0,
    i_13_448_898_0, i_13_448_1069_0, i_13_448_1088_0, i_13_448_1120_0,
    i_13_448_1210_0, i_13_448_1276_0, i_13_448_1303_0, i_13_448_1321_0,
    i_13_448_1329_0, i_13_448_1362_0, i_13_448_1473_0, i_13_448_1474_0,
    i_13_448_1492_0, i_13_448_1519_0, i_13_448_1520_0, i_13_448_1555_0,
    i_13_448_1789_0, i_13_448_1795_0, i_13_448_1807_0, i_13_448_1885_0,
    i_13_448_1921_0, i_13_448_1930_0, i_13_448_1933_0, i_13_448_1934_0,
    i_13_448_1960_0, i_13_448_2122_0, i_13_448_2244_0, i_13_448_2309_0,
    i_13_448_2365_0, i_13_448_2381_0, i_13_448_2473_0, i_13_448_2506_0,
    i_13_448_2695_0, i_13_448_2698_0, i_13_448_2941_0, i_13_448_2942_0,
    i_13_448_3002_0, i_13_448_3005_0, i_13_448_3022_0, i_13_448_3023_0,
    i_13_448_3064_0, i_13_448_3067_0, i_13_448_3103_0, i_13_448_3119_0,
    i_13_448_3122_0, i_13_448_3166_0, i_13_448_3210_0, i_13_448_3211_0,
    i_13_448_3346_0, i_13_448_3451_0, i_13_448_3490_0, i_13_448_3526_0,
    i_13_448_3527_0, i_13_448_3541_0, i_13_448_3544_0, i_13_448_3561_0,
    i_13_448_3631_0, i_13_448_3766_0, i_13_448_3796_0, i_13_448_3804_0,
    i_13_448_3806_0, i_13_448_3874_0, i_13_448_3910_0, i_13_448_4021_0,
    i_13_448_4048_0, i_13_448_4049_0, i_13_448_4057_0, i_13_448_4084_0,
    i_13_448_4090_0, i_13_448_4120_0, i_13_448_4273_0, i_13_448_4274_0,
    i_13_448_4353_0, i_13_448_4359_0, i_13_448_4381_0, i_13_448_4399_0,
    i_13_448_4417_0, i_13_448_4432_0, i_13_448_4593_0, i_13_448_4597_0;
  output o_13_448_0_0;
  assign o_13_448_0_0 = ~(i_13_448_697_0 | (i_13_448_1210_0 & i_13_448_4432_0) | (~i_13_448_106_0 & ~i_13_448_3103_0 & ~i_13_448_4057_0) | (~i_13_448_898_0 & ~i_13_448_3346_0 & ~i_13_448_3874_0) | (~i_13_448_537_0 & ~i_13_448_845_0 & ~i_13_448_1088_0 & ~i_13_448_4048_0));
endmodule



// Benchmark "kernel_13_449" written by ABC on Sun Jul 19 10:51:37 2020

module kernel_13_449 ( 
    i_13_449_41_0, i_13_449_62_0, i_13_449_74_0, i_13_449_77_0,
    i_13_449_137_0, i_13_449_167_0, i_13_449_227_0, i_13_449_274_0,
    i_13_449_337_0, i_13_449_537_0, i_13_449_571_0, i_13_449_582_0,
    i_13_449_641_0, i_13_449_681_0, i_13_449_689_0, i_13_449_690_0,
    i_13_449_694_0, i_13_449_695_0, i_13_449_697_0, i_13_449_814_0,
    i_13_449_820_0, i_13_449_821_0, i_13_449_824_0, i_13_449_825_0,
    i_13_449_887_0, i_13_449_1066_0, i_13_449_1067_0, i_13_449_1068_0,
    i_13_449_1211_0, i_13_449_1220_0, i_13_449_1271_0, i_13_449_1381_0,
    i_13_449_1388_0, i_13_449_1423_0, i_13_449_1444_0, i_13_449_1490_0,
    i_13_449_1594_0, i_13_449_1640_0, i_13_449_1670_0, i_13_449_1712_0,
    i_13_449_1793_0, i_13_449_1882_0, i_13_449_1883_0, i_13_449_1885_0,
    i_13_449_1886_0, i_13_449_1889_0, i_13_449_2364_0, i_13_449_2470_0,
    i_13_449_2549_0, i_13_449_2552_0, i_13_449_2611_0, i_13_449_2647_0,
    i_13_449_2651_0, i_13_449_2845_0, i_13_449_2848_0, i_13_449_2873_0,
    i_13_449_2885_0, i_13_449_2983_0, i_13_449_3011_0, i_13_449_3028_0,
    i_13_449_3109_0, i_13_449_3127_0, i_13_449_3173_0, i_13_449_3208_0,
    i_13_449_3269_0, i_13_449_3311_0, i_13_449_3343_0, i_13_449_3367_0,
    i_13_449_3376_0, i_13_449_3382_0, i_13_449_3383_0, i_13_449_3397_0,
    i_13_449_3415_0, i_13_449_3449_0, i_13_449_3487_0, i_13_449_3502_0,
    i_13_449_3503_0, i_13_449_3505_0, i_13_449_3728_0, i_13_449_3736_0,
    i_13_449_3740_0, i_13_449_3791_0, i_13_449_3836_0, i_13_449_3847_0,
    i_13_449_3871_0, i_13_449_4063_0, i_13_449_4064_0, i_13_449_4079_0,
    i_13_449_4187_0, i_13_449_4253_0, i_13_449_4262_0, i_13_449_4270_0,
    i_13_449_4295_0, i_13_449_4339_0, i_13_449_4342_0, i_13_449_4351_0,
    i_13_449_4441_0, i_13_449_4498_0, i_13_449_4591_0, i_13_449_4592_0,
    o_13_449_0_0  );
  input  i_13_449_41_0, i_13_449_62_0, i_13_449_74_0, i_13_449_77_0,
    i_13_449_137_0, i_13_449_167_0, i_13_449_227_0, i_13_449_274_0,
    i_13_449_337_0, i_13_449_537_0, i_13_449_571_0, i_13_449_582_0,
    i_13_449_641_0, i_13_449_681_0, i_13_449_689_0, i_13_449_690_0,
    i_13_449_694_0, i_13_449_695_0, i_13_449_697_0, i_13_449_814_0,
    i_13_449_820_0, i_13_449_821_0, i_13_449_824_0, i_13_449_825_0,
    i_13_449_887_0, i_13_449_1066_0, i_13_449_1067_0, i_13_449_1068_0,
    i_13_449_1211_0, i_13_449_1220_0, i_13_449_1271_0, i_13_449_1381_0,
    i_13_449_1388_0, i_13_449_1423_0, i_13_449_1444_0, i_13_449_1490_0,
    i_13_449_1594_0, i_13_449_1640_0, i_13_449_1670_0, i_13_449_1712_0,
    i_13_449_1793_0, i_13_449_1882_0, i_13_449_1883_0, i_13_449_1885_0,
    i_13_449_1886_0, i_13_449_1889_0, i_13_449_2364_0, i_13_449_2470_0,
    i_13_449_2549_0, i_13_449_2552_0, i_13_449_2611_0, i_13_449_2647_0,
    i_13_449_2651_0, i_13_449_2845_0, i_13_449_2848_0, i_13_449_2873_0,
    i_13_449_2885_0, i_13_449_2983_0, i_13_449_3011_0, i_13_449_3028_0,
    i_13_449_3109_0, i_13_449_3127_0, i_13_449_3173_0, i_13_449_3208_0,
    i_13_449_3269_0, i_13_449_3311_0, i_13_449_3343_0, i_13_449_3367_0,
    i_13_449_3376_0, i_13_449_3382_0, i_13_449_3383_0, i_13_449_3397_0,
    i_13_449_3415_0, i_13_449_3449_0, i_13_449_3487_0, i_13_449_3502_0,
    i_13_449_3503_0, i_13_449_3505_0, i_13_449_3728_0, i_13_449_3736_0,
    i_13_449_3740_0, i_13_449_3791_0, i_13_449_3836_0, i_13_449_3847_0,
    i_13_449_3871_0, i_13_449_4063_0, i_13_449_4064_0, i_13_449_4079_0,
    i_13_449_4187_0, i_13_449_4253_0, i_13_449_4262_0, i_13_449_4270_0,
    i_13_449_4295_0, i_13_449_4339_0, i_13_449_4342_0, i_13_449_4351_0,
    i_13_449_4441_0, i_13_449_4498_0, i_13_449_4591_0, i_13_449_4592_0;
  output o_13_449_0_0;
  assign o_13_449_0_0 = ~((~i_13_449_1490_0 & ((~i_13_449_824_0 & ~i_13_449_3487_0 & ~i_13_449_3736_0) | (i_13_449_3208_0 & i_13_449_3847_0))) | (~i_13_449_824_0 & ((~i_13_449_887_0 & ~i_13_449_3502_0) | (~i_13_449_820_0 & ~i_13_449_3740_0))) | (~i_13_449_1793_0 & ~i_13_449_1883_0 & i_13_449_3397_0 & ~i_13_449_3503_0) | (~i_13_449_1886_0 & ~i_13_449_2848_0 & ~i_13_449_3728_0 & i_13_449_3847_0 & ~i_13_449_4262_0) | (i_13_449_3871_0 & ~i_13_449_4351_0));
endmodule



// Benchmark "kernel_13_450" written by ABC on Sun Jul 19 10:51:38 2020

module kernel_13_450 ( 
    i_13_450_60_0, i_13_450_67_0, i_13_450_229_0, i_13_450_418_0,
    i_13_450_463_0, i_13_450_526_0, i_13_450_554_0, i_13_450_608_0,
    i_13_450_628_0, i_13_450_658_0, i_13_450_660_0, i_13_450_661_0,
    i_13_450_733_0, i_13_450_831_0, i_13_450_888_0, i_13_450_889_0,
    i_13_450_959_0, i_13_450_988_0, i_13_450_1071_0, i_13_450_1078_0,
    i_13_450_1087_0, i_13_450_1099_0, i_13_450_1108_0, i_13_450_1112_0,
    i_13_450_1120_0, i_13_450_1143_0, i_13_450_1279_0, i_13_450_1300_0,
    i_13_450_1330_0, i_13_450_1345_0, i_13_450_1466_0, i_13_450_1476_0,
    i_13_450_1516_0, i_13_450_1660_0, i_13_450_1678_0, i_13_450_1681_0,
    i_13_450_1744_0, i_13_450_2002_0, i_13_450_2019_0, i_13_450_2020_0,
    i_13_450_2021_0, i_13_450_2022_0, i_13_450_2023_0, i_13_450_2024_0,
    i_13_450_2077_0, i_13_450_2097_0, i_13_450_2137_0, i_13_450_2425_0,
    i_13_450_2453_0, i_13_450_2466_0, i_13_450_2470_0, i_13_450_2511_0,
    i_13_450_2614_0, i_13_450_2708_0, i_13_450_2723_0, i_13_450_2740_0,
    i_13_450_2741_0, i_13_450_2857_0, i_13_450_2935_0, i_13_450_2998_0,
    i_13_450_3004_0, i_13_450_3056_0, i_13_450_3089_0, i_13_450_3152_0,
    i_13_450_3272_0, i_13_450_3352_0, i_13_450_3483_0, i_13_450_3484_0,
    i_13_450_3490_0, i_13_450_3550_0, i_13_450_3553_0, i_13_450_3568_0,
    i_13_450_3621_0, i_13_450_3730_0, i_13_450_3766_0, i_13_450_3823_0,
    i_13_450_3861_0, i_13_450_3864_0, i_13_450_3866_0, i_13_450_3989_0,
    i_13_450_4027_0, i_13_450_4048_0, i_13_450_4051_0, i_13_450_4054_0,
    i_13_450_4160_0, i_13_450_4162_0, i_13_450_4163_0, i_13_450_4252_0,
    i_13_450_4253_0, i_13_450_4369_0, i_13_450_4370_0, i_13_450_4377_0,
    i_13_450_4388_0, i_13_450_4394_0, i_13_450_4396_0, i_13_450_4431_0,
    i_13_450_4517_0, i_13_450_4560_0, i_13_450_4603_0, i_13_450_4604_0,
    o_13_450_0_0  );
  input  i_13_450_60_0, i_13_450_67_0, i_13_450_229_0, i_13_450_418_0,
    i_13_450_463_0, i_13_450_526_0, i_13_450_554_0, i_13_450_608_0,
    i_13_450_628_0, i_13_450_658_0, i_13_450_660_0, i_13_450_661_0,
    i_13_450_733_0, i_13_450_831_0, i_13_450_888_0, i_13_450_889_0,
    i_13_450_959_0, i_13_450_988_0, i_13_450_1071_0, i_13_450_1078_0,
    i_13_450_1087_0, i_13_450_1099_0, i_13_450_1108_0, i_13_450_1112_0,
    i_13_450_1120_0, i_13_450_1143_0, i_13_450_1279_0, i_13_450_1300_0,
    i_13_450_1330_0, i_13_450_1345_0, i_13_450_1466_0, i_13_450_1476_0,
    i_13_450_1516_0, i_13_450_1660_0, i_13_450_1678_0, i_13_450_1681_0,
    i_13_450_1744_0, i_13_450_2002_0, i_13_450_2019_0, i_13_450_2020_0,
    i_13_450_2021_0, i_13_450_2022_0, i_13_450_2023_0, i_13_450_2024_0,
    i_13_450_2077_0, i_13_450_2097_0, i_13_450_2137_0, i_13_450_2425_0,
    i_13_450_2453_0, i_13_450_2466_0, i_13_450_2470_0, i_13_450_2511_0,
    i_13_450_2614_0, i_13_450_2708_0, i_13_450_2723_0, i_13_450_2740_0,
    i_13_450_2741_0, i_13_450_2857_0, i_13_450_2935_0, i_13_450_2998_0,
    i_13_450_3004_0, i_13_450_3056_0, i_13_450_3089_0, i_13_450_3152_0,
    i_13_450_3272_0, i_13_450_3352_0, i_13_450_3483_0, i_13_450_3484_0,
    i_13_450_3490_0, i_13_450_3550_0, i_13_450_3553_0, i_13_450_3568_0,
    i_13_450_3621_0, i_13_450_3730_0, i_13_450_3766_0, i_13_450_3823_0,
    i_13_450_3861_0, i_13_450_3864_0, i_13_450_3866_0, i_13_450_3989_0,
    i_13_450_4027_0, i_13_450_4048_0, i_13_450_4051_0, i_13_450_4054_0,
    i_13_450_4160_0, i_13_450_4162_0, i_13_450_4163_0, i_13_450_4252_0,
    i_13_450_4253_0, i_13_450_4369_0, i_13_450_4370_0, i_13_450_4377_0,
    i_13_450_4388_0, i_13_450_4394_0, i_13_450_4396_0, i_13_450_4431_0,
    i_13_450_4517_0, i_13_450_4560_0, i_13_450_4603_0, i_13_450_4604_0;
  output o_13_450_0_0;
  assign o_13_450_0_0 = ~((~i_13_450_1330_0 & ((i_13_450_526_0 & ~i_13_450_2740_0) | (~i_13_450_60_0 & ~i_13_450_831_0 & ~i_13_450_3866_0))) | ~i_13_450_2020_0 | (i_13_450_229_0 & ~i_13_450_2019_0 & ~i_13_450_2740_0 & ~i_13_450_3550_0) | (~i_13_450_2723_0 & ~i_13_450_3864_0) | (i_13_450_1345_0 & ~i_13_450_2741_0 & ~i_13_450_4370_0) | (~i_13_450_4252_0 & i_13_450_4396_0));
endmodule



// Benchmark "kernel_13_451" written by ABC on Sun Jul 19 10:51:39 2020

module kernel_13_451 ( 
    i_13_451_71_0, i_13_451_94_0, i_13_451_140_0, i_13_451_179_0,
    i_13_451_259_0, i_13_451_266_0, i_13_451_287_0, i_13_451_327_0,
    i_13_451_328_0, i_13_451_329_0, i_13_451_418_0, i_13_451_468_0,
    i_13_451_494_0, i_13_451_562_0, i_13_451_563_0, i_13_451_607_0,
    i_13_451_628_0, i_13_451_667_0, i_13_451_670_0, i_13_451_671_0,
    i_13_451_683_0, i_13_451_700_0, i_13_451_701_0, i_13_451_891_0,
    i_13_451_943_0, i_13_451_1021_0, i_13_451_1024_0, i_13_451_1078_0,
    i_13_451_1079_0, i_13_451_1314_0, i_13_451_1327_0, i_13_451_1403_0,
    i_13_451_1430_0, i_13_451_1444_0, i_13_451_1447_0, i_13_451_1479_0,
    i_13_451_1480_0, i_13_451_1484_0, i_13_451_1687_0, i_13_451_1780_0,
    i_13_451_1781_0, i_13_451_1789_0, i_13_451_1840_0, i_13_451_1885_0,
    i_13_451_1889_0, i_13_451_1906_0, i_13_451_1923_0, i_13_451_1935_0,
    i_13_451_2022_0, i_13_451_2059_0, i_13_451_2124_0, i_13_451_2125_0,
    i_13_451_2173_0, i_13_451_2197_0, i_13_451_2201_0, i_13_451_2245_0,
    i_13_451_2344_0, i_13_451_2384_0, i_13_451_2434_0, i_13_451_2561_0,
    i_13_451_2617_0, i_13_451_2618_0, i_13_451_2629_0, i_13_451_2746_0,
    i_13_451_2852_0, i_13_451_2875_0, i_13_451_2898_0, i_13_451_2902_0,
    i_13_451_2967_0, i_13_451_3043_0, i_13_451_3100_0, i_13_451_3175_0,
    i_13_451_3244_0, i_13_451_3381_0, i_13_451_3415_0, i_13_451_3429_0,
    i_13_451_3455_0, i_13_451_3460_0, i_13_451_3464_0, i_13_451_3482_0,
    i_13_451_3507_0, i_13_451_3535_0, i_13_451_3536_0, i_13_451_3596_0,
    i_13_451_3701_0, i_13_451_3731_0, i_13_451_3869_0, i_13_451_3911_0,
    i_13_451_3920_0, i_13_451_4100_0, i_13_451_4257_0, i_13_451_4342_0,
    i_13_451_4346_0, i_13_451_4350_0, i_13_451_4351_0, i_13_451_4354_0,
    i_13_451_4396_0, i_13_451_4451_0, i_13_451_4522_0, i_13_451_4606_0,
    o_13_451_0_0  );
  input  i_13_451_71_0, i_13_451_94_0, i_13_451_140_0, i_13_451_179_0,
    i_13_451_259_0, i_13_451_266_0, i_13_451_287_0, i_13_451_327_0,
    i_13_451_328_0, i_13_451_329_0, i_13_451_418_0, i_13_451_468_0,
    i_13_451_494_0, i_13_451_562_0, i_13_451_563_0, i_13_451_607_0,
    i_13_451_628_0, i_13_451_667_0, i_13_451_670_0, i_13_451_671_0,
    i_13_451_683_0, i_13_451_700_0, i_13_451_701_0, i_13_451_891_0,
    i_13_451_943_0, i_13_451_1021_0, i_13_451_1024_0, i_13_451_1078_0,
    i_13_451_1079_0, i_13_451_1314_0, i_13_451_1327_0, i_13_451_1403_0,
    i_13_451_1430_0, i_13_451_1444_0, i_13_451_1447_0, i_13_451_1479_0,
    i_13_451_1480_0, i_13_451_1484_0, i_13_451_1687_0, i_13_451_1780_0,
    i_13_451_1781_0, i_13_451_1789_0, i_13_451_1840_0, i_13_451_1885_0,
    i_13_451_1889_0, i_13_451_1906_0, i_13_451_1923_0, i_13_451_1935_0,
    i_13_451_2022_0, i_13_451_2059_0, i_13_451_2124_0, i_13_451_2125_0,
    i_13_451_2173_0, i_13_451_2197_0, i_13_451_2201_0, i_13_451_2245_0,
    i_13_451_2344_0, i_13_451_2384_0, i_13_451_2434_0, i_13_451_2561_0,
    i_13_451_2617_0, i_13_451_2618_0, i_13_451_2629_0, i_13_451_2746_0,
    i_13_451_2852_0, i_13_451_2875_0, i_13_451_2898_0, i_13_451_2902_0,
    i_13_451_2967_0, i_13_451_3043_0, i_13_451_3100_0, i_13_451_3175_0,
    i_13_451_3244_0, i_13_451_3381_0, i_13_451_3415_0, i_13_451_3429_0,
    i_13_451_3455_0, i_13_451_3460_0, i_13_451_3464_0, i_13_451_3482_0,
    i_13_451_3507_0, i_13_451_3535_0, i_13_451_3536_0, i_13_451_3596_0,
    i_13_451_3701_0, i_13_451_3731_0, i_13_451_3869_0, i_13_451_3911_0,
    i_13_451_3920_0, i_13_451_4100_0, i_13_451_4257_0, i_13_451_4342_0,
    i_13_451_4346_0, i_13_451_4350_0, i_13_451_4351_0, i_13_451_4354_0,
    i_13_451_4396_0, i_13_451_4451_0, i_13_451_4522_0, i_13_451_4606_0;
  output o_13_451_0_0;
  assign o_13_451_0_0 = ~((~i_13_451_2618_0 & ~i_13_451_3535_0) | (~i_13_451_700_0 & ~i_13_451_3911_0 & ~i_13_451_4396_0) | (~i_13_451_328_0 & i_13_451_2434_0 & ~i_13_451_3464_0) | (~i_13_451_1479_0 & ~i_13_451_1781_0 & i_13_451_3460_0) | (~i_13_451_943_0 & i_13_451_1021_0 & i_13_451_2022_0));
endmodule



// Benchmark "kernel_13_452" written by ABC on Sun Jul 19 10:51:39 2020

module kernel_13_452 ( 
    i_13_452_7_0, i_13_452_33_0, i_13_452_34_0, i_13_452_35_0,
    i_13_452_41_0, i_13_452_109_0, i_13_452_160_0, i_13_452_188_0,
    i_13_452_232_0, i_13_452_374_0, i_13_452_385_0, i_13_452_447_0,
    i_13_452_538_0, i_13_452_572_0, i_13_452_669_0, i_13_452_763_0,
    i_13_452_860_0, i_13_452_942_0, i_13_452_1075_0, i_13_452_1088_0,
    i_13_452_1215_0, i_13_452_1218_0, i_13_452_1219_0, i_13_452_1302_0,
    i_13_452_1348_0, i_13_452_1398_0, i_13_452_1473_0, i_13_452_1474_0,
    i_13_452_1475_0, i_13_452_1492_0, i_13_452_1545_0, i_13_452_1599_0,
    i_13_452_1636_0, i_13_452_1724_0, i_13_452_1789_0, i_13_452_1795_0,
    i_13_452_1992_0, i_13_452_1995_0, i_13_452_2002_0, i_13_452_2010_0,
    i_13_452_2046_0, i_13_452_2194_0, i_13_452_2209_0, i_13_452_2231_0,
    i_13_452_2242_0, i_13_452_2364_0, i_13_452_2365_0, i_13_452_2424_0,
    i_13_452_2426_0, i_13_452_2455_0, i_13_452_2472_0, i_13_452_2501_0,
    i_13_452_2532_0, i_13_452_2679_0, i_13_452_2904_0, i_13_452_2938_0,
    i_13_452_2958_0, i_13_452_3003_0, i_13_452_3004_0, i_13_452_3022_0,
    i_13_452_3023_0, i_13_452_3028_0, i_13_452_3066_0, i_13_452_3067_0,
    i_13_452_3112_0, i_13_452_3148_0, i_13_452_3163_0, i_13_452_3207_0,
    i_13_452_3210_0, i_13_452_3229_0, i_13_452_3234_0, i_13_452_3289_0,
    i_13_452_3308_0, i_13_452_3346_0, i_13_452_3382_0, i_13_452_3390_0,
    i_13_452_3423_0, i_13_452_3426_0, i_13_452_3490_0, i_13_452_3544_0,
    i_13_452_3580_0, i_13_452_3639_0, i_13_452_3648_0, i_13_452_3702_0,
    i_13_452_3796_0, i_13_452_3847_0, i_13_452_3873_0, i_13_452_3874_0,
    i_13_452_4008_0, i_13_452_4009_0, i_13_452_4035_0, i_13_452_4057_0,
    i_13_452_4120_0, i_13_452_4208_0, i_13_452_4354_0, i_13_452_4355_0,
    i_13_452_4399_0, i_13_452_4417_0, i_13_452_4418_0, i_13_452_4603_0,
    o_13_452_0_0  );
  input  i_13_452_7_0, i_13_452_33_0, i_13_452_34_0, i_13_452_35_0,
    i_13_452_41_0, i_13_452_109_0, i_13_452_160_0, i_13_452_188_0,
    i_13_452_232_0, i_13_452_374_0, i_13_452_385_0, i_13_452_447_0,
    i_13_452_538_0, i_13_452_572_0, i_13_452_669_0, i_13_452_763_0,
    i_13_452_860_0, i_13_452_942_0, i_13_452_1075_0, i_13_452_1088_0,
    i_13_452_1215_0, i_13_452_1218_0, i_13_452_1219_0, i_13_452_1302_0,
    i_13_452_1348_0, i_13_452_1398_0, i_13_452_1473_0, i_13_452_1474_0,
    i_13_452_1475_0, i_13_452_1492_0, i_13_452_1545_0, i_13_452_1599_0,
    i_13_452_1636_0, i_13_452_1724_0, i_13_452_1789_0, i_13_452_1795_0,
    i_13_452_1992_0, i_13_452_1995_0, i_13_452_2002_0, i_13_452_2010_0,
    i_13_452_2046_0, i_13_452_2194_0, i_13_452_2209_0, i_13_452_2231_0,
    i_13_452_2242_0, i_13_452_2364_0, i_13_452_2365_0, i_13_452_2424_0,
    i_13_452_2426_0, i_13_452_2455_0, i_13_452_2472_0, i_13_452_2501_0,
    i_13_452_2532_0, i_13_452_2679_0, i_13_452_2904_0, i_13_452_2938_0,
    i_13_452_2958_0, i_13_452_3003_0, i_13_452_3004_0, i_13_452_3022_0,
    i_13_452_3023_0, i_13_452_3028_0, i_13_452_3066_0, i_13_452_3067_0,
    i_13_452_3112_0, i_13_452_3148_0, i_13_452_3163_0, i_13_452_3207_0,
    i_13_452_3210_0, i_13_452_3229_0, i_13_452_3234_0, i_13_452_3289_0,
    i_13_452_3308_0, i_13_452_3346_0, i_13_452_3382_0, i_13_452_3390_0,
    i_13_452_3423_0, i_13_452_3426_0, i_13_452_3490_0, i_13_452_3544_0,
    i_13_452_3580_0, i_13_452_3639_0, i_13_452_3648_0, i_13_452_3702_0,
    i_13_452_3796_0, i_13_452_3847_0, i_13_452_3873_0, i_13_452_3874_0,
    i_13_452_4008_0, i_13_452_4009_0, i_13_452_4035_0, i_13_452_4057_0,
    i_13_452_4120_0, i_13_452_4208_0, i_13_452_4354_0, i_13_452_4355_0,
    i_13_452_4399_0, i_13_452_4417_0, i_13_452_4418_0, i_13_452_4603_0;
  output o_13_452_0_0;
  assign o_13_452_0_0 = ~((~i_13_452_3067_0 & ~i_13_452_4008_0) | (~i_13_452_385_0 & i_13_452_3289_0) | (~i_13_452_1218_0 & ~i_13_452_2426_0 & ~i_13_452_3346_0));
endmodule



// Benchmark "kernel_13_453" written by ABC on Sun Jul 19 10:51:40 2020

module kernel_13_453 ( 
    i_13_453_94_0, i_13_453_103_0, i_13_453_140_0, i_13_453_166_0,
    i_13_453_431_0, i_13_453_536_0, i_13_453_574_0, i_13_453_644_0,
    i_13_453_647_0, i_13_453_668_0, i_13_453_686_0, i_13_453_691_0,
    i_13_453_694_0, i_13_453_697_0, i_13_453_698_0, i_13_453_700_0,
    i_13_453_707_0, i_13_453_823_0, i_13_453_827_0, i_13_453_977_0,
    i_13_453_1033_0, i_13_453_1079_0, i_13_453_1115_0, i_13_453_1118_0,
    i_13_453_1121_0, i_13_453_1124_0, i_13_453_1138_0, i_13_453_1249_0,
    i_13_453_1277_0, i_13_453_1318_0, i_13_453_1319_0, i_13_453_1333_0,
    i_13_453_1388_0, i_13_453_1391_0, i_13_453_1447_0, i_13_453_1462_0,
    i_13_453_1465_0, i_13_453_1468_0, i_13_453_1469_0, i_13_453_1483_0,
    i_13_453_1484_0, i_13_453_1534_0, i_13_453_1586_0, i_13_453_1597_0,
    i_13_453_1711_0, i_13_453_1778_0, i_13_453_1781_0, i_13_453_1828_0,
    i_13_453_1849_0, i_13_453_1850_0, i_13_453_1886_0, i_13_453_1888_0,
    i_13_453_1889_0, i_13_453_1945_0, i_13_453_2102_0, i_13_453_2150_0,
    i_13_453_2206_0, i_13_453_2425_0, i_13_453_2567_0, i_13_453_2650_0,
    i_13_453_2651_0, i_13_453_2654_0, i_13_453_2689_0, i_13_453_2848_0,
    i_13_453_2849_0, i_13_453_2853_0, i_13_453_2875_0, i_13_453_2876_0,
    i_13_453_2888_0, i_13_453_3089_0, i_13_453_3217_0, i_13_453_3235_0,
    i_13_453_3244_0, i_13_453_3245_0, i_13_453_3299_0, i_13_453_3356_0,
    i_13_453_3398_0, i_13_453_3406_0, i_13_453_3448_0, i_13_453_3449_0,
    i_13_453_3501_0, i_13_453_3506_0, i_13_453_3526_0, i_13_453_3785_0,
    i_13_453_3794_0, i_13_453_3847_0, i_13_453_3854_0, i_13_453_3863_0,
    i_13_453_3982_0, i_13_453_3995_0, i_13_453_4090_0, i_13_453_4100_0,
    i_13_453_4187_0, i_13_453_4189_0, i_13_453_4190_0, i_13_453_4310_0,
    i_13_453_4364_0, i_13_453_4391_0, i_13_453_4481_0, i_13_453_4598_0,
    o_13_453_0_0  );
  input  i_13_453_94_0, i_13_453_103_0, i_13_453_140_0, i_13_453_166_0,
    i_13_453_431_0, i_13_453_536_0, i_13_453_574_0, i_13_453_644_0,
    i_13_453_647_0, i_13_453_668_0, i_13_453_686_0, i_13_453_691_0,
    i_13_453_694_0, i_13_453_697_0, i_13_453_698_0, i_13_453_700_0,
    i_13_453_707_0, i_13_453_823_0, i_13_453_827_0, i_13_453_977_0,
    i_13_453_1033_0, i_13_453_1079_0, i_13_453_1115_0, i_13_453_1118_0,
    i_13_453_1121_0, i_13_453_1124_0, i_13_453_1138_0, i_13_453_1249_0,
    i_13_453_1277_0, i_13_453_1318_0, i_13_453_1319_0, i_13_453_1333_0,
    i_13_453_1388_0, i_13_453_1391_0, i_13_453_1447_0, i_13_453_1462_0,
    i_13_453_1465_0, i_13_453_1468_0, i_13_453_1469_0, i_13_453_1483_0,
    i_13_453_1484_0, i_13_453_1534_0, i_13_453_1586_0, i_13_453_1597_0,
    i_13_453_1711_0, i_13_453_1778_0, i_13_453_1781_0, i_13_453_1828_0,
    i_13_453_1849_0, i_13_453_1850_0, i_13_453_1886_0, i_13_453_1888_0,
    i_13_453_1889_0, i_13_453_1945_0, i_13_453_2102_0, i_13_453_2150_0,
    i_13_453_2206_0, i_13_453_2425_0, i_13_453_2567_0, i_13_453_2650_0,
    i_13_453_2651_0, i_13_453_2654_0, i_13_453_2689_0, i_13_453_2848_0,
    i_13_453_2849_0, i_13_453_2853_0, i_13_453_2875_0, i_13_453_2876_0,
    i_13_453_2888_0, i_13_453_3089_0, i_13_453_3217_0, i_13_453_3235_0,
    i_13_453_3244_0, i_13_453_3245_0, i_13_453_3299_0, i_13_453_3356_0,
    i_13_453_3398_0, i_13_453_3406_0, i_13_453_3448_0, i_13_453_3449_0,
    i_13_453_3501_0, i_13_453_3506_0, i_13_453_3526_0, i_13_453_3785_0,
    i_13_453_3794_0, i_13_453_3847_0, i_13_453_3854_0, i_13_453_3863_0,
    i_13_453_3982_0, i_13_453_3995_0, i_13_453_4090_0, i_13_453_4100_0,
    i_13_453_4187_0, i_13_453_4189_0, i_13_453_4190_0, i_13_453_4310_0,
    i_13_453_4364_0, i_13_453_4391_0, i_13_453_4481_0, i_13_453_4598_0;
  output o_13_453_0_0;
  assign o_13_453_0_0 = ~((~i_13_453_140_0 & ~i_13_453_4189_0) | (~i_13_453_691_0 & ~i_13_453_1889_0 & ~i_13_453_3448_0) | (~i_13_453_1124_0 & ~i_13_453_1277_0 & ~i_13_453_2849_0) | (~i_13_453_1483_0 & ~i_13_453_1484_0 & ~i_13_453_1888_0 & ~i_13_453_1945_0));
endmodule



// Benchmark "kernel_13_454" written by ABC on Sun Jul 19 10:51:41 2020

module kernel_13_454 ( 
    i_13_454_44_0, i_13_454_49_0, i_13_454_56_0, i_13_454_70_0,
    i_13_454_78_0, i_13_454_172_0, i_13_454_176_0, i_13_454_177_0,
    i_13_454_282_0, i_13_454_317_0, i_13_454_321_0, i_13_454_447_0,
    i_13_454_448_0, i_13_454_457_0, i_13_454_461_0, i_13_454_525_0,
    i_13_454_555_0, i_13_454_568_0, i_13_454_645_0, i_13_454_651_0,
    i_13_454_670_0, i_13_454_673_0, i_13_454_679_0, i_13_454_681_0,
    i_13_454_682_0, i_13_454_688_0, i_13_454_740_0, i_13_454_757_0,
    i_13_454_994_0, i_13_454_1104_0, i_13_454_1150_0, i_13_454_1275_0,
    i_13_454_1276_0, i_13_454_1401_0, i_13_454_1402_0, i_13_454_1426_0,
    i_13_454_1510_0, i_13_454_1514_0, i_13_454_1548_0, i_13_454_1567_0,
    i_13_454_1599_0, i_13_454_1633_0, i_13_454_1645_0, i_13_454_1663_0,
    i_13_454_1725_0, i_13_454_1734_0, i_13_454_1798_0, i_13_454_1920_0,
    i_13_454_1945_0, i_13_454_1946_0, i_13_454_1948_0, i_13_454_1996_0,
    i_13_454_2029_0, i_13_454_2032_0, i_13_454_2191_0, i_13_454_2263_0,
    i_13_454_2265_0, i_13_454_2266_0, i_13_454_2407_0, i_13_454_2461_0,
    i_13_454_2472_0, i_13_454_2545_0, i_13_454_2587_0, i_13_454_2677_0,
    i_13_454_2680_0, i_13_454_2695_0, i_13_454_2697_0, i_13_454_2742_0,
    i_13_454_2748_0, i_13_454_2901_0, i_13_454_2902_0, i_13_454_2905_0,
    i_13_454_2922_0, i_13_454_2923_0, i_13_454_2940_0, i_13_454_2981_0,
    i_13_454_3030_0, i_13_454_3111_0, i_13_454_3269_0, i_13_454_3273_0,
    i_13_454_3367_0, i_13_454_3418_0, i_13_454_3525_0, i_13_454_3561_0,
    i_13_454_3592_0, i_13_454_3651_0, i_13_454_3730_0, i_13_454_3732_0,
    i_13_454_3787_0, i_13_454_3928_0, i_13_454_3940_0, i_13_454_3992_0,
    i_13_454_3993_0, i_13_454_3994_0, i_13_454_4053_0, i_13_454_4251_0,
    i_13_454_4308_0, i_13_454_4323_0, i_13_454_4566_0, i_13_454_4603_0,
    o_13_454_0_0  );
  input  i_13_454_44_0, i_13_454_49_0, i_13_454_56_0, i_13_454_70_0,
    i_13_454_78_0, i_13_454_172_0, i_13_454_176_0, i_13_454_177_0,
    i_13_454_282_0, i_13_454_317_0, i_13_454_321_0, i_13_454_447_0,
    i_13_454_448_0, i_13_454_457_0, i_13_454_461_0, i_13_454_525_0,
    i_13_454_555_0, i_13_454_568_0, i_13_454_645_0, i_13_454_651_0,
    i_13_454_670_0, i_13_454_673_0, i_13_454_679_0, i_13_454_681_0,
    i_13_454_682_0, i_13_454_688_0, i_13_454_740_0, i_13_454_757_0,
    i_13_454_994_0, i_13_454_1104_0, i_13_454_1150_0, i_13_454_1275_0,
    i_13_454_1276_0, i_13_454_1401_0, i_13_454_1402_0, i_13_454_1426_0,
    i_13_454_1510_0, i_13_454_1514_0, i_13_454_1548_0, i_13_454_1567_0,
    i_13_454_1599_0, i_13_454_1633_0, i_13_454_1645_0, i_13_454_1663_0,
    i_13_454_1725_0, i_13_454_1734_0, i_13_454_1798_0, i_13_454_1920_0,
    i_13_454_1945_0, i_13_454_1946_0, i_13_454_1948_0, i_13_454_1996_0,
    i_13_454_2029_0, i_13_454_2032_0, i_13_454_2191_0, i_13_454_2263_0,
    i_13_454_2265_0, i_13_454_2266_0, i_13_454_2407_0, i_13_454_2461_0,
    i_13_454_2472_0, i_13_454_2545_0, i_13_454_2587_0, i_13_454_2677_0,
    i_13_454_2680_0, i_13_454_2695_0, i_13_454_2697_0, i_13_454_2742_0,
    i_13_454_2748_0, i_13_454_2901_0, i_13_454_2902_0, i_13_454_2905_0,
    i_13_454_2922_0, i_13_454_2923_0, i_13_454_2940_0, i_13_454_2981_0,
    i_13_454_3030_0, i_13_454_3111_0, i_13_454_3269_0, i_13_454_3273_0,
    i_13_454_3367_0, i_13_454_3418_0, i_13_454_3525_0, i_13_454_3561_0,
    i_13_454_3592_0, i_13_454_3651_0, i_13_454_3730_0, i_13_454_3732_0,
    i_13_454_3787_0, i_13_454_3928_0, i_13_454_3940_0, i_13_454_3992_0,
    i_13_454_3993_0, i_13_454_3994_0, i_13_454_4053_0, i_13_454_4251_0,
    i_13_454_4308_0, i_13_454_4323_0, i_13_454_4566_0, i_13_454_4603_0;
  output o_13_454_0_0;
  assign o_13_454_0_0 = ~((~i_13_454_3993_0 & ((~i_13_454_282_0 & ~i_13_454_321_0) | (~i_13_454_70_0 & ~i_13_454_2697_0))) | (~i_13_454_1734_0 & i_13_454_3730_0));
endmodule



// Benchmark "kernel_13_455" written by ABC on Sun Jul 19 10:51:42 2020

module kernel_13_455 ( 
    i_13_455_2_0, i_13_455_156_0, i_13_455_164_0, i_13_455_166_0,
    i_13_455_191_0, i_13_455_241_0, i_13_455_269_0, i_13_455_278_0,
    i_13_455_287_0, i_13_455_314_0, i_13_455_340_0, i_13_455_358_0,
    i_13_455_385_0, i_13_455_386_0, i_13_455_466_0, i_13_455_470_0,
    i_13_455_592_0, i_13_455_593_0, i_13_455_745_0, i_13_455_746_0,
    i_13_455_768_0, i_13_455_823_0, i_13_455_824_0, i_13_455_827_0,
    i_13_455_851_0, i_13_455_916_0, i_13_455_947_0, i_13_455_952_0,
    i_13_455_985_0, i_13_455_1111_0, i_13_455_1120_0, i_13_455_1303_0,
    i_13_455_1304_0, i_13_455_1348_0, i_13_455_1435_0, i_13_455_1439_0,
    i_13_455_1447_0, i_13_455_1499_0, i_13_455_1501_0, i_13_455_1516_0,
    i_13_455_1541_0, i_13_455_1573_0, i_13_455_1574_0, i_13_455_1634_0,
    i_13_455_1682_0, i_13_455_1817_0, i_13_455_1867_0, i_13_455_1951_0,
    i_13_455_1952_0, i_13_455_1996_0, i_13_455_2033_0, i_13_455_2059_0,
    i_13_455_2060_0, i_13_455_2114_0, i_13_455_2123_0, i_13_455_2141_0,
    i_13_455_2284_0, i_13_455_2285_0, i_13_455_2401_0, i_13_455_2410_0,
    i_13_455_2411_0, i_13_455_2561_0, i_13_455_2570_0, i_13_455_2582_0,
    i_13_455_2590_0, i_13_455_2591_0, i_13_455_2617_0, i_13_455_2662_0,
    i_13_455_2720_0, i_13_455_2771_0, i_13_455_2824_0, i_13_455_2825_0,
    i_13_455_3064_0, i_13_455_3157_0, i_13_455_3221_0, i_13_455_3238_0,
    i_13_455_3240_0, i_13_455_3346_0, i_13_455_3347_0, i_13_455_3374_0,
    i_13_455_3419_0, i_13_455_3598_0, i_13_455_3599_0, i_13_455_3618_0,
    i_13_455_3623_0, i_13_455_3628_0, i_13_455_3634_0, i_13_455_3731_0,
    i_13_455_3733_0, i_13_455_3838_0, i_13_455_3923_0, i_13_455_3928_0,
    i_13_455_4048_0, i_13_455_4058_0, i_13_455_4237_0, i_13_455_4273_0,
    i_13_455_4274_0, i_13_455_4336_0, i_13_455_4400_0, i_13_455_4454_0,
    o_13_455_0_0  );
  input  i_13_455_2_0, i_13_455_156_0, i_13_455_164_0, i_13_455_166_0,
    i_13_455_191_0, i_13_455_241_0, i_13_455_269_0, i_13_455_278_0,
    i_13_455_287_0, i_13_455_314_0, i_13_455_340_0, i_13_455_358_0,
    i_13_455_385_0, i_13_455_386_0, i_13_455_466_0, i_13_455_470_0,
    i_13_455_592_0, i_13_455_593_0, i_13_455_745_0, i_13_455_746_0,
    i_13_455_768_0, i_13_455_823_0, i_13_455_824_0, i_13_455_827_0,
    i_13_455_851_0, i_13_455_916_0, i_13_455_947_0, i_13_455_952_0,
    i_13_455_985_0, i_13_455_1111_0, i_13_455_1120_0, i_13_455_1303_0,
    i_13_455_1304_0, i_13_455_1348_0, i_13_455_1435_0, i_13_455_1439_0,
    i_13_455_1447_0, i_13_455_1499_0, i_13_455_1501_0, i_13_455_1516_0,
    i_13_455_1541_0, i_13_455_1573_0, i_13_455_1574_0, i_13_455_1634_0,
    i_13_455_1682_0, i_13_455_1817_0, i_13_455_1867_0, i_13_455_1951_0,
    i_13_455_1952_0, i_13_455_1996_0, i_13_455_2033_0, i_13_455_2059_0,
    i_13_455_2060_0, i_13_455_2114_0, i_13_455_2123_0, i_13_455_2141_0,
    i_13_455_2284_0, i_13_455_2285_0, i_13_455_2401_0, i_13_455_2410_0,
    i_13_455_2411_0, i_13_455_2561_0, i_13_455_2570_0, i_13_455_2582_0,
    i_13_455_2590_0, i_13_455_2591_0, i_13_455_2617_0, i_13_455_2662_0,
    i_13_455_2720_0, i_13_455_2771_0, i_13_455_2824_0, i_13_455_2825_0,
    i_13_455_3064_0, i_13_455_3157_0, i_13_455_3221_0, i_13_455_3238_0,
    i_13_455_3240_0, i_13_455_3346_0, i_13_455_3347_0, i_13_455_3374_0,
    i_13_455_3419_0, i_13_455_3598_0, i_13_455_3599_0, i_13_455_3618_0,
    i_13_455_3623_0, i_13_455_3628_0, i_13_455_3634_0, i_13_455_3731_0,
    i_13_455_3733_0, i_13_455_3838_0, i_13_455_3923_0, i_13_455_3928_0,
    i_13_455_4048_0, i_13_455_4058_0, i_13_455_4237_0, i_13_455_4273_0,
    i_13_455_4274_0, i_13_455_4336_0, i_13_455_4400_0, i_13_455_4454_0;
  output o_13_455_0_0;
  assign o_13_455_0_0 = ~((~i_13_455_385_0 & ~i_13_455_3221_0 & ~i_13_455_3623_0) | (~i_13_455_340_0 & ~i_13_455_3238_0 & ~i_13_455_3599_0) | (~i_13_455_466_0 & ~i_13_455_2060_0 & ~i_13_455_2771_0));
endmodule



// Benchmark "kernel_13_456" written by ABC on Sun Jul 19 10:51:43 2020

module kernel_13_456 ( 
    i_13_456_39_0, i_13_456_40_0, i_13_456_48_0, i_13_456_49_0,
    i_13_456_68_0, i_13_456_70_0, i_13_456_159_0, i_13_456_259_0,
    i_13_456_277_0, i_13_456_351_0, i_13_456_411_0, i_13_456_453_0,
    i_13_456_520_0, i_13_456_535_0, i_13_456_628_0, i_13_456_673_0,
    i_13_456_760_0, i_13_456_834_0, i_13_456_900_0, i_13_456_934_0,
    i_13_456_939_0, i_13_456_1023_0, i_13_456_1104_0, i_13_456_1105_0,
    i_13_456_1150_0, i_13_456_1231_0, i_13_456_1330_0, i_13_456_1349_0,
    i_13_456_1363_0, i_13_456_1399_0, i_13_456_1402_0, i_13_456_1521_0,
    i_13_456_1596_0, i_13_456_1626_0, i_13_456_1644_0, i_13_456_1663_0,
    i_13_456_1668_0, i_13_456_1735_0, i_13_456_1780_0, i_13_456_1798_0,
    i_13_456_1884_0, i_13_456_1892_0, i_13_456_1894_0, i_13_456_1947_0,
    i_13_456_1948_0, i_13_456_2029_0, i_13_456_2058_0, i_13_456_2121_0,
    i_13_456_2148_0, i_13_456_2184_0, i_13_456_2228_0, i_13_456_2265_0,
    i_13_456_2299_0, i_13_456_2380_0, i_13_456_2399_0, i_13_456_2400_0,
    i_13_456_2436_0, i_13_456_2472_0, i_13_456_2517_0, i_13_456_2553_0,
    i_13_456_2571_0, i_13_456_2595_0, i_13_456_2614_0, i_13_456_2724_0,
    i_13_456_2742_0, i_13_456_2743_0, i_13_456_2874_0, i_13_456_2912_0,
    i_13_456_2915_0, i_13_456_2968_0, i_13_456_3030_0, i_13_456_3031_0,
    i_13_456_3111_0, i_13_456_3112_0, i_13_456_3135_0, i_13_456_3315_0,
    i_13_456_3355_0, i_13_456_3370_0, i_13_456_3399_0, i_13_456_3481_0,
    i_13_456_3489_0, i_13_456_3534_0, i_13_456_3739_0, i_13_456_3765_0,
    i_13_456_3767_0, i_13_456_3838_0, i_13_456_3842_0, i_13_456_3892_0,
    i_13_456_3900_0, i_13_456_3930_0, i_13_456_4002_0, i_13_456_4022_0,
    i_13_456_4055_0, i_13_456_4164_0, i_13_456_4174_0, i_13_456_4233_0,
    i_13_456_4254_0, i_13_456_4362_0, i_13_456_4478_0, i_13_456_4606_0,
    o_13_456_0_0  );
  input  i_13_456_39_0, i_13_456_40_0, i_13_456_48_0, i_13_456_49_0,
    i_13_456_68_0, i_13_456_70_0, i_13_456_159_0, i_13_456_259_0,
    i_13_456_277_0, i_13_456_351_0, i_13_456_411_0, i_13_456_453_0,
    i_13_456_520_0, i_13_456_535_0, i_13_456_628_0, i_13_456_673_0,
    i_13_456_760_0, i_13_456_834_0, i_13_456_900_0, i_13_456_934_0,
    i_13_456_939_0, i_13_456_1023_0, i_13_456_1104_0, i_13_456_1105_0,
    i_13_456_1150_0, i_13_456_1231_0, i_13_456_1330_0, i_13_456_1349_0,
    i_13_456_1363_0, i_13_456_1399_0, i_13_456_1402_0, i_13_456_1521_0,
    i_13_456_1596_0, i_13_456_1626_0, i_13_456_1644_0, i_13_456_1663_0,
    i_13_456_1668_0, i_13_456_1735_0, i_13_456_1780_0, i_13_456_1798_0,
    i_13_456_1884_0, i_13_456_1892_0, i_13_456_1894_0, i_13_456_1947_0,
    i_13_456_1948_0, i_13_456_2029_0, i_13_456_2058_0, i_13_456_2121_0,
    i_13_456_2148_0, i_13_456_2184_0, i_13_456_2228_0, i_13_456_2265_0,
    i_13_456_2299_0, i_13_456_2380_0, i_13_456_2399_0, i_13_456_2400_0,
    i_13_456_2436_0, i_13_456_2472_0, i_13_456_2517_0, i_13_456_2553_0,
    i_13_456_2571_0, i_13_456_2595_0, i_13_456_2614_0, i_13_456_2724_0,
    i_13_456_2742_0, i_13_456_2743_0, i_13_456_2874_0, i_13_456_2912_0,
    i_13_456_2915_0, i_13_456_2968_0, i_13_456_3030_0, i_13_456_3031_0,
    i_13_456_3111_0, i_13_456_3112_0, i_13_456_3135_0, i_13_456_3315_0,
    i_13_456_3355_0, i_13_456_3370_0, i_13_456_3399_0, i_13_456_3481_0,
    i_13_456_3489_0, i_13_456_3534_0, i_13_456_3739_0, i_13_456_3765_0,
    i_13_456_3767_0, i_13_456_3838_0, i_13_456_3842_0, i_13_456_3892_0,
    i_13_456_3900_0, i_13_456_3930_0, i_13_456_4002_0, i_13_456_4022_0,
    i_13_456_4055_0, i_13_456_4164_0, i_13_456_4174_0, i_13_456_4233_0,
    i_13_456_4254_0, i_13_456_4362_0, i_13_456_4478_0, i_13_456_4606_0;
  output o_13_456_0_0;
  assign o_13_456_0_0 = ~((~i_13_456_3900_0 & (~i_13_456_277_0 | ~i_13_456_2148_0)) | (i_13_456_535_0 & ~i_13_456_1330_0) | ~i_13_456_1735_0 | (~i_13_456_834_0 & ~i_13_456_3111_0));
endmodule



// Benchmark "kernel_13_457" written by ABC on Sun Jul 19 10:51:44 2020

module kernel_13_457 ( 
    i_13_457_51_0, i_13_457_52_0, i_13_457_97_0, i_13_457_106_0,
    i_13_457_159_0, i_13_457_196_0, i_13_457_286_0, i_13_457_340_0,
    i_13_457_385_0, i_13_457_467_0, i_13_457_574_0, i_13_457_592_0,
    i_13_457_625_0, i_13_457_688_0, i_13_457_700_0, i_13_457_745_0,
    i_13_457_817_0, i_13_457_948_0, i_13_457_962_0, i_13_457_985_0,
    i_13_457_1068_0, i_13_457_1069_0, i_13_457_1123_0, i_13_457_1150_0,
    i_13_457_1210_0, i_13_457_1258_0, i_13_457_1281_0, i_13_457_1308_0,
    i_13_457_1330_0, i_13_457_1574_0, i_13_457_1715_0, i_13_457_1780_0,
    i_13_457_1795_0, i_13_457_1806_0, i_13_457_1807_0, i_13_457_1808_0,
    i_13_457_1851_0, i_13_457_1852_0, i_13_457_1876_0, i_13_457_1932_0,
    i_13_457_1997_0, i_13_457_2002_0, i_13_457_2058_0, i_13_457_2059_0,
    i_13_457_2121_0, i_13_457_2123_0, i_13_457_2174_0, i_13_457_2194_0,
    i_13_457_2238_0, i_13_457_2266_0, i_13_457_2283_0, i_13_457_2284_0,
    i_13_457_2293_0, i_13_457_2343_0, i_13_457_2410_0, i_13_457_2429_0,
    i_13_457_2473_0, i_13_457_2498_0, i_13_457_2536_0, i_13_457_2573_0,
    i_13_457_2617_0, i_13_457_2752_0, i_13_457_2914_0, i_13_457_2920_0,
    i_13_457_2941_0, i_13_457_2986_0, i_13_457_3022_0, i_13_457_3023_0,
    i_13_457_3028_0, i_13_457_3109_0, i_13_457_3210_0, i_13_457_3211_0,
    i_13_457_3303_0, i_13_457_3346_0, i_13_457_3351_0, i_13_457_3391_0,
    i_13_457_3399_0, i_13_457_3401_0, i_13_457_3451_0, i_13_457_3504_0,
    i_13_457_3525_0, i_13_457_3526_0, i_13_457_3766_0, i_13_457_3850_0,
    i_13_457_3909_0, i_13_457_3911_0, i_13_457_4021_0, i_13_457_4047_0,
    i_13_457_4048_0, i_13_457_4049_0, i_13_457_4066_0, i_13_457_4084_0,
    i_13_457_4184_0, i_13_457_4234_0, i_13_457_4297_0, i_13_457_4308_0,
    i_13_457_4309_0, i_13_457_4318_0, i_13_457_4345_0, i_13_457_4346_0,
    o_13_457_0_0  );
  input  i_13_457_51_0, i_13_457_52_0, i_13_457_97_0, i_13_457_106_0,
    i_13_457_159_0, i_13_457_196_0, i_13_457_286_0, i_13_457_340_0,
    i_13_457_385_0, i_13_457_467_0, i_13_457_574_0, i_13_457_592_0,
    i_13_457_625_0, i_13_457_688_0, i_13_457_700_0, i_13_457_745_0,
    i_13_457_817_0, i_13_457_948_0, i_13_457_962_0, i_13_457_985_0,
    i_13_457_1068_0, i_13_457_1069_0, i_13_457_1123_0, i_13_457_1150_0,
    i_13_457_1210_0, i_13_457_1258_0, i_13_457_1281_0, i_13_457_1308_0,
    i_13_457_1330_0, i_13_457_1574_0, i_13_457_1715_0, i_13_457_1780_0,
    i_13_457_1795_0, i_13_457_1806_0, i_13_457_1807_0, i_13_457_1808_0,
    i_13_457_1851_0, i_13_457_1852_0, i_13_457_1876_0, i_13_457_1932_0,
    i_13_457_1997_0, i_13_457_2002_0, i_13_457_2058_0, i_13_457_2059_0,
    i_13_457_2121_0, i_13_457_2123_0, i_13_457_2174_0, i_13_457_2194_0,
    i_13_457_2238_0, i_13_457_2266_0, i_13_457_2283_0, i_13_457_2284_0,
    i_13_457_2293_0, i_13_457_2343_0, i_13_457_2410_0, i_13_457_2429_0,
    i_13_457_2473_0, i_13_457_2498_0, i_13_457_2536_0, i_13_457_2573_0,
    i_13_457_2617_0, i_13_457_2752_0, i_13_457_2914_0, i_13_457_2920_0,
    i_13_457_2941_0, i_13_457_2986_0, i_13_457_3022_0, i_13_457_3023_0,
    i_13_457_3028_0, i_13_457_3109_0, i_13_457_3210_0, i_13_457_3211_0,
    i_13_457_3303_0, i_13_457_3346_0, i_13_457_3351_0, i_13_457_3391_0,
    i_13_457_3399_0, i_13_457_3401_0, i_13_457_3451_0, i_13_457_3504_0,
    i_13_457_3525_0, i_13_457_3526_0, i_13_457_3766_0, i_13_457_3850_0,
    i_13_457_3909_0, i_13_457_3911_0, i_13_457_4021_0, i_13_457_4047_0,
    i_13_457_4048_0, i_13_457_4049_0, i_13_457_4066_0, i_13_457_4084_0,
    i_13_457_4184_0, i_13_457_4234_0, i_13_457_4297_0, i_13_457_4308_0,
    i_13_457_4309_0, i_13_457_4318_0, i_13_457_4345_0, i_13_457_4346_0;
  output o_13_457_0_0;
  assign o_13_457_0_0 = ~((i_13_457_1258_0 & ((~i_13_457_1308_0 & ~i_13_457_2941_0 & ~i_13_457_3346_0) | (~i_13_457_1932_0 & i_13_457_3850_0 & ~i_13_457_4309_0))) | (~i_13_457_3399_0 & ((~i_13_457_1330_0 & ~i_13_457_2002_0) | (~i_13_457_106_0 & ~i_13_457_286_0 & i_13_457_1210_0 & ~i_13_457_3911_0))) | (~i_13_457_286_0 & ((~i_13_457_385_0 & ~i_13_457_1069_0 & i_13_457_1795_0 & ~i_13_457_2986_0) | (~i_13_457_340_0 & ~i_13_457_1807_0 & ~i_13_457_3766_0))) | (~i_13_457_1808_0 & ~i_13_457_3109_0 & ~i_13_457_3210_0 & ~i_13_457_3211_0 & ~i_13_457_4048_0) | (~i_13_457_1123_0 & ~i_13_457_2284_0 & ~i_13_457_3346_0 & ~i_13_457_4318_0));
endmodule



// Benchmark "kernel_13_458" written by ABC on Sun Jul 19 10:51:45 2020

module kernel_13_458 ( 
    i_13_458_136_0, i_13_458_138_0, i_13_458_139_0, i_13_458_172_0,
    i_13_458_229_0, i_13_458_257_0, i_13_458_308_0, i_13_458_370_0,
    i_13_458_409_0, i_13_458_512_0, i_13_458_535_0, i_13_458_554_0,
    i_13_458_568_0, i_13_458_657_0, i_13_458_661_0, i_13_458_675_0,
    i_13_458_676_0, i_13_458_697_0, i_13_458_793_0, i_13_458_842_0,
    i_13_458_851_0, i_13_458_937_0, i_13_458_981_0, i_13_458_983_0,
    i_13_458_985_0, i_13_458_986_0, i_13_458_1066_0, i_13_458_1119_0,
    i_13_458_1134_0, i_13_458_1202_0, i_13_458_1219_0, i_13_458_1274_0,
    i_13_458_1324_0, i_13_458_1327_0, i_13_458_1328_0, i_13_458_1526_0,
    i_13_458_1629_0, i_13_458_1828_0, i_13_458_1885_0, i_13_458_1913_0,
    i_13_458_2020_0, i_13_458_2107_0, i_13_458_2182_0, i_13_458_2233_0,
    i_13_458_2242_0, i_13_458_2296_0, i_13_458_2299_0, i_13_458_2347_0,
    i_13_458_2430_0, i_13_458_2461_0, i_13_458_2467_0, i_13_458_2469_0,
    i_13_458_2470_0, i_13_458_2592_0, i_13_458_2695_0, i_13_458_2848_0,
    i_13_458_2850_0, i_13_458_2872_0, i_13_458_2875_0, i_13_458_2914_0,
    i_13_458_2980_0, i_13_458_2983_0, i_13_458_3006_0, i_13_458_3010_0,
    i_13_458_3073_0, i_13_458_3105_0, i_13_458_3106_0, i_13_458_3108_0,
    i_13_458_3151_0, i_13_458_3205_0, i_13_458_3207_0, i_13_458_3212_0,
    i_13_458_3335_0, i_13_458_3388_0, i_13_458_3397_0, i_13_458_3406_0,
    i_13_458_3442_0, i_13_458_3465_0, i_13_458_3479_0, i_13_458_3547_0,
    i_13_458_3763_0, i_13_458_3764_0, i_13_458_3817_0, i_13_458_3820_0,
    i_13_458_3826_0, i_13_458_3862_0, i_13_458_3916_0, i_13_458_3979_0,
    i_13_458_4072_0, i_13_458_4123_0, i_13_458_4159_0, i_13_458_4163_0,
    i_13_458_4203_0, i_13_458_4254_0, i_13_458_4327_0, i_13_458_4554_0,
    i_13_458_4563_0, i_13_458_4565_0, i_13_458_4567_0, i_13_458_4600_0,
    o_13_458_0_0  );
  input  i_13_458_136_0, i_13_458_138_0, i_13_458_139_0, i_13_458_172_0,
    i_13_458_229_0, i_13_458_257_0, i_13_458_308_0, i_13_458_370_0,
    i_13_458_409_0, i_13_458_512_0, i_13_458_535_0, i_13_458_554_0,
    i_13_458_568_0, i_13_458_657_0, i_13_458_661_0, i_13_458_675_0,
    i_13_458_676_0, i_13_458_697_0, i_13_458_793_0, i_13_458_842_0,
    i_13_458_851_0, i_13_458_937_0, i_13_458_981_0, i_13_458_983_0,
    i_13_458_985_0, i_13_458_986_0, i_13_458_1066_0, i_13_458_1119_0,
    i_13_458_1134_0, i_13_458_1202_0, i_13_458_1219_0, i_13_458_1274_0,
    i_13_458_1324_0, i_13_458_1327_0, i_13_458_1328_0, i_13_458_1526_0,
    i_13_458_1629_0, i_13_458_1828_0, i_13_458_1885_0, i_13_458_1913_0,
    i_13_458_2020_0, i_13_458_2107_0, i_13_458_2182_0, i_13_458_2233_0,
    i_13_458_2242_0, i_13_458_2296_0, i_13_458_2299_0, i_13_458_2347_0,
    i_13_458_2430_0, i_13_458_2461_0, i_13_458_2467_0, i_13_458_2469_0,
    i_13_458_2470_0, i_13_458_2592_0, i_13_458_2695_0, i_13_458_2848_0,
    i_13_458_2850_0, i_13_458_2872_0, i_13_458_2875_0, i_13_458_2914_0,
    i_13_458_2980_0, i_13_458_2983_0, i_13_458_3006_0, i_13_458_3010_0,
    i_13_458_3073_0, i_13_458_3105_0, i_13_458_3106_0, i_13_458_3108_0,
    i_13_458_3151_0, i_13_458_3205_0, i_13_458_3207_0, i_13_458_3212_0,
    i_13_458_3335_0, i_13_458_3388_0, i_13_458_3397_0, i_13_458_3406_0,
    i_13_458_3442_0, i_13_458_3465_0, i_13_458_3479_0, i_13_458_3547_0,
    i_13_458_3763_0, i_13_458_3764_0, i_13_458_3817_0, i_13_458_3820_0,
    i_13_458_3826_0, i_13_458_3862_0, i_13_458_3916_0, i_13_458_3979_0,
    i_13_458_4072_0, i_13_458_4123_0, i_13_458_4159_0, i_13_458_4163_0,
    i_13_458_4203_0, i_13_458_4254_0, i_13_458_4327_0, i_13_458_4554_0,
    i_13_458_4563_0, i_13_458_4565_0, i_13_458_4567_0, i_13_458_4600_0;
  output o_13_458_0_0;
  assign o_13_458_0_0 = ~((i_13_458_139_0 & ((~i_13_458_370_0 & ~i_13_458_2020_0) | (~i_13_458_676_0 & ~i_13_458_1324_0 & ~i_13_458_2983_0))) | (~i_13_458_3820_0 & ((~i_13_458_172_0 & ~i_13_458_2299_0 & ((~i_13_458_2430_0 & i_13_458_3388_0) | (~i_13_458_3105_0 & ~i_13_458_3108_0 & ~i_13_458_3212_0 & ~i_13_458_3547_0))) | (~i_13_458_1526_0 & ~i_13_458_1828_0 & ~i_13_458_3106_0 & ~i_13_458_3207_0 & ~i_13_458_3764_0 & ~i_13_458_3979_0 & ~i_13_458_4567_0))) | (~i_13_458_1324_0 & ((~i_13_458_568_0 & i_13_458_2872_0 & i_13_458_3205_0) | (i_13_458_697_0 & ~i_13_458_1202_0 & ~i_13_458_2983_0 & ~i_13_458_3763_0))) | (~i_13_458_3207_0 & i_13_458_4254_0 & (i_13_458_2875_0 | i_13_458_3820_0)) | (~i_13_458_2983_0 & ~i_13_458_3010_0 & i_13_458_3388_0) | (~i_13_458_981_0 & ~i_13_458_1328_0 & ~i_13_458_2242_0 & ~i_13_458_3108_0 & ~i_13_458_3205_0 & ~i_13_458_3764_0 & ~i_13_458_3817_0) | (~i_13_458_1327_0 & i_13_458_1885_0 & i_13_458_3862_0));
endmodule



// Benchmark "kernel_13_459" written by ABC on Sun Jul 19 10:51:46 2020

module kernel_13_459 ( 
    i_13_459_59_0, i_13_459_136_0, i_13_459_137_0, i_13_459_173_0,
    i_13_459_203_0, i_13_459_256_0, i_13_459_284_0, i_13_459_311_0,
    i_13_459_334_0, i_13_459_352_0, i_13_459_518_0, i_13_459_523_0,
    i_13_459_613_0, i_13_459_622_0, i_13_459_626_0, i_13_459_641_0,
    i_13_459_644_0, i_13_459_685_0, i_13_459_686_0, i_13_459_695_0,
    i_13_459_824_0, i_13_459_976_0, i_13_459_1117_0, i_13_459_1118_0,
    i_13_459_1201_0, i_13_459_1208_0, i_13_459_1270_0, i_13_459_1271_0,
    i_13_459_1273_0, i_13_459_1274_0, i_13_459_1282_0, i_13_459_1315_0,
    i_13_459_1388_0, i_13_459_1444_0, i_13_459_1468_0, i_13_459_1469_0,
    i_13_459_1481_0, i_13_459_1625_0, i_13_459_1640_0, i_13_459_1643_0,
    i_13_459_1667_0, i_13_459_1678_0, i_13_459_1711_0, i_13_459_1712_0,
    i_13_459_1732_0, i_13_459_1793_0, i_13_459_1802_0, i_13_459_1882_0,
    i_13_459_1883_0, i_13_459_1945_0, i_13_459_1991_0, i_13_459_2044_0,
    i_13_459_2134_0, i_13_459_2135_0, i_13_459_2245_0, i_13_459_2314_0,
    i_13_459_2351_0, i_13_459_2377_0, i_13_459_2378_0, i_13_459_2380_0,
    i_13_459_2542_0, i_13_459_2549_0, i_13_459_2551_0, i_13_459_2567_0,
    i_13_459_2592_0, i_13_459_2647_0, i_13_459_2648_0, i_13_459_2651_0,
    i_13_459_2669_0, i_13_459_2728_0, i_13_459_2747_0, i_13_459_2750_0,
    i_13_459_2845_0, i_13_459_2846_0, i_13_459_2848_0, i_13_459_2849_0,
    i_13_459_2873_0, i_13_459_2875_0, i_13_459_2903_0, i_13_459_3199_0,
    i_13_459_3235_0, i_13_459_3385_0, i_13_459_3403_0, i_13_459_3430_0,
    i_13_459_3556_0, i_13_459_3559_0, i_13_459_3568_0, i_13_459_3791_0,
    i_13_459_4018_0, i_13_459_4034_0, i_13_459_4186_0, i_13_459_4187_0,
    i_13_459_4234_0, i_13_459_4262_0, i_13_459_4294_0, i_13_459_4295_0,
    i_13_459_4351_0, i_13_459_4352_0, i_13_459_4376_0, i_13_459_4495_0,
    o_13_459_0_0  );
  input  i_13_459_59_0, i_13_459_136_0, i_13_459_137_0, i_13_459_173_0,
    i_13_459_203_0, i_13_459_256_0, i_13_459_284_0, i_13_459_311_0,
    i_13_459_334_0, i_13_459_352_0, i_13_459_518_0, i_13_459_523_0,
    i_13_459_613_0, i_13_459_622_0, i_13_459_626_0, i_13_459_641_0,
    i_13_459_644_0, i_13_459_685_0, i_13_459_686_0, i_13_459_695_0,
    i_13_459_824_0, i_13_459_976_0, i_13_459_1117_0, i_13_459_1118_0,
    i_13_459_1201_0, i_13_459_1208_0, i_13_459_1270_0, i_13_459_1271_0,
    i_13_459_1273_0, i_13_459_1274_0, i_13_459_1282_0, i_13_459_1315_0,
    i_13_459_1388_0, i_13_459_1444_0, i_13_459_1468_0, i_13_459_1469_0,
    i_13_459_1481_0, i_13_459_1625_0, i_13_459_1640_0, i_13_459_1643_0,
    i_13_459_1667_0, i_13_459_1678_0, i_13_459_1711_0, i_13_459_1712_0,
    i_13_459_1732_0, i_13_459_1793_0, i_13_459_1802_0, i_13_459_1882_0,
    i_13_459_1883_0, i_13_459_1945_0, i_13_459_1991_0, i_13_459_2044_0,
    i_13_459_2134_0, i_13_459_2135_0, i_13_459_2245_0, i_13_459_2314_0,
    i_13_459_2351_0, i_13_459_2377_0, i_13_459_2378_0, i_13_459_2380_0,
    i_13_459_2542_0, i_13_459_2549_0, i_13_459_2551_0, i_13_459_2567_0,
    i_13_459_2592_0, i_13_459_2647_0, i_13_459_2648_0, i_13_459_2651_0,
    i_13_459_2669_0, i_13_459_2728_0, i_13_459_2747_0, i_13_459_2750_0,
    i_13_459_2845_0, i_13_459_2846_0, i_13_459_2848_0, i_13_459_2849_0,
    i_13_459_2873_0, i_13_459_2875_0, i_13_459_2903_0, i_13_459_3199_0,
    i_13_459_3235_0, i_13_459_3385_0, i_13_459_3403_0, i_13_459_3430_0,
    i_13_459_3556_0, i_13_459_3559_0, i_13_459_3568_0, i_13_459_3791_0,
    i_13_459_4018_0, i_13_459_4034_0, i_13_459_4186_0, i_13_459_4187_0,
    i_13_459_4234_0, i_13_459_4262_0, i_13_459_4294_0, i_13_459_4295_0,
    i_13_459_4351_0, i_13_459_4352_0, i_13_459_4376_0, i_13_459_4495_0;
  output o_13_459_0_0;
  assign o_13_459_0_0 = ~(~i_13_459_2377_0 | (~i_13_459_1991_0 & ~i_13_459_2849_0) | (~i_13_459_1643_0 & ~i_13_459_1882_0));
endmodule



// Benchmark "kernel_13_460" written by ABC on Sun Jul 19 10:51:46 2020

module kernel_13_460 ( 
    i_13_460_40_0, i_13_460_61_0, i_13_460_79_0, i_13_460_105_0,
    i_13_460_115_0, i_13_460_124_0, i_13_460_169_0, i_13_460_268_0,
    i_13_460_269_0, i_13_460_391_0, i_13_460_465_0, i_13_460_466_0,
    i_13_460_509_0, i_13_460_673_0, i_13_460_689_0, i_13_460_734_0,
    i_13_460_813_0, i_13_460_815_0, i_13_460_816_0, i_13_460_817_0,
    i_13_460_935_0, i_13_460_952_0, i_13_460_1201_0, i_13_460_1210_0,
    i_13_460_1302_0, i_13_460_1303_0, i_13_460_1304_0, i_13_460_1331_0,
    i_13_460_1348_0, i_13_460_1447_0, i_13_460_1464_0, i_13_460_1554_0,
    i_13_460_1607_0, i_13_460_1713_0, i_13_460_1753_0, i_13_460_1789_0,
    i_13_460_1806_0, i_13_460_1807_0, i_13_460_1857_0, i_13_460_1858_0,
    i_13_460_1906_0, i_13_460_1943_0, i_13_460_1995_0, i_13_460_2114_0,
    i_13_460_2122_0, i_13_460_2139_0, i_13_460_2140_0, i_13_460_2141_0,
    i_13_460_2202_0, i_13_460_2224_0, i_13_460_2239_0, i_13_460_2247_0,
    i_13_460_2410_0, i_13_460_2446_0, i_13_460_2463_0, i_13_460_2496_0,
    i_13_460_2694_0, i_13_460_2696_0, i_13_460_2798_0, i_13_460_2823_0,
    i_13_460_2824_0, i_13_460_2825_0, i_13_460_2912_0, i_13_460_2920_0,
    i_13_460_2938_0, i_13_460_2941_0, i_13_460_2986_0, i_13_460_3022_0,
    i_13_460_3092_0, i_13_460_3244_0, i_13_460_3273_0, i_13_460_3346_0,
    i_13_460_3347_0, i_13_460_3373_0, i_13_460_3374_0, i_13_460_3391_0,
    i_13_460_3418_0, i_13_460_3427_0, i_13_460_3455_0, i_13_460_3505_0,
    i_13_460_3622_0, i_13_460_3633_0, i_13_460_3793_0, i_13_460_3824_0,
    i_13_460_3913_0, i_13_460_3991_0, i_13_460_3992_0, i_13_460_4046_0,
    i_13_460_4047_0, i_13_460_4058_0, i_13_460_4081_0, i_13_460_4162_0,
    i_13_460_4237_0, i_13_460_4308_0, i_13_460_4342_0, i_13_460_4344_0,
    i_13_460_4372_0, i_13_460_4380_0, i_13_460_4381_0, i_13_460_4526_0,
    o_13_460_0_0  );
  input  i_13_460_40_0, i_13_460_61_0, i_13_460_79_0, i_13_460_105_0,
    i_13_460_115_0, i_13_460_124_0, i_13_460_169_0, i_13_460_268_0,
    i_13_460_269_0, i_13_460_391_0, i_13_460_465_0, i_13_460_466_0,
    i_13_460_509_0, i_13_460_673_0, i_13_460_689_0, i_13_460_734_0,
    i_13_460_813_0, i_13_460_815_0, i_13_460_816_0, i_13_460_817_0,
    i_13_460_935_0, i_13_460_952_0, i_13_460_1201_0, i_13_460_1210_0,
    i_13_460_1302_0, i_13_460_1303_0, i_13_460_1304_0, i_13_460_1331_0,
    i_13_460_1348_0, i_13_460_1447_0, i_13_460_1464_0, i_13_460_1554_0,
    i_13_460_1607_0, i_13_460_1713_0, i_13_460_1753_0, i_13_460_1789_0,
    i_13_460_1806_0, i_13_460_1807_0, i_13_460_1857_0, i_13_460_1858_0,
    i_13_460_1906_0, i_13_460_1943_0, i_13_460_1995_0, i_13_460_2114_0,
    i_13_460_2122_0, i_13_460_2139_0, i_13_460_2140_0, i_13_460_2141_0,
    i_13_460_2202_0, i_13_460_2224_0, i_13_460_2239_0, i_13_460_2247_0,
    i_13_460_2410_0, i_13_460_2446_0, i_13_460_2463_0, i_13_460_2496_0,
    i_13_460_2694_0, i_13_460_2696_0, i_13_460_2798_0, i_13_460_2823_0,
    i_13_460_2824_0, i_13_460_2825_0, i_13_460_2912_0, i_13_460_2920_0,
    i_13_460_2938_0, i_13_460_2941_0, i_13_460_2986_0, i_13_460_3022_0,
    i_13_460_3092_0, i_13_460_3244_0, i_13_460_3273_0, i_13_460_3346_0,
    i_13_460_3347_0, i_13_460_3373_0, i_13_460_3374_0, i_13_460_3391_0,
    i_13_460_3418_0, i_13_460_3427_0, i_13_460_3455_0, i_13_460_3505_0,
    i_13_460_3622_0, i_13_460_3633_0, i_13_460_3793_0, i_13_460_3824_0,
    i_13_460_3913_0, i_13_460_3991_0, i_13_460_3992_0, i_13_460_4046_0,
    i_13_460_4047_0, i_13_460_4058_0, i_13_460_4081_0, i_13_460_4162_0,
    i_13_460_4237_0, i_13_460_4308_0, i_13_460_4342_0, i_13_460_4344_0,
    i_13_460_4372_0, i_13_460_4380_0, i_13_460_4381_0, i_13_460_4526_0;
  output o_13_460_0_0;
  assign o_13_460_0_0 = ~((i_13_460_3244_0 & (~i_13_460_4237_0 | (~i_13_460_79_0 & i_13_460_952_0))) | (~i_13_460_2139_0 & ~i_13_460_2140_0 & ~i_13_460_2141_0 & ~i_13_460_2239_0) | (~i_13_460_3427_0 & i_13_460_3455_0));
endmodule



// Benchmark "kernel_13_461" written by ABC on Sun Jul 19 10:51:47 2020

module kernel_13_461 ( 
    i_13_461_28_0, i_13_461_30_0, i_13_461_64_0, i_13_461_65_0,
    i_13_461_74_0, i_13_461_113_0, i_13_461_122_0, i_13_461_157_0,
    i_13_461_266_0, i_13_461_382_0, i_13_461_441_0, i_13_461_551_0,
    i_13_461_651_0, i_13_461_658_0, i_13_461_659_0, i_13_461_814_0,
    i_13_461_815_0, i_13_461_829_0, i_13_461_887_0, i_13_461_929_0,
    i_13_461_940_0, i_13_461_941_0, i_13_461_1082_0, i_13_461_1119_0,
    i_13_461_1125_0, i_13_461_1145_0, i_13_461_1208_0, i_13_461_1307_0,
    i_13_461_1344_0, i_13_461_1388_0, i_13_461_1389_0, i_13_461_1404_0,
    i_13_461_1424_0, i_13_461_1470_0, i_13_461_1593_0, i_13_461_1597_0,
    i_13_461_1657_0, i_13_461_1668_0, i_13_461_1712_0, i_13_461_1730_0,
    i_13_461_1755_0, i_13_461_1837_0, i_13_461_1838_0, i_13_461_1929_0,
    i_13_461_1993_0, i_13_461_1994_0, i_13_461_2016_0, i_13_461_2137_0,
    i_13_461_2170_0, i_13_461_2192_0, i_13_461_2405_0, i_13_461_2468_0,
    i_13_461_2610_0, i_13_461_2712_0, i_13_461_2845_0, i_13_461_2846_0,
    i_13_461_2847_0, i_13_461_2884_0, i_13_461_2939_0, i_13_461_3028_0,
    i_13_461_3063_0, i_13_461_3106_0, i_13_461_3157_0, i_13_461_3204_0,
    i_13_461_3240_0, i_13_461_3261_0, i_13_461_3387_0, i_13_461_3487_0,
    i_13_461_3502_0, i_13_461_3503_0, i_13_461_3569_0, i_13_461_3577_0,
    i_13_461_3618_0, i_13_461_3636_0, i_13_461_3646_0, i_13_461_3648_0,
    i_13_461_3667_0, i_13_461_3736_0, i_13_461_3738_0, i_13_461_3767_0,
    i_13_461_3889_0, i_13_461_3907_0, i_13_461_3915_0, i_13_461_4054_0,
    i_13_461_4078_0, i_13_461_4088_0, i_13_461_4160_0, i_13_461_4162_0,
    i_13_461_4164_0, i_13_461_4187_0, i_13_461_4233_0, i_13_461_4276_0,
    i_13_461_4330_0, i_13_461_4340_0, i_13_461_4365_0, i_13_461_4430_0,
    i_13_461_4540_0, i_13_461_4592_0, i_13_461_4600_0, i_13_461_4601_0,
    o_13_461_0_0  );
  input  i_13_461_28_0, i_13_461_30_0, i_13_461_64_0, i_13_461_65_0,
    i_13_461_74_0, i_13_461_113_0, i_13_461_122_0, i_13_461_157_0,
    i_13_461_266_0, i_13_461_382_0, i_13_461_441_0, i_13_461_551_0,
    i_13_461_651_0, i_13_461_658_0, i_13_461_659_0, i_13_461_814_0,
    i_13_461_815_0, i_13_461_829_0, i_13_461_887_0, i_13_461_929_0,
    i_13_461_940_0, i_13_461_941_0, i_13_461_1082_0, i_13_461_1119_0,
    i_13_461_1125_0, i_13_461_1145_0, i_13_461_1208_0, i_13_461_1307_0,
    i_13_461_1344_0, i_13_461_1388_0, i_13_461_1389_0, i_13_461_1404_0,
    i_13_461_1424_0, i_13_461_1470_0, i_13_461_1593_0, i_13_461_1597_0,
    i_13_461_1657_0, i_13_461_1668_0, i_13_461_1712_0, i_13_461_1730_0,
    i_13_461_1755_0, i_13_461_1837_0, i_13_461_1838_0, i_13_461_1929_0,
    i_13_461_1993_0, i_13_461_1994_0, i_13_461_2016_0, i_13_461_2137_0,
    i_13_461_2170_0, i_13_461_2192_0, i_13_461_2405_0, i_13_461_2468_0,
    i_13_461_2610_0, i_13_461_2712_0, i_13_461_2845_0, i_13_461_2846_0,
    i_13_461_2847_0, i_13_461_2884_0, i_13_461_2939_0, i_13_461_3028_0,
    i_13_461_3063_0, i_13_461_3106_0, i_13_461_3157_0, i_13_461_3204_0,
    i_13_461_3240_0, i_13_461_3261_0, i_13_461_3387_0, i_13_461_3487_0,
    i_13_461_3502_0, i_13_461_3503_0, i_13_461_3569_0, i_13_461_3577_0,
    i_13_461_3618_0, i_13_461_3636_0, i_13_461_3646_0, i_13_461_3648_0,
    i_13_461_3667_0, i_13_461_3736_0, i_13_461_3738_0, i_13_461_3767_0,
    i_13_461_3889_0, i_13_461_3907_0, i_13_461_3915_0, i_13_461_4054_0,
    i_13_461_4078_0, i_13_461_4088_0, i_13_461_4160_0, i_13_461_4162_0,
    i_13_461_4164_0, i_13_461_4187_0, i_13_461_4233_0, i_13_461_4276_0,
    i_13_461_4330_0, i_13_461_4340_0, i_13_461_4365_0, i_13_461_4430_0,
    i_13_461_4540_0, i_13_461_4592_0, i_13_461_4600_0, i_13_461_4601_0;
  output o_13_461_0_0;
  assign o_13_461_0_0 = ~(~i_13_461_4430_0 | ~i_13_461_1838_0 | ~i_13_461_3503_0);
endmodule



// Benchmark "kernel_13_462" written by ABC on Sun Jul 19 10:51:48 2020

module kernel_13_462 ( 
    i_13_462_49_0, i_13_462_50_0, i_13_462_138_0, i_13_462_139_0,
    i_13_462_231_0, i_13_462_256_0, i_13_462_268_0, i_13_462_447_0,
    i_13_462_492_0, i_13_462_517_0, i_13_462_537_0, i_13_462_589_0,
    i_13_462_615_0, i_13_462_626_0, i_13_462_643_0, i_13_462_644_0,
    i_13_462_645_0, i_13_462_686_0, i_13_462_688_0, i_13_462_690_0,
    i_13_462_699_0, i_13_462_822_0, i_13_462_897_0, i_13_462_976_0,
    i_13_462_1118_0, i_13_462_1120_0, i_13_462_1123_0, i_13_462_1197_0,
    i_13_462_1221_0, i_13_462_1273_0, i_13_462_1274_0, i_13_462_1389_0,
    i_13_462_1390_0, i_13_462_1392_0, i_13_462_1480_0, i_13_462_1644_0,
    i_13_462_1645_0, i_13_462_1649_0, i_13_462_1713_0, i_13_462_1725_0,
    i_13_462_1726_0, i_13_462_1735_0, i_13_462_1762_0, i_13_462_1779_0,
    i_13_462_1795_0, i_13_462_1796_0, i_13_462_1797_0, i_13_462_1798_0,
    i_13_462_1803_0, i_13_462_1831_0, i_13_462_1849_0, i_13_462_1885_0,
    i_13_462_1992_0, i_13_462_1994_0, i_13_462_2137_0, i_13_462_2191_0,
    i_13_462_2379_0, i_13_462_2616_0, i_13_462_2648_0, i_13_462_2748_0,
    i_13_462_2751_0, i_13_462_2757_0, i_13_462_2847_0, i_13_462_2848_0,
    i_13_462_2849_0, i_13_462_2851_0, i_13_462_2875_0, i_13_462_3039_0,
    i_13_462_3270_0, i_13_462_3368_0, i_13_462_3407_0, i_13_462_3432_0,
    i_13_462_3523_0, i_13_462_3534_0, i_13_462_3575_0, i_13_462_3670_0,
    i_13_462_3724_0, i_13_462_3730_0, i_13_462_3759_0, i_13_462_3838_0,
    i_13_462_3897_0, i_13_462_3930_0, i_13_462_3994_0, i_13_462_4054_0,
    i_13_462_4063_0, i_13_462_4099_0, i_13_462_4101_0, i_13_462_4125_0,
    i_13_462_4187_0, i_13_462_4189_0, i_13_462_4294_0, i_13_462_4297_0,
    i_13_462_4306_0, i_13_462_4341_0, i_13_462_4369_0, i_13_462_4396_0,
    i_13_462_4414_0, i_13_462_4449_0, i_13_462_4584_0, i_13_462_4597_0,
    o_13_462_0_0  );
  input  i_13_462_49_0, i_13_462_50_0, i_13_462_138_0, i_13_462_139_0,
    i_13_462_231_0, i_13_462_256_0, i_13_462_268_0, i_13_462_447_0,
    i_13_462_492_0, i_13_462_517_0, i_13_462_537_0, i_13_462_589_0,
    i_13_462_615_0, i_13_462_626_0, i_13_462_643_0, i_13_462_644_0,
    i_13_462_645_0, i_13_462_686_0, i_13_462_688_0, i_13_462_690_0,
    i_13_462_699_0, i_13_462_822_0, i_13_462_897_0, i_13_462_976_0,
    i_13_462_1118_0, i_13_462_1120_0, i_13_462_1123_0, i_13_462_1197_0,
    i_13_462_1221_0, i_13_462_1273_0, i_13_462_1274_0, i_13_462_1389_0,
    i_13_462_1390_0, i_13_462_1392_0, i_13_462_1480_0, i_13_462_1644_0,
    i_13_462_1645_0, i_13_462_1649_0, i_13_462_1713_0, i_13_462_1725_0,
    i_13_462_1726_0, i_13_462_1735_0, i_13_462_1762_0, i_13_462_1779_0,
    i_13_462_1795_0, i_13_462_1796_0, i_13_462_1797_0, i_13_462_1798_0,
    i_13_462_1803_0, i_13_462_1831_0, i_13_462_1849_0, i_13_462_1885_0,
    i_13_462_1992_0, i_13_462_1994_0, i_13_462_2137_0, i_13_462_2191_0,
    i_13_462_2379_0, i_13_462_2616_0, i_13_462_2648_0, i_13_462_2748_0,
    i_13_462_2751_0, i_13_462_2757_0, i_13_462_2847_0, i_13_462_2848_0,
    i_13_462_2849_0, i_13_462_2851_0, i_13_462_2875_0, i_13_462_3039_0,
    i_13_462_3270_0, i_13_462_3368_0, i_13_462_3407_0, i_13_462_3432_0,
    i_13_462_3523_0, i_13_462_3534_0, i_13_462_3575_0, i_13_462_3670_0,
    i_13_462_3724_0, i_13_462_3730_0, i_13_462_3759_0, i_13_462_3838_0,
    i_13_462_3897_0, i_13_462_3930_0, i_13_462_3994_0, i_13_462_4054_0,
    i_13_462_4063_0, i_13_462_4099_0, i_13_462_4101_0, i_13_462_4125_0,
    i_13_462_4187_0, i_13_462_4189_0, i_13_462_4294_0, i_13_462_4297_0,
    i_13_462_4306_0, i_13_462_4341_0, i_13_462_4369_0, i_13_462_4396_0,
    i_13_462_4414_0, i_13_462_4449_0, i_13_462_4584_0, i_13_462_4597_0;
  output o_13_462_0_0;
  assign o_13_462_0_0 = ~((~i_13_462_1713_0 & (i_13_462_4063_0 | (~i_13_462_1994_0 & ~i_13_462_4306_0))) | (~i_13_462_2849_0 & ((~i_13_462_231_0 & ~i_13_462_897_0 & ~i_13_462_1795_0 & ~i_13_462_2847_0) | (~i_13_462_1992_0 & ~i_13_462_4449_0))) | (~i_13_462_4449_0 & (i_13_462_517_0 | (~i_13_462_4054_0 & ~i_13_462_4306_0))) | (~i_13_462_4306_0 & ((~i_13_462_256_0 & ~i_13_462_3759_0) | (~i_13_462_2851_0 & ~i_13_462_4187_0))) | (~i_13_462_1735_0 & ~i_13_462_2379_0 & ~i_13_462_2648_0 & ~i_13_462_4369_0) | (~i_13_462_1273_0 & i_13_462_4396_0));
endmodule



// Benchmark "kernel_13_463" written by ABC on Sun Jul 19 10:51:49 2020

module kernel_13_463 ( 
    i_13_463_76_0, i_13_463_105_0, i_13_463_112_0, i_13_463_184_0,
    i_13_463_186_0, i_13_463_193_0, i_13_463_195_0, i_13_463_327_0,
    i_13_463_445_0, i_13_463_510_0, i_13_463_562_0, i_13_463_573_0,
    i_13_463_574_0, i_13_463_579_0, i_13_463_626_0, i_13_463_646_0,
    i_13_463_666_0, i_13_463_697_0, i_13_463_717_0, i_13_463_780_0,
    i_13_463_854_0, i_13_463_861_0, i_13_463_894_0, i_13_463_949_0,
    i_13_463_958_0, i_13_463_994_0, i_13_463_1059_0, i_13_463_1084_0,
    i_13_463_1231_0, i_13_463_1258_0, i_13_463_1285_0, i_13_463_1321_0,
    i_13_463_1393_0, i_13_463_1407_0, i_13_463_1410_0, i_13_463_1483_0,
    i_13_463_1484_0, i_13_463_1488_0, i_13_463_1633_0, i_13_463_1677_0,
    i_13_463_1680_0, i_13_463_1690_0, i_13_463_1723_0, i_13_463_1749_0,
    i_13_463_1750_0, i_13_463_1752_0, i_13_463_1753_0, i_13_463_1788_0,
    i_13_463_1803_0, i_13_463_1804_0, i_13_463_1807_0, i_13_463_1858_0,
    i_13_463_1860_0, i_13_463_1861_0, i_13_463_2266_0, i_13_463_2310_0,
    i_13_463_2314_0, i_13_463_2519_0, i_13_463_2635_0, i_13_463_2652_0,
    i_13_463_2653_0, i_13_463_2673_0, i_13_463_2713_0, i_13_463_2715_0,
    i_13_463_2787_0, i_13_463_2850_0, i_13_463_2856_0, i_13_463_2857_0,
    i_13_463_2920_0, i_13_463_2983_0, i_13_463_3063_0, i_13_463_3144_0,
    i_13_463_3208_0, i_13_463_3309_0, i_13_463_3310_0, i_13_463_3372_0,
    i_13_463_3435_0, i_13_463_3451_0, i_13_463_3562_0, i_13_463_3595_0,
    i_13_463_3642_0, i_13_463_3685_0, i_13_463_3688_0, i_13_463_3739_0,
    i_13_463_3888_0, i_13_463_3909_0, i_13_463_3912_0, i_13_463_3913_0,
    i_13_463_3922_0, i_13_463_3938_0, i_13_463_3984_0, i_13_463_3994_0,
    i_13_463_4011_0, i_13_463_4012_0, i_13_463_4054_0, i_13_463_4077_0,
    i_13_463_4378_0, i_13_463_4443_0, i_13_463_4587_0, i_13_463_4591_0,
    o_13_463_0_0  );
  input  i_13_463_76_0, i_13_463_105_0, i_13_463_112_0, i_13_463_184_0,
    i_13_463_186_0, i_13_463_193_0, i_13_463_195_0, i_13_463_327_0,
    i_13_463_445_0, i_13_463_510_0, i_13_463_562_0, i_13_463_573_0,
    i_13_463_574_0, i_13_463_579_0, i_13_463_626_0, i_13_463_646_0,
    i_13_463_666_0, i_13_463_697_0, i_13_463_717_0, i_13_463_780_0,
    i_13_463_854_0, i_13_463_861_0, i_13_463_894_0, i_13_463_949_0,
    i_13_463_958_0, i_13_463_994_0, i_13_463_1059_0, i_13_463_1084_0,
    i_13_463_1231_0, i_13_463_1258_0, i_13_463_1285_0, i_13_463_1321_0,
    i_13_463_1393_0, i_13_463_1407_0, i_13_463_1410_0, i_13_463_1483_0,
    i_13_463_1484_0, i_13_463_1488_0, i_13_463_1633_0, i_13_463_1677_0,
    i_13_463_1680_0, i_13_463_1690_0, i_13_463_1723_0, i_13_463_1749_0,
    i_13_463_1750_0, i_13_463_1752_0, i_13_463_1753_0, i_13_463_1788_0,
    i_13_463_1803_0, i_13_463_1804_0, i_13_463_1807_0, i_13_463_1858_0,
    i_13_463_1860_0, i_13_463_1861_0, i_13_463_2266_0, i_13_463_2310_0,
    i_13_463_2314_0, i_13_463_2519_0, i_13_463_2635_0, i_13_463_2652_0,
    i_13_463_2653_0, i_13_463_2673_0, i_13_463_2713_0, i_13_463_2715_0,
    i_13_463_2787_0, i_13_463_2850_0, i_13_463_2856_0, i_13_463_2857_0,
    i_13_463_2920_0, i_13_463_2983_0, i_13_463_3063_0, i_13_463_3144_0,
    i_13_463_3208_0, i_13_463_3309_0, i_13_463_3310_0, i_13_463_3372_0,
    i_13_463_3435_0, i_13_463_3451_0, i_13_463_3562_0, i_13_463_3595_0,
    i_13_463_3642_0, i_13_463_3685_0, i_13_463_3688_0, i_13_463_3739_0,
    i_13_463_3888_0, i_13_463_3909_0, i_13_463_3912_0, i_13_463_3913_0,
    i_13_463_3922_0, i_13_463_3938_0, i_13_463_3984_0, i_13_463_3994_0,
    i_13_463_4011_0, i_13_463_4012_0, i_13_463_4054_0, i_13_463_4077_0,
    i_13_463_4378_0, i_13_463_4443_0, i_13_463_4587_0, i_13_463_4591_0;
  output o_13_463_0_0;
  assign o_13_463_0_0 = ~((~i_13_463_1750_0 & ((~i_13_463_1410_0 & ~i_13_463_1861_0 & ~i_13_463_2653_0) | (~i_13_463_1803_0 & ~i_13_463_1858_0 & i_13_463_2920_0))) | (~i_13_463_861_0 & i_13_463_1084_0) | (~i_13_463_894_0 & i_13_463_2673_0) | (i_13_463_697_0 & ~i_13_463_1803_0 & i_13_463_1858_0 & i_13_463_3595_0) | (~i_13_463_1861_0 & i_13_463_3685_0) | (~i_13_463_195_0 & ~i_13_463_574_0 & ~i_13_463_3994_0 & ~i_13_463_4077_0));
endmodule



// Benchmark "kernel_13_464" written by ABC on Sun Jul 19 10:51:49 2020

module kernel_13_464 ( 
    i_13_464_173_0, i_13_464_325_0, i_13_464_370_0, i_13_464_414_0,
    i_13_464_523_0, i_13_464_568_0, i_13_464_657_0, i_13_464_658_0,
    i_13_464_659_0, i_13_464_660_0, i_13_464_661_0, i_13_464_662_0,
    i_13_464_677_0, i_13_464_685_0, i_13_464_724_0, i_13_464_812_0,
    i_13_464_846_0, i_13_464_847_0, i_13_464_848_0, i_13_464_850_0,
    i_13_464_851_0, i_13_464_858_0, i_13_464_937_0, i_13_464_1017_0,
    i_13_464_1018_0, i_13_464_1073_0, i_13_464_1200_0, i_13_464_1225_0,
    i_13_464_1228_0, i_13_464_1305_0, i_13_464_1315_0, i_13_464_1345_0,
    i_13_464_1396_0, i_13_464_1454_0, i_13_464_1486_0, i_13_464_1549_0,
    i_13_464_1607_0, i_13_464_1630_0, i_13_464_1751_0, i_13_464_1764_0,
    i_13_464_1854_0, i_13_464_1855_0, i_13_464_1858_0, i_13_464_1926_0,
    i_13_464_1948_0, i_13_464_1954_0, i_13_464_1955_0, i_13_464_2197_0,
    i_13_464_2297_0, i_13_464_2417_0, i_13_464_2444_0, i_13_464_2448_0,
    i_13_464_2449_0, i_13_464_2541_0, i_13_464_2910_0, i_13_464_3006_0,
    i_13_464_3007_0, i_13_464_3061_0, i_13_464_3217_0, i_13_464_3235_0,
    i_13_464_3305_0, i_13_464_3370_0, i_13_464_3377_0, i_13_464_3414_0,
    i_13_464_3456_0, i_13_464_3457_0, i_13_464_3468_0, i_13_464_3475_0,
    i_13_464_3483_0, i_13_464_3484_0, i_13_464_3537_0, i_13_464_3538_0,
    i_13_464_3542_0, i_13_464_3557_0, i_13_464_3573_0, i_13_464_3574_0,
    i_13_464_3575_0, i_13_464_3647_0, i_13_464_3648_0, i_13_464_3727_0,
    i_13_464_3780_0, i_13_464_3852_0, i_13_464_3864_0, i_13_464_3892_0,
    i_13_464_3909_0, i_13_464_3929_0, i_13_464_4124_0, i_13_464_4249_0,
    i_13_464_4253_0, i_13_464_4257_0, i_13_464_4302_0, i_13_464_4338_0,
    i_13_464_4368_0, i_13_464_4369_0, i_13_464_4374_0, i_13_464_4375_0,
    i_13_464_4376_0, i_13_464_4458_0, i_13_464_4554_0, i_13_464_4595_0,
    o_13_464_0_0  );
  input  i_13_464_173_0, i_13_464_325_0, i_13_464_370_0, i_13_464_414_0,
    i_13_464_523_0, i_13_464_568_0, i_13_464_657_0, i_13_464_658_0,
    i_13_464_659_0, i_13_464_660_0, i_13_464_661_0, i_13_464_662_0,
    i_13_464_677_0, i_13_464_685_0, i_13_464_724_0, i_13_464_812_0,
    i_13_464_846_0, i_13_464_847_0, i_13_464_848_0, i_13_464_850_0,
    i_13_464_851_0, i_13_464_858_0, i_13_464_937_0, i_13_464_1017_0,
    i_13_464_1018_0, i_13_464_1073_0, i_13_464_1200_0, i_13_464_1225_0,
    i_13_464_1228_0, i_13_464_1305_0, i_13_464_1315_0, i_13_464_1345_0,
    i_13_464_1396_0, i_13_464_1454_0, i_13_464_1486_0, i_13_464_1549_0,
    i_13_464_1607_0, i_13_464_1630_0, i_13_464_1751_0, i_13_464_1764_0,
    i_13_464_1854_0, i_13_464_1855_0, i_13_464_1858_0, i_13_464_1926_0,
    i_13_464_1948_0, i_13_464_1954_0, i_13_464_1955_0, i_13_464_2197_0,
    i_13_464_2297_0, i_13_464_2417_0, i_13_464_2444_0, i_13_464_2448_0,
    i_13_464_2449_0, i_13_464_2541_0, i_13_464_2910_0, i_13_464_3006_0,
    i_13_464_3007_0, i_13_464_3061_0, i_13_464_3217_0, i_13_464_3235_0,
    i_13_464_3305_0, i_13_464_3370_0, i_13_464_3377_0, i_13_464_3414_0,
    i_13_464_3456_0, i_13_464_3457_0, i_13_464_3468_0, i_13_464_3475_0,
    i_13_464_3483_0, i_13_464_3484_0, i_13_464_3537_0, i_13_464_3538_0,
    i_13_464_3542_0, i_13_464_3557_0, i_13_464_3573_0, i_13_464_3574_0,
    i_13_464_3575_0, i_13_464_3647_0, i_13_464_3648_0, i_13_464_3727_0,
    i_13_464_3780_0, i_13_464_3852_0, i_13_464_3864_0, i_13_464_3892_0,
    i_13_464_3909_0, i_13_464_3929_0, i_13_464_4124_0, i_13_464_4249_0,
    i_13_464_4253_0, i_13_464_4257_0, i_13_464_4302_0, i_13_464_4338_0,
    i_13_464_4368_0, i_13_464_4369_0, i_13_464_4374_0, i_13_464_4375_0,
    i_13_464_4376_0, i_13_464_4458_0, i_13_464_4554_0, i_13_464_4595_0;
  output o_13_464_0_0;
  assign o_13_464_0_0 = ~((~i_13_464_1549_0 & ~i_13_464_4375_0) | (~i_13_464_3483_0 & ~i_13_464_3574_0));
endmodule



// Benchmark "kernel_13_465" written by ABC on Sun Jul 19 10:51:50 2020

module kernel_13_465 ( 
    i_13_465_22_0, i_13_465_48_0, i_13_465_59_0, i_13_465_68_0,
    i_13_465_94_0, i_13_465_112_0, i_13_465_165_0, i_13_465_195_0,
    i_13_465_202_0, i_13_465_237_0, i_13_465_238_0, i_13_465_255_0,
    i_13_465_274_0, i_13_465_283_0, i_13_465_309_0, i_13_465_333_0,
    i_13_465_336_0, i_13_465_337_0, i_13_465_383_0, i_13_465_454_0,
    i_13_465_585_0, i_13_465_586_0, i_13_465_588_0, i_13_465_615_0,
    i_13_465_620_0, i_13_465_665_0, i_13_465_771_0, i_13_465_781_0,
    i_13_465_833_0, i_13_465_856_0, i_13_465_980_0, i_13_465_1265_0,
    i_13_465_1310_0, i_13_465_1341_0, i_13_465_1342_0, i_13_465_1471_0,
    i_13_465_1488_0, i_13_465_1567_0, i_13_465_1670_0, i_13_465_1767_0,
    i_13_465_1803_0, i_13_465_1804_0, i_13_465_1931_0, i_13_465_1990_0,
    i_13_465_1992_0, i_13_465_2145_0, i_13_465_2179_0, i_13_465_2209_0,
    i_13_465_2376_0, i_13_465_2506_0, i_13_465_2535_0, i_13_465_2569_0,
    i_13_465_2571_0, i_13_465_2595_0, i_13_465_2678_0, i_13_465_2898_0,
    i_13_465_2903_0, i_13_465_2934_0, i_13_465_3016_0, i_13_465_3027_0,
    i_13_465_3028_0, i_13_465_3036_0, i_13_465_3037_0, i_13_465_3040_0,
    i_13_465_3122_0, i_13_465_3145_0, i_13_465_3210_0, i_13_465_3216_0,
    i_13_465_3220_0, i_13_465_3221_0, i_13_465_3285_0, i_13_465_3289_0,
    i_13_465_3315_0, i_13_465_3339_0, i_13_465_3342_0, i_13_465_3344_0,
    i_13_465_3393_0, i_13_465_3421_0, i_13_465_3468_0, i_13_465_3523_0,
    i_13_465_3599_0, i_13_465_3601_0, i_13_465_3639_0, i_13_465_3640_0,
    i_13_465_3643_0, i_13_465_3768_0, i_13_465_3784_0, i_13_465_3889_0,
    i_13_465_3982_0, i_13_465_4193_0, i_13_465_4230_0, i_13_465_4231_0,
    i_13_465_4315_0, i_13_465_4392_0, i_13_465_4408_0, i_13_465_4446_0,
    i_13_465_4512_0, i_13_465_4530_0, i_13_465_4534_0, i_13_465_4594_0,
    o_13_465_0_0  );
  input  i_13_465_22_0, i_13_465_48_0, i_13_465_59_0, i_13_465_68_0,
    i_13_465_94_0, i_13_465_112_0, i_13_465_165_0, i_13_465_195_0,
    i_13_465_202_0, i_13_465_237_0, i_13_465_238_0, i_13_465_255_0,
    i_13_465_274_0, i_13_465_283_0, i_13_465_309_0, i_13_465_333_0,
    i_13_465_336_0, i_13_465_337_0, i_13_465_383_0, i_13_465_454_0,
    i_13_465_585_0, i_13_465_586_0, i_13_465_588_0, i_13_465_615_0,
    i_13_465_620_0, i_13_465_665_0, i_13_465_771_0, i_13_465_781_0,
    i_13_465_833_0, i_13_465_856_0, i_13_465_980_0, i_13_465_1265_0,
    i_13_465_1310_0, i_13_465_1341_0, i_13_465_1342_0, i_13_465_1471_0,
    i_13_465_1488_0, i_13_465_1567_0, i_13_465_1670_0, i_13_465_1767_0,
    i_13_465_1803_0, i_13_465_1804_0, i_13_465_1931_0, i_13_465_1990_0,
    i_13_465_1992_0, i_13_465_2145_0, i_13_465_2179_0, i_13_465_2209_0,
    i_13_465_2376_0, i_13_465_2506_0, i_13_465_2535_0, i_13_465_2569_0,
    i_13_465_2571_0, i_13_465_2595_0, i_13_465_2678_0, i_13_465_2898_0,
    i_13_465_2903_0, i_13_465_2934_0, i_13_465_3016_0, i_13_465_3027_0,
    i_13_465_3028_0, i_13_465_3036_0, i_13_465_3037_0, i_13_465_3040_0,
    i_13_465_3122_0, i_13_465_3145_0, i_13_465_3210_0, i_13_465_3216_0,
    i_13_465_3220_0, i_13_465_3221_0, i_13_465_3285_0, i_13_465_3289_0,
    i_13_465_3315_0, i_13_465_3339_0, i_13_465_3342_0, i_13_465_3344_0,
    i_13_465_3393_0, i_13_465_3421_0, i_13_465_3468_0, i_13_465_3523_0,
    i_13_465_3599_0, i_13_465_3601_0, i_13_465_3639_0, i_13_465_3640_0,
    i_13_465_3643_0, i_13_465_3768_0, i_13_465_3784_0, i_13_465_3889_0,
    i_13_465_3982_0, i_13_465_4193_0, i_13_465_4230_0, i_13_465_4231_0,
    i_13_465_4315_0, i_13_465_4392_0, i_13_465_4408_0, i_13_465_4446_0,
    i_13_465_4512_0, i_13_465_4530_0, i_13_465_4534_0, i_13_465_4594_0;
  output o_13_465_0_0;
  assign o_13_465_0_0 = ~((~i_13_465_3315_0 & ((~i_13_465_3339_0 & ~i_13_465_3784_0) | (~i_13_465_1341_0 & ~i_13_465_3285_0 & ~i_13_465_4512_0))) | (~i_13_465_4392_0 & ((~i_13_465_94_0 & ~i_13_465_238_0 & ~i_13_465_2179_0) | (~i_13_465_2376_0 & ~i_13_465_3210_0 & ~i_13_465_4315_0))) | (i_13_465_238_0 & ~i_13_465_255_0) | (~i_13_465_1471_0 & ~i_13_465_3289_0 & ~i_13_465_3421_0 & i_13_465_4512_0));
endmodule



// Benchmark "kernel_13_466" written by ABC on Sun Jul 19 10:51:51 2020

module kernel_13_466 ( 
    i_13_466_20_0, i_13_466_65_0, i_13_466_121_0, i_13_466_207_0,
    i_13_466_208_0, i_13_466_211_0, i_13_466_265_0, i_13_466_266_0,
    i_13_466_373_0, i_13_466_384_0, i_13_466_414_0, i_13_466_415_0,
    i_13_466_423_0, i_13_466_503_0, i_13_466_521_0, i_13_466_522_0,
    i_13_466_664_0, i_13_466_715_0, i_13_466_746_0, i_13_466_763_0,
    i_13_466_764_0, i_13_466_833_0, i_13_466_849_0, i_13_466_850_0,
    i_13_466_852_0, i_13_466_982_0, i_13_466_1081_0, i_13_466_1084_0,
    i_13_466_1131_0, i_13_466_1133_0, i_13_466_1151_0, i_13_466_1200_0,
    i_13_466_1219_0, i_13_466_1309_0, i_13_466_1312_0, i_13_466_1397_0,
    i_13_466_1436_0, i_13_466_1467_0, i_13_466_1522_0, i_13_466_1549_0,
    i_13_466_1550_0, i_13_466_1551_0, i_13_466_1552_0, i_13_466_1599_0,
    i_13_466_1604_0, i_13_466_1630_0, i_13_466_1723_0, i_13_466_1732_0,
    i_13_466_1750_0, i_13_466_1751_0, i_13_466_1952_0, i_13_466_1999_0,
    i_13_466_2048_0, i_13_466_2121_0, i_13_466_2125_0, i_13_466_2295_0,
    i_13_466_2434_0, i_13_466_2709_0, i_13_466_2723_0, i_13_466_3087_0,
    i_13_466_3088_0, i_13_466_3100_0, i_13_466_3125_0, i_13_466_3163_0,
    i_13_466_3271_0, i_13_466_3289_0, i_13_466_3345_0, i_13_466_3346_0,
    i_13_466_3383_0, i_13_466_3405_0, i_13_466_3414_0, i_13_466_3423_0,
    i_13_466_3483_0, i_13_466_3486_0, i_13_466_3524_0, i_13_466_3537_0,
    i_13_466_3538_0, i_13_466_3539_0, i_13_466_3541_0, i_13_466_3542_0,
    i_13_466_3619_0, i_13_466_3666_0, i_13_466_3667_0, i_13_466_3726_0,
    i_13_466_3728_0, i_13_466_3765_0, i_13_466_3798_0, i_13_466_3843_0,
    i_13_466_3906_0, i_13_466_3920_0, i_13_466_3985_0, i_13_466_4038_0,
    i_13_466_4039_0, i_13_466_4059_0, i_13_466_4204_0, i_13_466_4256_0,
    i_13_466_4336_0, i_13_466_4378_0, i_13_466_4447_0, i_13_466_4523_0,
    o_13_466_0_0  );
  input  i_13_466_20_0, i_13_466_65_0, i_13_466_121_0, i_13_466_207_0,
    i_13_466_208_0, i_13_466_211_0, i_13_466_265_0, i_13_466_266_0,
    i_13_466_373_0, i_13_466_384_0, i_13_466_414_0, i_13_466_415_0,
    i_13_466_423_0, i_13_466_503_0, i_13_466_521_0, i_13_466_522_0,
    i_13_466_664_0, i_13_466_715_0, i_13_466_746_0, i_13_466_763_0,
    i_13_466_764_0, i_13_466_833_0, i_13_466_849_0, i_13_466_850_0,
    i_13_466_852_0, i_13_466_982_0, i_13_466_1081_0, i_13_466_1084_0,
    i_13_466_1131_0, i_13_466_1133_0, i_13_466_1151_0, i_13_466_1200_0,
    i_13_466_1219_0, i_13_466_1309_0, i_13_466_1312_0, i_13_466_1397_0,
    i_13_466_1436_0, i_13_466_1467_0, i_13_466_1522_0, i_13_466_1549_0,
    i_13_466_1550_0, i_13_466_1551_0, i_13_466_1552_0, i_13_466_1599_0,
    i_13_466_1604_0, i_13_466_1630_0, i_13_466_1723_0, i_13_466_1732_0,
    i_13_466_1750_0, i_13_466_1751_0, i_13_466_1952_0, i_13_466_1999_0,
    i_13_466_2048_0, i_13_466_2121_0, i_13_466_2125_0, i_13_466_2295_0,
    i_13_466_2434_0, i_13_466_2709_0, i_13_466_2723_0, i_13_466_3087_0,
    i_13_466_3088_0, i_13_466_3100_0, i_13_466_3125_0, i_13_466_3163_0,
    i_13_466_3271_0, i_13_466_3289_0, i_13_466_3345_0, i_13_466_3346_0,
    i_13_466_3383_0, i_13_466_3405_0, i_13_466_3414_0, i_13_466_3423_0,
    i_13_466_3483_0, i_13_466_3486_0, i_13_466_3524_0, i_13_466_3537_0,
    i_13_466_3538_0, i_13_466_3539_0, i_13_466_3541_0, i_13_466_3542_0,
    i_13_466_3619_0, i_13_466_3666_0, i_13_466_3667_0, i_13_466_3726_0,
    i_13_466_3728_0, i_13_466_3765_0, i_13_466_3798_0, i_13_466_3843_0,
    i_13_466_3906_0, i_13_466_3920_0, i_13_466_3985_0, i_13_466_4038_0,
    i_13_466_4039_0, i_13_466_4059_0, i_13_466_4204_0, i_13_466_4256_0,
    i_13_466_4336_0, i_13_466_4378_0, i_13_466_4447_0, i_13_466_4523_0;
  output o_13_466_0_0;
  assign o_13_466_0_0 = ~((~i_13_466_4038_0 & ((~i_13_466_415_0 & ~i_13_466_3542_0) | (~i_13_466_3920_0 & i_13_466_3985_0))) | (i_13_466_1732_0 & ~i_13_466_1750_0) | (~i_13_466_384_0 & ~i_13_466_764_0 & ~i_13_466_1549_0 & ~i_13_466_1550_0 & ~i_13_466_3537_0) | (i_13_466_3289_0 & i_13_466_4038_0) | (i_13_466_2434_0 & i_13_466_4039_0));
endmodule



// Benchmark "kernel_13_467" written by ABC on Sun Jul 19 10:51:52 2020

module kernel_13_467 ( 
    i_13_467_56_0, i_13_467_131_0, i_13_467_166_0, i_13_467_187_0,
    i_13_467_202_0, i_13_467_211_0, i_13_467_284_0, i_13_467_319_0,
    i_13_467_355_0, i_13_467_365_0, i_13_467_392_0, i_13_467_520_0,
    i_13_467_521_0, i_13_467_527_0, i_13_467_545_0, i_13_467_563_0,
    i_13_467_589_0, i_13_467_616_0, i_13_467_652_0, i_13_467_688_0,
    i_13_467_833_0, i_13_467_1003_0, i_13_467_1066_0, i_13_467_1067_0,
    i_13_467_1069_0, i_13_467_1075_0, i_13_467_1108_0, i_13_467_1112_0,
    i_13_467_1129_0, i_13_467_1225_0, i_13_467_1278_0, i_13_467_1391_0,
    i_13_467_1454_0, i_13_467_1498_0, i_13_467_1523_0, i_13_467_1534_0,
    i_13_467_1598_0, i_13_467_1669_0, i_13_467_1687_0, i_13_467_1717_0,
    i_13_467_1723_0, i_13_467_1771_0, i_13_467_1781_0, i_13_467_1799_0,
    i_13_467_1930_0, i_13_467_1975_0, i_13_467_1984_0, i_13_467_1993_0,
    i_13_467_2023_0, i_13_467_2024_0, i_13_467_2087_0, i_13_467_2102_0,
    i_13_467_2137_0, i_13_467_2173_0, i_13_467_2200_0, i_13_467_2362_0,
    i_13_467_2363_0, i_13_467_2371_0, i_13_467_2386_0, i_13_467_2393_0,
    i_13_467_2425_0, i_13_467_2572_0, i_13_467_2606_0, i_13_467_2615_0,
    i_13_467_2618_0, i_13_467_2654_0, i_13_467_2681_0, i_13_467_2785_0,
    i_13_467_2815_0, i_13_467_2888_0, i_13_467_2969_0, i_13_467_2971_0,
    i_13_467_2974_0, i_13_467_3014_0, i_13_467_3032_0, i_13_467_3056_0,
    i_13_467_3181_0, i_13_467_3209_0, i_13_467_3212_0, i_13_467_3266_0,
    i_13_467_3487_0, i_13_467_3730_0, i_13_467_3778_0, i_13_467_3823_0,
    i_13_467_3901_0, i_13_467_3938_0, i_13_467_3941_0, i_13_467_4015_0,
    i_13_467_4031_0, i_13_467_4159_0, i_13_467_4165_0, i_13_467_4166_0,
    i_13_467_4225_0, i_13_467_4369_0, i_13_467_4373_0, i_13_467_4384_0,
    i_13_467_4451_0, i_13_467_4496_0, i_13_467_4507_0, i_13_467_4517_0,
    o_13_467_0_0  );
  input  i_13_467_56_0, i_13_467_131_0, i_13_467_166_0, i_13_467_187_0,
    i_13_467_202_0, i_13_467_211_0, i_13_467_284_0, i_13_467_319_0,
    i_13_467_355_0, i_13_467_365_0, i_13_467_392_0, i_13_467_520_0,
    i_13_467_521_0, i_13_467_527_0, i_13_467_545_0, i_13_467_563_0,
    i_13_467_589_0, i_13_467_616_0, i_13_467_652_0, i_13_467_688_0,
    i_13_467_833_0, i_13_467_1003_0, i_13_467_1066_0, i_13_467_1067_0,
    i_13_467_1069_0, i_13_467_1075_0, i_13_467_1108_0, i_13_467_1112_0,
    i_13_467_1129_0, i_13_467_1225_0, i_13_467_1278_0, i_13_467_1391_0,
    i_13_467_1454_0, i_13_467_1498_0, i_13_467_1523_0, i_13_467_1534_0,
    i_13_467_1598_0, i_13_467_1669_0, i_13_467_1687_0, i_13_467_1717_0,
    i_13_467_1723_0, i_13_467_1771_0, i_13_467_1781_0, i_13_467_1799_0,
    i_13_467_1930_0, i_13_467_1975_0, i_13_467_1984_0, i_13_467_1993_0,
    i_13_467_2023_0, i_13_467_2024_0, i_13_467_2087_0, i_13_467_2102_0,
    i_13_467_2137_0, i_13_467_2173_0, i_13_467_2200_0, i_13_467_2362_0,
    i_13_467_2363_0, i_13_467_2371_0, i_13_467_2386_0, i_13_467_2393_0,
    i_13_467_2425_0, i_13_467_2572_0, i_13_467_2606_0, i_13_467_2615_0,
    i_13_467_2618_0, i_13_467_2654_0, i_13_467_2681_0, i_13_467_2785_0,
    i_13_467_2815_0, i_13_467_2888_0, i_13_467_2969_0, i_13_467_2971_0,
    i_13_467_2974_0, i_13_467_3014_0, i_13_467_3032_0, i_13_467_3056_0,
    i_13_467_3181_0, i_13_467_3209_0, i_13_467_3212_0, i_13_467_3266_0,
    i_13_467_3487_0, i_13_467_3730_0, i_13_467_3778_0, i_13_467_3823_0,
    i_13_467_3901_0, i_13_467_3938_0, i_13_467_3941_0, i_13_467_4015_0,
    i_13_467_4031_0, i_13_467_4159_0, i_13_467_4165_0, i_13_467_4166_0,
    i_13_467_4225_0, i_13_467_4369_0, i_13_467_4373_0, i_13_467_4384_0,
    i_13_467_4451_0, i_13_467_4496_0, i_13_467_4507_0, i_13_467_4517_0;
  output o_13_467_0_0;
  assign o_13_467_0_0 = 0;
endmodule



// Benchmark "kernel_13_468" written by ABC on Sun Jul 19 10:51:52 2020

module kernel_13_468 ( 
    i_13_468_45_0, i_13_468_46_0, i_13_468_79_0, i_13_468_121_0,
    i_13_468_122_0, i_13_468_173_0, i_13_468_184_0, i_13_468_226_0,
    i_13_468_238_0, i_13_468_313_0, i_13_468_337_0, i_13_468_408_0,
    i_13_468_444_0, i_13_468_518_0, i_13_468_523_0, i_13_468_533_0,
    i_13_468_554_0, i_13_468_649_0, i_13_468_684_0, i_13_468_723_0,
    i_13_468_734_0, i_13_468_760_0, i_13_468_848_0, i_13_468_922_0,
    i_13_468_938_0, i_13_468_976_0, i_13_468_1017_0, i_13_468_1031_0,
    i_13_468_1071_0, i_13_468_1073_0, i_13_468_1101_0, i_13_468_1136_0,
    i_13_468_1148_0, i_13_468_1207_0, i_13_468_1225_0, i_13_468_1301_0,
    i_13_468_1306_0, i_13_468_1315_0, i_13_468_1372_0, i_13_468_1389_0,
    i_13_468_1427_0, i_13_468_1444_0, i_13_468_1445_0, i_13_468_1510_0,
    i_13_468_1549_0, i_13_468_1720_0, i_13_468_1728_0, i_13_468_1859_0,
    i_13_468_1945_0, i_13_468_2026_0, i_13_468_2027_0, i_13_468_2045_0,
    i_13_468_2126_0, i_13_468_2197_0, i_13_468_2198_0, i_13_468_2209_0,
    i_13_468_2262_0, i_13_468_2448_0, i_13_468_2469_0, i_13_468_2705_0,
    i_13_468_2763_0, i_13_468_2852_0, i_13_468_2918_0, i_13_468_3006_0,
    i_13_468_3007_0, i_13_468_3027_0, i_13_468_3128_0, i_13_468_3217_0,
    i_13_468_3218_0, i_13_468_3227_0, i_13_468_3235_0, i_13_468_3457_0,
    i_13_468_3458_0, i_13_468_3484_0, i_13_468_3485_0, i_13_468_3575_0,
    i_13_468_3781_0, i_13_468_3782_0, i_13_468_3800_0, i_13_468_3853_0,
    i_13_468_3915_0, i_13_468_3983_0, i_13_468_3990_0, i_13_468_4017_0,
    i_13_468_4080_0, i_13_468_4150_0, i_13_468_4193_0, i_13_468_4234_0,
    i_13_468_4249_0, i_13_468_4250_0, i_13_468_4258_0, i_13_468_4259_0,
    i_13_468_4262_0, i_13_468_4301_0, i_13_468_4369_0, i_13_468_4376_0,
    i_13_468_4447_0, i_13_468_4448_0, i_13_468_4593_0, i_13_468_4604_0,
    o_13_468_0_0  );
  input  i_13_468_45_0, i_13_468_46_0, i_13_468_79_0, i_13_468_121_0,
    i_13_468_122_0, i_13_468_173_0, i_13_468_184_0, i_13_468_226_0,
    i_13_468_238_0, i_13_468_313_0, i_13_468_337_0, i_13_468_408_0,
    i_13_468_444_0, i_13_468_518_0, i_13_468_523_0, i_13_468_533_0,
    i_13_468_554_0, i_13_468_649_0, i_13_468_684_0, i_13_468_723_0,
    i_13_468_734_0, i_13_468_760_0, i_13_468_848_0, i_13_468_922_0,
    i_13_468_938_0, i_13_468_976_0, i_13_468_1017_0, i_13_468_1031_0,
    i_13_468_1071_0, i_13_468_1073_0, i_13_468_1101_0, i_13_468_1136_0,
    i_13_468_1148_0, i_13_468_1207_0, i_13_468_1225_0, i_13_468_1301_0,
    i_13_468_1306_0, i_13_468_1315_0, i_13_468_1372_0, i_13_468_1389_0,
    i_13_468_1427_0, i_13_468_1444_0, i_13_468_1445_0, i_13_468_1510_0,
    i_13_468_1549_0, i_13_468_1720_0, i_13_468_1728_0, i_13_468_1859_0,
    i_13_468_1945_0, i_13_468_2026_0, i_13_468_2027_0, i_13_468_2045_0,
    i_13_468_2126_0, i_13_468_2197_0, i_13_468_2198_0, i_13_468_2209_0,
    i_13_468_2262_0, i_13_468_2448_0, i_13_468_2469_0, i_13_468_2705_0,
    i_13_468_2763_0, i_13_468_2852_0, i_13_468_2918_0, i_13_468_3006_0,
    i_13_468_3007_0, i_13_468_3027_0, i_13_468_3128_0, i_13_468_3217_0,
    i_13_468_3218_0, i_13_468_3227_0, i_13_468_3235_0, i_13_468_3457_0,
    i_13_468_3458_0, i_13_468_3484_0, i_13_468_3485_0, i_13_468_3575_0,
    i_13_468_3781_0, i_13_468_3782_0, i_13_468_3800_0, i_13_468_3853_0,
    i_13_468_3915_0, i_13_468_3983_0, i_13_468_3990_0, i_13_468_4017_0,
    i_13_468_4080_0, i_13_468_4150_0, i_13_468_4193_0, i_13_468_4234_0,
    i_13_468_4249_0, i_13_468_4250_0, i_13_468_4258_0, i_13_468_4259_0,
    i_13_468_4262_0, i_13_468_4301_0, i_13_468_4369_0, i_13_468_4376_0,
    i_13_468_4447_0, i_13_468_4448_0, i_13_468_4593_0, i_13_468_4604_0;
  output o_13_468_0_0;
  assign o_13_468_0_0 = ~(~i_13_468_3484_0 | (~i_13_468_2026_0 & ~i_13_468_4448_0) | (i_13_468_684_0 & ~i_13_468_4369_0) | (i_13_468_734_0 & ~i_13_468_938_0));
endmodule



// Benchmark "kernel_13_469" written by ABC on Sun Jul 19 10:51:53 2020

module kernel_13_469 ( 
    i_13_469_90_0, i_13_469_91_0, i_13_469_130_0, i_13_469_141_0,
    i_13_469_172_0, i_13_469_370_0, i_13_469_389_0, i_13_469_423_0,
    i_13_469_430_0, i_13_469_450_0, i_13_469_553_0, i_13_469_585_0,
    i_13_469_657_0, i_13_469_660_0, i_13_469_688_0, i_13_469_726_0,
    i_13_469_828_0, i_13_469_829_0, i_13_469_831_0, i_13_469_933_0,
    i_13_469_934_0, i_13_469_955_0, i_13_469_1063_0, i_13_469_1066_0,
    i_13_469_1075_0, i_13_469_1096_0, i_13_469_1116_0, i_13_469_1147_0,
    i_13_469_1224_0, i_13_469_1306_0, i_13_469_1324_0, i_13_469_1428_0,
    i_13_469_1471_0, i_13_469_1488_0, i_13_469_1494_0, i_13_469_1510_0,
    i_13_469_1552_0, i_13_469_1570_0, i_13_469_1696_0, i_13_469_1697_0,
    i_13_469_1726_0, i_13_469_1764_0, i_13_469_1786_0, i_13_469_1801_0,
    i_13_469_1846_0, i_13_469_1887_0, i_13_469_1892_0, i_13_469_1926_0,
    i_13_469_1927_0, i_13_469_1957_0, i_13_469_2044_0, i_13_469_2107_0,
    i_13_469_2119_0, i_13_469_2142_0, i_13_469_2143_0, i_13_469_2175_0,
    i_13_469_2265_0, i_13_469_2266_0, i_13_469_2296_0, i_13_469_2461_0,
    i_13_469_2877_0, i_13_469_2935_0, i_13_469_2938_0, i_13_469_3006_0,
    i_13_469_3016_0, i_13_469_3039_0, i_13_469_3043_0, i_13_469_3064_0,
    i_13_469_3225_0, i_13_469_3231_0, i_13_469_3241_0, i_13_469_3264_0,
    i_13_469_3274_0, i_13_469_3454_0, i_13_469_3457_0, i_13_469_3487_0,
    i_13_469_3523_0, i_13_469_3538_0, i_13_469_3637_0, i_13_469_3645_0,
    i_13_469_3742_0, i_13_469_3753_0, i_13_469_3754_0, i_13_469_3856_0,
    i_13_469_3916_0, i_13_469_3979_0, i_13_469_4018_0, i_13_469_4267_0,
    i_13_469_4268_0, i_13_469_4308_0, i_13_469_4312_0, i_13_469_4341_0,
    i_13_469_4368_0, i_13_469_4369_0, i_13_469_4429_0, i_13_469_4509_0,
    i_13_469_4510_0, i_13_469_4511_0, i_13_469_4524_0, i_13_469_4567_0,
    o_13_469_0_0  );
  input  i_13_469_90_0, i_13_469_91_0, i_13_469_130_0, i_13_469_141_0,
    i_13_469_172_0, i_13_469_370_0, i_13_469_389_0, i_13_469_423_0,
    i_13_469_430_0, i_13_469_450_0, i_13_469_553_0, i_13_469_585_0,
    i_13_469_657_0, i_13_469_660_0, i_13_469_688_0, i_13_469_726_0,
    i_13_469_828_0, i_13_469_829_0, i_13_469_831_0, i_13_469_933_0,
    i_13_469_934_0, i_13_469_955_0, i_13_469_1063_0, i_13_469_1066_0,
    i_13_469_1075_0, i_13_469_1096_0, i_13_469_1116_0, i_13_469_1147_0,
    i_13_469_1224_0, i_13_469_1306_0, i_13_469_1324_0, i_13_469_1428_0,
    i_13_469_1471_0, i_13_469_1488_0, i_13_469_1494_0, i_13_469_1510_0,
    i_13_469_1552_0, i_13_469_1570_0, i_13_469_1696_0, i_13_469_1697_0,
    i_13_469_1726_0, i_13_469_1764_0, i_13_469_1786_0, i_13_469_1801_0,
    i_13_469_1846_0, i_13_469_1887_0, i_13_469_1892_0, i_13_469_1926_0,
    i_13_469_1927_0, i_13_469_1957_0, i_13_469_2044_0, i_13_469_2107_0,
    i_13_469_2119_0, i_13_469_2142_0, i_13_469_2143_0, i_13_469_2175_0,
    i_13_469_2265_0, i_13_469_2266_0, i_13_469_2296_0, i_13_469_2461_0,
    i_13_469_2877_0, i_13_469_2935_0, i_13_469_2938_0, i_13_469_3006_0,
    i_13_469_3016_0, i_13_469_3039_0, i_13_469_3043_0, i_13_469_3064_0,
    i_13_469_3225_0, i_13_469_3231_0, i_13_469_3241_0, i_13_469_3264_0,
    i_13_469_3274_0, i_13_469_3454_0, i_13_469_3457_0, i_13_469_3487_0,
    i_13_469_3523_0, i_13_469_3538_0, i_13_469_3637_0, i_13_469_3645_0,
    i_13_469_3742_0, i_13_469_3753_0, i_13_469_3754_0, i_13_469_3856_0,
    i_13_469_3916_0, i_13_469_3979_0, i_13_469_4018_0, i_13_469_4267_0,
    i_13_469_4268_0, i_13_469_4308_0, i_13_469_4312_0, i_13_469_4341_0,
    i_13_469_4368_0, i_13_469_4369_0, i_13_469_4429_0, i_13_469_4509_0,
    i_13_469_4510_0, i_13_469_4511_0, i_13_469_4524_0, i_13_469_4567_0;
  output o_13_469_0_0;
  assign o_13_469_0_0 = ~((i_13_469_4511_0 & (~i_13_469_1552_0 | ~i_13_469_4312_0 | (~i_13_469_1075_0 & ~i_13_469_2935_0))) | ~i_13_469_3754_0 | (~i_13_469_1846_0 & ~i_13_469_4368_0 & ~i_13_469_4429_0) | (~i_13_469_3457_0 & ~i_13_469_4268_0 & ~i_13_469_4509_0));
endmodule



// Benchmark "kernel_13_470" written by ABC on Sun Jul 19 10:51:54 2020

module kernel_13_470 ( 
    i_13_470_51_0, i_13_470_124_0, i_13_470_186_0, i_13_470_229_0,
    i_13_470_250_0, i_13_470_258_0, i_13_470_276_0, i_13_470_277_0,
    i_13_470_309_0, i_13_470_375_0, i_13_470_376_0, i_13_470_420_0,
    i_13_470_430_0, i_13_470_561_0, i_13_470_588_0, i_13_470_618_0,
    i_13_470_619_0, i_13_470_642_0, i_13_470_654_0, i_13_470_672_0,
    i_13_470_699_0, i_13_470_738_0, i_13_470_771_0, i_13_470_823_0,
    i_13_470_840_0, i_13_470_942_0, i_13_470_979_0, i_13_470_1065_0,
    i_13_470_1069_0, i_13_470_1077_0, i_13_470_1078_0, i_13_470_1218_0,
    i_13_470_1230_0, i_13_470_1297_0, i_13_470_1327_0, i_13_470_1329_0,
    i_13_470_1443_0, i_13_470_1528_0, i_13_470_1569_0, i_13_470_1572_0,
    i_13_470_1596_0, i_13_470_1734_0, i_13_470_1735_0, i_13_470_1834_0,
    i_13_470_1852_0, i_13_470_1992_0, i_13_470_2002_0, i_13_470_2107_0,
    i_13_470_2185_0, i_13_470_2229_0, i_13_470_2230_0, i_13_470_2302_0,
    i_13_470_2313_0, i_13_470_2314_0, i_13_470_2362_0, i_13_470_2454_0,
    i_13_470_2572_0, i_13_470_2581_0, i_13_470_2694_0, i_13_470_2697_0,
    i_13_470_2742_0, i_13_470_2752_0, i_13_470_2769_0, i_13_470_2886_0,
    i_13_470_2887_0, i_13_470_2922_0, i_13_470_2958_0, i_13_470_2967_0,
    i_13_470_3006_0, i_13_470_3291_0, i_13_470_3315_0, i_13_470_3372_0,
    i_13_470_3522_0, i_13_470_3525_0, i_13_470_3549_0, i_13_470_3552_0,
    i_13_470_3553_0, i_13_470_3603_0, i_13_470_3612_0, i_13_470_3687_0,
    i_13_470_3714_0, i_13_470_3729_0, i_13_470_3730_0, i_13_470_3733_0,
    i_13_470_3748_0, i_13_470_3817_0, i_13_470_3822_0, i_13_470_3885_0,
    i_13_470_3903_0, i_13_470_3904_0, i_13_470_4047_0, i_13_470_4089_0,
    i_13_470_4164_0, i_13_470_4236_0, i_13_470_4282_0, i_13_470_4332_0,
    i_13_470_4387_0, i_13_470_4390_0, i_13_470_4461_0, i_13_470_4603_0,
    o_13_470_0_0  );
  input  i_13_470_51_0, i_13_470_124_0, i_13_470_186_0, i_13_470_229_0,
    i_13_470_250_0, i_13_470_258_0, i_13_470_276_0, i_13_470_277_0,
    i_13_470_309_0, i_13_470_375_0, i_13_470_376_0, i_13_470_420_0,
    i_13_470_430_0, i_13_470_561_0, i_13_470_588_0, i_13_470_618_0,
    i_13_470_619_0, i_13_470_642_0, i_13_470_654_0, i_13_470_672_0,
    i_13_470_699_0, i_13_470_738_0, i_13_470_771_0, i_13_470_823_0,
    i_13_470_840_0, i_13_470_942_0, i_13_470_979_0, i_13_470_1065_0,
    i_13_470_1069_0, i_13_470_1077_0, i_13_470_1078_0, i_13_470_1218_0,
    i_13_470_1230_0, i_13_470_1297_0, i_13_470_1327_0, i_13_470_1329_0,
    i_13_470_1443_0, i_13_470_1528_0, i_13_470_1569_0, i_13_470_1572_0,
    i_13_470_1596_0, i_13_470_1734_0, i_13_470_1735_0, i_13_470_1834_0,
    i_13_470_1852_0, i_13_470_1992_0, i_13_470_2002_0, i_13_470_2107_0,
    i_13_470_2185_0, i_13_470_2229_0, i_13_470_2230_0, i_13_470_2302_0,
    i_13_470_2313_0, i_13_470_2314_0, i_13_470_2362_0, i_13_470_2454_0,
    i_13_470_2572_0, i_13_470_2581_0, i_13_470_2694_0, i_13_470_2697_0,
    i_13_470_2742_0, i_13_470_2752_0, i_13_470_2769_0, i_13_470_2886_0,
    i_13_470_2887_0, i_13_470_2922_0, i_13_470_2958_0, i_13_470_2967_0,
    i_13_470_3006_0, i_13_470_3291_0, i_13_470_3315_0, i_13_470_3372_0,
    i_13_470_3522_0, i_13_470_3525_0, i_13_470_3549_0, i_13_470_3552_0,
    i_13_470_3553_0, i_13_470_3603_0, i_13_470_3612_0, i_13_470_3687_0,
    i_13_470_3714_0, i_13_470_3729_0, i_13_470_3730_0, i_13_470_3733_0,
    i_13_470_3748_0, i_13_470_3817_0, i_13_470_3822_0, i_13_470_3885_0,
    i_13_470_3903_0, i_13_470_3904_0, i_13_470_4047_0, i_13_470_4089_0,
    i_13_470_4164_0, i_13_470_4236_0, i_13_470_4282_0, i_13_470_4332_0,
    i_13_470_4387_0, i_13_470_4390_0, i_13_470_4461_0, i_13_470_4603_0;
  output o_13_470_0_0;
  assign o_13_470_0_0 = ~((~i_13_470_2742_0 & (~i_13_470_654_0 | (~i_13_470_51_0 & ~i_13_470_618_0 & ~i_13_470_3903_0))) | (~i_13_470_2302_0 & ((i_13_470_4236_0 & (~i_13_470_699_0 | ~i_13_470_3315_0)) | (i_13_470_1065_0 & ~i_13_470_3553_0))) | (~i_13_470_840_0 & ~i_13_470_2697_0 & ~i_13_470_3904_0) | (~i_13_470_1834_0 & ~i_13_470_4047_0));
endmodule



// Benchmark "kernel_13_471" written by ABC on Sun Jul 19 10:51:55 2020

module kernel_13_471 ( 
    i_13_471_49_0, i_13_471_66_0, i_13_471_133_0, i_13_471_195_0,
    i_13_471_327_0, i_13_471_381_0, i_13_471_483_0, i_13_471_528_0,
    i_13_471_529_0, i_13_471_673_0, i_13_471_717_0, i_13_471_799_0,
    i_13_471_842_0, i_13_471_844_0, i_13_471_861_0, i_13_471_951_0,
    i_13_471_1204_0, i_13_471_1222_0, i_13_471_1228_0, i_13_471_1230_0,
    i_13_471_1257_0, i_13_471_1258_0, i_13_471_1302_0, i_13_471_1320_0,
    i_13_471_1326_0, i_13_471_1384_0, i_13_471_1428_0, i_13_471_1437_0,
    i_13_471_1446_0, i_13_471_1491_0, i_13_471_1492_0, i_13_471_1501_0,
    i_13_471_1554_0, i_13_471_1555_0, i_13_471_1556_0, i_13_471_1699_0,
    i_13_471_1722_0, i_13_471_1795_0, i_13_471_1834_0, i_13_471_1884_0,
    i_13_471_1902_0, i_13_471_1930_0, i_13_471_1941_0, i_13_471_1960_0,
    i_13_471_2002_0, i_13_471_2005_0, i_13_471_2014_0, i_13_471_2033_0,
    i_13_471_2103_0, i_13_471_2128_0, i_13_471_2139_0, i_13_471_2148_0,
    i_13_471_2202_0, i_13_471_2203_0, i_13_471_2299_0, i_13_471_2302_0,
    i_13_471_2446_0, i_13_471_2535_0, i_13_471_2722_0, i_13_471_2743_0,
    i_13_471_2850_0, i_13_471_2937_0, i_13_471_2938_0, i_13_471_3027_0,
    i_13_471_3136_0, i_13_471_3174_0, i_13_471_3238_0, i_13_471_3244_0,
    i_13_471_3309_0, i_13_471_3310_0, i_13_471_3423_0, i_13_471_3445_0,
    i_13_471_3525_0, i_13_471_3543_0, i_13_471_3552_0, i_13_471_3597_0,
    i_13_471_3616_0, i_13_471_3706_0, i_13_471_3731_0, i_13_471_3732_0,
    i_13_471_3786_0, i_13_471_3805_0, i_13_471_3831_0, i_13_471_3849_0,
    i_13_471_3858_0, i_13_471_3859_0, i_13_471_3912_0, i_13_471_3913_0,
    i_13_471_3994_0, i_13_471_4011_0, i_13_471_4012_0, i_13_471_4117_0,
    i_13_471_4161_0, i_13_471_4254_0, i_13_471_4369_0, i_13_471_4380_0,
    i_13_471_4381_0, i_13_471_4443_0, i_13_471_4587_0, i_13_471_4588_0,
    o_13_471_0_0  );
  input  i_13_471_49_0, i_13_471_66_0, i_13_471_133_0, i_13_471_195_0,
    i_13_471_327_0, i_13_471_381_0, i_13_471_483_0, i_13_471_528_0,
    i_13_471_529_0, i_13_471_673_0, i_13_471_717_0, i_13_471_799_0,
    i_13_471_842_0, i_13_471_844_0, i_13_471_861_0, i_13_471_951_0,
    i_13_471_1204_0, i_13_471_1222_0, i_13_471_1228_0, i_13_471_1230_0,
    i_13_471_1257_0, i_13_471_1258_0, i_13_471_1302_0, i_13_471_1320_0,
    i_13_471_1326_0, i_13_471_1384_0, i_13_471_1428_0, i_13_471_1437_0,
    i_13_471_1446_0, i_13_471_1491_0, i_13_471_1492_0, i_13_471_1501_0,
    i_13_471_1554_0, i_13_471_1555_0, i_13_471_1556_0, i_13_471_1699_0,
    i_13_471_1722_0, i_13_471_1795_0, i_13_471_1834_0, i_13_471_1884_0,
    i_13_471_1902_0, i_13_471_1930_0, i_13_471_1941_0, i_13_471_1960_0,
    i_13_471_2002_0, i_13_471_2005_0, i_13_471_2014_0, i_13_471_2033_0,
    i_13_471_2103_0, i_13_471_2128_0, i_13_471_2139_0, i_13_471_2148_0,
    i_13_471_2202_0, i_13_471_2203_0, i_13_471_2299_0, i_13_471_2302_0,
    i_13_471_2446_0, i_13_471_2535_0, i_13_471_2722_0, i_13_471_2743_0,
    i_13_471_2850_0, i_13_471_2937_0, i_13_471_2938_0, i_13_471_3027_0,
    i_13_471_3136_0, i_13_471_3174_0, i_13_471_3238_0, i_13_471_3244_0,
    i_13_471_3309_0, i_13_471_3310_0, i_13_471_3423_0, i_13_471_3445_0,
    i_13_471_3525_0, i_13_471_3543_0, i_13_471_3552_0, i_13_471_3597_0,
    i_13_471_3616_0, i_13_471_3706_0, i_13_471_3731_0, i_13_471_3732_0,
    i_13_471_3786_0, i_13_471_3805_0, i_13_471_3831_0, i_13_471_3849_0,
    i_13_471_3858_0, i_13_471_3859_0, i_13_471_3912_0, i_13_471_3913_0,
    i_13_471_3994_0, i_13_471_4011_0, i_13_471_4012_0, i_13_471_4117_0,
    i_13_471_4161_0, i_13_471_4254_0, i_13_471_4369_0, i_13_471_4380_0,
    i_13_471_4381_0, i_13_471_4443_0, i_13_471_4587_0, i_13_471_4588_0;
  output o_13_471_0_0;
  assign o_13_471_0_0 = ~((~i_13_471_3912_0 & (~i_13_471_1501_0 | ~i_13_471_1555_0)) | (~i_13_471_483_0 & i_13_471_2005_0 & ~i_13_471_2299_0) | (~i_13_471_529_0 & ~i_13_471_3552_0) | (~i_13_471_1258_0 & ~i_13_471_3786_0) | (~i_13_471_2203_0 & ~i_13_471_2535_0 & ~i_13_471_3174_0 & ~i_13_471_4012_0) | (~i_13_471_1795_0 & i_13_471_1834_0 & ~i_13_471_4380_0) | (i_13_471_1556_0 & ~i_13_471_4381_0));
endmodule



// Benchmark "kernel_13_472" written by ABC on Sun Jul 19 10:51:56 2020

module kernel_13_472 ( 
    i_13_472_37_0, i_13_472_135_0, i_13_472_136_0, i_13_472_140_0,
    i_13_472_225_0, i_13_472_279_0, i_13_472_280_0, i_13_472_563_0,
    i_13_472_594_0, i_13_472_640_0, i_13_472_643_0, i_13_472_670_0,
    i_13_472_685_0, i_13_472_714_0, i_13_472_812_0, i_13_472_891_0,
    i_13_472_892_0, i_13_472_1025_0, i_13_472_1075_0, i_13_472_1093_0,
    i_13_472_1117_0, i_13_472_1200_0, i_13_472_1213_0, i_13_472_1214_0,
    i_13_472_1273_0, i_13_472_1314_0, i_13_472_1384_0, i_13_472_1387_0,
    i_13_472_1469_0, i_13_472_1480_0, i_13_472_1481_0, i_13_472_1669_0,
    i_13_472_1710_0, i_13_472_1711_0, i_13_472_1757_0, i_13_472_1778_0,
    i_13_472_1793_0, i_13_472_1828_0, i_13_472_1855_0, i_13_472_1881_0,
    i_13_472_1882_0, i_13_472_1885_0, i_13_472_1886_0, i_13_472_1915_0,
    i_13_472_2050_0, i_13_472_2380_0, i_13_472_2443_0, i_13_472_2585_0,
    i_13_472_2629_0, i_13_472_2630_0, i_13_472_2647_0, i_13_472_2649_0,
    i_13_472_2650_0, i_13_472_2651_0, i_13_472_2653_0, i_13_472_2656_0,
    i_13_472_2752_0, i_13_472_2844_0, i_13_472_2845_0, i_13_472_2849_0,
    i_13_472_2872_0, i_13_472_2874_0, i_13_472_2983_0, i_13_472_3109_0,
    i_13_472_3123_0, i_13_472_3208_0, i_13_472_3287_0, i_13_472_3311_0,
    i_13_472_3407_0, i_13_472_3429_0, i_13_472_3430_0, i_13_472_3448_0,
    i_13_472_3598_0, i_13_472_3757_0, i_13_472_3761_0, i_13_472_3781_0,
    i_13_472_3790_0, i_13_472_3791_0, i_13_472_3793_0, i_13_472_3835_0,
    i_13_472_3836_0, i_13_472_3871_0, i_13_472_3901_0, i_13_472_3923_0,
    i_13_472_3933_0, i_13_472_4042_0, i_13_472_4043_0, i_13_472_4054_0,
    i_13_472_4055_0, i_13_472_4096_0, i_13_472_4114_0, i_13_472_4198_0,
    i_13_472_4237_0, i_13_472_4351_0, i_13_472_4369_0, i_13_472_4388_0,
    i_13_472_4396_0, i_13_472_4441_0, i_13_472_4519_0, i_13_472_4567_0,
    o_13_472_0_0  );
  input  i_13_472_37_0, i_13_472_135_0, i_13_472_136_0, i_13_472_140_0,
    i_13_472_225_0, i_13_472_279_0, i_13_472_280_0, i_13_472_563_0,
    i_13_472_594_0, i_13_472_640_0, i_13_472_643_0, i_13_472_670_0,
    i_13_472_685_0, i_13_472_714_0, i_13_472_812_0, i_13_472_891_0,
    i_13_472_892_0, i_13_472_1025_0, i_13_472_1075_0, i_13_472_1093_0,
    i_13_472_1117_0, i_13_472_1200_0, i_13_472_1213_0, i_13_472_1214_0,
    i_13_472_1273_0, i_13_472_1314_0, i_13_472_1384_0, i_13_472_1387_0,
    i_13_472_1469_0, i_13_472_1480_0, i_13_472_1481_0, i_13_472_1669_0,
    i_13_472_1710_0, i_13_472_1711_0, i_13_472_1757_0, i_13_472_1778_0,
    i_13_472_1793_0, i_13_472_1828_0, i_13_472_1855_0, i_13_472_1881_0,
    i_13_472_1882_0, i_13_472_1885_0, i_13_472_1886_0, i_13_472_1915_0,
    i_13_472_2050_0, i_13_472_2380_0, i_13_472_2443_0, i_13_472_2585_0,
    i_13_472_2629_0, i_13_472_2630_0, i_13_472_2647_0, i_13_472_2649_0,
    i_13_472_2650_0, i_13_472_2651_0, i_13_472_2653_0, i_13_472_2656_0,
    i_13_472_2752_0, i_13_472_2844_0, i_13_472_2845_0, i_13_472_2849_0,
    i_13_472_2872_0, i_13_472_2874_0, i_13_472_2983_0, i_13_472_3109_0,
    i_13_472_3123_0, i_13_472_3208_0, i_13_472_3287_0, i_13_472_3311_0,
    i_13_472_3407_0, i_13_472_3429_0, i_13_472_3430_0, i_13_472_3448_0,
    i_13_472_3598_0, i_13_472_3757_0, i_13_472_3761_0, i_13_472_3781_0,
    i_13_472_3790_0, i_13_472_3791_0, i_13_472_3793_0, i_13_472_3835_0,
    i_13_472_3836_0, i_13_472_3871_0, i_13_472_3901_0, i_13_472_3923_0,
    i_13_472_3933_0, i_13_472_4042_0, i_13_472_4043_0, i_13_472_4054_0,
    i_13_472_4055_0, i_13_472_4096_0, i_13_472_4114_0, i_13_472_4198_0,
    i_13_472_4237_0, i_13_472_4351_0, i_13_472_4369_0, i_13_472_4388_0,
    i_13_472_4396_0, i_13_472_4441_0, i_13_472_4519_0, i_13_472_4567_0;
  output o_13_472_0_0;
  assign o_13_472_0_0 = ~(i_13_472_4369_0 | (~i_13_472_1710_0 & ~i_13_472_1711_0 & ~i_13_472_3781_0) | (~i_13_472_892_0 & ~i_13_472_1881_0 & ~i_13_472_2845_0));
endmodule



// Benchmark "kernel_13_473" written by ABC on Sun Jul 19 10:51:56 2020

module kernel_13_473 ( 
    i_13_473_48_0, i_13_473_51_0, i_13_473_52_0, i_13_473_72_0,
    i_13_473_73_0, i_13_473_166_0, i_13_473_169_0, i_13_473_285_0,
    i_13_473_339_0, i_13_473_384_0, i_13_473_618_0, i_13_473_619_0,
    i_13_473_678_0, i_13_473_690_0, i_13_473_771_0, i_13_473_816_0,
    i_13_473_817_0, i_13_473_840_0, i_13_473_844_0, i_13_473_856_0,
    i_13_473_1021_0, i_13_473_1069_0, i_13_473_1074_0, i_13_473_1258_0,
    i_13_473_1300_0, i_13_473_1390_0, i_13_473_1411_0, i_13_473_1572_0,
    i_13_473_1573_0, i_13_473_1623_0, i_13_473_1627_0, i_13_473_1629_0,
    i_13_473_1635_0, i_13_473_1636_0, i_13_473_1806_0, i_13_473_1807_0,
    i_13_473_1950_0, i_13_473_2014_0, i_13_473_2058_0, i_13_473_2059_0,
    i_13_473_2266_0, i_13_473_2283_0, i_13_473_2284_0, i_13_473_2346_0,
    i_13_473_2353_0, i_13_473_2380_0, i_13_473_2399_0, i_13_473_2410_0,
    i_13_473_2472_0, i_13_473_2536_0, i_13_473_2538_0, i_13_473_2590_0,
    i_13_473_2617_0, i_13_473_2650_0, i_13_473_2715_0, i_13_473_2751_0,
    i_13_473_2752_0, i_13_473_2759_0, i_13_473_2762_0, i_13_473_2787_0,
    i_13_473_2903_0, i_13_473_2941_0, i_13_473_3031_0, i_13_473_3042_0,
    i_13_473_3043_0, i_13_473_3109_0, i_13_473_3136_0, i_13_473_3141_0,
    i_13_473_3144_0, i_13_473_3147_0, i_13_473_3220_0, i_13_473_3292_0,
    i_13_473_3372_0, i_13_473_3373_0, i_13_473_3399_0, i_13_473_3526_0,
    i_13_473_3721_0, i_13_473_3730_0, i_13_473_3732_0, i_13_473_3850_0,
    i_13_473_3891_0, i_13_473_3915_0, i_13_473_4018_0, i_13_473_4020_0,
    i_13_473_4021_0, i_13_473_4047_0, i_13_473_4048_0, i_13_473_4131_0,
    i_13_473_4132_0, i_13_473_4234_0, i_13_473_4252_0, i_13_473_4255_0,
    i_13_473_4263_0, i_13_473_4300_0, i_13_473_4308_0, i_13_473_4318_0,
    i_13_473_4339_0, i_13_473_4554_0, i_13_473_4560_0, i_13_473_4561_0,
    o_13_473_0_0  );
  input  i_13_473_48_0, i_13_473_51_0, i_13_473_52_0, i_13_473_72_0,
    i_13_473_73_0, i_13_473_166_0, i_13_473_169_0, i_13_473_285_0,
    i_13_473_339_0, i_13_473_384_0, i_13_473_618_0, i_13_473_619_0,
    i_13_473_678_0, i_13_473_690_0, i_13_473_771_0, i_13_473_816_0,
    i_13_473_817_0, i_13_473_840_0, i_13_473_844_0, i_13_473_856_0,
    i_13_473_1021_0, i_13_473_1069_0, i_13_473_1074_0, i_13_473_1258_0,
    i_13_473_1300_0, i_13_473_1390_0, i_13_473_1411_0, i_13_473_1572_0,
    i_13_473_1573_0, i_13_473_1623_0, i_13_473_1627_0, i_13_473_1629_0,
    i_13_473_1635_0, i_13_473_1636_0, i_13_473_1806_0, i_13_473_1807_0,
    i_13_473_1950_0, i_13_473_2014_0, i_13_473_2058_0, i_13_473_2059_0,
    i_13_473_2266_0, i_13_473_2283_0, i_13_473_2284_0, i_13_473_2346_0,
    i_13_473_2353_0, i_13_473_2380_0, i_13_473_2399_0, i_13_473_2410_0,
    i_13_473_2472_0, i_13_473_2536_0, i_13_473_2538_0, i_13_473_2590_0,
    i_13_473_2617_0, i_13_473_2650_0, i_13_473_2715_0, i_13_473_2751_0,
    i_13_473_2752_0, i_13_473_2759_0, i_13_473_2762_0, i_13_473_2787_0,
    i_13_473_2903_0, i_13_473_2941_0, i_13_473_3031_0, i_13_473_3042_0,
    i_13_473_3043_0, i_13_473_3109_0, i_13_473_3136_0, i_13_473_3141_0,
    i_13_473_3144_0, i_13_473_3147_0, i_13_473_3220_0, i_13_473_3292_0,
    i_13_473_3372_0, i_13_473_3373_0, i_13_473_3399_0, i_13_473_3526_0,
    i_13_473_3721_0, i_13_473_3730_0, i_13_473_3732_0, i_13_473_3850_0,
    i_13_473_3891_0, i_13_473_3915_0, i_13_473_4018_0, i_13_473_4020_0,
    i_13_473_4021_0, i_13_473_4047_0, i_13_473_4048_0, i_13_473_4131_0,
    i_13_473_4132_0, i_13_473_4234_0, i_13_473_4252_0, i_13_473_4255_0,
    i_13_473_4263_0, i_13_473_4300_0, i_13_473_4308_0, i_13_473_4318_0,
    i_13_473_4339_0, i_13_473_4554_0, i_13_473_4560_0, i_13_473_4561_0;
  output o_13_473_0_0;
  assign o_13_473_0_0 = ~((~i_13_473_3147_0 & ((~i_13_473_816_0 & ~i_13_473_1573_0 & ~i_13_473_4255_0) | (~i_13_473_4048_0 & ~i_13_473_4560_0))) | (~i_13_473_52_0 & ~i_13_473_384_0 & ~i_13_473_817_0 & ~i_13_473_2283_0 & ~i_13_473_4047_0) | (i_13_473_1627_0 & ~i_13_473_4308_0) | (~i_13_473_1069_0 & ~i_13_473_3144_0 & ~i_13_473_4263_0 & ~i_13_473_4561_0));
endmodule



// Benchmark "kernel_13_474" written by ABC on Sun Jul 19 10:51:57 2020

module kernel_13_474 ( 
    i_13_474_95_0, i_13_474_98_0, i_13_474_134_0, i_13_474_139_0,
    i_13_474_170_0, i_13_474_175_0, i_13_474_176_0, i_13_474_178_0,
    i_13_474_233_0, i_13_474_311_0, i_13_474_374_0, i_13_474_428_0,
    i_13_474_464_0, i_13_474_527_0, i_13_474_575_0, i_13_474_599_0,
    i_13_474_646_0, i_13_474_664_0, i_13_474_671_0, i_13_474_818_0,
    i_13_474_851_0, i_13_474_854_0, i_13_474_985_0, i_13_474_986_0,
    i_13_474_989_0, i_13_474_1024_0, i_13_474_1070_0, i_13_474_1232_0,
    i_13_474_1300_0, i_13_474_1309_0, i_13_474_1327_0, i_13_474_1408_0,
    i_13_474_1436_0, i_13_474_1571_0, i_13_474_1723_0, i_13_474_1754_0,
    i_13_474_1765_0, i_13_474_1805_0, i_13_474_1831_0, i_13_474_1832_0,
    i_13_474_1850_0, i_13_474_1852_0, i_13_474_1853_0, i_13_474_1862_0,
    i_13_474_1885_0, i_13_474_1921_0, i_13_474_2300_0, i_13_474_2308_0,
    i_13_474_2366_0, i_13_474_2408_0, i_13_474_2461_0, i_13_474_2471_0,
    i_13_474_2473_0, i_13_474_2510_0, i_13_474_2633_0, i_13_474_2662_0,
    i_13_474_2680_0, i_13_474_2698_0, i_13_474_2848_0, i_13_474_2983_0,
    i_13_474_2987_0, i_13_474_3001_0, i_13_474_3013_0, i_13_474_3106_0,
    i_13_474_3109_0, i_13_474_3110_0, i_13_474_3112_0, i_13_474_3113_0,
    i_13_474_3116_0, i_13_474_3137_0, i_13_474_3157_0, i_13_474_3272_0,
    i_13_474_3404_0, i_13_474_3410_0, i_13_474_3419_0, i_13_474_3425_0,
    i_13_474_3427_0, i_13_474_3481_0, i_13_474_3490_0, i_13_474_3637_0,
    i_13_474_3686_0, i_13_474_3769_0, i_13_474_3799_0, i_13_474_3800_0,
    i_13_474_3820_0, i_13_474_3821_0, i_13_474_3860_0, i_13_474_3977_0,
    i_13_474_4022_0, i_13_474_4064_0, i_13_474_4067_0, i_13_474_4127_0,
    i_13_474_4354_0, i_13_474_4378_0, i_13_474_4444_0, i_13_474_4460_0,
    i_13_474_4513_0, i_13_474_4567_0, i_13_474_4568_0, i_13_474_4570_0,
    o_13_474_0_0  );
  input  i_13_474_95_0, i_13_474_98_0, i_13_474_134_0, i_13_474_139_0,
    i_13_474_170_0, i_13_474_175_0, i_13_474_176_0, i_13_474_178_0,
    i_13_474_233_0, i_13_474_311_0, i_13_474_374_0, i_13_474_428_0,
    i_13_474_464_0, i_13_474_527_0, i_13_474_575_0, i_13_474_599_0,
    i_13_474_646_0, i_13_474_664_0, i_13_474_671_0, i_13_474_818_0,
    i_13_474_851_0, i_13_474_854_0, i_13_474_985_0, i_13_474_986_0,
    i_13_474_989_0, i_13_474_1024_0, i_13_474_1070_0, i_13_474_1232_0,
    i_13_474_1300_0, i_13_474_1309_0, i_13_474_1327_0, i_13_474_1408_0,
    i_13_474_1436_0, i_13_474_1571_0, i_13_474_1723_0, i_13_474_1754_0,
    i_13_474_1765_0, i_13_474_1805_0, i_13_474_1831_0, i_13_474_1832_0,
    i_13_474_1850_0, i_13_474_1852_0, i_13_474_1853_0, i_13_474_1862_0,
    i_13_474_1885_0, i_13_474_1921_0, i_13_474_2300_0, i_13_474_2308_0,
    i_13_474_2366_0, i_13_474_2408_0, i_13_474_2461_0, i_13_474_2471_0,
    i_13_474_2473_0, i_13_474_2510_0, i_13_474_2633_0, i_13_474_2662_0,
    i_13_474_2680_0, i_13_474_2698_0, i_13_474_2848_0, i_13_474_2983_0,
    i_13_474_2987_0, i_13_474_3001_0, i_13_474_3013_0, i_13_474_3106_0,
    i_13_474_3109_0, i_13_474_3110_0, i_13_474_3112_0, i_13_474_3113_0,
    i_13_474_3116_0, i_13_474_3137_0, i_13_474_3157_0, i_13_474_3272_0,
    i_13_474_3404_0, i_13_474_3410_0, i_13_474_3419_0, i_13_474_3425_0,
    i_13_474_3427_0, i_13_474_3481_0, i_13_474_3490_0, i_13_474_3637_0,
    i_13_474_3686_0, i_13_474_3769_0, i_13_474_3799_0, i_13_474_3800_0,
    i_13_474_3820_0, i_13_474_3821_0, i_13_474_3860_0, i_13_474_3977_0,
    i_13_474_4022_0, i_13_474_4064_0, i_13_474_4067_0, i_13_474_4127_0,
    i_13_474_4354_0, i_13_474_4378_0, i_13_474_4444_0, i_13_474_4460_0,
    i_13_474_4513_0, i_13_474_4567_0, i_13_474_4568_0, i_13_474_4570_0;
  output o_13_474_0_0;
  assign o_13_474_0_0 = ~((~i_13_474_986_0 & ((~i_13_474_178_0 & ~i_13_474_3013_0) | (~i_13_474_1832_0 & ~i_13_474_2300_0 & ~i_13_474_4570_0))) | (~i_13_474_1832_0 & ((~i_13_474_1232_0 & ~i_13_474_2680_0 & ~i_13_474_3427_0) | (~i_13_474_1408_0 & ~i_13_474_1754_0 & ~i_13_474_4067_0 & ~i_13_474_4354_0))) | (~i_13_474_3112_0 & ((~i_13_474_2408_0 & ~i_13_474_3110_0 & ~i_13_474_3490_0 & ~i_13_474_3821_0) | (~i_13_474_4513_0 & ~i_13_474_4568_0))) | (~i_13_474_464_0 & i_13_474_1885_0 & ~i_13_474_3109_0 & ~i_13_474_3425_0 & ~i_13_474_4513_0) | (~i_13_474_311_0 & i_13_474_2461_0 & ~i_13_474_3427_0 & ~i_13_474_3860_0 & ~i_13_474_4354_0));
endmodule



// Benchmark "kernel_13_475" written by ABC on Sun Jul 19 10:51:58 2020

module kernel_13_475 ( 
    i_13_475_273_0, i_13_475_283_0, i_13_475_354_0, i_13_475_355_0,
    i_13_475_364_0, i_13_475_469_0, i_13_475_490_0, i_13_475_598_0,
    i_13_475_640_0, i_13_475_651_0, i_13_475_658_0, i_13_475_660_0,
    i_13_475_765_0, i_13_475_767_0, i_13_475_927_0, i_13_475_928_0,
    i_13_475_939_0, i_13_475_940_0, i_13_475_948_0, i_13_475_1037_0,
    i_13_475_1071_0, i_13_475_1080_0, i_13_475_1081_0, i_13_475_1082_0,
    i_13_475_1098_0, i_13_475_1099_0, i_13_475_1116_0, i_13_475_1225_0,
    i_13_475_1227_0, i_13_475_1306_0, i_13_475_1307_0, i_13_475_1443_0,
    i_13_475_1486_0, i_13_475_1497_0, i_13_475_1498_0, i_13_475_1566_0,
    i_13_475_1567_0, i_13_475_1620_0, i_13_475_1639_0, i_13_475_1710_0,
    i_13_475_1719_0, i_13_475_1720_0, i_13_475_1729_0, i_13_475_1765_0,
    i_13_475_1774_0, i_13_475_1782_0, i_13_475_1837_0, i_13_475_1840_0,
    i_13_475_1846_0, i_13_475_1927_0, i_13_475_1971_0, i_13_475_2100_0,
    i_13_475_2205_0, i_13_475_2259_0, i_13_475_2324_0, i_13_475_2358_0,
    i_13_475_2424_0, i_13_475_2467_0, i_13_475_2485_0, i_13_475_2587_0,
    i_13_475_2673_0, i_13_475_2684_0, i_13_475_2781_0, i_13_475_2844_0,
    i_13_475_2845_0, i_13_475_2884_0, i_13_475_3025_0, i_13_475_3163_0,
    i_13_475_3258_0, i_13_475_3285_0, i_13_475_3286_0, i_13_475_3361_0,
    i_13_475_3388_0, i_13_475_3420_0, i_13_475_3423_0, i_13_475_3424_0,
    i_13_475_3457_0, i_13_475_3487_0, i_13_475_3600_0, i_13_475_3601_0,
    i_13_475_3619_0, i_13_475_3754_0, i_13_475_3924_0, i_13_475_3933_0,
    i_13_475_3988_0, i_13_475_4008_0, i_13_475_4009_0, i_13_475_4050_0,
    i_13_475_4051_0, i_13_475_4077_0, i_13_475_4086_0, i_13_475_4088_0,
    i_13_475_4104_0, i_13_475_4195_0, i_13_475_4312_0, i_13_475_4377_0,
    i_13_475_4428_0, i_13_475_4429_0, i_13_475_4540_0, i_13_475_4582_0,
    o_13_475_0_0  );
  input  i_13_475_273_0, i_13_475_283_0, i_13_475_354_0, i_13_475_355_0,
    i_13_475_364_0, i_13_475_469_0, i_13_475_490_0, i_13_475_598_0,
    i_13_475_640_0, i_13_475_651_0, i_13_475_658_0, i_13_475_660_0,
    i_13_475_765_0, i_13_475_767_0, i_13_475_927_0, i_13_475_928_0,
    i_13_475_939_0, i_13_475_940_0, i_13_475_948_0, i_13_475_1037_0,
    i_13_475_1071_0, i_13_475_1080_0, i_13_475_1081_0, i_13_475_1082_0,
    i_13_475_1098_0, i_13_475_1099_0, i_13_475_1116_0, i_13_475_1225_0,
    i_13_475_1227_0, i_13_475_1306_0, i_13_475_1307_0, i_13_475_1443_0,
    i_13_475_1486_0, i_13_475_1497_0, i_13_475_1498_0, i_13_475_1566_0,
    i_13_475_1567_0, i_13_475_1620_0, i_13_475_1639_0, i_13_475_1710_0,
    i_13_475_1719_0, i_13_475_1720_0, i_13_475_1729_0, i_13_475_1765_0,
    i_13_475_1774_0, i_13_475_1782_0, i_13_475_1837_0, i_13_475_1840_0,
    i_13_475_1846_0, i_13_475_1927_0, i_13_475_1971_0, i_13_475_2100_0,
    i_13_475_2205_0, i_13_475_2259_0, i_13_475_2324_0, i_13_475_2358_0,
    i_13_475_2424_0, i_13_475_2467_0, i_13_475_2485_0, i_13_475_2587_0,
    i_13_475_2673_0, i_13_475_2684_0, i_13_475_2781_0, i_13_475_2844_0,
    i_13_475_2845_0, i_13_475_2884_0, i_13_475_3025_0, i_13_475_3163_0,
    i_13_475_3258_0, i_13_475_3285_0, i_13_475_3286_0, i_13_475_3361_0,
    i_13_475_3388_0, i_13_475_3420_0, i_13_475_3423_0, i_13_475_3424_0,
    i_13_475_3457_0, i_13_475_3487_0, i_13_475_3600_0, i_13_475_3601_0,
    i_13_475_3619_0, i_13_475_3754_0, i_13_475_3924_0, i_13_475_3933_0,
    i_13_475_3988_0, i_13_475_4008_0, i_13_475_4009_0, i_13_475_4050_0,
    i_13_475_4051_0, i_13_475_4077_0, i_13_475_4086_0, i_13_475_4088_0,
    i_13_475_4104_0, i_13_475_4195_0, i_13_475_4312_0, i_13_475_4377_0,
    i_13_475_4428_0, i_13_475_4429_0, i_13_475_4540_0, i_13_475_4582_0;
  output o_13_475_0_0;
  assign o_13_475_0_0 = ~(~i_13_475_928_0 | (~i_13_475_2673_0 & ~i_13_475_2844_0));
endmodule



// Benchmark "kernel_13_476" written by ABC on Sun Jul 19 10:51:59 2020

module kernel_13_476 ( 
    i_13_476_182_0, i_13_476_193_0, i_13_476_319_0, i_13_476_325_0,
    i_13_476_328_0, i_13_476_349_0, i_13_476_415_0, i_13_476_416_0,
    i_13_476_424_0, i_13_476_658_0, i_13_476_715_0, i_13_476_716_0,
    i_13_476_813_0, i_13_476_814_0, i_13_476_826_0, i_13_476_848_0,
    i_13_476_859_0, i_13_476_860_0, i_13_476_863_0, i_13_476_895_0,
    i_13_476_1072_0, i_13_476_1219_0, i_13_476_1224_0, i_13_476_1225_0,
    i_13_476_1226_0, i_13_476_1228_0, i_13_476_1229_0, i_13_476_1252_0,
    i_13_476_1255_0, i_13_476_1259_0, i_13_476_1315_0, i_13_476_1316_0,
    i_13_476_1318_0, i_13_476_1319_0, i_13_476_1345_0, i_13_476_1391_0,
    i_13_476_1404_0, i_13_476_1405_0, i_13_476_1411_0, i_13_476_1432_0,
    i_13_476_1444_0, i_13_476_1451_0, i_13_476_1484_0, i_13_476_1486_0,
    i_13_476_1490_0, i_13_476_1492_0, i_13_476_1541_0, i_13_476_1549_0,
    i_13_476_1553_0, i_13_476_1597_0, i_13_476_1677_0, i_13_476_1714_0,
    i_13_476_1750_0, i_13_476_1774_0, i_13_476_1778_0, i_13_476_1855_0,
    i_13_476_1871_0, i_13_476_1904_0, i_13_476_1922_0, i_13_476_1954_0,
    i_13_476_1955_0, i_13_476_1957_0, i_13_476_2056_0, i_13_476_2059_0,
    i_13_476_2137_0, i_13_476_2268_0, i_13_476_2506_0, i_13_476_2543_0,
    i_13_476_2611_0, i_13_476_2613_0, i_13_476_2614_0, i_13_476_2618_0,
    i_13_476_2633_0, i_13_476_2659_0, i_13_476_2660_0, i_13_476_2698_0,
    i_13_476_2705_0, i_13_476_2979_0, i_13_476_3005_0, i_13_476_3114_0,
    i_13_476_3119_0, i_13_476_3175_0, i_13_476_3287_0, i_13_476_3352_0,
    i_13_476_3369_0, i_13_476_3370_0, i_13_476_3421_0, i_13_476_3485_0,
    i_13_476_3506_0, i_13_476_3538_0, i_13_476_3539_0, i_13_476_3574_0,
    i_13_476_3595_0, i_13_476_3853_0, i_13_476_3979_0, i_13_476_4036_0,
    i_13_476_4249_0, i_13_476_4369_0, i_13_476_4376_0, i_13_476_4589_0,
    o_13_476_0_0  );
  input  i_13_476_182_0, i_13_476_193_0, i_13_476_319_0, i_13_476_325_0,
    i_13_476_328_0, i_13_476_349_0, i_13_476_415_0, i_13_476_416_0,
    i_13_476_424_0, i_13_476_658_0, i_13_476_715_0, i_13_476_716_0,
    i_13_476_813_0, i_13_476_814_0, i_13_476_826_0, i_13_476_848_0,
    i_13_476_859_0, i_13_476_860_0, i_13_476_863_0, i_13_476_895_0,
    i_13_476_1072_0, i_13_476_1219_0, i_13_476_1224_0, i_13_476_1225_0,
    i_13_476_1226_0, i_13_476_1228_0, i_13_476_1229_0, i_13_476_1252_0,
    i_13_476_1255_0, i_13_476_1259_0, i_13_476_1315_0, i_13_476_1316_0,
    i_13_476_1318_0, i_13_476_1319_0, i_13_476_1345_0, i_13_476_1391_0,
    i_13_476_1404_0, i_13_476_1405_0, i_13_476_1411_0, i_13_476_1432_0,
    i_13_476_1444_0, i_13_476_1451_0, i_13_476_1484_0, i_13_476_1486_0,
    i_13_476_1490_0, i_13_476_1492_0, i_13_476_1541_0, i_13_476_1549_0,
    i_13_476_1553_0, i_13_476_1597_0, i_13_476_1677_0, i_13_476_1714_0,
    i_13_476_1750_0, i_13_476_1774_0, i_13_476_1778_0, i_13_476_1855_0,
    i_13_476_1871_0, i_13_476_1904_0, i_13_476_1922_0, i_13_476_1954_0,
    i_13_476_1955_0, i_13_476_1957_0, i_13_476_2056_0, i_13_476_2059_0,
    i_13_476_2137_0, i_13_476_2268_0, i_13_476_2506_0, i_13_476_2543_0,
    i_13_476_2611_0, i_13_476_2613_0, i_13_476_2614_0, i_13_476_2618_0,
    i_13_476_2633_0, i_13_476_2659_0, i_13_476_2660_0, i_13_476_2698_0,
    i_13_476_2705_0, i_13_476_2979_0, i_13_476_3005_0, i_13_476_3114_0,
    i_13_476_3119_0, i_13_476_3175_0, i_13_476_3287_0, i_13_476_3352_0,
    i_13_476_3369_0, i_13_476_3370_0, i_13_476_3421_0, i_13_476_3485_0,
    i_13_476_3506_0, i_13_476_3538_0, i_13_476_3539_0, i_13_476_3574_0,
    i_13_476_3595_0, i_13_476_3853_0, i_13_476_3979_0, i_13_476_4036_0,
    i_13_476_4249_0, i_13_476_4369_0, i_13_476_4376_0, i_13_476_4589_0;
  output o_13_476_0_0;
  assign o_13_476_0_0 = ~((~i_13_476_4376_0 & (i_13_476_1219_0 | (~i_13_476_1490_0 & ~i_13_476_4369_0))) | (~i_13_476_416_0 & i_13_476_859_0 & i_13_476_1597_0) | (~i_13_476_1316_0 & ~i_13_476_1486_0 & ~i_13_476_1714_0) | (~i_13_476_193_0 & ~i_13_476_1855_0) | (~i_13_476_1255_0 & ~i_13_476_1774_0 & ~i_13_476_3539_0) | (~i_13_476_1405_0 & ~i_13_476_1677_0 & ~i_13_476_1955_0 & ~i_13_476_3979_0));
endmodule



// Benchmark "kernel_13_477" written by ABC on Sun Jul 19 10:51:59 2020

module kernel_13_477 ( 
    i_13_477_35_0, i_13_477_40_0, i_13_477_48_0, i_13_477_63_0,
    i_13_477_71_0, i_13_477_121_0, i_13_477_135_0, i_13_477_230_0,
    i_13_477_241_0, i_13_477_306_0, i_13_477_310_0, i_13_477_316_0,
    i_13_477_319_0, i_13_477_414_0, i_13_477_550_0, i_13_477_557_0,
    i_13_477_588_0, i_13_477_598_0, i_13_477_604_0, i_13_477_609_0,
    i_13_477_612_0, i_13_477_613_0, i_13_477_671_0, i_13_477_679_0,
    i_13_477_680_0, i_13_477_685_0, i_13_477_688_0, i_13_477_764_0,
    i_13_477_819_0, i_13_477_953_0, i_13_477_1116_0, i_13_477_1132_0,
    i_13_477_1207_0, i_13_477_1224_0, i_13_477_1269_0, i_13_477_1308_0,
    i_13_477_1422_0, i_13_477_1440_0, i_13_477_1441_0, i_13_477_1507_0,
    i_13_477_1526_0, i_13_477_1548_0, i_13_477_1596_0, i_13_477_1609_0,
    i_13_477_1673_0, i_13_477_1699_0, i_13_477_1700_0, i_13_477_1729_0,
    i_13_477_1764_0, i_13_477_1799_0, i_13_477_1847_0, i_13_477_1926_0,
    i_13_477_1927_0, i_13_477_1930_0, i_13_477_1944_0, i_13_477_2426_0,
    i_13_477_2461_0, i_13_477_2550_0, i_13_477_2557_0, i_13_477_2584_0,
    i_13_477_2673_0, i_13_477_2676_0, i_13_477_2718_0, i_13_477_2749_0,
    i_13_477_2771_0, i_13_477_3000_0, i_13_477_3217_0, i_13_477_3245_0,
    i_13_477_3267_0, i_13_477_3367_0, i_13_477_3483_0, i_13_477_3558_0,
    i_13_477_3637_0, i_13_477_3641_0, i_13_477_3653_0, i_13_477_3743_0,
    i_13_477_3754_0, i_13_477_3816_0, i_13_477_3871_0, i_13_477_3924_0,
    i_13_477_3937_0, i_13_477_3986_0, i_13_477_4032_0, i_13_477_4033_0,
    i_13_477_4035_0, i_13_477_4039_0, i_13_477_4217_0, i_13_477_4248_0,
    i_13_477_4250_0, i_13_477_4251_0, i_13_477_4293_0, i_13_477_4294_0,
    i_13_477_4298_0, i_13_477_4367_0, i_13_477_4521_0, i_13_477_4522_0,
    i_13_477_4565_0, i_13_477_4591_0, i_13_477_4593_0, i_13_477_4594_0,
    o_13_477_0_0  );
  input  i_13_477_35_0, i_13_477_40_0, i_13_477_48_0, i_13_477_63_0,
    i_13_477_71_0, i_13_477_121_0, i_13_477_135_0, i_13_477_230_0,
    i_13_477_241_0, i_13_477_306_0, i_13_477_310_0, i_13_477_316_0,
    i_13_477_319_0, i_13_477_414_0, i_13_477_550_0, i_13_477_557_0,
    i_13_477_588_0, i_13_477_598_0, i_13_477_604_0, i_13_477_609_0,
    i_13_477_612_0, i_13_477_613_0, i_13_477_671_0, i_13_477_679_0,
    i_13_477_680_0, i_13_477_685_0, i_13_477_688_0, i_13_477_764_0,
    i_13_477_819_0, i_13_477_953_0, i_13_477_1116_0, i_13_477_1132_0,
    i_13_477_1207_0, i_13_477_1224_0, i_13_477_1269_0, i_13_477_1308_0,
    i_13_477_1422_0, i_13_477_1440_0, i_13_477_1441_0, i_13_477_1507_0,
    i_13_477_1526_0, i_13_477_1548_0, i_13_477_1596_0, i_13_477_1609_0,
    i_13_477_1673_0, i_13_477_1699_0, i_13_477_1700_0, i_13_477_1729_0,
    i_13_477_1764_0, i_13_477_1799_0, i_13_477_1847_0, i_13_477_1926_0,
    i_13_477_1927_0, i_13_477_1930_0, i_13_477_1944_0, i_13_477_2426_0,
    i_13_477_2461_0, i_13_477_2550_0, i_13_477_2557_0, i_13_477_2584_0,
    i_13_477_2673_0, i_13_477_2676_0, i_13_477_2718_0, i_13_477_2749_0,
    i_13_477_2771_0, i_13_477_3000_0, i_13_477_3217_0, i_13_477_3245_0,
    i_13_477_3267_0, i_13_477_3367_0, i_13_477_3483_0, i_13_477_3558_0,
    i_13_477_3637_0, i_13_477_3641_0, i_13_477_3653_0, i_13_477_3743_0,
    i_13_477_3754_0, i_13_477_3816_0, i_13_477_3871_0, i_13_477_3924_0,
    i_13_477_3937_0, i_13_477_3986_0, i_13_477_4032_0, i_13_477_4033_0,
    i_13_477_4035_0, i_13_477_4039_0, i_13_477_4217_0, i_13_477_4248_0,
    i_13_477_4250_0, i_13_477_4251_0, i_13_477_4293_0, i_13_477_4294_0,
    i_13_477_4298_0, i_13_477_4367_0, i_13_477_4521_0, i_13_477_4522_0,
    i_13_477_4565_0, i_13_477_4591_0, i_13_477_4593_0, i_13_477_4594_0;
  output o_13_477_0_0;
  assign o_13_477_0_0 = ~((~i_13_477_1422_0 & (~i_13_477_1116_0 | (~i_13_477_1729_0 & i_13_477_3754_0))) | ~i_13_477_319_0 | ~i_13_477_1207_0 | (~i_13_477_685_0 & i_13_477_1422_0 & i_13_477_4251_0));
endmodule



// Benchmark "kernel_13_478" written by ABC on Sun Jul 19 10:52:00 2020

module kernel_13_478 ( 
    i_13_478_61_0, i_13_478_168_0, i_13_478_170_0, i_13_478_195_0,
    i_13_478_327_0, i_13_478_391_0, i_13_478_422_0, i_13_478_528_0,
    i_13_478_535_0, i_13_478_572_0, i_13_478_598_0, i_13_478_664_0,
    i_13_478_734_0, i_13_478_798_0, i_13_478_799_0, i_13_478_800_0,
    i_13_478_812_0, i_13_478_826_0, i_13_478_853_0, i_13_478_861_0,
    i_13_478_862_0, i_13_478_909_0, i_13_478_951_0, i_13_478_958_0,
    i_13_478_1069_0, i_13_478_1087_0, i_13_478_1119_0, i_13_478_1219_0,
    i_13_478_1226_0, i_13_478_1227_0, i_13_478_1228_0, i_13_478_1230_0,
    i_13_478_1231_0, i_13_478_1257_0, i_13_478_1258_0, i_13_478_1285_0,
    i_13_478_1300_0, i_13_478_1301_0, i_13_478_1302_0, i_13_478_1410_0,
    i_13_478_1437_0, i_13_478_1446_0, i_13_478_1482_0, i_13_478_1491_0,
    i_13_478_1492_0, i_13_478_1496_0, i_13_478_1523_0, i_13_478_1552_0,
    i_13_478_1554_0, i_13_478_1555_0, i_13_478_1755_0, i_13_478_1804_0,
    i_13_478_1829_0, i_13_478_1860_0, i_13_478_1959_0, i_13_478_1960_0,
    i_13_478_2008_0, i_13_478_2014_0, i_13_478_2103_0, i_13_478_2225_0,
    i_13_478_2239_0, i_13_478_2317_0, i_13_478_2347_0, i_13_478_2491_0,
    i_13_478_2535_0, i_13_478_2571_0, i_13_478_2707_0, i_13_478_2857_0,
    i_13_478_2972_0, i_13_478_2976_0, i_13_478_3121_0, i_13_478_3136_0,
    i_13_478_3145_0, i_13_478_3219_0, i_13_478_3233_0, i_13_478_3310_0,
    i_13_478_3410_0, i_13_478_3422_0, i_13_478_3423_0, i_13_478_3487_0,
    i_13_478_3489_0, i_13_478_3490_0, i_13_478_3531_0, i_13_478_3543_0,
    i_13_478_3639_0, i_13_478_3688_0, i_13_478_3739_0, i_13_478_3805_0,
    i_13_478_3858_0, i_13_478_3859_0, i_13_478_3984_0, i_13_478_3985_0,
    i_13_478_4380_0, i_13_478_4381_0, i_13_478_4396_0, i_13_478_4416_0,
    i_13_478_4454_0, i_13_478_4512_0, i_13_478_4528_0, i_13_478_4587_0,
    o_13_478_0_0  );
  input  i_13_478_61_0, i_13_478_168_0, i_13_478_170_0, i_13_478_195_0,
    i_13_478_327_0, i_13_478_391_0, i_13_478_422_0, i_13_478_528_0,
    i_13_478_535_0, i_13_478_572_0, i_13_478_598_0, i_13_478_664_0,
    i_13_478_734_0, i_13_478_798_0, i_13_478_799_0, i_13_478_800_0,
    i_13_478_812_0, i_13_478_826_0, i_13_478_853_0, i_13_478_861_0,
    i_13_478_862_0, i_13_478_909_0, i_13_478_951_0, i_13_478_958_0,
    i_13_478_1069_0, i_13_478_1087_0, i_13_478_1119_0, i_13_478_1219_0,
    i_13_478_1226_0, i_13_478_1227_0, i_13_478_1228_0, i_13_478_1230_0,
    i_13_478_1231_0, i_13_478_1257_0, i_13_478_1258_0, i_13_478_1285_0,
    i_13_478_1300_0, i_13_478_1301_0, i_13_478_1302_0, i_13_478_1410_0,
    i_13_478_1437_0, i_13_478_1446_0, i_13_478_1482_0, i_13_478_1491_0,
    i_13_478_1492_0, i_13_478_1496_0, i_13_478_1523_0, i_13_478_1552_0,
    i_13_478_1554_0, i_13_478_1555_0, i_13_478_1755_0, i_13_478_1804_0,
    i_13_478_1829_0, i_13_478_1860_0, i_13_478_1959_0, i_13_478_1960_0,
    i_13_478_2008_0, i_13_478_2014_0, i_13_478_2103_0, i_13_478_2225_0,
    i_13_478_2239_0, i_13_478_2317_0, i_13_478_2347_0, i_13_478_2491_0,
    i_13_478_2535_0, i_13_478_2571_0, i_13_478_2707_0, i_13_478_2857_0,
    i_13_478_2972_0, i_13_478_2976_0, i_13_478_3121_0, i_13_478_3136_0,
    i_13_478_3145_0, i_13_478_3219_0, i_13_478_3233_0, i_13_478_3310_0,
    i_13_478_3410_0, i_13_478_3422_0, i_13_478_3423_0, i_13_478_3487_0,
    i_13_478_3489_0, i_13_478_3490_0, i_13_478_3531_0, i_13_478_3543_0,
    i_13_478_3639_0, i_13_478_3688_0, i_13_478_3739_0, i_13_478_3805_0,
    i_13_478_3858_0, i_13_478_3859_0, i_13_478_3984_0, i_13_478_3985_0,
    i_13_478_4380_0, i_13_478_4381_0, i_13_478_4396_0, i_13_478_4416_0,
    i_13_478_4454_0, i_13_478_4512_0, i_13_478_4528_0, i_13_478_4587_0;
  output o_13_478_0_0;
  assign o_13_478_0_0 = ~((~i_13_478_3489_0 & ((~i_13_478_3219_0 & ~i_13_478_3487_0) | (~i_13_478_3145_0 & ~i_13_478_4454_0))) | (~i_13_478_3858_0 & (~i_13_478_1804_0 | (~i_13_478_1230_0 & ~i_13_478_1258_0))) | (i_13_478_422_0 & ~i_13_478_4381_0));
endmodule



// Benchmark "kernel_13_479" written by ABC on Sun Jul 19 10:52:01 2020

module kernel_13_479 ( 
    i_13_479_51_0, i_13_479_159_0, i_13_479_209_0, i_13_479_245_0,
    i_13_479_323_0, i_13_479_339_0, i_13_479_358_0, i_13_479_384_0,
    i_13_479_385_0, i_13_479_466_0, i_13_479_511_0, i_13_479_520_0,
    i_13_479_527_0, i_13_479_591_0, i_13_479_643_0, i_13_479_674_0,
    i_13_479_678_0, i_13_479_728_0, i_13_479_744_0, i_13_479_745_0,
    i_13_479_762_0, i_13_479_763_0, i_13_479_940_0, i_13_479_962_0,
    i_13_479_1066_0, i_13_479_1074_0, i_13_479_1130_0, i_13_479_1131_0,
    i_13_479_1213_0, i_13_479_1245_0, i_13_479_1301_0, i_13_479_1302_0,
    i_13_479_1303_0, i_13_479_1313_0, i_13_479_1346_0, i_13_479_1390_0,
    i_13_479_1403_0, i_13_479_1606_0, i_13_479_1632_0, i_13_479_1633_0,
    i_13_479_1634_0, i_13_479_1816_0, i_13_479_1835_0, i_13_479_1995_0,
    i_13_479_1996_0, i_13_479_2057_0, i_13_479_2058_0, i_13_479_2059_0,
    i_13_479_2121_0, i_13_479_2122_0, i_13_479_2204_0, i_13_479_2239_0,
    i_13_479_2265_0, i_13_479_2266_0, i_13_479_2267_0, i_13_479_2436_0,
    i_13_479_2460_0, i_13_479_2543_0, i_13_479_2617_0, i_13_479_2699_0,
    i_13_479_2847_0, i_13_479_2848_0, i_13_479_2859_0, i_13_479_2921_0,
    i_13_479_2941_0, i_13_479_3009_0, i_13_479_3011_0, i_13_479_3021_0,
    i_13_479_3022_0, i_13_479_3154_0, i_13_479_3273_0, i_13_479_3345_0,
    i_13_479_3346_0, i_13_479_3390_0, i_13_479_3399_0, i_13_479_3536_0,
    i_13_479_3542_0, i_13_479_3578_0, i_13_479_3619_0, i_13_479_3634_0,
    i_13_479_3669_0, i_13_479_3670_0, i_13_479_3692_0, i_13_479_3729_0,
    i_13_479_3731_0, i_13_479_3738_0, i_13_479_3739_0, i_13_479_3844_0,
    i_13_479_3846_0, i_13_479_3847_0, i_13_479_3892_0, i_13_479_3909_0,
    i_13_479_3911_0, i_13_479_4056_0, i_13_479_4217_0, i_13_479_4236_0,
    i_13_479_4255_0, i_13_479_4273_0, i_13_479_4399_0, i_13_479_4546_0,
    o_13_479_0_0  );
  input  i_13_479_51_0, i_13_479_159_0, i_13_479_209_0, i_13_479_245_0,
    i_13_479_323_0, i_13_479_339_0, i_13_479_358_0, i_13_479_384_0,
    i_13_479_385_0, i_13_479_466_0, i_13_479_511_0, i_13_479_520_0,
    i_13_479_527_0, i_13_479_591_0, i_13_479_643_0, i_13_479_674_0,
    i_13_479_678_0, i_13_479_728_0, i_13_479_744_0, i_13_479_745_0,
    i_13_479_762_0, i_13_479_763_0, i_13_479_940_0, i_13_479_962_0,
    i_13_479_1066_0, i_13_479_1074_0, i_13_479_1130_0, i_13_479_1131_0,
    i_13_479_1213_0, i_13_479_1245_0, i_13_479_1301_0, i_13_479_1302_0,
    i_13_479_1303_0, i_13_479_1313_0, i_13_479_1346_0, i_13_479_1390_0,
    i_13_479_1403_0, i_13_479_1606_0, i_13_479_1632_0, i_13_479_1633_0,
    i_13_479_1634_0, i_13_479_1816_0, i_13_479_1835_0, i_13_479_1995_0,
    i_13_479_1996_0, i_13_479_2057_0, i_13_479_2058_0, i_13_479_2059_0,
    i_13_479_2121_0, i_13_479_2122_0, i_13_479_2204_0, i_13_479_2239_0,
    i_13_479_2265_0, i_13_479_2266_0, i_13_479_2267_0, i_13_479_2436_0,
    i_13_479_2460_0, i_13_479_2543_0, i_13_479_2617_0, i_13_479_2699_0,
    i_13_479_2847_0, i_13_479_2848_0, i_13_479_2859_0, i_13_479_2921_0,
    i_13_479_2941_0, i_13_479_3009_0, i_13_479_3011_0, i_13_479_3021_0,
    i_13_479_3022_0, i_13_479_3154_0, i_13_479_3273_0, i_13_479_3345_0,
    i_13_479_3346_0, i_13_479_3390_0, i_13_479_3399_0, i_13_479_3536_0,
    i_13_479_3542_0, i_13_479_3578_0, i_13_479_3619_0, i_13_479_3634_0,
    i_13_479_3669_0, i_13_479_3670_0, i_13_479_3692_0, i_13_479_3729_0,
    i_13_479_3731_0, i_13_479_3738_0, i_13_479_3739_0, i_13_479_3844_0,
    i_13_479_3846_0, i_13_479_3847_0, i_13_479_3892_0, i_13_479_3909_0,
    i_13_479_3911_0, i_13_479_4056_0, i_13_479_4217_0, i_13_479_4236_0,
    i_13_479_4255_0, i_13_479_4273_0, i_13_479_4399_0, i_13_479_4546_0;
  output o_13_479_0_0;
  assign o_13_479_0_0 = ~((~i_13_479_3345_0 & ((~i_13_479_385_0 & ~i_13_479_466_0 & ~i_13_479_1995_0 & ~i_13_479_2058_0) | (~i_13_479_940_0 & i_13_479_2617_0 & ~i_13_479_3399_0))) | (~i_13_479_3346_0 & ~i_13_479_4056_0 & i_13_479_4236_0) | (i_13_479_940_0 & ~i_13_479_4273_0));
endmodule



// Benchmark "kernel_13_480" written by ABC on Sun Jul 19 10:52:02 2020

module kernel_13_480 ( 
    i_13_480_283_0, i_13_480_287_0, i_13_480_371_0, i_13_480_382_0,
    i_13_480_383_0, i_13_480_385_0, i_13_480_443_0, i_13_480_524_0,
    i_13_480_583_0, i_13_480_655_0, i_13_480_692_0, i_13_480_794_0,
    i_13_480_839_0, i_13_480_848_0, i_13_480_935_0, i_13_480_1018_0,
    i_13_480_1019_0, i_13_480_1088_0, i_13_480_1099_0, i_13_480_1136_0,
    i_13_480_1138_0, i_13_480_1331_0, i_13_480_1424_0, i_13_480_1441_0,
    i_13_480_1442_0, i_13_480_1496_0, i_13_480_1508_0, i_13_480_1520_0,
    i_13_480_1594_0, i_13_480_1630_0, i_13_480_1631_0, i_13_480_1639_0,
    i_13_480_1742_0, i_13_480_1792_0, i_13_480_1793_0, i_13_480_1799_0,
    i_13_480_1834_0, i_13_480_1999_0, i_13_480_2000_0, i_13_480_2003_0,
    i_13_480_2008_0, i_13_480_2050_0, i_13_480_2197_0, i_13_480_2198_0,
    i_13_480_2231_0, i_13_480_2233_0, i_13_480_2234_0, i_13_480_2269_0,
    i_13_480_2273_0, i_13_480_2411_0, i_13_480_2422_0, i_13_480_2459_0,
    i_13_480_2461_0, i_13_480_2462_0, i_13_480_2539_0, i_13_480_2540_0,
    i_13_480_2615_0, i_13_480_2852_0, i_13_480_2917_0, i_13_480_2918_0,
    i_13_480_2959_0, i_13_480_2987_0, i_13_480_3023_0, i_13_480_3032_0,
    i_13_480_3076_0, i_13_480_3134_0, i_13_480_3143_0, i_13_480_3169_0,
    i_13_480_3215_0, i_13_480_3247_0, i_13_480_3262_0, i_13_480_3304_0,
    i_13_480_3329_0, i_13_480_3350_0, i_13_480_3401_0, i_13_480_3686_0,
    i_13_480_3727_0, i_13_480_3728_0, i_13_480_3731_0, i_13_480_3871_0,
    i_13_480_3872_0, i_13_480_3907_0, i_13_480_3908_0, i_13_480_4007_0,
    i_13_480_4016_0, i_13_480_4018_0, i_13_480_4093_0, i_13_480_4100_0,
    i_13_480_4121_0, i_13_480_4204_0, i_13_480_4259_0, i_13_480_4339_0,
    i_13_480_4417_0, i_13_480_4513_0, i_13_480_4556_0, i_13_480_4558_0,
    i_13_480_4559_0, i_13_480_4571_0, i_13_480_4600_0, i_13_480_4601_0,
    o_13_480_0_0  );
  input  i_13_480_283_0, i_13_480_287_0, i_13_480_371_0, i_13_480_382_0,
    i_13_480_383_0, i_13_480_385_0, i_13_480_443_0, i_13_480_524_0,
    i_13_480_583_0, i_13_480_655_0, i_13_480_692_0, i_13_480_794_0,
    i_13_480_839_0, i_13_480_848_0, i_13_480_935_0, i_13_480_1018_0,
    i_13_480_1019_0, i_13_480_1088_0, i_13_480_1099_0, i_13_480_1136_0,
    i_13_480_1138_0, i_13_480_1331_0, i_13_480_1424_0, i_13_480_1441_0,
    i_13_480_1442_0, i_13_480_1496_0, i_13_480_1508_0, i_13_480_1520_0,
    i_13_480_1594_0, i_13_480_1630_0, i_13_480_1631_0, i_13_480_1639_0,
    i_13_480_1742_0, i_13_480_1792_0, i_13_480_1793_0, i_13_480_1799_0,
    i_13_480_1834_0, i_13_480_1999_0, i_13_480_2000_0, i_13_480_2003_0,
    i_13_480_2008_0, i_13_480_2050_0, i_13_480_2197_0, i_13_480_2198_0,
    i_13_480_2231_0, i_13_480_2233_0, i_13_480_2234_0, i_13_480_2269_0,
    i_13_480_2273_0, i_13_480_2411_0, i_13_480_2422_0, i_13_480_2459_0,
    i_13_480_2461_0, i_13_480_2462_0, i_13_480_2539_0, i_13_480_2540_0,
    i_13_480_2615_0, i_13_480_2852_0, i_13_480_2917_0, i_13_480_2918_0,
    i_13_480_2959_0, i_13_480_2987_0, i_13_480_3023_0, i_13_480_3032_0,
    i_13_480_3076_0, i_13_480_3134_0, i_13_480_3143_0, i_13_480_3169_0,
    i_13_480_3215_0, i_13_480_3247_0, i_13_480_3262_0, i_13_480_3304_0,
    i_13_480_3329_0, i_13_480_3350_0, i_13_480_3401_0, i_13_480_3686_0,
    i_13_480_3727_0, i_13_480_3728_0, i_13_480_3731_0, i_13_480_3871_0,
    i_13_480_3872_0, i_13_480_3907_0, i_13_480_3908_0, i_13_480_4007_0,
    i_13_480_4016_0, i_13_480_4018_0, i_13_480_4093_0, i_13_480_4100_0,
    i_13_480_4121_0, i_13_480_4204_0, i_13_480_4259_0, i_13_480_4339_0,
    i_13_480_4417_0, i_13_480_4513_0, i_13_480_4556_0, i_13_480_4558_0,
    i_13_480_4559_0, i_13_480_4571_0, i_13_480_4600_0, i_13_480_4601_0;
  output o_13_480_0_0;
  assign o_13_480_0_0 = ~((~i_13_480_2539_0 & ~i_13_480_4556_0) | (~i_13_480_3215_0 & ~i_13_480_3908_0) | (~i_13_480_2459_0 & ~i_13_480_2917_0) | (~i_13_480_2918_0 & ~i_13_480_3871_0 & ~i_13_480_4558_0));
endmodule



// Benchmark "kernel_13_481" written by ABC on Sun Jul 19 10:52:02 2020

module kernel_13_481 ( 
    i_13_481_61_0, i_13_481_118_0, i_13_481_130_0, i_13_481_136_0,
    i_13_481_168_0, i_13_481_282_0, i_13_481_312_0, i_13_481_357_0,
    i_13_481_364_0, i_13_481_492_0, i_13_481_528_0, i_13_481_645_0,
    i_13_481_646_0, i_13_481_663_0, i_13_481_717_0, i_13_481_726_0,
    i_13_481_826_0, i_13_481_888_0, i_13_481_958_0, i_13_481_1021_0,
    i_13_481_1101_0, i_13_481_1228_0, i_13_481_1230_0, i_13_481_1257_0,
    i_13_481_1258_0, i_13_481_1303_0, i_13_481_1308_0, i_13_481_1320_0,
    i_13_481_1407_0, i_13_481_1446_0, i_13_481_1491_0, i_13_481_1492_0,
    i_13_481_1500_0, i_13_481_1501_0, i_13_481_1554_0, i_13_481_1555_0,
    i_13_481_1572_0, i_13_481_1599_0, i_13_481_1641_0, i_13_481_1642_0,
    i_13_481_1699_0, i_13_481_1759_0, i_13_481_1795_0, i_13_481_1804_0,
    i_13_481_1806_0, i_13_481_1807_0, i_13_481_1959_0, i_13_481_1960_0,
    i_13_481_2014_0, i_13_481_2103_0, i_13_481_2145_0, i_13_481_2175_0,
    i_13_481_2193_0, i_13_481_2202_0, i_13_481_2205_0, i_13_481_2238_0,
    i_13_481_2239_0, i_13_481_2247_0, i_13_481_2430_0, i_13_481_2431_0,
    i_13_481_2445_0, i_13_481_2446_0, i_13_481_2508_0, i_13_481_2509_0,
    i_13_481_2514_0, i_13_481_2536_0, i_13_481_2608_0, i_13_481_2698_0,
    i_13_481_2818_0, i_13_481_2824_0, i_13_481_2937_0, i_13_481_2938_0,
    i_13_481_3244_0, i_13_481_3310_0, i_13_481_3420_0, i_13_481_3423_0,
    i_13_481_3426_0, i_13_481_3489_0, i_13_481_3543_0, i_13_481_3612_0,
    i_13_481_3639_0, i_13_481_3756_0, i_13_481_3805_0, i_13_481_3858_0,
    i_13_481_3859_0, i_13_481_3919_0, i_13_481_3936_0, i_13_481_3984_0,
    i_13_481_3985_0, i_13_481_4012_0, i_13_481_4065_0, i_13_481_4066_0,
    i_13_481_4215_0, i_13_481_4234_0, i_13_481_4272_0, i_13_481_4315_0,
    i_13_481_4380_0, i_13_481_4432_0, i_13_481_4512_0, i_13_481_4536_0,
    o_13_481_0_0  );
  input  i_13_481_61_0, i_13_481_118_0, i_13_481_130_0, i_13_481_136_0,
    i_13_481_168_0, i_13_481_282_0, i_13_481_312_0, i_13_481_357_0,
    i_13_481_364_0, i_13_481_492_0, i_13_481_528_0, i_13_481_645_0,
    i_13_481_646_0, i_13_481_663_0, i_13_481_717_0, i_13_481_726_0,
    i_13_481_826_0, i_13_481_888_0, i_13_481_958_0, i_13_481_1021_0,
    i_13_481_1101_0, i_13_481_1228_0, i_13_481_1230_0, i_13_481_1257_0,
    i_13_481_1258_0, i_13_481_1303_0, i_13_481_1308_0, i_13_481_1320_0,
    i_13_481_1407_0, i_13_481_1446_0, i_13_481_1491_0, i_13_481_1492_0,
    i_13_481_1500_0, i_13_481_1501_0, i_13_481_1554_0, i_13_481_1555_0,
    i_13_481_1572_0, i_13_481_1599_0, i_13_481_1641_0, i_13_481_1642_0,
    i_13_481_1699_0, i_13_481_1759_0, i_13_481_1795_0, i_13_481_1804_0,
    i_13_481_1806_0, i_13_481_1807_0, i_13_481_1959_0, i_13_481_1960_0,
    i_13_481_2014_0, i_13_481_2103_0, i_13_481_2145_0, i_13_481_2175_0,
    i_13_481_2193_0, i_13_481_2202_0, i_13_481_2205_0, i_13_481_2238_0,
    i_13_481_2239_0, i_13_481_2247_0, i_13_481_2430_0, i_13_481_2431_0,
    i_13_481_2445_0, i_13_481_2446_0, i_13_481_2508_0, i_13_481_2509_0,
    i_13_481_2514_0, i_13_481_2536_0, i_13_481_2608_0, i_13_481_2698_0,
    i_13_481_2818_0, i_13_481_2824_0, i_13_481_2937_0, i_13_481_2938_0,
    i_13_481_3244_0, i_13_481_3310_0, i_13_481_3420_0, i_13_481_3423_0,
    i_13_481_3426_0, i_13_481_3489_0, i_13_481_3543_0, i_13_481_3612_0,
    i_13_481_3639_0, i_13_481_3756_0, i_13_481_3805_0, i_13_481_3858_0,
    i_13_481_3859_0, i_13_481_3919_0, i_13_481_3936_0, i_13_481_3984_0,
    i_13_481_3985_0, i_13_481_4012_0, i_13_481_4065_0, i_13_481_4066_0,
    i_13_481_4215_0, i_13_481_4234_0, i_13_481_4272_0, i_13_481_4315_0,
    i_13_481_4380_0, i_13_481_4432_0, i_13_481_4512_0, i_13_481_4536_0;
  output o_13_481_0_0;
  assign o_13_481_0_0 = ~((~i_13_481_2938_0 & ~i_13_481_3984_0) | (~i_13_481_1257_0 & ~i_13_481_1554_0) | (~i_13_481_1491_0 & ~i_13_481_1795_0 & ~i_13_481_3859_0));
endmodule



// Benchmark "kernel_13_482" written by ABC on Sun Jul 19 10:52:03 2020

module kernel_13_482 ( 
    i_13_482_30_0, i_13_482_73_0, i_13_482_90_0, i_13_482_103_0,
    i_13_482_108_0, i_13_482_265_0, i_13_482_270_0, i_13_482_363_0,
    i_13_482_561_0, i_13_482_603_0, i_13_482_669_0, i_13_482_670_0,
    i_13_482_675_0, i_13_482_679_0, i_13_482_685_0, i_13_482_742_0,
    i_13_482_814_0, i_13_482_865_0, i_13_482_945_0, i_13_482_1083_0,
    i_13_482_1143_0, i_13_482_1215_0, i_13_482_1216_0, i_13_482_1284_0,
    i_13_482_1285_0, i_13_482_1324_0, i_13_482_1470_0, i_13_482_1515_0,
    i_13_482_1516_0, i_13_482_1620_0, i_13_482_1623_0, i_13_482_1801_0,
    i_13_482_1836_0, i_13_482_1837_0, i_13_482_1839_0, i_13_482_1840_0,
    i_13_482_1857_0, i_13_482_1912_0, i_13_482_2019_0, i_13_482_2133_0,
    i_13_482_2169_0, i_13_482_2275_0, i_13_482_2344_0, i_13_482_2434_0,
    i_13_482_2493_0, i_13_482_2496_0, i_13_482_2497_0, i_13_482_2529_0,
    i_13_482_2559_0, i_13_482_2610_0, i_13_482_2712_0, i_13_482_2934_0,
    i_13_482_2935_0, i_13_482_2955_0, i_13_482_3043_0, i_13_482_3096_0,
    i_13_482_3097_0, i_13_482_3099_0, i_13_482_3100_0, i_13_482_3142_0,
    i_13_482_3144_0, i_13_482_3149_0, i_13_482_3160_0, i_13_482_3162_0,
    i_13_482_3289_0, i_13_482_3415_0, i_13_482_3455_0, i_13_482_3475_0,
    i_13_482_3535_0, i_13_482_3546_0, i_13_482_3549_0, i_13_482_3567_0,
    i_13_482_3684_0, i_13_482_3738_0, i_13_482_3762_0, i_13_482_3763_0,
    i_13_482_3792_0, i_13_482_3802_0, i_13_482_3870_0, i_13_482_3936_0,
    i_13_482_3981_0, i_13_482_4005_0, i_13_482_4042_0, i_13_482_4045_0,
    i_13_482_4116_0, i_13_482_4123_0, i_13_482_4159_0, i_13_482_4188_0,
    i_13_482_4249_0, i_13_482_4260_0, i_13_482_4266_0, i_13_482_4324_0,
    i_13_482_4350_0, i_13_482_4365_0, i_13_482_4378_0, i_13_482_4413_0,
    i_13_482_4491_0, i_13_482_4512_0, i_13_482_4539_0, i_13_482_4557_0,
    o_13_482_0_0  );
  input  i_13_482_30_0, i_13_482_73_0, i_13_482_90_0, i_13_482_103_0,
    i_13_482_108_0, i_13_482_265_0, i_13_482_270_0, i_13_482_363_0,
    i_13_482_561_0, i_13_482_603_0, i_13_482_669_0, i_13_482_670_0,
    i_13_482_675_0, i_13_482_679_0, i_13_482_685_0, i_13_482_742_0,
    i_13_482_814_0, i_13_482_865_0, i_13_482_945_0, i_13_482_1083_0,
    i_13_482_1143_0, i_13_482_1215_0, i_13_482_1216_0, i_13_482_1284_0,
    i_13_482_1285_0, i_13_482_1324_0, i_13_482_1470_0, i_13_482_1515_0,
    i_13_482_1516_0, i_13_482_1620_0, i_13_482_1623_0, i_13_482_1801_0,
    i_13_482_1836_0, i_13_482_1837_0, i_13_482_1839_0, i_13_482_1840_0,
    i_13_482_1857_0, i_13_482_1912_0, i_13_482_2019_0, i_13_482_2133_0,
    i_13_482_2169_0, i_13_482_2275_0, i_13_482_2344_0, i_13_482_2434_0,
    i_13_482_2493_0, i_13_482_2496_0, i_13_482_2497_0, i_13_482_2529_0,
    i_13_482_2559_0, i_13_482_2610_0, i_13_482_2712_0, i_13_482_2934_0,
    i_13_482_2935_0, i_13_482_2955_0, i_13_482_3043_0, i_13_482_3096_0,
    i_13_482_3097_0, i_13_482_3099_0, i_13_482_3100_0, i_13_482_3142_0,
    i_13_482_3144_0, i_13_482_3149_0, i_13_482_3160_0, i_13_482_3162_0,
    i_13_482_3289_0, i_13_482_3415_0, i_13_482_3455_0, i_13_482_3475_0,
    i_13_482_3535_0, i_13_482_3546_0, i_13_482_3549_0, i_13_482_3567_0,
    i_13_482_3684_0, i_13_482_3738_0, i_13_482_3762_0, i_13_482_3763_0,
    i_13_482_3792_0, i_13_482_3802_0, i_13_482_3870_0, i_13_482_3936_0,
    i_13_482_3981_0, i_13_482_4005_0, i_13_482_4042_0, i_13_482_4045_0,
    i_13_482_4116_0, i_13_482_4123_0, i_13_482_4159_0, i_13_482_4188_0,
    i_13_482_4249_0, i_13_482_4260_0, i_13_482_4266_0, i_13_482_4324_0,
    i_13_482_4350_0, i_13_482_4365_0, i_13_482_4378_0, i_13_482_4413_0,
    i_13_482_4491_0, i_13_482_4512_0, i_13_482_4539_0, i_13_482_4557_0;
  output o_13_482_0_0;
  assign o_13_482_0_0 = ~(~i_13_482_3100_0 | (~i_13_482_1143_0 & ~i_13_482_4005_0) | (~i_13_482_1620_0 & ~i_13_482_3144_0));
endmodule



// Benchmark "kernel_13_483" written by ABC on Sun Jul 19 10:52:04 2020

module kernel_13_483 ( 
    i_13_483_22_0, i_13_483_45_0, i_13_483_48_0, i_13_483_240_0,
    i_13_483_319_0, i_13_483_370_0, i_13_483_450_0, i_13_483_451_0,
    i_13_483_453_0, i_13_483_561_0, i_13_483_587_0, i_13_483_598_0,
    i_13_483_622_0, i_13_483_928_0, i_13_483_940_0, i_13_483_1063_0,
    i_13_483_1064_0, i_13_483_1091_0, i_13_483_1244_0, i_13_483_1265_0,
    i_13_483_1297_0, i_13_483_1319_0, i_13_483_1342_0, i_13_483_1460_0,
    i_13_483_1468_0, i_13_483_1486_0, i_13_483_1495_0, i_13_483_1530_0,
    i_13_483_1566_0, i_13_483_1568_0, i_13_483_1569_0, i_13_483_1593_0,
    i_13_483_1594_0, i_13_483_1764_0, i_13_483_1774_0, i_13_483_1809_0,
    i_13_483_1810_0, i_13_483_1848_0, i_13_483_1884_0, i_13_483_1927_0,
    i_13_483_1959_0, i_13_483_1999_0, i_13_483_2107_0, i_13_483_2233_0,
    i_13_483_2278_0, i_13_483_2451_0, i_13_483_2452_0, i_13_483_2488_0,
    i_13_483_2543_0, i_13_483_2544_0, i_13_483_2617_0, i_13_483_2709_0,
    i_13_483_2710_0, i_13_483_2784_0, i_13_483_2882_0, i_13_483_2885_0,
    i_13_483_2886_0, i_13_483_2935_0, i_13_483_3016_0, i_13_483_3121_0,
    i_13_483_3213_0, i_13_483_3214_0, i_13_483_3216_0, i_13_483_3231_0,
    i_13_483_3244_0, i_13_483_3268_0, i_13_483_3286_0, i_13_483_3308_0,
    i_13_483_3340_0, i_13_483_3366_0, i_13_483_3367_0, i_13_483_3378_0,
    i_13_483_3388_0, i_13_483_3460_0, i_13_483_3532_0, i_13_483_3612_0,
    i_13_483_3688_0, i_13_483_3731_0, i_13_483_3763_0, i_13_483_3803_0,
    i_13_483_3817_0, i_13_483_3820_0, i_13_483_3876_0, i_13_483_3891_0,
    i_13_483_3999_0, i_13_483_4042_0, i_13_483_4063_0, i_13_483_4086_0,
    i_13_483_4087_0, i_13_483_4214_0, i_13_483_4266_0, i_13_483_4267_0,
    i_13_483_4269_0, i_13_483_4270_0, i_13_483_4313_0, i_13_483_4362_0,
    i_13_483_4371_0, i_13_483_4415_0, i_13_483_4459_0, i_13_483_4560_0,
    o_13_483_0_0  );
  input  i_13_483_22_0, i_13_483_45_0, i_13_483_48_0, i_13_483_240_0,
    i_13_483_319_0, i_13_483_370_0, i_13_483_450_0, i_13_483_451_0,
    i_13_483_453_0, i_13_483_561_0, i_13_483_587_0, i_13_483_598_0,
    i_13_483_622_0, i_13_483_928_0, i_13_483_940_0, i_13_483_1063_0,
    i_13_483_1064_0, i_13_483_1091_0, i_13_483_1244_0, i_13_483_1265_0,
    i_13_483_1297_0, i_13_483_1319_0, i_13_483_1342_0, i_13_483_1460_0,
    i_13_483_1468_0, i_13_483_1486_0, i_13_483_1495_0, i_13_483_1530_0,
    i_13_483_1566_0, i_13_483_1568_0, i_13_483_1569_0, i_13_483_1593_0,
    i_13_483_1594_0, i_13_483_1764_0, i_13_483_1774_0, i_13_483_1809_0,
    i_13_483_1810_0, i_13_483_1848_0, i_13_483_1884_0, i_13_483_1927_0,
    i_13_483_1959_0, i_13_483_1999_0, i_13_483_2107_0, i_13_483_2233_0,
    i_13_483_2278_0, i_13_483_2451_0, i_13_483_2452_0, i_13_483_2488_0,
    i_13_483_2543_0, i_13_483_2544_0, i_13_483_2617_0, i_13_483_2709_0,
    i_13_483_2710_0, i_13_483_2784_0, i_13_483_2882_0, i_13_483_2885_0,
    i_13_483_2886_0, i_13_483_2935_0, i_13_483_3016_0, i_13_483_3121_0,
    i_13_483_3213_0, i_13_483_3214_0, i_13_483_3216_0, i_13_483_3231_0,
    i_13_483_3244_0, i_13_483_3268_0, i_13_483_3286_0, i_13_483_3308_0,
    i_13_483_3340_0, i_13_483_3366_0, i_13_483_3367_0, i_13_483_3378_0,
    i_13_483_3388_0, i_13_483_3460_0, i_13_483_3532_0, i_13_483_3612_0,
    i_13_483_3688_0, i_13_483_3731_0, i_13_483_3763_0, i_13_483_3803_0,
    i_13_483_3817_0, i_13_483_3820_0, i_13_483_3876_0, i_13_483_3891_0,
    i_13_483_3999_0, i_13_483_4042_0, i_13_483_4063_0, i_13_483_4086_0,
    i_13_483_4087_0, i_13_483_4214_0, i_13_483_4266_0, i_13_483_4267_0,
    i_13_483_4269_0, i_13_483_4270_0, i_13_483_4313_0, i_13_483_4362_0,
    i_13_483_4371_0, i_13_483_4415_0, i_13_483_4459_0, i_13_483_4560_0;
  output o_13_483_0_0;
  assign o_13_483_0_0 = ~(~i_13_483_3817_0 | (~i_13_483_1566_0 & ~i_13_483_3244_0));
endmodule



// Benchmark "kernel_13_484" written by ABC on Sun Jul 19 10:52:04 2020

module kernel_13_484 ( 
    i_13_484_11_0, i_13_484_46_0, i_13_484_47_0, i_13_484_67_0,
    i_13_484_70_0, i_13_484_71_0, i_13_484_155_0, i_13_484_184_0,
    i_13_484_185_0, i_13_484_211_0, i_13_484_235_0, i_13_484_403_0,
    i_13_484_466_0, i_13_484_518_0, i_13_484_521_0, i_13_484_599_0,
    i_13_484_678_0, i_13_484_695_0, i_13_484_698_0, i_13_484_745_0,
    i_13_484_760_0, i_13_484_763_0, i_13_484_764_0, i_13_484_812_0,
    i_13_484_1062_0, i_13_484_1129_0, i_13_484_1132_0, i_13_484_1133_0,
    i_13_484_1189_0, i_13_484_1208_0, i_13_484_1210_0, i_13_484_1211_0,
    i_13_484_1310_0, i_13_484_1313_0, i_13_484_1394_0, i_13_484_1403_0,
    i_13_484_1506_0, i_13_484_1522_0, i_13_484_1548_0, i_13_484_1604_0,
    i_13_484_1659_0, i_13_484_1661_0, i_13_484_1673_0, i_13_484_1727_0,
    i_13_484_1927_0, i_13_484_1931_0, i_13_484_1945_0, i_13_484_1964_0,
    i_13_484_1967_0, i_13_484_2025_0, i_13_484_2097_0, i_13_484_2115_0,
    i_13_484_2132_0, i_13_484_2143_0, i_13_484_2316_0, i_13_484_2402_0,
    i_13_484_2552_0, i_13_484_2722_0, i_13_484_2767_0, i_13_484_2783_0,
    i_13_484_2848_0, i_13_484_2881_0, i_13_484_2884_0, i_13_484_3077_0,
    i_13_484_3091_0, i_13_484_3172_0, i_13_484_3251_0, i_13_484_3289_0,
    i_13_484_3308_0, i_13_484_3366_0, i_13_484_3370_0, i_13_484_3458_0,
    i_13_484_3542_0, i_13_484_3547_0, i_13_484_3591_0, i_13_484_3595_0,
    i_13_484_3611_0, i_13_484_3631_0, i_13_484_3636_0, i_13_484_3638_0,
    i_13_484_3641_0, i_13_484_3668_0, i_13_484_3752_0, i_13_484_3780_0,
    i_13_484_3890_0, i_13_484_3895_0, i_13_484_3898_0, i_13_484_3919_0,
    i_13_484_4036_0, i_13_484_4039_0, i_13_484_4214_0, i_13_484_4230_0,
    i_13_484_4270_0, i_13_484_4322_0, i_13_484_4332_0, i_13_484_4368_0,
    i_13_484_4397_0, i_13_484_4594_0, i_13_484_4595_0, i_13_484_4607_0,
    o_13_484_0_0  );
  input  i_13_484_11_0, i_13_484_46_0, i_13_484_47_0, i_13_484_67_0,
    i_13_484_70_0, i_13_484_71_0, i_13_484_155_0, i_13_484_184_0,
    i_13_484_185_0, i_13_484_211_0, i_13_484_235_0, i_13_484_403_0,
    i_13_484_466_0, i_13_484_518_0, i_13_484_521_0, i_13_484_599_0,
    i_13_484_678_0, i_13_484_695_0, i_13_484_698_0, i_13_484_745_0,
    i_13_484_760_0, i_13_484_763_0, i_13_484_764_0, i_13_484_812_0,
    i_13_484_1062_0, i_13_484_1129_0, i_13_484_1132_0, i_13_484_1133_0,
    i_13_484_1189_0, i_13_484_1208_0, i_13_484_1210_0, i_13_484_1211_0,
    i_13_484_1310_0, i_13_484_1313_0, i_13_484_1394_0, i_13_484_1403_0,
    i_13_484_1506_0, i_13_484_1522_0, i_13_484_1548_0, i_13_484_1604_0,
    i_13_484_1659_0, i_13_484_1661_0, i_13_484_1673_0, i_13_484_1727_0,
    i_13_484_1927_0, i_13_484_1931_0, i_13_484_1945_0, i_13_484_1964_0,
    i_13_484_1967_0, i_13_484_2025_0, i_13_484_2097_0, i_13_484_2115_0,
    i_13_484_2132_0, i_13_484_2143_0, i_13_484_2316_0, i_13_484_2402_0,
    i_13_484_2552_0, i_13_484_2722_0, i_13_484_2767_0, i_13_484_2783_0,
    i_13_484_2848_0, i_13_484_2881_0, i_13_484_2884_0, i_13_484_3077_0,
    i_13_484_3091_0, i_13_484_3172_0, i_13_484_3251_0, i_13_484_3289_0,
    i_13_484_3308_0, i_13_484_3366_0, i_13_484_3370_0, i_13_484_3458_0,
    i_13_484_3542_0, i_13_484_3547_0, i_13_484_3591_0, i_13_484_3595_0,
    i_13_484_3611_0, i_13_484_3631_0, i_13_484_3636_0, i_13_484_3638_0,
    i_13_484_3641_0, i_13_484_3668_0, i_13_484_3752_0, i_13_484_3780_0,
    i_13_484_3890_0, i_13_484_3895_0, i_13_484_3898_0, i_13_484_3919_0,
    i_13_484_4036_0, i_13_484_4039_0, i_13_484_4214_0, i_13_484_4230_0,
    i_13_484_4270_0, i_13_484_4322_0, i_13_484_4332_0, i_13_484_4368_0,
    i_13_484_4397_0, i_13_484_4594_0, i_13_484_4595_0, i_13_484_4607_0;
  output o_13_484_0_0;
  assign o_13_484_0_0 = ~((~i_13_484_518_0 & ((i_13_484_184_0 & ~i_13_484_1661_0) | (~i_13_484_812_0 & ~i_13_484_1945_0 & i_13_484_2881_0))) | (~i_13_484_764_0 & ~i_13_484_2783_0 & ((i_13_484_3289_0 & ~i_13_484_3542_0 & ~i_13_484_3547_0) | (i_13_484_3172_0 & ~i_13_484_4214_0))) | (~i_13_484_521_0 & i_13_484_1210_0 & i_13_484_2132_0) | (~i_13_484_1211_0 & ~i_13_484_2767_0) | (~i_13_484_698_0 & ~i_13_484_3289_0 & ~i_13_484_3898_0 & ~i_13_484_4214_0 & ~i_13_484_4397_0));
endmodule



// Benchmark "kernel_13_485" written by ABC on Sun Jul 19 10:52:05 2020

module kernel_13_485 ( 
    i_13_485_52_0, i_13_485_53_0, i_13_485_71_0, i_13_485_130_0,
    i_13_485_175_0, i_13_485_176_0, i_13_485_251_0, i_13_485_276_0,
    i_13_485_373_0, i_13_485_479_0, i_13_485_518_0, i_13_485_520_0,
    i_13_485_521_0, i_13_485_527_0, i_13_485_584_0, i_13_485_616_0,
    i_13_485_655_0, i_13_485_656_0, i_13_485_679_0, i_13_485_680_0,
    i_13_485_692_0, i_13_485_718_0, i_13_485_841_0, i_13_485_844_0,
    i_13_485_985_0, i_13_485_1084_0, i_13_485_1268_0, i_13_485_1330_0,
    i_13_485_1331_0, i_13_485_1435_0, i_13_485_1492_0, i_13_485_1573_0,
    i_13_485_1574_0, i_13_485_1663_0, i_13_485_1723_0, i_13_485_1754_0,
    i_13_485_1786_0, i_13_485_1814_0, i_13_485_1943_0, i_13_485_2024_0,
    i_13_485_2056_0, i_13_485_2057_0, i_13_485_2059_0, i_13_485_2060_0,
    i_13_485_2185_0, i_13_485_2186_0, i_13_485_2209_0, i_13_485_2239_0,
    i_13_485_2321_0, i_13_485_2455_0, i_13_485_2461_0, i_13_485_2507_0,
    i_13_485_2509_0, i_13_485_2510_0, i_13_485_2651_0, i_13_485_2698_0,
    i_13_485_2699_0, i_13_485_2733_0, i_13_485_2752_0, i_13_485_2753_0,
    i_13_485_2959_0, i_13_485_3068_0, i_13_485_3077_0, i_13_485_3100_0,
    i_13_485_3112_0, i_13_485_3163_0, i_13_485_3217_0, i_13_485_3256_0,
    i_13_485_3292_0, i_13_485_3373_0, i_13_485_3374_0, i_13_485_3406_0,
    i_13_485_3526_0, i_13_485_3571_0, i_13_485_3572_0, i_13_485_3613_0,
    i_13_485_3662_0, i_13_485_3725_0, i_13_485_3749_0, i_13_485_3767_0,
    i_13_485_3769_0, i_13_485_3830_0, i_13_485_3847_0, i_13_485_3874_0,
    i_13_485_3877_0, i_13_485_3991_0, i_13_485_3995_0, i_13_485_4009_0,
    i_13_485_4021_0, i_13_485_4022_0, i_13_485_4048_0, i_13_485_4127_0,
    i_13_485_4157_0, i_13_485_4189_0, i_13_485_4318_0, i_13_485_4319_0,
    i_13_485_4558_0, i_13_485_4598_0, i_13_485_4603_0, i_13_485_4604_0,
    o_13_485_0_0  );
  input  i_13_485_52_0, i_13_485_53_0, i_13_485_71_0, i_13_485_130_0,
    i_13_485_175_0, i_13_485_176_0, i_13_485_251_0, i_13_485_276_0,
    i_13_485_373_0, i_13_485_479_0, i_13_485_518_0, i_13_485_520_0,
    i_13_485_521_0, i_13_485_527_0, i_13_485_584_0, i_13_485_616_0,
    i_13_485_655_0, i_13_485_656_0, i_13_485_679_0, i_13_485_680_0,
    i_13_485_692_0, i_13_485_718_0, i_13_485_841_0, i_13_485_844_0,
    i_13_485_985_0, i_13_485_1084_0, i_13_485_1268_0, i_13_485_1330_0,
    i_13_485_1331_0, i_13_485_1435_0, i_13_485_1492_0, i_13_485_1573_0,
    i_13_485_1574_0, i_13_485_1663_0, i_13_485_1723_0, i_13_485_1754_0,
    i_13_485_1786_0, i_13_485_1814_0, i_13_485_1943_0, i_13_485_2024_0,
    i_13_485_2056_0, i_13_485_2057_0, i_13_485_2059_0, i_13_485_2060_0,
    i_13_485_2185_0, i_13_485_2186_0, i_13_485_2209_0, i_13_485_2239_0,
    i_13_485_2321_0, i_13_485_2455_0, i_13_485_2461_0, i_13_485_2507_0,
    i_13_485_2509_0, i_13_485_2510_0, i_13_485_2651_0, i_13_485_2698_0,
    i_13_485_2699_0, i_13_485_2733_0, i_13_485_2752_0, i_13_485_2753_0,
    i_13_485_2959_0, i_13_485_3068_0, i_13_485_3077_0, i_13_485_3100_0,
    i_13_485_3112_0, i_13_485_3163_0, i_13_485_3217_0, i_13_485_3256_0,
    i_13_485_3292_0, i_13_485_3373_0, i_13_485_3374_0, i_13_485_3406_0,
    i_13_485_3526_0, i_13_485_3571_0, i_13_485_3572_0, i_13_485_3613_0,
    i_13_485_3662_0, i_13_485_3725_0, i_13_485_3749_0, i_13_485_3767_0,
    i_13_485_3769_0, i_13_485_3830_0, i_13_485_3847_0, i_13_485_3874_0,
    i_13_485_3877_0, i_13_485_3991_0, i_13_485_3995_0, i_13_485_4009_0,
    i_13_485_4021_0, i_13_485_4022_0, i_13_485_4048_0, i_13_485_4127_0,
    i_13_485_4157_0, i_13_485_4189_0, i_13_485_4318_0, i_13_485_4319_0,
    i_13_485_4558_0, i_13_485_4598_0, i_13_485_4603_0, i_13_485_4604_0;
  output o_13_485_0_0;
  assign o_13_485_0_0 = ~((~i_13_485_53_0 & ~i_13_485_2698_0) | (~i_13_485_2056_0 & ~i_13_485_4157_0 & ~i_13_485_4189_0) | (~i_13_485_521_0 & ~i_13_485_1573_0 & ~i_13_485_2060_0 & ~i_13_485_4319_0));
endmodule



// Benchmark "kernel_13_486" written by ABC on Sun Jul 19 10:52:06 2020

module kernel_13_486 ( 
    i_13_486_70_0, i_13_486_75_0, i_13_486_120_0, i_13_486_121_0,
    i_13_486_184_0, i_13_486_244_0, i_13_486_333_0, i_13_486_414_0,
    i_13_486_423_0, i_13_486_459_0, i_13_486_517_0, i_13_486_522_0,
    i_13_486_523_0, i_13_486_524_0, i_13_486_525_0, i_13_486_526_0,
    i_13_486_532_0, i_13_486_571_0, i_13_486_585_0, i_13_486_588_0,
    i_13_486_670_0, i_13_486_697_0, i_13_486_759_0, i_13_486_1057_0,
    i_13_486_1066_0, i_13_486_1116_0, i_13_486_1207_0, i_13_486_1216_0,
    i_13_486_1306_0, i_13_486_1307_0, i_13_486_1314_0, i_13_486_1317_0,
    i_13_486_1341_0, i_13_486_1342_0, i_13_486_1389_0, i_13_486_1399_0,
    i_13_486_1440_0, i_13_486_1441_0, i_13_486_1444_0, i_13_486_1494_0,
    i_13_486_1515_0, i_13_486_1602_0, i_13_486_1603_0, i_13_486_1774_0,
    i_13_486_1887_0, i_13_486_1930_0, i_13_486_1944_0, i_13_486_1945_0,
    i_13_486_1998_0, i_13_486_2001_0, i_13_486_2025_0, i_13_486_2026_0,
    i_13_486_2124_0, i_13_486_2125_0, i_13_486_2196_0, i_13_486_2197_0,
    i_13_486_2278_0, i_13_486_2445_0, i_13_486_2533_0, i_13_486_2710_0,
    i_13_486_2766_0, i_13_486_2781_0, i_13_486_2902_0, i_13_486_2916_0,
    i_13_486_2917_0, i_13_486_2918_0, i_13_486_2983_0, i_13_486_3007_0,
    i_13_486_3046_0, i_13_486_3163_0, i_13_486_3208_0, i_13_486_3366_0,
    i_13_486_3367_0, i_13_486_3396_0, i_13_486_3406_0, i_13_486_3414_0,
    i_13_486_3438_0, i_13_486_3460_0, i_13_486_3541_0, i_13_486_3559_0,
    i_13_486_3573_0, i_13_486_3575_0, i_13_486_3592_0, i_13_486_3637_0,
    i_13_486_3666_0, i_13_486_3667_0, i_13_486_3726_0, i_13_486_3766_0,
    i_13_486_3907_0, i_13_486_4096_0, i_13_486_4105_0, i_13_486_4149_0,
    i_13_486_4204_0, i_13_486_4350_0, i_13_486_4351_0, i_13_486_4392_0,
    i_13_486_4441_0, i_13_486_4446_0, i_13_486_4447_0, i_13_486_4567_0,
    o_13_486_0_0  );
  input  i_13_486_70_0, i_13_486_75_0, i_13_486_120_0, i_13_486_121_0,
    i_13_486_184_0, i_13_486_244_0, i_13_486_333_0, i_13_486_414_0,
    i_13_486_423_0, i_13_486_459_0, i_13_486_517_0, i_13_486_522_0,
    i_13_486_523_0, i_13_486_524_0, i_13_486_525_0, i_13_486_526_0,
    i_13_486_532_0, i_13_486_571_0, i_13_486_585_0, i_13_486_588_0,
    i_13_486_670_0, i_13_486_697_0, i_13_486_759_0, i_13_486_1057_0,
    i_13_486_1066_0, i_13_486_1116_0, i_13_486_1207_0, i_13_486_1216_0,
    i_13_486_1306_0, i_13_486_1307_0, i_13_486_1314_0, i_13_486_1317_0,
    i_13_486_1341_0, i_13_486_1342_0, i_13_486_1389_0, i_13_486_1399_0,
    i_13_486_1440_0, i_13_486_1441_0, i_13_486_1444_0, i_13_486_1494_0,
    i_13_486_1515_0, i_13_486_1602_0, i_13_486_1603_0, i_13_486_1774_0,
    i_13_486_1887_0, i_13_486_1930_0, i_13_486_1944_0, i_13_486_1945_0,
    i_13_486_1998_0, i_13_486_2001_0, i_13_486_2025_0, i_13_486_2026_0,
    i_13_486_2124_0, i_13_486_2125_0, i_13_486_2196_0, i_13_486_2197_0,
    i_13_486_2278_0, i_13_486_2445_0, i_13_486_2533_0, i_13_486_2710_0,
    i_13_486_2766_0, i_13_486_2781_0, i_13_486_2902_0, i_13_486_2916_0,
    i_13_486_2917_0, i_13_486_2918_0, i_13_486_2983_0, i_13_486_3007_0,
    i_13_486_3046_0, i_13_486_3163_0, i_13_486_3208_0, i_13_486_3366_0,
    i_13_486_3367_0, i_13_486_3396_0, i_13_486_3406_0, i_13_486_3414_0,
    i_13_486_3438_0, i_13_486_3460_0, i_13_486_3541_0, i_13_486_3559_0,
    i_13_486_3573_0, i_13_486_3575_0, i_13_486_3592_0, i_13_486_3637_0,
    i_13_486_3666_0, i_13_486_3667_0, i_13_486_3726_0, i_13_486_3766_0,
    i_13_486_3907_0, i_13_486_4096_0, i_13_486_4105_0, i_13_486_4149_0,
    i_13_486_4204_0, i_13_486_4350_0, i_13_486_4351_0, i_13_486_4392_0,
    i_13_486_4441_0, i_13_486_4446_0, i_13_486_4447_0, i_13_486_4567_0;
  output o_13_486_0_0;
  assign o_13_486_0_0 = ~(~i_13_486_4446_0 & ((~i_13_486_517_0 & ~i_13_486_2125_0) | (~i_13_486_1494_0 & ~i_13_486_2124_0 & ~i_13_486_2278_0) | (~i_13_486_2197_0 & ~i_13_486_3541_0 & ~i_13_486_3573_0)));
endmodule



// Benchmark "kernel_13_487" written by ABC on Sun Jul 19 10:52:07 2020

module kernel_13_487 ( 
    i_13_487_40_0, i_13_487_110_0, i_13_487_126_0, i_13_487_132_0,
    i_13_487_273_0, i_13_487_282_0, i_13_487_283_0, i_13_487_284_0,
    i_13_487_335_0, i_13_487_357_0, i_13_487_360_0, i_13_487_361_0,
    i_13_487_472_0, i_13_487_519_0, i_13_487_538_0, i_13_487_689_0,
    i_13_487_838_0, i_13_487_866_0, i_13_487_867_0, i_13_487_869_0,
    i_13_487_1096_0, i_13_487_1111_0, i_13_487_1112_0, i_13_487_1114_0,
    i_13_487_1119_0, i_13_487_1132_0, i_13_487_1243_0, i_13_487_1329_0,
    i_13_487_1430_0, i_13_487_1501_0, i_13_487_1549_0, i_13_487_1745_0,
    i_13_487_1770_0, i_13_487_1792_0, i_13_487_1795_0, i_13_487_1834_0,
    i_13_487_1858_0, i_13_487_1884_0, i_13_487_1896_0, i_13_487_2004_0,
    i_13_487_2008_0, i_13_487_2010_0, i_13_487_2017_0, i_13_487_2097_0,
    i_13_487_2113_0, i_13_487_2145_0, i_13_487_2148_0, i_13_487_2223_0,
    i_13_487_2260_0, i_13_487_2384_0, i_13_487_2461_0, i_13_487_2514_0,
    i_13_487_2537_0, i_13_487_2733_0, i_13_487_2798_0, i_13_487_2883_0,
    i_13_487_2890_0, i_13_487_3048_0, i_13_487_3057_0, i_13_487_3059_0,
    i_13_487_3076_0, i_13_487_3077_0, i_13_487_3097_0, i_13_487_3145_0,
    i_13_487_3219_0, i_13_487_3266_0, i_13_487_3286_0, i_13_487_3315_0,
    i_13_487_3348_0, i_13_487_3489_0, i_13_487_3490_0, i_13_487_3549_0,
    i_13_487_3550_0, i_13_487_3604_0, i_13_487_3671_0, i_13_487_3730_0,
    i_13_487_3735_0, i_13_487_3748_0, i_13_487_3822_0, i_13_487_3869_0,
    i_13_487_3881_0, i_13_487_3909_0, i_13_487_3910_0, i_13_487_3952_0,
    i_13_487_4018_0, i_13_487_4125_0, i_13_487_4126_0, i_13_487_4165_0,
    i_13_487_4261_0, i_13_487_4272_0, i_13_487_4330_0, i_13_487_4333_0,
    i_13_487_4362_0, i_13_487_4433_0, i_13_487_4454_0, i_13_487_4467_0,
    i_13_487_4471_0, i_13_487_4516_0, i_13_487_4565_0, i_13_487_4578_0,
    o_13_487_0_0  );
  input  i_13_487_40_0, i_13_487_110_0, i_13_487_126_0, i_13_487_132_0,
    i_13_487_273_0, i_13_487_282_0, i_13_487_283_0, i_13_487_284_0,
    i_13_487_335_0, i_13_487_357_0, i_13_487_360_0, i_13_487_361_0,
    i_13_487_472_0, i_13_487_519_0, i_13_487_538_0, i_13_487_689_0,
    i_13_487_838_0, i_13_487_866_0, i_13_487_867_0, i_13_487_869_0,
    i_13_487_1096_0, i_13_487_1111_0, i_13_487_1112_0, i_13_487_1114_0,
    i_13_487_1119_0, i_13_487_1132_0, i_13_487_1243_0, i_13_487_1329_0,
    i_13_487_1430_0, i_13_487_1501_0, i_13_487_1549_0, i_13_487_1745_0,
    i_13_487_1770_0, i_13_487_1792_0, i_13_487_1795_0, i_13_487_1834_0,
    i_13_487_1858_0, i_13_487_1884_0, i_13_487_1896_0, i_13_487_2004_0,
    i_13_487_2008_0, i_13_487_2010_0, i_13_487_2017_0, i_13_487_2097_0,
    i_13_487_2113_0, i_13_487_2145_0, i_13_487_2148_0, i_13_487_2223_0,
    i_13_487_2260_0, i_13_487_2384_0, i_13_487_2461_0, i_13_487_2514_0,
    i_13_487_2537_0, i_13_487_2733_0, i_13_487_2798_0, i_13_487_2883_0,
    i_13_487_2890_0, i_13_487_3048_0, i_13_487_3057_0, i_13_487_3059_0,
    i_13_487_3076_0, i_13_487_3077_0, i_13_487_3097_0, i_13_487_3145_0,
    i_13_487_3219_0, i_13_487_3266_0, i_13_487_3286_0, i_13_487_3315_0,
    i_13_487_3348_0, i_13_487_3489_0, i_13_487_3490_0, i_13_487_3549_0,
    i_13_487_3550_0, i_13_487_3604_0, i_13_487_3671_0, i_13_487_3730_0,
    i_13_487_3735_0, i_13_487_3748_0, i_13_487_3822_0, i_13_487_3869_0,
    i_13_487_3881_0, i_13_487_3909_0, i_13_487_3910_0, i_13_487_3952_0,
    i_13_487_4018_0, i_13_487_4125_0, i_13_487_4126_0, i_13_487_4165_0,
    i_13_487_4261_0, i_13_487_4272_0, i_13_487_4330_0, i_13_487_4333_0,
    i_13_487_4362_0, i_13_487_4433_0, i_13_487_4454_0, i_13_487_4467_0,
    i_13_487_4471_0, i_13_487_4516_0, i_13_487_4565_0, i_13_487_4578_0;
  output o_13_487_0_0;
  assign o_13_487_0_0 = ~((~i_13_487_4272_0 & ((~i_13_487_3315_0 & ~i_13_487_3490_0) | (~i_13_487_4333_0 & ~i_13_487_4433_0))) | (~i_13_487_4362_0 & (i_13_487_283_0 | (~i_13_487_472_0 & ~i_13_487_2113_0 & ~i_13_487_4516_0))) | (~i_13_487_3489_0 & ~i_13_487_3550_0 & ~i_13_487_4165_0) | (~i_13_487_2537_0 & ~i_13_487_3822_0 & ~i_13_487_4333_0 & ~i_13_487_4516_0));
endmodule



// Benchmark "kernel_13_488" written by ABC on Sun Jul 19 10:52:08 2020

module kernel_13_488 ( 
    i_13_488_45_0, i_13_488_46_0, i_13_488_100_0, i_13_488_127_0,
    i_13_488_154_0, i_13_488_193_0, i_13_488_252_0, i_13_488_270_0,
    i_13_488_271_0, i_13_488_374_0, i_13_488_378_0, i_13_488_379_0,
    i_13_488_425_0, i_13_488_428_0, i_13_488_451_0, i_13_488_523_0,
    i_13_488_569_0, i_13_488_570_0, i_13_488_688_0, i_13_488_817_0,
    i_13_488_927_0, i_13_488_949_0, i_13_488_1063_0, i_13_488_1087_0,
    i_13_488_1147_0, i_13_488_1219_0, i_13_488_1271_0, i_13_488_1345_0,
    i_13_488_1379_0, i_13_488_1435_0, i_13_488_1458_0, i_13_488_1496_0,
    i_13_488_1539_0, i_13_488_1566_0, i_13_488_1567_0, i_13_488_1733_0,
    i_13_488_1749_0, i_13_488_1800_0, i_13_488_1801_0, i_13_488_1802_0,
    i_13_488_1810_0, i_13_488_1848_0, i_13_488_1891_0, i_13_488_2026_0,
    i_13_488_2107_0, i_13_488_2108_0, i_13_488_2146_0, i_13_488_2197_0,
    i_13_488_2233_0, i_13_488_2260_0, i_13_488_2435_0, i_13_488_2525_0,
    i_13_488_2576_0, i_13_488_2614_0, i_13_488_2618_0, i_13_488_2713_0,
    i_13_488_2740_0, i_13_488_2745_0, i_13_488_2747_0, i_13_488_2763_0,
    i_13_488_2917_0, i_13_488_2935_0, i_13_488_2987_0, i_13_488_3008_0,
    i_13_488_3016_0, i_13_488_3056_0, i_13_488_3214_0, i_13_488_3215_0,
    i_13_488_3367_0, i_13_488_3376_0, i_13_488_3377_0, i_13_488_3528_0,
    i_13_488_3547_0, i_13_488_3591_0, i_13_488_3722_0, i_13_488_3742_0,
    i_13_488_3763_0, i_13_488_3769_0, i_13_488_3770_0, i_13_488_3817_0,
    i_13_488_3821_0, i_13_488_3905_0, i_13_488_3978_0, i_13_488_4042_0,
    i_13_488_4064_0, i_13_488_4086_0, i_13_488_4087_0, i_13_488_4234_0,
    i_13_488_4250_0, i_13_488_4258_0, i_13_488_4266_0, i_13_488_4267_0,
    i_13_488_4268_0, i_13_488_4312_0, i_13_488_4322_0, i_13_488_4358_0,
    i_13_488_4385_0, i_13_488_4447_0, i_13_488_4562_0, i_13_488_4564_0,
    o_13_488_0_0  );
  input  i_13_488_45_0, i_13_488_46_0, i_13_488_100_0, i_13_488_127_0,
    i_13_488_154_0, i_13_488_193_0, i_13_488_252_0, i_13_488_270_0,
    i_13_488_271_0, i_13_488_374_0, i_13_488_378_0, i_13_488_379_0,
    i_13_488_425_0, i_13_488_428_0, i_13_488_451_0, i_13_488_523_0,
    i_13_488_569_0, i_13_488_570_0, i_13_488_688_0, i_13_488_817_0,
    i_13_488_927_0, i_13_488_949_0, i_13_488_1063_0, i_13_488_1087_0,
    i_13_488_1147_0, i_13_488_1219_0, i_13_488_1271_0, i_13_488_1345_0,
    i_13_488_1379_0, i_13_488_1435_0, i_13_488_1458_0, i_13_488_1496_0,
    i_13_488_1539_0, i_13_488_1566_0, i_13_488_1567_0, i_13_488_1733_0,
    i_13_488_1749_0, i_13_488_1800_0, i_13_488_1801_0, i_13_488_1802_0,
    i_13_488_1810_0, i_13_488_1848_0, i_13_488_1891_0, i_13_488_2026_0,
    i_13_488_2107_0, i_13_488_2108_0, i_13_488_2146_0, i_13_488_2197_0,
    i_13_488_2233_0, i_13_488_2260_0, i_13_488_2435_0, i_13_488_2525_0,
    i_13_488_2576_0, i_13_488_2614_0, i_13_488_2618_0, i_13_488_2713_0,
    i_13_488_2740_0, i_13_488_2745_0, i_13_488_2747_0, i_13_488_2763_0,
    i_13_488_2917_0, i_13_488_2935_0, i_13_488_2987_0, i_13_488_3008_0,
    i_13_488_3016_0, i_13_488_3056_0, i_13_488_3214_0, i_13_488_3215_0,
    i_13_488_3367_0, i_13_488_3376_0, i_13_488_3377_0, i_13_488_3528_0,
    i_13_488_3547_0, i_13_488_3591_0, i_13_488_3722_0, i_13_488_3742_0,
    i_13_488_3763_0, i_13_488_3769_0, i_13_488_3770_0, i_13_488_3817_0,
    i_13_488_3821_0, i_13_488_3905_0, i_13_488_3978_0, i_13_488_4042_0,
    i_13_488_4064_0, i_13_488_4086_0, i_13_488_4087_0, i_13_488_4234_0,
    i_13_488_4250_0, i_13_488_4258_0, i_13_488_4266_0, i_13_488_4267_0,
    i_13_488_4268_0, i_13_488_4312_0, i_13_488_4322_0, i_13_488_4358_0,
    i_13_488_4385_0, i_13_488_4447_0, i_13_488_4562_0, i_13_488_4564_0;
  output o_13_488_0_0;
  assign o_13_488_0_0 = ~((~i_13_488_4087_0 & ~i_13_488_4564_0) | (~i_13_488_1800_0 & ~i_13_488_2108_0) | (~i_13_488_1733_0 & ~i_13_488_3591_0 & ~i_13_488_4267_0 & ~i_13_488_4312_0));
endmodule



// Benchmark "kernel_13_489" written by ABC on Sun Jul 19 10:52:09 2020

module kernel_13_489 ( 
    i_13_489_73_0, i_13_489_108_0, i_13_489_111_0, i_13_489_112_0,
    i_13_489_136_0, i_13_489_261_0, i_13_489_363_0, i_13_489_387_0,
    i_13_489_442_0, i_13_489_581_0, i_13_489_603_0, i_13_489_604_0,
    i_13_489_666_0, i_13_489_669_0, i_13_489_810_0, i_13_489_813_0,
    i_13_489_814_0, i_13_489_855_0, i_13_489_856_0, i_13_489_1017_0,
    i_13_489_1081_0, i_13_489_1144_0, i_13_489_1211_0, i_13_489_1215_0,
    i_13_489_1216_0, i_13_489_1422_0, i_13_489_1423_0, i_13_489_1426_0,
    i_13_489_1454_0, i_13_489_1485_0, i_13_489_1486_0, i_13_489_1494_0,
    i_13_489_1566_0, i_13_489_1597_0, i_13_489_1620_0, i_13_489_1622_0,
    i_13_489_1629_0, i_13_489_1719_0, i_13_489_1774_0, i_13_489_1794_0,
    i_13_489_1812_0, i_13_489_1836_0, i_13_489_1837_0, i_13_489_1840_0,
    i_13_489_1849_0, i_13_489_1938_0, i_13_489_1989_0, i_13_489_2011_0,
    i_13_489_2137_0, i_13_489_2169_0, i_13_489_2404_0, i_13_489_2407_0,
    i_13_489_2434_0, i_13_489_2448_0, i_13_489_2451_0, i_13_489_2452_0,
    i_13_489_2497_0, i_13_489_2538_0, i_13_489_2610_0, i_13_489_2858_0,
    i_13_489_2907_0, i_13_489_2916_0, i_13_489_2917_0, i_13_489_2935_0,
    i_13_489_2938_0, i_13_489_3000_0, i_13_489_3100_0, i_13_489_3144_0,
    i_13_489_3213_0, i_13_489_3288_0, i_13_489_3315_0, i_13_489_3340_0,
    i_13_489_3384_0, i_13_489_3385_0, i_13_489_3393_0, i_13_489_3474_0,
    i_13_489_3475_0, i_13_489_3501_0, i_13_489_3502_0, i_13_489_3528_0,
    i_13_489_3529_0, i_13_489_3702_0, i_13_489_3738_0, i_13_489_3739_0,
    i_13_489_3888_0, i_13_489_3891_0, i_13_489_4055_0, i_13_489_4060_0,
    i_13_489_4063_0, i_13_489_4159_0, i_13_489_4204_0, i_13_489_4248_0,
    i_13_489_4251_0, i_13_489_4315_0, i_13_489_4338_0, i_13_489_4342_0,
    i_13_489_4365_0, i_13_489_4366_0, i_13_489_4368_0, i_13_489_4540_0,
    o_13_489_0_0  );
  input  i_13_489_73_0, i_13_489_108_0, i_13_489_111_0, i_13_489_112_0,
    i_13_489_136_0, i_13_489_261_0, i_13_489_363_0, i_13_489_387_0,
    i_13_489_442_0, i_13_489_581_0, i_13_489_603_0, i_13_489_604_0,
    i_13_489_666_0, i_13_489_669_0, i_13_489_810_0, i_13_489_813_0,
    i_13_489_814_0, i_13_489_855_0, i_13_489_856_0, i_13_489_1017_0,
    i_13_489_1081_0, i_13_489_1144_0, i_13_489_1211_0, i_13_489_1215_0,
    i_13_489_1216_0, i_13_489_1422_0, i_13_489_1423_0, i_13_489_1426_0,
    i_13_489_1454_0, i_13_489_1485_0, i_13_489_1486_0, i_13_489_1494_0,
    i_13_489_1566_0, i_13_489_1597_0, i_13_489_1620_0, i_13_489_1622_0,
    i_13_489_1629_0, i_13_489_1719_0, i_13_489_1774_0, i_13_489_1794_0,
    i_13_489_1812_0, i_13_489_1836_0, i_13_489_1837_0, i_13_489_1840_0,
    i_13_489_1849_0, i_13_489_1938_0, i_13_489_1989_0, i_13_489_2011_0,
    i_13_489_2137_0, i_13_489_2169_0, i_13_489_2404_0, i_13_489_2407_0,
    i_13_489_2434_0, i_13_489_2448_0, i_13_489_2451_0, i_13_489_2452_0,
    i_13_489_2497_0, i_13_489_2538_0, i_13_489_2610_0, i_13_489_2858_0,
    i_13_489_2907_0, i_13_489_2916_0, i_13_489_2917_0, i_13_489_2935_0,
    i_13_489_2938_0, i_13_489_3000_0, i_13_489_3100_0, i_13_489_3144_0,
    i_13_489_3213_0, i_13_489_3288_0, i_13_489_3315_0, i_13_489_3340_0,
    i_13_489_3384_0, i_13_489_3385_0, i_13_489_3393_0, i_13_489_3474_0,
    i_13_489_3475_0, i_13_489_3501_0, i_13_489_3502_0, i_13_489_3528_0,
    i_13_489_3529_0, i_13_489_3702_0, i_13_489_3738_0, i_13_489_3739_0,
    i_13_489_3888_0, i_13_489_3891_0, i_13_489_4055_0, i_13_489_4060_0,
    i_13_489_4063_0, i_13_489_4159_0, i_13_489_4204_0, i_13_489_4248_0,
    i_13_489_4251_0, i_13_489_4315_0, i_13_489_4338_0, i_13_489_4342_0,
    i_13_489_4365_0, i_13_489_4366_0, i_13_489_4368_0, i_13_489_4540_0;
  output o_13_489_0_0;
  assign o_13_489_0_0 = ~((~i_13_489_1485_0 & (i_13_489_2404_0 | (~i_13_489_1794_0 & ~i_13_489_3144_0))) | (~i_13_489_111_0 & i_13_489_3393_0) | (~i_13_489_3393_0 & ~i_13_489_3501_0) | (~i_13_489_1017_0 & ~i_13_489_2917_0 & ~i_13_489_4159_0));
endmodule



// Benchmark "kernel_13_490" written by ABC on Sun Jul 19 10:52:09 2020

module kernel_13_490 ( 
    i_13_490_19_0, i_13_490_31_0, i_13_490_99_0, i_13_490_112_0,
    i_13_490_162_0, i_13_490_165_0, i_13_490_166_0, i_13_490_180_0,
    i_13_490_183_0, i_13_490_184_0, i_13_490_185_0, i_13_490_216_0,
    i_13_490_217_0, i_13_490_256_0, i_13_490_393_0, i_13_490_639_0,
    i_13_490_796_0, i_13_490_837_0, i_13_490_1063_0, i_13_490_1078_0,
    i_13_490_1116_0, i_13_490_1118_0, i_13_490_1121_0, i_13_490_1146_0,
    i_13_490_1219_0, i_13_490_1231_0, i_13_490_1263_0, i_13_490_1323_0,
    i_13_490_1326_0, i_13_490_1426_0, i_13_490_1458_0, i_13_490_1480_0,
    i_13_490_1513_0, i_13_490_1521_0, i_13_490_1525_0, i_13_490_1677_0,
    i_13_490_1746_0, i_13_490_1764_0, i_13_490_1784_0, i_13_490_1804_0,
    i_13_490_1831_0, i_13_490_1840_0, i_13_490_1857_0, i_13_490_1909_0,
    i_13_490_1938_0, i_13_490_1940_0, i_13_490_1989_0, i_13_490_1999_0,
    i_13_490_2002_0, i_13_490_2043_0, i_13_490_2106_0, i_13_490_2107_0,
    i_13_490_2116_0, i_13_490_2145_0, i_13_490_2146_0, i_13_490_2185_0,
    i_13_490_2233_0, i_13_490_2260_0, i_13_490_2277_0, i_13_490_2340_0,
    i_13_490_2395_0, i_13_490_2466_0, i_13_490_2476_0, i_13_490_2564_0,
    i_13_490_2748_0, i_13_490_2761_0, i_13_490_2937_0, i_13_490_2979_0,
    i_13_490_2980_0, i_13_490_2997_0, i_13_490_3024_0, i_13_490_3026_0,
    i_13_490_3027_0, i_13_490_3108_0, i_13_490_3111_0, i_13_490_3115_0,
    i_13_490_3144_0, i_13_490_3145_0, i_13_490_3196_0, i_13_490_3208_0,
    i_13_490_3286_0, i_13_490_3289_0, i_13_490_3471_0, i_13_490_3558_0,
    i_13_490_3650_0, i_13_490_3730_0, i_13_490_3763_0, i_13_490_3892_0,
    i_13_490_4042_0, i_13_490_4077_0, i_13_490_4187_0, i_13_490_4203_0,
    i_13_490_4204_0, i_13_490_4268_0, i_13_490_4314_0, i_13_490_4396_0,
    i_13_490_4501_0, i_13_490_4558_0, i_13_490_4564_0, i_13_490_4600_0,
    o_13_490_0_0  );
  input  i_13_490_19_0, i_13_490_31_0, i_13_490_99_0, i_13_490_112_0,
    i_13_490_162_0, i_13_490_165_0, i_13_490_166_0, i_13_490_180_0,
    i_13_490_183_0, i_13_490_184_0, i_13_490_185_0, i_13_490_216_0,
    i_13_490_217_0, i_13_490_256_0, i_13_490_393_0, i_13_490_639_0,
    i_13_490_796_0, i_13_490_837_0, i_13_490_1063_0, i_13_490_1078_0,
    i_13_490_1116_0, i_13_490_1118_0, i_13_490_1121_0, i_13_490_1146_0,
    i_13_490_1219_0, i_13_490_1231_0, i_13_490_1263_0, i_13_490_1323_0,
    i_13_490_1326_0, i_13_490_1426_0, i_13_490_1458_0, i_13_490_1480_0,
    i_13_490_1513_0, i_13_490_1521_0, i_13_490_1525_0, i_13_490_1677_0,
    i_13_490_1746_0, i_13_490_1764_0, i_13_490_1784_0, i_13_490_1804_0,
    i_13_490_1831_0, i_13_490_1840_0, i_13_490_1857_0, i_13_490_1909_0,
    i_13_490_1938_0, i_13_490_1940_0, i_13_490_1989_0, i_13_490_1999_0,
    i_13_490_2002_0, i_13_490_2043_0, i_13_490_2106_0, i_13_490_2107_0,
    i_13_490_2116_0, i_13_490_2145_0, i_13_490_2146_0, i_13_490_2185_0,
    i_13_490_2233_0, i_13_490_2260_0, i_13_490_2277_0, i_13_490_2340_0,
    i_13_490_2395_0, i_13_490_2466_0, i_13_490_2476_0, i_13_490_2564_0,
    i_13_490_2748_0, i_13_490_2761_0, i_13_490_2937_0, i_13_490_2979_0,
    i_13_490_2980_0, i_13_490_2997_0, i_13_490_3024_0, i_13_490_3026_0,
    i_13_490_3027_0, i_13_490_3108_0, i_13_490_3111_0, i_13_490_3115_0,
    i_13_490_3144_0, i_13_490_3145_0, i_13_490_3196_0, i_13_490_3208_0,
    i_13_490_3286_0, i_13_490_3289_0, i_13_490_3471_0, i_13_490_3558_0,
    i_13_490_3650_0, i_13_490_3730_0, i_13_490_3763_0, i_13_490_3892_0,
    i_13_490_4042_0, i_13_490_4077_0, i_13_490_4187_0, i_13_490_4203_0,
    i_13_490_4204_0, i_13_490_4268_0, i_13_490_4314_0, i_13_490_4396_0,
    i_13_490_4501_0, i_13_490_4558_0, i_13_490_4564_0, i_13_490_4600_0;
  output o_13_490_0_0;
  assign o_13_490_0_0 = ~((~i_13_490_1525_0 & ((i_13_490_1146_0 & i_13_490_3111_0) | (i_13_490_31_0 & i_13_490_1840_0 & ~i_13_490_4077_0 & ~i_13_490_4314_0))) | (~i_13_490_4314_0 & ((~i_13_490_183_0 & ~i_13_490_2980_0) | (~i_13_490_1326_0 & i_13_490_4558_0))) | (~i_13_490_1118_0 & ~i_13_490_1677_0 & ~i_13_490_2277_0) | (~i_13_490_1480_0 & i_13_490_2761_0) | (~i_13_490_185_0 & ~i_13_490_1146_0 & ~i_13_490_1840_0 & ~i_13_490_2107_0 & ~i_13_490_2185_0 & ~i_13_490_4077_0) | (~i_13_490_1831_0 & i_13_490_4187_0) | (i_13_490_3144_0 & ~i_13_490_4564_0));
endmodule



// Benchmark "kernel_13_491" written by ABC on Sun Jul 19 10:52:10 2020

module kernel_13_491 ( 
    i_13_491_27_0, i_13_491_64_0, i_13_491_104_0, i_13_491_131_0,
    i_13_491_157_0, i_13_491_174_0, i_13_491_208_0, i_13_491_209_0,
    i_13_491_218_0, i_13_491_225_0, i_13_491_266_0, i_13_491_307_0,
    i_13_491_355_0, i_13_491_356_0, i_13_491_441_0, i_13_491_463_0,
    i_13_491_464_0, i_13_491_526_0, i_13_491_531_0, i_13_491_549_0,
    i_13_491_613_0, i_13_491_639_0, i_13_491_666_0, i_13_491_667_0,
    i_13_491_742_0, i_13_491_812_0, i_13_491_839_0, i_13_491_841_0,
    i_13_491_961_0, i_13_491_1019_0, i_13_491_1073_0, i_13_491_1129_0,
    i_13_491_1301_0, i_13_491_1307_0, i_13_491_1444_0, i_13_491_1535_0,
    i_13_491_1594_0, i_13_491_1595_0, i_13_491_1604_0, i_13_491_1624_0,
    i_13_491_1632_0, i_13_491_1639_0, i_13_491_1697_0, i_13_491_1723_0,
    i_13_491_1774_0, i_13_491_1846_0, i_13_491_1847_0, i_13_491_1909_0,
    i_13_491_2030_0, i_13_491_2091_0, i_13_491_2101_0, i_13_491_2143_0,
    i_13_491_2199_0, i_13_491_2200_0, i_13_491_2237_0, i_13_491_2263_0,
    i_13_491_2297_0, i_13_491_2444_0, i_13_491_2504_0, i_13_491_2507_0,
    i_13_491_2512_0, i_13_491_2551_0, i_13_491_2673_0, i_13_491_2691_0,
    i_13_491_2822_0, i_13_491_2885_0, i_13_491_2936_0, i_13_491_3070_0,
    i_13_491_3089_0, i_13_491_3143_0, i_13_491_3241_0, i_13_491_3242_0,
    i_13_491_3343_0, i_13_491_3389_0, i_13_491_3460_0, i_13_491_3469_0,
    i_13_491_3472_0, i_13_491_3530_0, i_13_491_3595_0, i_13_491_3599_0,
    i_13_491_3619_0, i_13_491_3631_0, i_13_491_3637_0, i_13_491_3667_0,
    i_13_491_3682_0, i_13_491_3719_0, i_13_491_3728_0, i_13_491_3793_0,
    i_13_491_3857_0, i_13_491_3924_0, i_13_491_3935_0, i_13_491_3989_0,
    i_13_491_4060_0, i_13_491_4061_0, i_13_491_4077_0, i_13_491_4122_0,
    i_13_491_4313_0, i_13_491_4342_0, i_13_491_4345_0, i_13_491_4379_0,
    o_13_491_0_0  );
  input  i_13_491_27_0, i_13_491_64_0, i_13_491_104_0, i_13_491_131_0,
    i_13_491_157_0, i_13_491_174_0, i_13_491_208_0, i_13_491_209_0,
    i_13_491_218_0, i_13_491_225_0, i_13_491_266_0, i_13_491_307_0,
    i_13_491_355_0, i_13_491_356_0, i_13_491_441_0, i_13_491_463_0,
    i_13_491_464_0, i_13_491_526_0, i_13_491_531_0, i_13_491_549_0,
    i_13_491_613_0, i_13_491_639_0, i_13_491_666_0, i_13_491_667_0,
    i_13_491_742_0, i_13_491_812_0, i_13_491_839_0, i_13_491_841_0,
    i_13_491_961_0, i_13_491_1019_0, i_13_491_1073_0, i_13_491_1129_0,
    i_13_491_1301_0, i_13_491_1307_0, i_13_491_1444_0, i_13_491_1535_0,
    i_13_491_1594_0, i_13_491_1595_0, i_13_491_1604_0, i_13_491_1624_0,
    i_13_491_1632_0, i_13_491_1639_0, i_13_491_1697_0, i_13_491_1723_0,
    i_13_491_1774_0, i_13_491_1846_0, i_13_491_1847_0, i_13_491_1909_0,
    i_13_491_2030_0, i_13_491_2091_0, i_13_491_2101_0, i_13_491_2143_0,
    i_13_491_2199_0, i_13_491_2200_0, i_13_491_2237_0, i_13_491_2263_0,
    i_13_491_2297_0, i_13_491_2444_0, i_13_491_2504_0, i_13_491_2507_0,
    i_13_491_2512_0, i_13_491_2551_0, i_13_491_2673_0, i_13_491_2691_0,
    i_13_491_2822_0, i_13_491_2885_0, i_13_491_2936_0, i_13_491_3070_0,
    i_13_491_3089_0, i_13_491_3143_0, i_13_491_3241_0, i_13_491_3242_0,
    i_13_491_3343_0, i_13_491_3389_0, i_13_491_3460_0, i_13_491_3469_0,
    i_13_491_3472_0, i_13_491_3530_0, i_13_491_3595_0, i_13_491_3599_0,
    i_13_491_3619_0, i_13_491_3631_0, i_13_491_3637_0, i_13_491_3667_0,
    i_13_491_3682_0, i_13_491_3719_0, i_13_491_3728_0, i_13_491_3793_0,
    i_13_491_3857_0, i_13_491_3924_0, i_13_491_3935_0, i_13_491_3989_0,
    i_13_491_4060_0, i_13_491_4061_0, i_13_491_4077_0, i_13_491_4122_0,
    i_13_491_4313_0, i_13_491_4342_0, i_13_491_4345_0, i_13_491_4379_0;
  output o_13_491_0_0;
  assign o_13_491_0_0 = ~(~i_13_491_3619_0 | (~i_13_491_463_0 & ~i_13_491_4313_0) | (i_13_491_441_0 & ~i_13_491_2551_0 & ~i_13_491_3682_0));
endmodule



// Benchmark "kernel_13_492" written by ABC on Sun Jul 19 10:52:11 2020

module kernel_13_492 ( 
    i_13_492_44_0, i_13_492_45_0, i_13_492_46_0, i_13_492_55_0,
    i_13_492_84_0, i_13_492_94_0, i_13_492_112_0, i_13_492_134_0,
    i_13_492_207_0, i_13_492_234_0, i_13_492_243_0, i_13_492_244_0,
    i_13_492_283_0, i_13_492_323_0, i_13_492_521_0, i_13_492_598_0,
    i_13_492_614_0, i_13_492_623_0, i_13_492_693_0, i_13_492_694_0,
    i_13_492_702_0, i_13_492_760_0, i_13_492_838_0, i_13_492_955_0,
    i_13_492_1071_0, i_13_492_1116_0, i_13_492_1119_0, i_13_492_1128_0,
    i_13_492_1129_0, i_13_492_1152_0, i_13_492_1219_0, i_13_492_1243_0,
    i_13_492_1317_0, i_13_492_1360_0, i_13_492_1405_0, i_13_492_1521_0,
    i_13_492_1533_0, i_13_492_1535_0, i_13_492_1647_0, i_13_492_1678_0,
    i_13_492_1777_0, i_13_492_1795_0, i_13_492_1804_0, i_13_492_1840_0,
    i_13_492_1929_0, i_13_492_1957_0, i_13_492_2002_0, i_13_492_2142_0,
    i_13_492_2208_0, i_13_492_2254_0, i_13_492_2460_0, i_13_492_2511_0,
    i_13_492_2512_0, i_13_492_2541_0, i_13_492_2578_0, i_13_492_2646_0,
    i_13_492_2666_0, i_13_492_2692_0, i_13_492_2845_0, i_13_492_2880_0,
    i_13_492_2910_0, i_13_492_3000_0, i_13_492_3002_0, i_13_492_3025_0,
    i_13_492_3113_0, i_13_492_3127_0, i_13_492_3367_0, i_13_492_3371_0,
    i_13_492_3420_0, i_13_492_3474_0, i_13_492_3475_0, i_13_492_3519_0,
    i_13_492_3528_0, i_13_492_3546_0, i_13_492_3636_0, i_13_492_3641_0,
    i_13_492_3753_0, i_13_492_3757_0, i_13_492_3819_0, i_13_492_3887_0,
    i_13_492_3898_0, i_13_492_3923_0, i_13_492_3987_0, i_13_492_4035_0,
    i_13_492_4036_0, i_13_492_4041_0, i_13_492_4167_0, i_13_492_4311_0,
    i_13_492_4329_0, i_13_492_4351_0, i_13_492_4377_0, i_13_492_4378_0,
    i_13_492_4414_0, i_13_492_4430_0, i_13_492_4450_0, i_13_492_4509_0,
    i_13_492_4510_0, i_13_492_4567_0, i_13_492_4593_0, i_13_492_4603_0,
    o_13_492_0_0  );
  input  i_13_492_44_0, i_13_492_45_0, i_13_492_46_0, i_13_492_55_0,
    i_13_492_84_0, i_13_492_94_0, i_13_492_112_0, i_13_492_134_0,
    i_13_492_207_0, i_13_492_234_0, i_13_492_243_0, i_13_492_244_0,
    i_13_492_283_0, i_13_492_323_0, i_13_492_521_0, i_13_492_598_0,
    i_13_492_614_0, i_13_492_623_0, i_13_492_693_0, i_13_492_694_0,
    i_13_492_702_0, i_13_492_760_0, i_13_492_838_0, i_13_492_955_0,
    i_13_492_1071_0, i_13_492_1116_0, i_13_492_1119_0, i_13_492_1128_0,
    i_13_492_1129_0, i_13_492_1152_0, i_13_492_1219_0, i_13_492_1243_0,
    i_13_492_1317_0, i_13_492_1360_0, i_13_492_1405_0, i_13_492_1521_0,
    i_13_492_1533_0, i_13_492_1535_0, i_13_492_1647_0, i_13_492_1678_0,
    i_13_492_1777_0, i_13_492_1795_0, i_13_492_1804_0, i_13_492_1840_0,
    i_13_492_1929_0, i_13_492_1957_0, i_13_492_2002_0, i_13_492_2142_0,
    i_13_492_2208_0, i_13_492_2254_0, i_13_492_2460_0, i_13_492_2511_0,
    i_13_492_2512_0, i_13_492_2541_0, i_13_492_2578_0, i_13_492_2646_0,
    i_13_492_2666_0, i_13_492_2692_0, i_13_492_2845_0, i_13_492_2880_0,
    i_13_492_2910_0, i_13_492_3000_0, i_13_492_3002_0, i_13_492_3025_0,
    i_13_492_3113_0, i_13_492_3127_0, i_13_492_3367_0, i_13_492_3371_0,
    i_13_492_3420_0, i_13_492_3474_0, i_13_492_3475_0, i_13_492_3519_0,
    i_13_492_3528_0, i_13_492_3546_0, i_13_492_3636_0, i_13_492_3641_0,
    i_13_492_3753_0, i_13_492_3757_0, i_13_492_3819_0, i_13_492_3887_0,
    i_13_492_3898_0, i_13_492_3923_0, i_13_492_3987_0, i_13_492_4035_0,
    i_13_492_4036_0, i_13_492_4041_0, i_13_492_4167_0, i_13_492_4311_0,
    i_13_492_4329_0, i_13_492_4351_0, i_13_492_4377_0, i_13_492_4378_0,
    i_13_492_4414_0, i_13_492_4430_0, i_13_492_4450_0, i_13_492_4509_0,
    i_13_492_4510_0, i_13_492_4567_0, i_13_492_4593_0, i_13_492_4603_0;
  output o_13_492_0_0;
  assign o_13_492_0_0 = ~(~i_13_492_4036_0 | (~i_13_492_1521_0 & (~i_13_492_234_0 | ~i_13_492_2880_0)));
endmodule



// Benchmark "kernel_13_493" written by ABC on Sun Jul 19 10:52:12 2020

module kernel_13_493 ( 
    i_13_493_30_0, i_13_493_38_0, i_13_493_158_0, i_13_493_161_0,
    i_13_493_172_0, i_13_493_173_0, i_13_493_175_0, i_13_493_190_0,
    i_13_493_247_0, i_13_493_280_0, i_13_493_281_0, i_13_493_283_0,
    i_13_493_284_0, i_13_493_316_0, i_13_493_334_0, i_13_493_488_0,
    i_13_493_525_0, i_13_493_527_0, i_13_493_577_0, i_13_493_640_0,
    i_13_493_685_0, i_13_493_688_0, i_13_493_689_0, i_13_493_797_0,
    i_13_493_820_0, i_13_493_821_0, i_13_493_822_0, i_13_493_847_0,
    i_13_493_1067_0, i_13_493_1120_0, i_13_493_1216_0, i_13_493_1219_0,
    i_13_493_1225_0, i_13_493_1306_0, i_13_493_1309_0, i_13_493_1504_0,
    i_13_493_1540_0, i_13_493_1594_0, i_13_493_1601_0, i_13_493_1730_0,
    i_13_493_1768_0, i_13_493_1813_0, i_13_493_1882_0, i_13_493_1926_0,
    i_13_493_2054_0, i_13_493_2092_0, i_13_493_2173_0, i_13_493_2188_0,
    i_13_493_2189_0, i_13_493_2236_0, i_13_493_2422_0, i_13_493_2425_0,
    i_13_493_2443_0, i_13_493_2475_0, i_13_493_2622_0, i_13_493_2674_0,
    i_13_493_2677_0, i_13_493_2702_0, i_13_493_3007_0, i_13_493_3069_0,
    i_13_493_3142_0, i_13_493_3214_0, i_13_493_3217_0, i_13_493_3250_0,
    i_13_493_3267_0, i_13_493_3268_0, i_13_493_3271_0, i_13_493_3272_0,
    i_13_493_3378_0, i_13_493_3386_0, i_13_493_3389_0, i_13_493_3421_0,
    i_13_493_3424_0, i_13_493_3451_0, i_13_493_3457_0, i_13_493_3722_0,
    i_13_493_3726_0, i_13_493_3730_0, i_13_493_3906_0, i_13_493_3910_0,
    i_13_493_3917_0, i_13_493_3982_0, i_13_493_3991_0, i_13_493_4014_0,
    i_13_493_4015_0, i_13_493_4016_0, i_13_493_4018_0, i_13_493_4062_0,
    i_13_493_4081_0, i_13_493_4180_0, i_13_493_4214_0, i_13_493_4249_0,
    i_13_493_4257_0, i_13_493_4261_0, i_13_493_4306_0, i_13_493_4374_0,
    i_13_493_4396_0, i_13_493_4424_0, i_13_493_4450_0, i_13_493_4544_0,
    o_13_493_0_0  );
  input  i_13_493_30_0, i_13_493_38_0, i_13_493_158_0, i_13_493_161_0,
    i_13_493_172_0, i_13_493_173_0, i_13_493_175_0, i_13_493_190_0,
    i_13_493_247_0, i_13_493_280_0, i_13_493_281_0, i_13_493_283_0,
    i_13_493_284_0, i_13_493_316_0, i_13_493_334_0, i_13_493_488_0,
    i_13_493_525_0, i_13_493_527_0, i_13_493_577_0, i_13_493_640_0,
    i_13_493_685_0, i_13_493_688_0, i_13_493_689_0, i_13_493_797_0,
    i_13_493_820_0, i_13_493_821_0, i_13_493_822_0, i_13_493_847_0,
    i_13_493_1067_0, i_13_493_1120_0, i_13_493_1216_0, i_13_493_1219_0,
    i_13_493_1225_0, i_13_493_1306_0, i_13_493_1309_0, i_13_493_1504_0,
    i_13_493_1540_0, i_13_493_1594_0, i_13_493_1601_0, i_13_493_1730_0,
    i_13_493_1768_0, i_13_493_1813_0, i_13_493_1882_0, i_13_493_1926_0,
    i_13_493_2054_0, i_13_493_2092_0, i_13_493_2173_0, i_13_493_2188_0,
    i_13_493_2189_0, i_13_493_2236_0, i_13_493_2422_0, i_13_493_2425_0,
    i_13_493_2443_0, i_13_493_2475_0, i_13_493_2622_0, i_13_493_2674_0,
    i_13_493_2677_0, i_13_493_2702_0, i_13_493_3007_0, i_13_493_3069_0,
    i_13_493_3142_0, i_13_493_3214_0, i_13_493_3217_0, i_13_493_3250_0,
    i_13_493_3267_0, i_13_493_3268_0, i_13_493_3271_0, i_13_493_3272_0,
    i_13_493_3378_0, i_13_493_3386_0, i_13_493_3389_0, i_13_493_3421_0,
    i_13_493_3424_0, i_13_493_3451_0, i_13_493_3457_0, i_13_493_3722_0,
    i_13_493_3726_0, i_13_493_3730_0, i_13_493_3906_0, i_13_493_3910_0,
    i_13_493_3917_0, i_13_493_3982_0, i_13_493_3991_0, i_13_493_4014_0,
    i_13_493_4015_0, i_13_493_4016_0, i_13_493_4018_0, i_13_493_4062_0,
    i_13_493_4081_0, i_13_493_4180_0, i_13_493_4214_0, i_13_493_4249_0,
    i_13_493_4257_0, i_13_493_4261_0, i_13_493_4306_0, i_13_493_4374_0,
    i_13_493_4396_0, i_13_493_4424_0, i_13_493_4450_0, i_13_493_4544_0;
  output o_13_493_0_0;
  assign o_13_493_0_0 = 0;
endmodule



// Benchmark "kernel_13_494" written by ABC on Sun Jul 19 10:52:12 2020

module kernel_13_494 ( 
    i_13_494_25_0, i_13_494_31_0, i_13_494_40_0, i_13_494_74_0,
    i_13_494_139_0, i_13_494_186_0, i_13_494_229_0, i_13_494_317_0,
    i_13_494_454_0, i_13_494_510_0, i_13_494_573_0, i_13_494_589_0,
    i_13_494_659_0, i_13_494_661_0, i_13_494_663_0, i_13_494_733_0,
    i_13_494_854_0, i_13_494_938_0, i_13_494_940_0, i_13_494_1021_0,
    i_13_494_1075_0, i_13_494_1144_0, i_13_494_1145_0, i_13_494_1282_0,
    i_13_494_1284_0, i_13_494_1320_0, i_13_494_1424_0, i_13_494_1437_0,
    i_13_494_1660_0, i_13_494_1669_0, i_13_494_1714_0, i_13_494_1723_0,
    i_13_494_1773_0, i_13_494_1775_0, i_13_494_2188_0, i_13_494_2297_0,
    i_13_494_2425_0, i_13_494_2611_0, i_13_494_2659_0, i_13_494_2705_0,
    i_13_494_2742_0, i_13_494_2857_0, i_13_494_2958_0, i_13_494_3009_0,
    i_13_494_3010_0, i_13_494_3013_0, i_13_494_3046_0, i_13_494_3050_0,
    i_13_494_3072_0, i_13_494_3108_0, i_13_494_3109_0, i_13_494_3111_0,
    i_13_494_3156_0, i_13_494_3157_0, i_13_494_3205_0, i_13_494_3388_0,
    i_13_494_3408_0, i_13_494_3442_0, i_13_494_3460_0, i_13_494_3463_0,
    i_13_494_3468_0, i_13_494_3483_0, i_13_494_3484_0, i_13_494_3487_0,
    i_13_494_3489_0, i_13_494_3504_0, i_13_494_3550_0, i_13_494_3552_0,
    i_13_494_3565_0, i_13_494_3566_0, i_13_494_3568_0, i_13_494_3577_0,
    i_13_494_3603_0, i_13_494_3648_0, i_13_494_3681_0, i_13_494_3763_0,
    i_13_494_3764_0, i_13_494_3803_0, i_13_494_3819_0, i_13_494_3822_0,
    i_13_494_3862_0, i_13_494_3865_0, i_13_494_3980_0, i_13_494_4054_0,
    i_13_494_4163_0, i_13_494_4251_0, i_13_494_4312_0, i_13_494_4325_0,
    i_13_494_4340_0, i_13_494_4366_0, i_13_494_4367_0, i_13_494_4369_0,
    i_13_494_4370_0, i_13_494_4372_0, i_13_494_4396_0, i_13_494_4479_0,
    i_13_494_4558_0, i_13_494_4560_0, i_13_494_4568_0, i_13_494_4600_0,
    o_13_494_0_0  );
  input  i_13_494_25_0, i_13_494_31_0, i_13_494_40_0, i_13_494_74_0,
    i_13_494_139_0, i_13_494_186_0, i_13_494_229_0, i_13_494_317_0,
    i_13_494_454_0, i_13_494_510_0, i_13_494_573_0, i_13_494_589_0,
    i_13_494_659_0, i_13_494_661_0, i_13_494_663_0, i_13_494_733_0,
    i_13_494_854_0, i_13_494_938_0, i_13_494_940_0, i_13_494_1021_0,
    i_13_494_1075_0, i_13_494_1144_0, i_13_494_1145_0, i_13_494_1282_0,
    i_13_494_1284_0, i_13_494_1320_0, i_13_494_1424_0, i_13_494_1437_0,
    i_13_494_1660_0, i_13_494_1669_0, i_13_494_1714_0, i_13_494_1723_0,
    i_13_494_1773_0, i_13_494_1775_0, i_13_494_2188_0, i_13_494_2297_0,
    i_13_494_2425_0, i_13_494_2611_0, i_13_494_2659_0, i_13_494_2705_0,
    i_13_494_2742_0, i_13_494_2857_0, i_13_494_2958_0, i_13_494_3009_0,
    i_13_494_3010_0, i_13_494_3013_0, i_13_494_3046_0, i_13_494_3050_0,
    i_13_494_3072_0, i_13_494_3108_0, i_13_494_3109_0, i_13_494_3111_0,
    i_13_494_3156_0, i_13_494_3157_0, i_13_494_3205_0, i_13_494_3388_0,
    i_13_494_3408_0, i_13_494_3442_0, i_13_494_3460_0, i_13_494_3463_0,
    i_13_494_3468_0, i_13_494_3483_0, i_13_494_3484_0, i_13_494_3487_0,
    i_13_494_3489_0, i_13_494_3504_0, i_13_494_3550_0, i_13_494_3552_0,
    i_13_494_3565_0, i_13_494_3566_0, i_13_494_3568_0, i_13_494_3577_0,
    i_13_494_3603_0, i_13_494_3648_0, i_13_494_3681_0, i_13_494_3763_0,
    i_13_494_3764_0, i_13_494_3803_0, i_13_494_3819_0, i_13_494_3822_0,
    i_13_494_3862_0, i_13_494_3865_0, i_13_494_3980_0, i_13_494_4054_0,
    i_13_494_4163_0, i_13_494_4251_0, i_13_494_4312_0, i_13_494_4325_0,
    i_13_494_4340_0, i_13_494_4366_0, i_13_494_4367_0, i_13_494_4369_0,
    i_13_494_4370_0, i_13_494_4372_0, i_13_494_4396_0, i_13_494_4479_0,
    i_13_494_4558_0, i_13_494_4560_0, i_13_494_4568_0, i_13_494_4600_0;
  output o_13_494_0_0;
  assign o_13_494_0_0 = ~((~i_13_494_4560_0 & ((~i_13_494_3577_0 & ((~i_13_494_3552_0 & ~i_13_494_3862_0 & ~i_13_494_4163_0) | (~i_13_494_1660_0 & ~i_13_494_4372_0 & ~i_13_494_4558_0))) | (~i_13_494_3013_0 & ~i_13_494_3484_0 & ~i_13_494_3565_0 & ~i_13_494_3822_0))) | (i_13_494_229_0 & ~i_13_494_940_0 & ~i_13_494_2742_0 & ~i_13_494_3460_0 & ~i_13_494_3463_0 & ~i_13_494_3483_0 & ~i_13_494_3566_0) | (~i_13_494_573_0 & ~i_13_494_938_0 & ~i_13_494_2425_0 & ~i_13_494_4325_0 & ~i_13_494_4366_0 & ~i_13_494_4372_0) | (~i_13_494_3550_0 & i_13_494_4163_0 & i_13_494_4372_0) | (~i_13_494_3865_0 & i_13_494_4396_0));
endmodule



// Benchmark "kernel_13_495" written by ABC on Sun Jul 19 10:52:13 2020

module kernel_13_495 ( 
    i_13_495_42_0, i_13_495_43_0, i_13_495_76_0, i_13_495_102_0,
    i_13_495_107_0, i_13_495_117_0, i_13_495_118_0, i_13_495_169_0,
    i_13_495_180_0, i_13_495_181_0, i_13_495_225_0, i_13_495_394_0,
    i_13_495_489_0, i_13_495_504_0, i_13_495_534_0, i_13_495_567_0,
    i_13_495_572_0, i_13_495_607_0, i_13_495_617_0, i_13_495_624_0,
    i_13_495_645_0, i_13_495_651_0, i_13_495_697_0, i_13_495_711_0,
    i_13_495_835_0, i_13_495_841_0, i_13_495_945_0, i_13_495_948_0,
    i_13_495_1072_0, i_13_495_1092_0, i_13_495_1115_0, i_13_495_1210_0,
    i_13_495_1225_0, i_13_495_1276_0, i_13_495_1300_0, i_13_495_1404_0,
    i_13_495_1522_0, i_13_495_1629_0, i_13_495_1719_0, i_13_495_1767_0,
    i_13_495_1782_0, i_13_495_1783_0, i_13_495_1785_0, i_13_495_1786_0,
    i_13_495_1801_0, i_13_495_2014_0, i_13_495_2056_0, i_13_495_2119_0,
    i_13_495_2182_0, i_13_495_2205_0, i_13_495_2206_0, i_13_495_2209_0,
    i_13_495_2280_0, i_13_495_2307_0, i_13_495_2321_0, i_13_495_2361_0,
    i_13_495_2394_0, i_13_495_2403_0, i_13_495_2427_0, i_13_495_2428_0,
    i_13_495_2452_0, i_13_495_2457_0, i_13_495_2458_0, i_13_495_2680_0,
    i_13_495_2879_0, i_13_495_2934_0, i_13_495_2938_0, i_13_495_3015_0,
    i_13_495_3019_0, i_13_495_3160_0, i_13_495_3163_0, i_13_495_3171_0,
    i_13_495_3204_0, i_13_495_3213_0, i_13_495_3214_0, i_13_495_3217_0,
    i_13_495_3231_0, i_13_495_3270_0, i_13_495_3420_0, i_13_495_3421_0,
    i_13_495_3426_0, i_13_495_3531_0, i_13_495_3532_0, i_13_495_3548_0,
    i_13_495_3562_0, i_13_495_3699_0, i_13_495_3745_0, i_13_495_3870_0,
    i_13_495_3873_0, i_13_495_3912_0, i_13_495_3981_0, i_13_495_3982_0,
    i_13_495_4005_0, i_13_495_4006_0, i_13_495_4017_0, i_13_495_4254_0,
    i_13_495_4302_0, i_13_495_4311_0, i_13_495_4413_0, i_13_495_4518_0,
    o_13_495_0_0  );
  input  i_13_495_42_0, i_13_495_43_0, i_13_495_76_0, i_13_495_102_0,
    i_13_495_107_0, i_13_495_117_0, i_13_495_118_0, i_13_495_169_0,
    i_13_495_180_0, i_13_495_181_0, i_13_495_225_0, i_13_495_394_0,
    i_13_495_489_0, i_13_495_504_0, i_13_495_534_0, i_13_495_567_0,
    i_13_495_572_0, i_13_495_607_0, i_13_495_617_0, i_13_495_624_0,
    i_13_495_645_0, i_13_495_651_0, i_13_495_697_0, i_13_495_711_0,
    i_13_495_835_0, i_13_495_841_0, i_13_495_945_0, i_13_495_948_0,
    i_13_495_1072_0, i_13_495_1092_0, i_13_495_1115_0, i_13_495_1210_0,
    i_13_495_1225_0, i_13_495_1276_0, i_13_495_1300_0, i_13_495_1404_0,
    i_13_495_1522_0, i_13_495_1629_0, i_13_495_1719_0, i_13_495_1767_0,
    i_13_495_1782_0, i_13_495_1783_0, i_13_495_1785_0, i_13_495_1786_0,
    i_13_495_1801_0, i_13_495_2014_0, i_13_495_2056_0, i_13_495_2119_0,
    i_13_495_2182_0, i_13_495_2205_0, i_13_495_2206_0, i_13_495_2209_0,
    i_13_495_2280_0, i_13_495_2307_0, i_13_495_2321_0, i_13_495_2361_0,
    i_13_495_2394_0, i_13_495_2403_0, i_13_495_2427_0, i_13_495_2428_0,
    i_13_495_2452_0, i_13_495_2457_0, i_13_495_2458_0, i_13_495_2680_0,
    i_13_495_2879_0, i_13_495_2934_0, i_13_495_2938_0, i_13_495_3015_0,
    i_13_495_3019_0, i_13_495_3160_0, i_13_495_3163_0, i_13_495_3171_0,
    i_13_495_3204_0, i_13_495_3213_0, i_13_495_3214_0, i_13_495_3217_0,
    i_13_495_3231_0, i_13_495_3270_0, i_13_495_3420_0, i_13_495_3421_0,
    i_13_495_3426_0, i_13_495_3531_0, i_13_495_3532_0, i_13_495_3548_0,
    i_13_495_3562_0, i_13_495_3699_0, i_13_495_3745_0, i_13_495_3870_0,
    i_13_495_3873_0, i_13_495_3912_0, i_13_495_3981_0, i_13_495_3982_0,
    i_13_495_4005_0, i_13_495_4006_0, i_13_495_4017_0, i_13_495_4254_0,
    i_13_495_4302_0, i_13_495_4311_0, i_13_495_4413_0, i_13_495_4518_0;
  output o_13_495_0_0;
  assign o_13_495_0_0 = ~((~i_13_495_3420_0 & ((~i_13_495_117_0 & i_13_495_2056_0) | (~i_13_495_3204_0 & ~i_13_495_3217_0))) | (~i_13_495_3981_0 & ~i_13_495_4006_0) | (~i_13_495_180_0 & ~i_13_495_2206_0 & ~i_13_495_4311_0));
endmodule



// Benchmark "kernel_13_496" written by ABC on Sun Jul 19 10:52:14 2020

module kernel_13_496 ( 
    i_13_496_71_0, i_13_496_79_0, i_13_496_169_0, i_13_496_171_0,
    i_13_496_175_0, i_13_496_216_0, i_13_496_233_0, i_13_496_246_0,
    i_13_496_325_0, i_13_496_397_0, i_13_496_604_0, i_13_496_613_0,
    i_13_496_624_0, i_13_496_643_0, i_13_496_679_0, i_13_496_683_0,
    i_13_496_685_0, i_13_496_694_0, i_13_496_697_0, i_13_496_819_0,
    i_13_496_822_0, i_13_496_826_0, i_13_496_841_0, i_13_496_854_0,
    i_13_496_855_0, i_13_496_878_0, i_13_496_937_0, i_13_496_973_0,
    i_13_496_1021_0, i_13_496_1062_0, i_13_496_1119_0, i_13_496_1120_0,
    i_13_496_1132_0, i_13_496_1224_0, i_13_496_1225_0, i_13_496_1308_0,
    i_13_496_1313_0, i_13_496_1315_0, i_13_496_1377_0, i_13_496_1485_0,
    i_13_496_1506_0, i_13_496_1525_0, i_13_496_1553_0, i_13_496_1663_0,
    i_13_496_1745_0, i_13_496_1771_0, i_13_496_1798_0, i_13_496_1799_0,
    i_13_496_1944_0, i_13_496_1948_0, i_13_496_1954_0, i_13_496_2000_0,
    i_13_496_2383_0, i_13_496_2452_0, i_13_496_2677_0, i_13_496_2749_0,
    i_13_496_2848_0, i_13_496_2878_0, i_13_496_3006_0, i_13_496_3007_0,
    i_13_496_3008_0, i_13_496_3094_0, i_13_496_3107_0, i_13_496_3168_0,
    i_13_496_3216_0, i_13_496_3352_0, i_13_496_3424_0, i_13_496_3429_0,
    i_13_496_3450_0, i_13_496_3487_0, i_13_496_3506_0, i_13_496_3538_0,
    i_13_496_3652_0, i_13_496_3728_0, i_13_496_3739_0, i_13_496_3742_0,
    i_13_496_3782_0, i_13_496_3895_0, i_13_496_3927_0, i_13_496_3937_0,
    i_13_496_3982_0, i_13_496_3994_0, i_13_496_4063_0, i_13_496_4096_0,
    i_13_496_4186_0, i_13_496_4188_0, i_13_496_4249_0, i_13_496_4252_0,
    i_13_496_4255_0, i_13_496_4256_0, i_13_496_4258_0, i_13_496_4261_0,
    i_13_496_4297_0, i_13_496_4300_0, i_13_496_4366_0, i_13_496_4372_0,
    i_13_496_4433_0, i_13_496_4447_0, i_13_496_4536_0, i_13_496_4598_0,
    o_13_496_0_0  );
  input  i_13_496_71_0, i_13_496_79_0, i_13_496_169_0, i_13_496_171_0,
    i_13_496_175_0, i_13_496_216_0, i_13_496_233_0, i_13_496_246_0,
    i_13_496_325_0, i_13_496_397_0, i_13_496_604_0, i_13_496_613_0,
    i_13_496_624_0, i_13_496_643_0, i_13_496_679_0, i_13_496_683_0,
    i_13_496_685_0, i_13_496_694_0, i_13_496_697_0, i_13_496_819_0,
    i_13_496_822_0, i_13_496_826_0, i_13_496_841_0, i_13_496_854_0,
    i_13_496_855_0, i_13_496_878_0, i_13_496_937_0, i_13_496_973_0,
    i_13_496_1021_0, i_13_496_1062_0, i_13_496_1119_0, i_13_496_1120_0,
    i_13_496_1132_0, i_13_496_1224_0, i_13_496_1225_0, i_13_496_1308_0,
    i_13_496_1313_0, i_13_496_1315_0, i_13_496_1377_0, i_13_496_1485_0,
    i_13_496_1506_0, i_13_496_1525_0, i_13_496_1553_0, i_13_496_1663_0,
    i_13_496_1745_0, i_13_496_1771_0, i_13_496_1798_0, i_13_496_1799_0,
    i_13_496_1944_0, i_13_496_1948_0, i_13_496_1954_0, i_13_496_2000_0,
    i_13_496_2383_0, i_13_496_2452_0, i_13_496_2677_0, i_13_496_2749_0,
    i_13_496_2848_0, i_13_496_2878_0, i_13_496_3006_0, i_13_496_3007_0,
    i_13_496_3008_0, i_13_496_3094_0, i_13_496_3107_0, i_13_496_3168_0,
    i_13_496_3216_0, i_13_496_3352_0, i_13_496_3424_0, i_13_496_3429_0,
    i_13_496_3450_0, i_13_496_3487_0, i_13_496_3506_0, i_13_496_3538_0,
    i_13_496_3652_0, i_13_496_3728_0, i_13_496_3739_0, i_13_496_3742_0,
    i_13_496_3782_0, i_13_496_3895_0, i_13_496_3927_0, i_13_496_3937_0,
    i_13_496_3982_0, i_13_496_3994_0, i_13_496_4063_0, i_13_496_4096_0,
    i_13_496_4186_0, i_13_496_4188_0, i_13_496_4249_0, i_13_496_4252_0,
    i_13_496_4255_0, i_13_496_4256_0, i_13_496_4258_0, i_13_496_4261_0,
    i_13_496_4297_0, i_13_496_4300_0, i_13_496_4366_0, i_13_496_4372_0,
    i_13_496_4433_0, i_13_496_4447_0, i_13_496_4536_0, i_13_496_4598_0;
  output o_13_496_0_0;
  assign o_13_496_0_0 = 0;
endmodule



// Benchmark "kernel_13_497" written by ABC on Sun Jul 19 10:52:15 2020

module kernel_13_497 ( 
    i_13_497_69_0, i_13_497_142_0, i_13_497_385_0, i_13_497_386_0,
    i_13_497_448_0, i_13_497_537_0, i_13_497_664_0, i_13_497_691_0,
    i_13_497_836_0, i_13_497_844_0, i_13_497_848_0, i_13_497_892_0,
    i_13_497_989_0, i_13_497_1102_0, i_13_497_1219_0, i_13_497_1228_0,
    i_13_497_1276_0, i_13_497_1287_0, i_13_497_1345_0, i_13_497_1402_0,
    i_13_497_1403_0, i_13_497_1444_0, i_13_497_1510_0, i_13_497_1600_0,
    i_13_497_1644_0, i_13_497_1678_0, i_13_497_1717_0, i_13_497_1725_0,
    i_13_497_1726_0, i_13_497_1748_0, i_13_497_1934_0, i_13_497_1948_0,
    i_13_497_1960_0, i_13_497_1995_0, i_13_497_1996_0, i_13_497_1999_0,
    i_13_497_2002_0, i_13_497_2060_0, i_13_497_2127_0, i_13_497_2194_0,
    i_13_497_2281_0, i_13_497_2311_0, i_13_497_2361_0, i_13_497_2379_0,
    i_13_497_2464_0, i_13_497_2470_0, i_13_497_2534_0, i_13_497_2698_0,
    i_13_497_2716_0, i_13_497_2726_0, i_13_497_2771_0, i_13_497_2857_0,
    i_13_497_2860_0, i_13_497_2887_0, i_13_497_2917_0, i_13_497_2949_0,
    i_13_497_3017_0, i_13_497_3028_0, i_13_497_3065_0, i_13_497_3066_0,
    i_13_497_3067_0, i_13_497_3068_0, i_13_497_3074_0, i_13_497_3329_0,
    i_13_497_3352_0, i_13_497_3446_0, i_13_497_3454_0, i_13_497_3490_0,
    i_13_497_3547_0, i_13_497_3595_0, i_13_497_3683_0, i_13_497_3686_0,
    i_13_497_3688_0, i_13_497_3689_0, i_13_497_3722_0, i_13_497_3737_0,
    i_13_497_3781_0, i_13_497_3900_0, i_13_497_3928_0, i_13_497_3988_0,
    i_13_497_3994_0, i_13_497_3995_0, i_13_497_4017_0, i_13_497_4054_0,
    i_13_497_4057_0, i_13_497_4094_0, i_13_497_4165_0, i_13_497_4214_0,
    i_13_497_4273_0, i_13_497_4304_0, i_13_497_4309_0, i_13_497_4393_0,
    i_13_497_4396_0, i_13_497_4399_0, i_13_497_4400_0, i_13_497_4411_0,
    i_13_497_4431_0, i_13_497_4432_0, i_13_497_4566_0, i_13_497_4597_0,
    o_13_497_0_0  );
  input  i_13_497_69_0, i_13_497_142_0, i_13_497_385_0, i_13_497_386_0,
    i_13_497_448_0, i_13_497_537_0, i_13_497_664_0, i_13_497_691_0,
    i_13_497_836_0, i_13_497_844_0, i_13_497_848_0, i_13_497_892_0,
    i_13_497_989_0, i_13_497_1102_0, i_13_497_1219_0, i_13_497_1228_0,
    i_13_497_1276_0, i_13_497_1287_0, i_13_497_1345_0, i_13_497_1402_0,
    i_13_497_1403_0, i_13_497_1444_0, i_13_497_1510_0, i_13_497_1600_0,
    i_13_497_1644_0, i_13_497_1678_0, i_13_497_1717_0, i_13_497_1725_0,
    i_13_497_1726_0, i_13_497_1748_0, i_13_497_1934_0, i_13_497_1948_0,
    i_13_497_1960_0, i_13_497_1995_0, i_13_497_1996_0, i_13_497_1999_0,
    i_13_497_2002_0, i_13_497_2060_0, i_13_497_2127_0, i_13_497_2194_0,
    i_13_497_2281_0, i_13_497_2311_0, i_13_497_2361_0, i_13_497_2379_0,
    i_13_497_2464_0, i_13_497_2470_0, i_13_497_2534_0, i_13_497_2698_0,
    i_13_497_2716_0, i_13_497_2726_0, i_13_497_2771_0, i_13_497_2857_0,
    i_13_497_2860_0, i_13_497_2887_0, i_13_497_2917_0, i_13_497_2949_0,
    i_13_497_3017_0, i_13_497_3028_0, i_13_497_3065_0, i_13_497_3066_0,
    i_13_497_3067_0, i_13_497_3068_0, i_13_497_3074_0, i_13_497_3329_0,
    i_13_497_3352_0, i_13_497_3446_0, i_13_497_3454_0, i_13_497_3490_0,
    i_13_497_3547_0, i_13_497_3595_0, i_13_497_3683_0, i_13_497_3686_0,
    i_13_497_3688_0, i_13_497_3689_0, i_13_497_3722_0, i_13_497_3737_0,
    i_13_497_3781_0, i_13_497_3900_0, i_13_497_3928_0, i_13_497_3988_0,
    i_13_497_3994_0, i_13_497_3995_0, i_13_497_4017_0, i_13_497_4054_0,
    i_13_497_4057_0, i_13_497_4094_0, i_13_497_4165_0, i_13_497_4214_0,
    i_13_497_4273_0, i_13_497_4304_0, i_13_497_4309_0, i_13_497_4393_0,
    i_13_497_4396_0, i_13_497_4399_0, i_13_497_4400_0, i_13_497_4411_0,
    i_13_497_4431_0, i_13_497_4432_0, i_13_497_4566_0, i_13_497_4597_0;
  output o_13_497_0_0;
  assign o_13_497_0_0 = ~((i_13_497_1228_0 & ~i_13_497_4165_0) | (~i_13_497_3067_0 & ~i_13_497_3688_0) | (~i_13_497_1510_0 & ~i_13_497_1717_0 & ~i_13_497_2857_0));
endmodule



// Benchmark "kernel_13_498" written by ABC on Sun Jul 19 10:52:15 2020

module kernel_13_498 ( 
    i_13_498_77_0, i_13_498_130_0, i_13_498_134_0, i_13_498_256_0,
    i_13_498_368_0, i_13_498_394_0, i_13_498_469_0, i_13_498_515_0,
    i_13_498_518_0, i_13_498_550_0, i_13_498_554_0, i_13_498_605_0,
    i_13_498_623_0, i_13_498_626_0, i_13_498_656_0, i_13_498_658_0,
    i_13_498_659_0, i_13_498_661_0, i_13_498_695_0, i_13_498_698_0,
    i_13_498_814_0, i_13_498_841_0, i_13_498_889_0, i_13_498_940_0,
    i_13_498_978_0, i_13_498_1063_0, i_13_498_1072_0, i_13_498_1073_0,
    i_13_498_1084_0, i_13_498_1088_0, i_13_498_1109_0, i_13_498_1144_0,
    i_13_498_1145_0, i_13_498_1153_0, i_13_498_1154_0, i_13_498_1214_0,
    i_13_498_1265_0, i_13_498_1424_0, i_13_498_1517_0, i_13_498_1535_0,
    i_13_498_1657_0, i_13_498_1658_0, i_13_498_1660_0, i_13_498_1730_0,
    i_13_498_1732_0, i_13_498_1733_0, i_13_498_1742_0, i_13_498_2017_0,
    i_13_498_2020_0, i_13_498_2021_0, i_13_498_2023_0, i_13_498_2131_0,
    i_13_498_2137_0, i_13_498_2209_0, i_13_498_2246_0, i_13_498_2297_0,
    i_13_498_2336_0, i_13_498_2401_0, i_13_498_2443_0, i_13_498_2461_0,
    i_13_498_2498_0, i_13_498_2513_0, i_13_498_2717_0, i_13_498_2740_0,
    i_13_498_2771_0, i_13_498_2882_0, i_13_498_2956_0, i_13_498_3044_0,
    i_13_498_3074_0, i_13_498_3075_0, i_13_498_3115_0, i_13_498_3154_0,
    i_13_498_3263_0, i_13_498_3476_0, i_13_498_3563_0, i_13_498_3568_0,
    i_13_498_3730_0, i_13_498_3740_0, i_13_498_3820_0, i_13_498_3910_0,
    i_13_498_4019_0, i_13_498_4091_0, i_13_498_4121_0, i_13_498_4160_0,
    i_13_498_4163_0, i_13_498_4187_0, i_13_498_4330_0, i_13_498_4333_0,
    i_13_498_4358_0, i_13_498_4360_0, i_13_498_4362_0, i_13_498_4363_0,
    i_13_498_4366_0, i_13_498_4367_0, i_13_498_4394_0, i_13_498_4429_0,
    i_13_498_4477_0, i_13_498_4514_0, i_13_498_4540_0, i_13_498_4603_0,
    o_13_498_0_0  );
  input  i_13_498_77_0, i_13_498_130_0, i_13_498_134_0, i_13_498_256_0,
    i_13_498_368_0, i_13_498_394_0, i_13_498_469_0, i_13_498_515_0,
    i_13_498_518_0, i_13_498_550_0, i_13_498_554_0, i_13_498_605_0,
    i_13_498_623_0, i_13_498_626_0, i_13_498_656_0, i_13_498_658_0,
    i_13_498_659_0, i_13_498_661_0, i_13_498_695_0, i_13_498_698_0,
    i_13_498_814_0, i_13_498_841_0, i_13_498_889_0, i_13_498_940_0,
    i_13_498_978_0, i_13_498_1063_0, i_13_498_1072_0, i_13_498_1073_0,
    i_13_498_1084_0, i_13_498_1088_0, i_13_498_1109_0, i_13_498_1144_0,
    i_13_498_1145_0, i_13_498_1153_0, i_13_498_1154_0, i_13_498_1214_0,
    i_13_498_1265_0, i_13_498_1424_0, i_13_498_1517_0, i_13_498_1535_0,
    i_13_498_1657_0, i_13_498_1658_0, i_13_498_1660_0, i_13_498_1730_0,
    i_13_498_1732_0, i_13_498_1733_0, i_13_498_1742_0, i_13_498_2017_0,
    i_13_498_2020_0, i_13_498_2021_0, i_13_498_2023_0, i_13_498_2131_0,
    i_13_498_2137_0, i_13_498_2209_0, i_13_498_2246_0, i_13_498_2297_0,
    i_13_498_2336_0, i_13_498_2401_0, i_13_498_2443_0, i_13_498_2461_0,
    i_13_498_2498_0, i_13_498_2513_0, i_13_498_2717_0, i_13_498_2740_0,
    i_13_498_2771_0, i_13_498_2882_0, i_13_498_2956_0, i_13_498_3044_0,
    i_13_498_3074_0, i_13_498_3075_0, i_13_498_3115_0, i_13_498_3154_0,
    i_13_498_3263_0, i_13_498_3476_0, i_13_498_3563_0, i_13_498_3568_0,
    i_13_498_3730_0, i_13_498_3740_0, i_13_498_3820_0, i_13_498_3910_0,
    i_13_498_4019_0, i_13_498_4091_0, i_13_498_4121_0, i_13_498_4160_0,
    i_13_498_4163_0, i_13_498_4187_0, i_13_498_4330_0, i_13_498_4333_0,
    i_13_498_4358_0, i_13_498_4360_0, i_13_498_4362_0, i_13_498_4363_0,
    i_13_498_4366_0, i_13_498_4367_0, i_13_498_4394_0, i_13_498_4429_0,
    i_13_498_4477_0, i_13_498_4514_0, i_13_498_4540_0, i_13_498_4603_0;
  output o_13_498_0_0;
  assign o_13_498_0_0 = ~((~i_13_498_1660_0 & ((~i_13_498_256_0 & ~i_13_498_1730_0) | (~i_13_498_1144_0 & ~i_13_498_2882_0))) | (~i_13_498_518_0 & ~i_13_498_2017_0 & ~i_13_498_2717_0) | (~i_13_498_656_0 & ~i_13_498_1730_0 & ~i_13_498_2740_0) | (~i_13_498_1084_0 & ~i_13_498_1265_0 & ~i_13_498_4360_0) | (~i_13_498_698_0 & ~i_13_498_1657_0 & ~i_13_498_2882_0 & ~i_13_498_3740_0 & ~i_13_498_4330_0 & ~i_13_498_4394_0));
endmodule



// Benchmark "kernel_13_499" written by ABC on Sun Jul 19 10:52:16 2020

module kernel_13_499 ( 
    i_13_499_46_0, i_13_499_139_0, i_13_499_185_0, i_13_499_331_0,
    i_13_499_334_0, i_13_499_335_0, i_13_499_352_0, i_13_499_362_0,
    i_13_499_409_0, i_13_499_449_0, i_13_499_451_0, i_13_499_506_0,
    i_13_499_568_0, i_13_499_626_0, i_13_499_649_0, i_13_499_658_0,
    i_13_499_769_0, i_13_499_884_0, i_13_499_932_0, i_13_499_935_0,
    i_13_499_937_0, i_13_499_1019_0, i_13_499_1024_0, i_13_499_1072_0,
    i_13_499_1073_0, i_13_499_1129_0, i_13_499_1130_0, i_13_499_1133_0,
    i_13_499_1148_0, i_13_499_1189_0, i_13_499_1244_0, i_13_499_1298_0,
    i_13_499_1328_0, i_13_499_1400_0, i_13_499_1406_0, i_13_499_1510_0,
    i_13_499_1523_0, i_13_499_1570_0, i_13_499_1649_0, i_13_499_1661_0,
    i_13_499_1679_0, i_13_499_1720_0, i_13_499_1727_0, i_13_499_1765_0,
    i_13_499_1888_0, i_13_499_1889_0, i_13_499_1933_0, i_13_499_1945_0,
    i_13_499_2026_0, i_13_499_2027_0, i_13_499_2135_0, i_13_499_2188_0,
    i_13_499_2197_0, i_13_499_2423_0, i_13_499_2470_0, i_13_499_2645_0,
    i_13_499_2694_0, i_13_499_2725_0, i_13_499_2741_0, i_13_499_2747_0,
    i_13_499_2801_0, i_13_499_2851_0, i_13_499_2899_0, i_13_499_2917_0,
    i_13_499_2966_0, i_13_499_2998_0, i_13_499_3028_0, i_13_499_3029_0,
    i_13_499_3073_0, i_13_499_3074_0, i_13_499_3163_0, i_13_499_3261_0,
    i_13_499_3262_0, i_13_499_3325_0, i_13_499_3378_0, i_13_499_3458_0,
    i_13_499_3484_0, i_13_499_3485_0, i_13_499_3547_0, i_13_499_3574_0,
    i_13_499_3575_0, i_13_499_3653_0, i_13_499_3728_0, i_13_499_3742_0,
    i_13_499_3760_0, i_13_499_3764_0, i_13_499_3781_0, i_13_499_3785_0,
    i_13_499_3853_0, i_13_499_3898_0, i_13_499_3899_0, i_13_499_4162_0,
    i_13_499_4231_0, i_13_499_4294_0, i_13_499_4298_0, i_13_499_4322_0,
    i_13_499_4360_0, i_13_499_4363_0, i_13_499_4537_0, i_13_499_4603_0,
    o_13_499_0_0  );
  input  i_13_499_46_0, i_13_499_139_0, i_13_499_185_0, i_13_499_331_0,
    i_13_499_334_0, i_13_499_335_0, i_13_499_352_0, i_13_499_362_0,
    i_13_499_409_0, i_13_499_449_0, i_13_499_451_0, i_13_499_506_0,
    i_13_499_568_0, i_13_499_626_0, i_13_499_649_0, i_13_499_658_0,
    i_13_499_769_0, i_13_499_884_0, i_13_499_932_0, i_13_499_935_0,
    i_13_499_937_0, i_13_499_1019_0, i_13_499_1024_0, i_13_499_1072_0,
    i_13_499_1073_0, i_13_499_1129_0, i_13_499_1130_0, i_13_499_1133_0,
    i_13_499_1148_0, i_13_499_1189_0, i_13_499_1244_0, i_13_499_1298_0,
    i_13_499_1328_0, i_13_499_1400_0, i_13_499_1406_0, i_13_499_1510_0,
    i_13_499_1523_0, i_13_499_1570_0, i_13_499_1649_0, i_13_499_1661_0,
    i_13_499_1679_0, i_13_499_1720_0, i_13_499_1727_0, i_13_499_1765_0,
    i_13_499_1888_0, i_13_499_1889_0, i_13_499_1933_0, i_13_499_1945_0,
    i_13_499_2026_0, i_13_499_2027_0, i_13_499_2135_0, i_13_499_2188_0,
    i_13_499_2197_0, i_13_499_2423_0, i_13_499_2470_0, i_13_499_2645_0,
    i_13_499_2694_0, i_13_499_2725_0, i_13_499_2741_0, i_13_499_2747_0,
    i_13_499_2801_0, i_13_499_2851_0, i_13_499_2899_0, i_13_499_2917_0,
    i_13_499_2966_0, i_13_499_2998_0, i_13_499_3028_0, i_13_499_3029_0,
    i_13_499_3073_0, i_13_499_3074_0, i_13_499_3163_0, i_13_499_3261_0,
    i_13_499_3262_0, i_13_499_3325_0, i_13_499_3378_0, i_13_499_3458_0,
    i_13_499_3484_0, i_13_499_3485_0, i_13_499_3547_0, i_13_499_3574_0,
    i_13_499_3575_0, i_13_499_3653_0, i_13_499_3728_0, i_13_499_3742_0,
    i_13_499_3760_0, i_13_499_3764_0, i_13_499_3781_0, i_13_499_3785_0,
    i_13_499_3853_0, i_13_499_3898_0, i_13_499_3899_0, i_13_499_4162_0,
    i_13_499_4231_0, i_13_499_4294_0, i_13_499_4298_0, i_13_499_4322_0,
    i_13_499_4360_0, i_13_499_4363_0, i_13_499_4537_0, i_13_499_4603_0;
  output o_13_499_0_0;
  assign o_13_499_0_0 = ~((~i_13_499_1523_0 & ((~i_13_499_1945_0 & ~i_13_499_2423_0 & ~i_13_499_3899_0) | (~i_13_499_3575_0 & ~i_13_499_3898_0 & ~i_13_499_4322_0))) | (~i_13_499_937_0 & ~i_13_499_1148_0) | (~i_13_499_1679_0 & ~i_13_499_3485_0 & ~i_13_499_3853_0 & ~i_13_499_4360_0));
endmodule



// Benchmark "kernel_13_500" written by ABC on Sun Jul 19 10:52:17 2020

module kernel_13_500 ( 
    i_13_500_46_0, i_13_500_47_0, i_13_500_121_0, i_13_500_226_0,
    i_13_500_357_0, i_13_500_407_0, i_13_500_447_0, i_13_500_514_0,
    i_13_500_532_0, i_13_500_568_0, i_13_500_794_0, i_13_500_833_0,
    i_13_500_847_0, i_13_500_848_0, i_13_500_931_0, i_13_500_937_0,
    i_13_500_947_0, i_13_500_1019_0, i_13_500_1072_0, i_13_500_1073_0,
    i_13_500_1136_0, i_13_500_1201_0, i_13_500_1225_0, i_13_500_1298_0,
    i_13_500_1315_0, i_13_500_1495_0, i_13_500_1496_0, i_13_500_1630_0,
    i_13_500_1631_0, i_13_500_1720_0, i_13_500_1724_0, i_13_500_1777_0,
    i_13_500_1779_0, i_13_500_1805_0, i_13_500_1855_0, i_13_500_1945_0,
    i_13_500_1946_0, i_13_500_1948_0, i_13_500_2020_0, i_13_500_2026_0,
    i_13_500_2027_0, i_13_500_2099_0, i_13_500_2134_0, i_13_500_2197_0,
    i_13_500_2198_0, i_13_500_2227_0, i_13_500_2449_0, i_13_500_2450_0,
    i_13_500_2452_0, i_13_500_2459_0, i_13_500_2477_0, i_13_500_2539_0,
    i_13_500_2540_0, i_13_500_2548_0, i_13_500_2740_0, i_13_500_2782_0,
    i_13_500_2917_0, i_13_500_2918_0, i_13_500_3010_0, i_13_500_3028_0,
    i_13_500_3097_0, i_13_500_3169_0, i_13_500_3268_0, i_13_500_3397_0,
    i_13_500_3412_0, i_13_500_3451_0, i_13_500_3457_0, i_13_500_3458_0,
    i_13_500_3484_0, i_13_500_3570_0, i_13_500_3574_0, i_13_500_3575_0,
    i_13_500_3593_0, i_13_500_3704_0, i_13_500_3728_0, i_13_500_3781_0,
    i_13_500_3782_0, i_13_500_3800_0, i_13_500_3853_0, i_13_500_3898_0,
    i_13_500_3907_0, i_13_500_3908_0, i_13_500_4001_0, i_13_500_4016_0,
    i_13_500_4249_0, i_13_500_4250_0, i_13_500_4252_0, i_13_500_4253_0,
    i_13_500_4259_0, i_13_500_4322_0, i_13_500_4339_0, i_13_500_4342_0,
    i_13_500_4365_0, i_13_500_4375_0, i_13_500_4376_0, i_13_500_4447_0,
    i_13_500_4511_0, i_13_500_4556_0, i_13_500_4558_0, i_13_500_4570_0,
    o_13_500_0_0  );
  input  i_13_500_46_0, i_13_500_47_0, i_13_500_121_0, i_13_500_226_0,
    i_13_500_357_0, i_13_500_407_0, i_13_500_447_0, i_13_500_514_0,
    i_13_500_532_0, i_13_500_568_0, i_13_500_794_0, i_13_500_833_0,
    i_13_500_847_0, i_13_500_848_0, i_13_500_931_0, i_13_500_937_0,
    i_13_500_947_0, i_13_500_1019_0, i_13_500_1072_0, i_13_500_1073_0,
    i_13_500_1136_0, i_13_500_1201_0, i_13_500_1225_0, i_13_500_1298_0,
    i_13_500_1315_0, i_13_500_1495_0, i_13_500_1496_0, i_13_500_1630_0,
    i_13_500_1631_0, i_13_500_1720_0, i_13_500_1724_0, i_13_500_1777_0,
    i_13_500_1779_0, i_13_500_1805_0, i_13_500_1855_0, i_13_500_1945_0,
    i_13_500_1946_0, i_13_500_1948_0, i_13_500_2020_0, i_13_500_2026_0,
    i_13_500_2027_0, i_13_500_2099_0, i_13_500_2134_0, i_13_500_2197_0,
    i_13_500_2198_0, i_13_500_2227_0, i_13_500_2449_0, i_13_500_2450_0,
    i_13_500_2452_0, i_13_500_2459_0, i_13_500_2477_0, i_13_500_2539_0,
    i_13_500_2540_0, i_13_500_2548_0, i_13_500_2740_0, i_13_500_2782_0,
    i_13_500_2917_0, i_13_500_2918_0, i_13_500_3010_0, i_13_500_3028_0,
    i_13_500_3097_0, i_13_500_3169_0, i_13_500_3268_0, i_13_500_3397_0,
    i_13_500_3412_0, i_13_500_3451_0, i_13_500_3457_0, i_13_500_3458_0,
    i_13_500_3484_0, i_13_500_3570_0, i_13_500_3574_0, i_13_500_3575_0,
    i_13_500_3593_0, i_13_500_3704_0, i_13_500_3728_0, i_13_500_3781_0,
    i_13_500_3782_0, i_13_500_3800_0, i_13_500_3853_0, i_13_500_3898_0,
    i_13_500_3907_0, i_13_500_3908_0, i_13_500_4001_0, i_13_500_4016_0,
    i_13_500_4249_0, i_13_500_4250_0, i_13_500_4252_0, i_13_500_4253_0,
    i_13_500_4259_0, i_13_500_4322_0, i_13_500_4339_0, i_13_500_4342_0,
    i_13_500_4365_0, i_13_500_4375_0, i_13_500_4376_0, i_13_500_4447_0,
    i_13_500_4511_0, i_13_500_4556_0, i_13_500_4558_0, i_13_500_4570_0;
  output o_13_500_0_0;
  assign o_13_500_0_0 = ~(~i_13_500_3593_0 | (~i_13_500_2197_0 & ~i_13_500_3574_0));
endmodule



// Benchmark "kernel_13_501" written by ABC on Sun Jul 19 10:52:18 2020

module kernel_13_501 ( 
    i_13_501_31_0, i_13_501_36_0, i_13_501_37_0, i_13_501_102_0,
    i_13_501_255_0, i_13_501_262_0, i_13_501_264_0, i_13_501_265_0,
    i_13_501_282_0, i_13_501_492_0, i_13_501_505_0, i_13_501_532_0,
    i_13_501_535_0, i_13_501_577_0, i_13_501_616_0, i_13_501_651_0,
    i_13_501_675_0, i_13_501_676_0, i_13_501_723_0, i_13_501_777_0,
    i_13_501_810_0, i_13_501_837_0, i_13_501_838_0, i_13_501_871_0,
    i_13_501_948_0, i_13_501_949_0, i_13_501_981_0, i_13_501_1116_0,
    i_13_501_1197_0, i_13_501_1198_0, i_13_501_1212_0, i_13_501_1242_0,
    i_13_501_1269_0, i_13_501_1278_0, i_13_501_1324_0, i_13_501_1326_0,
    i_13_501_1380_0, i_13_501_1396_0, i_13_501_1446_0, i_13_501_1456_0,
    i_13_501_1504_0, i_13_501_1552_0, i_13_501_1746_0, i_13_501_1786_0,
    i_13_501_1803_0, i_13_501_1840_0, i_13_501_1857_0, i_13_501_1908_0,
    i_13_501_2010_0, i_13_501_2029_0, i_13_501_2046_0, i_13_501_2055_0,
    i_13_501_2056_0, i_13_501_2116_0, i_13_501_2136_0, i_13_501_2137_0,
    i_13_501_2172_0, i_13_501_2187_0, i_13_501_2224_0, i_13_501_2230_0,
    i_13_501_2311_0, i_13_501_2379_0, i_13_501_2394_0, i_13_501_2406_0,
    i_13_501_2425_0, i_13_501_2461_0, i_13_501_2502_0, i_13_501_2511_0,
    i_13_501_2664_0, i_13_501_2673_0, i_13_501_2691_0, i_13_501_2692_0,
    i_13_501_2715_0, i_13_501_2748_0, i_13_501_3024_0, i_13_501_3025_0,
    i_13_501_3114_0, i_13_501_3145_0, i_13_501_3153_0, i_13_501_3342_0,
    i_13_501_3369_0, i_13_501_3370_0, i_13_501_3373_0, i_13_501_3405_0,
    i_13_501_3412_0, i_13_501_3532_0, i_13_501_3579_0, i_13_501_3619_0,
    i_13_501_3871_0, i_13_501_3874_0, i_13_501_3987_0, i_13_501_3988_0,
    i_13_501_4032_0, i_13_501_4204_0, i_13_501_4305_0, i_13_501_4522_0,
    i_13_501_4524_0, i_13_501_4582_0, i_13_501_4590_0, i_13_501_4600_0,
    o_13_501_0_0  );
  input  i_13_501_31_0, i_13_501_36_0, i_13_501_37_0, i_13_501_102_0,
    i_13_501_255_0, i_13_501_262_0, i_13_501_264_0, i_13_501_265_0,
    i_13_501_282_0, i_13_501_492_0, i_13_501_505_0, i_13_501_532_0,
    i_13_501_535_0, i_13_501_577_0, i_13_501_616_0, i_13_501_651_0,
    i_13_501_675_0, i_13_501_676_0, i_13_501_723_0, i_13_501_777_0,
    i_13_501_810_0, i_13_501_837_0, i_13_501_838_0, i_13_501_871_0,
    i_13_501_948_0, i_13_501_949_0, i_13_501_981_0, i_13_501_1116_0,
    i_13_501_1197_0, i_13_501_1198_0, i_13_501_1212_0, i_13_501_1242_0,
    i_13_501_1269_0, i_13_501_1278_0, i_13_501_1324_0, i_13_501_1326_0,
    i_13_501_1380_0, i_13_501_1396_0, i_13_501_1446_0, i_13_501_1456_0,
    i_13_501_1504_0, i_13_501_1552_0, i_13_501_1746_0, i_13_501_1786_0,
    i_13_501_1803_0, i_13_501_1840_0, i_13_501_1857_0, i_13_501_1908_0,
    i_13_501_2010_0, i_13_501_2029_0, i_13_501_2046_0, i_13_501_2055_0,
    i_13_501_2056_0, i_13_501_2116_0, i_13_501_2136_0, i_13_501_2137_0,
    i_13_501_2172_0, i_13_501_2187_0, i_13_501_2224_0, i_13_501_2230_0,
    i_13_501_2311_0, i_13_501_2379_0, i_13_501_2394_0, i_13_501_2406_0,
    i_13_501_2425_0, i_13_501_2461_0, i_13_501_2502_0, i_13_501_2511_0,
    i_13_501_2664_0, i_13_501_2673_0, i_13_501_2691_0, i_13_501_2692_0,
    i_13_501_2715_0, i_13_501_2748_0, i_13_501_3024_0, i_13_501_3025_0,
    i_13_501_3114_0, i_13_501_3145_0, i_13_501_3153_0, i_13_501_3342_0,
    i_13_501_3369_0, i_13_501_3370_0, i_13_501_3373_0, i_13_501_3405_0,
    i_13_501_3412_0, i_13_501_3532_0, i_13_501_3579_0, i_13_501_3619_0,
    i_13_501_3871_0, i_13_501_3874_0, i_13_501_3987_0, i_13_501_3988_0,
    i_13_501_4032_0, i_13_501_4204_0, i_13_501_4305_0, i_13_501_4522_0,
    i_13_501_4524_0, i_13_501_4582_0, i_13_501_4590_0, i_13_501_4600_0;
  output o_13_501_0_0;
  assign o_13_501_0_0 = ~((i_13_501_948_0 & ((~i_13_501_2029_0 & i_13_501_3145_0 & ~i_13_501_3987_0) | (~i_13_501_3342_0 & ~i_13_501_3988_0 & ~i_13_501_4032_0))) | (~i_13_501_676_0 & ~i_13_501_1269_0 & ~i_13_501_2029_0 & ~i_13_501_2136_0) | (~i_13_501_2055_0 & ~i_13_501_2379_0 & ~i_13_501_2692_0) | (~i_13_501_837_0 & ~i_13_501_1552_0 & ~i_13_501_2406_0 & ~i_13_501_3145_0 & ~i_13_501_3988_0) | (i_13_501_492_0 & ~i_13_501_4305_0));
endmodule



// Benchmark "kernel_13_502" written by ABC on Sun Jul 19 10:52:19 2020

module kernel_13_502 ( 
    i_13_502_45_0, i_13_502_63_0, i_13_502_73_0, i_13_502_93_0,
    i_13_502_100_0, i_13_502_102_0, i_13_502_130_0, i_13_502_207_0,
    i_13_502_319_0, i_13_502_396_0, i_13_502_468_0, i_13_502_469_0,
    i_13_502_532_0, i_13_502_570_0, i_13_502_603_0, i_13_502_666_0,
    i_13_502_667_0, i_13_502_675_0, i_13_502_676_0, i_13_502_684_0,
    i_13_502_837_0, i_13_502_838_0, i_13_502_927_0, i_13_502_945_0,
    i_13_502_946_0, i_13_502_1024_0, i_13_502_1071_0, i_13_502_1098_0,
    i_13_502_1129_0, i_13_502_1144_0, i_13_502_1305_0, i_13_502_1306_0,
    i_13_502_1344_0, i_13_502_1399_0, i_13_502_1461_0, i_13_502_1503_0,
    i_13_502_1504_0, i_13_502_1593_0, i_13_502_1594_0, i_13_502_1620_0,
    i_13_502_1719_0, i_13_502_1720_0, i_13_502_1777_0, i_13_502_1791_0,
    i_13_502_1803_0, i_13_502_1804_0, i_13_502_1812_0, i_13_502_1837_0,
    i_13_502_1894_0, i_13_502_1908_0, i_13_502_1927_0, i_13_502_2016_0,
    i_13_502_2056_0, i_13_502_2137_0, i_13_502_2169_0, i_13_502_2197_0,
    i_13_502_2280_0, i_13_502_2344_0, i_13_502_2400_0, i_13_502_2431_0,
    i_13_502_2458_0, i_13_502_2479_0, i_13_502_2511_0, i_13_502_2547_0,
    i_13_502_2613_0, i_13_502_2614_0, i_13_502_2691_0, i_13_502_2692_0,
    i_13_502_2797_0, i_13_502_2820_0, i_13_502_2874_0, i_13_502_3019_0,
    i_13_502_3043_0, i_13_502_3088_0, i_13_502_3387_0, i_13_502_3423_0,
    i_13_502_3468_0, i_13_502_3475_0, i_13_502_3502_0, i_13_502_3531_0,
    i_13_502_3532_0, i_13_502_3618_0, i_13_502_3619_0, i_13_502_3687_0,
    i_13_502_3862_0, i_13_502_3934_0, i_13_502_3987_0, i_13_502_3988_0,
    i_13_502_4123_0, i_13_502_4260_0, i_13_502_4269_0, i_13_502_4311_0,
    i_13_502_4329_0, i_13_502_4392_0, i_13_502_4429_0, i_13_502_4446_0,
    i_13_502_4510_0, i_13_502_4518_0, i_13_502_4590_0, i_13_502_4600_0,
    o_13_502_0_0  );
  input  i_13_502_45_0, i_13_502_63_0, i_13_502_73_0, i_13_502_93_0,
    i_13_502_100_0, i_13_502_102_0, i_13_502_130_0, i_13_502_207_0,
    i_13_502_319_0, i_13_502_396_0, i_13_502_468_0, i_13_502_469_0,
    i_13_502_532_0, i_13_502_570_0, i_13_502_603_0, i_13_502_666_0,
    i_13_502_667_0, i_13_502_675_0, i_13_502_676_0, i_13_502_684_0,
    i_13_502_837_0, i_13_502_838_0, i_13_502_927_0, i_13_502_945_0,
    i_13_502_946_0, i_13_502_1024_0, i_13_502_1071_0, i_13_502_1098_0,
    i_13_502_1129_0, i_13_502_1144_0, i_13_502_1305_0, i_13_502_1306_0,
    i_13_502_1344_0, i_13_502_1399_0, i_13_502_1461_0, i_13_502_1503_0,
    i_13_502_1504_0, i_13_502_1593_0, i_13_502_1594_0, i_13_502_1620_0,
    i_13_502_1719_0, i_13_502_1720_0, i_13_502_1777_0, i_13_502_1791_0,
    i_13_502_1803_0, i_13_502_1804_0, i_13_502_1812_0, i_13_502_1837_0,
    i_13_502_1894_0, i_13_502_1908_0, i_13_502_1927_0, i_13_502_2016_0,
    i_13_502_2056_0, i_13_502_2137_0, i_13_502_2169_0, i_13_502_2197_0,
    i_13_502_2280_0, i_13_502_2344_0, i_13_502_2400_0, i_13_502_2431_0,
    i_13_502_2458_0, i_13_502_2479_0, i_13_502_2511_0, i_13_502_2547_0,
    i_13_502_2613_0, i_13_502_2614_0, i_13_502_2691_0, i_13_502_2692_0,
    i_13_502_2797_0, i_13_502_2820_0, i_13_502_2874_0, i_13_502_3019_0,
    i_13_502_3043_0, i_13_502_3088_0, i_13_502_3387_0, i_13_502_3423_0,
    i_13_502_3468_0, i_13_502_3475_0, i_13_502_3502_0, i_13_502_3531_0,
    i_13_502_3532_0, i_13_502_3618_0, i_13_502_3619_0, i_13_502_3687_0,
    i_13_502_3862_0, i_13_502_3934_0, i_13_502_3987_0, i_13_502_3988_0,
    i_13_502_4123_0, i_13_502_4260_0, i_13_502_4269_0, i_13_502_4311_0,
    i_13_502_4329_0, i_13_502_4392_0, i_13_502_4429_0, i_13_502_4446_0,
    i_13_502_4510_0, i_13_502_4518_0, i_13_502_4590_0, i_13_502_4600_0;
  output o_13_502_0_0;
  assign o_13_502_0_0 = ~((~i_13_502_1791_0 & ((~i_13_502_676_0 & ~i_13_502_2280_0 & ~i_13_502_3987_0) | (~i_13_502_675_0 & ~i_13_502_1071_0 & ~i_13_502_4429_0))) | ~i_13_502_838_0 | (~i_13_502_532_0 & ~i_13_502_1593_0));
endmodule



// Benchmark "kernel_13_503" written by ABC on Sun Jul 19 10:52:19 2020

module kernel_13_503 ( 
    i_13_503_92_0, i_13_503_139_0, i_13_503_176_0, i_13_503_184_0,
    i_13_503_185_0, i_13_503_193_0, i_13_503_364_0, i_13_503_407_0,
    i_13_503_482_0, i_13_503_589_0, i_13_503_604_0, i_13_503_607_0,
    i_13_503_608_0, i_13_503_658_0, i_13_503_659_0, i_13_503_661_0,
    i_13_503_662_0, i_13_503_686_0, i_13_503_712_0, i_13_503_814_0,
    i_13_503_851_0, i_13_503_859_0, i_13_503_868_0, i_13_503_949_0,
    i_13_503_956_0, i_13_503_982_0, i_13_503_1138_0, i_13_503_1148_0,
    i_13_503_1150_0, i_13_503_1210_0, i_13_503_1211_0, i_13_503_1226_0,
    i_13_503_1229_0, i_13_503_1244_0, i_13_503_1253_0, i_13_503_1301_0,
    i_13_503_1321_0, i_13_503_1487_0, i_13_503_1730_0, i_13_503_1765_0,
    i_13_503_1766_0, i_13_503_1804_0, i_13_503_1813_0, i_13_503_1829_0,
    i_13_503_1840_0, i_13_503_1892_0, i_13_503_1904_0, i_13_503_1961_0,
    i_13_503_2012_0, i_13_503_2020_0, i_13_503_2137_0, i_13_503_2182_0,
    i_13_503_2207_0, i_13_503_2281_0, i_13_503_2341_0, i_13_503_2435_0,
    i_13_503_2593_0, i_13_503_2857_0, i_13_503_2858_0, i_13_503_2938_0,
    i_13_503_2981_0, i_13_503_3047_0, i_13_503_3053_0, i_13_503_3110_0,
    i_13_503_3164_0, i_13_503_3254_0, i_13_503_3260_0, i_13_503_3268_0,
    i_13_503_3289_0, i_13_503_3349_0, i_13_503_3352_0, i_13_503_3442_0,
    i_13_503_3476_0, i_13_503_3484_0, i_13_503_3485_0, i_13_503_3491_0,
    i_13_503_3530_0, i_13_503_3547_0, i_13_503_3664_0, i_13_503_3667_0,
    i_13_503_3754_0, i_13_503_3764_0, i_13_503_3817_0, i_13_503_3821_0,
    i_13_503_3872_0, i_13_503_3875_0, i_13_503_3979_0, i_13_503_4006_0,
    i_13_503_4055_0, i_13_503_4160_0, i_13_503_4163_0, i_13_503_4249_0,
    i_13_503_4333_0, i_13_503_4358_0, i_13_503_4369_0, i_13_503_4370_0,
    i_13_503_4430_0, i_13_503_4537_0, i_13_503_4538_0, i_13_503_4565_0,
    o_13_503_0_0  );
  input  i_13_503_92_0, i_13_503_139_0, i_13_503_176_0, i_13_503_184_0,
    i_13_503_185_0, i_13_503_193_0, i_13_503_364_0, i_13_503_407_0,
    i_13_503_482_0, i_13_503_589_0, i_13_503_604_0, i_13_503_607_0,
    i_13_503_608_0, i_13_503_658_0, i_13_503_659_0, i_13_503_661_0,
    i_13_503_662_0, i_13_503_686_0, i_13_503_712_0, i_13_503_814_0,
    i_13_503_851_0, i_13_503_859_0, i_13_503_868_0, i_13_503_949_0,
    i_13_503_956_0, i_13_503_982_0, i_13_503_1138_0, i_13_503_1148_0,
    i_13_503_1150_0, i_13_503_1210_0, i_13_503_1211_0, i_13_503_1226_0,
    i_13_503_1229_0, i_13_503_1244_0, i_13_503_1253_0, i_13_503_1301_0,
    i_13_503_1321_0, i_13_503_1487_0, i_13_503_1730_0, i_13_503_1765_0,
    i_13_503_1766_0, i_13_503_1804_0, i_13_503_1813_0, i_13_503_1829_0,
    i_13_503_1840_0, i_13_503_1892_0, i_13_503_1904_0, i_13_503_1961_0,
    i_13_503_2012_0, i_13_503_2020_0, i_13_503_2137_0, i_13_503_2182_0,
    i_13_503_2207_0, i_13_503_2281_0, i_13_503_2341_0, i_13_503_2435_0,
    i_13_503_2593_0, i_13_503_2857_0, i_13_503_2858_0, i_13_503_2938_0,
    i_13_503_2981_0, i_13_503_3047_0, i_13_503_3053_0, i_13_503_3110_0,
    i_13_503_3164_0, i_13_503_3254_0, i_13_503_3260_0, i_13_503_3268_0,
    i_13_503_3289_0, i_13_503_3349_0, i_13_503_3352_0, i_13_503_3442_0,
    i_13_503_3476_0, i_13_503_3484_0, i_13_503_3485_0, i_13_503_3491_0,
    i_13_503_3530_0, i_13_503_3547_0, i_13_503_3664_0, i_13_503_3667_0,
    i_13_503_3754_0, i_13_503_3764_0, i_13_503_3817_0, i_13_503_3821_0,
    i_13_503_3872_0, i_13_503_3875_0, i_13_503_3979_0, i_13_503_4006_0,
    i_13_503_4055_0, i_13_503_4160_0, i_13_503_4163_0, i_13_503_4249_0,
    i_13_503_4333_0, i_13_503_4358_0, i_13_503_4369_0, i_13_503_4370_0,
    i_13_503_4430_0, i_13_503_4537_0, i_13_503_4538_0, i_13_503_4565_0;
  output o_13_503_0_0;
  assign o_13_503_0_0 = ~((~i_13_503_4163_0 & (i_13_503_1210_0 | ~i_13_503_3530_0)) | ~i_13_503_1148_0 | (~i_13_503_3484_0 & ~i_13_503_4565_0));
endmodule



// Benchmark "kernel_13_504" written by ABC on Sun Jul 19 10:52:20 2020

module kernel_13_504 ( 
    i_13_504_34_0, i_13_504_44_0, i_13_504_67_0, i_13_504_70_0,
    i_13_504_94_0, i_13_504_95_0, i_13_504_418_0, i_13_504_435_0,
    i_13_504_447_0, i_13_504_449_0, i_13_504_592_0, i_13_504_593_0,
    i_13_504_607_0, i_13_504_665_0, i_13_504_679_0, i_13_504_681_0,
    i_13_504_698_0, i_13_504_763_0, i_13_504_764_0, i_13_504_1048_0,
    i_13_504_1075_0, i_13_504_1103_0, i_13_504_1106_0, i_13_504_1123_0,
    i_13_504_1131_0, i_13_504_1132_0, i_13_504_1213_0, i_13_504_1273_0,
    i_13_504_1312_0, i_13_504_1321_0, i_13_504_1349_0, i_13_504_1428_0,
    i_13_504_1544_0, i_13_504_1605_0, i_13_504_1606_0, i_13_504_1644_0,
    i_13_504_1672_0, i_13_504_1753_0, i_13_504_1780_0, i_13_504_1786_0,
    i_13_504_1796_0, i_13_504_1797_0, i_13_504_1798_0, i_13_504_1888_0,
    i_13_504_2004_0, i_13_504_2024_0, i_13_504_2120_0, i_13_504_2173_0,
    i_13_504_2382_0, i_13_504_2383_0, i_13_504_2455_0, i_13_504_2464_0,
    i_13_504_2570_0, i_13_504_2600_0, i_13_504_2679_0, i_13_504_2680_0,
    i_13_504_2725_0, i_13_504_2850_0, i_13_504_2851_0, i_13_504_2852_0,
    i_13_504_3003_0, i_13_504_3032_0, i_13_504_3076_0, i_13_504_3094_0,
    i_13_504_3163_0, i_13_504_3166_0, i_13_504_3265_0, i_13_504_3273_0,
    i_13_504_3311_0, i_13_504_3370_0, i_13_504_3391_0, i_13_504_3540_0,
    i_13_504_3541_0, i_13_504_3543_0, i_13_504_3545_0, i_13_504_3560_0,
    i_13_504_3651_0, i_13_504_3722_0, i_13_504_3741_0, i_13_504_3742_0,
    i_13_504_3757_0, i_13_504_3806_0, i_13_504_3900_0, i_13_504_3918_0,
    i_13_504_3940_0, i_13_504_4040_0, i_13_504_4083_0, i_13_504_4099_0,
    i_13_504_4297_0, i_13_504_4345_0, i_13_504_4381_0, i_13_504_4399_0,
    i_13_504_4417_0, i_13_504_4433_0, i_13_504_4561_0, i_13_504_4594_0,
    i_13_504_4595_0, i_13_504_4597_0, i_13_504_4598_0, i_13_504_4607_0,
    o_13_504_0_0  );
  input  i_13_504_34_0, i_13_504_44_0, i_13_504_67_0, i_13_504_70_0,
    i_13_504_94_0, i_13_504_95_0, i_13_504_418_0, i_13_504_435_0,
    i_13_504_447_0, i_13_504_449_0, i_13_504_592_0, i_13_504_593_0,
    i_13_504_607_0, i_13_504_665_0, i_13_504_679_0, i_13_504_681_0,
    i_13_504_698_0, i_13_504_763_0, i_13_504_764_0, i_13_504_1048_0,
    i_13_504_1075_0, i_13_504_1103_0, i_13_504_1106_0, i_13_504_1123_0,
    i_13_504_1131_0, i_13_504_1132_0, i_13_504_1213_0, i_13_504_1273_0,
    i_13_504_1312_0, i_13_504_1321_0, i_13_504_1349_0, i_13_504_1428_0,
    i_13_504_1544_0, i_13_504_1605_0, i_13_504_1606_0, i_13_504_1644_0,
    i_13_504_1672_0, i_13_504_1753_0, i_13_504_1780_0, i_13_504_1786_0,
    i_13_504_1796_0, i_13_504_1797_0, i_13_504_1798_0, i_13_504_1888_0,
    i_13_504_2004_0, i_13_504_2024_0, i_13_504_2120_0, i_13_504_2173_0,
    i_13_504_2382_0, i_13_504_2383_0, i_13_504_2455_0, i_13_504_2464_0,
    i_13_504_2570_0, i_13_504_2600_0, i_13_504_2679_0, i_13_504_2680_0,
    i_13_504_2725_0, i_13_504_2850_0, i_13_504_2851_0, i_13_504_2852_0,
    i_13_504_3003_0, i_13_504_3032_0, i_13_504_3076_0, i_13_504_3094_0,
    i_13_504_3163_0, i_13_504_3166_0, i_13_504_3265_0, i_13_504_3273_0,
    i_13_504_3311_0, i_13_504_3370_0, i_13_504_3391_0, i_13_504_3540_0,
    i_13_504_3541_0, i_13_504_3543_0, i_13_504_3545_0, i_13_504_3560_0,
    i_13_504_3651_0, i_13_504_3722_0, i_13_504_3741_0, i_13_504_3742_0,
    i_13_504_3757_0, i_13_504_3806_0, i_13_504_3900_0, i_13_504_3918_0,
    i_13_504_3940_0, i_13_504_4040_0, i_13_504_4083_0, i_13_504_4099_0,
    i_13_504_4297_0, i_13_504_4345_0, i_13_504_4381_0, i_13_504_4399_0,
    i_13_504_4417_0, i_13_504_4433_0, i_13_504_4561_0, i_13_504_4594_0,
    i_13_504_4595_0, i_13_504_4597_0, i_13_504_4598_0, i_13_504_4607_0;
  output o_13_504_0_0;
  assign o_13_504_0_0 = ~((~i_13_504_2680_0 & (i_13_504_94_0 | (~i_13_504_418_0 & ~i_13_504_3918_0))) | (~i_13_504_681_0 & ~i_13_504_1075_0 & ~i_13_504_1213_0 & ~i_13_504_3540_0) | (i_13_504_3545_0 & ~i_13_504_4040_0) | (~i_13_504_1798_0 & ~i_13_504_2383_0 & ~i_13_504_4083_0 & ~i_13_504_4381_0));
endmodule



// Benchmark "kernel_13_505" written by ABC on Sun Jul 19 10:52:21 2020

module kernel_13_505 ( 
    i_13_505_32_0, i_13_505_91_0, i_13_505_92_0, i_13_505_281_0,
    i_13_505_307_0, i_13_505_308_0, i_13_505_317_0, i_13_505_361_0,
    i_13_505_367_0, i_13_505_383_0, i_13_505_384_0, i_13_505_528_0,
    i_13_505_535_0, i_13_505_551_0, i_13_505_569_0, i_13_505_584_0,
    i_13_505_604_0, i_13_505_626_0, i_13_505_643_0, i_13_505_686_0,
    i_13_505_688_0, i_13_505_704_0, i_13_505_724_0, i_13_505_796_0,
    i_13_505_815_0, i_13_505_949_0, i_13_505_1067_0, i_13_505_1111_0,
    i_13_505_1216_0, i_13_505_1217_0, i_13_505_1219_0, i_13_505_1255_0,
    i_13_505_1321_0, i_13_505_1402_0, i_13_505_1432_0, i_13_505_1443_0,
    i_13_505_1471_0, i_13_505_1487_0, i_13_505_1552_0, i_13_505_1597_0,
    i_13_505_1635_0, i_13_505_1644_0, i_13_505_1657_0, i_13_505_1705_0,
    i_13_505_1721_0, i_13_505_1837_0, i_13_505_1900_0, i_13_505_1910_0,
    i_13_505_1922_0, i_13_505_1931_0, i_13_505_1999_0, i_13_505_2000_0,
    i_13_505_2002_0, i_13_505_2006_0, i_13_505_2056_0, i_13_505_2057_0,
    i_13_505_2173_0, i_13_505_2176_0, i_13_505_2231_0, i_13_505_2422_0,
    i_13_505_2423_0, i_13_505_2424_0, i_13_505_2452_0, i_13_505_2678_0,
    i_13_505_2767_0, i_13_505_2965_0, i_13_505_3039_0, i_13_505_3056_0,
    i_13_505_3064_0, i_13_505_3065_0, i_13_505_3127_0, i_13_505_3142_0,
    i_13_505_3145_0, i_13_505_3218_0, i_13_505_3372_0, i_13_505_3379_0,
    i_13_505_3415_0, i_13_505_3487_0, i_13_505_3524_0, i_13_505_3541_0,
    i_13_505_3700_0, i_13_505_3712_0, i_13_505_3794_0, i_13_505_3865_0,
    i_13_505_3871_0, i_13_505_4018_0, i_13_505_4037_0, i_13_505_4082_0,
    i_13_505_4118_0, i_13_505_4150_0, i_13_505_4217_0, i_13_505_4279_0,
    i_13_505_4306_0, i_13_505_4307_0, i_13_505_4339_0, i_13_505_4342_0,
    i_13_505_4350_0, i_13_505_4351_0, i_13_505_4397_0, i_13_505_4415_0,
    o_13_505_0_0  );
  input  i_13_505_32_0, i_13_505_91_0, i_13_505_92_0, i_13_505_281_0,
    i_13_505_307_0, i_13_505_308_0, i_13_505_317_0, i_13_505_361_0,
    i_13_505_367_0, i_13_505_383_0, i_13_505_384_0, i_13_505_528_0,
    i_13_505_535_0, i_13_505_551_0, i_13_505_569_0, i_13_505_584_0,
    i_13_505_604_0, i_13_505_626_0, i_13_505_643_0, i_13_505_686_0,
    i_13_505_688_0, i_13_505_704_0, i_13_505_724_0, i_13_505_796_0,
    i_13_505_815_0, i_13_505_949_0, i_13_505_1067_0, i_13_505_1111_0,
    i_13_505_1216_0, i_13_505_1217_0, i_13_505_1219_0, i_13_505_1255_0,
    i_13_505_1321_0, i_13_505_1402_0, i_13_505_1432_0, i_13_505_1443_0,
    i_13_505_1471_0, i_13_505_1487_0, i_13_505_1552_0, i_13_505_1597_0,
    i_13_505_1635_0, i_13_505_1644_0, i_13_505_1657_0, i_13_505_1705_0,
    i_13_505_1721_0, i_13_505_1837_0, i_13_505_1900_0, i_13_505_1910_0,
    i_13_505_1922_0, i_13_505_1931_0, i_13_505_1999_0, i_13_505_2000_0,
    i_13_505_2002_0, i_13_505_2006_0, i_13_505_2056_0, i_13_505_2057_0,
    i_13_505_2173_0, i_13_505_2176_0, i_13_505_2231_0, i_13_505_2422_0,
    i_13_505_2423_0, i_13_505_2424_0, i_13_505_2452_0, i_13_505_2678_0,
    i_13_505_2767_0, i_13_505_2965_0, i_13_505_3039_0, i_13_505_3056_0,
    i_13_505_3064_0, i_13_505_3065_0, i_13_505_3127_0, i_13_505_3142_0,
    i_13_505_3145_0, i_13_505_3218_0, i_13_505_3372_0, i_13_505_3379_0,
    i_13_505_3415_0, i_13_505_3487_0, i_13_505_3524_0, i_13_505_3541_0,
    i_13_505_3700_0, i_13_505_3712_0, i_13_505_3794_0, i_13_505_3865_0,
    i_13_505_3871_0, i_13_505_4018_0, i_13_505_4037_0, i_13_505_4082_0,
    i_13_505_4118_0, i_13_505_4150_0, i_13_505_4217_0, i_13_505_4279_0,
    i_13_505_4306_0, i_13_505_4307_0, i_13_505_4339_0, i_13_505_4342_0,
    i_13_505_4350_0, i_13_505_4351_0, i_13_505_4397_0, i_13_505_4415_0;
  output o_13_505_0_0;
  assign o_13_505_0_0 = ~((~i_13_505_4415_0 & (~i_13_505_3064_0 | (~i_13_505_535_0 & ~i_13_505_2231_0))) | i_13_505_2452_0 | (~i_13_505_1217_0 & ~i_13_505_3065_0) | ~i_13_505_4082_0 | (~i_13_505_688_0 & ~i_13_505_2006_0 & ~i_13_505_4150_0) | (~i_13_505_3145_0 & i_13_505_4351_0));
endmodule



// Benchmark "kernel_13_506" written by ABC on Sun Jul 19 10:52:22 2020

module kernel_13_506 ( 
    i_13_506_31_0, i_13_506_32_0, i_13_506_46_0, i_13_506_67_0,
    i_13_506_77_0, i_13_506_92_0, i_13_506_110_0, i_13_506_118_0,
    i_13_506_119_0, i_13_506_136_0, i_13_506_229_0, i_13_506_334_0,
    i_13_506_490_0, i_13_506_535_0, i_13_506_562_0, i_13_506_563_0,
    i_13_506_604_0, i_13_506_605_0, i_13_506_730_0, i_13_506_760_0,
    i_13_506_947_0, i_13_506_1084_0, i_13_506_1210_0, i_13_506_1216_0,
    i_13_506_1217_0, i_13_506_1315_0, i_13_506_1441_0, i_13_506_1442_0,
    i_13_506_1471_0, i_13_506_1486_0, i_13_506_1487_0, i_13_506_1507_0,
    i_13_506_1589_0, i_13_506_1606_0, i_13_506_1625_0, i_13_506_1633_0,
    i_13_506_1659_0, i_13_506_1678_0, i_13_506_1694_0, i_13_506_1731_0,
    i_13_506_1733_0, i_13_506_1787_0, i_13_506_1837_0, i_13_506_1840_0,
    i_13_506_1841_0, i_13_506_1886_0, i_13_506_1930_0, i_13_506_1931_0,
    i_13_506_1937_0, i_13_506_2000_0, i_13_506_2128_0, i_13_506_2173_0,
    i_13_506_2264_0, i_13_506_2362_0, i_13_506_2422_0, i_13_506_2423_0,
    i_13_506_2425_0, i_13_506_2426_0, i_13_506_2432_0, i_13_506_2452_0,
    i_13_506_2498_0, i_13_506_2747_0, i_13_506_3020_0, i_13_506_3035_0,
    i_13_506_3044_0, i_13_506_3100_0, i_13_506_3101_0, i_13_506_3127_0,
    i_13_506_3161_0, i_13_506_3214_0, i_13_506_3227_0, i_13_506_3375_0,
    i_13_506_3459_0, i_13_506_3461_0, i_13_506_3488_0, i_13_506_3577_0,
    i_13_506_3613_0, i_13_506_3700_0, i_13_506_3703_0, i_13_506_3756_0,
    i_13_506_3764_0, i_13_506_3784_0, i_13_506_3794_0, i_13_506_3844_0,
    i_13_506_3871_0, i_13_506_3872_0, i_13_506_4007_0, i_13_506_4081_0,
    i_13_506_4105_0, i_13_506_4117_0, i_13_506_4118_0, i_13_506_4159_0,
    i_13_506_4160_0, i_13_506_4163_0, i_13_506_4172_0, i_13_506_4295_0,
    i_13_506_4325_0, i_13_506_4348_0, i_13_506_4349_0, i_13_506_4474_0,
    o_13_506_0_0  );
  input  i_13_506_31_0, i_13_506_32_0, i_13_506_46_0, i_13_506_67_0,
    i_13_506_77_0, i_13_506_92_0, i_13_506_110_0, i_13_506_118_0,
    i_13_506_119_0, i_13_506_136_0, i_13_506_229_0, i_13_506_334_0,
    i_13_506_490_0, i_13_506_535_0, i_13_506_562_0, i_13_506_563_0,
    i_13_506_604_0, i_13_506_605_0, i_13_506_730_0, i_13_506_760_0,
    i_13_506_947_0, i_13_506_1084_0, i_13_506_1210_0, i_13_506_1216_0,
    i_13_506_1217_0, i_13_506_1315_0, i_13_506_1441_0, i_13_506_1442_0,
    i_13_506_1471_0, i_13_506_1486_0, i_13_506_1487_0, i_13_506_1507_0,
    i_13_506_1589_0, i_13_506_1606_0, i_13_506_1625_0, i_13_506_1633_0,
    i_13_506_1659_0, i_13_506_1678_0, i_13_506_1694_0, i_13_506_1731_0,
    i_13_506_1733_0, i_13_506_1787_0, i_13_506_1837_0, i_13_506_1840_0,
    i_13_506_1841_0, i_13_506_1886_0, i_13_506_1930_0, i_13_506_1931_0,
    i_13_506_1937_0, i_13_506_2000_0, i_13_506_2128_0, i_13_506_2173_0,
    i_13_506_2264_0, i_13_506_2362_0, i_13_506_2422_0, i_13_506_2423_0,
    i_13_506_2425_0, i_13_506_2426_0, i_13_506_2432_0, i_13_506_2452_0,
    i_13_506_2498_0, i_13_506_2747_0, i_13_506_3020_0, i_13_506_3035_0,
    i_13_506_3044_0, i_13_506_3100_0, i_13_506_3101_0, i_13_506_3127_0,
    i_13_506_3161_0, i_13_506_3214_0, i_13_506_3227_0, i_13_506_3375_0,
    i_13_506_3459_0, i_13_506_3461_0, i_13_506_3488_0, i_13_506_3577_0,
    i_13_506_3613_0, i_13_506_3700_0, i_13_506_3703_0, i_13_506_3756_0,
    i_13_506_3764_0, i_13_506_3784_0, i_13_506_3794_0, i_13_506_3844_0,
    i_13_506_3871_0, i_13_506_3872_0, i_13_506_4007_0, i_13_506_4081_0,
    i_13_506_4105_0, i_13_506_4117_0, i_13_506_4118_0, i_13_506_4159_0,
    i_13_506_4160_0, i_13_506_4163_0, i_13_506_4172_0, i_13_506_4295_0,
    i_13_506_4325_0, i_13_506_4348_0, i_13_506_4349_0, i_13_506_4474_0;
  output o_13_506_0_0;
  assign o_13_506_0_0 = ~(~i_13_506_3101_0 | (~i_13_506_1217_0 & i_13_506_3784_0) | (~i_13_506_1487_0 & ~i_13_506_2423_0) | (~i_13_506_92_0 & ~i_13_506_2422_0));
endmodule



// Benchmark "kernel_13_507" written by ABC on Sun Jul 19 10:52:23 2020

module kernel_13_507 ( 
    i_13_507_46_0, i_13_507_102_0, i_13_507_163_0, i_13_507_312_0,
    i_13_507_321_0, i_13_507_322_0, i_13_507_342_0, i_13_507_379_0,
    i_13_507_408_0, i_13_507_442_0, i_13_507_604_0, i_13_507_624_0,
    i_13_507_625_0, i_13_507_657_0, i_13_507_671_0, i_13_507_680_0,
    i_13_507_757_0, i_13_507_846_0, i_13_507_883_0, i_13_507_885_0,
    i_13_507_936_0, i_13_507_1018_0, i_13_507_1147_0, i_13_507_1266_0,
    i_13_507_1362_0, i_13_507_1434_0, i_13_507_1498_0, i_13_507_1513_0,
    i_13_507_1515_0, i_13_507_1563_0, i_13_507_1582_0, i_13_507_1593_0,
    i_13_507_1594_0, i_13_507_1605_0, i_13_507_1701_0, i_13_507_1828_0,
    i_13_507_1944_0, i_13_507_2002_0, i_13_507_2012_0, i_13_507_2019_0,
    i_13_507_2025_0, i_13_507_2248_0, i_13_507_2268_0, i_13_507_2296_0,
    i_13_507_2463_0, i_13_507_2469_0, i_13_507_2498_0, i_13_507_2524_0,
    i_13_507_2601_0, i_13_507_2606_0, i_13_507_2673_0, i_13_507_2917_0,
    i_13_507_2966_0, i_13_507_2968_0, i_13_507_3003_0, i_13_507_3007_0,
    i_13_507_3030_0, i_13_507_3032_0, i_13_507_3099_0, i_13_507_3105_0,
    i_13_507_3214_0, i_13_507_3261_0, i_13_507_3325_0, i_13_507_3352_0,
    i_13_507_3400_0, i_13_507_3452_0, i_13_507_3483_0, i_13_507_3484_0,
    i_13_507_3541_0, i_13_507_3549_0, i_13_507_3566_0, i_13_507_3575_0,
    i_13_507_3699_0, i_13_507_3717_0, i_13_507_3730_0, i_13_507_3763_0,
    i_13_507_3765_0, i_13_507_3781_0, i_13_507_3784_0, i_13_507_3819_0,
    i_13_507_3823_0, i_13_507_3861_0, i_13_507_3898_0, i_13_507_3910_0,
    i_13_507_3970_0, i_13_507_4116_0, i_13_507_4159_0, i_13_507_4321_0,
    i_13_507_4335_0, i_13_507_4365_0, i_13_507_4366_0, i_13_507_4422_0,
    i_13_507_4448_0, i_13_507_4537_0, i_13_507_4558_0, i_13_507_4563_0,
    i_13_507_4564_0, i_13_507_4565_0, i_13_507_4599_0, i_13_507_4607_0,
    o_13_507_0_0  );
  input  i_13_507_46_0, i_13_507_102_0, i_13_507_163_0, i_13_507_312_0,
    i_13_507_321_0, i_13_507_322_0, i_13_507_342_0, i_13_507_379_0,
    i_13_507_408_0, i_13_507_442_0, i_13_507_604_0, i_13_507_624_0,
    i_13_507_625_0, i_13_507_657_0, i_13_507_671_0, i_13_507_680_0,
    i_13_507_757_0, i_13_507_846_0, i_13_507_883_0, i_13_507_885_0,
    i_13_507_936_0, i_13_507_1018_0, i_13_507_1147_0, i_13_507_1266_0,
    i_13_507_1362_0, i_13_507_1434_0, i_13_507_1498_0, i_13_507_1513_0,
    i_13_507_1515_0, i_13_507_1563_0, i_13_507_1582_0, i_13_507_1593_0,
    i_13_507_1594_0, i_13_507_1605_0, i_13_507_1701_0, i_13_507_1828_0,
    i_13_507_1944_0, i_13_507_2002_0, i_13_507_2012_0, i_13_507_2019_0,
    i_13_507_2025_0, i_13_507_2248_0, i_13_507_2268_0, i_13_507_2296_0,
    i_13_507_2463_0, i_13_507_2469_0, i_13_507_2498_0, i_13_507_2524_0,
    i_13_507_2601_0, i_13_507_2606_0, i_13_507_2673_0, i_13_507_2917_0,
    i_13_507_2966_0, i_13_507_2968_0, i_13_507_3003_0, i_13_507_3007_0,
    i_13_507_3030_0, i_13_507_3032_0, i_13_507_3099_0, i_13_507_3105_0,
    i_13_507_3214_0, i_13_507_3261_0, i_13_507_3325_0, i_13_507_3352_0,
    i_13_507_3400_0, i_13_507_3452_0, i_13_507_3483_0, i_13_507_3484_0,
    i_13_507_3541_0, i_13_507_3549_0, i_13_507_3566_0, i_13_507_3575_0,
    i_13_507_3699_0, i_13_507_3717_0, i_13_507_3730_0, i_13_507_3763_0,
    i_13_507_3765_0, i_13_507_3781_0, i_13_507_3784_0, i_13_507_3819_0,
    i_13_507_3823_0, i_13_507_3861_0, i_13_507_3898_0, i_13_507_3910_0,
    i_13_507_3970_0, i_13_507_4116_0, i_13_507_4159_0, i_13_507_4321_0,
    i_13_507_4335_0, i_13_507_4365_0, i_13_507_4366_0, i_13_507_4422_0,
    i_13_507_4448_0, i_13_507_4537_0, i_13_507_4558_0, i_13_507_4563_0,
    i_13_507_4564_0, i_13_507_4565_0, i_13_507_4599_0, i_13_507_4607_0;
  output o_13_507_0_0;
  assign o_13_507_0_0 = ~((~i_13_507_3549_0 & (~i_13_507_4159_0 | (i_13_507_1594_0 & ~i_13_507_3898_0))) | (i_13_507_1266_0 & i_13_507_3730_0) | (~i_13_507_885_0 & ~i_13_507_1498_0 & i_13_507_3765_0) | (~i_13_507_1944_0 & i_13_507_3105_0 & ~i_13_507_3819_0 & ~i_13_507_3898_0) | (i_13_507_3784_0 & ~i_13_507_4321_0) | (~i_13_507_3261_0 & ~i_13_507_4565_0));
endmodule



// Benchmark "kernel_13_508" written by ABC on Sun Jul 19 10:52:23 2020

module kernel_13_508 ( 
    i_13_508_98_0, i_13_508_107_0, i_13_508_108_0, i_13_508_112_0,
    i_13_508_113_0, i_13_508_116_0, i_13_508_125_0, i_13_508_211_0,
    i_13_508_265_0, i_13_508_283_0, i_13_508_310_0, i_13_508_368_0,
    i_13_508_558_0, i_13_508_589_0, i_13_508_662_0, i_13_508_746_0,
    i_13_508_814_0, i_13_508_859_0, i_13_508_949_0, i_13_508_1017_0,
    i_13_508_1087_0, i_13_508_1088_0, i_13_508_1144_0, i_13_508_1219_0,
    i_13_508_1220_0, i_13_508_1474_0, i_13_508_1490_0, i_13_508_1520_0,
    i_13_508_1570_0, i_13_508_1574_0, i_13_508_1789_0, i_13_508_1790_0,
    i_13_508_1804_0, i_13_508_1841_0, i_13_508_1844_0, i_13_508_1915_0,
    i_13_508_1934_0, i_13_508_1993_0, i_13_508_2023_0, i_13_508_2173_0,
    i_13_508_2177_0, i_13_508_2276_0, i_13_508_2348_0, i_13_508_2421_0,
    i_13_508_2425_0, i_13_508_2434_0, i_13_508_2435_0, i_13_508_2438_0,
    i_13_508_2501_0, i_13_508_2542_0, i_13_508_2543_0, i_13_508_2561_0,
    i_13_508_2713_0, i_13_508_2716_0, i_13_508_2717_0, i_13_508_3047_0,
    i_13_508_3099_0, i_13_508_3146_0, i_13_508_3148_0, i_13_508_3149_0,
    i_13_508_3164_0, i_13_508_3167_0, i_13_508_3254_0, i_13_508_3344_0,
    i_13_508_3388_0, i_13_508_3413_0, i_13_508_3418_0, i_13_508_3419_0,
    i_13_508_3454_0, i_13_508_3455_0, i_13_508_3526_0, i_13_508_3527_0,
    i_13_508_3545_0, i_13_508_3640_0, i_13_508_3738_0, i_13_508_3742_0,
    i_13_508_3752_0, i_13_508_3766_0, i_13_508_3874_0, i_13_508_3875_0,
    i_13_508_3938_0, i_13_508_3994_0, i_13_508_4048_0, i_13_508_4077_0,
    i_13_508_4121_0, i_13_508_4163_0, i_13_508_4234_0, i_13_508_4252_0,
    i_13_508_4255_0, i_13_508_4264_0, i_13_508_4271_0, i_13_508_4309_0,
    i_13_508_4316_0, i_13_508_4328_0, i_13_508_4343_0, i_13_508_4354_0,
    i_13_508_4418_0, i_13_508_4518_0, i_13_508_4543_0, i_13_508_4544_0,
    o_13_508_0_0  );
  input  i_13_508_98_0, i_13_508_107_0, i_13_508_108_0, i_13_508_112_0,
    i_13_508_113_0, i_13_508_116_0, i_13_508_125_0, i_13_508_211_0,
    i_13_508_265_0, i_13_508_283_0, i_13_508_310_0, i_13_508_368_0,
    i_13_508_558_0, i_13_508_589_0, i_13_508_662_0, i_13_508_746_0,
    i_13_508_814_0, i_13_508_859_0, i_13_508_949_0, i_13_508_1017_0,
    i_13_508_1087_0, i_13_508_1088_0, i_13_508_1144_0, i_13_508_1219_0,
    i_13_508_1220_0, i_13_508_1474_0, i_13_508_1490_0, i_13_508_1520_0,
    i_13_508_1570_0, i_13_508_1574_0, i_13_508_1789_0, i_13_508_1790_0,
    i_13_508_1804_0, i_13_508_1841_0, i_13_508_1844_0, i_13_508_1915_0,
    i_13_508_1934_0, i_13_508_1993_0, i_13_508_2023_0, i_13_508_2173_0,
    i_13_508_2177_0, i_13_508_2276_0, i_13_508_2348_0, i_13_508_2421_0,
    i_13_508_2425_0, i_13_508_2434_0, i_13_508_2435_0, i_13_508_2438_0,
    i_13_508_2501_0, i_13_508_2542_0, i_13_508_2543_0, i_13_508_2561_0,
    i_13_508_2713_0, i_13_508_2716_0, i_13_508_2717_0, i_13_508_3047_0,
    i_13_508_3099_0, i_13_508_3146_0, i_13_508_3148_0, i_13_508_3149_0,
    i_13_508_3164_0, i_13_508_3167_0, i_13_508_3254_0, i_13_508_3344_0,
    i_13_508_3388_0, i_13_508_3413_0, i_13_508_3418_0, i_13_508_3419_0,
    i_13_508_3454_0, i_13_508_3455_0, i_13_508_3526_0, i_13_508_3527_0,
    i_13_508_3545_0, i_13_508_3640_0, i_13_508_3738_0, i_13_508_3742_0,
    i_13_508_3752_0, i_13_508_3766_0, i_13_508_3874_0, i_13_508_3875_0,
    i_13_508_3938_0, i_13_508_3994_0, i_13_508_4048_0, i_13_508_4077_0,
    i_13_508_4121_0, i_13_508_4163_0, i_13_508_4234_0, i_13_508_4252_0,
    i_13_508_4255_0, i_13_508_4264_0, i_13_508_4271_0, i_13_508_4309_0,
    i_13_508_4316_0, i_13_508_4328_0, i_13_508_4343_0, i_13_508_4354_0,
    i_13_508_4418_0, i_13_508_4518_0, i_13_508_4543_0, i_13_508_4544_0;
  output o_13_508_0_0;
  assign o_13_508_0_0 = ~(~i_13_508_1088_0 | ~i_13_508_4328_0);
endmodule



// Benchmark "kernel_13_509" written by ABC on Sun Jul 19 10:52:24 2020

module kernel_13_509 ( 
    i_13_509_31_0, i_13_509_32_0, i_13_509_35_0, i_13_509_94_0,
    i_13_509_95_0, i_13_509_97_0, i_13_509_98_0, i_13_509_113_0,
    i_13_509_115_0, i_13_509_116_0, i_13_509_121_0, i_13_509_122_0,
    i_13_509_178_0, i_13_509_229_0, i_13_509_232_0, i_13_509_260_0,
    i_13_509_313_0, i_13_509_386_0, i_13_509_448_0, i_13_509_449_0,
    i_13_509_538_0, i_13_509_539_0, i_13_509_565_0, i_13_509_607_0,
    i_13_509_730_0, i_13_509_733_0, i_13_509_800_0, i_13_509_868_0,
    i_13_509_943_0, i_13_509_953_0, i_13_509_1123_0, i_13_509_1193_0,
    i_13_509_1219_0, i_13_509_1313_0, i_13_509_1409_0, i_13_509_1440_0,
    i_13_509_1444_0, i_13_509_1445_0, i_13_509_1448_0, i_13_509_1628_0,
    i_13_509_1631_0, i_13_509_1787_0, i_13_509_1788_0, i_13_509_1799_0,
    i_13_509_1840_0, i_13_509_1841_0, i_13_509_1843_0, i_13_509_1844_0,
    i_13_509_1846_0, i_13_509_1912_0, i_13_509_1940_0, i_13_509_1943_0,
    i_13_509_2005_0, i_13_509_2021_0, i_13_509_2173_0, i_13_509_2176_0,
    i_13_509_2177_0, i_13_509_2279_0, i_13_509_2422_0, i_13_509_2425_0,
    i_13_509_2426_0, i_13_509_2428_0, i_13_509_2429_0, i_13_509_2447_0,
    i_13_509_2617_0, i_13_509_2677_0, i_13_509_2680_0, i_13_509_2681_0,
    i_13_509_2740_0, i_13_509_2749_0, i_13_509_2923_0, i_13_509_3002_0,
    i_13_509_3023_0, i_13_509_3037_0, i_13_509_3038_0, i_13_509_3064_0,
    i_13_509_3068_0, i_13_509_3146_0, i_13_509_3163_0, i_13_509_3164_0,
    i_13_509_3418_0, i_13_509_3419_0, i_13_509_3424_0, i_13_509_3425_0,
    i_13_509_3427_0, i_13_509_3428_0, i_13_509_3460_0, i_13_509_3487_0,
    i_13_509_3505_0, i_13_509_3580_0, i_13_509_3700_0, i_13_509_3865_0,
    i_13_509_3874_0, i_13_509_3875_0, i_13_509_4085_0, i_13_509_4351_0,
    i_13_509_4352_0, i_13_509_4453_0, i_13_509_4594_0, i_13_509_4598_0,
    o_13_509_0_0  );
  input  i_13_509_31_0, i_13_509_32_0, i_13_509_35_0, i_13_509_94_0,
    i_13_509_95_0, i_13_509_97_0, i_13_509_98_0, i_13_509_113_0,
    i_13_509_115_0, i_13_509_116_0, i_13_509_121_0, i_13_509_122_0,
    i_13_509_178_0, i_13_509_229_0, i_13_509_232_0, i_13_509_260_0,
    i_13_509_313_0, i_13_509_386_0, i_13_509_448_0, i_13_509_449_0,
    i_13_509_538_0, i_13_509_539_0, i_13_509_565_0, i_13_509_607_0,
    i_13_509_730_0, i_13_509_733_0, i_13_509_800_0, i_13_509_868_0,
    i_13_509_943_0, i_13_509_953_0, i_13_509_1123_0, i_13_509_1193_0,
    i_13_509_1219_0, i_13_509_1313_0, i_13_509_1409_0, i_13_509_1440_0,
    i_13_509_1444_0, i_13_509_1445_0, i_13_509_1448_0, i_13_509_1628_0,
    i_13_509_1631_0, i_13_509_1787_0, i_13_509_1788_0, i_13_509_1799_0,
    i_13_509_1840_0, i_13_509_1841_0, i_13_509_1843_0, i_13_509_1844_0,
    i_13_509_1846_0, i_13_509_1912_0, i_13_509_1940_0, i_13_509_1943_0,
    i_13_509_2005_0, i_13_509_2021_0, i_13_509_2173_0, i_13_509_2176_0,
    i_13_509_2177_0, i_13_509_2279_0, i_13_509_2422_0, i_13_509_2425_0,
    i_13_509_2426_0, i_13_509_2428_0, i_13_509_2429_0, i_13_509_2447_0,
    i_13_509_2617_0, i_13_509_2677_0, i_13_509_2680_0, i_13_509_2681_0,
    i_13_509_2740_0, i_13_509_2749_0, i_13_509_2923_0, i_13_509_3002_0,
    i_13_509_3023_0, i_13_509_3037_0, i_13_509_3038_0, i_13_509_3064_0,
    i_13_509_3068_0, i_13_509_3146_0, i_13_509_3163_0, i_13_509_3164_0,
    i_13_509_3418_0, i_13_509_3419_0, i_13_509_3424_0, i_13_509_3425_0,
    i_13_509_3427_0, i_13_509_3428_0, i_13_509_3460_0, i_13_509_3487_0,
    i_13_509_3505_0, i_13_509_3580_0, i_13_509_3700_0, i_13_509_3865_0,
    i_13_509_3874_0, i_13_509_3875_0, i_13_509_4085_0, i_13_509_4351_0,
    i_13_509_4352_0, i_13_509_4453_0, i_13_509_4594_0, i_13_509_4598_0;
  output o_13_509_0_0;
  assign o_13_509_0_0 = ~((~i_13_509_539_0 & ((~i_13_509_31_0 & ~i_13_509_2428_0) | (~i_13_509_1843_0 & ~i_13_509_3146_0))) | (~i_13_509_2425_0 & ~i_13_509_2426_0 & ((~i_13_509_1123_0 & ~i_13_509_1628_0) | (~i_13_509_116_0 & ~i_13_509_2428_0 & ~i_13_509_3038_0 & ~i_13_509_3068_0))) | (~i_13_509_32_0 & ~i_13_509_448_0 & ~i_13_509_538_0 & ~i_13_509_2005_0 & ~i_13_509_2680_0) | (i_13_509_3460_0 & i_13_509_3580_0));
endmodule



// Benchmark "kernel_13_510" written by ABC on Sun Jul 19 10:52:25 2020

module kernel_13_510 ( 
    i_13_510_130_0, i_13_510_170_0, i_13_510_187_0, i_13_510_188_0,
    i_13_510_202_0, i_13_510_266_0, i_13_510_269_0, i_13_510_311_0,
    i_13_510_446_0, i_13_510_464_0, i_13_510_583_0, i_13_510_644_0,
    i_13_510_646_0, i_13_510_647_0, i_13_510_697_0, i_13_510_815_0,
    i_13_510_817_0, i_13_510_818_0, i_13_510_844_0, i_13_510_845_0,
    i_13_510_916_0, i_13_510_931_0, i_13_510_950_0, i_13_510_986_0,
    i_13_510_1067_0, i_13_510_1070_0, i_13_510_1123_0, i_13_510_1124_0,
    i_13_510_1247_0, i_13_510_1274_0, i_13_510_1327_0, i_13_510_1331_0,
    i_13_510_1436_0, i_13_510_1490_0, i_13_510_1529_0, i_13_510_1601_0,
    i_13_510_1778_0, i_13_510_1807_0, i_13_510_1808_0, i_13_510_1835_0,
    i_13_510_1849_0, i_13_510_1850_0, i_13_510_1852_0, i_13_510_1853_0,
    i_13_510_1861_0, i_13_510_1933_0, i_13_510_1934_0, i_13_510_2050_0,
    i_13_510_2120_0, i_13_510_2149_0, i_13_510_2201_0, i_13_510_2213_0,
    i_13_510_2263_0, i_13_510_2264_0, i_13_510_2266_0, i_13_510_2267_0,
    i_13_510_2299_0, i_13_510_2345_0, i_13_510_2405_0, i_13_510_2407_0,
    i_13_510_2408_0, i_13_510_2410_0, i_13_510_2411_0, i_13_510_2446_0,
    i_13_510_2462_0, i_13_510_2545_0, i_13_510_2549_0, i_13_510_2600_0,
    i_13_510_2614_0, i_13_510_2698_0, i_13_510_2699_0, i_13_510_2749_0,
    i_13_510_2762_0, i_13_510_2795_0, i_13_510_2798_0, i_13_510_2899_0,
    i_13_510_2941_0, i_13_510_3004_0, i_13_510_3029_0, i_13_510_3094_0,
    i_13_510_3110_0, i_13_510_3112_0, i_13_510_3113_0, i_13_510_3292_0,
    i_13_510_3392_0, i_13_510_3478_0, i_13_510_3526_0, i_13_510_3553_0,
    i_13_510_3580_0, i_13_510_3821_0, i_13_510_3995_0, i_13_510_4066_0,
    i_13_510_4067_0, i_13_510_4171_0, i_13_510_4316_0, i_13_510_4318_0,
    i_13_510_4319_0, i_13_510_4342_0, i_13_510_4568_0, i_13_510_4598_0,
    o_13_510_0_0  );
  input  i_13_510_130_0, i_13_510_170_0, i_13_510_187_0, i_13_510_188_0,
    i_13_510_202_0, i_13_510_266_0, i_13_510_269_0, i_13_510_311_0,
    i_13_510_446_0, i_13_510_464_0, i_13_510_583_0, i_13_510_644_0,
    i_13_510_646_0, i_13_510_647_0, i_13_510_697_0, i_13_510_815_0,
    i_13_510_817_0, i_13_510_818_0, i_13_510_844_0, i_13_510_845_0,
    i_13_510_916_0, i_13_510_931_0, i_13_510_950_0, i_13_510_986_0,
    i_13_510_1067_0, i_13_510_1070_0, i_13_510_1123_0, i_13_510_1124_0,
    i_13_510_1247_0, i_13_510_1274_0, i_13_510_1327_0, i_13_510_1331_0,
    i_13_510_1436_0, i_13_510_1490_0, i_13_510_1529_0, i_13_510_1601_0,
    i_13_510_1778_0, i_13_510_1807_0, i_13_510_1808_0, i_13_510_1835_0,
    i_13_510_1849_0, i_13_510_1850_0, i_13_510_1852_0, i_13_510_1853_0,
    i_13_510_1861_0, i_13_510_1933_0, i_13_510_1934_0, i_13_510_2050_0,
    i_13_510_2120_0, i_13_510_2149_0, i_13_510_2201_0, i_13_510_2213_0,
    i_13_510_2263_0, i_13_510_2264_0, i_13_510_2266_0, i_13_510_2267_0,
    i_13_510_2299_0, i_13_510_2345_0, i_13_510_2405_0, i_13_510_2407_0,
    i_13_510_2408_0, i_13_510_2410_0, i_13_510_2411_0, i_13_510_2446_0,
    i_13_510_2462_0, i_13_510_2545_0, i_13_510_2549_0, i_13_510_2600_0,
    i_13_510_2614_0, i_13_510_2698_0, i_13_510_2699_0, i_13_510_2749_0,
    i_13_510_2762_0, i_13_510_2795_0, i_13_510_2798_0, i_13_510_2899_0,
    i_13_510_2941_0, i_13_510_3004_0, i_13_510_3029_0, i_13_510_3094_0,
    i_13_510_3110_0, i_13_510_3112_0, i_13_510_3113_0, i_13_510_3292_0,
    i_13_510_3392_0, i_13_510_3478_0, i_13_510_3526_0, i_13_510_3553_0,
    i_13_510_3580_0, i_13_510_3821_0, i_13_510_3995_0, i_13_510_4066_0,
    i_13_510_4067_0, i_13_510_4171_0, i_13_510_4316_0, i_13_510_4318_0,
    i_13_510_4319_0, i_13_510_4342_0, i_13_510_4568_0, i_13_510_4598_0;
  output o_13_510_0_0;
  assign o_13_510_0_0 = ~((~i_13_510_2698_0 & (~i_13_510_2762_0 | (~i_13_510_2149_0 & ~i_13_510_4318_0))) | (~i_13_510_1067_0 & ~i_13_510_3995_0 & ~i_13_510_4318_0));
endmodule



// Benchmark "kernel_13_511" written by ABC on Sun Jul 19 10:52:26 2020

module kernel_13_511 ( 
    i_13_511_43_0, i_13_511_48_0, i_13_511_69_0, i_13_511_70_0,
    i_13_511_79_0, i_13_511_141_0, i_13_511_244_0, i_13_511_305_0,
    i_13_511_321_0, i_13_511_322_0, i_13_511_328_0, i_13_511_411_0,
    i_13_511_417_0, i_13_511_448_0, i_13_511_522_0, i_13_511_570_0,
    i_13_511_589_0, i_13_511_591_0, i_13_511_598_0, i_13_511_615_0,
    i_13_511_784_0, i_13_511_924_0, i_13_511_937_0, i_13_511_951_0,
    i_13_511_1023_0, i_13_511_1105_0, i_13_511_1109_0, i_13_511_1122_0,
    i_13_511_1131_0, i_13_511_1132_0, i_13_511_1150_0, i_13_511_1230_0,
    i_13_511_1272_0, i_13_511_1284_0, i_13_511_1329_0, i_13_511_1402_0,
    i_13_511_1510_0, i_13_511_1511_0, i_13_511_1551_0, i_13_511_1644_0,
    i_13_511_1670_0, i_13_511_1722_0, i_13_511_1770_0, i_13_511_1797_0,
    i_13_511_1798_0, i_13_511_1806_0, i_13_511_1831_0, i_13_511_2028_0,
    i_13_511_2118_0, i_13_511_2265_0, i_13_511_2287_0, i_13_511_2296_0,
    i_13_511_2446_0, i_13_511_2461_0, i_13_511_2472_0, i_13_511_2473_0,
    i_13_511_2478_0, i_13_511_2505_0, i_13_511_2514_0, i_13_511_2560_0,
    i_13_511_2581_0, i_13_511_2677_0, i_13_511_2679_0, i_13_511_2680_0,
    i_13_511_2695_0, i_13_511_2698_0, i_13_511_2852_0, i_13_511_2999_0,
    i_13_511_3175_0, i_13_511_3264_0, i_13_511_3273_0, i_13_511_3274_0,
    i_13_511_3432_0, i_13_511_3478_0, i_13_511_3558_0, i_13_511_3561_0,
    i_13_511_3594_0, i_13_511_3640_0, i_13_511_3651_0, i_13_511_3702_0,
    i_13_511_3751_0, i_13_511_3759_0, i_13_511_3787_0, i_13_511_3822_0,
    i_13_511_3864_0, i_13_511_3899_0, i_13_511_3930_0, i_13_511_3940_0,
    i_13_511_4002_0, i_13_511_4036_0, i_13_511_4038_0, i_13_511_4174_0,
    i_13_511_4216_0, i_13_511_4407_0, i_13_511_4435_0, i_13_511_4448_0,
    i_13_511_4450_0, i_13_511_4513_0, i_13_511_4596_0, i_13_511_4597_0,
    o_13_511_0_0  );
  input  i_13_511_43_0, i_13_511_48_0, i_13_511_69_0, i_13_511_70_0,
    i_13_511_79_0, i_13_511_141_0, i_13_511_244_0, i_13_511_305_0,
    i_13_511_321_0, i_13_511_322_0, i_13_511_328_0, i_13_511_411_0,
    i_13_511_417_0, i_13_511_448_0, i_13_511_522_0, i_13_511_570_0,
    i_13_511_589_0, i_13_511_591_0, i_13_511_598_0, i_13_511_615_0,
    i_13_511_784_0, i_13_511_924_0, i_13_511_937_0, i_13_511_951_0,
    i_13_511_1023_0, i_13_511_1105_0, i_13_511_1109_0, i_13_511_1122_0,
    i_13_511_1131_0, i_13_511_1132_0, i_13_511_1150_0, i_13_511_1230_0,
    i_13_511_1272_0, i_13_511_1284_0, i_13_511_1329_0, i_13_511_1402_0,
    i_13_511_1510_0, i_13_511_1511_0, i_13_511_1551_0, i_13_511_1644_0,
    i_13_511_1670_0, i_13_511_1722_0, i_13_511_1770_0, i_13_511_1797_0,
    i_13_511_1798_0, i_13_511_1806_0, i_13_511_1831_0, i_13_511_2028_0,
    i_13_511_2118_0, i_13_511_2265_0, i_13_511_2287_0, i_13_511_2296_0,
    i_13_511_2446_0, i_13_511_2461_0, i_13_511_2472_0, i_13_511_2473_0,
    i_13_511_2478_0, i_13_511_2505_0, i_13_511_2514_0, i_13_511_2560_0,
    i_13_511_2581_0, i_13_511_2677_0, i_13_511_2679_0, i_13_511_2680_0,
    i_13_511_2695_0, i_13_511_2698_0, i_13_511_2852_0, i_13_511_2999_0,
    i_13_511_3175_0, i_13_511_3264_0, i_13_511_3273_0, i_13_511_3274_0,
    i_13_511_3432_0, i_13_511_3478_0, i_13_511_3558_0, i_13_511_3561_0,
    i_13_511_3594_0, i_13_511_3640_0, i_13_511_3651_0, i_13_511_3702_0,
    i_13_511_3751_0, i_13_511_3759_0, i_13_511_3787_0, i_13_511_3822_0,
    i_13_511_3864_0, i_13_511_3899_0, i_13_511_3930_0, i_13_511_3940_0,
    i_13_511_4002_0, i_13_511_4036_0, i_13_511_4038_0, i_13_511_4174_0,
    i_13_511_4216_0, i_13_511_4407_0, i_13_511_4435_0, i_13_511_4448_0,
    i_13_511_4450_0, i_13_511_4513_0, i_13_511_4596_0, i_13_511_4597_0;
  output o_13_511_0_0;
  assign o_13_511_0_0 = ~(~i_13_511_1644_0 | (~i_13_511_70_0 & ~i_13_511_1510_0));
endmodule



module kernel_13 (i_13_0, i_13_1, i_13_2, i_13_3, i_13_4, i_13_5, i_13_6, i_13_7, i_13_8, i_13_9, i_13_10, i_13_11, i_13_12, i_13_13, i_13_14, i_13_15, i_13_16, i_13_17, i_13_18, i_13_19, i_13_20, i_13_21, i_13_22, i_13_23, i_13_24, i_13_25, i_13_26, i_13_27, i_13_28, i_13_29, i_13_30, i_13_31, i_13_32, i_13_33, i_13_34, i_13_35, i_13_36, i_13_37, i_13_38, i_13_39, i_13_40, i_13_41, i_13_42, i_13_43, i_13_44, i_13_45, i_13_46, i_13_47, i_13_48, i_13_49, i_13_50, i_13_51, i_13_52, i_13_53, i_13_54, i_13_55, i_13_56, i_13_57, i_13_58, i_13_59, i_13_60, i_13_61, i_13_62, i_13_63, i_13_64, i_13_65, i_13_66, i_13_67, i_13_68, i_13_69, i_13_70, i_13_71, i_13_72, i_13_73, i_13_74, i_13_75, i_13_76, i_13_77, i_13_78, i_13_79, i_13_80, i_13_81, i_13_82, i_13_83, i_13_84, i_13_85, i_13_86, i_13_87, i_13_88, i_13_89, i_13_90, i_13_91, i_13_92, i_13_93, i_13_94, i_13_95, i_13_96, i_13_97, i_13_98, i_13_99, i_13_100, i_13_101, i_13_102, i_13_103, i_13_104, i_13_105, i_13_106, i_13_107, i_13_108, i_13_109, i_13_110, i_13_111, i_13_112, i_13_113, i_13_114, i_13_115, i_13_116, i_13_117, i_13_118, i_13_119, i_13_120, i_13_121, i_13_122, i_13_123, i_13_124, i_13_125, i_13_126, i_13_127, i_13_128, i_13_129, i_13_130, i_13_131, i_13_132, i_13_133, i_13_134, i_13_135, i_13_136, i_13_137, i_13_138, i_13_139, i_13_140, i_13_141, i_13_142, i_13_143, i_13_144, i_13_145, i_13_146, i_13_147, i_13_148, i_13_149, i_13_150, i_13_151, i_13_152, i_13_153, i_13_154, i_13_155, i_13_156, i_13_157, i_13_158, i_13_159, i_13_160, i_13_161, i_13_162, i_13_163, i_13_164, i_13_165, i_13_166, i_13_167, i_13_168, i_13_169, i_13_170, i_13_171, i_13_172, i_13_173, i_13_174, i_13_175, i_13_176, i_13_177, i_13_178, i_13_179, i_13_180, i_13_181, i_13_182, i_13_183, i_13_184, i_13_185, i_13_186, i_13_187, i_13_188, i_13_189, i_13_190, i_13_191, i_13_192, i_13_193, i_13_194, i_13_195, i_13_196, i_13_197, i_13_198, i_13_199, i_13_200, i_13_201, i_13_202, i_13_203, i_13_204, i_13_205, i_13_206, i_13_207, i_13_208, i_13_209, i_13_210, i_13_211, i_13_212, i_13_213, i_13_214, i_13_215, i_13_216, i_13_217, i_13_218, i_13_219, i_13_220, i_13_221, i_13_222, i_13_223, i_13_224, i_13_225, i_13_226, i_13_227, i_13_228, i_13_229, i_13_230, i_13_231, i_13_232, i_13_233, i_13_234, i_13_235, i_13_236, i_13_237, i_13_238, i_13_239, i_13_240, i_13_241, i_13_242, i_13_243, i_13_244, i_13_245, i_13_246, i_13_247, i_13_248, i_13_249, i_13_250, i_13_251, i_13_252, i_13_253, i_13_254, i_13_255, i_13_256, i_13_257, i_13_258, i_13_259, i_13_260, i_13_261, i_13_262, i_13_263, i_13_264, i_13_265, i_13_266, i_13_267, i_13_268, i_13_269, i_13_270, i_13_271, i_13_272, i_13_273, i_13_274, i_13_275, i_13_276, i_13_277, i_13_278, i_13_279, i_13_280, i_13_281, i_13_282, i_13_283, i_13_284, i_13_285, i_13_286, i_13_287, i_13_288, i_13_289, i_13_290, i_13_291, i_13_292, i_13_293, i_13_294, i_13_295, i_13_296, i_13_297, i_13_298, i_13_299, i_13_300, i_13_301, i_13_302, i_13_303, i_13_304, i_13_305, i_13_306, i_13_307, i_13_308, i_13_309, i_13_310, i_13_311, i_13_312, i_13_313, i_13_314, i_13_315, i_13_316, i_13_317, i_13_318, i_13_319, i_13_320, i_13_321, i_13_322, i_13_323, i_13_324, i_13_325, i_13_326, i_13_327, i_13_328, i_13_329, i_13_330, i_13_331, i_13_332, i_13_333, i_13_334, i_13_335, i_13_336, i_13_337, i_13_338, i_13_339, i_13_340, i_13_341, i_13_342, i_13_343, i_13_344, i_13_345, i_13_346, i_13_347, i_13_348, i_13_349, i_13_350, i_13_351, i_13_352, i_13_353, i_13_354, i_13_355, i_13_356, i_13_357, i_13_358, i_13_359, i_13_360, i_13_361, i_13_362, i_13_363, i_13_364, i_13_365, i_13_366, i_13_367, i_13_368, i_13_369, i_13_370, i_13_371, i_13_372, i_13_373, i_13_374, i_13_375, i_13_376, i_13_377, i_13_378, i_13_379, i_13_380, i_13_381, i_13_382, i_13_383, i_13_384, i_13_385, i_13_386, i_13_387, i_13_388, i_13_389, i_13_390, i_13_391, i_13_392, i_13_393, i_13_394, i_13_395, i_13_396, i_13_397, i_13_398, i_13_399, i_13_400, i_13_401, i_13_402, i_13_403, i_13_404, i_13_405, i_13_406, i_13_407, i_13_408, i_13_409, i_13_410, i_13_411, i_13_412, i_13_413, i_13_414, i_13_415, i_13_416, i_13_417, i_13_418, i_13_419, i_13_420, i_13_421, i_13_422, i_13_423, i_13_424, i_13_425, i_13_426, i_13_427, i_13_428, i_13_429, i_13_430, i_13_431, i_13_432, i_13_433, i_13_434, i_13_435, i_13_436, i_13_437, i_13_438, i_13_439, i_13_440, i_13_441, i_13_442, i_13_443, i_13_444, i_13_445, i_13_446, i_13_447, i_13_448, i_13_449, i_13_450, i_13_451, i_13_452, i_13_453, i_13_454, i_13_455, i_13_456, i_13_457, i_13_458, i_13_459, i_13_460, i_13_461, i_13_462, i_13_463, i_13_464, i_13_465, i_13_466, i_13_467, i_13_468, i_13_469, i_13_470, i_13_471, i_13_472, i_13_473, i_13_474, i_13_475, i_13_476, i_13_477, i_13_478, i_13_479, i_13_480, i_13_481, i_13_482, i_13_483, i_13_484, i_13_485, i_13_486, i_13_487, i_13_488, i_13_489, i_13_490, i_13_491, i_13_492, i_13_493, i_13_494, i_13_495, i_13_496, i_13_497, i_13_498, i_13_499, i_13_500, i_13_501, i_13_502, i_13_503, i_13_504, i_13_505, i_13_506, i_13_507, i_13_508, i_13_509, i_13_510, i_13_511, i_13_512, i_13_513, i_13_514, i_13_515, i_13_516, i_13_517, i_13_518, i_13_519, i_13_520, i_13_521, i_13_522, i_13_523, i_13_524, i_13_525, i_13_526, i_13_527, i_13_528, i_13_529, i_13_530, i_13_531, i_13_532, i_13_533, i_13_534, i_13_535, i_13_536, i_13_537, i_13_538, i_13_539, i_13_540, i_13_541, i_13_542, i_13_543, i_13_544, i_13_545, i_13_546, i_13_547, i_13_548, i_13_549, i_13_550, i_13_551, i_13_552, i_13_553, i_13_554, i_13_555, i_13_556, i_13_557, i_13_558, i_13_559, i_13_560, i_13_561, i_13_562, i_13_563, i_13_564, i_13_565, i_13_566, i_13_567, i_13_568, i_13_569, i_13_570, i_13_571, i_13_572, i_13_573, i_13_574, i_13_575, i_13_576, i_13_577, i_13_578, i_13_579, i_13_580, i_13_581, i_13_582, i_13_583, i_13_584, i_13_585, i_13_586, i_13_587, i_13_588, i_13_589, i_13_590, i_13_591, i_13_592, i_13_593, i_13_594, i_13_595, i_13_596, i_13_597, i_13_598, i_13_599, i_13_600, i_13_601, i_13_602, i_13_603, i_13_604, i_13_605, i_13_606, i_13_607, i_13_608, i_13_609, i_13_610, i_13_611, i_13_612, i_13_613, i_13_614, i_13_615, i_13_616, i_13_617, i_13_618, i_13_619, i_13_620, i_13_621, i_13_622, i_13_623, i_13_624, i_13_625, i_13_626, i_13_627, i_13_628, i_13_629, i_13_630, i_13_631, i_13_632, i_13_633, i_13_634, i_13_635, i_13_636, i_13_637, i_13_638, i_13_639, i_13_640, i_13_641, i_13_642, i_13_643, i_13_644, i_13_645, i_13_646, i_13_647, i_13_648, i_13_649, i_13_650, i_13_651, i_13_652, i_13_653, i_13_654, i_13_655, i_13_656, i_13_657, i_13_658, i_13_659, i_13_660, i_13_661, i_13_662, i_13_663, i_13_664, i_13_665, i_13_666, i_13_667, i_13_668, i_13_669, i_13_670, i_13_671, i_13_672, i_13_673, i_13_674, i_13_675, i_13_676, i_13_677, i_13_678, i_13_679, i_13_680, i_13_681, i_13_682, i_13_683, i_13_684, i_13_685, i_13_686, i_13_687, i_13_688, i_13_689, i_13_690, i_13_691, i_13_692, i_13_693, i_13_694, i_13_695, i_13_696, i_13_697, i_13_698, i_13_699, i_13_700, i_13_701, i_13_702, i_13_703, i_13_704, i_13_705, i_13_706, i_13_707, i_13_708, i_13_709, i_13_710, i_13_711, i_13_712, i_13_713, i_13_714, i_13_715, i_13_716, i_13_717, i_13_718, i_13_719, i_13_720, i_13_721, i_13_722, i_13_723, i_13_724, i_13_725, i_13_726, i_13_727, i_13_728, i_13_729, i_13_730, i_13_731, i_13_732, i_13_733, i_13_734, i_13_735, i_13_736, i_13_737, i_13_738, i_13_739, i_13_740, i_13_741, i_13_742, i_13_743, i_13_744, i_13_745, i_13_746, i_13_747, i_13_748, i_13_749, i_13_750, i_13_751, i_13_752, i_13_753, i_13_754, i_13_755, i_13_756, i_13_757, i_13_758, i_13_759, i_13_760, i_13_761, i_13_762, i_13_763, i_13_764, i_13_765, i_13_766, i_13_767, i_13_768, i_13_769, i_13_770, i_13_771, i_13_772, i_13_773, i_13_774, i_13_775, i_13_776, i_13_777, i_13_778, i_13_779, i_13_780, i_13_781, i_13_782, i_13_783, i_13_784, i_13_785, i_13_786, i_13_787, i_13_788, i_13_789, i_13_790, i_13_791, i_13_792, i_13_793, i_13_794, i_13_795, i_13_796, i_13_797, i_13_798, i_13_799, i_13_800, i_13_801, i_13_802, i_13_803, i_13_804, i_13_805, i_13_806, i_13_807, i_13_808, i_13_809, i_13_810, i_13_811, i_13_812, i_13_813, i_13_814, i_13_815, i_13_816, i_13_817, i_13_818, i_13_819, i_13_820, i_13_821, i_13_822, i_13_823, i_13_824, i_13_825, i_13_826, i_13_827, i_13_828, i_13_829, i_13_830, i_13_831, i_13_832, i_13_833, i_13_834, i_13_835, i_13_836, i_13_837, i_13_838, i_13_839, i_13_840, i_13_841, i_13_842, i_13_843, i_13_844, i_13_845, i_13_846, i_13_847, i_13_848, i_13_849, i_13_850, i_13_851, i_13_852, i_13_853, i_13_854, i_13_855, i_13_856, i_13_857, i_13_858, i_13_859, i_13_860, i_13_861, i_13_862, i_13_863, i_13_864, i_13_865, i_13_866, i_13_867, i_13_868, i_13_869, i_13_870, i_13_871, i_13_872, i_13_873, i_13_874, i_13_875, i_13_876, i_13_877, i_13_878, i_13_879, i_13_880, i_13_881, i_13_882, i_13_883, i_13_884, i_13_885, i_13_886, i_13_887, i_13_888, i_13_889, i_13_890, i_13_891, i_13_892, i_13_893, i_13_894, i_13_895, i_13_896, i_13_897, i_13_898, i_13_899, i_13_900, i_13_901, i_13_902, i_13_903, i_13_904, i_13_905, i_13_906, i_13_907, i_13_908, i_13_909, i_13_910, i_13_911, i_13_912, i_13_913, i_13_914, i_13_915, i_13_916, i_13_917, i_13_918, i_13_919, i_13_920, i_13_921, i_13_922, i_13_923, i_13_924, i_13_925, i_13_926, i_13_927, i_13_928, i_13_929, i_13_930, i_13_931, i_13_932, i_13_933, i_13_934, i_13_935, i_13_936, i_13_937, i_13_938, i_13_939, i_13_940, i_13_941, i_13_942, i_13_943, i_13_944, i_13_945, i_13_946, i_13_947, i_13_948, i_13_949, i_13_950, i_13_951, i_13_952, i_13_953, i_13_954, i_13_955, i_13_956, i_13_957, i_13_958, i_13_959, i_13_960, i_13_961, i_13_962, i_13_963, i_13_964, i_13_965, i_13_966, i_13_967, i_13_968, i_13_969, i_13_970, i_13_971, i_13_972, i_13_973, i_13_974, i_13_975, i_13_976, i_13_977, i_13_978, i_13_979, i_13_980, i_13_981, i_13_982, i_13_983, i_13_984, i_13_985, i_13_986, i_13_987, i_13_988, i_13_989, i_13_990, i_13_991, i_13_992, i_13_993, i_13_994, i_13_995, i_13_996, i_13_997, i_13_998, i_13_999, i_13_1000, i_13_1001, i_13_1002, i_13_1003, i_13_1004, i_13_1005, i_13_1006, i_13_1007, i_13_1008, i_13_1009, i_13_1010, i_13_1011, i_13_1012, i_13_1013, i_13_1014, i_13_1015, i_13_1016, i_13_1017, i_13_1018, i_13_1019, i_13_1020, i_13_1021, i_13_1022, i_13_1023, i_13_1024, i_13_1025, i_13_1026, i_13_1027, i_13_1028, i_13_1029, i_13_1030, i_13_1031, i_13_1032, i_13_1033, i_13_1034, i_13_1035, i_13_1036, i_13_1037, i_13_1038, i_13_1039, i_13_1040, i_13_1041, i_13_1042, i_13_1043, i_13_1044, i_13_1045, i_13_1046, i_13_1047, i_13_1048, i_13_1049, i_13_1050, i_13_1051, i_13_1052, i_13_1053, i_13_1054, i_13_1055, i_13_1056, i_13_1057, i_13_1058, i_13_1059, i_13_1060, i_13_1061, i_13_1062, i_13_1063, i_13_1064, i_13_1065, i_13_1066, i_13_1067, i_13_1068, i_13_1069, i_13_1070, i_13_1071, i_13_1072, i_13_1073, i_13_1074, i_13_1075, i_13_1076, i_13_1077, i_13_1078, i_13_1079, i_13_1080, i_13_1081, i_13_1082, i_13_1083, i_13_1084, i_13_1085, i_13_1086, i_13_1087, i_13_1088, i_13_1089, i_13_1090, i_13_1091, i_13_1092, i_13_1093, i_13_1094, i_13_1095, i_13_1096, i_13_1097, i_13_1098, i_13_1099, i_13_1100, i_13_1101, i_13_1102, i_13_1103, i_13_1104, i_13_1105, i_13_1106, i_13_1107, i_13_1108, i_13_1109, i_13_1110, i_13_1111, i_13_1112, i_13_1113, i_13_1114, i_13_1115, i_13_1116, i_13_1117, i_13_1118, i_13_1119, i_13_1120, i_13_1121, i_13_1122, i_13_1123, i_13_1124, i_13_1125, i_13_1126, i_13_1127, i_13_1128, i_13_1129, i_13_1130, i_13_1131, i_13_1132, i_13_1133, i_13_1134, i_13_1135, i_13_1136, i_13_1137, i_13_1138, i_13_1139, i_13_1140, i_13_1141, i_13_1142, i_13_1143, i_13_1144, i_13_1145, i_13_1146, i_13_1147, i_13_1148, i_13_1149, i_13_1150, i_13_1151, i_13_1152, i_13_1153, i_13_1154, i_13_1155, i_13_1156, i_13_1157, i_13_1158, i_13_1159, i_13_1160, i_13_1161, i_13_1162, i_13_1163, i_13_1164, i_13_1165, i_13_1166, i_13_1167, i_13_1168, i_13_1169, i_13_1170, i_13_1171, i_13_1172, i_13_1173, i_13_1174, i_13_1175, i_13_1176, i_13_1177, i_13_1178, i_13_1179, i_13_1180, i_13_1181, i_13_1182, i_13_1183, i_13_1184, i_13_1185, i_13_1186, i_13_1187, i_13_1188, i_13_1189, i_13_1190, i_13_1191, i_13_1192, i_13_1193, i_13_1194, i_13_1195, i_13_1196, i_13_1197, i_13_1198, i_13_1199, i_13_1200, i_13_1201, i_13_1202, i_13_1203, i_13_1204, i_13_1205, i_13_1206, i_13_1207, i_13_1208, i_13_1209, i_13_1210, i_13_1211, i_13_1212, i_13_1213, i_13_1214, i_13_1215, i_13_1216, i_13_1217, i_13_1218, i_13_1219, i_13_1220, i_13_1221, i_13_1222, i_13_1223, i_13_1224, i_13_1225, i_13_1226, i_13_1227, i_13_1228, i_13_1229, i_13_1230, i_13_1231, i_13_1232, i_13_1233, i_13_1234, i_13_1235, i_13_1236, i_13_1237, i_13_1238, i_13_1239, i_13_1240, i_13_1241, i_13_1242, i_13_1243, i_13_1244, i_13_1245, i_13_1246, i_13_1247, i_13_1248, i_13_1249, i_13_1250, i_13_1251, i_13_1252, i_13_1253, i_13_1254, i_13_1255, i_13_1256, i_13_1257, i_13_1258, i_13_1259, i_13_1260, i_13_1261, i_13_1262, i_13_1263, i_13_1264, i_13_1265, i_13_1266, i_13_1267, i_13_1268, i_13_1269, i_13_1270, i_13_1271, i_13_1272, i_13_1273, i_13_1274, i_13_1275, i_13_1276, i_13_1277, i_13_1278, i_13_1279, i_13_1280, i_13_1281, i_13_1282, i_13_1283, i_13_1284, i_13_1285, i_13_1286, i_13_1287, i_13_1288, i_13_1289, i_13_1290, i_13_1291, i_13_1292, i_13_1293, i_13_1294, i_13_1295, i_13_1296, i_13_1297, i_13_1298, i_13_1299, i_13_1300, i_13_1301, i_13_1302, i_13_1303, i_13_1304, i_13_1305, i_13_1306, i_13_1307, i_13_1308, i_13_1309, i_13_1310, i_13_1311, i_13_1312, i_13_1313, i_13_1314, i_13_1315, i_13_1316, i_13_1317, i_13_1318, i_13_1319, i_13_1320, i_13_1321, i_13_1322, i_13_1323, i_13_1324, i_13_1325, i_13_1326, i_13_1327, i_13_1328, i_13_1329, i_13_1330, i_13_1331, i_13_1332, i_13_1333, i_13_1334, i_13_1335, i_13_1336, i_13_1337, i_13_1338, i_13_1339, i_13_1340, i_13_1341, i_13_1342, i_13_1343, i_13_1344, i_13_1345, i_13_1346, i_13_1347, i_13_1348, i_13_1349, i_13_1350, i_13_1351, i_13_1352, i_13_1353, i_13_1354, i_13_1355, i_13_1356, i_13_1357, i_13_1358, i_13_1359, i_13_1360, i_13_1361, i_13_1362, i_13_1363, i_13_1364, i_13_1365, i_13_1366, i_13_1367, i_13_1368, i_13_1369, i_13_1370, i_13_1371, i_13_1372, i_13_1373, i_13_1374, i_13_1375, i_13_1376, i_13_1377, i_13_1378, i_13_1379, i_13_1380, i_13_1381, i_13_1382, i_13_1383, i_13_1384, i_13_1385, i_13_1386, i_13_1387, i_13_1388, i_13_1389, i_13_1390, i_13_1391, i_13_1392, i_13_1393, i_13_1394, i_13_1395, i_13_1396, i_13_1397, i_13_1398, i_13_1399, i_13_1400, i_13_1401, i_13_1402, i_13_1403, i_13_1404, i_13_1405, i_13_1406, i_13_1407, i_13_1408, i_13_1409, i_13_1410, i_13_1411, i_13_1412, i_13_1413, i_13_1414, i_13_1415, i_13_1416, i_13_1417, i_13_1418, i_13_1419, i_13_1420, i_13_1421, i_13_1422, i_13_1423, i_13_1424, i_13_1425, i_13_1426, i_13_1427, i_13_1428, i_13_1429, i_13_1430, i_13_1431, i_13_1432, i_13_1433, i_13_1434, i_13_1435, i_13_1436, i_13_1437, i_13_1438, i_13_1439, i_13_1440, i_13_1441, i_13_1442, i_13_1443, i_13_1444, i_13_1445, i_13_1446, i_13_1447, i_13_1448, i_13_1449, i_13_1450, i_13_1451, i_13_1452, i_13_1453, i_13_1454, i_13_1455, i_13_1456, i_13_1457, i_13_1458, i_13_1459, i_13_1460, i_13_1461, i_13_1462, i_13_1463, i_13_1464, i_13_1465, i_13_1466, i_13_1467, i_13_1468, i_13_1469, i_13_1470, i_13_1471, i_13_1472, i_13_1473, i_13_1474, i_13_1475, i_13_1476, i_13_1477, i_13_1478, i_13_1479, i_13_1480, i_13_1481, i_13_1482, i_13_1483, i_13_1484, i_13_1485, i_13_1486, i_13_1487, i_13_1488, i_13_1489, i_13_1490, i_13_1491, i_13_1492, i_13_1493, i_13_1494, i_13_1495, i_13_1496, i_13_1497, i_13_1498, i_13_1499, i_13_1500, i_13_1501, i_13_1502, i_13_1503, i_13_1504, i_13_1505, i_13_1506, i_13_1507, i_13_1508, i_13_1509, i_13_1510, i_13_1511, i_13_1512, i_13_1513, i_13_1514, i_13_1515, i_13_1516, i_13_1517, i_13_1518, i_13_1519, i_13_1520, i_13_1521, i_13_1522, i_13_1523, i_13_1524, i_13_1525, i_13_1526, i_13_1527, i_13_1528, i_13_1529, i_13_1530, i_13_1531, i_13_1532, i_13_1533, i_13_1534, i_13_1535, i_13_1536, i_13_1537, i_13_1538, i_13_1539, i_13_1540, i_13_1541, i_13_1542, i_13_1543, i_13_1544, i_13_1545, i_13_1546, i_13_1547, i_13_1548, i_13_1549, i_13_1550, i_13_1551, i_13_1552, i_13_1553, i_13_1554, i_13_1555, i_13_1556, i_13_1557, i_13_1558, i_13_1559, i_13_1560, i_13_1561, i_13_1562, i_13_1563, i_13_1564, i_13_1565, i_13_1566, i_13_1567, i_13_1568, i_13_1569, i_13_1570, i_13_1571, i_13_1572, i_13_1573, i_13_1574, i_13_1575, i_13_1576, i_13_1577, i_13_1578, i_13_1579, i_13_1580, i_13_1581, i_13_1582, i_13_1583, i_13_1584, i_13_1585, i_13_1586, i_13_1587, i_13_1588, i_13_1589, i_13_1590, i_13_1591, i_13_1592, i_13_1593, i_13_1594, i_13_1595, i_13_1596, i_13_1597, i_13_1598, i_13_1599, i_13_1600, i_13_1601, i_13_1602, i_13_1603, i_13_1604, i_13_1605, i_13_1606, i_13_1607, i_13_1608, i_13_1609, i_13_1610, i_13_1611, i_13_1612, i_13_1613, i_13_1614, i_13_1615, i_13_1616, i_13_1617, i_13_1618, i_13_1619, i_13_1620, i_13_1621, i_13_1622, i_13_1623, i_13_1624, i_13_1625, i_13_1626, i_13_1627, i_13_1628, i_13_1629, i_13_1630, i_13_1631, i_13_1632, i_13_1633, i_13_1634, i_13_1635, i_13_1636, i_13_1637, i_13_1638, i_13_1639, i_13_1640, i_13_1641, i_13_1642, i_13_1643, i_13_1644, i_13_1645, i_13_1646, i_13_1647, i_13_1648, i_13_1649, i_13_1650, i_13_1651, i_13_1652, i_13_1653, i_13_1654, i_13_1655, i_13_1656, i_13_1657, i_13_1658, i_13_1659, i_13_1660, i_13_1661, i_13_1662, i_13_1663, i_13_1664, i_13_1665, i_13_1666, i_13_1667, i_13_1668, i_13_1669, i_13_1670, i_13_1671, i_13_1672, i_13_1673, i_13_1674, i_13_1675, i_13_1676, i_13_1677, i_13_1678, i_13_1679, i_13_1680, i_13_1681, i_13_1682, i_13_1683, i_13_1684, i_13_1685, i_13_1686, i_13_1687, i_13_1688, i_13_1689, i_13_1690, i_13_1691, i_13_1692, i_13_1693, i_13_1694, i_13_1695, i_13_1696, i_13_1697, i_13_1698, i_13_1699, i_13_1700, i_13_1701, i_13_1702, i_13_1703, i_13_1704, i_13_1705, i_13_1706, i_13_1707, i_13_1708, i_13_1709, i_13_1710, i_13_1711, i_13_1712, i_13_1713, i_13_1714, i_13_1715, i_13_1716, i_13_1717, i_13_1718, i_13_1719, i_13_1720, i_13_1721, i_13_1722, i_13_1723, i_13_1724, i_13_1725, i_13_1726, i_13_1727, i_13_1728, i_13_1729, i_13_1730, i_13_1731, i_13_1732, i_13_1733, i_13_1734, i_13_1735, i_13_1736, i_13_1737, i_13_1738, i_13_1739, i_13_1740, i_13_1741, i_13_1742, i_13_1743, i_13_1744, i_13_1745, i_13_1746, i_13_1747, i_13_1748, i_13_1749, i_13_1750, i_13_1751, i_13_1752, i_13_1753, i_13_1754, i_13_1755, i_13_1756, i_13_1757, i_13_1758, i_13_1759, i_13_1760, i_13_1761, i_13_1762, i_13_1763, i_13_1764, i_13_1765, i_13_1766, i_13_1767, i_13_1768, i_13_1769, i_13_1770, i_13_1771, i_13_1772, i_13_1773, i_13_1774, i_13_1775, i_13_1776, i_13_1777, i_13_1778, i_13_1779, i_13_1780, i_13_1781, i_13_1782, i_13_1783, i_13_1784, i_13_1785, i_13_1786, i_13_1787, i_13_1788, i_13_1789, i_13_1790, i_13_1791, i_13_1792, i_13_1793, i_13_1794, i_13_1795, i_13_1796, i_13_1797, i_13_1798, i_13_1799, i_13_1800, i_13_1801, i_13_1802, i_13_1803, i_13_1804, i_13_1805, i_13_1806, i_13_1807, i_13_1808, i_13_1809, i_13_1810, i_13_1811, i_13_1812, i_13_1813, i_13_1814, i_13_1815, i_13_1816, i_13_1817, i_13_1818, i_13_1819, i_13_1820, i_13_1821, i_13_1822, i_13_1823, i_13_1824, i_13_1825, i_13_1826, i_13_1827, i_13_1828, i_13_1829, i_13_1830, i_13_1831, i_13_1832, i_13_1833, i_13_1834, i_13_1835, i_13_1836, i_13_1837, i_13_1838, i_13_1839, i_13_1840, i_13_1841, i_13_1842, i_13_1843, i_13_1844, i_13_1845, i_13_1846, i_13_1847, i_13_1848, i_13_1849, i_13_1850, i_13_1851, i_13_1852, i_13_1853, i_13_1854, i_13_1855, i_13_1856, i_13_1857, i_13_1858, i_13_1859, i_13_1860, i_13_1861, i_13_1862, i_13_1863, i_13_1864, i_13_1865, i_13_1866, i_13_1867, i_13_1868, i_13_1869, i_13_1870, i_13_1871, i_13_1872, i_13_1873, i_13_1874, i_13_1875, i_13_1876, i_13_1877, i_13_1878, i_13_1879, i_13_1880, i_13_1881, i_13_1882, i_13_1883, i_13_1884, i_13_1885, i_13_1886, i_13_1887, i_13_1888, i_13_1889, i_13_1890, i_13_1891, i_13_1892, i_13_1893, i_13_1894, i_13_1895, i_13_1896, i_13_1897, i_13_1898, i_13_1899, i_13_1900, i_13_1901, i_13_1902, i_13_1903, i_13_1904, i_13_1905, i_13_1906, i_13_1907, i_13_1908, i_13_1909, i_13_1910, i_13_1911, i_13_1912, i_13_1913, i_13_1914, i_13_1915, i_13_1916, i_13_1917, i_13_1918, i_13_1919, i_13_1920, i_13_1921, i_13_1922, i_13_1923, i_13_1924, i_13_1925, i_13_1926, i_13_1927, i_13_1928, i_13_1929, i_13_1930, i_13_1931, i_13_1932, i_13_1933, i_13_1934, i_13_1935, i_13_1936, i_13_1937, i_13_1938, i_13_1939, i_13_1940, i_13_1941, i_13_1942, i_13_1943, i_13_1944, i_13_1945, i_13_1946, i_13_1947, i_13_1948, i_13_1949, i_13_1950, i_13_1951, i_13_1952, i_13_1953, i_13_1954, i_13_1955, i_13_1956, i_13_1957, i_13_1958, i_13_1959, i_13_1960, i_13_1961, i_13_1962, i_13_1963, i_13_1964, i_13_1965, i_13_1966, i_13_1967, i_13_1968, i_13_1969, i_13_1970, i_13_1971, i_13_1972, i_13_1973, i_13_1974, i_13_1975, i_13_1976, i_13_1977, i_13_1978, i_13_1979, i_13_1980, i_13_1981, i_13_1982, i_13_1983, i_13_1984, i_13_1985, i_13_1986, i_13_1987, i_13_1988, i_13_1989, i_13_1990, i_13_1991, i_13_1992, i_13_1993, i_13_1994, i_13_1995, i_13_1996, i_13_1997, i_13_1998, i_13_1999, i_13_2000, i_13_2001, i_13_2002, i_13_2003, i_13_2004, i_13_2005, i_13_2006, i_13_2007, i_13_2008, i_13_2009, i_13_2010, i_13_2011, i_13_2012, i_13_2013, i_13_2014, i_13_2015, i_13_2016, i_13_2017, i_13_2018, i_13_2019, i_13_2020, i_13_2021, i_13_2022, i_13_2023, i_13_2024, i_13_2025, i_13_2026, i_13_2027, i_13_2028, i_13_2029, i_13_2030, i_13_2031, i_13_2032, i_13_2033, i_13_2034, i_13_2035, i_13_2036, i_13_2037, i_13_2038, i_13_2039, i_13_2040, i_13_2041, i_13_2042, i_13_2043, i_13_2044, i_13_2045, i_13_2046, i_13_2047, i_13_2048, i_13_2049, i_13_2050, i_13_2051, i_13_2052, i_13_2053, i_13_2054, i_13_2055, i_13_2056, i_13_2057, i_13_2058, i_13_2059, i_13_2060, i_13_2061, i_13_2062, i_13_2063, i_13_2064, i_13_2065, i_13_2066, i_13_2067, i_13_2068, i_13_2069, i_13_2070, i_13_2071, i_13_2072, i_13_2073, i_13_2074, i_13_2075, i_13_2076, i_13_2077, i_13_2078, i_13_2079, i_13_2080, i_13_2081, i_13_2082, i_13_2083, i_13_2084, i_13_2085, i_13_2086, i_13_2087, i_13_2088, i_13_2089, i_13_2090, i_13_2091, i_13_2092, i_13_2093, i_13_2094, i_13_2095, i_13_2096, i_13_2097, i_13_2098, i_13_2099, i_13_2100, i_13_2101, i_13_2102, i_13_2103, i_13_2104, i_13_2105, i_13_2106, i_13_2107, i_13_2108, i_13_2109, i_13_2110, i_13_2111, i_13_2112, i_13_2113, i_13_2114, i_13_2115, i_13_2116, i_13_2117, i_13_2118, i_13_2119, i_13_2120, i_13_2121, i_13_2122, i_13_2123, i_13_2124, i_13_2125, i_13_2126, i_13_2127, i_13_2128, i_13_2129, i_13_2130, i_13_2131, i_13_2132, i_13_2133, i_13_2134, i_13_2135, i_13_2136, i_13_2137, i_13_2138, i_13_2139, i_13_2140, i_13_2141, i_13_2142, i_13_2143, i_13_2144, i_13_2145, i_13_2146, i_13_2147, i_13_2148, i_13_2149, i_13_2150, i_13_2151, i_13_2152, i_13_2153, i_13_2154, i_13_2155, i_13_2156, i_13_2157, i_13_2158, i_13_2159, i_13_2160, i_13_2161, i_13_2162, i_13_2163, i_13_2164, i_13_2165, i_13_2166, i_13_2167, i_13_2168, i_13_2169, i_13_2170, i_13_2171, i_13_2172, i_13_2173, i_13_2174, i_13_2175, i_13_2176, i_13_2177, i_13_2178, i_13_2179, i_13_2180, i_13_2181, i_13_2182, i_13_2183, i_13_2184, i_13_2185, i_13_2186, i_13_2187, i_13_2188, i_13_2189, i_13_2190, i_13_2191, i_13_2192, i_13_2193, i_13_2194, i_13_2195, i_13_2196, i_13_2197, i_13_2198, i_13_2199, i_13_2200, i_13_2201, i_13_2202, i_13_2203, i_13_2204, i_13_2205, i_13_2206, i_13_2207, i_13_2208, i_13_2209, i_13_2210, i_13_2211, i_13_2212, i_13_2213, i_13_2214, i_13_2215, i_13_2216, i_13_2217, i_13_2218, i_13_2219, i_13_2220, i_13_2221, i_13_2222, i_13_2223, i_13_2224, i_13_2225, i_13_2226, i_13_2227, i_13_2228, i_13_2229, i_13_2230, i_13_2231, i_13_2232, i_13_2233, i_13_2234, i_13_2235, i_13_2236, i_13_2237, i_13_2238, i_13_2239, i_13_2240, i_13_2241, i_13_2242, i_13_2243, i_13_2244, i_13_2245, i_13_2246, i_13_2247, i_13_2248, i_13_2249, i_13_2250, i_13_2251, i_13_2252, i_13_2253, i_13_2254, i_13_2255, i_13_2256, i_13_2257, i_13_2258, i_13_2259, i_13_2260, i_13_2261, i_13_2262, i_13_2263, i_13_2264, i_13_2265, i_13_2266, i_13_2267, i_13_2268, i_13_2269, i_13_2270, i_13_2271, i_13_2272, i_13_2273, i_13_2274, i_13_2275, i_13_2276, i_13_2277, i_13_2278, i_13_2279, i_13_2280, i_13_2281, i_13_2282, i_13_2283, i_13_2284, i_13_2285, i_13_2286, i_13_2287, i_13_2288, i_13_2289, i_13_2290, i_13_2291, i_13_2292, i_13_2293, i_13_2294, i_13_2295, i_13_2296, i_13_2297, i_13_2298, i_13_2299, i_13_2300, i_13_2301, i_13_2302, i_13_2303, i_13_2304, i_13_2305, i_13_2306, i_13_2307, i_13_2308, i_13_2309, i_13_2310, i_13_2311, i_13_2312, i_13_2313, i_13_2314, i_13_2315, i_13_2316, i_13_2317, i_13_2318, i_13_2319, i_13_2320, i_13_2321, i_13_2322, i_13_2323, i_13_2324, i_13_2325, i_13_2326, i_13_2327, i_13_2328, i_13_2329, i_13_2330, i_13_2331, i_13_2332, i_13_2333, i_13_2334, i_13_2335, i_13_2336, i_13_2337, i_13_2338, i_13_2339, i_13_2340, i_13_2341, i_13_2342, i_13_2343, i_13_2344, i_13_2345, i_13_2346, i_13_2347, i_13_2348, i_13_2349, i_13_2350, i_13_2351, i_13_2352, i_13_2353, i_13_2354, i_13_2355, i_13_2356, i_13_2357, i_13_2358, i_13_2359, i_13_2360, i_13_2361, i_13_2362, i_13_2363, i_13_2364, i_13_2365, i_13_2366, i_13_2367, i_13_2368, i_13_2369, i_13_2370, i_13_2371, i_13_2372, i_13_2373, i_13_2374, i_13_2375, i_13_2376, i_13_2377, i_13_2378, i_13_2379, i_13_2380, i_13_2381, i_13_2382, i_13_2383, i_13_2384, i_13_2385, i_13_2386, i_13_2387, i_13_2388, i_13_2389, i_13_2390, i_13_2391, i_13_2392, i_13_2393, i_13_2394, i_13_2395, i_13_2396, i_13_2397, i_13_2398, i_13_2399, i_13_2400, i_13_2401, i_13_2402, i_13_2403, i_13_2404, i_13_2405, i_13_2406, i_13_2407, i_13_2408, i_13_2409, i_13_2410, i_13_2411, i_13_2412, i_13_2413, i_13_2414, i_13_2415, i_13_2416, i_13_2417, i_13_2418, i_13_2419, i_13_2420, i_13_2421, i_13_2422, i_13_2423, i_13_2424, i_13_2425, i_13_2426, i_13_2427, i_13_2428, i_13_2429, i_13_2430, i_13_2431, i_13_2432, i_13_2433, i_13_2434, i_13_2435, i_13_2436, i_13_2437, i_13_2438, i_13_2439, i_13_2440, i_13_2441, i_13_2442, i_13_2443, i_13_2444, i_13_2445, i_13_2446, i_13_2447, i_13_2448, i_13_2449, i_13_2450, i_13_2451, i_13_2452, i_13_2453, i_13_2454, i_13_2455, i_13_2456, i_13_2457, i_13_2458, i_13_2459, i_13_2460, i_13_2461, i_13_2462, i_13_2463, i_13_2464, i_13_2465, i_13_2466, i_13_2467, i_13_2468, i_13_2469, i_13_2470, i_13_2471, i_13_2472, i_13_2473, i_13_2474, i_13_2475, i_13_2476, i_13_2477, i_13_2478, i_13_2479, i_13_2480, i_13_2481, i_13_2482, i_13_2483, i_13_2484, i_13_2485, i_13_2486, i_13_2487, i_13_2488, i_13_2489, i_13_2490, i_13_2491, i_13_2492, i_13_2493, i_13_2494, i_13_2495, i_13_2496, i_13_2497, i_13_2498, i_13_2499, i_13_2500, i_13_2501, i_13_2502, i_13_2503, i_13_2504, i_13_2505, i_13_2506, i_13_2507, i_13_2508, i_13_2509, i_13_2510, i_13_2511, i_13_2512, i_13_2513, i_13_2514, i_13_2515, i_13_2516, i_13_2517, i_13_2518, i_13_2519, i_13_2520, i_13_2521, i_13_2522, i_13_2523, i_13_2524, i_13_2525, i_13_2526, i_13_2527, i_13_2528, i_13_2529, i_13_2530, i_13_2531, i_13_2532, i_13_2533, i_13_2534, i_13_2535, i_13_2536, i_13_2537, i_13_2538, i_13_2539, i_13_2540, i_13_2541, i_13_2542, i_13_2543, i_13_2544, i_13_2545, i_13_2546, i_13_2547, i_13_2548, i_13_2549, i_13_2550, i_13_2551, i_13_2552, i_13_2553, i_13_2554, i_13_2555, i_13_2556, i_13_2557, i_13_2558, i_13_2559, i_13_2560, i_13_2561, i_13_2562, i_13_2563, i_13_2564, i_13_2565, i_13_2566, i_13_2567, i_13_2568, i_13_2569, i_13_2570, i_13_2571, i_13_2572, i_13_2573, i_13_2574, i_13_2575, i_13_2576, i_13_2577, i_13_2578, i_13_2579, i_13_2580, i_13_2581, i_13_2582, i_13_2583, i_13_2584, i_13_2585, i_13_2586, i_13_2587, i_13_2588, i_13_2589, i_13_2590, i_13_2591, i_13_2592, i_13_2593, i_13_2594, i_13_2595, i_13_2596, i_13_2597, i_13_2598, i_13_2599, i_13_2600, i_13_2601, i_13_2602, i_13_2603, i_13_2604, i_13_2605, i_13_2606, i_13_2607, i_13_2608, i_13_2609, i_13_2610, i_13_2611, i_13_2612, i_13_2613, i_13_2614, i_13_2615, i_13_2616, i_13_2617, i_13_2618, i_13_2619, i_13_2620, i_13_2621, i_13_2622, i_13_2623, i_13_2624, i_13_2625, i_13_2626, i_13_2627, i_13_2628, i_13_2629, i_13_2630, i_13_2631, i_13_2632, i_13_2633, i_13_2634, i_13_2635, i_13_2636, i_13_2637, i_13_2638, i_13_2639, i_13_2640, i_13_2641, i_13_2642, i_13_2643, i_13_2644, i_13_2645, i_13_2646, i_13_2647, i_13_2648, i_13_2649, i_13_2650, i_13_2651, i_13_2652, i_13_2653, i_13_2654, i_13_2655, i_13_2656, i_13_2657, i_13_2658, i_13_2659, i_13_2660, i_13_2661, i_13_2662, i_13_2663, i_13_2664, i_13_2665, i_13_2666, i_13_2667, i_13_2668, i_13_2669, i_13_2670, i_13_2671, i_13_2672, i_13_2673, i_13_2674, i_13_2675, i_13_2676, i_13_2677, i_13_2678, i_13_2679, i_13_2680, i_13_2681, i_13_2682, i_13_2683, i_13_2684, i_13_2685, i_13_2686, i_13_2687, i_13_2688, i_13_2689, i_13_2690, i_13_2691, i_13_2692, i_13_2693, i_13_2694, i_13_2695, i_13_2696, i_13_2697, i_13_2698, i_13_2699, i_13_2700, i_13_2701, i_13_2702, i_13_2703, i_13_2704, i_13_2705, i_13_2706, i_13_2707, i_13_2708, i_13_2709, i_13_2710, i_13_2711, i_13_2712, i_13_2713, i_13_2714, i_13_2715, i_13_2716, i_13_2717, i_13_2718, i_13_2719, i_13_2720, i_13_2721, i_13_2722, i_13_2723, i_13_2724, i_13_2725, i_13_2726, i_13_2727, i_13_2728, i_13_2729, i_13_2730, i_13_2731, i_13_2732, i_13_2733, i_13_2734, i_13_2735, i_13_2736, i_13_2737, i_13_2738, i_13_2739, i_13_2740, i_13_2741, i_13_2742, i_13_2743, i_13_2744, i_13_2745, i_13_2746, i_13_2747, i_13_2748, i_13_2749, i_13_2750, i_13_2751, i_13_2752, i_13_2753, i_13_2754, i_13_2755, i_13_2756, i_13_2757, i_13_2758, i_13_2759, i_13_2760, i_13_2761, i_13_2762, i_13_2763, i_13_2764, i_13_2765, i_13_2766, i_13_2767, i_13_2768, i_13_2769, i_13_2770, i_13_2771, i_13_2772, i_13_2773, i_13_2774, i_13_2775, i_13_2776, i_13_2777, i_13_2778, i_13_2779, i_13_2780, i_13_2781, i_13_2782, i_13_2783, i_13_2784, i_13_2785, i_13_2786, i_13_2787, i_13_2788, i_13_2789, i_13_2790, i_13_2791, i_13_2792, i_13_2793, i_13_2794, i_13_2795, i_13_2796, i_13_2797, i_13_2798, i_13_2799, i_13_2800, i_13_2801, i_13_2802, i_13_2803, i_13_2804, i_13_2805, i_13_2806, i_13_2807, i_13_2808, i_13_2809, i_13_2810, i_13_2811, i_13_2812, i_13_2813, i_13_2814, i_13_2815, i_13_2816, i_13_2817, i_13_2818, i_13_2819, i_13_2820, i_13_2821, i_13_2822, i_13_2823, i_13_2824, i_13_2825, i_13_2826, i_13_2827, i_13_2828, i_13_2829, i_13_2830, i_13_2831, i_13_2832, i_13_2833, i_13_2834, i_13_2835, i_13_2836, i_13_2837, i_13_2838, i_13_2839, i_13_2840, i_13_2841, i_13_2842, i_13_2843, i_13_2844, i_13_2845, i_13_2846, i_13_2847, i_13_2848, i_13_2849, i_13_2850, i_13_2851, i_13_2852, i_13_2853, i_13_2854, i_13_2855, i_13_2856, i_13_2857, i_13_2858, i_13_2859, i_13_2860, i_13_2861, i_13_2862, i_13_2863, i_13_2864, i_13_2865, i_13_2866, i_13_2867, i_13_2868, i_13_2869, i_13_2870, i_13_2871, i_13_2872, i_13_2873, i_13_2874, i_13_2875, i_13_2876, i_13_2877, i_13_2878, i_13_2879, i_13_2880, i_13_2881, i_13_2882, i_13_2883, i_13_2884, i_13_2885, i_13_2886, i_13_2887, i_13_2888, i_13_2889, i_13_2890, i_13_2891, i_13_2892, i_13_2893, i_13_2894, i_13_2895, i_13_2896, i_13_2897, i_13_2898, i_13_2899, i_13_2900, i_13_2901, i_13_2902, i_13_2903, i_13_2904, i_13_2905, i_13_2906, i_13_2907, i_13_2908, i_13_2909, i_13_2910, i_13_2911, i_13_2912, i_13_2913, i_13_2914, i_13_2915, i_13_2916, i_13_2917, i_13_2918, i_13_2919, i_13_2920, i_13_2921, i_13_2922, i_13_2923, i_13_2924, i_13_2925, i_13_2926, i_13_2927, i_13_2928, i_13_2929, i_13_2930, i_13_2931, i_13_2932, i_13_2933, i_13_2934, i_13_2935, i_13_2936, i_13_2937, i_13_2938, i_13_2939, i_13_2940, i_13_2941, i_13_2942, i_13_2943, i_13_2944, i_13_2945, i_13_2946, i_13_2947, i_13_2948, i_13_2949, i_13_2950, i_13_2951, i_13_2952, i_13_2953, i_13_2954, i_13_2955, i_13_2956, i_13_2957, i_13_2958, i_13_2959, i_13_2960, i_13_2961, i_13_2962, i_13_2963, i_13_2964, i_13_2965, i_13_2966, i_13_2967, i_13_2968, i_13_2969, i_13_2970, i_13_2971, i_13_2972, i_13_2973, i_13_2974, i_13_2975, i_13_2976, i_13_2977, i_13_2978, i_13_2979, i_13_2980, i_13_2981, i_13_2982, i_13_2983, i_13_2984, i_13_2985, i_13_2986, i_13_2987, i_13_2988, i_13_2989, i_13_2990, i_13_2991, i_13_2992, i_13_2993, i_13_2994, i_13_2995, i_13_2996, i_13_2997, i_13_2998, i_13_2999, i_13_3000, i_13_3001, i_13_3002, i_13_3003, i_13_3004, i_13_3005, i_13_3006, i_13_3007, i_13_3008, i_13_3009, i_13_3010, i_13_3011, i_13_3012, i_13_3013, i_13_3014, i_13_3015, i_13_3016, i_13_3017, i_13_3018, i_13_3019, i_13_3020, i_13_3021, i_13_3022, i_13_3023, i_13_3024, i_13_3025, i_13_3026, i_13_3027, i_13_3028, i_13_3029, i_13_3030, i_13_3031, i_13_3032, i_13_3033, i_13_3034, i_13_3035, i_13_3036, i_13_3037, i_13_3038, i_13_3039, i_13_3040, i_13_3041, i_13_3042, i_13_3043, i_13_3044, i_13_3045, i_13_3046, i_13_3047, i_13_3048, i_13_3049, i_13_3050, i_13_3051, i_13_3052, i_13_3053, i_13_3054, i_13_3055, i_13_3056, i_13_3057, i_13_3058, i_13_3059, i_13_3060, i_13_3061, i_13_3062, i_13_3063, i_13_3064, i_13_3065, i_13_3066, i_13_3067, i_13_3068, i_13_3069, i_13_3070, i_13_3071, i_13_3072, i_13_3073, i_13_3074, i_13_3075, i_13_3076, i_13_3077, i_13_3078, i_13_3079, i_13_3080, i_13_3081, i_13_3082, i_13_3083, i_13_3084, i_13_3085, i_13_3086, i_13_3087, i_13_3088, i_13_3089, i_13_3090, i_13_3091, i_13_3092, i_13_3093, i_13_3094, i_13_3095, i_13_3096, i_13_3097, i_13_3098, i_13_3099, i_13_3100, i_13_3101, i_13_3102, i_13_3103, i_13_3104, i_13_3105, i_13_3106, i_13_3107, i_13_3108, i_13_3109, i_13_3110, i_13_3111, i_13_3112, i_13_3113, i_13_3114, i_13_3115, i_13_3116, i_13_3117, i_13_3118, i_13_3119, i_13_3120, i_13_3121, i_13_3122, i_13_3123, i_13_3124, i_13_3125, i_13_3126, i_13_3127, i_13_3128, i_13_3129, i_13_3130, i_13_3131, i_13_3132, i_13_3133, i_13_3134, i_13_3135, i_13_3136, i_13_3137, i_13_3138, i_13_3139, i_13_3140, i_13_3141, i_13_3142, i_13_3143, i_13_3144, i_13_3145, i_13_3146, i_13_3147, i_13_3148, i_13_3149, i_13_3150, i_13_3151, i_13_3152, i_13_3153, i_13_3154, i_13_3155, i_13_3156, i_13_3157, i_13_3158, i_13_3159, i_13_3160, i_13_3161, i_13_3162, i_13_3163, i_13_3164, i_13_3165, i_13_3166, i_13_3167, i_13_3168, i_13_3169, i_13_3170, i_13_3171, i_13_3172, i_13_3173, i_13_3174, i_13_3175, i_13_3176, i_13_3177, i_13_3178, i_13_3179, i_13_3180, i_13_3181, i_13_3182, i_13_3183, i_13_3184, i_13_3185, i_13_3186, i_13_3187, i_13_3188, i_13_3189, i_13_3190, i_13_3191, i_13_3192, i_13_3193, i_13_3194, i_13_3195, i_13_3196, i_13_3197, i_13_3198, i_13_3199, i_13_3200, i_13_3201, i_13_3202, i_13_3203, i_13_3204, i_13_3205, i_13_3206, i_13_3207, i_13_3208, i_13_3209, i_13_3210, i_13_3211, i_13_3212, i_13_3213, i_13_3214, i_13_3215, i_13_3216, i_13_3217, i_13_3218, i_13_3219, i_13_3220, i_13_3221, i_13_3222, i_13_3223, i_13_3224, i_13_3225, i_13_3226, i_13_3227, i_13_3228, i_13_3229, i_13_3230, i_13_3231, i_13_3232, i_13_3233, i_13_3234, i_13_3235, i_13_3236, i_13_3237, i_13_3238, i_13_3239, i_13_3240, i_13_3241, i_13_3242, i_13_3243, i_13_3244, i_13_3245, i_13_3246, i_13_3247, i_13_3248, i_13_3249, i_13_3250, i_13_3251, i_13_3252, i_13_3253, i_13_3254, i_13_3255, i_13_3256, i_13_3257, i_13_3258, i_13_3259, i_13_3260, i_13_3261, i_13_3262, i_13_3263, i_13_3264, i_13_3265, i_13_3266, i_13_3267, i_13_3268, i_13_3269, i_13_3270, i_13_3271, i_13_3272, i_13_3273, i_13_3274, i_13_3275, i_13_3276, i_13_3277, i_13_3278, i_13_3279, i_13_3280, i_13_3281, i_13_3282, i_13_3283, i_13_3284, i_13_3285, i_13_3286, i_13_3287, i_13_3288, i_13_3289, i_13_3290, i_13_3291, i_13_3292, i_13_3293, i_13_3294, i_13_3295, i_13_3296, i_13_3297, i_13_3298, i_13_3299, i_13_3300, i_13_3301, i_13_3302, i_13_3303, i_13_3304, i_13_3305, i_13_3306, i_13_3307, i_13_3308, i_13_3309, i_13_3310, i_13_3311, i_13_3312, i_13_3313, i_13_3314, i_13_3315, i_13_3316, i_13_3317, i_13_3318, i_13_3319, i_13_3320, i_13_3321, i_13_3322, i_13_3323, i_13_3324, i_13_3325, i_13_3326, i_13_3327, i_13_3328, i_13_3329, i_13_3330, i_13_3331, i_13_3332, i_13_3333, i_13_3334, i_13_3335, i_13_3336, i_13_3337, i_13_3338, i_13_3339, i_13_3340, i_13_3341, i_13_3342, i_13_3343, i_13_3344, i_13_3345, i_13_3346, i_13_3347, i_13_3348, i_13_3349, i_13_3350, i_13_3351, i_13_3352, i_13_3353, i_13_3354, i_13_3355, i_13_3356, i_13_3357, i_13_3358, i_13_3359, i_13_3360, i_13_3361, i_13_3362, i_13_3363, i_13_3364, i_13_3365, i_13_3366, i_13_3367, i_13_3368, i_13_3369, i_13_3370, i_13_3371, i_13_3372, i_13_3373, i_13_3374, i_13_3375, i_13_3376, i_13_3377, i_13_3378, i_13_3379, i_13_3380, i_13_3381, i_13_3382, i_13_3383, i_13_3384, i_13_3385, i_13_3386, i_13_3387, i_13_3388, i_13_3389, i_13_3390, i_13_3391, i_13_3392, i_13_3393, i_13_3394, i_13_3395, i_13_3396, i_13_3397, i_13_3398, i_13_3399, i_13_3400, i_13_3401, i_13_3402, i_13_3403, i_13_3404, i_13_3405, i_13_3406, i_13_3407, i_13_3408, i_13_3409, i_13_3410, i_13_3411, i_13_3412, i_13_3413, i_13_3414, i_13_3415, i_13_3416, i_13_3417, i_13_3418, i_13_3419, i_13_3420, i_13_3421, i_13_3422, i_13_3423, i_13_3424, i_13_3425, i_13_3426, i_13_3427, i_13_3428, i_13_3429, i_13_3430, i_13_3431, i_13_3432, i_13_3433, i_13_3434, i_13_3435, i_13_3436, i_13_3437, i_13_3438, i_13_3439, i_13_3440, i_13_3441, i_13_3442, i_13_3443, i_13_3444, i_13_3445, i_13_3446, i_13_3447, i_13_3448, i_13_3449, i_13_3450, i_13_3451, i_13_3452, i_13_3453, i_13_3454, i_13_3455, i_13_3456, i_13_3457, i_13_3458, i_13_3459, i_13_3460, i_13_3461, i_13_3462, i_13_3463, i_13_3464, i_13_3465, i_13_3466, i_13_3467, i_13_3468, i_13_3469, i_13_3470, i_13_3471, i_13_3472, i_13_3473, i_13_3474, i_13_3475, i_13_3476, i_13_3477, i_13_3478, i_13_3479, i_13_3480, i_13_3481, i_13_3482, i_13_3483, i_13_3484, i_13_3485, i_13_3486, i_13_3487, i_13_3488, i_13_3489, i_13_3490, i_13_3491, i_13_3492, i_13_3493, i_13_3494, i_13_3495, i_13_3496, i_13_3497, i_13_3498, i_13_3499, i_13_3500, i_13_3501, i_13_3502, i_13_3503, i_13_3504, i_13_3505, i_13_3506, i_13_3507, i_13_3508, i_13_3509, i_13_3510, i_13_3511, i_13_3512, i_13_3513, i_13_3514, i_13_3515, i_13_3516, i_13_3517, i_13_3518, i_13_3519, i_13_3520, i_13_3521, i_13_3522, i_13_3523, i_13_3524, i_13_3525, i_13_3526, i_13_3527, i_13_3528, i_13_3529, i_13_3530, i_13_3531, i_13_3532, i_13_3533, i_13_3534, i_13_3535, i_13_3536, i_13_3537, i_13_3538, i_13_3539, i_13_3540, i_13_3541, i_13_3542, i_13_3543, i_13_3544, i_13_3545, i_13_3546, i_13_3547, i_13_3548, i_13_3549, i_13_3550, i_13_3551, i_13_3552, i_13_3553, i_13_3554, i_13_3555, i_13_3556, i_13_3557, i_13_3558, i_13_3559, i_13_3560, i_13_3561, i_13_3562, i_13_3563, i_13_3564, i_13_3565, i_13_3566, i_13_3567, i_13_3568, i_13_3569, i_13_3570, i_13_3571, i_13_3572, i_13_3573, i_13_3574, i_13_3575, i_13_3576, i_13_3577, i_13_3578, i_13_3579, i_13_3580, i_13_3581, i_13_3582, i_13_3583, i_13_3584, i_13_3585, i_13_3586, i_13_3587, i_13_3588, i_13_3589, i_13_3590, i_13_3591, i_13_3592, i_13_3593, i_13_3594, i_13_3595, i_13_3596, i_13_3597, i_13_3598, i_13_3599, i_13_3600, i_13_3601, i_13_3602, i_13_3603, i_13_3604, i_13_3605, i_13_3606, i_13_3607, i_13_3608, i_13_3609, i_13_3610, i_13_3611, i_13_3612, i_13_3613, i_13_3614, i_13_3615, i_13_3616, i_13_3617, i_13_3618, i_13_3619, i_13_3620, i_13_3621, i_13_3622, i_13_3623, i_13_3624, i_13_3625, i_13_3626, i_13_3627, i_13_3628, i_13_3629, i_13_3630, i_13_3631, i_13_3632, i_13_3633, i_13_3634, i_13_3635, i_13_3636, i_13_3637, i_13_3638, i_13_3639, i_13_3640, i_13_3641, i_13_3642, i_13_3643, i_13_3644, i_13_3645, i_13_3646, i_13_3647, i_13_3648, i_13_3649, i_13_3650, i_13_3651, i_13_3652, i_13_3653, i_13_3654, i_13_3655, i_13_3656, i_13_3657, i_13_3658, i_13_3659, i_13_3660, i_13_3661, i_13_3662, i_13_3663, i_13_3664, i_13_3665, i_13_3666, i_13_3667, i_13_3668, i_13_3669, i_13_3670, i_13_3671, i_13_3672, i_13_3673, i_13_3674, i_13_3675, i_13_3676, i_13_3677, i_13_3678, i_13_3679, i_13_3680, i_13_3681, i_13_3682, i_13_3683, i_13_3684, i_13_3685, i_13_3686, i_13_3687, i_13_3688, i_13_3689, i_13_3690, i_13_3691, i_13_3692, i_13_3693, i_13_3694, i_13_3695, i_13_3696, i_13_3697, i_13_3698, i_13_3699, i_13_3700, i_13_3701, i_13_3702, i_13_3703, i_13_3704, i_13_3705, i_13_3706, i_13_3707, i_13_3708, i_13_3709, i_13_3710, i_13_3711, i_13_3712, i_13_3713, i_13_3714, i_13_3715, i_13_3716, i_13_3717, i_13_3718, i_13_3719, i_13_3720, i_13_3721, i_13_3722, i_13_3723, i_13_3724, i_13_3725, i_13_3726, i_13_3727, i_13_3728, i_13_3729, i_13_3730, i_13_3731, i_13_3732, i_13_3733, i_13_3734, i_13_3735, i_13_3736, i_13_3737, i_13_3738, i_13_3739, i_13_3740, i_13_3741, i_13_3742, i_13_3743, i_13_3744, i_13_3745, i_13_3746, i_13_3747, i_13_3748, i_13_3749, i_13_3750, i_13_3751, i_13_3752, i_13_3753, i_13_3754, i_13_3755, i_13_3756, i_13_3757, i_13_3758, i_13_3759, i_13_3760, i_13_3761, i_13_3762, i_13_3763, i_13_3764, i_13_3765, i_13_3766, i_13_3767, i_13_3768, i_13_3769, i_13_3770, i_13_3771, i_13_3772, i_13_3773, i_13_3774, i_13_3775, i_13_3776, i_13_3777, i_13_3778, i_13_3779, i_13_3780, i_13_3781, i_13_3782, i_13_3783, i_13_3784, i_13_3785, i_13_3786, i_13_3787, i_13_3788, i_13_3789, i_13_3790, i_13_3791, i_13_3792, i_13_3793, i_13_3794, i_13_3795, i_13_3796, i_13_3797, i_13_3798, i_13_3799, i_13_3800, i_13_3801, i_13_3802, i_13_3803, i_13_3804, i_13_3805, i_13_3806, i_13_3807, i_13_3808, i_13_3809, i_13_3810, i_13_3811, i_13_3812, i_13_3813, i_13_3814, i_13_3815, i_13_3816, i_13_3817, i_13_3818, i_13_3819, i_13_3820, i_13_3821, i_13_3822, i_13_3823, i_13_3824, i_13_3825, i_13_3826, i_13_3827, i_13_3828, i_13_3829, i_13_3830, i_13_3831, i_13_3832, i_13_3833, i_13_3834, i_13_3835, i_13_3836, i_13_3837, i_13_3838, i_13_3839, i_13_3840, i_13_3841, i_13_3842, i_13_3843, i_13_3844, i_13_3845, i_13_3846, i_13_3847, i_13_3848, i_13_3849, i_13_3850, i_13_3851, i_13_3852, i_13_3853, i_13_3854, i_13_3855, i_13_3856, i_13_3857, i_13_3858, i_13_3859, i_13_3860, i_13_3861, i_13_3862, i_13_3863, i_13_3864, i_13_3865, i_13_3866, i_13_3867, i_13_3868, i_13_3869, i_13_3870, i_13_3871, i_13_3872, i_13_3873, i_13_3874, i_13_3875, i_13_3876, i_13_3877, i_13_3878, i_13_3879, i_13_3880, i_13_3881, i_13_3882, i_13_3883, i_13_3884, i_13_3885, i_13_3886, i_13_3887, i_13_3888, i_13_3889, i_13_3890, i_13_3891, i_13_3892, i_13_3893, i_13_3894, i_13_3895, i_13_3896, i_13_3897, i_13_3898, i_13_3899, i_13_3900, i_13_3901, i_13_3902, i_13_3903, i_13_3904, i_13_3905, i_13_3906, i_13_3907, i_13_3908, i_13_3909, i_13_3910, i_13_3911, i_13_3912, i_13_3913, i_13_3914, i_13_3915, i_13_3916, i_13_3917, i_13_3918, i_13_3919, i_13_3920, i_13_3921, i_13_3922, i_13_3923, i_13_3924, i_13_3925, i_13_3926, i_13_3927, i_13_3928, i_13_3929, i_13_3930, i_13_3931, i_13_3932, i_13_3933, i_13_3934, i_13_3935, i_13_3936, i_13_3937, i_13_3938, i_13_3939, i_13_3940, i_13_3941, i_13_3942, i_13_3943, i_13_3944, i_13_3945, i_13_3946, i_13_3947, i_13_3948, i_13_3949, i_13_3950, i_13_3951, i_13_3952, i_13_3953, i_13_3954, i_13_3955, i_13_3956, i_13_3957, i_13_3958, i_13_3959, i_13_3960, i_13_3961, i_13_3962, i_13_3963, i_13_3964, i_13_3965, i_13_3966, i_13_3967, i_13_3968, i_13_3969, i_13_3970, i_13_3971, i_13_3972, i_13_3973, i_13_3974, i_13_3975, i_13_3976, i_13_3977, i_13_3978, i_13_3979, i_13_3980, i_13_3981, i_13_3982, i_13_3983, i_13_3984, i_13_3985, i_13_3986, i_13_3987, i_13_3988, i_13_3989, i_13_3990, i_13_3991, i_13_3992, i_13_3993, i_13_3994, i_13_3995, i_13_3996, i_13_3997, i_13_3998, i_13_3999, i_13_4000, i_13_4001, i_13_4002, i_13_4003, i_13_4004, i_13_4005, i_13_4006, i_13_4007, i_13_4008, i_13_4009, i_13_4010, i_13_4011, i_13_4012, i_13_4013, i_13_4014, i_13_4015, i_13_4016, i_13_4017, i_13_4018, i_13_4019, i_13_4020, i_13_4021, i_13_4022, i_13_4023, i_13_4024, i_13_4025, i_13_4026, i_13_4027, i_13_4028, i_13_4029, i_13_4030, i_13_4031, i_13_4032, i_13_4033, i_13_4034, i_13_4035, i_13_4036, i_13_4037, i_13_4038, i_13_4039, i_13_4040, i_13_4041, i_13_4042, i_13_4043, i_13_4044, i_13_4045, i_13_4046, i_13_4047, i_13_4048, i_13_4049, i_13_4050, i_13_4051, i_13_4052, i_13_4053, i_13_4054, i_13_4055, i_13_4056, i_13_4057, i_13_4058, i_13_4059, i_13_4060, i_13_4061, i_13_4062, i_13_4063, i_13_4064, i_13_4065, i_13_4066, i_13_4067, i_13_4068, i_13_4069, i_13_4070, i_13_4071, i_13_4072, i_13_4073, i_13_4074, i_13_4075, i_13_4076, i_13_4077, i_13_4078, i_13_4079, i_13_4080, i_13_4081, i_13_4082, i_13_4083, i_13_4084, i_13_4085, i_13_4086, i_13_4087, i_13_4088, i_13_4089, i_13_4090, i_13_4091, i_13_4092, i_13_4093, i_13_4094, i_13_4095, i_13_4096, i_13_4097, i_13_4098, i_13_4099, i_13_4100, i_13_4101, i_13_4102, i_13_4103, i_13_4104, i_13_4105, i_13_4106, i_13_4107, i_13_4108, i_13_4109, i_13_4110, i_13_4111, i_13_4112, i_13_4113, i_13_4114, i_13_4115, i_13_4116, i_13_4117, i_13_4118, i_13_4119, i_13_4120, i_13_4121, i_13_4122, i_13_4123, i_13_4124, i_13_4125, i_13_4126, i_13_4127, i_13_4128, i_13_4129, i_13_4130, i_13_4131, i_13_4132, i_13_4133, i_13_4134, i_13_4135, i_13_4136, i_13_4137, i_13_4138, i_13_4139, i_13_4140, i_13_4141, i_13_4142, i_13_4143, i_13_4144, i_13_4145, i_13_4146, i_13_4147, i_13_4148, i_13_4149, i_13_4150, i_13_4151, i_13_4152, i_13_4153, i_13_4154, i_13_4155, i_13_4156, i_13_4157, i_13_4158, i_13_4159, i_13_4160, i_13_4161, i_13_4162, i_13_4163, i_13_4164, i_13_4165, i_13_4166, i_13_4167, i_13_4168, i_13_4169, i_13_4170, i_13_4171, i_13_4172, i_13_4173, i_13_4174, i_13_4175, i_13_4176, i_13_4177, i_13_4178, i_13_4179, i_13_4180, i_13_4181, i_13_4182, i_13_4183, i_13_4184, i_13_4185, i_13_4186, i_13_4187, i_13_4188, i_13_4189, i_13_4190, i_13_4191, i_13_4192, i_13_4193, i_13_4194, i_13_4195, i_13_4196, i_13_4197, i_13_4198, i_13_4199, i_13_4200, i_13_4201, i_13_4202, i_13_4203, i_13_4204, i_13_4205, i_13_4206, i_13_4207, i_13_4208, i_13_4209, i_13_4210, i_13_4211, i_13_4212, i_13_4213, i_13_4214, i_13_4215, i_13_4216, i_13_4217, i_13_4218, i_13_4219, i_13_4220, i_13_4221, i_13_4222, i_13_4223, i_13_4224, i_13_4225, i_13_4226, i_13_4227, i_13_4228, i_13_4229, i_13_4230, i_13_4231, i_13_4232, i_13_4233, i_13_4234, i_13_4235, i_13_4236, i_13_4237, i_13_4238, i_13_4239, i_13_4240, i_13_4241, i_13_4242, i_13_4243, i_13_4244, i_13_4245, i_13_4246, i_13_4247, i_13_4248, i_13_4249, i_13_4250, i_13_4251, i_13_4252, i_13_4253, i_13_4254, i_13_4255, i_13_4256, i_13_4257, i_13_4258, i_13_4259, i_13_4260, i_13_4261, i_13_4262, i_13_4263, i_13_4264, i_13_4265, i_13_4266, i_13_4267, i_13_4268, i_13_4269, i_13_4270, i_13_4271, i_13_4272, i_13_4273, i_13_4274, i_13_4275, i_13_4276, i_13_4277, i_13_4278, i_13_4279, i_13_4280, i_13_4281, i_13_4282, i_13_4283, i_13_4284, i_13_4285, i_13_4286, i_13_4287, i_13_4288, i_13_4289, i_13_4290, i_13_4291, i_13_4292, i_13_4293, i_13_4294, i_13_4295, i_13_4296, i_13_4297, i_13_4298, i_13_4299, i_13_4300, i_13_4301, i_13_4302, i_13_4303, i_13_4304, i_13_4305, i_13_4306, i_13_4307, i_13_4308, i_13_4309, i_13_4310, i_13_4311, i_13_4312, i_13_4313, i_13_4314, i_13_4315, i_13_4316, i_13_4317, i_13_4318, i_13_4319, i_13_4320, i_13_4321, i_13_4322, i_13_4323, i_13_4324, i_13_4325, i_13_4326, i_13_4327, i_13_4328, i_13_4329, i_13_4330, i_13_4331, i_13_4332, i_13_4333, i_13_4334, i_13_4335, i_13_4336, i_13_4337, i_13_4338, i_13_4339, i_13_4340, i_13_4341, i_13_4342, i_13_4343, i_13_4344, i_13_4345, i_13_4346, i_13_4347, i_13_4348, i_13_4349, i_13_4350, i_13_4351, i_13_4352, i_13_4353, i_13_4354, i_13_4355, i_13_4356, i_13_4357, i_13_4358, i_13_4359, i_13_4360, i_13_4361, i_13_4362, i_13_4363, i_13_4364, i_13_4365, i_13_4366, i_13_4367, i_13_4368, i_13_4369, i_13_4370, i_13_4371, i_13_4372, i_13_4373, i_13_4374, i_13_4375, i_13_4376, i_13_4377, i_13_4378, i_13_4379, i_13_4380, i_13_4381, i_13_4382, i_13_4383, i_13_4384, i_13_4385, i_13_4386, i_13_4387, i_13_4388, i_13_4389, i_13_4390, i_13_4391, i_13_4392, i_13_4393, i_13_4394, i_13_4395, i_13_4396, i_13_4397, i_13_4398, i_13_4399, i_13_4400, i_13_4401, i_13_4402, i_13_4403, i_13_4404, i_13_4405, i_13_4406, i_13_4407, i_13_4408, i_13_4409, i_13_4410, i_13_4411, i_13_4412, i_13_4413, i_13_4414, i_13_4415, i_13_4416, i_13_4417, i_13_4418, i_13_4419, i_13_4420, i_13_4421, i_13_4422, i_13_4423, i_13_4424, i_13_4425, i_13_4426, i_13_4427, i_13_4428, i_13_4429, i_13_4430, i_13_4431, i_13_4432, i_13_4433, i_13_4434, i_13_4435, i_13_4436, i_13_4437, i_13_4438, i_13_4439, i_13_4440, i_13_4441, i_13_4442, i_13_4443, i_13_4444, i_13_4445, i_13_4446, i_13_4447, i_13_4448, i_13_4449, i_13_4450, i_13_4451, i_13_4452, i_13_4453, i_13_4454, i_13_4455, i_13_4456, i_13_4457, i_13_4458, i_13_4459, i_13_4460, i_13_4461, i_13_4462, i_13_4463, i_13_4464, i_13_4465, i_13_4466, i_13_4467, i_13_4468, i_13_4469, i_13_4470, i_13_4471, i_13_4472, i_13_4473, i_13_4474, i_13_4475, i_13_4476, i_13_4477, i_13_4478, i_13_4479, i_13_4480, i_13_4481, i_13_4482, i_13_4483, i_13_4484, i_13_4485, i_13_4486, i_13_4487, i_13_4488, i_13_4489, i_13_4490, i_13_4491, i_13_4492, i_13_4493, i_13_4494, i_13_4495, i_13_4496, i_13_4497, i_13_4498, i_13_4499, i_13_4500, i_13_4501, i_13_4502, i_13_4503, i_13_4504, i_13_4505, i_13_4506, i_13_4507, i_13_4508, i_13_4509, i_13_4510, i_13_4511, i_13_4512, i_13_4513, i_13_4514, i_13_4515, i_13_4516, i_13_4517, i_13_4518, i_13_4519, i_13_4520, i_13_4521, i_13_4522, i_13_4523, i_13_4524, i_13_4525, i_13_4526, i_13_4527, i_13_4528, i_13_4529, i_13_4530, i_13_4531, i_13_4532, i_13_4533, i_13_4534, i_13_4535, i_13_4536, i_13_4537, i_13_4538, i_13_4539, i_13_4540, i_13_4541, i_13_4542, i_13_4543, i_13_4544, i_13_4545, i_13_4546, i_13_4547, i_13_4548, i_13_4549, i_13_4550, i_13_4551, i_13_4552, i_13_4553, i_13_4554, i_13_4555, i_13_4556, i_13_4557, i_13_4558, i_13_4559, i_13_4560, i_13_4561, i_13_4562, i_13_4563, i_13_4564, i_13_4565, i_13_4566, i_13_4567, i_13_4568, i_13_4569, i_13_4570, i_13_4571, i_13_4572, i_13_4573, i_13_4574, i_13_4575, i_13_4576, i_13_4577, i_13_4578, i_13_4579, i_13_4580, i_13_4581, i_13_4582, i_13_4583, i_13_4584, i_13_4585, i_13_4586, i_13_4587, i_13_4588, i_13_4589, i_13_4590, i_13_4591, i_13_4592, i_13_4593, i_13_4594, i_13_4595, i_13_4596, i_13_4597, i_13_4598, i_13_4599, i_13_4600, i_13_4601, i_13_4602, i_13_4603, i_13_4604, i_13_4605, i_13_4606, i_13_4607, o_13_0, o_13_1, o_13_2, o_13_3, o_13_4, o_13_5, o_13_6, o_13_7, o_13_8, o_13_9, o_13_10, o_13_11, o_13_12, o_13_13, o_13_14, o_13_15, o_13_16, o_13_17, o_13_18, o_13_19, o_13_20, o_13_21, o_13_22, o_13_23, o_13_24, o_13_25, o_13_26, o_13_27, o_13_28, o_13_29, o_13_30, o_13_31, o_13_32, o_13_33, o_13_34, o_13_35, o_13_36, o_13_37, o_13_38, o_13_39, o_13_40, o_13_41, o_13_42, o_13_43, o_13_44, o_13_45, o_13_46, o_13_47, o_13_48, o_13_49, o_13_50, o_13_51, o_13_52, o_13_53, o_13_54, o_13_55, o_13_56, o_13_57, o_13_58, o_13_59, o_13_60, o_13_61, o_13_62, o_13_63, o_13_64, o_13_65, o_13_66, o_13_67, o_13_68, o_13_69, o_13_70, o_13_71, o_13_72, o_13_73, o_13_74, o_13_75, o_13_76, o_13_77, o_13_78, o_13_79, o_13_80, o_13_81, o_13_82, o_13_83, o_13_84, o_13_85, o_13_86, o_13_87, o_13_88, o_13_89, o_13_90, o_13_91, o_13_92, o_13_93, o_13_94, o_13_95, o_13_96, o_13_97, o_13_98, o_13_99, o_13_100, o_13_101, o_13_102, o_13_103, o_13_104, o_13_105, o_13_106, o_13_107, o_13_108, o_13_109, o_13_110, o_13_111, o_13_112, o_13_113, o_13_114, o_13_115, o_13_116, o_13_117, o_13_118, o_13_119, o_13_120, o_13_121, o_13_122, o_13_123, o_13_124, o_13_125, o_13_126, o_13_127, o_13_128, o_13_129, o_13_130, o_13_131, o_13_132, o_13_133, o_13_134, o_13_135, o_13_136, o_13_137, o_13_138, o_13_139, o_13_140, o_13_141, o_13_142, o_13_143, o_13_144, o_13_145, o_13_146, o_13_147, o_13_148, o_13_149, o_13_150, o_13_151, o_13_152, o_13_153, o_13_154, o_13_155, o_13_156, o_13_157, o_13_158, o_13_159, o_13_160, o_13_161, o_13_162, o_13_163, o_13_164, o_13_165, o_13_166, o_13_167, o_13_168, o_13_169, o_13_170, o_13_171, o_13_172, o_13_173, o_13_174, o_13_175, o_13_176, o_13_177, o_13_178, o_13_179, o_13_180, o_13_181, o_13_182, o_13_183, o_13_184, o_13_185, o_13_186, o_13_187, o_13_188, o_13_189, o_13_190, o_13_191, o_13_192, o_13_193, o_13_194, o_13_195, o_13_196, o_13_197, o_13_198, o_13_199, o_13_200, o_13_201, o_13_202, o_13_203, o_13_204, o_13_205, o_13_206, o_13_207, o_13_208, o_13_209, o_13_210, o_13_211, o_13_212, o_13_213, o_13_214, o_13_215, o_13_216, o_13_217, o_13_218, o_13_219, o_13_220, o_13_221, o_13_222, o_13_223, o_13_224, o_13_225, o_13_226, o_13_227, o_13_228, o_13_229, o_13_230, o_13_231, o_13_232, o_13_233, o_13_234, o_13_235, o_13_236, o_13_237, o_13_238, o_13_239, o_13_240, o_13_241, o_13_242, o_13_243, o_13_244, o_13_245, o_13_246, o_13_247, o_13_248, o_13_249, o_13_250, o_13_251, o_13_252, o_13_253, o_13_254, o_13_255, o_13_256, o_13_257, o_13_258, o_13_259, o_13_260, o_13_261, o_13_262, o_13_263, o_13_264, o_13_265, o_13_266, o_13_267, o_13_268, o_13_269, o_13_270, o_13_271, o_13_272, o_13_273, o_13_274, o_13_275, o_13_276, o_13_277, o_13_278, o_13_279, o_13_280, o_13_281, o_13_282, o_13_283, o_13_284, o_13_285, o_13_286, o_13_287, o_13_288, o_13_289, o_13_290, o_13_291, o_13_292, o_13_293, o_13_294, o_13_295, o_13_296, o_13_297, o_13_298, o_13_299, o_13_300, o_13_301, o_13_302, o_13_303, o_13_304, o_13_305, o_13_306, o_13_307, o_13_308, o_13_309, o_13_310, o_13_311, o_13_312, o_13_313, o_13_314, o_13_315, o_13_316, o_13_317, o_13_318, o_13_319, o_13_320, o_13_321, o_13_322, o_13_323, o_13_324, o_13_325, o_13_326, o_13_327, o_13_328, o_13_329, o_13_330, o_13_331, o_13_332, o_13_333, o_13_334, o_13_335, o_13_336, o_13_337, o_13_338, o_13_339, o_13_340, o_13_341, o_13_342, o_13_343, o_13_344, o_13_345, o_13_346, o_13_347, o_13_348, o_13_349, o_13_350, o_13_351, o_13_352, o_13_353, o_13_354, o_13_355, o_13_356, o_13_357, o_13_358, o_13_359, o_13_360, o_13_361, o_13_362, o_13_363, o_13_364, o_13_365, o_13_366, o_13_367, o_13_368, o_13_369, o_13_370, o_13_371, o_13_372, o_13_373, o_13_374, o_13_375, o_13_376, o_13_377, o_13_378, o_13_379, o_13_380, o_13_381, o_13_382, o_13_383, o_13_384, o_13_385, o_13_386, o_13_387, o_13_388, o_13_389, o_13_390, o_13_391, o_13_392, o_13_393, o_13_394, o_13_395, o_13_396, o_13_397, o_13_398, o_13_399, o_13_400, o_13_401, o_13_402, o_13_403, o_13_404, o_13_405, o_13_406, o_13_407, o_13_408, o_13_409, o_13_410, o_13_411, o_13_412, o_13_413, o_13_414, o_13_415, o_13_416, o_13_417, o_13_418, o_13_419, o_13_420, o_13_421, o_13_422, o_13_423, o_13_424, o_13_425, o_13_426, o_13_427, o_13_428, o_13_429, o_13_430, o_13_431, o_13_432, o_13_433, o_13_434, o_13_435, o_13_436, o_13_437, o_13_438, o_13_439, o_13_440, o_13_441, o_13_442, o_13_443, o_13_444, o_13_445, o_13_446, o_13_447, o_13_448, o_13_449, o_13_450, o_13_451, o_13_452, o_13_453, o_13_454, o_13_455, o_13_456, o_13_457, o_13_458, o_13_459, o_13_460, o_13_461, o_13_462, o_13_463, o_13_464, o_13_465, o_13_466, o_13_467, o_13_468, o_13_469, o_13_470, o_13_471, o_13_472, o_13_473, o_13_474, o_13_475, o_13_476, o_13_477, o_13_478, o_13_479, o_13_480, o_13_481, o_13_482, o_13_483, o_13_484, o_13_485, o_13_486, o_13_487, o_13_488, o_13_489, o_13_490, o_13_491, o_13_492, o_13_493, o_13_494, o_13_495, o_13_496, o_13_497, o_13_498, o_13_499, o_13_500, o_13_501, o_13_502, o_13_503, o_13_504, o_13_505, o_13_506, o_13_507, o_13_508, o_13_509, o_13_510, o_13_511);
input i_13_0, i_13_1, i_13_2, i_13_3, i_13_4, i_13_5, i_13_6, i_13_7, i_13_8, i_13_9, i_13_10, i_13_11, i_13_12, i_13_13, i_13_14, i_13_15, i_13_16, i_13_17, i_13_18, i_13_19, i_13_20, i_13_21, i_13_22, i_13_23, i_13_24, i_13_25, i_13_26, i_13_27, i_13_28, i_13_29, i_13_30, i_13_31, i_13_32, i_13_33, i_13_34, i_13_35, i_13_36, i_13_37, i_13_38, i_13_39, i_13_40, i_13_41, i_13_42, i_13_43, i_13_44, i_13_45, i_13_46, i_13_47, i_13_48, i_13_49, i_13_50, i_13_51, i_13_52, i_13_53, i_13_54, i_13_55, i_13_56, i_13_57, i_13_58, i_13_59, i_13_60, i_13_61, i_13_62, i_13_63, i_13_64, i_13_65, i_13_66, i_13_67, i_13_68, i_13_69, i_13_70, i_13_71, i_13_72, i_13_73, i_13_74, i_13_75, i_13_76, i_13_77, i_13_78, i_13_79, i_13_80, i_13_81, i_13_82, i_13_83, i_13_84, i_13_85, i_13_86, i_13_87, i_13_88, i_13_89, i_13_90, i_13_91, i_13_92, i_13_93, i_13_94, i_13_95, i_13_96, i_13_97, i_13_98, i_13_99, i_13_100, i_13_101, i_13_102, i_13_103, i_13_104, i_13_105, i_13_106, i_13_107, i_13_108, i_13_109, i_13_110, i_13_111, i_13_112, i_13_113, i_13_114, i_13_115, i_13_116, i_13_117, i_13_118, i_13_119, i_13_120, i_13_121, i_13_122, i_13_123, i_13_124, i_13_125, i_13_126, i_13_127, i_13_128, i_13_129, i_13_130, i_13_131, i_13_132, i_13_133, i_13_134, i_13_135, i_13_136, i_13_137, i_13_138, i_13_139, i_13_140, i_13_141, i_13_142, i_13_143, i_13_144, i_13_145, i_13_146, i_13_147, i_13_148, i_13_149, i_13_150, i_13_151, i_13_152, i_13_153, i_13_154, i_13_155, i_13_156, i_13_157, i_13_158, i_13_159, i_13_160, i_13_161, i_13_162, i_13_163, i_13_164, i_13_165, i_13_166, i_13_167, i_13_168, i_13_169, i_13_170, i_13_171, i_13_172, i_13_173, i_13_174, i_13_175, i_13_176, i_13_177, i_13_178, i_13_179, i_13_180, i_13_181, i_13_182, i_13_183, i_13_184, i_13_185, i_13_186, i_13_187, i_13_188, i_13_189, i_13_190, i_13_191, i_13_192, i_13_193, i_13_194, i_13_195, i_13_196, i_13_197, i_13_198, i_13_199, i_13_200, i_13_201, i_13_202, i_13_203, i_13_204, i_13_205, i_13_206, i_13_207, i_13_208, i_13_209, i_13_210, i_13_211, i_13_212, i_13_213, i_13_214, i_13_215, i_13_216, i_13_217, i_13_218, i_13_219, i_13_220, i_13_221, i_13_222, i_13_223, i_13_224, i_13_225, i_13_226, i_13_227, i_13_228, i_13_229, i_13_230, i_13_231, i_13_232, i_13_233, i_13_234, i_13_235, i_13_236, i_13_237, i_13_238, i_13_239, i_13_240, i_13_241, i_13_242, i_13_243, i_13_244, i_13_245, i_13_246, i_13_247, i_13_248, i_13_249, i_13_250, i_13_251, i_13_252, i_13_253, i_13_254, i_13_255, i_13_256, i_13_257, i_13_258, i_13_259, i_13_260, i_13_261, i_13_262, i_13_263, i_13_264, i_13_265, i_13_266, i_13_267, i_13_268, i_13_269, i_13_270, i_13_271, i_13_272, i_13_273, i_13_274, i_13_275, i_13_276, i_13_277, i_13_278, i_13_279, i_13_280, i_13_281, i_13_282, i_13_283, i_13_284, i_13_285, i_13_286, i_13_287, i_13_288, i_13_289, i_13_290, i_13_291, i_13_292, i_13_293, i_13_294, i_13_295, i_13_296, i_13_297, i_13_298, i_13_299, i_13_300, i_13_301, i_13_302, i_13_303, i_13_304, i_13_305, i_13_306, i_13_307, i_13_308, i_13_309, i_13_310, i_13_311, i_13_312, i_13_313, i_13_314, i_13_315, i_13_316, i_13_317, i_13_318, i_13_319, i_13_320, i_13_321, i_13_322, i_13_323, i_13_324, i_13_325, i_13_326, i_13_327, i_13_328, i_13_329, i_13_330, i_13_331, i_13_332, i_13_333, i_13_334, i_13_335, i_13_336, i_13_337, i_13_338, i_13_339, i_13_340, i_13_341, i_13_342, i_13_343, i_13_344, i_13_345, i_13_346, i_13_347, i_13_348, i_13_349, i_13_350, i_13_351, i_13_352, i_13_353, i_13_354, i_13_355, i_13_356, i_13_357, i_13_358, i_13_359, i_13_360, i_13_361, i_13_362, i_13_363, i_13_364, i_13_365, i_13_366, i_13_367, i_13_368, i_13_369, i_13_370, i_13_371, i_13_372, i_13_373, i_13_374, i_13_375, i_13_376, i_13_377, i_13_378, i_13_379, i_13_380, i_13_381, i_13_382, i_13_383, i_13_384, i_13_385, i_13_386, i_13_387, i_13_388, i_13_389, i_13_390, i_13_391, i_13_392, i_13_393, i_13_394, i_13_395, i_13_396, i_13_397, i_13_398, i_13_399, i_13_400, i_13_401, i_13_402, i_13_403, i_13_404, i_13_405, i_13_406, i_13_407, i_13_408, i_13_409, i_13_410, i_13_411, i_13_412, i_13_413, i_13_414, i_13_415, i_13_416, i_13_417, i_13_418, i_13_419, i_13_420, i_13_421, i_13_422, i_13_423, i_13_424, i_13_425, i_13_426, i_13_427, i_13_428, i_13_429, i_13_430, i_13_431, i_13_432, i_13_433, i_13_434, i_13_435, i_13_436, i_13_437, i_13_438, i_13_439, i_13_440, i_13_441, i_13_442, i_13_443, i_13_444, i_13_445, i_13_446, i_13_447, i_13_448, i_13_449, i_13_450, i_13_451, i_13_452, i_13_453, i_13_454, i_13_455, i_13_456, i_13_457, i_13_458, i_13_459, i_13_460, i_13_461, i_13_462, i_13_463, i_13_464, i_13_465, i_13_466, i_13_467, i_13_468, i_13_469, i_13_470, i_13_471, i_13_472, i_13_473, i_13_474, i_13_475, i_13_476, i_13_477, i_13_478, i_13_479, i_13_480, i_13_481, i_13_482, i_13_483, i_13_484, i_13_485, i_13_486, i_13_487, i_13_488, i_13_489, i_13_490, i_13_491, i_13_492, i_13_493, i_13_494, i_13_495, i_13_496, i_13_497, i_13_498, i_13_499, i_13_500, i_13_501, i_13_502, i_13_503, i_13_504, i_13_505, i_13_506, i_13_507, i_13_508, i_13_509, i_13_510, i_13_511, i_13_512, i_13_513, i_13_514, i_13_515, i_13_516, i_13_517, i_13_518, i_13_519, i_13_520, i_13_521, i_13_522, i_13_523, i_13_524, i_13_525, i_13_526, i_13_527, i_13_528, i_13_529, i_13_530, i_13_531, i_13_532, i_13_533, i_13_534, i_13_535, i_13_536, i_13_537, i_13_538, i_13_539, i_13_540, i_13_541, i_13_542, i_13_543, i_13_544, i_13_545, i_13_546, i_13_547, i_13_548, i_13_549, i_13_550, i_13_551, i_13_552, i_13_553, i_13_554, i_13_555, i_13_556, i_13_557, i_13_558, i_13_559, i_13_560, i_13_561, i_13_562, i_13_563, i_13_564, i_13_565, i_13_566, i_13_567, i_13_568, i_13_569, i_13_570, i_13_571, i_13_572, i_13_573, i_13_574, i_13_575, i_13_576, i_13_577, i_13_578, i_13_579, i_13_580, i_13_581, i_13_582, i_13_583, i_13_584, i_13_585, i_13_586, i_13_587, i_13_588, i_13_589, i_13_590, i_13_591, i_13_592, i_13_593, i_13_594, i_13_595, i_13_596, i_13_597, i_13_598, i_13_599, i_13_600, i_13_601, i_13_602, i_13_603, i_13_604, i_13_605, i_13_606, i_13_607, i_13_608, i_13_609, i_13_610, i_13_611, i_13_612, i_13_613, i_13_614, i_13_615, i_13_616, i_13_617, i_13_618, i_13_619, i_13_620, i_13_621, i_13_622, i_13_623, i_13_624, i_13_625, i_13_626, i_13_627, i_13_628, i_13_629, i_13_630, i_13_631, i_13_632, i_13_633, i_13_634, i_13_635, i_13_636, i_13_637, i_13_638, i_13_639, i_13_640, i_13_641, i_13_642, i_13_643, i_13_644, i_13_645, i_13_646, i_13_647, i_13_648, i_13_649, i_13_650, i_13_651, i_13_652, i_13_653, i_13_654, i_13_655, i_13_656, i_13_657, i_13_658, i_13_659, i_13_660, i_13_661, i_13_662, i_13_663, i_13_664, i_13_665, i_13_666, i_13_667, i_13_668, i_13_669, i_13_670, i_13_671, i_13_672, i_13_673, i_13_674, i_13_675, i_13_676, i_13_677, i_13_678, i_13_679, i_13_680, i_13_681, i_13_682, i_13_683, i_13_684, i_13_685, i_13_686, i_13_687, i_13_688, i_13_689, i_13_690, i_13_691, i_13_692, i_13_693, i_13_694, i_13_695, i_13_696, i_13_697, i_13_698, i_13_699, i_13_700, i_13_701, i_13_702, i_13_703, i_13_704, i_13_705, i_13_706, i_13_707, i_13_708, i_13_709, i_13_710, i_13_711, i_13_712, i_13_713, i_13_714, i_13_715, i_13_716, i_13_717, i_13_718, i_13_719, i_13_720, i_13_721, i_13_722, i_13_723, i_13_724, i_13_725, i_13_726, i_13_727, i_13_728, i_13_729, i_13_730, i_13_731, i_13_732, i_13_733, i_13_734, i_13_735, i_13_736, i_13_737, i_13_738, i_13_739, i_13_740, i_13_741, i_13_742, i_13_743, i_13_744, i_13_745, i_13_746, i_13_747, i_13_748, i_13_749, i_13_750, i_13_751, i_13_752, i_13_753, i_13_754, i_13_755, i_13_756, i_13_757, i_13_758, i_13_759, i_13_760, i_13_761, i_13_762, i_13_763, i_13_764, i_13_765, i_13_766, i_13_767, i_13_768, i_13_769, i_13_770, i_13_771, i_13_772, i_13_773, i_13_774, i_13_775, i_13_776, i_13_777, i_13_778, i_13_779, i_13_780, i_13_781, i_13_782, i_13_783, i_13_784, i_13_785, i_13_786, i_13_787, i_13_788, i_13_789, i_13_790, i_13_791, i_13_792, i_13_793, i_13_794, i_13_795, i_13_796, i_13_797, i_13_798, i_13_799, i_13_800, i_13_801, i_13_802, i_13_803, i_13_804, i_13_805, i_13_806, i_13_807, i_13_808, i_13_809, i_13_810, i_13_811, i_13_812, i_13_813, i_13_814, i_13_815, i_13_816, i_13_817, i_13_818, i_13_819, i_13_820, i_13_821, i_13_822, i_13_823, i_13_824, i_13_825, i_13_826, i_13_827, i_13_828, i_13_829, i_13_830, i_13_831, i_13_832, i_13_833, i_13_834, i_13_835, i_13_836, i_13_837, i_13_838, i_13_839, i_13_840, i_13_841, i_13_842, i_13_843, i_13_844, i_13_845, i_13_846, i_13_847, i_13_848, i_13_849, i_13_850, i_13_851, i_13_852, i_13_853, i_13_854, i_13_855, i_13_856, i_13_857, i_13_858, i_13_859, i_13_860, i_13_861, i_13_862, i_13_863, i_13_864, i_13_865, i_13_866, i_13_867, i_13_868, i_13_869, i_13_870, i_13_871, i_13_872, i_13_873, i_13_874, i_13_875, i_13_876, i_13_877, i_13_878, i_13_879, i_13_880, i_13_881, i_13_882, i_13_883, i_13_884, i_13_885, i_13_886, i_13_887, i_13_888, i_13_889, i_13_890, i_13_891, i_13_892, i_13_893, i_13_894, i_13_895, i_13_896, i_13_897, i_13_898, i_13_899, i_13_900, i_13_901, i_13_902, i_13_903, i_13_904, i_13_905, i_13_906, i_13_907, i_13_908, i_13_909, i_13_910, i_13_911, i_13_912, i_13_913, i_13_914, i_13_915, i_13_916, i_13_917, i_13_918, i_13_919, i_13_920, i_13_921, i_13_922, i_13_923, i_13_924, i_13_925, i_13_926, i_13_927, i_13_928, i_13_929, i_13_930, i_13_931, i_13_932, i_13_933, i_13_934, i_13_935, i_13_936, i_13_937, i_13_938, i_13_939, i_13_940, i_13_941, i_13_942, i_13_943, i_13_944, i_13_945, i_13_946, i_13_947, i_13_948, i_13_949, i_13_950, i_13_951, i_13_952, i_13_953, i_13_954, i_13_955, i_13_956, i_13_957, i_13_958, i_13_959, i_13_960, i_13_961, i_13_962, i_13_963, i_13_964, i_13_965, i_13_966, i_13_967, i_13_968, i_13_969, i_13_970, i_13_971, i_13_972, i_13_973, i_13_974, i_13_975, i_13_976, i_13_977, i_13_978, i_13_979, i_13_980, i_13_981, i_13_982, i_13_983, i_13_984, i_13_985, i_13_986, i_13_987, i_13_988, i_13_989, i_13_990, i_13_991, i_13_992, i_13_993, i_13_994, i_13_995, i_13_996, i_13_997, i_13_998, i_13_999, i_13_1000, i_13_1001, i_13_1002, i_13_1003, i_13_1004, i_13_1005, i_13_1006, i_13_1007, i_13_1008, i_13_1009, i_13_1010, i_13_1011, i_13_1012, i_13_1013, i_13_1014, i_13_1015, i_13_1016, i_13_1017, i_13_1018, i_13_1019, i_13_1020, i_13_1021, i_13_1022, i_13_1023, i_13_1024, i_13_1025, i_13_1026, i_13_1027, i_13_1028, i_13_1029, i_13_1030, i_13_1031, i_13_1032, i_13_1033, i_13_1034, i_13_1035, i_13_1036, i_13_1037, i_13_1038, i_13_1039, i_13_1040, i_13_1041, i_13_1042, i_13_1043, i_13_1044, i_13_1045, i_13_1046, i_13_1047, i_13_1048, i_13_1049, i_13_1050, i_13_1051, i_13_1052, i_13_1053, i_13_1054, i_13_1055, i_13_1056, i_13_1057, i_13_1058, i_13_1059, i_13_1060, i_13_1061, i_13_1062, i_13_1063, i_13_1064, i_13_1065, i_13_1066, i_13_1067, i_13_1068, i_13_1069, i_13_1070, i_13_1071, i_13_1072, i_13_1073, i_13_1074, i_13_1075, i_13_1076, i_13_1077, i_13_1078, i_13_1079, i_13_1080, i_13_1081, i_13_1082, i_13_1083, i_13_1084, i_13_1085, i_13_1086, i_13_1087, i_13_1088, i_13_1089, i_13_1090, i_13_1091, i_13_1092, i_13_1093, i_13_1094, i_13_1095, i_13_1096, i_13_1097, i_13_1098, i_13_1099, i_13_1100, i_13_1101, i_13_1102, i_13_1103, i_13_1104, i_13_1105, i_13_1106, i_13_1107, i_13_1108, i_13_1109, i_13_1110, i_13_1111, i_13_1112, i_13_1113, i_13_1114, i_13_1115, i_13_1116, i_13_1117, i_13_1118, i_13_1119, i_13_1120, i_13_1121, i_13_1122, i_13_1123, i_13_1124, i_13_1125, i_13_1126, i_13_1127, i_13_1128, i_13_1129, i_13_1130, i_13_1131, i_13_1132, i_13_1133, i_13_1134, i_13_1135, i_13_1136, i_13_1137, i_13_1138, i_13_1139, i_13_1140, i_13_1141, i_13_1142, i_13_1143, i_13_1144, i_13_1145, i_13_1146, i_13_1147, i_13_1148, i_13_1149, i_13_1150, i_13_1151, i_13_1152, i_13_1153, i_13_1154, i_13_1155, i_13_1156, i_13_1157, i_13_1158, i_13_1159, i_13_1160, i_13_1161, i_13_1162, i_13_1163, i_13_1164, i_13_1165, i_13_1166, i_13_1167, i_13_1168, i_13_1169, i_13_1170, i_13_1171, i_13_1172, i_13_1173, i_13_1174, i_13_1175, i_13_1176, i_13_1177, i_13_1178, i_13_1179, i_13_1180, i_13_1181, i_13_1182, i_13_1183, i_13_1184, i_13_1185, i_13_1186, i_13_1187, i_13_1188, i_13_1189, i_13_1190, i_13_1191, i_13_1192, i_13_1193, i_13_1194, i_13_1195, i_13_1196, i_13_1197, i_13_1198, i_13_1199, i_13_1200, i_13_1201, i_13_1202, i_13_1203, i_13_1204, i_13_1205, i_13_1206, i_13_1207, i_13_1208, i_13_1209, i_13_1210, i_13_1211, i_13_1212, i_13_1213, i_13_1214, i_13_1215, i_13_1216, i_13_1217, i_13_1218, i_13_1219, i_13_1220, i_13_1221, i_13_1222, i_13_1223, i_13_1224, i_13_1225, i_13_1226, i_13_1227, i_13_1228, i_13_1229, i_13_1230, i_13_1231, i_13_1232, i_13_1233, i_13_1234, i_13_1235, i_13_1236, i_13_1237, i_13_1238, i_13_1239, i_13_1240, i_13_1241, i_13_1242, i_13_1243, i_13_1244, i_13_1245, i_13_1246, i_13_1247, i_13_1248, i_13_1249, i_13_1250, i_13_1251, i_13_1252, i_13_1253, i_13_1254, i_13_1255, i_13_1256, i_13_1257, i_13_1258, i_13_1259, i_13_1260, i_13_1261, i_13_1262, i_13_1263, i_13_1264, i_13_1265, i_13_1266, i_13_1267, i_13_1268, i_13_1269, i_13_1270, i_13_1271, i_13_1272, i_13_1273, i_13_1274, i_13_1275, i_13_1276, i_13_1277, i_13_1278, i_13_1279, i_13_1280, i_13_1281, i_13_1282, i_13_1283, i_13_1284, i_13_1285, i_13_1286, i_13_1287, i_13_1288, i_13_1289, i_13_1290, i_13_1291, i_13_1292, i_13_1293, i_13_1294, i_13_1295, i_13_1296, i_13_1297, i_13_1298, i_13_1299, i_13_1300, i_13_1301, i_13_1302, i_13_1303, i_13_1304, i_13_1305, i_13_1306, i_13_1307, i_13_1308, i_13_1309, i_13_1310, i_13_1311, i_13_1312, i_13_1313, i_13_1314, i_13_1315, i_13_1316, i_13_1317, i_13_1318, i_13_1319, i_13_1320, i_13_1321, i_13_1322, i_13_1323, i_13_1324, i_13_1325, i_13_1326, i_13_1327, i_13_1328, i_13_1329, i_13_1330, i_13_1331, i_13_1332, i_13_1333, i_13_1334, i_13_1335, i_13_1336, i_13_1337, i_13_1338, i_13_1339, i_13_1340, i_13_1341, i_13_1342, i_13_1343, i_13_1344, i_13_1345, i_13_1346, i_13_1347, i_13_1348, i_13_1349, i_13_1350, i_13_1351, i_13_1352, i_13_1353, i_13_1354, i_13_1355, i_13_1356, i_13_1357, i_13_1358, i_13_1359, i_13_1360, i_13_1361, i_13_1362, i_13_1363, i_13_1364, i_13_1365, i_13_1366, i_13_1367, i_13_1368, i_13_1369, i_13_1370, i_13_1371, i_13_1372, i_13_1373, i_13_1374, i_13_1375, i_13_1376, i_13_1377, i_13_1378, i_13_1379, i_13_1380, i_13_1381, i_13_1382, i_13_1383, i_13_1384, i_13_1385, i_13_1386, i_13_1387, i_13_1388, i_13_1389, i_13_1390, i_13_1391, i_13_1392, i_13_1393, i_13_1394, i_13_1395, i_13_1396, i_13_1397, i_13_1398, i_13_1399, i_13_1400, i_13_1401, i_13_1402, i_13_1403, i_13_1404, i_13_1405, i_13_1406, i_13_1407, i_13_1408, i_13_1409, i_13_1410, i_13_1411, i_13_1412, i_13_1413, i_13_1414, i_13_1415, i_13_1416, i_13_1417, i_13_1418, i_13_1419, i_13_1420, i_13_1421, i_13_1422, i_13_1423, i_13_1424, i_13_1425, i_13_1426, i_13_1427, i_13_1428, i_13_1429, i_13_1430, i_13_1431, i_13_1432, i_13_1433, i_13_1434, i_13_1435, i_13_1436, i_13_1437, i_13_1438, i_13_1439, i_13_1440, i_13_1441, i_13_1442, i_13_1443, i_13_1444, i_13_1445, i_13_1446, i_13_1447, i_13_1448, i_13_1449, i_13_1450, i_13_1451, i_13_1452, i_13_1453, i_13_1454, i_13_1455, i_13_1456, i_13_1457, i_13_1458, i_13_1459, i_13_1460, i_13_1461, i_13_1462, i_13_1463, i_13_1464, i_13_1465, i_13_1466, i_13_1467, i_13_1468, i_13_1469, i_13_1470, i_13_1471, i_13_1472, i_13_1473, i_13_1474, i_13_1475, i_13_1476, i_13_1477, i_13_1478, i_13_1479, i_13_1480, i_13_1481, i_13_1482, i_13_1483, i_13_1484, i_13_1485, i_13_1486, i_13_1487, i_13_1488, i_13_1489, i_13_1490, i_13_1491, i_13_1492, i_13_1493, i_13_1494, i_13_1495, i_13_1496, i_13_1497, i_13_1498, i_13_1499, i_13_1500, i_13_1501, i_13_1502, i_13_1503, i_13_1504, i_13_1505, i_13_1506, i_13_1507, i_13_1508, i_13_1509, i_13_1510, i_13_1511, i_13_1512, i_13_1513, i_13_1514, i_13_1515, i_13_1516, i_13_1517, i_13_1518, i_13_1519, i_13_1520, i_13_1521, i_13_1522, i_13_1523, i_13_1524, i_13_1525, i_13_1526, i_13_1527, i_13_1528, i_13_1529, i_13_1530, i_13_1531, i_13_1532, i_13_1533, i_13_1534, i_13_1535, i_13_1536, i_13_1537, i_13_1538, i_13_1539, i_13_1540, i_13_1541, i_13_1542, i_13_1543, i_13_1544, i_13_1545, i_13_1546, i_13_1547, i_13_1548, i_13_1549, i_13_1550, i_13_1551, i_13_1552, i_13_1553, i_13_1554, i_13_1555, i_13_1556, i_13_1557, i_13_1558, i_13_1559, i_13_1560, i_13_1561, i_13_1562, i_13_1563, i_13_1564, i_13_1565, i_13_1566, i_13_1567, i_13_1568, i_13_1569, i_13_1570, i_13_1571, i_13_1572, i_13_1573, i_13_1574, i_13_1575, i_13_1576, i_13_1577, i_13_1578, i_13_1579, i_13_1580, i_13_1581, i_13_1582, i_13_1583, i_13_1584, i_13_1585, i_13_1586, i_13_1587, i_13_1588, i_13_1589, i_13_1590, i_13_1591, i_13_1592, i_13_1593, i_13_1594, i_13_1595, i_13_1596, i_13_1597, i_13_1598, i_13_1599, i_13_1600, i_13_1601, i_13_1602, i_13_1603, i_13_1604, i_13_1605, i_13_1606, i_13_1607, i_13_1608, i_13_1609, i_13_1610, i_13_1611, i_13_1612, i_13_1613, i_13_1614, i_13_1615, i_13_1616, i_13_1617, i_13_1618, i_13_1619, i_13_1620, i_13_1621, i_13_1622, i_13_1623, i_13_1624, i_13_1625, i_13_1626, i_13_1627, i_13_1628, i_13_1629, i_13_1630, i_13_1631, i_13_1632, i_13_1633, i_13_1634, i_13_1635, i_13_1636, i_13_1637, i_13_1638, i_13_1639, i_13_1640, i_13_1641, i_13_1642, i_13_1643, i_13_1644, i_13_1645, i_13_1646, i_13_1647, i_13_1648, i_13_1649, i_13_1650, i_13_1651, i_13_1652, i_13_1653, i_13_1654, i_13_1655, i_13_1656, i_13_1657, i_13_1658, i_13_1659, i_13_1660, i_13_1661, i_13_1662, i_13_1663, i_13_1664, i_13_1665, i_13_1666, i_13_1667, i_13_1668, i_13_1669, i_13_1670, i_13_1671, i_13_1672, i_13_1673, i_13_1674, i_13_1675, i_13_1676, i_13_1677, i_13_1678, i_13_1679, i_13_1680, i_13_1681, i_13_1682, i_13_1683, i_13_1684, i_13_1685, i_13_1686, i_13_1687, i_13_1688, i_13_1689, i_13_1690, i_13_1691, i_13_1692, i_13_1693, i_13_1694, i_13_1695, i_13_1696, i_13_1697, i_13_1698, i_13_1699, i_13_1700, i_13_1701, i_13_1702, i_13_1703, i_13_1704, i_13_1705, i_13_1706, i_13_1707, i_13_1708, i_13_1709, i_13_1710, i_13_1711, i_13_1712, i_13_1713, i_13_1714, i_13_1715, i_13_1716, i_13_1717, i_13_1718, i_13_1719, i_13_1720, i_13_1721, i_13_1722, i_13_1723, i_13_1724, i_13_1725, i_13_1726, i_13_1727, i_13_1728, i_13_1729, i_13_1730, i_13_1731, i_13_1732, i_13_1733, i_13_1734, i_13_1735, i_13_1736, i_13_1737, i_13_1738, i_13_1739, i_13_1740, i_13_1741, i_13_1742, i_13_1743, i_13_1744, i_13_1745, i_13_1746, i_13_1747, i_13_1748, i_13_1749, i_13_1750, i_13_1751, i_13_1752, i_13_1753, i_13_1754, i_13_1755, i_13_1756, i_13_1757, i_13_1758, i_13_1759, i_13_1760, i_13_1761, i_13_1762, i_13_1763, i_13_1764, i_13_1765, i_13_1766, i_13_1767, i_13_1768, i_13_1769, i_13_1770, i_13_1771, i_13_1772, i_13_1773, i_13_1774, i_13_1775, i_13_1776, i_13_1777, i_13_1778, i_13_1779, i_13_1780, i_13_1781, i_13_1782, i_13_1783, i_13_1784, i_13_1785, i_13_1786, i_13_1787, i_13_1788, i_13_1789, i_13_1790, i_13_1791, i_13_1792, i_13_1793, i_13_1794, i_13_1795, i_13_1796, i_13_1797, i_13_1798, i_13_1799, i_13_1800, i_13_1801, i_13_1802, i_13_1803, i_13_1804, i_13_1805, i_13_1806, i_13_1807, i_13_1808, i_13_1809, i_13_1810, i_13_1811, i_13_1812, i_13_1813, i_13_1814, i_13_1815, i_13_1816, i_13_1817, i_13_1818, i_13_1819, i_13_1820, i_13_1821, i_13_1822, i_13_1823, i_13_1824, i_13_1825, i_13_1826, i_13_1827, i_13_1828, i_13_1829, i_13_1830, i_13_1831, i_13_1832, i_13_1833, i_13_1834, i_13_1835, i_13_1836, i_13_1837, i_13_1838, i_13_1839, i_13_1840, i_13_1841, i_13_1842, i_13_1843, i_13_1844, i_13_1845, i_13_1846, i_13_1847, i_13_1848, i_13_1849, i_13_1850, i_13_1851, i_13_1852, i_13_1853, i_13_1854, i_13_1855, i_13_1856, i_13_1857, i_13_1858, i_13_1859, i_13_1860, i_13_1861, i_13_1862, i_13_1863, i_13_1864, i_13_1865, i_13_1866, i_13_1867, i_13_1868, i_13_1869, i_13_1870, i_13_1871, i_13_1872, i_13_1873, i_13_1874, i_13_1875, i_13_1876, i_13_1877, i_13_1878, i_13_1879, i_13_1880, i_13_1881, i_13_1882, i_13_1883, i_13_1884, i_13_1885, i_13_1886, i_13_1887, i_13_1888, i_13_1889, i_13_1890, i_13_1891, i_13_1892, i_13_1893, i_13_1894, i_13_1895, i_13_1896, i_13_1897, i_13_1898, i_13_1899, i_13_1900, i_13_1901, i_13_1902, i_13_1903, i_13_1904, i_13_1905, i_13_1906, i_13_1907, i_13_1908, i_13_1909, i_13_1910, i_13_1911, i_13_1912, i_13_1913, i_13_1914, i_13_1915, i_13_1916, i_13_1917, i_13_1918, i_13_1919, i_13_1920, i_13_1921, i_13_1922, i_13_1923, i_13_1924, i_13_1925, i_13_1926, i_13_1927, i_13_1928, i_13_1929, i_13_1930, i_13_1931, i_13_1932, i_13_1933, i_13_1934, i_13_1935, i_13_1936, i_13_1937, i_13_1938, i_13_1939, i_13_1940, i_13_1941, i_13_1942, i_13_1943, i_13_1944, i_13_1945, i_13_1946, i_13_1947, i_13_1948, i_13_1949, i_13_1950, i_13_1951, i_13_1952, i_13_1953, i_13_1954, i_13_1955, i_13_1956, i_13_1957, i_13_1958, i_13_1959, i_13_1960, i_13_1961, i_13_1962, i_13_1963, i_13_1964, i_13_1965, i_13_1966, i_13_1967, i_13_1968, i_13_1969, i_13_1970, i_13_1971, i_13_1972, i_13_1973, i_13_1974, i_13_1975, i_13_1976, i_13_1977, i_13_1978, i_13_1979, i_13_1980, i_13_1981, i_13_1982, i_13_1983, i_13_1984, i_13_1985, i_13_1986, i_13_1987, i_13_1988, i_13_1989, i_13_1990, i_13_1991, i_13_1992, i_13_1993, i_13_1994, i_13_1995, i_13_1996, i_13_1997, i_13_1998, i_13_1999, i_13_2000, i_13_2001, i_13_2002, i_13_2003, i_13_2004, i_13_2005, i_13_2006, i_13_2007, i_13_2008, i_13_2009, i_13_2010, i_13_2011, i_13_2012, i_13_2013, i_13_2014, i_13_2015, i_13_2016, i_13_2017, i_13_2018, i_13_2019, i_13_2020, i_13_2021, i_13_2022, i_13_2023, i_13_2024, i_13_2025, i_13_2026, i_13_2027, i_13_2028, i_13_2029, i_13_2030, i_13_2031, i_13_2032, i_13_2033, i_13_2034, i_13_2035, i_13_2036, i_13_2037, i_13_2038, i_13_2039, i_13_2040, i_13_2041, i_13_2042, i_13_2043, i_13_2044, i_13_2045, i_13_2046, i_13_2047, i_13_2048, i_13_2049, i_13_2050, i_13_2051, i_13_2052, i_13_2053, i_13_2054, i_13_2055, i_13_2056, i_13_2057, i_13_2058, i_13_2059, i_13_2060, i_13_2061, i_13_2062, i_13_2063, i_13_2064, i_13_2065, i_13_2066, i_13_2067, i_13_2068, i_13_2069, i_13_2070, i_13_2071, i_13_2072, i_13_2073, i_13_2074, i_13_2075, i_13_2076, i_13_2077, i_13_2078, i_13_2079, i_13_2080, i_13_2081, i_13_2082, i_13_2083, i_13_2084, i_13_2085, i_13_2086, i_13_2087, i_13_2088, i_13_2089, i_13_2090, i_13_2091, i_13_2092, i_13_2093, i_13_2094, i_13_2095, i_13_2096, i_13_2097, i_13_2098, i_13_2099, i_13_2100, i_13_2101, i_13_2102, i_13_2103, i_13_2104, i_13_2105, i_13_2106, i_13_2107, i_13_2108, i_13_2109, i_13_2110, i_13_2111, i_13_2112, i_13_2113, i_13_2114, i_13_2115, i_13_2116, i_13_2117, i_13_2118, i_13_2119, i_13_2120, i_13_2121, i_13_2122, i_13_2123, i_13_2124, i_13_2125, i_13_2126, i_13_2127, i_13_2128, i_13_2129, i_13_2130, i_13_2131, i_13_2132, i_13_2133, i_13_2134, i_13_2135, i_13_2136, i_13_2137, i_13_2138, i_13_2139, i_13_2140, i_13_2141, i_13_2142, i_13_2143, i_13_2144, i_13_2145, i_13_2146, i_13_2147, i_13_2148, i_13_2149, i_13_2150, i_13_2151, i_13_2152, i_13_2153, i_13_2154, i_13_2155, i_13_2156, i_13_2157, i_13_2158, i_13_2159, i_13_2160, i_13_2161, i_13_2162, i_13_2163, i_13_2164, i_13_2165, i_13_2166, i_13_2167, i_13_2168, i_13_2169, i_13_2170, i_13_2171, i_13_2172, i_13_2173, i_13_2174, i_13_2175, i_13_2176, i_13_2177, i_13_2178, i_13_2179, i_13_2180, i_13_2181, i_13_2182, i_13_2183, i_13_2184, i_13_2185, i_13_2186, i_13_2187, i_13_2188, i_13_2189, i_13_2190, i_13_2191, i_13_2192, i_13_2193, i_13_2194, i_13_2195, i_13_2196, i_13_2197, i_13_2198, i_13_2199, i_13_2200, i_13_2201, i_13_2202, i_13_2203, i_13_2204, i_13_2205, i_13_2206, i_13_2207, i_13_2208, i_13_2209, i_13_2210, i_13_2211, i_13_2212, i_13_2213, i_13_2214, i_13_2215, i_13_2216, i_13_2217, i_13_2218, i_13_2219, i_13_2220, i_13_2221, i_13_2222, i_13_2223, i_13_2224, i_13_2225, i_13_2226, i_13_2227, i_13_2228, i_13_2229, i_13_2230, i_13_2231, i_13_2232, i_13_2233, i_13_2234, i_13_2235, i_13_2236, i_13_2237, i_13_2238, i_13_2239, i_13_2240, i_13_2241, i_13_2242, i_13_2243, i_13_2244, i_13_2245, i_13_2246, i_13_2247, i_13_2248, i_13_2249, i_13_2250, i_13_2251, i_13_2252, i_13_2253, i_13_2254, i_13_2255, i_13_2256, i_13_2257, i_13_2258, i_13_2259, i_13_2260, i_13_2261, i_13_2262, i_13_2263, i_13_2264, i_13_2265, i_13_2266, i_13_2267, i_13_2268, i_13_2269, i_13_2270, i_13_2271, i_13_2272, i_13_2273, i_13_2274, i_13_2275, i_13_2276, i_13_2277, i_13_2278, i_13_2279, i_13_2280, i_13_2281, i_13_2282, i_13_2283, i_13_2284, i_13_2285, i_13_2286, i_13_2287, i_13_2288, i_13_2289, i_13_2290, i_13_2291, i_13_2292, i_13_2293, i_13_2294, i_13_2295, i_13_2296, i_13_2297, i_13_2298, i_13_2299, i_13_2300, i_13_2301, i_13_2302, i_13_2303, i_13_2304, i_13_2305, i_13_2306, i_13_2307, i_13_2308, i_13_2309, i_13_2310, i_13_2311, i_13_2312, i_13_2313, i_13_2314, i_13_2315, i_13_2316, i_13_2317, i_13_2318, i_13_2319, i_13_2320, i_13_2321, i_13_2322, i_13_2323, i_13_2324, i_13_2325, i_13_2326, i_13_2327, i_13_2328, i_13_2329, i_13_2330, i_13_2331, i_13_2332, i_13_2333, i_13_2334, i_13_2335, i_13_2336, i_13_2337, i_13_2338, i_13_2339, i_13_2340, i_13_2341, i_13_2342, i_13_2343, i_13_2344, i_13_2345, i_13_2346, i_13_2347, i_13_2348, i_13_2349, i_13_2350, i_13_2351, i_13_2352, i_13_2353, i_13_2354, i_13_2355, i_13_2356, i_13_2357, i_13_2358, i_13_2359, i_13_2360, i_13_2361, i_13_2362, i_13_2363, i_13_2364, i_13_2365, i_13_2366, i_13_2367, i_13_2368, i_13_2369, i_13_2370, i_13_2371, i_13_2372, i_13_2373, i_13_2374, i_13_2375, i_13_2376, i_13_2377, i_13_2378, i_13_2379, i_13_2380, i_13_2381, i_13_2382, i_13_2383, i_13_2384, i_13_2385, i_13_2386, i_13_2387, i_13_2388, i_13_2389, i_13_2390, i_13_2391, i_13_2392, i_13_2393, i_13_2394, i_13_2395, i_13_2396, i_13_2397, i_13_2398, i_13_2399, i_13_2400, i_13_2401, i_13_2402, i_13_2403, i_13_2404, i_13_2405, i_13_2406, i_13_2407, i_13_2408, i_13_2409, i_13_2410, i_13_2411, i_13_2412, i_13_2413, i_13_2414, i_13_2415, i_13_2416, i_13_2417, i_13_2418, i_13_2419, i_13_2420, i_13_2421, i_13_2422, i_13_2423, i_13_2424, i_13_2425, i_13_2426, i_13_2427, i_13_2428, i_13_2429, i_13_2430, i_13_2431, i_13_2432, i_13_2433, i_13_2434, i_13_2435, i_13_2436, i_13_2437, i_13_2438, i_13_2439, i_13_2440, i_13_2441, i_13_2442, i_13_2443, i_13_2444, i_13_2445, i_13_2446, i_13_2447, i_13_2448, i_13_2449, i_13_2450, i_13_2451, i_13_2452, i_13_2453, i_13_2454, i_13_2455, i_13_2456, i_13_2457, i_13_2458, i_13_2459, i_13_2460, i_13_2461, i_13_2462, i_13_2463, i_13_2464, i_13_2465, i_13_2466, i_13_2467, i_13_2468, i_13_2469, i_13_2470, i_13_2471, i_13_2472, i_13_2473, i_13_2474, i_13_2475, i_13_2476, i_13_2477, i_13_2478, i_13_2479, i_13_2480, i_13_2481, i_13_2482, i_13_2483, i_13_2484, i_13_2485, i_13_2486, i_13_2487, i_13_2488, i_13_2489, i_13_2490, i_13_2491, i_13_2492, i_13_2493, i_13_2494, i_13_2495, i_13_2496, i_13_2497, i_13_2498, i_13_2499, i_13_2500, i_13_2501, i_13_2502, i_13_2503, i_13_2504, i_13_2505, i_13_2506, i_13_2507, i_13_2508, i_13_2509, i_13_2510, i_13_2511, i_13_2512, i_13_2513, i_13_2514, i_13_2515, i_13_2516, i_13_2517, i_13_2518, i_13_2519, i_13_2520, i_13_2521, i_13_2522, i_13_2523, i_13_2524, i_13_2525, i_13_2526, i_13_2527, i_13_2528, i_13_2529, i_13_2530, i_13_2531, i_13_2532, i_13_2533, i_13_2534, i_13_2535, i_13_2536, i_13_2537, i_13_2538, i_13_2539, i_13_2540, i_13_2541, i_13_2542, i_13_2543, i_13_2544, i_13_2545, i_13_2546, i_13_2547, i_13_2548, i_13_2549, i_13_2550, i_13_2551, i_13_2552, i_13_2553, i_13_2554, i_13_2555, i_13_2556, i_13_2557, i_13_2558, i_13_2559, i_13_2560, i_13_2561, i_13_2562, i_13_2563, i_13_2564, i_13_2565, i_13_2566, i_13_2567, i_13_2568, i_13_2569, i_13_2570, i_13_2571, i_13_2572, i_13_2573, i_13_2574, i_13_2575, i_13_2576, i_13_2577, i_13_2578, i_13_2579, i_13_2580, i_13_2581, i_13_2582, i_13_2583, i_13_2584, i_13_2585, i_13_2586, i_13_2587, i_13_2588, i_13_2589, i_13_2590, i_13_2591, i_13_2592, i_13_2593, i_13_2594, i_13_2595, i_13_2596, i_13_2597, i_13_2598, i_13_2599, i_13_2600, i_13_2601, i_13_2602, i_13_2603, i_13_2604, i_13_2605, i_13_2606, i_13_2607, i_13_2608, i_13_2609, i_13_2610, i_13_2611, i_13_2612, i_13_2613, i_13_2614, i_13_2615, i_13_2616, i_13_2617, i_13_2618, i_13_2619, i_13_2620, i_13_2621, i_13_2622, i_13_2623, i_13_2624, i_13_2625, i_13_2626, i_13_2627, i_13_2628, i_13_2629, i_13_2630, i_13_2631, i_13_2632, i_13_2633, i_13_2634, i_13_2635, i_13_2636, i_13_2637, i_13_2638, i_13_2639, i_13_2640, i_13_2641, i_13_2642, i_13_2643, i_13_2644, i_13_2645, i_13_2646, i_13_2647, i_13_2648, i_13_2649, i_13_2650, i_13_2651, i_13_2652, i_13_2653, i_13_2654, i_13_2655, i_13_2656, i_13_2657, i_13_2658, i_13_2659, i_13_2660, i_13_2661, i_13_2662, i_13_2663, i_13_2664, i_13_2665, i_13_2666, i_13_2667, i_13_2668, i_13_2669, i_13_2670, i_13_2671, i_13_2672, i_13_2673, i_13_2674, i_13_2675, i_13_2676, i_13_2677, i_13_2678, i_13_2679, i_13_2680, i_13_2681, i_13_2682, i_13_2683, i_13_2684, i_13_2685, i_13_2686, i_13_2687, i_13_2688, i_13_2689, i_13_2690, i_13_2691, i_13_2692, i_13_2693, i_13_2694, i_13_2695, i_13_2696, i_13_2697, i_13_2698, i_13_2699, i_13_2700, i_13_2701, i_13_2702, i_13_2703, i_13_2704, i_13_2705, i_13_2706, i_13_2707, i_13_2708, i_13_2709, i_13_2710, i_13_2711, i_13_2712, i_13_2713, i_13_2714, i_13_2715, i_13_2716, i_13_2717, i_13_2718, i_13_2719, i_13_2720, i_13_2721, i_13_2722, i_13_2723, i_13_2724, i_13_2725, i_13_2726, i_13_2727, i_13_2728, i_13_2729, i_13_2730, i_13_2731, i_13_2732, i_13_2733, i_13_2734, i_13_2735, i_13_2736, i_13_2737, i_13_2738, i_13_2739, i_13_2740, i_13_2741, i_13_2742, i_13_2743, i_13_2744, i_13_2745, i_13_2746, i_13_2747, i_13_2748, i_13_2749, i_13_2750, i_13_2751, i_13_2752, i_13_2753, i_13_2754, i_13_2755, i_13_2756, i_13_2757, i_13_2758, i_13_2759, i_13_2760, i_13_2761, i_13_2762, i_13_2763, i_13_2764, i_13_2765, i_13_2766, i_13_2767, i_13_2768, i_13_2769, i_13_2770, i_13_2771, i_13_2772, i_13_2773, i_13_2774, i_13_2775, i_13_2776, i_13_2777, i_13_2778, i_13_2779, i_13_2780, i_13_2781, i_13_2782, i_13_2783, i_13_2784, i_13_2785, i_13_2786, i_13_2787, i_13_2788, i_13_2789, i_13_2790, i_13_2791, i_13_2792, i_13_2793, i_13_2794, i_13_2795, i_13_2796, i_13_2797, i_13_2798, i_13_2799, i_13_2800, i_13_2801, i_13_2802, i_13_2803, i_13_2804, i_13_2805, i_13_2806, i_13_2807, i_13_2808, i_13_2809, i_13_2810, i_13_2811, i_13_2812, i_13_2813, i_13_2814, i_13_2815, i_13_2816, i_13_2817, i_13_2818, i_13_2819, i_13_2820, i_13_2821, i_13_2822, i_13_2823, i_13_2824, i_13_2825, i_13_2826, i_13_2827, i_13_2828, i_13_2829, i_13_2830, i_13_2831, i_13_2832, i_13_2833, i_13_2834, i_13_2835, i_13_2836, i_13_2837, i_13_2838, i_13_2839, i_13_2840, i_13_2841, i_13_2842, i_13_2843, i_13_2844, i_13_2845, i_13_2846, i_13_2847, i_13_2848, i_13_2849, i_13_2850, i_13_2851, i_13_2852, i_13_2853, i_13_2854, i_13_2855, i_13_2856, i_13_2857, i_13_2858, i_13_2859, i_13_2860, i_13_2861, i_13_2862, i_13_2863, i_13_2864, i_13_2865, i_13_2866, i_13_2867, i_13_2868, i_13_2869, i_13_2870, i_13_2871, i_13_2872, i_13_2873, i_13_2874, i_13_2875, i_13_2876, i_13_2877, i_13_2878, i_13_2879, i_13_2880, i_13_2881, i_13_2882, i_13_2883, i_13_2884, i_13_2885, i_13_2886, i_13_2887, i_13_2888, i_13_2889, i_13_2890, i_13_2891, i_13_2892, i_13_2893, i_13_2894, i_13_2895, i_13_2896, i_13_2897, i_13_2898, i_13_2899, i_13_2900, i_13_2901, i_13_2902, i_13_2903, i_13_2904, i_13_2905, i_13_2906, i_13_2907, i_13_2908, i_13_2909, i_13_2910, i_13_2911, i_13_2912, i_13_2913, i_13_2914, i_13_2915, i_13_2916, i_13_2917, i_13_2918, i_13_2919, i_13_2920, i_13_2921, i_13_2922, i_13_2923, i_13_2924, i_13_2925, i_13_2926, i_13_2927, i_13_2928, i_13_2929, i_13_2930, i_13_2931, i_13_2932, i_13_2933, i_13_2934, i_13_2935, i_13_2936, i_13_2937, i_13_2938, i_13_2939, i_13_2940, i_13_2941, i_13_2942, i_13_2943, i_13_2944, i_13_2945, i_13_2946, i_13_2947, i_13_2948, i_13_2949, i_13_2950, i_13_2951, i_13_2952, i_13_2953, i_13_2954, i_13_2955, i_13_2956, i_13_2957, i_13_2958, i_13_2959, i_13_2960, i_13_2961, i_13_2962, i_13_2963, i_13_2964, i_13_2965, i_13_2966, i_13_2967, i_13_2968, i_13_2969, i_13_2970, i_13_2971, i_13_2972, i_13_2973, i_13_2974, i_13_2975, i_13_2976, i_13_2977, i_13_2978, i_13_2979, i_13_2980, i_13_2981, i_13_2982, i_13_2983, i_13_2984, i_13_2985, i_13_2986, i_13_2987, i_13_2988, i_13_2989, i_13_2990, i_13_2991, i_13_2992, i_13_2993, i_13_2994, i_13_2995, i_13_2996, i_13_2997, i_13_2998, i_13_2999, i_13_3000, i_13_3001, i_13_3002, i_13_3003, i_13_3004, i_13_3005, i_13_3006, i_13_3007, i_13_3008, i_13_3009, i_13_3010, i_13_3011, i_13_3012, i_13_3013, i_13_3014, i_13_3015, i_13_3016, i_13_3017, i_13_3018, i_13_3019, i_13_3020, i_13_3021, i_13_3022, i_13_3023, i_13_3024, i_13_3025, i_13_3026, i_13_3027, i_13_3028, i_13_3029, i_13_3030, i_13_3031, i_13_3032, i_13_3033, i_13_3034, i_13_3035, i_13_3036, i_13_3037, i_13_3038, i_13_3039, i_13_3040, i_13_3041, i_13_3042, i_13_3043, i_13_3044, i_13_3045, i_13_3046, i_13_3047, i_13_3048, i_13_3049, i_13_3050, i_13_3051, i_13_3052, i_13_3053, i_13_3054, i_13_3055, i_13_3056, i_13_3057, i_13_3058, i_13_3059, i_13_3060, i_13_3061, i_13_3062, i_13_3063, i_13_3064, i_13_3065, i_13_3066, i_13_3067, i_13_3068, i_13_3069, i_13_3070, i_13_3071, i_13_3072, i_13_3073, i_13_3074, i_13_3075, i_13_3076, i_13_3077, i_13_3078, i_13_3079, i_13_3080, i_13_3081, i_13_3082, i_13_3083, i_13_3084, i_13_3085, i_13_3086, i_13_3087, i_13_3088, i_13_3089, i_13_3090, i_13_3091, i_13_3092, i_13_3093, i_13_3094, i_13_3095, i_13_3096, i_13_3097, i_13_3098, i_13_3099, i_13_3100, i_13_3101, i_13_3102, i_13_3103, i_13_3104, i_13_3105, i_13_3106, i_13_3107, i_13_3108, i_13_3109, i_13_3110, i_13_3111, i_13_3112, i_13_3113, i_13_3114, i_13_3115, i_13_3116, i_13_3117, i_13_3118, i_13_3119, i_13_3120, i_13_3121, i_13_3122, i_13_3123, i_13_3124, i_13_3125, i_13_3126, i_13_3127, i_13_3128, i_13_3129, i_13_3130, i_13_3131, i_13_3132, i_13_3133, i_13_3134, i_13_3135, i_13_3136, i_13_3137, i_13_3138, i_13_3139, i_13_3140, i_13_3141, i_13_3142, i_13_3143, i_13_3144, i_13_3145, i_13_3146, i_13_3147, i_13_3148, i_13_3149, i_13_3150, i_13_3151, i_13_3152, i_13_3153, i_13_3154, i_13_3155, i_13_3156, i_13_3157, i_13_3158, i_13_3159, i_13_3160, i_13_3161, i_13_3162, i_13_3163, i_13_3164, i_13_3165, i_13_3166, i_13_3167, i_13_3168, i_13_3169, i_13_3170, i_13_3171, i_13_3172, i_13_3173, i_13_3174, i_13_3175, i_13_3176, i_13_3177, i_13_3178, i_13_3179, i_13_3180, i_13_3181, i_13_3182, i_13_3183, i_13_3184, i_13_3185, i_13_3186, i_13_3187, i_13_3188, i_13_3189, i_13_3190, i_13_3191, i_13_3192, i_13_3193, i_13_3194, i_13_3195, i_13_3196, i_13_3197, i_13_3198, i_13_3199, i_13_3200, i_13_3201, i_13_3202, i_13_3203, i_13_3204, i_13_3205, i_13_3206, i_13_3207, i_13_3208, i_13_3209, i_13_3210, i_13_3211, i_13_3212, i_13_3213, i_13_3214, i_13_3215, i_13_3216, i_13_3217, i_13_3218, i_13_3219, i_13_3220, i_13_3221, i_13_3222, i_13_3223, i_13_3224, i_13_3225, i_13_3226, i_13_3227, i_13_3228, i_13_3229, i_13_3230, i_13_3231, i_13_3232, i_13_3233, i_13_3234, i_13_3235, i_13_3236, i_13_3237, i_13_3238, i_13_3239, i_13_3240, i_13_3241, i_13_3242, i_13_3243, i_13_3244, i_13_3245, i_13_3246, i_13_3247, i_13_3248, i_13_3249, i_13_3250, i_13_3251, i_13_3252, i_13_3253, i_13_3254, i_13_3255, i_13_3256, i_13_3257, i_13_3258, i_13_3259, i_13_3260, i_13_3261, i_13_3262, i_13_3263, i_13_3264, i_13_3265, i_13_3266, i_13_3267, i_13_3268, i_13_3269, i_13_3270, i_13_3271, i_13_3272, i_13_3273, i_13_3274, i_13_3275, i_13_3276, i_13_3277, i_13_3278, i_13_3279, i_13_3280, i_13_3281, i_13_3282, i_13_3283, i_13_3284, i_13_3285, i_13_3286, i_13_3287, i_13_3288, i_13_3289, i_13_3290, i_13_3291, i_13_3292, i_13_3293, i_13_3294, i_13_3295, i_13_3296, i_13_3297, i_13_3298, i_13_3299, i_13_3300, i_13_3301, i_13_3302, i_13_3303, i_13_3304, i_13_3305, i_13_3306, i_13_3307, i_13_3308, i_13_3309, i_13_3310, i_13_3311, i_13_3312, i_13_3313, i_13_3314, i_13_3315, i_13_3316, i_13_3317, i_13_3318, i_13_3319, i_13_3320, i_13_3321, i_13_3322, i_13_3323, i_13_3324, i_13_3325, i_13_3326, i_13_3327, i_13_3328, i_13_3329, i_13_3330, i_13_3331, i_13_3332, i_13_3333, i_13_3334, i_13_3335, i_13_3336, i_13_3337, i_13_3338, i_13_3339, i_13_3340, i_13_3341, i_13_3342, i_13_3343, i_13_3344, i_13_3345, i_13_3346, i_13_3347, i_13_3348, i_13_3349, i_13_3350, i_13_3351, i_13_3352, i_13_3353, i_13_3354, i_13_3355, i_13_3356, i_13_3357, i_13_3358, i_13_3359, i_13_3360, i_13_3361, i_13_3362, i_13_3363, i_13_3364, i_13_3365, i_13_3366, i_13_3367, i_13_3368, i_13_3369, i_13_3370, i_13_3371, i_13_3372, i_13_3373, i_13_3374, i_13_3375, i_13_3376, i_13_3377, i_13_3378, i_13_3379, i_13_3380, i_13_3381, i_13_3382, i_13_3383, i_13_3384, i_13_3385, i_13_3386, i_13_3387, i_13_3388, i_13_3389, i_13_3390, i_13_3391, i_13_3392, i_13_3393, i_13_3394, i_13_3395, i_13_3396, i_13_3397, i_13_3398, i_13_3399, i_13_3400, i_13_3401, i_13_3402, i_13_3403, i_13_3404, i_13_3405, i_13_3406, i_13_3407, i_13_3408, i_13_3409, i_13_3410, i_13_3411, i_13_3412, i_13_3413, i_13_3414, i_13_3415, i_13_3416, i_13_3417, i_13_3418, i_13_3419, i_13_3420, i_13_3421, i_13_3422, i_13_3423, i_13_3424, i_13_3425, i_13_3426, i_13_3427, i_13_3428, i_13_3429, i_13_3430, i_13_3431, i_13_3432, i_13_3433, i_13_3434, i_13_3435, i_13_3436, i_13_3437, i_13_3438, i_13_3439, i_13_3440, i_13_3441, i_13_3442, i_13_3443, i_13_3444, i_13_3445, i_13_3446, i_13_3447, i_13_3448, i_13_3449, i_13_3450, i_13_3451, i_13_3452, i_13_3453, i_13_3454, i_13_3455, i_13_3456, i_13_3457, i_13_3458, i_13_3459, i_13_3460, i_13_3461, i_13_3462, i_13_3463, i_13_3464, i_13_3465, i_13_3466, i_13_3467, i_13_3468, i_13_3469, i_13_3470, i_13_3471, i_13_3472, i_13_3473, i_13_3474, i_13_3475, i_13_3476, i_13_3477, i_13_3478, i_13_3479, i_13_3480, i_13_3481, i_13_3482, i_13_3483, i_13_3484, i_13_3485, i_13_3486, i_13_3487, i_13_3488, i_13_3489, i_13_3490, i_13_3491, i_13_3492, i_13_3493, i_13_3494, i_13_3495, i_13_3496, i_13_3497, i_13_3498, i_13_3499, i_13_3500, i_13_3501, i_13_3502, i_13_3503, i_13_3504, i_13_3505, i_13_3506, i_13_3507, i_13_3508, i_13_3509, i_13_3510, i_13_3511, i_13_3512, i_13_3513, i_13_3514, i_13_3515, i_13_3516, i_13_3517, i_13_3518, i_13_3519, i_13_3520, i_13_3521, i_13_3522, i_13_3523, i_13_3524, i_13_3525, i_13_3526, i_13_3527, i_13_3528, i_13_3529, i_13_3530, i_13_3531, i_13_3532, i_13_3533, i_13_3534, i_13_3535, i_13_3536, i_13_3537, i_13_3538, i_13_3539, i_13_3540, i_13_3541, i_13_3542, i_13_3543, i_13_3544, i_13_3545, i_13_3546, i_13_3547, i_13_3548, i_13_3549, i_13_3550, i_13_3551, i_13_3552, i_13_3553, i_13_3554, i_13_3555, i_13_3556, i_13_3557, i_13_3558, i_13_3559, i_13_3560, i_13_3561, i_13_3562, i_13_3563, i_13_3564, i_13_3565, i_13_3566, i_13_3567, i_13_3568, i_13_3569, i_13_3570, i_13_3571, i_13_3572, i_13_3573, i_13_3574, i_13_3575, i_13_3576, i_13_3577, i_13_3578, i_13_3579, i_13_3580, i_13_3581, i_13_3582, i_13_3583, i_13_3584, i_13_3585, i_13_3586, i_13_3587, i_13_3588, i_13_3589, i_13_3590, i_13_3591, i_13_3592, i_13_3593, i_13_3594, i_13_3595, i_13_3596, i_13_3597, i_13_3598, i_13_3599, i_13_3600, i_13_3601, i_13_3602, i_13_3603, i_13_3604, i_13_3605, i_13_3606, i_13_3607, i_13_3608, i_13_3609, i_13_3610, i_13_3611, i_13_3612, i_13_3613, i_13_3614, i_13_3615, i_13_3616, i_13_3617, i_13_3618, i_13_3619, i_13_3620, i_13_3621, i_13_3622, i_13_3623, i_13_3624, i_13_3625, i_13_3626, i_13_3627, i_13_3628, i_13_3629, i_13_3630, i_13_3631, i_13_3632, i_13_3633, i_13_3634, i_13_3635, i_13_3636, i_13_3637, i_13_3638, i_13_3639, i_13_3640, i_13_3641, i_13_3642, i_13_3643, i_13_3644, i_13_3645, i_13_3646, i_13_3647, i_13_3648, i_13_3649, i_13_3650, i_13_3651, i_13_3652, i_13_3653, i_13_3654, i_13_3655, i_13_3656, i_13_3657, i_13_3658, i_13_3659, i_13_3660, i_13_3661, i_13_3662, i_13_3663, i_13_3664, i_13_3665, i_13_3666, i_13_3667, i_13_3668, i_13_3669, i_13_3670, i_13_3671, i_13_3672, i_13_3673, i_13_3674, i_13_3675, i_13_3676, i_13_3677, i_13_3678, i_13_3679, i_13_3680, i_13_3681, i_13_3682, i_13_3683, i_13_3684, i_13_3685, i_13_3686, i_13_3687, i_13_3688, i_13_3689, i_13_3690, i_13_3691, i_13_3692, i_13_3693, i_13_3694, i_13_3695, i_13_3696, i_13_3697, i_13_3698, i_13_3699, i_13_3700, i_13_3701, i_13_3702, i_13_3703, i_13_3704, i_13_3705, i_13_3706, i_13_3707, i_13_3708, i_13_3709, i_13_3710, i_13_3711, i_13_3712, i_13_3713, i_13_3714, i_13_3715, i_13_3716, i_13_3717, i_13_3718, i_13_3719, i_13_3720, i_13_3721, i_13_3722, i_13_3723, i_13_3724, i_13_3725, i_13_3726, i_13_3727, i_13_3728, i_13_3729, i_13_3730, i_13_3731, i_13_3732, i_13_3733, i_13_3734, i_13_3735, i_13_3736, i_13_3737, i_13_3738, i_13_3739, i_13_3740, i_13_3741, i_13_3742, i_13_3743, i_13_3744, i_13_3745, i_13_3746, i_13_3747, i_13_3748, i_13_3749, i_13_3750, i_13_3751, i_13_3752, i_13_3753, i_13_3754, i_13_3755, i_13_3756, i_13_3757, i_13_3758, i_13_3759, i_13_3760, i_13_3761, i_13_3762, i_13_3763, i_13_3764, i_13_3765, i_13_3766, i_13_3767, i_13_3768, i_13_3769, i_13_3770, i_13_3771, i_13_3772, i_13_3773, i_13_3774, i_13_3775, i_13_3776, i_13_3777, i_13_3778, i_13_3779, i_13_3780, i_13_3781, i_13_3782, i_13_3783, i_13_3784, i_13_3785, i_13_3786, i_13_3787, i_13_3788, i_13_3789, i_13_3790, i_13_3791, i_13_3792, i_13_3793, i_13_3794, i_13_3795, i_13_3796, i_13_3797, i_13_3798, i_13_3799, i_13_3800, i_13_3801, i_13_3802, i_13_3803, i_13_3804, i_13_3805, i_13_3806, i_13_3807, i_13_3808, i_13_3809, i_13_3810, i_13_3811, i_13_3812, i_13_3813, i_13_3814, i_13_3815, i_13_3816, i_13_3817, i_13_3818, i_13_3819, i_13_3820, i_13_3821, i_13_3822, i_13_3823, i_13_3824, i_13_3825, i_13_3826, i_13_3827, i_13_3828, i_13_3829, i_13_3830, i_13_3831, i_13_3832, i_13_3833, i_13_3834, i_13_3835, i_13_3836, i_13_3837, i_13_3838, i_13_3839, i_13_3840, i_13_3841, i_13_3842, i_13_3843, i_13_3844, i_13_3845, i_13_3846, i_13_3847, i_13_3848, i_13_3849, i_13_3850, i_13_3851, i_13_3852, i_13_3853, i_13_3854, i_13_3855, i_13_3856, i_13_3857, i_13_3858, i_13_3859, i_13_3860, i_13_3861, i_13_3862, i_13_3863, i_13_3864, i_13_3865, i_13_3866, i_13_3867, i_13_3868, i_13_3869, i_13_3870, i_13_3871, i_13_3872, i_13_3873, i_13_3874, i_13_3875, i_13_3876, i_13_3877, i_13_3878, i_13_3879, i_13_3880, i_13_3881, i_13_3882, i_13_3883, i_13_3884, i_13_3885, i_13_3886, i_13_3887, i_13_3888, i_13_3889, i_13_3890, i_13_3891, i_13_3892, i_13_3893, i_13_3894, i_13_3895, i_13_3896, i_13_3897, i_13_3898, i_13_3899, i_13_3900, i_13_3901, i_13_3902, i_13_3903, i_13_3904, i_13_3905, i_13_3906, i_13_3907, i_13_3908, i_13_3909, i_13_3910, i_13_3911, i_13_3912, i_13_3913, i_13_3914, i_13_3915, i_13_3916, i_13_3917, i_13_3918, i_13_3919, i_13_3920, i_13_3921, i_13_3922, i_13_3923, i_13_3924, i_13_3925, i_13_3926, i_13_3927, i_13_3928, i_13_3929, i_13_3930, i_13_3931, i_13_3932, i_13_3933, i_13_3934, i_13_3935, i_13_3936, i_13_3937, i_13_3938, i_13_3939, i_13_3940, i_13_3941, i_13_3942, i_13_3943, i_13_3944, i_13_3945, i_13_3946, i_13_3947, i_13_3948, i_13_3949, i_13_3950, i_13_3951, i_13_3952, i_13_3953, i_13_3954, i_13_3955, i_13_3956, i_13_3957, i_13_3958, i_13_3959, i_13_3960, i_13_3961, i_13_3962, i_13_3963, i_13_3964, i_13_3965, i_13_3966, i_13_3967, i_13_3968, i_13_3969, i_13_3970, i_13_3971, i_13_3972, i_13_3973, i_13_3974, i_13_3975, i_13_3976, i_13_3977, i_13_3978, i_13_3979, i_13_3980, i_13_3981, i_13_3982, i_13_3983, i_13_3984, i_13_3985, i_13_3986, i_13_3987, i_13_3988, i_13_3989, i_13_3990, i_13_3991, i_13_3992, i_13_3993, i_13_3994, i_13_3995, i_13_3996, i_13_3997, i_13_3998, i_13_3999, i_13_4000, i_13_4001, i_13_4002, i_13_4003, i_13_4004, i_13_4005, i_13_4006, i_13_4007, i_13_4008, i_13_4009, i_13_4010, i_13_4011, i_13_4012, i_13_4013, i_13_4014, i_13_4015, i_13_4016, i_13_4017, i_13_4018, i_13_4019, i_13_4020, i_13_4021, i_13_4022, i_13_4023, i_13_4024, i_13_4025, i_13_4026, i_13_4027, i_13_4028, i_13_4029, i_13_4030, i_13_4031, i_13_4032, i_13_4033, i_13_4034, i_13_4035, i_13_4036, i_13_4037, i_13_4038, i_13_4039, i_13_4040, i_13_4041, i_13_4042, i_13_4043, i_13_4044, i_13_4045, i_13_4046, i_13_4047, i_13_4048, i_13_4049, i_13_4050, i_13_4051, i_13_4052, i_13_4053, i_13_4054, i_13_4055, i_13_4056, i_13_4057, i_13_4058, i_13_4059, i_13_4060, i_13_4061, i_13_4062, i_13_4063, i_13_4064, i_13_4065, i_13_4066, i_13_4067, i_13_4068, i_13_4069, i_13_4070, i_13_4071, i_13_4072, i_13_4073, i_13_4074, i_13_4075, i_13_4076, i_13_4077, i_13_4078, i_13_4079, i_13_4080, i_13_4081, i_13_4082, i_13_4083, i_13_4084, i_13_4085, i_13_4086, i_13_4087, i_13_4088, i_13_4089, i_13_4090, i_13_4091, i_13_4092, i_13_4093, i_13_4094, i_13_4095, i_13_4096, i_13_4097, i_13_4098, i_13_4099, i_13_4100, i_13_4101, i_13_4102, i_13_4103, i_13_4104, i_13_4105, i_13_4106, i_13_4107, i_13_4108, i_13_4109, i_13_4110, i_13_4111, i_13_4112, i_13_4113, i_13_4114, i_13_4115, i_13_4116, i_13_4117, i_13_4118, i_13_4119, i_13_4120, i_13_4121, i_13_4122, i_13_4123, i_13_4124, i_13_4125, i_13_4126, i_13_4127, i_13_4128, i_13_4129, i_13_4130, i_13_4131, i_13_4132, i_13_4133, i_13_4134, i_13_4135, i_13_4136, i_13_4137, i_13_4138, i_13_4139, i_13_4140, i_13_4141, i_13_4142, i_13_4143, i_13_4144, i_13_4145, i_13_4146, i_13_4147, i_13_4148, i_13_4149, i_13_4150, i_13_4151, i_13_4152, i_13_4153, i_13_4154, i_13_4155, i_13_4156, i_13_4157, i_13_4158, i_13_4159, i_13_4160, i_13_4161, i_13_4162, i_13_4163, i_13_4164, i_13_4165, i_13_4166, i_13_4167, i_13_4168, i_13_4169, i_13_4170, i_13_4171, i_13_4172, i_13_4173, i_13_4174, i_13_4175, i_13_4176, i_13_4177, i_13_4178, i_13_4179, i_13_4180, i_13_4181, i_13_4182, i_13_4183, i_13_4184, i_13_4185, i_13_4186, i_13_4187, i_13_4188, i_13_4189, i_13_4190, i_13_4191, i_13_4192, i_13_4193, i_13_4194, i_13_4195, i_13_4196, i_13_4197, i_13_4198, i_13_4199, i_13_4200, i_13_4201, i_13_4202, i_13_4203, i_13_4204, i_13_4205, i_13_4206, i_13_4207, i_13_4208, i_13_4209, i_13_4210, i_13_4211, i_13_4212, i_13_4213, i_13_4214, i_13_4215, i_13_4216, i_13_4217, i_13_4218, i_13_4219, i_13_4220, i_13_4221, i_13_4222, i_13_4223, i_13_4224, i_13_4225, i_13_4226, i_13_4227, i_13_4228, i_13_4229, i_13_4230, i_13_4231, i_13_4232, i_13_4233, i_13_4234, i_13_4235, i_13_4236, i_13_4237, i_13_4238, i_13_4239, i_13_4240, i_13_4241, i_13_4242, i_13_4243, i_13_4244, i_13_4245, i_13_4246, i_13_4247, i_13_4248, i_13_4249, i_13_4250, i_13_4251, i_13_4252, i_13_4253, i_13_4254, i_13_4255, i_13_4256, i_13_4257, i_13_4258, i_13_4259, i_13_4260, i_13_4261, i_13_4262, i_13_4263, i_13_4264, i_13_4265, i_13_4266, i_13_4267, i_13_4268, i_13_4269, i_13_4270, i_13_4271, i_13_4272, i_13_4273, i_13_4274, i_13_4275, i_13_4276, i_13_4277, i_13_4278, i_13_4279, i_13_4280, i_13_4281, i_13_4282, i_13_4283, i_13_4284, i_13_4285, i_13_4286, i_13_4287, i_13_4288, i_13_4289, i_13_4290, i_13_4291, i_13_4292, i_13_4293, i_13_4294, i_13_4295, i_13_4296, i_13_4297, i_13_4298, i_13_4299, i_13_4300, i_13_4301, i_13_4302, i_13_4303, i_13_4304, i_13_4305, i_13_4306, i_13_4307, i_13_4308, i_13_4309, i_13_4310, i_13_4311, i_13_4312, i_13_4313, i_13_4314, i_13_4315, i_13_4316, i_13_4317, i_13_4318, i_13_4319, i_13_4320, i_13_4321, i_13_4322, i_13_4323, i_13_4324, i_13_4325, i_13_4326, i_13_4327, i_13_4328, i_13_4329, i_13_4330, i_13_4331, i_13_4332, i_13_4333, i_13_4334, i_13_4335, i_13_4336, i_13_4337, i_13_4338, i_13_4339, i_13_4340, i_13_4341, i_13_4342, i_13_4343, i_13_4344, i_13_4345, i_13_4346, i_13_4347, i_13_4348, i_13_4349, i_13_4350, i_13_4351, i_13_4352, i_13_4353, i_13_4354, i_13_4355, i_13_4356, i_13_4357, i_13_4358, i_13_4359, i_13_4360, i_13_4361, i_13_4362, i_13_4363, i_13_4364, i_13_4365, i_13_4366, i_13_4367, i_13_4368, i_13_4369, i_13_4370, i_13_4371, i_13_4372, i_13_4373, i_13_4374, i_13_4375, i_13_4376, i_13_4377, i_13_4378, i_13_4379, i_13_4380, i_13_4381, i_13_4382, i_13_4383, i_13_4384, i_13_4385, i_13_4386, i_13_4387, i_13_4388, i_13_4389, i_13_4390, i_13_4391, i_13_4392, i_13_4393, i_13_4394, i_13_4395, i_13_4396, i_13_4397, i_13_4398, i_13_4399, i_13_4400, i_13_4401, i_13_4402, i_13_4403, i_13_4404, i_13_4405, i_13_4406, i_13_4407, i_13_4408, i_13_4409, i_13_4410, i_13_4411, i_13_4412, i_13_4413, i_13_4414, i_13_4415, i_13_4416, i_13_4417, i_13_4418, i_13_4419, i_13_4420, i_13_4421, i_13_4422, i_13_4423, i_13_4424, i_13_4425, i_13_4426, i_13_4427, i_13_4428, i_13_4429, i_13_4430, i_13_4431, i_13_4432, i_13_4433, i_13_4434, i_13_4435, i_13_4436, i_13_4437, i_13_4438, i_13_4439, i_13_4440, i_13_4441, i_13_4442, i_13_4443, i_13_4444, i_13_4445, i_13_4446, i_13_4447, i_13_4448, i_13_4449, i_13_4450, i_13_4451, i_13_4452, i_13_4453, i_13_4454, i_13_4455, i_13_4456, i_13_4457, i_13_4458, i_13_4459, i_13_4460, i_13_4461, i_13_4462, i_13_4463, i_13_4464, i_13_4465, i_13_4466, i_13_4467, i_13_4468, i_13_4469, i_13_4470, i_13_4471, i_13_4472, i_13_4473, i_13_4474, i_13_4475, i_13_4476, i_13_4477, i_13_4478, i_13_4479, i_13_4480, i_13_4481, i_13_4482, i_13_4483, i_13_4484, i_13_4485, i_13_4486, i_13_4487, i_13_4488, i_13_4489, i_13_4490, i_13_4491, i_13_4492, i_13_4493, i_13_4494, i_13_4495, i_13_4496, i_13_4497, i_13_4498, i_13_4499, i_13_4500, i_13_4501, i_13_4502, i_13_4503, i_13_4504, i_13_4505, i_13_4506, i_13_4507, i_13_4508, i_13_4509, i_13_4510, i_13_4511, i_13_4512, i_13_4513, i_13_4514, i_13_4515, i_13_4516, i_13_4517, i_13_4518, i_13_4519, i_13_4520, i_13_4521, i_13_4522, i_13_4523, i_13_4524, i_13_4525, i_13_4526, i_13_4527, i_13_4528, i_13_4529, i_13_4530, i_13_4531, i_13_4532, i_13_4533, i_13_4534, i_13_4535, i_13_4536, i_13_4537, i_13_4538, i_13_4539, i_13_4540, i_13_4541, i_13_4542, i_13_4543, i_13_4544, i_13_4545, i_13_4546, i_13_4547, i_13_4548, i_13_4549, i_13_4550, i_13_4551, i_13_4552, i_13_4553, i_13_4554, i_13_4555, i_13_4556, i_13_4557, i_13_4558, i_13_4559, i_13_4560, i_13_4561, i_13_4562, i_13_4563, i_13_4564, i_13_4565, i_13_4566, i_13_4567, i_13_4568, i_13_4569, i_13_4570, i_13_4571, i_13_4572, i_13_4573, i_13_4574, i_13_4575, i_13_4576, i_13_4577, i_13_4578, i_13_4579, i_13_4580, i_13_4581, i_13_4582, i_13_4583, i_13_4584, i_13_4585, i_13_4586, i_13_4587, i_13_4588, i_13_4589, i_13_4590, i_13_4591, i_13_4592, i_13_4593, i_13_4594, i_13_4595, i_13_4596, i_13_4597, i_13_4598, i_13_4599, i_13_4600, i_13_4601, i_13_4602, i_13_4603, i_13_4604, i_13_4605, i_13_4606, i_13_4607;
output o_13_0, o_13_1, o_13_2, o_13_3, o_13_4, o_13_5, o_13_6, o_13_7, o_13_8, o_13_9, o_13_10, o_13_11, o_13_12, o_13_13, o_13_14, o_13_15, o_13_16, o_13_17, o_13_18, o_13_19, o_13_20, o_13_21, o_13_22, o_13_23, o_13_24, o_13_25, o_13_26, o_13_27, o_13_28, o_13_29, o_13_30, o_13_31, o_13_32, o_13_33, o_13_34, o_13_35, o_13_36, o_13_37, o_13_38, o_13_39, o_13_40, o_13_41, o_13_42, o_13_43, o_13_44, o_13_45, o_13_46, o_13_47, o_13_48, o_13_49, o_13_50, o_13_51, o_13_52, o_13_53, o_13_54, o_13_55, o_13_56, o_13_57, o_13_58, o_13_59, o_13_60, o_13_61, o_13_62, o_13_63, o_13_64, o_13_65, o_13_66, o_13_67, o_13_68, o_13_69, o_13_70, o_13_71, o_13_72, o_13_73, o_13_74, o_13_75, o_13_76, o_13_77, o_13_78, o_13_79, o_13_80, o_13_81, o_13_82, o_13_83, o_13_84, o_13_85, o_13_86, o_13_87, o_13_88, o_13_89, o_13_90, o_13_91, o_13_92, o_13_93, o_13_94, o_13_95, o_13_96, o_13_97, o_13_98, o_13_99, o_13_100, o_13_101, o_13_102, o_13_103, o_13_104, o_13_105, o_13_106, o_13_107, o_13_108, o_13_109, o_13_110, o_13_111, o_13_112, o_13_113, o_13_114, o_13_115, o_13_116, o_13_117, o_13_118, o_13_119, o_13_120, o_13_121, o_13_122, o_13_123, o_13_124, o_13_125, o_13_126, o_13_127, o_13_128, o_13_129, o_13_130, o_13_131, o_13_132, o_13_133, o_13_134, o_13_135, o_13_136, o_13_137, o_13_138, o_13_139, o_13_140, o_13_141, o_13_142, o_13_143, o_13_144, o_13_145, o_13_146, o_13_147, o_13_148, o_13_149, o_13_150, o_13_151, o_13_152, o_13_153, o_13_154, o_13_155, o_13_156, o_13_157, o_13_158, o_13_159, o_13_160, o_13_161, o_13_162, o_13_163, o_13_164, o_13_165, o_13_166, o_13_167, o_13_168, o_13_169, o_13_170, o_13_171, o_13_172, o_13_173, o_13_174, o_13_175, o_13_176, o_13_177, o_13_178, o_13_179, o_13_180, o_13_181, o_13_182, o_13_183, o_13_184, o_13_185, o_13_186, o_13_187, o_13_188, o_13_189, o_13_190, o_13_191, o_13_192, o_13_193, o_13_194, o_13_195, o_13_196, o_13_197, o_13_198, o_13_199, o_13_200, o_13_201, o_13_202, o_13_203, o_13_204, o_13_205, o_13_206, o_13_207, o_13_208, o_13_209, o_13_210, o_13_211, o_13_212, o_13_213, o_13_214, o_13_215, o_13_216, o_13_217, o_13_218, o_13_219, o_13_220, o_13_221, o_13_222, o_13_223, o_13_224, o_13_225, o_13_226, o_13_227, o_13_228, o_13_229, o_13_230, o_13_231, o_13_232, o_13_233, o_13_234, o_13_235, o_13_236, o_13_237, o_13_238, o_13_239, o_13_240, o_13_241, o_13_242, o_13_243, o_13_244, o_13_245, o_13_246, o_13_247, o_13_248, o_13_249, o_13_250, o_13_251, o_13_252, o_13_253, o_13_254, o_13_255, o_13_256, o_13_257, o_13_258, o_13_259, o_13_260, o_13_261, o_13_262, o_13_263, o_13_264, o_13_265, o_13_266, o_13_267, o_13_268, o_13_269, o_13_270, o_13_271, o_13_272, o_13_273, o_13_274, o_13_275, o_13_276, o_13_277, o_13_278, o_13_279, o_13_280, o_13_281, o_13_282, o_13_283, o_13_284, o_13_285, o_13_286, o_13_287, o_13_288, o_13_289, o_13_290, o_13_291, o_13_292, o_13_293, o_13_294, o_13_295, o_13_296, o_13_297, o_13_298, o_13_299, o_13_300, o_13_301, o_13_302, o_13_303, o_13_304, o_13_305, o_13_306, o_13_307, o_13_308, o_13_309, o_13_310, o_13_311, o_13_312, o_13_313, o_13_314, o_13_315, o_13_316, o_13_317, o_13_318, o_13_319, o_13_320, o_13_321, o_13_322, o_13_323, o_13_324, o_13_325, o_13_326, o_13_327, o_13_328, o_13_329, o_13_330, o_13_331, o_13_332, o_13_333, o_13_334, o_13_335, o_13_336, o_13_337, o_13_338, o_13_339, o_13_340, o_13_341, o_13_342, o_13_343, o_13_344, o_13_345, o_13_346, o_13_347, o_13_348, o_13_349, o_13_350, o_13_351, o_13_352, o_13_353, o_13_354, o_13_355, o_13_356, o_13_357, o_13_358, o_13_359, o_13_360, o_13_361, o_13_362, o_13_363, o_13_364, o_13_365, o_13_366, o_13_367, o_13_368, o_13_369, o_13_370, o_13_371, o_13_372, o_13_373, o_13_374, o_13_375, o_13_376, o_13_377, o_13_378, o_13_379, o_13_380, o_13_381, o_13_382, o_13_383, o_13_384, o_13_385, o_13_386, o_13_387, o_13_388, o_13_389, o_13_390, o_13_391, o_13_392, o_13_393, o_13_394, o_13_395, o_13_396, o_13_397, o_13_398, o_13_399, o_13_400, o_13_401, o_13_402, o_13_403, o_13_404, o_13_405, o_13_406, o_13_407, o_13_408, o_13_409, o_13_410, o_13_411, o_13_412, o_13_413, o_13_414, o_13_415, o_13_416, o_13_417, o_13_418, o_13_419, o_13_420, o_13_421, o_13_422, o_13_423, o_13_424, o_13_425, o_13_426, o_13_427, o_13_428, o_13_429, o_13_430, o_13_431, o_13_432, o_13_433, o_13_434, o_13_435, o_13_436, o_13_437, o_13_438, o_13_439, o_13_440, o_13_441, o_13_442, o_13_443, o_13_444, o_13_445, o_13_446, o_13_447, o_13_448, o_13_449, o_13_450, o_13_451, o_13_452, o_13_453, o_13_454, o_13_455, o_13_456, o_13_457, o_13_458, o_13_459, o_13_460, o_13_461, o_13_462, o_13_463, o_13_464, o_13_465, o_13_466, o_13_467, o_13_468, o_13_469, o_13_470, o_13_471, o_13_472, o_13_473, o_13_474, o_13_475, o_13_476, o_13_477, o_13_478, o_13_479, o_13_480, o_13_481, o_13_482, o_13_483, o_13_484, o_13_485, o_13_486, o_13_487, o_13_488, o_13_489, o_13_490, o_13_491, o_13_492, o_13_493, o_13_494, o_13_495, o_13_496, o_13_497, o_13_498, o_13_499, o_13_500, o_13_501, o_13_502, o_13_503, o_13_504, o_13_505, o_13_506, o_13_507, o_13_508, o_13_509, o_13_510, o_13_511;
	kernel_13_0 k_13_0(i_13_20, i_13_59, i_13_74, i_13_76, i_13_182, i_13_187, i_13_232, i_13_283, i_13_286, i_13_338, i_13_445, i_13_448, i_13_535, i_13_548, i_13_574, i_13_617, i_13_629, i_13_643, i_13_644, i_13_646, i_13_647, i_13_652, i_13_689, i_13_718, i_13_781, i_13_782, i_13_827, i_13_835, i_13_895, i_13_977, i_13_980, i_13_1120, i_13_1124, i_13_1132, i_13_1142, i_13_1151, i_13_1231, i_13_1258, i_13_1277, i_13_1286, i_13_1394, i_13_1411, i_13_1435, i_13_1465, i_13_1483, i_13_1484, i_13_1627, i_13_1642, i_13_1646, i_13_1673, i_13_1753, i_13_1790, i_13_1796, i_13_1799, i_13_1802, i_13_1804, i_13_1840, i_13_1862, i_13_2000, i_13_2150, i_13_2168, i_13_2201, i_13_2239, i_13_2276, i_13_2311, i_13_2383, i_13_2545, i_13_2570, i_13_2848, i_13_2851, i_13_2852, i_13_2878, i_13_2879, i_13_2885, i_13_3028, i_13_3047, i_13_3095, i_13_3122, i_13_3293, i_13_3356, i_13_3389, i_13_3406, i_13_3433, i_13_3446, i_13_3482, i_13_3722, i_13_3734, i_13_3794, i_13_3839, i_13_3887, i_13_3985, i_13_4012, i_13_4013, i_13_4046, i_13_4189, i_13_4301, i_13_4315, i_13_4435, i_13_4481, i_13_4541, o_13_0);
	kernel_13_1 k_13_1(i_13_40, i_13_73, i_13_90, i_13_91, i_13_93, i_13_94, i_13_97, i_13_111, i_13_118, i_13_160, i_13_177, i_13_273, i_13_306, i_13_310, i_13_364, i_13_411, i_13_561, i_13_567, i_13_568, i_13_571, i_13_604, i_13_694, i_13_697, i_13_729, i_13_730, i_13_733, i_13_793, i_13_855, i_13_861, i_13_863, i_13_942, i_13_1058, i_13_1210, i_13_1405, i_13_1440, i_13_1486, i_13_1491, i_13_1681, i_13_1781, i_13_1828, i_13_1836, i_13_1837, i_13_1862, i_13_1918, i_13_2172, i_13_2173, i_13_2205, i_13_2206, i_13_2316, i_13_2365, i_13_2421, i_13_2422, i_13_2433, i_13_2434, i_13_2437, i_13_2452, i_13_2464, i_13_2551, i_13_2677, i_13_2888, i_13_2985, i_13_3023, i_13_3064, i_13_3102, i_13_3149, i_13_3164, i_13_3166, i_13_3208, i_13_3423, i_13_3424, i_13_3489, i_13_3490, i_13_3535, i_13_3541, i_13_3568, i_13_3577, i_13_3682, i_13_3699, i_13_3762, i_13_3856, i_13_3870, i_13_3871, i_13_3872, i_13_3877, i_13_3972, i_13_3982, i_13_4118, i_13_4155, i_13_4278, i_13_4335, i_13_4350, i_13_4351, i_13_4354, i_13_4378, i_13_4390, i_13_4425, i_13_4536, i_13_4540, i_13_4567, i_13_4591, o_13_1);
	kernel_13_2 k_13_2(i_13_94, i_13_103, i_13_104, i_13_143, i_13_157, i_13_280, i_13_316, i_13_379, i_13_523, i_13_586, i_13_604, i_13_666, i_13_671, i_13_696, i_13_768, i_13_802, i_13_850, i_13_959, i_13_1081, i_13_1142, i_13_1206, i_13_1207, i_13_1274, i_13_1277, i_13_1300, i_13_1341, i_13_1342, i_13_1343, i_13_1363, i_13_1403, i_13_1435, i_13_1440, i_13_1467, i_13_1515, i_13_1594, i_13_1692, i_13_1714, i_13_1750, i_13_1781, i_13_1802, i_13_1810, i_13_1840, i_13_1882, i_13_1900, i_13_1926, i_13_1927, i_13_1939, i_13_2002, i_13_2011, i_13_2052, i_13_2053, i_13_2054, i_13_2173, i_13_2189, i_13_2197, i_13_2236, i_13_2278, i_13_2396, i_13_2423, i_13_2450, i_13_2548, i_13_2592, i_13_2614, i_13_2615, i_13_2695, i_13_2710, i_13_2853, i_13_2854, i_13_3019, i_13_3109, i_13_3329, i_13_3343, i_13_3366, i_13_3367, i_13_3386, i_13_3398, i_13_3404, i_13_3439, i_13_3487, i_13_3502, i_13_3611, i_13_3619, i_13_3650, i_13_3736, i_13_3910, i_13_3931, i_13_3994, i_13_3995, i_13_4015, i_13_4087, i_13_4104, i_13_4230, i_13_4231, i_13_4232, i_13_4267, i_13_4392, i_13_4393, i_13_4394, i_13_4554, i_13_4559, o_13_2);
	kernel_13_3 k_13_3(i_13_46, i_13_74, i_13_100, i_13_108, i_13_110, i_13_127, i_13_166, i_13_280, i_13_281, i_13_284, i_13_486, i_13_677, i_13_723, i_13_758, i_13_760, i_13_794, i_13_820, i_13_821, i_13_856, i_13_946, i_13_1215, i_13_1216, i_13_1217, i_13_1219, i_13_1317, i_13_1341, i_13_1388, i_13_1422, i_13_1424, i_13_1486, i_13_1487, i_13_1494, i_13_1566, i_13_1605, i_13_1630, i_13_1732, i_13_1774, i_13_1804, i_13_1837, i_13_1838, i_13_1841, i_13_1883, i_13_1911, i_13_1940, i_13_1945, i_13_1999, i_13_2000, i_13_2055, i_13_2146, i_13_2170, i_13_2236, i_13_2263, i_13_2335, i_13_2422, i_13_2435, i_13_2448, i_13_2532, i_13_2611, i_13_2612, i_13_2614, i_13_2709, i_13_2716, i_13_2746, i_13_2767, i_13_2782, i_13_2882, i_13_2955, i_13_2961, i_13_3034, i_13_3051, i_13_3145, i_13_3146, i_13_3379, i_13_3422, i_13_3438, i_13_3452, i_13_3502, i_13_3503, i_13_3529, i_13_3530, i_13_3610, i_13_3726, i_13_3729, i_13_3735, i_13_3736, i_13_3739, i_13_3872, i_13_3889, i_13_3890, i_13_3980, i_13_4053, i_13_4121, i_13_4158, i_13_4248, i_13_4252, i_13_4262, i_13_4322, i_13_4340, i_13_4415, i_13_4557, o_13_3);
	kernel_13_4 k_13_4(i_13_192, i_13_199, i_13_225, i_13_324, i_13_378, i_13_531, i_13_532, i_13_573, i_13_577, i_13_639, i_13_640, i_13_658, i_13_660, i_13_661, i_13_714, i_13_768, i_13_849, i_13_927, i_13_945, i_13_1062, i_13_1080, i_13_1084, i_13_1116, i_13_1188, i_13_1206, i_13_1254, i_13_1407, i_13_1423, i_13_1506, i_13_1513, i_13_1539, i_13_1593, i_13_1594, i_13_1638, i_13_1639, i_13_1710, i_13_1719, i_13_1782, i_13_1783, i_13_1792, i_13_1800, i_13_1801, i_13_1881, i_13_1882, i_13_1929, i_13_1989, i_13_1990, i_13_2055, i_13_2092, i_13_2100, i_13_2116, i_13_2341, i_13_2358, i_13_2376, i_13_2424, i_13_2460, i_13_2524, i_13_2532, i_13_2569, i_13_2673, i_13_2817, i_13_2844, i_13_2845, i_13_2934, i_13_2935, i_13_3024, i_13_3114, i_13_3141, i_13_3258, i_13_3259, i_13_3267, i_13_3285, i_13_3286, i_13_3381, i_13_3384, i_13_3394, i_13_3415, i_13_3420, i_13_3421, i_13_3423, i_13_3424, i_13_3447, i_13_3451, i_13_3472, i_13_3753, i_13_3790, i_13_3873, i_13_3919, i_13_3924, i_13_3982, i_13_4008, i_13_4009, i_13_4018, i_13_4050, i_13_4077, i_13_4078, i_13_4207, i_13_4249, i_13_4420, i_13_4521, o_13_4);
	kernel_13_5 k_13_5(i_13_71, i_13_76, i_13_175, i_13_178, i_13_209, i_13_245, i_13_283, i_13_284, i_13_286, i_13_287, i_13_374, i_13_410, i_13_517, i_13_526, i_13_527, i_13_625, i_13_689, i_13_691, i_13_800, i_13_814, i_13_818, i_13_826, i_13_851, i_13_923, i_13_1073, i_13_1097, i_13_1147, i_13_1312, i_13_1313, i_13_1499, i_13_1502, i_13_1543, i_13_1633, i_13_1634, i_13_1636, i_13_1637, i_13_1678, i_13_1681, i_13_1696, i_13_2005, i_13_2146, i_13_2194, i_13_2195, i_13_2291, i_13_2426, i_13_2438, i_13_2453, i_13_2462, i_13_2465, i_13_2527, i_13_2543, i_13_2677, i_13_2906, i_13_3025, i_13_3029, i_13_3050, i_13_3145, i_13_3146, i_13_3148, i_13_3172, i_13_3175, i_13_3272, i_13_3274, i_13_3275, i_13_3418, i_13_3425, i_13_3427, i_13_3428, i_13_3485, i_13_3490, i_13_3548, i_13_3616, i_13_3730, i_13_3731, i_13_3733, i_13_3734, i_13_3866, i_13_3892, i_13_3911, i_13_3913, i_13_3937, i_13_3995, i_13_4018, i_13_4019, i_13_4021, i_13_4022, i_13_4252, i_13_4253, i_13_4255, i_13_4256, i_13_4262, i_13_4264, i_13_4265, i_13_4342, i_13_4511, i_13_4559, i_13_4561, i_13_4562, i_13_4565, i_13_4586, o_13_5);
	kernel_13_6 k_13_6(i_13_139, i_13_229, i_13_280, i_13_282, i_13_285, i_13_410, i_13_418, i_13_475, i_13_561, i_13_562, i_13_574, i_13_849, i_13_850, i_13_853, i_13_924, i_13_981, i_13_988, i_13_1018, i_13_1021, i_13_1075, i_13_1219, i_13_1262, i_13_1308, i_13_1342, i_13_1345, i_13_1488, i_13_1496, i_13_1498, i_13_1515, i_13_1520, i_13_1630, i_13_1669, i_13_1678, i_13_1730, i_13_1753, i_13_1773, i_13_1809, i_13_1829, i_13_1854, i_13_1857, i_13_1858, i_13_1861, i_13_2002, i_13_2008, i_13_2028, i_13_2191, i_13_2226, i_13_2452, i_13_2455, i_13_2461, i_13_2539, i_13_2542, i_13_2544, i_13_2590, i_13_2722, i_13_2767, i_13_2857, i_13_3007, i_13_3010, i_13_3012, i_13_3037, i_13_3061, i_13_3064, i_13_3111, i_13_3127, i_13_3211, i_13_3235, i_13_3271, i_13_3442, i_13_3487, i_13_3490, i_13_3508, i_13_3541, i_13_3577, i_13_3640, i_13_3645, i_13_3729, i_13_3787, i_13_3817, i_13_3820, i_13_3838, i_13_3856, i_13_3888, i_13_3889, i_13_3907, i_13_3909, i_13_3910, i_13_3912, i_13_4078, i_13_4086, i_13_4250, i_13_4252, i_13_4254, i_13_4255, i_13_4375, i_13_4378, i_13_4380, i_13_4420, i_13_4426, i_13_4531, o_13_6);
	kernel_13_7 k_13_7(i_13_20, i_13_38, i_13_76, i_13_77, i_13_158, i_13_166, i_13_185, i_13_334, i_13_337, i_13_338, i_13_354, i_13_379, i_13_407, i_13_418, i_13_516, i_13_532, i_13_545, i_13_571, i_13_596, i_13_597, i_13_641, i_13_697, i_13_698, i_13_699, i_13_715, i_13_757, i_13_778, i_13_834, i_13_892, i_13_911, i_13_1067, i_13_1120, i_13_1219, i_13_1224, i_13_1297, i_13_1298, i_13_1301, i_13_1426, i_13_1499, i_13_1504, i_13_1523, i_13_1550, i_13_1558, i_13_1623, i_13_1747, i_13_1757, i_13_1783, i_13_1814, i_13_1840, i_13_1856, i_13_1904, i_13_1940, i_13_2116, i_13_2165, i_13_2169, i_13_2207, i_13_2209, i_13_2210, i_13_2225, i_13_2236, i_13_2261, i_13_2452, i_13_2458, i_13_2459, i_13_2549, i_13_2585, i_13_2639, i_13_2884, i_13_2935, i_13_2939, i_13_2980, i_13_2981, i_13_2985, i_13_3037, i_13_3170, i_13_3206, i_13_3217, i_13_3241, i_13_3290, i_13_3308, i_13_3415, i_13_3424, i_13_3568, i_13_3640, i_13_3700, i_13_3718, i_13_3755, i_13_3874, i_13_3908, i_13_3925, i_13_3987, i_13_4009, i_13_4010, i_13_4052, i_13_4054, i_13_4060, i_13_4261, i_13_4313, i_13_4333, i_13_4335, o_13_7);
	kernel_13_8 k_13_8(i_13_65, i_13_101, i_13_207, i_13_208, i_13_209, i_13_266, i_13_273, i_13_355, i_13_371, i_13_415, i_13_416, i_13_463, i_13_464, i_13_567, i_13_614, i_13_671, i_13_761, i_13_948, i_13_950, i_13_956, i_13_1081, i_13_1129, i_13_1319, i_13_1372, i_13_1504, i_13_1522, i_13_1523, i_13_1553, i_13_1604, i_13_1640, i_13_1687, i_13_1697, i_13_1786, i_13_1827, i_13_1830, i_13_1840, i_13_1841, i_13_1846, i_13_1847, i_13_1930, i_13_1931, i_13_1958, i_13_2056, i_13_2143, i_13_2200, i_13_2201, i_13_2237, i_13_2297, i_13_2399, i_13_2403, i_13_2444, i_13_2563, i_13_2692, i_13_2821, i_13_2822, i_13_3001, i_13_3045, i_13_3062, i_13_3164, i_13_3234, i_13_3240, i_13_3241, i_13_3242, i_13_3259, i_13_3261, i_13_3308, i_13_3343, i_13_3344, i_13_3388, i_13_3519, i_13_3538, i_13_3618, i_13_3619, i_13_3620, i_13_3631, i_13_3632, i_13_3637, i_13_3638, i_13_3857, i_13_3873, i_13_3904, i_13_3916, i_13_3928, i_13_3935, i_13_3988, i_13_3989, i_13_3992, i_13_4008, i_13_4061, i_13_4118, i_13_4205, i_13_4270, i_13_4271, i_13_4302, i_13_4312, i_13_4313, i_13_4339, i_13_4378, i_13_4477, i_13_4536, o_13_8);
	kernel_13_9 k_13_9(i_13_48, i_13_73, i_13_94, i_13_173, i_13_193, i_13_225, i_13_280, i_13_391, i_13_443, i_13_451, i_13_515, i_13_533, i_13_550, i_13_551, i_13_553, i_13_645, i_13_651, i_13_652, i_13_655, i_13_656, i_13_658, i_13_668, i_13_675, i_13_676, i_13_685, i_13_688, i_13_691, i_13_830, i_13_841, i_13_949, i_13_1098, i_13_1117, i_13_1144, i_13_1191, i_13_1267, i_13_1270, i_13_1305, i_13_1347, i_13_1383, i_13_1384, i_13_1404, i_13_1465, i_13_1515, i_13_1518, i_13_1773, i_13_1774, i_13_1777, i_13_1836, i_13_1858, i_13_1909, i_13_2046, i_13_2049, i_13_2058, i_13_2191, i_13_2351, i_13_2503, i_13_2511, i_13_2581, i_13_2627, i_13_2650, i_13_2749, i_13_2857, i_13_2999, i_13_3000, i_13_3037, i_13_3062, i_13_3087, i_13_3101, i_13_3214, i_13_3216, i_13_3235, i_13_3367, i_13_3371, i_13_3418, i_13_3532, i_13_3646, i_13_3863, i_13_3865, i_13_3888, i_13_3889, i_13_3890, i_13_3987, i_13_3988, i_13_3989, i_13_4018, i_13_4051, i_13_4054, i_13_4117, i_13_4122, i_13_4189, i_13_4233, i_13_4263, i_13_4305, i_13_4330, i_13_4366, i_13_4539, i_13_4594, i_13_4600, i_13_4601, i_13_4603, o_13_9);
	kernel_13_10 k_13_10(i_13_34, i_13_43, i_13_69, i_13_70, i_13_322, i_13_384, i_13_411, i_13_421, i_13_426, i_13_448, i_13_463, i_13_467, i_13_493, i_13_525, i_13_538, i_13_591, i_13_619, i_13_628, i_13_646, i_13_679, i_13_762, i_13_763, i_13_931, i_13_934, i_13_943, i_13_1021, i_13_1083, i_13_1096, i_13_1104, i_13_1105, i_13_1123, i_13_1131, i_13_1132, i_13_1347, i_13_1473, i_13_1510, i_13_1536, i_13_1537, i_13_1795, i_13_1797, i_13_1798, i_13_1803, i_13_1912, i_13_2001, i_13_2002, i_13_2023, i_13_2044, i_13_2048, i_13_2055, i_13_2231, i_13_2472, i_13_2508, i_13_2551, i_13_2599, i_13_2680, i_13_2724, i_13_2850, i_13_2859, i_13_2860, i_13_2904, i_13_2998, i_13_3030, i_13_3094, i_13_3127, i_13_3131, i_13_3155, i_13_3262, i_13_3264, i_13_3370, i_13_3390, i_13_3391, i_13_3417, i_13_3445, i_13_3558, i_13_3639, i_13_3640, i_13_3643, i_13_3649, i_13_3652, i_13_3680, i_13_3730, i_13_3769, i_13_3799, i_13_3847, i_13_3892, i_13_4021, i_13_4038, i_13_4039, i_13_4057, i_13_4084, i_13_4117, i_13_4166, i_13_4398, i_13_4408, i_13_4435, i_13_4541, i_13_4586, i_13_4596, i_13_4597, i_13_4606, o_13_10);
	kernel_13_11 k_13_11(i_13_45, i_13_69, i_13_76, i_13_93, i_13_127, i_13_384, i_13_385, i_13_411, i_13_462, i_13_537, i_13_564, i_13_603, i_13_645, i_13_682, i_13_825, i_13_882, i_13_933, i_13_1080, i_13_1086, i_13_1104, i_13_1341, i_13_1342, i_13_1401, i_13_1402, i_13_1468, i_13_1473, i_13_1479, i_13_1509, i_13_1510, i_13_1599, i_13_1600, i_13_1644, i_13_1657, i_13_1716, i_13_1717, i_13_1725, i_13_1728, i_13_1780, i_13_1797, i_13_1941, i_13_1995, i_13_1996, i_13_2053, i_13_2058, i_13_2176, i_13_2187, i_13_2188, i_13_2193, i_13_2265, i_13_2275, i_13_2277, i_13_2278, i_13_2304, i_13_2305, i_13_2340, i_13_2341, i_13_2424, i_13_2679, i_13_2725, i_13_2919, i_13_3066, i_13_3067, i_13_3102, i_13_3103, i_13_3147, i_13_3234, i_13_3289, i_13_3366, i_13_3394, i_13_3410, i_13_3441, i_13_3525, i_13_3555, i_13_3556, i_13_3580, i_13_3687, i_13_3688, i_13_3729, i_13_3730, i_13_3742, i_13_3786, i_13_3787, i_13_3796, i_13_3805, i_13_3816, i_13_3817, i_13_3894, i_13_3930, i_13_3991, i_13_3993, i_13_3994, i_13_4056, i_13_4057, i_13_4065, i_13_4093, i_13_4119, i_13_4166, i_13_4257, i_13_4393, i_13_4399, o_13_11);
	kernel_13_12 k_13_12(i_13_60, i_13_90, i_13_91, i_13_93, i_13_94, i_13_97, i_13_126, i_13_174, i_13_175, i_13_184, i_13_280, i_13_282, i_13_307, i_13_310, i_13_315, i_13_316, i_13_328, i_13_516, i_13_570, i_13_571, i_13_599, i_13_616, i_13_661, i_13_667, i_13_697, i_13_759, i_13_981, i_13_982, i_13_1020, i_13_1226, i_13_1256, i_13_1305, i_13_1323, i_13_1404, i_13_1426, i_13_1440, i_13_1441, i_13_1446, i_13_1494, i_13_1515, i_13_1629, i_13_1669, i_13_1769, i_13_1777, i_13_1828, i_13_1848, i_13_1849, i_13_1859, i_13_1885, i_13_1908, i_13_1921, i_13_1998, i_13_2003, i_13_2116, i_13_2172, i_13_2173, i_13_2407, i_13_2421, i_13_2676, i_13_2692, i_13_2875, i_13_2983, i_13_3026, i_13_3109, i_13_3163, i_13_3207, i_13_3241, i_13_3263, i_13_3327, i_13_3420, i_13_3421, i_13_3471, i_13_3478, i_13_3529, i_13_3556, i_13_3568, i_13_3575, i_13_3756, i_13_3765, i_13_3766, i_13_3782, i_13_3817, i_13_3844, i_13_3864, i_13_3871, i_13_3888, i_13_4037, i_13_4060, i_13_4066, i_13_4080, i_13_4163, i_13_4252, i_13_4316, i_13_4350, i_13_4351, i_13_4452, i_13_4469, i_13_4566, i_13_4567, i_13_4601, o_13_12);
	kernel_13_13 k_13_13(i_13_48, i_13_49, i_13_70, i_13_76, i_13_106, i_13_127, i_13_229, i_13_270, i_13_271, i_13_313, i_13_369, i_13_411, i_13_447, i_13_475, i_13_561, i_13_564, i_13_565, i_13_620, i_13_663, i_13_673, i_13_732, i_13_736, i_13_745, i_13_834, i_13_835, i_13_934, i_13_946, i_13_952, i_13_1043, i_13_1087, i_13_1104, i_13_1131, i_13_1150, i_13_1231, i_13_1232, i_13_1246, i_13_1402, i_13_1431, i_13_1465, i_13_1468, i_13_1497, i_13_1537, i_13_1566, i_13_1626, i_13_1657, i_13_1663, i_13_1729, i_13_1732, i_13_1735, i_13_1764, i_13_1765, i_13_1767, i_13_1797, i_13_1798, i_13_1805, i_13_1894, i_13_1947, i_13_2022, i_13_2029, i_13_2107, i_13_2175, i_13_2208, i_13_2223, i_13_2224, i_13_2436, i_13_2564, i_13_2709, i_13_2724, i_13_2754, i_13_2955, i_13_2968, i_13_3217, i_13_3258, i_13_3259, i_13_3264, i_13_3283, i_13_3354, i_13_3370, i_13_3478, i_13_3520, i_13_3536, i_13_3551, i_13_3757, i_13_3783, i_13_3900, i_13_3918, i_13_3930, i_13_4038, i_13_4045, i_13_4083, i_13_4164, i_13_4165, i_13_4189, i_13_4233, i_13_4269, i_13_4296, i_13_4324, i_13_4372, i_13_4513, i_13_4606, o_13_13);
	kernel_13_14 k_13_14(i_13_51, i_13_76, i_13_112, i_13_123, i_13_124, i_13_169, i_13_178, i_13_186, i_13_187, i_13_195, i_13_283, i_13_339, i_13_520, i_13_535, i_13_573, i_13_574, i_13_618, i_13_642, i_13_643, i_13_644, i_13_646, i_13_690, i_13_691, i_13_697, i_13_717, i_13_756, i_13_816, i_13_859, i_13_932, i_13_1068, i_13_1069, i_13_1123, i_13_1138, i_13_1258, i_13_1273, i_13_1282, i_13_1297, i_13_1384, i_13_1407, i_13_1426, i_13_1461, i_13_1552, i_13_1610, i_13_1642, i_13_1804, i_13_1839, i_13_1851, i_13_1852, i_13_1861, i_13_1990, i_13_1993, i_13_2118, i_13_2128, i_13_2133, i_13_2136, i_13_2149, i_13_2212, i_13_2227, i_13_2262, i_13_2263, i_13_2275, i_13_2379, i_13_2410, i_13_2451, i_13_2536, i_13_2636, i_13_2709, i_13_2847, i_13_2920, i_13_2986, i_13_3030, i_13_3112, i_13_3166, i_13_3174, i_13_3211, i_13_3220, i_13_3303, i_13_3339, i_13_3424, i_13_3426, i_13_3427, i_13_3541, i_13_3706, i_13_3768, i_13_3769, i_13_3823, i_13_3918, i_13_3995, i_13_4011, i_13_4012, i_13_4066, i_13_4081, i_13_4189, i_13_4282, i_13_4314, i_13_4317, i_13_4318, i_13_4566, i_13_4569, i_13_4594, o_13_14);
	kernel_13_15 k_13_15(i_13_235, i_13_328, i_13_329, i_13_527, i_13_530, i_13_599, i_13_611, i_13_646, i_13_671, i_13_676, i_13_700, i_13_718, i_13_777, i_13_799, i_13_826, i_13_827, i_13_862, i_13_863, i_13_895, i_13_941, i_13_1024, i_13_1025, i_13_1078, i_13_1079, i_13_1231, i_13_1258, i_13_1259, i_13_1318, i_13_1411, i_13_1430, i_13_1486, i_13_1492, i_13_1493, i_13_1609, i_13_1636, i_13_1651, i_13_1691, i_13_1736, i_13_1780, i_13_1781, i_13_1858, i_13_1861, i_13_1862, i_13_1921, i_13_2021, i_13_2023, i_13_2059, i_13_2194, i_13_2201, i_13_2239, i_13_2266, i_13_2294, i_13_2404, i_13_2405, i_13_2455, i_13_2464, i_13_2465, i_13_2545, i_13_2546, i_13_2617, i_13_2618, i_13_2633, i_13_2654, i_13_2708, i_13_2876, i_13_3017, i_13_3172, i_13_3173, i_13_3175, i_13_3176, i_13_3233, i_13_3367, i_13_3373, i_13_3464, i_13_3482, i_13_3536, i_13_3542, i_13_3544, i_13_3563, i_13_3622, i_13_3788, i_13_3806, i_13_3847, i_13_3859, i_13_3877, i_13_3890, i_13_3896, i_13_3914, i_13_4013, i_13_4019, i_13_4100, i_13_4118, i_13_4126, i_13_4162, i_13_4192, i_13_4262, i_13_4280, i_13_4373, i_13_4396, i_13_4444, o_13_15);
	kernel_13_16 k_13_16(i_13_35, i_13_106, i_13_178, i_13_187, i_13_284, i_13_322, i_13_325, i_13_326, i_13_355, i_13_454, i_13_480, i_13_496, i_13_521, i_13_562, i_13_574, i_13_575, i_13_599, i_13_644, i_13_646, i_13_647, i_13_685, i_13_718, i_13_849, i_13_850, i_13_851, i_13_914, i_13_1210, i_13_1229, i_13_1255, i_13_1282, i_13_1345, i_13_1410, i_13_1444, i_13_1471, i_13_1552, i_13_1646, i_13_1678, i_13_1683, i_13_1691, i_13_1740, i_13_1750, i_13_1753, i_13_1788, i_13_1807, i_13_1857, i_13_1858, i_13_1859, i_13_1861, i_13_1862, i_13_1958, i_13_1993, i_13_2050, i_13_2103, i_13_2141, i_13_2159, i_13_2182, i_13_2281, i_13_2302, i_13_2311, i_13_2459, i_13_2463, i_13_2551, i_13_2588, i_13_2653, i_13_2654, i_13_2722, i_13_2752, i_13_2790, i_13_3064, i_13_3170, i_13_3172, i_13_3175, i_13_3209, i_13_3235, i_13_3271, i_13_3272, i_13_3274, i_13_3275, i_13_3309, i_13_3401, i_13_3426, i_13_3433, i_13_3562, i_13_3563, i_13_3847, i_13_3856, i_13_3892, i_13_3911, i_13_3912, i_13_3913, i_13_3914, i_13_4016, i_13_4047, i_13_4098, i_13_4149, i_13_4262, i_13_4378, i_13_4379, i_13_4382, i_13_4581, o_13_16);
	kernel_13_17 k_13_17(i_13_27, i_13_28, i_13_31, i_13_63, i_13_67, i_13_90, i_13_100, i_13_111, i_13_130, i_13_174, i_13_196, i_13_225, i_13_226, i_13_255, i_13_306, i_13_307, i_13_372, i_13_462, i_13_612, i_13_616, i_13_666, i_13_667, i_13_670, i_13_729, i_13_796, i_13_828, i_13_853, i_13_855, i_13_858, i_13_1075, i_13_1120, i_13_1128, i_13_1200, i_13_1215, i_13_1225, i_13_1231, i_13_1306, i_13_1321, i_13_1344, i_13_1398, i_13_1440, i_13_1480, i_13_1620, i_13_1689, i_13_1696, i_13_1846, i_13_1927, i_13_1998, i_13_1999, i_13_2100, i_13_2200, i_13_2205, i_13_2206, i_13_2422, i_13_2430, i_13_2431, i_13_2538, i_13_2718, i_13_2719, i_13_2739, i_13_2740, i_13_2766, i_13_2781, i_13_2796, i_13_2797, i_13_2880, i_13_3066, i_13_3126, i_13_3133, i_13_3231, i_13_3240, i_13_3241, i_13_3309, i_13_3388, i_13_3414, i_13_3420, i_13_3460, i_13_3619, i_13_3636, i_13_3637, i_13_3682, i_13_3699, i_13_3717, i_13_3760, i_13_3762, i_13_3795, i_13_3843, i_13_3844, i_13_3862, i_13_3870, i_13_3906, i_13_3934, i_13_4050, i_13_4212, i_13_4326, i_13_4347, i_13_4350, i_13_4360, i_13_4387, i_13_4470, o_13_17);
	kernel_13_18 k_13_18(i_13_38, i_13_41, i_13_91, i_13_109, i_13_210, i_13_227, i_13_279, i_13_282, i_13_405, i_13_459, i_13_643, i_13_651, i_13_686, i_13_734, i_13_792, i_13_793, i_13_847, i_13_855, i_13_902, i_13_955, i_13_1017, i_13_1018, i_13_1020, i_13_1021, i_13_1120, i_13_1200, i_13_1270, i_13_1273, i_13_1308, i_13_1440, i_13_1459, i_13_1485, i_13_1486, i_13_1535, i_13_1548, i_13_1603, i_13_1629, i_13_1630, i_13_1639, i_13_1792, i_13_1813, i_13_1828, i_13_1832, i_13_1854, i_13_1998, i_13_2197, i_13_2205, i_13_2421, i_13_2435, i_13_2457, i_13_2458, i_13_2461, i_13_2467, i_13_2529, i_13_2538, i_13_2539, i_13_2542, i_13_2551, i_13_2712, i_13_2848, i_13_2916, i_13_2917, i_13_2918, i_13_3126, i_13_3160, i_13_3169, i_13_3268, i_13_3404, i_13_3407, i_13_3450, i_13_3460, i_13_3537, i_13_3551, i_13_3577, i_13_3663, i_13_3684, i_13_3726, i_13_3728, i_13_3754, i_13_3843, i_13_3853, i_13_3907, i_13_3910, i_13_3928, i_13_3987, i_13_4015, i_13_4033, i_13_4123, i_13_4186, i_13_4252, i_13_4322, i_13_4338, i_13_4341, i_13_4519, i_13_4522, i_13_4534, i_13_4558, i_13_4559, i_13_4591, i_13_4600, o_13_18);
	kernel_13_19 k_13_19(i_13_41, i_13_59, i_13_76, i_13_100, i_13_106, i_13_136, i_13_190, i_13_193, i_13_218, i_13_256, i_13_328, i_13_376, i_13_416, i_13_428, i_13_533, i_13_577, i_13_599, i_13_614, i_13_622, i_13_626, i_13_628, i_13_629, i_13_644, i_13_685, i_13_715, i_13_725, i_13_778, i_13_854, i_13_884, i_13_892, i_13_895, i_13_911, i_13_980, i_13_1022, i_13_1096, i_13_1124, i_13_1249, i_13_1256, i_13_1280, i_13_1391, i_13_1445, i_13_1462, i_13_1471, i_13_1483, i_13_1484, i_13_1541, i_13_1597, i_13_1643, i_13_1676, i_13_1678, i_13_1688, i_13_1691, i_13_1748, i_13_1757, i_13_1849, i_13_1855, i_13_1856, i_13_1858, i_13_1862, i_13_1883, i_13_2053, i_13_2209, i_13_2245, i_13_2434, i_13_2506, i_13_2507, i_13_2630, i_13_2717, i_13_2818, i_13_2845, i_13_2848, i_13_2849, i_13_2851, i_13_2857, i_13_2875, i_13_2878, i_13_2909, i_13_2911, i_13_2921, i_13_3064, i_13_3065, i_13_3118, i_13_3170, i_13_3265, i_13_3305, i_13_3433, i_13_3436, i_13_3766, i_13_3791, i_13_3818, i_13_3832, i_13_3869, i_13_3884, i_13_4297, i_13_4328, i_13_4379, i_13_4421, i_13_4441, i_13_4508, i_13_4607, o_13_19);
	kernel_13_20 k_13_20(i_13_45, i_13_75, i_13_117, i_13_139, i_13_162, i_13_167, i_13_178, i_13_184, i_13_211, i_13_336, i_13_419, i_13_517, i_13_562, i_13_571, i_13_574, i_13_607, i_13_746, i_13_814, i_13_815, i_13_875, i_13_910, i_13_955, i_13_1080, i_13_1084, i_13_1132, i_13_1192, i_13_1219, i_13_1220, i_13_1345, i_13_1404, i_13_1409, i_13_1465, i_13_1496, i_13_1525, i_13_1526, i_13_1552, i_13_1555, i_13_1642, i_13_1699, i_13_1782, i_13_1800, i_13_1857, i_13_1858, i_13_1886, i_13_1960, i_13_1961, i_13_2201, i_13_2209, i_13_2223, i_13_2239, i_13_2240, i_13_2259, i_13_2277, i_13_2296, i_13_2381, i_13_2407, i_13_2428, i_13_2508, i_13_2552, i_13_2712, i_13_2848, i_13_2857, i_13_2898, i_13_2938, i_13_3100, i_13_3101, i_13_3146, i_13_3169, i_13_3208, i_13_3244, i_13_3347, i_13_3419, i_13_3473, i_13_3490, i_13_3505, i_13_3542, i_13_3555, i_13_3592, i_13_3618, i_13_3641, i_13_3670, i_13_3739, i_13_3804, i_13_3859, i_13_3860, i_13_3899, i_13_3909, i_13_3911, i_13_3913, i_13_4012, i_13_4081, i_13_4096, i_13_4097, i_13_4147, i_13_4189, i_13_4237, i_13_4293, i_13_4315, i_13_4322, i_13_4433, o_13_20);
	kernel_13_21 k_13_21(i_13_69, i_13_70, i_13_78, i_13_124, i_13_286, i_13_313, i_13_375, i_13_385, i_13_411, i_13_448, i_13_520, i_13_535, i_13_588, i_13_646, i_13_672, i_13_673, i_13_682, i_13_699, i_13_700, i_13_843, i_13_844, i_13_886, i_13_934, i_13_980, i_13_1102, i_13_1104, i_13_1105, i_13_1122, i_13_1222, i_13_1275, i_13_1276, i_13_1302, i_13_1311, i_13_1312, i_13_1402, i_13_1403, i_13_1428, i_13_1437, i_13_1438, i_13_1510, i_13_1600, i_13_1663, i_13_1665, i_13_1723, i_13_1725, i_13_1735, i_13_1777, i_13_1779, i_13_1798, i_13_1887, i_13_1888, i_13_1933, i_13_1935, i_13_1936, i_13_1947, i_13_1948, i_13_1995, i_13_1996, i_13_2004, i_13_2014, i_13_2029, i_13_2139, i_13_2140, i_13_2379, i_13_2383, i_13_2480, i_13_2551, i_13_2569, i_13_2599, i_13_2616, i_13_2650, i_13_2679, i_13_2697, i_13_2698, i_13_2712, i_13_2770, i_13_2824, i_13_2851, i_13_2901, i_13_2923, i_13_2958, i_13_3031, i_13_3208, i_13_3595, i_13_3596, i_13_3613, i_13_3742, i_13_3787, i_13_3930, i_13_3931, i_13_4063, i_13_4260, i_13_4302, i_13_4308, i_13_4309, i_13_4450, i_13_4596, i_13_4597, i_13_4606, i_13_4607, o_13_21);
	kernel_13_22 k_13_22(i_13_142, i_13_169, i_13_224, i_13_240, i_13_310, i_13_327, i_13_328, i_13_340, i_13_367, i_13_472, i_13_529, i_13_553, i_13_599, i_13_607, i_13_618, i_13_619, i_13_620, i_13_670, i_13_689, i_13_699, i_13_725, i_13_780, i_13_824, i_13_912, i_13_980, i_13_1024, i_13_1078, i_13_1214, i_13_1259, i_13_1273, i_13_1483, i_13_1636, i_13_1687, i_13_1726, i_13_1749, i_13_1780, i_13_1781, i_13_1852, i_13_1888, i_13_1996, i_13_2020, i_13_2186, i_13_2200, i_13_2293, i_13_2391, i_13_2455, i_13_2461, i_13_2462, i_13_2464, i_13_2465, i_13_2470, i_13_2507, i_13_2509, i_13_2545, i_13_2633, i_13_2789, i_13_3109, i_13_3172, i_13_3174, i_13_3175, i_13_3262, i_13_3388, i_13_3409, i_13_3414, i_13_3415, i_13_3419, i_13_3432, i_13_3463, i_13_3477, i_13_3482, i_13_3535, i_13_3536, i_13_3544, i_13_3545, i_13_3562, i_13_3643, i_13_3666, i_13_3723, i_13_3734, i_13_3766, i_13_3910, i_13_3913, i_13_3914, i_13_3927, i_13_3928, i_13_4019, i_13_4099, i_13_4100, i_13_4126, i_13_4255, i_13_4333, i_13_4354, i_13_4381, i_13_4391, i_13_4396, i_13_4440, i_13_4449, i_13_4525, i_13_4534, i_13_4561, o_13_22);
	kernel_13_23 k_13_23(i_13_48, i_13_52, i_13_53, i_13_118, i_13_167, i_13_183, i_13_287, i_13_319, i_13_320, i_13_337, i_13_518, i_13_532, i_13_574, i_13_575, i_13_602, i_13_625, i_13_644, i_13_647, i_13_651, i_13_655, i_13_676, i_13_679, i_13_680, i_13_688, i_13_689, i_13_844, i_13_981, i_13_986, i_13_1048, i_13_1049, i_13_1070, i_13_1123, i_13_1124, i_13_1151, i_13_1228, i_13_1256, i_13_1385, i_13_1441, i_13_1465, i_13_1515, i_13_1519, i_13_1574, i_13_1712, i_13_1746, i_13_1751, i_13_1852, i_13_1857, i_13_1862, i_13_1888, i_13_2009, i_13_2050, i_13_2101, i_13_2136, i_13_2264, i_13_2267, i_13_2411, i_13_2556, i_13_2649, i_13_2651, i_13_2653, i_13_2654, i_13_2677, i_13_2678, i_13_2699, i_13_2722, i_13_2752, i_13_2753, i_13_2849, i_13_2984, i_13_3001, i_13_3146, i_13_3214, i_13_3217, i_13_3259, i_13_3260, i_13_3293, i_13_3398, i_13_3401, i_13_3437, i_13_3523, i_13_3734, i_13_3866, i_13_3888, i_13_3893, i_13_3909, i_13_3914, i_13_3991, i_13_3992, i_13_3995, i_13_4021, i_13_4067, i_13_4117, i_13_4307, i_13_4310, i_13_4318, i_13_4319, i_13_4513, i_13_4514, i_13_4556, i_13_4598, o_13_23);
	kernel_13_24 k_13_24(i_13_40, i_13_52, i_13_94, i_13_101, i_13_241, i_13_251, i_13_259, i_13_278, i_13_310, i_13_334, i_13_377, i_13_519, i_13_607, i_13_619, i_13_620, i_13_663, i_13_700, i_13_701, i_13_858, i_13_868, i_13_871, i_13_886, i_13_929, i_13_980, i_13_1024, i_13_1075, i_13_1078, i_13_1079, i_13_1213, i_13_1214, i_13_1265, i_13_1282, i_13_1283, i_13_1397, i_13_1408, i_13_1426, i_13_1441, i_13_1480, i_13_1535, i_13_1561, i_13_1573, i_13_1609, i_13_1637, i_13_1642, i_13_1715, i_13_1776, i_13_1921, i_13_2104, i_13_2149, i_13_2150, i_13_2201, i_13_2260, i_13_2294, i_13_2455, i_13_2456, i_13_2546, i_13_2596, i_13_2647, i_13_2707, i_13_2768, i_13_2788, i_13_2789, i_13_2901, i_13_2959, i_13_3002, i_13_3005, i_13_3037, i_13_3292, i_13_3410, i_13_3419, i_13_3435, i_13_3449, i_13_3462, i_13_3464, i_13_3520, i_13_3559, i_13_3647, i_13_3650, i_13_3688, i_13_3689, i_13_3712, i_13_3847, i_13_3904, i_13_3918, i_13_3966, i_13_3994, i_13_4030, i_13_4090, i_13_4091, i_13_4157, i_13_4218, i_13_4250, i_13_4256, i_13_4271, i_13_4354, i_13_4361, i_13_4396, i_13_4450, i_13_4526, i_13_4541, o_13_24);
	kernel_13_25 k_13_25(i_13_17, i_13_64, i_13_111, i_13_139, i_13_160, i_13_169, i_13_170, i_13_188, i_13_251, i_13_259, i_13_310, i_13_320, i_13_340, i_13_341, i_13_457, i_13_458, i_13_493, i_13_494, i_13_619, i_13_657, i_13_728, i_13_814, i_13_817, i_13_818, i_13_945, i_13_980, i_13_1070, i_13_1079, i_13_1129, i_13_1142, i_13_1273, i_13_1303, i_13_1304, i_13_1305, i_13_1349, i_13_1364, i_13_1440, i_13_1441, i_13_1492, i_13_1565, i_13_1623, i_13_1640, i_13_1786, i_13_1808, i_13_1816, i_13_1817, i_13_1831, i_13_1839, i_13_1943, i_13_1989, i_13_1996, i_13_2123, i_13_2140, i_13_2150, i_13_2232, i_13_2267, i_13_2430, i_13_2431, i_13_2470, i_13_2519, i_13_2719, i_13_2752, i_13_2788, i_13_2789, i_13_2860, i_13_2941, i_13_2942, i_13_2969, i_13_3032, i_13_3040, i_13_3112, i_13_3141, i_13_3162, i_13_3220, i_13_3221, i_13_3428, i_13_3527, i_13_3541, i_13_3689, i_13_3769, i_13_3816, i_13_3892, i_13_4049, i_13_4057, i_13_4058, i_13_4066, i_13_4077, i_13_4081, i_13_4094, i_13_4237, i_13_4274, i_13_4319, i_13_4350, i_13_4363, i_13_4391, i_13_4512, i_13_4519, i_13_4534, i_13_4594, i_13_4604, o_13_25);
	kernel_13_26 k_13_26(i_13_40, i_13_45, i_13_48, i_13_76, i_13_90, i_13_91, i_13_118, i_13_121, i_13_163, i_13_333, i_13_336, i_13_337, i_13_374, i_13_377, i_13_379, i_13_410, i_13_450, i_13_567, i_13_643, i_13_667, i_13_688, i_13_694, i_13_729, i_13_822, i_13_823, i_13_850, i_13_1063, i_13_1115, i_13_1120, i_13_1243, i_13_1267, i_13_1269, i_13_1341, i_13_1440, i_13_1441, i_13_1498, i_13_1782, i_13_1845, i_13_1924, i_13_1947, i_13_2116, i_13_2173, i_13_2197, i_13_2205, i_13_2206, i_13_2233, i_13_2235, i_13_2317, i_13_2421, i_13_2424, i_13_2539, i_13_2584, i_13_2613, i_13_2746, i_13_2781, i_13_2790, i_13_2853, i_13_2906, i_13_2916, i_13_2935, i_13_2966, i_13_2969, i_13_3016, i_13_3060, i_13_3108, i_13_3204, i_13_3213, i_13_3214, i_13_3217, i_13_3231, i_13_3234, i_13_3239, i_13_3241, i_13_3367, i_13_3398, i_13_3475, i_13_3477, i_13_3609, i_13_3717, i_13_3754, i_13_3817, i_13_3862, i_13_3870, i_13_3873, i_13_3889, i_13_3925, i_13_4014, i_13_4060, i_13_4158, i_13_4186, i_13_4189, i_13_4266, i_13_4267, i_13_4347, i_13_4348, i_13_4423, i_13_4530, i_13_4588, i_13_4594, i_13_4600, o_13_26);
	kernel_13_27 k_13_27(i_13_23, i_13_28, i_13_29, i_13_41, i_13_92, i_13_112, i_13_244, i_13_257, i_13_266, i_13_367, i_13_370, i_13_373, i_13_376, i_13_384, i_13_391, i_13_442, i_13_443, i_13_463, i_13_483, i_13_526, i_13_604, i_13_605, i_13_608, i_13_613, i_13_668, i_13_730, i_13_797, i_13_830, i_13_832, i_13_947, i_13_1082, i_13_1085, i_13_1145, i_13_1226, i_13_1271, i_13_1318, i_13_1423, i_13_1424, i_13_1473, i_13_1487, i_13_1496, i_13_1514, i_13_1571, i_13_1621, i_13_1721, i_13_1730, i_13_1750, i_13_1804, i_13_1837, i_13_1838, i_13_1840, i_13_1841, i_13_1851, i_13_2017, i_13_2112, i_13_2137, i_13_2170, i_13_2171, i_13_2173, i_13_2207, i_13_2380, i_13_2422, i_13_2423, i_13_2426, i_13_2431, i_13_2432, i_13_2435, i_13_2471, i_13_2579, i_13_2938, i_13_3018, i_13_3034, i_13_3127, i_13_3237, i_13_3260, i_13_3422, i_13_3425, i_13_3433, i_13_3503, i_13_3547, i_13_3622, i_13_3667, i_13_3763, i_13_3767, i_13_3871, i_13_3872, i_13_3875, i_13_3889, i_13_3964, i_13_4033, i_13_4047, i_13_4079, i_13_4089, i_13_4118, i_13_4343, i_13_4349, i_13_4351, i_13_4352, i_13_4541, i_13_4558, o_13_27);
	kernel_13_28 k_13_28(i_13_72, i_13_318, i_13_342, i_13_406, i_13_433, i_13_469, i_13_531, i_13_532, i_13_536, i_13_550, i_13_553, i_13_562, i_13_651, i_13_660, i_13_661, i_13_666, i_13_669, i_13_676, i_13_693, i_13_694, i_13_696, i_13_700, i_13_828, i_13_843, i_13_885, i_13_930, i_13_942, i_13_1098, i_13_1116, i_13_1117, i_13_1144, i_13_1263, i_13_1269, i_13_1279, i_13_1656, i_13_1657, i_13_1659, i_13_1660, i_13_1693, i_13_1719, i_13_1731, i_13_1774, i_13_1791, i_13_1836, i_13_1915, i_13_2016, i_13_2017, i_13_2339, i_13_2398, i_13_2413, i_13_2442, i_13_2460, i_13_2466, i_13_2467, i_13_2692, i_13_2844, i_13_2845, i_13_2881, i_13_2888, i_13_2925, i_13_2958, i_13_2983, i_13_3025, i_13_3061, i_13_3101, i_13_3114, i_13_3153, i_13_3207, i_13_3216, i_13_3258, i_13_3372, i_13_3531, i_13_3549, i_13_3579, i_13_3592, i_13_3639, i_13_3654, i_13_3703, i_13_3738, i_13_3739, i_13_3862, i_13_3875, i_13_3906, i_13_3987, i_13_4015, i_13_4077, i_13_4123, i_13_4185, i_13_4186, i_13_4212, i_13_4279, i_13_4323, i_13_4329, i_13_4339, i_13_4368, i_13_4512, i_13_4590, i_13_4599, i_13_4600, i_13_4602, o_13_28);
	kernel_13_29 k_13_29(i_13_49, i_13_69, i_13_94, i_13_282, i_13_321, i_13_327, i_13_328, i_13_375, i_13_411, i_13_529, i_13_547, i_13_598, i_13_624, i_13_717, i_13_745, i_13_780, i_13_796, i_13_825, i_13_826, i_13_861, i_13_862, i_13_894, i_13_912, i_13_922, i_13_1023, i_13_1077, i_13_1257, i_13_1258, i_13_1320, i_13_1321, i_13_1383, i_13_1410, i_13_1491, i_13_1501, i_13_1608, i_13_1635, i_13_1643, i_13_1762, i_13_1770, i_13_1777, i_13_1861, i_13_2032, i_13_2059, i_13_2060, i_13_2139, i_13_2185, i_13_2240, i_13_2310, i_13_2427, i_13_2454, i_13_2461, i_13_2613, i_13_2632, i_13_2653, i_13_2654, i_13_2679, i_13_2749, i_13_2762, i_13_2848, i_13_2883, i_13_2886, i_13_2966, i_13_3056, i_13_3145, i_13_3174, i_13_3175, i_13_3219, i_13_3347, i_13_3392, i_13_3417, i_13_3418, i_13_3432, i_13_3450, i_13_3463, i_13_3490, i_13_3535, i_13_3550, i_13_3562, i_13_3571, i_13_3579, i_13_3640, i_13_3702, i_13_3723, i_13_3733, i_13_3786, i_13_3793, i_13_3846, i_13_3876, i_13_3912, i_13_3913, i_13_3948, i_13_4012, i_13_4238, i_13_4274, i_13_4380, i_13_4381, i_13_4443, i_13_4560, i_13_4561, i_13_4597, o_13_29);
	kernel_13_30 k_13_30(i_13_108, i_13_121, i_13_274, i_13_275, i_13_309, i_13_310, i_13_337, i_13_357, i_13_454, i_13_558, i_13_559, i_13_562, i_13_618, i_13_633, i_13_658, i_13_850, i_13_851, i_13_1064, i_13_1081, i_13_1085, i_13_1228, i_13_1266, i_13_1309, i_13_1336, i_13_1396, i_13_1407, i_13_1471, i_13_1525, i_13_1549, i_13_1597, i_13_1621, i_13_1624, i_13_1629, i_13_1678, i_13_1719, i_13_1783, i_13_1787, i_13_1813, i_13_1841, i_13_1858, i_13_1914, i_13_1929, i_13_1936, i_13_1937, i_13_2110, i_13_2170, i_13_2202, i_13_2431, i_13_2542, i_13_2563, i_13_2564, i_13_2592, i_13_2709, i_13_2712, i_13_2768, i_13_2855, i_13_2859, i_13_2903, i_13_2916, i_13_2984, i_13_3061, i_13_3062, i_13_3096, i_13_3097, i_13_3100, i_13_3106, i_13_3153, i_13_3160, i_13_3217, i_13_3231, i_13_3232, i_13_3234, i_13_3235, i_13_3276, i_13_3285, i_13_3450, i_13_3496, i_13_3520, i_13_3537, i_13_3538, i_13_3600, i_13_3614, i_13_3682, i_13_3684, i_13_3685, i_13_3720, i_13_3753, i_13_3865, i_13_3878, i_13_3904, i_13_3937, i_13_4090, i_13_4091, i_13_4189, i_13_4249, i_13_4302, i_13_4351, i_13_4385, i_13_4517, i_13_4554, o_13_30);
	kernel_13_31 k_13_31(i_13_34, i_13_44, i_13_71, i_13_79, i_13_114, i_13_138, i_13_142, i_13_231, i_13_232, i_13_411, i_13_447, i_13_448, i_13_480, i_13_537, i_13_538, i_13_556, i_13_584, i_13_589, i_13_593, i_13_600, i_13_606, i_13_609, i_13_610, i_13_646, i_13_660, i_13_673, i_13_681, i_13_682, i_13_688, i_13_760, i_13_763, i_13_952, i_13_1119, i_13_1150, i_13_1275, i_13_1308, i_13_1311, i_13_1312, i_13_1344, i_13_1402, i_13_1428, i_13_1510, i_13_1626, i_13_1663, i_13_1672, i_13_1713, i_13_1725, i_13_1726, i_13_1734, i_13_1780, i_13_1798, i_13_1887, i_13_1911, i_13_1912, i_13_1923, i_13_1934, i_13_1947, i_13_1948, i_13_2175, i_13_2321, i_13_2379, i_13_2552, i_13_2598, i_13_2599, i_13_2679, i_13_2712, i_13_2752, i_13_2847, i_13_2850, i_13_2851, i_13_2856, i_13_2877, i_13_2923, i_13_3046, i_13_3067, i_13_3103, i_13_3129, i_13_3370, i_13_3371, i_13_3652, i_13_3668, i_13_3786, i_13_3930, i_13_3931, i_13_3940, i_13_4154, i_13_4188, i_13_4189, i_13_4219, i_13_4296, i_13_4297, i_13_4306, i_13_4308, i_13_4325, i_13_4336, i_13_4435, i_13_4450, i_13_4539, i_13_4596, i_13_4597, o_13_31);
	kernel_13_32 k_13_32(i_13_258, i_13_259, i_13_276, i_13_382, i_13_515, i_13_516, i_13_519, i_13_526, i_13_546, i_13_551, i_13_578, i_13_580, i_13_627, i_13_640, i_13_663, i_13_797, i_13_838, i_13_843, i_13_844, i_13_885, i_13_888, i_13_932, i_13_939, i_13_942, i_13_1077, i_13_1111, i_13_1119, i_13_1149, i_13_1222, i_13_1224, i_13_1230, i_13_1323, i_13_1404, i_13_1444, i_13_1464, i_13_1469, i_13_1483, i_13_1516, i_13_1552, i_13_1660, i_13_1677, i_13_1732, i_13_1734, i_13_1744, i_13_1745, i_13_1770, i_13_1830, i_13_1914, i_13_1915, i_13_1923, i_13_1947, i_13_1959, i_13_2002, i_13_2004, i_13_2019, i_13_2020, i_13_2022, i_13_2025, i_13_2197, i_13_2209, i_13_2320, i_13_2425, i_13_2722, i_13_2742, i_13_2860, i_13_2898, i_13_2938, i_13_2959, i_13_3030, i_13_3117, i_13_3156, i_13_3315, i_13_3351, i_13_3354, i_13_3355, i_13_3412, i_13_3418, i_13_3478, i_13_3525, i_13_3570, i_13_3684, i_13_3759, i_13_3763, i_13_3822, i_13_3864, i_13_3901, i_13_4029, i_13_4054, i_13_4063, i_13_4124, i_13_4161, i_13_4165, i_13_4230, i_13_4300, i_13_4303, i_13_4362, i_13_4567, i_13_4602, i_13_4605, i_13_4606, o_13_32);
	kernel_13_33 k_13_33(i_13_45, i_13_67, i_13_117, i_13_135, i_13_136, i_13_138, i_13_192, i_13_228, i_13_333, i_13_418, i_13_534, i_13_535, i_13_604, i_13_607, i_13_612, i_13_624, i_13_625, i_13_642, i_13_643, i_13_676, i_13_822, i_13_894, i_13_976, i_13_1116, i_13_1119, i_13_1120, i_13_1147, i_13_1272, i_13_1273, i_13_1390, i_13_1479, i_13_1642, i_13_1648, i_13_1669, i_13_1777, i_13_1795, i_13_1885, i_13_1886, i_13_1903, i_13_1944, i_13_1993, i_13_2230, i_13_2313, i_13_2361, i_13_2376, i_13_2379, i_13_2380, i_13_2397, i_13_2400, i_13_2401, i_13_2541, i_13_2578, i_13_2646, i_13_2647, i_13_2782, i_13_2847, i_13_2848, i_13_2874, i_13_2878, i_13_2898, i_13_2899, i_13_3036, i_13_3090, i_13_3091, i_13_3103, i_13_3117, i_13_3126, i_13_3250, i_13_3256, i_13_3261, i_13_3262, i_13_3352, i_13_3367, i_13_3384, i_13_3388, i_13_3508, i_13_3546, i_13_3547, i_13_3729, i_13_3730, i_13_3738, i_13_3835, i_13_3889, i_13_3919, i_13_4018, i_13_4060, i_13_4063, i_13_4185, i_13_4186, i_13_4209, i_13_4210, i_13_4293, i_13_4294, i_13_4320, i_13_4351, i_13_4480, i_13_4500, i_13_4537, i_13_4567, i_13_4594, o_13_33);
	kernel_13_34 k_13_34(i_13_53, i_13_76, i_13_121, i_13_134, i_13_184, i_13_232, i_13_251, i_13_286, i_13_357, i_13_358, i_13_359, i_13_466, i_13_467, i_13_468, i_13_592, i_13_680, i_13_745, i_13_842, i_13_916, i_13_1021, i_13_1025, i_13_1348, i_13_1349, i_13_1400, i_13_1501, i_13_1507, i_13_1516, i_13_1637, i_13_1644, i_13_1671, i_13_1727, i_13_1768, i_13_1816, i_13_1844, i_13_1951, i_13_1952, i_13_1961, i_13_2032, i_13_2033, i_13_2059, i_13_2060, i_13_2113, i_13_2203, i_13_2204, i_13_2284, i_13_2285, i_13_2321, i_13_2382, i_13_2398, i_13_2399, i_13_2509, i_13_2515, i_13_2554, i_13_2555, i_13_2570, i_13_2691, i_13_2752, i_13_2753, i_13_2902, i_13_2923, i_13_2924, i_13_2959, i_13_3013, i_13_3040, i_13_3131, i_13_3155, i_13_3163, i_13_3266, i_13_3373, i_13_3374, i_13_3392, i_13_3419, i_13_3580, i_13_3581, i_13_3598, i_13_3599, i_13_3622, i_13_3623, i_13_3634, i_13_3725, i_13_3787, i_13_3874, i_13_3877, i_13_3915, i_13_3923, i_13_3968, i_13_3991, i_13_3992, i_13_4175, i_13_4216, i_13_4256, i_13_4265, i_13_4316, i_13_4333, i_13_4334, i_13_4433, i_13_4453, i_13_4454, i_13_4507, i_13_4589, o_13_34);
	kernel_13_35 k_13_35(i_13_16, i_13_43, i_13_133, i_13_141, i_13_168, i_13_186, i_13_231, i_13_258, i_13_472, i_13_531, i_13_537, i_13_618, i_13_642, i_13_643, i_13_645, i_13_646, i_13_681, i_13_688, i_13_690, i_13_780, i_13_816, i_13_817, i_13_823, i_13_847, i_13_897, i_13_979, i_13_1122, i_13_1123, i_13_1128, i_13_1225, i_13_1275, i_13_1276, i_13_1464, i_13_1470, i_13_1552, i_13_1600, i_13_1645, i_13_1723, i_13_1725, i_13_1734, i_13_1780, i_13_1851, i_13_1887, i_13_1995, i_13_1996, i_13_2136, i_13_2196, i_13_2262, i_13_2266, i_13_2379, i_13_2382, i_13_2407, i_13_2409, i_13_2410, i_13_2422, i_13_2434, i_13_2542, i_13_2550, i_13_2587, i_13_2616, i_13_2650, i_13_2653, i_13_2698, i_13_2751, i_13_2760, i_13_2797, i_13_2877, i_13_2940, i_13_2941, i_13_3030, i_13_3039, i_13_3067, i_13_3112, i_13_3291, i_13_3423, i_13_3438, i_13_3484, i_13_3487, i_13_3526, i_13_3534, i_13_3724, i_13_3834, i_13_3874, i_13_3921, i_13_3994, i_13_4015, i_13_4099, i_13_4146, i_13_4216, i_13_4308, i_13_4309, i_13_4317, i_13_4318, i_13_4344, i_13_4354, i_13_4375, i_13_4432, i_13_4554, i_13_4563, i_13_4597, o_13_35);
	kernel_13_36 k_13_36(i_13_96, i_13_105, i_13_115, i_13_160, i_13_286, i_13_453, i_13_551, i_13_575, i_13_591, i_13_592, i_13_673, i_13_692, i_13_717, i_13_832, i_13_863, i_13_871, i_13_959, i_13_1024, i_13_1084, i_13_1132, i_13_1150, i_13_1232, i_13_1302, i_13_1303, i_13_1320, i_13_1464, i_13_1501, i_13_1556, i_13_1641, i_13_1732, i_13_1754, i_13_1759, i_13_1768, i_13_1772, i_13_1806, i_13_1807, i_13_1815, i_13_1816, i_13_1859, i_13_1886, i_13_1905, i_13_1961, i_13_2059, i_13_2103, i_13_2123, i_13_2139, i_13_2140, i_13_2141, i_13_2202, i_13_2284, i_13_2310, i_13_2366, i_13_2445, i_13_2446, i_13_2470, i_13_2545, i_13_2617, i_13_2640, i_13_2652, i_13_2654, i_13_2660, i_13_2663, i_13_2704, i_13_2711, i_13_2823, i_13_2824, i_13_2858, i_13_2910, i_13_2941, i_13_3049, i_13_3209, i_13_3219, i_13_3273, i_13_3374, i_13_3390, i_13_3391, i_13_3621, i_13_3622, i_13_3633, i_13_3661, i_13_3740, i_13_3786, i_13_3805, i_13_3868, i_13_3914, i_13_3991, i_13_4049, i_13_4057, i_13_4162, i_13_4233, i_13_4236, i_13_4371, i_13_4372, i_13_4380, i_13_4381, i_13_4382, i_13_4398, i_13_4399, i_13_4443, i_13_4452, o_13_36);
	kernel_13_37 k_13_37(i_13_30, i_13_37, i_13_116, i_13_120, i_13_126, i_13_133, i_13_135, i_13_136, i_13_324, i_13_327, i_13_454, i_13_487, i_13_544, i_13_570, i_13_576, i_13_594, i_13_595, i_13_597, i_13_616, i_13_684, i_13_714, i_13_777, i_13_828, i_13_891, i_13_910, i_13_1092, i_13_1246, i_13_1296, i_13_1300, i_13_1306, i_13_1369, i_13_1380, i_13_1461, i_13_1479, i_13_1480, i_13_1495, i_13_1552, i_13_1693, i_13_1710, i_13_1723, i_13_1746, i_13_1756, i_13_1782, i_13_1804, i_13_1869, i_13_1881, i_13_1903, i_13_1938, i_13_1939, i_13_2058, i_13_2136, i_13_2289, i_13_2307, i_13_2316, i_13_2317, i_13_2358, i_13_2454, i_13_2457, i_13_2458, i_13_2506, i_13_2596, i_13_2629, i_13_2646, i_13_2649, i_13_2748, i_13_2755, i_13_2820, i_13_2848, i_13_2907, i_13_2908, i_13_3010, i_13_3012, i_13_3013, i_13_3142, i_13_3171, i_13_3205, i_13_3216, i_13_3217, i_13_3234, i_13_3388, i_13_3406, i_13_3415, i_13_3429, i_13_3555, i_13_3556, i_13_3559, i_13_3610, i_13_3790, i_13_3910, i_13_3918, i_13_3988, i_13_4008, i_13_4009, i_13_4054, i_13_4078, i_13_4261, i_13_4263, i_13_4410, i_13_4440, i_13_4584, o_13_37);
	kernel_13_38 k_13_38(i_13_52, i_13_53, i_13_163, i_13_170, i_13_175, i_13_176, i_13_178, i_13_179, i_13_188, i_13_283, i_13_284, i_13_286, i_13_287, i_13_319, i_13_529, i_13_572, i_13_574, i_13_575, i_13_613, i_13_692, i_13_718, i_13_797, i_13_812, i_13_826, i_13_827, i_13_859, i_13_887, i_13_955, i_13_1019, i_13_1067, i_13_1070, i_13_1072, i_13_1252, i_13_1310, i_13_1313, i_13_1316, i_13_1447, i_13_1499, i_13_1501, i_13_1502, i_13_1523, i_13_1634, i_13_1636, i_13_1673, i_13_1676, i_13_1808, i_13_1849, i_13_1855, i_13_1861, i_13_2242, i_13_2263, i_13_2297, i_13_2410, i_13_2411, i_13_2428, i_13_2429, i_13_2465, i_13_2555, i_13_2612, i_13_2677, i_13_2681, i_13_2695, i_13_3110, i_13_3113, i_13_3209, i_13_3245, i_13_3272, i_13_3274, i_13_3275, i_13_3424, i_13_3425, i_13_3427, i_13_3428, i_13_3458, i_13_3485, i_13_3731, i_13_3733, i_13_3734, i_13_3770, i_13_3821, i_13_3838, i_13_3853, i_13_3854, i_13_3857, i_13_3875, i_13_3992, i_13_4018, i_13_4019, i_13_4021, i_13_4022, i_13_4085, i_13_4090, i_13_4253, i_13_4256, i_13_4264, i_13_4354, i_13_4510, i_13_4561, i_13_4562, i_13_4598, o_13_38);
	kernel_13_39 k_13_39(i_13_62, i_13_76, i_13_77, i_13_326, i_13_416, i_13_562, i_13_571, i_13_622, i_13_688, i_13_697, i_13_707, i_13_719, i_13_827, i_13_841, i_13_863, i_13_925, i_13_938, i_13_958, i_13_1022, i_13_1072, i_13_1073, i_13_1077, i_13_1219, i_13_1225, i_13_1228, i_13_1256, i_13_1259, i_13_1262, i_13_1280, i_13_1300, i_13_1315, i_13_1318, i_13_1319, i_13_1444, i_13_1445, i_13_1465, i_13_1553, i_13_1589, i_13_1606, i_13_1679, i_13_1774, i_13_1775, i_13_1778, i_13_1855, i_13_1858, i_13_1859, i_13_1914, i_13_1922, i_13_1982, i_13_1989, i_13_2000, i_13_2002, i_13_2056, i_13_2159, i_13_2173, i_13_2270, i_13_2461, i_13_2540, i_13_2630, i_13_2657, i_13_2677, i_13_2705, i_13_2774, i_13_2858, i_13_3010, i_13_3064, i_13_3091, i_13_3145, i_13_3173, i_13_3269, i_13_3308, i_13_3416, i_13_3449, i_13_3484, i_13_3487, i_13_3507, i_13_3541, i_13_3542, i_13_3544, i_13_3578, i_13_3634, i_13_3761, i_13_3803, i_13_3814, i_13_3863, i_13_4013, i_13_4018, i_13_4054, i_13_4253, i_13_4279, i_13_4333, i_13_4351, i_13_4370, i_13_4372, i_13_4376, i_13_4378, i_13_4379, i_13_4519, i_13_4520, i_13_4567, o_13_39);
	kernel_13_40 k_13_40(i_13_31, i_13_44, i_13_77, i_13_103, i_13_275, i_13_469, i_13_497, i_13_527, i_13_557, i_13_562, i_13_563, i_13_611, i_13_664, i_13_827, i_13_941, i_13_953, i_13_1021, i_13_1022, i_13_1025, i_13_1060, i_13_1075, i_13_1076, i_13_1139, i_13_1151, i_13_1256, i_13_1259, i_13_1270, i_13_1313, i_13_1318, i_13_1319, i_13_1333, i_13_1339, i_13_1372, i_13_1377, i_13_1553, i_13_1634, i_13_1691, i_13_1717, i_13_1723, i_13_1786, i_13_1804, i_13_1858, i_13_1861, i_13_1862, i_13_1942, i_13_1958, i_13_2026, i_13_2158, i_13_2197, i_13_2455, i_13_2476, i_13_2552, i_13_2618, i_13_2702, i_13_2744, i_13_2750, i_13_2921, i_13_2966, i_13_3010, i_13_3011, i_13_3014, i_13_3037, i_13_3163, i_13_3173, i_13_3226, i_13_3235, i_13_3245, i_13_3272, i_13_3443, i_13_3461, i_13_3479, i_13_3482, i_13_3487, i_13_3488, i_13_3491, i_13_3541, i_13_3542, i_13_3569, i_13_3571, i_13_3572, i_13_3574, i_13_3577, i_13_3578, i_13_3784, i_13_3785, i_13_3859, i_13_3895, i_13_3911, i_13_3960, i_13_4252, i_13_4253, i_13_4256, i_13_4258, i_13_4261, i_13_4262, i_13_4351, i_13_4372, i_13_4378, i_13_4447, i_13_4567, o_13_40);
	kernel_13_41 k_13_41(i_13_27, i_13_105, i_13_183, i_13_185, i_13_186, i_13_187, i_13_205, i_13_229, i_13_256, i_13_376, i_13_382, i_13_388, i_13_439, i_13_526, i_13_550, i_13_589, i_13_600, i_13_610, i_13_624, i_13_625, i_13_658, i_13_669, i_13_673, i_13_676, i_13_681, i_13_765, i_13_796, i_13_887, i_13_1111, i_13_1123, i_13_1144, i_13_1150, i_13_1195, i_13_1201, i_13_1270, i_13_1326, i_13_1327, i_13_1363, i_13_1404, i_13_1497, i_13_1503, i_13_1515, i_13_1516, i_13_1653, i_13_1677, i_13_1678, i_13_1680, i_13_1714, i_13_1729, i_13_1733, i_13_1741, i_13_1834, i_13_1839, i_13_1857, i_13_1860, i_13_1909, i_13_1911, i_13_1912, i_13_1999, i_13_2001, i_13_2002, i_13_2020, i_13_2175, i_13_2176, i_13_2200, i_13_2363, i_13_2556, i_13_2616, i_13_2722, i_13_2727, i_13_2760, i_13_2793, i_13_2857, i_13_2860, i_13_2973, i_13_3000, i_13_3028, i_13_3087, i_13_3090, i_13_3121, i_13_3382, i_13_3460, i_13_3522, i_13_3546, i_13_3552, i_13_3685, i_13_3730, i_13_3766, i_13_3864, i_13_3925, i_13_4054, i_13_4080, i_13_4186, i_13_4200, i_13_4393, i_13_4480, i_13_4567, i_13_4581, i_13_4600, i_13_4602, o_13_41);
	kernel_13_42 k_13_42(i_13_40, i_13_90, i_13_129, i_13_130, i_13_156, i_13_190, i_13_270, i_13_273, i_13_336, i_13_418, i_13_453, i_13_468, i_13_490, i_13_526, i_13_558, i_13_561, i_13_562, i_13_633, i_13_657, i_13_724, i_13_732, i_13_742, i_13_823, i_13_838, i_13_945, i_13_1083, i_13_1084, i_13_1143, i_13_1147, i_13_1242, i_13_1350, i_13_1470, i_13_1620, i_13_1650, i_13_1768, i_13_1785, i_13_1812, i_13_1840, i_13_1857, i_13_1936, i_13_2001, i_13_2205, i_13_2430, i_13_2497, i_13_2529, i_13_2546, i_13_2649, i_13_2650, i_13_2664, i_13_2709, i_13_2784, i_13_2982, i_13_3019, i_13_3043, i_13_3046, i_13_3070, i_13_3097, i_13_3099, i_13_3100, i_13_3135, i_13_3141, i_13_3213, i_13_3231, i_13_3234, i_13_3252, i_13_3351, i_13_3388, i_13_3415, i_13_3487, i_13_3541, i_13_3549, i_13_3603, i_13_3636, i_13_3640, i_13_3655, i_13_3682, i_13_3685, i_13_3699, i_13_3730, i_13_3747, i_13_3762, i_13_3870, i_13_3897, i_13_3909, i_13_3979, i_13_3981, i_13_3982, i_13_4158, i_13_4159, i_13_4161, i_13_4162, i_13_4164, i_13_4177, i_13_4194, i_13_4195, i_13_4269, i_13_4321, i_13_4324, i_13_4428, i_13_4539, o_13_42);
	kernel_13_43 k_13_43(i_13_31, i_13_49, i_13_63, i_13_66, i_13_67, i_13_136, i_13_140, i_13_211, i_13_227, i_13_228, i_13_285, i_13_409, i_13_447, i_13_490, i_13_537, i_13_609, i_13_612, i_13_614, i_13_645, i_13_649, i_13_672, i_13_684, i_13_686, i_13_699, i_13_771, i_13_814, i_13_820, i_13_982, i_13_1066, i_13_1116, i_13_1117, i_13_1118, i_13_1119, i_13_1225, i_13_1226, i_13_1270, i_13_1274, i_13_1307, i_13_1327, i_13_1388, i_13_1411, i_13_1427, i_13_1489, i_13_1513, i_13_1539, i_13_1570, i_13_1639, i_13_1672, i_13_1723, i_13_1732, i_13_1793, i_13_1795, i_13_1801, i_13_1849, i_13_1885, i_13_1909, i_13_2056, i_13_2128, i_13_2135, i_13_2297, i_13_2407, i_13_2408, i_13_2423, i_13_2433, i_13_2434, i_13_2635, i_13_2719, i_13_2722, i_13_2847, i_13_2848, i_13_2850, i_13_2875, i_13_3037, i_13_3093, i_13_3165, i_13_3268, i_13_3387, i_13_3400, i_13_3520, i_13_3537, i_13_3539, i_13_3577, i_13_3741, i_13_3766, i_13_3793, i_13_3836, i_13_3837, i_13_3894, i_13_3924, i_13_3965, i_13_4033, i_13_4043, i_13_4053, i_13_4078, i_13_4216, i_13_4294, i_13_4295, i_13_4296, i_13_4297, i_13_4376, o_13_43);
	kernel_13_44 k_13_44(i_13_31, i_13_61, i_13_99, i_13_116, i_13_184, i_13_186, i_13_187, i_13_229, i_13_258, i_13_259, i_13_426, i_13_431, i_13_526, i_13_601, i_13_618, i_13_619, i_13_620, i_13_628, i_13_670, i_13_691, i_13_756, i_13_799, i_13_800, i_13_840, i_13_962, i_13_1024, i_13_1077, i_13_1079, i_13_1123, i_13_1184, i_13_1187, i_13_1411, i_13_1444, i_13_1457, i_13_1482, i_13_1483, i_13_1519, i_13_1529, i_13_1573, i_13_1637, i_13_1677, i_13_1681, i_13_1747, i_13_1753, i_13_1771, i_13_1806, i_13_1807, i_13_1817, i_13_1861, i_13_1908, i_13_1912, i_13_1930, i_13_2001, i_13_2002, i_13_2003, i_13_2005, i_13_2024, i_13_2139, i_13_2140, i_13_2223, i_13_2224, i_13_2248, i_13_2259, i_13_2425, i_13_2446, i_13_2482, i_13_2653, i_13_2722, i_13_2743, i_13_2745, i_13_2751, i_13_2789, i_13_2798, i_13_2807, i_13_2857, i_13_3030, i_13_3122, i_13_3221, i_13_3244, i_13_3291, i_13_3293, i_13_3405, i_13_3439, i_13_3464, i_13_3525, i_13_3532, i_13_3552, i_13_3553, i_13_3759, i_13_3869, i_13_3905, i_13_4044, i_13_4054, i_13_4094, i_13_4152, i_13_4189, i_13_4317, i_13_4363, i_13_4387, i_13_4390, o_13_44);
	kernel_13_45 k_13_45(i_13_36, i_13_37, i_13_80, i_13_179, i_13_314, i_13_324, i_13_431, i_13_525, i_13_531, i_13_544, i_13_553, i_13_554, i_13_557, i_13_570, i_13_576, i_13_595, i_13_611, i_13_662, i_13_682, i_13_683, i_13_701, i_13_714, i_13_724, i_13_777, i_13_845, i_13_891, i_13_895, i_13_927, i_13_1041, i_13_1092, i_13_1151, i_13_1214, i_13_1369, i_13_1380, i_13_1399, i_13_1430, i_13_1461, i_13_1479, i_13_1480, i_13_1484, i_13_1596, i_13_1634, i_13_1710, i_13_1719, i_13_1720, i_13_1736, i_13_1767, i_13_1781, i_13_1782, i_13_1792, i_13_1881, i_13_1882, i_13_1952, i_13_2048, i_13_2129, i_13_2164, i_13_2210, i_13_2224, i_13_2236, i_13_2277, i_13_2307, i_13_2457, i_13_2600, i_13_2610, i_13_2629, i_13_2646, i_13_2649, i_13_2726, i_13_2820, i_13_2844, i_13_2845, i_13_2871, i_13_2885, i_13_3216, i_13_3420, i_13_3429, i_13_3448, i_13_3599, i_13_3743, i_13_3758, i_13_3784, i_13_3790, i_13_3866, i_13_3902, i_13_3924, i_13_3941, i_13_4014, i_13_4077, i_13_4114, i_13_4257, i_13_4265, i_13_4337, i_13_4360, i_13_4361, i_13_4436, i_13_4440, i_13_4540, i_13_4594, i_13_4598, i_13_4607, o_13_45);
	kernel_13_46 k_13_46(i_13_114, i_13_127, i_13_159, i_13_160, i_13_166, i_13_211, i_13_241, i_13_247, i_13_268, i_13_269, i_13_275, i_13_319, i_13_340, i_13_357, i_13_375, i_13_443, i_13_465, i_13_466, i_13_519, i_13_520, i_13_536, i_13_643, i_13_699, i_13_714, i_13_744, i_13_745, i_13_762, i_13_862, i_13_947, i_13_1123, i_13_1212, i_13_1213, i_13_1255, i_13_1303, i_13_1347, i_13_1400, i_13_1411, i_13_1428, i_13_1456, i_13_1482, i_13_1483, i_13_1774, i_13_1775, i_13_1813, i_13_1816, i_13_1945, i_13_1946, i_13_2059, i_13_2132, i_13_2181, i_13_2202, i_13_2283, i_13_2284, i_13_2285, i_13_2354, i_13_2417, i_13_2496, i_13_2715, i_13_2724, i_13_2725, i_13_2770, i_13_2771, i_13_2788, i_13_2792, i_13_2938, i_13_3048, i_13_3056, i_13_3063, i_13_3068, i_13_3122, i_13_3144, i_13_3220, i_13_3235, i_13_3271, i_13_3373, i_13_3419, i_13_3441, i_13_3453, i_13_3523, i_13_3530, i_13_3597, i_13_3598, i_13_3617, i_13_3621, i_13_3635, i_13_3666, i_13_3685, i_13_3824, i_13_3875, i_13_3922, i_13_4057, i_13_4081, i_13_4093, i_13_4184, i_13_4197, i_13_4261, i_13_4272, i_13_4273, i_13_4274, i_13_4399, o_13_46);
	kernel_13_47 k_13_47(i_13_63, i_13_97, i_13_124, i_13_125, i_13_140, i_13_187, i_13_188, i_13_196, i_13_328, i_13_374, i_13_520, i_13_536, i_13_552, i_13_574, i_13_577, i_13_580, i_13_583, i_13_592, i_13_603, i_13_641, i_13_664, i_13_715, i_13_718, i_13_729, i_13_745, i_13_781, i_13_793, i_13_800, i_13_862, i_13_863, i_13_886, i_13_989, i_13_1025, i_13_1135, i_13_1193, i_13_1258, i_13_1411, i_13_1447, i_13_1457, i_13_1493, i_13_1502, i_13_1573, i_13_1627, i_13_1636, i_13_1744, i_13_1751, i_13_1787, i_13_1831, i_13_1836, i_13_1859, i_13_1871, i_13_1885, i_13_1952, i_13_2015, i_13_2029, i_13_2168, i_13_2177, i_13_2267, i_13_2362, i_13_2383, i_13_2428, i_13_2465, i_13_2503, i_13_2536, i_13_2537, i_13_2633, i_13_2770, i_13_2825, i_13_2984, i_13_3004, i_13_3040, i_13_3159, i_13_3167, i_13_3175, i_13_3246, i_13_3290, i_13_3322, i_13_3323, i_13_3427, i_13_3428, i_13_3466, i_13_3581, i_13_3617, i_13_3699, i_13_3748, i_13_3787, i_13_3794, i_13_3806, i_13_3839, i_13_3877, i_13_3914, i_13_3922, i_13_4012, i_13_4013, i_13_4081, i_13_4171, i_13_4522, i_13_4566, i_13_4586, i_13_4588, o_13_47);
	kernel_13_48 k_13_48(i_13_37, i_13_59, i_13_136, i_13_167, i_13_230, i_13_260, i_13_283, i_13_308, i_13_545, i_13_577, i_13_596, i_13_617, i_13_625, i_13_626, i_13_646, i_13_671, i_13_717, i_13_728, i_13_778, i_13_779, i_13_838, i_13_839, i_13_852, i_13_865, i_13_911, i_13_956, i_13_1022, i_13_1094, i_13_1097, i_13_1118, i_13_1121, i_13_1146, i_13_1228, i_13_1281, i_13_1301, i_13_1318, i_13_1462, i_13_1464, i_13_1480, i_13_1481, i_13_1484, i_13_1522, i_13_1643, i_13_1675, i_13_1678, i_13_1688, i_13_1691, i_13_1721, i_13_1747, i_13_1750, i_13_1757, i_13_1768, i_13_1804, i_13_1805, i_13_1857, i_13_1858, i_13_1860, i_13_2002, i_13_2120, i_13_2138, i_13_2139, i_13_2165, i_13_2225, i_13_2308, i_13_2380, i_13_2425, i_13_2443, i_13_2444, i_13_2446, i_13_2447, i_13_2647, i_13_2650, i_13_2692, i_13_2693, i_13_2822, i_13_2999, i_13_3012, i_13_3076, i_13_3094, i_13_3110, i_13_3197, i_13_3290, i_13_3320, i_13_3353, i_13_3430, i_13_3560, i_13_3741, i_13_3911, i_13_3989, i_13_4115, i_13_4187, i_13_4189, i_13_4235, i_13_4263, i_13_4300, i_13_4351, i_13_4352, i_13_4379, i_13_4396, i_13_4441, o_13_48);
	kernel_13_49 k_13_49(i_13_22, i_13_61, i_13_79, i_13_94, i_13_95, i_13_259, i_13_261, i_13_319, i_13_322, i_13_336, i_13_492, i_13_521, i_13_619, i_13_697, i_13_700, i_13_745, i_13_823, i_13_835, i_13_837, i_13_870, i_13_960, i_13_970, i_13_978, i_13_979, i_13_980, i_13_1025, i_13_1075, i_13_1076, i_13_1095, i_13_1213, i_13_1281, i_13_1283, i_13_1302, i_13_1320, i_13_1321, i_13_1364, i_13_1384, i_13_1434, i_13_1438, i_13_1444, i_13_1464, i_13_1483, i_13_1568, i_13_1658, i_13_1813, i_13_1816, i_13_1817, i_13_1830, i_13_1870, i_13_1921, i_13_1943, i_13_1951, i_13_2082, i_13_2176, i_13_2209, i_13_2248, i_13_2425, i_13_2445, i_13_2446, i_13_2447, i_13_2460, i_13_2511, i_13_2516, i_13_2542, i_13_2554, i_13_2619, i_13_2923, i_13_3004, i_13_3056, i_13_3077, i_13_3094, i_13_3130, i_13_3220, i_13_3306, i_13_3418, i_13_3419, i_13_3433, i_13_3444, i_13_3482, i_13_3490, i_13_3550, i_13_3598, i_13_3737, i_13_3821, i_13_3874, i_13_3888, i_13_3992, i_13_4004, i_13_4018, i_13_4087, i_13_4188, i_13_4273, i_13_4333, i_13_4347, i_13_4351, i_13_4354, i_13_4381, i_13_4382, i_13_4390, i_13_4586, o_13_49);
	kernel_13_50 k_13_50(i_13_72, i_13_75, i_13_78, i_13_112, i_13_141, i_13_240, i_13_250, i_13_258, i_13_282, i_13_310, i_13_372, i_13_559, i_13_579, i_13_618, i_13_619, i_13_697, i_13_699, i_13_816, i_13_843, i_13_931, i_13_1023, i_13_1024, i_13_1077, i_13_1078, i_13_1084, i_13_1143, i_13_1204, i_13_1212, i_13_1255, i_13_1273, i_13_1284, i_13_1317, i_13_1332, i_13_1348, i_13_1427, i_13_1468, i_13_1513, i_13_1521, i_13_1572, i_13_1573, i_13_1597, i_13_1609, i_13_1633, i_13_1635, i_13_1725, i_13_1812, i_13_1843, i_13_1849, i_13_1881, i_13_1888, i_13_2103, i_13_2198, i_13_2278, i_13_2404, i_13_2442, i_13_2454, i_13_2563, i_13_2710, i_13_2712, i_13_2715, i_13_2742, i_13_2887, i_13_2955, i_13_2958, i_13_3036, i_13_3169, i_13_3204, i_13_3208, i_13_3241, i_13_3244, i_13_3291, i_13_3379, i_13_3412, i_13_3450, i_13_3451, i_13_3453, i_13_3454, i_13_3462, i_13_3525, i_13_3532, i_13_3570, i_13_3571, i_13_3649, i_13_3684, i_13_3685, i_13_3687, i_13_3688, i_13_3708, i_13_3756, i_13_3757, i_13_3781, i_13_3982, i_13_4020, i_13_4188, i_13_4233, i_13_4260, i_13_4312, i_13_4393, i_13_4497, i_13_4509, o_13_50);
	kernel_13_51 k_13_51(i_13_35, i_13_76, i_13_94, i_13_121, i_13_184, i_13_193, i_13_241, i_13_251, i_13_260, i_13_278, i_13_358, i_13_361, i_13_521, i_13_527, i_13_535, i_13_616, i_13_652, i_13_664, i_13_715, i_13_896, i_13_898, i_13_1024, i_13_1025, i_13_1078, i_13_1079, i_13_1211, i_13_1213, i_13_1244, i_13_1259, i_13_1286, i_13_1331, i_13_1349, i_13_1400, i_13_1408, i_13_1424, i_13_1427, i_13_1430, i_13_1483, i_13_1501, i_13_1502, i_13_1508, i_13_1609, i_13_1637, i_13_1696, i_13_1817, i_13_1835, i_13_1841, i_13_1921, i_13_1943, i_13_1961, i_13_2005, i_13_2006, i_13_2033, i_13_2131, i_13_2201, i_13_2315, i_13_2360, i_13_2455, i_13_2456, i_13_2471, i_13_2546, i_13_2573, i_13_2651, i_13_2716, i_13_2717, i_13_2726, i_13_2768, i_13_2923, i_13_2924, i_13_2959, i_13_2965, i_13_3163, i_13_3373, i_13_3374, i_13_3419, i_13_3565, i_13_3580, i_13_3599, i_13_3650, i_13_3731, i_13_3733, i_13_3734, i_13_3787, i_13_3905, i_13_3910, i_13_3919, i_13_3923, i_13_3985, i_13_4253, i_13_4255, i_13_4256, i_13_4262, i_13_4265, i_13_4453, i_13_4454, i_13_4526, i_13_4541, i_13_4558, i_13_4559, i_13_4561, o_13_51);
	kernel_13_52 k_13_52(i_13_2, i_13_78, i_13_180, i_13_184, i_13_185, i_13_187, i_13_189, i_13_192, i_13_193, i_13_283, i_13_324, i_13_370, i_13_509, i_13_517, i_13_533, i_13_570, i_13_571, i_13_594, i_13_640, i_13_641, i_13_714, i_13_715, i_13_718, i_13_798, i_13_858, i_13_887, i_13_939, i_13_958, i_13_1116, i_13_1193, i_13_1219, i_13_1228, i_13_1229, i_13_1254, i_13_1299, i_13_1314, i_13_1407, i_13_1408, i_13_1435, i_13_1464, i_13_1479, i_13_1530, i_13_1597, i_13_1639, i_13_1674, i_13_1713, i_13_1732, i_13_1741, i_13_1761, i_13_1762, i_13_1764, i_13_1769, i_13_1782, i_13_1785, i_13_1786, i_13_1801, i_13_1804, i_13_1957, i_13_2017, i_13_2055, i_13_2210, i_13_2280, i_13_2365, i_13_2397, i_13_2502, i_13_2567, i_13_2619, i_13_2693, i_13_2713, i_13_2857, i_13_3025, i_13_3030, i_13_3034, i_13_3045, i_13_3046, i_13_3163, i_13_3168, i_13_3259, i_13_3265, i_13_3286, i_13_3287, i_13_3352, i_13_3403, i_13_3423, i_13_3424, i_13_3754, i_13_3756, i_13_3759, i_13_3972, i_13_3979, i_13_3981, i_13_3984, i_13_4042, i_13_4086, i_13_4187, i_13_4199, i_13_4363, i_13_4434, i_13_4537, i_13_4565, o_13_52);
	kernel_13_53 k_13_53(i_13_172, i_13_192, i_13_199, i_13_280, i_13_324, i_13_361, i_13_378, i_13_525, i_13_570, i_13_576, i_13_639, i_13_640, i_13_685, i_13_714, i_13_777, i_13_810, i_13_858, i_13_891, i_13_927, i_13_948, i_13_954, i_13_1020, i_13_1026, i_13_1059, i_13_1063, i_13_1098, i_13_1209, i_13_1224, i_13_1225, i_13_1227, i_13_1254, i_13_1263, i_13_1296, i_13_1297, i_13_1407, i_13_1443, i_13_1498, i_13_1539, i_13_1594, i_13_1632, i_13_1710, i_13_1719, i_13_1747, i_13_1767, i_13_1782, i_13_1792, i_13_1800, i_13_1801, i_13_1857, i_13_1881, i_13_1926, i_13_1990, i_13_2011, i_13_2100, i_13_2116, i_13_2259, i_13_2358, i_13_2403, i_13_2460, i_13_2514, i_13_2532, i_13_2629, i_13_2646, i_13_2844, i_13_2853, i_13_2899, i_13_2934, i_13_2980, i_13_3105, i_13_3171, i_13_3241, i_13_3259, i_13_3267, i_13_3268, i_13_3285, i_13_3286, i_13_3325, i_13_3420, i_13_3421, i_13_3423, i_13_3447, i_13_3790, i_13_3873, i_13_3970, i_13_3991, i_13_4008, i_13_4009, i_13_4041, i_13_4042, i_13_4077, i_13_4086, i_13_4087, i_13_4153, i_13_4231, i_13_4248, i_13_4267, i_13_4278, i_13_4293, i_13_4410, i_13_4584, o_13_53);
	kernel_13_54 k_13_54(i_13_31, i_13_58, i_13_67, i_13_130, i_13_139, i_13_183, i_13_184, i_13_192, i_13_219, i_13_255, i_13_361, i_13_373, i_13_382, i_13_390, i_13_549, i_13_624, i_13_685, i_13_717, i_13_777, i_13_822, i_13_891, i_13_894, i_13_897, i_13_975, i_13_976, i_13_1093, i_13_1108, i_13_1116, i_13_1120, i_13_1145, i_13_1308, i_13_1314, i_13_1345, i_13_1380, i_13_1386, i_13_1387, i_13_1393, i_13_1407, i_13_1461, i_13_1476, i_13_1479, i_13_1480, i_13_1487, i_13_1498, i_13_1513, i_13_1526, i_13_1585, i_13_1597, i_13_1669, i_13_1674, i_13_1677, i_13_1690, i_13_1731, i_13_1749, i_13_1752, i_13_1756, i_13_1803, i_13_1956, i_13_2017, i_13_2190, i_13_2191, i_13_2442, i_13_2443, i_13_2449, i_13_2461, i_13_2479, i_13_2539, i_13_2559, i_13_2632, i_13_2676, i_13_2686, i_13_2739, i_13_2751, i_13_2895, i_13_2967, i_13_2997, i_13_3001, i_13_3114, i_13_3199, i_13_3261, i_13_3348, i_13_3352, i_13_3433, i_13_3468, i_13_3478, i_13_3520, i_13_3522, i_13_3525, i_13_3561, i_13_3567, i_13_3756, i_13_3865, i_13_3981, i_13_4294, i_13_4348, i_13_4351, i_13_4363, i_13_4413, i_13_4532, i_13_4591, o_13_54);
	kernel_13_55 k_13_55(i_13_47, i_13_92, i_13_94, i_13_95, i_13_139, i_13_170, i_13_173, i_13_175, i_13_178, i_13_214, i_13_215, i_13_311, i_13_362, i_13_441, i_13_452, i_13_535, i_13_555, i_13_569, i_13_571, i_13_572, i_13_609, i_13_659, i_13_662, i_13_686, i_13_847, i_13_851, i_13_854, i_13_951, i_13_956, i_13_986, i_13_1120, i_13_1229, i_13_1250, i_13_1260, i_13_1307, i_13_1311, i_13_1408, i_13_1422, i_13_1513, i_13_1514, i_13_1527, i_13_1540, i_13_1567, i_13_1723, i_13_1766, i_13_1791, i_13_1802, i_13_1829, i_13_1832, i_13_1847, i_13_1850, i_13_1858, i_13_1885, i_13_2108, i_13_2150, i_13_2227, i_13_2234, i_13_2297, i_13_2410, i_13_2467, i_13_2677, i_13_2680, i_13_2696, i_13_2713, i_13_2740, i_13_2934, i_13_2980, i_13_2985, i_13_3007, i_13_3011, i_13_3012, i_13_3025, i_13_3026, i_13_3064, i_13_3109, i_13_3110, i_13_3113, i_13_3208, i_13_3217, i_13_3268, i_13_3269, i_13_3386, i_13_3519, i_13_3739, i_13_3755, i_13_3764, i_13_3818, i_13_3879, i_13_3987, i_13_4061, i_13_4064, i_13_4371, i_13_4375, i_13_4432, i_13_4472, i_13_4514, i_13_4565, i_13_4568, i_13_4569, i_13_4591, o_13_55);
	kernel_13_56 k_13_56(i_13_40, i_13_76, i_13_133, i_13_192, i_13_251, i_13_283, i_13_318, i_13_334, i_13_336, i_13_358, i_13_457, i_13_492, i_13_493, i_13_620, i_13_715, i_13_758, i_13_813, i_13_829, i_13_876, i_13_956, i_13_1025, i_13_1100, i_13_1102, i_13_1230, i_13_1257, i_13_1300, i_13_1303, i_13_1327, i_13_1405, i_13_1446, i_13_1447, i_13_1502, i_13_1525, i_13_1640, i_13_1641, i_13_1698, i_13_1722, i_13_1723, i_13_1742, i_13_1785, i_13_1793, i_13_1794, i_13_1835, i_13_1937, i_13_2014, i_13_2056, i_13_2060, i_13_2103, i_13_2118, i_13_2146, i_13_2185, i_13_2236, i_13_2237, i_13_2239, i_13_2365, i_13_2407, i_13_2427, i_13_2445, i_13_2452, i_13_2535, i_13_2587, i_13_2617, i_13_2721, i_13_2922, i_13_2924, i_13_2937, i_13_3032, i_13_3036, i_13_3217, i_13_3219, i_13_3220, i_13_3234, i_13_3243, i_13_3244, i_13_3343, i_13_3424, i_13_3480, i_13_3550, i_13_3639, i_13_3649, i_13_3700, i_13_3702, i_13_3757, i_13_3766, i_13_3846, i_13_3865, i_13_3878, i_13_3889, i_13_3984, i_13_3985, i_13_4054, i_13_4213, i_13_4237, i_13_4273, i_13_4315, i_13_4400, i_13_4510, i_13_4513, i_13_4561, i_13_4587, o_13_56);
	kernel_13_57 k_13_57(i_13_63, i_13_76, i_13_136, i_13_339, i_13_340, i_13_357, i_13_358, i_13_534, i_13_535, i_13_546, i_13_579, i_13_645, i_13_687, i_13_690, i_13_697, i_13_825, i_13_915, i_13_1066, i_13_1213, i_13_1303, i_13_1306, i_13_1321, i_13_1347, i_13_1383, i_13_1446, i_13_1465, i_13_1501, i_13_1518, i_13_1642, i_13_1722, i_13_1723, i_13_1740, i_13_1815, i_13_1845, i_13_1950, i_13_1951, i_13_1960, i_13_2005, i_13_2023, i_13_2032, i_13_2058, i_13_2106, i_13_2110, i_13_2320, i_13_2428, i_13_2446, i_13_2514, i_13_2554, i_13_2640, i_13_2644, i_13_2649, i_13_2652, i_13_2677, i_13_2692, i_13_2751, i_13_2763, i_13_2847, i_13_2848, i_13_2913, i_13_2920, i_13_2922, i_13_2923, i_13_2958, i_13_2962, i_13_3028, i_13_3144, i_13_3219, i_13_3372, i_13_3373, i_13_3391, i_13_3393, i_13_3418, i_13_3444, i_13_3577, i_13_3595, i_13_3597, i_13_3598, i_13_3621, i_13_3669, i_13_3721, i_13_3741, i_13_3787, i_13_3793, i_13_3928, i_13_3990, i_13_3991, i_13_4021, i_13_4191, i_13_4237, i_13_4263, i_13_4264, i_13_4315, i_13_4332, i_13_4333, i_13_4350, i_13_4381, i_13_4398, i_13_4435, i_13_4452, i_13_4453, o_13_57);
	kernel_13_58 k_13_58(i_13_42, i_13_78, i_13_111, i_13_194, i_13_199, i_13_276, i_13_282, i_13_285, i_13_310, i_13_384, i_13_417, i_13_418, i_13_448, i_13_519, i_13_520, i_13_535, i_13_553, i_13_643, i_13_670, i_13_838, i_13_873, i_13_935, i_13_952, i_13_1020, i_13_1021, i_13_1023, i_13_1024, i_13_1075, i_13_1203, i_13_1254, i_13_1317, i_13_1390, i_13_1428, i_13_1429, i_13_1600, i_13_1605, i_13_1626, i_13_1632, i_13_1642, i_13_1777, i_13_1779, i_13_1780, i_13_1807, i_13_1813, i_13_1933, i_13_1940, i_13_2159, i_13_2199, i_13_2356, i_13_2454, i_13_2464, i_13_2541, i_13_2542, i_13_2575, i_13_2583, i_13_2617, i_13_2708, i_13_2769, i_13_2770, i_13_2847, i_13_2904, i_13_2919, i_13_2920, i_13_3031, i_13_3045, i_13_3246, i_13_3261, i_13_3353, i_13_3415, i_13_3453, i_13_3454, i_13_3456, i_13_3457, i_13_3459, i_13_3460, i_13_3462, i_13_3463, i_13_3534, i_13_3535, i_13_3541, i_13_3544, i_13_3558, i_13_3576, i_13_3619, i_13_3739, i_13_3783, i_13_3822, i_13_3868, i_13_3927, i_13_3975, i_13_3999, i_13_4080, i_13_4081, i_13_4252, i_13_4254, i_13_4255, i_13_4371, i_13_4449, i_13_4450, i_13_4602, o_13_58);
	kernel_13_59 k_13_59(i_13_33, i_13_61, i_13_192, i_13_195, i_13_205, i_13_253, i_13_260, i_13_282, i_13_309, i_13_310, i_13_375, i_13_382, i_13_463, i_13_466, i_13_578, i_13_589, i_13_617, i_13_618, i_13_619, i_13_624, i_13_625, i_13_672, i_13_673, i_13_760, i_13_768, i_13_816, i_13_942, i_13_976, i_13_979, i_13_1023, i_13_1081, i_13_1082, i_13_1087, i_13_1088, i_13_1096, i_13_1106, i_13_1147, i_13_1214, i_13_1270, i_13_1282, i_13_1309, i_13_1411, i_13_1514, i_13_1518, i_13_1561, i_13_1597, i_13_1680, i_13_1734, i_13_1741, i_13_1780, i_13_1849, i_13_1860, i_13_2002, i_13_2056, i_13_2191, i_13_2225, i_13_2383, i_13_2622, i_13_2769, i_13_2851, i_13_2878, i_13_2887, i_13_2907, i_13_2959, i_13_3028, i_13_3049, i_13_3113, i_13_3118, i_13_3156, i_13_3349, i_13_3352, i_13_3355, i_13_3382, i_13_3464, i_13_3534, i_13_3552, i_13_3571, i_13_3667, i_13_3730, i_13_3742, i_13_3984, i_13_3994, i_13_4063, i_13_4070, i_13_4108, i_13_4128, i_13_4155, i_13_4162, i_13_4165, i_13_4187, i_13_4299, i_13_4325, i_13_4335, i_13_4363, i_13_4369, i_13_4372, i_13_4418, i_13_4434, i_13_4532, i_13_4539, o_13_59);
	kernel_13_60 k_13_60(i_13_48, i_13_70, i_13_76, i_13_177, i_13_193, i_13_197, i_13_204, i_13_411, i_13_445, i_13_482, i_13_570, i_13_610, i_13_628, i_13_660, i_13_663, i_13_672, i_13_682, i_13_853, i_13_939, i_13_980, i_13_989, i_13_1084, i_13_1105, i_13_1224, i_13_1227, i_13_1228, i_13_1231, i_13_1232, i_13_1246, i_13_1275, i_13_1317, i_13_1385, i_13_1483, i_13_1515, i_13_1525, i_13_1626, i_13_1645, i_13_1677, i_13_1727, i_13_1732, i_13_1764, i_13_1767, i_13_1768, i_13_1830, i_13_1894, i_13_1914, i_13_1929, i_13_1933, i_13_1936, i_13_2022, i_13_2137, i_13_2199, i_13_2298, i_13_2301, i_13_2366, i_13_2473, i_13_2518, i_13_2707, i_13_2851, i_13_3031, i_13_3117, i_13_3135, i_13_3176, i_13_3264, i_13_3274, i_13_3354, i_13_3426, i_13_3483, i_13_3486, i_13_3489, i_13_3549, i_13_3576, i_13_3577, i_13_3651, i_13_3729, i_13_3730, i_13_3756, i_13_3785, i_13_3822, i_13_3869, i_13_3900, i_13_3901, i_13_3932, i_13_3981, i_13_3994, i_13_4017, i_13_4164, i_13_4297, i_13_4321, i_13_4324, i_13_4336, i_13_4368, i_13_4371, i_13_4372, i_13_4379, i_13_4435, i_13_4506, i_13_4540, i_13_4566, i_13_4606, o_13_60);
	kernel_13_61 k_13_61(i_13_91, i_13_92, i_13_94, i_13_175, i_13_176, i_13_186, i_13_231, i_13_238, i_13_256, i_13_308, i_13_316, i_13_317, i_13_375, i_13_381, i_13_382, i_13_558, i_13_572, i_13_582, i_13_604, i_13_605, i_13_607, i_13_609, i_13_613, i_13_641, i_13_644, i_13_658, i_13_659, i_13_668, i_13_689, i_13_743, i_13_758, i_13_829, i_13_986, i_13_1060, i_13_1100, i_13_1119, i_13_1226, i_13_1228, i_13_1273, i_13_1391, i_13_1398, i_13_1399, i_13_1408, i_13_1442, i_13_1518, i_13_1568, i_13_1595, i_13_1638, i_13_1639, i_13_1765, i_13_1805, i_13_1813, i_13_1828, i_13_1831, i_13_1840, i_13_1918, i_13_2012, i_13_2128, i_13_2173, i_13_2281, i_13_2423, i_13_2431, i_13_2677, i_13_2767, i_13_3047, i_13_3107, i_13_3164, i_13_3235, i_13_3241, i_13_3291, i_13_3416, i_13_3423, i_13_3426, i_13_3451, i_13_3547, i_13_3631, i_13_3686, i_13_3709, i_13_3754, i_13_3767, i_13_3817, i_13_3872, i_13_3893, i_13_3919, i_13_3928, i_13_3992, i_13_4164, i_13_4186, i_13_4273, i_13_4376, i_13_4396, i_13_4430, i_13_4487, i_13_4511, i_13_4523, i_13_4538, i_13_4566, i_13_4567, i_13_4568, i_13_4591, o_13_61);
	kernel_13_62 k_13_62(i_13_41, i_13_113, i_13_115, i_13_137, i_13_166, i_13_167, i_13_189, i_13_227, i_13_266, i_13_279, i_13_367, i_13_390, i_13_534, i_13_572, i_13_606, i_13_608, i_13_660, i_13_679, i_13_811, i_13_814, i_13_856, i_13_947, i_13_1084, i_13_1085, i_13_1094, i_13_1211, i_13_1217, i_13_1219, i_13_1352, i_13_1427, i_13_1462, i_13_1621, i_13_1622, i_13_1634, i_13_1640, i_13_1778, i_13_1788, i_13_1837, i_13_1838, i_13_1840, i_13_1841, i_13_1849, i_13_1939, i_13_1998, i_13_2021, i_13_2128, i_13_2135, i_13_2170, i_13_2172, i_13_2173, i_13_2209, i_13_2264, i_13_2404, i_13_2405, i_13_2407, i_13_2408, i_13_2421, i_13_2426, i_13_2432, i_13_2435, i_13_2448, i_13_2458, i_13_2495, i_13_2498, i_13_2564, i_13_2713, i_13_2714, i_13_2791, i_13_2846, i_13_2880, i_13_2907, i_13_2920, i_13_3044, i_13_3128, i_13_3141, i_13_3145, i_13_3146, i_13_3149, i_13_3407, i_13_3451, i_13_3452, i_13_3505, i_13_3509, i_13_3515, i_13_3529, i_13_3605, i_13_3613, i_13_3699, i_13_3737, i_13_3739, i_13_3763, i_13_3891, i_13_3892, i_13_4007, i_13_4160, i_13_4315, i_13_4325, i_13_4542, i_13_4555, i_13_4559, o_13_62);
	kernel_13_63 k_13_63(i_13_49, i_13_67, i_13_71, i_13_77, i_13_183, i_13_314, i_13_319, i_13_412, i_13_439, i_13_445, i_13_456, i_13_459, i_13_611, i_13_616, i_13_619, i_13_661, i_13_664, i_13_683, i_13_760, i_13_761, i_13_763, i_13_833, i_13_846, i_13_912, i_13_934, i_13_935, i_13_1096, i_13_1097, i_13_1102, i_13_1105, i_13_1132, i_13_1133, i_13_1155, i_13_1247, i_13_1258, i_13_1409, i_13_1483, i_13_1511, i_13_1525, i_13_1597, i_13_1645, i_13_1679, i_13_1733, i_13_1736, i_13_1754, i_13_1768, i_13_1771, i_13_1798, i_13_1799, i_13_1808, i_13_1885, i_13_1915, i_13_2023, i_13_2024, i_13_2029, i_13_2056, i_13_2149, i_13_2473, i_13_2474, i_13_2677, i_13_2708, i_13_2744, i_13_2857, i_13_2898, i_13_2902, i_13_2941, i_13_3031, i_13_3032, i_13_3077, i_13_3121, i_13_3231, i_13_3246, i_13_3265, i_13_3266, i_13_3346, i_13_3356, i_13_3397, i_13_3436, i_13_3461, i_13_3550, i_13_3551, i_13_3702, i_13_3739, i_13_3760, i_13_3784, i_13_3823, i_13_3847, i_13_3902, i_13_3911, i_13_3928, i_13_4085, i_13_4165, i_13_4245, i_13_4274, i_13_4325, i_13_4374, i_13_4397, i_13_4558, i_13_4606, i_13_4607, o_13_63);
	kernel_13_64 k_13_64(i_13_46, i_13_48, i_13_166, i_13_506, i_13_551, i_13_837, i_13_840, i_13_870, i_13_936, i_13_1058, i_13_1066, i_13_1119, i_13_1188, i_13_1189, i_13_1219, i_13_1245, i_13_1262, i_13_1323, i_13_1324, i_13_1326, i_13_1327, i_13_1405, i_13_1458, i_13_1512, i_13_1527, i_13_1628, i_13_1664, i_13_1777, i_13_1803, i_13_1805, i_13_1828, i_13_1831, i_13_1848, i_13_1849, i_13_1850, i_13_1855, i_13_1884, i_13_1885, i_13_1892, i_13_1896, i_13_2009, i_13_2043, i_13_2107, i_13_2145, i_13_2262, i_13_2299, i_13_2302, i_13_2351, i_13_2403, i_13_2469, i_13_2470, i_13_2472, i_13_2694, i_13_2697, i_13_2735, i_13_2740, i_13_2745, i_13_2980, i_13_2981, i_13_2982, i_13_2985, i_13_3028, i_13_3029, i_13_3055, i_13_3068, i_13_3105, i_13_3107, i_13_3108, i_13_3126, i_13_3211, i_13_3343, i_13_3503, i_13_3512, i_13_3523, i_13_3547, i_13_3548, i_13_3549, i_13_3604, i_13_3739, i_13_3763, i_13_3785, i_13_3816, i_13_3817, i_13_3820, i_13_3908, i_13_3930, i_13_4045, i_13_4059, i_13_4062, i_13_4063, i_13_4126, i_13_4162, i_13_4218, i_13_4315, i_13_4322, i_13_4376, i_13_4441, i_13_4497, i_13_4563, i_13_4567, o_13_64);
	kernel_13_65 k_13_65(i_13_137, i_13_164, i_13_166, i_13_167, i_13_169, i_13_172, i_13_229, i_13_263, i_13_266, i_13_281, i_13_380, i_13_460, i_13_530, i_13_607, i_13_640, i_13_676, i_13_688, i_13_794, i_13_811, i_13_814, i_13_815, i_13_821, i_13_823, i_13_824, i_13_913, i_13_961, i_13_982, i_13_1063, i_13_1064, i_13_1249, i_13_1324, i_13_1332, i_13_1495, i_13_1499, i_13_1502, i_13_1655, i_13_1846, i_13_1847, i_13_1849, i_13_1850, i_13_1852, i_13_1909, i_13_1958, i_13_1962, i_13_2107, i_13_2108, i_13_2116, i_13_2117, i_13_2134, i_13_2146, i_13_2227, i_13_2234, i_13_2247, i_13_2260, i_13_2261, i_13_2404, i_13_2405, i_13_2407, i_13_2408, i_13_2419, i_13_2449, i_13_2674, i_13_2678, i_13_2753, i_13_2848, i_13_2935, i_13_2936, i_13_3011, i_13_3148, i_13_3268, i_13_3374, i_13_3394, i_13_3438, i_13_3503, i_13_3505, i_13_3523, i_13_3595, i_13_3641, i_13_3739, i_13_3762, i_13_3817, i_13_3818, i_13_3862, i_13_3977, i_13_4015, i_13_4042, i_13_4060, i_13_4061, i_13_4063, i_13_4064, i_13_4123, i_13_4268, i_13_4303, i_13_4304, i_13_4315, i_13_4316, i_13_4319, i_13_4335, i_13_4405, i_13_4466, o_13_65);
	kernel_13_66 k_13_66(i_13_40, i_13_59, i_13_121, i_13_139, i_13_192, i_13_229, i_13_236, i_13_383, i_13_398, i_13_576, i_13_589, i_13_658, i_13_660, i_13_661, i_13_829, i_13_832, i_13_886, i_13_928, i_13_939, i_13_1000, i_13_1063, i_13_1098, i_13_1117, i_13_1118, i_13_1147, i_13_1225, i_13_1226, i_13_1227, i_13_1228, i_13_1244, i_13_1407, i_13_1408, i_13_1410, i_13_1479, i_13_1481, i_13_1513, i_13_1539, i_13_1552, i_13_1596, i_13_1652, i_13_1657, i_13_1675, i_13_1678, i_13_1733, i_13_1764, i_13_1765, i_13_1801, i_13_1802, i_13_1892, i_13_1927, i_13_1999, i_13_2002, i_13_2016, i_13_2296, i_13_2359, i_13_2443, i_13_2467, i_13_2569, i_13_2702, i_13_2705, i_13_2835, i_13_2857, i_13_2859, i_13_2874, i_13_2907, i_13_2980, i_13_2982, i_13_3017, i_13_3109, i_13_3133, i_13_3145, i_13_3371, i_13_3421, i_13_3475, i_13_3476, i_13_3486, i_13_3546, i_13_3547, i_13_3667, i_13_3730, i_13_3754, i_13_3757, i_13_3862, i_13_3979, i_13_3980, i_13_4086, i_13_4162, i_13_4186, i_13_4195, i_13_4295, i_13_4369, i_13_4393, i_13_4396, i_13_4428, i_13_4510, i_13_4511, i_13_4538, i_13_4599, i_13_4600, i_13_4603, o_13_66);
	kernel_13_67 k_13_67(i_13_64, i_13_90, i_13_91, i_13_139, i_13_174, i_13_175, i_13_204, i_13_228, i_13_229, i_13_282, i_13_283, i_13_284, i_13_336, i_13_337, i_13_341, i_13_393, i_13_414, i_13_417, i_13_450, i_13_522, i_13_535, i_13_567, i_13_657, i_13_661, i_13_733, i_13_796, i_13_823, i_13_824, i_13_846, i_13_847, i_13_849, i_13_850, i_13_981, i_13_985, i_13_1219, i_13_1224, i_13_1252, i_13_1263, i_13_1309, i_13_1312, i_13_1317, i_13_1462, i_13_1485, i_13_1549, i_13_1551, i_13_1552, i_13_1624, i_13_1644, i_13_1710, i_13_1803, i_13_1857, i_13_1858, i_13_1860, i_13_2197, i_13_2431, i_13_2452, i_13_2454, i_13_2517, i_13_2566, i_13_3006, i_13_3009, i_13_3012, i_13_3037, i_13_3061, i_13_3099, i_13_3100, i_13_3108, i_13_3168, i_13_3173, i_13_3217, i_13_3274, i_13_3343, i_13_3403, i_13_3456, i_13_3486, i_13_3487, i_13_3537, i_13_3540, i_13_3541, i_13_3574, i_13_3763, i_13_3799, i_13_3855, i_13_3856, i_13_3864, i_13_3867, i_13_3892, i_13_3937, i_13_4116, i_13_4200, i_13_4252, i_13_4254, i_13_4255, i_13_4257, i_13_4258, i_13_4260, i_13_4377, i_13_4378, i_13_4557, i_13_4560, o_13_67);
	kernel_13_68 k_13_68(i_13_28, i_13_48, i_13_63, i_13_64, i_13_73, i_13_142, i_13_144, i_13_226, i_13_279, i_13_282, i_13_307, i_13_315, i_13_316, i_13_405, i_13_532, i_13_550, i_13_604, i_13_639, i_13_651, i_13_666, i_13_667, i_13_675, i_13_676, i_13_688, i_13_757, i_13_868, i_13_875, i_13_931, i_13_940, i_13_947, i_13_1021, i_13_1099, i_13_1116, i_13_1207, i_13_1216, i_13_1278, i_13_1319, i_13_1467, i_13_1504, i_13_1522, i_13_1593, i_13_1594, i_13_1595, i_13_1602, i_13_1711, i_13_1839, i_13_1881, i_13_1990, i_13_2052, i_13_2053, i_13_2127, i_13_2169, i_13_2209, i_13_2260, i_13_2264, i_13_2277, i_13_2278, i_13_2380, i_13_2467, i_13_2470, i_13_2505, i_13_2578, i_13_2630, i_13_2674, i_13_2844, i_13_2845, i_13_2853, i_13_2908, i_13_2938, i_13_3001, i_13_3087, i_13_3096, i_13_3097, i_13_3108, i_13_3142, i_13_3260, i_13_3343, i_13_3349, i_13_3385, i_13_3501, i_13_3502, i_13_3525, i_13_3532, i_13_3646, i_13_3765, i_13_3767, i_13_3817, i_13_3888, i_13_3898, i_13_3907, i_13_3910, i_13_3925, i_13_4006, i_13_4033, i_13_4077, i_13_4107, i_13_4159, i_13_4186, i_13_4591, i_13_4600, o_13_68);
	kernel_13_69 k_13_69(i_13_48, i_13_52, i_13_75, i_13_158, i_13_182, i_13_213, i_13_214, i_13_277, i_13_286, i_13_383, i_13_526, i_13_577, i_13_578, i_13_582, i_13_599, i_13_618, i_13_619, i_13_661, i_13_697, i_13_715, i_13_792, i_13_937, i_13_949, i_13_1022, i_13_1076, i_13_1085, i_13_1141, i_13_1302, i_13_1304, i_13_1330, i_13_1362, i_13_1404, i_13_1492, i_13_1498, i_13_1500, i_13_1572, i_13_1623, i_13_1636, i_13_1807, i_13_1816, i_13_1817, i_13_2023, i_13_2107, i_13_2128, i_13_2141, i_13_2173, i_13_2284, i_13_2428, i_13_2440, i_13_2449, i_13_2452, i_13_2455, i_13_2459, i_13_2462, i_13_2668, i_13_2716, i_13_2753, i_13_2785, i_13_2787, i_13_2940, i_13_2958, i_13_3020, i_13_3105, i_13_3110, i_13_3143, i_13_3148, i_13_3231, i_13_3327, i_13_3428, i_13_3444, i_13_3454, i_13_3522, i_13_3523, i_13_3527, i_13_3553, i_13_3687, i_13_3688, i_13_3730, i_13_3733, i_13_3734, i_13_3757, i_13_3876, i_13_3911, i_13_4019, i_13_4020, i_13_4021, i_13_4047, i_13_4090, i_13_4093, i_13_4130, i_13_4254, i_13_4255, i_13_4270, i_13_4307, i_13_4416, i_13_4526, i_13_4539, i_13_4557, i_13_4559, i_13_4561, o_13_69);
	kernel_13_70 k_13_70(i_13_31, i_13_51, i_13_52, i_13_78, i_13_105, i_13_129, i_13_173, i_13_177, i_13_279, i_13_280, i_13_281, i_13_282, i_13_283, i_13_316, i_13_445, i_13_490, i_13_514, i_13_562, i_13_577, i_13_600, i_13_676, i_13_724, i_13_757, i_13_823, i_13_856, i_13_1018, i_13_1019, i_13_1022, i_13_1063, i_13_1082, i_13_1093, i_13_1143, i_13_1147, i_13_1526, i_13_1631, i_13_1634, i_13_1653, i_13_1654, i_13_1691, i_13_1786, i_13_1851, i_13_1940, i_13_2053, i_13_2055, i_13_2108, i_13_2116, i_13_2134, i_13_2198, i_13_2234, i_13_2236, i_13_2260, i_13_2335, i_13_2408, i_13_2443, i_13_2444, i_13_2506, i_13_2532, i_13_2543, i_13_2748, i_13_2752, i_13_3025, i_13_3093, i_13_3152, i_13_3165, i_13_3166, i_13_3175, i_13_3210, i_13_3262, i_13_3291, i_13_3461, i_13_3525, i_13_3539, i_13_3665, i_13_3727, i_13_3729, i_13_3731, i_13_3768, i_13_3817, i_13_3841, i_13_3854, i_13_3877, i_13_3889, i_13_3890, i_13_3910, i_13_3911, i_13_3971, i_13_3982, i_13_4015, i_13_4016, i_13_4063, i_13_4065, i_13_4216, i_13_4237, i_13_4258, i_13_4259, i_13_4297, i_13_4351, i_13_4375, i_13_4417, i_13_4524, o_13_70);
	kernel_13_71 k_13_71(i_13_51, i_13_52, i_13_107, i_13_111, i_13_117, i_13_277, i_13_340, i_13_418, i_13_511, i_13_561, i_13_565, i_13_618, i_13_628, i_13_651, i_13_745, i_13_835, i_13_855, i_13_915, i_13_1069, i_13_1083, i_13_1086, i_13_1120, i_13_1231, i_13_1335, i_13_1347, i_13_1363, i_13_1412, i_13_1467, i_13_1491, i_13_1492, i_13_1525, i_13_1572, i_13_1573, i_13_1623, i_13_1642, i_13_1654, i_13_1672, i_13_1785, i_13_1795, i_13_1806, i_13_1815, i_13_1906, i_13_1950, i_13_2008, i_13_2058, i_13_2059, i_13_2184, i_13_2283, i_13_2341, i_13_2353, i_13_2707, i_13_2712, i_13_2713, i_13_2715, i_13_2716, i_13_2787, i_13_2958, i_13_3010, i_13_3019, i_13_3063, i_13_3066, i_13_3099, i_13_3100, i_13_3156, i_13_3160, i_13_3165, i_13_3219, i_13_3220, i_13_3237, i_13_3238, i_13_3273, i_13_3291, i_13_3328, i_13_3346, i_13_3489, i_13_3525, i_13_3526, i_13_3540, i_13_3550, i_13_3552, i_13_3553, i_13_3598, i_13_3684, i_13_3687, i_13_3688, i_13_3922, i_13_4021, i_13_4047, i_13_4057, i_13_4065, i_13_4119, i_13_4120, i_13_4206, i_13_4216, i_13_4273, i_13_4387, i_13_4416, i_13_4452, i_13_4521, i_13_4560, o_13_71);
	kernel_13_72 k_13_72(i_13_68, i_13_134, i_13_138, i_13_283, i_13_358, i_13_359, i_13_363, i_13_400, i_13_472, i_13_529, i_13_661, i_13_662, i_13_664, i_13_665, i_13_745, i_13_827, i_13_835, i_13_842, i_13_854, i_13_887, i_13_943, i_13_949, i_13_959, i_13_1098, i_13_1123, i_13_1222, i_13_1229, i_13_1232, i_13_1259, i_13_1447, i_13_1501, i_13_1502, i_13_1508, i_13_1726, i_13_1745, i_13_1754, i_13_1951, i_13_1961, i_13_2002, i_13_2006, i_13_2020, i_13_2024, i_13_2033, i_13_2060, i_13_2104, i_13_2146, i_13_2181, i_13_2203, i_13_2240, i_13_2258, i_13_2284, i_13_2285, i_13_2344, i_13_2429, i_13_2447, i_13_2455, i_13_2515, i_13_2555, i_13_2696, i_13_2860, i_13_2885, i_13_2891, i_13_2920, i_13_3004, i_13_3013, i_13_3076, i_13_3172, i_13_3272, i_13_3404, i_13_3419, i_13_3490, i_13_3491, i_13_3580, i_13_3598, i_13_3599, i_13_3623, i_13_3757, i_13_3758, i_13_3787, i_13_3919, i_13_3959, i_13_3991, i_13_4122, i_13_4165, i_13_4166, i_13_4264, i_13_4265, i_13_4273, i_13_4333, i_13_4345, i_13_4382, i_13_4405, i_13_4433, i_13_4453, i_13_4454, i_13_4513, i_13_4571, i_13_4595, i_13_4597, i_13_4604, o_13_72);
	kernel_13_73 k_13_73(i_13_33, i_13_34, i_13_40, i_13_67, i_13_138, i_13_139, i_13_228, i_13_232, i_13_447, i_13_448, i_13_457, i_13_511, i_13_529, i_13_535, i_13_591, i_13_615, i_13_678, i_13_679, i_13_695, i_13_867, i_13_872, i_13_985, i_13_1110, i_13_1201, i_13_1301, i_13_1303, i_13_1348, i_13_1409, i_13_1435, i_13_1438, i_13_1447, i_13_1471, i_13_1714, i_13_1715, i_13_1717, i_13_1723, i_13_1725, i_13_1740, i_13_1783, i_13_1816, i_13_1832, i_13_1852, i_13_1888, i_13_1889, i_13_1928, i_13_1938, i_13_2044, i_13_2209, i_13_2228, i_13_2239, i_13_2361, i_13_2380, i_13_2427, i_13_2938, i_13_2949, i_13_2983, i_13_3001, i_13_3036, i_13_3039, i_13_3104, i_13_3109, i_13_3111, i_13_3112, i_13_3211, i_13_3217, i_13_3347, i_13_3388, i_13_3390, i_13_3391, i_13_3598, i_13_3612, i_13_3640, i_13_3683, i_13_3687, i_13_3703, i_13_3741, i_13_3746, i_13_3766, i_13_3793, i_13_3820, i_13_3836, i_13_3838, i_13_3847, i_13_3848, i_13_3984, i_13_4038, i_13_4054, i_13_4055, i_13_4110, i_13_4236, i_13_4237, i_13_4318, i_13_4352, i_13_4369, i_13_4397, i_13_4398, i_13_4399, i_13_4502, i_13_4536, i_13_4567, o_13_73);
	kernel_13_74 k_13_74(i_13_64, i_13_120, i_13_192, i_13_199, i_13_324, i_13_361, i_13_378, i_13_379, i_13_441, i_13_517, i_13_531, i_13_532, i_13_570, i_13_571, i_13_575, i_13_576, i_13_588, i_13_615, i_13_639, i_13_640, i_13_676, i_13_678, i_13_697, i_13_698, i_13_714, i_13_756, i_13_820, i_13_891, i_13_927, i_13_928, i_13_930, i_13_931, i_13_1063, i_13_1080, i_13_1098, i_13_1099, i_13_1101, i_13_1227, i_13_1257, i_13_1270, i_13_1407, i_13_1503, i_13_1504, i_13_1596, i_13_1597, i_13_1638, i_13_1719, i_13_1746, i_13_1747, i_13_1782, i_13_1792, i_13_1795, i_13_1800, i_13_1881, i_13_1989, i_13_1990, i_13_2011, i_13_2116, i_13_2118, i_13_2191, i_13_2259, i_13_2260, i_13_2358, i_13_2458, i_13_2466, i_13_2505, i_13_2609, i_13_2722, i_13_2848, i_13_2881, i_13_2901, i_13_2934, i_13_3000, i_13_3024, i_13_3027, i_13_3060, i_13_3114, i_13_3204, i_13_3259, i_13_3286, i_13_3420, i_13_3421, i_13_3448, i_13_3537, i_13_3753, i_13_3781, i_13_3790, i_13_3808, i_13_3811, i_13_3873, i_13_3924, i_13_3925, i_13_3928, i_13_3936, i_13_4008, i_13_4009, i_13_4077, i_13_4078, i_13_4086, i_13_4231, o_13_74);
	kernel_13_75 k_13_75(i_13_49, i_13_166, i_13_245, i_13_262, i_13_266, i_13_375, i_13_382, i_13_417, i_13_446, i_13_464, i_13_490, i_13_571, i_13_589, i_13_607, i_13_760, i_13_761, i_13_771, i_13_812, i_13_814, i_13_823, i_13_862, i_13_987, i_13_1066, i_13_1137, i_13_1147, i_13_1196, i_13_1228, i_13_1343, i_13_1489, i_13_1502, i_13_1558, i_13_1598, i_13_1760, i_13_1840, i_13_1841, i_13_1849, i_13_1853, i_13_1859, i_13_1931, i_13_1994, i_13_2137, i_13_2149, i_13_2179, i_13_2183, i_13_2192, i_13_2207, i_13_2263, i_13_2266, i_13_2346, i_13_2380, i_13_2396, i_13_2400, i_13_2408, i_13_2411, i_13_2469, i_13_2533, i_13_2696, i_13_2722, i_13_2749, i_13_2760, i_13_2769, i_13_2786, i_13_2857, i_13_2884, i_13_2938, i_13_2941, i_13_3028, i_13_3034, i_13_3047, i_13_3068, i_13_3218, i_13_3262, i_13_3316, i_13_3341, i_13_3343, i_13_3371, i_13_3394, i_13_3413, i_13_3442, i_13_3475, i_13_3506, i_13_3542, i_13_3630, i_13_3664, i_13_3667, i_13_3668, i_13_3750, i_13_3920, i_13_4009, i_13_4015, i_13_4061, i_13_4063, i_13_4162, i_13_4171, i_13_4315, i_13_4316, i_13_4317, i_13_4318, i_13_4369, i_13_4396, o_13_75);
	kernel_13_76 k_13_76(i_13_19, i_13_80, i_13_111, i_13_113, i_13_125, i_13_241, i_13_242, i_13_277, i_13_278, i_13_336, i_13_386, i_13_418, i_13_558, i_13_619, i_13_643, i_13_696, i_13_718, i_13_741, i_13_779, i_13_855, i_13_910, i_13_1017, i_13_1083, i_13_1084, i_13_1085, i_13_1087, i_13_1092, i_13_1381, i_13_1569, i_13_1620, i_13_1623, i_13_1624, i_13_1637, i_13_1642, i_13_1710, i_13_1774, i_13_1817, i_13_1840, i_13_1918, i_13_1952, i_13_1990, i_13_2174, i_13_2185, i_13_2348, i_13_2358, i_13_2433, i_13_2497, i_13_2548, i_13_2610, i_13_2712, i_13_2713, i_13_2716, i_13_2717, i_13_2739, i_13_2788, i_13_2921, i_13_2959, i_13_3047, i_13_3067, i_13_3097, i_13_3100, i_13_3101, i_13_3141, i_13_3145, i_13_3167, i_13_3221, i_13_3302, i_13_3312, i_13_3329, i_13_3374, i_13_3450, i_13_3454, i_13_3484, i_13_3486, i_13_3549, i_13_3553, i_13_3576, i_13_3684, i_13_3685, i_13_3688, i_13_3689, i_13_3736, i_13_3738, i_13_3878, i_13_3913, i_13_4022, i_13_4036, i_13_4050, i_13_4066, i_13_4081, i_13_4174, i_13_4269, i_13_4274, i_13_4328, i_13_4356, i_13_4363, i_13_4417, i_13_4522, i_13_4526, i_13_4536, o_13_76);
	kernel_13_77 k_13_77(i_13_43, i_13_49, i_13_80, i_13_115, i_13_196, i_13_265, i_13_277, i_13_278, i_13_310, i_13_352, i_13_377, i_13_405, i_13_454, i_13_476, i_13_520, i_13_562, i_13_563, i_13_578, i_13_582, i_13_661, i_13_664, i_13_665, i_13_673, i_13_741, i_13_823, i_13_833, i_13_850, i_13_935, i_13_1145, i_13_1327, i_13_1333, i_13_1364, i_13_1473, i_13_1508, i_13_1552, i_13_1627, i_13_1730, i_13_1732, i_13_1735, i_13_1754, i_13_1768, i_13_1841, i_13_1844, i_13_1864, i_13_2003, i_13_2018, i_13_2019, i_13_2020, i_13_2024, i_13_2098, i_13_2149, i_13_2265, i_13_2300, i_13_2452, i_13_2471, i_13_2519, i_13_2653, i_13_2708, i_13_2712, i_13_2743, i_13_2744, i_13_2898, i_13_2955, i_13_3007, i_13_3050, i_13_3100, i_13_3118, i_13_3234, i_13_3266, i_13_3316, i_13_3351, i_13_3418, i_13_3453, i_13_3464, i_13_3479, i_13_3553, i_13_3571, i_13_3604, i_13_3730, i_13_3757, i_13_3781, i_13_3799, i_13_3823, i_13_3904, i_13_3905, i_13_3972, i_13_4056, i_13_4122, i_13_4130, i_13_4162, i_13_4163, i_13_4165, i_13_4166, i_13_4237, i_13_4370, i_13_4432, i_13_4513, i_13_4517, i_13_4555, i_13_4607, o_13_77);
	kernel_13_78 k_13_78(i_13_39, i_13_49, i_13_79, i_13_285, i_13_327, i_13_340, i_13_528, i_13_530, i_13_672, i_13_673, i_13_717, i_13_797, i_13_825, i_13_862, i_13_894, i_13_1023, i_13_1024, i_13_1029, i_13_1258, i_13_1300, i_13_1320, i_13_1321, i_13_1383, i_13_1489, i_13_1500, i_13_1543, i_13_1552, i_13_1732, i_13_1743, i_13_1857, i_13_1884, i_13_1933, i_13_1947, i_13_1960, i_13_2014, i_13_2015, i_13_2032, i_13_2136, i_13_2139, i_13_2190, i_13_2204, i_13_2229, i_13_2460, i_13_2461, i_13_2463, i_13_2464, i_13_2595, i_13_2613, i_13_2652, i_13_2824, i_13_2874, i_13_2922, i_13_2923, i_13_2983, i_13_3174, i_13_3321, i_13_3322, i_13_3406, i_13_3417, i_13_3418, i_13_3432, i_13_3498, i_13_3522, i_13_3540, i_13_3541, i_13_3543, i_13_3550, i_13_3579, i_13_3613, i_13_3730, i_13_3731, i_13_3732, i_13_3733, i_13_3768, i_13_3769, i_13_3786, i_13_3787, i_13_3805, i_13_3831, i_13_3858, i_13_3912, i_13_3913, i_13_3931, i_13_3994, i_13_4117, i_13_4161, i_13_4188, i_13_4237, i_13_4255, i_13_4263, i_13_4296, i_13_4341, i_13_4380, i_13_4381, i_13_4414, i_13_4443, i_13_4567, i_13_4587, i_13_4597, i_13_4602, o_13_78);
	kernel_13_79 k_13_79(i_13_94, i_13_95, i_13_98, i_13_106, i_13_107, i_13_179, i_13_187, i_13_278, i_13_283, i_13_310, i_13_311, i_13_313, i_13_314, i_13_316, i_13_318, i_13_319, i_13_320, i_13_323, i_13_508, i_13_554, i_13_567, i_13_575, i_13_607, i_13_647, i_13_689, i_13_692, i_13_707, i_13_821, i_13_837, i_13_973, i_13_981, i_13_982, i_13_1024, i_13_1070, i_13_1101, i_13_1115, i_13_1123, i_13_1124, i_13_1184, i_13_1327, i_13_1394, i_13_1408, i_13_1471, i_13_1574, i_13_1609, i_13_1754, i_13_1773, i_13_1796, i_13_1859, i_13_1889, i_13_1931, i_13_1992, i_13_2123, i_13_2266, i_13_2267, i_13_2277, i_13_2403, i_13_2411, i_13_2494, i_13_2503, i_13_2545, i_13_2614, i_13_2680, i_13_2681, i_13_2699, i_13_2768, i_13_2824, i_13_2986, i_13_3065, i_13_3068, i_13_3130, i_13_3157, i_13_3167, i_13_3211, i_13_3212, i_13_3275, i_13_3339, i_13_3347, i_13_3392, i_13_3410, i_13_3416, i_13_3460, i_13_3544, i_13_3646, i_13_3685, i_13_3689, i_13_3799, i_13_3928, i_13_3931, i_13_4037, i_13_4080, i_13_4085, i_13_4270, i_13_4309, i_13_4342, i_13_4354, i_13_4369, i_13_4534, i_13_4570, i_13_4598, o_13_79);
	kernel_13_80 k_13_80(i_13_93, i_13_94, i_13_170, i_13_179, i_13_188, i_13_258, i_13_307, i_13_310, i_13_319, i_13_451, i_13_575, i_13_670, i_13_697, i_13_812, i_13_822, i_13_979, i_13_1020, i_13_1021, i_13_1023, i_13_1024, i_13_1077, i_13_1078, i_13_1138, i_13_1179, i_13_1219, i_13_1228, i_13_1273, i_13_1317, i_13_1318, i_13_1320, i_13_1429, i_13_1438, i_13_1608, i_13_1631, i_13_1633, i_13_1779, i_13_1780, i_13_1840, i_13_1853, i_13_1857, i_13_1920, i_13_2026, i_13_2136, i_13_2172, i_13_2200, i_13_2213, i_13_2245, i_13_2267, i_13_2399, i_13_2434, i_13_2454, i_13_2509, i_13_2571, i_13_2616, i_13_2617, i_13_2707, i_13_2749, i_13_2767, i_13_2787, i_13_2912, i_13_2983, i_13_3002, i_13_3094, i_13_3113, i_13_3171, i_13_3172, i_13_3209, i_13_3271, i_13_3326, i_13_3460, i_13_3463, i_13_3464, i_13_3534, i_13_3541, i_13_3544, i_13_3576, i_13_3664, i_13_3784, i_13_3821, i_13_3850, i_13_3855, i_13_3877, i_13_3894, i_13_3913, i_13_3927, i_13_4036, i_13_4067, i_13_4099, i_13_4178, i_13_4219, i_13_4255, i_13_4351, i_13_4353, i_13_4354, i_13_4381, i_13_4395, i_13_4431, i_13_4450, i_13_4556, i_13_4567, o_13_80);
	kernel_13_81 k_13_81(i_13_51, i_13_52, i_13_75, i_13_120, i_13_121, i_13_138, i_13_183, i_13_240, i_13_250, i_13_338, i_13_339, i_13_357, i_13_373, i_13_392, i_13_465, i_13_529, i_13_561, i_13_596, i_13_655, i_13_663, i_13_714, i_13_743, i_13_937, i_13_941, i_13_942, i_13_1077, i_13_1100, i_13_1211, i_13_1212, i_13_1397, i_13_1407, i_13_1408, i_13_1424, i_13_1469, i_13_1500, i_13_1501, i_13_1507, i_13_1523, i_13_1572, i_13_1608, i_13_1635, i_13_1636, i_13_1695, i_13_1722, i_13_1730, i_13_1775, i_13_1920, i_13_1951, i_13_1992, i_13_2031, i_13_2032, i_13_2058, i_13_2117, i_13_2169, i_13_2284, i_13_2343, i_13_2425, i_13_2455, i_13_2545, i_13_2724, i_13_2767, i_13_2787, i_13_2882, i_13_2923, i_13_2958, i_13_3061, i_13_3087, i_13_3088, i_13_3291, i_13_3372, i_13_3373, i_13_3417, i_13_3418, i_13_3427, i_13_3448, i_13_3463, i_13_3469, i_13_3489, i_13_3579, i_13_3597, i_13_3598, i_13_3633, i_13_3647, i_13_3649, i_13_3682, i_13_3687, i_13_3733, i_13_3767, i_13_3903, i_13_3990, i_13_4191, i_13_4249, i_13_4250, i_13_4263, i_13_4264, i_13_4412, i_13_4430, i_13_4452, i_13_4453, i_13_4541, o_13_81);
	kernel_13_82 k_13_82(i_13_40, i_13_46, i_13_76, i_13_172, i_13_264, i_13_279, i_13_282, i_13_283, i_13_337, i_13_378, i_13_525, i_13_693, i_13_697, i_13_1021, i_13_1066, i_13_1081, i_13_1082, i_13_1120, i_13_1224, i_13_1270, i_13_1306, i_13_1323, i_13_1401, i_13_1444, i_13_1495, i_13_1497, i_13_1498, i_13_1541, i_13_1566, i_13_1569, i_13_1633, i_13_1634, i_13_1783, i_13_1802, i_13_1916, i_13_1921, i_13_1927, i_13_1984, i_13_1990, i_13_1991, i_13_2001, i_13_2034, i_13_2037, i_13_2092, i_13_2117, i_13_2128, i_13_2177, i_13_2363, i_13_2424, i_13_2425, i_13_2430, i_13_2431, i_13_2449, i_13_2461, i_13_2548, i_13_2551, i_13_2601, i_13_2660, i_13_2674, i_13_2675, i_13_2934, i_13_2936, i_13_3004, i_13_3127, i_13_3142, i_13_3268, i_13_3269, i_13_3272, i_13_3393, i_13_3406, i_13_3421, i_13_3424, i_13_3582, i_13_3647, i_13_3727, i_13_3728, i_13_3730, i_13_3872, i_13_3987, i_13_4010, i_13_4014, i_13_4015, i_13_4016, i_13_4051, i_13_4087, i_13_4088, i_13_4120, i_13_4171, i_13_4224, i_13_4225, i_13_4249, i_13_4252, i_13_4261, i_13_4268, i_13_4297, i_13_4305, i_13_4393, i_13_4404, i_13_4475, i_13_4558, o_13_82);
	kernel_13_83 k_13_83(i_13_73, i_13_74, i_13_76, i_13_104, i_13_109, i_13_110, i_13_112, i_13_116, i_13_122, i_13_193, i_13_284, i_13_287, i_13_320, i_13_368, i_13_376, i_13_407, i_13_559, i_13_586, i_13_589, i_13_605, i_13_652, i_13_757, i_13_856, i_13_859, i_13_1021, i_13_1076, i_13_1086, i_13_1087, i_13_1217, i_13_1219, i_13_1273, i_13_1274, i_13_1474, i_13_1486, i_13_1567, i_13_1574, i_13_1630, i_13_1634, i_13_1678, i_13_1719, i_13_1775, i_13_1778, i_13_1837, i_13_1841, i_13_1849, i_13_1945, i_13_2137, i_13_2175, i_13_2192, i_13_2263, i_13_2423, i_13_2434, i_13_2435, i_13_2437, i_13_2438, i_13_2462, i_13_2465, i_13_2501, i_13_2535, i_13_2542, i_13_2716, i_13_2722, i_13_2920, i_13_3098, i_13_3101, i_13_3102, i_13_3143, i_13_3145, i_13_3146, i_13_3167, i_13_3290, i_13_3385, i_13_3452, i_13_3453, i_13_3478, i_13_3530, i_13_3532, i_13_3570, i_13_3578, i_13_3734, i_13_3764, i_13_3874, i_13_3938, i_13_4021, i_13_4036, i_13_4051, i_13_4093, i_13_4120, i_13_4121, i_13_4254, i_13_4255, i_13_4282, i_13_4283, i_13_4325, i_13_4366, i_13_4379, i_13_4524, i_13_4541, i_13_4559, i_13_4562, o_13_83);
	kernel_13_84 k_13_84(i_13_35, i_13_171, i_13_192, i_13_193, i_13_199, i_13_256, i_13_382, i_13_450, i_13_567, i_13_585, i_13_626, i_13_639, i_13_640, i_13_660, i_13_927, i_13_939, i_13_955, i_13_1062, i_13_1116, i_13_1121, i_13_1147, i_13_1192, i_13_1224, i_13_1225, i_13_1227, i_13_1228, i_13_1255, i_13_1314, i_13_1341, i_13_1407, i_13_1488, i_13_1494, i_13_1512, i_13_1521, i_13_1534, i_13_1552, i_13_1567, i_13_1570, i_13_1677, i_13_1724, i_13_1764, i_13_1765, i_13_1767, i_13_1801, i_13_1890, i_13_1891, i_13_1926, i_13_1956, i_13_1990, i_13_2044, i_13_2055, i_13_2056, i_13_2092, i_13_2240, i_13_2300, i_13_2568, i_13_2614, i_13_2646, i_13_2691, i_13_2781, i_13_2899, i_13_2934, i_13_2935, i_13_3006, i_13_3025, i_13_3118, i_13_3136, i_13_3144, i_13_3164, i_13_3214, i_13_3230, i_13_3267, i_13_3285, i_13_3286, i_13_3312, i_13_3339, i_13_3420, i_13_3421, i_13_3478, i_13_3531, i_13_3537, i_13_3901, i_13_3918, i_13_3978, i_13_3986, i_13_4009, i_13_4042, i_13_4077, i_13_4086, i_13_4087, i_13_4185, i_13_4248, i_13_4266, i_13_4267, i_13_4293, i_13_4302, i_13_4351, i_13_4368, i_13_4375, i_13_4468, o_13_84);
	kernel_13_85 k_13_85(i_13_67, i_13_282, i_13_285, i_13_384, i_13_385, i_13_448, i_13_456, i_13_625, i_13_669, i_13_745, i_13_796, i_13_816, i_13_852, i_13_865, i_13_889, i_13_948, i_13_1068, i_13_1101, i_13_1120, i_13_1259, i_13_1272, i_13_1273, i_13_1302, i_13_1303, i_13_1312, i_13_1390, i_13_1402, i_13_1484, i_13_1507, i_13_1573, i_13_1632, i_13_1642, i_13_1768, i_13_1777, i_13_1794, i_13_1795, i_13_1851, i_13_1933, i_13_1995, i_13_1996, i_13_2001, i_13_2014, i_13_2122, i_13_2211, i_13_2256, i_13_2266, i_13_2380, i_13_2427, i_13_2433, i_13_2434, i_13_2461, i_13_2463, i_13_2464, i_13_2470, i_13_2541, i_13_2754, i_13_2796, i_13_2884, i_13_2905, i_13_2916, i_13_2919, i_13_2940, i_13_2941, i_13_3021, i_13_3022, i_13_3039, i_13_3127, i_13_3273, i_13_3291, i_13_3307, i_13_3345, i_13_3399, i_13_3418, i_13_3427, i_13_3453, i_13_3454, i_13_3526, i_13_3534, i_13_3729, i_13_3730, i_13_3780, i_13_3788, i_13_3874, i_13_3927, i_13_3967, i_13_3990, i_13_4036, i_13_4065, i_13_4092, i_13_4189, i_13_4273, i_13_4297, i_13_4318, i_13_4341, i_13_4525, i_13_4560, i_13_4561, i_13_4567, i_13_4594, i_13_4603, o_13_85);
	kernel_13_86 k_13_86(i_13_51, i_13_52, i_13_66, i_13_75, i_13_76, i_13_110, i_13_111, i_13_119, i_13_123, i_13_182, i_13_183, i_13_250, i_13_277, i_13_451, i_13_507, i_13_528, i_13_554, i_13_559, i_13_561, i_13_562, i_13_563, i_13_605, i_13_618, i_13_655, i_13_679, i_13_697, i_13_699, i_13_730, i_13_942, i_13_1078, i_13_1081, i_13_1082, i_13_1084, i_13_1147, i_13_1210, i_13_1213, i_13_1284, i_13_1495, i_13_1573, i_13_1622, i_13_1645, i_13_1659, i_13_1660, i_13_1783, i_13_1784, i_13_1858, i_13_1920, i_13_1938, i_13_2002, i_13_2023, i_13_2170, i_13_2234, i_13_2320, i_13_2423, i_13_2436, i_13_2454, i_13_2455, i_13_2545, i_13_2616, i_13_2715, i_13_2752, i_13_2886, i_13_2887, i_13_2958, i_13_2959, i_13_3035, i_13_3062, i_13_3112, i_13_3129, i_13_3207, i_13_3214, i_13_3291, i_13_3372, i_13_3373, i_13_3390, i_13_3405, i_13_3417, i_13_3418, i_13_3454, i_13_3521, i_13_3526, i_13_3552, i_13_3571, i_13_3598, i_13_3649, i_13_3682, i_13_3687, i_13_3700, i_13_3769, i_13_3903, i_13_3904, i_13_3910, i_13_4332, i_13_4348, i_13_4349, i_13_4362, i_13_4371, i_13_4454, i_13_4538, i_13_4603, o_13_86);
	kernel_13_87 k_13_87(i_13_51, i_13_52, i_13_62, i_13_79, i_13_105, i_13_114, i_13_139, i_13_143, i_13_169, i_13_229, i_13_268, i_13_269, i_13_281, i_13_285, i_13_339, i_13_340, i_13_462, i_13_573, i_13_574, i_13_610, i_13_679, i_13_690, i_13_759, i_13_813, i_13_816, i_13_817, i_13_821, i_13_984, i_13_985, i_13_1142, i_13_1147, i_13_1274, i_13_1326, i_13_1476, i_13_1492, i_13_1599, i_13_1626, i_13_1749, i_13_1780, i_13_1807, i_13_1851, i_13_1852, i_13_1911, i_13_1950, i_13_2055, i_13_2058, i_13_2059, i_13_2110, i_13_2119, i_13_2139, i_13_2184, i_13_2283, i_13_2284, i_13_2409, i_13_2410, i_13_2579, i_13_2652, i_13_2696, i_13_2714, i_13_2752, i_13_2859, i_13_2879, i_13_2940, i_13_3049, i_13_3144, i_13_3211, i_13_3266, i_13_3291, i_13_3372, i_13_3373, i_13_3452, i_13_3480, i_13_3505, i_13_3535, i_13_3563, i_13_3646, i_13_3732, i_13_3820, i_13_3912, i_13_4018, i_13_4020, i_13_4045, i_13_4047, i_13_4062, i_13_4065, i_13_4066, i_13_4116, i_13_4117, i_13_4234, i_13_4262, i_13_4263, i_13_4296, i_13_4297, i_13_4309, i_13_4318, i_13_4380, i_13_4391, i_13_4453, i_13_4560, i_13_4564, o_13_87);
	kernel_13_88 k_13_88(i_13_35, i_13_66, i_13_130, i_13_133, i_13_177, i_13_236, i_13_253, i_13_357, i_13_444, i_13_455, i_13_465, i_13_466, i_13_528, i_13_582, i_13_606, i_13_720, i_13_744, i_13_915, i_13_1085, i_13_1276, i_13_1321, i_13_1329, i_13_1363, i_13_1396, i_13_1444, i_13_1446, i_13_1492, i_13_1500, i_13_1501, i_13_1507, i_13_1554, i_13_1555, i_13_1573, i_13_1604, i_13_1641, i_13_1644, i_13_1699, i_13_1700, i_13_1802, i_13_1848, i_13_1849, i_13_1929, i_13_2028, i_13_2032, i_13_2103, i_13_2143, i_13_2202, i_13_2203, i_13_2297, i_13_2346, i_13_2424, i_13_2425, i_13_2427, i_13_2468, i_13_2498, i_13_2499, i_13_2524, i_13_2559, i_13_2569, i_13_2720, i_13_2755, i_13_2767, i_13_2796, i_13_2887, i_13_2938, i_13_3027, i_13_3136, i_13_3232, i_13_3242, i_13_3243, i_13_3244, i_13_3470, i_13_3507, i_13_3541, i_13_3548, i_13_3596, i_13_3597, i_13_3613, i_13_3621, i_13_3633, i_13_3794, i_13_3840, i_13_3847, i_13_3849, i_13_3859, i_13_3994, i_13_4061, i_13_4063, i_13_4092, i_13_4125, i_13_4254, i_13_4265, i_13_4297, i_13_4315, i_13_4325, i_13_4398, i_13_4471, i_13_4512, i_13_4557, i_13_4603, o_13_88);
	kernel_13_89 k_13_89(i_13_95, i_13_121, i_13_139, i_13_140, i_13_335, i_13_362, i_13_370, i_13_380, i_13_461, i_13_586, i_13_587, i_13_659, i_13_685, i_13_812, i_13_856, i_13_1063, i_13_1064, i_13_1082, i_13_1090, i_13_1189, i_13_1217, i_13_1252, i_13_1273, i_13_1277, i_13_1298, i_13_1342, i_13_1343, i_13_1441, i_13_1468, i_13_1487, i_13_1568, i_13_1598, i_13_1678, i_13_1712, i_13_1778, i_13_1802, i_13_1811, i_13_1859, i_13_1928, i_13_1954, i_13_1958, i_13_1990, i_13_1994, i_13_2003, i_13_2053, i_13_2056, i_13_2189, i_13_2207, i_13_2260, i_13_2278, i_13_2279, i_13_2377, i_13_2404, i_13_2494, i_13_2548, i_13_2611, i_13_2612, i_13_2615, i_13_2633, i_13_2709, i_13_2710, i_13_2711, i_13_2746, i_13_2794, i_13_2855, i_13_2984, i_13_3110, i_13_3125, i_13_3136, i_13_3206, i_13_3217, i_13_3341, i_13_3367, i_13_3379, i_13_3385, i_13_3386, i_13_3407, i_13_3415, i_13_3416, i_13_3461, i_13_3476, i_13_3478, i_13_3532, i_13_3652, i_13_3664, i_13_3682, i_13_3703, i_13_3704, i_13_3818, i_13_3862, i_13_4051, i_13_4052, i_13_4097, i_13_4231, i_13_4268, i_13_4315, i_13_4393, i_13_4394, i_13_4405, i_13_4411, o_13_89);
	kernel_13_90 k_13_90(i_13_40, i_13_49, i_13_95, i_13_96, i_13_274, i_13_279, i_13_443, i_13_446, i_13_454, i_13_497, i_13_536, i_13_562, i_13_565, i_13_697, i_13_910, i_13_931, i_13_949, i_13_1067, i_13_1069, i_13_1214, i_13_1273, i_13_1391, i_13_1426, i_13_1480, i_13_1499, i_13_1532, i_13_1624, i_13_1636, i_13_1637, i_13_1642, i_13_1752, i_13_1783, i_13_1784, i_13_1840, i_13_1885, i_13_1932, i_13_2137, i_13_2170, i_13_2174, i_13_2209, i_13_2211, i_13_2233, i_13_2288, i_13_2434, i_13_2437, i_13_2438, i_13_2446, i_13_2486, i_13_2544, i_13_2545, i_13_2576, i_13_2650, i_13_2713, i_13_2716, i_13_2764, i_13_3020, i_13_3064, i_13_3091, i_13_3093, i_13_3109, i_13_3110, i_13_3143, i_13_3145, i_13_3164, i_13_3218, i_13_3271, i_13_3308, i_13_3371, i_13_3394, i_13_3424, i_13_3425, i_13_3692, i_13_3721, i_13_3750, i_13_3766, i_13_3767, i_13_3821, i_13_3856, i_13_3874, i_13_3875, i_13_3878, i_13_3905, i_13_4018, i_13_4019, i_13_4066, i_13_4087, i_13_4090, i_13_4091, i_13_4162, i_13_4205, i_13_4253, i_13_4271, i_13_4351, i_13_4352, i_13_4354, i_13_4361, i_13_4526, i_13_4561, i_13_4562, i_13_4567, o_13_90);
	kernel_13_91 k_13_91(i_13_51, i_13_52, i_13_53, i_13_94, i_13_106, i_13_125, i_13_149, i_13_166, i_13_168, i_13_169, i_13_188, i_13_241, i_13_251, i_13_261, i_13_264, i_13_340, i_13_370, i_13_374, i_13_418, i_13_459, i_13_531, i_13_574, i_13_619, i_13_620, i_13_679, i_13_680, i_13_772, i_13_842, i_13_889, i_13_895, i_13_952, i_13_976, i_13_980, i_13_1024, i_13_1048, i_13_1078, i_13_1079, i_13_1092, i_13_1142, i_13_1204, i_13_1255, i_13_1318, i_13_1465, i_13_1479, i_13_1502, i_13_1573, i_13_1574, i_13_1589, i_13_1609, i_13_1636, i_13_1637, i_13_1710, i_13_1749, i_13_1750, i_13_1751, i_13_1761, i_13_1808, i_13_1817, i_13_2033, i_13_2050, i_13_2411, i_13_2447, i_13_2722, i_13_2736, i_13_2752, i_13_2753, i_13_2788, i_13_2941, i_13_2942, i_13_2959, i_13_3220, i_13_3221, i_13_3373, i_13_3374, i_13_3418, i_13_3419, i_13_3423, i_13_3452, i_13_3550, i_13_3554, i_13_3559, i_13_3652, i_13_3653, i_13_3688, i_13_3719, i_13_3847, i_13_3965, i_13_3991, i_13_4000, i_13_4009, i_13_4021, i_13_4048, i_13_4066, i_13_4094, i_13_4318, i_13_4319, i_13_4364, i_13_4382, i_13_4391, i_13_4525, o_13_91);
	kernel_13_92 k_13_92(i_13_31, i_13_45, i_13_49, i_13_139, i_13_160, i_13_175, i_13_214, i_13_514, i_13_550, i_13_617, i_13_648, i_13_654, i_13_656, i_13_659, i_13_679, i_13_683, i_13_823, i_13_847, i_13_850, i_13_981, i_13_984, i_13_985, i_13_1115, i_13_1148, i_13_1326, i_13_1327, i_13_1331, i_13_1456, i_13_1516, i_13_1517, i_13_1519, i_13_1573, i_13_1660, i_13_1749, i_13_1807, i_13_1885, i_13_2021, i_13_2024, i_13_2059, i_13_2091, i_13_2097, i_13_2107, i_13_2185, i_13_2195, i_13_2230, i_13_2277, i_13_2469, i_13_2470, i_13_2473, i_13_2474, i_13_2519, i_13_2556, i_13_2642, i_13_2691, i_13_2699, i_13_2722, i_13_2749, i_13_2766, i_13_2889, i_13_3009, i_13_3031, i_13_3032, i_13_3037, i_13_3077, i_13_3112, i_13_3113, i_13_3138, i_13_3274, i_13_3378, i_13_3388, i_13_3474, i_13_3483, i_13_3522, i_13_3547, i_13_3558, i_13_3649, i_13_3662, i_13_3781, i_13_3819, i_13_3820, i_13_3823, i_13_3861, i_13_3973, i_13_3978, i_13_4055, i_13_4120, i_13_4123, i_13_4162, i_13_4165, i_13_4166, i_13_4365, i_13_4366, i_13_4370, i_13_4396, i_13_4557, i_13_4564, i_13_4567, i_13_4597, i_13_4600, i_13_4603, o_13_92);
	kernel_13_93 k_13_93(i_13_78, i_13_92, i_13_157, i_13_166, i_13_176, i_13_317, i_13_382, i_13_383, i_13_449, i_13_536, i_13_551, i_13_605, i_13_644, i_13_652, i_13_653, i_13_659, i_13_668, i_13_676, i_13_679, i_13_683, i_13_689, i_13_699, i_13_701, i_13_841, i_13_842, i_13_910, i_13_1106, i_13_1120, i_13_1121, i_13_1145, i_13_1207, i_13_1208, i_13_1310, i_13_1330, i_13_1423, i_13_1507, i_13_1516, i_13_1517, i_13_1570, i_13_1571, i_13_1664, i_13_1733, i_13_1742, i_13_1749, i_13_1924, i_13_1925, i_13_1937, i_13_2021, i_13_2054, i_13_2092, i_13_2208, i_13_2209, i_13_2318, i_13_2398, i_13_2468, i_13_2549, i_13_2552, i_13_2567, i_13_2582, i_13_2693, i_13_2699, i_13_3044, i_13_3077, i_13_3089, i_13_3101, i_13_3214, i_13_3217, i_13_3269, i_13_3532, i_13_3536, i_13_3559, i_13_3568, i_13_3569, i_13_3730, i_13_3731, i_13_3857, i_13_3863, i_13_3866, i_13_3874, i_13_3928, i_13_3991, i_13_3995, i_13_4033, i_13_4187, i_13_4190, i_13_4276, i_13_4280, i_13_4307, i_13_4335, i_13_4364, i_13_4435, i_13_4531, i_13_4565, i_13_4568, i_13_4585, i_13_4591, i_13_4592, i_13_4595, i_13_4600, i_13_4601, o_13_93);
	kernel_13_94 k_13_94(i_13_80, i_13_176, i_13_263, i_13_280, i_13_310, i_13_311, i_13_316, i_13_317, i_13_320, i_13_338, i_13_355, i_13_425, i_13_454, i_13_490, i_13_550, i_13_569, i_13_640, i_13_641, i_13_644, i_13_655, i_13_670, i_13_671, i_13_685, i_13_686, i_13_688, i_13_689, i_13_820, i_13_841, i_13_848, i_13_949, i_13_1072, i_13_1120, i_13_1121, i_13_1123, i_13_1136, i_13_1228, i_13_1273, i_13_1274, i_13_1276, i_13_1328, i_13_1361, i_13_1598, i_13_1661, i_13_1739, i_13_1786, i_13_1940, i_13_2027, i_13_2053, i_13_2054, i_13_2057, i_13_2173, i_13_2264, i_13_2345, i_13_2377, i_13_2398, i_13_2405, i_13_2453, i_13_2462, i_13_2507, i_13_2548, i_13_2549, i_13_2570, i_13_2579, i_13_2599, i_13_2651, i_13_2677, i_13_2693, i_13_2695, i_13_2696, i_13_2699, i_13_2747, i_13_3004, i_13_3008, i_13_3217, i_13_3340, i_13_3479, i_13_3538, i_13_3592, i_13_3721, i_13_3782, i_13_3862, i_13_3875, i_13_3893, i_13_3931, i_13_3982, i_13_3991, i_13_3992, i_13_3994, i_13_4019, i_13_4033, i_13_4186, i_13_4258, i_13_4259, i_13_4262, i_13_4375, i_13_4540, i_13_4565, i_13_4592, i_13_4595, i_13_4601, o_13_94);
	kernel_13_95 k_13_95(i_13_48, i_13_53, i_13_93, i_13_188, i_13_316, i_13_351, i_13_444, i_13_454, i_13_549, i_13_550, i_13_612, i_13_620, i_13_640, i_13_643, i_13_651, i_13_652, i_13_667, i_13_675, i_13_676, i_13_692, i_13_742, i_13_839, i_13_844, i_13_981, i_13_982, i_13_985, i_13_1117, i_13_1179, i_13_1181, i_13_1210, i_13_1498, i_13_1513, i_13_1515, i_13_1516, i_13_1519, i_13_1574, i_13_1641, i_13_1747, i_13_1792, i_13_1808, i_13_1810, i_13_1852, i_13_1853, i_13_1912, i_13_2003, i_13_2017, i_13_2050, i_13_2060, i_13_2169, i_13_2170, i_13_2243, i_13_2278, i_13_2348, i_13_2467, i_13_2511, i_13_2614, i_13_2674, i_13_2857, i_13_2935, i_13_2980, i_13_3208, i_13_3212, i_13_3214, i_13_3367, i_13_3369, i_13_3374, i_13_3401, i_13_3413, i_13_3416, i_13_3428, i_13_3491, i_13_3532, i_13_3541, i_13_3550, i_13_3554, i_13_3592, i_13_3645, i_13_3727, i_13_3730, i_13_3736, i_13_3765, i_13_3770, i_13_3862, i_13_3866, i_13_3888, i_13_3889, i_13_3890, i_13_3925, i_13_3987, i_13_3988, i_13_4049, i_13_4123, i_13_4265, i_13_4361, i_13_4544, i_13_4564, i_13_4566, i_13_4591, i_13_4599, i_13_4600, o_13_95);
	kernel_13_96 k_13_96(i_13_33, i_13_40, i_13_61, i_13_105, i_13_142, i_13_184, i_13_186, i_13_187, i_13_231, i_13_237, i_13_274, i_13_282, i_13_310, i_13_313, i_13_318, i_13_319, i_13_445, i_13_453, i_13_537, i_13_564, i_13_573, i_13_574, i_13_601, i_13_643, i_13_645, i_13_646, i_13_688, i_13_690, i_13_691, i_13_700, i_13_714, i_13_823, i_13_897, i_13_898, i_13_940, i_13_1069, i_13_1119, i_13_1123, i_13_1221, i_13_1275, i_13_1276, i_13_1383, i_13_1498, i_13_1635, i_13_1641, i_13_1642, i_13_1671, i_13_1716, i_13_1745, i_13_1852, i_13_1862, i_13_2047, i_13_2103, i_13_2140, i_13_2239, i_13_2299, i_13_2316, i_13_2321, i_13_2407, i_13_2509, i_13_2514, i_13_2635, i_13_2650, i_13_2652, i_13_2653, i_13_2679, i_13_2698, i_13_2722, i_13_2767, i_13_2770, i_13_2847, i_13_2848, i_13_2851, i_13_2984, i_13_3129, i_13_3210, i_13_3274, i_13_3292, i_13_3387, i_13_3390, i_13_3391, i_13_3408, i_13_3426, i_13_3460, i_13_3487, i_13_3606, i_13_3838, i_13_3892, i_13_3921, i_13_3927, i_13_3930, i_13_4018, i_13_4080, i_13_4084, i_13_4201, i_13_4344, i_13_4372, i_13_4570, i_13_4584, i_13_4597, o_13_96);
	kernel_13_97 k_13_97(i_13_52, i_13_103, i_13_106, i_13_107, i_13_158, i_13_166, i_13_233, i_13_287, i_13_310, i_13_337, i_13_454, i_13_470, i_13_537, i_13_553, i_13_584, i_13_607, i_13_608, i_13_646, i_13_647, i_13_679, i_13_688, i_13_691, i_13_692, i_13_843, i_13_844, i_13_1070, i_13_1086, i_13_1087, i_13_1106, i_13_1123, i_13_1131, i_13_1300, i_13_1331, i_13_1519, i_13_1554, i_13_1572, i_13_1573, i_13_1780, i_13_1804, i_13_1840, i_13_1915, i_13_1930, i_13_2024, i_13_2059, i_13_2060, i_13_2172, i_13_2173, i_13_2194, i_13_2284, i_13_2316, i_13_2380, i_13_2455, i_13_2624, i_13_2680, i_13_2698, i_13_2715, i_13_2798, i_13_2852, i_13_2902, i_13_2923, i_13_2938, i_13_3046, i_13_3066, i_13_3067, i_13_3103, i_13_3147, i_13_3148, i_13_3209, i_13_3289, i_13_3346, i_13_3383, i_13_3391, i_13_3392, i_13_3397, i_13_3446, i_13_3526, i_13_3530, i_13_3535, i_13_3544, i_13_3687, i_13_3742, i_13_3748, i_13_3865, i_13_3930, i_13_4020, i_13_4021, i_13_4048, i_13_4085, i_13_4119, i_13_4120, i_13_4121, i_13_4214, i_13_4308, i_13_4417, i_13_4450, i_13_4568, i_13_4570, i_13_4597, i_13_4598, i_13_4604, o_13_97);
	kernel_13_98 k_13_98(i_13_67, i_13_122, i_13_162, i_13_185, i_13_193, i_13_277, i_13_333, i_13_363, i_13_367, i_13_412, i_13_444, i_13_457, i_13_493, i_13_565, i_13_571, i_13_572, i_13_608, i_13_661, i_13_715, i_13_760, i_13_935, i_13_949, i_13_952, i_13_953, i_13_1210, i_13_1232, i_13_1267, i_13_1408, i_13_1443, i_13_1507, i_13_1625, i_13_1627, i_13_1628, i_13_1634, i_13_1637, i_13_1717, i_13_1736, i_13_1768, i_13_1771, i_13_1789, i_13_1790, i_13_1805, i_13_1808, i_13_1832, i_13_1912, i_13_1921, i_13_1940, i_13_2003, i_13_2012, i_13_2056, i_13_2123, i_13_2209, i_13_2240, i_13_2314, i_13_2426, i_13_2437, i_13_2533, i_13_2534, i_13_2538, i_13_2620, i_13_2987, i_13_3023, i_13_3032, i_13_3047, i_13_3104, i_13_3105, i_13_3166, i_13_3167, i_13_3231, i_13_3253, i_13_3265, i_13_3329, i_13_3397, i_13_3416, i_13_3420, i_13_3527, i_13_3550, i_13_3616, i_13_3681, i_13_3703, i_13_3847, i_13_3870, i_13_3874, i_13_3875, i_13_3878, i_13_3892, i_13_3982, i_13_3985, i_13_3986, i_13_4009, i_13_4198, i_13_4248, i_13_4311, i_13_4325, i_13_4327, i_13_4347, i_13_4351, i_13_4509, i_13_4514, i_13_4541, o_13_98);
	kernel_13_99 k_13_99(i_13_31, i_13_67, i_13_94, i_13_229, i_13_258, i_13_276, i_13_310, i_13_311, i_13_319, i_13_320, i_13_418, i_13_425, i_13_515, i_13_517, i_13_520, i_13_628, i_13_662, i_13_688, i_13_868, i_13_915, i_13_941, i_13_980, i_13_1021, i_13_1077, i_13_1202, i_13_1330, i_13_1331, i_13_1424, i_13_1444, i_13_1596, i_13_1598, i_13_1642, i_13_1663, i_13_1723, i_13_1734, i_13_1745, i_13_1824, i_13_1832, i_13_2008, i_13_2027, i_13_2132, i_13_2272, i_13_2317, i_13_2374, i_13_2450, i_13_2453, i_13_2497, i_13_2541, i_13_2542, i_13_2593, i_13_2666, i_13_2677, i_13_2740, i_13_2743, i_13_2744, i_13_2904, i_13_2915, i_13_2920, i_13_2968, i_13_3002, i_13_3121, i_13_3139, i_13_3176, i_13_3245, i_13_3312, i_13_3316, i_13_3414, i_13_3454, i_13_3455, i_13_3460, i_13_3463, i_13_3464, i_13_3479, i_13_3486, i_13_3488, i_13_3523, i_13_3569, i_13_3570, i_13_3571, i_13_3572, i_13_3577, i_13_3578, i_13_3593, i_13_3767, i_13_3831, i_13_3866, i_13_3942, i_13_4054, i_13_4094, i_13_4153, i_13_4164, i_13_4255, i_13_4256, i_13_4336, i_13_4352, i_13_4368, i_13_4372, i_13_4373, i_13_4517, i_13_4557, o_13_99);
	kernel_13_100 k_13_100(i_13_48, i_13_49, i_13_70, i_13_163, i_13_175, i_13_258, i_13_259, i_13_266, i_13_285, i_13_310, i_13_336, i_13_373, i_13_448, i_13_474, i_13_616, i_13_625, i_13_669, i_13_697, i_13_834, i_13_930, i_13_933, i_13_1071, i_13_1104, i_13_1105, i_13_1402, i_13_1648, i_13_1726, i_13_1735, i_13_1780, i_13_1797, i_13_1798, i_13_1804, i_13_1816, i_13_1818, i_13_1950, i_13_1995, i_13_1996, i_13_2004, i_13_2022, i_13_2148, i_13_2212, i_13_2356, i_13_2407, i_13_2409, i_13_2472, i_13_2473, i_13_2501, i_13_2617, i_13_2652, i_13_2673, i_13_2907, i_13_2915, i_13_2940, i_13_2941, i_13_2987, i_13_2997, i_13_3000, i_13_3030, i_13_3031, i_13_3127, i_13_3129, i_13_3130, i_13_3135, i_13_3217, i_13_3220, i_13_3265, i_13_3291, i_13_3312, i_13_3315, i_13_3376, i_13_3399, i_13_3417, i_13_3453, i_13_3639, i_13_3702, i_13_3741, i_13_3822, i_13_3834, i_13_3892, i_13_3940, i_13_3994, i_13_4045, i_13_4056, i_13_4057, i_13_4065, i_13_4083, i_13_4094, i_13_4153, i_13_4164, i_13_4188, i_13_4234, i_13_4251, i_13_4269, i_13_4273, i_13_4274, i_13_4324, i_13_4360, i_13_4526, i_13_4533, i_13_4606, o_13_100);
	kernel_13_101 k_13_101(i_13_51, i_13_52, i_13_105, i_13_106, i_13_312, i_13_381, i_13_508, i_13_537, i_13_552, i_13_553, i_13_655, i_13_679, i_13_691, i_13_817, i_13_843, i_13_983, i_13_984, i_13_985, i_13_1068, i_13_1069, i_13_1258, i_13_1300, i_13_1326, i_13_1329, i_13_1330, i_13_1345, i_13_1429, i_13_1492, i_13_1511, i_13_1516, i_13_1518, i_13_1519, i_13_1572, i_13_1573, i_13_1714, i_13_1778, i_13_1779, i_13_1803, i_13_1861, i_13_1885, i_13_1906, i_13_1911, i_13_1912, i_13_2002, i_13_2049, i_13_2059, i_13_2109, i_13_2175, i_13_2242, i_13_2243, i_13_2361, i_13_2409, i_13_2410, i_13_2464, i_13_2469, i_13_2470, i_13_2472, i_13_2533, i_13_2617, i_13_2693, i_13_2698, i_13_2725, i_13_2901, i_13_2919, i_13_2920, i_13_2982, i_13_2983, i_13_3030, i_13_3099, i_13_3111, i_13_3118, i_13_3130, i_13_3209, i_13_3346, i_13_3417, i_13_3418, i_13_3490, i_13_3525, i_13_3526, i_13_3535, i_13_3729, i_13_3769, i_13_3822, i_13_3864, i_13_3865, i_13_3891, i_13_3999, i_13_4038, i_13_4047, i_13_4048, i_13_4066, i_13_4119, i_13_4125, i_13_4126, i_13_4270, i_13_4323, i_13_4332, i_13_4353, i_13_4530, i_13_4569, o_13_101);
	kernel_13_102 k_13_102(i_13_48, i_13_79, i_13_251, i_13_277, i_13_310, i_13_319, i_13_340, i_13_409, i_13_597, i_13_643, i_13_664, i_13_745, i_13_760, i_13_1023, i_13_1024, i_13_1075, i_13_1096, i_13_1120, i_13_1140, i_13_1213, i_13_1266, i_13_1329, i_13_1403, i_13_1429, i_13_1430, i_13_1437, i_13_1482, i_13_1507, i_13_1573, i_13_1597, i_13_1626, i_13_1627, i_13_1634, i_13_1642, i_13_1686, i_13_1726, i_13_1780, i_13_1795, i_13_1844, i_13_2030, i_13_2106, i_13_2200, i_13_2272, i_13_2451, i_13_2454, i_13_2455, i_13_2541, i_13_2542, i_13_2545, i_13_2650, i_13_2708, i_13_2715, i_13_2716, i_13_2743, i_13_2770, i_13_2794, i_13_2904, i_13_2914, i_13_2919, i_13_2920, i_13_2921, i_13_3030, i_13_3105, i_13_3145, i_13_3244, i_13_3383, i_13_3388, i_13_3411, i_13_3412, i_13_3417, i_13_3418, i_13_3454, i_13_3463, i_13_3490, i_13_3535, i_13_3559, i_13_3568, i_13_3572, i_13_3574, i_13_3577, i_13_3688, i_13_3699, i_13_3877, i_13_3922, i_13_3928, i_13_3937, i_13_4036, i_13_4063, i_13_4255, i_13_4338, i_13_4352, i_13_4372, i_13_4373, i_13_4449, i_13_4522, i_13_4523, i_13_4525, i_13_4540, i_13_4558, i_13_4561, o_13_102);
	kernel_13_103 k_13_103(i_13_23, i_13_49, i_13_50, i_13_73, i_13_74, i_13_118, i_13_163, i_13_198, i_13_230, i_13_248, i_13_275, i_13_338, i_13_515, i_13_518, i_13_535, i_13_578, i_13_676, i_13_695, i_13_712, i_13_742, i_13_839, i_13_977, i_13_1082, i_13_1208, i_13_1210, i_13_1243, i_13_1262, i_13_1307, i_13_1397, i_13_1424, i_13_1505, i_13_1570, i_13_1658, i_13_1900, i_13_1918, i_13_1919, i_13_1928, i_13_1936, i_13_1954, i_13_1991, i_13_2030, i_13_2057, i_13_2173, i_13_2187, i_13_2261, i_13_2362, i_13_2395, i_13_2450, i_13_2452, i_13_2453, i_13_2512, i_13_2531, i_13_2549, i_13_2552, i_13_2576, i_13_2711, i_13_2741, i_13_2749, i_13_2764, i_13_2765, i_13_2785, i_13_2956, i_13_2963, i_13_3026, i_13_3061, i_13_3062, i_13_3128, i_13_3313, i_13_3370, i_13_3371, i_13_3376, i_13_3377, i_13_3415, i_13_3416, i_13_3475, i_13_3506, i_13_3533, i_13_3596, i_13_3613, i_13_3646, i_13_3647, i_13_3656, i_13_3671, i_13_3710, i_13_3719, i_13_3793, i_13_3872, i_13_3902, i_13_3920, i_13_4086, i_13_4123, i_13_4262, i_13_4331, i_13_4351, i_13_4367, i_13_4430, i_13_4450, i_13_4451, i_13_4557, i_13_4591, o_13_103);
	kernel_13_104 k_13_104(i_13_49, i_13_52, i_13_53, i_13_94, i_13_95, i_13_98, i_13_106, i_13_107, i_13_139, i_13_166, i_13_179, i_13_283, i_13_311, i_13_319, i_13_337, i_13_367, i_13_512, i_13_554, i_13_575, i_13_655, i_13_656, i_13_670, i_13_671, i_13_679, i_13_680, i_13_688, i_13_691, i_13_692, i_13_823, i_13_844, i_13_845, i_13_889, i_13_962, i_13_974, i_13_985, i_13_986, i_13_1052, i_13_1222, i_13_1331, i_13_1519, i_13_1520, i_13_1627, i_13_1636, i_13_1697, i_13_1789, i_13_1839, i_13_1861, i_13_1942, i_13_2032, i_13_2173, i_13_2182, i_13_2438, i_13_2618, i_13_2680, i_13_2725, i_13_2753, i_13_2905, i_13_2938, i_13_3002, i_13_3028, i_13_3112, i_13_3130, i_13_3155, i_13_3166, i_13_3167, i_13_3217, i_13_3218, i_13_3227, i_13_3280, i_13_3374, i_13_3418, i_13_3479, i_13_3505, i_13_3526, i_13_3536, i_13_3685, i_13_3719, i_13_3739, i_13_3769, i_13_3770, i_13_3865, i_13_3866, i_13_3892, i_13_3893, i_13_4021, i_13_4022, i_13_4049, i_13_4120, i_13_4121, i_13_4126, i_13_4127, i_13_4265, i_13_4270, i_13_4339, i_13_4340, i_13_4354, i_13_4534, i_13_4561, i_13_4570, i_13_4571, o_13_104);
	kernel_13_105 k_13_105(i_13_31, i_13_33, i_13_38, i_13_67, i_13_76, i_13_121, i_13_138, i_13_139, i_13_165, i_13_184, i_13_229, i_13_230, i_13_254, i_13_284, i_13_382, i_13_401, i_13_415, i_13_443, i_13_474, i_13_516, i_13_535, i_13_537, i_13_571, i_13_578, i_13_636, i_13_661, i_13_673, i_13_677, i_13_698, i_13_704, i_13_760, i_13_797, i_13_822, i_13_850, i_13_884, i_13_944, i_13_950, i_13_959, i_13_1042, i_13_1135, i_13_1218, i_13_1286, i_13_1339, i_13_1394, i_13_1472, i_13_1723, i_13_1725, i_13_1734, i_13_1794, i_13_1858, i_13_1943, i_13_1993, i_13_1994, i_13_1999, i_13_2000, i_13_2012, i_13_2060, i_13_2170, i_13_2407, i_13_2418, i_13_2434, i_13_2501, i_13_2509, i_13_2668, i_13_2679, i_13_2722, i_13_2749, i_13_2805, i_13_2858, i_13_2872, i_13_2897, i_13_3036, i_13_3064, i_13_3108, i_13_3109, i_13_3329, i_13_3374, i_13_3395, i_13_3444, i_13_3604, i_13_3622, i_13_3637, i_13_3651, i_13_3786, i_13_3794, i_13_3894, i_13_3974, i_13_3984, i_13_3988, i_13_4050, i_13_4064, i_13_4078, i_13_4094, i_13_4121, i_13_4195, i_13_4265, i_13_4336, i_13_4370, i_13_4454, i_13_4567, o_13_105);
	kernel_13_106 k_13_106(i_13_45, i_13_48, i_13_121, i_13_172, i_13_226, i_13_234, i_13_279, i_13_333, i_13_414, i_13_553, i_13_607, i_13_612, i_13_613, i_13_640, i_13_643, i_13_657, i_13_658, i_13_660, i_13_666, i_13_684, i_13_685, i_13_711, i_13_760, i_13_828, i_13_939, i_13_955, i_13_1071, i_13_1072, i_13_1116, i_13_1117, i_13_1225, i_13_1228, i_13_1232, i_13_1286, i_13_1390, i_13_1440, i_13_1493, i_13_1521, i_13_1522, i_13_1554, i_13_1638, i_13_1639, i_13_1696, i_13_1729, i_13_1736, i_13_1764, i_13_1792, i_13_1795, i_13_1801, i_13_1891, i_13_1926, i_13_1927, i_13_1944, i_13_2100, i_13_2115, i_13_2142, i_13_2211, i_13_2254, i_13_2299, i_13_2303, i_13_2313, i_13_2340, i_13_2376, i_13_2461, i_13_2595, i_13_2676, i_13_2677, i_13_2678, i_13_2721, i_13_2847, i_13_2848, i_13_2880, i_13_2881, i_13_3114, i_13_3261, i_13_3267, i_13_3367, i_13_3420, i_13_3421, i_13_3423, i_13_3546, i_13_3555, i_13_3564, i_13_3636, i_13_3753, i_13_3754, i_13_3892, i_13_3910, i_13_3924, i_13_4063, i_13_4186, i_13_4266, i_13_4280, i_13_4293, i_13_4294, i_13_4311, i_13_4467, i_13_4509, i_13_4593, i_13_4594, o_13_106);
	kernel_13_107 k_13_107(i_13_46, i_13_64, i_13_172, i_13_279, i_13_355, i_13_516, i_13_522, i_13_523, i_13_626, i_13_657, i_13_658, i_13_667, i_13_723, i_13_724, i_13_793, i_13_847, i_13_930, i_13_937, i_13_938, i_13_1017, i_13_1018, i_13_1071, i_13_1072, i_13_1093, i_13_1094, i_13_1099, i_13_1201, i_13_1225, i_13_1226, i_13_1279, i_13_1282, i_13_1315, i_13_1389, i_13_1423, i_13_1480, i_13_1486, i_13_1495, i_13_1523, i_13_1549, i_13_1630, i_13_1639, i_13_1792, i_13_1855, i_13_1884, i_13_1937, i_13_1955, i_13_2019, i_13_2020, i_13_2026, i_13_2127, i_13_2196, i_13_2197, i_13_2287, i_13_2317, i_13_2449, i_13_2452, i_13_2498, i_13_2539, i_13_2540, i_13_2592, i_13_2746, i_13_2917, i_13_2918, i_13_3029, i_13_3127, i_13_3241, i_13_3421, i_13_3422, i_13_3457, i_13_3458, i_13_3479, i_13_3483, i_13_3484, i_13_3485, i_13_3538, i_13_3574, i_13_3575, i_13_3595, i_13_3648, i_13_3738, i_13_3780, i_13_3781, i_13_3782, i_13_3820, i_13_3837, i_13_3918, i_13_4249, i_13_4250, i_13_4252, i_13_4257, i_13_4259, i_13_4321, i_13_4356, i_13_4366, i_13_4376, i_13_4446, i_13_4448, i_13_4450, i_13_4555, i_13_4604, o_13_107);
	kernel_13_108 k_13_108(i_13_25, i_13_34, i_13_156, i_13_160, i_13_224, i_13_228, i_13_231, i_13_273, i_13_278, i_13_328, i_13_382, i_13_411, i_13_417, i_13_534, i_13_565, i_13_603, i_13_604, i_13_665, i_13_688, i_13_732, i_13_741, i_13_933, i_13_945, i_13_946, i_13_1083, i_13_1084, i_13_1120, i_13_1218, i_13_1269, i_13_1344, i_13_1354, i_13_1443, i_13_1444, i_13_1473, i_13_1569, i_13_1605, i_13_1620, i_13_1687, i_13_1769, i_13_1836, i_13_1857, i_13_1957, i_13_2001, i_13_2047, i_13_2056, i_13_2150, i_13_2275, i_13_2280, i_13_2421, i_13_2424, i_13_2430, i_13_2497, i_13_2584, i_13_2712, i_13_2721, i_13_2722, i_13_2725, i_13_2784, i_13_2786, i_13_2856, i_13_2857, i_13_2859, i_13_2860, i_13_3010, i_13_3063, i_13_3064, i_13_3066, i_13_3097, i_13_3100, i_13_3103, i_13_3213, i_13_3234, i_13_3238, i_13_3255, i_13_3334, i_13_3428, i_13_3442, i_13_3487, i_13_3541, i_13_3554, i_13_3684, i_13_3691, i_13_3702, i_13_3717, i_13_3865, i_13_3871, i_13_3931, i_13_3977, i_13_4020, i_13_4252, i_13_4270, i_13_4328, i_13_4337, i_13_4350, i_13_4351, i_13_4395, i_13_4398, i_13_4413, i_13_4517, i_13_4593, o_13_108);
	kernel_13_109 k_13_109(i_13_118, i_13_127, i_13_181, i_13_182, i_13_260, i_13_280, i_13_281, i_13_283, i_13_325, i_13_355, i_13_535, i_13_569, i_13_596, i_13_598, i_13_599, i_13_667, i_13_697, i_13_712, i_13_728, i_13_742, i_13_745, i_13_778, i_13_821, i_13_847, i_13_853, i_13_856, i_13_863, i_13_898, i_13_946, i_13_986, i_13_1082, i_13_1094, i_13_1279, i_13_1280, i_13_1486, i_13_1487, i_13_1507, i_13_1669, i_13_1688, i_13_1724, i_13_1747, i_13_1751, i_13_1787, i_13_1808, i_13_1855, i_13_1856, i_13_1921, i_13_1940, i_13_1955, i_13_2056, i_13_2120, i_13_2146, i_13_2227, i_13_2305, i_13_2308, i_13_2314, i_13_2363, i_13_2425, i_13_2458, i_13_2459, i_13_2462, i_13_2467, i_13_2539, i_13_2540, i_13_2611, i_13_2612, i_13_2630, i_13_2765, i_13_2824, i_13_2882, i_13_2942, i_13_2981, i_13_3014, i_13_3020, i_13_3146, i_13_3148, i_13_3164, i_13_3169, i_13_3170, i_13_3173, i_13_3268, i_13_3290, i_13_3313, i_13_3370, i_13_3380, i_13_3425, i_13_3529, i_13_3782, i_13_3854, i_13_3871, i_13_3872, i_13_3875, i_13_3907, i_13_3908, i_13_3911, i_13_3941, i_13_4015, i_13_4261, i_13_4441, i_13_4519, o_13_109);
	kernel_13_110 k_13_110(i_13_31, i_13_34, i_13_35, i_13_39, i_13_64, i_13_67, i_13_122, i_13_134, i_13_161, i_13_225, i_13_232, i_13_233, i_13_272, i_13_306, i_13_386, i_13_449, i_13_490, i_13_493, i_13_538, i_13_607, i_13_612, i_13_648, i_13_746, i_13_759, i_13_762, i_13_763, i_13_764, i_13_868, i_13_1078, i_13_1128, i_13_1132, i_13_1186, i_13_1230, i_13_1303, i_13_1349, i_13_1444, i_13_1445, i_13_1447, i_13_1609, i_13_1700, i_13_1723, i_13_1724, i_13_1799, i_13_1817, i_13_1844, i_13_1912, i_13_1934, i_13_2142, i_13_2177, i_13_2194, i_13_2240, i_13_2318, i_13_2399, i_13_2430, i_13_2560, i_13_2681, i_13_2721, i_13_2722, i_13_2723, i_13_2726, i_13_2762, i_13_2825, i_13_2856, i_13_2860, i_13_2861, i_13_3002, i_13_3037, i_13_3130, i_13_3139, i_13_3213, i_13_3233, i_13_3366, i_13_3392, i_13_3415, i_13_3418, i_13_3438, i_13_3443, i_13_3618, i_13_3636, i_13_3637, i_13_3641, i_13_3650, i_13_3683, i_13_3686, i_13_3719, i_13_3725, i_13_3731, i_13_3843, i_13_3847, i_13_3848, i_13_3892, i_13_3991, i_13_4039, i_13_4040, i_13_4054, i_13_4237, i_13_4273, i_13_4347, i_13_4399, i_13_4400, o_13_110);
	kernel_13_111 k_13_111(i_13_38, i_13_103, i_13_112, i_13_185, i_13_280, i_13_281, i_13_284, i_13_320, i_13_338, i_13_373, i_13_376, i_13_454, i_13_533, i_13_571, i_13_590, i_13_596, i_13_598, i_13_599, i_13_641, i_13_677, i_13_685, i_13_686, i_13_715, i_13_761, i_13_814, i_13_815, i_13_820, i_13_821, i_13_832, i_13_896, i_13_1067, i_13_1076, i_13_1084, i_13_1129, i_13_1381, i_13_1438, i_13_1694, i_13_1714, i_13_1747, i_13_1748, i_13_1814, i_13_1856, i_13_1859, i_13_1909, i_13_1991, i_13_2138, i_13_2308, i_13_2366, i_13_2407, i_13_2458, i_13_2459, i_13_2461, i_13_2479, i_13_2506, i_13_2615, i_13_2633, i_13_2647, i_13_2650, i_13_2651, i_13_2722, i_13_2732, i_13_2749, i_13_2876, i_13_2938, i_13_2981, i_13_3142, i_13_3169, i_13_3206, i_13_3290, i_13_3376, i_13_3398, i_13_3415, i_13_3422, i_13_3524, i_13_3647, i_13_3692, i_13_3791, i_13_3844, i_13_3889, i_13_3890, i_13_3910, i_13_3911, i_13_3937, i_13_3989, i_13_3992, i_13_4015, i_13_4019, i_13_4036, i_13_4045, i_13_4052, i_13_4064, i_13_4078, i_13_4090, i_13_4097, i_13_4217, i_13_4259, i_13_4369, i_13_4559, i_13_4594, i_13_4603, o_13_111);
	kernel_13_112 k_13_112(i_13_3, i_13_37, i_13_180, i_13_181, i_13_183, i_13_185, i_13_187, i_13_193, i_13_210, i_13_244, i_13_255, i_13_360, i_13_382, i_13_446, i_13_526, i_13_550, i_13_596, i_13_597, i_13_625, i_13_640, i_13_642, i_13_643, i_13_646, i_13_647, i_13_685, i_13_692, i_13_851, i_13_894, i_13_898, i_13_975, i_13_1021, i_13_1093, i_13_1119, i_13_1120, i_13_1124, i_13_1276, i_13_1277, i_13_1391, i_13_1394, i_13_1407, i_13_1408, i_13_1461, i_13_1479, i_13_1488, i_13_1516, i_13_1643, i_13_1646, i_13_1668, i_13_1673, i_13_1813, i_13_1871, i_13_1990, i_13_2002, i_13_2046, i_13_2231, i_13_2361, i_13_2442, i_13_2542, i_13_2570, i_13_2676, i_13_2696, i_13_2767, i_13_2848, i_13_2852, i_13_2874, i_13_2920, i_13_2923, i_13_3092, i_13_3200, i_13_3291, i_13_3352, i_13_3419, i_13_3519, i_13_3523, i_13_3532, i_13_3541, i_13_3622, i_13_3730, i_13_3796, i_13_3900, i_13_3909, i_13_3918, i_13_3927, i_13_3928, i_13_3931, i_13_3993, i_13_3995, i_13_4083, i_13_4186, i_13_4189, i_13_4190, i_13_4192, i_13_4270, i_13_4297, i_13_4298, i_13_4341, i_13_4417, i_13_4596, i_13_4598, i_13_4599, o_13_112);
	kernel_13_113 k_13_113(i_13_26, i_13_52, i_13_167, i_13_170, i_13_248, i_13_263, i_13_278, i_13_320, i_13_340, i_13_376, i_13_452, i_13_454, i_13_460, i_13_607, i_13_732, i_13_811, i_13_815, i_13_1078, i_13_1079, i_13_1217, i_13_1304, i_13_1313, i_13_1343, i_13_1346, i_13_1402, i_13_1403, i_13_1408, i_13_1468, i_13_1529, i_13_1781, i_13_1805, i_13_1814, i_13_1835, i_13_1851, i_13_1852, i_13_1853, i_13_1912, i_13_1957, i_13_2006, i_13_2111, i_13_2128, i_13_2150, i_13_2174, i_13_2201, i_13_2234, i_13_2278, i_13_2279, i_13_2303, i_13_2318, i_13_2453, i_13_2618, i_13_2746, i_13_2765, i_13_2767, i_13_2788, i_13_2789, i_13_2848, i_13_2858, i_13_2872, i_13_3001, i_13_3002, i_13_3020, i_13_3091, i_13_3124, i_13_3131, i_13_3154, i_13_3215, i_13_3218, i_13_3232, i_13_3238, i_13_3305, i_13_3371, i_13_3442, i_13_3464, i_13_3505, i_13_3532, i_13_3545, i_13_3613, i_13_3616, i_13_3644, i_13_3689, i_13_3706, i_13_3712, i_13_3739, i_13_3892, i_13_3904, i_13_3961, i_13_4063, i_13_4231, i_13_4268, i_13_4271, i_13_4316, i_13_4367, i_13_4384, i_13_4393, i_13_4413, i_13_4450, i_13_4523, i_13_4532, i_13_4595, o_13_113);
	kernel_13_114 k_13_114(i_13_67, i_13_68, i_13_76, i_13_100, i_13_115, i_13_121, i_13_135, i_13_136, i_13_372, i_13_550, i_13_553, i_13_587, i_13_598, i_13_604, i_13_625, i_13_643, i_13_658, i_13_667, i_13_679, i_13_685, i_13_694, i_13_703, i_13_711, i_13_760, i_13_819, i_13_825, i_13_1116, i_13_1117, i_13_1153, i_13_1206, i_13_1207, i_13_1211, i_13_1273, i_13_1314, i_13_1390, i_13_1440, i_13_1507, i_13_1660, i_13_1668, i_13_1725, i_13_1729, i_13_1732, i_13_1735, i_13_1742, i_13_1774, i_13_1795, i_13_1796, i_13_1831, i_13_1944, i_13_1945, i_13_1999, i_13_2115, i_13_2201, i_13_2377, i_13_2380, i_13_2381, i_13_2422, i_13_2461, i_13_2548, i_13_2584, i_13_2646, i_13_2676, i_13_2718, i_13_2749, i_13_2847, i_13_2848, i_13_2881, i_13_2962, i_13_3090, i_13_3092, i_13_3094, i_13_3153, i_13_3352, i_13_3367, i_13_3414, i_13_3445, i_13_3637, i_13_3649, i_13_3865, i_13_3892, i_13_3893, i_13_3910, i_13_3927, i_13_3928, i_13_3990, i_13_4060, i_13_4063, i_13_4186, i_13_4192, i_13_4216, i_13_4293, i_13_4295, i_13_4297, i_13_4303, i_13_4305, i_13_4329, i_13_4432, i_13_4447, i_13_4558, i_13_4593, o_13_114);
	kernel_13_115 k_13_115(i_13_45, i_13_50, i_13_174, i_13_251, i_13_279, i_13_280, i_13_282, i_13_285, i_13_286, i_13_373, i_13_516, i_13_531, i_13_665, i_13_670, i_13_688, i_13_762, i_13_769, i_13_851, i_13_1020, i_13_1021, i_13_1024, i_13_1071, i_13_1272, i_13_1273, i_13_1425, i_13_1529, i_13_1601, i_13_1632, i_13_1633, i_13_1635, i_13_1636, i_13_1637, i_13_1693, i_13_1780, i_13_1932, i_13_2001, i_13_2034, i_13_2352, i_13_2380, i_13_2448, i_13_2449, i_13_2454, i_13_2455, i_13_2461, i_13_2464, i_13_2475, i_13_2545, i_13_2617, i_13_2641, i_13_2677, i_13_2762, i_13_2839, i_13_2844, i_13_2961, i_13_3105, i_13_3118, i_13_3129, i_13_3167, i_13_3198, i_13_3417, i_13_3421, i_13_3424, i_13_3447, i_13_3450, i_13_3460, i_13_3535, i_13_3612, i_13_3727, i_13_3729, i_13_3730, i_13_3731, i_13_3733, i_13_3793, i_13_3838, i_13_3909, i_13_3913, i_13_4014, i_13_4017, i_13_4018, i_13_4248, i_13_4251, i_13_4252, i_13_4253, i_13_4255, i_13_4256, i_13_4258, i_13_4260, i_13_4350, i_13_4407, i_13_4461, i_13_4513, i_13_4524, i_13_4554, i_13_4555, i_13_4557, i_13_4558, i_13_4560, i_13_4561, i_13_4562, i_13_4579, o_13_115);
	kernel_13_116 k_13_116(i_13_56, i_13_128, i_13_139, i_13_168, i_13_173, i_13_175, i_13_176, i_13_193, i_13_317, i_13_355, i_13_418, i_13_420, i_13_454, i_13_515, i_13_571, i_13_572, i_13_608, i_13_647, i_13_812, i_13_947, i_13_959, i_13_986, i_13_988, i_13_1216, i_13_1300, i_13_1345, i_13_1399, i_13_1405, i_13_1410, i_13_1453, i_13_1516, i_13_1552, i_13_1602, i_13_1714, i_13_1765, i_13_1767, i_13_1777, i_13_1793, i_13_1804, i_13_1828, i_13_1829, i_13_1831, i_13_1833, i_13_1885, i_13_2018, i_13_2019, i_13_2108, i_13_2146, i_13_2300, i_13_2335, i_13_2408, i_13_2470, i_13_2472, i_13_2474, i_13_2697, i_13_2705, i_13_2713, i_13_2746, i_13_2857, i_13_2858, i_13_2952, i_13_2980, i_13_2981, i_13_2982, i_13_2983, i_13_2985, i_13_3007, i_13_3027, i_13_3110, i_13_3154, i_13_3160, i_13_3211, i_13_3233, i_13_3386, i_13_3451, i_13_3549, i_13_3619, i_13_3710, i_13_3739, i_13_3763, i_13_3782, i_13_3817, i_13_3818, i_13_3872, i_13_4018, i_13_4054, i_13_4079, i_13_4084, i_13_4198, i_13_4258, i_13_4259, i_13_4376, i_13_4396, i_13_4511, i_13_4513, i_13_4522, i_13_4564, i_13_4565, i_13_4567, i_13_4570, o_13_116);
	kernel_13_117 k_13_117(i_13_70, i_13_71, i_13_80, i_13_260, i_13_262, i_13_377, i_13_386, i_13_448, i_13_449, i_13_464, i_13_523, i_13_527, i_13_592, i_13_674, i_13_687, i_13_701, i_13_763, i_13_845, i_13_887, i_13_935, i_13_979, i_13_1070, i_13_1214, i_13_1346, i_13_1402, i_13_1403, i_13_1430, i_13_1439, i_13_1492, i_13_1538, i_13_1600, i_13_1601, i_13_1645, i_13_1722, i_13_1727, i_13_1731, i_13_1733, i_13_1736, i_13_1781, i_13_1798, i_13_1799, i_13_1810, i_13_1889, i_13_1934, i_13_1948, i_13_1993, i_13_2001, i_13_2002, i_13_2020, i_13_2030, i_13_2059, i_13_2177, i_13_2194, i_13_2197, i_13_2285, i_13_2376, i_13_2381, i_13_2384, i_13_2507, i_13_2552, i_13_2680, i_13_2699, i_13_2723, i_13_2726, i_13_2744, i_13_2770, i_13_2771, i_13_2888, i_13_2916, i_13_2917, i_13_2973, i_13_3032, i_13_3064, i_13_3140, i_13_3262, i_13_3367, i_13_3371, i_13_3418, i_13_3438, i_13_3442, i_13_3536, i_13_3596, i_13_3639, i_13_3641, i_13_3684, i_13_3689, i_13_3780, i_13_3842, i_13_3896, i_13_3928, i_13_3994, i_13_3995, i_13_4058, i_13_4096, i_13_4392, i_13_4429, i_13_4451, i_13_4501, i_13_4598, i_13_4599, o_13_117);
	kernel_13_118 k_13_118(i_13_14, i_13_31, i_13_32, i_13_62, i_13_67, i_13_100, i_13_187, i_13_193, i_13_196, i_13_224, i_13_240, i_13_258, i_13_259, i_13_260, i_13_263, i_13_276, i_13_310, i_13_311, i_13_377, i_13_618, i_13_620, i_13_622, i_13_626, i_13_628, i_13_629, i_13_778, i_13_781, i_13_782, i_13_895, i_13_979, i_13_980, i_13_1077, i_13_1096, i_13_1112, i_13_1124, i_13_1140, i_13_1255, i_13_1256, i_13_1318, i_13_1391, i_13_1411, i_13_1469, i_13_1480, i_13_1483, i_13_1484, i_13_1558, i_13_1565, i_13_1643, i_13_1678, i_13_1688, i_13_1691, i_13_1745, i_13_1771, i_13_1805, i_13_1862, i_13_1991, i_13_2002, i_13_2120, i_13_2150, i_13_2291, i_13_2314, i_13_2365, i_13_2400, i_13_2425, i_13_2446, i_13_2447, i_13_2454, i_13_2677, i_13_2743, i_13_2857, i_13_2858, i_13_3005, i_13_3040, i_13_3131, i_13_3156, i_13_3292, i_13_3299, i_13_3356, i_13_3380, i_13_3383, i_13_3413, i_13_3419, i_13_3482, i_13_3523, i_13_3525, i_13_3526, i_13_3553, i_13_3554, i_13_3562, i_13_3570, i_13_3571, i_13_3642, i_13_4022, i_13_4254, i_13_4261, i_13_4364, i_13_4379, i_13_4391, i_13_4412, i_13_4508, o_13_118);
	kernel_13_119 k_13_119(i_13_76, i_13_249, i_13_258, i_13_324, i_13_372, i_13_531, i_13_576, i_13_580, i_13_595, i_13_670, i_13_699, i_13_714, i_13_718, i_13_719, i_13_777, i_13_781, i_13_811, i_13_838, i_13_843, i_13_891, i_13_942, i_13_1036, i_13_1092, i_13_1098, i_13_1116, i_13_1192, i_13_1321, i_13_1380, i_13_1461, i_13_1462, i_13_1479, i_13_1500, i_13_1664, i_13_1710, i_13_1743, i_13_1746, i_13_1756, i_13_1884, i_13_1887, i_13_1979, i_13_2140, i_13_2223, i_13_2224, i_13_2388, i_13_2404, i_13_2442, i_13_2452, i_13_2457, i_13_2499, i_13_2502, i_13_2565, i_13_2616, i_13_2633, i_13_2646, i_13_2667, i_13_2752, i_13_2820, i_13_2821, i_13_2824, i_13_3034, i_13_3046, i_13_3108, i_13_3171, i_13_3172, i_13_3216, i_13_3286, i_13_3289, i_13_3294, i_13_3306, i_13_3324, i_13_3372, i_13_3379, i_13_3433, i_13_3447, i_13_3462, i_13_3525, i_13_3559, i_13_3613, i_13_3639, i_13_3733, i_13_3790, i_13_3794, i_13_3798, i_13_3873, i_13_3913, i_13_3988, i_13_3992, i_13_4008, i_13_4212, i_13_4238, i_13_4377, i_13_4382, i_13_4387, i_13_4389, i_13_4410, i_13_4411, i_13_4440, i_13_4518, i_13_4557, i_13_4561, o_13_119);
	kernel_13_120 k_13_120(i_13_49, i_13_70, i_13_142, i_13_187, i_13_428, i_13_447, i_13_448, i_13_571, i_13_612, i_13_639, i_13_646, i_13_672, i_13_682, i_13_683, i_13_688, i_13_701, i_13_818, i_13_823, i_13_843, i_13_1105, i_13_1116, i_13_1123, i_13_1124, i_13_1269, i_13_1276, i_13_1277, i_13_1313, i_13_1374, i_13_1403, i_13_1474, i_13_1510, i_13_1511, i_13_1599, i_13_1600, i_13_1601, i_13_1638, i_13_1644, i_13_1645, i_13_1672, i_13_1726, i_13_1727, i_13_1736, i_13_1798, i_13_1925, i_13_1933, i_13_1996, i_13_2005, i_13_2052, i_13_2057, i_13_2107, i_13_2116, i_13_2133, i_13_2194, i_13_2266, i_13_2278, i_13_2403, i_13_2455, i_13_2456, i_13_2614, i_13_2679, i_13_2680, i_13_2697, i_13_2698, i_13_2699, i_13_2746, i_13_2887, i_13_2934, i_13_2940, i_13_3024, i_13_3113, i_13_3285, i_13_3393, i_13_3519, i_13_3595, i_13_3596, i_13_3652, i_13_3653, i_13_3733, i_13_3753, i_13_3797, i_13_3930, i_13_3940, i_13_3994, i_13_3995, i_13_4018, i_13_4019, i_13_4039, i_13_4085, i_13_4121, i_13_4252, i_13_4255, i_13_4262, i_13_4309, i_13_4310, i_13_4311, i_13_4318, i_13_4396, i_13_4559, i_13_4597, i_13_4598, o_13_120);
	kernel_13_121 k_13_121(i_13_1, i_13_31, i_13_36, i_13_37, i_13_76, i_13_99, i_13_163, i_13_165, i_13_167, i_13_168, i_13_183, i_13_184, i_13_217, i_13_336, i_13_372, i_13_526, i_13_532, i_13_570, i_13_676, i_13_686, i_13_714, i_13_718, i_13_813, i_13_814, i_13_1027, i_13_1067, i_13_1210, i_13_1272, i_13_1426, i_13_1495, i_13_1515, i_13_1525, i_13_1597, i_13_1677, i_13_1683, i_13_1731, i_13_1746, i_13_1747, i_13_1749, i_13_1756, i_13_1782, i_13_1801, i_13_1804, i_13_1805, i_13_1831, i_13_1832, i_13_1909, i_13_1911, i_13_2043, i_13_2046, i_13_2115, i_13_2116, i_13_2233, i_13_2263, i_13_2277, i_13_2407, i_13_2434, i_13_2476, i_13_2556, i_13_2722, i_13_2736, i_13_2748, i_13_2857, i_13_2889, i_13_2937, i_13_2980, i_13_3024, i_13_3027, i_13_3091, i_13_3126, i_13_3142, i_13_3196, i_13_3205, i_13_3216, i_13_3249, i_13_3289, i_13_3414, i_13_3444, i_13_3445, i_13_3472, i_13_3519, i_13_3549, i_13_3607, i_13_3661, i_13_3720, i_13_3739, i_13_3817, i_13_3918, i_13_3919, i_13_3988, i_13_4036, i_13_4044, i_13_4045, i_13_4059, i_13_4404, i_13_4413, i_13_4425, i_13_4497, i_13_4521, i_13_4593, o_13_121);
	kernel_13_122 k_13_122(i_13_40, i_13_50, i_13_112, i_13_115, i_13_121, i_13_192, i_13_251, i_13_274, i_13_277, i_13_415, i_13_457, i_13_561, i_13_562, i_13_607, i_13_616, i_13_688, i_13_928, i_13_951, i_13_952, i_13_1084, i_13_1085, i_13_1134, i_13_1141, i_13_1163, i_13_1273, i_13_1318, i_13_1444, i_13_1502, i_13_1573, i_13_1624, i_13_1633, i_13_1636, i_13_1642, i_13_1669, i_13_1678, i_13_1750, i_13_1839, i_13_1840, i_13_1858, i_13_1885, i_13_1930, i_13_2116, i_13_2175, i_13_2206, i_13_2233, i_13_2380, i_13_2433, i_13_2434, i_13_2435, i_13_2437, i_13_2438, i_13_2465, i_13_2505, i_13_2541, i_13_2590, i_13_2650, i_13_2716, i_13_2875, i_13_3004, i_13_3016, i_13_3047, i_13_3098, i_13_3101, i_13_3145, i_13_3146, i_13_3160, i_13_3162, i_13_3163, i_13_3166, i_13_3379, i_13_3455, i_13_3473, i_13_3527, i_13_3541, i_13_3604, i_13_3686, i_13_3688, i_13_3689, i_13_3784, i_13_3871, i_13_3872, i_13_3874, i_13_3904, i_13_3938, i_13_3991, i_13_4036, i_13_4057, i_13_4094, i_13_4158, i_13_4207, i_13_4253, i_13_4324, i_13_4350, i_13_4351, i_13_4352, i_13_4378, i_13_4379, i_13_4429, i_13_4468, i_13_4593, o_13_122);
	kernel_13_123 k_13_123(i_13_46, i_13_91, i_13_100, i_13_121, i_13_167, i_13_169, i_13_219, i_13_280, i_13_284, i_13_379, i_13_380, i_13_425, i_13_523, i_13_535, i_13_571, i_13_697, i_13_730, i_13_731, i_13_928, i_13_949, i_13_954, i_13_1063, i_13_1064, i_13_1093, i_13_1156, i_13_1297, i_13_1323, i_13_1324, i_13_1381, i_13_1441, i_13_1443, i_13_1471, i_13_1495, i_13_1525, i_13_1783, i_13_1800, i_13_1810, i_13_1828, i_13_1829, i_13_1846, i_13_1848, i_13_1849, i_13_1850, i_13_1928, i_13_2053, i_13_2107, i_13_2108, i_13_2116, i_13_2133, i_13_2134, i_13_2205, i_13_2232, i_13_2233, i_13_2234, i_13_2342, i_13_2404, i_13_2544, i_13_2746, i_13_2793, i_13_2848, i_13_2854, i_13_2872, i_13_2925, i_13_2935, i_13_3007, i_13_3053, i_13_3091, i_13_3108, i_13_3109, i_13_3110, i_13_3232, i_13_3242, i_13_3244, i_13_3306, i_13_3386, i_13_3394, i_13_3431, i_13_3612, i_13_3613, i_13_3739, i_13_3762, i_13_3765, i_13_3769, i_13_3817, i_13_3818, i_13_3820, i_13_3996, i_13_4015, i_13_4016, i_13_4042, i_13_4060, i_13_4061, i_13_4063, i_13_4064, i_13_4231, i_13_4249, i_13_4250, i_13_4267, i_13_4268, i_13_4567, o_13_123);
	kernel_13_124 k_13_124(i_13_63, i_13_64, i_13_73, i_13_130, i_13_139, i_13_175, i_13_191, i_13_283, i_13_354, i_13_355, i_13_356, i_13_357, i_13_450, i_13_468, i_13_469, i_13_470, i_13_485, i_13_507, i_13_668, i_13_694, i_13_831, i_13_883, i_13_946, i_13_947, i_13_1099, i_13_1208, i_13_1219, i_13_1337, i_13_1393, i_13_1395, i_13_1396, i_13_1517, i_13_1554, i_13_1696, i_13_1719, i_13_1721, i_13_1729, i_13_1730, i_13_1774, i_13_1777, i_13_1838, i_13_1846, i_13_1927, i_13_2143, i_13_2202, i_13_2230, i_13_2231, i_13_2366, i_13_2426, i_13_2430, i_13_2443, i_13_2444, i_13_2461, i_13_2466, i_13_2477, i_13_2511, i_13_2512, i_13_2538, i_13_2608, i_13_2692, i_13_2719, i_13_2755, i_13_2845, i_13_2881, i_13_2882, i_13_2920, i_13_2921, i_13_2938, i_13_3012, i_13_3087, i_13_3128, i_13_3133, i_13_3208, i_13_3370, i_13_3375, i_13_3532, i_13_3547, i_13_3595, i_13_3596, i_13_3619, i_13_3620, i_13_3632, i_13_3754, i_13_3781, i_13_3793, i_13_3924, i_13_3935, i_13_3982, i_13_3987, i_13_4162, i_13_4213, i_13_4214, i_13_4312, i_13_4329, i_13_4330, i_13_4331, i_13_4429, i_13_4450, i_13_4513, i_13_4540, o_13_124);
	kernel_13_125 k_13_125(i_13_52, i_13_71, i_13_80, i_13_140, i_13_232, i_13_323, i_13_419, i_13_448, i_13_521, i_13_526, i_13_539, i_13_557, i_13_629, i_13_646, i_13_647, i_13_681, i_13_683, i_13_698, i_13_718, i_13_745, i_13_814, i_13_823, i_13_827, i_13_871, i_13_872, i_13_985, i_13_1066, i_13_1075, i_13_1103, i_13_1133, i_13_1214, i_13_1219, i_13_1398, i_13_1430, i_13_1454, i_13_1510, i_13_1511, i_13_1529, i_13_1538, i_13_1664, i_13_1668, i_13_1673, i_13_1736, i_13_1750, i_13_1798, i_13_1799, i_13_1835, i_13_1889, i_13_1898, i_13_1912, i_13_1948, i_13_2046, i_13_2110, i_13_2181, i_13_2236, i_13_2555, i_13_2561, i_13_2680, i_13_2725, i_13_2726, i_13_2748, i_13_2851, i_13_2852, i_13_2884, i_13_2885, i_13_2938, i_13_3094, i_13_3243, i_13_3265, i_13_3381, i_13_3392, i_13_3541, i_13_3597, i_13_3742, i_13_3743, i_13_3759, i_13_3797, i_13_3821, i_13_3895, i_13_3896, i_13_3931, i_13_3994, i_13_4040, i_13_4063, i_13_4084, i_13_4190, i_13_4193, i_13_4219, i_13_4297, i_13_4298, i_13_4301, i_13_4325, i_13_4342, i_13_4377, i_13_4399, i_13_4400, i_13_4436, i_13_4597, i_13_4598, i_13_4607, o_13_125);
	kernel_13_126 k_13_126(i_13_34, i_13_121, i_13_126, i_13_191, i_13_205, i_13_231, i_13_324, i_13_416, i_13_493, i_13_494, i_13_529, i_13_534, i_13_538, i_13_576, i_13_602, i_13_715, i_13_728, i_13_782, i_13_832, i_13_841, i_13_930, i_13_1074, i_13_1096, i_13_1097, i_13_1204, i_13_1220, i_13_1304, i_13_1309, i_13_1474, i_13_1508, i_13_1627, i_13_1674, i_13_1723, i_13_1726, i_13_1727, i_13_1772, i_13_1784, i_13_1785, i_13_1786, i_13_1787, i_13_1790, i_13_1930, i_13_2056, i_13_2119, i_13_2123, i_13_2239, i_13_2248, i_13_2312, i_13_2340, i_13_2365, i_13_2461, i_13_2467, i_13_2501, i_13_2547, i_13_2646, i_13_2717, i_13_2898, i_13_2941, i_13_2942, i_13_3019, i_13_3023, i_13_3027, i_13_3034, i_13_3036, i_13_3104, i_13_3159, i_13_3160, i_13_3215, i_13_3254, i_13_3396, i_13_3409, i_13_3416, i_13_3506, i_13_3535, i_13_3616, i_13_3687, i_13_3703, i_13_3769, i_13_3794, i_13_3910, i_13_3951, i_13_3986, i_13_4008, i_13_4009, i_13_4036, i_13_4057, i_13_4063, i_13_4109, i_13_4193, i_13_4238, i_13_4261, i_13_4310, i_13_4328, i_13_4408, i_13_4416, i_13_4518, i_13_4519, i_13_4522, i_13_4523, i_13_4594, o_13_126);
	kernel_13_127 k_13_127(i_13_4, i_13_38, i_13_64, i_13_65, i_13_73, i_13_74, i_13_76, i_13_208, i_13_226, i_13_229, i_13_308, i_13_355, i_13_356, i_13_469, i_13_470, i_13_509, i_13_533, i_13_541, i_13_668, i_13_676, i_13_677, i_13_829, i_13_839, i_13_887, i_13_1100, i_13_1144, i_13_1145, i_13_1192, i_13_1246, i_13_1279, i_13_1307, i_13_1397, i_13_1400, i_13_1408, i_13_1445, i_13_1505, i_13_1621, i_13_1720, i_13_1721, i_13_1724, i_13_1730, i_13_1777, i_13_1778, i_13_1792, i_13_1909, i_13_1919, i_13_1928, i_13_2027, i_13_2056, i_13_2057, i_13_2237, i_13_2281, i_13_2282, i_13_2318, i_13_2354, i_13_2378, i_13_2468, i_13_2512, i_13_2534, i_13_2639, i_13_2656, i_13_2674, i_13_2692, i_13_2693, i_13_2720, i_13_2875, i_13_2882, i_13_2908, i_13_2974, i_13_3025, i_13_3034, i_13_3062, i_13_3136, i_13_3242, i_13_3251, i_13_3254, i_13_3371, i_13_3529, i_13_3532, i_13_3533, i_13_3593, i_13_3596, i_13_3619, i_13_3620, i_13_3631, i_13_3794, i_13_3935, i_13_3965, i_13_3988, i_13_3989, i_13_4034, i_13_4124, i_13_4187, i_13_4213, i_13_4214, i_13_4330, i_13_4331, i_13_4405, i_13_4430, i_13_4591, o_13_127);
	kernel_13_128 k_13_128(i_13_101, i_13_196, i_13_340, i_13_379, i_13_380, i_13_452, i_13_454, i_13_504, i_13_553, i_13_623, i_13_825, i_13_928, i_13_985, i_13_1063, i_13_1081, i_13_1082, i_13_1232, i_13_1297, i_13_1298, i_13_1320, i_13_1342, i_13_1410, i_13_1411, i_13_1412, i_13_1489, i_13_1491, i_13_1499, i_13_1502, i_13_1516, i_13_1517, i_13_1553, i_13_1554, i_13_1566, i_13_1627, i_13_1637, i_13_1801, i_13_1810, i_13_1926, i_13_1959, i_13_1990, i_13_2002, i_13_2107, i_13_2116, i_13_2134, i_13_2135, i_13_2201, i_13_2233, i_13_2234, i_13_2237, i_13_2294, i_13_2401, i_13_2461, i_13_2463, i_13_2515, i_13_2535, i_13_2572, i_13_2618, i_13_2934, i_13_2935, i_13_2936, i_13_2939, i_13_2977, i_13_3039, i_13_3172, i_13_3174, i_13_3218, i_13_3259, i_13_3285, i_13_3287, i_13_3339, i_13_3340, i_13_3341, i_13_3385, i_13_3421, i_13_3464, i_13_3521, i_13_3536, i_13_3579, i_13_3865, i_13_3877, i_13_3905, i_13_3912, i_13_4012, i_13_4013, i_13_4043, i_13_4051, i_13_4087, i_13_4162, i_13_4189, i_13_4266, i_13_4267, i_13_4271, i_13_4362, i_13_4393, i_13_4394, i_13_4396, i_13_4414, i_13_4443, i_13_4531, i_13_4594, o_13_128);
	kernel_13_129 k_13_129(i_13_116, i_13_121, i_13_122, i_13_139, i_13_173, i_13_175, i_13_226, i_13_229, i_13_280, i_13_281, i_13_311, i_13_319, i_13_337, i_13_373, i_13_416, i_13_523, i_13_526, i_13_563, i_13_590, i_13_658, i_13_733, i_13_847, i_13_848, i_13_850, i_13_851, i_13_938, i_13_986, i_13_1073, i_13_1201, i_13_1225, i_13_1280, i_13_1306, i_13_1345, i_13_1471, i_13_1549, i_13_1550, i_13_1712, i_13_1723, i_13_1751, i_13_1783, i_13_1855, i_13_1857, i_13_1858, i_13_1859, i_13_1901, i_13_1928, i_13_2125, i_13_2126, i_13_2169, i_13_2209, i_13_2238, i_13_2468, i_13_2510, i_13_2570, i_13_2692, i_13_2713, i_13_3001, i_13_3007, i_13_3008, i_13_3010, i_13_3037, i_13_3128, i_13_3133, i_13_3196, i_13_3217, i_13_3262, i_13_3269, i_13_3394, i_13_3412, i_13_3439, i_13_3442, i_13_3484, i_13_3485, i_13_3538, i_13_3539, i_13_3575, i_13_3685, i_13_3686, i_13_3820, i_13_3854, i_13_3862, i_13_3863, i_13_3868, i_13_3890, i_13_3908, i_13_4045, i_13_4106, i_13_4250, i_13_4253, i_13_4259, i_13_4276, i_13_4352, i_13_4369, i_13_4376, i_13_4379, i_13_4411, i_13_4522, i_13_4523, i_13_4531, i_13_4595, o_13_129);
	kernel_13_130 k_13_130(i_13_73, i_13_77, i_13_95, i_13_121, i_13_122, i_13_126, i_13_184, i_13_207, i_13_208, i_13_238, i_13_243, i_13_297, i_13_415, i_13_418, i_13_473, i_13_516, i_13_517, i_13_520, i_13_697, i_13_721, i_13_850, i_13_853, i_13_855, i_13_933, i_13_936, i_13_937, i_13_949, i_13_985, i_13_990, i_13_1071, i_13_1080, i_13_1128, i_13_1203, i_13_1209, i_13_1222, i_13_1252, i_13_1305, i_13_1317, i_13_1404, i_13_1521, i_13_1522, i_13_1548, i_13_1549, i_13_1552, i_13_1553, i_13_1602, i_13_1603, i_13_1699, i_13_1700, i_13_1711, i_13_1719, i_13_1723, i_13_1750, i_13_1786, i_13_1840, i_13_1843, i_13_1943, i_13_1957, i_13_1962, i_13_2033, i_13_2101, i_13_2113, i_13_2124, i_13_2125, i_13_2244, i_13_2248, i_13_2263, i_13_2333, i_13_2365, i_13_2442, i_13_2539, i_13_2581, i_13_2969, i_13_3007, i_13_3009, i_13_3040, i_13_3163, i_13_3268, i_13_3456, i_13_3461, i_13_3541, i_13_3577, i_13_3635, i_13_3739, i_13_3791, i_13_3796, i_13_3854, i_13_3898, i_13_3919, i_13_3921, i_13_3971, i_13_4078, i_13_4101, i_13_4261, i_13_4321, i_13_4334, i_13_4363, i_13_4380, i_13_4472, i_13_4509, o_13_130);
	kernel_13_131 k_13_131(i_13_37, i_13_91, i_13_92, i_13_94, i_13_95, i_13_112, i_13_230, i_13_238, i_13_256, i_13_260, i_13_263, i_13_274, i_13_277, i_13_315, i_13_316, i_13_326, i_13_364, i_13_374, i_13_518, i_13_607, i_13_670, i_13_694, i_13_697, i_13_698, i_13_778, i_13_832, i_13_943, i_13_976, i_13_977, i_13_979, i_13_1076, i_13_1082, i_13_1231, i_13_1262, i_13_1315, i_13_1336, i_13_1427, i_13_1433, i_13_1444, i_13_1468, i_13_1469, i_13_1512, i_13_1516, i_13_1669, i_13_1840, i_13_1861, i_13_1862, i_13_1886, i_13_1918, i_13_2140, i_13_2147, i_13_2198, i_13_2245, i_13_2298, i_13_2434, i_13_2521, i_13_2647, i_13_2651, i_13_2677, i_13_2702, i_13_2734, i_13_2735, i_13_2740, i_13_2899, i_13_2983, i_13_3143, i_13_3172, i_13_3208, i_13_3313, i_13_3341, i_13_3370, i_13_3373, i_13_3430, i_13_3448, i_13_3452, i_13_3593, i_13_3763, i_13_3806, i_13_3871, i_13_3907, i_13_4097, i_13_4118, i_13_4162, i_13_4177, i_13_4185, i_13_4278, i_13_4307, i_13_4351, i_13_4379, i_13_4387, i_13_4388, i_13_4390, i_13_4393, i_13_4441, i_13_4447, i_13_4448, i_13_4451, i_13_4518, i_13_4523, i_13_4567, o_13_131);
	kernel_13_132 k_13_132(i_13_46, i_13_78, i_13_103, i_13_154, i_13_245, i_13_379, i_13_411, i_13_421, i_13_443, i_13_450, i_13_451, i_13_460, i_13_461, i_13_552, i_13_658, i_13_661, i_13_698, i_13_820, i_13_897, i_13_940, i_13_1193, i_13_1251, i_13_1285, i_13_1297, i_13_1331, i_13_1342, i_13_1422, i_13_1432, i_13_1441, i_13_1442, i_13_1495, i_13_1567, i_13_1568, i_13_1601, i_13_1632, i_13_1633, i_13_1786, i_13_1801, i_13_1835, i_13_1858, i_13_1921, i_13_1928, i_13_1944, i_13_1945, i_13_1957, i_13_1959, i_13_2002, i_13_2098, i_13_2134, i_13_2135, i_13_2150, i_13_2197, i_13_2198, i_13_2278, i_13_2302, i_13_2316, i_13_2357, i_13_2380, i_13_2381, i_13_2405, i_13_2452, i_13_2544, i_13_2579, i_13_2614, i_13_2821, i_13_2983, i_13_2987, i_13_3010, i_13_3014, i_13_3017, i_13_3212, i_13_3268, i_13_3269, i_13_3341, i_13_3366, i_13_3375, i_13_3422, i_13_3485, i_13_3593, i_13_3727, i_13_3817, i_13_4015, i_13_4051, i_13_4086, i_13_4087, i_13_4208, i_13_4230, i_13_4231, i_13_4234, i_13_4249, i_13_4251, i_13_4252, i_13_4259, i_13_4261, i_13_4267, i_13_4268, i_13_4274, i_13_4393, i_13_4414, i_13_4447, o_13_132);
	kernel_13_133 k_13_133(i_13_25, i_13_168, i_13_229, i_13_318, i_13_463, i_13_517, i_13_523, i_13_526, i_13_535, i_13_538, i_13_571, i_13_601, i_13_717, i_13_759, i_13_850, i_13_895, i_13_1018, i_13_1120, i_13_1144, i_13_1210, i_13_1219, i_13_1273, i_13_1279, i_13_1426, i_13_1495, i_13_1497, i_13_1498, i_13_1528, i_13_1549, i_13_1606, i_13_1630, i_13_1631, i_13_1632, i_13_2001, i_13_2197, i_13_2198, i_13_2200, i_13_2365, i_13_2384, i_13_2457, i_13_2538, i_13_2541, i_13_2542, i_13_2764, i_13_2765, i_13_2767, i_13_2919, i_13_2935, i_13_3010, i_13_3037, i_13_3052, i_13_3100, i_13_3108, i_13_3119, i_13_3122, i_13_3141, i_13_3163, i_13_3169, i_13_3247, i_13_3262, i_13_3342, i_13_3459, i_13_3460, i_13_3540, i_13_3541, i_13_3612, i_13_3666, i_13_3722, i_13_3726, i_13_3727, i_13_3729, i_13_3730, i_13_3731, i_13_3838, i_13_3855, i_13_3859, i_13_3907, i_13_3916, i_13_3996, i_13_4014, i_13_4059, i_13_4060, i_13_4081, i_13_4162, i_13_4189, i_13_4207, i_13_4208, i_13_4251, i_13_4252, i_13_4255, i_13_4260, i_13_4266, i_13_4311, i_13_4341, i_13_4353, i_13_4465, i_13_4530, i_13_4555, i_13_4600, i_13_4603, o_13_133);
	kernel_13_134 k_13_134(i_13_65, i_13_94, i_13_95, i_13_173, i_13_175, i_13_176, i_13_202, i_13_235, i_13_307, i_13_308, i_13_442, i_13_443, i_13_485, i_13_572, i_13_604, i_13_605, i_13_658, i_13_662, i_13_667, i_13_668, i_13_676, i_13_677, i_13_698, i_13_934, i_13_946, i_13_1066, i_13_1217, i_13_1267, i_13_1306, i_13_1310, i_13_1388, i_13_1499, i_13_1504, i_13_1505, i_13_1561, i_13_1621, i_13_1630, i_13_1670, i_13_1720, i_13_1730, i_13_1802, i_13_1837, i_13_1838, i_13_1840, i_13_1841, i_13_1904, i_13_2170, i_13_2173, i_13_2230, i_13_2422, i_13_2423, i_13_2424, i_13_2425, i_13_2426, i_13_2431, i_13_2432, i_13_2435, i_13_2503, i_13_2593, i_13_2674, i_13_2675, i_13_2677, i_13_2678, i_13_2702, i_13_2912, i_13_2950, i_13_2951, i_13_3142, i_13_3143, i_13_3145, i_13_3242, i_13_3260, i_13_3269, i_13_3304, i_13_3305, i_13_3421, i_13_3422, i_13_3424, i_13_3425, i_13_3446, i_13_3529, i_13_3592, i_13_3726, i_13_3871, i_13_4016, i_13_4018, i_13_4019, i_13_4078, i_13_4079, i_13_4249, i_13_4253, i_13_4258, i_13_4351, i_13_4430, i_13_4447, i_13_4541, i_13_4555, i_13_4556, i_13_4559, i_13_4591, o_13_134);
	kernel_13_135 k_13_135(i_13_90, i_13_91, i_13_94, i_13_117, i_13_118, i_13_165, i_13_168, i_13_180, i_13_181, i_13_183, i_13_201, i_13_306, i_13_561, i_13_567, i_13_685, i_13_694, i_13_697, i_13_729, i_13_732, i_13_822, i_13_855, i_13_945, i_13_949, i_13_1065, i_13_1075, i_13_1251, i_13_1263, i_13_1297, i_13_1341, i_13_1344, i_13_1363, i_13_1404, i_13_1405, i_13_1440, i_13_1485, i_13_1515, i_13_1620, i_13_1624, i_13_1629, i_13_1633, i_13_1828, i_13_1836, i_13_1885, i_13_1888, i_13_1917, i_13_1921, i_13_1936, i_13_2004, i_13_2107, i_13_2170, i_13_2172, i_13_2205, i_13_2208, i_13_2233, i_13_2421, i_13_2424, i_13_2433, i_13_2452, i_13_2467, i_13_2614, i_13_2676, i_13_2725, i_13_2910, i_13_3019, i_13_3034, i_13_3063, i_13_3099, i_13_3106, i_13_3108, i_13_3126, i_13_3144, i_13_3162, i_13_3163, i_13_3172, i_13_3207, i_13_3208, i_13_3213, i_13_3240, i_13_3396, i_13_3414, i_13_3415, i_13_3486, i_13_3699, i_13_3717, i_13_3762, i_13_3783, i_13_3834, i_13_3843, i_13_3870, i_13_3871, i_13_4005, i_13_4006, i_13_4044, i_13_4117, i_13_4350, i_13_4374, i_13_4401, i_13_4440, i_13_4452, i_13_4564, o_13_135);
	kernel_13_136 k_13_136(i_13_49, i_13_73, i_13_76, i_13_157, i_13_228, i_13_229, i_13_282, i_13_283, i_13_515, i_13_517, i_13_535, i_13_657, i_13_659, i_13_660, i_13_724, i_13_821, i_13_850, i_13_1017, i_13_1019, i_13_1053, i_13_1074, i_13_1075, i_13_1286, i_13_1422, i_13_1425, i_13_1426, i_13_1570, i_13_1632, i_13_1633, i_13_1634, i_13_1635, i_13_1773, i_13_1786, i_13_1795, i_13_1841, i_13_2026, i_13_2029, i_13_2209, i_13_2236, i_13_2396, i_13_2426, i_13_2448, i_13_2449, i_13_2451, i_13_2452, i_13_2453, i_13_2454, i_13_2707, i_13_2722, i_13_3009, i_13_3010, i_13_3037, i_13_3269, i_13_3388, i_13_3450, i_13_3459, i_13_3460, i_13_3467, i_13_3484, i_13_3551, i_13_3567, i_13_3568, i_13_3573, i_13_3576, i_13_3577, i_13_3636, i_13_3645, i_13_3646, i_13_3647, i_13_3648, i_13_3684, i_13_3702, i_13_3729, i_13_3730, i_13_3838, i_13_3852, i_13_3862, i_13_3889, i_13_3890, i_13_3893, i_13_3988, i_13_4015, i_13_4017, i_13_4018, i_13_4079, i_13_4189, i_13_4251, i_13_4252, i_13_4253, i_13_4261, i_13_4262, i_13_4305, i_13_4358, i_13_4361, i_13_4513, i_13_4556, i_13_4557, i_13_4558, i_13_4559, i_13_4591, o_13_136);
	kernel_13_137 k_13_137(i_13_31, i_13_48, i_13_55, i_13_75, i_13_139, i_13_205, i_13_210, i_13_214, i_13_228, i_13_229, i_13_230, i_13_379, i_13_422, i_13_514, i_13_517, i_13_520, i_13_572, i_13_625, i_13_659, i_13_705, i_13_710, i_13_813, i_13_848, i_13_850, i_13_856, i_13_865, i_13_949, i_13_981, i_13_985, i_13_1018, i_13_1200, i_13_1219, i_13_1300, i_13_1327, i_13_1334, i_13_1438, i_13_1569, i_13_1570, i_13_1630, i_13_1678, i_13_1682, i_13_1831, i_13_1840, i_13_1853, i_13_1861, i_13_1908, i_13_1909, i_13_1923, i_13_2027, i_13_2107, i_13_2197, i_13_2239, i_13_2406, i_13_2407, i_13_2452, i_13_2455, i_13_2698, i_13_2699, i_13_2721, i_13_2722, i_13_2753, i_13_2794, i_13_2942, i_13_3010, i_13_3011, i_13_3014, i_13_3027, i_13_3037, i_13_3109, i_13_3288, i_13_3397, i_13_3403, i_13_3464, i_13_3488, i_13_3526, i_13_3546, i_13_3646, i_13_3763, i_13_3764, i_13_3788, i_13_3864, i_13_3865, i_13_3888, i_13_3907, i_13_3910, i_13_3914, i_13_4009, i_13_4018, i_13_4022, i_13_4157, i_13_4249, i_13_4252, i_13_4255, i_13_4265, i_13_4382, i_13_4432, i_13_4557, i_13_4561, i_13_4562, i_13_4589, o_13_137);
	kernel_13_138 k_13_138(i_13_40, i_13_76, i_13_121, i_13_122, i_13_226, i_13_372, i_13_442, i_13_456, i_13_490, i_13_517, i_13_531, i_13_532, i_13_533, i_13_572, i_13_715, i_13_722, i_13_930, i_13_948, i_13_951, i_13_1099, i_13_1100, i_13_1280, i_13_1303, i_13_1327, i_13_1408, i_13_1426, i_13_1433, i_13_1446, i_13_1468, i_13_1623, i_13_1666, i_13_1720, i_13_1723, i_13_1758, i_13_1783, i_13_1785, i_13_1786, i_13_1787, i_13_1837, i_13_1904, i_13_1940, i_13_2014, i_13_2103, i_13_2207, i_13_2209, i_13_2225, i_13_2236, i_13_2238, i_13_2242, i_13_2243, i_13_2343, i_13_2358, i_13_2425, i_13_2428, i_13_2533, i_13_2677, i_13_2695, i_13_2845, i_13_3018, i_13_3037, i_13_3038, i_13_3163, i_13_3164, i_13_3217, i_13_3218, i_13_3219, i_13_3259, i_13_3281, i_13_3286, i_13_3287, i_13_3322, i_13_3422, i_13_3426, i_13_3649, i_13_3739, i_13_3754, i_13_3791, i_13_3873, i_13_3874, i_13_3875, i_13_3876, i_13_3919, i_13_3925, i_13_3984, i_13_3985, i_13_3998, i_13_4009, i_13_4010, i_13_4051, i_13_4078, i_13_4079, i_13_4106, i_13_4162, i_13_4213, i_13_4261, i_13_4519, i_13_4524, i_13_4531, i_13_4540, i_13_4558, o_13_138);
	kernel_13_139 k_13_139(i_13_135, i_13_136, i_13_181, i_13_255, i_13_264, i_13_418, i_13_517, i_13_535, i_13_577, i_13_624, i_13_640, i_13_643, i_13_685, i_13_689, i_13_696, i_13_718, i_13_777, i_13_778, i_13_891, i_13_894, i_13_928, i_13_975, i_13_976, i_13_1079, i_13_1120, i_13_1152, i_13_1210, i_13_1257, i_13_1269, i_13_1277, i_13_1359, i_13_1386, i_13_1387, i_13_1390, i_13_1407, i_13_1412, i_13_1462, i_13_1465, i_13_1479, i_13_1480, i_13_1484, i_13_1669, i_13_1677, i_13_1683, i_13_1687, i_13_1711, i_13_1756, i_13_1792, i_13_1800, i_13_1858, i_13_1861, i_13_1907, i_13_2191, i_13_2379, i_13_2404, i_13_2442, i_13_2503, i_13_2542, i_13_2586, i_13_2646, i_13_2647, i_13_2687, i_13_2718, i_13_2746, i_13_2844, i_13_2845, i_13_2872, i_13_2874, i_13_2875, i_13_2884, i_13_3224, i_13_3343, i_13_3352, i_13_3384, i_13_3392, i_13_3402, i_13_3415, i_13_3429, i_13_3558, i_13_3567, i_13_3735, i_13_3766, i_13_3790, i_13_3791, i_13_3836, i_13_3933, i_13_4063, i_13_4077, i_13_4086, i_13_4097, i_13_4185, i_13_4186, i_13_4216, i_13_4294, i_13_4296, i_13_4306, i_13_4375, i_13_4433, i_13_4444, i_13_4599, o_13_139);
	kernel_13_140 k_13_140(i_13_39, i_13_80, i_13_105, i_13_159, i_13_169, i_13_247, i_13_268, i_13_337, i_13_339, i_13_340, i_13_373, i_13_386, i_13_466, i_13_490, i_13_607, i_13_610, i_13_618, i_13_661, i_13_780, i_13_816, i_13_817, i_13_886, i_13_931, i_13_979, i_13_1084, i_13_1147, i_13_1150, i_13_1185, i_13_1210, i_13_1248, i_13_1255, i_13_1265, i_13_1302, i_13_1303, i_13_1304, i_13_1313, i_13_1464, i_13_1600, i_13_1725, i_13_1750, i_13_1763, i_13_1806, i_13_1807, i_13_1815, i_13_1816, i_13_1934, i_13_2106, i_13_2130, i_13_2139, i_13_2140, i_13_2141, i_13_2266, i_13_2267, i_13_2410, i_13_2446, i_13_2463, i_13_2484, i_13_2657, i_13_2705, i_13_2752, i_13_2759, i_13_2824, i_13_2859, i_13_2918, i_13_2941, i_13_3001, i_13_3219, i_13_3220, i_13_3250, i_13_3272, i_13_3292, i_13_3308, i_13_3392, i_13_3416, i_13_3476, i_13_3479, i_13_3482, i_13_3505, i_13_3733, i_13_3874, i_13_3910, i_13_3913, i_13_3931, i_13_3991, i_13_4015, i_13_4016, i_13_4066, i_13_4136, i_13_4162, i_13_4232, i_13_4237, i_13_4273, i_13_4309, i_13_4310, i_13_4317, i_13_4319, i_13_4371, i_13_4372, i_13_4381, i_13_4497, o_13_140);
	kernel_13_141 k_13_141(i_13_45, i_13_91, i_13_95, i_13_116, i_13_139, i_13_164, i_13_165, i_13_167, i_13_175, i_13_180, i_13_185, i_13_310, i_13_319, i_13_412, i_13_455, i_13_568, i_13_648, i_13_696, i_13_697, i_13_698, i_13_743, i_13_763, i_13_813, i_13_853, i_13_858, i_13_898, i_13_961, i_13_978, i_13_981, i_13_982, i_13_984, i_13_1065, i_13_1067, i_13_1133, i_13_1219, i_13_1360, i_13_1394, i_13_1405, i_13_1408, i_13_1515, i_13_1517, i_13_1526, i_13_1664, i_13_1695, i_13_1777, i_13_1790, i_13_1831, i_13_1832, i_13_1849, i_13_1852, i_13_1885, i_13_2046, i_13_2097, i_13_2246, i_13_2265, i_13_2356, i_13_2404, i_13_2407, i_13_2437, i_13_2469, i_13_2473, i_13_2532, i_13_2544, i_13_2691, i_13_2921, i_13_2982, i_13_2983, i_13_2984, i_13_3000, i_13_3006, i_13_3059, i_13_3108, i_13_3110, i_13_3145, i_13_3159, i_13_3205, i_13_3207, i_13_3208, i_13_3209, i_13_3210, i_13_3211, i_13_3343, i_13_3355, i_13_3406, i_13_3428, i_13_3511, i_13_3764, i_13_3793, i_13_3819, i_13_3907, i_13_3911, i_13_3931, i_13_3995, i_13_4063, i_13_4066, i_13_4182, i_13_4375, i_13_4519, i_13_4564, i_13_4567, o_13_141);
	kernel_13_142 k_13_142(i_13_106, i_13_107, i_13_112, i_13_124, i_13_367, i_13_607, i_13_624, i_13_625, i_13_858, i_13_870, i_13_948, i_13_1069, i_13_1070, i_13_1075, i_13_1086, i_13_1087, i_13_1203, i_13_1348, i_13_1473, i_13_1474, i_13_1518, i_13_1519, i_13_1571, i_13_1572, i_13_1573, i_13_1574, i_13_1623, i_13_1632, i_13_1642, i_13_1780, i_13_1789, i_13_1795, i_13_1804, i_13_1840, i_13_1843, i_13_1869, i_13_1993, i_13_2024, i_13_2059, i_13_2060, i_13_2120, i_13_2137, i_13_2173, i_13_2191, i_13_2267, i_13_2348, i_13_2380, i_13_2407, i_13_2417, i_13_2429, i_13_2434, i_13_2437, i_13_2536, i_13_2563, i_13_2705, i_13_2715, i_13_2716, i_13_2767, i_13_2986, i_13_2998, i_13_3103, i_13_3126, i_13_3145, i_13_3147, i_13_3148, i_13_3166, i_13_3238, i_13_3274, i_13_3343, i_13_3346, i_13_3373, i_13_3378, i_13_3392, i_13_3418, i_13_3419, i_13_3423, i_13_3427, i_13_3454, i_13_3527, i_13_3544, i_13_3554, i_13_3561, i_13_3767, i_13_3874, i_13_3937, i_13_3994, i_13_4021, i_13_4045, i_13_4048, i_13_4093, i_13_4119, i_13_4120, i_13_4237, i_13_4328, i_13_4342, i_13_4353, i_13_4399, i_13_4417, i_13_4544, i_13_4561, o_13_142);
	kernel_13_143 k_13_143(i_13_41, i_13_52, i_13_53, i_13_142, i_13_194, i_13_196, i_13_283, i_13_314, i_13_319, i_13_320, i_13_325, i_13_326, i_13_463, i_13_464, i_13_580, i_13_592, i_13_647, i_13_661, i_13_688, i_13_689, i_13_691, i_13_692, i_13_707, i_13_817, i_13_818, i_13_826, i_13_844, i_13_848, i_13_862, i_13_1019, i_13_1124, i_13_1255, i_13_1316, i_13_1358, i_13_1445, i_13_1471, i_13_1489, i_13_1492, i_13_1574, i_13_1600, i_13_1672, i_13_1852, i_13_1876, i_13_1955, i_13_1997, i_13_2173, i_13_2177, i_13_2185, i_13_2195, i_13_2264, i_13_2266, i_13_2267, i_13_2383, i_13_2408, i_13_2410, i_13_2411, i_13_2591, i_13_2600, i_13_2653, i_13_2654, i_13_2699, i_13_2860, i_13_2914, i_13_2918, i_13_2941, i_13_3067, i_13_3068, i_13_3077, i_13_3145, i_13_3146, i_13_3292, i_13_3373, i_13_3374, i_13_3392, i_13_3479, i_13_3527, i_13_3541, i_13_3595, i_13_3722, i_13_3733, i_13_3770, i_13_3781, i_13_3821, i_13_3982, i_13_3985, i_13_3995, i_13_4021, i_13_4022, i_13_4066, i_13_4067, i_13_4171, i_13_4318, i_13_4319, i_13_4369, i_13_4372, i_13_4448, i_13_4513, i_13_4540, i_13_4559, i_13_4598, o_13_143);
	kernel_13_144 k_13_144(i_13_20, i_13_77, i_13_78, i_13_107, i_13_113, i_13_174, i_13_195, i_13_368, i_13_386, i_13_454, i_13_460, i_13_502, i_13_528, i_13_725, i_13_814, i_13_859, i_13_949, i_13_1087, i_13_1088, i_13_1148, i_13_1211, i_13_1219, i_13_1348, i_13_1394, i_13_1399, i_13_1410, i_13_1426, i_13_1474, i_13_1509, i_13_1570, i_13_1573, i_13_1622, i_13_1624, i_13_1633, i_13_1741, i_13_1789, i_13_1804, i_13_1840, i_13_1841, i_13_1844, i_13_1942, i_13_2001, i_13_2024, i_13_2059, i_13_2123, i_13_2128, i_13_2137, i_13_2230, i_13_2283, i_13_2284, i_13_2317, i_13_2348, i_13_2383, i_13_2399, i_13_2435, i_13_2437, i_13_2438, i_13_2501, i_13_2716, i_13_2717, i_13_2749, i_13_2856, i_13_3023, i_13_3066, i_13_3067, i_13_3127, i_13_3137, i_13_3144, i_13_3147, i_13_3148, i_13_3149, i_13_3166, i_13_3167, i_13_3329, i_13_3343, i_13_3374, i_13_3392, i_13_3413, i_13_3428, i_13_3432, i_13_3455, i_13_3553, i_13_3599, i_13_3923, i_13_4111, i_13_4120, i_13_4121, i_13_4192, i_13_4256, i_13_4263, i_13_4264, i_13_4328, i_13_4333, i_13_4400, i_13_4417, i_13_4418, i_13_4469, i_13_4526, i_13_4544, i_13_4596, o_13_144);
	kernel_13_145 k_13_145(i_13_106, i_13_187, i_13_284, i_13_337, i_13_339, i_13_427, i_13_454, i_13_513, i_13_526, i_13_553, i_13_589, i_13_607, i_13_646, i_13_651, i_13_673, i_13_679, i_13_688, i_13_691, i_13_694, i_13_699, i_13_733, i_13_823, i_13_840, i_13_898, i_13_925, i_13_1033, i_13_1101, i_13_1123, i_13_1144, i_13_1148, i_13_1179, i_13_1180, i_13_1226, i_13_1270, i_13_1272, i_13_1273, i_13_1318, i_13_1345, i_13_1384, i_13_1449, i_13_1519, i_13_1570, i_13_1633, i_13_1656, i_13_1657, i_13_1750, i_13_1840, i_13_1858, i_13_1915, i_13_1930, i_13_1933, i_13_1935, i_13_2002, i_13_2029, i_13_2088, i_13_2200, i_13_2209, i_13_2461, i_13_2494, i_13_2496, i_13_2542, i_13_2600, i_13_2653, i_13_2736, i_13_2767, i_13_2770, i_13_2845, i_13_2848, i_13_2886, i_13_3055, i_13_3145, i_13_3151, i_13_3258, i_13_3316, i_13_3370, i_13_3378, i_13_3382, i_13_3418, i_13_3431, i_13_3505, i_13_3535, i_13_3561, i_13_3730, i_13_3736, i_13_3739, i_13_3756, i_13_3846, i_13_3892, i_13_3927, i_13_4021, i_13_4036, i_13_4081, i_13_4158, i_13_4188, i_13_4189, i_13_4315, i_13_4417, i_13_4578, i_13_4594, i_13_4602, o_13_145);
	kernel_13_146 k_13_146(i_13_28, i_13_32, i_13_46, i_13_49, i_13_65, i_13_91, i_13_92, i_13_118, i_13_122, i_13_157, i_13_163, i_13_317, i_13_320, i_13_454, i_13_562, i_13_568, i_13_671, i_13_676, i_13_697, i_13_722, i_13_730, i_13_758, i_13_946, i_13_1075, i_13_1076, i_13_1381, i_13_1405, i_13_1442, i_13_1454, i_13_1526, i_13_1606, i_13_1621, i_13_1630, i_13_1633, i_13_1837, i_13_1846, i_13_1955, i_13_1999, i_13_2000, i_13_2173, i_13_2174, i_13_2206, i_13_2207, i_13_2422, i_13_2431, i_13_2432, i_13_2452, i_13_2548, i_13_2559, i_13_2719, i_13_2750, i_13_2793, i_13_2846, i_13_2884, i_13_3019, i_13_3034, i_13_3035, i_13_3126, i_13_3127, i_13_3161, i_13_3164, i_13_3214, i_13_3242, i_13_3272, i_13_3415, i_13_3421, i_13_3422, i_13_3434, i_13_3449, i_13_3477, i_13_3528, i_13_3530, i_13_3637, i_13_3638, i_13_3646, i_13_3647, i_13_3699, i_13_3700, i_13_3718, i_13_3837, i_13_3843, i_13_3844, i_13_3857, i_13_3871, i_13_3872, i_13_3889, i_13_3901, i_13_4006, i_13_4007, i_13_4042, i_13_4043, i_13_4105, i_13_4177, i_13_4304, i_13_4312, i_13_4348, i_13_4349, i_13_4351, i_13_4387, i_13_4510, o_13_146);
	kernel_13_147 k_13_147(i_13_26, i_13_34, i_13_76, i_13_79, i_13_102, i_13_115, i_13_127, i_13_128, i_13_140, i_13_142, i_13_230, i_13_232, i_13_233, i_13_268, i_13_362, i_13_538, i_13_539, i_13_573, i_13_620, i_13_690, i_13_691, i_13_696, i_13_697, i_13_699, i_13_700, i_13_768, i_13_814, i_13_826, i_13_827, i_13_857, i_13_885, i_13_1066, i_13_1123, i_13_1219, i_13_1220, i_13_1222, i_13_1275, i_13_1391, i_13_1440, i_13_1629, i_13_1714, i_13_1718, i_13_1726, i_13_1777, i_13_1795, i_13_1804, i_13_1807, i_13_1843, i_13_1888, i_13_2006, i_13_2101, i_13_2119, i_13_2317, i_13_2342, i_13_2410, i_13_2434, i_13_2469, i_13_2472, i_13_2654, i_13_2657, i_13_2713, i_13_2722, i_13_2726, i_13_2851, i_13_3028, i_13_3038, i_13_3067, i_13_3100, i_13_3145, i_13_3146, i_13_3148, i_13_3208, i_13_3211, i_13_3313, i_13_3419, i_13_3443, i_13_3490, i_13_3501, i_13_3505, i_13_3506, i_13_3557, i_13_3571, i_13_3572, i_13_3685, i_13_3741, i_13_3742, i_13_3743, i_13_4063, i_13_4084, i_13_4092, i_13_4208, i_13_4256, i_13_4269, i_13_4297, i_13_4298, i_13_4316, i_13_4367, i_13_4399, i_13_4513, i_13_4538, o_13_147);
	kernel_13_148 k_13_148(i_13_61, i_13_71, i_13_179, i_13_274, i_13_275, i_13_280, i_13_286, i_13_493, i_13_529, i_13_530, i_13_553, i_13_562, i_13_599, i_13_673, i_13_797, i_13_841, i_13_853, i_13_854, i_13_965, i_13_1025, i_13_1075, i_13_1147, i_13_1282, i_13_1303, i_13_1304, i_13_1321, i_13_1327, i_13_1490, i_13_1502, i_13_1516, i_13_1552, i_13_1553, i_13_1660, i_13_1700, i_13_1817, i_13_1858, i_13_2002, i_13_2003, i_13_2020, i_13_2021, i_13_2050, i_13_2201, i_13_2240, i_13_2263, i_13_2275, i_13_2366, i_13_2461, i_13_2462, i_13_2470, i_13_2471, i_13_2509, i_13_2543, i_13_2551, i_13_2615, i_13_2653, i_13_2824, i_13_2825, i_13_2860, i_13_2920, i_13_2984, i_13_3173, i_13_3274, i_13_3347, i_13_3418, i_13_3424, i_13_3428, i_13_3482, i_13_3533, i_13_3541, i_13_3542, i_13_3544, i_13_3545, i_13_3580, i_13_3614, i_13_3622, i_13_3634, i_13_3730, i_13_3731, i_13_3743, i_13_3787, i_13_3788, i_13_3910, i_13_3911, i_13_3913, i_13_3914, i_13_4118, i_13_4126, i_13_4162, i_13_4189, i_13_4237, i_13_4238, i_13_4256, i_13_4282, i_13_4378, i_13_4381, i_13_4382, i_13_4400, i_13_4567, i_13_4594, i_13_4604, o_13_148);
	kernel_13_149 k_13_149(i_13_63, i_13_207, i_13_265, i_13_306, i_13_354, i_13_370, i_13_372, i_13_381, i_13_409, i_13_414, i_13_462, i_13_463, i_13_466, i_13_467, i_13_588, i_13_589, i_13_595, i_13_660, i_13_666, i_13_670, i_13_697, i_13_759, i_13_948, i_13_1179, i_13_1344, i_13_1349, i_13_1549, i_13_1569, i_13_1594, i_13_1603, i_13_1767, i_13_1845, i_13_1846, i_13_1854, i_13_1947, i_13_1959, i_13_1993, i_13_2028, i_13_2029, i_13_2100, i_13_2137, i_13_2142, i_13_2199, i_13_2200, i_13_2204, i_13_2263, i_13_2280, i_13_2434, i_13_2457, i_13_2503, i_13_2506, i_13_2511, i_13_2554, i_13_2559, i_13_2820, i_13_2821, i_13_2856, i_13_2880, i_13_2982, i_13_3000, i_13_3001, i_13_3046, i_13_3130, i_13_3144, i_13_3213, i_13_3240, i_13_3241, i_13_3343, i_13_3387, i_13_3392, i_13_3411, i_13_3412, i_13_3480, i_13_3537, i_13_3538, i_13_3567, i_13_3592, i_13_3594, i_13_3595, i_13_3618, i_13_3619, i_13_3630, i_13_3631, i_13_3634, i_13_3636, i_13_3637, i_13_3666, i_13_3670, i_13_3766, i_13_3846, i_13_3906, i_13_3915, i_13_4060, i_13_4162, i_13_4269, i_13_4316, i_13_4324, i_13_4327, i_13_4368, i_13_4443, o_13_149);
	kernel_13_150 k_13_150(i_13_136, i_13_139, i_13_166, i_13_190, i_13_229, i_13_251, i_13_374, i_13_419, i_13_508, i_13_536, i_13_545, i_13_556, i_13_613, i_13_614, i_13_622, i_13_646, i_13_665, i_13_695, i_13_698, i_13_713, i_13_793, i_13_814, i_13_895, i_13_939, i_13_952, i_13_979, i_13_1021, i_13_1094, i_13_1117, i_13_1120, i_13_1130, i_13_1228, i_13_1249, i_13_1252, i_13_1273, i_13_1390, i_13_1467, i_13_1480, i_13_1484, i_13_1502, i_13_1642, i_13_1670, i_13_1675, i_13_1757, i_13_1759, i_13_1778, i_13_1795, i_13_1796, i_13_1825, i_13_1947, i_13_1960, i_13_2004, i_13_2030, i_13_2111, i_13_2245, i_13_2288, i_13_2380, i_13_2407, i_13_2408, i_13_2464, i_13_2552, i_13_2615, i_13_2747, i_13_2750, i_13_2767, i_13_2848, i_13_2849, i_13_2850, i_13_2851, i_13_2875, i_13_2882, i_13_2976, i_13_3088, i_13_3092, i_13_3116, i_13_3256, i_13_3368, i_13_3371, i_13_3460, i_13_3556, i_13_3638, i_13_3730, i_13_3794, i_13_3839, i_13_3929, i_13_3997, i_13_4055, i_13_4064, i_13_4117, i_13_4138, i_13_4186, i_13_4189, i_13_4190, i_13_4197, i_13_4294, i_13_4296, i_13_4297, i_13_4337, i_13_4344, i_13_4515, o_13_150);
	kernel_13_151 k_13_151(i_13_113, i_13_121, i_13_137, i_13_138, i_13_139, i_13_140, i_13_143, i_13_175, i_13_229, i_13_231, i_13_260, i_13_340, i_13_380, i_13_473, i_13_535, i_13_536, i_13_537, i_13_573, i_13_574, i_13_725, i_13_832, i_13_850, i_13_853, i_13_868, i_13_869, i_13_985, i_13_1216, i_13_1219, i_13_1228, i_13_1470, i_13_1475, i_13_1540, i_13_1546, i_13_1547, i_13_1552, i_13_1667, i_13_1711, i_13_1714, i_13_1715, i_13_1723, i_13_1724, i_13_1725, i_13_1726, i_13_1734, i_13_1787, i_13_1831, i_13_1840, i_13_1841, i_13_1849, i_13_1858, i_13_1940, i_13_1993, i_13_2128, i_13_2156, i_13_2158, i_13_2345, i_13_2467, i_13_2570, i_13_2692, i_13_2695, i_13_2701, i_13_2712, i_13_2845, i_13_2848, i_13_3010, i_13_3011, i_13_3037, i_13_3064, i_13_3065, i_13_3066, i_13_3109, i_13_3146, i_13_3174, i_13_3229, i_13_3293, i_13_3444, i_13_3452, i_13_3478, i_13_3487, i_13_3524, i_13_3541, i_13_3570, i_13_3686, i_13_3688, i_13_3701, i_13_3739, i_13_3799, i_13_3836, i_13_4054, i_13_4058, i_13_4063, i_13_4151, i_13_4193, i_13_4234, i_13_4369, i_13_4378, i_13_4394, i_13_4411, i_13_4415, i_13_4523, o_13_151);
	kernel_13_152 k_13_152(i_13_50, i_13_73, i_13_102, i_13_137, i_13_189, i_13_252, i_13_280, i_13_407, i_13_434, i_13_441, i_13_515, i_13_559, i_13_617, i_13_623, i_13_659, i_13_661, i_13_666, i_13_693, i_13_694, i_13_695, i_13_696, i_13_838, i_13_839, i_13_921, i_13_975, i_13_1072, i_13_1073, i_13_1109, i_13_1116, i_13_1117, i_13_1118, i_13_1145, i_13_1270, i_13_1423, i_13_1424, i_13_1427, i_13_1657, i_13_1658, i_13_1730, i_13_1742, i_13_1791, i_13_1858, i_13_2016, i_13_2017, i_13_2020, i_13_2021, i_13_2207, i_13_2209, i_13_2324, i_13_2344, i_13_2443, i_13_2452, i_13_2453, i_13_2461, i_13_2467, i_13_2512, i_13_2513, i_13_2551, i_13_2552, i_13_2718, i_13_2741, i_13_2880, i_13_2881, i_13_2882, i_13_2883, i_13_2956, i_13_3001, i_13_3074, i_13_3089, i_13_3091, i_13_3107, i_13_3269, i_13_3371, i_13_3416, i_13_3424, i_13_3476, i_13_3487, i_13_3532, i_13_3547, i_13_3646, i_13_3740, i_13_3820, i_13_3862, i_13_3919, i_13_3987, i_13_3989, i_13_4252, i_13_4293, i_13_4315, i_13_4324, i_13_4330, i_13_4331, i_13_4429, i_13_4450, i_13_4451, i_13_4455, i_13_4591, i_13_4592, i_13_4600, i_13_4601, o_13_152);
	kernel_13_153 k_13_153(i_13_138, i_13_139, i_13_184, i_13_226, i_13_280, i_13_380, i_13_415, i_13_524, i_13_585, i_13_651, i_13_675, i_13_832, i_13_1074, i_13_1182, i_13_1200, i_13_1206, i_13_1207, i_13_1252, i_13_1296, i_13_1297, i_13_1341, i_13_1342, i_13_1468, i_13_1515, i_13_1516, i_13_1711, i_13_1712, i_13_1720, i_13_1722, i_13_1723, i_13_1777, i_13_1778, i_13_1881, i_13_1882, i_13_1884, i_13_1923, i_13_1924, i_13_1926, i_13_1989, i_13_1990, i_13_1999, i_13_2001, i_13_2020, i_13_2052, i_13_2133, i_13_2134, i_13_2169, i_13_2277, i_13_2377, i_13_2470, i_13_2548, i_13_2646, i_13_2647, i_13_2676, i_13_2694, i_13_2710, i_13_2787, i_13_2853, i_13_2872, i_13_2934, i_13_2983, i_13_3037, i_13_3132, i_13_3208, i_13_3343, i_13_3384, i_13_3414, i_13_3415, i_13_3438, i_13_3445, i_13_3447, i_13_3448, i_13_3474, i_13_3475, i_13_3547, i_13_3592, i_13_3615, i_13_3616, i_13_3645, i_13_3646, i_13_3663, i_13_3684, i_13_3736, i_13_3820, i_13_3987, i_13_3988, i_13_4050, i_13_4053, i_13_4077, i_13_4117, i_13_4159, i_13_4203, i_13_4270, i_13_4338, i_13_4392, i_13_4393, i_13_4410, i_13_4411, i_13_4554, i_13_4567, o_13_153);
	kernel_13_154 k_13_154(i_13_34, i_13_67, i_13_78, i_13_114, i_13_135, i_13_138, i_13_141, i_13_156, i_13_178, i_13_189, i_13_192, i_13_282, i_13_285, i_13_373, i_13_381, i_13_385, i_13_508, i_13_585, i_13_588, i_13_589, i_13_1119, i_13_1209, i_13_1281, i_13_1300, i_13_1312, i_13_1344, i_13_1399, i_13_1402, i_13_1407, i_13_1429, i_13_1443, i_13_1482, i_13_1515, i_13_1725, i_13_1770, i_13_1771, i_13_1778, i_13_1779, i_13_1812, i_13_1813, i_13_1884, i_13_1885, i_13_1888, i_13_1903, i_13_1924, i_13_1992, i_13_1995, i_13_2002, i_13_2004, i_13_2005, i_13_2020, i_13_2055, i_13_2118, i_13_2190, i_13_2193, i_13_2199, i_13_2235, i_13_2280, i_13_2281, i_13_2454, i_13_2595, i_13_2712, i_13_2721, i_13_2725, i_13_2726, i_13_2856, i_13_2857, i_13_2860, i_13_2899, i_13_2937, i_13_2959, i_13_3236, i_13_3274, i_13_3417, i_13_3418, i_13_3441, i_13_3453, i_13_3466, i_13_3477, i_13_3478, i_13_3481, i_13_3523, i_13_3595, i_13_3613, i_13_3666, i_13_3721, i_13_3729, i_13_3758, i_13_3769, i_13_3860, i_13_3897, i_13_3986, i_13_4017, i_13_4054, i_13_4217, i_13_4233, i_13_4395, i_13_4396, i_13_4399, i_13_4567, o_13_154);
	kernel_13_155 k_13_155(i_13_44, i_13_67, i_13_70, i_13_75, i_13_95, i_13_124, i_13_269, i_13_271, i_13_310, i_13_314, i_13_322, i_13_346, i_13_361, i_13_410, i_13_412, i_13_445, i_13_466, i_13_590, i_13_592, i_13_593, i_13_622, i_13_646, i_13_647, i_13_657, i_13_688, i_13_689, i_13_700, i_13_763, i_13_764, i_13_811, i_13_842, i_13_955, i_13_1120, i_13_1124, i_13_1132, i_13_1207, i_13_1261, i_13_1283, i_13_1285, i_13_1286, i_13_1312, i_13_1349, i_13_1511, i_13_1513, i_13_1601, i_13_1636, i_13_1728, i_13_1741, i_13_1754, i_13_1781, i_13_1799, i_13_1807, i_13_1997, i_13_2056, i_13_2057, i_13_2059, i_13_2060, i_13_2104, i_13_2123, i_13_2141, i_13_2195, i_13_2266, i_13_2267, i_13_2272, i_13_2377, i_13_2384, i_13_2426, i_13_2455, i_13_2512, i_13_2545, i_13_2555, i_13_2653, i_13_2680, i_13_2851, i_13_2939, i_13_3043, i_13_3175, i_13_3274, i_13_3346, i_13_3347, i_13_3391, i_13_3392, i_13_3640, i_13_3641, i_13_3722, i_13_3877, i_13_3905, i_13_3940, i_13_3994, i_13_4036, i_13_4037, i_13_4039, i_13_4040, i_13_4085, i_13_4144, i_13_4342, i_13_4382, i_13_4595, i_13_4597, i_13_4598, o_13_155);
	kernel_13_156 k_13_156(i_13_73, i_13_103, i_13_109, i_13_184, i_13_193, i_13_248, i_13_379, i_13_446, i_13_454, i_13_524, i_13_554, i_13_571, i_13_572, i_13_589, i_13_590, i_13_715, i_13_742, i_13_743, i_13_859, i_13_946, i_13_947, i_13_1021, i_13_1085, i_13_1140, i_13_1209, i_13_1228, i_13_1248, i_13_1255, i_13_1286, i_13_1345, i_13_1346, i_13_1397, i_13_1408, i_13_1427, i_13_1444, i_13_1571, i_13_1597, i_13_1607, i_13_1629, i_13_1678, i_13_1750, i_13_1777, i_13_1831, i_13_1858, i_13_1918, i_13_1930, i_13_1931, i_13_1940, i_13_1941, i_13_1948, i_13_1954, i_13_2002, i_13_2056, i_13_2057, i_13_2188, i_13_2281, i_13_2282, i_13_2299, i_13_2506, i_13_2512, i_13_2515, i_13_2614, i_13_2710, i_13_2713, i_13_2714, i_13_2719, i_13_2720, i_13_2723, i_13_2750, i_13_2768, i_13_2784, i_13_2785, i_13_2857, i_13_2858, i_13_2916, i_13_3065, i_13_3145, i_13_3154, i_13_3344, i_13_3370, i_13_3439, i_13_3596, i_13_3616, i_13_3617, i_13_3631, i_13_3681, i_13_3683, i_13_3685, i_13_3727, i_13_3920, i_13_3956, i_13_4037, i_13_4046, i_13_4091, i_13_4280, i_13_4330, i_13_4385, i_13_4396, i_13_4426, i_13_4555, o_13_156);
	kernel_13_157 k_13_157(i_13_40, i_13_51, i_13_74, i_13_91, i_13_94, i_13_139, i_13_142, i_13_164, i_13_172, i_13_241, i_13_248, i_13_251, i_13_338, i_13_365, i_13_371, i_13_420, i_13_480, i_13_533, i_13_580, i_13_581, i_13_620, i_13_640, i_13_641, i_13_663, i_13_677, i_13_699, i_13_861, i_13_977, i_13_979, i_13_985, i_13_1098, i_13_1281, i_13_1284, i_13_1428, i_13_1462, i_13_1468, i_13_1487, i_13_1499, i_13_1553, i_13_1633, i_13_1634, i_13_1658, i_13_1720, i_13_1775, i_13_1885, i_13_1918, i_13_1990, i_13_1994, i_13_2050, i_13_2174, i_13_2348, i_13_2457, i_13_2507, i_13_2544, i_13_2552, i_13_2650, i_13_2788, i_13_2845, i_13_2846, i_13_2885, i_13_2888, i_13_2910, i_13_2924, i_13_2936, i_13_2949, i_13_2956, i_13_3208, i_13_3448, i_13_3449, i_13_3511, i_13_3524, i_13_3568, i_13_3572, i_13_3581, i_13_3638, i_13_3647, i_13_3652, i_13_3685, i_13_3686, i_13_3689, i_13_3736, i_13_3769, i_13_3847, i_13_3853, i_13_3905, i_13_3917, i_13_3988, i_13_4021, i_13_4036, i_13_4079, i_13_4088, i_13_4117, i_13_4260, i_13_4351, i_13_4352, i_13_4371, i_13_4391, i_13_4568, i_13_4576, i_13_4601, o_13_157);
	kernel_13_158 k_13_158(i_13_28, i_13_36, i_13_37, i_13_138, i_13_171, i_13_174, i_13_280, i_13_313, i_13_333, i_13_562, i_13_639, i_13_642, i_13_643, i_13_646, i_13_675, i_13_679, i_13_684, i_13_685, i_13_687, i_13_688, i_13_778, i_13_820, i_13_823, i_13_849, i_13_1119, i_13_1224, i_13_1269, i_13_1273, i_13_1305, i_13_1461, i_13_1521, i_13_1636, i_13_1668, i_13_1713, i_13_1749, i_13_1839, i_13_1855, i_13_1858, i_13_1881, i_13_1882, i_13_1884, i_13_2424, i_13_2457, i_13_2505, i_13_2559, i_13_2584, i_13_2646, i_13_2649, i_13_2650, i_13_2673, i_13_2677, i_13_2694, i_13_2730, i_13_2844, i_13_2847, i_13_2848, i_13_2874, i_13_2919, i_13_3088, i_13_3093, i_13_3094, i_13_3144, i_13_3234, i_13_3261, i_13_3270, i_13_3271, i_13_3304, i_13_3378, i_13_3387, i_13_3388, i_13_3420, i_13_3421, i_13_3423, i_13_3424, i_13_3429, i_13_3523, i_13_3561, i_13_3648, i_13_3721, i_13_3738, i_13_3798, i_13_3819, i_13_3924, i_13_3930, i_13_3987, i_13_4017, i_13_4036, i_13_4077, i_13_4080, i_13_4081, i_13_4185, i_13_4186, i_13_4257, i_13_4293, i_13_4339, i_13_4350, i_13_4465, i_13_4593, i_13_4594, i_13_4597, o_13_158);
	kernel_13_159 k_13_159(i_13_67, i_13_74, i_13_121, i_13_122, i_13_140, i_13_281, i_13_325, i_13_373, i_13_379, i_13_406, i_13_442, i_13_443, i_13_463, i_13_532, i_13_589, i_13_622, i_13_641, i_13_677, i_13_715, i_13_742, i_13_760, i_13_769, i_13_814, i_13_820, i_13_821, i_13_824, i_13_859, i_13_860, i_13_919, i_13_928, i_13_929, i_13_959, i_13_1030, i_13_1066, i_13_1082, i_13_1100, i_13_1129, i_13_1196, i_13_1226, i_13_1250, i_13_1256, i_13_1301, i_13_1331, i_13_1489, i_13_1490, i_13_1642, i_13_1712, i_13_1751, i_13_1793, i_13_1804, i_13_1883, i_13_1942, i_13_1990, i_13_1991, i_13_2012, i_13_2056, i_13_2117, i_13_2260, i_13_2263, i_13_2344, i_13_2380, i_13_2470, i_13_2542, i_13_2611, i_13_2675, i_13_2767, i_13_2768, i_13_2846, i_13_2920, i_13_2983, i_13_3004, i_13_3019, i_13_3110, i_13_3164, i_13_3259, i_13_3286, i_13_3287, i_13_3343, i_13_3386, i_13_3416, i_13_3421, i_13_3422, i_13_3430, i_13_3434, i_13_3502, i_13_3503, i_13_3731, i_13_3736, i_13_3740, i_13_3794, i_13_3802, i_13_3874, i_13_3890, i_13_3892, i_13_3898, i_13_3919, i_13_4078, i_13_4079, i_13_4270, i_13_4595, o_13_159);
	kernel_13_160 k_13_160(i_13_38, i_13_71, i_13_95, i_13_201, i_13_233, i_13_263, i_13_308, i_13_337, i_13_344, i_13_412, i_13_527, i_13_533, i_13_556, i_13_628, i_13_643, i_13_646, i_13_653, i_13_666, i_13_683, i_13_712, i_13_827, i_13_845, i_13_897, i_13_956, i_13_979, i_13_1120, i_13_1123, i_13_1155, i_13_1275, i_13_1276, i_13_1312, i_13_1333, i_13_1381, i_13_1390, i_13_1447, i_13_1462, i_13_1482, i_13_1499, i_13_1561, i_13_1570, i_13_1600, i_13_1645, i_13_1646, i_13_1664, i_13_1670, i_13_1678, i_13_1727, i_13_1753, i_13_1797, i_13_1882, i_13_1953, i_13_2040, i_13_2074, i_13_2231, i_13_2277, i_13_2310, i_13_2315, i_13_2378, i_13_2381, i_13_2384, i_13_2434, i_13_2548, i_13_2549, i_13_2570, i_13_2616, i_13_2634, i_13_2686, i_13_2687, i_13_2887, i_13_3082, i_13_3087, i_13_3197, i_13_3214, i_13_3241, i_13_3296, i_13_3355, i_13_3435, i_13_3597, i_13_3652, i_13_3739, i_13_3743, i_13_3781, i_13_3786, i_13_3838, i_13_3994, i_13_4063, i_13_4083, i_13_4097, i_13_4187, i_13_4296, i_13_4351, i_13_4369, i_13_4381, i_13_4418, i_13_4502, i_13_4558, i_13_4590, i_13_4595, i_13_4601, i_13_4605, o_13_160);
	kernel_13_161 k_13_161(i_13_57, i_13_76, i_13_79, i_13_111, i_13_177, i_13_243, i_13_265, i_13_411, i_13_606, i_13_607, i_13_609, i_13_628, i_13_657, i_13_660, i_13_661, i_13_663, i_13_669, i_13_850, i_13_915, i_13_942, i_13_947, i_13_1018, i_13_1020, i_13_1023, i_13_1060, i_13_1075, i_13_1134, i_13_1150, i_13_1213, i_13_1317, i_13_1425, i_13_1426, i_13_1428, i_13_1429, i_13_1571, i_13_1597, i_13_1632, i_13_1732, i_13_1849, i_13_1857, i_13_1858, i_13_2022, i_13_2023, i_13_2373, i_13_2407, i_13_2451, i_13_2454, i_13_2455, i_13_2498, i_13_2572, i_13_2740, i_13_2908, i_13_2938, i_13_3009, i_13_3012, i_13_3016, i_13_3124, i_13_3145, i_13_3148, i_13_3175, i_13_3250, i_13_3264, i_13_3273, i_13_3321, i_13_3403, i_13_3459, i_13_3486, i_13_3487, i_13_3530, i_13_3570, i_13_3640, i_13_3706, i_13_3783, i_13_3790, i_13_3864, i_13_3865, i_13_3894, i_13_3990, i_13_4021, i_13_4054, i_13_4057, i_13_4083, i_13_4095, i_13_4117, i_13_4119, i_13_4189, i_13_4252, i_13_4254, i_13_4255, i_13_4261, i_13_4263, i_13_4327, i_13_4368, i_13_4369, i_13_4370, i_13_4371, i_13_4471, i_13_4557, i_13_4560, i_13_4596, o_13_161);
	kernel_13_162 k_13_162(i_13_91, i_13_92, i_13_94, i_13_95, i_13_102, i_13_120, i_13_185, i_13_200, i_13_308, i_13_316, i_13_317, i_13_335, i_13_571, i_13_572, i_13_617, i_13_651, i_13_668, i_13_671, i_13_730, i_13_794, i_13_947, i_13_950, i_13_1064, i_13_1067, i_13_1093, i_13_1202, i_13_1210, i_13_1211, i_13_1229, i_13_1307, i_13_1318, i_13_1324, i_13_1325, i_13_1405, i_13_1426, i_13_1497, i_13_1514, i_13_1526, i_13_1595, i_13_1631, i_13_1642, i_13_1730, i_13_1757, i_13_1765, i_13_1802, i_13_1812, i_13_1828, i_13_1829, i_13_1850, i_13_1885, i_13_2108, i_13_2117, i_13_2128, i_13_2136, i_13_2206, i_13_2234, i_13_2261, i_13_2264, i_13_2444, i_13_2506, i_13_2539, i_13_2674, i_13_2919, i_13_3109, i_13_3110, i_13_3116, i_13_3164, i_13_3208, i_13_3209, i_13_3242, i_13_3258, i_13_3286, i_13_3395, i_13_3407, i_13_3415, i_13_3416, i_13_3422, i_13_3530, i_13_3766, i_13_3767, i_13_3783, i_13_3785, i_13_3817, i_13_3818, i_13_3872, i_13_3924, i_13_3925, i_13_3987, i_13_3988, i_13_4061, i_13_4132, i_13_4280, i_13_4339, i_13_4342, i_13_4351, i_13_4352, i_13_4379, i_13_4567, i_13_4568, i_13_4591, o_13_162);
	kernel_13_163 k_13_163(i_13_48, i_13_69, i_13_71, i_13_79, i_13_176, i_13_181, i_13_258, i_13_411, i_13_452, i_13_535, i_13_609, i_13_628, i_13_642, i_13_650, i_13_660, i_13_663, i_13_682, i_13_690, i_13_745, i_13_760, i_13_762, i_13_812, i_13_850, i_13_979, i_13_1067, i_13_1119, i_13_1121, i_13_1122, i_13_1132, i_13_1136, i_13_1149, i_13_1271, i_13_1275, i_13_1276, i_13_1311, i_13_1316, i_13_1402, i_13_1506, i_13_1510, i_13_1514, i_13_1516, i_13_1551, i_13_1563, i_13_1572, i_13_1596, i_13_1597, i_13_1676, i_13_1714, i_13_1797, i_13_1798, i_13_1807, i_13_2028, i_13_2057, i_13_2194, i_13_2199, i_13_2425, i_13_2454, i_13_2676, i_13_2678, i_13_2679, i_13_2697, i_13_2724, i_13_2742, i_13_2940, i_13_2953, i_13_2967, i_13_2976, i_13_3094, i_13_3118, i_13_3209, i_13_3264, i_13_3273, i_13_3354, i_13_3368, i_13_3399, i_13_3459, i_13_3487, i_13_3549, i_13_3651, i_13_3652, i_13_3697, i_13_3759, i_13_3764, i_13_3822, i_13_3864, i_13_3930, i_13_3939, i_13_4018, i_13_4037, i_13_4082, i_13_4255, i_13_4272, i_13_4300, i_13_4306, i_13_4335, i_13_4377, i_13_4447, i_13_4515, i_13_4565, i_13_4606, o_13_163);
	kernel_13_164 k_13_164(i_13_3, i_13_40, i_13_62, i_13_94, i_13_112, i_13_115, i_13_127, i_13_184, i_13_187, i_13_207, i_13_225, i_13_234, i_13_244, i_13_266, i_13_268, i_13_333, i_13_538, i_13_607, i_13_670, i_13_769, i_13_814, i_13_1084, i_13_1191, i_13_1205, i_13_1219, i_13_1274, i_13_1321, i_13_1482, i_13_1489, i_13_1538, i_13_1680, i_13_1749, i_13_1750, i_13_1752, i_13_1804, i_13_1807, i_13_1840, i_13_1843, i_13_1845, i_13_1995, i_13_1996, i_13_2128, i_13_2138, i_13_2140, i_13_2142, i_13_2173, i_13_2176, i_13_2304, i_13_2407, i_13_2409, i_13_2425, i_13_2434, i_13_2446, i_13_2494, i_13_2506, i_13_2576, i_13_2581, i_13_2694, i_13_2742, i_13_2745, i_13_2749, i_13_2940, i_13_2965, i_13_3030, i_13_3031, i_13_3100, i_13_3120, i_13_3123, i_13_3135, i_13_3145, i_13_3148, i_13_3163, i_13_3273, i_13_3343, i_13_3373, i_13_3402, i_13_3418, i_13_3504, i_13_3505, i_13_3537, i_13_3569, i_13_3637, i_13_3669, i_13_3739, i_13_3746, i_13_3874, i_13_3878, i_13_3892, i_13_3909, i_13_3912, i_13_3991, i_13_4104, i_13_4120, i_13_4341, i_13_4354, i_13_4378, i_13_4380, i_13_4390, i_13_4461, i_13_4583, o_13_164);
	kernel_13_165 k_13_165(i_13_51, i_13_76, i_13_96, i_13_129, i_13_157, i_13_159, i_13_164, i_13_167, i_13_169, i_13_170, i_13_266, i_13_282, i_13_375, i_13_377, i_13_384, i_13_568, i_13_598, i_13_683, i_13_697, i_13_714, i_13_814, i_13_816, i_13_817, i_13_844, i_13_858, i_13_984, i_13_1068, i_13_1106, i_13_1301, i_13_1511, i_13_1570, i_13_1749, i_13_1777, i_13_1795, i_13_1807, i_13_1829, i_13_1851, i_13_1852, i_13_1857, i_13_1912, i_13_1924, i_13_2108, i_13_2110, i_13_2122, i_13_2139, i_13_2208, i_13_2241, i_13_2264, i_13_2266, i_13_2407, i_13_2425, i_13_2437, i_13_2497, i_13_2554, i_13_2567, i_13_2570, i_13_2679, i_13_2698, i_13_2797, i_13_2848, i_13_2884, i_13_2921, i_13_2940, i_13_2941, i_13_2983, i_13_3030, i_13_3031, i_13_3038, i_13_3110, i_13_3116, i_13_3147, i_13_3208, i_13_3210, i_13_3212, i_13_3239, i_13_3327, i_13_3345, i_13_3400, i_13_3408, i_13_3505, i_13_3732, i_13_3739, i_13_3741, i_13_3767, i_13_3820, i_13_3941, i_13_3994, i_13_4045, i_13_4048, i_13_4061, i_13_4063, i_13_4064, i_13_4066, i_13_4080, i_13_4119, i_13_4309, i_13_4318, i_13_4333, i_13_4397, i_13_4607, o_13_165);
	kernel_13_166 k_13_166(i_13_235, i_13_238, i_13_414, i_13_415, i_13_416, i_13_432, i_13_446, i_13_507, i_13_523, i_13_526, i_13_535, i_13_562, i_13_568, i_13_694, i_13_797, i_13_823, i_13_841, i_13_842, i_13_946, i_13_1018, i_13_1073, i_13_1076, i_13_1129, i_13_1132, i_13_1190, i_13_1193, i_13_1214, i_13_1228, i_13_1252, i_13_1256, i_13_1268, i_13_1400, i_13_1411, i_13_1531, i_13_1548, i_13_1549, i_13_1550, i_13_1552, i_13_1553, i_13_1603, i_13_1696, i_13_1846, i_13_1934, i_13_1957, i_13_1958, i_13_2043, i_13_2109, i_13_2203, i_13_2289, i_13_2334, i_13_2380, i_13_2449, i_13_2539, i_13_2555, i_13_2611, i_13_2713, i_13_2754, i_13_2900, i_13_3010, i_13_3013, i_13_3014, i_13_3064, i_13_3065, i_13_3070, i_13_3101, i_13_3172, i_13_3272, i_13_3382, i_13_3416, i_13_3451, i_13_3461, i_13_3484, i_13_3487, i_13_3488, i_13_3523, i_13_3537, i_13_3538, i_13_3539, i_13_3541, i_13_3542, i_13_3544, i_13_3545, i_13_3686, i_13_3730, i_13_3766, i_13_3852, i_13_3856, i_13_3857, i_13_3880, i_13_3895, i_13_3908, i_13_3915, i_13_3916, i_13_4252, i_13_4256, i_13_4369, i_13_4378, i_13_4379, i_13_4382, i_13_4536, o_13_166);
	kernel_13_167 k_13_167(i_13_80, i_13_139, i_13_232, i_13_283, i_13_332, i_13_358, i_13_376, i_13_428, i_13_447, i_13_457, i_13_538, i_13_599, i_13_607, i_13_646, i_13_647, i_13_688, i_13_689, i_13_691, i_13_692, i_13_718, i_13_728, i_13_940, i_13_979, i_13_1120, i_13_1204, i_13_1263, i_13_1275, i_13_1276, i_13_1277, i_13_1348, i_13_1393, i_13_1484, i_13_1493, i_13_1570, i_13_1642, i_13_1645, i_13_1646, i_13_1672, i_13_1673, i_13_1691, i_13_1713, i_13_1723, i_13_1726, i_13_1727, i_13_1741, i_13_1780, i_13_1781, i_13_1885, i_13_1888, i_13_1933, i_13_1996, i_13_2113, i_13_2137, i_13_2150, i_13_2191, i_13_2194, i_13_2282, i_13_2379, i_13_2383, i_13_2533, i_13_2542, i_13_2552, i_13_2617, i_13_2649, i_13_2650, i_13_2651, i_13_2653, i_13_2654, i_13_2661, i_13_2671, i_13_2690, i_13_2742, i_13_2751, i_13_2847, i_13_2848, i_13_2851, i_13_2852, i_13_2875, i_13_2878, i_13_3139, i_13_3392, i_13_3535, i_13_3581, i_13_3760, i_13_3797, i_13_3874, i_13_3995, i_13_4045, i_13_4162, i_13_4190, i_13_4193, i_13_4219, i_13_4234, i_13_4354, i_13_4377, i_13_4423, i_13_4432, i_13_4444, i_13_4597, i_13_4598, o_13_167);
	kernel_13_168 k_13_168(i_13_52, i_13_116, i_13_167, i_13_185, i_13_199, i_13_251, i_13_286, i_13_287, i_13_418, i_13_441, i_13_517, i_13_556, i_13_559, i_13_576, i_13_619, i_13_620, i_13_655, i_13_675, i_13_715, i_13_928, i_13_929, i_13_944, i_13_1018, i_13_1085, i_13_1098, i_13_1310, i_13_1364, i_13_1397, i_13_1426, i_13_1471, i_13_1498, i_13_1501, i_13_1502, i_13_1505, i_13_1606, i_13_1609, i_13_1633, i_13_1634, i_13_1636, i_13_1637, i_13_1731, i_13_1735, i_13_1754, i_13_1917, i_13_1949, i_13_2171, i_13_2276, i_13_2342, i_13_2369, i_13_2455, i_13_2492, i_13_2545, i_13_2581, i_13_2673, i_13_2708, i_13_2714, i_13_2753, i_13_2788, i_13_2888, i_13_2922, i_13_2923, i_13_2956, i_13_2959, i_13_3130, i_13_3145, i_13_3146, i_13_3149, i_13_3253, i_13_3373, i_13_3409, i_13_3418, i_13_3419, i_13_3447, i_13_3464, i_13_3486, i_13_3581, i_13_3599, i_13_3647, i_13_3650, i_13_3724, i_13_3734, i_13_3765, i_13_3770, i_13_3787, i_13_3816, i_13_3904, i_13_3905, i_13_4015, i_13_4019, i_13_4077, i_13_4087, i_13_4088, i_13_4253, i_13_4255, i_13_4256, i_13_4391, i_13_4531, i_13_4562, i_13_4567, i_13_4590, o_13_168);
	kernel_13_169 k_13_169(i_13_112, i_13_136, i_13_158, i_13_163, i_13_226, i_13_229, i_13_336, i_13_380, i_13_382, i_13_418, i_13_445, i_13_453, i_13_517, i_13_569, i_13_571, i_13_577, i_13_596, i_13_614, i_13_641, i_13_652, i_13_686, i_13_715, i_13_733, i_13_778, i_13_779, i_13_841, i_13_873, i_13_1101, i_13_1300, i_13_1327, i_13_1444, i_13_1462, i_13_1503, i_13_1517, i_13_1521, i_13_1625, i_13_1711, i_13_1713, i_13_1720, i_13_1721, i_13_1730, i_13_1783, i_13_1786, i_13_1787, i_13_1802, i_13_1811, i_13_1882, i_13_1884, i_13_1999, i_13_2018, i_13_2097, i_13_2120, i_13_2170, i_13_2192, i_13_2210, i_13_2260, i_13_2425, i_13_2458, i_13_2541, i_13_2647, i_13_2712, i_13_2722, i_13_2845, i_13_2935, i_13_2939, i_13_3015, i_13_3020, i_13_3033, i_13_3034, i_13_3036, i_13_3037, i_13_3124, i_13_3142, i_13_3143, i_13_3164, i_13_3213, i_13_3270, i_13_3290, i_13_3421, i_13_3422, i_13_3424, i_13_3425, i_13_3430, i_13_3449, i_13_3547, i_13_3568, i_13_3791, i_13_3862, i_13_3865, i_13_3983, i_13_4009, i_13_4010, i_13_4015, i_13_4016, i_13_4054, i_13_4086, i_13_4234, i_13_4306, i_13_4311, i_13_4369, o_13_169);
	kernel_13_170 k_13_170(i_13_48, i_13_136, i_13_144, i_13_211, i_13_229, i_13_271, i_13_283, i_13_300, i_13_382, i_13_517, i_13_571, i_13_585, i_13_639, i_13_705, i_13_711, i_13_738, i_13_796, i_13_940, i_13_999, i_13_1044, i_13_1101, i_13_1344, i_13_1377, i_13_1390, i_13_1399, i_13_1408, i_13_1432, i_13_1513, i_13_1632, i_13_1633, i_13_1639, i_13_1768, i_13_1776, i_13_1795, i_13_1848, i_13_1893, i_13_1936, i_13_1945, i_13_2029, i_13_2030, i_13_2053, i_13_2250, i_13_2251, i_13_2253, i_13_2278, i_13_2413, i_13_2424, i_13_2433, i_13_2497, i_13_2515, i_13_2542, i_13_2547, i_13_2614, i_13_2668, i_13_2674, i_13_2712, i_13_2713, i_13_2755, i_13_2953, i_13_2980, i_13_3051, i_13_3123, i_13_3235, i_13_3250, i_13_3334, i_13_3352, i_13_3487, i_13_3574, i_13_3592, i_13_3595, i_13_3684, i_13_3700, i_13_3729, i_13_3730, i_13_3816, i_13_3856, i_13_3901, i_13_3927, i_13_3928, i_13_3982, i_13_4009, i_13_4018, i_13_4045, i_13_4054, i_13_4081, i_13_4090, i_13_4096, i_13_4189, i_13_4215, i_13_4230, i_13_4234, i_13_4251, i_13_4252, i_13_4267, i_13_4296, i_13_4297, i_13_4405, i_13_4432, i_13_4558, i_13_4590, o_13_170);
	kernel_13_171 k_13_171(i_13_48, i_13_63, i_13_64, i_13_71, i_13_158, i_13_172, i_13_176, i_13_207, i_13_209, i_13_227, i_13_245, i_13_256, i_13_304, i_13_415, i_13_526, i_13_605, i_13_612, i_13_613, i_13_616, i_13_764, i_13_828, i_13_838, i_13_854, i_13_1075, i_13_1132, i_13_1227, i_13_1304, i_13_1305, i_13_1309, i_13_1360, i_13_1441, i_13_1443, i_13_1495, i_13_1521, i_13_1522, i_13_1523, i_13_1525, i_13_1548, i_13_1549, i_13_1593, i_13_1604, i_13_1638, i_13_1639, i_13_1696, i_13_1721, i_13_1728, i_13_1730, i_13_1799, i_13_1846, i_13_1926, i_13_1930, i_13_1931, i_13_2142, i_13_2182, i_13_2199, i_13_2243, i_13_2297, i_13_2407, i_13_2421, i_13_2430, i_13_2505, i_13_2554, i_13_2673, i_13_2675, i_13_2722, i_13_2748, i_13_2881, i_13_2883, i_13_3240, i_13_3241, i_13_3288, i_13_3367, i_13_3395, i_13_3414, i_13_3420, i_13_3538, i_13_3539, i_13_3548, i_13_3636, i_13_3637, i_13_3638, i_13_3640, i_13_3758, i_13_3766, i_13_3843, i_13_3845, i_13_3889, i_13_3898, i_13_3913, i_13_3916, i_13_3934, i_13_4217, i_13_4312, i_13_4322, i_13_4472, i_13_4509, i_13_4511, i_13_4522, i_13_4590, i_13_4607, o_13_171);
	kernel_13_172 k_13_172(i_13_35, i_13_52, i_13_69, i_13_70, i_13_71, i_13_78, i_13_90, i_13_127, i_13_314, i_13_402, i_13_449, i_13_537, i_13_565, i_13_641, i_13_673, i_13_679, i_13_737, i_13_763, i_13_823, i_13_843, i_13_933, i_13_1021, i_13_1101, i_13_1102, i_13_1105, i_13_1106, i_13_1151, i_13_1228, i_13_1263, i_13_1276, i_13_1345, i_13_1363, i_13_1401, i_13_1402, i_13_1519, i_13_1599, i_13_1627, i_13_1644, i_13_1725, i_13_1726, i_13_1777, i_13_1780, i_13_1781, i_13_1797, i_13_1799, i_13_1827, i_13_1853, i_13_1858, i_13_1925, i_13_1948, i_13_1995, i_13_2054, i_13_2176, i_13_2208, i_13_2312, i_13_2617, i_13_2638, i_13_2695, i_13_2698, i_13_2715, i_13_2725, i_13_2752, i_13_2760, i_13_2770, i_13_2851, i_13_2878, i_13_2901, i_13_2905, i_13_3039, i_13_3067, i_13_3128, i_13_3367, i_13_3370, i_13_3417, i_13_3418, i_13_3441, i_13_3534, i_13_3580, i_13_3595, i_13_3640, i_13_3648, i_13_3684, i_13_3685, i_13_3739, i_13_3757, i_13_3767, i_13_3787, i_13_3796, i_13_3869, i_13_3895, i_13_3913, i_13_3928, i_13_3931, i_13_3991, i_13_3994, i_13_4264, i_13_4335, i_13_4434, i_13_4450, i_13_4451, o_13_172);
	kernel_13_173 k_13_173(i_13_41, i_13_74, i_13_104, i_13_109, i_13_110, i_13_280, i_13_283, i_13_320, i_13_406, i_13_452, i_13_506, i_13_553, i_13_581, i_13_599, i_13_604, i_13_622, i_13_677, i_13_680, i_13_794, i_13_856, i_13_859, i_13_946, i_13_947, i_13_1019, i_13_1022, i_13_1084, i_13_1282, i_13_1424, i_13_1436, i_13_1444, i_13_1472, i_13_1486, i_13_1487, i_13_1543, i_13_1553, i_13_1621, i_13_1630, i_13_1670, i_13_1838, i_13_1841, i_13_1856, i_13_1927, i_13_1999, i_13_2047, i_13_2053, i_13_2146, i_13_2263, i_13_2314, i_13_2396, i_13_2432, i_13_2435, i_13_2458, i_13_2459, i_13_2462, i_13_2501, i_13_2503, i_13_2504, i_13_2506, i_13_2507, i_13_2521, i_13_2529, i_13_2539, i_13_2540, i_13_2611, i_13_2612, i_13_2714, i_13_2746, i_13_2911, i_13_2920, i_13_3071, i_13_3124, i_13_3143, i_13_3145, i_13_3146, i_13_3154, i_13_3340, i_13_3422, i_13_3523, i_13_3529, i_13_3530, i_13_3542, i_13_3577, i_13_3661, i_13_3757, i_13_3844, i_13_3871, i_13_3889, i_13_3890, i_13_3928, i_13_4046, i_13_4063, i_13_4223, i_13_4252, i_13_4253, i_13_4325, i_13_4366, i_13_4424, i_13_4519, i_13_4520, i_13_4556, o_13_173);
	kernel_13_174 k_13_174(i_13_67, i_13_106, i_13_123, i_13_138, i_13_139, i_13_161, i_13_166, i_13_232, i_13_247, i_13_310, i_13_327, i_13_328, i_13_430, i_13_526, i_13_537, i_13_571, i_13_598, i_13_670, i_13_717, i_13_780, i_13_825, i_13_832, i_13_841, i_13_861, i_13_890, i_13_894, i_13_1023, i_13_1024, i_13_1095, i_13_1096, i_13_1111, i_13_1281, i_13_1299, i_13_1303, i_13_1326, i_13_1464, i_13_1488, i_13_1489, i_13_1490, i_13_1515, i_13_1777, i_13_1785, i_13_1786, i_13_1788, i_13_1857, i_13_1858, i_13_1884, i_13_1887, i_13_1930, i_13_2056, i_13_2146, i_13_2175, i_13_2190, i_13_2263, i_13_2309, i_13_2310, i_13_2311, i_13_2316, i_13_2460, i_13_2461, i_13_2462, i_13_2464, i_13_2500, i_13_2506, i_13_2532, i_13_2565, i_13_2566, i_13_2613, i_13_2632, i_13_2885, i_13_2941, i_13_3087, i_13_3148, i_13_3171, i_13_3173, i_13_3174, i_13_3348, i_13_3432, i_13_3481, i_13_3532, i_13_3534, i_13_3535, i_13_3661, i_13_3732, i_13_3741, i_13_3783, i_13_3797, i_13_3820, i_13_3913, i_13_3923, i_13_3932, i_13_4012, i_13_4210, i_13_4237, i_13_4341, i_13_4443, i_13_4514, i_13_4521, i_13_4522, i_13_4567, o_13_174);
	kernel_13_175 k_13_175(i_13_76, i_13_77, i_13_88, i_13_94, i_13_130, i_13_134, i_13_256, i_13_269, i_13_332, i_13_358, i_13_359, i_13_370, i_13_371, i_13_400, i_13_458, i_13_520, i_13_571, i_13_611, i_13_617, i_13_667, i_13_671, i_13_823, i_13_842, i_13_980, i_13_1091, i_13_1115, i_13_1213, i_13_1282, i_13_1348, i_13_1400, i_13_1402, i_13_1403, i_13_1508, i_13_1519, i_13_1660, i_13_1750, i_13_1763, i_13_1778, i_13_1951, i_13_1952, i_13_2032, i_13_2033, i_13_2059, i_13_2060, i_13_2141, i_13_2191, i_13_2203, i_13_2240, i_13_2284, i_13_2285, i_13_2321, i_13_2348, i_13_2408, i_13_2410, i_13_2447, i_13_2497, i_13_2503, i_13_2510, i_13_2515, i_13_2516, i_13_2555, i_13_2590, i_13_2696, i_13_2705, i_13_2902, i_13_2920, i_13_2923, i_13_2924, i_13_2959, i_13_3013, i_13_3073, i_13_3218, i_13_3373, i_13_3374, i_13_3419, i_13_3580, i_13_3581, i_13_3598, i_13_3599, i_13_3622, i_13_3623, i_13_3634, i_13_3635, i_13_3784, i_13_3788, i_13_3988, i_13_3991, i_13_4076, i_13_4190, i_13_4208, i_13_4216, i_13_4237, i_13_4264, i_13_4265, i_13_4333, i_13_4334, i_13_4378, i_13_4433, i_13_4453, i_13_4454, o_13_175);
	kernel_13_176 k_13_176(i_13_68, i_13_94, i_13_112, i_13_139, i_13_140, i_13_237, i_13_320, i_13_380, i_13_445, i_13_524, i_13_553, i_13_586, i_13_587, i_13_607, i_13_614, i_13_686, i_13_696, i_13_698, i_13_739, i_13_796, i_13_883, i_13_1075, i_13_1103, i_13_1117, i_13_1208, i_13_1268, i_13_1273, i_13_1274, i_13_1298, i_13_1342, i_13_1343, i_13_1400, i_13_1441, i_13_1442, i_13_1468, i_13_1507, i_13_1516, i_13_1568, i_13_1598, i_13_1712, i_13_1775, i_13_1778, i_13_1810, i_13_1811, i_13_1921, i_13_1928, i_13_1945, i_13_1990, i_13_1991, i_13_2053, i_13_2054, i_13_2189, i_13_2197, i_13_2236, i_13_2260, i_13_2278, i_13_2279, i_13_2320, i_13_2377, i_13_2503, i_13_2593, i_13_2647, i_13_2675, i_13_2696, i_13_2710, i_13_2720, i_13_2723, i_13_2782, i_13_2899, i_13_2921, i_13_2998, i_13_3001, i_13_3058, i_13_3059, i_13_3061, i_13_3064, i_13_3065, i_13_3136, i_13_3208, i_13_3367, i_13_3368, i_13_3386, i_13_3415, i_13_3439, i_13_3593, i_13_3650, i_13_3856, i_13_4096, i_13_4187, i_13_4231, i_13_4258, i_13_4259, i_13_4268, i_13_4339, i_13_4393, i_13_4394, i_13_4405, i_13_4429, i_13_4447, i_13_4448, o_13_176);
	kernel_13_177 k_13_177(i_13_52, i_13_73, i_13_76, i_13_121, i_13_158, i_13_205, i_13_259, i_13_275, i_13_277, i_13_310, i_13_355, i_13_450, i_13_451, i_13_452, i_13_454, i_13_661, i_13_665, i_13_674, i_13_716, i_13_874, i_13_929, i_13_952, i_13_1063, i_13_1139, i_13_1151, i_13_1228, i_13_1229, i_13_1256, i_13_1258, i_13_1408, i_13_1411, i_13_1412, i_13_1469, i_13_1516, i_13_1528, i_13_1679, i_13_1681, i_13_1732, i_13_1736, i_13_1768, i_13_1769, i_13_1781, i_13_1805, i_13_1895, i_13_2021, i_13_2056, i_13_2111, i_13_2149, i_13_2284, i_13_2299, i_13_2300, i_13_2354, i_13_2572, i_13_2596, i_13_2597, i_13_2614, i_13_2615, i_13_2617, i_13_2665, i_13_2708, i_13_2782, i_13_2891, i_13_2900, i_13_2983, i_13_2987, i_13_3029, i_13_3032, i_13_3114, i_13_3130, i_13_3157, i_13_3215, i_13_3218, i_13_3287, i_13_3313, i_13_3355, i_13_3461, i_13_3467, i_13_3488, i_13_3521, i_13_3598, i_13_3687, i_13_3730, i_13_3757, i_13_3784, i_13_3875, i_13_3979, i_13_4055, i_13_4073, i_13_4088, i_13_4102, i_13_4162, i_13_4163, i_13_4228, i_13_4237, i_13_4268, i_13_4372, i_13_4448, i_13_4517, i_13_4559, i_13_4607, o_13_177);
	kernel_13_178 k_13_178(i_13_40, i_13_109, i_13_113, i_13_116, i_13_129, i_13_162, i_13_286, i_13_322, i_13_325, i_13_535, i_13_571, i_13_687, i_13_691, i_13_855, i_13_946, i_13_1012, i_13_1080, i_13_1081, i_13_1087, i_13_1120, i_13_1220, i_13_1395, i_13_1423, i_13_1424, i_13_1494, i_13_1569, i_13_1574, i_13_1629, i_13_1630, i_13_1632, i_13_1633, i_13_1634, i_13_1637, i_13_1773, i_13_1795, i_13_1938, i_13_1998, i_13_2059, i_13_2080, i_13_2081, i_13_2237, i_13_2342, i_13_2433, i_13_2438, i_13_2452, i_13_2462, i_13_2464, i_13_2498, i_13_2539, i_13_2541, i_13_2545, i_13_2546, i_13_2716, i_13_2905, i_13_2917, i_13_2920, i_13_2921, i_13_2955, i_13_3064, i_13_3065, i_13_3141, i_13_3143, i_13_3145, i_13_3146, i_13_3148, i_13_3338, i_13_3454, i_13_3455, i_13_3463, i_13_3464, i_13_3466, i_13_3688, i_13_3689, i_13_3727, i_13_3730, i_13_3734, i_13_3767, i_13_3770, i_13_3919, i_13_3968, i_13_3995, i_13_4018, i_13_4021, i_13_4022, i_13_4036, i_13_4049, i_13_4091, i_13_4253, i_13_4255, i_13_4256, i_13_4309, i_13_4354, i_13_4469, i_13_4513, i_13_4522, i_13_4523, i_13_4526, i_13_4558, i_13_4561, i_13_4562, o_13_178);
	kernel_13_179 k_13_179(i_13_31, i_13_79, i_13_111, i_13_112, i_13_114, i_13_166, i_13_168, i_13_169, i_13_229, i_13_318, i_13_327, i_13_490, i_13_525, i_13_526, i_13_564, i_13_643, i_13_822, i_13_850, i_13_858, i_13_862, i_13_924, i_13_940, i_13_960, i_13_1021, i_13_1075, i_13_1077, i_13_1200, i_13_1281, i_13_1419, i_13_1426, i_13_1428, i_13_1488, i_13_1498, i_13_1552, i_13_1632, i_13_1633, i_13_1642, i_13_1645, i_13_1704, i_13_1731, i_13_1831, i_13_1843, i_13_1950, i_13_1957, i_13_1986, i_13_2004, i_13_2026, i_13_2029, i_13_2193, i_13_2211, i_13_2271, i_13_2370, i_13_2452, i_13_2454, i_13_2455, i_13_2463, i_13_2541, i_13_2613, i_13_2707, i_13_2766, i_13_2778, i_13_2919, i_13_2920, i_13_2973, i_13_3030, i_13_3037, i_13_3090, i_13_3117, i_13_3148, i_13_3172, i_13_3180, i_13_3414, i_13_3453, i_13_3454, i_13_3459, i_13_3460, i_13_3462, i_13_3481, i_13_3483, i_13_3505, i_13_3540, i_13_3541, i_13_3561, i_13_3567, i_13_3574, i_13_3721, i_13_3867, i_13_3892, i_13_3936, i_13_4018, i_13_4063, i_13_4071, i_13_4164, i_13_4251, i_13_4255, i_13_4324, i_13_4341, i_13_4372, i_13_4378, i_13_4558, o_13_179);
	kernel_13_180 k_13_180(i_13_49, i_13_50, i_13_104, i_13_164, i_13_268, i_13_308, i_13_316, i_13_317, i_13_334, i_13_373, i_13_374, i_13_376, i_13_445, i_13_533, i_13_551, i_13_605, i_13_641, i_13_652, i_13_668, i_13_676, i_13_677, i_13_689, i_13_698, i_13_757, i_13_772, i_13_896, i_13_982, i_13_983, i_13_1121, i_13_1148, i_13_1250, i_13_1348, i_13_1412, i_13_1442, i_13_1516, i_13_1573, i_13_1648, i_13_1721, i_13_1750, i_13_1760, i_13_1789, i_13_1814, i_13_1832, i_13_1885, i_13_1909, i_13_1934, i_13_1957, i_13_2018, i_13_2032, i_13_2053, i_13_2113, i_13_2170, i_13_2281, i_13_2320, i_13_2348, i_13_2363, i_13_2468, i_13_2506, i_13_2507, i_13_2555, i_13_2716, i_13_2999, i_13_3047, i_13_3139, i_13_3215, i_13_3328, i_13_3352, i_13_3370, i_13_3376, i_13_3433, i_13_3437, i_13_3524, i_13_3533, i_13_3541, i_13_3565, i_13_3646, i_13_3686, i_13_3767, i_13_3865, i_13_3889, i_13_3890, i_13_3983, i_13_3988, i_13_4018, i_13_4019, i_13_4033, i_13_4046, i_13_4048, i_13_4079, i_13_4121, i_13_4124, i_13_4178, i_13_4447, i_13_4459, i_13_4471, i_13_4544, i_13_4591, i_13_4592, i_13_4600, i_13_4601, o_13_180);
	kernel_13_181 k_13_181(i_13_76, i_13_93, i_13_117, i_13_180, i_13_181, i_13_226, i_13_228, i_13_394, i_13_517, i_13_534, i_13_594, i_13_680, i_13_696, i_13_711, i_13_728, i_13_732, i_13_737, i_13_861, i_13_894, i_13_1075, i_13_1121, i_13_1207, i_13_1209, i_13_1252, i_13_1299, i_13_1408, i_13_1495, i_13_1507, i_13_1602, i_13_1632, i_13_1640, i_13_1700, i_13_1721, i_13_1723, i_13_1747, i_13_1782, i_13_1783, i_13_1785, i_13_1786, i_13_1921, i_13_1949, i_13_1955, i_13_1991, i_13_2055, i_13_2056, i_13_2096, i_13_2119, i_13_2182, i_13_2201, i_13_2204, i_13_2205, i_13_2208, i_13_2209, i_13_2235, i_13_2361, i_13_2452, i_13_2465, i_13_2560, i_13_2641, i_13_2789, i_13_2938, i_13_3019, i_13_3037, i_13_3062, i_13_3162, i_13_3163, i_13_3176, i_13_3204, i_13_3213, i_13_3285, i_13_3289, i_13_3353, i_13_3420, i_13_3423, i_13_3424, i_13_3531, i_13_3596, i_13_3620, i_13_3766, i_13_3782, i_13_3794, i_13_3870, i_13_3871, i_13_3981, i_13_4006, i_13_4008, i_13_4014, i_13_4022, i_13_4050, i_13_4058, i_13_4184, i_13_4214, i_13_4238, i_13_4261, i_13_4302, i_13_4397, i_13_4413, i_13_4451, i_13_4518, i_13_4540, o_13_181);
	kernel_13_182 k_13_182(i_13_45, i_13_48, i_13_76, i_13_94, i_13_247, i_13_411, i_13_450, i_13_534, i_13_556, i_13_601, i_13_625, i_13_626, i_13_660, i_13_661, i_13_812, i_13_834, i_13_835, i_13_850, i_13_909, i_13_940, i_13_1075, i_13_1147, i_13_1204, i_13_1227, i_13_1228, i_13_1230, i_13_1255, i_13_1271, i_13_1305, i_13_1314, i_13_1329, i_13_1345, i_13_1404, i_13_1463, i_13_1480, i_13_1497, i_13_1515, i_13_1522, i_13_1551, i_13_1647, i_13_1732, i_13_1744, i_13_1757, i_13_1767, i_13_1768, i_13_1803, i_13_1804, i_13_1884, i_13_1885, i_13_1944, i_13_1954, i_13_2001, i_13_2002, i_13_2100, i_13_2135, i_13_2145, i_13_2148, i_13_2199, i_13_2244, i_13_2469, i_13_2470, i_13_2472, i_13_2571, i_13_2625, i_13_2679, i_13_2854, i_13_2857, i_13_2896, i_13_2911, i_13_2968, i_13_2982, i_13_2985, i_13_3013, i_13_3031, i_13_3145, i_13_3258, i_13_3399, i_13_3423, i_13_3486, i_13_3549, i_13_3739, i_13_3803, i_13_3819, i_13_3850, i_13_3864, i_13_3868, i_13_3981, i_13_4126, i_13_4164, i_13_4252, i_13_4267, i_13_4269, i_13_4295, i_13_4369, i_13_4455, i_13_4467, i_13_4512, i_13_4513, i_13_4539, i_13_4566, o_13_182);
	kernel_13_183 k_13_183(i_13_39, i_13_40, i_13_46, i_13_154, i_13_156, i_13_229, i_13_238, i_13_274, i_13_275, i_13_280, i_13_306, i_13_310, i_13_311, i_13_319, i_13_335, i_13_351, i_13_362, i_13_409, i_13_451, i_13_452, i_13_517, i_13_567, i_13_568, i_13_644, i_13_739, i_13_837, i_13_928, i_13_929, i_13_937, i_13_1082, i_13_1368, i_13_1432, i_13_1469, i_13_1496, i_13_1661, i_13_1765, i_13_1766, i_13_1829, i_13_1892, i_13_1945, i_13_2098, i_13_2227, i_13_2233, i_13_2234, i_13_2297, i_13_2434, i_13_2452, i_13_2542, i_13_2650, i_13_2677, i_13_2744, i_13_2746, i_13_2765, i_13_2767, i_13_2875, i_13_2981, i_13_3017, i_13_3029, i_13_3056, i_13_3107, i_13_3164, i_13_3214, i_13_3218, i_13_3232, i_13_3235, i_13_3286, i_13_3312, i_13_3313, i_13_3485, i_13_3487, i_13_3488, i_13_3523, i_13_3684, i_13_3698, i_13_3764, i_13_3766, i_13_3869, i_13_3898, i_13_3899, i_13_3901, i_13_4041, i_13_4063, i_13_4087, i_13_4088, i_13_4159, i_13_4162, i_13_4231, i_13_4250, i_13_4253, i_13_4267, i_13_4268, i_13_4270, i_13_4325, i_13_4359, i_13_4369, i_13_4370, i_13_4392, i_13_4447, i_13_4448, i_13_4559, o_13_183);
	kernel_13_184 k_13_184(i_13_19, i_13_40, i_13_55, i_13_73, i_13_94, i_13_103, i_13_157, i_13_211, i_13_280, i_13_425, i_13_451, i_13_463, i_13_524, i_13_586, i_13_697, i_13_715, i_13_824, i_13_868, i_13_928, i_13_1017, i_13_1021, i_13_1066, i_13_1075, i_13_1204, i_13_1205, i_13_1207, i_13_1228, i_13_1274, i_13_1297, i_13_1342, i_13_1343, i_13_1405, i_13_1426, i_13_1427, i_13_1435, i_13_1468, i_13_1568, i_13_1634, i_13_1642, i_13_1711, i_13_1777, i_13_1811, i_13_1831, i_13_1882, i_13_1918, i_13_1940, i_13_1990, i_13_2004, i_13_2053, i_13_2110, i_13_2197, i_13_2236, i_13_2311, i_13_2362, i_13_2376, i_13_2452, i_13_2453, i_13_2504, i_13_2542, i_13_2549, i_13_2615, i_13_2710, i_13_2749, i_13_2854, i_13_2855, i_13_2912, i_13_2917, i_13_2918, i_13_3142, i_13_3143, i_13_3163, i_13_3208, i_13_3343, i_13_3441, i_13_3460, i_13_3467, i_13_3502, i_13_3503, i_13_3576, i_13_3637, i_13_3646, i_13_3764, i_13_3966, i_13_3982, i_13_4087, i_13_4088, i_13_4231, i_13_4258, i_13_4259, i_13_4392, i_13_4393, i_13_4394, i_13_4446, i_13_4447, i_13_4448, i_13_4511, i_13_4513, i_13_4555, i_13_4559, i_13_4564, o_13_184);
	kernel_13_185 k_13_185(i_13_27, i_13_49, i_13_64, i_13_67, i_13_120, i_13_121, i_13_192, i_13_193, i_13_201, i_13_225, i_13_270, i_13_324, i_13_378, i_13_379, i_13_441, i_13_507, i_13_553, i_13_570, i_13_571, i_13_576, i_13_694, i_13_697, i_13_714, i_13_715, i_13_717, i_13_768, i_13_858, i_13_948, i_13_1120, i_13_1200, i_13_1228, i_13_1372, i_13_1407, i_13_1426, i_13_1443, i_13_1467, i_13_1507, i_13_1516, i_13_1552, i_13_1623, i_13_1782, i_13_1783, i_13_1800, i_13_1801, i_13_1990, i_13_2011, i_13_2055, i_13_2056, i_13_2116, i_13_2128, i_13_2134, i_13_2206, i_13_2208, i_13_2209, i_13_2260, i_13_2358, i_13_2404, i_13_2424, i_13_2430, i_13_2452, i_13_2532, i_13_2589, i_13_2593, i_13_2710, i_13_2718, i_13_2934, i_13_2935, i_13_3015, i_13_3016, i_13_3151, i_13_3171, i_13_3208, i_13_3214, i_13_3241, i_13_3258, i_13_3267, i_13_3286, i_13_3342, i_13_3415, i_13_3420, i_13_3421, i_13_3423, i_13_3424, i_13_3532, i_13_3610, i_13_3846, i_13_3847, i_13_3871, i_13_3873, i_13_3874, i_13_3981, i_13_4009, i_13_4050, i_13_4051, i_13_4123, i_13_4150, i_13_4188, i_13_4404, i_13_4410, i_13_4594, o_13_185);
	kernel_13_186 k_13_186(i_13_78, i_13_96, i_13_106, i_13_327, i_13_529, i_13_598, i_13_627, i_13_672, i_13_673, i_13_717, i_13_727, i_13_780, i_13_781, i_13_815, i_13_825, i_13_841, i_13_850, i_13_894, i_13_949, i_13_979, i_13_1095, i_13_1141, i_13_1259, i_13_1302, i_13_1303, i_13_1320, i_13_1327, i_13_1383, i_13_1464, i_13_1465, i_13_1466, i_13_1482, i_13_1483, i_13_1484, i_13_1643, i_13_1751, i_13_1759, i_13_1789, i_13_1806, i_13_1807, i_13_1808, i_13_1815, i_13_1885, i_13_1887, i_13_1905, i_13_1906, i_13_2033, i_13_2122, i_13_2123, i_13_2139, i_13_2140, i_13_2167, i_13_2177, i_13_2247, i_13_2310, i_13_2380, i_13_2445, i_13_2446, i_13_2470, i_13_2474, i_13_2652, i_13_2698, i_13_2751, i_13_2823, i_13_2824, i_13_2861, i_13_3009, i_13_3112, i_13_3174, i_13_3219, i_13_3220, i_13_3293, i_13_3391, i_13_3398, i_13_3432, i_13_3451, i_13_3452, i_13_3564, i_13_3577, i_13_3579, i_13_3734, i_13_3793, i_13_3820, i_13_3855, i_13_3874, i_13_3883, i_13_3927, i_13_3929, i_13_3991, i_13_3992, i_13_4049, i_13_4237, i_13_4308, i_13_4318, i_13_4365, i_13_4380, i_13_4414, i_13_4443, i_13_4453, i_13_4521, o_13_186);
	kernel_13_187 k_13_187(i_13_31, i_13_101, i_13_235, i_13_238, i_13_248, i_13_251, i_13_256, i_13_263, i_13_275, i_13_278, i_13_338, i_13_407, i_13_411, i_13_447, i_13_451, i_13_485, i_13_535, i_13_559, i_13_563, i_13_577, i_13_578, i_13_616, i_13_619, i_13_620, i_13_644, i_13_793, i_13_813, i_13_832, i_13_841, i_13_941, i_13_942, i_13_977, i_13_979, i_13_1095, i_13_1112, i_13_1262, i_13_1333, i_13_1342, i_13_1396, i_13_1397, i_13_1477, i_13_1494, i_13_1541, i_13_1570, i_13_1647, i_13_1658, i_13_1722, i_13_1729, i_13_1814, i_13_1835, i_13_1842, i_13_1858, i_13_1920, i_13_1947, i_13_2106, i_13_2108, i_13_2113, i_13_2230, i_13_2233, i_13_2261, i_13_2280, i_13_2445, i_13_2713, i_13_2721, i_13_2737, i_13_2740, i_13_2765, i_13_2785, i_13_2888, i_13_2951, i_13_3018, i_13_3056, i_13_3115, i_13_3135, i_13_3152, i_13_3208, i_13_3217, i_13_3218, i_13_3313, i_13_3316, i_13_3403, i_13_3412, i_13_3435, i_13_3461, i_13_3601, i_13_3602, i_13_3616, i_13_3617, i_13_3709, i_13_3764, i_13_3858, i_13_3901, i_13_3902, i_13_4124, i_13_4178, i_13_4207, i_13_4268, i_13_4360, i_13_4391, i_13_4483, o_13_187);
	kernel_13_188 k_13_188(i_13_44, i_13_91, i_13_98, i_13_175, i_13_176, i_13_179, i_13_181, i_13_229, i_13_280, i_13_283, i_13_308, i_13_309, i_13_313, i_13_314, i_13_317, i_13_320, i_13_549, i_13_554, i_13_571, i_13_657, i_13_697, i_13_710, i_13_758, i_13_846, i_13_847, i_13_855, i_13_981, i_13_985, i_13_986, i_13_1105, i_13_1106, i_13_1260, i_13_1327, i_13_1471, i_13_1486, i_13_1511, i_13_1532, i_13_1714, i_13_1799, i_13_1832, i_13_1852, i_13_1853, i_13_1858, i_13_1859, i_13_1861, i_13_1996, i_13_2096, i_13_2406, i_13_2411, i_13_2447, i_13_2452, i_13_2460, i_13_2473, i_13_2475, i_13_2565, i_13_2676, i_13_2699, i_13_2798, i_13_2849, i_13_2983, i_13_3006, i_13_3008, i_13_3009, i_13_3032, i_13_3061, i_13_3108, i_13_3109, i_13_3112, i_13_3141, i_13_3204, i_13_3205, i_13_3208, i_13_3211, i_13_3212, i_13_3335, i_13_3343, i_13_3382, i_13_3397, i_13_3405, i_13_3765, i_13_3766, i_13_3816, i_13_3817, i_13_3818, i_13_3823, i_13_3865, i_13_3866, i_13_3910, i_13_4043, i_13_4063, i_13_4067, i_13_4084, i_13_4085, i_13_4304, i_13_4350, i_13_4379, i_13_4414, i_13_4522, i_13_4581, i_13_4598, o_13_188);
	kernel_13_189 k_13_189(i_13_29, i_13_36, i_13_37, i_13_46, i_13_64, i_13_121, i_13_136, i_13_311, i_13_334, i_13_370, i_13_412, i_13_414, i_13_415, i_13_585, i_13_612, i_13_613, i_13_654, i_13_684, i_13_685, i_13_693, i_13_694, i_13_760, i_13_837, i_13_838, i_13_841, i_13_889, i_13_955, i_13_1071, i_13_1072, i_13_1081, i_13_1117, i_13_1121, i_13_1270, i_13_1285, i_13_1299, i_13_1317, i_13_1360, i_13_1390, i_13_1516, i_13_1521, i_13_1522, i_13_1534, i_13_1633, i_13_1639, i_13_1668, i_13_1750, i_13_1756, i_13_1792, i_13_1885, i_13_1914, i_13_2125, i_13_2191, i_13_2244, i_13_2379, i_13_2380, i_13_2434, i_13_2457, i_13_2541, i_13_2646, i_13_2647, i_13_2650, i_13_2820, i_13_2821, i_13_2847, i_13_2848, i_13_3091, i_13_3109, i_13_3269, i_13_3306, i_13_3307, i_13_3372, i_13_3387, i_13_3388, i_13_3429, i_13_3451, i_13_3538, i_13_3547, i_13_3555, i_13_3636, i_13_3637, i_13_3766, i_13_3836, i_13_3889, i_13_3906, i_13_3910, i_13_3934, i_13_3936, i_13_3988, i_13_4017, i_13_4032, i_13_4033, i_13_4036, i_13_4164, i_13_4269, i_13_4294, i_13_4327, i_13_4378, i_13_4396, i_13_4510, i_13_4593, o_13_189);
	kernel_13_190 k_13_190(i_13_76, i_13_184, i_13_189, i_13_229, i_13_408, i_13_415, i_13_418, i_13_517, i_13_549, i_13_571, i_13_604, i_13_657, i_13_658, i_13_665, i_13_761, i_13_793, i_13_847, i_13_855, i_13_856, i_13_885, i_13_936, i_13_937, i_13_1129, i_13_1144, i_13_1266, i_13_1420, i_13_1513, i_13_1518, i_13_1710, i_13_1711, i_13_1741, i_13_1742, i_13_1885, i_13_2019, i_13_2020, i_13_2024, i_13_2159, i_13_2224, i_13_2263, i_13_2321, i_13_2442, i_13_2448, i_13_2462, i_13_2466, i_13_2467, i_13_2470, i_13_2501, i_13_2512, i_13_2514, i_13_2538, i_13_2595, i_13_2611, i_13_2647, i_13_2692, i_13_2708, i_13_2730, i_13_2734, i_13_2881, i_13_2907, i_13_2908, i_13_2938, i_13_3037, i_13_3105, i_13_3325, i_13_3478, i_13_3483, i_13_3484, i_13_3486, i_13_3487, i_13_3565, i_13_3639, i_13_3640, i_13_3763, i_13_3861, i_13_3865, i_13_3868, i_13_3965, i_13_3992, i_13_4008, i_13_4009, i_13_4018, i_13_4098, i_13_4116, i_13_4127, i_13_4158, i_13_4159, i_13_4161, i_13_4198, i_13_4321, i_13_4324, i_13_4330, i_13_4333, i_13_4335, i_13_4365, i_13_4366, i_13_4369, i_13_4454, i_13_4458, i_13_4535, i_13_4599, o_13_190);
	kernel_13_191 k_13_191(i_13_46, i_13_47, i_13_66, i_13_100, i_13_262, i_13_567, i_13_585, i_13_587, i_13_639, i_13_640, i_13_675, i_13_689, i_13_946, i_13_1063, i_13_1064, i_13_1207, i_13_1260, i_13_1272, i_13_1282, i_13_1323, i_13_1343, i_13_1435, i_13_1468, i_13_1505, i_13_1507, i_13_1567, i_13_1568, i_13_1596, i_13_1597, i_13_1802, i_13_1810, i_13_1855, i_13_1927, i_13_1935, i_13_1945, i_13_1992, i_13_2017, i_13_2053, i_13_2054, i_13_2107, i_13_2117, i_13_2135, i_13_2146, i_13_2153, i_13_2189, i_13_2244, i_13_2261, i_13_2278, i_13_2279, i_13_2351, i_13_2404, i_13_2405, i_13_2417, i_13_2585, i_13_2611, i_13_2615, i_13_2694, i_13_2713, i_13_2745, i_13_2746, i_13_2782, i_13_2898, i_13_2934, i_13_2935, i_13_3025, i_13_3054, i_13_3145, i_13_3313, i_13_3339, i_13_3340, i_13_3341, i_13_3367, i_13_3368, i_13_3385, i_13_3386, i_13_3414, i_13_3415, i_13_3456, i_13_3481, i_13_3529, i_13_3548, i_13_3592, i_13_3627, i_13_3754, i_13_3817, i_13_3818, i_13_3889, i_13_3901, i_13_3909, i_13_3936, i_13_4041, i_13_4042, i_13_4230, i_13_4231, i_13_4232, i_13_4258, i_13_4268, i_13_4304, i_13_4324, i_13_4394, o_13_191);
	kernel_13_192 k_13_192(i_13_45, i_13_112, i_13_138, i_13_139, i_13_172, i_13_174, i_13_279, i_13_405, i_13_406, i_13_414, i_13_441, i_13_505, i_13_567, i_13_633, i_13_657, i_13_658, i_13_660, i_13_666, i_13_667, i_13_669, i_13_828, i_13_831, i_13_940, i_13_945, i_13_1071, i_13_1072, i_13_1081, i_13_1147, i_13_1228, i_13_1284, i_13_1305, i_13_1306, i_13_1326, i_13_1423, i_13_1494, i_13_1497, i_13_1498, i_13_1504, i_13_1522, i_13_1548, i_13_1593, i_13_1620, i_13_1633, i_13_1684, i_13_1695, i_13_1729, i_13_1737, i_13_1764, i_13_1777, i_13_1837, i_13_1858, i_13_1926, i_13_1938, i_13_2019, i_13_2020, i_13_2296, i_13_2316, i_13_2344, i_13_2395, i_13_2430, i_13_2431, i_13_2448, i_13_2469, i_13_2511, i_13_2610, i_13_2637, i_13_2719, i_13_2757, i_13_2781, i_13_3070, i_13_3108, i_13_3126, i_13_3172, i_13_3241, i_13_3258, i_13_3261, i_13_3268, i_13_3271, i_13_3406, i_13_3420, i_13_3423, i_13_3546, i_13_3637, i_13_3640, i_13_3667, i_13_3897, i_13_3910, i_13_4035, i_13_4051, i_13_4086, i_13_4248, i_13_4251, i_13_4252, i_13_4260, i_13_4321, i_13_4429, i_13_4458, i_13_4503, i_13_4564, i_13_4593, o_13_192);
	kernel_13_193 k_13_193(i_13_28, i_13_91, i_13_92, i_13_176, i_13_181, i_13_256, i_13_274, i_13_307, i_13_308, i_13_310, i_13_315, i_13_316, i_13_317, i_13_337, i_13_371, i_13_379, i_13_407, i_13_408, i_13_551, i_13_589, i_13_604, i_13_639, i_13_640, i_13_666, i_13_668, i_13_670, i_13_676, i_13_723, i_13_757, i_13_769, i_13_842, i_13_867, i_13_875, i_13_981, i_13_1021, i_13_1063, i_13_1093, i_13_1218, i_13_1300, i_13_1318, i_13_1324, i_13_1325, i_13_1480, i_13_1595, i_13_1602, i_13_1699, i_13_1828, i_13_1840, i_13_1909, i_13_1926, i_13_2116, i_13_2245, i_13_2260, i_13_2280, i_13_2407, i_13_2511, i_13_2648, i_13_2660, i_13_2673, i_13_2675, i_13_2678, i_13_2767, i_13_2781, i_13_2785, i_13_2981, i_13_3100, i_13_3128, i_13_3416, i_13_3469, i_13_3479, i_13_3482, i_13_3529, i_13_3541, i_13_3631, i_13_3682, i_13_3738, i_13_3766, i_13_3767, i_13_3817, i_13_3818, i_13_3889, i_13_3925, i_13_3991, i_13_3992, i_13_4033, i_13_4034, i_13_4041, i_13_4078, i_13_4086, i_13_4234, i_13_4252, i_13_4262, i_13_4270, i_13_4305, i_13_4351, i_13_4519, i_13_4522, i_13_4565, i_13_4567, i_13_4591, o_13_193);
	kernel_13_194 k_13_194(i_13_51, i_13_123, i_13_124, i_13_141, i_13_169, i_13_240, i_13_241, i_13_250, i_13_375, i_13_456, i_13_467, i_13_588, i_13_618, i_13_619, i_13_654, i_13_682, i_13_699, i_13_763, i_13_850, i_13_931, i_13_943, i_13_979, i_13_980, i_13_1033, i_13_1058, i_13_1059, i_13_1077, i_13_1078, i_13_1079, i_13_1084, i_13_1401, i_13_1448, i_13_1470, i_13_1501, i_13_1502, i_13_1507, i_13_1525, i_13_1528, i_13_1599, i_13_1608, i_13_1609, i_13_1635, i_13_1636, i_13_1637, i_13_1777, i_13_1815, i_13_2002, i_13_2014, i_13_2140, i_13_2211, i_13_2226, i_13_2284, i_13_2294, i_13_2319, i_13_2454, i_13_2544, i_13_2616, i_13_2787, i_13_2788, i_13_2887, i_13_2922, i_13_2923, i_13_2959, i_13_3003, i_13_3023, i_13_3219, i_13_3220, i_13_3372, i_13_3382, i_13_3406, i_13_3417, i_13_3418, i_13_3428, i_13_3463, i_13_3464, i_13_3471, i_13_3541, i_13_3553, i_13_3569, i_13_3577, i_13_3643, i_13_3723, i_13_3730, i_13_3769, i_13_3788, i_13_3877, i_13_3903, i_13_3904, i_13_4011, i_13_4012, i_13_4020, i_13_4082, i_13_4089, i_13_4091, i_13_4389, i_13_4396, i_13_4418, i_13_4533, i_13_4557, i_13_4589, o_13_194);
	kernel_13_195 k_13_195(i_13_64, i_13_65, i_13_76, i_13_131, i_13_158, i_13_160, i_13_163, i_13_164, i_13_307, i_13_355, i_13_358, i_13_463, i_13_465, i_13_466, i_13_469, i_13_490, i_13_492, i_13_537, i_13_564, i_13_580, i_13_697, i_13_812, i_13_829, i_13_831, i_13_839, i_13_1100, i_13_1121, i_13_1131, i_13_1302, i_13_1307, i_13_1345, i_13_1389, i_13_1396, i_13_1397, i_13_1400, i_13_1434, i_13_1471, i_13_1504, i_13_1594, i_13_1609, i_13_1696, i_13_1697, i_13_1783, i_13_1784, i_13_1793, i_13_1794, i_13_1840, i_13_1846, i_13_1847, i_13_1859, i_13_1928, i_13_1990, i_13_1995, i_13_2032, i_13_2101, i_13_2108, i_13_2111, i_13_2143, i_13_2187, i_13_2200, i_13_2202, i_13_2203, i_13_2206, i_13_2237, i_13_2297, i_13_2379, i_13_2404, i_13_2405, i_13_2506, i_13_2585, i_13_2692, i_13_2881, i_13_2884, i_13_2936, i_13_3165, i_13_3241, i_13_3242, i_13_3309, i_13_3380, i_13_3415, i_13_3422, i_13_3539, i_13_3568, i_13_3596, i_13_3597, i_13_3598, i_13_3619, i_13_3631, i_13_3633, i_13_3638, i_13_3686, i_13_3845, i_13_3856, i_13_3912, i_13_4060, i_13_4189, i_13_4313, i_13_4416, i_13_4453, i_13_4510, o_13_195);
	kernel_13_196 k_13_196(i_13_64, i_13_77, i_13_121, i_13_179, i_13_184, i_13_229, i_13_232, i_13_358, i_13_374, i_13_415, i_13_527, i_13_530, i_13_557, i_13_599, i_13_608, i_13_611, i_13_661, i_13_662, i_13_664, i_13_665, i_13_800, i_13_829, i_13_832, i_13_833, i_13_850, i_13_895, i_13_1066, i_13_1121, i_13_1213, i_13_1228, i_13_1229, i_13_1307, i_13_1309, i_13_1310, i_13_1313, i_13_1427, i_13_1430, i_13_1498, i_13_1499, i_13_1505, i_13_1553, i_13_1556, i_13_1568, i_13_1726, i_13_1811, i_13_1919, i_13_1922, i_13_1930, i_13_1961, i_13_1991, i_13_1993, i_13_2033, i_13_2297, i_13_2399, i_13_2452, i_13_2456, i_13_2467, i_13_2678, i_13_2693, i_13_2708, i_13_2768, i_13_2924, i_13_3010, i_13_3013, i_13_3037, i_13_3061, i_13_3062, i_13_3149, i_13_3217, i_13_3242, i_13_3260, i_13_3269, i_13_3289, i_13_3307, i_13_3394, i_13_3406, i_13_3461, i_13_3490, i_13_3523, i_13_3541, i_13_3542, i_13_3545, i_13_3580, i_13_3581, i_13_3734, i_13_3788, i_13_3806, i_13_3859, i_13_3860, i_13_3892, i_13_3895, i_13_3919, i_13_3983, i_13_4253, i_13_4256, i_13_4265, i_13_4430, i_13_4558, i_13_4559, i_13_4580, o_13_196);
	kernel_13_197 k_13_197(i_13_41, i_13_71, i_13_138, i_13_139, i_13_141, i_13_142, i_13_231, i_13_232, i_13_310, i_13_418, i_13_471, i_13_472, i_13_517, i_13_537, i_13_538, i_13_764, i_13_826, i_13_832, i_13_1029, i_13_1086, i_13_1214, i_13_1218, i_13_1219, i_13_1221, i_13_1222, i_13_1266, i_13_1276, i_13_1362, i_13_1392, i_13_1426, i_13_1473, i_13_1722, i_13_1725, i_13_1726, i_13_1734, i_13_1785, i_13_1788, i_13_1789, i_13_1842, i_13_1849, i_13_1857, i_13_1883, i_13_1884, i_13_1887, i_13_1889, i_13_2004, i_13_2122, i_13_2145, i_13_2146, i_13_2175, i_13_2231, i_13_2299, i_13_2464, i_13_2543, i_13_2616, i_13_2649, i_13_2650, i_13_2695, i_13_2766, i_13_2847, i_13_2851, i_13_2861, i_13_2877, i_13_3039, i_13_3067, i_13_3095, i_13_3103, i_13_3129, i_13_3148, i_13_3165, i_13_3173, i_13_3292, i_13_3391, i_13_3423, i_13_3427, i_13_3432, i_13_3472, i_13_3507, i_13_3534, i_13_3607, i_13_3688, i_13_3706, i_13_3796, i_13_3852, i_13_3869, i_13_3912, i_13_4017, i_13_4063, i_13_4094, i_13_4110, i_13_4188, i_13_4220, i_13_4256, i_13_4309, i_13_4315, i_13_4333, i_13_4381, i_13_4417, i_13_4593, i_13_4597, o_13_197);
	kernel_13_198 k_13_198(i_13_79, i_13_95, i_13_140, i_13_187, i_13_275, i_13_322, i_13_328, i_13_329, i_13_365, i_13_370, i_13_431, i_13_445, i_13_511, i_13_562, i_13_599, i_13_602, i_13_610, i_13_674, i_13_718, i_13_728, i_13_781, i_13_832, i_13_861, i_13_862, i_13_895, i_13_1023, i_13_1078, i_13_1096, i_13_1195, i_13_1258, i_13_1321, i_13_1343, i_13_1384, i_13_1516, i_13_1637, i_13_1687, i_13_1726, i_13_1751, i_13_1768, i_13_1849, i_13_1859, i_13_1886, i_13_1888, i_13_1907, i_13_1913, i_13_1954, i_13_2101, i_13_2123, i_13_2168, i_13_2290, i_13_2311, i_13_2399, i_13_2428, i_13_2462, i_13_2492, i_13_2633, i_13_2650, i_13_2651, i_13_2653, i_13_2654, i_13_2722, i_13_2852, i_13_2884, i_13_2887, i_13_2922, i_13_2941, i_13_2942, i_13_2983, i_13_3023, i_13_3056, i_13_3127, i_13_3146, i_13_3154, i_13_3172, i_13_3173, i_13_3175, i_13_3176, i_13_3235, i_13_3238, i_13_3392, i_13_3433, i_13_3544, i_13_3563, i_13_3732, i_13_3785, i_13_3794, i_13_3847, i_13_3876, i_13_3913, i_13_3914, i_13_3965, i_13_4021, i_13_4100, i_13_4162, i_13_4238, i_13_4342, i_13_4382, i_13_4409, i_13_4444, i_13_4513, o_13_198);
	kernel_13_199 k_13_199(i_13_74, i_13_121, i_13_122, i_13_125, i_13_142, i_13_175, i_13_176, i_13_227, i_13_229, i_13_311, i_13_338, i_13_341, i_13_517, i_13_524, i_13_533, i_13_535, i_13_536, i_13_596, i_13_599, i_13_617, i_13_766, i_13_830, i_13_850, i_13_911, i_13_977, i_13_1084, i_13_1085, i_13_1093, i_13_1139, i_13_1216, i_13_1433, i_13_1469, i_13_1496, i_13_1597, i_13_1598, i_13_1622, i_13_1721, i_13_1741, i_13_1757, i_13_1783, i_13_1784, i_13_1814, i_13_1817, i_13_1958, i_13_2012, i_13_2021, i_13_2120, i_13_2168, i_13_2210, i_13_2225, i_13_2309, i_13_2341, i_13_2432, i_13_2458, i_13_2462, i_13_2465, i_13_2500, i_13_2612, i_13_2630, i_13_2657, i_13_2714, i_13_2738, i_13_2818, i_13_2824, i_13_2885, i_13_3010, i_13_3019, i_13_3035, i_13_3037, i_13_3044, i_13_3128, i_13_3143, i_13_3169, i_13_3215, i_13_3217, i_13_3218, i_13_3221, i_13_3290, i_13_3413, i_13_3416, i_13_3449, i_13_3452, i_13_3524, i_13_3527, i_13_3737, i_13_3854, i_13_3865, i_13_3884, i_13_3998, i_13_4036, i_13_4055, i_13_4097, i_13_4238, i_13_4391, i_13_4414, i_13_4415, i_13_4519, i_13_4520, i_13_4523, i_13_4538, o_13_199);
	kernel_13_200 k_13_200(i_13_31, i_13_271, i_13_273, i_13_274, i_13_275, i_13_279, i_13_310, i_13_322, i_13_426, i_13_442, i_13_450, i_13_451, i_13_589, i_13_592, i_13_643, i_13_657, i_13_660, i_13_760, i_13_831, i_13_838, i_13_858, i_13_867, i_13_868, i_13_894, i_13_928, i_13_939, i_13_940, i_13_944, i_13_1017, i_13_1080, i_13_1081, i_13_1148, i_13_1150, i_13_1444, i_13_1470, i_13_1492, i_13_1497, i_13_1597, i_13_1632, i_13_1642, i_13_1733, i_13_1750, i_13_1765, i_13_1854, i_13_1947, i_13_2011, i_13_2140, i_13_2191, i_13_2226, i_13_2233, i_13_2380, i_13_2421, i_13_2449, i_13_2451, i_13_2467, i_13_2506, i_13_2541, i_13_2542, i_13_2544, i_13_2545, i_13_2568, i_13_2857, i_13_2884, i_13_2924, i_13_2955, i_13_3109, i_13_3142, i_13_3388, i_13_3414, i_13_3415, i_13_3451, i_13_3459, i_13_3460, i_13_3463, i_13_3475, i_13_3477, i_13_3486, i_13_3549, i_13_3567, i_13_3570, i_13_3576, i_13_3627, i_13_3900, i_13_3919, i_13_3928, i_13_3991, i_13_4054, i_13_4086, i_13_4162, i_13_4166, i_13_4265, i_13_4266, i_13_4368, i_13_4369, i_13_4433, i_13_4514, i_13_4537, i_13_4554, i_13_4555, i_13_4593, o_13_200);
	kernel_13_201 k_13_201(i_13_38, i_13_92, i_13_95, i_13_107, i_13_113, i_13_118, i_13_274, i_13_361, i_13_406, i_13_407, i_13_446, i_13_448, i_13_449, i_13_562, i_13_565, i_13_572, i_13_607, i_13_608, i_13_610, i_13_733, i_13_796, i_13_797, i_13_895, i_13_949, i_13_950, i_13_952, i_13_1034, i_13_1084, i_13_1087, i_13_1096, i_13_1186, i_13_1244, i_13_1253, i_13_1262, i_13_1409, i_13_1432, i_13_1441, i_13_1510, i_13_1541, i_13_1589, i_13_1633, i_13_1730, i_13_1750, i_13_1765, i_13_1787, i_13_1832, i_13_1841, i_13_1885, i_13_1954, i_13_2003, i_13_2120, i_13_2137, i_13_2173, i_13_2174, i_13_2177, i_13_2209, i_13_2435, i_13_2498, i_13_2564, i_13_2702, i_13_2875, i_13_2939, i_13_3035, i_13_3044, i_13_3047, i_13_3101, i_13_3104, i_13_3161, i_13_3163, i_13_3164, i_13_3209, i_13_3235, i_13_3344, i_13_3511, i_13_3703, i_13_3764, i_13_3803, i_13_3844, i_13_3847, i_13_3871, i_13_3872, i_13_3874, i_13_3875, i_13_3979, i_13_3980, i_13_4010, i_13_4081, i_13_4090, i_13_4118, i_13_4120, i_13_4121, i_13_4162, i_13_4163, i_13_4349, i_13_4351, i_13_4352, i_13_4354, i_13_4541, i_13_4568, i_13_4598, o_13_201);
	kernel_13_202 k_13_202(i_13_112, i_13_131, i_13_133, i_13_134, i_13_160, i_13_169, i_13_170, i_13_358, i_13_457, i_13_466, i_13_664, i_13_799, i_13_831, i_13_853, i_13_956, i_13_959, i_13_1078, i_13_1132, i_13_1231, i_13_1303, i_13_1310, i_13_1364, i_13_1400, i_13_1407, i_13_1446, i_13_1447, i_13_1471, i_13_1501, i_13_1507, i_13_1555, i_13_1556, i_13_1639, i_13_1699, i_13_1847, i_13_1849, i_13_1850, i_13_1896, i_13_1930, i_13_1961, i_13_2103, i_13_2104, i_13_2111, i_13_2143, i_13_2145, i_13_2146, i_13_2156, i_13_2202, i_13_2203, i_13_2204, i_13_2209, i_13_2237, i_13_2398, i_13_2407, i_13_2428, i_13_2429, i_13_2595, i_13_2681, i_13_2882, i_13_2936, i_13_2938, i_13_2939, i_13_2986, i_13_3028, i_13_3101, i_13_3146, i_13_3232, i_13_3242, i_13_3244, i_13_3245, i_13_3341, i_13_3406, i_13_3410, i_13_3637, i_13_3638, i_13_3644, i_13_3739, i_13_3755, i_13_3757, i_13_3758, i_13_3805, i_13_3812, i_13_3859, i_13_3860, i_13_3919, i_13_3935, i_13_4054, i_13_4061, i_13_4063, i_13_4214, i_13_4220, i_13_4270, i_13_4273, i_13_4313, i_13_4316, i_13_4423, i_13_4432, i_13_4453, i_13_4481, i_13_4510, i_13_4512, o_13_202);
	kernel_13_203 k_13_203(i_13_28, i_13_64, i_13_65, i_13_74, i_13_308, i_13_355, i_13_442, i_13_443, i_13_445, i_13_446, i_13_667, i_13_668, i_13_676, i_13_677, i_13_743, i_13_829, i_13_931, i_13_947, i_13_1081, i_13_1099, i_13_1100, i_13_1102, i_13_1274, i_13_1279, i_13_1306, i_13_1307, i_13_1397, i_13_1424, i_13_1435, i_13_1444, i_13_1499, i_13_1504, i_13_1505, i_13_1594, i_13_1595, i_13_1621, i_13_1634, i_13_1639, i_13_1642, i_13_1723, i_13_1768, i_13_1773, i_13_1774, i_13_1783, i_13_1793, i_13_1838, i_13_1847, i_13_1903, i_13_1921, i_13_1957, i_13_1958, i_13_1993, i_13_2002, i_13_2030, i_13_2200, i_13_2209, i_13_2317, i_13_2468, i_13_2512, i_13_2567, i_13_2656, i_13_2673, i_13_2675, i_13_2999, i_13_3061, i_13_3065, i_13_3073, i_13_3089, i_13_3109, i_13_3127, i_13_3128, i_13_3242, i_13_3397, i_13_3448, i_13_3449, i_13_3524, i_13_3551, i_13_3574, i_13_3595, i_13_3596, i_13_3619, i_13_3646, i_13_3781, i_13_3782, i_13_3857, i_13_3863, i_13_3890, i_13_3924, i_13_3925, i_13_3988, i_13_4061, i_13_4078, i_13_4087, i_13_4330, i_13_4342, i_13_4430, i_13_4433, i_13_4447, i_13_4520, i_13_4556, o_13_203);
	kernel_13_204 k_13_204(i_13_163, i_13_173, i_13_175, i_13_176, i_13_177, i_13_178, i_13_280, i_13_307, i_13_379, i_13_380, i_13_452, i_13_526, i_13_527, i_13_617, i_13_625, i_13_735, i_13_742, i_13_766, i_13_797, i_13_814, i_13_817, i_13_829, i_13_976, i_13_977, i_13_1063, i_13_1076, i_13_1093, i_13_1094, i_13_1204, i_13_1297, i_13_1309, i_13_1319, i_13_1327, i_13_1442, i_13_1445, i_13_1446, i_13_1460, i_13_1498, i_13_1499, i_13_1502, i_13_1594, i_13_1595, i_13_1601, i_13_1687, i_13_1732, i_13_1846, i_13_1850, i_13_1927, i_13_1931, i_13_1990, i_13_2020, i_13_2119, i_13_2135, i_13_2191, i_13_2246, i_13_2264, i_13_2405, i_13_2413, i_13_2425, i_13_2431, i_13_2505, i_13_2578, i_13_2849, i_13_2875, i_13_2935, i_13_2938, i_13_3011, i_13_3053, i_13_3109, i_13_3110, i_13_3130, i_13_3244, i_13_3373, i_13_3399, i_13_3416, i_13_3421, i_13_3423, i_13_3425, i_13_3428, i_13_3437, i_13_3523, i_13_3649, i_13_3728, i_13_3731, i_13_3794, i_13_3865, i_13_4018, i_13_4019, i_13_4051, i_13_4060, i_13_4061, i_13_4063, i_13_4136, i_13_4267, i_13_4268, i_13_4306, i_13_4312, i_13_4314, i_13_4342, i_13_4568, o_13_204);
	kernel_13_205 k_13_205(i_13_31, i_13_184, i_13_196, i_13_259, i_13_325, i_13_327, i_13_328, i_13_382, i_13_526, i_13_624, i_13_660, i_13_661, i_13_742, i_13_820, i_13_840, i_13_850, i_13_852, i_13_854, i_13_858, i_13_861, i_13_1020, i_13_1074, i_13_1093, i_13_1097, i_13_1227, i_13_1228, i_13_1229, i_13_1254, i_13_1255, i_13_1256, i_13_1258, i_13_1314, i_13_1317, i_13_1383, i_13_1428, i_13_1443, i_13_1444, i_13_1447, i_13_1483, i_13_1488, i_13_1645, i_13_1675, i_13_1691, i_13_1753, i_13_1848, i_13_1849, i_13_1854, i_13_1857, i_13_1858, i_13_1861, i_13_1953, i_13_1957, i_13_1993, i_13_2042, i_13_2247, i_13_2248, i_13_2281, i_13_2394, i_13_2407, i_13_2412, i_13_2434, i_13_2488, i_13_2614, i_13_2617, i_13_2701, i_13_2712, i_13_2857, i_13_2878, i_13_2978, i_13_3064, i_13_3118, i_13_3122, i_13_3153, i_13_3172, i_13_3307, i_13_3338, i_13_3355, i_13_3418, i_13_3436, i_13_3456, i_13_3460, i_13_3478, i_13_3484, i_13_3486, i_13_3487, i_13_3489, i_13_3537, i_13_3562, i_13_3689, i_13_3783, i_13_3802, i_13_3868, i_13_3907, i_13_4063, i_13_4351, i_13_4365, i_13_4372, i_13_4378, i_13_4396, i_13_4518, o_13_205);
	kernel_13_206 k_13_206(i_13_13, i_13_28, i_13_31, i_13_43, i_13_64, i_13_66, i_13_173, i_13_310, i_13_399, i_13_575, i_13_598, i_13_604, i_13_607, i_13_641, i_13_661, i_13_670, i_13_672, i_13_676, i_13_772, i_13_814, i_13_829, i_13_830, i_13_832, i_13_833, i_13_851, i_13_885, i_13_1066, i_13_1102, i_13_1113, i_13_1225, i_13_1232, i_13_1259, i_13_1306, i_13_1307, i_13_1309, i_13_1385, i_13_1442, i_13_1466, i_13_1491, i_13_1523, i_13_1549, i_13_1554, i_13_1639, i_13_1697, i_13_1729, i_13_1795, i_13_1927, i_13_1928, i_13_1965, i_13_2103, i_13_2135, i_13_2229, i_13_2297, i_13_2298, i_13_2381, i_13_2535, i_13_2552, i_13_2677, i_13_2720, i_13_2721, i_13_2740, i_13_2749, i_13_2802, i_13_2806, i_13_2879, i_13_2882, i_13_2963, i_13_3000, i_13_3047, i_13_3255, i_13_3308, i_13_3367, i_13_3368, i_13_3479, i_13_3537, i_13_3539, i_13_3544, i_13_3545, i_13_3556, i_13_3637, i_13_3730, i_13_3754, i_13_3755, i_13_3894, i_13_3910, i_13_3921, i_13_3935, i_13_4036, i_13_4063, i_13_4249, i_13_4294, i_13_4313, i_13_4342, i_13_4349, i_13_4371, i_13_4406, i_13_4414, i_13_4432, i_13_4592, i_13_4594, o_13_206);
	kernel_13_207 k_13_207(i_13_112, i_13_143, i_13_205, i_13_210, i_13_223, i_13_251, i_13_277, i_13_278, i_13_287, i_13_322, i_13_340, i_13_341, i_13_386, i_13_447, i_13_457, i_13_512, i_13_562, i_13_563, i_13_619, i_13_746, i_13_781, i_13_1024, i_13_1085, i_13_1087, i_13_1088, i_13_1411, i_13_1429, i_13_1430, i_13_1443, i_13_1475, i_13_1484, i_13_1573, i_13_1574, i_13_1623, i_13_1624, i_13_1625, i_13_1634, i_13_1651, i_13_1659, i_13_1736, i_13_1786, i_13_1816, i_13_1817, i_13_1844, i_13_1915, i_13_1939, i_13_2005, i_13_2123, i_13_2137, i_13_2276, i_13_2347, i_13_2348, i_13_2437, i_13_2455, i_13_2489, i_13_2501, i_13_2543, i_13_2555, i_13_2712, i_13_2715, i_13_2716, i_13_2717, i_13_2725, i_13_2726, i_13_2788, i_13_2858, i_13_2876, i_13_3047, i_13_3068, i_13_3148, i_13_3149, i_13_3166, i_13_3221, i_13_3238, i_13_3274, i_13_3328, i_13_3419, i_13_3454, i_13_3455, i_13_3525, i_13_3527, i_13_3554, i_13_3685, i_13_3688, i_13_3689, i_13_3724, i_13_3922, i_13_3932, i_13_3939, i_13_4036, i_13_4057, i_13_4094, i_13_4184, i_13_4274, i_13_4328, i_13_4400, i_13_4408, i_13_4522, i_13_4525, i_13_4544, o_13_207);
	kernel_13_208 k_13_208(i_13_32, i_13_49, i_13_104, i_13_106, i_13_117, i_13_175, i_13_185, i_13_189, i_13_193, i_13_196, i_13_216, i_13_337, i_13_526, i_13_569, i_13_575, i_13_602, i_13_616, i_13_625, i_13_626, i_13_643, i_13_711, i_13_742, i_13_746, i_13_757, i_13_780, i_13_839, i_13_845, i_13_895, i_13_897, i_13_1018, i_13_1093, i_13_1099, i_13_1226, i_13_1251, i_13_1310, i_13_1360, i_13_1381, i_13_1405, i_13_1464, i_13_1478, i_13_1480, i_13_1481, i_13_1499, i_13_1507, i_13_1643, i_13_1667, i_13_1678, i_13_1714, i_13_1720, i_13_1748, i_13_1750, i_13_1754, i_13_1760, i_13_1805, i_13_1808, i_13_1858, i_13_1930, i_13_2002, i_13_2119, i_13_2120, i_13_2138, i_13_2274, i_13_2309, i_13_2395, i_13_2408, i_13_2447, i_13_2458, i_13_2470, i_13_2506, i_13_2542, i_13_2621, i_13_2747, i_13_2751, i_13_2825, i_13_2848, i_13_2876, i_13_2999, i_13_3173, i_13_3220, i_13_3221, i_13_3260, i_13_3379, i_13_3380, i_13_3466, i_13_3721, i_13_3782, i_13_3790, i_13_3791, i_13_3937, i_13_3942, i_13_3989, i_13_4046, i_13_4101, i_13_4121, i_13_4238, i_13_4295, i_13_4315, i_13_4519, i_13_4523, i_13_4525, o_13_208);
	kernel_13_209 k_13_209(i_13_19, i_13_69, i_13_77, i_13_107, i_13_109, i_13_112, i_13_113, i_13_124, i_13_125, i_13_130, i_13_132, i_13_211, i_13_368, i_13_463, i_13_525, i_13_589, i_13_680, i_13_949, i_13_950, i_13_1061, i_13_1085, i_13_1087, i_13_1284, i_13_1311, i_13_1327, i_13_1428, i_13_1489, i_13_1490, i_13_1519, i_13_1525, i_13_1571, i_13_1574, i_13_1633, i_13_1634, i_13_1637, i_13_1643, i_13_1815, i_13_1840, i_13_1841, i_13_2045, i_13_2128, i_13_2137, i_13_2173, i_13_2266, i_13_2337, i_13_2380, i_13_2407, i_13_2435, i_13_2438, i_13_2501, i_13_2512, i_13_2542, i_13_2543, i_13_2713, i_13_2716, i_13_2717, i_13_2785, i_13_2923, i_13_3100, i_13_3144, i_13_3146, i_13_3148, i_13_3149, i_13_3166, i_13_3167, i_13_3227, i_13_3370, i_13_3371, i_13_3406, i_13_3418, i_13_3419, i_13_3455, i_13_3506, i_13_3530, i_13_3553, i_13_3623, i_13_3686, i_13_3688, i_13_3734, i_13_3770, i_13_3878, i_13_3892, i_13_3912, i_13_3919, i_13_4021, i_13_4048, i_13_4120, i_13_4174, i_13_4256, i_13_4355, i_13_4409, i_13_4417, i_13_4418, i_13_4513, i_13_4522, i_13_4523, i_13_4525, i_13_4544, i_13_4555, i_13_4561, o_13_209);
	kernel_13_210 k_13_210(i_13_35, i_13_77, i_13_103, i_13_107, i_13_121, i_13_140, i_13_161, i_13_358, i_13_368, i_13_382, i_13_383, i_13_386, i_13_458, i_13_584, i_13_592, i_13_737, i_13_745, i_13_746, i_13_934, i_13_950, i_13_953, i_13_1066, i_13_1087, i_13_1132, i_13_1214, i_13_1220, i_13_1304, i_13_1348, i_13_1349, i_13_1411, i_13_1438, i_13_1462, i_13_1474, i_13_1624, i_13_1724, i_13_1726, i_13_1768, i_13_1772, i_13_1840, i_13_1934, i_13_1942, i_13_2059, i_13_2060, i_13_2284, i_13_2285, i_13_2348, i_13_2408, i_13_2515, i_13_2518, i_13_2555, i_13_2617, i_13_2716, i_13_2717, i_13_2860, i_13_2861, i_13_2884, i_13_3130, i_13_3139, i_13_3148, i_13_3325, i_13_3326, i_13_3388, i_13_3391, i_13_3392, i_13_3526, i_13_3551, i_13_3562, i_13_3598, i_13_3599, i_13_3622, i_13_3623, i_13_3634, i_13_3635, i_13_3686, i_13_3734, i_13_3742, i_13_3743, i_13_3847, i_13_3923, i_13_4055, i_13_4085, i_13_4093, i_13_4100, i_13_4103, i_13_4121, i_13_4165, i_13_4166, i_13_4237, i_13_4255, i_13_4333, i_13_4345, i_13_4346, i_13_4388, i_13_4399, i_13_4400, i_13_4418, i_13_4454, i_13_4514, i_13_4525, i_13_4568, o_13_210);
	kernel_13_211 k_13_211(i_13_14, i_13_38, i_13_112, i_13_120, i_13_127, i_13_128, i_13_180, i_13_236, i_13_248, i_13_260, i_13_319, i_13_320, i_13_418, i_13_527, i_13_531, i_13_533, i_13_576, i_13_577, i_13_596, i_13_607, i_13_615, i_13_671, i_13_695, i_13_769, i_13_892, i_13_928, i_13_945, i_13_977, i_13_1022, i_13_1089, i_13_1117, i_13_1121, i_13_1301, i_13_1318, i_13_1396, i_13_1397, i_13_1462, i_13_1480, i_13_1674, i_13_1706, i_13_1714, i_13_1757, i_13_1760, i_13_1777, i_13_1805, i_13_1814, i_13_1904, i_13_1918, i_13_2137, i_13_2138, i_13_2141, i_13_2147, i_13_2165, i_13_2173, i_13_2181, i_13_2225, i_13_2300, i_13_2443, i_13_2444, i_13_2458, i_13_2459, i_13_2630, i_13_2748, i_13_2749, i_13_2755, i_13_2785, i_13_2786, i_13_2821, i_13_2822, i_13_2921, i_13_2935, i_13_3105, i_13_3128, i_13_3206, i_13_3218, i_13_3254, i_13_3371, i_13_3560, i_13_3593, i_13_3619, i_13_3620, i_13_3631, i_13_3721, i_13_3791, i_13_3911, i_13_3928, i_13_3929, i_13_3988, i_13_3989, i_13_4015, i_13_4082, i_13_4207, i_13_4312, i_13_4369, i_13_4379, i_13_4391, i_13_4519, i_13_4522, i_13_4525, i_13_4566, o_13_211);
	kernel_13_212 k_13_212(i_13_94, i_13_95, i_13_139, i_13_140, i_13_175, i_13_177, i_13_178, i_13_187, i_13_310, i_13_319, i_13_321, i_13_415, i_13_457, i_13_510, i_13_553, i_13_555, i_13_571, i_13_574, i_13_580, i_13_607, i_13_609, i_13_610, i_13_646, i_13_660, i_13_668, i_13_714, i_13_771, i_13_796, i_13_850, i_13_853, i_13_952, i_13_987, i_13_988, i_13_1080, i_13_1123, i_13_1184, i_13_1203, i_13_1226, i_13_1264, i_13_1282, i_13_1300, i_13_1302, i_13_1432, i_13_1457, i_13_1650, i_13_1818, i_13_1828, i_13_1831, i_13_1861, i_13_2092, i_13_2100, i_13_2140, i_13_2172, i_13_2175, i_13_2176, i_13_2177, i_13_2346, i_13_2425, i_13_2427, i_13_2446, i_13_2470, i_13_2624, i_13_2676, i_13_2695, i_13_2860, i_13_2887, i_13_2901, i_13_3014, i_13_3108, i_13_3109, i_13_3112, i_13_3208, i_13_3217, i_13_3271, i_13_3415, i_13_3418, i_13_3423, i_13_3426, i_13_3488, i_13_3615, i_13_3616, i_13_3641, i_13_3685, i_13_3819, i_13_3820, i_13_3874, i_13_3994, i_13_4054, i_13_4080, i_13_4084, i_13_4251, i_13_4359, i_13_4436, i_13_4522, i_13_4523, i_13_4566, i_13_4567, i_13_4569, i_13_4570, i_13_4593, o_13_212);
	kernel_13_213 k_13_213(i_13_70, i_13_71, i_13_78, i_13_79, i_13_176, i_13_223, i_13_313, i_13_338, i_13_448, i_13_601, i_13_608, i_13_610, i_13_611, i_13_661, i_13_662, i_13_664, i_13_682, i_13_689, i_13_760, i_13_764, i_13_823, i_13_953, i_13_985, i_13_1103, i_13_1105, i_13_1123, i_13_1151, i_13_1232, i_13_1275, i_13_1276, i_13_1313, i_13_1318, i_13_1399, i_13_1511, i_13_1542, i_13_1601, i_13_1627, i_13_1645, i_13_1733, i_13_1736, i_13_1764, i_13_1768, i_13_1797, i_13_1798, i_13_1799, i_13_1843, i_13_1888, i_13_1947, i_13_1948, i_13_1996, i_13_2023, i_13_2024, i_13_2177, i_13_2426, i_13_2437, i_13_2507, i_13_2679, i_13_2680, i_13_2681, i_13_2697, i_13_2788, i_13_2851, i_13_2929, i_13_2930, i_13_3001, i_13_3130, i_13_3146, i_13_3220, i_13_3274, i_13_3370, i_13_3418, i_13_3652, i_13_3656, i_13_3761, i_13_3822, i_13_3823, i_13_3847, i_13_3895, i_13_3931, i_13_3941, i_13_3970, i_13_3994, i_13_4019, i_13_4040, i_13_4063, i_13_4084, i_13_4175, i_13_4189, i_13_4252, i_13_4297, i_13_4325, i_13_4450, i_13_4453, i_13_4517, i_13_4522, i_13_4597, i_13_4598, i_13_4602, i_13_4606, i_13_4607, o_13_213);
	kernel_13_214 k_13_214(i_13_4, i_13_70, i_13_111, i_13_139, i_13_193, i_13_229, i_13_382, i_13_480, i_13_519, i_13_607, i_13_610, i_13_628, i_13_655, i_13_661, i_13_663, i_13_682, i_13_683, i_13_886, i_13_934, i_13_939, i_13_940, i_13_988, i_13_1065, i_13_1086, i_13_1087, i_13_1132, i_13_1147, i_13_1156, i_13_1321, i_13_1330, i_13_1335, i_13_1519, i_13_1573, i_13_1660, i_13_1678, i_13_1735, i_13_1744, i_13_1745, i_13_1798, i_13_1994, i_13_2020, i_13_2022, i_13_2023, i_13_2024, i_13_2027, i_13_2198, i_13_2274, i_13_2338, i_13_2345, i_13_2455, i_13_2471, i_13_2482, i_13_2501, i_13_2507, i_13_2573, i_13_2715, i_13_2743, i_13_2765, i_13_2939, i_13_3031, i_13_3075, i_13_3076, i_13_3094, i_13_3234, i_13_3244, i_13_3265, i_13_3355, i_13_3452, i_13_3453, i_13_3454, i_13_3455, i_13_3549, i_13_3616, i_13_3635, i_13_3643, i_13_3647, i_13_3649, i_13_3670, i_13_3742, i_13_3822, i_13_3823, i_13_3939, i_13_4063, i_13_4126, i_13_4164, i_13_4165, i_13_4166, i_13_4171, i_13_4175, i_13_4189, i_13_4192, i_13_4201, i_13_4209, i_13_4324, i_13_4370, i_13_4596, i_13_4597, i_13_4603, i_13_4606, i_13_4607, o_13_214);
	kernel_13_215 k_13_215(i_13_40, i_13_136, i_13_193, i_13_228, i_13_229, i_13_265, i_13_378, i_13_445, i_13_586, i_13_639, i_13_643, i_13_680, i_13_692, i_13_711, i_13_738, i_13_768, i_13_975, i_13_1117, i_13_1124, i_13_1246, i_13_1269, i_13_1270, i_13_1314, i_13_1341, i_13_1342, i_13_1387, i_13_1388, i_13_1390, i_13_1440, i_13_1467, i_13_1468, i_13_1512, i_13_1513, i_13_1520, i_13_1567, i_13_1587, i_13_1633, i_13_1638, i_13_1722, i_13_1723, i_13_1726, i_13_1740, i_13_1767, i_13_1792, i_13_1793, i_13_1801, i_13_1903, i_13_1926, i_13_1944, i_13_1945, i_13_2029, i_13_2056, i_13_2134, i_13_2277, i_13_2278, i_13_2377, i_13_2411, i_13_2458, i_13_2461, i_13_2646, i_13_2721, i_13_2745, i_13_2746, i_13_2847, i_13_2874, i_13_3123, i_13_3135, i_13_3221, i_13_3340, i_13_3343, i_13_3366, i_13_3367, i_13_3384, i_13_3385, i_13_3439, i_13_3443, i_13_3636, i_13_3730, i_13_3784, i_13_3790, i_13_3793, i_13_3927, i_13_3928, i_13_4017, i_13_4018, i_13_4041, i_13_4042, i_13_4186, i_13_4216, i_13_4230, i_13_4231, i_13_4266, i_13_4293, i_13_4294, i_13_4338, i_13_4375, i_13_4410, i_13_4411, i_13_4447, i_13_4538, o_13_215);
	kernel_13_216 k_13_216(i_13_75, i_13_132, i_13_240, i_13_250, i_13_258, i_13_274, i_13_277, i_13_321, i_13_339, i_13_357, i_13_456, i_13_561, i_13_588, i_13_618, i_13_642, i_13_699, i_13_844, i_13_850, i_13_858, i_13_943, i_13_1077, i_13_1084, i_13_1105, i_13_1326, i_13_1363, i_13_1399, i_13_1431, i_13_1437, i_13_1470, i_13_1488, i_13_1489, i_13_1507, i_13_1527, i_13_1528, i_13_1552, i_13_1570, i_13_1591, i_13_1608, i_13_1693, i_13_1807, i_13_1908, i_13_1917, i_13_1920, i_13_2002, i_13_2004, i_13_2016, i_13_2032, i_13_2110, i_13_2302, i_13_2437, i_13_2502, i_13_2535, i_13_2544, i_13_2545, i_13_2589, i_13_2751, i_13_2766, i_13_2769, i_13_2787, i_13_2937, i_13_3024, i_13_3025, i_13_3064, i_13_3070, i_13_3129, i_13_3130, i_13_3220, i_13_3315, i_13_3372, i_13_3417, i_13_3418, i_13_3448, i_13_3471, i_13_3489, i_13_3552, i_13_3598, i_13_3613, i_13_3643, i_13_3646, i_13_3687, i_13_3705, i_13_3711, i_13_3714, i_13_3856, i_13_3876, i_13_3903, i_13_3904, i_13_4083, i_13_4084, i_13_4090, i_13_4117, i_13_4160, i_13_4189, i_13_4360, i_13_4362, i_13_4378, i_13_4452, i_13_4540, i_13_4543, i_13_4588, o_13_216);
	kernel_13_217 k_13_217(i_13_97, i_13_116, i_13_117, i_13_121, i_13_122, i_13_124, i_13_125, i_13_171, i_13_229, i_13_279, i_13_340, i_13_427, i_13_575, i_13_589, i_13_602, i_13_657, i_13_728, i_13_741, i_13_800, i_13_823, i_13_931, i_13_949, i_13_951, i_13_985, i_13_1024, i_13_1096, i_13_1123, i_13_1224, i_13_1282, i_13_1283, i_13_1304, i_13_1489, i_13_1490, i_13_1597, i_13_1600, i_13_1713, i_13_1787, i_13_1817, i_13_1844, i_13_1848, i_13_2056, i_13_2090, i_13_2118, i_13_2205, i_13_2209, i_13_2404, i_13_2429, i_13_2458, i_13_2461, i_13_2465, i_13_2614, i_13_2615, i_13_2639, i_13_2698, i_13_2785, i_13_2884, i_13_2980, i_13_3023, i_13_3047, i_13_3105, i_13_3146, i_13_3166, i_13_3167, i_13_3176, i_13_3208, i_13_3214, i_13_3220, i_13_3221, i_13_3267, i_13_3418, i_13_3420, i_13_3421, i_13_3425, i_13_3506, i_13_3532, i_13_3535, i_13_3553, i_13_3688, i_13_3699, i_13_3700, i_13_3788, i_13_3875, i_13_3877, i_13_3878, i_13_3928, i_13_3981, i_13_3985, i_13_4008, i_13_4013, i_13_4018, i_13_4036, i_13_4261, i_13_4328, i_13_4522, i_13_4523, i_13_4543, i_13_4544, i_13_4554, i_13_4561, i_13_4597, o_13_217);
	kernel_13_218 k_13_218(i_13_58, i_13_121, i_13_183, i_13_185, i_13_192, i_13_199, i_13_225, i_13_324, i_13_325, i_13_378, i_13_380, i_13_396, i_13_441, i_13_486, i_13_526, i_13_570, i_13_576, i_13_588, i_13_589, i_13_640, i_13_660, i_13_669, i_13_697, i_13_714, i_13_715, i_13_741, i_13_756, i_13_828, i_13_829, i_13_858, i_13_859, i_13_893, i_13_927, i_13_929, i_13_948, i_13_1084, i_13_1102, i_13_1118, i_13_1210, i_13_1219, i_13_1224, i_13_1225, i_13_1227, i_13_1254, i_13_1296, i_13_1369, i_13_1408, i_13_1413, i_13_1434, i_13_1488, i_13_1489, i_13_1507, i_13_1629, i_13_1719, i_13_1720, i_13_1782, i_13_1800, i_13_1818, i_13_1819, i_13_1882, i_13_1990, i_13_2011, i_13_2055, i_13_2128, i_13_2210, i_13_2224, i_13_2262, i_13_2343, i_13_2358, i_13_2503, i_13_2532, i_13_2722, i_13_2757, i_13_2766, i_13_2980, i_13_2981, i_13_3024, i_13_3114, i_13_3171, i_13_3259, i_13_3285, i_13_3286, i_13_3287, i_13_3420, i_13_3421, i_13_3423, i_13_3424, i_13_3451, i_13_3577, i_13_3649, i_13_3873, i_13_4008, i_13_4009, i_13_4050, i_13_4077, i_13_4087, i_13_4167, i_13_4232, i_13_4557, i_13_4582, o_13_218);
	kernel_13_219 k_13_219(i_13_49, i_13_101, i_13_109, i_13_112, i_13_141, i_13_175, i_13_210, i_13_220, i_13_279, i_13_281, i_13_284, i_13_287, i_13_317, i_13_337, i_13_382, i_13_425, i_13_445, i_13_534, i_13_550, i_13_551, i_13_554, i_13_613, i_13_652, i_13_653, i_13_654, i_13_655, i_13_658, i_13_668, i_13_676, i_13_677, i_13_679, i_13_688, i_13_844, i_13_852, i_13_853, i_13_1018, i_13_1144, i_13_1216, i_13_1300, i_13_1400, i_13_1423, i_13_1424, i_13_1516, i_13_1624, i_13_1643, i_13_1658, i_13_1668, i_13_1671, i_13_1748, i_13_1774, i_13_1801, i_13_1804, i_13_1840, i_13_1842, i_13_1921, i_13_1945, i_13_2000, i_13_2101, i_13_2146, i_13_2170, i_13_2331, i_13_2380, i_13_2433, i_13_2472, i_13_2473, i_13_2611, i_13_2674, i_13_2693, i_13_2697, i_13_2722, i_13_2767, i_13_2847, i_13_2850, i_13_2938, i_13_2956, i_13_2999, i_13_3054, i_13_3108, i_13_3368, i_13_3502, i_13_3523, i_13_3524, i_13_3637, i_13_3640, i_13_3767, i_13_3863, i_13_3889, i_13_3890, i_13_4034, i_13_4045, i_13_4117, i_13_4121, i_13_4270, i_13_4314, i_13_4377, i_13_4413, i_13_4556, i_13_4558, i_13_4600, i_13_4601, o_13_219);
	kernel_13_220 k_13_220(i_13_48, i_13_134, i_13_184, i_13_234, i_13_238, i_13_322, i_13_351, i_13_354, i_13_357, i_13_358, i_13_374, i_13_455, i_13_480, i_13_525, i_13_529, i_13_530, i_13_558, i_13_1024, i_13_1053, i_13_1079, i_13_1080, i_13_1085, i_13_1210, i_13_1371, i_13_1396, i_13_1399, i_13_1422, i_13_1426, i_13_1430, i_13_1458, i_13_1497, i_13_1498, i_13_1501, i_13_1502, i_13_1504, i_13_1555, i_13_1556, i_13_1620, i_13_1629, i_13_1637, i_13_1917, i_13_1921, i_13_1950, i_13_2006, i_13_2031, i_13_2033, i_13_2109, i_13_2203, i_13_2300, i_13_2368, i_13_2510, i_13_2511, i_13_2542, i_13_2691, i_13_2723, i_13_2767, i_13_2768, i_13_2788, i_13_2924, i_13_2934, i_13_2939, i_13_2955, i_13_2959, i_13_3014, i_13_3065, i_13_3069, i_13_3110, i_13_3123, i_13_3221, i_13_3235, i_13_3316, i_13_3373, i_13_3374, i_13_3403, i_13_3405, i_13_3432, i_13_3439, i_13_3464, i_13_3491, i_13_3576, i_13_3581, i_13_3594, i_13_3598, i_13_3599, i_13_3618, i_13_3646, i_13_3733, i_13_3781, i_13_3860, i_13_3904, i_13_3987, i_13_4067, i_13_4108, i_13_4212, i_13_4249, i_13_4271, i_13_4329, i_13_4453, i_13_4454, i_13_4561, o_13_220);
	kernel_13_221 k_13_221(i_13_37, i_13_73, i_13_74, i_13_109, i_13_110, i_13_113, i_13_116, i_13_122, i_13_157, i_13_262, i_13_365, i_13_366, i_13_551, i_13_559, i_13_562, i_13_604, i_13_605, i_13_613, i_13_639, i_13_676, i_13_677, i_13_814, i_13_821, i_13_947, i_13_992, i_13_1081, i_13_1084, i_13_1085, i_13_1120, i_13_1144, i_13_1217, i_13_1220, i_13_1283, i_13_1408, i_13_1424, i_13_1521, i_13_1541, i_13_1567, i_13_1621, i_13_1631, i_13_1720, i_13_1721, i_13_1775, i_13_1837, i_13_1838, i_13_1840, i_13_1841, i_13_1898, i_13_1945, i_13_1957, i_13_2021, i_13_2054, i_13_2134, i_13_2170, i_13_2171, i_13_2341, i_13_2345, i_13_2404, i_13_2432, i_13_2498, i_13_2611, i_13_2702, i_13_2746, i_13_2767, i_13_2818, i_13_2845, i_13_2846, i_13_2956, i_13_2958, i_13_3044, i_13_3098, i_13_3099, i_13_3100, i_13_3110, i_13_3125, i_13_3142, i_13_3146, i_13_3148, i_13_3152, i_13_3376, i_13_3377, i_13_3404, i_13_3452, i_13_3503, i_13_3524, i_13_3552, i_13_3686, i_13_3731, i_13_3736, i_13_3737, i_13_3802, i_13_3836, i_13_3910, i_13_3917, i_13_4051, i_13_4118, i_13_4160, i_13_4339, i_13_4541, i_13_4542, o_13_221);
	kernel_13_222 k_13_222(i_13_40, i_13_100, i_13_106, i_13_115, i_13_116, i_13_125, i_13_184, i_13_197, i_13_269, i_13_278, i_13_602, i_13_610, i_13_611, i_13_664, i_13_665, i_13_700, i_13_701, i_13_763, i_13_772, i_13_832, i_13_862, i_13_863, i_13_872, i_13_932, i_13_943, i_13_944, i_13_950, i_13_953, i_13_1075, i_13_1085, i_13_1262, i_13_1277, i_13_1286, i_13_1298, i_13_1411, i_13_1438, i_13_1481, i_13_1501, i_13_1539, i_13_1625, i_13_1636, i_13_1637, i_13_1660, i_13_1661, i_13_1682, i_13_1734, i_13_1843, i_13_1844, i_13_1931, i_13_1961, i_13_1996, i_13_2003, i_13_2006, i_13_2140, i_13_2303, i_13_2320, i_13_2438, i_13_2456, i_13_2536, i_13_2544, i_13_2545, i_13_2546, i_13_2616, i_13_2617, i_13_2618, i_13_2663, i_13_2798, i_13_2887, i_13_2888, i_13_2959, i_13_3004, i_13_3050, i_13_3113, i_13_3262, i_13_3316, i_13_3464, i_13_3490, i_13_3535, i_13_3571, i_13_3604, i_13_3731, i_13_3733, i_13_3769, i_13_3770, i_13_3878, i_13_3904, i_13_3905, i_13_3910, i_13_4090, i_13_4091, i_13_4166, i_13_4211, i_13_4343, i_13_4358, i_13_4372, i_13_4373, i_13_4391, i_13_4433, i_13_4517, i_13_4586, o_13_222);
	kernel_13_223 k_13_223(i_13_76, i_13_118, i_13_156, i_13_162, i_13_163, i_13_244, i_13_310, i_13_319, i_13_336, i_13_337, i_13_381, i_13_453, i_13_561, i_13_567, i_13_615, i_13_633, i_13_654, i_13_757, i_13_841, i_13_855, i_13_960, i_13_1063, i_13_1120, i_13_1218, i_13_1219, i_13_1300, i_13_1344, i_13_1434, i_13_1458, i_13_1522, i_13_1566, i_13_1593, i_13_1620, i_13_1693, i_13_1734, i_13_1783, i_13_1785, i_13_1786, i_13_1803, i_13_1813, i_13_1815, i_13_1816, i_13_1854, i_13_1992, i_13_2115, i_13_2116, i_13_2133, i_13_2205, i_13_2208, i_13_2212, i_13_2213, i_13_2403, i_13_2404, i_13_2421, i_13_2556, i_13_2584, i_13_2712, i_13_2935, i_13_2937, i_13_2938, i_13_3015, i_13_3034, i_13_3036, i_13_3060, i_13_3106, i_13_3145, i_13_3160, i_13_3213, i_13_3214, i_13_3216, i_13_3217, i_13_3220, i_13_3234, i_13_3268, i_13_3325, i_13_3438, i_13_3717, i_13_3741, i_13_3745, i_13_3816, i_13_3817, i_13_3843, i_13_3870, i_13_3884, i_13_3891, i_13_3982, i_13_4006, i_13_4041, i_13_4053, i_13_4207, i_13_4261, i_13_4302, i_13_4314, i_13_4321, i_13_4522, i_13_4530, i_13_4533, i_13_4582, i_13_4591, i_13_4600, o_13_223);
	kernel_13_224 k_13_224(i_13_41, i_13_74, i_13_76, i_13_103, i_13_112, i_13_113, i_13_184, i_13_185, i_13_193, i_13_208, i_13_316, i_13_317, i_13_374, i_13_571, i_13_572, i_13_575, i_13_643, i_13_644, i_13_685, i_13_689, i_13_715, i_13_778, i_13_811, i_13_814, i_13_895, i_13_982, i_13_983, i_13_1064, i_13_1067, i_13_1096, i_13_1102, i_13_1120, i_13_1121, i_13_1282, i_13_1507, i_13_1525, i_13_1678, i_13_1747, i_13_1750, i_13_1751, i_13_1804, i_13_1805, i_13_1829, i_13_1832, i_13_1834, i_13_1858, i_13_1907, i_13_1912, i_13_1921, i_13_2002, i_13_2044, i_13_2116, i_13_2120, i_13_2135, i_13_2137, i_13_2180, i_13_2264, i_13_2273, i_13_2404, i_13_2408, i_13_2434, i_13_2470, i_13_2542, i_13_2567, i_13_2651, i_13_2677, i_13_2692, i_13_2693, i_13_2696, i_13_2713, i_13_2737, i_13_2746, i_13_2747, i_13_2798, i_13_2920, i_13_2936, i_13_3206, i_13_3208, i_13_3209, i_13_3272, i_13_3406, i_13_3407, i_13_3427, i_13_3478, i_13_3607, i_13_3650, i_13_3686, i_13_3719, i_13_3817, i_13_3818, i_13_3854, i_13_3892, i_13_3989, i_13_4033, i_13_4036, i_13_4042, i_13_4141, i_13_4396, i_13_4421, i_13_4567, o_13_224);
	kernel_13_225 k_13_225(i_13_51, i_13_69, i_13_153, i_13_169, i_13_186, i_13_283, i_13_285, i_13_286, i_13_310, i_13_318, i_13_319, i_13_328, i_13_364, i_13_384, i_13_385, i_13_448, i_13_569, i_13_625, i_13_642, i_13_646, i_13_673, i_13_681, i_13_688, i_13_690, i_13_697, i_13_759, i_13_816, i_13_817, i_13_844, i_13_1122, i_13_1254, i_13_1255, i_13_1303, i_13_1438, i_13_1542, i_13_1572, i_13_1599, i_13_1644, i_13_1677, i_13_1723, i_13_1777, i_13_1851, i_13_1852, i_13_1933, i_13_1954, i_13_2001, i_13_2055, i_13_2058, i_13_2119, i_13_2184, i_13_2280, i_13_2319, i_13_2407, i_13_2409, i_13_2410, i_13_2578, i_13_2614, i_13_2626, i_13_2679, i_13_2697, i_13_2698, i_13_2923, i_13_2940, i_13_2941, i_13_3112, i_13_3117, i_13_3129, i_13_3145, i_13_3210, i_13_3291, i_13_3399, i_13_3400, i_13_3417, i_13_3460, i_13_3541, i_13_3613, i_13_3705, i_13_3768, i_13_3820, i_13_3858, i_13_3993, i_13_3994, i_13_4021, i_13_4038, i_13_4056, i_13_4065, i_13_4066, i_13_4162, i_13_4308, i_13_4309, i_13_4317, i_13_4318, i_13_4341, i_13_4344, i_13_4378, i_13_4381, i_13_4440, i_13_4461, i_13_4594, i_13_4597, o_13_225);
	kernel_13_226 k_13_226(i_13_91, i_13_94, i_13_114, i_13_118, i_13_121, i_13_123, i_13_136, i_13_190, i_13_231, i_13_276, i_13_376, i_13_396, i_13_474, i_13_517, i_13_597, i_13_609, i_13_732, i_13_793, i_13_832, i_13_840, i_13_841, i_13_861, i_13_862, i_13_879, i_13_913, i_13_950, i_13_1257, i_13_1272, i_13_1309, i_13_1491, i_13_1532, i_13_1599, i_13_1626, i_13_1736, i_13_1748, i_13_1786, i_13_1831, i_13_1839, i_13_1840, i_13_1842, i_13_1843, i_13_1930, i_13_1993, i_13_2117, i_13_2175, i_13_2206, i_13_2208, i_13_2211, i_13_2306, i_13_2361, i_13_2424, i_13_2426, i_13_2431, i_13_2436, i_13_2437, i_13_2459, i_13_2461, i_13_2463, i_13_2470, i_13_2541, i_13_2544, i_13_2616, i_13_2727, i_13_2744, i_13_3037, i_13_3163, i_13_3206, i_13_3369, i_13_3377, i_13_3422, i_13_3423, i_13_3426, i_13_3455, i_13_3530, i_13_3534, i_13_3651, i_13_3702, i_13_3849, i_13_3870, i_13_3871, i_13_3873, i_13_3874, i_13_3876, i_13_3877, i_13_3912, i_13_3991, i_13_4036, i_13_4086, i_13_4115, i_13_4180, i_13_4192, i_13_4206, i_13_4258, i_13_4271, i_13_4325, i_13_4349, i_13_4350, i_13_4351, i_13_4415, i_13_4582, o_13_226);
	kernel_13_227 k_13_227(i_13_31, i_13_45, i_13_174, i_13_262, i_13_352, i_13_373, i_13_489, i_13_507, i_13_553, i_13_567, i_13_606, i_13_607, i_13_625, i_13_627, i_13_657, i_13_658, i_13_679, i_13_697, i_13_819, i_13_823, i_13_850, i_13_931, i_13_936, i_13_960, i_13_981, i_13_1021, i_13_1129, i_13_1224, i_13_1225, i_13_1228, i_13_1327, i_13_1359, i_13_1515, i_13_1522, i_13_1609, i_13_1677, i_13_1729, i_13_1732, i_13_1764, i_13_1767, i_13_1768, i_13_1771, i_13_1794, i_13_1795, i_13_1831, i_13_1832, i_13_2019, i_13_2020, i_13_2113, i_13_2120, i_13_2146, i_13_2237, i_13_2469, i_13_2470, i_13_2473, i_13_2541, i_13_2562, i_13_2566, i_13_2592, i_13_2767, i_13_2835, i_13_2848, i_13_2901, i_13_2908, i_13_2983, i_13_3028, i_13_3087, i_13_3123, i_13_3132, i_13_3208, i_13_3220, i_13_3234, i_13_3261, i_13_3262, i_13_3264, i_13_3270, i_13_3381, i_13_3417, i_13_3418, i_13_3483, i_13_3546, i_13_3613, i_13_3651, i_13_3720, i_13_3729, i_13_3730, i_13_3819, i_13_3820, i_13_3897, i_13_3901, i_13_3978, i_13_4035, i_13_4161, i_13_4162, i_13_4164, i_13_4321, i_13_4344, i_13_4350, i_13_4476, i_13_4603, o_13_227);
	kernel_13_228 k_13_228(i_13_73, i_13_94, i_13_96, i_13_120, i_13_192, i_13_199, i_13_228, i_13_323, i_13_373, i_13_380, i_13_441, i_13_485, i_13_492, i_13_526, i_13_570, i_13_588, i_13_593, i_13_647, i_13_661, i_13_712, i_13_714, i_13_735, i_13_819, i_13_841, i_13_858, i_13_899, i_13_917, i_13_948, i_13_950, i_13_1066, i_13_1080, i_13_1298, i_13_1327, i_13_1394, i_13_1400, i_13_1407, i_13_1443, i_13_1569, i_13_1570, i_13_1627, i_13_1639, i_13_1673, i_13_1691, i_13_1722, i_13_1800, i_13_1831, i_13_1956, i_13_2011, i_13_2141, i_13_2210, i_13_2238, i_13_2239, i_13_2281, i_13_2407, i_13_2424, i_13_2425, i_13_2474, i_13_2532, i_13_2589, i_13_2636, i_13_2705, i_13_2739, i_13_2874, i_13_2935, i_13_2955, i_13_2986, i_13_3024, i_13_3026, i_13_3240, i_13_3241, i_13_3258, i_13_3370, i_13_3395, i_13_3421, i_13_3424, i_13_3426, i_13_3450, i_13_3463, i_13_3521, i_13_3595, i_13_3666, i_13_3753, i_13_3791, i_13_3797, i_13_3842, i_13_3846, i_13_3873, i_13_3893, i_13_3918, i_13_3919, i_13_3932, i_13_3981, i_13_4008, i_13_4009, i_13_4043, i_13_4077, i_13_4090, i_13_4193, i_13_4353, i_13_4584, o_13_228);
	kernel_13_229 k_13_229(i_13_48, i_13_66, i_13_67, i_13_105, i_13_136, i_13_447, i_13_469, i_13_529, i_13_568, i_13_609, i_13_615, i_13_619, i_13_627, i_13_628, i_13_645, i_13_646, i_13_669, i_13_760, i_13_763, i_13_781, i_13_933, i_13_994, i_13_1074, i_13_1084, i_13_1086, i_13_1095, i_13_1122, i_13_1131, i_13_1132, i_13_1167, i_13_1317, i_13_1482, i_13_1483, i_13_1501, i_13_1525, i_13_1634, i_13_1645, i_13_1716, i_13_1752, i_13_1770, i_13_1788, i_13_1798, i_13_1806, i_13_1807, i_13_1857, i_13_1914, i_13_1995, i_13_2022, i_13_2023, i_13_2091, i_13_2122, i_13_2134, i_13_2291, i_13_2364, i_13_2462, i_13_2472, i_13_2473, i_13_2488, i_13_2515, i_13_2569, i_13_2581, i_13_2676, i_13_2722, i_13_2857, i_13_2909, i_13_2912, i_13_2940, i_13_2981, i_13_3030, i_13_3031, i_13_3076, i_13_3211, i_13_3264, i_13_3435, i_13_3459, i_13_3479, i_13_3487, i_13_3505, i_13_3669, i_13_3759, i_13_3783, i_13_3822, i_13_3856, i_13_3900, i_13_3901, i_13_3907, i_13_4017, i_13_4063, i_13_4101, i_13_4161, i_13_4164, i_13_4165, i_13_4270, i_13_4272, i_13_4296, i_13_4324, i_13_4416, i_13_4521, i_13_4523, i_13_4606, o_13_229);
	kernel_13_230 k_13_230(i_13_26, i_13_38, i_13_40, i_13_79, i_13_103, i_13_105, i_13_266, i_13_431, i_13_599, i_13_607, i_13_677, i_13_679, i_13_685, i_13_686, i_13_717, i_13_761, i_13_778, i_13_815, i_13_816, i_13_839, i_13_895, i_13_924, i_13_983, i_13_1088, i_13_1150, i_13_1187, i_13_1270, i_13_1271, i_13_1437, i_13_1456, i_13_1462, i_13_1490, i_13_1518, i_13_1571, i_13_1594, i_13_1655, i_13_1747, i_13_1748, i_13_1750, i_13_1751, i_13_1805, i_13_1806, i_13_1815, i_13_1841, i_13_1856, i_13_1858, i_13_1909, i_13_1914, i_13_2047, i_13_2049, i_13_2112, i_13_2137, i_13_2138, i_13_2139, i_13_2140, i_13_2141, i_13_2224, i_13_2354, i_13_2357, i_13_2407, i_13_2408, i_13_2557, i_13_2562, i_13_2579, i_13_2650, i_13_2651, i_13_2652, i_13_2692, i_13_2722, i_13_2749, i_13_2750, i_13_2751, i_13_2752, i_13_2822, i_13_2823, i_13_2939, i_13_2999, i_13_3206, i_13_3208, i_13_3273, i_13_3290, i_13_3374, i_13_3430, i_13_3449, i_13_3533, i_13_3534, i_13_3556, i_13_3876, i_13_3911, i_13_3912, i_13_3943, i_13_3989, i_13_3991, i_13_4048, i_13_4161, i_13_4187, i_13_4309, i_13_4369, i_13_4381, i_13_4426, o_13_230);
	kernel_13_231 k_13_231(i_13_76, i_13_106, i_13_107, i_13_139, i_13_170, i_13_229, i_13_232, i_13_269, i_13_313, i_13_340, i_13_357, i_13_395, i_13_510, i_13_515, i_13_524, i_13_667, i_13_691, i_13_695, i_13_817, i_13_818, i_13_820, i_13_911, i_13_980, i_13_1069, i_13_1070, i_13_1208, i_13_1217, i_13_1222, i_13_1307, i_13_1316, i_13_1329, i_13_1330, i_13_1489, i_13_1573, i_13_1750, i_13_1807, i_13_1808, i_13_1815, i_13_1852, i_13_1882, i_13_1912, i_13_1999, i_13_2000, i_13_2059, i_13_2125, i_13_2126, i_13_2135, i_13_2139, i_13_2140, i_13_2185, i_13_2188, i_13_2225, i_13_2380, i_13_2409, i_13_2410, i_13_2411, i_13_2536, i_13_2586, i_13_2614, i_13_2656, i_13_2698, i_13_2722, i_13_2744, i_13_2751, i_13_2752, i_13_2797, i_13_2941, i_13_3003, i_13_3208, i_13_3220, i_13_3237, i_13_3238, i_13_3269, i_13_3273, i_13_3291, i_13_3292, i_13_3346, i_13_3372, i_13_3373, i_13_3505, i_13_3532, i_13_3538, i_13_3539, i_13_3727, i_13_3728, i_13_3853, i_13_3877, i_13_3895, i_13_3910, i_13_4021, i_13_4048, i_13_4063, i_13_4065, i_13_4066, i_13_4088, i_13_4252, i_13_4274, i_13_4318, i_13_4319, i_13_4448, o_13_231);
	kernel_13_232 k_13_232(i_13_39, i_13_40, i_13_43, i_13_105, i_13_114, i_13_186, i_13_187, i_13_373, i_13_445, i_13_529, i_13_533, i_13_547, i_13_556, i_13_573, i_13_600, i_13_607, i_13_629, i_13_682, i_13_717, i_13_732, i_13_780, i_13_817, i_13_897, i_13_940, i_13_1069, i_13_1084, i_13_1123, i_13_1159, i_13_1210, i_13_1266, i_13_1276, i_13_1464, i_13_1465, i_13_1482, i_13_1483, i_13_1501, i_13_1502, i_13_1645, i_13_1677, i_13_1690, i_13_1732, i_13_1749, i_13_1750, i_13_1752, i_13_1753, i_13_1770, i_13_1776, i_13_1788, i_13_1806, i_13_1807, i_13_1826, i_13_1862, i_13_1914, i_13_2051, i_13_2122, i_13_2139, i_13_2140, i_13_2149, i_13_2266, i_13_2310, i_13_2365, i_13_2582, i_13_2653, i_13_2722, i_13_2751, i_13_2752, i_13_2823, i_13_2824, i_13_2874, i_13_2883, i_13_2940, i_13_2941, i_13_2983, i_13_3030, i_13_3032, i_13_3119, i_13_3121, i_13_3122, i_13_3293, i_13_3345, i_13_3373, i_13_3400, i_13_3417, i_13_3418, i_13_3471, i_13_3525, i_13_3526, i_13_3562, i_13_3864, i_13_3895, i_13_3994, i_13_4047, i_13_4049, i_13_4080, i_13_4101, i_13_4156, i_13_4272, i_13_4318, i_13_4381, i_13_4443, o_13_232);
	kernel_13_233 k_13_233(i_13_48, i_13_165, i_13_211, i_13_217, i_13_441, i_13_531, i_13_532, i_13_558, i_13_570, i_13_640, i_13_676, i_13_679, i_13_837, i_13_928, i_13_931, i_13_945, i_13_1098, i_13_1117, i_13_1270, i_13_1380, i_13_1381, i_13_1396, i_13_1399, i_13_1434, i_13_1471, i_13_1530, i_13_1593, i_13_1657, i_13_1674, i_13_1719, i_13_1746, i_13_1777, i_13_1791, i_13_1792, i_13_1795, i_13_1908, i_13_1917, i_13_1930, i_13_2011, i_13_2016, i_13_2046, i_13_2115, i_13_2191, i_13_2259, i_13_2397, i_13_2466, i_13_2505, i_13_2673, i_13_2722, i_13_2748, i_13_2749, i_13_2818, i_13_2844, i_13_2857, i_13_2901, i_13_2911, i_13_2916, i_13_3024, i_13_3025, i_13_3060, i_13_3069, i_13_3090, i_13_3258, i_13_3348, i_13_3349, i_13_3375, i_13_3414, i_13_3415, i_13_3421, i_13_3532, i_13_3573, i_13_3685, i_13_3735, i_13_3765, i_13_3766, i_13_3783, i_13_3784, i_13_3846, i_13_3855, i_13_3862, i_13_3888, i_13_3924, i_13_3925, i_13_3987, i_13_3988, i_13_4054, i_13_4077, i_13_4086, i_13_4122, i_13_4123, i_13_4203, i_13_4204, i_13_4212, i_13_4447, i_13_4590, i_13_4591, i_13_4594, i_13_4599, i_13_4600, i_13_4604, o_13_233);
	kernel_13_234 k_13_234(i_13_81, i_13_137, i_13_140, i_13_142, i_13_143, i_13_166, i_13_232, i_13_279, i_13_280, i_13_355, i_13_454, i_13_534, i_13_539, i_13_582, i_13_595, i_13_603, i_13_611, i_13_620, i_13_691, i_13_700, i_13_725, i_13_726, i_13_780, i_13_824, i_13_894, i_13_1215, i_13_1222, i_13_1276, i_13_1277, i_13_1486, i_13_1498, i_13_1552, i_13_1678, i_13_1710, i_13_1711, i_13_1714, i_13_1715, i_13_1722, i_13_1725, i_13_1726, i_13_1727, i_13_1731, i_13_1761, i_13_1780, i_13_1781, i_13_1846, i_13_1881, i_13_1884, i_13_1885, i_13_1886, i_13_1888, i_13_1889, i_13_1999, i_13_2009, i_13_2158, i_13_2380, i_13_2461, i_13_2462, i_13_2470, i_13_2629, i_13_2647, i_13_2650, i_13_2651, i_13_2714, i_13_2848, i_13_2849, i_13_2875, i_13_2878, i_13_2887, i_13_2916, i_13_2917, i_13_3004, i_13_3040, i_13_3041, i_13_3109, i_13_3145, i_13_3146, i_13_3293, i_13_3406, i_13_3429, i_13_3689, i_13_3707, i_13_3781, i_13_3794, i_13_3964, i_13_4083, i_13_4095, i_13_4096, i_13_4100, i_13_4153, i_13_4190, i_13_4253, i_13_4390, i_13_4414, i_13_4426, i_13_4437, i_13_4440, i_13_4513, i_13_4519, i_13_4526, o_13_234);
	kernel_13_235 k_13_235(i_13_67, i_13_68, i_13_70, i_13_97, i_13_173, i_13_233, i_13_234, i_13_311, i_13_319, i_13_349, i_13_389, i_13_412, i_13_444, i_13_534, i_13_538, i_13_539, i_13_643, i_13_644, i_13_646, i_13_682, i_13_797, i_13_841, i_13_898, i_13_930, i_13_932, i_13_938, i_13_1105, i_13_1120, i_13_1121, i_13_1222, i_13_1259, i_13_1274, i_13_1281, i_13_1390, i_13_1391, i_13_1400, i_13_1428, i_13_1461, i_13_1491, i_13_1511, i_13_1512, i_13_1552, i_13_1642, i_13_1733, i_13_1765, i_13_1795, i_13_1796, i_13_1798, i_13_1804, i_13_1867, i_13_1881, i_13_1886, i_13_1924, i_13_1945, i_13_1946, i_13_2017, i_13_2021, i_13_2032, i_13_2056, i_13_2142, i_13_2315, i_13_2461, i_13_2542, i_13_2594, i_13_2678, i_13_2847, i_13_2848, i_13_2849, i_13_2878, i_13_2884, i_13_2966, i_13_3040, i_13_3075, i_13_3101, i_13_3172, i_13_3176, i_13_3367, i_13_3523, i_13_3730, i_13_3736, i_13_3740, i_13_3757, i_13_3784, i_13_3889, i_13_3910, i_13_3928, i_13_3930, i_13_3931, i_13_4038, i_13_4186, i_13_4187, i_13_4189, i_13_4294, i_13_4297, i_13_4303, i_13_4351, i_13_4453, i_13_4595, i_13_4597, i_13_4606, o_13_235);
	kernel_13_236 k_13_236(i_13_76, i_13_77, i_13_79, i_13_94, i_13_116, i_13_251, i_13_329, i_13_431, i_13_450, i_13_494, i_13_518, i_13_571, i_13_604, i_13_605, i_13_619, i_13_658, i_13_670, i_13_697, i_13_698, i_13_700, i_13_845, i_13_928, i_13_940, i_13_1024, i_13_1078, i_13_1079, i_13_1081, i_13_1082, i_13_1213, i_13_1276, i_13_1277, i_13_1317, i_13_1318, i_13_1341, i_13_1408, i_13_1427, i_13_1429, i_13_1430, i_13_1444, i_13_1573, i_13_1629, i_13_1637, i_13_1711, i_13_1731, i_13_1736, i_13_1781, i_13_1888, i_13_2027, i_13_2029, i_13_2060, i_13_2104, i_13_2198, i_13_2209, i_13_2236, i_13_2448, i_13_2453, i_13_2455, i_13_2511, i_13_2617, i_13_2632, i_13_2710, i_13_2726, i_13_2764, i_13_2809, i_13_2821, i_13_2854, i_13_2887, i_13_2888, i_13_2959, i_13_2986, i_13_3061, i_13_3208, i_13_3343, i_13_3392, i_13_3419, i_13_3452, i_13_3454, i_13_3460, i_13_3464, i_13_3490, i_13_3536, i_13_3571, i_13_3572, i_13_3593, i_13_3601, i_13_3662, i_13_3688, i_13_3717, i_13_3847, i_13_3850, i_13_4009, i_13_4063, i_13_4087, i_13_4094, i_13_4252, i_13_4264, i_13_4267, i_13_4330, i_13_4365, i_13_4562, o_13_236);
	kernel_13_237 k_13_237(i_13_97, i_13_106, i_13_125, i_13_134, i_13_233, i_13_358, i_13_376, i_13_409, i_13_512, i_13_529, i_13_530, i_13_573, i_13_574, i_13_575, i_13_607, i_13_718, i_13_799, i_13_800, i_13_845, i_13_1101, i_13_1304, i_13_1322, i_13_1410, i_13_1447, i_13_1492, i_13_1493, i_13_1501, i_13_1502, i_13_1511, i_13_1538, i_13_1543, i_13_1555, i_13_1556, i_13_1642, i_13_1643, i_13_1711, i_13_1744, i_13_1760, i_13_1796, i_13_1840, i_13_1933, i_13_1951, i_13_1990, i_13_1991, i_13_2015, i_13_2104, i_13_2239, i_13_2240, i_13_2246, i_13_2266, i_13_2318, i_13_2362, i_13_2428, i_13_2429, i_13_2458, i_13_2483, i_13_2536, i_13_2825, i_13_2906, i_13_2935, i_13_2936, i_13_2938, i_13_2947, i_13_2971, i_13_2983, i_13_3028, i_13_3065, i_13_3100, i_13_3117, i_13_3127, i_13_3207, i_13_3208, i_13_3244, i_13_3245, i_13_3425, i_13_3427, i_13_3428, i_13_3455, i_13_3478, i_13_3544, i_13_3722, i_13_3788, i_13_3794, i_13_3806, i_13_3859, i_13_3860, i_13_3914, i_13_3968, i_13_3985, i_13_4012, i_13_4013, i_13_4120, i_13_4219, i_13_4308, i_13_4313, i_13_4433, i_13_4444, i_13_4541, i_13_4567, i_13_4588, o_13_237);
	kernel_13_238 k_13_238(i_13_49, i_13_93, i_13_117, i_13_180, i_13_181, i_13_183, i_13_184, i_13_190, i_13_193, i_13_381, i_13_382, i_13_489, i_13_527, i_13_531, i_13_567, i_13_589, i_13_621, i_13_624, i_13_689, i_13_712, i_13_713, i_13_715, i_13_858, i_13_948, i_13_1099, i_13_1116, i_13_1117, i_13_1146, i_13_1219, i_13_1225, i_13_1251, i_13_1254, i_13_1255, i_13_1280, i_13_1387, i_13_1404, i_13_1407, i_13_1408, i_13_1488, i_13_1489, i_13_1512, i_13_1513, i_13_1677, i_13_1680, i_13_1760, i_13_1765, i_13_1786, i_13_1792, i_13_1801, i_13_1857, i_13_1862, i_13_1991, i_13_2002, i_13_2123, i_13_2242, i_13_2263, i_13_2281, i_13_2314, i_13_2533, i_13_2690, i_13_2836, i_13_2848, i_13_2856, i_13_2857, i_13_2908, i_13_2967, i_13_3025, i_13_3064, i_13_3126, i_13_3148, i_13_3153, i_13_3260, i_13_3262, i_13_3348, i_13_3352, i_13_3427, i_13_3456, i_13_3466, i_13_3478, i_13_3486, i_13_3489, i_13_3612, i_13_3638, i_13_3685, i_13_3699, i_13_3753, i_13_3754, i_13_3756, i_13_3757, i_13_3762, i_13_3874, i_13_3890, i_13_3978, i_13_4045, i_13_4261, i_13_4404, i_13_4509, i_13_4510, i_13_4538, i_13_4563, o_13_238);
	kernel_13_239 k_13_239(i_13_24, i_13_44, i_13_66, i_13_112, i_13_115, i_13_183, i_13_210, i_13_268, i_13_357, i_13_391, i_13_465, i_13_466, i_13_527, i_13_529, i_13_552, i_13_591, i_13_744, i_13_762, i_13_795, i_13_831, i_13_859, i_13_1083, i_13_1084, i_13_1131, i_13_1302, i_13_1303, i_13_1321, i_13_1419, i_13_1434, i_13_1474, i_13_1565, i_13_1597, i_13_1605, i_13_1607, i_13_1627, i_13_1677, i_13_1753, i_13_1806, i_13_1842, i_13_1843, i_13_1849, i_13_1914, i_13_1960, i_13_2029, i_13_2139, i_13_2145, i_13_2202, i_13_2203, i_13_2239, i_13_2284, i_13_2397, i_13_2401, i_13_2472, i_13_2506, i_13_2544, i_13_2545, i_13_2553, i_13_2578, i_13_2699, i_13_2704, i_13_2759, i_13_2762, i_13_2824, i_13_3003, i_13_3075, i_13_3092, i_13_3166, i_13_3243, i_13_3326, i_13_3345, i_13_3346, i_13_3373, i_13_3391, i_13_3477, i_13_3481, i_13_3579, i_13_3597, i_13_3633, i_13_3669, i_13_3724, i_13_3768, i_13_3805, i_13_3823, i_13_3859, i_13_3860, i_13_3894, i_13_3939, i_13_4038, i_13_4099, i_13_4164, i_13_4254, i_13_4264, i_13_4265, i_13_4272, i_13_4309, i_13_4315, i_13_4380, i_13_4381, i_13_4452, i_13_4453, o_13_239);
	kernel_13_240 k_13_240(i_13_65, i_13_131, i_13_163, i_13_252, i_13_256, i_13_266, i_13_269, i_13_272, i_13_308, i_13_340, i_13_354, i_13_379, i_13_380, i_13_458, i_13_463, i_13_466, i_13_467, i_13_475, i_13_535, i_13_592, i_13_684, i_13_821, i_13_829, i_13_895, i_13_1116, i_13_1120, i_13_1121, i_13_1307, i_13_1397, i_13_1444, i_13_1448, i_13_1467, i_13_1480, i_13_1496, i_13_1553, i_13_1594, i_13_1595, i_13_1697, i_13_1710, i_13_1723, i_13_1802, i_13_1844, i_13_1846, i_13_1847, i_13_1885, i_13_1908, i_13_1927, i_13_1928, i_13_1958, i_13_1989, i_13_1991, i_13_2101, i_13_2108, i_13_2261, i_13_2297, i_13_2366, i_13_2650, i_13_2677, i_13_2848, i_13_2849, i_13_2871, i_13_2935, i_13_2936, i_13_3035, i_13_3050, i_13_3167, i_13_3232, i_13_3241, i_13_3242, i_13_3415, i_13_3447, i_13_3519, i_13_3523, i_13_3569, i_13_3597, i_13_3598, i_13_3667, i_13_3730, i_13_3818, i_13_3857, i_13_3859, i_13_4017, i_13_4052, i_13_4060, i_13_4061, i_13_4063, i_13_4088, i_13_4165, i_13_4187, i_13_4189, i_13_4204, i_13_4205, i_13_4214, i_13_4267, i_13_4268, i_13_4313, i_13_4413, i_13_4430, i_13_4530, i_13_4562, o_13_240);
	kernel_13_241 k_13_241(i_13_69, i_13_101, i_13_230, i_13_326, i_13_336, i_13_379, i_13_505, i_13_573, i_13_578, i_13_623, i_13_641, i_13_690, i_13_717, i_13_780, i_13_1063, i_13_1064, i_13_1297, i_13_1298, i_13_1342, i_13_1410, i_13_1499, i_13_1529, i_13_1609, i_13_1627, i_13_1635, i_13_1712, i_13_1723, i_13_1777, i_13_1778, i_13_1801, i_13_1802, i_13_1810, i_13_1900, i_13_1906, i_13_1939, i_13_1990, i_13_1991, i_13_1993, i_13_2003, i_13_2012, i_13_2107, i_13_2134, i_13_2135, i_13_2209, i_13_2260, i_13_2261, i_13_2302, i_13_2309, i_13_2341, i_13_2359, i_13_2396, i_13_2404, i_13_2512, i_13_2522, i_13_2576, i_13_2614, i_13_2648, i_13_2746, i_13_2859, i_13_2935, i_13_2936, i_13_2939, i_13_2980, i_13_3012, i_13_3037, i_13_3143, i_13_3213, i_13_3286, i_13_3287, i_13_3340, i_13_3385, i_13_3386, i_13_3416, i_13_3421, i_13_3466, i_13_3476, i_13_3532, i_13_3642, i_13_3665, i_13_3729, i_13_3739, i_13_3747, i_13_3791, i_13_3876, i_13_4009, i_13_4011, i_13_4012, i_13_4015, i_13_4043, i_13_4055, i_13_4209, i_13_4230, i_13_4231, i_13_4232, i_13_4393, i_13_4398, i_13_4412, i_13_4531, i_13_4533, i_13_4587, o_13_241);
	kernel_13_242 k_13_242(i_13_94, i_13_121, i_13_229, i_13_230, i_13_232, i_13_518, i_13_520, i_13_521, i_13_535, i_13_645, i_13_661, i_13_739, i_13_756, i_13_820, i_13_850, i_13_851, i_13_870, i_13_938, i_13_1072, i_13_1073, i_13_1075, i_13_1201, i_13_1219, i_13_1262, i_13_1423, i_13_1424, i_13_1549, i_13_1550, i_13_1624, i_13_1630, i_13_1723, i_13_1758, i_13_1774, i_13_1787, i_13_1858, i_13_1939, i_13_1970, i_13_2027, i_13_2029, i_13_2033, i_13_2201, i_13_2209, i_13_2425, i_13_2451, i_13_2452, i_13_2454, i_13_2455, i_13_2558, i_13_2567, i_13_2612, i_13_2693, i_13_2764, i_13_2848, i_13_2850, i_13_3010, i_13_3011, i_13_3014, i_13_3037, i_13_3040, i_13_3143, i_13_3163, i_13_3217, i_13_3251, i_13_3272, i_13_3424, i_13_3442, i_13_3467, i_13_3472, i_13_3473, i_13_3485, i_13_3487, i_13_3488, i_13_3539, i_13_3541, i_13_3575, i_13_3731, i_13_3784, i_13_3853, i_13_3856, i_13_3863, i_13_3866, i_13_3893, i_13_3991, i_13_4038, i_13_4210, i_13_4216, i_13_4252, i_13_4253, i_13_4261, i_13_4262, i_13_4264, i_13_4265, i_13_4355, i_13_4370, i_13_4372, i_13_4379, i_13_4380, i_13_4511, i_13_4540, i_13_4558, o_13_242);
	kernel_13_243 k_13_243(i_13_37, i_13_77, i_13_104, i_13_112, i_13_117, i_13_337, i_13_379, i_13_451, i_13_452, i_13_461, i_13_561, i_13_583, i_13_586, i_13_589, i_13_643, i_13_676, i_13_724, i_13_769, i_13_914, i_13_949, i_13_950, i_13_1062, i_13_1064, i_13_1208, i_13_1243, i_13_1270, i_13_1297, i_13_1341, i_13_1342, i_13_1423, i_13_1427, i_13_1441, i_13_1495, i_13_1516, i_13_1594, i_13_1633, i_13_1693, i_13_1764, i_13_1811, i_13_1893, i_13_1945, i_13_2003, i_13_2099, i_13_2107, i_13_2108, i_13_2147, i_13_2197, i_13_2233, i_13_2234, i_13_2278, i_13_2542, i_13_2615, i_13_2650, i_13_2705, i_13_2710, i_13_2765, i_13_2782, i_13_2854, i_13_2898, i_13_2917, i_13_2918, i_13_2921, i_13_2926, i_13_3016, i_13_3017, i_13_3037, i_13_3064, i_13_3092, i_13_3136, i_13_3154, i_13_3199, i_13_3215, i_13_3218, i_13_3232, i_13_3289, i_13_3367, i_13_3415, i_13_3416, i_13_3532, i_13_3593, i_13_3739, i_13_3818, i_13_3874, i_13_3925, i_13_4019, i_13_4051, i_13_4087, i_13_4088, i_13_4106, i_13_4231, i_13_4232, i_13_4234, i_13_4250, i_13_4258, i_13_4267, i_13_4268, i_13_4393, i_13_4394, i_13_4448, i_13_4591, o_13_243);
	kernel_13_244 k_13_244(i_13_37, i_13_53, i_13_61, i_13_180, i_13_227, i_13_279, i_13_280, i_13_325, i_13_414, i_13_558, i_13_595, i_13_598, i_13_642, i_13_670, i_13_690, i_13_777, i_13_794, i_13_846, i_13_847, i_13_848, i_13_855, i_13_1073, i_13_1225, i_13_1252, i_13_1302, i_13_1314, i_13_1322, i_13_1404, i_13_1405, i_13_1444, i_13_1465, i_13_1479, i_13_1481, i_13_1483, i_13_1486, i_13_1548, i_13_1549, i_13_1574, i_13_1660, i_13_1746, i_13_1749, i_13_1776, i_13_1807, i_13_1854, i_13_1855, i_13_1856, i_13_1857, i_13_1858, i_13_1954, i_13_2022, i_13_2113, i_13_2134, i_13_2278, i_13_2281, i_13_2304, i_13_2307, i_13_2310, i_13_2311, i_13_2457, i_13_2458, i_13_2459, i_13_2553, i_13_2610, i_13_2629, i_13_2630, i_13_2636, i_13_2710, i_13_2877, i_13_2926, i_13_2937, i_13_3007, i_13_3019, i_13_3097, i_13_3129, i_13_3169, i_13_3170, i_13_3429, i_13_3448, i_13_3539, i_13_3579, i_13_3633, i_13_3741, i_13_3781, i_13_3791, i_13_3853, i_13_3907, i_13_3908, i_13_3910, i_13_3915, i_13_3987, i_13_4036, i_13_4059, i_13_4237, i_13_4267, i_13_4374, i_13_4375, i_13_4378, i_13_4381, i_13_4413, i_13_4518, o_13_244);
	kernel_13_245 k_13_245(i_13_41, i_13_45, i_13_46, i_13_59, i_13_163, i_13_213, i_13_234, i_13_236, i_13_241, i_13_274, i_13_333, i_13_355, i_13_370, i_13_384, i_13_450, i_13_453, i_13_457, i_13_535, i_13_586, i_13_612, i_13_810, i_13_816, i_13_832, i_13_894, i_13_954, i_13_956, i_13_1219, i_13_1342, i_13_1459, i_13_1509, i_13_1521, i_13_1522, i_13_1524, i_13_1551, i_13_1552, i_13_1568, i_13_1696, i_13_1750, i_13_1765, i_13_1767, i_13_1891, i_13_1903, i_13_1927, i_13_2121, i_13_2142, i_13_2143, i_13_2144, i_13_2296, i_13_2394, i_13_2461, i_13_2560, i_13_2565, i_13_2568, i_13_2613, i_13_2691, i_13_2715, i_13_2716, i_13_2764, i_13_2766, i_13_2781, i_13_2782, i_13_2845, i_13_2881, i_13_2935, i_13_3028, i_13_3108, i_13_3142, i_13_3145, i_13_3146, i_13_3207, i_13_3231, i_13_3238, i_13_3274, i_13_3342, i_13_3366, i_13_3382, i_13_3546, i_13_3636, i_13_3754, i_13_3836, i_13_3856, i_13_3889, i_13_3900, i_13_3902, i_13_3916, i_13_3921, i_13_3982, i_13_4017, i_13_4052, i_13_4081, i_13_4086, i_13_4249, i_13_4269, i_13_4270, i_13_4311, i_13_4312, i_13_4428, i_13_4509, i_13_4510, i_13_4533, o_13_245);
	kernel_13_246 k_13_246(i_13_53, i_13_76, i_13_77, i_13_116, i_13_166, i_13_184, i_13_193, i_13_203, i_13_446, i_13_530, i_13_554, i_13_561, i_13_571, i_13_592, i_13_655, i_13_656, i_13_671, i_13_697, i_13_698, i_13_700, i_13_826, i_13_944, i_13_1084, i_13_1085, i_13_1147, i_13_1148, i_13_1211, i_13_1223, i_13_1267, i_13_1285, i_13_1430, i_13_1502, i_13_1508, i_13_1517, i_13_1525, i_13_1552, i_13_1636, i_13_1637, i_13_1660, i_13_1661, i_13_1664, i_13_1741, i_13_1831, i_13_1840, i_13_1843, i_13_1844, i_13_1885, i_13_1886, i_13_2033, i_13_2172, i_13_2245, i_13_2314, i_13_2321, i_13_2354, i_13_2398, i_13_2438, i_13_2455, i_13_2456, i_13_2510, i_13_2762, i_13_2848, i_13_2849, i_13_2887, i_13_2924, i_13_2959, i_13_2983, i_13_3001, i_13_3002, i_13_3004, i_13_3050, i_13_3130, i_13_3383, i_13_3436, i_13_3467, i_13_3476, i_13_3505, i_13_3571, i_13_3572, i_13_3599, i_13_3602, i_13_3649, i_13_3650, i_13_3689, i_13_3740, i_13_3742, i_13_3866, i_13_3875, i_13_4021, i_13_4045, i_13_4063, i_13_4190, i_13_4264, i_13_4279, i_13_4301, i_13_4333, i_13_4378, i_13_4417, i_13_4594, i_13_4603, i_13_4604, o_13_246);
	kernel_13_247 k_13_247(i_13_74, i_13_91, i_13_94, i_13_103, i_13_104, i_13_109, i_13_112, i_13_118, i_13_166, i_13_201, i_13_263, i_13_364, i_13_607, i_13_643, i_13_730, i_13_733, i_13_768, i_13_793, i_13_794, i_13_856, i_13_946, i_13_1084, i_13_1086, i_13_1102, i_13_1144, i_13_1217, i_13_1273, i_13_1486, i_13_1487, i_13_1552, i_13_1621, i_13_1630, i_13_1692, i_13_1774, i_13_1775, i_13_1836, i_13_1837, i_13_1839, i_13_1846, i_13_2000, i_13_2009, i_13_2137, i_13_2170, i_13_2172, i_13_2173, i_13_2201, i_13_2381, i_13_2407, i_13_2422, i_13_2430, i_13_2431, i_13_2434, i_13_2497, i_13_2498, i_13_2539, i_13_2542, i_13_2569, i_13_2579, i_13_2611, i_13_2875, i_13_2943, i_13_2958, i_13_3024, i_13_3054, i_13_3100, i_13_3143, i_13_3145, i_13_3146, i_13_3370, i_13_3375, i_13_3452, i_13_3525, i_13_3529, i_13_3530, i_13_3646, i_13_3696, i_13_3739, i_13_3864, i_13_3871, i_13_3872, i_13_3891, i_13_4036, i_13_4063, i_13_4091, i_13_4106, i_13_4118, i_13_4119, i_13_4122, i_13_4234, i_13_4252, i_13_4263, i_13_4339, i_13_4351, i_13_4367, i_13_4413, i_13_4417, i_13_4431, i_13_4542, i_13_4559, i_13_4560, o_13_247);
	kernel_13_248 k_13_248(i_13_97, i_13_154, i_13_164, i_13_217, i_13_251, i_13_272, i_13_319, i_13_355, i_13_451, i_13_559, i_13_688, i_13_895, i_13_928, i_13_929, i_13_966, i_13_974, i_13_1081, i_13_1099, i_13_1120, i_13_1252, i_13_1262, i_13_1283, i_13_1298, i_13_1340, i_13_1372, i_13_1396, i_13_1397, i_13_1468, i_13_1502, i_13_1505, i_13_1568, i_13_1606, i_13_1628, i_13_1633, i_13_1786, i_13_1811, i_13_1855, i_13_1858, i_13_1891, i_13_1910, i_13_1928, i_13_1990, i_13_2003, i_13_2108, i_13_2117, i_13_2180, i_13_2234, i_13_2314, i_13_2333, i_13_2430, i_13_2467, i_13_2483, i_13_2542, i_13_2543, i_13_2696, i_13_2711, i_13_2755, i_13_2764, i_13_2765, i_13_2785, i_13_2786, i_13_2935, i_13_2936, i_13_2958, i_13_3016, i_13_3017, i_13_3061, i_13_3062, i_13_3206, i_13_3218, i_13_3231, i_13_3234, i_13_3239, i_13_3242, i_13_3271, i_13_3312, i_13_3313, i_13_3340, i_13_3341, i_13_3532, i_13_3601, i_13_3683, i_13_3709, i_13_3723, i_13_3851, i_13_3920, i_13_4081, i_13_4082, i_13_4087, i_13_4160, i_13_4214, i_13_4266, i_13_4268, i_13_4313, i_13_4361, i_13_4430, i_13_4453, i_13_4462, i_13_4466, i_13_4595, o_13_248);
	kernel_13_249 k_13_249(i_13_34, i_13_47, i_13_139, i_13_143, i_13_184, i_13_233, i_13_380, i_13_383, i_13_385, i_13_386, i_13_529, i_13_649, i_13_666, i_13_675, i_13_701, i_13_763, i_13_824, i_13_871, i_13_883, i_13_985, i_13_1082, i_13_1206, i_13_1220, i_13_1281, i_13_1326, i_13_1403, i_13_1442, i_13_1445, i_13_1502, i_13_1511, i_13_1516, i_13_1600, i_13_1664, i_13_1678, i_13_1684, i_13_1750, i_13_1780, i_13_1787, i_13_1817, i_13_1861, i_13_1912, i_13_1930, i_13_2002, i_13_2003, i_13_2005, i_13_2006, i_13_2054, i_13_2177, i_13_2189, i_13_2196, i_13_2210, i_13_2246, i_13_2259, i_13_2266, i_13_2279, i_13_2351, i_13_2537, i_13_2543, i_13_2677, i_13_2708, i_13_2719, i_13_2722, i_13_2723, i_13_2725, i_13_2726, i_13_2854, i_13_2855, i_13_2858, i_13_2861, i_13_2969, i_13_3218, i_13_3347, i_13_3379, i_13_3392, i_13_3418, i_13_3419, i_13_3442, i_13_3577, i_13_3593, i_13_3614, i_13_3653, i_13_3686, i_13_3730, i_13_3844, i_13_3865, i_13_3873, i_13_3892, i_13_3917, i_13_4052, i_13_4057, i_13_4058, i_13_4171, i_13_4268, i_13_4273, i_13_4282, i_13_4345, i_13_4394, i_13_4400, i_13_4568, i_13_4583, o_13_249);
	kernel_13_250 k_13_250(i_13_47, i_13_65, i_13_169, i_13_170, i_13_319, i_13_438, i_13_463, i_13_524, i_13_538, i_13_623, i_13_659, i_13_667, i_13_848, i_13_937, i_13_938, i_13_1018, i_13_1019, i_13_1072, i_13_1073, i_13_1086, i_13_1095, i_13_1096, i_13_1100, i_13_1252, i_13_1253, i_13_1315, i_13_1365, i_13_1400, i_13_1428, i_13_1488, i_13_1550, i_13_1596, i_13_1662, i_13_1694, i_13_1778, i_13_1792, i_13_1825, i_13_1913, i_13_1947, i_13_2026, i_13_2027, i_13_2056, i_13_2103, i_13_2122, i_13_2197, i_13_2227, i_13_2360, i_13_2364, i_13_2373, i_13_2770, i_13_2910, i_13_2915, i_13_2918, i_13_2975, i_13_3001, i_13_3008, i_13_3010, i_13_3103, i_13_3120, i_13_3166, i_13_3265, i_13_3352, i_13_3353, i_13_3382, i_13_3432, i_13_3452, i_13_3454, i_13_3459, i_13_3484, i_13_3534, i_13_3538, i_13_3539, i_13_3574, i_13_3575, i_13_3727, i_13_3741, i_13_3781, i_13_3782, i_13_3783, i_13_3820, i_13_3840, i_13_3847, i_13_3853, i_13_3859, i_13_3893, i_13_3908, i_13_3918, i_13_4063, i_13_4108, i_13_4150, i_13_4250, i_13_4253, i_13_4259, i_13_4335, i_13_4336, i_13_4344, i_13_4448, i_13_4583, i_13_4604, i_13_4605, o_13_250);
	kernel_13_251 k_13_251(i_13_37, i_13_38, i_13_51, i_13_75, i_13_76, i_13_103, i_13_112, i_13_165, i_13_173, i_13_181, i_13_184, i_13_240, i_13_252, i_13_280, i_13_281, i_13_324, i_13_325, i_13_339, i_13_571, i_13_577, i_13_596, i_13_597, i_13_598, i_13_618, i_13_640, i_13_643, i_13_685, i_13_715, i_13_744, i_13_778, i_13_814, i_13_840, i_13_891, i_13_892, i_13_894, i_13_896, i_13_1031, i_13_1093, i_13_1248, i_13_1249, i_13_1462, i_13_1480, i_13_1541, i_13_1711, i_13_1746, i_13_1747, i_13_1786, i_13_1804, i_13_1805, i_13_1806, i_13_1854, i_13_1855, i_13_1856, i_13_1858, i_13_2119, i_13_2121, i_13_2137, i_13_2138, i_13_2165, i_13_2344, i_13_2360, i_13_2403, i_13_2452, i_13_2557, i_13_2559, i_13_2630, i_13_2647, i_13_2650, i_13_2719, i_13_2722, i_13_2749, i_13_2751, i_13_2821, i_13_2881, i_13_2896, i_13_2938, i_13_3019, i_13_3064, i_13_3205, i_13_3290, i_13_3325, i_13_3372, i_13_3430, i_13_3439, i_13_3520, i_13_3524, i_13_3525, i_13_3910, i_13_3919, i_13_3925, i_13_3926, i_13_3974, i_13_3987, i_13_3992, i_13_4032, i_13_4078, i_13_4183, i_13_4270, i_13_4294, i_13_4369, o_13_251);
	kernel_13_252 k_13_252(i_13_37, i_13_49, i_13_100, i_13_127, i_13_136, i_13_154, i_13_166, i_13_167, i_13_269, i_13_271, i_13_280, i_13_283, i_13_316, i_13_379, i_13_385, i_13_386, i_13_415, i_13_450, i_13_451, i_13_558, i_13_571, i_13_639, i_13_640, i_13_658, i_13_676, i_13_677, i_13_720, i_13_758, i_13_869, i_13_940, i_13_982, i_13_1062, i_13_1063, i_13_1082, i_13_1093, i_13_1210, i_13_1300, i_13_1324, i_13_1390, i_13_1423, i_13_1436, i_13_1494, i_13_1525, i_13_1567, i_13_1633, i_13_1714, i_13_1807, i_13_1850, i_13_1909, i_13_1991, i_13_2054, i_13_2107, i_13_2108, i_13_2116, i_13_2233, i_13_2234, i_13_2297, i_13_2313, i_13_2361, i_13_2398, i_13_2467, i_13_2507, i_13_2542, i_13_2547, i_13_2663, i_13_2692, i_13_2766, i_13_2848, i_13_2872, i_13_3016, i_13_3106, i_13_3107, i_13_3109, i_13_3110, i_13_3307, i_13_3406, i_13_3433, i_13_3522, i_13_3528, i_13_3646, i_13_3708, i_13_3763, i_13_3766, i_13_3768, i_13_3817, i_13_3818, i_13_3901, i_13_4015, i_13_4078, i_13_4087, i_13_4117, i_13_4207, i_13_4230, i_13_4259, i_13_4266, i_13_4267, i_13_4302, i_13_4510, i_13_4555, i_13_4564, o_13_252);
	kernel_13_253 k_13_253(i_13_93, i_13_94, i_13_112, i_13_121, i_13_165, i_13_192, i_13_193, i_13_199, i_13_225, i_13_504, i_13_531, i_13_570, i_13_571, i_13_588, i_13_639, i_13_714, i_13_715, i_13_729, i_13_814, i_13_891, i_13_927, i_13_948, i_13_999, i_13_1053, i_13_1200, i_13_1209, i_13_1210, i_13_1227, i_13_1317, i_13_1386, i_13_1407, i_13_1426, i_13_1467, i_13_1488, i_13_1512, i_13_1720, i_13_1764, i_13_1767, i_13_1782, i_13_1783, i_13_1785, i_13_1800, i_13_1801, i_13_1908, i_13_1990, i_13_1992, i_13_2011, i_13_2056, i_13_2109, i_13_2116, i_13_2128, i_13_2164, i_13_2206, i_13_2209, i_13_2225, i_13_2235, i_13_2452, i_13_2505, i_13_2532, i_13_2568, i_13_2623, i_13_2722, i_13_2875, i_13_2889, i_13_2934, i_13_3024, i_13_3046, i_13_3087, i_13_3154, i_13_3162, i_13_3163, i_13_3214, i_13_3286, i_13_3304, i_13_3375, i_13_3420, i_13_3421, i_13_3423, i_13_3451, i_13_3522, i_13_3753, i_13_3790, i_13_3873, i_13_3883, i_13_3918, i_13_3924, i_13_3981, i_13_4008, i_13_4009, i_13_4077, i_13_4167, i_13_4194, i_13_4212, i_13_4305, i_13_4320, i_13_4497, i_13_4530, i_13_4539, i_13_4584, i_13_4594, o_13_253);
	kernel_13_254 k_13_254(i_13_0, i_13_46, i_13_55, i_13_121, i_13_164, i_13_172, i_13_208, i_13_243, i_13_346, i_13_416, i_13_482, i_13_490, i_13_606, i_13_625, i_13_644, i_13_676, i_13_695, i_13_712, i_13_764, i_13_782, i_13_841, i_13_850, i_13_882, i_13_884, i_13_936, i_13_982, i_13_983, i_13_1242, i_13_1252, i_13_1263, i_13_1307, i_13_1484, i_13_1489, i_13_1507, i_13_1521, i_13_1525, i_13_1564, i_13_1570, i_13_1611, i_13_1643, i_13_1750, i_13_1751, i_13_1757, i_13_1841, i_13_1940, i_13_1943, i_13_1953, i_13_2024, i_13_2047, i_13_2097, i_13_2389, i_13_2443, i_13_2515, i_13_2539, i_13_2542, i_13_2605, i_13_2614, i_13_2692, i_13_2763, i_13_2782, i_13_2880, i_13_2963, i_13_3073, i_13_3077, i_13_3091, i_13_3106, i_13_3172, i_13_3261, i_13_3320, i_13_3352, i_13_3412, i_13_3566, i_13_3638, i_13_3657, i_13_3753, i_13_3781, i_13_3838, i_13_3845, i_13_3852, i_13_3865, i_13_3898, i_13_3983, i_13_3988, i_13_3991, i_13_3996, i_13_4036, i_13_4187, i_13_4214, i_13_4242, i_13_4270, i_13_4272, i_13_4295, i_13_4297, i_13_4307, i_13_4311, i_13_4375, i_13_4378, i_13_4511, i_13_4513, i_13_4603, o_13_254);
	kernel_13_255 k_13_255(i_13_0, i_13_1, i_13_136, i_13_298, i_13_326, i_13_364, i_13_544, i_13_550, i_13_568, i_13_625, i_13_626, i_13_712, i_13_730, i_13_847, i_13_850, i_13_901, i_13_941, i_13_1044, i_13_1125, i_13_1129, i_13_1225, i_13_1226, i_13_1252, i_13_1270, i_13_1279, i_13_1310, i_13_1480, i_13_1486, i_13_1522, i_13_1552, i_13_1584, i_13_1585, i_13_1604, i_13_1749, i_13_1765, i_13_1810, i_13_1828, i_13_1854, i_13_1891, i_13_2020, i_13_2098, i_13_2116, i_13_2119, i_13_2214, i_13_2395, i_13_2422, i_13_2566, i_13_2593, i_13_2642, i_13_2647, i_13_2740, i_13_2755, i_13_2803, i_13_2875, i_13_2876, i_13_2917, i_13_2971, i_13_2972, i_13_2974, i_13_3019, i_13_3044, i_13_3091, i_13_3100, i_13_3101, i_13_3115, i_13_3127, i_13_3133, i_13_3145, i_13_3190, i_13_3213, i_13_3214, i_13_3262, i_13_3304, i_13_3331, i_13_3380, i_13_3416, i_13_3460, i_13_3485, i_13_3573, i_13_3822, i_13_3853, i_13_3899, i_13_3916, i_13_3944, i_13_3964, i_13_3979, i_13_3981, i_13_4033, i_13_4078, i_13_4091, i_13_4160, i_13_4266, i_13_4270, i_13_4303, i_13_4320, i_13_4325, i_13_4460, i_13_4475, i_13_4504, i_13_4529, o_13_255);
	kernel_13_256 k_13_256(i_13_27, i_13_30, i_13_63, i_13_64, i_13_130, i_13_135, i_13_136, i_13_156, i_13_202, i_13_207, i_13_208, i_13_225, i_13_354, i_13_355, i_13_378, i_13_453, i_13_454, i_13_468, i_13_469, i_13_489, i_13_549, i_13_612, i_13_643, i_13_675, i_13_730, i_13_732, i_13_793, i_13_796, i_13_810, i_13_831, i_13_840, i_13_946, i_13_954, i_13_1021, i_13_1063, i_13_1120, i_13_1128, i_13_1273, i_13_1300, i_13_1344, i_13_1486, i_13_1522, i_13_1525, i_13_1620, i_13_1621, i_13_1677, i_13_1692, i_13_1696, i_13_1719, i_13_1720, i_13_1836, i_13_1846, i_13_2002, i_13_2100, i_13_2173, i_13_2296, i_13_2316, i_13_2340, i_13_2341, i_13_2421, i_13_2431, i_13_2538, i_13_2550, i_13_2676, i_13_2677, i_13_2694, i_13_2718, i_13_2719, i_13_2748, i_13_2880, i_13_2946, i_13_3033, i_13_3072, i_13_3109, i_13_3231, i_13_3241, i_13_3421, i_13_3466, i_13_3528, i_13_3594, i_13_3610, i_13_3618, i_13_3619, i_13_3636, i_13_3637, i_13_3666, i_13_3681, i_13_3726, i_13_3843, i_13_3982, i_13_4233, i_13_4261, i_13_4269, i_13_4279, i_13_4315, i_13_4329, i_13_4396, i_13_4509, i_13_4519, i_13_4537, o_13_256);
	kernel_13_257 k_13_257(i_13_171, i_13_172, i_13_174, i_13_175, i_13_279, i_13_280, i_13_283, i_13_465, i_13_472, i_13_523, i_13_525, i_13_562, i_13_612, i_13_657, i_13_661, i_13_793, i_13_820, i_13_822, i_13_823, i_13_847, i_13_849, i_13_1017, i_13_1071, i_13_1072, i_13_1224, i_13_1225, i_13_1227, i_13_1308, i_13_1309, i_13_1363, i_13_1422, i_13_1425, i_13_1485, i_13_1489, i_13_1494, i_13_1495, i_13_1549, i_13_1629, i_13_1641, i_13_1855, i_13_1858, i_13_1881, i_13_1999, i_13_2070, i_13_2190, i_13_2206, i_13_2314, i_13_2347, i_13_2422, i_13_2448, i_13_2449, i_13_2539, i_13_2658, i_13_2673, i_13_2676, i_13_2692, i_13_2746, i_13_3007, i_13_3009, i_13_3096, i_13_3133, i_13_3216, i_13_3235, i_13_3267, i_13_3268, i_13_3270, i_13_3271, i_13_3414, i_13_3420, i_13_3421, i_13_3423, i_13_3523, i_13_3537, i_13_3538, i_13_3540, i_13_3643, i_13_3730, i_13_3741, i_13_3781, i_13_3798, i_13_3834, i_13_4015, i_13_4080, i_13_4195, i_13_4248, i_13_4249, i_13_4251, i_13_4252, i_13_4257, i_13_4258, i_13_4260, i_13_4275, i_13_4293, i_13_4338, i_13_4351, i_13_4375, i_13_4381, i_13_4414, i_13_4494, i_13_4555, o_13_257);
	kernel_13_258 k_13_258(i_13_105, i_13_106, i_13_213, i_13_420, i_13_600, i_13_609, i_13_619, i_13_742, i_13_745, i_13_858, i_13_1024, i_13_1068, i_13_1069, i_13_1086, i_13_1087, i_13_1095, i_13_1347, i_13_1488, i_13_1500, i_13_1507, i_13_1518, i_13_1519, i_13_1536, i_13_1561, i_13_1570, i_13_1572, i_13_1795, i_13_1813, i_13_1860, i_13_1930, i_13_2058, i_13_2059, i_13_2095, i_13_2149, i_13_2265, i_13_2280, i_13_2380, i_13_2400, i_13_2496, i_13_2500, i_13_2541, i_13_2551, i_13_2598, i_13_2599, i_13_2617, i_13_2679, i_13_2707, i_13_2715, i_13_2751, i_13_2851, i_13_2938, i_13_2985, i_13_2986, i_13_3012, i_13_3019, i_13_3031, i_13_3067, i_13_3073, i_13_3147, i_13_3148, i_13_3210, i_13_3211, i_13_3217, i_13_3328, i_13_3343, i_13_3346, i_13_3388, i_13_3400, i_13_3417, i_13_3418, i_13_3453, i_13_3454, i_13_3478, i_13_3525, i_13_3526, i_13_3531, i_13_3532, i_13_3732, i_13_3769, i_13_3891, i_13_4020, i_13_4039, i_13_4047, i_13_4048, i_13_4093, i_13_4119, i_13_4120, i_13_4234, i_13_4236, i_13_4254, i_13_4270, i_13_4317, i_13_4327, i_13_4353, i_13_4396, i_13_4416, i_13_4417, i_13_4476, i_13_4543, i_13_4557, o_13_258);
	kernel_13_259 k_13_259(i_13_49, i_13_64, i_13_118, i_13_166, i_13_233, i_13_238, i_13_308, i_13_311, i_13_317, i_13_328, i_13_569, i_13_586, i_13_587, i_13_640, i_13_641, i_13_712, i_13_739, i_13_740, i_13_757, i_13_838, i_13_839, i_13_856, i_13_929, i_13_1017, i_13_1082, i_13_1201, i_13_1253, i_13_1324, i_13_1325, i_13_1350, i_13_1442, i_13_1468, i_13_1486, i_13_1505, i_13_1526, i_13_1550, i_13_1568, i_13_1830, i_13_1832, i_13_1908, i_13_1990, i_13_2002, i_13_2045, i_13_2053, i_13_2054, i_13_2056, i_13_2108, i_13_2117, i_13_2234, i_13_2245, i_13_2259, i_13_2260, i_13_2261, i_13_2263, i_13_2264, i_13_2277, i_13_2278, i_13_2279, i_13_2407, i_13_2709, i_13_2711, i_13_2722, i_13_2750, i_13_2855, i_13_2945, i_13_3037, i_13_3061, i_13_3064, i_13_3065, i_13_3109, i_13_3110, i_13_3288, i_13_3388, i_13_3438, i_13_3439, i_13_3476, i_13_3483, i_13_3611, i_13_3614, i_13_3688, i_13_3703, i_13_3757, i_13_3766, i_13_3817, i_13_3818, i_13_3901, i_13_3928, i_13_3993, i_13_4007, i_13_4033, i_13_4186, i_13_4187, i_13_4276, i_13_4303, i_13_4304, i_13_4306, i_13_4315, i_13_4339, i_13_4394, i_13_4601, o_13_259);
	kernel_13_260 k_13_260(i_13_20, i_13_39, i_13_64, i_13_65, i_13_73, i_13_173, i_13_356, i_13_357, i_13_379, i_13_406, i_13_443, i_13_469, i_13_526, i_13_527, i_13_530, i_13_667, i_13_668, i_13_676, i_13_677, i_13_695, i_13_700, i_13_758, i_13_829, i_13_830, i_13_838, i_13_839, i_13_853, i_13_854, i_13_947, i_13_949, i_13_950, i_13_1024, i_13_1099, i_13_1118, i_13_1397, i_13_1438, i_13_1487, i_13_1499, i_13_1505, i_13_1594, i_13_1658, i_13_1720, i_13_1742, i_13_1744, i_13_1751, i_13_1792, i_13_1883, i_13_1913, i_13_1928, i_13_1950, i_13_2030, i_13_2032, i_13_2224, i_13_2242, i_13_2341, i_13_2454, i_13_2467, i_13_2468, i_13_2512, i_13_2514, i_13_2692, i_13_2693, i_13_2720, i_13_2750, i_13_2764, i_13_2912, i_13_3010, i_13_3026, i_13_3044, i_13_3061, i_13_3062, i_13_3128, i_13_3134, i_13_3146, i_13_3370, i_13_3371, i_13_3373, i_13_3382, i_13_3533, i_13_3596, i_13_3597, i_13_3598, i_13_3620, i_13_3632, i_13_3633, i_13_3638, i_13_3733, i_13_3783, i_13_3860, i_13_3925, i_13_3926, i_13_3988, i_13_4264, i_13_4312, i_13_4330, i_13_4331, i_13_4332, i_13_4414, i_13_4430, i_13_4451, o_13_260);
	kernel_13_261 k_13_261(i_13_31, i_13_116, i_13_197, i_13_219, i_13_226, i_13_359, i_13_370, i_13_382, i_13_396, i_13_405, i_13_441, i_13_450, i_13_473, i_13_553, i_13_558, i_13_607, i_13_651, i_13_666, i_13_667, i_13_671, i_13_675, i_13_676, i_13_823, i_13_828, i_13_829, i_13_833, i_13_1062, i_13_1098, i_13_1116, i_13_1147, i_13_1148, i_13_1454, i_13_1492, i_13_1507, i_13_1530, i_13_1624, i_13_1642, i_13_1729, i_13_1754, i_13_1777, i_13_1795, i_13_1837, i_13_1840, i_13_1858, i_13_1908, i_13_1993, i_13_2020, i_13_2024, i_13_2045, i_13_2186, i_13_2280, i_13_2281, i_13_2307, i_13_2413, i_13_2431, i_13_2438, i_13_2456, i_13_2461, i_13_2466, i_13_2471, i_13_2709, i_13_2938, i_13_3097, i_13_3098, i_13_3104, i_13_3267, i_13_3388, i_13_3490, i_13_3505, i_13_3541, i_13_3599, i_13_3670, i_13_3725, i_13_3740, i_13_3753, i_13_3766, i_13_3769, i_13_3819, i_13_3910, i_13_3925, i_13_3987, i_13_4086, i_13_4096, i_13_4126, i_13_4158, i_13_4162, i_13_4165, i_13_4212, i_13_4213, i_13_4343, i_13_4354, i_13_4355, i_13_4394, i_13_4429, i_13_4433, i_13_4514, i_13_4540, i_13_4571, i_13_4590, i_13_4600, o_13_261);
	kernel_13_262 k_13_262(i_13_58, i_13_61, i_13_136, i_13_220, i_13_283, i_13_310, i_13_493, i_13_554, i_13_577, i_13_628, i_13_684, i_13_698, i_13_891, i_13_897, i_13_917, i_13_1071, i_13_1096, i_13_1111, i_13_1129, i_13_1142, i_13_1263, i_13_1271, i_13_1282, i_13_1299, i_13_1302, i_13_1304, i_13_1317, i_13_1321, i_13_1322, i_13_1380, i_13_1441, i_13_1462, i_13_1464, i_13_1480, i_13_1484, i_13_1498, i_13_1633, i_13_1673, i_13_1742, i_13_1756, i_13_1770, i_13_1774, i_13_1781, i_13_1796, i_13_1806, i_13_1840, i_13_1849, i_13_2002, i_13_2380, i_13_2382, i_13_2407, i_13_2409, i_13_2425, i_13_2442, i_13_2443, i_13_2446, i_13_2447, i_13_2498, i_13_2650, i_13_2749, i_13_2785, i_13_2820, i_13_2835, i_13_2871, i_13_2872, i_13_3035, i_13_3056, i_13_3093, i_13_3094, i_13_3113, i_13_3118, i_13_3145, i_13_3253, i_13_3311, i_13_3312, i_13_3356, i_13_3390, i_13_3418, i_13_3419, i_13_3516, i_13_3542, i_13_3766, i_13_3817, i_13_3855, i_13_3869, i_13_3887, i_13_3960, i_13_3963, i_13_3981, i_13_4018, i_13_4019, i_13_4026, i_13_4238, i_13_4336, i_13_4349, i_13_4377, i_13_4382, i_13_4407, i_13_4519, i_13_4567, o_13_262);
	kernel_13_263 k_13_263(i_13_104, i_13_124, i_13_169, i_13_197, i_13_203, i_13_217, i_13_382, i_13_383, i_13_590, i_13_607, i_13_619, i_13_626, i_13_718, i_13_719, i_13_838, i_13_862, i_13_863, i_13_932, i_13_952, i_13_1024, i_13_1025, i_13_1033, i_13_1147, i_13_1232, i_13_1243, i_13_1259, i_13_1301, i_13_1411, i_13_1412, i_13_1493, i_13_1529, i_13_1628, i_13_1711, i_13_1780, i_13_1786, i_13_1789, i_13_1814, i_13_1961, i_13_1990, i_13_1994, i_13_2006, i_13_2015, i_13_2021, i_13_2104, i_13_2126, i_13_2212, i_13_2213, i_13_2237, i_13_2246, i_13_2264, i_13_2434, i_13_2464, i_13_2465, i_13_2507, i_13_2536, i_13_2537, i_13_2545, i_13_2617, i_13_2618, i_13_2714, i_13_2923, i_13_2934, i_13_2938, i_13_2939, i_13_3040, i_13_3041, i_13_3176, i_13_3218, i_13_3220, i_13_3286, i_13_3290, i_13_3344, i_13_3388, i_13_3395, i_13_3424, i_13_3425, i_13_3467, i_13_3536, i_13_3613, i_13_3643, i_13_3644, i_13_3790, i_13_3796, i_13_3806, i_13_3865, i_13_3877, i_13_3878, i_13_4008, i_13_4012, i_13_4013, i_13_4022, i_13_4078, i_13_4091, i_13_4162, i_13_4333, i_13_4369, i_13_4410, i_13_4414, i_13_4534, i_13_4600, o_13_263);
	kernel_13_264 k_13_264(i_13_76, i_13_118, i_13_119, i_13_122, i_13_181, i_13_182, i_13_184, i_13_202, i_13_226, i_13_227, i_13_229, i_13_380, i_13_418, i_13_491, i_13_518, i_13_524, i_13_532, i_13_533, i_13_562, i_13_572, i_13_715, i_13_725, i_13_831, i_13_833, i_13_841, i_13_911, i_13_946, i_13_1046, i_13_1109, i_13_1112, i_13_1128, i_13_1226, i_13_1406, i_13_1523, i_13_1540, i_13_1690, i_13_1720, i_13_1721, i_13_1723, i_13_1757, i_13_1783, i_13_1784, i_13_1786, i_13_1787, i_13_1837, i_13_1838, i_13_1921, i_13_1940, i_13_1967, i_13_2054, i_13_2056, i_13_2110, i_13_2116, i_13_2120, i_13_2165, i_13_2206, i_13_2207, i_13_2210, i_13_2213, i_13_2225, i_13_2236, i_13_2295, i_13_2426, i_13_2563, i_13_2579, i_13_2630, i_13_2639, i_13_2786, i_13_3010, i_13_3020, i_13_3037, i_13_3044, i_13_3163, i_13_3164, i_13_3214, i_13_3260, i_13_3278, i_13_3422, i_13_3425, i_13_3524, i_13_3533, i_13_3700, i_13_3791, i_13_3836, i_13_3871, i_13_3872, i_13_3874, i_13_3884, i_13_3919, i_13_3983, i_13_4010, i_13_4087, i_13_4111, i_13_4258, i_13_4276, i_13_4448, i_13_4519, i_13_4531, i_13_4537, i_13_4583, o_13_264);
	kernel_13_265 k_13_265(i_13_64, i_13_94, i_13_183, i_13_184, i_13_279, i_13_280, i_13_306, i_13_307, i_13_315, i_13_316, i_13_324, i_13_372, i_13_517, i_13_531, i_13_554, i_13_570, i_13_571, i_13_573, i_13_639, i_13_640, i_13_642, i_13_643, i_13_684, i_13_685, i_13_688, i_13_697, i_13_714, i_13_741, i_13_819, i_13_825, i_13_978, i_13_1089, i_13_1120, i_13_1206, i_13_1246, i_13_1269, i_13_1270, i_13_1380, i_13_1387, i_13_1426, i_13_1438, i_13_1503, i_13_1593, i_13_1594, i_13_1638, i_13_1639, i_13_1677, i_13_1693, i_13_1710, i_13_1720, i_13_1752, i_13_1804, i_13_1857, i_13_1858, i_13_1873, i_13_1914, i_13_1915, i_13_1959, i_13_2022, i_13_2023, i_13_2133, i_13_2134, i_13_2259, i_13_2260, i_13_2268, i_13_2272, i_13_2452, i_13_2472, i_13_2550, i_13_2646, i_13_2650, i_13_2673, i_13_2674, i_13_2845, i_13_2916, i_13_3024, i_13_3198, i_13_3205, i_13_3208, i_13_3267, i_13_3270, i_13_3384, i_13_3423, i_13_3735, i_13_3760, i_13_3817, i_13_3924, i_13_4032, i_13_4077, i_13_4078, i_13_4252, i_13_4344, i_13_4357, i_13_4369, i_13_4411, i_13_4566, i_13_4587, i_13_4590, i_13_4591, i_13_4592, o_13_265);
	kernel_13_266 k_13_266(i_13_40, i_13_48, i_13_49, i_13_51, i_13_101, i_13_112, i_13_139, i_13_165, i_13_166, i_13_216, i_13_229, i_13_265, i_13_282, i_13_328, i_13_365, i_13_452, i_13_488, i_13_500, i_13_570, i_13_676, i_13_737, i_13_813, i_13_814, i_13_815, i_13_823, i_13_840, i_13_869, i_13_960, i_13_1063, i_13_1166, i_13_1226, i_13_1242, i_13_1524, i_13_1525, i_13_1570, i_13_1624, i_13_1741, i_13_1753, i_13_1776, i_13_1811, i_13_1831, i_13_1848, i_13_1849, i_13_1882, i_13_1885, i_13_1943, i_13_1997, i_13_2029, i_13_2056, i_13_2136, i_13_2184, i_13_2201, i_13_2380, i_13_2403, i_13_2404, i_13_2407, i_13_2408, i_13_2465, i_13_2551, i_13_2693, i_13_2695, i_13_2756, i_13_2760, i_13_2848, i_13_2938, i_13_3003, i_13_3010, i_13_3092, i_13_3108, i_13_3109, i_13_3274, i_13_3352, i_13_3370, i_13_3440, i_13_3502, i_13_3505, i_13_3506, i_13_3640, i_13_3738, i_13_3739, i_13_3817, i_13_3838, i_13_3889, i_13_3892, i_13_3980, i_13_4017, i_13_4018, i_13_4063, i_13_4064, i_13_4085, i_13_4297, i_13_4315, i_13_4316, i_13_4318, i_13_4319, i_13_4378, i_13_4418, i_13_4425, i_13_4432, i_13_4544, o_13_266);
	kernel_13_267 k_13_267(i_13_28, i_13_31, i_13_63, i_13_64, i_13_90, i_13_91, i_13_94, i_13_95, i_13_225, i_13_226, i_13_287, i_13_306, i_13_307, i_13_355, i_13_367, i_13_369, i_13_380, i_13_468, i_13_538, i_13_606, i_13_607, i_13_616, i_13_649, i_13_667, i_13_729, i_13_756, i_13_757, i_13_814, i_13_829, i_13_945, i_13_946, i_13_953, i_13_1075, i_13_1076, i_13_1099, i_13_1215, i_13_1218, i_13_1219, i_13_1228, i_13_1306, i_13_1318, i_13_1444, i_13_1462, i_13_1594, i_13_1678, i_13_1719, i_13_1720, i_13_1777, i_13_1790, i_13_1840, i_13_1843, i_13_1844, i_13_1858, i_13_1926, i_13_1999, i_13_2001, i_13_2172, i_13_2176, i_13_2407, i_13_2421, i_13_2478, i_13_2534, i_13_2676, i_13_2718, i_13_2719, i_13_2749, i_13_2785, i_13_2821, i_13_2881, i_13_3028, i_13_3060, i_13_3063, i_13_3109, i_13_3116, i_13_3119, i_13_3149, i_13_3241, i_13_3316, i_13_3416, i_13_3460, i_13_3464, i_13_3636, i_13_3712, i_13_3738, i_13_3760, i_13_3797, i_13_3875, i_13_3910, i_13_3925, i_13_3929, i_13_3932, i_13_3979, i_13_4060, i_13_4093, i_13_4120, i_13_4212, i_13_4213, i_13_4351, i_13_4354, i_13_4544, o_13_267);
	kernel_13_268 k_13_268(i_13_103, i_13_133, i_13_134, i_13_139, i_13_237, i_13_252, i_13_280, i_13_319, i_13_326, i_13_429, i_13_469, i_13_524, i_13_588, i_13_608, i_13_668, i_13_821, i_13_852, i_13_951, i_13_1021, i_13_1066, i_13_1076, i_13_1122, i_13_1230, i_13_1275, i_13_1311, i_13_1343, i_13_1401, i_13_1426, i_13_1428, i_13_1468, i_13_1499, i_13_1509, i_13_1599, i_13_1634, i_13_1644, i_13_1651, i_13_1680, i_13_1691, i_13_1696, i_13_1712, i_13_1777, i_13_1778, i_13_1794, i_13_1797, i_13_1811, i_13_1882, i_13_1883, i_13_1914, i_13_1929, i_13_1990, i_13_1991, i_13_1999, i_13_2000, i_13_2002, i_13_2003, i_13_2115, i_13_2134, i_13_2198, i_13_2237, i_13_2265, i_13_2377, i_13_2461, i_13_2470, i_13_2647, i_13_2711, i_13_2763, i_13_2845, i_13_2854, i_13_2935, i_13_2983, i_13_3142, i_13_3143, i_13_3172, i_13_3273, i_13_3448, i_13_3461, i_13_3503, i_13_3727, i_13_3728, i_13_3731, i_13_3783, i_13_3816, i_13_3838, i_13_3874, i_13_4015, i_13_4016, i_13_4038, i_13_4083, i_13_4097, i_13_4162, i_13_4259, i_13_4268, i_13_4270, i_13_4314, i_13_4393, i_13_4411, i_13_4554, i_13_4558, i_13_4567, i_13_4568, o_13_268);
	kernel_13_269 k_13_269(i_13_30, i_13_75, i_13_111, i_13_114, i_13_115, i_13_123, i_13_124, i_13_247, i_13_265, i_13_276, i_13_363, i_13_366, i_13_418, i_13_444, i_13_561, i_13_564, i_13_606, i_13_607, i_13_609, i_13_654, i_13_663, i_13_670, i_13_672, i_13_688, i_13_814, i_13_817, i_13_939, i_13_949, i_13_1083, i_13_1084, i_13_1086, i_13_1114, i_13_1408, i_13_1434, i_13_1446, i_13_1470, i_13_1626, i_13_1653, i_13_1750, i_13_1776, i_13_1804, i_13_1839, i_13_1840, i_13_1842, i_13_1843, i_13_2056, i_13_2130, i_13_2136, i_13_2157, i_13_2172, i_13_2173, i_13_2175, i_13_2247, i_13_2299, i_13_2347, i_13_2407, i_13_2425, i_13_2434, i_13_2436, i_13_2437, i_13_2452, i_13_2497, i_13_2581, i_13_2704, i_13_2748, i_13_2938, i_13_3031, i_13_3049, i_13_3099, i_13_3100, i_13_3103, i_13_3147, i_13_3148, i_13_3156, i_13_3165, i_13_3261, i_13_3504, i_13_3505, i_13_3541, i_13_3615, i_13_3688, i_13_3741, i_13_3760, i_13_3769, i_13_3784, i_13_3877, i_13_3891, i_13_3909, i_13_3910, i_13_4044, i_13_4084, i_13_4119, i_13_4120, i_13_4162, i_13_4327, i_13_4353, i_13_4354, i_13_4449, i_13_4528, i_13_4543, o_13_269);
	kernel_13_270 k_13_270(i_13_25, i_13_61, i_13_76, i_13_119, i_13_163, i_13_164, i_13_177, i_13_182, i_13_184, i_13_185, i_13_186, i_13_187, i_13_192, i_13_193, i_13_194, i_13_196, i_13_347, i_13_382, i_13_419, i_13_518, i_13_571, i_13_573, i_13_574, i_13_625, i_13_628, i_13_661, i_13_697, i_13_715, i_13_717, i_13_811, i_13_837, i_13_841, i_13_850, i_13_853, i_13_1151, i_13_1210, i_13_1211, i_13_1285, i_13_1406, i_13_1407, i_13_1408, i_13_1409, i_13_1411, i_13_1416, i_13_1426, i_13_1471, i_13_1516, i_13_1525, i_13_1681, i_13_1770, i_13_1771, i_13_1805, i_13_1831, i_13_1832, i_13_1834, i_13_1908, i_13_1912, i_13_1959, i_13_1960, i_13_2002, i_13_2146, i_13_2178, i_13_2403, i_13_2452, i_13_2504, i_13_2563, i_13_2572, i_13_2612, i_13_2723, i_13_2736, i_13_2857, i_13_2983, i_13_3049, i_13_3064, i_13_3065, i_13_3108, i_13_3145, i_13_3164, i_13_3165, i_13_3166, i_13_3208, i_13_3209, i_13_3212, i_13_3215, i_13_3261, i_13_3446, i_13_3602, i_13_3604, i_13_3616, i_13_3685, i_13_3730, i_13_3733, i_13_3901, i_13_3979, i_13_4073, i_13_4162, i_13_4261, i_13_4396, i_13_4421, i_13_4569, o_13_270);
	kernel_13_271 k_13_271(i_13_46, i_13_48, i_13_117, i_13_118, i_13_127, i_13_164, i_13_189, i_13_323, i_13_409, i_13_504, i_13_532, i_13_572, i_13_604, i_13_616, i_13_711, i_13_712, i_13_832, i_13_909, i_13_918, i_13_935, i_13_1081, i_13_1147, i_13_1226, i_13_1252, i_13_1378, i_13_1404, i_13_1426, i_13_1435, i_13_1440, i_13_1495, i_13_1503, i_13_1513, i_13_1514, i_13_1534, i_13_1548, i_13_1549, i_13_1595, i_13_1664, i_13_1695, i_13_1711, i_13_1728, i_13_1764, i_13_1766, i_13_1768, i_13_1795, i_13_1906, i_13_1916, i_13_2025, i_13_2056, i_13_2097, i_13_2143, i_13_2149, i_13_2172, i_13_2286, i_13_2296, i_13_2360, i_13_2379, i_13_2430, i_13_2529, i_13_2744, i_13_2901, i_13_2978, i_13_3106, i_13_3113, i_13_3123, i_13_3132, i_13_3214, i_13_3261, i_13_3367, i_13_3547, i_13_3565, i_13_3574, i_13_3637, i_13_3645, i_13_3782, i_13_3843, i_13_3844, i_13_3888, i_13_3897, i_13_3898, i_13_3908, i_13_3910, i_13_3913, i_13_3916, i_13_3979, i_13_3982, i_13_4019, i_13_4042, i_13_4097, i_13_4159, i_13_4230, i_13_4266, i_13_4293, i_13_4321, i_13_4331, i_13_4401, i_13_4509, i_13_4510, i_13_4536, i_13_4606, o_13_271);
	kernel_13_272 k_13_272(i_13_29, i_13_47, i_13_71, i_13_155, i_13_209, i_13_231, i_13_269, i_13_300, i_13_314, i_13_352, i_13_416, i_13_445, i_13_583, i_13_610, i_13_628, i_13_646, i_13_647, i_13_689, i_13_713, i_13_764, i_13_854, i_13_953, i_13_985, i_13_986, i_13_1086, i_13_1106, i_13_1132, i_13_1136, i_13_1226, i_13_1303, i_13_1408, i_13_1495, i_13_1511, i_13_1525, i_13_1551, i_13_1606, i_13_1644, i_13_1717, i_13_1753, i_13_1754, i_13_1799, i_13_1802, i_13_1808, i_13_1918, i_13_1945, i_13_1996, i_13_2122, i_13_2123, i_13_2193, i_13_2195, i_13_2240, i_13_2294, i_13_2373, i_13_2390, i_13_2473, i_13_2515, i_13_2518, i_13_2545, i_13_2567, i_13_2680, i_13_2695, i_13_2698, i_13_2699, i_13_2715, i_13_2786, i_13_2816, i_13_2911, i_13_2941, i_13_3014, i_13_3021, i_13_3031, i_13_3032, i_13_3128, i_13_3133, i_13_3134, i_13_3212, i_13_3232, i_13_3262, i_13_3264, i_13_3347, i_13_3355, i_13_3399, i_13_3453, i_13_3589, i_13_3700, i_13_3760, i_13_3782, i_13_3853, i_13_3916, i_13_4038, i_13_4046, i_13_4085, i_13_4254, i_13_4273, i_13_4326, i_13_4396, i_13_4398, i_13_4557, i_13_4597, i_13_4607, o_13_272);
	kernel_13_273 k_13_273(i_13_106, i_13_107, i_13_124, i_13_142, i_13_170, i_13_184, i_13_269, i_13_320, i_13_340, i_13_341, i_13_380, i_13_449, i_13_458, i_13_511, i_13_618, i_13_746, i_13_781, i_13_817, i_13_818, i_13_836, i_13_934, i_13_980, i_13_1055, i_13_1220, i_13_1222, i_13_1303, i_13_1304, i_13_1309, i_13_1349, i_13_1465, i_13_1573, i_13_1574, i_13_1723, i_13_1789, i_13_1808, i_13_1817, i_13_1825, i_13_1996, i_13_1997, i_13_2053, i_13_2060, i_13_2122, i_13_2123, i_13_2140, i_13_2141, i_13_2411, i_13_2438, i_13_2461, i_13_2506, i_13_2573, i_13_2582, i_13_2728, i_13_2729, i_13_2752, i_13_2861, i_13_2940, i_13_2941, i_13_2942, i_13_3001, i_13_3022, i_13_3023, i_13_3030, i_13_3220, i_13_3221, i_13_3238, i_13_3272, i_13_3292, i_13_3293, i_13_3346, i_13_3347, i_13_3386, i_13_3391, i_13_3392, i_13_3400, i_13_3401, i_13_3418, i_13_3419, i_13_3437, i_13_3505, i_13_3526, i_13_3527, i_13_3560, i_13_3670, i_13_3824, i_13_3881, i_13_3911, i_13_3926, i_13_4049, i_13_4058, i_13_4067, i_13_4166, i_13_4273, i_13_4318, i_13_4319, i_13_4332, i_13_4372, i_13_4396, i_13_4400, i_13_4416, i_13_4594, o_13_273);
	kernel_13_274 k_13_274(i_13_177, i_13_274, i_13_281, i_13_310, i_13_312, i_13_313, i_13_314, i_13_315, i_13_318, i_13_320, i_13_554, i_13_587, i_13_642, i_13_643, i_13_645, i_13_647, i_13_688, i_13_689, i_13_691, i_13_692, i_13_820, i_13_840, i_13_854, i_13_871, i_13_1106, i_13_1119, i_13_1123, i_13_1124, i_13_1211, i_13_1223, i_13_1276, i_13_1277, i_13_1283, i_13_1308, i_13_1311, i_13_1343, i_13_1391, i_13_1394, i_13_1399, i_13_1442, i_13_1511, i_13_1593, i_13_1597, i_13_1600, i_13_1633, i_13_1642, i_13_1649, i_13_1791, i_13_1798, i_13_1799, i_13_1853, i_13_1997, i_13_2000, i_13_2001, i_13_2003, i_13_2004, i_13_2055, i_13_2057, i_13_2194, i_13_2262, i_13_2270, i_13_2272, i_13_2303, i_13_2434, i_13_2555, i_13_2588, i_13_2651, i_13_2680, i_13_2681, i_13_2711, i_13_3011, i_13_3037, i_13_3246, i_13_3272, i_13_3368, i_13_3415, i_13_3419, i_13_3653, i_13_3666, i_13_3736, i_13_3743, i_13_3782, i_13_3868, i_13_3931, i_13_3990, i_13_3995, i_13_4043, i_13_4081, i_13_4085, i_13_4090, i_13_4190, i_13_4193, i_13_4207, i_13_4232, i_13_4297, i_13_4531, i_13_4594, i_13_4595, i_13_4598, i_13_4604, o_13_274);
	kernel_13_275 k_13_275(i_13_63, i_13_64, i_13_75, i_13_103, i_13_174, i_13_184, i_13_211, i_13_379, i_13_453, i_13_523, i_13_558, i_13_567, i_13_585, i_13_696, i_13_707, i_13_738, i_13_741, i_13_759, i_13_840, i_13_855, i_13_1092, i_13_1093, i_13_1137, i_13_1180, i_13_1192, i_13_1200, i_13_1206, i_13_1207, i_13_1209, i_13_1341, i_13_1342, i_13_1425, i_13_1441, i_13_1467, i_13_1468, i_13_1569, i_13_1604, i_13_1649, i_13_1755, i_13_1810, i_13_1855, i_13_1857, i_13_1858, i_13_1920, i_13_1927, i_13_1944, i_13_1946, i_13_2001, i_13_2052, i_13_2053, i_13_2055, i_13_2187, i_13_2262, i_13_2277, i_13_2278, i_13_2341, i_13_2350, i_13_2376, i_13_2563, i_13_2596, i_13_2676, i_13_2709, i_13_2719, i_13_2722, i_13_2766, i_13_2767, i_13_2856, i_13_2857, i_13_2934, i_13_3060, i_13_3061, i_13_3063, i_13_3098, i_13_3126, i_13_3366, i_13_3369, i_13_3414, i_13_3415, i_13_3438, i_13_3439, i_13_3592, i_13_3627, i_13_3681, i_13_3684, i_13_3726, i_13_3910, i_13_4015, i_13_4033, i_13_4152, i_13_4203, i_13_4230, i_13_4302, i_13_4305, i_13_4306, i_13_4348, i_13_4393, i_13_4395, i_13_4410, i_13_4441, i_13_4554, o_13_275);
	kernel_13_276 k_13_276(i_13_37, i_13_61, i_13_117, i_13_189, i_13_190, i_13_222, i_13_223, i_13_226, i_13_273, i_13_333, i_13_387, i_13_396, i_13_408, i_13_561, i_13_567, i_13_585, i_13_603, i_13_604, i_13_607, i_13_608, i_13_629, i_13_657, i_13_669, i_13_742, i_13_855, i_13_945, i_13_1083, i_13_1112, i_13_1368, i_13_1404, i_13_1440, i_13_1486, i_13_1516, i_13_1620, i_13_1623, i_13_1729, i_13_1745, i_13_1785, i_13_1813, i_13_1836, i_13_1837, i_13_1840, i_13_1844, i_13_1924, i_13_2019, i_13_2020, i_13_2023, i_13_2137, i_13_2214, i_13_2359, i_13_2422, i_13_2431, i_13_2497, i_13_2529, i_13_2622, i_13_2650, i_13_2907, i_13_3043, i_13_3099, i_13_3101, i_13_3114, i_13_3126, i_13_3160, i_13_3163, i_13_3261, i_13_3274, i_13_3307, i_13_3322, i_13_3465, i_13_3475, i_13_3523, i_13_3565, i_13_3567, i_13_3598, i_13_3600, i_13_3648, i_13_3730, i_13_3738, i_13_3762, i_13_3763, i_13_3784, i_13_3819, i_13_3843, i_13_3897, i_13_3978, i_13_4005, i_13_4116, i_13_4117, i_13_4158, i_13_4159, i_13_4161, i_13_4162, i_13_4260, i_13_4315, i_13_4324, i_13_4355, i_13_4366, i_13_4467, i_13_4507, i_13_4537, o_13_276);
	kernel_13_277 k_13_277(i_13_130, i_13_170, i_13_286, i_13_352, i_13_383, i_13_422, i_13_461, i_13_466, i_13_467, i_13_512, i_13_526, i_13_527, i_13_529, i_13_530, i_13_535, i_13_547, i_13_625, i_13_800, i_13_817, i_13_881, i_13_1025, i_13_1148, i_13_1273, i_13_1313, i_13_1516, i_13_1553, i_13_1556, i_13_1600, i_13_1634, i_13_1636, i_13_1678, i_13_1849, i_13_1940, i_13_2005, i_13_2006, i_13_2033, i_13_2105, i_13_2131, i_13_2137, i_13_2200, i_13_2203, i_13_2204, i_13_2267, i_13_2278, i_13_2363, i_13_2408, i_13_2462, i_13_2465, i_13_2474, i_13_2510, i_13_2545, i_13_2546, i_13_2557, i_13_2618, i_13_2690, i_13_2711, i_13_2747, i_13_2806, i_13_2852, i_13_2939, i_13_3100, i_13_3118, i_13_3125, i_13_3235, i_13_3265, i_13_3346, i_13_3368, i_13_3461, i_13_3541, i_13_3598, i_13_3644, i_13_3667, i_13_3670, i_13_3730, i_13_3731, i_13_3733, i_13_3734, i_13_3742, i_13_3787, i_13_3860, i_13_3910, i_13_3913, i_13_3914, i_13_3920, i_13_4018, i_13_4019, i_13_4063, i_13_4064, i_13_4210, i_13_4255, i_13_4256, i_13_4265, i_13_4298, i_13_4316, i_13_4342, i_13_4393, i_13_4423, i_13_4543, i_13_4561, i_13_4603, o_13_277);
	kernel_13_278 k_13_278(i_13_0, i_13_14, i_13_22, i_13_64, i_13_76, i_13_168, i_13_182, i_13_199, i_13_225, i_13_228, i_13_247, i_13_280, i_13_336, i_13_339, i_13_378, i_13_381, i_13_531, i_13_536, i_13_573, i_13_585, i_13_586, i_13_639, i_13_640, i_13_717, i_13_781, i_13_927, i_13_1004, i_13_1064, i_13_1081, i_13_1116, i_13_1117, i_13_1141, i_13_1142, i_13_1181, i_13_1296, i_13_1467, i_13_1468, i_13_1470, i_13_1497, i_13_1503, i_13_1647, i_13_1648, i_13_1710, i_13_1711, i_13_1719, i_13_1731, i_13_1782, i_13_1786, i_13_1791, i_13_1792, i_13_1800, i_13_1802, i_13_1851, i_13_1989, i_13_1990, i_13_1993, i_13_2115, i_13_2116, i_13_2259, i_13_2265, i_13_2290, i_13_2358, i_13_2377, i_13_2379, i_13_2536, i_13_2667, i_13_2672, i_13_2673, i_13_2709, i_13_2844, i_13_2845, i_13_2934, i_13_3036, i_13_3040, i_13_3061, i_13_3123, i_13_3153, i_13_3215, i_13_3285, i_13_3286, i_13_3468, i_13_3475, i_13_3550, i_13_3554, i_13_3581, i_13_3610, i_13_3639, i_13_3818, i_13_3924, i_13_4008, i_13_4011, i_13_4042, i_13_4230, i_13_4232, i_13_4302, i_13_4303, i_13_4390, i_13_4391, i_13_4410, i_13_4411, o_13_278);
	kernel_13_279 k_13_279(i_13_46, i_13_53, i_13_80, i_13_91, i_13_114, i_13_140, i_13_161, i_13_171, i_13_178, i_13_216, i_13_228, i_13_237, i_13_251, i_13_273, i_13_278, i_13_441, i_13_455, i_13_518, i_13_544, i_13_562, i_13_576, i_13_619, i_13_700, i_13_723, i_13_885, i_13_888, i_13_936, i_13_944, i_13_945, i_13_1071, i_13_1131, i_13_1262, i_13_1265, i_13_1329, i_13_1483, i_13_1515, i_13_1517, i_13_1569, i_13_1626, i_13_1642, i_13_1643, i_13_1742, i_13_1757, i_13_1777, i_13_1921, i_13_1948, i_13_1953, i_13_2020, i_13_2024, i_13_2087, i_13_2185, i_13_2294, i_13_2302, i_13_2321, i_13_2370, i_13_2424, i_13_2442, i_13_2446, i_13_2447, i_13_2455, i_13_2466, i_13_2716, i_13_2742, i_13_2743, i_13_2744, i_13_2955, i_13_2959, i_13_3042, i_13_3043, i_13_3208, i_13_3316, i_13_3374, i_13_3490, i_13_3541, i_13_3546, i_13_3599, i_13_3604, i_13_3683, i_13_3767, i_13_3769, i_13_3870, i_13_3904, i_13_4110, i_13_4158, i_13_4159, i_13_4161, i_13_4166, i_13_4249, i_13_4321, i_13_4364, i_13_4365, i_13_4432, i_13_4451, i_13_4454, i_13_4495, i_13_4516, i_13_4518, i_13_4536, i_13_4542, i_13_4575, o_13_279);
	kernel_13_280 k_13_280(i_13_32, i_13_52, i_13_70, i_13_71, i_13_79, i_13_80, i_13_140, i_13_176, i_13_230, i_13_314, i_13_322, i_13_323, i_13_377, i_13_526, i_13_527, i_13_557, i_13_589, i_13_608, i_13_610, i_13_647, i_13_674, i_13_683, i_13_734, i_13_853, i_13_986, i_13_1105, i_13_1202, i_13_1222, i_13_1228, i_13_1229, i_13_1231, i_13_1277, i_13_1283, i_13_1312, i_13_1313, i_13_1336, i_13_1394, i_13_1426, i_13_1430, i_13_1510, i_13_1511, i_13_1664, i_13_1724, i_13_1736, i_13_1750, i_13_1751, i_13_1781, i_13_1799, i_13_1843, i_13_1844, i_13_1858, i_13_1886, i_13_1912, i_13_1931, i_13_1934, i_13_1948, i_13_2119, i_13_2194, i_13_2195, i_13_2287, i_13_2426, i_13_2462, i_13_2509, i_13_2552, i_13_2600, i_13_2722, i_13_2851, i_13_2852, i_13_3095, i_13_3104, i_13_3118, i_13_3146, i_13_3271, i_13_3272, i_13_3398, i_13_3418, i_13_3419, i_13_3433, i_13_3439, i_13_3479, i_13_3548, i_13_3614, i_13_3743, i_13_3761, i_13_3769, i_13_3869, i_13_3896, i_13_3932, i_13_3994, i_13_4040, i_13_4063, i_13_4085, i_13_4190, i_13_4252, i_13_4297, i_13_4298, i_13_4382, i_13_4534, i_13_4597, i_13_4598, o_13_280);
	kernel_13_281 k_13_281(i_13_31, i_13_58, i_13_94, i_13_184, i_13_192, i_13_310, i_13_324, i_13_463, i_13_570, i_13_575, i_13_628, i_13_660, i_13_661, i_13_714, i_13_760, i_13_796, i_13_840, i_13_858, i_13_859, i_13_861, i_13_927, i_13_1224, i_13_1225, i_13_1227, i_13_1228, i_13_1230, i_13_1231, i_13_1254, i_13_1255, i_13_1345, i_13_1407, i_13_1408, i_13_1452, i_13_1470, i_13_1488, i_13_1489, i_13_1507, i_13_1596, i_13_1597, i_13_1632, i_13_1686, i_13_1687, i_13_1714, i_13_1740, i_13_1758, i_13_1769, i_13_1854, i_13_1857, i_13_1858, i_13_1917, i_13_1918, i_13_1930, i_13_1957, i_13_2011, i_13_2055, i_13_2056, i_13_2226, i_13_2312, i_13_2425, i_13_2458, i_13_2568, i_13_2618, i_13_2629, i_13_2676, i_13_2695, i_13_2856, i_13_2857, i_13_2946, i_13_3031, i_13_3063, i_13_3064, i_13_3100, i_13_3114, i_13_3171, i_13_3172, i_13_3204, i_13_3414, i_13_3421, i_13_3459, i_13_3460, i_13_3487, i_13_3531, i_13_3532, i_13_3718, i_13_3802, i_13_3854, i_13_3855, i_13_3856, i_13_3873, i_13_3874, i_13_3982, i_13_4050, i_13_4216, i_13_4306, i_13_4341, i_13_4363, i_13_4396, i_13_4423, i_13_4446, i_13_4507, o_13_281);
	kernel_13_282 k_13_282(i_13_92, i_13_96, i_13_97, i_13_105, i_13_112, i_13_175, i_13_237, i_13_310, i_13_319, i_13_519, i_13_578, i_13_604, i_13_618, i_13_643, i_13_652, i_13_653, i_13_740, i_13_771, i_13_816, i_13_884, i_13_913, i_13_921, i_13_929, i_13_940, i_13_979, i_13_1077, i_13_1084, i_13_1109, i_13_1280, i_13_1329, i_13_1337, i_13_1441, i_13_1464, i_13_1480, i_13_1535, i_13_1597, i_13_1607, i_13_1609, i_13_1667, i_13_1776, i_13_1786, i_13_1816, i_13_1841, i_13_1894, i_13_1924, i_13_1948, i_13_2020, i_13_2029, i_13_2144, i_13_2156, i_13_2173, i_13_2317, i_13_2425, i_13_2444, i_13_2468, i_13_2498, i_13_2667, i_13_2749, i_13_2750, i_13_2813, i_13_2838, i_13_2884, i_13_2940, i_13_3110, i_13_3155, i_13_3218, i_13_3230, i_13_3268, i_13_3315, i_13_3350, i_13_3380, i_13_3460, i_13_3491, i_13_3504, i_13_3522, i_13_3620, i_13_3649, i_13_3746, i_13_3757, i_13_3824, i_13_3874, i_13_3910, i_13_3913, i_13_4036, i_13_4089, i_13_4091, i_13_4124, i_13_4126, i_13_4187, i_13_4360, i_13_4361, i_13_4366, i_13_4372, i_13_4396, i_13_4412, i_13_4416, i_13_4465, i_13_4492, i_13_4519, i_13_4523, o_13_282);
	kernel_13_283 k_13_283(i_13_27, i_13_28, i_13_102, i_13_103, i_13_126, i_13_153, i_13_154, i_13_190, i_13_282, i_13_585, i_13_586, i_13_669, i_13_846, i_13_856, i_13_914, i_13_949, i_13_1080, i_13_1081, i_13_1206, i_13_1305, i_13_1341, i_13_1342, i_13_1422, i_13_1434, i_13_1441, i_13_1443, i_13_1467, i_13_1504, i_13_1540, i_13_1632, i_13_1678, i_13_1750, i_13_1782, i_13_1803, i_13_1810, i_13_1839, i_13_1840, i_13_1926, i_13_1927, i_13_1999, i_13_2001, i_13_2052, i_13_2053, i_13_2054, i_13_2109, i_13_2119, i_13_2197, i_13_2259, i_13_2277, i_13_2278, i_13_2341, i_13_2407, i_13_2433, i_13_2443, i_13_2512, i_13_2541, i_13_2542, i_13_2550, i_13_2614, i_13_2619, i_13_2629, i_13_2686, i_13_2709, i_13_2710, i_13_2853, i_13_2854, i_13_2858, i_13_2917, i_13_2946, i_13_3061, i_13_3150, i_13_3205, i_13_3307, i_13_3315, i_13_3415, i_13_3432, i_13_3528, i_13_3532, i_13_3610, i_13_3627, i_13_3730, i_13_3862, i_13_3979, i_13_4014, i_13_4050, i_13_4059, i_13_4087, i_13_4114, i_13_4230, i_13_4231, i_13_4248, i_13_4257, i_13_4268, i_13_4270, i_13_4338, i_13_4342, i_13_4392, i_13_4393, i_13_4394, i_13_4536, o_13_283);
	kernel_13_284 k_13_284(i_13_39, i_13_40, i_13_66, i_13_125, i_13_178, i_13_268, i_13_308, i_13_310, i_13_318, i_13_319, i_13_463, i_13_466, i_13_489, i_13_536, i_13_589, i_13_591, i_13_592, i_13_625, i_13_640, i_13_645, i_13_646, i_13_690, i_13_691, i_13_763, i_13_817, i_13_841, i_13_933, i_13_1122, i_13_1228, i_13_1284, i_13_1347, i_13_1348, i_13_1411, i_13_1437, i_13_1542, i_13_1596, i_13_1597, i_13_1599, i_13_1671, i_13_1754, i_13_1852, i_13_1941, i_13_1959, i_13_2001, i_13_2002, i_13_2058, i_13_2059, i_13_2139, i_13_2181, i_13_2182, i_13_2193, i_13_2265, i_13_2275, i_13_2283, i_13_2284, i_13_2410, i_13_2554, i_13_2614, i_13_2617, i_13_2652, i_13_2653, i_13_2673, i_13_2679, i_13_2697, i_13_2698, i_13_2760, i_13_2823, i_13_2856, i_13_2859, i_13_2860, i_13_2997, i_13_3004, i_13_3212, i_13_3275, i_13_3372, i_13_3390, i_13_3391, i_13_3392, i_13_3415, i_13_3487, i_13_3532, i_13_3535, i_13_3616, i_13_3721, i_13_3877, i_13_3930, i_13_4034, i_13_4035, i_13_4207, i_13_4218, i_13_4308, i_13_4309, i_13_4341, i_13_4363, i_13_4372, i_13_4399, i_13_4540, i_13_4543, i_13_4585, i_13_4597, o_13_284);
	kernel_13_285 k_13_285(i_13_25, i_13_40, i_13_67, i_13_70, i_13_87, i_13_276, i_13_310, i_13_319, i_13_382, i_13_411, i_13_492, i_13_520, i_13_609, i_13_628, i_13_660, i_13_663, i_13_744, i_13_746, i_13_805, i_13_835, i_13_912, i_13_934, i_13_939, i_13_1020, i_13_1021, i_13_1074, i_13_1086, i_13_1087, i_13_1095, i_13_1096, i_13_1111, i_13_1147, i_13_1156, i_13_1330, i_13_1403, i_13_1470, i_13_1474, i_13_1597, i_13_1716, i_13_1735, i_13_1744, i_13_1750, i_13_1767, i_13_1795, i_13_1798, i_13_1857, i_13_1965, i_13_2022, i_13_2023, i_13_2028, i_13_2059, i_13_2060, i_13_2199, i_13_2235, i_13_2454, i_13_2472, i_13_2473, i_13_2500, i_13_2617, i_13_2676, i_13_2715, i_13_2733, i_13_2743, i_13_2769, i_13_2884, i_13_3030, i_13_3031, i_13_3076, i_13_3093, i_13_3121, i_13_3144, i_13_3264, i_13_3265, i_13_3306, i_13_3355, i_13_3435, i_13_3453, i_13_3454, i_13_3486, i_13_3527, i_13_3549, i_13_3576, i_13_3613, i_13_3741, i_13_3742, i_13_3822, i_13_3823, i_13_3927, i_13_3981, i_13_4092, i_13_4093, i_13_4119, i_13_4161, i_13_4164, i_13_4165, i_13_4254, i_13_4417, i_13_4461, i_13_4596, i_13_4606, o_13_285);
	kernel_13_286 k_13_286(i_13_24, i_13_87, i_13_133, i_13_165, i_13_168, i_13_183, i_13_192, i_13_318, i_13_319, i_13_334, i_13_336, i_13_447, i_13_468, i_13_469, i_13_492, i_13_516, i_13_594, i_13_615, i_13_619, i_13_627, i_13_628, i_13_648, i_13_762, i_13_945, i_13_946, i_13_951, i_13_999, i_13_1018, i_13_1095, i_13_1227, i_13_1257, i_13_1314, i_13_1482, i_13_1483, i_13_1495, i_13_1525, i_13_1537, i_13_1542, i_13_1548, i_13_1620, i_13_1626, i_13_1627, i_13_1633, i_13_1723, i_13_1725, i_13_1734, i_13_1770, i_13_1806, i_13_1924, i_13_1941, i_13_1959, i_13_2002, i_13_2052, i_13_2103, i_13_2142, i_13_2238, i_13_2258, i_13_2364, i_13_2382, i_13_2445, i_13_2538, i_13_2727, i_13_2730, i_13_2850, i_13_2940, i_13_2985, i_13_2998, i_13_3021, i_13_3075, i_13_3220, i_13_3240, i_13_3241, i_13_3246, i_13_3264, i_13_3265, i_13_3282, i_13_3310, i_13_3345, i_13_3355, i_13_3528, i_13_3534, i_13_3535, i_13_3639, i_13_3702, i_13_3733, i_13_3759, i_13_3877, i_13_3889, i_13_3891, i_13_3892, i_13_3984, i_13_3985, i_13_4018, i_13_4044, i_13_4137, i_13_4185, i_13_4272, i_13_4294, i_13_4296, i_13_4425, o_13_286);
	kernel_13_287 k_13_287(i_13_40, i_13_53, i_13_95, i_13_96, i_13_143, i_13_274, i_13_287, i_13_341, i_13_476, i_13_521, i_13_529, i_13_565, i_13_592, i_13_644, i_13_646, i_13_647, i_13_688, i_13_689, i_13_691, i_13_692, i_13_797, i_13_980, i_13_1025, i_13_1101, i_13_1121, i_13_1123, i_13_1124, i_13_1204, i_13_1256, i_13_1273, i_13_1277, i_13_1384, i_13_1391, i_13_1444, i_13_1445, i_13_1465, i_13_1484, i_13_1489, i_13_1502, i_13_1627, i_13_1643, i_13_1714, i_13_1715, i_13_1885, i_13_1886, i_13_1888, i_13_1991, i_13_2059, i_13_2140, i_13_2267, i_13_2285, i_13_2354, i_13_2428, i_13_2447, i_13_2464, i_13_2497, i_13_2506, i_13_2509, i_13_2510, i_13_2511, i_13_2533, i_13_2542, i_13_2569, i_13_2648, i_13_2650, i_13_2651, i_13_2653, i_13_2654, i_13_2677, i_13_2752, i_13_2753, i_13_2825, i_13_2848, i_13_2849, i_13_2920, i_13_3004, i_13_3126, i_13_3146, i_13_3217, i_13_3391, i_13_3392, i_13_3424, i_13_3445, i_13_3550, i_13_3794, i_13_3874, i_13_3914, i_13_3982, i_13_3991, i_13_3992, i_13_3995, i_13_4057, i_13_4081, i_13_4085, i_13_4153, i_13_4162, i_13_4318, i_13_4372, i_13_4381, i_13_4444, o_13_287);
	kernel_13_288 k_13_288(i_13_49, i_13_167, i_13_173, i_13_190, i_13_211, i_13_255, i_13_280, i_13_283, i_13_314, i_13_379, i_13_380, i_13_472, i_13_526, i_13_530, i_13_571, i_13_640, i_13_641, i_13_659, i_13_661, i_13_662, i_13_668, i_13_676, i_13_677, i_13_810, i_13_928, i_13_941, i_13_992, i_13_1063, i_13_1081, i_13_1082, i_13_1306, i_13_1307, i_13_1411, i_13_1444, i_13_1498, i_13_1499, i_13_1504, i_13_1505, i_13_1633, i_13_1636, i_13_1730, i_13_1783, i_13_1801, i_13_1838, i_13_1846, i_13_1880, i_13_1927, i_13_1942, i_13_2054, i_13_2170, i_13_2315, i_13_2425, i_13_2431, i_13_2432, i_13_2674, i_13_2923, i_13_3107, i_13_3142, i_13_3143, i_13_3242, i_13_3267, i_13_3269, i_13_3271, i_13_3371, i_13_3420, i_13_3421, i_13_3422, i_13_3424, i_13_3425, i_13_3545, i_13_3646, i_13_3730, i_13_3731, i_13_3767, i_13_3817, i_13_3818, i_13_3925, i_13_3971, i_13_3989, i_13_4015, i_13_4016, i_13_4018, i_13_4019, i_13_4044, i_13_4060, i_13_4061, i_13_4078, i_13_4214, i_13_4249, i_13_4250, i_13_4253, i_13_4261, i_13_4313, i_13_4340, i_13_4351, i_13_4430, i_13_4556, i_13_4558, i_13_4567, i_13_4591, o_13_288);
	kernel_13_289 k_13_289(i_13_120, i_13_139, i_13_140, i_13_142, i_13_175, i_13_177, i_13_227, i_13_228, i_13_281, i_13_310, i_13_338, i_13_371, i_13_418, i_13_532, i_13_538, i_13_617, i_13_654, i_13_700, i_13_769, i_13_817, i_13_821, i_13_892, i_13_897, i_13_918, i_13_982, i_13_985, i_13_1114, i_13_1219, i_13_1220, i_13_1228, i_13_1327, i_13_1424, i_13_1473, i_13_1525, i_13_1599, i_13_1627, i_13_1711, i_13_1714, i_13_1720, i_13_1723, i_13_1724, i_13_1831, i_13_1841, i_13_1844, i_13_1849, i_13_1882, i_13_1883, i_13_1885, i_13_1888, i_13_2104, i_13_2110, i_13_2206, i_13_2407, i_13_2410, i_13_2424, i_13_2463, i_13_2499, i_13_2663, i_13_2678, i_13_2695, i_13_2845, i_13_2846, i_13_2857, i_13_2875, i_13_2983, i_13_3005, i_13_3010, i_13_3109, i_13_3142, i_13_3143, i_13_3165, i_13_3444, i_13_3450, i_13_3451, i_13_3482, i_13_3503, i_13_3505, i_13_3506, i_13_3524, i_13_3571, i_13_3685, i_13_3686, i_13_3688, i_13_3736, i_13_3737, i_13_3740, i_13_3820, i_13_3836, i_13_3900, i_13_3928, i_13_4015, i_13_4066, i_13_4082, i_13_4204, i_13_4315, i_13_4388, i_13_4412, i_13_4459, i_13_4520, i_13_4567, o_13_289);
	kernel_13_290 k_13_290(i_13_127, i_13_130, i_13_131, i_13_272, i_13_280, i_13_329, i_13_354, i_13_355, i_13_364, i_13_442, i_13_469, i_13_490, i_13_667, i_13_668, i_13_694, i_13_820, i_13_828, i_13_829, i_13_830, i_13_939, i_13_946, i_13_1022, i_13_1081, i_13_1100, i_13_1256, i_13_1271, i_13_1306, i_13_1307, i_13_1397, i_13_1435, i_13_1499, i_13_1504, i_13_1620, i_13_1639, i_13_1640, i_13_1657, i_13_1696, i_13_1697, i_13_1721, i_13_1777, i_13_1792, i_13_1793, i_13_1846, i_13_2029, i_13_2142, i_13_2143, i_13_2191, i_13_2296, i_13_2297, i_13_2317, i_13_2431, i_13_2432, i_13_2444, i_13_2468, i_13_2511, i_13_2512, i_13_2549, i_13_2552, i_13_2692, i_13_2719, i_13_2720, i_13_2880, i_13_2881, i_13_2882, i_13_2921, i_13_2935, i_13_3097, i_13_3136, i_13_3241, i_13_3242, i_13_3416, i_13_3421, i_13_3523, i_13_3595, i_13_3619, i_13_3620, i_13_3631, i_13_3632, i_13_3731, i_13_3754, i_13_3780, i_13_3802, i_13_3925, i_13_3935, i_13_3989, i_13_3991, i_13_3992, i_13_4198, i_13_4212, i_13_4214, i_13_4311, i_13_4313, i_13_4329, i_13_4330, i_13_4331, i_13_4339, i_13_4429, i_13_4430, i_13_4450, i_13_4510, o_13_290);
	kernel_13_291 k_13_291(i_13_31, i_13_48, i_13_49, i_13_51, i_13_94, i_13_121, i_13_137, i_13_166, i_13_229, i_13_316, i_13_514, i_13_550, i_13_558, i_13_640, i_13_652, i_13_657, i_13_676, i_13_677, i_13_678, i_13_756, i_13_757, i_13_838, i_13_839, i_13_855, i_13_928, i_13_939, i_13_940, i_13_981, i_13_982, i_13_1063, i_13_1072, i_13_1080, i_13_1098, i_13_1323, i_13_1324, i_13_1327, i_13_1486, i_13_1570, i_13_1647, i_13_1747, i_13_1809, i_13_1831, i_13_1908, i_13_1911, i_13_2016, i_13_2017, i_13_2052, i_13_2055, i_13_2107, i_13_2116, i_13_2260, i_13_2380, i_13_2407, i_13_2433, i_13_2448, i_13_2449, i_13_2467, i_13_2505, i_13_2506, i_13_2592, i_13_2674, i_13_2702, i_13_2710, i_13_2749, i_13_2817, i_13_2908, i_13_2939, i_13_2979, i_13_2980, i_13_3025, i_13_3096, i_13_3109, i_13_3110, i_13_3142, i_13_3291, i_13_3519, i_13_3532, i_13_3541, i_13_3549, i_13_3550, i_13_3646, i_13_3737, i_13_3765, i_13_3766, i_13_3817, i_13_3818, i_13_3862, i_13_3889, i_13_3987, i_13_3988, i_13_4063, i_13_4087, i_13_4122, i_13_4158, i_13_4185, i_13_4279, i_13_4320, i_13_4393, i_13_4591, i_13_4600, o_13_291);
	kernel_13_292 k_13_292(i_13_49, i_13_70, i_13_71, i_13_78, i_13_79, i_13_80, i_13_105, i_13_232, i_13_312, i_13_313, i_13_314, i_13_319, i_13_320, i_13_358, i_13_448, i_13_457, i_13_525, i_13_553, i_13_624, i_13_644, i_13_646, i_13_673, i_13_682, i_13_688, i_13_689, i_13_692, i_13_844, i_13_935, i_13_969, i_13_1050, i_13_1104, i_13_1105, i_13_1110, i_13_1123, i_13_1274, i_13_1311, i_13_1312, i_13_1330, i_13_1402, i_13_1403, i_13_1429, i_13_1508, i_13_1510, i_13_1541, i_13_1645, i_13_1646, i_13_1798, i_13_1799, i_13_1843, i_13_1853, i_13_1887, i_13_1912, i_13_1945, i_13_1946, i_13_1948, i_13_2027, i_13_2104, i_13_2203, i_13_2229, i_13_2245, i_13_2291, i_13_2415, i_13_2680, i_13_2697, i_13_2698, i_13_2699, i_13_2852, i_13_2853, i_13_2858, i_13_2923, i_13_3031, i_13_3054, i_13_3067, i_13_3130, i_13_3138, i_13_3245, i_13_3370, i_13_3373, i_13_3418, i_13_3561, i_13_3595, i_13_3622, i_13_3623, i_13_3652, i_13_3787, i_13_3895, i_13_3931, i_13_3940, i_13_3994, i_13_3995, i_13_4068, i_13_4084, i_13_4111, i_13_4156, i_13_4435, i_13_4454, i_13_4595, i_13_4596, i_13_4597, i_13_4598, o_13_292);
	kernel_13_293 k_13_293(i_13_49, i_13_74, i_13_77, i_13_113, i_13_166, i_13_172, i_13_175, i_13_176, i_13_200, i_13_326, i_13_337, i_13_523, i_13_544, i_13_658, i_13_661, i_13_662, i_13_694, i_13_824, i_13_839, i_13_841, i_13_848, i_13_853, i_13_859, i_13_1018, i_13_1019, i_13_1072, i_13_1073, i_13_1148, i_13_1225, i_13_1226, i_13_1229, i_13_1231, i_13_1253, i_13_1310, i_13_1315, i_13_1316, i_13_1324, i_13_1378, i_13_1424, i_13_1427, i_13_1441, i_13_1486, i_13_1487, i_13_1549, i_13_1550, i_13_1630, i_13_1778, i_13_1849, i_13_1883, i_13_1885, i_13_1886, i_13_1909, i_13_2021, i_13_2137, i_13_2173, i_13_2371, i_13_2452, i_13_2453, i_13_2462, i_13_2539, i_13_2540, i_13_2561, i_13_2611, i_13_2749, i_13_2917, i_13_2984, i_13_3269, i_13_3367, i_13_3370, i_13_3395, i_13_3484, i_13_3485, i_13_3488, i_13_3502, i_13_3503, i_13_3530, i_13_3538, i_13_3539, i_13_3541, i_13_3542, i_13_3548, i_13_3574, i_13_3575, i_13_3703, i_13_3740, i_13_3812, i_13_3854, i_13_3866, i_13_3892, i_13_3916, i_13_4063, i_13_4064, i_13_4249, i_13_4250, i_13_4252, i_13_4253, i_13_4366, i_13_4369, i_13_4376, i_13_4448, o_13_293);
	kernel_13_294 k_13_294(i_13_28, i_13_29, i_13_52, i_13_65, i_13_103, i_13_124, i_13_140, i_13_175, i_13_211, i_13_257, i_13_266, i_13_308, i_13_316, i_13_340, i_13_358, i_13_359, i_13_371, i_13_418, i_13_419, i_13_584, i_13_587, i_13_604, i_13_640, i_13_641, i_13_668, i_13_679, i_13_757, i_13_758, i_13_856, i_13_928, i_13_1081, i_13_1082, i_13_1117, i_13_1300, i_13_1342, i_13_1343, i_13_1345, i_13_1501, i_13_1502, i_13_1567, i_13_1637, i_13_1793, i_13_1804, i_13_1813, i_13_1840, i_13_1841, i_13_1928, i_13_1991, i_13_2002, i_13_2032, i_13_2033, i_13_2054, i_13_2119, i_13_2137, i_13_2260, i_13_2432, i_13_2549, i_13_2554, i_13_2674, i_13_2675, i_13_2710, i_13_2719, i_13_2846, i_13_2848, i_13_2924, i_13_2938, i_13_2960, i_13_3061, i_13_3073, i_13_3088, i_13_3217, i_13_3289, i_13_3343, i_13_3386, i_13_3415, i_13_3416, i_13_3440, i_13_3485, i_13_3501, i_13_3502, i_13_3503, i_13_3634, i_13_3737, i_13_3788, i_13_3800, i_13_3806, i_13_3851, i_13_3893, i_13_4018, i_13_4034, i_13_4078, i_13_4234, i_13_4267, i_13_4268, i_13_4270, i_13_4274, i_13_4411, i_13_4454, i_13_4591, i_13_4592, o_13_294);
	kernel_13_295 k_13_295(i_13_39, i_13_94, i_13_95, i_13_97, i_13_102, i_13_176, i_13_178, i_13_179, i_13_241, i_13_310, i_13_311, i_13_313, i_13_314, i_13_318, i_13_319, i_13_320, i_13_337, i_13_418, i_13_510, i_13_527, i_13_574, i_13_575, i_13_580, i_13_643, i_13_646, i_13_647, i_13_674, i_13_689, i_13_872, i_13_931, i_13_985, i_13_988, i_13_989, i_13_1123, i_13_1124, i_13_1186, i_13_1444, i_13_1516, i_13_1526, i_13_1598, i_13_1641, i_13_1642, i_13_1813, i_13_1850, i_13_1934, i_13_2137, i_13_2176, i_13_2177, i_13_2264, i_13_2314, i_13_2408, i_13_2567, i_13_2614, i_13_2678, i_13_2680, i_13_2681, i_13_2698, i_13_2699, i_13_2788, i_13_2887, i_13_2923, i_13_2983, i_13_3010, i_13_3113, i_13_3127, i_13_3128, i_13_3212, i_13_3217, i_13_3274, i_13_3370, i_13_3379, i_13_3408, i_13_3409, i_13_3410, i_13_3415, i_13_3426, i_13_3469, i_13_3554, i_13_3688, i_13_3821, i_13_3901, i_13_3931, i_13_3932, i_13_4034, i_13_4036, i_13_4037, i_13_4084, i_13_4208, i_13_4261, i_13_4327, i_13_4342, i_13_4354, i_13_4522, i_13_4523, i_13_4568, i_13_4569, i_13_4570, i_13_4571, i_13_4595, i_13_4598, o_13_295);
	kernel_13_296 k_13_296(i_13_106, i_13_116, i_13_139, i_13_213, i_13_229, i_13_241, i_13_319, i_13_326, i_13_359, i_13_492, i_13_744, i_13_745, i_13_826, i_13_948, i_13_1066, i_13_1071, i_13_1087, i_13_1095, i_13_1096, i_13_1097, i_13_1131, i_13_1239, i_13_1267, i_13_1274, i_13_1302, i_13_1303, i_13_1347, i_13_1348, i_13_1349, i_13_1402, i_13_1435, i_13_1438, i_13_1446, i_13_1464, i_13_1529, i_13_1721, i_13_1722, i_13_1723, i_13_1755, i_13_1803, i_13_1815, i_13_1816, i_13_1817, i_13_1916, i_13_2023, i_13_2111, i_13_2123, i_13_2199, i_13_2238, i_13_2239, i_13_2273, i_13_2347, i_13_2348, i_13_2447, i_13_2500, i_13_2550, i_13_2715, i_13_2716, i_13_2717, i_13_2760, i_13_2789, i_13_2814, i_13_2822, i_13_2825, i_13_2853, i_13_2875, i_13_3023, i_13_3028, i_13_3036, i_13_3112, i_13_3328, i_13_3391, i_13_3422, i_13_3443, i_13_3446, i_13_3479, i_13_3482, i_13_3532, i_13_3594, i_13_3595, i_13_3622, i_13_3742, i_13_3817, i_13_3820, i_13_3830, i_13_3893, i_13_3921, i_13_3984, i_13_3985, i_13_4093, i_13_4120, i_13_4237, i_13_4252, i_13_4261, i_13_4272, i_13_4327, i_13_4328, i_13_4396, i_13_4399, i_13_4417, o_13_296);
	kernel_13_297 k_13_297(i_13_69, i_13_124, i_13_154, i_13_166, i_13_178, i_13_195, i_13_210, i_13_211, i_13_228, i_13_231, i_13_232, i_13_247, i_13_376, i_13_528, i_13_534, i_13_640, i_13_642, i_13_646, i_13_714, i_13_717, i_13_771, i_13_826, i_13_861, i_13_862, i_13_895, i_13_951, i_13_952, i_13_1066, i_13_1075, i_13_1221, i_13_1222, i_13_1275, i_13_1293, i_13_1390, i_13_1410, i_13_1432, i_13_1491, i_13_1492, i_13_1627, i_13_1635, i_13_1641, i_13_1713, i_13_1726, i_13_1795, i_13_1842, i_13_1843, i_13_1884, i_13_1885, i_13_1929, i_13_1989, i_13_1993, i_13_2014, i_13_2028, i_13_2110, i_13_2175, i_13_2262, i_13_2410, i_13_2425, i_13_2463, i_13_2506, i_13_2535, i_13_2536, i_13_2616, i_13_2760, i_13_2847, i_13_2850, i_13_2851, i_13_3097, i_13_3345, i_13_3384, i_13_3387, i_13_3418, i_13_3426, i_13_3504, i_13_3505, i_13_3594, i_13_3669, i_13_3706, i_13_3766, i_13_3838, i_13_3876, i_13_3895, i_13_3931, i_13_4003, i_13_4011, i_13_4048, i_13_4080, i_13_4081, i_13_4086, i_13_4087, i_13_4114, i_13_4189, i_13_4210, i_13_4218, i_13_4273, i_13_4296, i_13_4297, i_13_4315, i_13_4543, i_13_4557, o_13_297);
	kernel_13_298 k_13_298(i_13_31, i_13_39, i_13_63, i_13_64, i_13_98, i_13_128, i_13_137, i_13_175, i_13_184, i_13_214, i_13_229, i_13_269, i_13_279, i_13_280, i_13_306, i_13_323, i_13_337, i_13_352, i_13_379, i_13_525, i_13_605, i_13_616, i_13_683, i_13_768, i_13_824, i_13_1066, i_13_1070, i_13_1142, i_13_1150, i_13_1216, i_13_1218, i_13_1306, i_13_1309, i_13_1326, i_13_1553, i_13_1561, i_13_1570, i_13_1593, i_13_1594, i_13_1604, i_13_1638, i_13_1720, i_13_1748, i_13_1792, i_13_1804, i_13_1831, i_13_1835, i_13_1847, i_13_1882, i_13_1930, i_13_1998, i_13_1999, i_13_2233, i_13_2267, i_13_2407, i_13_2426, i_13_2429, i_13_2505, i_13_2657, i_13_2673, i_13_2677, i_13_2718, i_13_2739, i_13_2740, i_13_2853, i_13_2856, i_13_2872, i_13_2986, i_13_3028, i_13_3073, i_13_3141, i_13_3149, i_13_3211, i_13_3446, i_13_3488, i_13_3501, i_13_3502, i_13_3523, i_13_3538, i_13_3539, i_13_3541, i_13_3609, i_13_3638, i_13_3641, i_13_3727, i_13_3728, i_13_3857, i_13_3860, i_13_3934, i_13_4022, i_13_4063, i_13_4085, i_13_4121, i_13_4126, i_13_4162, i_13_4315, i_13_4318, i_13_4355, i_13_4395, i_13_4570, o_13_298);
	kernel_13_299 k_13_299(i_13_31, i_13_58, i_13_64, i_13_103, i_13_104, i_13_130, i_13_162, i_13_184, i_13_237, i_13_307, i_13_553, i_13_556, i_13_586, i_13_598, i_13_612, i_13_684, i_13_693, i_13_814, i_13_822, i_13_828, i_13_837, i_13_1065, i_13_1066, i_13_1117, i_13_1120, i_13_1206, i_13_1213, i_13_1305, i_13_1306, i_13_1309, i_13_1387, i_13_1390, i_13_1425, i_13_1507, i_13_1624, i_13_1639, i_13_1644, i_13_1648, i_13_1669, i_13_1741, i_13_1846, i_13_1926, i_13_1927, i_13_1957, i_13_2008, i_13_2100, i_13_2142, i_13_2143, i_13_2188, i_13_2199, i_13_2377, i_13_2380, i_13_2407, i_13_2461, i_13_2462, i_13_2676, i_13_2692, i_13_2718, i_13_2754, i_13_2848, i_13_2858, i_13_2881, i_13_2935, i_13_2938, i_13_3009, i_13_3047, i_13_3205, i_13_3208, i_13_3486, i_13_3537, i_13_3637, i_13_3719, i_13_3738, i_13_3753, i_13_3754, i_13_3853, i_13_3907, i_13_3910, i_13_3924, i_13_3927, i_13_3928, i_13_3936, i_13_4032, i_13_4033, i_13_4034, i_13_4035, i_13_4063, i_13_4214, i_13_4216, i_13_4294, i_13_4311, i_13_4315, i_13_4318, i_13_4325, i_13_4330, i_13_4341, i_13_4509, i_13_4522, i_13_4591, i_13_4593, o_13_299);
	kernel_13_300 k_13_300(i_13_91, i_13_93, i_13_94, i_13_95, i_13_121, i_13_125, i_13_165, i_13_184, i_13_238, i_13_309, i_13_367, i_13_564, i_13_571, i_13_572, i_13_697, i_13_730, i_13_733, i_13_793, i_13_797, i_13_859, i_13_1120, i_13_1179, i_13_1180, i_13_1188, i_13_1210, i_13_1218, i_13_1273, i_13_1390, i_13_1408, i_13_1441, i_13_1489, i_13_1624, i_13_1632, i_13_1660, i_13_1683, i_13_1786, i_13_1832, i_13_1843, i_13_1844, i_13_1921, i_13_2088, i_13_2127, i_13_2128, i_13_2169, i_13_2173, i_13_2175, i_13_2176, i_13_2208, i_13_2209, i_13_2237, i_13_2380, i_13_2424, i_13_2425, i_13_2426, i_13_2427, i_13_2428, i_13_2446, i_13_2533, i_13_2541, i_13_2542, i_13_2551, i_13_2567, i_13_2614, i_13_2652, i_13_2722, i_13_2848, i_13_2884, i_13_2985, i_13_3109, i_13_3112, i_13_3147, i_13_3163, i_13_3165, i_13_3211, i_13_3216, i_13_3348, i_13_3373, i_13_3388, i_13_3390, i_13_3424, i_13_3425, i_13_3532, i_13_3732, i_13_3767, i_13_3846, i_13_3870, i_13_3872, i_13_3874, i_13_3875, i_13_4006, i_13_4008, i_13_4121, i_13_4189, i_13_4346, i_13_4351, i_13_4353, i_13_4354, i_13_4355, i_13_4570, i_13_4579, o_13_300);
	kernel_13_301 k_13_301(i_13_124, i_13_143, i_13_187, i_13_188, i_13_229, i_13_283, i_13_287, i_13_340, i_13_374, i_13_446, i_13_508, i_13_535, i_13_536, i_13_543, i_13_548, i_13_571, i_13_574, i_13_580, i_13_594, i_13_599, i_13_616, i_13_644, i_13_718, i_13_728, i_13_777, i_13_781, i_13_845, i_13_895, i_13_914, i_13_941, i_13_1069, i_13_1231, i_13_1249, i_13_1435, i_13_1439, i_13_1444, i_13_1465, i_13_1484, i_13_1499, i_13_1502, i_13_1543, i_13_1634, i_13_1636, i_13_1643, i_13_1694, i_13_1724, i_13_1742, i_13_1750, i_13_1762, i_13_1771, i_13_1772, i_13_1796, i_13_1804, i_13_1827, i_13_1853, i_13_1912, i_13_1930, i_13_2150, i_13_2168, i_13_2183, i_13_2200, i_13_2201, i_13_2228, i_13_2264, i_13_2311, i_13_2425, i_13_2510, i_13_2542, i_13_2554, i_13_2579, i_13_2633, i_13_2650, i_13_2660, i_13_2695, i_13_2848, i_13_2917, i_13_2920, i_13_3131, i_13_3169, i_13_3220, i_13_3221, i_13_3433, i_13_3523, i_13_3536, i_13_3636, i_13_3722, i_13_3794, i_13_3839, i_13_3901, i_13_4012, i_13_4013, i_13_4193, i_13_4238, i_13_4271, i_13_4408, i_13_4444, i_13_4526, i_13_4544, i_13_4586, i_13_4588, o_13_301);
	kernel_13_302 k_13_302(i_13_29, i_13_48, i_13_69, i_13_70, i_13_124, i_13_140, i_13_160, i_13_231, i_13_240, i_13_245, i_13_313, i_13_380, i_13_385, i_13_447, i_13_610, i_13_645, i_13_688, i_13_742, i_13_762, i_13_870, i_13_1020, i_13_1069, i_13_1084, i_13_1086, i_13_1104, i_13_1123, i_13_1132, i_13_1218, i_13_1221, i_13_1257, i_13_1276, i_13_1312, i_13_1441, i_13_1444, i_13_1507, i_13_1510, i_13_1522, i_13_1529, i_13_1598, i_13_1609, i_13_1626, i_13_1716, i_13_1726, i_13_1798, i_13_1803, i_13_1887, i_13_1932, i_13_1933, i_13_1939, i_13_1947, i_13_1995, i_13_2001, i_13_2032, i_13_2122, i_13_2175, i_13_2193, i_13_2194, i_13_2235, i_13_2236, i_13_2266, i_13_2459, i_13_2472, i_13_2679, i_13_2680, i_13_2697, i_13_2724, i_13_2748, i_13_2757, i_13_2810, i_13_2855, i_13_2929, i_13_3003, i_13_3031, i_13_3044, i_13_3147, i_13_3211, i_13_3290, i_13_3370, i_13_3417, i_13_3418, i_13_3553, i_13_3616, i_13_3637, i_13_3640, i_13_3796, i_13_3822, i_13_3823, i_13_3891, i_13_3892, i_13_3930, i_13_4038, i_13_4039, i_13_4056, i_13_4083, i_13_4084, i_13_4308, i_13_4312, i_13_4596, i_13_4597, i_13_4606, o_13_302);
	kernel_13_303 k_13_303(i_13_103, i_13_105, i_13_106, i_13_159, i_13_160, i_13_175, i_13_227, i_13_339, i_13_357, i_13_372, i_13_421, i_13_456, i_13_457, i_13_471, i_13_486, i_13_492, i_13_696, i_13_697, i_13_735, i_13_797, i_13_825, i_13_949, i_13_1086, i_13_1131, i_13_1213, i_13_1299, i_13_1302, i_13_1303, i_13_1346, i_13_1347, i_13_1348, i_13_1437, i_13_1446, i_13_1463, i_13_1464, i_13_1473, i_13_1474, i_13_1528, i_13_1609, i_13_1721, i_13_1722, i_13_1743, i_13_1771, i_13_1815, i_13_1816, i_13_1883, i_13_1951, i_13_2031, i_13_2045, i_13_2056, i_13_2103, i_13_2110, i_13_2223, i_13_2238, i_13_2239, i_13_2378, i_13_2404, i_13_2407, i_13_2422, i_13_2445, i_13_2446, i_13_2553, i_13_2697, i_13_2715, i_13_2716, i_13_2823, i_13_2824, i_13_2846, i_13_2911, i_13_2922, i_13_3009, i_13_3058, i_13_3112, i_13_3219, i_13_3220, i_13_3255, i_13_3390, i_13_3391, i_13_3418, i_13_3420, i_13_3531, i_13_3595, i_13_3612, i_13_3621, i_13_3622, i_13_3706, i_13_3741, i_13_3985, i_13_3999, i_13_4042, i_13_4083, i_13_4092, i_13_4236, i_13_4237, i_13_4326, i_13_4327, i_13_4398, i_13_4512, i_13_4521, i_13_4567, o_13_303);
	kernel_13_304 k_13_304(i_13_59, i_13_70, i_13_112, i_13_119, i_13_157, i_13_171, i_13_172, i_13_175, i_13_184, i_13_280, i_13_282, i_13_283, i_13_313, i_13_319, i_13_370, i_13_489, i_13_523, i_13_532, i_13_598, i_13_607, i_13_657, i_13_658, i_13_660, i_13_675, i_13_694, i_13_695, i_13_939, i_13_1018, i_13_1020, i_13_1066, i_13_1072, i_13_1074, i_13_1075, i_13_1206, i_13_1224, i_13_1225, i_13_1300, i_13_1305, i_13_1422, i_13_1423, i_13_1444, i_13_1494, i_13_1630, i_13_1631, i_13_1632, i_13_1633, i_13_1639, i_13_1657, i_13_1720, i_13_1729, i_13_1732, i_13_1779, i_13_1838, i_13_1936, i_13_1954, i_13_2196, i_13_2235, i_13_2377, i_13_2448, i_13_2449, i_13_2451, i_13_2452, i_13_3141, i_13_3142, i_13_3217, i_13_3244, i_13_3264, i_13_3388, i_13_3447, i_13_3483, i_13_3484, i_13_3538, i_13_3568, i_13_3574, i_13_3612, i_13_3726, i_13_3880, i_13_3888, i_13_3889, i_13_3994, i_13_4017, i_13_4086, i_13_4087, i_13_4186, i_13_4248, i_13_4249, i_13_4251, i_13_4252, i_13_4254, i_13_4258, i_13_4260, i_13_4261, i_13_4393, i_13_4415, i_13_4455, i_13_4521, i_13_4541, i_13_4554, i_13_4558, i_13_4591, o_13_304);
	kernel_13_305 k_13_305(i_13_70, i_13_98, i_13_229, i_13_268, i_13_359, i_13_562, i_13_607, i_13_608, i_13_610, i_13_611, i_13_646, i_13_655, i_13_661, i_13_662, i_13_671, i_13_673, i_13_701, i_13_814, i_13_825, i_13_950, i_13_1024, i_13_1085, i_13_1102, i_13_1120, i_13_1123, i_13_1148, i_13_1167, i_13_1220, i_13_1430, i_13_1660, i_13_1661, i_13_1672, i_13_1727, i_13_1733, i_13_1735, i_13_1736, i_13_1745, i_13_1840, i_13_1841, i_13_1843, i_13_1844, i_13_1858, i_13_2020, i_13_2021, i_13_2024, i_13_2099, i_13_2137, i_13_2173, i_13_2348, i_13_2435, i_13_2471, i_13_2716, i_13_2787, i_13_2885, i_13_2902, i_13_2959, i_13_3029, i_13_3047, i_13_3050, i_13_3092, i_13_3100, i_13_3101, i_13_3145, i_13_3262, i_13_3352, i_13_3417, i_13_3479, i_13_3527, i_13_3613, i_13_3649, i_13_3662, i_13_3667, i_13_3730, i_13_3743, i_13_3751, i_13_3866, i_13_3896, i_13_3910, i_13_3911, i_13_3931, i_13_4063, i_13_4162, i_13_4163, i_13_4166, i_13_4189, i_13_4190, i_13_4192, i_13_4193, i_13_4294, i_13_4296, i_13_4297, i_13_4328, i_13_4343, i_13_4364, i_13_4530, i_13_4594, i_13_4597, i_13_4603, i_13_4604, i_13_4607, o_13_305);
	kernel_13_306 k_13_306(i_13_53, i_13_71, i_13_108, i_13_173, i_13_193, i_13_241, i_13_311, i_13_314, i_13_466, i_13_538, i_13_557, i_13_620, i_13_628, i_13_629, i_13_644, i_13_646, i_13_647, i_13_683, i_13_686, i_13_689, i_13_698, i_13_758, i_13_827, i_13_859, i_13_985, i_13_1066, i_13_1124, i_13_1133, i_13_1151, i_13_1228, i_13_1274, i_13_1277, i_13_1378, i_13_1394, i_13_1459, i_13_1484, i_13_1511, i_13_1549, i_13_1624, i_13_1645, i_13_1646, i_13_1660, i_13_1670, i_13_1673, i_13_1727, i_13_1745, i_13_1796, i_13_1798, i_13_1799, i_13_1889, i_13_1912, i_13_2119, i_13_2134, i_13_2384, i_13_2651, i_13_2654, i_13_2690, i_13_2851, i_13_2852, i_13_2876, i_13_2878, i_13_2906, i_13_2983, i_13_3095, i_13_3097, i_13_3131, i_13_3157, i_13_3265, i_13_3274, i_13_3343, i_13_3356, i_13_3397, i_13_3479, i_13_3575, i_13_3663, i_13_3742, i_13_3743, i_13_3785, i_13_3797, i_13_3842, i_13_3869, i_13_3896, i_13_3931, i_13_3941, i_13_3995, i_13_4033, i_13_4055, i_13_4059, i_13_4084, i_13_4085, i_13_4190, i_13_4297, i_13_4298, i_13_4301, i_13_4436, i_13_4448, i_13_4463, i_13_4530, i_13_4598, i_13_4607, o_13_306);
	kernel_13_307 k_13_307(i_13_31, i_13_32, i_13_64, i_13_121, i_13_207, i_13_208, i_13_307, i_13_374, i_13_399, i_13_412, i_13_489, i_13_524, i_13_586, i_13_598, i_13_612, i_13_613, i_13_671, i_13_715, i_13_738, i_13_759, i_13_760, i_13_796, i_13_829, i_13_1066, i_13_1121, i_13_1128, i_13_1129, i_13_1207, i_13_1223, i_13_1281, i_13_1286, i_13_1306, i_13_1372, i_13_1423, i_13_1441, i_13_1507, i_13_1523, i_13_1559, i_13_1562, i_13_1639, i_13_1696, i_13_1697, i_13_1720, i_13_1792, i_13_1795, i_13_1927, i_13_1928, i_13_1945, i_13_1964, i_13_2101, i_13_2126, i_13_2172, i_13_2200, i_13_2237, i_13_2351, i_13_2365, i_13_2377, i_13_2438, i_13_2542, i_13_2552, i_13_2593, i_13_2677, i_13_2719, i_13_2749, i_13_2759, i_13_2771, i_13_2857, i_13_2881, i_13_2882, i_13_3127, i_13_3172, i_13_3242, i_13_3269, i_13_3367, i_13_3438, i_13_3446, i_13_3572, i_13_3591, i_13_3605, i_13_3637, i_13_3638, i_13_3889, i_13_3910, i_13_3916, i_13_3925, i_13_3928, i_13_3934, i_13_4033, i_13_4034, i_13_4036, i_13_4042, i_13_4045, i_13_4052, i_13_4166, i_13_4313, i_13_4337, i_13_4494, i_13_4510, i_13_4522, i_13_4591, o_13_307);
	kernel_13_308 k_13_308(i_13_64, i_13_65, i_13_118, i_13_188, i_13_190, i_13_226, i_13_274, i_13_308, i_13_320, i_13_357, i_13_359, i_13_373, i_13_464, i_13_544, i_13_589, i_13_601, i_13_695, i_13_712, i_13_758, i_13_839, i_13_890, i_13_949, i_13_1100, i_13_1190, i_13_1207, i_13_1208, i_13_1271, i_13_1306, i_13_1307, i_13_1319, i_13_1345, i_13_1346, i_13_1436, i_13_1486, i_13_1504, i_13_1505, i_13_1594, i_13_1595, i_13_1639, i_13_1640, i_13_1688, i_13_1768, i_13_1792, i_13_1831, i_13_1913, i_13_1928, i_13_1948, i_13_2003, i_13_2030, i_13_2053, i_13_2054, i_13_2056, i_13_2099, i_13_2101, i_13_2189, i_13_2281, i_13_2282, i_13_2345, i_13_2398, i_13_2494, i_13_2552, i_13_2674, i_13_2675, i_13_2720, i_13_2846, i_13_2854, i_13_2861, i_13_2900, i_13_2917, i_13_2918, i_13_2983, i_13_3062, i_13_3089, i_13_3136, i_13_3169, i_13_3377, i_13_3380, i_13_3389, i_13_3479, i_13_3595, i_13_3596, i_13_3631, i_13_3730, i_13_3781, i_13_3916, i_13_3935, i_13_3979, i_13_3989, i_13_4034, i_13_4052, i_13_4097, i_13_4127, i_13_4204, i_13_4262, i_13_4394, i_13_4447, i_13_4555, i_13_4586, i_13_4591, i_13_4592, o_13_308);
	kernel_13_309 k_13_309(i_13_72, i_13_121, i_13_156, i_13_175, i_13_192, i_13_207, i_13_244, i_13_264, i_13_265, i_13_336, i_13_354, i_13_367, i_13_372, i_13_381, i_13_462, i_13_463, i_13_516, i_13_588, i_13_607, i_13_660, i_13_670, i_13_768, i_13_811, i_13_813, i_13_831, i_13_1072, i_13_1116, i_13_1200, i_13_1203, i_13_1227, i_13_1228, i_13_1252, i_13_1306, i_13_1344, i_13_1345, i_13_1407, i_13_1488, i_13_1593, i_13_1602, i_13_1633, i_13_1723, i_13_1813, i_13_1839, i_13_1840, i_13_1845, i_13_1846, i_13_1996, i_13_2029, i_13_2055, i_13_2124, i_13_2133, i_13_2136, i_13_2142, i_13_2190, i_13_2199, i_13_2200, i_13_2208, i_13_2280, i_13_2281, i_13_2395, i_13_2469, i_13_2506, i_13_2538, i_13_2613, i_13_2820, i_13_2934, i_13_3136, i_13_3241, i_13_3342, i_13_3343, i_13_3370, i_13_3387, i_13_3486, i_13_3502, i_13_3532, i_13_3549, i_13_3550, i_13_3567, i_13_3594, i_13_3595, i_13_3618, i_13_3619, i_13_3630, i_13_3663, i_13_3666, i_13_3667, i_13_3670, i_13_3691, i_13_3934, i_13_3988, i_13_4059, i_13_4060, i_13_4162, i_13_4233, i_13_4311, i_13_4312, i_13_4408, i_13_4449, i_13_4545, i_13_4599, o_13_309);
	kernel_13_310 k_13_310(i_13_71, i_13_79, i_13_125, i_13_139, i_13_172, i_13_175, i_13_179, i_13_205, i_13_279, i_13_285, i_13_310, i_13_313, i_13_358, i_13_373, i_13_448, i_13_522, i_13_538, i_13_604, i_13_607, i_13_646, i_13_657, i_13_672, i_13_682, i_13_683, i_13_685, i_13_688, i_13_691, i_13_820, i_13_844, i_13_1123, i_13_1124, i_13_1215, i_13_1224, i_13_1275, i_13_1276, i_13_1277, i_13_1286, i_13_1305, i_13_1311, i_13_1501, i_13_1511, i_13_1599, i_13_1645, i_13_1672, i_13_1732, i_13_1771, i_13_1799, i_13_1881, i_13_1886, i_13_1934, i_13_2175, i_13_2481, i_13_2646, i_13_2650, i_13_2677, i_13_2680, i_13_2698, i_13_2851, i_13_2878, i_13_2916, i_13_2938, i_13_3014, i_13_3204, i_13_3217, i_13_3235, i_13_3270, i_13_3271, i_13_3275, i_13_3356, i_13_3392, i_13_3418, i_13_3421, i_13_3574, i_13_3652, i_13_3742, i_13_3761, i_13_3895, i_13_3994, i_13_4083, i_13_4084, i_13_4186, i_13_4248, i_13_4251, i_13_4252, i_13_4260, i_13_4293, i_13_4296, i_13_4306, i_13_4307, i_13_4309, i_13_4400, i_13_4435, i_13_4446, i_13_4447, i_13_4557, i_13_4590, i_13_4593, i_13_4594, i_13_4597, i_13_4598, o_13_310);
	kernel_13_311 k_13_311(i_13_75, i_13_76, i_13_79, i_13_94, i_13_95, i_13_122, i_13_143, i_13_166, i_13_193, i_13_322, i_13_406, i_13_518, i_13_586, i_13_698, i_13_700, i_13_701, i_13_827, i_13_841, i_13_932, i_13_943, i_13_979, i_13_1025, i_13_1078, i_13_1079, i_13_1084, i_13_1115, i_13_1209, i_13_1276, i_13_1330, i_13_1408, i_13_1429, i_13_1430, i_13_1439, i_13_1546, i_13_1596, i_13_1610, i_13_1632, i_13_1636, i_13_1675, i_13_1777, i_13_1778, i_13_1831, i_13_1888, i_13_1908, i_13_1947, i_13_2028, i_13_2119, i_13_2343, i_13_2450, i_13_2455, i_13_2610, i_13_2618, i_13_2709, i_13_2788, i_13_2858, i_13_2880, i_13_2887, i_13_2888, i_13_2919, i_13_2955, i_13_2959, i_13_2983, i_13_3141, i_13_3208, i_13_3211, i_13_3244, i_13_3437, i_13_3448, i_13_3451, i_13_3454, i_13_3455, i_13_3464, i_13_3482, i_13_3486, i_13_3526, i_13_3528, i_13_3532, i_13_3571, i_13_3572, i_13_3576, i_13_3618, i_13_3640, i_13_3649, i_13_3688, i_13_3767, i_13_3783, i_13_3799, i_13_3837, i_13_3846, i_13_3888, i_13_3967, i_13_4009, i_13_4086, i_13_4170, i_13_4190, i_13_4248, i_13_4252, i_13_4265, i_13_4301, i_13_4451, o_13_311);
	kernel_13_312 k_13_312(i_13_25, i_13_30, i_13_48, i_13_69, i_13_70, i_13_177, i_13_186, i_13_193, i_13_321, i_13_381, i_13_411, i_13_417, i_13_492, i_13_498, i_13_570, i_13_609, i_13_645, i_13_678, i_13_699, i_13_759, i_13_760, i_13_762, i_13_763, i_13_870, i_13_933, i_13_994, i_13_1021, i_13_1083, i_13_1084, i_13_1086, i_13_1095, i_13_1104, i_13_1131, i_13_1132, i_13_1224, i_13_1302, i_13_1303, i_13_1308, i_13_1347, i_13_1407, i_13_1525, i_13_1528, i_13_1551, i_13_1605, i_13_1632, i_13_1644, i_13_1714, i_13_1716, i_13_1789, i_13_1797, i_13_1798, i_13_1806, i_13_1807, i_13_1843, i_13_1942, i_13_1992, i_13_1995, i_13_2023, i_13_2055, i_13_2122, i_13_2224, i_13_2472, i_13_2473, i_13_2505, i_13_2536, i_13_2541, i_13_2542, i_13_2722, i_13_2757, i_13_2955, i_13_3022, i_13_3030, i_13_3031, i_13_3118, i_13_3121, i_13_3198, i_13_3264, i_13_3346, i_13_3375, i_13_3399, i_13_3453, i_13_3702, i_13_3739, i_13_3804, i_13_3822, i_13_4038, i_13_4081, i_13_4090, i_13_4093, i_13_4117, i_13_4189, i_13_4233, i_13_4255, i_13_4272, i_13_4273, i_13_4308, i_13_4336, i_13_4596, i_13_4605, i_13_4606, o_13_312);
	kernel_13_313 k_13_313(i_13_136, i_13_137, i_13_139, i_13_140, i_13_175, i_13_226, i_13_227, i_13_230, i_13_268, i_13_362, i_13_419, i_13_533, i_13_536, i_13_641, i_13_695, i_13_824, i_13_850, i_13_892, i_13_976, i_13_982, i_13_985, i_13_1201, i_13_1217, i_13_1219, i_13_1220, i_13_1274, i_13_1283, i_13_1343, i_13_1467, i_13_1607, i_13_1711, i_13_1712, i_13_1722, i_13_1723, i_13_1778, i_13_1882, i_13_1883, i_13_1885, i_13_1886, i_13_1958, i_13_2003, i_13_2098, i_13_2189, i_13_2210, i_13_2297, i_13_2426, i_13_2549, i_13_2647, i_13_2648, i_13_2708, i_13_2747, i_13_2846, i_13_2848, i_13_2855, i_13_2858, i_13_2872, i_13_2885, i_13_2909, i_13_2935, i_13_2956, i_13_2983, i_13_3001, i_13_3004, i_13_3005, i_13_3010, i_13_3037, i_13_3038, i_13_3056, i_13_3109, i_13_3143, i_13_3322, i_13_3370, i_13_3382, i_13_3385, i_13_3386, i_13_3425, i_13_3439, i_13_3449, i_13_3487, i_13_3503, i_13_3542, i_13_3743, i_13_3820, i_13_3836, i_13_3839, i_13_3865, i_13_4016, i_13_4054, i_13_4060, i_13_4063, i_13_4181, i_13_4190, i_13_4211, i_13_4342, i_13_4388, i_13_4394, i_13_4411, i_13_4414, i_13_4522, i_13_4531, o_13_313);
	kernel_13_314 k_13_314(i_13_45, i_13_99, i_13_102, i_13_157, i_13_192, i_13_193, i_13_195, i_13_333, i_13_442, i_13_450, i_13_451, i_13_577, i_13_612, i_13_624, i_13_640, i_13_657, i_13_714, i_13_721, i_13_858, i_13_946, i_13_948, i_13_955, i_13_982, i_13_1062, i_13_1116, i_13_1147, i_13_1224, i_13_1225, i_13_1227, i_13_1231, i_13_1282, i_13_1297, i_13_1314, i_13_1345, i_13_1407, i_13_1435, i_13_1443, i_13_1458, i_13_1468, i_13_1488, i_13_1494, i_13_1566, i_13_1567, i_13_1764, i_13_1776, i_13_1800, i_13_1801, i_13_1803, i_13_1891, i_13_1926, i_13_1990, i_13_1999, i_13_2056, i_13_2107, i_13_2137, i_13_2145, i_13_2205, i_13_2209, i_13_2296, i_13_2425, i_13_2532, i_13_2568, i_13_2613, i_13_2614, i_13_2691, i_13_2745, i_13_2820, i_13_3006, i_13_3024, i_13_3052, i_13_3055, i_13_3144, i_13_3214, i_13_3267, i_13_3286, i_13_3339, i_13_3342, i_13_3420, i_13_3421, i_13_3474, i_13_3486, i_13_3753, i_13_3873, i_13_3978, i_13_4017, i_13_4086, i_13_4087, i_13_4230, i_13_4231, i_13_4233, i_13_4266, i_13_4267, i_13_4302, i_13_4339, i_13_4341, i_13_4404, i_13_4431, i_13_4468, i_13_4509, i_13_4513, o_13_314);
	kernel_13_315 k_13_315(i_13_26, i_13_69, i_13_93, i_13_96, i_13_97, i_13_106, i_13_107, i_13_117, i_13_121, i_13_159, i_13_180, i_13_183, i_13_352, i_13_386, i_13_409, i_13_410, i_13_415, i_13_457, i_13_529, i_13_565, i_13_654, i_13_697, i_13_746, i_13_760, i_13_800, i_13_832, i_13_933, i_13_944, i_13_1086, i_13_1087, i_13_1088, i_13_1097, i_13_1303, i_13_1491, i_13_1507, i_13_1529, i_13_1725, i_13_1789, i_13_1790, i_13_1797, i_13_1807, i_13_1815, i_13_1995, i_13_1996, i_13_2122, i_13_2177, i_13_2211, i_13_2212, i_13_2239, i_13_2240, i_13_2303, i_13_2429, i_13_2614, i_13_2713, i_13_2716, i_13_2760, i_13_2848, i_13_2942, i_13_3022, i_13_3030, i_13_3066, i_13_3103, i_13_3147, i_13_3153, i_13_3237, i_13_3326, i_13_3345, i_13_3391, i_13_3399, i_13_3400, i_13_3525, i_13_3527, i_13_3580, i_13_3607, i_13_3686, i_13_3702, i_13_3739, i_13_3797, i_13_3846, i_13_3985, i_13_3986, i_13_4006, i_13_4008, i_13_4009, i_13_4046, i_13_4047, i_13_4094, i_13_4193, i_13_4235, i_13_4238, i_13_4261, i_13_4264, i_13_4273, i_13_4310, i_13_4327, i_13_4343, i_13_4399, i_13_4416, i_13_4417, i_13_4463, o_13_315);
	kernel_13_316 k_13_316(i_13_40, i_13_58, i_13_259, i_13_276, i_13_369, i_13_450, i_13_513, i_13_526, i_13_552, i_13_604, i_13_606, i_13_607, i_13_610, i_13_657, i_13_658, i_13_660, i_13_661, i_13_663, i_13_670, i_13_678, i_13_829, i_13_840, i_13_931, i_13_936, i_13_939, i_13_1056, i_13_1059, i_13_1060, i_13_1072, i_13_1102, i_13_1119, i_13_1147, i_13_1516, i_13_1534, i_13_1606, i_13_1659, i_13_1660, i_13_1663, i_13_1729, i_13_1731, i_13_1732, i_13_1764, i_13_1767, i_13_1891, i_13_1897, i_13_1911, i_13_1998, i_13_1999, i_13_2001, i_13_2019, i_13_2020, i_13_2148, i_13_2425, i_13_2437, i_13_2448, i_13_2467, i_13_2469, i_13_2514, i_13_2515, i_13_2626, i_13_2740, i_13_2910, i_13_2955, i_13_2958, i_13_3027, i_13_3046, i_13_3072, i_13_3073, i_13_3108, i_13_3127, i_13_3261, i_13_3262, i_13_3486, i_13_3549, i_13_3550, i_13_3565, i_13_3567, i_13_3573, i_13_3648, i_13_3819, i_13_3891, i_13_3897, i_13_3909, i_13_3910, i_13_3990, i_13_4158, i_13_4159, i_13_4161, i_13_4162, i_13_4251, i_13_4293, i_13_4333, i_13_4336, i_13_4365, i_13_4368, i_13_4369, i_13_4434, i_13_4510, i_13_4602, i_13_4603, o_13_316);
	kernel_13_317 k_13_317(i_13_32, i_13_69, i_13_93, i_13_94, i_13_120, i_13_121, i_13_157, i_13_229, i_13_276, i_13_382, i_13_446, i_13_447, i_13_508, i_13_542, i_13_564, i_13_672, i_13_697, i_13_732, i_13_733, i_13_886, i_13_951, i_13_952, i_13_1185, i_13_1226, i_13_1231, i_13_1303, i_13_1318, i_13_1443, i_13_1444, i_13_1446, i_13_1498, i_13_1602, i_13_1626, i_13_1632, i_13_1758, i_13_1786, i_13_1813, i_13_2012, i_13_2173, i_13_2175, i_13_2176, i_13_2189, i_13_2208, i_13_2209, i_13_2262, i_13_2424, i_13_2425, i_13_2427, i_13_2436, i_13_2463, i_13_2541, i_13_2565, i_13_2581, i_13_2698, i_13_2749, i_13_2857, i_13_2939, i_13_3000, i_13_3004, i_13_3019, i_13_3020, i_13_3037, i_13_3063, i_13_3066, i_13_3067, i_13_3102, i_13_3129, i_13_3130, i_13_3147, i_13_3160, i_13_3165, i_13_3274, i_13_3287, i_13_3307, i_13_3399, i_13_3417, i_13_3418, i_13_3424, i_13_3426, i_13_3427, i_13_3441, i_13_3534, i_13_3541, i_13_3702, i_13_3739, i_13_3801, i_13_3843, i_13_3844, i_13_3980, i_13_3990, i_13_4008, i_13_4009, i_13_4021, i_13_4054, i_13_4251, i_13_4341, i_13_4353, i_13_4380, i_13_4560, i_13_4561, o_13_317);
	kernel_13_318 k_13_318(i_13_73, i_13_74, i_13_121, i_13_139, i_13_182, i_13_184, i_13_185, i_13_193, i_13_229, i_13_235, i_13_253, i_13_355, i_13_415, i_13_469, i_13_470, i_13_590, i_13_668, i_13_694, i_13_695, i_13_743, i_13_829, i_13_947, i_13_1072, i_13_1073, i_13_1118, i_13_1145, i_13_1208, i_13_1247, i_13_1307, i_13_1408, i_13_1424, i_13_1522, i_13_1523, i_13_1536, i_13_1549, i_13_1658, i_13_1667, i_13_1723, i_13_1742, i_13_1774, i_13_1849, i_13_1919, i_13_1998, i_13_2000, i_13_2017, i_13_2021, i_13_2056, i_13_2057, i_13_2126, i_13_2143, i_13_2144, i_13_2308, i_13_2425, i_13_2444, i_13_2449, i_13_2450, i_13_2512, i_13_2513, i_13_2539, i_13_2660, i_13_2692, i_13_2855, i_13_2881, i_13_2882, i_13_2907, i_13_3010, i_13_3025, i_13_3037, i_13_3128, i_13_3254, i_13_3269, i_13_3415, i_13_3416, i_13_3610, i_13_3620, i_13_3683, i_13_3863, i_13_3865, i_13_3874, i_13_3916, i_13_3919, i_13_3921, i_13_3988, i_13_4009, i_13_4118, i_13_4180, i_13_4253, i_13_4262, i_13_4271, i_13_4330, i_13_4331, i_13_4366, i_13_4430, i_13_4529, i_13_4538, i_13_4583, i_13_4591, i_13_4592, i_13_4601, i_13_4604, o_13_318);
	kernel_13_319 k_13_319(i_13_95, i_13_136, i_13_137, i_13_139, i_13_140, i_13_202, i_13_226, i_13_230, i_13_262, i_13_383, i_13_384, i_13_418, i_13_607, i_13_618, i_13_686, i_13_688, i_13_725, i_13_779, i_13_824, i_13_985, i_13_1094, i_13_1217, i_13_1265, i_13_1270, i_13_1274, i_13_1282, i_13_1442, i_13_1462, i_13_1499, i_13_1552, i_13_1712, i_13_1723, i_13_1778, i_13_1802, i_13_1832, i_13_1837, i_13_1882, i_13_1883, i_13_1885, i_13_1886, i_13_1993, i_13_1994, i_13_1999, i_13_2000, i_13_2018, i_13_2054, i_13_2120, i_13_2170, i_13_2192, i_13_2207, i_13_2224, i_13_2314, i_13_2426, i_13_2593, i_13_2647, i_13_2648, i_13_2651, i_13_2845, i_13_2848, i_13_2849, i_13_2857, i_13_2875, i_13_2885, i_13_3044, i_13_3065, i_13_3091, i_13_3143, i_13_3154, i_13_3164, i_13_3322, i_13_3368, i_13_3389, i_13_3424, i_13_3425, i_13_3444, i_13_3478, i_13_3487, i_13_3488, i_13_3556, i_13_3686, i_13_3791, i_13_3794, i_13_3799, i_13_3836, i_13_3841, i_13_3992, i_13_4025, i_13_4051, i_13_4097, i_13_4124, i_13_4186, i_13_4187, i_13_4235, i_13_4295, i_13_4301, i_13_4369, i_13_4394, i_13_4397, i_13_4501, i_13_4568, o_13_319);
	kernel_13_320 k_13_320(i_13_61, i_13_65, i_13_76, i_13_111, i_13_112, i_13_186, i_13_187, i_13_283, i_13_309, i_13_382, i_13_406, i_13_473, i_13_532, i_13_571, i_13_573, i_13_574, i_13_623, i_13_643, i_13_646, i_13_717, i_13_780, i_13_814, i_13_889, i_13_1073, i_13_1201, i_13_1210, i_13_1271, i_13_1388, i_13_1390, i_13_1426, i_13_1492, i_13_1525, i_13_1528, i_13_1542, i_13_1633, i_13_1640, i_13_1641, i_13_1642, i_13_1677, i_13_1680, i_13_1721, i_13_1749, i_13_1793, i_13_1803, i_13_1804, i_13_1870, i_13_1993, i_13_2014, i_13_2103, i_13_2197, i_13_2211, i_13_2212, i_13_2262, i_13_2272, i_13_2407, i_13_2428, i_13_2452, i_13_2535, i_13_2616, i_13_2649, i_13_2653, i_13_2679, i_13_2846, i_13_3027, i_13_3028, i_13_3089, i_13_3166, i_13_3207, i_13_3208, i_13_3292, i_13_3378, i_13_3387, i_13_3424, i_13_3426, i_13_3476, i_13_3480, i_13_3561, i_13_3610, i_13_3649, i_13_3755, i_13_3836, i_13_3859, i_13_3904, i_13_3991, i_13_3994, i_13_4011, i_13_4012, i_13_4021, i_13_4073, i_13_4079, i_13_4080, i_13_4083, i_13_4183, i_13_4188, i_13_4264, i_13_4295, i_13_4411, i_13_4558, i_13_4587, i_13_4596, o_13_320);
	kernel_13_321 k_13_321(i_13_36, i_13_39, i_13_40, i_13_42, i_13_49, i_13_70, i_13_137, i_13_306, i_13_454, i_13_492, i_13_585, i_13_643, i_13_688, i_13_689, i_13_690, i_13_697, i_13_726, i_13_823, i_13_826, i_13_1084, i_13_1271, i_13_1272, i_13_1278, i_13_1279, i_13_1299, i_13_1303, i_13_1347, i_13_1391, i_13_1465, i_13_1593, i_13_1600, i_13_1638, i_13_1642, i_13_1669, i_13_1672, i_13_1759, i_13_1792, i_13_1831, i_13_1837, i_13_1845, i_13_1884, i_13_1885, i_13_2059, i_13_2082, i_13_2104, i_13_2140, i_13_2161, i_13_2199, i_13_2239, i_13_2378, i_13_2380, i_13_2434, i_13_2554, i_13_2589, i_13_2650, i_13_2652, i_13_2653, i_13_2694, i_13_2761, i_13_2823, i_13_2824, i_13_2848, i_13_2871, i_13_3001, i_13_3006, i_13_3114, i_13_3130, i_13_3151, i_13_3156, i_13_3387, i_13_3388, i_13_3390, i_13_3391, i_13_3394, i_13_3538, i_13_3541, i_13_3597, i_13_3633, i_13_3766, i_13_3816, i_13_3874, i_13_3877, i_13_3895, i_13_3912, i_13_3925, i_13_4014, i_13_4039, i_13_4162, i_13_4187, i_13_4197, i_13_4203, i_13_4297, i_13_4341, i_13_4351, i_13_4356, i_13_4368, i_13_4369, i_13_4381, i_13_4429, i_13_4554, o_13_321);
	kernel_13_322 k_13_322(i_13_45, i_13_103, i_13_120, i_13_139, i_13_172, i_13_189, i_13_202, i_13_229, i_13_408, i_13_414, i_13_549, i_13_568, i_13_604, i_13_606, i_13_625, i_13_642, i_13_643, i_13_648, i_13_657, i_13_684, i_13_685, i_13_796, i_13_936, i_13_982, i_13_1071, i_13_1191, i_13_1225, i_13_1228, i_13_1272, i_13_1282, i_13_1300, i_13_1404, i_13_1432, i_13_1498, i_13_1521, i_13_1548, i_13_1560, i_13_1629, i_13_1674, i_13_1677, i_13_1729, i_13_1750, i_13_1767, i_13_1768, i_13_1795, i_13_1803, i_13_1804, i_13_1808, i_13_1854, i_13_1896, i_13_1911, i_13_2001, i_13_2019, i_13_2020, i_13_2047, i_13_2119, i_13_2286, i_13_2314, i_13_2361, i_13_2469, i_13_2470, i_13_2542, i_13_2578, i_13_2691, i_13_2979, i_13_3000, i_13_3006, i_13_3009, i_13_3027, i_13_3028, i_13_3105, i_13_3204, i_13_3205, i_13_3208, i_13_3261, i_13_3396, i_13_3420, i_13_3475, i_13_3483, i_13_3522, i_13_3546, i_13_3573, i_13_3657, i_13_3811, i_13_3819, i_13_3820, i_13_3897, i_13_3898, i_13_3907, i_13_3978, i_13_3990, i_13_4248, i_13_4251, i_13_4269, i_13_4332, i_13_4392, i_13_4404, i_13_4582, i_13_4594, i_13_4603, o_13_322);
	kernel_13_323 k_13_323(i_13_112, i_13_142, i_13_143, i_13_188, i_13_203, i_13_229, i_13_232, i_13_233, i_13_283, i_13_341, i_13_428, i_13_607, i_13_619, i_13_643, i_13_644, i_13_647, i_13_689, i_13_692, i_13_827, i_13_859, i_13_887, i_13_931, i_13_941, i_13_1079, i_13_1120, i_13_1121, i_13_1124, i_13_1147, i_13_1204, i_13_1276, i_13_1277, i_13_1283, i_13_1346, i_13_1411, i_13_1426, i_13_1448, i_13_1502, i_13_1520, i_13_1637, i_13_1714, i_13_1715, i_13_1726, i_13_1786, i_13_1790, i_13_1796, i_13_1885, i_13_1994, i_13_2005, i_13_2056, i_13_2137, i_13_2138, i_13_2186, i_13_2212, i_13_2213, i_13_2263, i_13_2408, i_13_2428, i_13_2429, i_13_2464, i_13_2542, i_13_2597, i_13_2614, i_13_2617, i_13_2650, i_13_2651, i_13_2654, i_13_2848, i_13_2857, i_13_3040, i_13_3041, i_13_3257, i_13_3308, i_13_3389, i_13_3392, i_13_3425, i_13_3427, i_13_3428, i_13_3482, i_13_3541, i_13_3661, i_13_3724, i_13_3725, i_13_3733, i_13_3856, i_13_3865, i_13_4012, i_13_4013, i_13_4018, i_13_4019, i_13_4057, i_13_4081, i_13_4235, i_13_4307, i_13_4333, i_13_4334, i_13_4369, i_13_4370, i_13_4415, i_13_4534, i_13_4595, o_13_323);
	kernel_13_324 k_13_324(i_13_37, i_13_64, i_13_121, i_13_274, i_13_280, i_13_331, i_13_338, i_13_401, i_13_463, i_13_526, i_13_561, i_13_562, i_13_589, i_13_608, i_13_662, i_13_694, i_13_724, i_13_823, i_13_914, i_13_1066, i_13_1256, i_13_1309, i_13_1310, i_13_1327, i_13_1483, i_13_1499, i_13_1561, i_13_1594, i_13_1595, i_13_1624, i_13_1639, i_13_1661, i_13_1684, i_13_1729, i_13_1732, i_13_1775, i_13_1778, i_13_1793, i_13_1795, i_13_1882, i_13_1883, i_13_1885, i_13_1925, i_13_1927, i_13_1942, i_13_1943, i_13_1999, i_13_2233, i_13_2380, i_13_2443, i_13_2558, i_13_2585, i_13_2650, i_13_2651, i_13_2821, i_13_2872, i_13_2900, i_13_2914, i_13_2983, i_13_3109, i_13_3142, i_13_3163, i_13_3215, i_13_3235, i_13_3271, i_13_3289, i_13_3388, i_13_3389, i_13_3395, i_13_3523, i_13_3538, i_13_3539, i_13_3542, i_13_3662, i_13_3667, i_13_3668, i_13_3728, i_13_3730, i_13_3731, i_13_3739, i_13_3740, i_13_3766, i_13_3792, i_13_3803, i_13_3901, i_13_3904, i_13_3916, i_13_3935, i_13_3989, i_13_4099, i_13_4162, i_13_4324, i_13_4351, i_13_4364, i_13_4369, i_13_4379, i_13_4396, i_13_4443, i_13_4540, i_13_4567, o_13_324);
	kernel_13_325 k_13_325(i_13_61, i_13_62, i_13_76, i_13_106, i_13_112, i_13_166, i_13_169, i_13_193, i_13_220, i_13_382, i_13_484, i_13_535, i_13_544, i_13_573, i_13_574, i_13_575, i_13_601, i_13_728, i_13_815, i_13_895, i_13_914, i_13_1040, i_13_1093, i_13_1120, i_13_1124, i_13_1258, i_13_1277, i_13_1393, i_13_1394, i_13_1411, i_13_1466, i_13_1483, i_13_1484, i_13_1537, i_13_1561, i_13_1628, i_13_1643, i_13_1660, i_13_1691, i_13_1723, i_13_1726, i_13_1727, i_13_1750, i_13_1760, i_13_1771, i_13_1781, i_13_1786, i_13_1789, i_13_1796, i_13_1804, i_13_1834, i_13_1858, i_13_1894, i_13_1907, i_13_2002, i_13_2005, i_13_2041, i_13_2049, i_13_2150, i_13_2168, i_13_2212, i_13_2213, i_13_2263, i_13_2408, i_13_2446, i_13_2542, i_13_2618, i_13_2633, i_13_2642, i_13_2650, i_13_2654, i_13_2687, i_13_2750, i_13_2767, i_13_2785, i_13_3001, i_13_3027, i_13_3041, i_13_3157, i_13_3158, i_13_3200, i_13_3238, i_13_3308, i_13_3427, i_13_3433, i_13_3469, i_13_3472, i_13_3522, i_13_3527, i_13_3562, i_13_3730, i_13_3794, i_13_3884, i_13_3887, i_13_3976, i_13_4012, i_13_4081, i_13_4156, i_13_4157, i_13_4325, o_13_325);
	kernel_13_326 k_13_326(i_13_48, i_13_72, i_13_73, i_13_77, i_13_162, i_13_217, i_13_226, i_13_286, i_13_370, i_13_406, i_13_463, i_13_480, i_13_558, i_13_582, i_13_583, i_13_651, i_13_652, i_13_659, i_13_675, i_13_676, i_13_696, i_13_811, i_13_939, i_13_1071, i_13_1074, i_13_1116, i_13_1141, i_13_1143, i_13_1144, i_13_1145, i_13_1200, i_13_1281, i_13_1362, i_13_1437, i_13_1549, i_13_1632, i_13_1656, i_13_1657, i_13_1658, i_13_1720, i_13_1837, i_13_1839, i_13_1841, i_13_2017, i_13_2047, i_13_2241, i_13_2317, i_13_2394, i_13_2404, i_13_2451, i_13_2452, i_13_2468, i_13_2511, i_13_2550, i_13_2745, i_13_2754, i_13_2791, i_13_2844, i_13_2845, i_13_2854, i_13_2883, i_13_2925, i_13_2944, i_13_2955, i_13_2959, i_13_2986, i_13_2997, i_13_2998, i_13_3096, i_13_3100, i_13_3105, i_13_3204, i_13_3447, i_13_3448, i_13_3501, i_13_3522, i_13_3549, i_13_3567, i_13_3568, i_13_3577, i_13_3645, i_13_3646, i_13_3663, i_13_3735, i_13_3847, i_13_3891, i_13_3907, i_13_3933, i_13_4017, i_13_4095, i_13_4160, i_13_4186, i_13_4258, i_13_4311, i_13_4329, i_13_4590, i_13_4591, i_13_4599, i_13_4600, i_13_4601, o_13_326);
	kernel_13_327 k_13_327(i_13_48, i_13_67, i_13_69, i_13_186, i_13_229, i_13_258, i_13_285, i_13_310, i_13_411, i_13_438, i_13_520, i_13_610, i_13_616, i_13_627, i_13_628, i_13_760, i_13_762, i_13_853, i_13_934, i_13_939, i_13_1023, i_13_1105, i_13_1132, i_13_1149, i_13_1150, i_13_1191, i_13_1227, i_13_1317, i_13_1381, i_13_1402, i_13_1429, i_13_1482, i_13_1509, i_13_1537, i_13_1563, i_13_1596, i_13_1597, i_13_1610, i_13_1644, i_13_1651, i_13_1744, i_13_1753, i_13_1770, i_13_1794, i_13_1798, i_13_1829, i_13_1838, i_13_1884, i_13_1922, i_13_1923, i_13_1947, i_13_2022, i_13_2122, i_13_2199, i_13_2311, i_13_2427, i_13_2428, i_13_2454, i_13_2472, i_13_2473, i_13_2506, i_13_2517, i_13_2742, i_13_2743, i_13_2770, i_13_2940, i_13_2968, i_13_3009, i_13_3012, i_13_3030, i_13_3031, i_13_3075, i_13_3076, i_13_3091, i_13_3093, i_13_3211, i_13_3264, i_13_3273, i_13_3292, i_13_3345, i_13_3354, i_13_3381, i_13_3382, i_13_3418, i_13_3435, i_13_3540, i_13_3576, i_13_3759, i_13_3822, i_13_3900, i_13_3929, i_13_4036, i_13_4083, i_13_4164, i_13_4272, i_13_4362, i_13_4450, i_13_4497, i_13_4605, i_13_4606, o_13_327);
	kernel_13_328 k_13_328(i_13_18, i_13_58, i_13_102, i_13_130, i_13_131, i_13_132, i_13_223, i_13_355, i_13_371, i_13_374, i_13_415, i_13_489, i_13_614, i_13_736, i_13_955, i_13_956, i_13_1084, i_13_1100, i_13_1128, i_13_1227, i_13_1256, i_13_1300, i_13_1302, i_13_1305, i_13_1306, i_13_1322, i_13_1409, i_13_1445, i_13_1451, i_13_1472, i_13_1494, i_13_1503, i_13_1517, i_13_1522, i_13_1551, i_13_1552, i_13_1553, i_13_1554, i_13_1638, i_13_1639, i_13_1736, i_13_1778, i_13_1801, i_13_1802, i_13_1814, i_13_1846, i_13_1957, i_13_2090, i_13_2093, i_13_2100, i_13_2101, i_13_2142, i_13_2199, i_13_2235, i_13_2236, i_13_2296, i_13_2297, i_13_2522, i_13_2744, i_13_2789, i_13_2821, i_13_2822, i_13_2935, i_13_2936, i_13_2997, i_13_3024, i_13_3064, i_13_3100, i_13_3119, i_13_3145, i_13_3206, i_13_3241, i_13_3242, i_13_3308, i_13_3383, i_13_3388, i_13_3420, i_13_3433, i_13_3451, i_13_3477, i_13_3523, i_13_3537, i_13_3539, i_13_3617, i_13_3638, i_13_3685, i_13_3686, i_13_3754, i_13_3855, i_13_3856, i_13_3857, i_13_3916, i_13_4018, i_13_4060, i_13_4311, i_13_4312, i_13_4378, i_13_4382, i_13_4509, i_13_4592, o_13_328);
	kernel_13_329 k_13_329(i_13_45, i_13_46, i_13_169, i_13_175, i_13_179, i_13_187, i_13_283, i_13_310, i_13_343, i_13_444, i_13_515, i_13_532, i_13_554, i_13_567, i_13_568, i_13_574, i_13_649, i_13_719, i_13_730, i_13_847, i_13_854, i_13_886, i_13_986, i_13_1037, i_13_1072, i_13_1105, i_13_1228, i_13_1232, i_13_1309, i_13_1316, i_13_1550, i_13_1729, i_13_1741, i_13_1765, i_13_1804, i_13_1805, i_13_1822, i_13_1832, i_13_1846, i_13_1850, i_13_1852, i_13_1895, i_13_1992, i_13_1996, i_13_2020, i_13_2288, i_13_2314, i_13_2365, i_13_2372, i_13_2408, i_13_2422, i_13_2434, i_13_2443, i_13_2449, i_13_2450, i_13_2470, i_13_2473, i_13_2479, i_13_2680, i_13_2681, i_13_2897, i_13_3010, i_13_3011, i_13_3032, i_13_3110, i_13_3168, i_13_3207, i_13_3208, i_13_3212, i_13_3272, i_13_3400, i_13_3420, i_13_3421, i_13_3483, i_13_3502, i_13_3578, i_13_3637, i_13_3748, i_13_3871, i_13_3872, i_13_3907, i_13_3914, i_13_3955, i_13_4015, i_13_4036, i_13_4041, i_13_4042, i_13_4095, i_13_4190, i_13_4248, i_13_4252, i_13_4253, i_13_4270, i_13_4368, i_13_4369, i_13_4374, i_13_4379, i_13_4441, i_13_4514, i_13_4607, o_13_329);
	kernel_13_330 k_13_330(i_13_50, i_13_80, i_13_201, i_13_203, i_13_229, i_13_286, i_13_421, i_13_535, i_13_626, i_13_661, i_13_792, i_13_823, i_13_847, i_13_850, i_13_851, i_13_867, i_13_869, i_13_941, i_13_1018, i_13_1021, i_13_1022, i_13_1060, i_13_1075, i_13_1076, i_13_1232, i_13_1318, i_13_1427, i_13_1530, i_13_1541, i_13_1549, i_13_1550, i_13_1551, i_13_1598, i_13_1679, i_13_1774, i_13_1780, i_13_1855, i_13_1858, i_13_2030, i_13_2197, i_13_2199, i_13_2200, i_13_2202, i_13_2452, i_13_2539, i_13_2543, i_13_2617, i_13_2703, i_13_2913, i_13_2920, i_13_2999, i_13_3007, i_13_3010, i_13_3011, i_13_3013, i_13_3064, i_13_3087, i_13_3104, i_13_3169, i_13_3172, i_13_3399, i_13_3453, i_13_3454, i_13_3461, i_13_3484, i_13_3486, i_13_3487, i_13_3488, i_13_3535, i_13_3539, i_13_3541, i_13_3542, i_13_3576, i_13_3577, i_13_3578, i_13_3616, i_13_3703, i_13_3730, i_13_3764, i_13_3781, i_13_3782, i_13_3784, i_13_3785, i_13_3854, i_13_3865, i_13_3866, i_13_3868, i_13_3885, i_13_3889, i_13_3892, i_13_3906, i_13_4176, i_13_4179, i_13_4249, i_13_4252, i_13_4256, i_13_4262, i_13_4378, i_13_4379, i_13_4561, o_13_330);
	kernel_13_331 k_13_331(i_13_28, i_13_29, i_13_31, i_13_32, i_13_64, i_13_65, i_13_91, i_13_136, i_13_137, i_13_184, i_13_226, i_13_227, i_13_228, i_13_307, i_13_308, i_13_309, i_13_316, i_13_317, i_13_380, i_13_418, i_13_419, i_13_459, i_13_535, i_13_553, i_13_639, i_13_718, i_13_873, i_13_950, i_13_1075, i_13_1143, i_13_1208, i_13_1216, i_13_1217, i_13_1308, i_13_1318, i_13_1341, i_13_1408, i_13_1422, i_13_1435, i_13_1445, i_13_1526, i_13_1594, i_13_1596, i_13_1678, i_13_1720, i_13_1785, i_13_1841, i_13_1848, i_13_1858, i_13_1922, i_13_1999, i_13_2000, i_13_2002, i_13_2003, i_13_2052, i_13_2055, i_13_2142, i_13_2146, i_13_2174, i_13_2189, i_13_2259, i_13_2280, i_13_2345, i_13_2403, i_13_2422, i_13_2423, i_13_2547, i_13_2552, i_13_2674, i_13_2694, i_13_2710, i_13_2719, i_13_2720, i_13_2740, i_13_2854, i_13_2855, i_13_2857, i_13_2884, i_13_2937, i_13_3034, i_13_3036, i_13_3127, i_13_3204, i_13_3207, i_13_3366, i_13_3487, i_13_3523, i_13_3529, i_13_3663, i_13_3727, i_13_3764, i_13_3902, i_13_3990, i_13_4034, i_13_4036, i_13_4082, i_13_4349, i_13_4351, i_13_4397, i_13_4514, o_13_331);
	kernel_13_332 k_13_332(i_13_16, i_13_40, i_13_119, i_13_138, i_13_139, i_13_141, i_13_225, i_13_231, i_13_273, i_13_369, i_13_431, i_13_447, i_13_469, i_13_537, i_13_613, i_13_646, i_13_690, i_13_691, i_13_717, i_13_727, i_13_760, i_13_780, i_13_811, i_13_894, i_13_940, i_13_984, i_13_1092, i_13_1203, i_13_1221, i_13_1249, i_13_1251, i_13_1260, i_13_1276, i_13_1299, i_13_1383, i_13_1386, i_13_1393, i_13_1464, i_13_1470, i_13_1567, i_13_1642, i_13_1671, i_13_1672, i_13_1713, i_13_1725, i_13_1726, i_13_1731, i_13_1884, i_13_1885, i_13_1887, i_13_1906, i_13_1990, i_13_1996, i_13_2136, i_13_2139, i_13_2167, i_13_2187, i_13_2464, i_13_2470, i_13_2577, i_13_2632, i_13_2649, i_13_2650, i_13_2652, i_13_2653, i_13_2680, i_13_2709, i_13_2755, i_13_2847, i_13_2877, i_13_2884, i_13_2914, i_13_3009, i_13_3108, i_13_3174, i_13_3219, i_13_3273, i_13_3279, i_13_3387, i_13_3391, i_13_3432, i_13_3474, i_13_3487, i_13_3528, i_13_3532, i_13_3682, i_13_3766, i_13_3793, i_13_3801, i_13_3838, i_13_3874, i_13_3906, i_13_4126, i_13_4156, i_13_4162, i_13_4308, i_13_4371, i_13_4443, i_13_4521, i_13_4533, o_13_332);
	kernel_13_333 k_13_333(i_13_34, i_13_35, i_13_74, i_13_104, i_13_117, i_13_118, i_13_122, i_13_137, i_13_139, i_13_175, i_13_190, i_13_226, i_13_227, i_13_374, i_13_377, i_13_460, i_13_463, i_13_490, i_13_526, i_13_527, i_13_533, i_13_535, i_13_536, i_13_617, i_13_667, i_13_715, i_13_895, i_13_946, i_13_1084, i_13_1093, i_13_1094, i_13_1313, i_13_1444, i_13_1471, i_13_1597, i_13_1621, i_13_1684, i_13_1720, i_13_1721, i_13_1724, i_13_1784, i_13_1786, i_13_1787, i_13_1838, i_13_1841, i_13_1844, i_13_1849, i_13_1931, i_13_2056, i_13_2120, i_13_2177, i_13_2197, i_13_2263, i_13_2345, i_13_2459, i_13_2501, i_13_2611, i_13_2705, i_13_2714, i_13_2872, i_13_3010, i_13_3034, i_13_3037, i_13_3044, i_13_3047, i_13_3101, i_13_3159, i_13_3161, i_13_3162, i_13_3163, i_13_3164, i_13_3275, i_13_3326, i_13_3353, i_13_3376, i_13_3407, i_13_3449, i_13_3524, i_13_3539, i_13_3653, i_13_3685, i_13_3731, i_13_3737, i_13_3740, i_13_3857, i_13_3917, i_13_3919, i_13_3982, i_13_4106, i_13_4234, i_13_4235, i_13_4258, i_13_4316, i_13_4325, i_13_4414, i_13_4415, i_13_4492, i_13_4519, i_13_4540, i_13_4541, o_13_333);
	kernel_13_334 k_13_334(i_13_41, i_13_274, i_13_283, i_13_284, i_13_383, i_13_422, i_13_454, i_13_529, i_13_553, i_13_554, i_13_558, i_13_565, i_13_599, i_13_607, i_13_666, i_13_820, i_13_821, i_13_896, i_13_1024, i_13_1099, i_13_1120, i_13_1147, i_13_1270, i_13_1314, i_13_1387, i_13_1433, i_13_1609, i_13_1635, i_13_1636, i_13_1637, i_13_1665, i_13_1687, i_13_1715, i_13_1716, i_13_1720, i_13_1732, i_13_1737, i_13_1774, i_13_1775, i_13_1788, i_13_1840, i_13_1859, i_13_1886, i_13_1960, i_13_1994, i_13_2005, i_13_2015, i_13_2121, i_13_2137, i_13_2302, i_13_2381, i_13_2459, i_13_2461, i_13_2462, i_13_2464, i_13_2493, i_13_2593, i_13_2630, i_13_2677, i_13_2678, i_13_2722, i_13_2839, i_13_2884, i_13_2983, i_13_3100, i_13_3172, i_13_3173, i_13_3175, i_13_3367, i_13_3448, i_13_3464, i_13_3545, i_13_3667, i_13_3730, i_13_3731, i_13_3733, i_13_3734, i_13_3787, i_13_3909, i_13_3910, i_13_3911, i_13_3913, i_13_3914, i_13_3931, i_13_4018, i_13_4091, i_13_4097, i_13_4162, i_13_4216, i_13_4255, i_13_4315, i_13_4351, i_13_4369, i_13_4372, i_13_4432, i_13_4514, i_13_4561, i_13_4568, i_13_4594, i_13_4603, o_13_334);
	kernel_13_335 k_13_335(i_13_77, i_13_92, i_13_203, i_13_259, i_13_265, i_13_266, i_13_353, i_13_374, i_13_382, i_13_413, i_13_451, i_13_520, i_13_569, i_13_605, i_13_607, i_13_608, i_13_658, i_13_661, i_13_670, i_13_671, i_13_680, i_13_929, i_13_940, i_13_943, i_13_950, i_13_1081, i_13_1082, i_13_1145, i_13_1148, i_13_1229, i_13_1300, i_13_1307, i_13_1385, i_13_1444, i_13_1454, i_13_1486, i_13_1663, i_13_1730, i_13_1733, i_13_1765, i_13_1766, i_13_1841, i_13_1865, i_13_1885, i_13_1892, i_13_1927, i_13_2020, i_13_2054, i_13_2137, i_13_2281, i_13_2300, i_13_2365, i_13_2423, i_13_2435, i_13_2468, i_13_2546, i_13_2570, i_13_2614, i_13_2615, i_13_2650, i_13_2858, i_13_2887, i_13_2980, i_13_3017, i_13_3047, i_13_3077, i_13_3142, i_13_3259, i_13_3269, i_13_3343, i_13_3359, i_13_3445, i_13_3449, i_13_3476, i_13_3484, i_13_3485, i_13_3646, i_13_3731, i_13_3764, i_13_3781, i_13_3872, i_13_3875, i_13_3979, i_13_4018, i_13_4054, i_13_4079, i_13_4160, i_13_4162, i_13_4163, i_13_4166, i_13_4199, i_13_4369, i_13_4370, i_13_4372, i_13_4394, i_13_4430, i_13_4441, i_13_4477, i_13_4555, i_13_4568, o_13_335);
	kernel_13_336 k_13_336(i_13_39, i_13_76, i_13_137, i_13_156, i_13_157, i_13_193, i_13_238, i_13_279, i_13_280, i_13_310, i_13_313, i_13_316, i_13_337, i_13_360, i_13_373, i_13_428, i_13_454, i_13_490, i_13_550, i_13_562, i_13_641, i_13_643, i_13_685, i_13_686, i_13_688, i_13_756, i_13_757, i_13_770, i_13_819, i_13_895, i_13_949, i_13_1057, i_13_1118, i_13_1120, i_13_1121, i_13_1122, i_13_1272, i_13_1273, i_13_1364, i_13_1371, i_13_1498, i_13_1552, i_13_1669, i_13_1722, i_13_1750, i_13_1813, i_13_1858, i_13_1884, i_13_1943, i_13_2053, i_13_2101, i_13_2153, i_13_2190, i_13_2200, i_13_2296, i_13_2548, i_13_2592, i_13_2614, i_13_2647, i_13_2650, i_13_2677, i_13_2695, i_13_2722, i_13_2767, i_13_2857, i_13_3002, i_13_3088, i_13_3127, i_13_3217, i_13_3235, i_13_3262, i_13_3303, i_13_3384, i_13_3403, i_13_3478, i_13_3847, i_13_3889, i_13_3928, i_13_3982, i_13_3990, i_13_3991, i_13_3992, i_13_4032, i_13_4033, i_13_4045, i_13_4075, i_13_4078, i_13_4081, i_13_4082, i_13_4153, i_13_4186, i_13_4187, i_13_4258, i_13_4270, i_13_4540, i_13_4560, i_13_4592, i_13_4594, i_13_4595, i_13_4600, o_13_336);
	kernel_13_337 k_13_337(i_13_102, i_13_103, i_13_276, i_13_307, i_13_448, i_13_450, i_13_460, i_13_585, i_13_586, i_13_598, i_13_610, i_13_704, i_13_828, i_13_843, i_13_844, i_13_940, i_13_1063, i_13_1081, i_13_1093, i_13_1095, i_13_1206, i_13_1305, i_13_1309, i_13_1341, i_13_1342, i_13_1380, i_13_1399, i_13_1402, i_13_1440, i_13_1441, i_13_1442, i_13_1473, i_13_1495, i_13_1529, i_13_1531, i_13_1652, i_13_1671, i_13_1698, i_13_1744, i_13_1765, i_13_1795, i_13_1810, i_13_1845, i_13_1927, i_13_1944, i_13_1990, i_13_1993, i_13_2001, i_13_2023, i_13_2197, i_13_2236, i_13_2260, i_13_2277, i_13_2278, i_13_2382, i_13_2448, i_13_2500, i_13_2547, i_13_2614, i_13_2650, i_13_2709, i_13_2718, i_13_2719, i_13_2722, i_13_2742, i_13_2766, i_13_2821, i_13_2919, i_13_2935, i_13_2949, i_13_2950, i_13_3016, i_13_3019, i_13_3061, i_13_3122, i_13_3345, i_13_3366, i_13_3367, i_13_3368, i_13_3390, i_13_3420, i_13_3454, i_13_3525, i_13_3592, i_13_3689, i_13_3730, i_13_3741, i_13_3754, i_13_3856, i_13_4051, i_13_4086, i_13_4165, i_13_4231, i_13_4257, i_13_4266, i_13_4267, i_13_4294, i_13_4302, i_13_4393, i_13_4448, o_13_337);
	kernel_13_338 k_13_338(i_13_76, i_13_118, i_13_121, i_13_158, i_13_184, i_13_186, i_13_376, i_13_508, i_13_517, i_13_526, i_13_535, i_13_557, i_13_600, i_13_616, i_13_617, i_13_661, i_13_670, i_13_737, i_13_778, i_13_850, i_13_931, i_13_945, i_13_946, i_13_1067, i_13_1069, i_13_1084, i_13_1191, i_13_1210, i_13_1276, i_13_1406, i_13_1424, i_13_1444, i_13_1545, i_13_1552, i_13_1558, i_13_1624, i_13_1631, i_13_1723, i_13_1725, i_13_1786, i_13_1814, i_13_1841, i_13_1938, i_13_1940, i_13_2120, i_13_2200, i_13_2209, i_13_2211, i_13_2212, i_13_2365, i_13_2427, i_13_2434, i_13_2459, i_13_2461, i_13_2713, i_13_2938, i_13_2939, i_13_3019, i_13_3020, i_13_3028, i_13_3029, i_13_3037, i_13_3039, i_13_3040, i_13_3044, i_13_3139, i_13_3160, i_13_3162, i_13_3163, i_13_3164, i_13_3165, i_13_3205, i_13_3209, i_13_3217, i_13_3218, i_13_3250, i_13_3289, i_13_3292, i_13_3413, i_13_3421, i_13_3424, i_13_3541, i_13_3545, i_13_3595, i_13_3874, i_13_3899, i_13_4009, i_13_4194, i_13_4233, i_13_4234, i_13_4271, i_13_4312, i_13_4333, i_13_4352, i_13_4360, i_13_4361, i_13_4414, i_13_4498, i_13_4526, i_13_4544, o_13_338);
	kernel_13_339 k_13_339(i_13_110, i_13_184, i_13_186, i_13_192, i_13_193, i_13_194, i_13_195, i_13_328, i_13_333, i_13_572, i_13_573, i_13_618, i_13_625, i_13_641, i_13_658, i_13_715, i_13_716, i_13_858, i_13_859, i_13_867, i_13_868, i_13_928, i_13_955, i_13_1116, i_13_1117, i_13_1148, i_13_1149, i_13_1210, i_13_1225, i_13_1226, i_13_1228, i_13_1229, i_13_1256, i_13_1258, i_13_1259, i_13_1329, i_13_1404, i_13_1405, i_13_1408, i_13_1411, i_13_1507, i_13_1513, i_13_1570, i_13_1597, i_13_1678, i_13_1680, i_13_1729, i_13_1734, i_13_1765, i_13_1768, i_13_1801, i_13_1802, i_13_1829, i_13_1956, i_13_1991, i_13_2002, i_13_2056, i_13_2059, i_13_2225, i_13_2281, i_13_2302, i_13_2341, i_13_2532, i_13_2614, i_13_2619, i_13_2648, i_13_2705, i_13_2746, i_13_2857, i_13_2981, i_13_3034, i_13_3064, i_13_3118, i_13_3145, i_13_3214, i_13_3258, i_13_3268, i_13_3269, i_13_3287, i_13_3291, i_13_3310, i_13_3386, i_13_3421, i_13_3424, i_13_3546, i_13_3562, i_13_3606, i_13_3755, i_13_3763, i_13_3764, i_13_3979, i_13_4018, i_13_4078, i_13_4201, i_13_4202, i_13_4213, i_13_4267, i_13_4297, i_13_4362, i_13_4515, o_13_339);
	kernel_13_340 k_13_340(i_13_45, i_13_46, i_13_55, i_13_103, i_13_138, i_13_154, i_13_186, i_13_255, i_13_258, i_13_259, i_13_307, i_13_309, i_13_352, i_13_408, i_13_450, i_13_505, i_13_644, i_13_660, i_13_667, i_13_848, i_13_894, i_13_930, i_13_936, i_13_937, i_13_1108, i_13_1227, i_13_1228, i_13_1243, i_13_1326, i_13_1328, i_13_1399, i_13_1479, i_13_1513, i_13_1623, i_13_1660, i_13_1677, i_13_1723, i_13_1764, i_13_1767, i_13_1801, i_13_1803, i_13_1804, i_13_1944, i_13_1945, i_13_1948, i_13_2025, i_13_2026, i_13_2053, i_13_2134, i_13_2145, i_13_2197, i_13_2206, i_13_2277, i_13_2297, i_13_2403, i_13_2404, i_13_2430, i_13_2471, i_13_2578, i_13_2611, i_13_2613, i_13_2622, i_13_2745, i_13_2793, i_13_2848, i_13_2916, i_13_2980, i_13_3001, i_13_3027, i_13_3028, i_13_3073, i_13_3133, i_13_3213, i_13_3352, i_13_3367, i_13_3378, i_13_3439, i_13_3591, i_13_3592, i_13_3703, i_13_3763, i_13_3780, i_13_3820, i_13_3898, i_13_3978, i_13_3979, i_13_4017, i_13_4158, i_13_4231, i_13_4249, i_13_4302, i_13_4332, i_13_4351, i_13_4360, i_13_4367, i_13_4387, i_13_4438, i_13_4446, i_13_4563, i_13_4602, o_13_340);
	kernel_13_341 k_13_341(i_13_97, i_13_107, i_13_119, i_13_121, i_13_122, i_13_181, i_13_285, i_13_286, i_13_311, i_13_320, i_13_430, i_13_535, i_13_538, i_13_569, i_13_599, i_13_697, i_13_712, i_13_746, i_13_781, i_13_850, i_13_934, i_13_976, i_13_985, i_13_1034, i_13_1093, i_13_1094, i_13_1216, i_13_1279, i_13_1283, i_13_1284, i_13_1300, i_13_1471, i_13_1526, i_13_1552, i_13_1714, i_13_1721, i_13_1726, i_13_1757, i_13_1760, i_13_1783, i_13_1786, i_13_1787, i_13_1789, i_13_1817, i_13_2072, i_13_2120, i_13_2123, i_13_2209, i_13_2308, i_13_2312, i_13_2365, i_13_2458, i_13_2459, i_13_2465, i_13_2551, i_13_2630, i_13_2633, i_13_2663, i_13_2939, i_13_3040, i_13_3148, i_13_3161, i_13_3163, i_13_3167, i_13_3211, i_13_3212, i_13_3218, i_13_3265, i_13_3271, i_13_3347, i_13_3424, i_13_3482, i_13_3483, i_13_3506, i_13_3523, i_13_3527, i_13_3688, i_13_3689, i_13_3700, i_13_3746, i_13_3844, i_13_3871, i_13_3878, i_13_3935, i_13_3962, i_13_4009, i_13_4012, i_13_4048, i_13_4093, i_13_4105, i_13_4106, i_13_4235, i_13_4237, i_13_4238, i_13_4261, i_13_4273, i_13_4414, i_13_4417, i_13_4450, i_13_4519, o_13_341);
	kernel_13_342 k_13_342(i_13_31, i_13_93, i_13_94, i_13_97, i_13_114, i_13_121, i_13_123, i_13_159, i_13_184, i_13_328, i_13_435, i_13_517, i_13_564, i_13_570, i_13_571, i_13_574, i_13_614, i_13_696, i_13_697, i_13_732, i_13_733, i_13_742, i_13_796, i_13_799, i_13_822, i_13_1210, i_13_1254, i_13_1390, i_13_1408, i_13_1446, i_13_1447, i_13_1456, i_13_1473, i_13_1489, i_13_1551, i_13_1552, i_13_1569, i_13_1642, i_13_1761, i_13_1786, i_13_1789, i_13_1860, i_13_1910, i_13_2018, i_13_2056, i_13_2103, i_13_2175, i_13_2176, i_13_2202, i_13_2208, i_13_2235, i_13_2238, i_13_2269, i_13_2427, i_13_2434, i_13_2541, i_13_2680, i_13_2767, i_13_2914, i_13_2985, i_13_3009, i_13_3022, i_13_3028, i_13_3053, i_13_3091, i_13_3163, i_13_3207, i_13_3243, i_13_3244, i_13_3415, i_13_3422, i_13_3423, i_13_3424, i_13_3426, i_13_3427, i_13_3432, i_13_3451, i_13_3521, i_13_3571, i_13_3649, i_13_3665, i_13_3702, i_13_3739, i_13_3846, i_13_3847, i_13_3850, i_13_3873, i_13_3874, i_13_3876, i_13_3967, i_13_4009, i_13_4038, i_13_4119, i_13_4188, i_13_4189, i_13_4195, i_13_4236, i_13_4351, i_13_4353, i_13_4569, o_13_342);
	kernel_13_343 k_13_343(i_13_39, i_13_48, i_13_139, i_13_163, i_13_174, i_13_274, i_13_279, i_13_280, i_13_307, i_13_310, i_13_315, i_13_316, i_13_514, i_13_549, i_13_550, i_13_639, i_13_640, i_13_646, i_13_667, i_13_670, i_13_675, i_13_676, i_13_684, i_13_685, i_13_687, i_13_688, i_13_691, i_13_757, i_13_875, i_13_981, i_13_1055, i_13_1099, i_13_1116, i_13_1270, i_13_1363, i_13_1438, i_13_1445, i_13_1449, i_13_1593, i_13_1594, i_13_1597, i_13_1632, i_13_1803, i_13_1813, i_13_1847, i_13_2053, i_13_2236, i_13_2274, i_13_2313, i_13_2396, i_13_2397, i_13_2422, i_13_2507, i_13_2614, i_13_2648, i_13_2649, i_13_2650, i_13_2673, i_13_2674, i_13_2693, i_13_2694, i_13_2695, i_13_2698, i_13_2929, i_13_3011, i_13_3034, i_13_3142, i_13_3145, i_13_3217, i_13_3385, i_13_3415, i_13_3532, i_13_3610, i_13_3685, i_13_3730, i_13_3736, i_13_3739, i_13_3816, i_13_3817, i_13_3888, i_13_3889, i_13_3987, i_13_3991, i_13_4017, i_13_4032, i_13_4033, i_13_4034, i_13_4077, i_13_4086, i_13_4187, i_13_4278, i_13_4306, i_13_4338, i_13_4458, i_13_4531, i_13_4540, i_13_4590, i_13_4591, i_13_4594, i_13_4600, o_13_343);
	kernel_13_344 k_13_344(i_13_112, i_13_121, i_13_122, i_13_139, i_13_193, i_13_230, i_13_267, i_13_274, i_13_275, i_13_320, i_13_382, i_13_409, i_13_410, i_13_418, i_13_454, i_13_466, i_13_528, i_13_562, i_13_589, i_13_590, i_13_591, i_13_597, i_13_625, i_13_646, i_13_688, i_13_718, i_13_760, i_13_761, i_13_824, i_13_839, i_13_843, i_13_915, i_13_949, i_13_1208, i_13_1211, i_13_1274, i_13_1307, i_13_1310, i_13_1348, i_13_1391, i_13_1531, i_13_1597, i_13_1598, i_13_1624, i_13_1640, i_13_1643, i_13_1646, i_13_1670, i_13_1886, i_13_1938, i_13_2138, i_13_2140, i_13_2192, i_13_2209, i_13_2248, i_13_2363, i_13_2434, i_13_2542, i_13_2550, i_13_2551, i_13_2552, i_13_2623, i_13_2651, i_13_2678, i_13_2821, i_13_2822, i_13_2857, i_13_2998, i_13_3108, i_13_3109, i_13_3110, i_13_3116, i_13_3163, i_13_3235, i_13_3269, i_13_3323, i_13_3361, i_13_3370, i_13_3388, i_13_3389, i_13_3391, i_13_3491, i_13_3595, i_13_3633, i_13_3668, i_13_3685, i_13_3767, i_13_3882, i_13_4036, i_13_4037, i_13_4055, i_13_4162, i_13_4262, i_13_4351, i_13_4372, i_13_4397, i_13_4451, i_13_4559, i_13_4567, i_13_4596, o_13_344);
	kernel_13_345 k_13_345(i_13_48, i_13_61, i_13_93, i_13_106, i_13_136, i_13_259, i_13_492, i_13_619, i_13_624, i_13_625, i_13_627, i_13_673, i_13_697, i_13_707, i_13_823, i_13_825, i_13_826, i_13_948, i_13_978, i_13_979, i_13_1024, i_13_1072, i_13_1095, i_13_1102, i_13_1200, i_13_1279, i_13_1303, i_13_1320, i_13_1321, i_13_1428, i_13_1434, i_13_1444, i_13_1464, i_13_1465, i_13_1480, i_13_1483, i_13_1547, i_13_1572, i_13_1752, i_13_1757, i_13_1786, i_13_1807, i_13_1911, i_13_1960, i_13_2010, i_13_2103, i_13_2238, i_13_2244, i_13_2245, i_13_2263, i_13_2343, i_13_2424, i_13_2442, i_13_2443, i_13_2445, i_13_2446, i_13_2454, i_13_2554, i_13_2743, i_13_2752, i_13_2823, i_13_2824, i_13_2857, i_13_2883, i_13_3073, i_13_3135, i_13_3153, i_13_3310, i_13_3345, i_13_3381, i_13_3418, i_13_3432, i_13_3437, i_13_3475, i_13_3489, i_13_3594, i_13_3618, i_13_3622, i_13_3766, i_13_3786, i_13_3874, i_13_3936, i_13_3937, i_13_4018, i_13_4209, i_13_4210, i_13_4237, i_13_4330, i_13_4332, i_13_4333, i_13_4341, i_13_4344, i_13_4351, i_13_4381, i_13_4396, i_13_4452, i_13_4453, i_13_4509, i_13_4567, i_13_4587, o_13_345);
	kernel_13_346 k_13_346(i_13_40, i_13_117, i_13_121, i_13_162, i_13_166, i_13_183, i_13_189, i_13_192, i_13_283, i_13_315, i_13_333, i_13_454, i_13_517, i_13_532, i_13_576, i_13_661, i_13_714, i_13_760, i_13_862, i_13_927, i_13_948, i_13_1098, i_13_1135, i_13_1227, i_13_1254, i_13_1259, i_13_1261, i_13_1279, i_13_1407, i_13_1430, i_13_1458, i_13_1468, i_13_1479, i_13_1488, i_13_1507, i_13_1522, i_13_1570, i_13_1597, i_13_1624, i_13_1647, i_13_1685, i_13_1710, i_13_1723, i_13_1767, i_13_1771, i_13_1782, i_13_1786, i_13_1800, i_13_1939, i_13_2011, i_13_2056, i_13_2100, i_13_2115, i_13_2208, i_13_2209, i_13_2223, i_13_2224, i_13_2235, i_13_2236, i_13_2358, i_13_2394, i_13_2407, i_13_2438, i_13_2457, i_13_2532, i_13_2565, i_13_2595, i_13_2835, i_13_2902, i_13_3036, i_13_3136, i_13_3216, i_13_3217, i_13_3221, i_13_3286, i_13_3339, i_13_3369, i_13_3414, i_13_3424, i_13_3429, i_13_3468, i_13_3549, i_13_3613, i_13_3699, i_13_3855, i_13_3873, i_13_3877, i_13_3883, i_13_3982, i_13_4008, i_13_4009, i_13_4260, i_13_4261, i_13_4297, i_13_4360, i_13_4518, i_13_4527, i_13_4530, i_13_4540, i_13_4594, o_13_346);
	kernel_13_347 k_13_347(i_13_161, i_13_232, i_13_242, i_13_285, i_13_359, i_13_412, i_13_469, i_13_503, i_13_526, i_13_528, i_13_529, i_13_535, i_13_706, i_13_843, i_13_853, i_13_882, i_13_895, i_13_897, i_13_1024, i_13_1203, i_13_1309, i_13_1310, i_13_1312, i_13_1390, i_13_1426, i_13_1428, i_13_1438, i_13_1496, i_13_1500, i_13_1501, i_13_1550, i_13_1552, i_13_1574, i_13_1631, i_13_1723, i_13_1726, i_13_1786, i_13_1834, i_13_1917, i_13_1950, i_13_2004, i_13_2033, i_13_2114, i_13_2200, i_13_2201, i_13_2202, i_13_2263, i_13_2407, i_13_2449, i_13_2452, i_13_2454, i_13_2455, i_13_2721, i_13_2764, i_13_2767, i_13_2924, i_13_3012, i_13_3163, i_13_3217, i_13_3323, i_13_3373, i_13_3460, i_13_3464, i_13_3533, i_13_3539, i_13_3545, i_13_3579, i_13_3581, i_13_3597, i_13_3623, i_13_3635, i_13_3646, i_13_3666, i_13_3669, i_13_3730, i_13_3731, i_13_3733, i_13_3734, i_13_3786, i_13_3787, i_13_3856, i_13_3865, i_13_3892, i_13_3931, i_13_4016, i_13_4081, i_13_4234, i_13_4252, i_13_4253, i_13_4261, i_13_4263, i_13_4264, i_13_4279, i_13_4369, i_13_4380, i_13_4435, i_13_4452, i_13_4554, i_13_4555, i_13_4558, o_13_347);
	kernel_13_348 k_13_348(i_13_49, i_13_76, i_13_77, i_13_100, i_13_329, i_13_353, i_13_356, i_13_409, i_13_410, i_13_419, i_13_529, i_13_530, i_13_562, i_13_611, i_13_698, i_13_742, i_13_827, i_13_853, i_13_854, i_13_953, i_13_1025, i_13_1076, i_13_1109, i_13_1142, i_13_1232, i_13_1305, i_13_1309, i_13_1310, i_13_1313, i_13_1321, i_13_1322, i_13_1330, i_13_1430, i_13_1444, i_13_1462, i_13_1493, i_13_1552, i_13_1553, i_13_1694, i_13_1723, i_13_1741, i_13_1771, i_13_1777, i_13_1846, i_13_1889, i_13_1948, i_13_1951, i_13_1961, i_13_2011, i_13_2033, i_13_2141, i_13_2203, i_13_2236, i_13_2237, i_13_2282, i_13_2354, i_13_2402, i_13_2428, i_13_2546, i_13_2596, i_13_2654, i_13_2923, i_13_2924, i_13_3013, i_13_3014, i_13_3016, i_13_3034, i_13_3071, i_13_3197, i_13_3274, i_13_3419, i_13_3427, i_13_3442, i_13_3542, i_13_3544, i_13_3580, i_13_3595, i_13_3726, i_13_3730, i_13_3734, i_13_3787, i_13_3788, i_13_3806, i_13_3896, i_13_3913, i_13_3914, i_13_3929, i_13_3938, i_13_4060, i_13_4238, i_13_4256, i_13_4264, i_13_4265, i_13_4334, i_13_4381, i_13_4382, i_13_4450, i_13_4454, i_13_4478, i_13_4600, o_13_348);
	kernel_13_349 k_13_349(i_13_205, i_13_210, i_13_285, i_13_363, i_13_417, i_13_465, i_13_520, i_13_525, i_13_528, i_13_529, i_13_537, i_13_690, i_13_736, i_13_825, i_13_852, i_13_853, i_13_1020, i_13_1023, i_13_1024, i_13_1075, i_13_1120, i_13_1131, i_13_1212, i_13_1311, i_13_1312, i_13_1317, i_13_1320, i_13_1461, i_13_1498, i_13_1551, i_13_1552, i_13_1554, i_13_1555, i_13_1605, i_13_1699, i_13_1749, i_13_1906, i_13_1920, i_13_1932, i_13_1941, i_13_1959, i_13_1960, i_13_2032, i_13_2127, i_13_2136, i_13_2139, i_13_2199, i_13_2202, i_13_2454, i_13_2491, i_13_2506, i_13_2572, i_13_2677, i_13_3012, i_13_3013, i_13_3103, i_13_3118, i_13_3156, i_13_3172, i_13_3271, i_13_3378, i_13_3432, i_13_3453, i_13_3460, i_13_3478, i_13_3505, i_13_3540, i_13_3541, i_13_3543, i_13_3571, i_13_3579, i_13_3580, i_13_3597, i_13_3633, i_13_3669, i_13_3670, i_13_3729, i_13_3732, i_13_3733, i_13_3786, i_13_3787, i_13_3805, i_13_3858, i_13_3912, i_13_3918, i_13_3919, i_13_3985, i_13_4039, i_13_4120, i_13_4164, i_13_4254, i_13_4255, i_13_4260, i_13_4341, i_13_4351, i_13_4354, i_13_4378, i_13_4380, i_13_4381, i_13_4578, o_13_349);
	kernel_13_350 k_13_350(i_13_31, i_13_46, i_13_47, i_13_163, i_13_164, i_13_173, i_13_174, i_13_245, i_13_273, i_13_299, i_13_326, i_13_415, i_13_416, i_13_518, i_13_533, i_13_568, i_13_626, i_13_658, i_13_659, i_13_688, i_13_721, i_13_757, i_13_758, i_13_761, i_13_848, i_13_856, i_13_937, i_13_938, i_13_1023, i_13_1072, i_13_1073, i_13_1129, i_13_1130, i_13_1201, i_13_1219, i_13_1252, i_13_1253, i_13_1280, i_13_1445, i_13_1495, i_13_1522, i_13_1523, i_13_1535, i_13_1549, i_13_1550, i_13_1603, i_13_1604, i_13_1725, i_13_1751, i_13_1946, i_13_1991, i_13_2026, i_13_2027, i_13_2116, i_13_2297, i_13_2425, i_13_2443, i_13_2471, i_13_2472, i_13_2539, i_13_2540, i_13_2722, i_13_2724, i_13_2801, i_13_2920, i_13_2981, i_13_3000, i_13_3001, i_13_3003, i_13_3007, i_13_3029, i_13_3124, i_13_3215, i_13_3218, i_13_3262, i_13_3457, i_13_3458, i_13_3485, i_13_3538, i_13_3539, i_13_3547, i_13_3575, i_13_3638, i_13_3818, i_13_3822, i_13_3844, i_13_3894, i_13_3898, i_13_3899, i_13_3908, i_13_4018, i_13_4053, i_13_4061, i_13_4102, i_13_4322, i_13_4331, i_13_4339, i_13_4511, i_13_4604, i_13_4605, o_13_350);
	kernel_13_351 k_13_351(i_13_33, i_13_46, i_13_160, i_13_167, i_13_175, i_13_200, i_13_238, i_13_248, i_13_274, i_13_275, i_13_277, i_13_278, i_13_283, i_13_284, i_13_315, i_13_340, i_13_376, i_13_454, i_13_457, i_13_492, i_13_494, i_13_521, i_13_565, i_13_566, i_13_575, i_13_584, i_13_615, i_13_644, i_13_688, i_13_713, i_13_741, i_13_742, i_13_745, i_13_823, i_13_824, i_13_960, i_13_1092, i_13_1201, i_13_1221, i_13_1349, i_13_1400, i_13_1494, i_13_1499, i_13_1715, i_13_1722, i_13_1770, i_13_1817, i_13_1858, i_13_1861, i_13_1890, i_13_1920, i_13_2147, i_13_2300, i_13_2524, i_13_2540, i_13_2651, i_13_2676, i_13_2721, i_13_2723, i_13_2725, i_13_2726, i_13_2771, i_13_2785, i_13_3036, i_13_3076, i_13_3214, i_13_3216, i_13_3218, i_13_3234, i_13_3235, i_13_3366, i_13_3423, i_13_3426, i_13_3432, i_13_3461, i_13_3477, i_13_3549, i_13_3639, i_13_3689, i_13_3723, i_13_3730, i_13_3858, i_13_3892, i_13_3897, i_13_3901, i_13_3904, i_13_3923, i_13_3981, i_13_3986, i_13_4011, i_13_4089, i_13_4163, i_13_4218, i_13_4261, i_13_4273, i_13_4363, i_13_4472, i_13_4512, i_13_4569, i_13_4598, o_13_351);
	kernel_13_352 k_13_352(i_13_74, i_13_77, i_13_137, i_13_170, i_13_265, i_13_266, i_13_283, i_13_319, i_13_337, i_13_492, i_13_518, i_13_571, i_13_582, i_13_662, i_13_688, i_13_697, i_13_814, i_13_886, i_13_888, i_13_935, i_13_939, i_13_1066, i_13_1112, i_13_1145, i_13_1148, i_13_1208, i_13_1210, i_13_1217, i_13_1226, i_13_1253, i_13_1266, i_13_1426, i_13_1530, i_13_1633, i_13_1660, i_13_1662, i_13_1730, i_13_1731, i_13_1733, i_13_1734, i_13_1849, i_13_1886, i_13_2020, i_13_2021, i_13_2031, i_13_2117, i_13_2137, i_13_2209, i_13_2263, i_13_2297, i_13_2407, i_13_2408, i_13_2432, i_13_2445, i_13_2498, i_13_2501, i_13_2517, i_13_2725, i_13_2812, i_13_2884, i_13_2938, i_13_3047, i_13_3076, i_13_3089, i_13_3115, i_13_3208, i_13_3209, i_13_3424, i_13_3476, i_13_3505, i_13_3565, i_13_3569, i_13_3597, i_13_3611, i_13_3614, i_13_3730, i_13_3739, i_13_3740, i_13_3741, i_13_3747, i_13_4036, i_13_4063, i_13_4064, i_13_4160, i_13_4163, i_13_4164, i_13_4202, i_13_4316, i_13_4327, i_13_4330, i_13_4331, i_13_4340, i_13_4367, i_13_4369, i_13_4370, i_13_4372, i_13_4517, i_13_4600, i_13_4604, i_13_4606, o_13_352);
	kernel_13_353 k_13_353(i_13_52, i_13_111, i_13_124, i_13_140, i_13_169, i_13_170, i_13_269, i_13_273, i_13_283, i_13_287, i_13_371, i_13_373, i_13_417, i_13_463, i_13_509, i_13_692, i_13_817, i_13_818, i_13_849, i_13_851, i_13_853, i_13_886, i_13_887, i_13_916, i_13_939, i_13_943, i_13_985, i_13_1053, i_13_1067, i_13_1110, i_13_1121, i_13_1122, i_13_1328, i_13_1329, i_13_1492, i_13_1573, i_13_1623, i_13_1808, i_13_1830, i_13_1840, i_13_1852, i_13_1853, i_13_1857, i_13_1924, i_13_2006, i_13_2051, i_13_2123, i_13_2136, i_13_2140, i_13_2141, i_13_2173, i_13_2237, i_13_2407, i_13_2408, i_13_2410, i_13_2411, i_13_2460, i_13_2552, i_13_2696, i_13_2823, i_13_2848, i_13_2875, i_13_2941, i_13_2942, i_13_3011, i_13_3031, i_13_3037, i_13_3050, i_13_3108, i_13_3346, i_13_3400, i_13_3424, i_13_3453, i_13_3478, i_13_3479, i_13_3505, i_13_3525, i_13_3526, i_13_3567, i_13_3741, i_13_3742, i_13_3765, i_13_3821, i_13_3867, i_13_3911, i_13_3928, i_13_3984, i_13_4022, i_13_4063, i_13_4064, i_13_4066, i_13_4067, i_13_4164, i_13_4209, i_13_4309, i_13_4318, i_13_4319, i_13_4434, i_13_4441, i_13_4451, o_13_353);
	kernel_13_354 k_13_354(i_13_73, i_13_74, i_13_123, i_13_186, i_13_235, i_13_280, i_13_284, i_13_442, i_13_523, i_13_532, i_13_533, i_13_640, i_13_668, i_13_676, i_13_677, i_13_680, i_13_717, i_13_832, i_13_839, i_13_958, i_13_982, i_13_1084, i_13_1099, i_13_1145, i_13_1256, i_13_1270, i_13_1271, i_13_1302, i_13_1400, i_13_1464, i_13_1504, i_13_1505, i_13_1594, i_13_1658, i_13_1720, i_13_1723, i_13_1744, i_13_1775, i_13_1792, i_13_1796, i_13_1881, i_13_1915, i_13_1989, i_13_2017, i_13_2026, i_13_2116, i_13_2223, i_13_2446, i_13_2511, i_13_2512, i_13_2539, i_13_2575, i_13_2576, i_13_2611, i_13_2750, i_13_2844, i_13_2845, i_13_2854, i_13_2921, i_13_2922, i_13_2935, i_13_3001, i_13_3135, i_13_3259, i_13_3260, i_13_3287, i_13_3289, i_13_3321, i_13_3350, i_13_3371, i_13_3396, i_13_3449, i_13_3452, i_13_3477, i_13_3578, i_13_3593, i_13_3647, i_13_3784, i_13_3865, i_13_3889, i_13_3907, i_13_3924, i_13_3925, i_13_3926, i_13_3984, i_13_3988, i_13_3989, i_13_4078, i_13_4079, i_13_4099, i_13_4106, i_13_4163, i_13_4186, i_13_4187, i_13_4331, i_13_4340, i_13_4430, i_13_4452, i_13_4543, i_13_4592, o_13_354);
	kernel_13_355 k_13_355(i_13_45, i_13_172, i_13_175, i_13_178, i_13_179, i_13_229, i_13_280, i_13_283, i_13_284, i_13_286, i_13_287, i_13_335, i_13_360, i_13_454, i_13_562, i_13_574, i_13_589, i_13_645, i_13_687, i_13_688, i_13_691, i_13_742, i_13_760, i_13_823, i_13_832, i_13_867, i_13_871, i_13_872, i_13_1078, i_13_1085, i_13_1122, i_13_1228, i_13_1229, i_13_1469, i_13_1573, i_13_1636, i_13_1710, i_13_1712, i_13_1716, i_13_1732, i_13_1747, i_13_1750, i_13_1751, i_13_1855, i_13_1858, i_13_1859, i_13_1861, i_13_1864, i_13_1933, i_13_2239, i_13_2341, i_13_2428, i_13_2624, i_13_2652, i_13_2653, i_13_2654, i_13_2708, i_13_2722, i_13_2731, i_13_2752, i_13_2785, i_13_2851, i_13_3092, i_13_3100, i_13_3113, i_13_3172, i_13_3174, i_13_3235, i_13_3267, i_13_3268, i_13_3271, i_13_3274, i_13_3293, i_13_3371, i_13_3400, i_13_3424, i_13_3426, i_13_3427, i_13_3428, i_13_3646, i_13_3686, i_13_3783, i_13_3890, i_13_3910, i_13_3911, i_13_3913, i_13_3914, i_13_3995, i_13_4017, i_13_4018, i_13_4019, i_13_4021, i_13_4090, i_13_4097, i_13_4295, i_13_4322, i_13_4556, i_13_4559, i_13_4561, i_13_4573, o_13_355);
	kernel_13_356 k_13_356(i_13_44, i_13_79, i_13_80, i_13_168, i_13_276, i_13_537, i_13_539, i_13_554, i_13_591, i_13_608, i_13_611, i_13_645, i_13_647, i_13_672, i_13_673, i_13_674, i_13_682, i_13_683, i_13_691, i_13_692, i_13_701, i_13_718, i_13_823, i_13_844, i_13_978, i_13_1065, i_13_1104, i_13_1123, i_13_1124, i_13_1218, i_13_1223, i_13_1283, i_13_1410, i_13_1423, i_13_1426, i_13_1429, i_13_1470, i_13_1659, i_13_1660, i_13_1663, i_13_1689, i_13_1727, i_13_1734, i_13_1736, i_13_1799, i_13_1803, i_13_1842, i_13_1849, i_13_1992, i_13_2022, i_13_2024, i_13_2058, i_13_2104, i_13_2450, i_13_2496, i_13_2570, i_13_2698, i_13_2715, i_13_2887, i_13_2938, i_13_2982, i_13_3027, i_13_3067, i_13_3068, i_13_3088, i_13_3089, i_13_3102, i_13_3104, i_13_3244, i_13_3289, i_13_3454, i_13_3525, i_13_3572, i_13_3653, i_13_3682, i_13_3739, i_13_3742, i_13_3743, i_13_3787, i_13_3797, i_13_3858, i_13_3930, i_13_3931, i_13_3932, i_13_3994, i_13_3995, i_13_4063, i_13_4084, i_13_4189, i_13_4190, i_13_4191, i_13_4193, i_13_4249, i_13_4368, i_13_4515, i_13_4533, i_13_4595, i_13_4596, i_13_4597, i_13_4598, o_13_356);
	kernel_13_357 k_13_357(i_13_27, i_13_28, i_13_35, i_13_37, i_13_54, i_13_63, i_13_64, i_13_80, i_13_135, i_13_172, i_13_178, i_13_306, i_13_307, i_13_316, i_13_325, i_13_379, i_13_383, i_13_588, i_13_612, i_13_639, i_13_642, i_13_647, i_13_694, i_13_772, i_13_944, i_13_1121, i_13_1131, i_13_1198, i_13_1206, i_13_1227, i_13_1269, i_13_1270, i_13_1272, i_13_1305, i_13_1309, i_13_1342, i_13_1351, i_13_1390, i_13_1396, i_13_1489, i_13_1504, i_13_1593, i_13_1594, i_13_1638, i_13_1639, i_13_1792, i_13_1828, i_13_1881, i_13_1882, i_13_1909, i_13_1918, i_13_1926, i_13_1927, i_13_1931, i_13_2008, i_13_2011, i_13_2126, i_13_2537, i_13_2596, i_13_2673, i_13_2674, i_13_2719, i_13_2848, i_13_2849, i_13_2875, i_13_2880, i_13_2881, i_13_2934, i_13_3040, i_13_3060, i_13_3061, i_13_3204, i_13_3208, i_13_3218, i_13_3241, i_13_3387, i_13_3397, i_13_3505, i_13_3636, i_13_3738, i_13_3853, i_13_3916, i_13_3925, i_13_3932, i_13_3934, i_13_3973, i_13_4033, i_13_4064, i_13_4091, i_13_4185, i_13_4213, i_13_4215, i_13_4260, i_13_4294, i_13_4302, i_13_4308, i_13_4315, i_13_4393, i_13_4396, i_13_4593, o_13_357);
	kernel_13_358 k_13_358(i_13_67, i_13_105, i_13_106, i_13_165, i_13_241, i_13_258, i_13_339, i_13_527, i_13_662, i_13_697, i_13_771, i_13_793, i_13_817, i_13_831, i_13_832, i_13_851, i_13_855, i_13_856, i_13_897, i_13_1068, i_13_1069, i_13_1076, i_13_1099, i_13_1279, i_13_1309, i_13_1464, i_13_1470, i_13_1485, i_13_1497, i_13_1572, i_13_1573, i_13_1597, i_13_1642, i_13_1679, i_13_1735, i_13_1788, i_13_1852, i_13_1914, i_13_1935, i_13_1996, i_13_2120, i_13_2122, i_13_2123, i_13_2139, i_13_2140, i_13_2184, i_13_2209, i_13_2280, i_13_2409, i_13_2453, i_13_2460, i_13_2461, i_13_2464, i_13_2536, i_13_2640, i_13_2722, i_13_2751, i_13_2757, i_13_2760, i_13_2940, i_13_2941, i_13_2942, i_13_2982, i_13_3014, i_13_3030, i_13_3031, i_13_3040, i_13_3106, i_13_3148, i_13_3244, i_13_3291, i_13_3292, i_13_3322, i_13_3346, i_13_3399, i_13_3400, i_13_3402, i_13_3417, i_13_3418, i_13_3423, i_13_3525, i_13_3526, i_13_3732, i_13_3785, i_13_3866, i_13_3909, i_13_3911, i_13_4047, i_13_4056, i_13_4066, i_13_4120, i_13_4216, i_13_4317, i_13_4318, i_13_4357, i_13_4366, i_13_4391, i_13_4524, i_13_4559, i_13_4562, o_13_358);
	kernel_13_359 k_13_359(i_13_40, i_13_48, i_13_64, i_13_72, i_13_139, i_13_163, i_13_174, i_13_237, i_13_241, i_13_273, i_13_274, i_13_336, i_13_378, i_13_379, i_13_450, i_13_453, i_13_513, i_13_558, i_13_559, i_13_561, i_13_586, i_13_817, i_13_840, i_13_849, i_13_850, i_13_889, i_13_927, i_13_928, i_13_1078, i_13_1080, i_13_1081, i_13_1200, i_13_1261, i_13_1327, i_13_1359, i_13_1371, i_13_1396, i_13_1494, i_13_1620, i_13_1623, i_13_1657, i_13_1731, i_13_1732, i_13_1750, i_13_1785, i_13_1809, i_13_1810, i_13_1917, i_13_1935, i_13_1936, i_13_2055, i_13_2091, i_13_2229, i_13_2388, i_13_2430, i_13_2506, i_13_2512, i_13_2560, i_13_2565, i_13_2650, i_13_2709, i_13_2938, i_13_2955, i_13_3016, i_13_3043, i_13_3060, i_13_3096, i_13_3097, i_13_3141, i_13_3150, i_13_3162, i_13_3204, i_13_3205, i_13_3213, i_13_3216, i_13_3217, i_13_3231, i_13_3234, i_13_3312, i_13_3519, i_13_3549, i_13_3600, i_13_3681, i_13_3684, i_13_3720, i_13_3853, i_13_3873, i_13_3900, i_13_4087, i_13_4159, i_13_4162, i_13_4170, i_13_4207, i_13_4339, i_13_4359, i_13_4410, i_13_4530, i_13_4554, i_13_4594, i_13_4603, o_13_359);
	kernel_13_360 k_13_360(i_13_66, i_13_108, i_13_121, i_13_124, i_13_125, i_13_140, i_13_229, i_13_230, i_13_232, i_13_268, i_13_282, i_13_341, i_13_353, i_13_381, i_13_387, i_13_418, i_13_449, i_13_517, i_13_532, i_13_535, i_13_538, i_13_539, i_13_575, i_13_637, i_13_729, i_13_734, i_13_792, i_13_855, i_13_949, i_13_985, i_13_1049, i_13_1215, i_13_1301, i_13_1318, i_13_1367, i_13_1376, i_13_1394, i_13_1448, i_13_1465, i_13_1485, i_13_1512, i_13_1723, i_13_1724, i_13_1783, i_13_1786, i_13_1787, i_13_1789, i_13_1790, i_13_1827, i_13_1840, i_13_1841, i_13_1843, i_13_1844, i_13_2128, i_13_2169, i_13_2224, i_13_2240, i_13_2429, i_13_2430, i_13_2435, i_13_2849, i_13_2861, i_13_2873, i_13_3023, i_13_3038, i_13_3047, i_13_3159, i_13_3166, i_13_3167, i_13_3220, i_13_3236, i_13_3266, i_13_3410, i_13_3420, i_13_3425, i_13_3428, i_13_3431, i_13_3487, i_13_3541, i_13_3616, i_13_3725, i_13_3794, i_13_3839, i_13_3878, i_13_3906, i_13_3978, i_13_3985, i_13_4005, i_13_4009, i_13_4011, i_13_4012, i_13_4013, i_13_4185, i_13_4237, i_13_4238, i_13_4328, i_13_4370, i_13_4418, i_13_4498, i_13_4536, o_13_360);
	kernel_13_361 k_13_361(i_13_49, i_13_50, i_13_52, i_13_71, i_13_94, i_13_97, i_13_98, i_13_248, i_13_251, i_13_259, i_13_278, i_13_310, i_13_319, i_13_364, i_13_521, i_13_575, i_13_619, i_13_620, i_13_700, i_13_800, i_13_889, i_13_979, i_13_980, i_13_1025, i_13_1079, i_13_1087, i_13_1265, i_13_1331, i_13_1403, i_13_1427, i_13_1429, i_13_1430, i_13_1435, i_13_1436, i_13_1573, i_13_1637, i_13_1652, i_13_1661, i_13_1664, i_13_1735, i_13_1736, i_13_1777, i_13_1808, i_13_1817, i_13_1921, i_13_1933, i_13_2023, i_13_2024, i_13_2030, i_13_2051, i_13_2059, i_13_2230, i_13_2344, i_13_2455, i_13_2456, i_13_2588, i_13_2716, i_13_2726, i_13_2743, i_13_2744, i_13_2788, i_13_2789, i_13_2959, i_13_3002, i_13_3032, i_13_3058, i_13_3076, i_13_3077, i_13_3119, i_13_3128, i_13_3272, i_13_3292, i_13_3316, i_13_3370, i_13_3380, i_13_3419, i_13_3452, i_13_3454, i_13_3464, i_13_3472, i_13_3481, i_13_3514, i_13_3653, i_13_3685, i_13_3689, i_13_3707, i_13_3802, i_13_3905, i_13_3923, i_13_4022, i_13_4031, i_13_4256, i_13_4265, i_13_4274, i_13_4336, i_13_4342, i_13_4391, i_13_4450, i_13_4451, i_13_4558, o_13_361);
	kernel_13_362 k_13_362(i_13_38, i_13_40, i_13_72, i_13_73, i_13_108, i_13_173, i_13_226, i_13_252, i_13_271, i_13_355, i_13_363, i_13_364, i_13_441, i_13_442, i_13_453, i_13_468, i_13_469, i_13_558, i_13_559, i_13_643, i_13_666, i_13_667, i_13_732, i_13_796, i_13_839, i_13_945, i_13_946, i_13_947, i_13_1081, i_13_1099, i_13_1100, i_13_1143, i_13_1144, i_13_1307, i_13_1344, i_13_1407, i_13_1443, i_13_1620, i_13_1621, i_13_1719, i_13_1720, i_13_1729, i_13_1773, i_13_1802, i_13_1836, i_13_1837, i_13_2016, i_13_2169, i_13_2210, i_13_2281, i_13_2299, i_13_2358, i_13_2430, i_13_2431, i_13_2433, i_13_2448, i_13_2468, i_13_2511, i_13_2610, i_13_2611, i_13_2712, i_13_2719, i_13_2757, i_13_2784, i_13_2874, i_13_2880, i_13_2920, i_13_2955, i_13_3026, i_13_3033, i_13_3048, i_13_3060, i_13_3097, i_13_3107, i_13_3127, i_13_3162, i_13_3216, i_13_3231, i_13_3369, i_13_3421, i_13_3467, i_13_3481, i_13_3521, i_13_3528, i_13_3550, i_13_3592, i_13_3595, i_13_3619, i_13_3720, i_13_3727, i_13_3908, i_13_4126, i_13_4215, i_13_4258, i_13_4329, i_13_4340, i_13_4350, i_13_4351, i_13_4446, i_13_4540, o_13_362);
	kernel_13_363 k_13_363(i_13_77, i_13_94, i_13_230, i_13_259, i_13_518, i_13_536, i_13_554, i_13_611, i_13_616, i_13_627, i_13_647, i_13_655, i_13_664, i_13_689, i_13_692, i_13_697, i_13_698, i_13_700, i_13_862, i_13_943, i_13_980, i_13_1025, i_13_1076, i_13_1079, i_13_1121, i_13_1124, i_13_1183, i_13_1214, i_13_1304, i_13_1330, i_13_1331, i_13_1483, i_13_1517, i_13_1519, i_13_1678, i_13_1682, i_13_1735, i_13_1745, i_13_1778, i_13_1795, i_13_1889, i_13_1922, i_13_2024, i_13_2113, i_13_2209, i_13_2212, i_13_2321, i_13_2447, i_13_2455, i_13_2651, i_13_2654, i_13_2696, i_13_2851, i_13_2887, i_13_2888, i_13_2894, i_13_2959, i_13_3030, i_13_3037, i_13_3073, i_13_3091, i_13_3157, i_13_3203, i_13_3208, i_13_3217, i_13_3238, i_13_3265, i_13_3310, i_13_3418, i_13_3482, i_13_3526, i_13_3527, i_13_3571, i_13_3572, i_13_3695, i_13_3742, i_13_3743, i_13_3847, i_13_3866, i_13_3874, i_13_3887, i_13_3930, i_13_4045, i_13_4064, i_13_4081, i_13_4091, i_13_4130, i_13_4162, i_13_4190, i_13_4192, i_13_4193, i_13_4256, i_13_4270, i_13_4336, i_13_4372, i_13_4382, i_13_4460, i_13_4598, i_13_4603, i_13_4604, o_13_363);
	kernel_13_364 k_13_364(i_13_34, i_13_51, i_13_52, i_13_75, i_13_93, i_13_129, i_13_130, i_13_141, i_13_240, i_13_250, i_13_258, i_13_340, i_13_561, i_13_570, i_13_585, i_13_618, i_13_619, i_13_642, i_13_699, i_13_700, i_13_714, i_13_763, i_13_840, i_13_843, i_13_844, i_13_931, i_13_1077, i_13_1078, i_13_1342, i_13_1399, i_13_1401, i_13_1408, i_13_1471, i_13_1482, i_13_1527, i_13_1552, i_13_1572, i_13_1608, i_13_1635, i_13_1636, i_13_1660, i_13_1710, i_13_1734, i_13_1912, i_13_1920, i_13_1921, i_13_1992, i_13_2019, i_13_2032, i_13_2055, i_13_2277, i_13_2280, i_13_2311, i_13_2454, i_13_2505, i_13_2551, i_13_2569, i_13_2670, i_13_2724, i_13_2787, i_13_2847, i_13_2854, i_13_2857, i_13_2886, i_13_2887, i_13_2958, i_13_2959, i_13_3063, i_13_3145, i_13_3244, i_13_3315, i_13_3322, i_13_3372, i_13_3379, i_13_3382, i_13_3451, i_13_3463, i_13_3525, i_13_3540, i_13_3552, i_13_3553, i_13_3613, i_13_3630, i_13_3643, i_13_3646, i_13_3649, i_13_3667, i_13_3687, i_13_3688, i_13_3694, i_13_3724, i_13_3739, i_13_4104, i_13_4162, i_13_4209, i_13_4254, i_13_4390, i_13_4392, i_13_4393, i_13_4395, o_13_364);
	kernel_13_365 k_13_365(i_13_39, i_13_66, i_13_75, i_13_96, i_13_106, i_13_168, i_13_268, i_13_284, i_13_357, i_13_410, i_13_411, i_13_465, i_13_466, i_13_515, i_13_529, i_13_569, i_13_591, i_13_592, i_13_654, i_13_794, i_13_824, i_13_914, i_13_1019, i_13_1021, i_13_1118, i_13_1212, i_13_1229, i_13_1347, i_13_1348, i_13_1391, i_13_1409, i_13_1443, i_13_1446, i_13_1490, i_13_1492, i_13_1501, i_13_1596, i_13_1713, i_13_1776, i_13_1777, i_13_1802, i_13_1884, i_13_1931, i_13_1950, i_13_1960, i_13_2032, i_13_2058, i_13_2059, i_13_2103, i_13_2110, i_13_2202, i_13_2283, i_13_2284, i_13_2347, i_13_2409, i_13_2410, i_13_2444, i_13_2446, i_13_2465, i_13_2514, i_13_2553, i_13_2554, i_13_3173, i_13_3215, i_13_3263, i_13_3353, i_13_3372, i_13_3373, i_13_3390, i_13_3391, i_13_3418, i_13_3425, i_13_3530, i_13_3535, i_13_3579, i_13_3597, i_13_3598, i_13_3621, i_13_3633, i_13_3638, i_13_3755, i_13_3783, i_13_3784, i_13_3785, i_13_3786, i_13_3787, i_13_3800, i_13_3874, i_13_3983, i_13_3990, i_13_4236, i_13_4250, i_13_4263, i_13_4264, i_13_4332, i_13_4367, i_13_4432, i_13_4452, i_13_4453, i_13_4543, o_13_365);
	kernel_13_366 k_13_366(i_13_46, i_13_119, i_13_154, i_13_157, i_13_164, i_13_167, i_13_214, i_13_259, i_13_269, i_13_275, i_13_278, i_13_334, i_13_352, i_13_353, i_13_451, i_13_455, i_13_506, i_13_518, i_13_617, i_13_667, i_13_814, i_13_815, i_13_841, i_13_845, i_13_932, i_13_961, i_13_977, i_13_1066, i_13_1103, i_13_1244, i_13_1327, i_13_1342, i_13_1400, i_13_1402, i_13_1445, i_13_1480, i_13_1508, i_13_1543, i_13_1570, i_13_1573, i_13_1594, i_13_1604, i_13_1649, i_13_1766, i_13_1801, i_13_1805, i_13_1807, i_13_1850, i_13_1852, i_13_1931, i_13_1946, i_13_2026, i_13_2146, i_13_2149, i_13_2201, i_13_2237, i_13_2278, i_13_2303, i_13_2408, i_13_2569, i_13_2585, i_13_2591, i_13_2600, i_13_2621, i_13_2768, i_13_2899, i_13_2965, i_13_2972, i_13_3106, i_13_3112, i_13_3127, i_13_3128, i_13_3215, i_13_3274, i_13_3313, i_13_3379, i_13_3397, i_13_3398, i_13_3400, i_13_3439, i_13_3521, i_13_3592, i_13_3628, i_13_3664, i_13_3739, i_13_3821, i_13_3889, i_13_3899, i_13_4042, i_13_4043, i_13_4061, i_13_4063, i_13_4231, i_13_4253, i_13_4318, i_13_4319, i_13_4348, i_13_4375, i_13_4534, i_13_4556, o_13_366);
	kernel_13_367 k_13_367(i_13_139, i_13_357, i_13_382, i_13_399, i_13_409, i_13_441, i_13_456, i_13_468, i_13_472, i_13_478, i_13_572, i_13_594, i_13_605, i_13_622, i_13_652, i_13_654, i_13_657, i_13_660, i_13_661, i_13_663, i_13_885, i_13_889, i_13_939, i_13_943, i_13_1076, i_13_1114, i_13_1119, i_13_1143, i_13_1144, i_13_1147, i_13_1270, i_13_1515, i_13_1656, i_13_1657, i_13_1660, i_13_1723, i_13_1734, i_13_1741, i_13_1768, i_13_1791, i_13_1792, i_13_1832, i_13_1922, i_13_2002, i_13_2016, i_13_2017, i_13_2019, i_13_2020, i_13_2023, i_13_2057, i_13_2131, i_13_2295, i_13_2320, i_13_2407, i_13_2461, i_13_2469, i_13_2470, i_13_2512, i_13_2534, i_13_2819, i_13_2847, i_13_2955, i_13_2958, i_13_3057, i_13_3075, i_13_3115, i_13_3259, i_13_3352, i_13_3418, i_13_3486, i_13_3489, i_13_3658, i_13_3666, i_13_3729, i_13_3730, i_13_3739, i_13_3742, i_13_3756, i_13_3865, i_13_3901, i_13_3903, i_13_3909, i_13_3910, i_13_3924, i_13_4161, i_13_4162, i_13_4165, i_13_4186, i_13_4217, i_13_4315, i_13_4330, i_13_4332, i_13_4363, i_13_4429, i_13_4432, i_13_4516, i_13_4591, i_13_4599, i_13_4600, i_13_4602, o_13_367);
	kernel_13_368 k_13_368(i_13_25, i_13_28, i_13_64, i_13_65, i_13_131, i_13_156, i_13_212, i_13_253, i_13_308, i_13_356, i_13_373, i_13_376, i_13_397, i_13_469, i_13_524, i_13_535, i_13_667, i_13_668, i_13_712, i_13_725, i_13_758, i_13_829, i_13_830, i_13_850, i_13_896, i_13_929, i_13_947, i_13_1081, i_13_1082, i_13_1099, i_13_1246, i_13_1273, i_13_1274, i_13_1306, i_13_1307, i_13_1397, i_13_1443, i_13_1504, i_13_1505, i_13_1550, i_13_1639, i_13_1714, i_13_1721, i_13_1723, i_13_1774, i_13_1786, i_13_1838, i_13_1847, i_13_1918, i_13_1927, i_13_1999, i_13_2000, i_13_2030, i_13_2101, i_13_2297, i_13_2378, i_13_2395, i_13_2468, i_13_2507, i_13_2512, i_13_2693, i_13_2764, i_13_2875, i_13_2881, i_13_2935, i_13_2936, i_13_2938, i_13_3001, i_13_3037, i_13_3241, i_13_3242, i_13_3251, i_13_3259, i_13_3290, i_13_3376, i_13_3377, i_13_3397, i_13_3415, i_13_3529, i_13_3596, i_13_3620, i_13_3728, i_13_3730, i_13_3754, i_13_3755, i_13_3857, i_13_3935, i_13_3988, i_13_4060, i_13_4213, i_13_4262, i_13_4313, i_13_4330, i_13_4340, i_13_4341, i_13_4429, i_13_4430, i_13_4448, i_13_4511, i_13_4592, o_13_368);
	kernel_13_369 k_13_369(i_13_48, i_13_126, i_13_127, i_13_159, i_13_162, i_13_188, i_13_210, i_13_275, i_13_318, i_13_431, i_13_456, i_13_465, i_13_519, i_13_520, i_13_535, i_13_665, i_13_679, i_13_744, i_13_762, i_13_763, i_13_823, i_13_939, i_13_944, i_13_1103, i_13_1131, i_13_1132, i_13_1230, i_13_1303, i_13_1320, i_13_1392, i_13_1524, i_13_1525, i_13_1551, i_13_1555, i_13_1556, i_13_1602, i_13_1605, i_13_1606, i_13_1698, i_13_1699, i_13_1753, i_13_1803, i_13_1806, i_13_1903, i_13_1961, i_13_1998, i_13_2025, i_13_2106, i_13_2145, i_13_2239, i_13_2277, i_13_2299, i_13_2400, i_13_2472, i_13_2473, i_13_2508, i_13_2709, i_13_2724, i_13_2787, i_13_3075, i_13_3076, i_13_3144, i_13_3198, i_13_3234, i_13_3263, i_13_3264, i_13_3345, i_13_3366, i_13_3368, i_13_3399, i_13_3402, i_13_3460, i_13_3553, i_13_3581, i_13_3639, i_13_3640, i_13_3744, i_13_3780, i_13_3788, i_13_3822, i_13_3823, i_13_3867, i_13_3891, i_13_3900, i_13_3914, i_13_3922, i_13_3933, i_13_4038, i_13_4062, i_13_4206, i_13_4252, i_13_4256, i_13_4272, i_13_4341, i_13_4342, i_13_4448, i_13_4514, i_13_4517, i_13_4576, i_13_4596, o_13_369);
	kernel_13_370 k_13_370(i_13_69, i_13_282, i_13_285, i_13_321, i_13_327, i_13_328, i_13_411, i_13_448, i_13_457, i_13_528, i_13_529, i_13_573, i_13_579, i_13_598, i_13_601, i_13_640, i_13_676, i_13_717, i_13_745, i_13_762, i_13_780, i_13_825, i_13_826, i_13_861, i_13_862, i_13_894, i_13_913, i_13_1023, i_13_1024, i_13_1095, i_13_1134, i_13_1182, i_13_1230, i_13_1258, i_13_1320, i_13_1326, i_13_1347, i_13_1410, i_13_1464, i_13_1635, i_13_1636, i_13_1690, i_13_1713, i_13_1732, i_13_1749, i_13_1816, i_13_1858, i_13_1861, i_13_1884, i_13_1923, i_13_2005, i_13_2110, i_13_2139, i_13_2310, i_13_2454, i_13_2461, i_13_2464, i_13_2502, i_13_2544, i_13_2545, i_13_2559, i_13_2616, i_13_2632, i_13_2652, i_13_2653, i_13_2770, i_13_2874, i_13_3001, i_13_3088, i_13_3174, i_13_3175, i_13_3219, i_13_3321, i_13_3370, i_13_3399, i_13_3432, i_13_3562, i_13_3565, i_13_3630, i_13_3640, i_13_3721, i_13_3732, i_13_3793, i_13_3858, i_13_3876, i_13_3912, i_13_3913, i_13_3922, i_13_3924, i_13_4015, i_13_4078, i_13_4237, i_13_4254, i_13_4255, i_13_4263, i_13_4350, i_13_4380, i_13_4381, i_13_4443, i_13_4567, o_13_370);
	kernel_13_371 k_13_371(i_13_69, i_13_70, i_13_94, i_13_258, i_13_372, i_13_373, i_13_645, i_13_673, i_13_686, i_13_797, i_13_820, i_13_921, i_13_1065, i_13_1103, i_13_1104, i_13_1148, i_13_1274, i_13_1275, i_13_1276, i_13_1297, i_13_1317, i_13_1401, i_13_1402, i_13_1428, i_13_1456, i_13_1469, i_13_1599, i_13_1600, i_13_1644, i_13_1649, i_13_1720, i_13_1722, i_13_1726, i_13_1777, i_13_1780, i_13_1807, i_13_1914, i_13_1923, i_13_1939, i_13_1945, i_13_1946, i_13_1947, i_13_1995, i_13_2026, i_13_2054, i_13_2107, i_13_2193, i_13_2197, i_13_2265, i_13_2279, i_13_2302, i_13_2406, i_13_2472, i_13_2548, i_13_2549, i_13_2568, i_13_2697, i_13_2742, i_13_2747, i_13_2755, i_13_2786, i_13_2884, i_13_2886, i_13_2887, i_13_2899, i_13_2901, i_13_2919, i_13_2940, i_13_2954, i_13_3030, i_13_3130, i_13_3291, i_13_3292, i_13_3367, i_13_3368, i_13_3399, i_13_3459, i_13_3525, i_13_3534, i_13_3570, i_13_3592, i_13_3593, i_13_3594, i_13_3595, i_13_3759, i_13_3785, i_13_3787, i_13_3822, i_13_3908, i_13_3927, i_13_3992, i_13_4037, i_13_4231, i_13_4305, i_13_4308, i_13_4317, i_13_4434, i_13_4448, i_13_4449, i_13_4450, o_13_371);
	kernel_13_372 k_13_372(i_13_118, i_13_125, i_13_179, i_13_191, i_13_195, i_13_196, i_13_197, i_13_303, i_13_575, i_13_614, i_13_664, i_13_712, i_13_719, i_13_772, i_13_800, i_13_862, i_13_863, i_13_932, i_13_943, i_13_952, i_13_953, i_13_1073, i_13_1079, i_13_1226, i_13_1228, i_13_1231, i_13_1232, i_13_1252, i_13_1253, i_13_1259, i_13_1285, i_13_1315, i_13_1318, i_13_1321, i_13_1322, i_13_1410, i_13_1411, i_13_1491, i_13_1492, i_13_1493, i_13_1502, i_13_1538, i_13_1550, i_13_1556, i_13_1573, i_13_1739, i_13_1741, i_13_1781, i_13_1919, i_13_1960, i_13_1961, i_13_2002, i_13_2015, i_13_2059, i_13_2195, i_13_2207, i_13_2242, i_13_2265, i_13_2300, i_13_2314, i_13_2359, i_13_2423, i_13_2536, i_13_2545, i_13_2573, i_13_2617, i_13_2618, i_13_2712, i_13_2918, i_13_3049, i_13_3050, i_13_3117, i_13_3170, i_13_3212, i_13_3220, i_13_3221, i_13_3290, i_13_3346, i_13_3391, i_13_3471, i_13_3475, i_13_3491, i_13_3535, i_13_3536, i_13_3560, i_13_3565, i_13_3575, i_13_3781, i_13_3782, i_13_3859, i_13_3878, i_13_4012, i_13_4013, i_13_4091, i_13_4094, i_13_4252, i_13_4372, i_13_4381, i_13_4520, i_13_4559, o_13_372);
	kernel_13_373 k_13_373(i_13_40, i_13_43, i_13_112, i_13_113, i_13_141, i_13_142, i_13_193, i_13_241, i_13_251, i_13_380, i_13_389, i_13_562, i_13_581, i_13_583, i_13_619, i_13_776, i_13_819, i_13_843, i_13_1083, i_13_1084, i_13_1087, i_13_1098, i_13_1212, i_13_1219, i_13_1273, i_13_1318, i_13_1427, i_13_1429, i_13_1444, i_13_1473, i_13_1474, i_13_1552, i_13_1572, i_13_1602, i_13_1624, i_13_1636, i_13_1681, i_13_1750, i_13_1800, i_13_1804, i_13_1817, i_13_1840, i_13_1924, i_13_1933, i_13_1943, i_13_1960, i_13_1996, i_13_2005, i_13_2006, i_13_2124, i_13_2187, i_13_2196, i_13_2276, i_13_2428, i_13_2434, i_13_2437, i_13_2455, i_13_2646, i_13_2713, i_13_2716, i_13_2717, i_13_2726, i_13_2858, i_13_2958, i_13_3010, i_13_3038, i_13_3064, i_13_3066, i_13_3067, i_13_3146, i_13_3227, i_13_3258, i_13_3326, i_13_3373, i_13_3374, i_13_3440, i_13_3442, i_13_3526, i_13_3537, i_13_3541, i_13_3559, i_13_3564, i_13_3573, i_13_3649, i_13_3653, i_13_3685, i_13_3686, i_13_3687, i_13_3688, i_13_3689, i_13_3726, i_13_3780, i_13_3852, i_13_3856, i_13_4021, i_13_4057, i_13_4093, i_13_4230, i_13_4257, i_13_4400, o_13_373);
	kernel_13_374 k_13_374(i_13_30, i_13_63, i_13_64, i_13_79, i_13_99, i_13_112, i_13_162, i_13_199, i_13_225, i_13_272, i_13_357, i_13_370, i_13_396, i_13_405, i_13_428, i_13_445, i_13_468, i_13_470, i_13_489, i_13_568, i_13_622, i_13_684, i_13_695, i_13_810, i_13_956, i_13_1017, i_13_1098, i_13_1263, i_13_1269, i_13_1296, i_13_1363, i_13_1424, i_13_1432, i_13_1478, i_13_1503, i_13_1504, i_13_1593, i_13_1638, i_13_1642, i_13_1643, i_13_1688, i_13_1719, i_13_1720, i_13_1791, i_13_1792, i_13_1828, i_13_1881, i_13_1927, i_13_2015, i_13_2100, i_13_2103, i_13_2111, i_13_2179, i_13_2235, i_13_2238, i_13_2246, i_13_2376, i_13_2377, i_13_2378, i_13_2444, i_13_2558, i_13_2720, i_13_2749, i_13_2917, i_13_2934, i_13_2935, i_13_3171, i_13_3241, i_13_3262, i_13_3305, i_13_3396, i_13_3450, i_13_3451, i_13_3479, i_13_3566, i_13_3648, i_13_3762, i_13_3763, i_13_3790, i_13_3859, i_13_3865, i_13_3893, i_13_3987, i_13_3988, i_13_4050, i_13_4051, i_13_4078, i_13_4159, i_13_4212, i_13_4215, i_13_4234, i_13_4303, i_13_4312, i_13_4369, i_13_4375, i_13_4379, i_13_4410, i_13_4432, i_13_4512, i_13_4582, o_13_374);
	kernel_13_375 k_13_375(i_13_46, i_13_49, i_13_71, i_13_136, i_13_190, i_13_316, i_13_338, i_13_362, i_13_373, i_13_412, i_13_415, i_13_550, i_13_568, i_13_626, i_13_651, i_13_662, i_13_811, i_13_836, i_13_851, i_13_934, i_13_937, i_13_939, i_13_940, i_13_1018, i_13_1022, i_13_1072, i_13_1101, i_13_1102, i_13_1104, i_13_1105, i_13_1119, i_13_1120, i_13_1230, i_13_1391, i_13_1407, i_13_1508, i_13_1544, i_13_1549, i_13_1603, i_13_1661, i_13_1668, i_13_1736, i_13_1768, i_13_1796, i_13_1798, i_13_1799, i_13_1858, i_13_2020, i_13_2021, i_13_2145, i_13_2301, i_13_2381, i_13_2461, i_13_2469, i_13_2470, i_13_2471, i_13_2473, i_13_2474, i_13_2677, i_13_2857, i_13_2858, i_13_2907, i_13_2966, i_13_2969, i_13_2986, i_13_3029, i_13_3031, i_13_3032, i_13_3077, i_13_3117, i_13_3128, i_13_3204, i_13_3210, i_13_3261, i_13_3265, i_13_3272, i_13_3380, i_13_3404, i_13_3457, i_13_3476, i_13_3482, i_13_3484, i_13_3505, i_13_3548, i_13_3568, i_13_3666, i_13_3823, i_13_3898, i_13_3899, i_13_3901, i_13_3964, i_13_4018, i_13_4069, i_13_4090, i_13_4116, i_13_4204, i_13_4298, i_13_4505, i_13_4604, i_13_4607, o_13_375);
	kernel_13_376 k_13_376(i_13_49, i_13_67, i_13_70, i_13_178, i_13_259, i_13_276, i_13_277, i_13_310, i_13_355, i_13_476, i_13_520, i_13_535, i_13_619, i_13_642, i_13_651, i_13_673, i_13_745, i_13_922, i_13_934, i_13_1024, i_13_1104, i_13_1105, i_13_1132, i_13_1276, i_13_1330, i_13_1401, i_13_1402, i_13_1481, i_13_1510, i_13_1564, i_13_1573, i_13_1574, i_13_1597, i_13_1641, i_13_1653, i_13_1659, i_13_1723, i_13_1735, i_13_1779, i_13_1835, i_13_1914, i_13_1923, i_13_1924, i_13_1932, i_13_1947, i_13_2019, i_13_2022, i_13_2028, i_13_2029, i_13_2185, i_13_2196, i_13_2199, i_13_2302, i_13_2436, i_13_2454, i_13_2469, i_13_2473, i_13_2518, i_13_2677, i_13_2697, i_13_2742, i_13_2743, i_13_2769, i_13_2770, i_13_2850, i_13_2923, i_13_2940, i_13_2968, i_13_3030, i_13_3031, i_13_3077, i_13_3110, i_13_3121, i_13_3130, i_13_3246, i_13_3291, i_13_3315, i_13_3381, i_13_3418, i_13_3453, i_13_3525, i_13_3577, i_13_3595, i_13_3625, i_13_3785, i_13_3786, i_13_3787, i_13_3819, i_13_3822, i_13_3901, i_13_3930, i_13_4029, i_13_4093, i_13_4323, i_13_4324, i_13_4325, i_13_4390, i_13_4434, i_13_4516, i_13_4606, o_13_376);
	kernel_13_377 k_13_377(i_13_98, i_13_107, i_13_113, i_13_140, i_13_251, i_13_262, i_13_368, i_13_370, i_13_538, i_13_554, i_13_562, i_13_608, i_13_620, i_13_647, i_13_655, i_13_661, i_13_671, i_13_680, i_13_845, i_13_949, i_13_1070, i_13_1087, i_13_1145, i_13_1148, i_13_1219, i_13_1220, i_13_1264, i_13_1318, i_13_1348, i_13_1474, i_13_1519, i_13_1520, i_13_1574, i_13_1624, i_13_1727, i_13_1742, i_13_1745, i_13_1789, i_13_1840, i_13_1841, i_13_2024, i_13_2137, i_13_2173, i_13_2284, i_13_2285, i_13_2348, i_13_2380, i_13_2417, i_13_2435, i_13_2437, i_13_2438, i_13_2501, i_13_2510, i_13_2599, i_13_2680, i_13_2716, i_13_2717, i_13_2749, i_13_2879, i_13_2906, i_13_2987, i_13_3047, i_13_3053, i_13_3059, i_13_3067, i_13_3100, i_13_3130, i_13_3131, i_13_3148, i_13_3149, i_13_3166, i_13_3167, i_13_3329, i_13_3343, i_13_3347, i_13_3373, i_13_3455, i_13_3464, i_13_3478, i_13_3527, i_13_3623, i_13_3632, i_13_4021, i_13_4049, i_13_4100, i_13_4120, i_13_4121, i_13_4192, i_13_4262, i_13_4264, i_13_4321, i_13_4328, i_13_4343, i_13_4354, i_13_4418, i_13_4460, i_13_4463, i_13_4543, i_13_4544, i_13_4604, o_13_377);
	kernel_13_378 k_13_378(i_13_31, i_13_99, i_13_139, i_13_155, i_13_210, i_13_228, i_13_229, i_13_237, i_13_247, i_13_372, i_13_513, i_13_514, i_13_517, i_13_535, i_13_569, i_13_606, i_13_652, i_13_823, i_13_840, i_13_983, i_13_984, i_13_985, i_13_1025, i_13_1063, i_13_1075, i_13_1112, i_13_1192, i_13_1219, i_13_1300, i_13_1324, i_13_1326, i_13_1327, i_13_1447, i_13_1476, i_13_1489, i_13_1525, i_13_1549, i_13_1569, i_13_1570, i_13_1584, i_13_1670, i_13_1714, i_13_1723, i_13_1746, i_13_1831, i_13_1848, i_13_1936, i_13_2002, i_13_2025, i_13_2029, i_13_2107, i_13_2108, i_13_2116, i_13_2182, i_13_2233, i_13_2259, i_13_2377, i_13_2406, i_13_2489, i_13_2557, i_13_2673, i_13_2677, i_13_2736, i_13_2848, i_13_2966, i_13_3006, i_13_3007, i_13_3108, i_13_3109, i_13_3150, i_13_3151, i_13_3209, i_13_3226, i_13_3313, i_13_3376, i_13_3388, i_13_3406, i_13_3439, i_13_3460, i_13_3485, i_13_3546, i_13_3554, i_13_3730, i_13_3763, i_13_3766, i_13_3817, i_13_3861, i_13_3900, i_13_3977, i_13_4063, i_13_4123, i_13_4158, i_13_4452, i_13_4455, i_13_4513, i_13_4554, i_13_4556, i_13_4564, i_13_4568, i_13_4600, o_13_378);
	kernel_13_379 k_13_379(i_13_28, i_13_100, i_13_109, i_13_163, i_13_184, i_13_298, i_13_317, i_13_382, i_13_415, i_13_416, i_13_470, i_13_568, i_13_640, i_13_686, i_13_743, i_13_794, i_13_797, i_13_856, i_13_886, i_13_947, i_13_1072, i_13_1073, i_13_1093, i_13_1129, i_13_1225, i_13_1252, i_13_1253, i_13_1268, i_13_1280, i_13_1301, i_13_1361, i_13_1424, i_13_1484, i_13_1486, i_13_1499, i_13_1526, i_13_1550, i_13_1603, i_13_1621, i_13_1631, i_13_1690, i_13_1691, i_13_1720, i_13_1814, i_13_2000, i_13_2237, i_13_2260, i_13_2444, i_13_2458, i_13_2459, i_13_2498, i_13_2503, i_13_2506, i_13_2530, i_13_2535, i_13_2539, i_13_2560, i_13_2567, i_13_2576, i_13_2600, i_13_2611, i_13_2612, i_13_2675, i_13_2882, i_13_2948, i_13_3136, i_13_3344, i_13_3349, i_13_3388, i_13_3457, i_13_3458, i_13_3476, i_13_3529, i_13_3539, i_13_3544, i_13_3566, i_13_3619, i_13_3620, i_13_3638, i_13_3683, i_13_3718, i_13_3739, i_13_3766, i_13_3818, i_13_3844, i_13_3845, i_13_3908, i_13_3920, i_13_3983, i_13_4007, i_13_4186, i_13_4204, i_13_4315, i_13_4330, i_13_4339, i_13_4340, i_13_4342, i_13_4519, i_13_4582, i_13_4595, o_13_379);
	kernel_13_380 k_13_380(i_13_48, i_13_78, i_13_102, i_13_121, i_13_157, i_13_169, i_13_188, i_13_197, i_13_259, i_13_274, i_13_275, i_13_283, i_13_337, i_13_338, i_13_431, i_13_454, i_13_556, i_13_588, i_13_612, i_13_616, i_13_620, i_13_664, i_13_669, i_13_709, i_13_850, i_13_926, i_13_953, i_13_1191, i_13_1301, i_13_1329, i_13_1346, i_13_1377, i_13_1399, i_13_1400, i_13_1469, i_13_1529, i_13_1571, i_13_1643, i_13_1678, i_13_1724, i_13_1727, i_13_1735, i_13_1736, i_13_1750, i_13_1852, i_13_1921, i_13_1993, i_13_2002, i_13_2081, i_13_2118, i_13_2137, i_13_2138, i_13_2148, i_13_2191, i_13_2210, i_13_2363, i_13_2408, i_13_2425, i_13_2542, i_13_2617, i_13_2618, i_13_2699, i_13_2708, i_13_2786, i_13_2885, i_13_2888, i_13_3027, i_13_3038, i_13_3039, i_13_3040, i_13_3041, i_13_3050, i_13_3145, i_13_3217, i_13_3386, i_13_3491, i_13_3536, i_13_3640, i_13_3641, i_13_3644, i_13_3702, i_13_3705, i_13_3730, i_13_3758, i_13_3787, i_13_3892, i_13_4089, i_13_4136, i_13_4230, i_13_4232, i_13_4234, i_13_4235, i_13_4261, i_13_4262, i_13_4305, i_13_4360, i_13_4436, i_13_4449, i_13_4513, i_13_4531, o_13_380);
	kernel_13_381 k_13_381(i_13_112, i_13_175, i_13_178, i_13_186, i_13_225, i_13_237, i_13_273, i_13_282, i_13_283, i_13_310, i_13_361, i_13_375, i_13_469, i_13_471, i_13_490, i_13_573, i_13_574, i_13_642, i_13_643, i_13_645, i_13_646, i_13_647, i_13_687, i_13_688, i_13_690, i_13_691, i_13_702, i_13_717, i_13_760, i_13_862, i_13_1123, i_13_1267, i_13_1308, i_13_1311, i_13_1313, i_13_1399, i_13_1597, i_13_1641, i_13_1642, i_13_1672, i_13_1804, i_13_1857, i_13_1860, i_13_1861, i_13_1884, i_13_1939, i_13_2002, i_13_2029, i_13_2055, i_13_2136, i_13_2137, i_13_2176, i_13_2193, i_13_2263, i_13_2310, i_13_2427, i_13_2586, i_13_2599, i_13_2649, i_13_2650, i_13_2652, i_13_2653, i_13_2654, i_13_2676, i_13_2677, i_13_2680, i_13_2770, i_13_2847, i_13_2851, i_13_2913, i_13_2964, i_13_3003, i_13_3270, i_13_3271, i_13_3273, i_13_3274, i_13_3315, i_13_3378, i_13_3387, i_13_3423, i_13_3424, i_13_3426, i_13_3427, i_13_3478, i_13_3535, i_13_3639, i_13_3732, i_13_3875, i_13_3913, i_13_4018, i_13_4020, i_13_4045, i_13_4077, i_13_4080, i_13_4084, i_13_4162, i_13_4174, i_13_4219, i_13_4426, i_13_4594, o_13_381);
	kernel_13_382 k_13_382(i_13_51, i_13_52, i_13_105, i_13_106, i_13_312, i_13_313, i_13_337, i_13_381, i_13_409, i_13_420, i_13_427, i_13_484, i_13_507, i_13_526, i_13_553, i_13_609, i_13_654, i_13_678, i_13_679, i_13_691, i_13_735, i_13_843, i_13_844, i_13_961, i_13_1042, i_13_1303, i_13_1311, i_13_1329, i_13_1330, i_13_1345, i_13_1407, i_13_1462, i_13_1518, i_13_1519, i_13_1572, i_13_1573, i_13_1677, i_13_1686, i_13_1813, i_13_1861, i_13_1911, i_13_2004, i_13_2023, i_13_2031, i_13_2049, i_13_2094, i_13_2131, i_13_2191, i_13_2209, i_13_2281, i_13_2596, i_13_2640, i_13_2695, i_13_2698, i_13_2722, i_13_2856, i_13_2928, i_13_2938, i_13_2982, i_13_2985, i_13_3090, i_13_3127, i_13_3217, i_13_3291, i_13_3364, i_13_3370, i_13_3372, i_13_3400, i_13_3417, i_13_3439, i_13_3490, i_13_3525, i_13_3526, i_13_3535, i_13_3549, i_13_3561, i_13_3616, i_13_3618, i_13_3648, i_13_3768, i_13_3769, i_13_3822, i_13_3864, i_13_3865, i_13_3891, i_13_3993, i_13_4035, i_13_4047, i_13_4119, i_13_4120, i_13_4161, i_13_4162, i_13_4191, i_13_4270, i_13_4369, i_13_4567, i_13_4597, i_13_4599, i_13_4602, i_13_4603, o_13_382);
	kernel_13_383 k_13_383(i_13_33, i_13_76, i_13_111, i_13_120, i_13_159, i_13_160, i_13_271, i_13_285, i_13_313, i_13_322, i_13_384, i_13_385, i_13_456, i_13_511, i_13_537, i_13_564, i_13_570, i_13_611, i_13_643, i_13_655, i_13_760, i_13_840, i_13_943, i_13_1086, i_13_1087, i_13_1218, i_13_1255, i_13_1302, i_13_1303, i_13_1443, i_13_1473, i_13_1477, i_13_1489, i_13_1509, i_13_1599, i_13_1635, i_13_1636, i_13_1650, i_13_1735, i_13_1789, i_13_1795, i_13_1995, i_13_2056, i_13_2112, i_13_2122, i_13_2173, i_13_2193, i_13_2208, i_13_2242, i_13_2400, i_13_2424, i_13_2436, i_13_2500, i_13_2532, i_13_2541, i_13_2715, i_13_2716, i_13_2847, i_13_2919, i_13_2941, i_13_3000, i_13_3004, i_13_3022, i_13_3028, i_13_3103, i_13_3129, i_13_3147, i_13_3163, i_13_3172, i_13_3261, i_13_3274, i_13_3321, i_13_3346, i_13_3382, i_13_3388, i_13_3580, i_13_3615, i_13_3616, i_13_3702, i_13_3720, i_13_3783, i_13_3796, i_13_3802, i_13_3846, i_13_3873, i_13_3874, i_13_3910, i_13_4008, i_13_4009, i_13_4036, i_13_4045, i_13_4083, i_13_4084, i_13_4093, i_13_4107, i_13_4120, i_13_4236, i_13_4282, i_13_4336, i_13_4417, o_13_383);
	kernel_13_384 k_13_384(i_13_66, i_13_69, i_13_70, i_13_133, i_13_205, i_13_208, i_13_209, i_13_357, i_13_466, i_13_535, i_13_588, i_13_591, i_13_616, i_13_653, i_13_745, i_13_762, i_13_763, i_13_814, i_13_1073, i_13_1131, i_13_1132, i_13_1302, i_13_1303, i_13_1312, i_13_1347, i_13_1445, i_13_1453, i_13_1523, i_13_1524, i_13_1525, i_13_1605, i_13_1649, i_13_1650, i_13_1699, i_13_1717, i_13_1930, i_13_1932, i_13_1933, i_13_1995, i_13_2103, i_13_2125, i_13_2128, i_13_2135, i_13_2145, i_13_2193, i_13_2194, i_13_2195, i_13_2239, i_13_2380, i_13_2418, i_13_2435, i_13_2472, i_13_2553, i_13_2697, i_13_2698, i_13_2699, i_13_2721, i_13_2770, i_13_3129, i_13_3244, i_13_3272, i_13_3308, i_13_3344, i_13_3403, i_13_3541, i_13_3634, i_13_3637, i_13_3639, i_13_3640, i_13_3666, i_13_3718, i_13_3742, i_13_3757, i_13_3766, i_13_3844, i_13_3847, i_13_3871, i_13_3900, i_13_3918, i_13_3940, i_13_3973, i_13_3985, i_13_3994, i_13_4010, i_13_4035, i_13_4036, i_13_4038, i_13_4039, i_13_4060, i_13_4225, i_13_4236, i_13_4272, i_13_4273, i_13_4295, i_13_4309, i_13_4312, i_13_4398, i_13_4593, i_13_4596, i_13_4606, o_13_384);
	kernel_13_385 k_13_385(i_13_76, i_13_79, i_13_115, i_13_285, i_13_409, i_13_471, i_13_520, i_13_525, i_13_597, i_13_609, i_13_660, i_13_663, i_13_664, i_13_700, i_13_798, i_13_825, i_13_831, i_13_841, i_13_852, i_13_940, i_13_942, i_13_1066, i_13_1104, i_13_1147, i_13_1150, i_13_1230, i_13_1231, i_13_1309, i_13_1311, i_13_1317, i_13_1492, i_13_1497, i_13_1524, i_13_1551, i_13_1599, i_13_1659, i_13_1660, i_13_1744, i_13_1794, i_13_1884, i_13_1921, i_13_1929, i_13_1959, i_13_1960, i_13_1965, i_13_2230, i_13_2299, i_13_2334, i_13_2356, i_13_2451, i_13_2454, i_13_2455, i_13_2469, i_13_2553, i_13_2724, i_13_2850, i_13_2883, i_13_2941, i_13_3012, i_13_3028, i_13_3049, i_13_3117, i_13_3135, i_13_3156, i_13_3388, i_13_3478, i_13_3486, i_13_3489, i_13_3490, i_13_3504, i_13_3541, i_13_3543, i_13_3544, i_13_3549, i_13_3579, i_13_3580, i_13_3648, i_13_3742, i_13_3894, i_13_4019, i_13_4054, i_13_4126, i_13_4164, i_13_4165, i_13_4201, i_13_4251, i_13_4254, i_13_4255, i_13_4263, i_13_4264, i_13_4269, i_13_4296, i_13_4318, i_13_4332, i_13_4333, i_13_4396, i_13_4431, i_13_4452, i_13_4461, i_13_4603, o_13_385);
	kernel_13_386 k_13_386(i_13_36, i_13_37, i_13_72, i_13_130, i_13_136, i_13_163, i_13_182, i_13_186, i_13_216, i_13_225, i_13_279, i_13_280, i_13_324, i_13_375, i_13_382, i_13_407, i_13_532, i_13_544, i_13_595, i_13_641, i_13_670, i_13_680, i_13_694, i_13_714, i_13_724, i_13_777, i_13_823, i_13_828, i_13_831, i_13_848, i_13_850, i_13_891, i_13_976, i_13_1022, i_13_1065, i_13_1117, i_13_1217, i_13_1309, i_13_1332, i_13_1380, i_13_1390, i_13_1404, i_13_1461, i_13_1487, i_13_1667, i_13_1710, i_13_1711, i_13_1746, i_13_1828, i_13_1829, i_13_1831, i_13_1858, i_13_1881, i_13_1882, i_13_1884, i_13_1903, i_13_2093, i_13_2120, i_13_2296, i_13_2307, i_13_2342, i_13_2423, i_13_2435, i_13_2629, i_13_2646, i_13_2647, i_13_2649, i_13_2650, i_13_2700, i_13_2745, i_13_2844, i_13_2845, i_13_2871, i_13_2872, i_13_3029, i_13_3109, i_13_3142, i_13_3161, i_13_3171, i_13_3216, i_13_3241, i_13_3384, i_13_3429, i_13_3447, i_13_3559, i_13_3641, i_13_3784, i_13_3790, i_13_3817, i_13_3821, i_13_3854, i_13_3893, i_13_4077, i_13_4096, i_13_4162, i_13_4207, i_13_4348, i_13_4412, i_13_4440, i_13_4567, o_13_386);
	kernel_13_387 k_13_387(i_13_32, i_13_49, i_13_56, i_13_71, i_13_77, i_13_80, i_13_153, i_13_412, i_13_611, i_13_629, i_13_661, i_13_662, i_13_664, i_13_674, i_13_683, i_13_686, i_13_716, i_13_851, i_13_854, i_13_940, i_13_1060, i_13_1071, i_13_1076, i_13_1101, i_13_1105, i_13_1106, i_13_1133, i_13_1151, i_13_1188, i_13_1224, i_13_1228, i_13_1229, i_13_1232, i_13_1244, i_13_1256, i_13_1318, i_13_1345, i_13_1484, i_13_1733, i_13_1765, i_13_1766, i_13_1768, i_13_1787, i_13_1799, i_13_1892, i_13_1927, i_13_1962, i_13_2005, i_13_2023, i_13_2024, i_13_2026, i_13_2212, i_13_2284, i_13_2288, i_13_2434, i_13_2518, i_13_2582, i_13_2852, i_13_2903, i_13_2975, i_13_2987, i_13_3010, i_13_3013, i_13_3027, i_13_3032, i_13_3050, i_13_3064, i_13_3122, i_13_3261, i_13_3355, i_13_3356, i_13_3487, i_13_3539, i_13_3542, i_13_3573, i_13_3574, i_13_3731, i_13_3734, i_13_3755, i_13_3866, i_13_3869, i_13_3928, i_13_3978, i_13_4166, i_13_4212, i_13_4255, i_13_4256, i_13_4302, i_13_4322, i_13_4336, i_13_4343, i_13_4372, i_13_4373, i_13_4382, i_13_4450, i_13_4514, i_13_4516, i_13_4598, i_13_4606, i_13_4607, o_13_387);
	kernel_13_388 k_13_388(i_13_31, i_13_53, i_13_103, i_13_125, i_13_142, i_13_143, i_13_241, i_13_251, i_13_278, i_13_322, i_13_340, i_13_449, i_13_508, i_13_575, i_13_619, i_13_620, i_13_728, i_13_781, i_13_850, i_13_980, i_13_1079, i_13_1084, i_13_1250, i_13_1265, i_13_1309, i_13_1364, i_13_1402, i_13_1436, i_13_1498, i_13_1502, i_13_1529, i_13_1566, i_13_1609, i_13_1636, i_13_1637, i_13_1726, i_13_1735, i_13_1796, i_13_1817, i_13_1907, i_13_1913, i_13_1921, i_13_1930, i_13_1989, i_13_2097, i_13_2120, i_13_2294, i_13_2358, i_13_2545, i_13_2564, i_13_2570, i_13_2596, i_13_2709, i_13_2768, i_13_2788, i_13_2789, i_13_2844, i_13_2848, i_13_2959, i_13_3004, i_13_3070, i_13_3130, i_13_3131, i_13_3167, i_13_3220, i_13_3221, i_13_3253, i_13_3374, i_13_3383, i_13_3411, i_13_3416, i_13_3418, i_13_3419, i_13_3447, i_13_3527, i_13_3554, i_13_3581, i_13_3641, i_13_3643, i_13_3662, i_13_3688, i_13_3740, i_13_3788, i_13_3847, i_13_3856, i_13_3874, i_13_3875, i_13_3914, i_13_4012, i_13_4057, i_13_4084, i_13_4090, i_13_4091, i_13_4108, i_13_4171, i_13_4271, i_13_4364, i_13_4391, i_13_4415, i_13_4526, o_13_388);
	kernel_13_389 k_13_389(i_13_28, i_13_37, i_13_48, i_13_63, i_13_64, i_13_65, i_13_198, i_13_352, i_13_354, i_13_361, i_13_378, i_13_462, i_13_588, i_13_668, i_13_685, i_13_694, i_13_712, i_13_756, i_13_823, i_13_828, i_13_838, i_13_859, i_13_909, i_13_1117, i_13_1137, i_13_1296, i_13_1304, i_13_1306, i_13_1309, i_13_1345, i_13_1372, i_13_1396, i_13_1405, i_13_1503, i_13_1504, i_13_1517, i_13_1543, i_13_1557, i_13_1593, i_13_1594, i_13_1638, i_13_1639, i_13_1669, i_13_1710, i_13_1732, i_13_1740, i_13_1858, i_13_1927, i_13_2056, i_13_2071, i_13_2124, i_13_2142, i_13_2189, i_13_2281, i_13_2317, i_13_2377, i_13_2395, i_13_2461, i_13_2478, i_13_2511, i_13_2539, i_13_2691, i_13_2718, i_13_2719, i_13_2720, i_13_2912, i_13_3052, i_13_3060, i_13_3109, i_13_3163, i_13_3172, i_13_3388, i_13_3414, i_13_3532, i_13_3594, i_13_3595, i_13_3609, i_13_3618, i_13_3637, i_13_3766, i_13_3863, i_13_3910, i_13_3916, i_13_3924, i_13_4032, i_13_4033, i_13_4036, i_13_4063, i_13_4213, i_13_4262, i_13_4302, i_13_4307, i_13_4312, i_13_4315, i_13_4330, i_13_4396, i_13_4429, i_13_4430, i_13_4477, i_13_4591, o_13_389);
	kernel_13_390 k_13_390(i_13_72, i_13_121, i_13_139, i_13_165, i_13_173, i_13_175, i_13_311, i_13_523, i_13_526, i_13_532, i_13_535, i_13_796, i_13_798, i_13_811, i_13_814, i_13_848, i_13_850, i_13_851, i_13_958, i_13_985, i_13_1073, i_13_1079, i_13_1225, i_13_1228, i_13_1258, i_13_1411, i_13_1468, i_13_1471, i_13_1497, i_13_1549, i_13_1550, i_13_1552, i_13_1624, i_13_1750, i_13_1803, i_13_1831, i_13_1846, i_13_1858, i_13_1922, i_13_1925, i_13_1957, i_13_2124, i_13_2133, i_13_2203, i_13_2303, i_13_2408, i_13_2458, i_13_2570, i_13_2614, i_13_2785, i_13_2884, i_13_2918, i_13_3007, i_13_3010, i_13_3037, i_13_3061, i_13_3100, i_13_3108, i_13_3109, i_13_3268, i_13_3271, i_13_3274, i_13_3342, i_13_3396, i_13_3402, i_13_3409, i_13_3464, i_13_3469, i_13_3539, i_13_3541, i_13_3568, i_13_3604, i_13_3663, i_13_3666, i_13_3727, i_13_3728, i_13_3729, i_13_3838, i_13_3856, i_13_3869, i_13_3907, i_13_3909, i_13_3911, i_13_3928, i_13_4018, i_13_4054, i_13_4099, i_13_4249, i_13_4251, i_13_4252, i_13_4253, i_13_4255, i_13_4256, i_13_4258, i_13_4259, i_13_4277, i_13_4375, i_13_4376, i_13_4540, i_13_4557, o_13_390);
	kernel_13_391 k_13_391(i_13_259, i_13_311, i_13_328, i_13_329, i_13_562, i_13_583, i_13_611, i_13_628, i_13_629, i_13_823, i_13_826, i_13_862, i_13_863, i_13_894, i_13_1024, i_13_1025, i_13_1033, i_13_1076, i_13_1096, i_13_1097, i_13_1228, i_13_1229, i_13_1232, i_13_1256, i_13_1258, i_13_1259, i_13_1320, i_13_1321, i_13_1327, i_13_1384, i_13_1439, i_13_1483, i_13_1484, i_13_1490, i_13_1492, i_13_1679, i_13_1691, i_13_1780, i_13_1781, i_13_1789, i_13_1858, i_13_1859, i_13_1861, i_13_1862, i_13_1886, i_13_1889, i_13_2030, i_13_2056, i_13_2123, i_13_2150, i_13_2230, i_13_2312, i_13_2461, i_13_2465, i_13_2509, i_13_2510, i_13_2570, i_13_2851, i_13_2852, i_13_2875, i_13_2876, i_13_2977, i_13_3001, i_13_3064, i_13_3094, i_13_3100, i_13_3101, i_13_3122, i_13_3157, i_13_3173, i_13_3176, i_13_3211, i_13_3432, i_13_3433, i_13_3460, i_13_3479, i_13_3488, i_13_3506, i_13_3524, i_13_3535, i_13_3536, i_13_3542, i_13_3545, i_13_3563, i_13_3707, i_13_3785, i_13_3835, i_13_3857, i_13_3895, i_13_3911, i_13_3914, i_13_4036, i_13_4207, i_13_4255, i_13_4342, i_13_4373, i_13_4378, i_13_4381, i_13_4382, i_13_4594, o_13_391);
	kernel_13_392 k_13_392(i_13_30, i_13_67, i_13_72, i_13_73, i_13_103, i_13_108, i_13_255, i_13_282, i_13_297, i_13_354, i_13_355, i_13_358, i_13_360, i_13_369, i_13_373, i_13_396, i_13_468, i_13_523, i_13_588, i_13_603, i_13_639, i_13_666, i_13_667, i_13_741, i_13_742, i_13_759, i_13_828, i_13_838, i_13_945, i_13_946, i_13_975, i_13_1084, i_13_1209, i_13_1304, i_13_1344, i_13_1504, i_13_1620, i_13_1683, i_13_1693, i_13_1774, i_13_1777, i_13_1947, i_13_1999, i_13_2055, i_13_2056, i_13_2169, i_13_2181, i_13_2280, i_13_2281, i_13_2298, i_13_2348, i_13_2350, i_13_2430, i_13_2431, i_13_2469, i_13_2511, i_13_2512, i_13_2539, i_13_2613, i_13_2614, i_13_2691, i_13_2692, i_13_2721, i_13_2880, i_13_2881, i_13_2907, i_13_2916, i_13_3007, i_13_3385, i_13_3387, i_13_3528, i_13_3558, i_13_3594, i_13_3595, i_13_3599, i_13_3613, i_13_3618, i_13_3619, i_13_3631, i_13_3634, i_13_3636, i_13_3685, i_13_3726, i_13_3978, i_13_3987, i_13_4041, i_13_4117, i_13_4123, i_13_4188, i_13_4202, i_13_4233, i_13_4260, i_13_4329, i_13_4330, i_13_4365, i_13_4366, i_13_4410, i_13_4428, i_13_4429, i_13_4450, o_13_392);
	kernel_13_393 k_13_393(i_13_19, i_13_73, i_13_94, i_13_355, i_13_443, i_13_530, i_13_628, i_13_695, i_13_697, i_13_706, i_13_831, i_13_886, i_13_1022, i_13_1066, i_13_1072, i_13_1073, i_13_1100, i_13_1112, i_13_1208, i_13_1210, i_13_1217, i_13_1258, i_13_1286, i_13_1337, i_13_1399, i_13_1419, i_13_1424, i_13_1427, i_13_1491, i_13_1499, i_13_1522, i_13_1658, i_13_1732, i_13_1774, i_13_1775, i_13_1837, i_13_1960, i_13_1966, i_13_2006, i_13_2020, i_13_2021, i_13_2029, i_13_2045, i_13_2144, i_13_2209, i_13_2232, i_13_2281, i_13_2297, i_13_2347, i_13_2425, i_13_2443, i_13_2444, i_13_2446, i_13_2449, i_13_2453, i_13_2454, i_13_2512, i_13_2515, i_13_2555, i_13_2693, i_13_2719, i_13_2822, i_13_2884, i_13_2896, i_13_3037, i_13_3074, i_13_3307, i_13_3370, i_13_3416, i_13_3442, i_13_3547, i_13_3568, i_13_3578, i_13_3579, i_13_3598, i_13_3620, i_13_3634, i_13_3682, i_13_3740, i_13_3756, i_13_3806, i_13_3958, i_13_3967, i_13_3989, i_13_4018, i_13_4039, i_13_4208, i_13_4263, i_13_4272, i_13_4330, i_13_4332, i_13_4333, i_13_4379, i_13_4430, i_13_4453, i_13_4510, i_13_4513, i_13_4594, i_13_4596, i_13_4604, o_13_393);
	kernel_13_394 k_13_394(i_13_58, i_13_59, i_13_140, i_13_190, i_13_256, i_13_259, i_13_334, i_13_428, i_13_484, i_13_485, i_13_612, i_13_625, i_13_626, i_13_628, i_13_629, i_13_657, i_13_685, i_13_779, i_13_781, i_13_913, i_13_914, i_13_977, i_13_980, i_13_1094, i_13_1115, i_13_1117, i_13_1228, i_13_1263, i_13_1274, i_13_1318, i_13_1343, i_13_1469, i_13_1480, i_13_1481, i_13_1484, i_13_1512, i_13_1561, i_13_1633, i_13_1639, i_13_1648, i_13_1649, i_13_1670, i_13_1673, i_13_1696, i_13_1733, i_13_1756, i_13_1778, i_13_1796, i_13_1801, i_13_1886, i_13_2180, i_13_2230, i_13_2307, i_13_2308, i_13_2366, i_13_2377, i_13_2380, i_13_2381, i_13_2425, i_13_2447, i_13_2461, i_13_2483, i_13_2647, i_13_2743, i_13_2781, i_13_2783, i_13_2849, i_13_2899, i_13_2950, i_13_2951, i_13_2953, i_13_3001, i_13_3005, i_13_3074, i_13_3091, i_13_3110, i_13_3135, i_13_3145, i_13_3153, i_13_3163, i_13_3308, i_13_3356, i_13_3433, i_13_3529, i_13_3637, i_13_3754, i_13_3766, i_13_3799, i_13_3842, i_13_3843, i_13_3874, i_13_4018, i_13_4187, i_13_4231, i_13_4294, i_13_4391, i_13_4448, i_13_4468, i_13_4481, i_13_4508, o_13_394);
	kernel_13_395 k_13_395(i_13_28, i_13_52, i_13_126, i_13_253, i_13_274, i_13_279, i_13_282, i_13_306, i_13_307, i_13_310, i_13_315, i_13_316, i_13_334, i_13_371, i_13_373, i_13_453, i_13_504, i_13_589, i_13_615, i_13_616, i_13_642, i_13_643, i_13_679, i_13_685, i_13_687, i_13_688, i_13_757, i_13_819, i_13_820, i_13_832, i_13_858, i_13_976, i_13_1075, i_13_1138, i_13_1222, i_13_1228, i_13_1284, i_13_1404, i_13_1422, i_13_1426, i_13_1518, i_13_1594, i_13_1597, i_13_1768, i_13_1813, i_13_1819, i_13_1827, i_13_1926, i_13_1999, i_13_2175, i_13_2200, i_13_2434, i_13_2436, i_13_2443, i_13_2497, i_13_2647, i_13_2673, i_13_2676, i_13_2695, i_13_2707, i_13_2713, i_13_2715, i_13_2740, i_13_2767, i_13_2845, i_13_2853, i_13_2883, i_13_2884, i_13_3087, i_13_3102, i_13_3106, i_13_3205, i_13_3207, i_13_3217, i_13_3415, i_13_3441, i_13_3457, i_13_3460, i_13_3486, i_13_3609, i_13_3688, i_13_3720, i_13_3726, i_13_3735, i_13_3736, i_13_3769, i_13_3888, i_13_3889, i_13_3919, i_13_4014, i_13_4015, i_13_4032, i_13_4033, i_13_4162, i_13_4269, i_13_4381, i_13_4392, i_13_4393, i_13_4513, i_13_4594, o_13_395);
	kernel_13_396 k_13_396(i_13_46, i_13_73, i_13_92, i_13_119, i_13_173, i_13_175, i_13_181, i_13_307, i_13_311, i_13_409, i_13_550, i_13_551, i_13_568, i_13_569, i_13_626, i_13_643, i_13_649, i_13_686, i_13_847, i_13_848, i_13_937, i_13_982, i_13_983, i_13_1120, i_13_1129, i_13_1130, i_13_1136, i_13_1253, i_13_1324, i_13_1328, i_13_1361, i_13_1372, i_13_1405, i_13_1406, i_13_1468, i_13_1523, i_13_1630, i_13_1750, i_13_1751, i_13_1778, i_13_1805, i_13_1936, i_13_2021, i_13_2098, i_13_2120, i_13_2264, i_13_2287, i_13_2384, i_13_2470, i_13_2507, i_13_2543, i_13_2567, i_13_2593, i_13_2692, i_13_2696, i_13_2851, i_13_2884, i_13_2900, i_13_2926, i_13_2980, i_13_2983, i_13_3002, i_13_3007, i_13_3029, i_13_3047, i_13_3106, i_13_3107, i_13_3172, i_13_3209, i_13_3262, i_13_3344, i_13_3403, i_13_3407, i_13_3485, i_13_3547, i_13_3568, i_13_3638, i_13_3640, i_13_3685, i_13_3754, i_13_3764, i_13_3802, i_13_3820, i_13_3821, i_13_3892, i_13_3898, i_13_3908, i_13_3992, i_13_4036, i_13_4081, i_13_4250, i_13_4262, i_13_4322, i_13_4399, i_13_4402, i_13_4495, i_13_4564, i_13_4565, i_13_4595, i_13_4604, o_13_396);
	kernel_13_397 k_13_397(i_13_30, i_13_31, i_13_58, i_13_90, i_13_91, i_13_108, i_13_228, i_13_459, i_13_534, i_13_660, i_13_685, i_13_732, i_13_742, i_13_757, i_13_793, i_13_811, i_13_850, i_13_855, i_13_957, i_13_958, i_13_1075, i_13_1083, i_13_1084, i_13_1117, i_13_1215, i_13_1228, i_13_1324, i_13_1462, i_13_1470, i_13_1485, i_13_1486, i_13_1677, i_13_1758, i_13_1813, i_13_1836, i_13_1899, i_13_1957, i_13_1998, i_13_1999, i_13_2043, i_13_2205, i_13_2227, i_13_2259, i_13_2286, i_13_2313, i_13_2421, i_13_2431, i_13_2497, i_13_2529, i_13_2538, i_13_2539, i_13_2563, i_13_2712, i_13_2731, i_13_2916, i_13_2917, i_13_2937, i_13_2979, i_13_3018, i_13_3019, i_13_3025, i_13_3043, i_13_3088, i_13_3099, i_13_3106, i_13_3126, i_13_3144, i_13_3145, i_13_3168, i_13_3325, i_13_3385, i_13_3457, i_13_3486, i_13_3487, i_13_3577, i_13_3609, i_13_3616, i_13_3622, i_13_3717, i_13_3802, i_13_3844, i_13_3846, i_13_3870, i_13_3871, i_13_3880, i_13_3906, i_13_3919, i_13_4006, i_13_4032, i_13_4054, i_13_4116, i_13_4121, i_13_4174, i_13_4186, i_13_4294, i_13_4347, i_13_4396, i_13_4521, i_13_4542, i_13_4557, o_13_397);
	kernel_13_398 k_13_398(i_13_124, i_13_139, i_13_165, i_13_169, i_13_179, i_13_229, i_13_258, i_13_283, i_13_284, i_13_285, i_13_286, i_13_414, i_13_512, i_13_517, i_13_572, i_13_662, i_13_768, i_13_817, i_13_849, i_13_850, i_13_853, i_13_984, i_13_985, i_13_1019, i_13_1021, i_13_1022, i_13_1037, i_13_1226, i_13_1310, i_13_1313, i_13_1334, i_13_1344, i_13_1506, i_13_1549, i_13_1550, i_13_1714, i_13_1723, i_13_1749, i_13_1786, i_13_1858, i_13_1859, i_13_1860, i_13_1861, i_13_1921, i_13_2014, i_13_2142, i_13_2298, i_13_2407, i_13_2657, i_13_2680, i_13_2852, i_13_2857, i_13_2967, i_13_3010, i_13_3011, i_13_3014, i_13_3030, i_13_3037, i_13_3040, i_13_3108, i_13_3109, i_13_3112, i_13_3122, i_13_3163, i_13_3217, i_13_3218, i_13_3400, i_13_3542, i_13_3577, i_13_3636, i_13_3785, i_13_3838, i_13_3847, i_13_3856, i_13_3861, i_13_3865, i_13_3866, i_13_3868, i_13_3892, i_13_3910, i_13_3911, i_13_3913, i_13_3916, i_13_3936, i_13_3982, i_13_4047, i_13_4066, i_13_4162, i_13_4170, i_13_4204, i_13_4207, i_13_4250, i_13_4253, i_13_4258, i_13_4261, i_13_4304, i_13_4345, i_13_4351, i_13_4358, i_13_4379, o_13_398);
	kernel_13_399 k_13_399(i_13_29, i_13_91, i_13_95, i_13_104, i_13_118, i_13_119, i_13_158, i_13_164, i_13_181, i_13_182, i_13_224, i_13_383, i_13_395, i_13_454, i_13_515, i_13_523, i_13_568, i_13_572, i_13_697, i_13_824, i_13_856, i_13_868, i_13_913, i_13_946, i_13_1076, i_13_1085, i_13_1118, i_13_1190, i_13_1216, i_13_1301, i_13_1360, i_13_1361, i_13_1406, i_13_1606, i_13_1621, i_13_1694, i_13_1723, i_13_1786, i_13_1787, i_13_1805, i_13_1906, i_13_1907, i_13_1918, i_13_2000, i_13_2173, i_13_2174, i_13_2206, i_13_2209, i_13_2422, i_13_2431, i_13_2432, i_13_2434, i_13_2435, i_13_2552, i_13_2956, i_13_2984, i_13_3020, i_13_3101, i_13_3145, i_13_3146, i_13_3161, i_13_3163, i_13_3164, i_13_3205, i_13_3209, i_13_3235, i_13_3344, i_13_3380, i_13_3421, i_13_3461, i_13_3487, i_13_3488, i_13_3530, i_13_3533, i_13_3541, i_13_3542, i_13_3577, i_13_3700, i_13_3718, i_13_3728, i_13_3764, i_13_3784, i_13_3794, i_13_3844, i_13_3871, i_13_3872, i_13_3983, i_13_4006, i_13_4007, i_13_4118, i_13_4132, i_13_4204, i_13_4325, i_13_4348, i_13_4349, i_13_4351, i_13_4415, i_13_4583, i_13_4588, i_13_4589, o_13_399);
	kernel_13_400 k_13_400(i_13_71, i_13_74, i_13_76, i_13_79, i_13_80, i_13_139, i_13_176, i_13_309, i_13_323, i_13_358, i_13_376, i_13_610, i_13_647, i_13_672, i_13_673, i_13_674, i_13_683, i_13_772, i_13_814, i_13_821, i_13_841, i_13_952, i_13_1103, i_13_1106, i_13_1123, i_13_1151, i_13_1210, i_13_1276, i_13_1277, i_13_1282, i_13_1312, i_13_1403, i_13_1430, i_13_1468, i_13_1496, i_13_1509, i_13_1511, i_13_1600, i_13_1645, i_13_1687, i_13_1690, i_13_1726, i_13_1736, i_13_1750, i_13_1781, i_13_1798, i_13_1799, i_13_1857, i_13_1889, i_13_1912, i_13_1925, i_13_2002, i_13_2030, i_13_2032, i_13_2176, i_13_2177, i_13_2232, i_13_2240, i_13_2344, i_13_2407, i_13_2513, i_13_2654, i_13_2679, i_13_2680, i_13_2681, i_13_2698, i_13_2817, i_13_2818, i_13_2851, i_13_2852, i_13_2924, i_13_3028, i_13_3142, i_13_3221, i_13_3355, i_13_3386, i_13_3406, i_13_3607, i_13_3622, i_13_3739, i_13_3743, i_13_3784, i_13_3787, i_13_3797, i_13_3816, i_13_3860, i_13_3896, i_13_3930, i_13_3931, i_13_3932, i_13_3994, i_13_3995, i_13_4219, i_13_4372, i_13_4447, i_13_4453, i_13_4454, i_13_4596, i_13_4597, i_13_4598, o_13_400);
	kernel_13_401 k_13_401(i_13_112, i_13_171, i_13_189, i_13_316, i_13_325, i_13_414, i_13_415, i_13_416, i_13_558, i_13_562, i_13_625, i_13_778, i_13_826, i_13_841, i_13_847, i_13_849, i_13_850, i_13_891, i_13_918, i_13_984, i_13_1021, i_13_1072, i_13_1081, i_13_1092, i_13_1096, i_13_1200, i_13_1224, i_13_1225, i_13_1230, i_13_1255, i_13_1278, i_13_1302, i_13_1317, i_13_1318, i_13_1480, i_13_1486, i_13_1491, i_13_1548, i_13_1549, i_13_1674, i_13_1728, i_13_1740, i_13_1746, i_13_1749, i_13_1756, i_13_1777, i_13_1854, i_13_1855, i_13_1857, i_13_1858, i_13_1954, i_13_2307, i_13_2308, i_13_2353, i_13_2395, i_13_2434, i_13_2457, i_13_2505, i_13_2539, i_13_2556, i_13_2586, i_13_2629, i_13_2691, i_13_2722, i_13_2820, i_13_2821, i_13_2850, i_13_2875, i_13_3000, i_13_3008, i_13_3064, i_13_3092, i_13_3118, i_13_3153, i_13_3163, i_13_3168, i_13_3234, i_13_3244, i_13_3267, i_13_3304, i_13_3429, i_13_3432, i_13_3484, i_13_3519, i_13_3537, i_13_3538, i_13_3574, i_13_3575, i_13_3781, i_13_3852, i_13_3906, i_13_3907, i_13_3909, i_13_4018, i_13_4366, i_13_4374, i_13_4375, i_13_4378, i_13_4393, i_13_4519, o_13_401);
	kernel_13_402 k_13_402(i_13_113, i_13_204, i_13_273, i_13_276, i_13_277, i_13_278, i_13_319, i_13_328, i_13_340, i_13_366, i_13_368, i_13_391, i_13_394, i_13_447, i_13_457, i_13_492, i_13_565, i_13_637, i_13_643, i_13_744, i_13_745, i_13_746, i_13_845, i_13_871, i_13_948, i_13_978, i_13_979, i_13_1023, i_13_1070, i_13_1086, i_13_1087, i_13_1088, i_13_1096, i_13_1141, i_13_1349, i_13_1465, i_13_1519, i_13_1623, i_13_1625, i_13_1815, i_13_1816, i_13_1943, i_13_1950, i_13_1951, i_13_2022, i_13_2060, i_13_2266, i_13_2347, i_13_2433, i_13_2437, i_13_2464, i_13_2480, i_13_2613, i_13_2677, i_13_2715, i_13_2716, i_13_2787, i_13_2788, i_13_2912, i_13_2921, i_13_2987, i_13_3003, i_13_3010, i_13_3068, i_13_3112, i_13_3127, i_13_3146, i_13_3166, i_13_3220, i_13_3229, i_13_3238, i_13_3417, i_13_3419, i_13_3451, i_13_3524, i_13_3568, i_13_3607, i_13_3658, i_13_3687, i_13_3688, i_13_3742, i_13_4001, i_13_4049, i_13_4093, i_13_4104, i_13_4120, i_13_4173, i_13_4237, i_13_4273, i_13_4297, i_13_4327, i_13_4333, i_13_4343, i_13_4399, i_13_4417, i_13_4495, i_13_4522, i_13_4533, i_13_4544, i_13_4578, o_13_402);
	kernel_13_403 k_13_403(i_13_33, i_13_34, i_13_61, i_13_70, i_13_121, i_13_136, i_13_159, i_13_160, i_13_166, i_13_226, i_13_319, i_13_385, i_13_386, i_13_414, i_13_448, i_13_456, i_13_457, i_13_492, i_13_515, i_13_565, i_13_629, i_13_646, i_13_717, i_13_735, i_13_745, i_13_938, i_13_983, i_13_985, i_13_1023, i_13_1066, i_13_1096, i_13_1116, i_13_1132, i_13_1182, i_13_1208, i_13_1216, i_13_1217, i_13_1266, i_13_1275, i_13_1302, i_13_1304, i_13_1348, i_13_1380, i_13_1489, i_13_1521, i_13_1525, i_13_1605, i_13_1743, i_13_1774, i_13_1792, i_13_1793, i_13_1808, i_13_1816, i_13_1967, i_13_2056, i_13_2123, i_13_2209, i_13_2244, i_13_2248, i_13_2281, i_13_2364, i_13_2407, i_13_2705, i_13_2749, i_13_2851, i_13_2859, i_13_2876, i_13_3022, i_13_3034, i_13_3036, i_13_3094, i_13_3095, i_13_3101, i_13_3207, i_13_3265, i_13_3354, i_13_3391, i_13_3551, i_13_3564, i_13_3759, i_13_3768, i_13_3769, i_13_3820, i_13_3821, i_13_3847, i_13_3848, i_13_3859, i_13_3954, i_13_3985, i_13_3989, i_13_4076, i_13_4084, i_13_4090, i_13_4238, i_13_4273, i_13_4299, i_13_4328, i_13_4399, i_13_4400, i_13_4594, o_13_403);
	kernel_13_404 k_13_404(i_13_22, i_13_59, i_13_91, i_13_92, i_13_139, i_13_215, i_13_316, i_13_317, i_13_418, i_13_419, i_13_456, i_13_484, i_13_550, i_13_554, i_13_607, i_13_671, i_13_727, i_13_793, i_13_843, i_13_847, i_13_851, i_13_860, i_13_986, i_13_1018, i_13_1019, i_13_1083, i_13_1122, i_13_1129, i_13_1210, i_13_1226, i_13_1256, i_13_1300, i_13_1301, i_13_1306, i_13_1345, i_13_1361, i_13_1486, i_13_1487, i_13_1550, i_13_1599, i_13_1631, i_13_1644, i_13_1721, i_13_1733, i_13_1763, i_13_1769, i_13_1813, i_13_1855, i_13_1858, i_13_1859, i_13_1911, i_13_2016, i_13_2028, i_13_2173, i_13_2179, i_13_2207, i_13_2290, i_13_2296, i_13_2422, i_13_2450, i_13_2593, i_13_2615, i_13_2679, i_13_2697, i_13_2748, i_13_2857, i_13_2981, i_13_3007, i_13_3008, i_13_3010, i_13_3037, i_13_3110, i_13_3217, i_13_3389, i_13_3404, i_13_3428, i_13_3481, i_13_3530, i_13_3563, i_13_3570, i_13_3574, i_13_3767, i_13_3853, i_13_3854, i_13_3874, i_13_3889, i_13_3890, i_13_3893, i_13_3939, i_13_4016, i_13_4018, i_13_4055, i_13_4163, i_13_4232, i_13_4258, i_13_4369, i_13_4370, i_13_4376, i_13_4565, i_13_4568, o_13_404);
	kernel_13_405 k_13_405(i_13_52, i_13_78, i_13_94, i_13_118, i_13_124, i_13_142, i_13_159, i_13_241, i_13_251, i_13_259, i_13_327, i_13_485, i_13_526, i_13_552, i_13_553, i_13_555, i_13_584, i_13_591, i_13_619, i_13_620, i_13_680, i_13_713, i_13_732, i_13_742, i_13_796, i_13_943, i_13_944, i_13_961, i_13_980, i_13_1030, i_13_1078, i_13_1079, i_13_1249, i_13_1313, i_13_1366, i_13_1403, i_13_1472, i_13_1502, i_13_1552, i_13_1553, i_13_1636, i_13_1637, i_13_1661, i_13_1817, i_13_1951, i_13_1995, i_13_2118, i_13_2211, i_13_2238, i_13_2321, i_13_2402, i_13_2451, i_13_2455, i_13_2476, i_13_2555, i_13_2570, i_13_2596, i_13_2726, i_13_2788, i_13_2789, i_13_2861, i_13_2888, i_13_2959, i_13_3026, i_13_3037, i_13_3063, i_13_3207, i_13_3219, i_13_3373, i_13_3374, i_13_3452, i_13_3464, i_13_3554, i_13_3571, i_13_3572, i_13_3581, i_13_3650, i_13_3651, i_13_3689, i_13_3738, i_13_3894, i_13_3904, i_13_3905, i_13_3938, i_13_4057, i_13_4091, i_13_4118, i_13_4125, i_13_4254, i_13_4306, i_13_4318, i_13_4345, i_13_4364, i_13_4391, i_13_4414, i_13_4415, i_13_4526, i_13_4534, i_13_4556, i_13_4604, o_13_405);
	kernel_13_406 k_13_406(i_13_76, i_13_111, i_13_129, i_13_179, i_13_266, i_13_277, i_13_282, i_13_283, i_13_302, i_13_358, i_13_366, i_13_471, i_13_472, i_13_509, i_13_510, i_13_545, i_13_591, i_13_598, i_13_664, i_13_726, i_13_799, i_13_832, i_13_854, i_13_862, i_13_894, i_13_1073, i_13_1203, i_13_1212, i_13_1213, i_13_1307, i_13_1308, i_13_1310, i_13_1390, i_13_1505, i_13_1623, i_13_1682, i_13_1698, i_13_1730, i_13_2020, i_13_2023, i_13_2024, i_13_2059, i_13_2285, i_13_2297, i_13_2299, i_13_2321, i_13_2445, i_13_2455, i_13_2456, i_13_2464, i_13_2554, i_13_2650, i_13_2715, i_13_2716, i_13_2722, i_13_2884, i_13_2897, i_13_2959, i_13_3046, i_13_3062, i_13_3076, i_13_3093, i_13_3145, i_13_3253, i_13_3327, i_13_3329, i_13_3374, i_13_3380, i_13_3388, i_13_3417, i_13_3418, i_13_3490, i_13_3550, i_13_3597, i_13_3599, i_13_3635, i_13_3659, i_13_3764, i_13_3846, i_13_3910, i_13_3923, i_13_3990, i_13_4119, i_13_4164, i_13_4192, i_13_4216, i_13_4255, i_13_4265, i_13_4332, i_13_4333, i_13_4334, i_13_4367, i_13_4369, i_13_4431, i_13_4433, i_13_4454, i_13_4461, i_13_4472, i_13_4510, i_13_4512, o_13_406);
	kernel_13_407 k_13_407(i_13_19, i_13_64, i_13_111, i_13_165, i_13_166, i_13_237, i_13_325, i_13_336, i_13_450, i_13_495, i_13_585, i_13_615, i_13_639, i_13_756, i_13_811, i_13_813, i_13_855, i_13_882, i_13_984, i_13_1062, i_13_1063, i_13_1216, i_13_1219, i_13_1251, i_13_1395, i_13_1458, i_13_1503, i_13_1513, i_13_1524, i_13_1608, i_13_1714, i_13_1848, i_13_1927, i_13_1990, i_13_2052, i_13_2053, i_13_2107, i_13_2116, i_13_2124, i_13_2127, i_13_2133, i_13_2134, i_13_2136, i_13_2145, i_13_2172, i_13_2233, i_13_2259, i_13_2260, i_13_2277, i_13_2278, i_13_2340, i_13_2364, i_13_2403, i_13_2404, i_13_2520, i_13_2614, i_13_2709, i_13_2713, i_13_2745, i_13_2757, i_13_2781, i_13_2934, i_13_2937, i_13_2938, i_13_3010, i_13_3024, i_13_3127, i_13_3339, i_13_3376, i_13_3394, i_13_3612, i_13_3627, i_13_3628, i_13_3639, i_13_3663, i_13_3703, i_13_3708, i_13_3738, i_13_3739, i_13_3793, i_13_3817, i_13_3891, i_13_4017, i_13_4059, i_13_4060, i_13_4062, i_13_4086, i_13_4102, i_13_4267, i_13_4276, i_13_4303, i_13_4315, i_13_4329, i_13_4338, i_13_4377, i_13_4392, i_13_4446, i_13_4447, i_13_4530, i_13_4568, o_13_407);
	kernel_13_408 k_13_408(i_13_64, i_13_97, i_13_121, i_13_131, i_13_158, i_13_208, i_13_236, i_13_245, i_13_251, i_13_415, i_13_416, i_13_463, i_13_464, i_13_571, i_13_589, i_13_596, i_13_761, i_13_829, i_13_1073, i_13_1129, i_13_1207, i_13_1211, i_13_1318, i_13_1346, i_13_1361, i_13_1466, i_13_1510, i_13_1511, i_13_1522, i_13_1550, i_13_1570, i_13_1604, i_13_1640, i_13_1696, i_13_1697, i_13_1700, i_13_1751, i_13_1840, i_13_1847, i_13_1853, i_13_1874, i_13_1928, i_13_1958, i_13_1964, i_13_1994, i_13_2057, i_13_2101, i_13_2102, i_13_2143, i_13_2200, i_13_2201, i_13_2209, i_13_2297, i_13_2315, i_13_2434, i_13_2444, i_13_2551, i_13_2612, i_13_2798, i_13_2881, i_13_2936, i_13_2939, i_13_3056, i_13_3113, i_13_3143, i_13_3208, i_13_3242, i_13_3254, i_13_3347, i_13_3370, i_13_3388, i_13_3458, i_13_3551, i_13_3596, i_13_3610, i_13_3619, i_13_3632, i_13_3637, i_13_3638, i_13_3667, i_13_3704, i_13_3766, i_13_3844, i_13_3857, i_13_3916, i_13_3935, i_13_4009, i_13_4019, i_13_4037, i_13_4045, i_13_4105, i_13_4208, i_13_4214, i_13_4330, i_13_4378, i_13_4430, i_13_4451, i_13_4510, i_13_4559, i_13_4582, o_13_408);
	kernel_13_409 k_13_409(i_13_20, i_13_91, i_13_92, i_13_100, i_13_155, i_13_166, i_13_169, i_13_174, i_13_203, i_13_280, i_13_284, i_13_316, i_13_381, i_13_490, i_13_517, i_13_571, i_13_607, i_13_697, i_13_931, i_13_1021, i_13_1063, i_13_1064, i_13_1066, i_13_1092, i_13_1093, i_13_1219, i_13_1268, i_13_1324, i_13_1364, i_13_1440, i_13_1496, i_13_1528, i_13_1570, i_13_1747, i_13_1810, i_13_1829, i_13_1848, i_13_1849, i_13_1870, i_13_1885, i_13_1909, i_13_2053, i_13_2107, i_13_2108, i_13_2116, i_13_2117, i_13_2233, i_13_2234, i_13_2260, i_13_2274, i_13_2332, i_13_2333, i_13_2396, i_13_2404, i_13_2406, i_13_2443, i_13_2597, i_13_2624, i_13_2701, i_13_2790, i_13_2793, i_13_2848, i_13_2853, i_13_2872, i_13_2935, i_13_2938, i_13_2980, i_13_3007, i_13_3089, i_13_3109, i_13_3143, i_13_3205, i_13_3339, i_13_3352, i_13_3397, i_13_3541, i_13_3603, i_13_3733, i_13_3739, i_13_3742, i_13_3764, i_13_3766, i_13_3816, i_13_3817, i_13_3818, i_13_3870, i_13_4012, i_13_4016, i_13_4018, i_13_4059, i_13_4060, i_13_4061, i_13_4062, i_13_4063, i_13_4143, i_13_4259, i_13_4267, i_13_4315, i_13_4352, i_13_4567, o_13_409);
	kernel_13_410 k_13_410(i_13_18, i_13_34, i_13_45, i_13_67, i_13_70, i_13_94, i_13_128, i_13_129, i_13_156, i_13_157, i_13_160, i_13_218, i_13_222, i_13_275, i_13_333, i_13_385, i_13_409, i_13_473, i_13_490, i_13_493, i_13_615, i_13_643, i_13_644, i_13_737, i_13_738, i_13_741, i_13_742, i_13_745, i_13_829, i_13_841, i_13_934, i_13_950, i_13_956, i_13_1120, i_13_1211, i_13_1263, i_13_1300, i_13_1302, i_13_1395, i_13_1447, i_13_1522, i_13_1570, i_13_1605, i_13_1720, i_13_1760, i_13_1815, i_13_1847, i_13_1903, i_13_1939, i_13_2002, i_13_2007, i_13_2021, i_13_2101, i_13_2142, i_13_2154, i_13_2193, i_13_2235, i_13_2242, i_13_2297, i_13_2397, i_13_2584, i_13_2620, i_13_2676, i_13_2695, i_13_2781, i_13_2891, i_13_2998, i_13_3033, i_13_3213, i_13_3217, i_13_3240, i_13_3241, i_13_3242, i_13_3265, i_13_3531, i_13_3599, i_13_3618, i_13_3636, i_13_3637, i_13_3692, i_13_3702, i_13_3723, i_13_3766, i_13_3843, i_13_3846, i_13_3847, i_13_3876, i_13_3892, i_13_3915, i_13_3982, i_13_3985, i_13_4081, i_13_4117, i_13_4214, i_13_4273, i_13_4281, i_13_4327, i_13_4352, i_13_4461, i_13_4509, o_13_410);
	kernel_13_411 k_13_411(i_13_112, i_13_119, i_13_124, i_13_125, i_13_142, i_13_197, i_13_208, i_13_241, i_13_277, i_13_319, i_13_337, i_13_377, i_13_416, i_13_454, i_13_562, i_13_565, i_13_646, i_13_665, i_13_727, i_13_733, i_13_857, i_13_931, i_13_943, i_13_953, i_13_1019, i_13_1085, i_13_1225, i_13_1301, i_13_1302, i_13_1345, i_13_1375, i_13_1486, i_13_1487, i_13_1529, i_13_1627, i_13_1631, i_13_1726, i_13_1768, i_13_1787, i_13_1844, i_13_2015, i_13_2206, i_13_2212, i_13_2237, i_13_2438, i_13_2546, i_13_2618, i_13_2653, i_13_2680, i_13_2825, i_13_2917, i_13_2918, i_13_2920, i_13_3011, i_13_3020, i_13_3040, i_13_3113, i_13_3161, i_13_3167, i_13_3170, i_13_3212, i_13_3215, i_13_3217, i_13_3218, i_13_3238, i_13_3261, i_13_3328, i_13_3391, i_13_3421, i_13_3422, i_13_3463, i_13_3535, i_13_3536, i_13_3553, i_13_3644, i_13_3688, i_13_3689, i_13_3700, i_13_3781, i_13_3799, i_13_3821, i_13_3850, i_13_3872, i_13_3877, i_13_3878, i_13_3890, i_13_3898, i_13_3907, i_13_3983, i_13_3991, i_13_4012, i_13_4066, i_13_4067, i_13_4090, i_13_4270, i_13_4346, i_13_4534, i_13_4535, i_13_4543, i_13_4594, o_13_411);
	kernel_13_412 k_13_412(i_13_70, i_13_174, i_13_326, i_13_355, i_13_409, i_13_522, i_13_527, i_13_561, i_13_661, i_13_663, i_13_762, i_13_796, i_13_822, i_13_826, i_13_850, i_13_851, i_13_853, i_13_887, i_13_940, i_13_952, i_13_1020, i_13_1023, i_13_1075, i_13_1077, i_13_1186, i_13_1224, i_13_1227, i_13_1228, i_13_1230, i_13_1255, i_13_1275, i_13_1279, i_13_1303, i_13_1312, i_13_1317, i_13_1321, i_13_1345, i_13_1498, i_13_1551, i_13_1552, i_13_1570, i_13_1770, i_13_1780, i_13_1798, i_13_1854, i_13_1858, i_13_1860, i_13_1956, i_13_1957, i_13_2056, i_13_2110, i_13_2265, i_13_2281, i_13_2366, i_13_2452, i_13_2454, i_13_2460, i_13_2473, i_13_2505, i_13_2539, i_13_2541, i_13_2613, i_13_2622, i_13_2647, i_13_3031, i_13_3100, i_13_3120, i_13_3170, i_13_3172, i_13_3273, i_13_3381, i_13_3427, i_13_3429, i_13_3460, i_13_3468, i_13_3483, i_13_3503, i_13_3505, i_13_3541, i_13_3559, i_13_3570, i_13_3651, i_13_3729, i_13_3783, i_13_3822, i_13_3829, i_13_3856, i_13_3896, i_13_3910, i_13_3911, i_13_4252, i_13_4254, i_13_4256, i_13_4261, i_13_4377, i_13_4396, i_13_4415, i_13_4579, i_13_4597, i_13_4606, o_13_412);
	kernel_13_413 k_13_413(i_13_78, i_13_79, i_13_103, i_13_157, i_13_158, i_13_185, i_13_219, i_13_374, i_13_379, i_13_515, i_13_533, i_13_536, i_13_550, i_13_551, i_13_644, i_13_648, i_13_652, i_13_653, i_13_676, i_13_685, i_13_689, i_13_823, i_13_833, i_13_839, i_13_842, i_13_1074, i_13_1104, i_13_1122, i_13_1145, i_13_1327, i_13_1514, i_13_1515, i_13_1516, i_13_1517, i_13_1632, i_13_1657, i_13_1675, i_13_1677, i_13_1678, i_13_1692, i_13_1739, i_13_1747, i_13_1752, i_13_1776, i_13_1792, i_13_1909, i_13_1912, i_13_1999, i_13_2002, i_13_2017, i_13_2025, i_13_2047, i_13_2101, i_13_2467, i_13_2468, i_13_2507, i_13_2512, i_13_2542, i_13_2547, i_13_2557, i_13_2570, i_13_2622, i_13_2722, i_13_2737, i_13_2740, i_13_2766, i_13_2850, i_13_2854, i_13_2898, i_13_2908, i_13_2917, i_13_2956, i_13_3052, i_13_3088, i_13_3235, i_13_3367, i_13_3377, i_13_3476, i_13_3486, i_13_3487, i_13_3523, i_13_3604, i_13_3727, i_13_3857, i_13_3862, i_13_3863, i_13_3925, i_13_3988, i_13_4123, i_13_4124, i_13_4160, i_13_4187, i_13_4188, i_13_4260, i_13_4512, i_13_4581, i_13_4591, i_13_4596, i_13_4600, i_13_4601, o_13_413);
	kernel_13_414 k_13_414(i_13_1, i_13_45, i_13_46, i_13_67, i_13_171, i_13_172, i_13_234, i_13_351, i_13_352, i_13_408, i_13_450, i_13_472, i_13_505, i_13_508, i_13_511, i_13_567, i_13_648, i_13_657, i_13_661, i_13_673, i_13_735, i_13_850, i_13_936, i_13_937, i_13_1071, i_13_1128, i_13_1129, i_13_1211, i_13_1243, i_13_1266, i_13_1272, i_13_1314, i_13_1326, i_13_1410, i_13_1422, i_13_1434, i_13_1480, i_13_1642, i_13_1663, i_13_1692, i_13_1729, i_13_1764, i_13_1786, i_13_1795, i_13_1915, i_13_1939, i_13_1944, i_13_1999, i_13_2019, i_13_2020, i_13_2026, i_13_2097, i_13_2176, i_13_2196, i_13_2299, i_13_2340, i_13_2448, i_13_2469, i_13_2470, i_13_2592, i_13_2637, i_13_2701, i_13_2704, i_13_3027, i_13_3028, i_13_3111, i_13_3112, i_13_3126, i_13_3127, i_13_3132, i_13_3261, i_13_3367, i_13_3418, i_13_3474, i_13_3478, i_13_3480, i_13_3481, i_13_3483, i_13_3484, i_13_3531, i_13_3546, i_13_3573, i_13_3574, i_13_3577, i_13_3726, i_13_3780, i_13_3781, i_13_3819, i_13_3897, i_13_3898, i_13_4015, i_13_4161, i_13_4230, i_13_4293, i_13_4321, i_13_4375, i_13_4521, i_13_4561, i_13_4563, i_13_4603, o_13_414);
	kernel_13_415 k_13_415(i_13_162, i_13_174, i_13_201, i_13_363, i_13_412, i_13_468, i_13_604, i_13_657, i_13_658, i_13_660, i_13_661, i_13_667, i_13_694, i_13_822, i_13_828, i_13_829, i_13_831, i_13_853, i_13_946, i_13_954, i_13_955, i_13_984, i_13_1071, i_13_1075, i_13_1098, i_13_1224, i_13_1225, i_13_1269, i_13_1270, i_13_1305, i_13_1423, i_13_1435, i_13_1497, i_13_1503, i_13_1522, i_13_1534, i_13_1548, i_13_1620, i_13_1657, i_13_1722, i_13_1729, i_13_1764, i_13_1767, i_13_1791, i_13_1837, i_13_2019, i_13_2020, i_13_2142, i_13_2172, i_13_2296, i_13_2340, i_13_2365, i_13_2394, i_13_2430, i_13_2431, i_13_2448, i_13_2550, i_13_2647, i_13_2691, i_13_2721, i_13_2880, i_13_2881, i_13_2907, i_13_3000, i_13_3001, i_13_3060, i_13_3231, i_13_3324, i_13_3370, i_13_3456, i_13_3478, i_13_3483, i_13_3484, i_13_3486, i_13_3546, i_13_3547, i_13_3613, i_13_3619, i_13_3636, i_13_3637, i_13_3753, i_13_3843, i_13_3853, i_13_3910, i_13_3982, i_13_4063, i_13_4123, i_13_4161, i_13_4162, i_13_4251, i_13_4315, i_13_4329, i_13_4339, i_13_4378, i_13_4429, i_13_4449, i_13_4458, i_13_4509, i_13_4510, i_13_4600, o_13_415);
	kernel_13_416 k_13_416(i_13_33, i_13_40, i_13_93, i_13_96, i_13_105, i_13_106, i_13_159, i_13_185, i_13_268, i_13_286, i_13_318, i_13_321, i_13_338, i_13_372, i_13_569, i_13_699, i_13_700, i_13_744, i_13_816, i_13_817, i_13_843, i_13_931, i_13_984, i_13_985, i_13_1069, i_13_1122, i_13_1210, i_13_1308, i_13_1407, i_13_1429, i_13_1446, i_13_1481, i_13_1499, i_13_1518, i_13_1645, i_13_1652, i_13_1730, i_13_1733, i_13_1752, i_13_1753, i_13_1787, i_13_1813, i_13_1851, i_13_1933, i_13_1992, i_13_1995, i_13_2017, i_13_2058, i_13_2122, i_13_2139, i_13_2172, i_13_2266, i_13_2409, i_13_2410, i_13_2459, i_13_2472, i_13_2545, i_13_2617, i_13_2679, i_13_2680, i_13_2741, i_13_2787, i_13_2940, i_13_2981, i_13_2985, i_13_3022, i_13_3210, i_13_3211, i_13_3345, i_13_3371, i_13_3381, i_13_3390, i_13_3399, i_13_3400, i_13_3422, i_13_3449, i_13_3451, i_13_3488, i_13_3489, i_13_3521, i_13_3535, i_13_3702, i_13_3720, i_13_3764, i_13_3791, i_13_3911, i_13_3983, i_13_4047, i_13_4066, i_13_4083, i_13_4084, i_13_4191, i_13_4295, i_13_4350, i_13_4353, i_13_4395, i_13_4396, i_13_4416, i_13_4451, i_13_4538, o_13_416);
	kernel_13_417 k_13_417(i_13_76, i_13_205, i_13_258, i_13_286, i_13_309, i_13_340, i_13_411, i_13_519, i_13_561, i_13_586, i_13_607, i_13_618, i_13_619, i_13_627, i_13_640, i_13_661, i_13_663, i_13_672, i_13_757, i_13_771, i_13_799, i_13_856, i_13_1021, i_13_1111, i_13_1147, i_13_1278, i_13_1279, i_13_1303, i_13_1329, i_13_1330, i_13_1429, i_13_1572, i_13_1596, i_13_1633, i_13_1659, i_13_1734, i_13_1735, i_13_1744, i_13_1767, i_13_1834, i_13_1843, i_13_1891, i_13_1932, i_13_1959, i_13_2019, i_13_2022, i_13_2023, i_13_2134, i_13_2211, i_13_2248, i_13_2260, i_13_2452, i_13_2454, i_13_2455, i_13_2469, i_13_2610, i_13_2707, i_13_2715, i_13_2742, i_13_2743, i_13_2746, i_13_2787, i_13_2886, i_13_2922, i_13_2958, i_13_3031, i_13_3075, i_13_3076, i_13_3102, i_13_3315, i_13_3448, i_13_3486, i_13_3489, i_13_3490, i_13_3519, i_13_3553, i_13_3570, i_13_3603, i_13_3822, i_13_3865, i_13_3901, i_13_4021, i_13_4119, i_13_4161, i_13_4164, i_13_4165, i_13_4179, i_13_4189, i_13_4191, i_13_4255, i_13_4293, i_13_4332, i_13_4333, i_13_4362, i_13_4374, i_13_4516, i_13_4600, i_13_4602, i_13_4605, i_13_4606, o_13_417);
	kernel_13_418 k_13_418(i_13_64, i_13_76, i_13_77, i_13_103, i_13_121, i_13_173, i_13_190, i_13_284, i_13_374, i_13_382, i_13_385, i_13_415, i_13_463, i_13_493, i_13_524, i_13_527, i_13_571, i_13_581, i_13_589, i_13_598, i_13_599, i_13_686, i_13_694, i_13_695, i_13_698, i_13_824, i_13_1207, i_13_1208, i_13_1211, i_13_1307, i_13_1309, i_13_1310, i_13_1343, i_13_1385, i_13_1403, i_13_1508, i_13_1516, i_13_1550, i_13_1594, i_13_1595, i_13_1597, i_13_1610, i_13_1685, i_13_1883, i_13_1886, i_13_1928, i_13_1931, i_13_1939, i_13_1945, i_13_2000, i_13_2002, i_13_2003, i_13_2125, i_13_2189, i_13_2201, i_13_2209, i_13_2239, i_13_2302, i_13_2449, i_13_2549, i_13_2657, i_13_2675, i_13_2719, i_13_2720, i_13_2824, i_13_2857, i_13_2858, i_13_2969, i_13_3010, i_13_3031, i_13_3062, i_13_3208, i_13_3217, i_13_3374, i_13_3400, i_13_3562, i_13_3563, i_13_3650, i_13_3667, i_13_3670, i_13_3727, i_13_3728, i_13_3731, i_13_3893, i_13_3916, i_13_3982, i_13_4015, i_13_4016, i_13_4019, i_13_4259, i_13_4261, i_13_4262, i_13_4303, i_13_4396, i_13_4397, i_13_4417, i_13_4447, i_13_4454, i_13_4540, i_13_4556, o_13_418);
	kernel_13_419 k_13_419(i_13_121, i_13_171, i_13_175, i_13_202, i_13_324, i_13_325, i_13_414, i_13_415, i_13_432, i_13_558, i_13_566, i_13_568, i_13_822, i_13_823, i_13_868, i_13_891, i_13_1020, i_13_1071, i_13_1072, i_13_1092, i_13_1224, i_13_1225, i_13_1227, i_13_1251, i_13_1255, i_13_1278, i_13_1314, i_13_1317, i_13_1380, i_13_1414, i_13_1469, i_13_1511, i_13_1534, i_13_1540, i_13_1548, i_13_1549, i_13_1602, i_13_1668, i_13_1767, i_13_1775, i_13_1809, i_13_1854, i_13_1855, i_13_1881, i_13_1885, i_13_2171, i_13_2244, i_13_2405, i_13_2448, i_13_2457, i_13_2458, i_13_2539, i_13_2560, i_13_2566, i_13_2610, i_13_2629, i_13_2659, i_13_2883, i_13_2919, i_13_3007, i_13_3091, i_13_3168, i_13_3176, i_13_3236, i_13_3261, i_13_3307, i_13_3322, i_13_3415, i_13_3429, i_13_3456, i_13_3457, i_13_3459, i_13_3531, i_13_3537, i_13_3538, i_13_3540, i_13_3573, i_13_3726, i_13_3766, i_13_3784, i_13_3817, i_13_3855, i_13_3907, i_13_3909, i_13_3983, i_13_3988, i_13_4014, i_13_4015, i_13_4096, i_13_4248, i_13_4304, i_13_4338, i_13_4351, i_13_4374, i_13_4375, i_13_4378, i_13_4440, i_13_4447, i_13_4554, i_13_4557, o_13_419);
	kernel_13_420 k_13_420(i_13_0, i_13_45, i_13_46, i_13_63, i_13_64, i_13_66, i_13_121, i_13_183, i_13_234, i_13_255, i_13_256, i_13_310, i_13_414, i_13_415, i_13_444, i_13_468, i_13_469, i_13_489, i_13_490, i_13_586, i_13_603, i_13_612, i_13_613, i_13_666, i_13_685, i_13_694, i_13_695, i_13_760, i_13_839, i_13_928, i_13_945, i_13_1073, i_13_1101, i_13_1116, i_13_1129, i_13_1269, i_13_1270, i_13_1342, i_13_1422, i_13_1494, i_13_1506, i_13_1549, i_13_1596, i_13_1597, i_13_1603, i_13_1641, i_13_1669, i_13_1751, i_13_1777, i_13_1795, i_13_1926, i_13_1927, i_13_1930, i_13_1944, i_13_1998, i_13_1999, i_13_2070, i_13_2299, i_13_2377, i_13_2460, i_13_2505, i_13_2547, i_13_2676, i_13_2721, i_13_2722, i_13_2749, i_13_2880, i_13_2881, i_13_3091, i_13_3127, i_13_3261, i_13_3334, i_13_3366, i_13_3414, i_13_3415, i_13_3546, i_13_3547, i_13_3550, i_13_3610, i_13_3636, i_13_3637, i_13_3638, i_13_3699, i_13_3765, i_13_3766, i_13_3767, i_13_3781, i_13_3784, i_13_3793, i_13_3897, i_13_3937, i_13_3990, i_13_4036, i_13_4042, i_13_4080, i_13_4248, i_13_4257, i_13_4293, i_13_4294, i_13_4347, o_13_420);
	kernel_13_421 k_13_421(i_13_76, i_13_184, i_13_187, i_13_188, i_13_193, i_13_322, i_13_382, i_13_509, i_13_567, i_13_571, i_13_572, i_13_575, i_13_628, i_13_647, i_13_658, i_13_689, i_13_692, i_13_818, i_13_879, i_13_898, i_13_959, i_13_995, i_13_1020, i_13_1075, i_13_1098, i_13_1121, i_13_1123, i_13_1124, i_13_1143, i_13_1166, i_13_1224, i_13_1228, i_13_1232, i_13_1277, i_13_1346, i_13_1408, i_13_1411, i_13_1484, i_13_1516, i_13_1519, i_13_1645, i_13_1671, i_13_1678, i_13_1728, i_13_1729, i_13_1751, i_13_1754, i_13_1771, i_13_1804, i_13_1805, i_13_1807, i_13_1808, i_13_1858, i_13_1859, i_13_1862, i_13_2123, i_13_2136, i_13_2195, i_13_2267, i_13_2357, i_13_2473, i_13_2474, i_13_2624, i_13_2679, i_13_2681, i_13_2723, i_13_2823, i_13_2825, i_13_2857, i_13_2942, i_13_2983, i_13_2986, i_13_2987, i_13_3031, i_13_3032, i_13_3064, i_13_3074, i_13_3208, i_13_3209, i_13_3235, i_13_3265, i_13_3293, i_13_3347, i_13_3382, i_13_3401, i_13_3427, i_13_3506, i_13_3526, i_13_3681, i_13_3824, i_13_3861, i_13_3911, i_13_3913, i_13_4338, i_13_4396, i_13_4514, i_13_4540, i_13_4567, i_13_4598, i_13_4607, o_13_421);
	kernel_13_422 k_13_422(i_13_37, i_13_38, i_13_51, i_13_76, i_13_77, i_13_371, i_13_382, i_13_518, i_13_603, i_13_625, i_13_660, i_13_661, i_13_663, i_13_771, i_13_792, i_13_794, i_13_825, i_13_861, i_13_910, i_13_942, i_13_983, i_13_1018, i_13_1066, i_13_1077, i_13_1082, i_13_1120, i_13_1227, i_13_1284, i_13_1397, i_13_1425, i_13_1428, i_13_1429, i_13_1433, i_13_1571, i_13_1605, i_13_1631, i_13_1659, i_13_1681, i_13_1695, i_13_1744, i_13_1776, i_13_1777, i_13_1919, i_13_2027, i_13_2137, i_13_2189, i_13_2197, i_13_2209, i_13_2263, i_13_2297, i_13_2407, i_13_2451, i_13_2454, i_13_2553, i_13_2614, i_13_2662, i_13_2765, i_13_2821, i_13_3011, i_13_3037, i_13_3049, i_13_3135, i_13_3217, i_13_3322, i_13_3345, i_13_3377, i_13_3389, i_13_3397, i_13_3418, i_13_3461, i_13_3489, i_13_3490, i_13_3504, i_13_3505, i_13_3508, i_13_3567, i_13_3568, i_13_3570, i_13_3612, i_13_3618, i_13_3638, i_13_3651, i_13_3739, i_13_3740, i_13_3741, i_13_3742, i_13_3866, i_13_3891, i_13_3894, i_13_3895, i_13_4054, i_13_4088, i_13_4233, i_13_4254, i_13_4282, i_13_4356, i_13_4366, i_13_4368, i_13_4369, i_13_4603, o_13_422);
	kernel_13_423 k_13_423(i_13_38, i_13_193, i_13_209, i_13_274, i_13_284, i_13_287, i_13_310, i_13_317, i_13_382, i_13_525, i_13_528, i_13_529, i_13_561, i_13_679, i_13_682, i_13_826, i_13_852, i_13_863, i_13_914, i_13_979, i_13_1021, i_13_1022, i_13_1212, i_13_1227, i_13_1311, i_13_1312, i_13_1317, i_13_1327, i_13_1363, i_13_1429, i_13_1528, i_13_1565, i_13_1678, i_13_1726, i_13_1740, i_13_1780, i_13_1781, i_13_1871, i_13_1885, i_13_1886, i_13_1888, i_13_1960, i_13_2005, i_13_2108, i_13_2136, i_13_2146, i_13_2173, i_13_2261, i_13_2267, i_13_2302, i_13_2350, i_13_2394, i_13_2420, i_13_2462, i_13_2464, i_13_2470, i_13_2561, i_13_2653, i_13_2676, i_13_2740, i_13_2904, i_13_2962, i_13_3005, i_13_3012, i_13_3058, i_13_3100, i_13_3128, i_13_3130, i_13_3146, i_13_3197, i_13_3199, i_13_3262, i_13_3352, i_13_3509, i_13_3526, i_13_3541, i_13_3613, i_13_3614, i_13_3649, i_13_3709, i_13_3729, i_13_3730, i_13_3731, i_13_3733, i_13_3769, i_13_3854, i_13_3895, i_13_3913, i_13_4017, i_13_4057, i_13_4126, i_13_4255, i_13_4263, i_13_4264, i_13_4399, i_13_4432, i_13_4513, i_13_4557, i_13_4567, i_13_4597, o_13_423);
	kernel_13_424 k_13_424(i_13_52, i_13_68, i_13_71, i_13_140, i_13_143, i_13_177, i_13_230, i_13_309, i_13_364, i_13_539, i_13_608, i_13_610, i_13_646, i_13_647, i_13_652, i_13_674, i_13_689, i_13_764, i_13_851, i_13_887, i_13_935, i_13_938, i_13_995, i_13_1117, i_13_1123, i_13_1124, i_13_1133, i_13_1145, i_13_1270, i_13_1277, i_13_1286, i_13_1342, i_13_1364, i_13_1403, i_13_1445, i_13_1472, i_13_1511, i_13_1660, i_13_1733, i_13_1735, i_13_1736, i_13_1768, i_13_1796, i_13_1798, i_13_1799, i_13_1809, i_13_1833, i_13_1920, i_13_1944, i_13_2052, i_13_2059, i_13_2115, i_13_2134, i_13_2265, i_13_2403, i_13_2406, i_13_2429, i_13_2462, i_13_2555, i_13_2679, i_13_2694, i_13_2725, i_13_2851, i_13_2852, i_13_2885, i_13_2983, i_13_3044, i_13_3050, i_13_3157, i_13_3208, i_13_3265, i_13_3339, i_13_3356, i_13_3371, i_13_3438, i_13_3451, i_13_3522, i_13_3532, i_13_3568, i_13_3569, i_13_3611, i_13_3653, i_13_3743, i_13_3787, i_13_3896, i_13_3913, i_13_3914, i_13_3927, i_13_3930, i_13_3931, i_13_3932, i_13_4040, i_13_4063, i_13_4190, i_13_4261, i_13_4279, i_13_4297, i_13_4298, i_13_4597, i_13_4598, o_13_424);
	kernel_13_425 k_13_425(i_13_28, i_13_31, i_13_67, i_13_136, i_13_157, i_13_184, i_13_193, i_13_206, i_13_266, i_13_316, i_13_335, i_13_338, i_13_373, i_13_381, i_13_383, i_13_459, i_13_543, i_13_581, i_13_590, i_13_715, i_13_742, i_13_746, i_13_795, i_13_813, i_13_870, i_13_1075, i_13_1120, i_13_1134, i_13_1216, i_13_1282, i_13_1300, i_13_1301, i_13_1327, i_13_1345, i_13_1400, i_13_1408, i_13_1444, i_13_1489, i_13_1495, i_13_1603, i_13_1633, i_13_1678, i_13_1717, i_13_1718, i_13_1811, i_13_1813, i_13_1831, i_13_1858, i_13_1993, i_13_1997, i_13_2056, i_13_2191, i_13_2208, i_13_2399, i_13_2480, i_13_2539, i_13_2540, i_13_2575, i_13_2632, i_13_2719, i_13_2721, i_13_2723, i_13_2857, i_13_2858, i_13_2860, i_13_2916, i_13_2970, i_13_2998, i_13_3016, i_13_3019, i_13_3061, i_13_3232, i_13_3235, i_13_3439, i_13_3441, i_13_3490, i_13_3615, i_13_3616, i_13_3619, i_13_3631, i_13_3666, i_13_3683, i_13_3685, i_13_3700, i_13_3727, i_13_3766, i_13_3844, i_13_3892, i_13_3921, i_13_3974, i_13_4055, i_13_4184, i_13_4186, i_13_4235, i_13_4369, i_13_4378, i_13_4395, i_13_4396, i_13_4397, i_13_4521, o_13_425);
	kernel_13_426 k_13_426(i_13_32, i_13_36, i_13_179, i_13_184, i_13_279, i_13_286, i_13_315, i_13_319, i_13_320, i_13_337, i_13_454, i_13_553, i_13_592, i_13_645, i_13_646, i_13_647, i_13_655, i_13_670, i_13_679, i_13_680, i_13_684, i_13_691, i_13_692, i_13_835, i_13_844, i_13_898, i_13_952, i_13_1116, i_13_1121, i_13_1123, i_13_1124, i_13_1260, i_13_1262, i_13_1267, i_13_1274, i_13_1301, i_13_1519, i_13_1532, i_13_1553, i_13_1597, i_13_1643, i_13_1743, i_13_1813, i_13_1854, i_13_2058, i_13_2059, i_13_2104, i_13_2133, i_13_2210, i_13_2284, i_13_2466, i_13_2617, i_13_2677, i_13_2678, i_13_2708, i_13_2756, i_13_2781, i_13_2845, i_13_3012, i_13_3113, i_13_3145, i_13_3217, i_13_3218, i_13_3322, i_13_3379, i_13_3383, i_13_3401, i_13_3412, i_13_3418, i_13_3476, i_13_3533, i_13_3535, i_13_3538, i_13_3574, i_13_3598, i_13_3701, i_13_3724, i_13_3735, i_13_3739, i_13_3769, i_13_3770, i_13_3867, i_13_3892, i_13_3928, i_13_3935, i_13_3992, i_13_4021, i_13_4022, i_13_4032, i_13_4077, i_13_4081, i_13_4085, i_13_4090, i_13_4185, i_13_4270, i_13_4534, i_13_4586, i_13_4594, i_13_4595, i_13_4598, o_13_426);
	kernel_13_427 k_13_427(i_13_44, i_13_61, i_13_76, i_13_113, i_13_184, i_13_187, i_13_231, i_13_313, i_13_314, i_13_321, i_13_382, i_13_538, i_13_556, i_13_574, i_13_643, i_13_645, i_13_646, i_13_647, i_13_687, i_13_745, i_13_840, i_13_853, i_13_897, i_13_898, i_13_956, i_13_1021, i_13_1058, i_13_1112, i_13_1120, i_13_1121, i_13_1122, i_13_1123, i_13_1135, i_13_1275, i_13_1276, i_13_1426, i_13_1472, i_13_1516, i_13_1624, i_13_1633, i_13_1642, i_13_1643, i_13_1646, i_13_1678, i_13_1680, i_13_1716, i_13_1752, i_13_1789, i_13_1790, i_13_1800, i_13_1802, i_13_1804, i_13_1807, i_13_1816, i_13_1834, i_13_1853, i_13_1858, i_13_1861, i_13_1862, i_13_2002, i_13_2005, i_13_2057, i_13_2200, i_13_2213, i_13_2266, i_13_2267, i_13_2407, i_13_2408, i_13_2452, i_13_2528, i_13_2535, i_13_2542, i_13_2617, i_13_2697, i_13_2722, i_13_2850, i_13_2851, i_13_2903, i_13_2923, i_13_2965, i_13_2981, i_13_3028, i_13_3031, i_13_3065, i_13_3156, i_13_3292, i_13_3419, i_13_3703, i_13_3931, i_13_3993, i_13_3995, i_13_4044, i_13_4189, i_13_4190, i_13_4266, i_13_4297, i_13_4312, i_13_4356, i_13_4435, i_13_4598, o_13_427);
	kernel_13_428 k_13_428(i_13_41, i_13_67, i_13_135, i_13_136, i_13_137, i_13_138, i_13_139, i_13_166, i_13_181, i_13_283, i_13_373, i_13_489, i_13_493, i_13_535, i_13_539, i_13_621, i_13_625, i_13_694, i_13_695, i_13_696, i_13_814, i_13_856, i_13_864, i_13_884, i_13_1020, i_13_1021, i_13_1092, i_13_1129, i_13_1137, i_13_1218, i_13_1232, i_13_1306, i_13_1307, i_13_1404, i_13_1428, i_13_1431, i_13_1484, i_13_1516, i_13_1742, i_13_1759, i_13_1769, i_13_1795, i_13_1849, i_13_1882, i_13_1904, i_13_1947, i_13_1954, i_13_2119, i_13_2170, i_13_2200, i_13_2310, i_13_2354, i_13_2377, i_13_2407, i_13_2410, i_13_2445, i_13_2493, i_13_2505, i_13_2542, i_13_2720, i_13_2848, i_13_2849, i_13_2854, i_13_2872, i_13_2882, i_13_2997, i_13_2998, i_13_3021, i_13_3065, i_13_3109, i_13_3110, i_13_3130, i_13_3170, i_13_3371, i_13_3381, i_13_3481, i_13_3555, i_13_3684, i_13_3703, i_13_3723, i_13_3739, i_13_3740, i_13_3766, i_13_3818, i_13_3820, i_13_3836, i_13_3910, i_13_4006, i_13_4018, i_13_4063, i_13_4078, i_13_4152, i_13_4250, i_13_4294, i_13_4295, i_13_4316, i_13_4328, i_13_4341, i_13_4567, i_13_4581, o_13_428);
	kernel_13_429 k_13_429(i_13_4, i_13_58, i_13_61, i_13_73, i_13_93, i_13_94, i_13_283, i_13_310, i_13_373, i_13_415, i_13_426, i_13_562, i_13_571, i_13_614, i_13_627, i_13_696, i_13_697, i_13_699, i_13_780, i_13_825, i_13_955, i_13_956, i_13_1006, i_13_1023, i_13_1071, i_13_1072, i_13_1098, i_13_1213, i_13_1225, i_13_1270, i_13_1301, i_13_1317, i_13_1318, i_13_1320, i_13_1380, i_13_1383, i_13_1428, i_13_1464, i_13_1479, i_13_1482, i_13_1483, i_13_1707, i_13_1721, i_13_1740, i_13_1759, i_13_1775, i_13_1795, i_13_1885, i_13_1888, i_13_1951, i_13_1957, i_13_2119, i_13_2244, i_13_2367, i_13_2407, i_13_2443, i_13_2444, i_13_2445, i_13_2446, i_13_2491, i_13_2512, i_13_2553, i_13_2554, i_13_2613, i_13_2676, i_13_2824, i_13_2857, i_13_2875, i_13_2964, i_13_2974, i_13_3093, i_13_3094, i_13_3119, i_13_3230, i_13_3235, i_13_3304, i_13_3307, i_13_3432, i_13_3479, i_13_3489, i_13_3540, i_13_3567, i_13_3580, i_13_3756, i_13_3820, i_13_3989, i_13_3991, i_13_4018, i_13_4205, i_13_4313, i_13_4315, i_13_4350, i_13_4353, i_13_4369, i_13_4378, i_13_4379, i_13_4380, i_13_4443, i_13_4498, i_13_4503, o_13_429);
	kernel_13_430 k_13_430(i_13_33, i_13_114, i_13_159, i_13_183, i_13_384, i_13_385, i_13_406, i_13_537, i_13_570, i_13_571, i_13_589, i_13_591, i_13_681, i_13_724, i_13_760, i_13_762, i_13_795, i_13_816, i_13_913, i_13_931, i_13_942, i_13_1068, i_13_1084, i_13_1086, i_13_1266, i_13_1302, i_13_1303, i_13_1390, i_13_1408, i_13_1473, i_13_1509, i_13_1716, i_13_1788, i_13_1789, i_13_1803, i_13_1807, i_13_1815, i_13_1816, i_13_1951, i_13_1992, i_13_1995, i_13_1996, i_13_2001, i_13_2002, i_13_2122, i_13_2208, i_13_2226, i_13_2266, i_13_2424, i_13_2455, i_13_2472, i_13_2535, i_13_2541, i_13_2560, i_13_2577, i_13_2632, i_13_2790, i_13_2847, i_13_2919, i_13_2941, i_13_3003, i_13_3022, i_13_3031, i_13_3102, i_13_3126, i_13_3129, i_13_3147, i_13_3163, i_13_3265, i_13_3274, i_13_3328, i_13_3346, i_13_3381, i_13_3391, i_13_3399, i_13_3441, i_13_3453, i_13_3522, i_13_3535, i_13_3615, i_13_3624, i_13_3661, i_13_3702, i_13_3796, i_13_3846, i_13_3873, i_13_3928, i_13_3993, i_13_4057, i_13_4119, i_13_4165, i_13_4207, i_13_4236, i_13_4272, i_13_4273, i_13_4341, i_13_4399, i_13_4416, i_13_4417, i_13_4540, o_13_430);
	kernel_13_431 k_13_431(i_13_37, i_13_93, i_13_102, i_13_138, i_13_139, i_13_174, i_13_229, i_13_267, i_13_373, i_13_505, i_13_549, i_13_550, i_13_603, i_13_604, i_13_657, i_13_660, i_13_661, i_13_663, i_13_669, i_13_675, i_13_676, i_13_855, i_13_1023, i_13_1072, i_13_1144, i_13_1219, i_13_1494, i_13_1515, i_13_1516, i_13_1521, i_13_1629, i_13_1630, i_13_1656, i_13_1711, i_13_1827, i_13_1828, i_13_1858, i_13_1881, i_13_1884, i_13_2001, i_13_2002, i_13_2016, i_13_2019, i_13_2020, i_13_2169, i_13_2340, i_13_2341, i_13_2362, i_13_2397, i_13_2398, i_13_2422, i_13_2448, i_13_2467, i_13_2497, i_13_2511, i_13_2611, i_13_2614, i_13_2718, i_13_2935, i_13_2982, i_13_3006, i_13_3009, i_13_3105, i_13_3108, i_13_3133, i_13_3159, i_13_3234, i_13_3385, i_13_3415, i_13_3475, i_13_3522, i_13_3639, i_13_3640, i_13_3738, i_13_3762, i_13_3763, i_13_3843, i_13_3861, i_13_3862, i_13_3889, i_13_3987, i_13_4077, i_13_4116, i_13_4159, i_13_4180, i_13_4186, i_13_4213, i_13_4248, i_13_4257, i_13_4320, i_13_4365, i_13_4366, i_13_4429, i_13_4521, i_13_4564, i_13_4566, i_13_4567, i_13_4590, i_13_4599, i_13_4600, o_13_431);
	kernel_13_432 k_13_432(i_13_49, i_13_75, i_13_76, i_13_94, i_13_133, i_13_139, i_13_183, i_13_187, i_13_192, i_13_193, i_13_195, i_13_207, i_13_321, i_13_526, i_13_542, i_13_570, i_13_574, i_13_612, i_13_663, i_13_668, i_13_697, i_13_714, i_13_798, i_13_831, i_13_847, i_13_853, i_13_854, i_13_985, i_13_988, i_13_1069, i_13_1149, i_13_1222, i_13_1230, i_13_1231, i_13_1321, i_13_1407, i_13_1408, i_13_1410, i_13_1521, i_13_1537, i_13_1548, i_13_1678, i_13_1732, i_13_1771, i_13_1804, i_13_1827, i_13_1834, i_13_1857, i_13_1860, i_13_1861, i_13_1885, i_13_2002, i_13_2100, i_13_2142, i_13_2145, i_13_2203, i_13_2299, i_13_2402, i_13_2422, i_13_2473, i_13_2680, i_13_2856, i_13_2857, i_13_2982, i_13_3000, i_13_3009, i_13_3064, i_13_3112, i_13_3159, i_13_3207, i_13_3208, i_13_3210, i_13_3212, i_13_3244, i_13_3409, i_13_3439, i_13_3442, i_13_3487, i_13_3531, i_13_3558, i_13_3667, i_13_3685, i_13_3730, i_13_3756, i_13_3763, i_13_3765, i_13_3979, i_13_3982, i_13_3984, i_13_4084, i_13_4357, i_13_4396, i_13_4432, i_13_4504, i_13_4512, i_13_4565, i_13_4566, i_13_4567, i_13_4569, i_13_4587, o_13_432);
	kernel_13_433 k_13_433(i_13_18, i_13_36, i_13_90, i_13_94, i_13_139, i_13_407, i_13_446, i_13_572, i_13_580, i_13_697, i_13_732, i_13_737, i_13_796, i_13_797, i_13_799, i_13_800, i_13_838, i_13_844, i_13_855, i_13_862, i_13_949, i_13_950, i_13_979, i_13_1030, i_13_1120, i_13_1196, i_13_1227, i_13_1303, i_13_1427, i_13_1445, i_13_1489, i_13_1492, i_13_1498, i_13_1499, i_13_1633, i_13_1732, i_13_1792, i_13_1854, i_13_1867, i_13_1996, i_13_2003, i_13_2005, i_13_2056, i_13_2208, i_13_2209, i_13_2272, i_13_2321, i_13_2357, i_13_2365, i_13_2425, i_13_2428, i_13_2434, i_13_2436, i_13_2437, i_13_2446, i_13_2461, i_13_2464, i_13_2465, i_13_2542, i_13_2544, i_13_2551, i_13_2614, i_13_2740, i_13_2749, i_13_2758, i_13_2919, i_13_2963, i_13_3001, i_13_3051, i_13_3059, i_13_3148, i_13_3163, i_13_3289, i_13_3424, i_13_3425, i_13_3476, i_13_3523, i_13_3531, i_13_3532, i_13_3535, i_13_3617, i_13_3726, i_13_3730, i_13_3733, i_13_3871, i_13_3873, i_13_3874, i_13_3877, i_13_3906, i_13_3910, i_13_4006, i_13_4036, i_13_4155, i_13_4189, i_13_4202, i_13_4236, i_13_4254, i_13_4450, i_13_4561, i_13_4603, o_13_433);
	kernel_13_434 k_13_434(i_13_94, i_13_141, i_13_142, i_13_168, i_13_240, i_13_258, i_13_264, i_13_310, i_13_322, i_13_339, i_13_340, i_13_373, i_13_430, i_13_526, i_13_553, i_13_582, i_13_598, i_13_607, i_13_618, i_13_619, i_13_717, i_13_727, i_13_780, i_13_799, i_13_979, i_13_1077, i_13_1078, i_13_1231, i_13_1276, i_13_1311, i_13_1402, i_13_1435, i_13_1470, i_13_1471, i_13_1483, i_13_1597, i_13_1626, i_13_1635, i_13_1650, i_13_1699, i_13_1725, i_13_1734, i_13_1776, i_13_1780, i_13_1783, i_13_1785, i_13_1816, i_13_1849, i_13_1960, i_13_1996, i_13_2059, i_13_2149, i_13_2293, i_13_2319, i_13_2347, i_13_2434, i_13_2649, i_13_2679, i_13_2742, i_13_2751, i_13_2787, i_13_2859, i_13_2886, i_13_2937, i_13_3013, i_13_3039, i_13_3291, i_13_3292, i_13_3414, i_13_3415, i_13_3444, i_13_3481, i_13_3525, i_13_3526, i_13_3532, i_13_3534, i_13_3541, i_13_3550, i_13_3642, i_13_3643, i_13_3687, i_13_3688, i_13_3706, i_13_3756, i_13_3757, i_13_4278, i_13_4318, i_13_4327, i_13_4335, i_13_4354, i_13_4360, i_13_4363, i_13_4389, i_13_4390, i_13_4395, i_13_4417, i_13_4432, i_13_4513, i_13_4525, i_13_4533, o_13_434);
	kernel_13_435 k_13_435(i_13_34, i_13_67, i_13_71, i_13_95, i_13_136, i_13_137, i_13_185, i_13_200, i_13_448, i_13_449, i_13_517, i_13_535, i_13_536, i_13_538, i_13_605, i_13_613, i_13_614, i_13_644, i_13_682, i_13_686, i_13_703, i_13_934, i_13_1077, i_13_1087, i_13_1105, i_13_1123, i_13_1196, i_13_1215, i_13_1216, i_13_1218, i_13_1232, i_13_1274, i_13_1276, i_13_1283, i_13_1402, i_13_1403, i_13_1441, i_13_1598, i_13_1606, i_13_1643, i_13_1674, i_13_1736, i_13_1767, i_13_1796, i_13_1798, i_13_1799, i_13_1858, i_13_1889, i_13_1931, i_13_1934, i_13_1945, i_13_1998, i_13_2075, i_13_2123, i_13_2174, i_13_2176, i_13_2267, i_13_2421, i_13_2422, i_13_2425, i_13_2426, i_13_2567, i_13_2648, i_13_2917, i_13_3031, i_13_3032, i_13_3064, i_13_3103, i_13_3104, i_13_3128, i_13_3130, i_13_3212, i_13_3216, i_13_3239, i_13_3265, i_13_3367, i_13_3368, i_13_3406, i_13_3418, i_13_3419, i_13_3439, i_13_3456, i_13_3638, i_13_3699, i_13_3745, i_13_3787, i_13_3876, i_13_3899, i_13_3931, i_13_3932, i_13_3994, i_13_3995, i_13_4015, i_13_4042, i_13_4046, i_13_4066, i_13_4084, i_13_4085, i_13_4297, i_13_4606, o_13_435);
	kernel_13_436 k_13_436(i_13_47, i_13_73, i_13_74, i_13_157, i_13_166, i_13_184, i_13_229, i_13_342, i_13_357, i_13_362, i_13_428, i_13_431, i_13_434, i_13_513, i_13_515, i_13_533, i_13_551, i_13_605, i_13_607, i_13_649, i_13_652, i_13_653, i_13_659, i_13_667, i_13_694, i_13_698, i_13_841, i_13_886, i_13_1110, i_13_1117, i_13_1144, i_13_1145, i_13_1207, i_13_1208, i_13_1658, i_13_1732, i_13_1742, i_13_1791, i_13_1792, i_13_1918, i_13_1920, i_13_1939, i_13_1950, i_13_1951, i_13_2017, i_13_2020, i_13_2030, i_13_2206, i_13_2209, i_13_2318, i_13_2377, i_13_2443, i_13_2452, i_13_2467, i_13_2514, i_13_2691, i_13_2785, i_13_2884, i_13_2906, i_13_2938, i_13_2939, i_13_2956, i_13_2958, i_13_3044, i_13_3101, i_13_3153, i_13_3241, i_13_3312, i_13_3313, i_13_3367, i_13_3476, i_13_3479, i_13_3488, i_13_3532, i_13_3550, i_13_3568, i_13_3569, i_13_3596, i_13_3598, i_13_3646, i_13_3739, i_13_3866, i_13_3910, i_13_4063, i_13_4158, i_13_4177, i_13_4186, i_13_4187, i_13_4190, i_13_4199, i_13_4257, i_13_4297, i_13_4306, i_13_4330, i_13_4331, i_13_4333, i_13_4448, i_13_4522, i_13_4540, i_13_4601, o_13_436);
	kernel_13_437 k_13_437(i_13_47, i_13_65, i_13_109, i_13_110, i_13_111, i_13_112, i_13_206, i_13_276, i_13_382, i_13_411, i_13_520, i_13_605, i_13_626, i_13_659, i_13_680, i_13_816, i_13_856, i_13_927, i_13_932, i_13_937, i_13_938, i_13_1054, i_13_1072, i_13_1077, i_13_1086, i_13_1096, i_13_1212, i_13_1316, i_13_1424, i_13_1481, i_13_1495, i_13_1498, i_13_1519, i_13_1626, i_13_1653, i_13_1662, i_13_1735, i_13_1742, i_13_1746, i_13_1747, i_13_2020, i_13_2023, i_13_2136, i_13_2191, i_13_2248, i_13_2263, i_13_2320, i_13_2407, i_13_2481, i_13_2500, i_13_2529, i_13_2539, i_13_2562, i_13_2595, i_13_2677, i_13_2723, i_13_2884, i_13_2913, i_13_2935, i_13_3047, i_13_3089, i_13_3095, i_13_3100, i_13_3102, i_13_3103, i_13_3315, i_13_3326, i_13_3339, i_13_3355, i_13_3451, i_13_3452, i_13_3478, i_13_3550, i_13_3564, i_13_3570, i_13_3602, i_13_3606, i_13_3661, i_13_3685, i_13_3688, i_13_3730, i_13_3741, i_13_3859, i_13_4119, i_13_4159, i_13_4160, i_13_4162, i_13_4165, i_13_4173, i_13_4181, i_13_4184, i_13_4325, i_13_4332, i_13_4334, i_13_4335, i_13_4365, i_13_4366, i_13_4370, i_13_4372, i_13_4544, o_13_437);
	kernel_13_438 k_13_438(i_13_29, i_13_45, i_13_107, i_13_271, i_13_300, i_13_352, i_13_374, i_13_422, i_13_451, i_13_559, i_13_561, i_13_562, i_13_569, i_13_604, i_13_605, i_13_607, i_13_608, i_13_610, i_13_658, i_13_659, i_13_661, i_13_662, i_13_670, i_13_680, i_13_829, i_13_832, i_13_833, i_13_882, i_13_885, i_13_886, i_13_946, i_13_1075, i_13_1084, i_13_1226, i_13_1281, i_13_1381, i_13_1404, i_13_1405, i_13_1467, i_13_1520, i_13_1522, i_13_1535, i_13_1660, i_13_1768, i_13_1787, i_13_1802, i_13_1838, i_13_1846, i_13_1885, i_13_1897, i_13_1927, i_13_2021, i_13_2137, i_13_2170, i_13_2297, i_13_2423, i_13_2431, i_13_2435, i_13_2647, i_13_2650, i_13_2749, i_13_2880, i_13_3047, i_13_3106, i_13_3117, i_13_3311, i_13_3457, i_13_3476, i_13_3547, i_13_3638, i_13_3664, i_13_3683, i_13_3740, i_13_3844, i_13_3871, i_13_3872, i_13_3889, i_13_3910, i_13_3932, i_13_3982, i_13_4006, i_13_4096, i_13_4115, i_13_4158, i_13_4160, i_13_4162, i_13_4163, i_13_4261, i_13_4313, i_13_4315, i_13_4324, i_13_4351, i_13_4369, i_13_4429, i_13_4441, i_13_4463, i_13_4510, i_13_4537, i_13_4540, i_13_4541, o_13_438);
	kernel_13_439 k_13_439(i_13_108, i_13_112, i_13_171, i_13_282, i_13_336, i_13_594, i_13_639, i_13_739, i_13_793, i_13_819, i_13_820, i_13_847, i_13_855, i_13_856, i_13_868, i_13_894, i_13_1017, i_13_1120, i_13_1215, i_13_1224, i_13_1251, i_13_1252, i_13_1278, i_13_1279, i_13_1299, i_13_1309, i_13_1395, i_13_1422, i_13_1440, i_13_1467, i_13_1485, i_13_1486, i_13_1490, i_13_1494, i_13_1548, i_13_1549, i_13_1570, i_13_1629, i_13_1630, i_13_1693, i_13_1792, i_13_1827, i_13_1855, i_13_1857, i_13_1954, i_13_1998, i_13_1999, i_13_2044, i_13_2060, i_13_2172, i_13_2196, i_13_2377, i_13_2380, i_13_2394, i_13_2421, i_13_2422, i_13_2457, i_13_2494, i_13_2501, i_13_2529, i_13_2530, i_13_2538, i_13_2539, i_13_2542, i_13_2543, i_13_2592, i_13_2610, i_13_2712, i_13_2716, i_13_2728, i_13_2817, i_13_2902, i_13_2916, i_13_2917, i_13_2997, i_13_3025, i_13_3123, i_13_3144, i_13_3145, i_13_3168, i_13_3370, i_13_3420, i_13_3442, i_13_3465, i_13_3475, i_13_3483, i_13_3780, i_13_3870, i_13_3871, i_13_3991, i_13_4005, i_13_4006, i_13_4114, i_13_4185, i_13_4230, i_13_4248, i_13_4249, i_13_4251, i_13_4342, i_13_4374, o_13_439);
	kernel_13_440 k_13_440(i_13_52, i_13_71, i_13_76, i_13_112, i_13_113, i_13_241, i_13_251, i_13_273, i_13_278, i_13_284, i_13_341, i_13_594, i_13_619, i_13_855, i_13_878, i_13_1102, i_13_1120, i_13_1273, i_13_1309, i_13_1364, i_13_1426, i_13_1474, i_13_1525, i_13_1573, i_13_1597, i_13_1629, i_13_1633, i_13_1634, i_13_1642, i_13_1669, i_13_1741, i_13_1753, i_13_1795, i_13_1796, i_13_1816, i_13_1817, i_13_1939, i_13_2452, i_13_2455, i_13_2465, i_13_2497, i_13_2501, i_13_2561, i_13_2570, i_13_2712, i_13_2713, i_13_2715, i_13_2716, i_13_2761, i_13_2884, i_13_2920, i_13_2942, i_13_2983, i_13_3004, i_13_3010, i_13_3067, i_13_3101, i_13_3145, i_13_3148, i_13_3201, i_13_3238, i_13_3292, i_13_3310, i_13_3328, i_13_3329, i_13_3391, i_13_3406, i_13_3417, i_13_3451, i_13_3454, i_13_3455, i_13_3477, i_13_3527, i_13_3541, i_13_3599, i_13_3646, i_13_3660, i_13_3684, i_13_3687, i_13_3688, i_13_3689, i_13_3730, i_13_3832, i_13_3874, i_13_3922, i_13_3982, i_13_4021, i_13_4036, i_13_4057, i_13_4093, i_13_4157, i_13_4158, i_13_4274, i_13_4408, i_13_4409, i_13_4427, i_13_4522, i_13_4543, i_13_4558, i_13_4594, o_13_440);
	kernel_13_441 k_13_441(i_13_31, i_13_48, i_13_49, i_13_51, i_13_67, i_13_124, i_13_139, i_13_229, i_13_247, i_13_257, i_13_492, i_13_493, i_13_515, i_13_652, i_13_672, i_13_678, i_13_816, i_13_840, i_13_843, i_13_853, i_13_942, i_13_979, i_13_984, i_13_985, i_13_1191, i_13_1267, i_13_1326, i_13_1327, i_13_1329, i_13_1330, i_13_1509, i_13_1572, i_13_1681, i_13_1686, i_13_1723, i_13_1852, i_13_1908, i_13_2002, i_13_2022, i_13_2028, i_13_2148, i_13_2184, i_13_2229, i_13_2265, i_13_2277, i_13_2302, i_13_2318, i_13_2472, i_13_2506, i_13_2508, i_13_2509, i_13_2697, i_13_2698, i_13_2742, i_13_2743, i_13_2748, i_13_2751, i_13_2752, i_13_2874, i_13_2875, i_13_2958, i_13_2967, i_13_2973, i_13_3013, i_13_3058, i_13_3108, i_13_3115, i_13_3118, i_13_3144, i_13_3172, i_13_3210, i_13_3291, i_13_3315, i_13_3349, i_13_3372, i_13_3405, i_13_3418, i_13_3453, i_13_3463, i_13_3489, i_13_3490, i_13_3522, i_13_3525, i_13_3546, i_13_3552, i_13_3706, i_13_3765, i_13_3766, i_13_3769, i_13_3865, i_13_3876, i_13_3903, i_13_3994, i_13_4089, i_13_4161, i_13_4174, i_13_4318, i_13_4331, i_13_4495, i_13_4560, o_13_441);
	kernel_13_442 k_13_442(i_13_184, i_13_259, i_13_285, i_13_286, i_13_310, i_13_357, i_13_454, i_13_466, i_13_503, i_13_592, i_13_636, i_13_683, i_13_690, i_13_841, i_13_952, i_13_1111, i_13_1213, i_13_1218, i_13_1219, i_13_1261, i_13_1263, i_13_1313, i_13_1318, i_13_1347, i_13_1348, i_13_1364, i_13_1427, i_13_1447, i_13_1462, i_13_1525, i_13_1529, i_13_1561, i_13_1678, i_13_1868, i_13_1894, i_13_1933, i_13_1941, i_13_1993, i_13_2001, i_13_2002, i_13_2003, i_13_2005, i_13_2058, i_13_2059, i_13_2060, i_13_2146, i_13_2149, i_13_2236, i_13_2283, i_13_2284, i_13_2285, i_13_2299, i_13_2407, i_13_2425, i_13_2456, i_13_2554, i_13_2589, i_13_2590, i_13_2610, i_13_2653, i_13_2654, i_13_2658, i_13_2681, i_13_2743, i_13_2824, i_13_2856, i_13_2860, i_13_2906, i_13_2956, i_13_3146, i_13_3148, i_13_3220, i_13_3316, i_13_3345, i_13_3391, i_13_3392, i_13_3482, i_13_3553, i_13_3580, i_13_3598, i_13_3633, i_13_3729, i_13_3732, i_13_3734, i_13_3787, i_13_3994, i_13_4020, i_13_4114, i_13_4237, i_13_4263, i_13_4264, i_13_4310, i_13_4333, i_13_4363, i_13_4398, i_13_4399, i_13_4400, i_13_4534, i_13_4567, i_13_4598, o_13_442);
	kernel_13_443 k_13_443(i_13_62, i_13_117, i_13_134, i_13_136, i_13_174, i_13_283, i_13_333, i_13_351, i_13_489, i_13_493, i_13_599, i_13_612, i_13_617, i_13_624, i_13_828, i_13_889, i_13_1098, i_13_1099, i_13_1100, i_13_1116, i_13_1123, i_13_1128, i_13_1132, i_13_1208, i_13_1256, i_13_1394, i_13_1429, i_13_1442, i_13_1517, i_13_1521, i_13_1522, i_13_1639, i_13_1699, i_13_1745, i_13_1754, i_13_1811, i_13_1958, i_13_2111, i_13_2142, i_13_2143, i_13_2208, i_13_2295, i_13_2296, i_13_2300, i_13_2380, i_13_2402, i_13_2423, i_13_2438, i_13_2442, i_13_2464, i_13_2511, i_13_2781, i_13_2880, i_13_2986, i_13_3015, i_13_3065, i_13_3090, i_13_3094, i_13_3133, i_13_3171, i_13_3196, i_13_3241, i_13_3269, i_13_3307, i_13_3339, i_13_3366, i_13_3368, i_13_3429, i_13_3474, i_13_3537, i_13_3547, i_13_3636, i_13_3637, i_13_3685, i_13_3699, i_13_3753, i_13_3754, i_13_3765, i_13_3855, i_13_3889, i_13_3896, i_13_3910, i_13_3978, i_13_3985, i_13_4017, i_13_4018, i_13_4216, i_13_4297, i_13_4311, i_13_4312, i_13_4315, i_13_4321, i_13_4336, i_13_4394, i_13_4414, i_13_4509, i_13_4513, i_13_4514, i_13_4568, i_13_4598, o_13_443);
	kernel_13_444 k_13_444(i_13_48, i_13_49, i_13_70, i_13_107, i_13_178, i_13_411, i_13_448, i_13_535, i_13_570, i_13_610, i_13_616, i_13_645, i_13_760, i_13_762, i_13_797, i_13_933, i_13_934, i_13_939, i_13_1083, i_13_1101, i_13_1104, i_13_1131, i_13_1132, i_13_1137, i_13_1276, i_13_1285, i_13_1428, i_13_1482, i_13_1506, i_13_1509, i_13_1510, i_13_1515, i_13_1574, i_13_1626, i_13_1634, i_13_1644, i_13_1651, i_13_1716, i_13_1735, i_13_1767, i_13_1768, i_13_1770, i_13_1797, i_13_1798, i_13_1804, i_13_1841, i_13_1884, i_13_1945, i_13_1957, i_13_1995, i_13_2022, i_13_2023, i_13_2049, i_13_2122, i_13_2348, i_13_2454, i_13_2472, i_13_2473, i_13_2483, i_13_2501, i_13_2615, i_13_2679, i_13_2724, i_13_2913, i_13_2937, i_13_3031, i_13_3076, i_13_3120, i_13_3164, i_13_3263, i_13_3264, i_13_3274, i_13_3351, i_13_3389, i_13_3399, i_13_3417, i_13_3418, i_13_3455, i_13_3570, i_13_3613, i_13_3640, i_13_3651, i_13_3783, i_13_3813, i_13_3822, i_13_3823, i_13_3900, i_13_3940, i_13_3982, i_13_4084, i_13_4164, i_13_4193, i_13_4300, i_13_4308, i_13_4324, i_13_4400, i_13_4596, i_13_4597, i_13_4605, i_13_4606, o_13_444);
	kernel_13_445 k_13_445(i_13_67, i_13_68, i_13_112, i_13_120, i_13_123, i_13_175, i_13_214, i_13_242, i_13_251, i_13_259, i_13_273, i_13_277, i_13_278, i_13_283, i_13_311, i_13_376, i_13_412, i_13_454, i_13_471, i_13_521, i_13_609, i_13_620, i_13_800, i_13_841, i_13_935, i_13_980, i_13_1070, i_13_1112, i_13_1330, i_13_1331, i_13_1389, i_13_1394, i_13_1398, i_13_1410, i_13_1455, i_13_1472, i_13_1483, i_13_1512, i_13_1520, i_13_1573, i_13_1597, i_13_1598, i_13_1642, i_13_1664, i_13_1674, i_13_1731, i_13_1807, i_13_1835, i_13_1836, i_13_1945, i_13_2023, i_13_2025, i_13_2029, i_13_2149, i_13_2186, i_13_2200, i_13_2303, i_13_2433, i_13_2456, i_13_2698, i_13_2743, i_13_2744, i_13_2789, i_13_2883, i_13_2888, i_13_2937, i_13_2942, i_13_2959, i_13_2969, i_13_3043, i_13_3050, i_13_3077, i_13_3212, i_13_3238, i_13_3292, i_13_3316, i_13_3329, i_13_3381, i_13_3419, i_13_3454, i_13_3526, i_13_3533, i_13_3553, i_13_3596, i_13_3613, i_13_3689, i_13_3730, i_13_3762, i_13_3928, i_13_4066, i_13_4173, i_13_4253, i_13_4274, i_13_4363, i_13_4446, i_13_4503, i_13_4506, i_13_4517, i_13_4526, i_13_4563, o_13_445);
	kernel_13_446 k_13_446(i_13_92, i_13_95, i_13_121, i_13_122, i_13_233, i_13_280, i_13_287, i_13_443, i_13_452, i_13_517, i_13_568, i_13_569, i_13_572, i_13_576, i_13_607, i_13_608, i_13_677, i_13_712, i_13_730, i_13_734, i_13_737, i_13_841, i_13_859, i_13_886, i_13_950, i_13_961, i_13_1058, i_13_1069, i_13_1225, i_13_1229, i_13_1327, i_13_1406, i_13_1448, i_13_1625, i_13_1720, i_13_1721, i_13_1783, i_13_1784, i_13_1787, i_13_1840, i_13_1855, i_13_1921, i_13_2056, i_13_2128, i_13_2129, i_13_2173, i_13_2206, i_13_2207, i_13_2359, i_13_2410, i_13_2422, i_13_2425, i_13_2426, i_13_2429, i_13_2458, i_13_2462, i_13_2465, i_13_2564, i_13_2654, i_13_2695, i_13_2741, i_13_2844, i_13_2941, i_13_2981, i_13_3015, i_13_3106, i_13_3142, i_13_3143, i_13_3161, i_13_3163, i_13_3164, i_13_3171, i_13_3214, i_13_3287, i_13_3421, i_13_3422, i_13_3424, i_13_3425, i_13_3428, i_13_3689, i_13_3769, i_13_3871, i_13_3874, i_13_3875, i_13_3878, i_13_3916, i_13_4006, i_13_4009, i_13_4010, i_13_4011, i_13_4015, i_13_4021, i_13_4048, i_13_4049, i_13_4066, i_13_4078, i_13_4318, i_13_4351, i_13_4357, i_13_4603, o_13_446);
	kernel_13_447 k_13_447(i_13_107, i_13_114, i_13_115, i_13_118, i_13_130, i_13_170, i_13_240, i_13_250, i_13_382, i_13_383, i_13_410, i_13_454, i_13_464, i_13_526, i_13_528, i_13_598, i_13_697, i_13_799, i_13_813, i_13_897, i_13_979, i_13_1066, i_13_1067, i_13_1085, i_13_1096, i_13_1300, i_13_1345, i_13_1444, i_13_1465, i_13_1500, i_13_1528, i_13_1544, i_13_1628, i_13_1636, i_13_1750, i_13_1813, i_13_1814, i_13_1851, i_13_1852, i_13_1867, i_13_1993, i_13_2005, i_13_2006, i_13_2045, i_13_2110, i_13_2200, i_13_2236, i_13_2435, i_13_2462, i_13_2464, i_13_2544, i_13_2545, i_13_2546, i_13_2572, i_13_2617, i_13_2618, i_13_2767, i_13_2825, i_13_2858, i_13_2938, i_13_2939, i_13_2985, i_13_3001, i_13_3014, i_13_3020, i_13_3112, i_13_3127, i_13_3140, i_13_3207, i_13_3234, i_13_3256, i_13_3262, i_13_3392, i_13_3418, i_13_3467, i_13_3526, i_13_3536, i_13_3643, i_13_3705, i_13_3722, i_13_3725, i_13_3733, i_13_3742, i_13_3850, i_13_3851, i_13_3865, i_13_3923, i_13_3963, i_13_4022, i_13_4063, i_13_4089, i_13_4090, i_13_4091, i_13_4234, i_13_4270, i_13_4271, i_13_4396, i_13_4533, i_13_4561, i_13_4579, o_13_447);
	kernel_13_448 k_13_448(i_13_93, i_13_106, i_13_121, i_13_183, i_13_184, i_13_285, i_13_322, i_13_410, i_13_445, i_13_466, i_13_490, i_13_537, i_13_571, i_13_588, i_13_645, i_13_646, i_13_691, i_13_697, i_13_832, i_13_845, i_13_898, i_13_1069, i_13_1088, i_13_1120, i_13_1210, i_13_1276, i_13_1303, i_13_1321, i_13_1329, i_13_1362, i_13_1473, i_13_1474, i_13_1492, i_13_1519, i_13_1520, i_13_1555, i_13_1789, i_13_1795, i_13_1807, i_13_1885, i_13_1921, i_13_1930, i_13_1933, i_13_1934, i_13_1960, i_13_2122, i_13_2244, i_13_2309, i_13_2365, i_13_2381, i_13_2473, i_13_2506, i_13_2695, i_13_2698, i_13_2941, i_13_2942, i_13_3002, i_13_3005, i_13_3022, i_13_3023, i_13_3064, i_13_3067, i_13_3103, i_13_3119, i_13_3122, i_13_3166, i_13_3210, i_13_3211, i_13_3346, i_13_3451, i_13_3490, i_13_3526, i_13_3527, i_13_3541, i_13_3544, i_13_3561, i_13_3631, i_13_3766, i_13_3796, i_13_3804, i_13_3806, i_13_3874, i_13_3910, i_13_4021, i_13_4048, i_13_4049, i_13_4057, i_13_4084, i_13_4090, i_13_4120, i_13_4273, i_13_4274, i_13_4353, i_13_4359, i_13_4381, i_13_4399, i_13_4417, i_13_4432, i_13_4593, i_13_4597, o_13_448);
	kernel_13_449 k_13_449(i_13_41, i_13_62, i_13_74, i_13_77, i_13_137, i_13_167, i_13_227, i_13_274, i_13_337, i_13_537, i_13_571, i_13_582, i_13_641, i_13_681, i_13_689, i_13_690, i_13_694, i_13_695, i_13_697, i_13_814, i_13_820, i_13_821, i_13_824, i_13_825, i_13_887, i_13_1066, i_13_1067, i_13_1068, i_13_1211, i_13_1220, i_13_1271, i_13_1381, i_13_1388, i_13_1423, i_13_1444, i_13_1490, i_13_1594, i_13_1640, i_13_1670, i_13_1712, i_13_1793, i_13_1882, i_13_1883, i_13_1885, i_13_1886, i_13_1889, i_13_2364, i_13_2470, i_13_2549, i_13_2552, i_13_2611, i_13_2647, i_13_2651, i_13_2845, i_13_2848, i_13_2873, i_13_2885, i_13_2983, i_13_3011, i_13_3028, i_13_3109, i_13_3127, i_13_3173, i_13_3208, i_13_3269, i_13_3311, i_13_3343, i_13_3367, i_13_3376, i_13_3382, i_13_3383, i_13_3397, i_13_3415, i_13_3449, i_13_3487, i_13_3502, i_13_3503, i_13_3505, i_13_3728, i_13_3736, i_13_3740, i_13_3791, i_13_3836, i_13_3847, i_13_3871, i_13_4063, i_13_4064, i_13_4079, i_13_4187, i_13_4253, i_13_4262, i_13_4270, i_13_4295, i_13_4339, i_13_4342, i_13_4351, i_13_4441, i_13_4498, i_13_4591, i_13_4592, o_13_449);
	kernel_13_450 k_13_450(i_13_60, i_13_67, i_13_229, i_13_418, i_13_463, i_13_526, i_13_554, i_13_608, i_13_628, i_13_658, i_13_660, i_13_661, i_13_733, i_13_831, i_13_888, i_13_889, i_13_959, i_13_988, i_13_1071, i_13_1078, i_13_1087, i_13_1099, i_13_1108, i_13_1112, i_13_1120, i_13_1143, i_13_1279, i_13_1300, i_13_1330, i_13_1345, i_13_1466, i_13_1476, i_13_1516, i_13_1660, i_13_1678, i_13_1681, i_13_1744, i_13_2002, i_13_2019, i_13_2020, i_13_2021, i_13_2022, i_13_2023, i_13_2024, i_13_2077, i_13_2097, i_13_2137, i_13_2425, i_13_2453, i_13_2466, i_13_2470, i_13_2511, i_13_2614, i_13_2708, i_13_2723, i_13_2740, i_13_2741, i_13_2857, i_13_2935, i_13_2998, i_13_3004, i_13_3056, i_13_3089, i_13_3152, i_13_3272, i_13_3352, i_13_3483, i_13_3484, i_13_3490, i_13_3550, i_13_3553, i_13_3568, i_13_3621, i_13_3730, i_13_3766, i_13_3823, i_13_3861, i_13_3864, i_13_3866, i_13_3989, i_13_4027, i_13_4048, i_13_4051, i_13_4054, i_13_4160, i_13_4162, i_13_4163, i_13_4252, i_13_4253, i_13_4369, i_13_4370, i_13_4377, i_13_4388, i_13_4394, i_13_4396, i_13_4431, i_13_4517, i_13_4560, i_13_4603, i_13_4604, o_13_450);
	kernel_13_451 k_13_451(i_13_71, i_13_94, i_13_140, i_13_179, i_13_259, i_13_266, i_13_287, i_13_327, i_13_328, i_13_329, i_13_418, i_13_468, i_13_494, i_13_562, i_13_563, i_13_607, i_13_628, i_13_667, i_13_670, i_13_671, i_13_683, i_13_700, i_13_701, i_13_891, i_13_943, i_13_1021, i_13_1024, i_13_1078, i_13_1079, i_13_1314, i_13_1327, i_13_1403, i_13_1430, i_13_1444, i_13_1447, i_13_1479, i_13_1480, i_13_1484, i_13_1687, i_13_1780, i_13_1781, i_13_1789, i_13_1840, i_13_1885, i_13_1889, i_13_1906, i_13_1923, i_13_1935, i_13_2022, i_13_2059, i_13_2124, i_13_2125, i_13_2173, i_13_2197, i_13_2201, i_13_2245, i_13_2344, i_13_2384, i_13_2434, i_13_2561, i_13_2617, i_13_2618, i_13_2629, i_13_2746, i_13_2852, i_13_2875, i_13_2898, i_13_2902, i_13_2967, i_13_3043, i_13_3100, i_13_3175, i_13_3244, i_13_3381, i_13_3415, i_13_3429, i_13_3455, i_13_3460, i_13_3464, i_13_3482, i_13_3507, i_13_3535, i_13_3536, i_13_3596, i_13_3701, i_13_3731, i_13_3869, i_13_3911, i_13_3920, i_13_4100, i_13_4257, i_13_4342, i_13_4346, i_13_4350, i_13_4351, i_13_4354, i_13_4396, i_13_4451, i_13_4522, i_13_4606, o_13_451);
	kernel_13_452 k_13_452(i_13_7, i_13_33, i_13_34, i_13_35, i_13_41, i_13_109, i_13_160, i_13_188, i_13_232, i_13_374, i_13_385, i_13_447, i_13_538, i_13_572, i_13_669, i_13_763, i_13_860, i_13_942, i_13_1075, i_13_1088, i_13_1215, i_13_1218, i_13_1219, i_13_1302, i_13_1348, i_13_1398, i_13_1473, i_13_1474, i_13_1475, i_13_1492, i_13_1545, i_13_1599, i_13_1636, i_13_1724, i_13_1789, i_13_1795, i_13_1992, i_13_1995, i_13_2002, i_13_2010, i_13_2046, i_13_2194, i_13_2209, i_13_2231, i_13_2242, i_13_2364, i_13_2365, i_13_2424, i_13_2426, i_13_2455, i_13_2472, i_13_2501, i_13_2532, i_13_2679, i_13_2904, i_13_2938, i_13_2958, i_13_3003, i_13_3004, i_13_3022, i_13_3023, i_13_3028, i_13_3066, i_13_3067, i_13_3112, i_13_3148, i_13_3163, i_13_3207, i_13_3210, i_13_3229, i_13_3234, i_13_3289, i_13_3308, i_13_3346, i_13_3382, i_13_3390, i_13_3423, i_13_3426, i_13_3490, i_13_3544, i_13_3580, i_13_3639, i_13_3648, i_13_3702, i_13_3796, i_13_3847, i_13_3873, i_13_3874, i_13_4008, i_13_4009, i_13_4035, i_13_4057, i_13_4120, i_13_4208, i_13_4354, i_13_4355, i_13_4399, i_13_4417, i_13_4418, i_13_4603, o_13_452);
	kernel_13_453 k_13_453(i_13_94, i_13_103, i_13_140, i_13_166, i_13_431, i_13_536, i_13_574, i_13_644, i_13_647, i_13_668, i_13_686, i_13_691, i_13_694, i_13_697, i_13_698, i_13_700, i_13_707, i_13_823, i_13_827, i_13_977, i_13_1033, i_13_1079, i_13_1115, i_13_1118, i_13_1121, i_13_1124, i_13_1138, i_13_1249, i_13_1277, i_13_1318, i_13_1319, i_13_1333, i_13_1388, i_13_1391, i_13_1447, i_13_1462, i_13_1465, i_13_1468, i_13_1469, i_13_1483, i_13_1484, i_13_1534, i_13_1586, i_13_1597, i_13_1711, i_13_1778, i_13_1781, i_13_1828, i_13_1849, i_13_1850, i_13_1886, i_13_1888, i_13_1889, i_13_1945, i_13_2102, i_13_2150, i_13_2206, i_13_2425, i_13_2567, i_13_2650, i_13_2651, i_13_2654, i_13_2689, i_13_2848, i_13_2849, i_13_2853, i_13_2875, i_13_2876, i_13_2888, i_13_3089, i_13_3217, i_13_3235, i_13_3244, i_13_3245, i_13_3299, i_13_3356, i_13_3398, i_13_3406, i_13_3448, i_13_3449, i_13_3501, i_13_3506, i_13_3526, i_13_3785, i_13_3794, i_13_3847, i_13_3854, i_13_3863, i_13_3982, i_13_3995, i_13_4090, i_13_4100, i_13_4187, i_13_4189, i_13_4190, i_13_4310, i_13_4364, i_13_4391, i_13_4481, i_13_4598, o_13_453);
	kernel_13_454 k_13_454(i_13_44, i_13_49, i_13_56, i_13_70, i_13_78, i_13_172, i_13_176, i_13_177, i_13_282, i_13_317, i_13_321, i_13_447, i_13_448, i_13_457, i_13_461, i_13_525, i_13_555, i_13_568, i_13_645, i_13_651, i_13_670, i_13_673, i_13_679, i_13_681, i_13_682, i_13_688, i_13_740, i_13_757, i_13_994, i_13_1104, i_13_1150, i_13_1275, i_13_1276, i_13_1401, i_13_1402, i_13_1426, i_13_1510, i_13_1514, i_13_1548, i_13_1567, i_13_1599, i_13_1633, i_13_1645, i_13_1663, i_13_1725, i_13_1734, i_13_1798, i_13_1920, i_13_1945, i_13_1946, i_13_1948, i_13_1996, i_13_2029, i_13_2032, i_13_2191, i_13_2263, i_13_2265, i_13_2266, i_13_2407, i_13_2461, i_13_2472, i_13_2545, i_13_2587, i_13_2677, i_13_2680, i_13_2695, i_13_2697, i_13_2742, i_13_2748, i_13_2901, i_13_2902, i_13_2905, i_13_2922, i_13_2923, i_13_2940, i_13_2981, i_13_3030, i_13_3111, i_13_3269, i_13_3273, i_13_3367, i_13_3418, i_13_3525, i_13_3561, i_13_3592, i_13_3651, i_13_3730, i_13_3732, i_13_3787, i_13_3928, i_13_3940, i_13_3992, i_13_3993, i_13_3994, i_13_4053, i_13_4251, i_13_4308, i_13_4323, i_13_4566, i_13_4603, o_13_454);
	kernel_13_455 k_13_455(i_13_2, i_13_156, i_13_164, i_13_166, i_13_191, i_13_241, i_13_269, i_13_278, i_13_287, i_13_314, i_13_340, i_13_358, i_13_385, i_13_386, i_13_466, i_13_470, i_13_592, i_13_593, i_13_745, i_13_746, i_13_768, i_13_823, i_13_824, i_13_827, i_13_851, i_13_916, i_13_947, i_13_952, i_13_985, i_13_1111, i_13_1120, i_13_1303, i_13_1304, i_13_1348, i_13_1435, i_13_1439, i_13_1447, i_13_1499, i_13_1501, i_13_1516, i_13_1541, i_13_1573, i_13_1574, i_13_1634, i_13_1682, i_13_1817, i_13_1867, i_13_1951, i_13_1952, i_13_1996, i_13_2033, i_13_2059, i_13_2060, i_13_2114, i_13_2123, i_13_2141, i_13_2284, i_13_2285, i_13_2401, i_13_2410, i_13_2411, i_13_2561, i_13_2570, i_13_2582, i_13_2590, i_13_2591, i_13_2617, i_13_2662, i_13_2720, i_13_2771, i_13_2824, i_13_2825, i_13_3064, i_13_3157, i_13_3221, i_13_3238, i_13_3240, i_13_3346, i_13_3347, i_13_3374, i_13_3419, i_13_3598, i_13_3599, i_13_3618, i_13_3623, i_13_3628, i_13_3634, i_13_3731, i_13_3733, i_13_3838, i_13_3923, i_13_3928, i_13_4048, i_13_4058, i_13_4237, i_13_4273, i_13_4274, i_13_4336, i_13_4400, i_13_4454, o_13_455);
	kernel_13_456 k_13_456(i_13_39, i_13_40, i_13_48, i_13_49, i_13_68, i_13_70, i_13_159, i_13_259, i_13_277, i_13_351, i_13_411, i_13_453, i_13_520, i_13_535, i_13_628, i_13_673, i_13_760, i_13_834, i_13_900, i_13_934, i_13_939, i_13_1023, i_13_1104, i_13_1105, i_13_1150, i_13_1231, i_13_1330, i_13_1349, i_13_1363, i_13_1399, i_13_1402, i_13_1521, i_13_1596, i_13_1626, i_13_1644, i_13_1663, i_13_1668, i_13_1735, i_13_1780, i_13_1798, i_13_1884, i_13_1892, i_13_1894, i_13_1947, i_13_1948, i_13_2029, i_13_2058, i_13_2121, i_13_2148, i_13_2184, i_13_2228, i_13_2265, i_13_2299, i_13_2380, i_13_2399, i_13_2400, i_13_2436, i_13_2472, i_13_2517, i_13_2553, i_13_2571, i_13_2595, i_13_2614, i_13_2724, i_13_2742, i_13_2743, i_13_2874, i_13_2912, i_13_2915, i_13_2968, i_13_3030, i_13_3031, i_13_3111, i_13_3112, i_13_3135, i_13_3315, i_13_3355, i_13_3370, i_13_3399, i_13_3481, i_13_3489, i_13_3534, i_13_3739, i_13_3765, i_13_3767, i_13_3838, i_13_3842, i_13_3892, i_13_3900, i_13_3930, i_13_4002, i_13_4022, i_13_4055, i_13_4164, i_13_4174, i_13_4233, i_13_4254, i_13_4362, i_13_4478, i_13_4606, o_13_456);
	kernel_13_457 k_13_457(i_13_51, i_13_52, i_13_97, i_13_106, i_13_159, i_13_196, i_13_286, i_13_340, i_13_385, i_13_467, i_13_574, i_13_592, i_13_625, i_13_688, i_13_700, i_13_745, i_13_817, i_13_948, i_13_962, i_13_985, i_13_1068, i_13_1069, i_13_1123, i_13_1150, i_13_1210, i_13_1258, i_13_1281, i_13_1308, i_13_1330, i_13_1574, i_13_1715, i_13_1780, i_13_1795, i_13_1806, i_13_1807, i_13_1808, i_13_1851, i_13_1852, i_13_1876, i_13_1932, i_13_1997, i_13_2002, i_13_2058, i_13_2059, i_13_2121, i_13_2123, i_13_2174, i_13_2194, i_13_2238, i_13_2266, i_13_2283, i_13_2284, i_13_2293, i_13_2343, i_13_2410, i_13_2429, i_13_2473, i_13_2498, i_13_2536, i_13_2573, i_13_2617, i_13_2752, i_13_2914, i_13_2920, i_13_2941, i_13_2986, i_13_3022, i_13_3023, i_13_3028, i_13_3109, i_13_3210, i_13_3211, i_13_3303, i_13_3346, i_13_3351, i_13_3391, i_13_3399, i_13_3401, i_13_3451, i_13_3504, i_13_3525, i_13_3526, i_13_3766, i_13_3850, i_13_3909, i_13_3911, i_13_4021, i_13_4047, i_13_4048, i_13_4049, i_13_4066, i_13_4084, i_13_4184, i_13_4234, i_13_4297, i_13_4308, i_13_4309, i_13_4318, i_13_4345, i_13_4346, o_13_457);
	kernel_13_458 k_13_458(i_13_136, i_13_138, i_13_139, i_13_172, i_13_229, i_13_257, i_13_308, i_13_370, i_13_409, i_13_512, i_13_535, i_13_554, i_13_568, i_13_657, i_13_661, i_13_675, i_13_676, i_13_697, i_13_793, i_13_842, i_13_851, i_13_937, i_13_981, i_13_983, i_13_985, i_13_986, i_13_1066, i_13_1119, i_13_1134, i_13_1202, i_13_1219, i_13_1274, i_13_1324, i_13_1327, i_13_1328, i_13_1526, i_13_1629, i_13_1828, i_13_1885, i_13_1913, i_13_2020, i_13_2107, i_13_2182, i_13_2233, i_13_2242, i_13_2296, i_13_2299, i_13_2347, i_13_2430, i_13_2461, i_13_2467, i_13_2469, i_13_2470, i_13_2592, i_13_2695, i_13_2848, i_13_2850, i_13_2872, i_13_2875, i_13_2914, i_13_2980, i_13_2983, i_13_3006, i_13_3010, i_13_3073, i_13_3105, i_13_3106, i_13_3108, i_13_3151, i_13_3205, i_13_3207, i_13_3212, i_13_3335, i_13_3388, i_13_3397, i_13_3406, i_13_3442, i_13_3465, i_13_3479, i_13_3547, i_13_3763, i_13_3764, i_13_3817, i_13_3820, i_13_3826, i_13_3862, i_13_3916, i_13_3979, i_13_4072, i_13_4123, i_13_4159, i_13_4163, i_13_4203, i_13_4254, i_13_4327, i_13_4554, i_13_4563, i_13_4565, i_13_4567, i_13_4600, o_13_458);
	kernel_13_459 k_13_459(i_13_59, i_13_136, i_13_137, i_13_173, i_13_203, i_13_256, i_13_284, i_13_311, i_13_334, i_13_352, i_13_518, i_13_523, i_13_613, i_13_622, i_13_626, i_13_641, i_13_644, i_13_685, i_13_686, i_13_695, i_13_824, i_13_976, i_13_1117, i_13_1118, i_13_1201, i_13_1208, i_13_1270, i_13_1271, i_13_1273, i_13_1274, i_13_1282, i_13_1315, i_13_1388, i_13_1444, i_13_1468, i_13_1469, i_13_1481, i_13_1625, i_13_1640, i_13_1643, i_13_1667, i_13_1678, i_13_1711, i_13_1712, i_13_1732, i_13_1793, i_13_1802, i_13_1882, i_13_1883, i_13_1945, i_13_1991, i_13_2044, i_13_2134, i_13_2135, i_13_2245, i_13_2314, i_13_2351, i_13_2377, i_13_2378, i_13_2380, i_13_2542, i_13_2549, i_13_2551, i_13_2567, i_13_2592, i_13_2647, i_13_2648, i_13_2651, i_13_2669, i_13_2728, i_13_2747, i_13_2750, i_13_2845, i_13_2846, i_13_2848, i_13_2849, i_13_2873, i_13_2875, i_13_2903, i_13_3199, i_13_3235, i_13_3385, i_13_3403, i_13_3430, i_13_3556, i_13_3559, i_13_3568, i_13_3791, i_13_4018, i_13_4034, i_13_4186, i_13_4187, i_13_4234, i_13_4262, i_13_4294, i_13_4295, i_13_4351, i_13_4352, i_13_4376, i_13_4495, o_13_459);
	kernel_13_460 k_13_460(i_13_40, i_13_61, i_13_79, i_13_105, i_13_115, i_13_124, i_13_169, i_13_268, i_13_269, i_13_391, i_13_465, i_13_466, i_13_509, i_13_673, i_13_689, i_13_734, i_13_813, i_13_815, i_13_816, i_13_817, i_13_935, i_13_952, i_13_1201, i_13_1210, i_13_1302, i_13_1303, i_13_1304, i_13_1331, i_13_1348, i_13_1447, i_13_1464, i_13_1554, i_13_1607, i_13_1713, i_13_1753, i_13_1789, i_13_1806, i_13_1807, i_13_1857, i_13_1858, i_13_1906, i_13_1943, i_13_1995, i_13_2114, i_13_2122, i_13_2139, i_13_2140, i_13_2141, i_13_2202, i_13_2224, i_13_2239, i_13_2247, i_13_2410, i_13_2446, i_13_2463, i_13_2496, i_13_2694, i_13_2696, i_13_2798, i_13_2823, i_13_2824, i_13_2825, i_13_2912, i_13_2920, i_13_2938, i_13_2941, i_13_2986, i_13_3022, i_13_3092, i_13_3244, i_13_3273, i_13_3346, i_13_3347, i_13_3373, i_13_3374, i_13_3391, i_13_3418, i_13_3427, i_13_3455, i_13_3505, i_13_3622, i_13_3633, i_13_3793, i_13_3824, i_13_3913, i_13_3991, i_13_3992, i_13_4046, i_13_4047, i_13_4058, i_13_4081, i_13_4162, i_13_4237, i_13_4308, i_13_4342, i_13_4344, i_13_4372, i_13_4380, i_13_4381, i_13_4526, o_13_460);
	kernel_13_461 k_13_461(i_13_28, i_13_30, i_13_64, i_13_65, i_13_74, i_13_113, i_13_122, i_13_157, i_13_266, i_13_382, i_13_441, i_13_551, i_13_651, i_13_658, i_13_659, i_13_814, i_13_815, i_13_829, i_13_887, i_13_929, i_13_940, i_13_941, i_13_1082, i_13_1119, i_13_1125, i_13_1145, i_13_1208, i_13_1307, i_13_1344, i_13_1388, i_13_1389, i_13_1404, i_13_1424, i_13_1470, i_13_1593, i_13_1597, i_13_1657, i_13_1668, i_13_1712, i_13_1730, i_13_1755, i_13_1837, i_13_1838, i_13_1929, i_13_1993, i_13_1994, i_13_2016, i_13_2137, i_13_2170, i_13_2192, i_13_2405, i_13_2468, i_13_2610, i_13_2712, i_13_2845, i_13_2846, i_13_2847, i_13_2884, i_13_2939, i_13_3028, i_13_3063, i_13_3106, i_13_3157, i_13_3204, i_13_3240, i_13_3261, i_13_3387, i_13_3487, i_13_3502, i_13_3503, i_13_3569, i_13_3577, i_13_3618, i_13_3636, i_13_3646, i_13_3648, i_13_3667, i_13_3736, i_13_3738, i_13_3767, i_13_3889, i_13_3907, i_13_3915, i_13_4054, i_13_4078, i_13_4088, i_13_4160, i_13_4162, i_13_4164, i_13_4187, i_13_4233, i_13_4276, i_13_4330, i_13_4340, i_13_4365, i_13_4430, i_13_4540, i_13_4592, i_13_4600, i_13_4601, o_13_461);
	kernel_13_462 k_13_462(i_13_49, i_13_50, i_13_138, i_13_139, i_13_231, i_13_256, i_13_268, i_13_447, i_13_492, i_13_517, i_13_537, i_13_589, i_13_615, i_13_626, i_13_643, i_13_644, i_13_645, i_13_686, i_13_688, i_13_690, i_13_699, i_13_822, i_13_897, i_13_976, i_13_1118, i_13_1120, i_13_1123, i_13_1197, i_13_1221, i_13_1273, i_13_1274, i_13_1389, i_13_1390, i_13_1392, i_13_1480, i_13_1644, i_13_1645, i_13_1649, i_13_1713, i_13_1725, i_13_1726, i_13_1735, i_13_1762, i_13_1779, i_13_1795, i_13_1796, i_13_1797, i_13_1798, i_13_1803, i_13_1831, i_13_1849, i_13_1885, i_13_1992, i_13_1994, i_13_2137, i_13_2191, i_13_2379, i_13_2616, i_13_2648, i_13_2748, i_13_2751, i_13_2757, i_13_2847, i_13_2848, i_13_2849, i_13_2851, i_13_2875, i_13_3039, i_13_3270, i_13_3368, i_13_3407, i_13_3432, i_13_3523, i_13_3534, i_13_3575, i_13_3670, i_13_3724, i_13_3730, i_13_3759, i_13_3838, i_13_3897, i_13_3930, i_13_3994, i_13_4054, i_13_4063, i_13_4099, i_13_4101, i_13_4125, i_13_4187, i_13_4189, i_13_4294, i_13_4297, i_13_4306, i_13_4341, i_13_4369, i_13_4396, i_13_4414, i_13_4449, i_13_4584, i_13_4597, o_13_462);
	kernel_13_463 k_13_463(i_13_76, i_13_105, i_13_112, i_13_184, i_13_186, i_13_193, i_13_195, i_13_327, i_13_445, i_13_510, i_13_562, i_13_573, i_13_574, i_13_579, i_13_626, i_13_646, i_13_666, i_13_697, i_13_717, i_13_780, i_13_854, i_13_861, i_13_894, i_13_949, i_13_958, i_13_994, i_13_1059, i_13_1084, i_13_1231, i_13_1258, i_13_1285, i_13_1321, i_13_1393, i_13_1407, i_13_1410, i_13_1483, i_13_1484, i_13_1488, i_13_1633, i_13_1677, i_13_1680, i_13_1690, i_13_1723, i_13_1749, i_13_1750, i_13_1752, i_13_1753, i_13_1788, i_13_1803, i_13_1804, i_13_1807, i_13_1858, i_13_1860, i_13_1861, i_13_2266, i_13_2310, i_13_2314, i_13_2519, i_13_2635, i_13_2652, i_13_2653, i_13_2673, i_13_2713, i_13_2715, i_13_2787, i_13_2850, i_13_2856, i_13_2857, i_13_2920, i_13_2983, i_13_3063, i_13_3144, i_13_3208, i_13_3309, i_13_3310, i_13_3372, i_13_3435, i_13_3451, i_13_3562, i_13_3595, i_13_3642, i_13_3685, i_13_3688, i_13_3739, i_13_3888, i_13_3909, i_13_3912, i_13_3913, i_13_3922, i_13_3938, i_13_3984, i_13_3994, i_13_4011, i_13_4012, i_13_4054, i_13_4077, i_13_4378, i_13_4443, i_13_4587, i_13_4591, o_13_463);
	kernel_13_464 k_13_464(i_13_173, i_13_325, i_13_370, i_13_414, i_13_523, i_13_568, i_13_657, i_13_658, i_13_659, i_13_660, i_13_661, i_13_662, i_13_677, i_13_685, i_13_724, i_13_812, i_13_846, i_13_847, i_13_848, i_13_850, i_13_851, i_13_858, i_13_937, i_13_1017, i_13_1018, i_13_1073, i_13_1200, i_13_1225, i_13_1228, i_13_1305, i_13_1315, i_13_1345, i_13_1396, i_13_1454, i_13_1486, i_13_1549, i_13_1607, i_13_1630, i_13_1751, i_13_1764, i_13_1854, i_13_1855, i_13_1858, i_13_1926, i_13_1948, i_13_1954, i_13_1955, i_13_2197, i_13_2297, i_13_2417, i_13_2444, i_13_2448, i_13_2449, i_13_2541, i_13_2910, i_13_3006, i_13_3007, i_13_3061, i_13_3217, i_13_3235, i_13_3305, i_13_3370, i_13_3377, i_13_3414, i_13_3456, i_13_3457, i_13_3468, i_13_3475, i_13_3483, i_13_3484, i_13_3537, i_13_3538, i_13_3542, i_13_3557, i_13_3573, i_13_3574, i_13_3575, i_13_3647, i_13_3648, i_13_3727, i_13_3780, i_13_3852, i_13_3864, i_13_3892, i_13_3909, i_13_3929, i_13_4124, i_13_4249, i_13_4253, i_13_4257, i_13_4302, i_13_4338, i_13_4368, i_13_4369, i_13_4374, i_13_4375, i_13_4376, i_13_4458, i_13_4554, i_13_4595, o_13_464);
	kernel_13_465 k_13_465(i_13_22, i_13_48, i_13_59, i_13_68, i_13_94, i_13_112, i_13_165, i_13_195, i_13_202, i_13_237, i_13_238, i_13_255, i_13_274, i_13_283, i_13_309, i_13_333, i_13_336, i_13_337, i_13_383, i_13_454, i_13_585, i_13_586, i_13_588, i_13_615, i_13_620, i_13_665, i_13_771, i_13_781, i_13_833, i_13_856, i_13_980, i_13_1265, i_13_1310, i_13_1341, i_13_1342, i_13_1471, i_13_1488, i_13_1567, i_13_1670, i_13_1767, i_13_1803, i_13_1804, i_13_1931, i_13_1990, i_13_1992, i_13_2145, i_13_2179, i_13_2209, i_13_2376, i_13_2506, i_13_2535, i_13_2569, i_13_2571, i_13_2595, i_13_2678, i_13_2898, i_13_2903, i_13_2934, i_13_3016, i_13_3027, i_13_3028, i_13_3036, i_13_3037, i_13_3040, i_13_3122, i_13_3145, i_13_3210, i_13_3216, i_13_3220, i_13_3221, i_13_3285, i_13_3289, i_13_3315, i_13_3339, i_13_3342, i_13_3344, i_13_3393, i_13_3421, i_13_3468, i_13_3523, i_13_3599, i_13_3601, i_13_3639, i_13_3640, i_13_3643, i_13_3768, i_13_3784, i_13_3889, i_13_3982, i_13_4193, i_13_4230, i_13_4231, i_13_4315, i_13_4392, i_13_4408, i_13_4446, i_13_4512, i_13_4530, i_13_4534, i_13_4594, o_13_465);
	kernel_13_466 k_13_466(i_13_20, i_13_65, i_13_121, i_13_207, i_13_208, i_13_211, i_13_265, i_13_266, i_13_373, i_13_384, i_13_414, i_13_415, i_13_423, i_13_503, i_13_521, i_13_522, i_13_664, i_13_715, i_13_746, i_13_763, i_13_764, i_13_833, i_13_849, i_13_850, i_13_852, i_13_982, i_13_1081, i_13_1084, i_13_1131, i_13_1133, i_13_1151, i_13_1200, i_13_1219, i_13_1309, i_13_1312, i_13_1397, i_13_1436, i_13_1467, i_13_1522, i_13_1549, i_13_1550, i_13_1551, i_13_1552, i_13_1599, i_13_1604, i_13_1630, i_13_1723, i_13_1732, i_13_1750, i_13_1751, i_13_1952, i_13_1999, i_13_2048, i_13_2121, i_13_2125, i_13_2295, i_13_2434, i_13_2709, i_13_2723, i_13_3087, i_13_3088, i_13_3100, i_13_3125, i_13_3163, i_13_3271, i_13_3289, i_13_3345, i_13_3346, i_13_3383, i_13_3405, i_13_3414, i_13_3423, i_13_3483, i_13_3486, i_13_3524, i_13_3537, i_13_3538, i_13_3539, i_13_3541, i_13_3542, i_13_3619, i_13_3666, i_13_3667, i_13_3726, i_13_3728, i_13_3765, i_13_3798, i_13_3843, i_13_3906, i_13_3920, i_13_3985, i_13_4038, i_13_4039, i_13_4059, i_13_4204, i_13_4256, i_13_4336, i_13_4378, i_13_4447, i_13_4523, o_13_466);
	kernel_13_467 k_13_467(i_13_56, i_13_131, i_13_166, i_13_187, i_13_202, i_13_211, i_13_284, i_13_319, i_13_355, i_13_365, i_13_392, i_13_520, i_13_521, i_13_527, i_13_545, i_13_563, i_13_589, i_13_616, i_13_652, i_13_688, i_13_833, i_13_1003, i_13_1066, i_13_1067, i_13_1069, i_13_1075, i_13_1108, i_13_1112, i_13_1129, i_13_1225, i_13_1278, i_13_1391, i_13_1454, i_13_1498, i_13_1523, i_13_1534, i_13_1598, i_13_1669, i_13_1687, i_13_1717, i_13_1723, i_13_1771, i_13_1781, i_13_1799, i_13_1930, i_13_1975, i_13_1984, i_13_1993, i_13_2023, i_13_2024, i_13_2087, i_13_2102, i_13_2137, i_13_2173, i_13_2200, i_13_2362, i_13_2363, i_13_2371, i_13_2386, i_13_2393, i_13_2425, i_13_2572, i_13_2606, i_13_2615, i_13_2618, i_13_2654, i_13_2681, i_13_2785, i_13_2815, i_13_2888, i_13_2969, i_13_2971, i_13_2974, i_13_3014, i_13_3032, i_13_3056, i_13_3181, i_13_3209, i_13_3212, i_13_3266, i_13_3487, i_13_3730, i_13_3778, i_13_3823, i_13_3901, i_13_3938, i_13_3941, i_13_4015, i_13_4031, i_13_4159, i_13_4165, i_13_4166, i_13_4225, i_13_4369, i_13_4373, i_13_4384, i_13_4451, i_13_4496, i_13_4507, i_13_4517, o_13_467);
	kernel_13_468 k_13_468(i_13_45, i_13_46, i_13_79, i_13_121, i_13_122, i_13_173, i_13_184, i_13_226, i_13_238, i_13_313, i_13_337, i_13_408, i_13_444, i_13_518, i_13_523, i_13_533, i_13_554, i_13_649, i_13_684, i_13_723, i_13_734, i_13_760, i_13_848, i_13_922, i_13_938, i_13_976, i_13_1017, i_13_1031, i_13_1071, i_13_1073, i_13_1101, i_13_1136, i_13_1148, i_13_1207, i_13_1225, i_13_1301, i_13_1306, i_13_1315, i_13_1372, i_13_1389, i_13_1427, i_13_1444, i_13_1445, i_13_1510, i_13_1549, i_13_1720, i_13_1728, i_13_1859, i_13_1945, i_13_2026, i_13_2027, i_13_2045, i_13_2126, i_13_2197, i_13_2198, i_13_2209, i_13_2262, i_13_2448, i_13_2469, i_13_2705, i_13_2763, i_13_2852, i_13_2918, i_13_3006, i_13_3007, i_13_3027, i_13_3128, i_13_3217, i_13_3218, i_13_3227, i_13_3235, i_13_3457, i_13_3458, i_13_3484, i_13_3485, i_13_3575, i_13_3781, i_13_3782, i_13_3800, i_13_3853, i_13_3915, i_13_3983, i_13_3990, i_13_4017, i_13_4080, i_13_4150, i_13_4193, i_13_4234, i_13_4249, i_13_4250, i_13_4258, i_13_4259, i_13_4262, i_13_4301, i_13_4369, i_13_4376, i_13_4447, i_13_4448, i_13_4593, i_13_4604, o_13_468);
	kernel_13_469 k_13_469(i_13_90, i_13_91, i_13_130, i_13_141, i_13_172, i_13_370, i_13_389, i_13_423, i_13_430, i_13_450, i_13_553, i_13_585, i_13_657, i_13_660, i_13_688, i_13_726, i_13_828, i_13_829, i_13_831, i_13_933, i_13_934, i_13_955, i_13_1063, i_13_1066, i_13_1075, i_13_1096, i_13_1116, i_13_1147, i_13_1224, i_13_1306, i_13_1324, i_13_1428, i_13_1471, i_13_1488, i_13_1494, i_13_1510, i_13_1552, i_13_1570, i_13_1696, i_13_1697, i_13_1726, i_13_1764, i_13_1786, i_13_1801, i_13_1846, i_13_1887, i_13_1892, i_13_1926, i_13_1927, i_13_1957, i_13_2044, i_13_2107, i_13_2119, i_13_2142, i_13_2143, i_13_2175, i_13_2265, i_13_2266, i_13_2296, i_13_2461, i_13_2877, i_13_2935, i_13_2938, i_13_3006, i_13_3016, i_13_3039, i_13_3043, i_13_3064, i_13_3225, i_13_3231, i_13_3241, i_13_3264, i_13_3274, i_13_3454, i_13_3457, i_13_3487, i_13_3523, i_13_3538, i_13_3637, i_13_3645, i_13_3742, i_13_3753, i_13_3754, i_13_3856, i_13_3916, i_13_3979, i_13_4018, i_13_4267, i_13_4268, i_13_4308, i_13_4312, i_13_4341, i_13_4368, i_13_4369, i_13_4429, i_13_4509, i_13_4510, i_13_4511, i_13_4524, i_13_4567, o_13_469);
	kernel_13_470 k_13_470(i_13_51, i_13_124, i_13_186, i_13_229, i_13_250, i_13_258, i_13_276, i_13_277, i_13_309, i_13_375, i_13_376, i_13_420, i_13_430, i_13_561, i_13_588, i_13_618, i_13_619, i_13_642, i_13_654, i_13_672, i_13_699, i_13_738, i_13_771, i_13_823, i_13_840, i_13_942, i_13_979, i_13_1065, i_13_1069, i_13_1077, i_13_1078, i_13_1218, i_13_1230, i_13_1297, i_13_1327, i_13_1329, i_13_1443, i_13_1528, i_13_1569, i_13_1572, i_13_1596, i_13_1734, i_13_1735, i_13_1834, i_13_1852, i_13_1992, i_13_2002, i_13_2107, i_13_2185, i_13_2229, i_13_2230, i_13_2302, i_13_2313, i_13_2314, i_13_2362, i_13_2454, i_13_2572, i_13_2581, i_13_2694, i_13_2697, i_13_2742, i_13_2752, i_13_2769, i_13_2886, i_13_2887, i_13_2922, i_13_2958, i_13_2967, i_13_3006, i_13_3291, i_13_3315, i_13_3372, i_13_3522, i_13_3525, i_13_3549, i_13_3552, i_13_3553, i_13_3603, i_13_3612, i_13_3687, i_13_3714, i_13_3729, i_13_3730, i_13_3733, i_13_3748, i_13_3817, i_13_3822, i_13_3885, i_13_3903, i_13_3904, i_13_4047, i_13_4089, i_13_4164, i_13_4236, i_13_4282, i_13_4332, i_13_4387, i_13_4390, i_13_4461, i_13_4603, o_13_470);
	kernel_13_471 k_13_471(i_13_49, i_13_66, i_13_133, i_13_195, i_13_327, i_13_381, i_13_483, i_13_528, i_13_529, i_13_673, i_13_717, i_13_799, i_13_842, i_13_844, i_13_861, i_13_951, i_13_1204, i_13_1222, i_13_1228, i_13_1230, i_13_1257, i_13_1258, i_13_1302, i_13_1320, i_13_1326, i_13_1384, i_13_1428, i_13_1437, i_13_1446, i_13_1491, i_13_1492, i_13_1501, i_13_1554, i_13_1555, i_13_1556, i_13_1699, i_13_1722, i_13_1795, i_13_1834, i_13_1884, i_13_1902, i_13_1930, i_13_1941, i_13_1960, i_13_2002, i_13_2005, i_13_2014, i_13_2033, i_13_2103, i_13_2128, i_13_2139, i_13_2148, i_13_2202, i_13_2203, i_13_2299, i_13_2302, i_13_2446, i_13_2535, i_13_2722, i_13_2743, i_13_2850, i_13_2937, i_13_2938, i_13_3027, i_13_3136, i_13_3174, i_13_3238, i_13_3244, i_13_3309, i_13_3310, i_13_3423, i_13_3445, i_13_3525, i_13_3543, i_13_3552, i_13_3597, i_13_3616, i_13_3706, i_13_3731, i_13_3732, i_13_3786, i_13_3805, i_13_3831, i_13_3849, i_13_3858, i_13_3859, i_13_3912, i_13_3913, i_13_3994, i_13_4011, i_13_4012, i_13_4117, i_13_4161, i_13_4254, i_13_4369, i_13_4380, i_13_4381, i_13_4443, i_13_4587, i_13_4588, o_13_471);
	kernel_13_472 k_13_472(i_13_37, i_13_135, i_13_136, i_13_140, i_13_225, i_13_279, i_13_280, i_13_563, i_13_594, i_13_640, i_13_643, i_13_670, i_13_685, i_13_714, i_13_812, i_13_891, i_13_892, i_13_1025, i_13_1075, i_13_1093, i_13_1117, i_13_1200, i_13_1213, i_13_1214, i_13_1273, i_13_1314, i_13_1384, i_13_1387, i_13_1469, i_13_1480, i_13_1481, i_13_1669, i_13_1710, i_13_1711, i_13_1757, i_13_1778, i_13_1793, i_13_1828, i_13_1855, i_13_1881, i_13_1882, i_13_1885, i_13_1886, i_13_1915, i_13_2050, i_13_2380, i_13_2443, i_13_2585, i_13_2629, i_13_2630, i_13_2647, i_13_2649, i_13_2650, i_13_2651, i_13_2653, i_13_2656, i_13_2752, i_13_2844, i_13_2845, i_13_2849, i_13_2872, i_13_2874, i_13_2983, i_13_3109, i_13_3123, i_13_3208, i_13_3287, i_13_3311, i_13_3407, i_13_3429, i_13_3430, i_13_3448, i_13_3598, i_13_3757, i_13_3761, i_13_3781, i_13_3790, i_13_3791, i_13_3793, i_13_3835, i_13_3836, i_13_3871, i_13_3901, i_13_3923, i_13_3933, i_13_4042, i_13_4043, i_13_4054, i_13_4055, i_13_4096, i_13_4114, i_13_4198, i_13_4237, i_13_4351, i_13_4369, i_13_4388, i_13_4396, i_13_4441, i_13_4519, i_13_4567, o_13_472);
	kernel_13_473 k_13_473(i_13_48, i_13_51, i_13_52, i_13_72, i_13_73, i_13_166, i_13_169, i_13_285, i_13_339, i_13_384, i_13_618, i_13_619, i_13_678, i_13_690, i_13_771, i_13_816, i_13_817, i_13_840, i_13_844, i_13_856, i_13_1021, i_13_1069, i_13_1074, i_13_1258, i_13_1300, i_13_1390, i_13_1411, i_13_1572, i_13_1573, i_13_1623, i_13_1627, i_13_1629, i_13_1635, i_13_1636, i_13_1806, i_13_1807, i_13_1950, i_13_2014, i_13_2058, i_13_2059, i_13_2266, i_13_2283, i_13_2284, i_13_2346, i_13_2353, i_13_2380, i_13_2399, i_13_2410, i_13_2472, i_13_2536, i_13_2538, i_13_2590, i_13_2617, i_13_2650, i_13_2715, i_13_2751, i_13_2752, i_13_2759, i_13_2762, i_13_2787, i_13_2903, i_13_2941, i_13_3031, i_13_3042, i_13_3043, i_13_3109, i_13_3136, i_13_3141, i_13_3144, i_13_3147, i_13_3220, i_13_3292, i_13_3372, i_13_3373, i_13_3399, i_13_3526, i_13_3721, i_13_3730, i_13_3732, i_13_3850, i_13_3891, i_13_3915, i_13_4018, i_13_4020, i_13_4021, i_13_4047, i_13_4048, i_13_4131, i_13_4132, i_13_4234, i_13_4252, i_13_4255, i_13_4263, i_13_4300, i_13_4308, i_13_4318, i_13_4339, i_13_4554, i_13_4560, i_13_4561, o_13_473);
	kernel_13_474 k_13_474(i_13_95, i_13_98, i_13_134, i_13_139, i_13_170, i_13_175, i_13_176, i_13_178, i_13_233, i_13_311, i_13_374, i_13_428, i_13_464, i_13_527, i_13_575, i_13_599, i_13_646, i_13_664, i_13_671, i_13_818, i_13_851, i_13_854, i_13_985, i_13_986, i_13_989, i_13_1024, i_13_1070, i_13_1232, i_13_1300, i_13_1309, i_13_1327, i_13_1408, i_13_1436, i_13_1571, i_13_1723, i_13_1754, i_13_1765, i_13_1805, i_13_1831, i_13_1832, i_13_1850, i_13_1852, i_13_1853, i_13_1862, i_13_1885, i_13_1921, i_13_2300, i_13_2308, i_13_2366, i_13_2408, i_13_2461, i_13_2471, i_13_2473, i_13_2510, i_13_2633, i_13_2662, i_13_2680, i_13_2698, i_13_2848, i_13_2983, i_13_2987, i_13_3001, i_13_3013, i_13_3106, i_13_3109, i_13_3110, i_13_3112, i_13_3113, i_13_3116, i_13_3137, i_13_3157, i_13_3272, i_13_3404, i_13_3410, i_13_3419, i_13_3425, i_13_3427, i_13_3481, i_13_3490, i_13_3637, i_13_3686, i_13_3769, i_13_3799, i_13_3800, i_13_3820, i_13_3821, i_13_3860, i_13_3977, i_13_4022, i_13_4064, i_13_4067, i_13_4127, i_13_4354, i_13_4378, i_13_4444, i_13_4460, i_13_4513, i_13_4567, i_13_4568, i_13_4570, o_13_474);
	kernel_13_475 k_13_475(i_13_273, i_13_283, i_13_354, i_13_355, i_13_364, i_13_469, i_13_490, i_13_598, i_13_640, i_13_651, i_13_658, i_13_660, i_13_765, i_13_767, i_13_927, i_13_928, i_13_939, i_13_940, i_13_948, i_13_1037, i_13_1071, i_13_1080, i_13_1081, i_13_1082, i_13_1098, i_13_1099, i_13_1116, i_13_1225, i_13_1227, i_13_1306, i_13_1307, i_13_1443, i_13_1486, i_13_1497, i_13_1498, i_13_1566, i_13_1567, i_13_1620, i_13_1639, i_13_1710, i_13_1719, i_13_1720, i_13_1729, i_13_1765, i_13_1774, i_13_1782, i_13_1837, i_13_1840, i_13_1846, i_13_1927, i_13_1971, i_13_2100, i_13_2205, i_13_2259, i_13_2324, i_13_2358, i_13_2424, i_13_2467, i_13_2485, i_13_2587, i_13_2673, i_13_2684, i_13_2781, i_13_2844, i_13_2845, i_13_2884, i_13_3025, i_13_3163, i_13_3258, i_13_3285, i_13_3286, i_13_3361, i_13_3388, i_13_3420, i_13_3423, i_13_3424, i_13_3457, i_13_3487, i_13_3600, i_13_3601, i_13_3619, i_13_3754, i_13_3924, i_13_3933, i_13_3988, i_13_4008, i_13_4009, i_13_4050, i_13_4051, i_13_4077, i_13_4086, i_13_4088, i_13_4104, i_13_4195, i_13_4312, i_13_4377, i_13_4428, i_13_4429, i_13_4540, i_13_4582, o_13_475);
	kernel_13_476 k_13_476(i_13_182, i_13_193, i_13_319, i_13_325, i_13_328, i_13_349, i_13_415, i_13_416, i_13_424, i_13_658, i_13_715, i_13_716, i_13_813, i_13_814, i_13_826, i_13_848, i_13_859, i_13_860, i_13_863, i_13_895, i_13_1072, i_13_1219, i_13_1224, i_13_1225, i_13_1226, i_13_1228, i_13_1229, i_13_1252, i_13_1255, i_13_1259, i_13_1315, i_13_1316, i_13_1318, i_13_1319, i_13_1345, i_13_1391, i_13_1404, i_13_1405, i_13_1411, i_13_1432, i_13_1444, i_13_1451, i_13_1484, i_13_1486, i_13_1490, i_13_1492, i_13_1541, i_13_1549, i_13_1553, i_13_1597, i_13_1677, i_13_1714, i_13_1750, i_13_1774, i_13_1778, i_13_1855, i_13_1871, i_13_1904, i_13_1922, i_13_1954, i_13_1955, i_13_1957, i_13_2056, i_13_2059, i_13_2137, i_13_2268, i_13_2506, i_13_2543, i_13_2611, i_13_2613, i_13_2614, i_13_2618, i_13_2633, i_13_2659, i_13_2660, i_13_2698, i_13_2705, i_13_2979, i_13_3005, i_13_3114, i_13_3119, i_13_3175, i_13_3287, i_13_3352, i_13_3369, i_13_3370, i_13_3421, i_13_3485, i_13_3506, i_13_3538, i_13_3539, i_13_3574, i_13_3595, i_13_3853, i_13_3979, i_13_4036, i_13_4249, i_13_4369, i_13_4376, i_13_4589, o_13_476);
	kernel_13_477 k_13_477(i_13_35, i_13_40, i_13_48, i_13_63, i_13_71, i_13_121, i_13_135, i_13_230, i_13_241, i_13_306, i_13_310, i_13_316, i_13_319, i_13_414, i_13_550, i_13_557, i_13_588, i_13_598, i_13_604, i_13_609, i_13_612, i_13_613, i_13_671, i_13_679, i_13_680, i_13_685, i_13_688, i_13_764, i_13_819, i_13_953, i_13_1116, i_13_1132, i_13_1207, i_13_1224, i_13_1269, i_13_1308, i_13_1422, i_13_1440, i_13_1441, i_13_1507, i_13_1526, i_13_1548, i_13_1596, i_13_1609, i_13_1673, i_13_1699, i_13_1700, i_13_1729, i_13_1764, i_13_1799, i_13_1847, i_13_1926, i_13_1927, i_13_1930, i_13_1944, i_13_2426, i_13_2461, i_13_2550, i_13_2557, i_13_2584, i_13_2673, i_13_2676, i_13_2718, i_13_2749, i_13_2771, i_13_3000, i_13_3217, i_13_3245, i_13_3267, i_13_3367, i_13_3483, i_13_3558, i_13_3637, i_13_3641, i_13_3653, i_13_3743, i_13_3754, i_13_3816, i_13_3871, i_13_3924, i_13_3937, i_13_3986, i_13_4032, i_13_4033, i_13_4035, i_13_4039, i_13_4217, i_13_4248, i_13_4250, i_13_4251, i_13_4293, i_13_4294, i_13_4298, i_13_4367, i_13_4521, i_13_4522, i_13_4565, i_13_4591, i_13_4593, i_13_4594, o_13_477);
	kernel_13_478 k_13_478(i_13_61, i_13_168, i_13_170, i_13_195, i_13_327, i_13_391, i_13_422, i_13_528, i_13_535, i_13_572, i_13_598, i_13_664, i_13_734, i_13_798, i_13_799, i_13_800, i_13_812, i_13_826, i_13_853, i_13_861, i_13_862, i_13_909, i_13_951, i_13_958, i_13_1069, i_13_1087, i_13_1119, i_13_1219, i_13_1226, i_13_1227, i_13_1228, i_13_1230, i_13_1231, i_13_1257, i_13_1258, i_13_1285, i_13_1300, i_13_1301, i_13_1302, i_13_1410, i_13_1437, i_13_1446, i_13_1482, i_13_1491, i_13_1492, i_13_1496, i_13_1523, i_13_1552, i_13_1554, i_13_1555, i_13_1755, i_13_1804, i_13_1829, i_13_1860, i_13_1959, i_13_1960, i_13_2008, i_13_2014, i_13_2103, i_13_2225, i_13_2239, i_13_2317, i_13_2347, i_13_2491, i_13_2535, i_13_2571, i_13_2707, i_13_2857, i_13_2972, i_13_2976, i_13_3121, i_13_3136, i_13_3145, i_13_3219, i_13_3233, i_13_3310, i_13_3410, i_13_3422, i_13_3423, i_13_3487, i_13_3489, i_13_3490, i_13_3531, i_13_3543, i_13_3639, i_13_3688, i_13_3739, i_13_3805, i_13_3858, i_13_3859, i_13_3984, i_13_3985, i_13_4380, i_13_4381, i_13_4396, i_13_4416, i_13_4454, i_13_4512, i_13_4528, i_13_4587, o_13_478);
	kernel_13_479 k_13_479(i_13_51, i_13_159, i_13_209, i_13_245, i_13_323, i_13_339, i_13_358, i_13_384, i_13_385, i_13_466, i_13_511, i_13_520, i_13_527, i_13_591, i_13_643, i_13_674, i_13_678, i_13_728, i_13_744, i_13_745, i_13_762, i_13_763, i_13_940, i_13_962, i_13_1066, i_13_1074, i_13_1130, i_13_1131, i_13_1213, i_13_1245, i_13_1301, i_13_1302, i_13_1303, i_13_1313, i_13_1346, i_13_1390, i_13_1403, i_13_1606, i_13_1632, i_13_1633, i_13_1634, i_13_1816, i_13_1835, i_13_1995, i_13_1996, i_13_2057, i_13_2058, i_13_2059, i_13_2121, i_13_2122, i_13_2204, i_13_2239, i_13_2265, i_13_2266, i_13_2267, i_13_2436, i_13_2460, i_13_2543, i_13_2617, i_13_2699, i_13_2847, i_13_2848, i_13_2859, i_13_2921, i_13_2941, i_13_3009, i_13_3011, i_13_3021, i_13_3022, i_13_3154, i_13_3273, i_13_3345, i_13_3346, i_13_3390, i_13_3399, i_13_3536, i_13_3542, i_13_3578, i_13_3619, i_13_3634, i_13_3669, i_13_3670, i_13_3692, i_13_3729, i_13_3731, i_13_3738, i_13_3739, i_13_3844, i_13_3846, i_13_3847, i_13_3892, i_13_3909, i_13_3911, i_13_4056, i_13_4217, i_13_4236, i_13_4255, i_13_4273, i_13_4399, i_13_4546, o_13_479);
	kernel_13_480 k_13_480(i_13_283, i_13_287, i_13_371, i_13_382, i_13_383, i_13_385, i_13_443, i_13_524, i_13_583, i_13_655, i_13_692, i_13_794, i_13_839, i_13_848, i_13_935, i_13_1018, i_13_1019, i_13_1088, i_13_1099, i_13_1136, i_13_1138, i_13_1331, i_13_1424, i_13_1441, i_13_1442, i_13_1496, i_13_1508, i_13_1520, i_13_1594, i_13_1630, i_13_1631, i_13_1639, i_13_1742, i_13_1792, i_13_1793, i_13_1799, i_13_1834, i_13_1999, i_13_2000, i_13_2003, i_13_2008, i_13_2050, i_13_2197, i_13_2198, i_13_2231, i_13_2233, i_13_2234, i_13_2269, i_13_2273, i_13_2411, i_13_2422, i_13_2459, i_13_2461, i_13_2462, i_13_2539, i_13_2540, i_13_2615, i_13_2852, i_13_2917, i_13_2918, i_13_2959, i_13_2987, i_13_3023, i_13_3032, i_13_3076, i_13_3134, i_13_3143, i_13_3169, i_13_3215, i_13_3247, i_13_3262, i_13_3304, i_13_3329, i_13_3350, i_13_3401, i_13_3686, i_13_3727, i_13_3728, i_13_3731, i_13_3871, i_13_3872, i_13_3907, i_13_3908, i_13_4007, i_13_4016, i_13_4018, i_13_4093, i_13_4100, i_13_4121, i_13_4204, i_13_4259, i_13_4339, i_13_4417, i_13_4513, i_13_4556, i_13_4558, i_13_4559, i_13_4571, i_13_4600, i_13_4601, o_13_480);
	kernel_13_481 k_13_481(i_13_61, i_13_118, i_13_130, i_13_136, i_13_168, i_13_282, i_13_312, i_13_357, i_13_364, i_13_492, i_13_528, i_13_645, i_13_646, i_13_663, i_13_717, i_13_726, i_13_826, i_13_888, i_13_958, i_13_1021, i_13_1101, i_13_1228, i_13_1230, i_13_1257, i_13_1258, i_13_1303, i_13_1308, i_13_1320, i_13_1407, i_13_1446, i_13_1491, i_13_1492, i_13_1500, i_13_1501, i_13_1554, i_13_1555, i_13_1572, i_13_1599, i_13_1641, i_13_1642, i_13_1699, i_13_1759, i_13_1795, i_13_1804, i_13_1806, i_13_1807, i_13_1959, i_13_1960, i_13_2014, i_13_2103, i_13_2145, i_13_2175, i_13_2193, i_13_2202, i_13_2205, i_13_2238, i_13_2239, i_13_2247, i_13_2430, i_13_2431, i_13_2445, i_13_2446, i_13_2508, i_13_2509, i_13_2514, i_13_2536, i_13_2608, i_13_2698, i_13_2818, i_13_2824, i_13_2937, i_13_2938, i_13_3244, i_13_3310, i_13_3420, i_13_3423, i_13_3426, i_13_3489, i_13_3543, i_13_3612, i_13_3639, i_13_3756, i_13_3805, i_13_3858, i_13_3859, i_13_3919, i_13_3936, i_13_3984, i_13_3985, i_13_4012, i_13_4065, i_13_4066, i_13_4215, i_13_4234, i_13_4272, i_13_4315, i_13_4380, i_13_4432, i_13_4512, i_13_4536, o_13_481);
	kernel_13_482 k_13_482(i_13_30, i_13_73, i_13_90, i_13_103, i_13_108, i_13_265, i_13_270, i_13_363, i_13_561, i_13_603, i_13_669, i_13_670, i_13_675, i_13_679, i_13_685, i_13_742, i_13_814, i_13_865, i_13_945, i_13_1083, i_13_1143, i_13_1215, i_13_1216, i_13_1284, i_13_1285, i_13_1324, i_13_1470, i_13_1515, i_13_1516, i_13_1620, i_13_1623, i_13_1801, i_13_1836, i_13_1837, i_13_1839, i_13_1840, i_13_1857, i_13_1912, i_13_2019, i_13_2133, i_13_2169, i_13_2275, i_13_2344, i_13_2434, i_13_2493, i_13_2496, i_13_2497, i_13_2529, i_13_2559, i_13_2610, i_13_2712, i_13_2934, i_13_2935, i_13_2955, i_13_3043, i_13_3096, i_13_3097, i_13_3099, i_13_3100, i_13_3142, i_13_3144, i_13_3149, i_13_3160, i_13_3162, i_13_3289, i_13_3415, i_13_3455, i_13_3475, i_13_3535, i_13_3546, i_13_3549, i_13_3567, i_13_3684, i_13_3738, i_13_3762, i_13_3763, i_13_3792, i_13_3802, i_13_3870, i_13_3936, i_13_3981, i_13_4005, i_13_4042, i_13_4045, i_13_4116, i_13_4123, i_13_4159, i_13_4188, i_13_4249, i_13_4260, i_13_4266, i_13_4324, i_13_4350, i_13_4365, i_13_4378, i_13_4413, i_13_4491, i_13_4512, i_13_4539, i_13_4557, o_13_482);
	kernel_13_483 k_13_483(i_13_22, i_13_45, i_13_48, i_13_240, i_13_319, i_13_370, i_13_450, i_13_451, i_13_453, i_13_561, i_13_587, i_13_598, i_13_622, i_13_928, i_13_940, i_13_1063, i_13_1064, i_13_1091, i_13_1244, i_13_1265, i_13_1297, i_13_1319, i_13_1342, i_13_1460, i_13_1468, i_13_1486, i_13_1495, i_13_1530, i_13_1566, i_13_1568, i_13_1569, i_13_1593, i_13_1594, i_13_1764, i_13_1774, i_13_1809, i_13_1810, i_13_1848, i_13_1884, i_13_1927, i_13_1959, i_13_1999, i_13_2107, i_13_2233, i_13_2278, i_13_2451, i_13_2452, i_13_2488, i_13_2543, i_13_2544, i_13_2617, i_13_2709, i_13_2710, i_13_2784, i_13_2882, i_13_2885, i_13_2886, i_13_2935, i_13_3016, i_13_3121, i_13_3213, i_13_3214, i_13_3216, i_13_3231, i_13_3244, i_13_3268, i_13_3286, i_13_3308, i_13_3340, i_13_3366, i_13_3367, i_13_3378, i_13_3388, i_13_3460, i_13_3532, i_13_3612, i_13_3688, i_13_3731, i_13_3763, i_13_3803, i_13_3817, i_13_3820, i_13_3876, i_13_3891, i_13_3999, i_13_4042, i_13_4063, i_13_4086, i_13_4087, i_13_4214, i_13_4266, i_13_4267, i_13_4269, i_13_4270, i_13_4313, i_13_4362, i_13_4371, i_13_4415, i_13_4459, i_13_4560, o_13_483);
	kernel_13_484 k_13_484(i_13_11, i_13_46, i_13_47, i_13_67, i_13_70, i_13_71, i_13_155, i_13_184, i_13_185, i_13_211, i_13_235, i_13_403, i_13_466, i_13_518, i_13_521, i_13_599, i_13_678, i_13_695, i_13_698, i_13_745, i_13_760, i_13_763, i_13_764, i_13_812, i_13_1062, i_13_1129, i_13_1132, i_13_1133, i_13_1189, i_13_1208, i_13_1210, i_13_1211, i_13_1310, i_13_1313, i_13_1394, i_13_1403, i_13_1506, i_13_1522, i_13_1548, i_13_1604, i_13_1659, i_13_1661, i_13_1673, i_13_1727, i_13_1927, i_13_1931, i_13_1945, i_13_1964, i_13_1967, i_13_2025, i_13_2097, i_13_2115, i_13_2132, i_13_2143, i_13_2316, i_13_2402, i_13_2552, i_13_2722, i_13_2767, i_13_2783, i_13_2848, i_13_2881, i_13_2884, i_13_3077, i_13_3091, i_13_3172, i_13_3251, i_13_3289, i_13_3308, i_13_3366, i_13_3370, i_13_3458, i_13_3542, i_13_3547, i_13_3591, i_13_3595, i_13_3611, i_13_3631, i_13_3636, i_13_3638, i_13_3641, i_13_3668, i_13_3752, i_13_3780, i_13_3890, i_13_3895, i_13_3898, i_13_3919, i_13_4036, i_13_4039, i_13_4214, i_13_4230, i_13_4270, i_13_4322, i_13_4332, i_13_4368, i_13_4397, i_13_4594, i_13_4595, i_13_4607, o_13_484);
	kernel_13_485 k_13_485(i_13_52, i_13_53, i_13_71, i_13_130, i_13_175, i_13_176, i_13_251, i_13_276, i_13_373, i_13_479, i_13_518, i_13_520, i_13_521, i_13_527, i_13_584, i_13_616, i_13_655, i_13_656, i_13_679, i_13_680, i_13_692, i_13_718, i_13_841, i_13_844, i_13_985, i_13_1084, i_13_1268, i_13_1330, i_13_1331, i_13_1435, i_13_1492, i_13_1573, i_13_1574, i_13_1663, i_13_1723, i_13_1754, i_13_1786, i_13_1814, i_13_1943, i_13_2024, i_13_2056, i_13_2057, i_13_2059, i_13_2060, i_13_2185, i_13_2186, i_13_2209, i_13_2239, i_13_2321, i_13_2455, i_13_2461, i_13_2507, i_13_2509, i_13_2510, i_13_2651, i_13_2698, i_13_2699, i_13_2733, i_13_2752, i_13_2753, i_13_2959, i_13_3068, i_13_3077, i_13_3100, i_13_3112, i_13_3163, i_13_3217, i_13_3256, i_13_3292, i_13_3373, i_13_3374, i_13_3406, i_13_3526, i_13_3571, i_13_3572, i_13_3613, i_13_3662, i_13_3725, i_13_3749, i_13_3767, i_13_3769, i_13_3830, i_13_3847, i_13_3874, i_13_3877, i_13_3991, i_13_3995, i_13_4009, i_13_4021, i_13_4022, i_13_4048, i_13_4127, i_13_4157, i_13_4189, i_13_4318, i_13_4319, i_13_4558, i_13_4598, i_13_4603, i_13_4604, o_13_485);
	kernel_13_486 k_13_486(i_13_70, i_13_75, i_13_120, i_13_121, i_13_184, i_13_244, i_13_333, i_13_414, i_13_423, i_13_459, i_13_517, i_13_522, i_13_523, i_13_524, i_13_525, i_13_526, i_13_532, i_13_571, i_13_585, i_13_588, i_13_670, i_13_697, i_13_759, i_13_1057, i_13_1066, i_13_1116, i_13_1207, i_13_1216, i_13_1306, i_13_1307, i_13_1314, i_13_1317, i_13_1341, i_13_1342, i_13_1389, i_13_1399, i_13_1440, i_13_1441, i_13_1444, i_13_1494, i_13_1515, i_13_1602, i_13_1603, i_13_1774, i_13_1887, i_13_1930, i_13_1944, i_13_1945, i_13_1998, i_13_2001, i_13_2025, i_13_2026, i_13_2124, i_13_2125, i_13_2196, i_13_2197, i_13_2278, i_13_2445, i_13_2533, i_13_2710, i_13_2766, i_13_2781, i_13_2902, i_13_2916, i_13_2917, i_13_2918, i_13_2983, i_13_3007, i_13_3046, i_13_3163, i_13_3208, i_13_3366, i_13_3367, i_13_3396, i_13_3406, i_13_3414, i_13_3438, i_13_3460, i_13_3541, i_13_3559, i_13_3573, i_13_3575, i_13_3592, i_13_3637, i_13_3666, i_13_3667, i_13_3726, i_13_3766, i_13_3907, i_13_4096, i_13_4105, i_13_4149, i_13_4204, i_13_4350, i_13_4351, i_13_4392, i_13_4441, i_13_4446, i_13_4447, i_13_4567, o_13_486);
	kernel_13_487 k_13_487(i_13_40, i_13_110, i_13_126, i_13_132, i_13_273, i_13_282, i_13_283, i_13_284, i_13_335, i_13_357, i_13_360, i_13_361, i_13_472, i_13_519, i_13_538, i_13_689, i_13_838, i_13_866, i_13_867, i_13_869, i_13_1096, i_13_1111, i_13_1112, i_13_1114, i_13_1119, i_13_1132, i_13_1243, i_13_1329, i_13_1430, i_13_1501, i_13_1549, i_13_1745, i_13_1770, i_13_1792, i_13_1795, i_13_1834, i_13_1858, i_13_1884, i_13_1896, i_13_2004, i_13_2008, i_13_2010, i_13_2017, i_13_2097, i_13_2113, i_13_2145, i_13_2148, i_13_2223, i_13_2260, i_13_2384, i_13_2461, i_13_2514, i_13_2537, i_13_2733, i_13_2798, i_13_2883, i_13_2890, i_13_3048, i_13_3057, i_13_3059, i_13_3076, i_13_3077, i_13_3097, i_13_3145, i_13_3219, i_13_3266, i_13_3286, i_13_3315, i_13_3348, i_13_3489, i_13_3490, i_13_3549, i_13_3550, i_13_3604, i_13_3671, i_13_3730, i_13_3735, i_13_3748, i_13_3822, i_13_3869, i_13_3881, i_13_3909, i_13_3910, i_13_3952, i_13_4018, i_13_4125, i_13_4126, i_13_4165, i_13_4261, i_13_4272, i_13_4330, i_13_4333, i_13_4362, i_13_4433, i_13_4454, i_13_4467, i_13_4471, i_13_4516, i_13_4565, i_13_4578, o_13_487);
	kernel_13_488 k_13_488(i_13_45, i_13_46, i_13_100, i_13_127, i_13_154, i_13_193, i_13_252, i_13_270, i_13_271, i_13_374, i_13_378, i_13_379, i_13_425, i_13_428, i_13_451, i_13_523, i_13_569, i_13_570, i_13_688, i_13_817, i_13_927, i_13_949, i_13_1063, i_13_1087, i_13_1147, i_13_1219, i_13_1271, i_13_1345, i_13_1379, i_13_1435, i_13_1458, i_13_1496, i_13_1539, i_13_1566, i_13_1567, i_13_1733, i_13_1749, i_13_1800, i_13_1801, i_13_1802, i_13_1810, i_13_1848, i_13_1891, i_13_2026, i_13_2107, i_13_2108, i_13_2146, i_13_2197, i_13_2233, i_13_2260, i_13_2435, i_13_2525, i_13_2576, i_13_2614, i_13_2618, i_13_2713, i_13_2740, i_13_2745, i_13_2747, i_13_2763, i_13_2917, i_13_2935, i_13_2987, i_13_3008, i_13_3016, i_13_3056, i_13_3214, i_13_3215, i_13_3367, i_13_3376, i_13_3377, i_13_3528, i_13_3547, i_13_3591, i_13_3722, i_13_3742, i_13_3763, i_13_3769, i_13_3770, i_13_3817, i_13_3821, i_13_3905, i_13_3978, i_13_4042, i_13_4064, i_13_4086, i_13_4087, i_13_4234, i_13_4250, i_13_4258, i_13_4266, i_13_4267, i_13_4268, i_13_4312, i_13_4322, i_13_4358, i_13_4385, i_13_4447, i_13_4562, i_13_4564, o_13_488);
	kernel_13_489 k_13_489(i_13_73, i_13_108, i_13_111, i_13_112, i_13_136, i_13_261, i_13_363, i_13_387, i_13_442, i_13_581, i_13_603, i_13_604, i_13_666, i_13_669, i_13_810, i_13_813, i_13_814, i_13_855, i_13_856, i_13_1017, i_13_1081, i_13_1144, i_13_1211, i_13_1215, i_13_1216, i_13_1422, i_13_1423, i_13_1426, i_13_1454, i_13_1485, i_13_1486, i_13_1494, i_13_1566, i_13_1597, i_13_1620, i_13_1622, i_13_1629, i_13_1719, i_13_1774, i_13_1794, i_13_1812, i_13_1836, i_13_1837, i_13_1840, i_13_1849, i_13_1938, i_13_1989, i_13_2011, i_13_2137, i_13_2169, i_13_2404, i_13_2407, i_13_2434, i_13_2448, i_13_2451, i_13_2452, i_13_2497, i_13_2538, i_13_2610, i_13_2858, i_13_2907, i_13_2916, i_13_2917, i_13_2935, i_13_2938, i_13_3000, i_13_3100, i_13_3144, i_13_3213, i_13_3288, i_13_3315, i_13_3340, i_13_3384, i_13_3385, i_13_3393, i_13_3474, i_13_3475, i_13_3501, i_13_3502, i_13_3528, i_13_3529, i_13_3702, i_13_3738, i_13_3739, i_13_3888, i_13_3891, i_13_4055, i_13_4060, i_13_4063, i_13_4159, i_13_4204, i_13_4248, i_13_4251, i_13_4315, i_13_4338, i_13_4342, i_13_4365, i_13_4366, i_13_4368, i_13_4540, o_13_489);
	kernel_13_490 k_13_490(i_13_19, i_13_31, i_13_99, i_13_112, i_13_162, i_13_165, i_13_166, i_13_180, i_13_183, i_13_184, i_13_185, i_13_216, i_13_217, i_13_256, i_13_393, i_13_639, i_13_796, i_13_837, i_13_1063, i_13_1078, i_13_1116, i_13_1118, i_13_1121, i_13_1146, i_13_1219, i_13_1231, i_13_1263, i_13_1323, i_13_1326, i_13_1426, i_13_1458, i_13_1480, i_13_1513, i_13_1521, i_13_1525, i_13_1677, i_13_1746, i_13_1764, i_13_1784, i_13_1804, i_13_1831, i_13_1840, i_13_1857, i_13_1909, i_13_1938, i_13_1940, i_13_1989, i_13_1999, i_13_2002, i_13_2043, i_13_2106, i_13_2107, i_13_2116, i_13_2145, i_13_2146, i_13_2185, i_13_2233, i_13_2260, i_13_2277, i_13_2340, i_13_2395, i_13_2466, i_13_2476, i_13_2564, i_13_2748, i_13_2761, i_13_2937, i_13_2979, i_13_2980, i_13_2997, i_13_3024, i_13_3026, i_13_3027, i_13_3108, i_13_3111, i_13_3115, i_13_3144, i_13_3145, i_13_3196, i_13_3208, i_13_3286, i_13_3289, i_13_3471, i_13_3558, i_13_3650, i_13_3730, i_13_3763, i_13_3892, i_13_4042, i_13_4077, i_13_4187, i_13_4203, i_13_4204, i_13_4268, i_13_4314, i_13_4396, i_13_4501, i_13_4558, i_13_4564, i_13_4600, o_13_490);
	kernel_13_491 k_13_491(i_13_27, i_13_64, i_13_104, i_13_131, i_13_157, i_13_174, i_13_208, i_13_209, i_13_218, i_13_225, i_13_266, i_13_307, i_13_355, i_13_356, i_13_441, i_13_463, i_13_464, i_13_526, i_13_531, i_13_549, i_13_613, i_13_639, i_13_666, i_13_667, i_13_742, i_13_812, i_13_839, i_13_841, i_13_961, i_13_1019, i_13_1073, i_13_1129, i_13_1301, i_13_1307, i_13_1444, i_13_1535, i_13_1594, i_13_1595, i_13_1604, i_13_1624, i_13_1632, i_13_1639, i_13_1697, i_13_1723, i_13_1774, i_13_1846, i_13_1847, i_13_1909, i_13_2030, i_13_2091, i_13_2101, i_13_2143, i_13_2199, i_13_2200, i_13_2237, i_13_2263, i_13_2297, i_13_2444, i_13_2504, i_13_2507, i_13_2512, i_13_2551, i_13_2673, i_13_2691, i_13_2822, i_13_2885, i_13_2936, i_13_3070, i_13_3089, i_13_3143, i_13_3241, i_13_3242, i_13_3343, i_13_3389, i_13_3460, i_13_3469, i_13_3472, i_13_3530, i_13_3595, i_13_3599, i_13_3619, i_13_3631, i_13_3637, i_13_3667, i_13_3682, i_13_3719, i_13_3728, i_13_3793, i_13_3857, i_13_3924, i_13_3935, i_13_3989, i_13_4060, i_13_4061, i_13_4077, i_13_4122, i_13_4313, i_13_4342, i_13_4345, i_13_4379, o_13_491);
	kernel_13_492 k_13_492(i_13_44, i_13_45, i_13_46, i_13_55, i_13_84, i_13_94, i_13_112, i_13_134, i_13_207, i_13_234, i_13_243, i_13_244, i_13_283, i_13_323, i_13_521, i_13_598, i_13_614, i_13_623, i_13_693, i_13_694, i_13_702, i_13_760, i_13_838, i_13_955, i_13_1071, i_13_1116, i_13_1119, i_13_1128, i_13_1129, i_13_1152, i_13_1219, i_13_1243, i_13_1317, i_13_1360, i_13_1405, i_13_1521, i_13_1533, i_13_1535, i_13_1647, i_13_1678, i_13_1777, i_13_1795, i_13_1804, i_13_1840, i_13_1929, i_13_1957, i_13_2002, i_13_2142, i_13_2208, i_13_2254, i_13_2460, i_13_2511, i_13_2512, i_13_2541, i_13_2578, i_13_2646, i_13_2666, i_13_2692, i_13_2845, i_13_2880, i_13_2910, i_13_3000, i_13_3002, i_13_3025, i_13_3113, i_13_3127, i_13_3367, i_13_3371, i_13_3420, i_13_3474, i_13_3475, i_13_3519, i_13_3528, i_13_3546, i_13_3636, i_13_3641, i_13_3753, i_13_3757, i_13_3819, i_13_3887, i_13_3898, i_13_3923, i_13_3987, i_13_4035, i_13_4036, i_13_4041, i_13_4167, i_13_4311, i_13_4329, i_13_4351, i_13_4377, i_13_4378, i_13_4414, i_13_4430, i_13_4450, i_13_4509, i_13_4510, i_13_4567, i_13_4593, i_13_4603, o_13_492);
	kernel_13_493 k_13_493(i_13_30, i_13_38, i_13_158, i_13_161, i_13_172, i_13_173, i_13_175, i_13_190, i_13_247, i_13_280, i_13_281, i_13_283, i_13_284, i_13_316, i_13_334, i_13_488, i_13_525, i_13_527, i_13_577, i_13_640, i_13_685, i_13_688, i_13_689, i_13_797, i_13_820, i_13_821, i_13_822, i_13_847, i_13_1067, i_13_1120, i_13_1216, i_13_1219, i_13_1225, i_13_1306, i_13_1309, i_13_1504, i_13_1540, i_13_1594, i_13_1601, i_13_1730, i_13_1768, i_13_1813, i_13_1882, i_13_1926, i_13_2054, i_13_2092, i_13_2173, i_13_2188, i_13_2189, i_13_2236, i_13_2422, i_13_2425, i_13_2443, i_13_2475, i_13_2622, i_13_2674, i_13_2677, i_13_2702, i_13_3007, i_13_3069, i_13_3142, i_13_3214, i_13_3217, i_13_3250, i_13_3267, i_13_3268, i_13_3271, i_13_3272, i_13_3378, i_13_3386, i_13_3389, i_13_3421, i_13_3424, i_13_3451, i_13_3457, i_13_3722, i_13_3726, i_13_3730, i_13_3906, i_13_3910, i_13_3917, i_13_3982, i_13_3991, i_13_4014, i_13_4015, i_13_4016, i_13_4018, i_13_4062, i_13_4081, i_13_4180, i_13_4214, i_13_4249, i_13_4257, i_13_4261, i_13_4306, i_13_4374, i_13_4396, i_13_4424, i_13_4450, i_13_4544, o_13_493);
	kernel_13_494 k_13_494(i_13_25, i_13_31, i_13_40, i_13_74, i_13_139, i_13_186, i_13_229, i_13_317, i_13_454, i_13_510, i_13_573, i_13_589, i_13_659, i_13_661, i_13_663, i_13_733, i_13_854, i_13_938, i_13_940, i_13_1021, i_13_1075, i_13_1144, i_13_1145, i_13_1282, i_13_1284, i_13_1320, i_13_1424, i_13_1437, i_13_1660, i_13_1669, i_13_1714, i_13_1723, i_13_1773, i_13_1775, i_13_2188, i_13_2297, i_13_2425, i_13_2611, i_13_2659, i_13_2705, i_13_2742, i_13_2857, i_13_2958, i_13_3009, i_13_3010, i_13_3013, i_13_3046, i_13_3050, i_13_3072, i_13_3108, i_13_3109, i_13_3111, i_13_3156, i_13_3157, i_13_3205, i_13_3388, i_13_3408, i_13_3442, i_13_3460, i_13_3463, i_13_3468, i_13_3483, i_13_3484, i_13_3487, i_13_3489, i_13_3504, i_13_3550, i_13_3552, i_13_3565, i_13_3566, i_13_3568, i_13_3577, i_13_3603, i_13_3648, i_13_3681, i_13_3763, i_13_3764, i_13_3803, i_13_3819, i_13_3822, i_13_3862, i_13_3865, i_13_3980, i_13_4054, i_13_4163, i_13_4251, i_13_4312, i_13_4325, i_13_4340, i_13_4366, i_13_4367, i_13_4369, i_13_4370, i_13_4372, i_13_4396, i_13_4479, i_13_4558, i_13_4560, i_13_4568, i_13_4600, o_13_494);
	kernel_13_495 k_13_495(i_13_42, i_13_43, i_13_76, i_13_102, i_13_107, i_13_117, i_13_118, i_13_169, i_13_180, i_13_181, i_13_225, i_13_394, i_13_489, i_13_504, i_13_534, i_13_567, i_13_572, i_13_607, i_13_617, i_13_624, i_13_645, i_13_651, i_13_697, i_13_711, i_13_835, i_13_841, i_13_945, i_13_948, i_13_1072, i_13_1092, i_13_1115, i_13_1210, i_13_1225, i_13_1276, i_13_1300, i_13_1404, i_13_1522, i_13_1629, i_13_1719, i_13_1767, i_13_1782, i_13_1783, i_13_1785, i_13_1786, i_13_1801, i_13_2014, i_13_2056, i_13_2119, i_13_2182, i_13_2205, i_13_2206, i_13_2209, i_13_2280, i_13_2307, i_13_2321, i_13_2361, i_13_2394, i_13_2403, i_13_2427, i_13_2428, i_13_2452, i_13_2457, i_13_2458, i_13_2680, i_13_2879, i_13_2934, i_13_2938, i_13_3015, i_13_3019, i_13_3160, i_13_3163, i_13_3171, i_13_3204, i_13_3213, i_13_3214, i_13_3217, i_13_3231, i_13_3270, i_13_3420, i_13_3421, i_13_3426, i_13_3531, i_13_3532, i_13_3548, i_13_3562, i_13_3699, i_13_3745, i_13_3870, i_13_3873, i_13_3912, i_13_3981, i_13_3982, i_13_4005, i_13_4006, i_13_4017, i_13_4254, i_13_4302, i_13_4311, i_13_4413, i_13_4518, o_13_495);
	kernel_13_496 k_13_496(i_13_71, i_13_79, i_13_169, i_13_171, i_13_175, i_13_216, i_13_233, i_13_246, i_13_325, i_13_397, i_13_604, i_13_613, i_13_624, i_13_643, i_13_679, i_13_683, i_13_685, i_13_694, i_13_697, i_13_819, i_13_822, i_13_826, i_13_841, i_13_854, i_13_855, i_13_878, i_13_937, i_13_973, i_13_1021, i_13_1062, i_13_1119, i_13_1120, i_13_1132, i_13_1224, i_13_1225, i_13_1308, i_13_1313, i_13_1315, i_13_1377, i_13_1485, i_13_1506, i_13_1525, i_13_1553, i_13_1663, i_13_1745, i_13_1771, i_13_1798, i_13_1799, i_13_1944, i_13_1948, i_13_1954, i_13_2000, i_13_2383, i_13_2452, i_13_2677, i_13_2749, i_13_2848, i_13_2878, i_13_3006, i_13_3007, i_13_3008, i_13_3094, i_13_3107, i_13_3168, i_13_3216, i_13_3352, i_13_3424, i_13_3429, i_13_3450, i_13_3487, i_13_3506, i_13_3538, i_13_3652, i_13_3728, i_13_3739, i_13_3742, i_13_3782, i_13_3895, i_13_3927, i_13_3937, i_13_3982, i_13_3994, i_13_4063, i_13_4096, i_13_4186, i_13_4188, i_13_4249, i_13_4252, i_13_4255, i_13_4256, i_13_4258, i_13_4261, i_13_4297, i_13_4300, i_13_4366, i_13_4372, i_13_4433, i_13_4447, i_13_4536, i_13_4598, o_13_496);
	kernel_13_497 k_13_497(i_13_69, i_13_142, i_13_385, i_13_386, i_13_448, i_13_537, i_13_664, i_13_691, i_13_836, i_13_844, i_13_848, i_13_892, i_13_989, i_13_1102, i_13_1219, i_13_1228, i_13_1276, i_13_1287, i_13_1345, i_13_1402, i_13_1403, i_13_1444, i_13_1510, i_13_1600, i_13_1644, i_13_1678, i_13_1717, i_13_1725, i_13_1726, i_13_1748, i_13_1934, i_13_1948, i_13_1960, i_13_1995, i_13_1996, i_13_1999, i_13_2002, i_13_2060, i_13_2127, i_13_2194, i_13_2281, i_13_2311, i_13_2361, i_13_2379, i_13_2464, i_13_2470, i_13_2534, i_13_2698, i_13_2716, i_13_2726, i_13_2771, i_13_2857, i_13_2860, i_13_2887, i_13_2917, i_13_2949, i_13_3017, i_13_3028, i_13_3065, i_13_3066, i_13_3067, i_13_3068, i_13_3074, i_13_3329, i_13_3352, i_13_3446, i_13_3454, i_13_3490, i_13_3547, i_13_3595, i_13_3683, i_13_3686, i_13_3688, i_13_3689, i_13_3722, i_13_3737, i_13_3781, i_13_3900, i_13_3928, i_13_3988, i_13_3994, i_13_3995, i_13_4017, i_13_4054, i_13_4057, i_13_4094, i_13_4165, i_13_4214, i_13_4273, i_13_4304, i_13_4309, i_13_4393, i_13_4396, i_13_4399, i_13_4400, i_13_4411, i_13_4431, i_13_4432, i_13_4566, i_13_4597, o_13_497);
	kernel_13_498 k_13_498(i_13_77, i_13_130, i_13_134, i_13_256, i_13_368, i_13_394, i_13_469, i_13_515, i_13_518, i_13_550, i_13_554, i_13_605, i_13_623, i_13_626, i_13_656, i_13_658, i_13_659, i_13_661, i_13_695, i_13_698, i_13_814, i_13_841, i_13_889, i_13_940, i_13_978, i_13_1063, i_13_1072, i_13_1073, i_13_1084, i_13_1088, i_13_1109, i_13_1144, i_13_1145, i_13_1153, i_13_1154, i_13_1214, i_13_1265, i_13_1424, i_13_1517, i_13_1535, i_13_1657, i_13_1658, i_13_1660, i_13_1730, i_13_1732, i_13_1733, i_13_1742, i_13_2017, i_13_2020, i_13_2021, i_13_2023, i_13_2131, i_13_2137, i_13_2209, i_13_2246, i_13_2297, i_13_2336, i_13_2401, i_13_2443, i_13_2461, i_13_2498, i_13_2513, i_13_2717, i_13_2740, i_13_2771, i_13_2882, i_13_2956, i_13_3044, i_13_3074, i_13_3075, i_13_3115, i_13_3154, i_13_3263, i_13_3476, i_13_3563, i_13_3568, i_13_3730, i_13_3740, i_13_3820, i_13_3910, i_13_4019, i_13_4091, i_13_4121, i_13_4160, i_13_4163, i_13_4187, i_13_4330, i_13_4333, i_13_4358, i_13_4360, i_13_4362, i_13_4363, i_13_4366, i_13_4367, i_13_4394, i_13_4429, i_13_4477, i_13_4514, i_13_4540, i_13_4603, o_13_498);
	kernel_13_499 k_13_499(i_13_46, i_13_139, i_13_185, i_13_331, i_13_334, i_13_335, i_13_352, i_13_362, i_13_409, i_13_449, i_13_451, i_13_506, i_13_568, i_13_626, i_13_649, i_13_658, i_13_769, i_13_884, i_13_932, i_13_935, i_13_937, i_13_1019, i_13_1024, i_13_1072, i_13_1073, i_13_1129, i_13_1130, i_13_1133, i_13_1148, i_13_1189, i_13_1244, i_13_1298, i_13_1328, i_13_1400, i_13_1406, i_13_1510, i_13_1523, i_13_1570, i_13_1649, i_13_1661, i_13_1679, i_13_1720, i_13_1727, i_13_1765, i_13_1888, i_13_1889, i_13_1933, i_13_1945, i_13_2026, i_13_2027, i_13_2135, i_13_2188, i_13_2197, i_13_2423, i_13_2470, i_13_2645, i_13_2694, i_13_2725, i_13_2741, i_13_2747, i_13_2801, i_13_2851, i_13_2899, i_13_2917, i_13_2966, i_13_2998, i_13_3028, i_13_3029, i_13_3073, i_13_3074, i_13_3163, i_13_3261, i_13_3262, i_13_3325, i_13_3378, i_13_3458, i_13_3484, i_13_3485, i_13_3547, i_13_3574, i_13_3575, i_13_3653, i_13_3728, i_13_3742, i_13_3760, i_13_3764, i_13_3781, i_13_3785, i_13_3853, i_13_3898, i_13_3899, i_13_4162, i_13_4231, i_13_4294, i_13_4298, i_13_4322, i_13_4360, i_13_4363, i_13_4537, i_13_4603, o_13_499);
	kernel_13_500 k_13_500(i_13_46, i_13_47, i_13_121, i_13_226, i_13_357, i_13_407, i_13_447, i_13_514, i_13_532, i_13_568, i_13_794, i_13_833, i_13_847, i_13_848, i_13_931, i_13_937, i_13_947, i_13_1019, i_13_1072, i_13_1073, i_13_1136, i_13_1201, i_13_1225, i_13_1298, i_13_1315, i_13_1495, i_13_1496, i_13_1630, i_13_1631, i_13_1720, i_13_1724, i_13_1777, i_13_1779, i_13_1805, i_13_1855, i_13_1945, i_13_1946, i_13_1948, i_13_2020, i_13_2026, i_13_2027, i_13_2099, i_13_2134, i_13_2197, i_13_2198, i_13_2227, i_13_2449, i_13_2450, i_13_2452, i_13_2459, i_13_2477, i_13_2539, i_13_2540, i_13_2548, i_13_2740, i_13_2782, i_13_2917, i_13_2918, i_13_3010, i_13_3028, i_13_3097, i_13_3169, i_13_3268, i_13_3397, i_13_3412, i_13_3451, i_13_3457, i_13_3458, i_13_3484, i_13_3570, i_13_3574, i_13_3575, i_13_3593, i_13_3704, i_13_3728, i_13_3781, i_13_3782, i_13_3800, i_13_3853, i_13_3898, i_13_3907, i_13_3908, i_13_4001, i_13_4016, i_13_4249, i_13_4250, i_13_4252, i_13_4253, i_13_4259, i_13_4322, i_13_4339, i_13_4342, i_13_4365, i_13_4375, i_13_4376, i_13_4447, i_13_4511, i_13_4556, i_13_4558, i_13_4570, o_13_500);
	kernel_13_501 k_13_501(i_13_31, i_13_36, i_13_37, i_13_102, i_13_255, i_13_262, i_13_264, i_13_265, i_13_282, i_13_492, i_13_505, i_13_532, i_13_535, i_13_577, i_13_616, i_13_651, i_13_675, i_13_676, i_13_723, i_13_777, i_13_810, i_13_837, i_13_838, i_13_871, i_13_948, i_13_949, i_13_981, i_13_1116, i_13_1197, i_13_1198, i_13_1212, i_13_1242, i_13_1269, i_13_1278, i_13_1324, i_13_1326, i_13_1380, i_13_1396, i_13_1446, i_13_1456, i_13_1504, i_13_1552, i_13_1746, i_13_1786, i_13_1803, i_13_1840, i_13_1857, i_13_1908, i_13_2010, i_13_2029, i_13_2046, i_13_2055, i_13_2056, i_13_2116, i_13_2136, i_13_2137, i_13_2172, i_13_2187, i_13_2224, i_13_2230, i_13_2311, i_13_2379, i_13_2394, i_13_2406, i_13_2425, i_13_2461, i_13_2502, i_13_2511, i_13_2664, i_13_2673, i_13_2691, i_13_2692, i_13_2715, i_13_2748, i_13_3024, i_13_3025, i_13_3114, i_13_3145, i_13_3153, i_13_3342, i_13_3369, i_13_3370, i_13_3373, i_13_3405, i_13_3412, i_13_3532, i_13_3579, i_13_3619, i_13_3871, i_13_3874, i_13_3987, i_13_3988, i_13_4032, i_13_4204, i_13_4305, i_13_4522, i_13_4524, i_13_4582, i_13_4590, i_13_4600, o_13_501);
	kernel_13_502 k_13_502(i_13_45, i_13_63, i_13_73, i_13_93, i_13_100, i_13_102, i_13_130, i_13_207, i_13_319, i_13_396, i_13_468, i_13_469, i_13_532, i_13_570, i_13_603, i_13_666, i_13_667, i_13_675, i_13_676, i_13_684, i_13_837, i_13_838, i_13_927, i_13_945, i_13_946, i_13_1024, i_13_1071, i_13_1098, i_13_1129, i_13_1144, i_13_1305, i_13_1306, i_13_1344, i_13_1399, i_13_1461, i_13_1503, i_13_1504, i_13_1593, i_13_1594, i_13_1620, i_13_1719, i_13_1720, i_13_1777, i_13_1791, i_13_1803, i_13_1804, i_13_1812, i_13_1837, i_13_1894, i_13_1908, i_13_1927, i_13_2016, i_13_2056, i_13_2137, i_13_2169, i_13_2197, i_13_2280, i_13_2344, i_13_2400, i_13_2431, i_13_2458, i_13_2479, i_13_2511, i_13_2547, i_13_2613, i_13_2614, i_13_2691, i_13_2692, i_13_2797, i_13_2820, i_13_2874, i_13_3019, i_13_3043, i_13_3088, i_13_3387, i_13_3423, i_13_3468, i_13_3475, i_13_3502, i_13_3531, i_13_3532, i_13_3618, i_13_3619, i_13_3687, i_13_3862, i_13_3934, i_13_3987, i_13_3988, i_13_4123, i_13_4260, i_13_4269, i_13_4311, i_13_4329, i_13_4392, i_13_4429, i_13_4446, i_13_4510, i_13_4518, i_13_4590, i_13_4600, o_13_502);
	kernel_13_503 k_13_503(i_13_92, i_13_139, i_13_176, i_13_184, i_13_185, i_13_193, i_13_364, i_13_407, i_13_482, i_13_589, i_13_604, i_13_607, i_13_608, i_13_658, i_13_659, i_13_661, i_13_662, i_13_686, i_13_712, i_13_814, i_13_851, i_13_859, i_13_868, i_13_949, i_13_956, i_13_982, i_13_1138, i_13_1148, i_13_1150, i_13_1210, i_13_1211, i_13_1226, i_13_1229, i_13_1244, i_13_1253, i_13_1301, i_13_1321, i_13_1487, i_13_1730, i_13_1765, i_13_1766, i_13_1804, i_13_1813, i_13_1829, i_13_1840, i_13_1892, i_13_1904, i_13_1961, i_13_2012, i_13_2020, i_13_2137, i_13_2182, i_13_2207, i_13_2281, i_13_2341, i_13_2435, i_13_2593, i_13_2857, i_13_2858, i_13_2938, i_13_2981, i_13_3047, i_13_3053, i_13_3110, i_13_3164, i_13_3254, i_13_3260, i_13_3268, i_13_3289, i_13_3349, i_13_3352, i_13_3442, i_13_3476, i_13_3484, i_13_3485, i_13_3491, i_13_3530, i_13_3547, i_13_3664, i_13_3667, i_13_3754, i_13_3764, i_13_3817, i_13_3821, i_13_3872, i_13_3875, i_13_3979, i_13_4006, i_13_4055, i_13_4160, i_13_4163, i_13_4249, i_13_4333, i_13_4358, i_13_4369, i_13_4370, i_13_4430, i_13_4537, i_13_4538, i_13_4565, o_13_503);
	kernel_13_504 k_13_504(i_13_34, i_13_44, i_13_67, i_13_70, i_13_94, i_13_95, i_13_418, i_13_435, i_13_447, i_13_449, i_13_592, i_13_593, i_13_607, i_13_665, i_13_679, i_13_681, i_13_698, i_13_763, i_13_764, i_13_1048, i_13_1075, i_13_1103, i_13_1106, i_13_1123, i_13_1131, i_13_1132, i_13_1213, i_13_1273, i_13_1312, i_13_1321, i_13_1349, i_13_1428, i_13_1544, i_13_1605, i_13_1606, i_13_1644, i_13_1672, i_13_1753, i_13_1780, i_13_1786, i_13_1796, i_13_1797, i_13_1798, i_13_1888, i_13_2004, i_13_2024, i_13_2120, i_13_2173, i_13_2382, i_13_2383, i_13_2455, i_13_2464, i_13_2570, i_13_2600, i_13_2679, i_13_2680, i_13_2725, i_13_2850, i_13_2851, i_13_2852, i_13_3003, i_13_3032, i_13_3076, i_13_3094, i_13_3163, i_13_3166, i_13_3265, i_13_3273, i_13_3311, i_13_3370, i_13_3391, i_13_3540, i_13_3541, i_13_3543, i_13_3545, i_13_3560, i_13_3651, i_13_3722, i_13_3741, i_13_3742, i_13_3757, i_13_3806, i_13_3900, i_13_3918, i_13_3940, i_13_4040, i_13_4083, i_13_4099, i_13_4297, i_13_4345, i_13_4381, i_13_4399, i_13_4417, i_13_4433, i_13_4561, i_13_4594, i_13_4595, i_13_4597, i_13_4598, i_13_4607, o_13_504);
	kernel_13_505 k_13_505(i_13_32, i_13_91, i_13_92, i_13_281, i_13_307, i_13_308, i_13_317, i_13_361, i_13_367, i_13_383, i_13_384, i_13_528, i_13_535, i_13_551, i_13_569, i_13_584, i_13_604, i_13_626, i_13_643, i_13_686, i_13_688, i_13_704, i_13_724, i_13_796, i_13_815, i_13_949, i_13_1067, i_13_1111, i_13_1216, i_13_1217, i_13_1219, i_13_1255, i_13_1321, i_13_1402, i_13_1432, i_13_1443, i_13_1471, i_13_1487, i_13_1552, i_13_1597, i_13_1635, i_13_1644, i_13_1657, i_13_1705, i_13_1721, i_13_1837, i_13_1900, i_13_1910, i_13_1922, i_13_1931, i_13_1999, i_13_2000, i_13_2002, i_13_2006, i_13_2056, i_13_2057, i_13_2173, i_13_2176, i_13_2231, i_13_2422, i_13_2423, i_13_2424, i_13_2452, i_13_2678, i_13_2767, i_13_2965, i_13_3039, i_13_3056, i_13_3064, i_13_3065, i_13_3127, i_13_3142, i_13_3145, i_13_3218, i_13_3372, i_13_3379, i_13_3415, i_13_3487, i_13_3524, i_13_3541, i_13_3700, i_13_3712, i_13_3794, i_13_3865, i_13_3871, i_13_4018, i_13_4037, i_13_4082, i_13_4118, i_13_4150, i_13_4217, i_13_4279, i_13_4306, i_13_4307, i_13_4339, i_13_4342, i_13_4350, i_13_4351, i_13_4397, i_13_4415, o_13_505);
	kernel_13_506 k_13_506(i_13_31, i_13_32, i_13_46, i_13_67, i_13_77, i_13_92, i_13_110, i_13_118, i_13_119, i_13_136, i_13_229, i_13_334, i_13_490, i_13_535, i_13_562, i_13_563, i_13_604, i_13_605, i_13_730, i_13_760, i_13_947, i_13_1084, i_13_1210, i_13_1216, i_13_1217, i_13_1315, i_13_1441, i_13_1442, i_13_1471, i_13_1486, i_13_1487, i_13_1507, i_13_1589, i_13_1606, i_13_1625, i_13_1633, i_13_1659, i_13_1678, i_13_1694, i_13_1731, i_13_1733, i_13_1787, i_13_1837, i_13_1840, i_13_1841, i_13_1886, i_13_1930, i_13_1931, i_13_1937, i_13_2000, i_13_2128, i_13_2173, i_13_2264, i_13_2362, i_13_2422, i_13_2423, i_13_2425, i_13_2426, i_13_2432, i_13_2452, i_13_2498, i_13_2747, i_13_3020, i_13_3035, i_13_3044, i_13_3100, i_13_3101, i_13_3127, i_13_3161, i_13_3214, i_13_3227, i_13_3375, i_13_3459, i_13_3461, i_13_3488, i_13_3577, i_13_3613, i_13_3700, i_13_3703, i_13_3756, i_13_3764, i_13_3784, i_13_3794, i_13_3844, i_13_3871, i_13_3872, i_13_4007, i_13_4081, i_13_4105, i_13_4117, i_13_4118, i_13_4159, i_13_4160, i_13_4163, i_13_4172, i_13_4295, i_13_4325, i_13_4348, i_13_4349, i_13_4474, o_13_506);
	kernel_13_507 k_13_507(i_13_46, i_13_102, i_13_163, i_13_312, i_13_321, i_13_322, i_13_342, i_13_379, i_13_408, i_13_442, i_13_604, i_13_624, i_13_625, i_13_657, i_13_671, i_13_680, i_13_757, i_13_846, i_13_883, i_13_885, i_13_936, i_13_1018, i_13_1147, i_13_1266, i_13_1362, i_13_1434, i_13_1498, i_13_1513, i_13_1515, i_13_1563, i_13_1582, i_13_1593, i_13_1594, i_13_1605, i_13_1701, i_13_1828, i_13_1944, i_13_2002, i_13_2012, i_13_2019, i_13_2025, i_13_2248, i_13_2268, i_13_2296, i_13_2463, i_13_2469, i_13_2498, i_13_2524, i_13_2601, i_13_2606, i_13_2673, i_13_2917, i_13_2966, i_13_2968, i_13_3003, i_13_3007, i_13_3030, i_13_3032, i_13_3099, i_13_3105, i_13_3214, i_13_3261, i_13_3325, i_13_3352, i_13_3400, i_13_3452, i_13_3483, i_13_3484, i_13_3541, i_13_3549, i_13_3566, i_13_3575, i_13_3699, i_13_3717, i_13_3730, i_13_3763, i_13_3765, i_13_3781, i_13_3784, i_13_3819, i_13_3823, i_13_3861, i_13_3898, i_13_3910, i_13_3970, i_13_4116, i_13_4159, i_13_4321, i_13_4335, i_13_4365, i_13_4366, i_13_4422, i_13_4448, i_13_4537, i_13_4558, i_13_4563, i_13_4564, i_13_4565, i_13_4599, i_13_4607, o_13_507);
	kernel_13_508 k_13_508(i_13_98, i_13_107, i_13_108, i_13_112, i_13_113, i_13_116, i_13_125, i_13_211, i_13_265, i_13_283, i_13_310, i_13_368, i_13_558, i_13_589, i_13_662, i_13_746, i_13_814, i_13_859, i_13_949, i_13_1017, i_13_1087, i_13_1088, i_13_1144, i_13_1219, i_13_1220, i_13_1474, i_13_1490, i_13_1520, i_13_1570, i_13_1574, i_13_1789, i_13_1790, i_13_1804, i_13_1841, i_13_1844, i_13_1915, i_13_1934, i_13_1993, i_13_2023, i_13_2173, i_13_2177, i_13_2276, i_13_2348, i_13_2421, i_13_2425, i_13_2434, i_13_2435, i_13_2438, i_13_2501, i_13_2542, i_13_2543, i_13_2561, i_13_2713, i_13_2716, i_13_2717, i_13_3047, i_13_3099, i_13_3146, i_13_3148, i_13_3149, i_13_3164, i_13_3167, i_13_3254, i_13_3344, i_13_3388, i_13_3413, i_13_3418, i_13_3419, i_13_3454, i_13_3455, i_13_3526, i_13_3527, i_13_3545, i_13_3640, i_13_3738, i_13_3742, i_13_3752, i_13_3766, i_13_3874, i_13_3875, i_13_3938, i_13_3994, i_13_4048, i_13_4077, i_13_4121, i_13_4163, i_13_4234, i_13_4252, i_13_4255, i_13_4264, i_13_4271, i_13_4309, i_13_4316, i_13_4328, i_13_4343, i_13_4354, i_13_4418, i_13_4518, i_13_4543, i_13_4544, o_13_508);
	kernel_13_509 k_13_509(i_13_31, i_13_32, i_13_35, i_13_94, i_13_95, i_13_97, i_13_98, i_13_113, i_13_115, i_13_116, i_13_121, i_13_122, i_13_178, i_13_229, i_13_232, i_13_260, i_13_313, i_13_386, i_13_448, i_13_449, i_13_538, i_13_539, i_13_565, i_13_607, i_13_730, i_13_733, i_13_800, i_13_868, i_13_943, i_13_953, i_13_1123, i_13_1193, i_13_1219, i_13_1313, i_13_1409, i_13_1440, i_13_1444, i_13_1445, i_13_1448, i_13_1628, i_13_1631, i_13_1787, i_13_1788, i_13_1799, i_13_1840, i_13_1841, i_13_1843, i_13_1844, i_13_1846, i_13_1912, i_13_1940, i_13_1943, i_13_2005, i_13_2021, i_13_2173, i_13_2176, i_13_2177, i_13_2279, i_13_2422, i_13_2425, i_13_2426, i_13_2428, i_13_2429, i_13_2447, i_13_2617, i_13_2677, i_13_2680, i_13_2681, i_13_2740, i_13_2749, i_13_2923, i_13_3002, i_13_3023, i_13_3037, i_13_3038, i_13_3064, i_13_3068, i_13_3146, i_13_3163, i_13_3164, i_13_3418, i_13_3419, i_13_3424, i_13_3425, i_13_3427, i_13_3428, i_13_3460, i_13_3487, i_13_3505, i_13_3580, i_13_3700, i_13_3865, i_13_3874, i_13_3875, i_13_4085, i_13_4351, i_13_4352, i_13_4453, i_13_4594, i_13_4598, o_13_509);
	kernel_13_510 k_13_510(i_13_130, i_13_170, i_13_187, i_13_188, i_13_202, i_13_266, i_13_269, i_13_311, i_13_446, i_13_464, i_13_583, i_13_644, i_13_646, i_13_647, i_13_697, i_13_815, i_13_817, i_13_818, i_13_844, i_13_845, i_13_916, i_13_931, i_13_950, i_13_986, i_13_1067, i_13_1070, i_13_1123, i_13_1124, i_13_1247, i_13_1274, i_13_1327, i_13_1331, i_13_1436, i_13_1490, i_13_1529, i_13_1601, i_13_1778, i_13_1807, i_13_1808, i_13_1835, i_13_1849, i_13_1850, i_13_1852, i_13_1853, i_13_1861, i_13_1933, i_13_1934, i_13_2050, i_13_2120, i_13_2149, i_13_2201, i_13_2213, i_13_2263, i_13_2264, i_13_2266, i_13_2267, i_13_2299, i_13_2345, i_13_2405, i_13_2407, i_13_2408, i_13_2410, i_13_2411, i_13_2446, i_13_2462, i_13_2545, i_13_2549, i_13_2600, i_13_2614, i_13_2698, i_13_2699, i_13_2749, i_13_2762, i_13_2795, i_13_2798, i_13_2899, i_13_2941, i_13_3004, i_13_3029, i_13_3094, i_13_3110, i_13_3112, i_13_3113, i_13_3292, i_13_3392, i_13_3478, i_13_3526, i_13_3553, i_13_3580, i_13_3821, i_13_3995, i_13_4066, i_13_4067, i_13_4171, i_13_4316, i_13_4318, i_13_4319, i_13_4342, i_13_4568, i_13_4598, o_13_510);
	kernel_13_511 k_13_511(i_13_43, i_13_48, i_13_69, i_13_70, i_13_79, i_13_141, i_13_244, i_13_305, i_13_321, i_13_322, i_13_328, i_13_411, i_13_417, i_13_448, i_13_522, i_13_570, i_13_589, i_13_591, i_13_598, i_13_615, i_13_784, i_13_924, i_13_937, i_13_951, i_13_1023, i_13_1105, i_13_1109, i_13_1122, i_13_1131, i_13_1132, i_13_1150, i_13_1230, i_13_1272, i_13_1284, i_13_1329, i_13_1402, i_13_1510, i_13_1511, i_13_1551, i_13_1644, i_13_1670, i_13_1722, i_13_1770, i_13_1797, i_13_1798, i_13_1806, i_13_1831, i_13_2028, i_13_2118, i_13_2265, i_13_2287, i_13_2296, i_13_2446, i_13_2461, i_13_2472, i_13_2473, i_13_2478, i_13_2505, i_13_2514, i_13_2560, i_13_2581, i_13_2677, i_13_2679, i_13_2680, i_13_2695, i_13_2698, i_13_2852, i_13_2999, i_13_3175, i_13_3264, i_13_3273, i_13_3274, i_13_3432, i_13_3478, i_13_3558, i_13_3561, i_13_3594, i_13_3640, i_13_3651, i_13_3702, i_13_3751, i_13_3759, i_13_3787, i_13_3822, i_13_3864, i_13_3899, i_13_3930, i_13_3940, i_13_4002, i_13_4036, i_13_4038, i_13_4174, i_13_4216, i_13_4407, i_13_4435, i_13_4448, i_13_4450, i_13_4513, i_13_4596, i_13_4597, o_13_511);
endmodule


module kernel_13_wrapper (input ap_clk, ap_rst, ap_ce, ap_start, ap_continue,
                        input [4607:0] in_reg,
                        output ap_idle, ap_done, ap_ready,
                        output out_reg_ap_vld,
                        output reg [511:0] out_reg);

  wire ce = ap_ce;
  reg i_13_0, i_13_1, i_13_2, i_13_3, i_13_4, i_13_5, i_13_6, i_13_7, i_13_8, i_13_9, i_13_10, i_13_11, i_13_12, i_13_13, i_13_14, i_13_15, i_13_16, i_13_17, i_13_18, i_13_19, i_13_20, i_13_21, i_13_22, i_13_23, i_13_24, i_13_25, i_13_26, i_13_27, i_13_28, i_13_29, i_13_30, i_13_31, i_13_32, i_13_33, i_13_34, i_13_35, i_13_36, i_13_37, i_13_38, i_13_39, i_13_40, i_13_41, i_13_42, i_13_43, i_13_44, i_13_45, i_13_46, i_13_47, i_13_48, i_13_49, i_13_50, i_13_51, i_13_52, i_13_53, i_13_54, i_13_55, i_13_56, i_13_57, i_13_58, i_13_59, i_13_60, i_13_61, i_13_62, i_13_63, i_13_64, i_13_65, i_13_66, i_13_67, i_13_68, i_13_69, i_13_70, i_13_71, i_13_72, i_13_73, i_13_74, i_13_75, i_13_76, i_13_77, i_13_78, i_13_79, i_13_80, i_13_81, i_13_82, i_13_83, i_13_84, i_13_85, i_13_86, i_13_87, i_13_88, i_13_89, i_13_90, i_13_91, i_13_92, i_13_93, i_13_94, i_13_95, i_13_96, i_13_97, i_13_98, i_13_99, i_13_100, i_13_101, i_13_102, i_13_103, i_13_104, i_13_105, i_13_106, i_13_107, i_13_108, i_13_109, i_13_110, i_13_111, i_13_112, i_13_113, i_13_114, i_13_115, i_13_116, i_13_117, i_13_118, i_13_119, i_13_120, i_13_121, i_13_122, i_13_123, i_13_124, i_13_125, i_13_126, i_13_127, i_13_128, i_13_129, i_13_130, i_13_131, i_13_132, i_13_133, i_13_134, i_13_135, i_13_136, i_13_137, i_13_138, i_13_139, i_13_140, i_13_141, i_13_142, i_13_143, i_13_144, i_13_145, i_13_146, i_13_147, i_13_148, i_13_149, i_13_150, i_13_151, i_13_152, i_13_153, i_13_154, i_13_155, i_13_156, i_13_157, i_13_158, i_13_159, i_13_160, i_13_161, i_13_162, i_13_163, i_13_164, i_13_165, i_13_166, i_13_167, i_13_168, i_13_169, i_13_170, i_13_171, i_13_172, i_13_173, i_13_174, i_13_175, i_13_176, i_13_177, i_13_178, i_13_179, i_13_180, i_13_181, i_13_182, i_13_183, i_13_184, i_13_185, i_13_186, i_13_187, i_13_188, i_13_189, i_13_190, i_13_191, i_13_192, i_13_193, i_13_194, i_13_195, i_13_196, i_13_197, i_13_198, i_13_199, i_13_200, i_13_201, i_13_202, i_13_203, i_13_204, i_13_205, i_13_206, i_13_207, i_13_208, i_13_209, i_13_210, i_13_211, i_13_212, i_13_213, i_13_214, i_13_215, i_13_216, i_13_217, i_13_218, i_13_219, i_13_220, i_13_221, i_13_222, i_13_223, i_13_224, i_13_225, i_13_226, i_13_227, i_13_228, i_13_229, i_13_230, i_13_231, i_13_232, i_13_233, i_13_234, i_13_235, i_13_236, i_13_237, i_13_238, i_13_239, i_13_240, i_13_241, i_13_242, i_13_243, i_13_244, i_13_245, i_13_246, i_13_247, i_13_248, i_13_249, i_13_250, i_13_251, i_13_252, i_13_253, i_13_254, i_13_255, i_13_256, i_13_257, i_13_258, i_13_259, i_13_260, i_13_261, i_13_262, i_13_263, i_13_264, i_13_265, i_13_266, i_13_267, i_13_268, i_13_269, i_13_270, i_13_271, i_13_272, i_13_273, i_13_274, i_13_275, i_13_276, i_13_277, i_13_278, i_13_279, i_13_280, i_13_281, i_13_282, i_13_283, i_13_284, i_13_285, i_13_286, i_13_287, i_13_288, i_13_289, i_13_290, i_13_291, i_13_292, i_13_293, i_13_294, i_13_295, i_13_296, i_13_297, i_13_298, i_13_299, i_13_300, i_13_301, i_13_302, i_13_303, i_13_304, i_13_305, i_13_306, i_13_307, i_13_308, i_13_309, i_13_310, i_13_311, i_13_312, i_13_313, i_13_314, i_13_315, i_13_316, i_13_317, i_13_318, i_13_319, i_13_320, i_13_321, i_13_322, i_13_323, i_13_324, i_13_325, i_13_326, i_13_327, i_13_328, i_13_329, i_13_330, i_13_331, i_13_332, i_13_333, i_13_334, i_13_335, i_13_336, i_13_337, i_13_338, i_13_339, i_13_340, i_13_341, i_13_342, i_13_343, i_13_344, i_13_345, i_13_346, i_13_347, i_13_348, i_13_349, i_13_350, i_13_351, i_13_352, i_13_353, i_13_354, i_13_355, i_13_356, i_13_357, i_13_358, i_13_359, i_13_360, i_13_361, i_13_362, i_13_363, i_13_364, i_13_365, i_13_366, i_13_367, i_13_368, i_13_369, i_13_370, i_13_371, i_13_372, i_13_373, i_13_374, i_13_375, i_13_376, i_13_377, i_13_378, i_13_379, i_13_380, i_13_381, i_13_382, i_13_383, i_13_384, i_13_385, i_13_386, i_13_387, i_13_388, i_13_389, i_13_390, i_13_391, i_13_392, i_13_393, i_13_394, i_13_395, i_13_396, i_13_397, i_13_398, i_13_399, i_13_400, i_13_401, i_13_402, i_13_403, i_13_404, i_13_405, i_13_406, i_13_407, i_13_408, i_13_409, i_13_410, i_13_411, i_13_412, i_13_413, i_13_414, i_13_415, i_13_416, i_13_417, i_13_418, i_13_419, i_13_420, i_13_421, i_13_422, i_13_423, i_13_424, i_13_425, i_13_426, i_13_427, i_13_428, i_13_429, i_13_430, i_13_431, i_13_432, i_13_433, i_13_434, i_13_435, i_13_436, i_13_437, i_13_438, i_13_439, i_13_440, i_13_441, i_13_442, i_13_443, i_13_444, i_13_445, i_13_446, i_13_447, i_13_448, i_13_449, i_13_450, i_13_451, i_13_452, i_13_453, i_13_454, i_13_455, i_13_456, i_13_457, i_13_458, i_13_459, i_13_460, i_13_461, i_13_462, i_13_463, i_13_464, i_13_465, i_13_466, i_13_467, i_13_468, i_13_469, i_13_470, i_13_471, i_13_472, i_13_473, i_13_474, i_13_475, i_13_476, i_13_477, i_13_478, i_13_479, i_13_480, i_13_481, i_13_482, i_13_483, i_13_484, i_13_485, i_13_486, i_13_487, i_13_488, i_13_489, i_13_490, i_13_491, i_13_492, i_13_493, i_13_494, i_13_495, i_13_496, i_13_497, i_13_498, i_13_499, i_13_500, i_13_501, i_13_502, i_13_503, i_13_504, i_13_505, i_13_506, i_13_507, i_13_508, i_13_509, i_13_510, i_13_511, i_13_512, i_13_513, i_13_514, i_13_515, i_13_516, i_13_517, i_13_518, i_13_519, i_13_520, i_13_521, i_13_522, i_13_523, i_13_524, i_13_525, i_13_526, i_13_527, i_13_528, i_13_529, i_13_530, i_13_531, i_13_532, i_13_533, i_13_534, i_13_535, i_13_536, i_13_537, i_13_538, i_13_539, i_13_540, i_13_541, i_13_542, i_13_543, i_13_544, i_13_545, i_13_546, i_13_547, i_13_548, i_13_549, i_13_550, i_13_551, i_13_552, i_13_553, i_13_554, i_13_555, i_13_556, i_13_557, i_13_558, i_13_559, i_13_560, i_13_561, i_13_562, i_13_563, i_13_564, i_13_565, i_13_566, i_13_567, i_13_568, i_13_569, i_13_570, i_13_571, i_13_572, i_13_573, i_13_574, i_13_575, i_13_576, i_13_577, i_13_578, i_13_579, i_13_580, i_13_581, i_13_582, i_13_583, i_13_584, i_13_585, i_13_586, i_13_587, i_13_588, i_13_589, i_13_590, i_13_591, i_13_592, i_13_593, i_13_594, i_13_595, i_13_596, i_13_597, i_13_598, i_13_599, i_13_600, i_13_601, i_13_602, i_13_603, i_13_604, i_13_605, i_13_606, i_13_607, i_13_608, i_13_609, i_13_610, i_13_611, i_13_612, i_13_613, i_13_614, i_13_615, i_13_616, i_13_617, i_13_618, i_13_619, i_13_620, i_13_621, i_13_622, i_13_623, i_13_624, i_13_625, i_13_626, i_13_627, i_13_628, i_13_629, i_13_630, i_13_631, i_13_632, i_13_633, i_13_634, i_13_635, i_13_636, i_13_637, i_13_638, i_13_639, i_13_640, i_13_641, i_13_642, i_13_643, i_13_644, i_13_645, i_13_646, i_13_647, i_13_648, i_13_649, i_13_650, i_13_651, i_13_652, i_13_653, i_13_654, i_13_655, i_13_656, i_13_657, i_13_658, i_13_659, i_13_660, i_13_661, i_13_662, i_13_663, i_13_664, i_13_665, i_13_666, i_13_667, i_13_668, i_13_669, i_13_670, i_13_671, i_13_672, i_13_673, i_13_674, i_13_675, i_13_676, i_13_677, i_13_678, i_13_679, i_13_680, i_13_681, i_13_682, i_13_683, i_13_684, i_13_685, i_13_686, i_13_687, i_13_688, i_13_689, i_13_690, i_13_691, i_13_692, i_13_693, i_13_694, i_13_695, i_13_696, i_13_697, i_13_698, i_13_699, i_13_700, i_13_701, i_13_702, i_13_703, i_13_704, i_13_705, i_13_706, i_13_707, i_13_708, i_13_709, i_13_710, i_13_711, i_13_712, i_13_713, i_13_714, i_13_715, i_13_716, i_13_717, i_13_718, i_13_719, i_13_720, i_13_721, i_13_722, i_13_723, i_13_724, i_13_725, i_13_726, i_13_727, i_13_728, i_13_729, i_13_730, i_13_731, i_13_732, i_13_733, i_13_734, i_13_735, i_13_736, i_13_737, i_13_738, i_13_739, i_13_740, i_13_741, i_13_742, i_13_743, i_13_744, i_13_745, i_13_746, i_13_747, i_13_748, i_13_749, i_13_750, i_13_751, i_13_752, i_13_753, i_13_754, i_13_755, i_13_756, i_13_757, i_13_758, i_13_759, i_13_760, i_13_761, i_13_762, i_13_763, i_13_764, i_13_765, i_13_766, i_13_767, i_13_768, i_13_769, i_13_770, i_13_771, i_13_772, i_13_773, i_13_774, i_13_775, i_13_776, i_13_777, i_13_778, i_13_779, i_13_780, i_13_781, i_13_782, i_13_783, i_13_784, i_13_785, i_13_786, i_13_787, i_13_788, i_13_789, i_13_790, i_13_791, i_13_792, i_13_793, i_13_794, i_13_795, i_13_796, i_13_797, i_13_798, i_13_799, i_13_800, i_13_801, i_13_802, i_13_803, i_13_804, i_13_805, i_13_806, i_13_807, i_13_808, i_13_809, i_13_810, i_13_811, i_13_812, i_13_813, i_13_814, i_13_815, i_13_816, i_13_817, i_13_818, i_13_819, i_13_820, i_13_821, i_13_822, i_13_823, i_13_824, i_13_825, i_13_826, i_13_827, i_13_828, i_13_829, i_13_830, i_13_831, i_13_832, i_13_833, i_13_834, i_13_835, i_13_836, i_13_837, i_13_838, i_13_839, i_13_840, i_13_841, i_13_842, i_13_843, i_13_844, i_13_845, i_13_846, i_13_847, i_13_848, i_13_849, i_13_850, i_13_851, i_13_852, i_13_853, i_13_854, i_13_855, i_13_856, i_13_857, i_13_858, i_13_859, i_13_860, i_13_861, i_13_862, i_13_863, i_13_864, i_13_865, i_13_866, i_13_867, i_13_868, i_13_869, i_13_870, i_13_871, i_13_872, i_13_873, i_13_874, i_13_875, i_13_876, i_13_877, i_13_878, i_13_879, i_13_880, i_13_881, i_13_882, i_13_883, i_13_884, i_13_885, i_13_886, i_13_887, i_13_888, i_13_889, i_13_890, i_13_891, i_13_892, i_13_893, i_13_894, i_13_895, i_13_896, i_13_897, i_13_898, i_13_899, i_13_900, i_13_901, i_13_902, i_13_903, i_13_904, i_13_905, i_13_906, i_13_907, i_13_908, i_13_909, i_13_910, i_13_911, i_13_912, i_13_913, i_13_914, i_13_915, i_13_916, i_13_917, i_13_918, i_13_919, i_13_920, i_13_921, i_13_922, i_13_923, i_13_924, i_13_925, i_13_926, i_13_927, i_13_928, i_13_929, i_13_930, i_13_931, i_13_932, i_13_933, i_13_934, i_13_935, i_13_936, i_13_937, i_13_938, i_13_939, i_13_940, i_13_941, i_13_942, i_13_943, i_13_944, i_13_945, i_13_946, i_13_947, i_13_948, i_13_949, i_13_950, i_13_951, i_13_952, i_13_953, i_13_954, i_13_955, i_13_956, i_13_957, i_13_958, i_13_959, i_13_960, i_13_961, i_13_962, i_13_963, i_13_964, i_13_965, i_13_966, i_13_967, i_13_968, i_13_969, i_13_970, i_13_971, i_13_972, i_13_973, i_13_974, i_13_975, i_13_976, i_13_977, i_13_978, i_13_979, i_13_980, i_13_981, i_13_982, i_13_983, i_13_984, i_13_985, i_13_986, i_13_987, i_13_988, i_13_989, i_13_990, i_13_991, i_13_992, i_13_993, i_13_994, i_13_995, i_13_996, i_13_997, i_13_998, i_13_999, i_13_1000, i_13_1001, i_13_1002, i_13_1003, i_13_1004, i_13_1005, i_13_1006, i_13_1007, i_13_1008, i_13_1009, i_13_1010, i_13_1011, i_13_1012, i_13_1013, i_13_1014, i_13_1015, i_13_1016, i_13_1017, i_13_1018, i_13_1019, i_13_1020, i_13_1021, i_13_1022, i_13_1023, i_13_1024, i_13_1025, i_13_1026, i_13_1027, i_13_1028, i_13_1029, i_13_1030, i_13_1031, i_13_1032, i_13_1033, i_13_1034, i_13_1035, i_13_1036, i_13_1037, i_13_1038, i_13_1039, i_13_1040, i_13_1041, i_13_1042, i_13_1043, i_13_1044, i_13_1045, i_13_1046, i_13_1047, i_13_1048, i_13_1049, i_13_1050, i_13_1051, i_13_1052, i_13_1053, i_13_1054, i_13_1055, i_13_1056, i_13_1057, i_13_1058, i_13_1059, i_13_1060, i_13_1061, i_13_1062, i_13_1063, i_13_1064, i_13_1065, i_13_1066, i_13_1067, i_13_1068, i_13_1069, i_13_1070, i_13_1071, i_13_1072, i_13_1073, i_13_1074, i_13_1075, i_13_1076, i_13_1077, i_13_1078, i_13_1079, i_13_1080, i_13_1081, i_13_1082, i_13_1083, i_13_1084, i_13_1085, i_13_1086, i_13_1087, i_13_1088, i_13_1089, i_13_1090, i_13_1091, i_13_1092, i_13_1093, i_13_1094, i_13_1095, i_13_1096, i_13_1097, i_13_1098, i_13_1099, i_13_1100, i_13_1101, i_13_1102, i_13_1103, i_13_1104, i_13_1105, i_13_1106, i_13_1107, i_13_1108, i_13_1109, i_13_1110, i_13_1111, i_13_1112, i_13_1113, i_13_1114, i_13_1115, i_13_1116, i_13_1117, i_13_1118, i_13_1119, i_13_1120, i_13_1121, i_13_1122, i_13_1123, i_13_1124, i_13_1125, i_13_1126, i_13_1127, i_13_1128, i_13_1129, i_13_1130, i_13_1131, i_13_1132, i_13_1133, i_13_1134, i_13_1135, i_13_1136, i_13_1137, i_13_1138, i_13_1139, i_13_1140, i_13_1141, i_13_1142, i_13_1143, i_13_1144, i_13_1145, i_13_1146, i_13_1147, i_13_1148, i_13_1149, i_13_1150, i_13_1151, i_13_1152, i_13_1153, i_13_1154, i_13_1155, i_13_1156, i_13_1157, i_13_1158, i_13_1159, i_13_1160, i_13_1161, i_13_1162, i_13_1163, i_13_1164, i_13_1165, i_13_1166, i_13_1167, i_13_1168, i_13_1169, i_13_1170, i_13_1171, i_13_1172, i_13_1173, i_13_1174, i_13_1175, i_13_1176, i_13_1177, i_13_1178, i_13_1179, i_13_1180, i_13_1181, i_13_1182, i_13_1183, i_13_1184, i_13_1185, i_13_1186, i_13_1187, i_13_1188, i_13_1189, i_13_1190, i_13_1191, i_13_1192, i_13_1193, i_13_1194, i_13_1195, i_13_1196, i_13_1197, i_13_1198, i_13_1199, i_13_1200, i_13_1201, i_13_1202, i_13_1203, i_13_1204, i_13_1205, i_13_1206, i_13_1207, i_13_1208, i_13_1209, i_13_1210, i_13_1211, i_13_1212, i_13_1213, i_13_1214, i_13_1215, i_13_1216, i_13_1217, i_13_1218, i_13_1219, i_13_1220, i_13_1221, i_13_1222, i_13_1223, i_13_1224, i_13_1225, i_13_1226, i_13_1227, i_13_1228, i_13_1229, i_13_1230, i_13_1231, i_13_1232, i_13_1233, i_13_1234, i_13_1235, i_13_1236, i_13_1237, i_13_1238, i_13_1239, i_13_1240, i_13_1241, i_13_1242, i_13_1243, i_13_1244, i_13_1245, i_13_1246, i_13_1247, i_13_1248, i_13_1249, i_13_1250, i_13_1251, i_13_1252, i_13_1253, i_13_1254, i_13_1255, i_13_1256, i_13_1257, i_13_1258, i_13_1259, i_13_1260, i_13_1261, i_13_1262, i_13_1263, i_13_1264, i_13_1265, i_13_1266, i_13_1267, i_13_1268, i_13_1269, i_13_1270, i_13_1271, i_13_1272, i_13_1273, i_13_1274, i_13_1275, i_13_1276, i_13_1277, i_13_1278, i_13_1279, i_13_1280, i_13_1281, i_13_1282, i_13_1283, i_13_1284, i_13_1285, i_13_1286, i_13_1287, i_13_1288, i_13_1289, i_13_1290, i_13_1291, i_13_1292, i_13_1293, i_13_1294, i_13_1295, i_13_1296, i_13_1297, i_13_1298, i_13_1299, i_13_1300, i_13_1301, i_13_1302, i_13_1303, i_13_1304, i_13_1305, i_13_1306, i_13_1307, i_13_1308, i_13_1309, i_13_1310, i_13_1311, i_13_1312, i_13_1313, i_13_1314, i_13_1315, i_13_1316, i_13_1317, i_13_1318, i_13_1319, i_13_1320, i_13_1321, i_13_1322, i_13_1323, i_13_1324, i_13_1325, i_13_1326, i_13_1327, i_13_1328, i_13_1329, i_13_1330, i_13_1331, i_13_1332, i_13_1333, i_13_1334, i_13_1335, i_13_1336, i_13_1337, i_13_1338, i_13_1339, i_13_1340, i_13_1341, i_13_1342, i_13_1343, i_13_1344, i_13_1345, i_13_1346, i_13_1347, i_13_1348, i_13_1349, i_13_1350, i_13_1351, i_13_1352, i_13_1353, i_13_1354, i_13_1355, i_13_1356, i_13_1357, i_13_1358, i_13_1359, i_13_1360, i_13_1361, i_13_1362, i_13_1363, i_13_1364, i_13_1365, i_13_1366, i_13_1367, i_13_1368, i_13_1369, i_13_1370, i_13_1371, i_13_1372, i_13_1373, i_13_1374, i_13_1375, i_13_1376, i_13_1377, i_13_1378, i_13_1379, i_13_1380, i_13_1381, i_13_1382, i_13_1383, i_13_1384, i_13_1385, i_13_1386, i_13_1387, i_13_1388, i_13_1389, i_13_1390, i_13_1391, i_13_1392, i_13_1393, i_13_1394, i_13_1395, i_13_1396, i_13_1397, i_13_1398, i_13_1399, i_13_1400, i_13_1401, i_13_1402, i_13_1403, i_13_1404, i_13_1405, i_13_1406, i_13_1407, i_13_1408, i_13_1409, i_13_1410, i_13_1411, i_13_1412, i_13_1413, i_13_1414, i_13_1415, i_13_1416, i_13_1417, i_13_1418, i_13_1419, i_13_1420, i_13_1421, i_13_1422, i_13_1423, i_13_1424, i_13_1425, i_13_1426, i_13_1427, i_13_1428, i_13_1429, i_13_1430, i_13_1431, i_13_1432, i_13_1433, i_13_1434, i_13_1435, i_13_1436, i_13_1437, i_13_1438, i_13_1439, i_13_1440, i_13_1441, i_13_1442, i_13_1443, i_13_1444, i_13_1445, i_13_1446, i_13_1447, i_13_1448, i_13_1449, i_13_1450, i_13_1451, i_13_1452, i_13_1453, i_13_1454, i_13_1455, i_13_1456, i_13_1457, i_13_1458, i_13_1459, i_13_1460, i_13_1461, i_13_1462, i_13_1463, i_13_1464, i_13_1465, i_13_1466, i_13_1467, i_13_1468, i_13_1469, i_13_1470, i_13_1471, i_13_1472, i_13_1473, i_13_1474, i_13_1475, i_13_1476, i_13_1477, i_13_1478, i_13_1479, i_13_1480, i_13_1481, i_13_1482, i_13_1483, i_13_1484, i_13_1485, i_13_1486, i_13_1487, i_13_1488, i_13_1489, i_13_1490, i_13_1491, i_13_1492, i_13_1493, i_13_1494, i_13_1495, i_13_1496, i_13_1497, i_13_1498, i_13_1499, i_13_1500, i_13_1501, i_13_1502, i_13_1503, i_13_1504, i_13_1505, i_13_1506, i_13_1507, i_13_1508, i_13_1509, i_13_1510, i_13_1511, i_13_1512, i_13_1513, i_13_1514, i_13_1515, i_13_1516, i_13_1517, i_13_1518, i_13_1519, i_13_1520, i_13_1521, i_13_1522, i_13_1523, i_13_1524, i_13_1525, i_13_1526, i_13_1527, i_13_1528, i_13_1529, i_13_1530, i_13_1531, i_13_1532, i_13_1533, i_13_1534, i_13_1535, i_13_1536, i_13_1537, i_13_1538, i_13_1539, i_13_1540, i_13_1541, i_13_1542, i_13_1543, i_13_1544, i_13_1545, i_13_1546, i_13_1547, i_13_1548, i_13_1549, i_13_1550, i_13_1551, i_13_1552, i_13_1553, i_13_1554, i_13_1555, i_13_1556, i_13_1557, i_13_1558, i_13_1559, i_13_1560, i_13_1561, i_13_1562, i_13_1563, i_13_1564, i_13_1565, i_13_1566, i_13_1567, i_13_1568, i_13_1569, i_13_1570, i_13_1571, i_13_1572, i_13_1573, i_13_1574, i_13_1575, i_13_1576, i_13_1577, i_13_1578, i_13_1579, i_13_1580, i_13_1581, i_13_1582, i_13_1583, i_13_1584, i_13_1585, i_13_1586, i_13_1587, i_13_1588, i_13_1589, i_13_1590, i_13_1591, i_13_1592, i_13_1593, i_13_1594, i_13_1595, i_13_1596, i_13_1597, i_13_1598, i_13_1599, i_13_1600, i_13_1601, i_13_1602, i_13_1603, i_13_1604, i_13_1605, i_13_1606, i_13_1607, i_13_1608, i_13_1609, i_13_1610, i_13_1611, i_13_1612, i_13_1613, i_13_1614, i_13_1615, i_13_1616, i_13_1617, i_13_1618, i_13_1619, i_13_1620, i_13_1621, i_13_1622, i_13_1623, i_13_1624, i_13_1625, i_13_1626, i_13_1627, i_13_1628, i_13_1629, i_13_1630, i_13_1631, i_13_1632, i_13_1633, i_13_1634, i_13_1635, i_13_1636, i_13_1637, i_13_1638, i_13_1639, i_13_1640, i_13_1641, i_13_1642, i_13_1643, i_13_1644, i_13_1645, i_13_1646, i_13_1647, i_13_1648, i_13_1649, i_13_1650, i_13_1651, i_13_1652, i_13_1653, i_13_1654, i_13_1655, i_13_1656, i_13_1657, i_13_1658, i_13_1659, i_13_1660, i_13_1661, i_13_1662, i_13_1663, i_13_1664, i_13_1665, i_13_1666, i_13_1667, i_13_1668, i_13_1669, i_13_1670, i_13_1671, i_13_1672, i_13_1673, i_13_1674, i_13_1675, i_13_1676, i_13_1677, i_13_1678, i_13_1679, i_13_1680, i_13_1681, i_13_1682, i_13_1683, i_13_1684, i_13_1685, i_13_1686, i_13_1687, i_13_1688, i_13_1689, i_13_1690, i_13_1691, i_13_1692, i_13_1693, i_13_1694, i_13_1695, i_13_1696, i_13_1697, i_13_1698, i_13_1699, i_13_1700, i_13_1701, i_13_1702, i_13_1703, i_13_1704, i_13_1705, i_13_1706, i_13_1707, i_13_1708, i_13_1709, i_13_1710, i_13_1711, i_13_1712, i_13_1713, i_13_1714, i_13_1715, i_13_1716, i_13_1717, i_13_1718, i_13_1719, i_13_1720, i_13_1721, i_13_1722, i_13_1723, i_13_1724, i_13_1725, i_13_1726, i_13_1727, i_13_1728, i_13_1729, i_13_1730, i_13_1731, i_13_1732, i_13_1733, i_13_1734, i_13_1735, i_13_1736, i_13_1737, i_13_1738, i_13_1739, i_13_1740, i_13_1741, i_13_1742, i_13_1743, i_13_1744, i_13_1745, i_13_1746, i_13_1747, i_13_1748, i_13_1749, i_13_1750, i_13_1751, i_13_1752, i_13_1753, i_13_1754, i_13_1755, i_13_1756, i_13_1757, i_13_1758, i_13_1759, i_13_1760, i_13_1761, i_13_1762, i_13_1763, i_13_1764, i_13_1765, i_13_1766, i_13_1767, i_13_1768, i_13_1769, i_13_1770, i_13_1771, i_13_1772, i_13_1773, i_13_1774, i_13_1775, i_13_1776, i_13_1777, i_13_1778, i_13_1779, i_13_1780, i_13_1781, i_13_1782, i_13_1783, i_13_1784, i_13_1785, i_13_1786, i_13_1787, i_13_1788, i_13_1789, i_13_1790, i_13_1791, i_13_1792, i_13_1793, i_13_1794, i_13_1795, i_13_1796, i_13_1797, i_13_1798, i_13_1799, i_13_1800, i_13_1801, i_13_1802, i_13_1803, i_13_1804, i_13_1805, i_13_1806, i_13_1807, i_13_1808, i_13_1809, i_13_1810, i_13_1811, i_13_1812, i_13_1813, i_13_1814, i_13_1815, i_13_1816, i_13_1817, i_13_1818, i_13_1819, i_13_1820, i_13_1821, i_13_1822, i_13_1823, i_13_1824, i_13_1825, i_13_1826, i_13_1827, i_13_1828, i_13_1829, i_13_1830, i_13_1831, i_13_1832, i_13_1833, i_13_1834, i_13_1835, i_13_1836, i_13_1837, i_13_1838, i_13_1839, i_13_1840, i_13_1841, i_13_1842, i_13_1843, i_13_1844, i_13_1845, i_13_1846, i_13_1847, i_13_1848, i_13_1849, i_13_1850, i_13_1851, i_13_1852, i_13_1853, i_13_1854, i_13_1855, i_13_1856, i_13_1857, i_13_1858, i_13_1859, i_13_1860, i_13_1861, i_13_1862, i_13_1863, i_13_1864, i_13_1865, i_13_1866, i_13_1867, i_13_1868, i_13_1869, i_13_1870, i_13_1871, i_13_1872, i_13_1873, i_13_1874, i_13_1875, i_13_1876, i_13_1877, i_13_1878, i_13_1879, i_13_1880, i_13_1881, i_13_1882, i_13_1883, i_13_1884, i_13_1885, i_13_1886, i_13_1887, i_13_1888, i_13_1889, i_13_1890, i_13_1891, i_13_1892, i_13_1893, i_13_1894, i_13_1895, i_13_1896, i_13_1897, i_13_1898, i_13_1899, i_13_1900, i_13_1901, i_13_1902, i_13_1903, i_13_1904, i_13_1905, i_13_1906, i_13_1907, i_13_1908, i_13_1909, i_13_1910, i_13_1911, i_13_1912, i_13_1913, i_13_1914, i_13_1915, i_13_1916, i_13_1917, i_13_1918, i_13_1919, i_13_1920, i_13_1921, i_13_1922, i_13_1923, i_13_1924, i_13_1925, i_13_1926, i_13_1927, i_13_1928, i_13_1929, i_13_1930, i_13_1931, i_13_1932, i_13_1933, i_13_1934, i_13_1935, i_13_1936, i_13_1937, i_13_1938, i_13_1939, i_13_1940, i_13_1941, i_13_1942, i_13_1943, i_13_1944, i_13_1945, i_13_1946, i_13_1947, i_13_1948, i_13_1949, i_13_1950, i_13_1951, i_13_1952, i_13_1953, i_13_1954, i_13_1955, i_13_1956, i_13_1957, i_13_1958, i_13_1959, i_13_1960, i_13_1961, i_13_1962, i_13_1963, i_13_1964, i_13_1965, i_13_1966, i_13_1967, i_13_1968, i_13_1969, i_13_1970, i_13_1971, i_13_1972, i_13_1973, i_13_1974, i_13_1975, i_13_1976, i_13_1977, i_13_1978, i_13_1979, i_13_1980, i_13_1981, i_13_1982, i_13_1983, i_13_1984, i_13_1985, i_13_1986, i_13_1987, i_13_1988, i_13_1989, i_13_1990, i_13_1991, i_13_1992, i_13_1993, i_13_1994, i_13_1995, i_13_1996, i_13_1997, i_13_1998, i_13_1999, i_13_2000, i_13_2001, i_13_2002, i_13_2003, i_13_2004, i_13_2005, i_13_2006, i_13_2007, i_13_2008, i_13_2009, i_13_2010, i_13_2011, i_13_2012, i_13_2013, i_13_2014, i_13_2015, i_13_2016, i_13_2017, i_13_2018, i_13_2019, i_13_2020, i_13_2021, i_13_2022, i_13_2023, i_13_2024, i_13_2025, i_13_2026, i_13_2027, i_13_2028, i_13_2029, i_13_2030, i_13_2031, i_13_2032, i_13_2033, i_13_2034, i_13_2035, i_13_2036, i_13_2037, i_13_2038, i_13_2039, i_13_2040, i_13_2041, i_13_2042, i_13_2043, i_13_2044, i_13_2045, i_13_2046, i_13_2047, i_13_2048, i_13_2049, i_13_2050, i_13_2051, i_13_2052, i_13_2053, i_13_2054, i_13_2055, i_13_2056, i_13_2057, i_13_2058, i_13_2059, i_13_2060, i_13_2061, i_13_2062, i_13_2063, i_13_2064, i_13_2065, i_13_2066, i_13_2067, i_13_2068, i_13_2069, i_13_2070, i_13_2071, i_13_2072, i_13_2073, i_13_2074, i_13_2075, i_13_2076, i_13_2077, i_13_2078, i_13_2079, i_13_2080, i_13_2081, i_13_2082, i_13_2083, i_13_2084, i_13_2085, i_13_2086, i_13_2087, i_13_2088, i_13_2089, i_13_2090, i_13_2091, i_13_2092, i_13_2093, i_13_2094, i_13_2095, i_13_2096, i_13_2097, i_13_2098, i_13_2099, i_13_2100, i_13_2101, i_13_2102, i_13_2103, i_13_2104, i_13_2105, i_13_2106, i_13_2107, i_13_2108, i_13_2109, i_13_2110, i_13_2111, i_13_2112, i_13_2113, i_13_2114, i_13_2115, i_13_2116, i_13_2117, i_13_2118, i_13_2119, i_13_2120, i_13_2121, i_13_2122, i_13_2123, i_13_2124, i_13_2125, i_13_2126, i_13_2127, i_13_2128, i_13_2129, i_13_2130, i_13_2131, i_13_2132, i_13_2133, i_13_2134, i_13_2135, i_13_2136, i_13_2137, i_13_2138, i_13_2139, i_13_2140, i_13_2141, i_13_2142, i_13_2143, i_13_2144, i_13_2145, i_13_2146, i_13_2147, i_13_2148, i_13_2149, i_13_2150, i_13_2151, i_13_2152, i_13_2153, i_13_2154, i_13_2155, i_13_2156, i_13_2157, i_13_2158, i_13_2159, i_13_2160, i_13_2161, i_13_2162, i_13_2163, i_13_2164, i_13_2165, i_13_2166, i_13_2167, i_13_2168, i_13_2169, i_13_2170, i_13_2171, i_13_2172, i_13_2173, i_13_2174, i_13_2175, i_13_2176, i_13_2177, i_13_2178, i_13_2179, i_13_2180, i_13_2181, i_13_2182, i_13_2183, i_13_2184, i_13_2185, i_13_2186, i_13_2187, i_13_2188, i_13_2189, i_13_2190, i_13_2191, i_13_2192, i_13_2193, i_13_2194, i_13_2195, i_13_2196, i_13_2197, i_13_2198, i_13_2199, i_13_2200, i_13_2201, i_13_2202, i_13_2203, i_13_2204, i_13_2205, i_13_2206, i_13_2207, i_13_2208, i_13_2209, i_13_2210, i_13_2211, i_13_2212, i_13_2213, i_13_2214, i_13_2215, i_13_2216, i_13_2217, i_13_2218, i_13_2219, i_13_2220, i_13_2221, i_13_2222, i_13_2223, i_13_2224, i_13_2225, i_13_2226, i_13_2227, i_13_2228, i_13_2229, i_13_2230, i_13_2231, i_13_2232, i_13_2233, i_13_2234, i_13_2235, i_13_2236, i_13_2237, i_13_2238, i_13_2239, i_13_2240, i_13_2241, i_13_2242, i_13_2243, i_13_2244, i_13_2245, i_13_2246, i_13_2247, i_13_2248, i_13_2249, i_13_2250, i_13_2251, i_13_2252, i_13_2253, i_13_2254, i_13_2255, i_13_2256, i_13_2257, i_13_2258, i_13_2259, i_13_2260, i_13_2261, i_13_2262, i_13_2263, i_13_2264, i_13_2265, i_13_2266, i_13_2267, i_13_2268, i_13_2269, i_13_2270, i_13_2271, i_13_2272, i_13_2273, i_13_2274, i_13_2275, i_13_2276, i_13_2277, i_13_2278, i_13_2279, i_13_2280, i_13_2281, i_13_2282, i_13_2283, i_13_2284, i_13_2285, i_13_2286, i_13_2287, i_13_2288, i_13_2289, i_13_2290, i_13_2291, i_13_2292, i_13_2293, i_13_2294, i_13_2295, i_13_2296, i_13_2297, i_13_2298, i_13_2299, i_13_2300, i_13_2301, i_13_2302, i_13_2303, i_13_2304, i_13_2305, i_13_2306, i_13_2307, i_13_2308, i_13_2309, i_13_2310, i_13_2311, i_13_2312, i_13_2313, i_13_2314, i_13_2315, i_13_2316, i_13_2317, i_13_2318, i_13_2319, i_13_2320, i_13_2321, i_13_2322, i_13_2323, i_13_2324, i_13_2325, i_13_2326, i_13_2327, i_13_2328, i_13_2329, i_13_2330, i_13_2331, i_13_2332, i_13_2333, i_13_2334, i_13_2335, i_13_2336, i_13_2337, i_13_2338, i_13_2339, i_13_2340, i_13_2341, i_13_2342, i_13_2343, i_13_2344, i_13_2345, i_13_2346, i_13_2347, i_13_2348, i_13_2349, i_13_2350, i_13_2351, i_13_2352, i_13_2353, i_13_2354, i_13_2355, i_13_2356, i_13_2357, i_13_2358, i_13_2359, i_13_2360, i_13_2361, i_13_2362, i_13_2363, i_13_2364, i_13_2365, i_13_2366, i_13_2367, i_13_2368, i_13_2369, i_13_2370, i_13_2371, i_13_2372, i_13_2373, i_13_2374, i_13_2375, i_13_2376, i_13_2377, i_13_2378, i_13_2379, i_13_2380, i_13_2381, i_13_2382, i_13_2383, i_13_2384, i_13_2385, i_13_2386, i_13_2387, i_13_2388, i_13_2389, i_13_2390, i_13_2391, i_13_2392, i_13_2393, i_13_2394, i_13_2395, i_13_2396, i_13_2397, i_13_2398, i_13_2399, i_13_2400, i_13_2401, i_13_2402, i_13_2403, i_13_2404, i_13_2405, i_13_2406, i_13_2407, i_13_2408, i_13_2409, i_13_2410, i_13_2411, i_13_2412, i_13_2413, i_13_2414, i_13_2415, i_13_2416, i_13_2417, i_13_2418, i_13_2419, i_13_2420, i_13_2421, i_13_2422, i_13_2423, i_13_2424, i_13_2425, i_13_2426, i_13_2427, i_13_2428, i_13_2429, i_13_2430, i_13_2431, i_13_2432, i_13_2433, i_13_2434, i_13_2435, i_13_2436, i_13_2437, i_13_2438, i_13_2439, i_13_2440, i_13_2441, i_13_2442, i_13_2443, i_13_2444, i_13_2445, i_13_2446, i_13_2447, i_13_2448, i_13_2449, i_13_2450, i_13_2451, i_13_2452, i_13_2453, i_13_2454, i_13_2455, i_13_2456, i_13_2457, i_13_2458, i_13_2459, i_13_2460, i_13_2461, i_13_2462, i_13_2463, i_13_2464, i_13_2465, i_13_2466, i_13_2467, i_13_2468, i_13_2469, i_13_2470, i_13_2471, i_13_2472, i_13_2473, i_13_2474, i_13_2475, i_13_2476, i_13_2477, i_13_2478, i_13_2479, i_13_2480, i_13_2481, i_13_2482, i_13_2483, i_13_2484, i_13_2485, i_13_2486, i_13_2487, i_13_2488, i_13_2489, i_13_2490, i_13_2491, i_13_2492, i_13_2493, i_13_2494, i_13_2495, i_13_2496, i_13_2497, i_13_2498, i_13_2499, i_13_2500, i_13_2501, i_13_2502, i_13_2503, i_13_2504, i_13_2505, i_13_2506, i_13_2507, i_13_2508, i_13_2509, i_13_2510, i_13_2511, i_13_2512, i_13_2513, i_13_2514, i_13_2515, i_13_2516, i_13_2517, i_13_2518, i_13_2519, i_13_2520, i_13_2521, i_13_2522, i_13_2523, i_13_2524, i_13_2525, i_13_2526, i_13_2527, i_13_2528, i_13_2529, i_13_2530, i_13_2531, i_13_2532, i_13_2533, i_13_2534, i_13_2535, i_13_2536, i_13_2537, i_13_2538, i_13_2539, i_13_2540, i_13_2541, i_13_2542, i_13_2543, i_13_2544, i_13_2545, i_13_2546, i_13_2547, i_13_2548, i_13_2549, i_13_2550, i_13_2551, i_13_2552, i_13_2553, i_13_2554, i_13_2555, i_13_2556, i_13_2557, i_13_2558, i_13_2559, i_13_2560, i_13_2561, i_13_2562, i_13_2563, i_13_2564, i_13_2565, i_13_2566, i_13_2567, i_13_2568, i_13_2569, i_13_2570, i_13_2571, i_13_2572, i_13_2573, i_13_2574, i_13_2575, i_13_2576, i_13_2577, i_13_2578, i_13_2579, i_13_2580, i_13_2581, i_13_2582, i_13_2583, i_13_2584, i_13_2585, i_13_2586, i_13_2587, i_13_2588, i_13_2589, i_13_2590, i_13_2591, i_13_2592, i_13_2593, i_13_2594, i_13_2595, i_13_2596, i_13_2597, i_13_2598, i_13_2599, i_13_2600, i_13_2601, i_13_2602, i_13_2603, i_13_2604, i_13_2605, i_13_2606, i_13_2607, i_13_2608, i_13_2609, i_13_2610, i_13_2611, i_13_2612, i_13_2613, i_13_2614, i_13_2615, i_13_2616, i_13_2617, i_13_2618, i_13_2619, i_13_2620, i_13_2621, i_13_2622, i_13_2623, i_13_2624, i_13_2625, i_13_2626, i_13_2627, i_13_2628, i_13_2629, i_13_2630, i_13_2631, i_13_2632, i_13_2633, i_13_2634, i_13_2635, i_13_2636, i_13_2637, i_13_2638, i_13_2639, i_13_2640, i_13_2641, i_13_2642, i_13_2643, i_13_2644, i_13_2645, i_13_2646, i_13_2647, i_13_2648, i_13_2649, i_13_2650, i_13_2651, i_13_2652, i_13_2653, i_13_2654, i_13_2655, i_13_2656, i_13_2657, i_13_2658, i_13_2659, i_13_2660, i_13_2661, i_13_2662, i_13_2663, i_13_2664, i_13_2665, i_13_2666, i_13_2667, i_13_2668, i_13_2669, i_13_2670, i_13_2671, i_13_2672, i_13_2673, i_13_2674, i_13_2675, i_13_2676, i_13_2677, i_13_2678, i_13_2679, i_13_2680, i_13_2681, i_13_2682, i_13_2683, i_13_2684, i_13_2685, i_13_2686, i_13_2687, i_13_2688, i_13_2689, i_13_2690, i_13_2691, i_13_2692, i_13_2693, i_13_2694, i_13_2695, i_13_2696, i_13_2697, i_13_2698, i_13_2699, i_13_2700, i_13_2701, i_13_2702, i_13_2703, i_13_2704, i_13_2705, i_13_2706, i_13_2707, i_13_2708, i_13_2709, i_13_2710, i_13_2711, i_13_2712, i_13_2713, i_13_2714, i_13_2715, i_13_2716, i_13_2717, i_13_2718, i_13_2719, i_13_2720, i_13_2721, i_13_2722, i_13_2723, i_13_2724, i_13_2725, i_13_2726, i_13_2727, i_13_2728, i_13_2729, i_13_2730, i_13_2731, i_13_2732, i_13_2733, i_13_2734, i_13_2735, i_13_2736, i_13_2737, i_13_2738, i_13_2739, i_13_2740, i_13_2741, i_13_2742, i_13_2743, i_13_2744, i_13_2745, i_13_2746, i_13_2747, i_13_2748, i_13_2749, i_13_2750, i_13_2751, i_13_2752, i_13_2753, i_13_2754, i_13_2755, i_13_2756, i_13_2757, i_13_2758, i_13_2759, i_13_2760, i_13_2761, i_13_2762, i_13_2763, i_13_2764, i_13_2765, i_13_2766, i_13_2767, i_13_2768, i_13_2769, i_13_2770, i_13_2771, i_13_2772, i_13_2773, i_13_2774, i_13_2775, i_13_2776, i_13_2777, i_13_2778, i_13_2779, i_13_2780, i_13_2781, i_13_2782, i_13_2783, i_13_2784, i_13_2785, i_13_2786, i_13_2787, i_13_2788, i_13_2789, i_13_2790, i_13_2791, i_13_2792, i_13_2793, i_13_2794, i_13_2795, i_13_2796, i_13_2797, i_13_2798, i_13_2799, i_13_2800, i_13_2801, i_13_2802, i_13_2803, i_13_2804, i_13_2805, i_13_2806, i_13_2807, i_13_2808, i_13_2809, i_13_2810, i_13_2811, i_13_2812, i_13_2813, i_13_2814, i_13_2815, i_13_2816, i_13_2817, i_13_2818, i_13_2819, i_13_2820, i_13_2821, i_13_2822, i_13_2823, i_13_2824, i_13_2825, i_13_2826, i_13_2827, i_13_2828, i_13_2829, i_13_2830, i_13_2831, i_13_2832, i_13_2833, i_13_2834, i_13_2835, i_13_2836, i_13_2837, i_13_2838, i_13_2839, i_13_2840, i_13_2841, i_13_2842, i_13_2843, i_13_2844, i_13_2845, i_13_2846, i_13_2847, i_13_2848, i_13_2849, i_13_2850, i_13_2851, i_13_2852, i_13_2853, i_13_2854, i_13_2855, i_13_2856, i_13_2857, i_13_2858, i_13_2859, i_13_2860, i_13_2861, i_13_2862, i_13_2863, i_13_2864, i_13_2865, i_13_2866, i_13_2867, i_13_2868, i_13_2869, i_13_2870, i_13_2871, i_13_2872, i_13_2873, i_13_2874, i_13_2875, i_13_2876, i_13_2877, i_13_2878, i_13_2879, i_13_2880, i_13_2881, i_13_2882, i_13_2883, i_13_2884, i_13_2885, i_13_2886, i_13_2887, i_13_2888, i_13_2889, i_13_2890, i_13_2891, i_13_2892, i_13_2893, i_13_2894, i_13_2895, i_13_2896, i_13_2897, i_13_2898, i_13_2899, i_13_2900, i_13_2901, i_13_2902, i_13_2903, i_13_2904, i_13_2905, i_13_2906, i_13_2907, i_13_2908, i_13_2909, i_13_2910, i_13_2911, i_13_2912, i_13_2913, i_13_2914, i_13_2915, i_13_2916, i_13_2917, i_13_2918, i_13_2919, i_13_2920, i_13_2921, i_13_2922, i_13_2923, i_13_2924, i_13_2925, i_13_2926, i_13_2927, i_13_2928, i_13_2929, i_13_2930, i_13_2931, i_13_2932, i_13_2933, i_13_2934, i_13_2935, i_13_2936, i_13_2937, i_13_2938, i_13_2939, i_13_2940, i_13_2941, i_13_2942, i_13_2943, i_13_2944, i_13_2945, i_13_2946, i_13_2947, i_13_2948, i_13_2949, i_13_2950, i_13_2951, i_13_2952, i_13_2953, i_13_2954, i_13_2955, i_13_2956, i_13_2957, i_13_2958, i_13_2959, i_13_2960, i_13_2961, i_13_2962, i_13_2963, i_13_2964, i_13_2965, i_13_2966, i_13_2967, i_13_2968, i_13_2969, i_13_2970, i_13_2971, i_13_2972, i_13_2973, i_13_2974, i_13_2975, i_13_2976, i_13_2977, i_13_2978, i_13_2979, i_13_2980, i_13_2981, i_13_2982, i_13_2983, i_13_2984, i_13_2985, i_13_2986, i_13_2987, i_13_2988, i_13_2989, i_13_2990, i_13_2991, i_13_2992, i_13_2993, i_13_2994, i_13_2995, i_13_2996, i_13_2997, i_13_2998, i_13_2999, i_13_3000, i_13_3001, i_13_3002, i_13_3003, i_13_3004, i_13_3005, i_13_3006, i_13_3007, i_13_3008, i_13_3009, i_13_3010, i_13_3011, i_13_3012, i_13_3013, i_13_3014, i_13_3015, i_13_3016, i_13_3017, i_13_3018, i_13_3019, i_13_3020, i_13_3021, i_13_3022, i_13_3023, i_13_3024, i_13_3025, i_13_3026, i_13_3027, i_13_3028, i_13_3029, i_13_3030, i_13_3031, i_13_3032, i_13_3033, i_13_3034, i_13_3035, i_13_3036, i_13_3037, i_13_3038, i_13_3039, i_13_3040, i_13_3041, i_13_3042, i_13_3043, i_13_3044, i_13_3045, i_13_3046, i_13_3047, i_13_3048, i_13_3049, i_13_3050, i_13_3051, i_13_3052, i_13_3053, i_13_3054, i_13_3055, i_13_3056, i_13_3057, i_13_3058, i_13_3059, i_13_3060, i_13_3061, i_13_3062, i_13_3063, i_13_3064, i_13_3065, i_13_3066, i_13_3067, i_13_3068, i_13_3069, i_13_3070, i_13_3071, i_13_3072, i_13_3073, i_13_3074, i_13_3075, i_13_3076, i_13_3077, i_13_3078, i_13_3079, i_13_3080, i_13_3081, i_13_3082, i_13_3083, i_13_3084, i_13_3085, i_13_3086, i_13_3087, i_13_3088, i_13_3089, i_13_3090, i_13_3091, i_13_3092, i_13_3093, i_13_3094, i_13_3095, i_13_3096, i_13_3097, i_13_3098, i_13_3099, i_13_3100, i_13_3101, i_13_3102, i_13_3103, i_13_3104, i_13_3105, i_13_3106, i_13_3107, i_13_3108, i_13_3109, i_13_3110, i_13_3111, i_13_3112, i_13_3113, i_13_3114, i_13_3115, i_13_3116, i_13_3117, i_13_3118, i_13_3119, i_13_3120, i_13_3121, i_13_3122, i_13_3123, i_13_3124, i_13_3125, i_13_3126, i_13_3127, i_13_3128, i_13_3129, i_13_3130, i_13_3131, i_13_3132, i_13_3133, i_13_3134, i_13_3135, i_13_3136, i_13_3137, i_13_3138, i_13_3139, i_13_3140, i_13_3141, i_13_3142, i_13_3143, i_13_3144, i_13_3145, i_13_3146, i_13_3147, i_13_3148, i_13_3149, i_13_3150, i_13_3151, i_13_3152, i_13_3153, i_13_3154, i_13_3155, i_13_3156, i_13_3157, i_13_3158, i_13_3159, i_13_3160, i_13_3161, i_13_3162, i_13_3163, i_13_3164, i_13_3165, i_13_3166, i_13_3167, i_13_3168, i_13_3169, i_13_3170, i_13_3171, i_13_3172, i_13_3173, i_13_3174, i_13_3175, i_13_3176, i_13_3177, i_13_3178, i_13_3179, i_13_3180, i_13_3181, i_13_3182, i_13_3183, i_13_3184, i_13_3185, i_13_3186, i_13_3187, i_13_3188, i_13_3189, i_13_3190, i_13_3191, i_13_3192, i_13_3193, i_13_3194, i_13_3195, i_13_3196, i_13_3197, i_13_3198, i_13_3199, i_13_3200, i_13_3201, i_13_3202, i_13_3203, i_13_3204, i_13_3205, i_13_3206, i_13_3207, i_13_3208, i_13_3209, i_13_3210, i_13_3211, i_13_3212, i_13_3213, i_13_3214, i_13_3215, i_13_3216, i_13_3217, i_13_3218, i_13_3219, i_13_3220, i_13_3221, i_13_3222, i_13_3223, i_13_3224, i_13_3225, i_13_3226, i_13_3227, i_13_3228, i_13_3229, i_13_3230, i_13_3231, i_13_3232, i_13_3233, i_13_3234, i_13_3235, i_13_3236, i_13_3237, i_13_3238, i_13_3239, i_13_3240, i_13_3241, i_13_3242, i_13_3243, i_13_3244, i_13_3245, i_13_3246, i_13_3247, i_13_3248, i_13_3249, i_13_3250, i_13_3251, i_13_3252, i_13_3253, i_13_3254, i_13_3255, i_13_3256, i_13_3257, i_13_3258, i_13_3259, i_13_3260, i_13_3261, i_13_3262, i_13_3263, i_13_3264, i_13_3265, i_13_3266, i_13_3267, i_13_3268, i_13_3269, i_13_3270, i_13_3271, i_13_3272, i_13_3273, i_13_3274, i_13_3275, i_13_3276, i_13_3277, i_13_3278, i_13_3279, i_13_3280, i_13_3281, i_13_3282, i_13_3283, i_13_3284, i_13_3285, i_13_3286, i_13_3287, i_13_3288, i_13_3289, i_13_3290, i_13_3291, i_13_3292, i_13_3293, i_13_3294, i_13_3295, i_13_3296, i_13_3297, i_13_3298, i_13_3299, i_13_3300, i_13_3301, i_13_3302, i_13_3303, i_13_3304, i_13_3305, i_13_3306, i_13_3307, i_13_3308, i_13_3309, i_13_3310, i_13_3311, i_13_3312, i_13_3313, i_13_3314, i_13_3315, i_13_3316, i_13_3317, i_13_3318, i_13_3319, i_13_3320, i_13_3321, i_13_3322, i_13_3323, i_13_3324, i_13_3325, i_13_3326, i_13_3327, i_13_3328, i_13_3329, i_13_3330, i_13_3331, i_13_3332, i_13_3333, i_13_3334, i_13_3335, i_13_3336, i_13_3337, i_13_3338, i_13_3339, i_13_3340, i_13_3341, i_13_3342, i_13_3343, i_13_3344, i_13_3345, i_13_3346, i_13_3347, i_13_3348, i_13_3349, i_13_3350, i_13_3351, i_13_3352, i_13_3353, i_13_3354, i_13_3355, i_13_3356, i_13_3357, i_13_3358, i_13_3359, i_13_3360, i_13_3361, i_13_3362, i_13_3363, i_13_3364, i_13_3365, i_13_3366, i_13_3367, i_13_3368, i_13_3369, i_13_3370, i_13_3371, i_13_3372, i_13_3373, i_13_3374, i_13_3375, i_13_3376, i_13_3377, i_13_3378, i_13_3379, i_13_3380, i_13_3381, i_13_3382, i_13_3383, i_13_3384, i_13_3385, i_13_3386, i_13_3387, i_13_3388, i_13_3389, i_13_3390, i_13_3391, i_13_3392, i_13_3393, i_13_3394, i_13_3395, i_13_3396, i_13_3397, i_13_3398, i_13_3399, i_13_3400, i_13_3401, i_13_3402, i_13_3403, i_13_3404, i_13_3405, i_13_3406, i_13_3407, i_13_3408, i_13_3409, i_13_3410, i_13_3411, i_13_3412, i_13_3413, i_13_3414, i_13_3415, i_13_3416, i_13_3417, i_13_3418, i_13_3419, i_13_3420, i_13_3421, i_13_3422, i_13_3423, i_13_3424, i_13_3425, i_13_3426, i_13_3427, i_13_3428, i_13_3429, i_13_3430, i_13_3431, i_13_3432, i_13_3433, i_13_3434, i_13_3435, i_13_3436, i_13_3437, i_13_3438, i_13_3439, i_13_3440, i_13_3441, i_13_3442, i_13_3443, i_13_3444, i_13_3445, i_13_3446, i_13_3447, i_13_3448, i_13_3449, i_13_3450, i_13_3451, i_13_3452, i_13_3453, i_13_3454, i_13_3455, i_13_3456, i_13_3457, i_13_3458, i_13_3459, i_13_3460, i_13_3461, i_13_3462, i_13_3463, i_13_3464, i_13_3465, i_13_3466, i_13_3467, i_13_3468, i_13_3469, i_13_3470, i_13_3471, i_13_3472, i_13_3473, i_13_3474, i_13_3475, i_13_3476, i_13_3477, i_13_3478, i_13_3479, i_13_3480, i_13_3481, i_13_3482, i_13_3483, i_13_3484, i_13_3485, i_13_3486, i_13_3487, i_13_3488, i_13_3489, i_13_3490, i_13_3491, i_13_3492, i_13_3493, i_13_3494, i_13_3495, i_13_3496, i_13_3497, i_13_3498, i_13_3499, i_13_3500, i_13_3501, i_13_3502, i_13_3503, i_13_3504, i_13_3505, i_13_3506, i_13_3507, i_13_3508, i_13_3509, i_13_3510, i_13_3511, i_13_3512, i_13_3513, i_13_3514, i_13_3515, i_13_3516, i_13_3517, i_13_3518, i_13_3519, i_13_3520, i_13_3521, i_13_3522, i_13_3523, i_13_3524, i_13_3525, i_13_3526, i_13_3527, i_13_3528, i_13_3529, i_13_3530, i_13_3531, i_13_3532, i_13_3533, i_13_3534, i_13_3535, i_13_3536, i_13_3537, i_13_3538, i_13_3539, i_13_3540, i_13_3541, i_13_3542, i_13_3543, i_13_3544, i_13_3545, i_13_3546, i_13_3547, i_13_3548, i_13_3549, i_13_3550, i_13_3551, i_13_3552, i_13_3553, i_13_3554, i_13_3555, i_13_3556, i_13_3557, i_13_3558, i_13_3559, i_13_3560, i_13_3561, i_13_3562, i_13_3563, i_13_3564, i_13_3565, i_13_3566, i_13_3567, i_13_3568, i_13_3569, i_13_3570, i_13_3571, i_13_3572, i_13_3573, i_13_3574, i_13_3575, i_13_3576, i_13_3577, i_13_3578, i_13_3579, i_13_3580, i_13_3581, i_13_3582, i_13_3583, i_13_3584, i_13_3585, i_13_3586, i_13_3587, i_13_3588, i_13_3589, i_13_3590, i_13_3591, i_13_3592, i_13_3593, i_13_3594, i_13_3595, i_13_3596, i_13_3597, i_13_3598, i_13_3599, i_13_3600, i_13_3601, i_13_3602, i_13_3603, i_13_3604, i_13_3605, i_13_3606, i_13_3607, i_13_3608, i_13_3609, i_13_3610, i_13_3611, i_13_3612, i_13_3613, i_13_3614, i_13_3615, i_13_3616, i_13_3617, i_13_3618, i_13_3619, i_13_3620, i_13_3621, i_13_3622, i_13_3623, i_13_3624, i_13_3625, i_13_3626, i_13_3627, i_13_3628, i_13_3629, i_13_3630, i_13_3631, i_13_3632, i_13_3633, i_13_3634, i_13_3635, i_13_3636, i_13_3637, i_13_3638, i_13_3639, i_13_3640, i_13_3641, i_13_3642, i_13_3643, i_13_3644, i_13_3645, i_13_3646, i_13_3647, i_13_3648, i_13_3649, i_13_3650, i_13_3651, i_13_3652, i_13_3653, i_13_3654, i_13_3655, i_13_3656, i_13_3657, i_13_3658, i_13_3659, i_13_3660, i_13_3661, i_13_3662, i_13_3663, i_13_3664, i_13_3665, i_13_3666, i_13_3667, i_13_3668, i_13_3669, i_13_3670, i_13_3671, i_13_3672, i_13_3673, i_13_3674, i_13_3675, i_13_3676, i_13_3677, i_13_3678, i_13_3679, i_13_3680, i_13_3681, i_13_3682, i_13_3683, i_13_3684, i_13_3685, i_13_3686, i_13_3687, i_13_3688, i_13_3689, i_13_3690, i_13_3691, i_13_3692, i_13_3693, i_13_3694, i_13_3695, i_13_3696, i_13_3697, i_13_3698, i_13_3699, i_13_3700, i_13_3701, i_13_3702, i_13_3703, i_13_3704, i_13_3705, i_13_3706, i_13_3707, i_13_3708, i_13_3709, i_13_3710, i_13_3711, i_13_3712, i_13_3713, i_13_3714, i_13_3715, i_13_3716, i_13_3717, i_13_3718, i_13_3719, i_13_3720, i_13_3721, i_13_3722, i_13_3723, i_13_3724, i_13_3725, i_13_3726, i_13_3727, i_13_3728, i_13_3729, i_13_3730, i_13_3731, i_13_3732, i_13_3733, i_13_3734, i_13_3735, i_13_3736, i_13_3737, i_13_3738, i_13_3739, i_13_3740, i_13_3741, i_13_3742, i_13_3743, i_13_3744, i_13_3745, i_13_3746, i_13_3747, i_13_3748, i_13_3749, i_13_3750, i_13_3751, i_13_3752, i_13_3753, i_13_3754, i_13_3755, i_13_3756, i_13_3757, i_13_3758, i_13_3759, i_13_3760, i_13_3761, i_13_3762, i_13_3763, i_13_3764, i_13_3765, i_13_3766, i_13_3767, i_13_3768, i_13_3769, i_13_3770, i_13_3771, i_13_3772, i_13_3773, i_13_3774, i_13_3775, i_13_3776, i_13_3777, i_13_3778, i_13_3779, i_13_3780, i_13_3781, i_13_3782, i_13_3783, i_13_3784, i_13_3785, i_13_3786, i_13_3787, i_13_3788, i_13_3789, i_13_3790, i_13_3791, i_13_3792, i_13_3793, i_13_3794, i_13_3795, i_13_3796, i_13_3797, i_13_3798, i_13_3799, i_13_3800, i_13_3801, i_13_3802, i_13_3803, i_13_3804, i_13_3805, i_13_3806, i_13_3807, i_13_3808, i_13_3809, i_13_3810, i_13_3811, i_13_3812, i_13_3813, i_13_3814, i_13_3815, i_13_3816, i_13_3817, i_13_3818, i_13_3819, i_13_3820, i_13_3821, i_13_3822, i_13_3823, i_13_3824, i_13_3825, i_13_3826, i_13_3827, i_13_3828, i_13_3829, i_13_3830, i_13_3831, i_13_3832, i_13_3833, i_13_3834, i_13_3835, i_13_3836, i_13_3837, i_13_3838, i_13_3839, i_13_3840, i_13_3841, i_13_3842, i_13_3843, i_13_3844, i_13_3845, i_13_3846, i_13_3847, i_13_3848, i_13_3849, i_13_3850, i_13_3851, i_13_3852, i_13_3853, i_13_3854, i_13_3855, i_13_3856, i_13_3857, i_13_3858, i_13_3859, i_13_3860, i_13_3861, i_13_3862, i_13_3863, i_13_3864, i_13_3865, i_13_3866, i_13_3867, i_13_3868, i_13_3869, i_13_3870, i_13_3871, i_13_3872, i_13_3873, i_13_3874, i_13_3875, i_13_3876, i_13_3877, i_13_3878, i_13_3879, i_13_3880, i_13_3881, i_13_3882, i_13_3883, i_13_3884, i_13_3885, i_13_3886, i_13_3887, i_13_3888, i_13_3889, i_13_3890, i_13_3891, i_13_3892, i_13_3893, i_13_3894, i_13_3895, i_13_3896, i_13_3897, i_13_3898, i_13_3899, i_13_3900, i_13_3901, i_13_3902, i_13_3903, i_13_3904, i_13_3905, i_13_3906, i_13_3907, i_13_3908, i_13_3909, i_13_3910, i_13_3911, i_13_3912, i_13_3913, i_13_3914, i_13_3915, i_13_3916, i_13_3917, i_13_3918, i_13_3919, i_13_3920, i_13_3921, i_13_3922, i_13_3923, i_13_3924, i_13_3925, i_13_3926, i_13_3927, i_13_3928, i_13_3929, i_13_3930, i_13_3931, i_13_3932, i_13_3933, i_13_3934, i_13_3935, i_13_3936, i_13_3937, i_13_3938, i_13_3939, i_13_3940, i_13_3941, i_13_3942, i_13_3943, i_13_3944, i_13_3945, i_13_3946, i_13_3947, i_13_3948, i_13_3949, i_13_3950, i_13_3951, i_13_3952, i_13_3953, i_13_3954, i_13_3955, i_13_3956, i_13_3957, i_13_3958, i_13_3959, i_13_3960, i_13_3961, i_13_3962, i_13_3963, i_13_3964, i_13_3965, i_13_3966, i_13_3967, i_13_3968, i_13_3969, i_13_3970, i_13_3971, i_13_3972, i_13_3973, i_13_3974, i_13_3975, i_13_3976, i_13_3977, i_13_3978, i_13_3979, i_13_3980, i_13_3981, i_13_3982, i_13_3983, i_13_3984, i_13_3985, i_13_3986, i_13_3987, i_13_3988, i_13_3989, i_13_3990, i_13_3991, i_13_3992, i_13_3993, i_13_3994, i_13_3995, i_13_3996, i_13_3997, i_13_3998, i_13_3999, i_13_4000, i_13_4001, i_13_4002, i_13_4003, i_13_4004, i_13_4005, i_13_4006, i_13_4007, i_13_4008, i_13_4009, i_13_4010, i_13_4011, i_13_4012, i_13_4013, i_13_4014, i_13_4015, i_13_4016, i_13_4017, i_13_4018, i_13_4019, i_13_4020, i_13_4021, i_13_4022, i_13_4023, i_13_4024, i_13_4025, i_13_4026, i_13_4027, i_13_4028, i_13_4029, i_13_4030, i_13_4031, i_13_4032, i_13_4033, i_13_4034, i_13_4035, i_13_4036, i_13_4037, i_13_4038, i_13_4039, i_13_4040, i_13_4041, i_13_4042, i_13_4043, i_13_4044, i_13_4045, i_13_4046, i_13_4047, i_13_4048, i_13_4049, i_13_4050, i_13_4051, i_13_4052, i_13_4053, i_13_4054, i_13_4055, i_13_4056, i_13_4057, i_13_4058, i_13_4059, i_13_4060, i_13_4061, i_13_4062, i_13_4063, i_13_4064, i_13_4065, i_13_4066, i_13_4067, i_13_4068, i_13_4069, i_13_4070, i_13_4071, i_13_4072, i_13_4073, i_13_4074, i_13_4075, i_13_4076, i_13_4077, i_13_4078, i_13_4079, i_13_4080, i_13_4081, i_13_4082, i_13_4083, i_13_4084, i_13_4085, i_13_4086, i_13_4087, i_13_4088, i_13_4089, i_13_4090, i_13_4091, i_13_4092, i_13_4093, i_13_4094, i_13_4095, i_13_4096, i_13_4097, i_13_4098, i_13_4099, i_13_4100, i_13_4101, i_13_4102, i_13_4103, i_13_4104, i_13_4105, i_13_4106, i_13_4107, i_13_4108, i_13_4109, i_13_4110, i_13_4111, i_13_4112, i_13_4113, i_13_4114, i_13_4115, i_13_4116, i_13_4117, i_13_4118, i_13_4119, i_13_4120, i_13_4121, i_13_4122, i_13_4123, i_13_4124, i_13_4125, i_13_4126, i_13_4127, i_13_4128, i_13_4129, i_13_4130, i_13_4131, i_13_4132, i_13_4133, i_13_4134, i_13_4135, i_13_4136, i_13_4137, i_13_4138, i_13_4139, i_13_4140, i_13_4141, i_13_4142, i_13_4143, i_13_4144, i_13_4145, i_13_4146, i_13_4147, i_13_4148, i_13_4149, i_13_4150, i_13_4151, i_13_4152, i_13_4153, i_13_4154, i_13_4155, i_13_4156, i_13_4157, i_13_4158, i_13_4159, i_13_4160, i_13_4161, i_13_4162, i_13_4163, i_13_4164, i_13_4165, i_13_4166, i_13_4167, i_13_4168, i_13_4169, i_13_4170, i_13_4171, i_13_4172, i_13_4173, i_13_4174, i_13_4175, i_13_4176, i_13_4177, i_13_4178, i_13_4179, i_13_4180, i_13_4181, i_13_4182, i_13_4183, i_13_4184, i_13_4185, i_13_4186, i_13_4187, i_13_4188, i_13_4189, i_13_4190, i_13_4191, i_13_4192, i_13_4193, i_13_4194, i_13_4195, i_13_4196, i_13_4197, i_13_4198, i_13_4199, i_13_4200, i_13_4201, i_13_4202, i_13_4203, i_13_4204, i_13_4205, i_13_4206, i_13_4207, i_13_4208, i_13_4209, i_13_4210, i_13_4211, i_13_4212, i_13_4213, i_13_4214, i_13_4215, i_13_4216, i_13_4217, i_13_4218, i_13_4219, i_13_4220, i_13_4221, i_13_4222, i_13_4223, i_13_4224, i_13_4225, i_13_4226, i_13_4227, i_13_4228, i_13_4229, i_13_4230, i_13_4231, i_13_4232, i_13_4233, i_13_4234, i_13_4235, i_13_4236, i_13_4237, i_13_4238, i_13_4239, i_13_4240, i_13_4241, i_13_4242, i_13_4243, i_13_4244, i_13_4245, i_13_4246, i_13_4247, i_13_4248, i_13_4249, i_13_4250, i_13_4251, i_13_4252, i_13_4253, i_13_4254, i_13_4255, i_13_4256, i_13_4257, i_13_4258, i_13_4259, i_13_4260, i_13_4261, i_13_4262, i_13_4263, i_13_4264, i_13_4265, i_13_4266, i_13_4267, i_13_4268, i_13_4269, i_13_4270, i_13_4271, i_13_4272, i_13_4273, i_13_4274, i_13_4275, i_13_4276, i_13_4277, i_13_4278, i_13_4279, i_13_4280, i_13_4281, i_13_4282, i_13_4283, i_13_4284, i_13_4285, i_13_4286, i_13_4287, i_13_4288, i_13_4289, i_13_4290, i_13_4291, i_13_4292, i_13_4293, i_13_4294, i_13_4295, i_13_4296, i_13_4297, i_13_4298, i_13_4299, i_13_4300, i_13_4301, i_13_4302, i_13_4303, i_13_4304, i_13_4305, i_13_4306, i_13_4307, i_13_4308, i_13_4309, i_13_4310, i_13_4311, i_13_4312, i_13_4313, i_13_4314, i_13_4315, i_13_4316, i_13_4317, i_13_4318, i_13_4319, i_13_4320, i_13_4321, i_13_4322, i_13_4323, i_13_4324, i_13_4325, i_13_4326, i_13_4327, i_13_4328, i_13_4329, i_13_4330, i_13_4331, i_13_4332, i_13_4333, i_13_4334, i_13_4335, i_13_4336, i_13_4337, i_13_4338, i_13_4339, i_13_4340, i_13_4341, i_13_4342, i_13_4343, i_13_4344, i_13_4345, i_13_4346, i_13_4347, i_13_4348, i_13_4349, i_13_4350, i_13_4351, i_13_4352, i_13_4353, i_13_4354, i_13_4355, i_13_4356, i_13_4357, i_13_4358, i_13_4359, i_13_4360, i_13_4361, i_13_4362, i_13_4363, i_13_4364, i_13_4365, i_13_4366, i_13_4367, i_13_4368, i_13_4369, i_13_4370, i_13_4371, i_13_4372, i_13_4373, i_13_4374, i_13_4375, i_13_4376, i_13_4377, i_13_4378, i_13_4379, i_13_4380, i_13_4381, i_13_4382, i_13_4383, i_13_4384, i_13_4385, i_13_4386, i_13_4387, i_13_4388, i_13_4389, i_13_4390, i_13_4391, i_13_4392, i_13_4393, i_13_4394, i_13_4395, i_13_4396, i_13_4397, i_13_4398, i_13_4399, i_13_4400, i_13_4401, i_13_4402, i_13_4403, i_13_4404, i_13_4405, i_13_4406, i_13_4407, i_13_4408, i_13_4409, i_13_4410, i_13_4411, i_13_4412, i_13_4413, i_13_4414, i_13_4415, i_13_4416, i_13_4417, i_13_4418, i_13_4419, i_13_4420, i_13_4421, i_13_4422, i_13_4423, i_13_4424, i_13_4425, i_13_4426, i_13_4427, i_13_4428, i_13_4429, i_13_4430, i_13_4431, i_13_4432, i_13_4433, i_13_4434, i_13_4435, i_13_4436, i_13_4437, i_13_4438, i_13_4439, i_13_4440, i_13_4441, i_13_4442, i_13_4443, i_13_4444, i_13_4445, i_13_4446, i_13_4447, i_13_4448, i_13_4449, i_13_4450, i_13_4451, i_13_4452, i_13_4453, i_13_4454, i_13_4455, i_13_4456, i_13_4457, i_13_4458, i_13_4459, i_13_4460, i_13_4461, i_13_4462, i_13_4463, i_13_4464, i_13_4465, i_13_4466, i_13_4467, i_13_4468, i_13_4469, i_13_4470, i_13_4471, i_13_4472, i_13_4473, i_13_4474, i_13_4475, i_13_4476, i_13_4477, i_13_4478, i_13_4479, i_13_4480, i_13_4481, i_13_4482, i_13_4483, i_13_4484, i_13_4485, i_13_4486, i_13_4487, i_13_4488, i_13_4489, i_13_4490, i_13_4491, i_13_4492, i_13_4493, i_13_4494, i_13_4495, i_13_4496, i_13_4497, i_13_4498, i_13_4499, i_13_4500, i_13_4501, i_13_4502, i_13_4503, i_13_4504, i_13_4505, i_13_4506, i_13_4507, i_13_4508, i_13_4509, i_13_4510, i_13_4511, i_13_4512, i_13_4513, i_13_4514, i_13_4515, i_13_4516, i_13_4517, i_13_4518, i_13_4519, i_13_4520, i_13_4521, i_13_4522, i_13_4523, i_13_4524, i_13_4525, i_13_4526, i_13_4527, i_13_4528, i_13_4529, i_13_4530, i_13_4531, i_13_4532, i_13_4533, i_13_4534, i_13_4535, i_13_4536, i_13_4537, i_13_4538, i_13_4539, i_13_4540, i_13_4541, i_13_4542, i_13_4543, i_13_4544, i_13_4545, i_13_4546, i_13_4547, i_13_4548, i_13_4549, i_13_4550, i_13_4551, i_13_4552, i_13_4553, i_13_4554, i_13_4555, i_13_4556, i_13_4557, i_13_4558, i_13_4559, i_13_4560, i_13_4561, i_13_4562, i_13_4563, i_13_4564, i_13_4565, i_13_4566, i_13_4567, i_13_4568, i_13_4569, i_13_4570, i_13_4571, i_13_4572, i_13_4573, i_13_4574, i_13_4575, i_13_4576, i_13_4577, i_13_4578, i_13_4579, i_13_4580, i_13_4581, i_13_4582, i_13_4583, i_13_4584, i_13_4585, i_13_4586, i_13_4587, i_13_4588, i_13_4589, i_13_4590, i_13_4591, i_13_4592, i_13_4593, i_13_4594, i_13_4595, i_13_4596, i_13_4597, i_13_4598, i_13_4599, i_13_4600, i_13_4601, i_13_4602, i_13_4603, i_13_4604, i_13_4605, i_13_4606, i_13_4607;
  reg dly1, dly2;
  wire o_13_0, o_13_1, o_13_2, o_13_3, o_13_4, o_13_5, o_13_6, o_13_7, o_13_8, o_13_9, o_13_10, o_13_11, o_13_12, o_13_13, o_13_14, o_13_15, o_13_16, o_13_17, o_13_18, o_13_19, o_13_20, o_13_21, o_13_22, o_13_23, o_13_24, o_13_25, o_13_26, o_13_27, o_13_28, o_13_29, o_13_30, o_13_31, o_13_32, o_13_33, o_13_34, o_13_35, o_13_36, o_13_37, o_13_38, o_13_39, o_13_40, o_13_41, o_13_42, o_13_43, o_13_44, o_13_45, o_13_46, o_13_47, o_13_48, o_13_49, o_13_50, o_13_51, o_13_52, o_13_53, o_13_54, o_13_55, o_13_56, o_13_57, o_13_58, o_13_59, o_13_60, o_13_61, o_13_62, o_13_63, o_13_64, o_13_65, o_13_66, o_13_67, o_13_68, o_13_69, o_13_70, o_13_71, o_13_72, o_13_73, o_13_74, o_13_75, o_13_76, o_13_77, o_13_78, o_13_79, o_13_80, o_13_81, o_13_82, o_13_83, o_13_84, o_13_85, o_13_86, o_13_87, o_13_88, o_13_89, o_13_90, o_13_91, o_13_92, o_13_93, o_13_94, o_13_95, o_13_96, o_13_97, o_13_98, o_13_99, o_13_100, o_13_101, o_13_102, o_13_103, o_13_104, o_13_105, o_13_106, o_13_107, o_13_108, o_13_109, o_13_110, o_13_111, o_13_112, o_13_113, o_13_114, o_13_115, o_13_116, o_13_117, o_13_118, o_13_119, o_13_120, o_13_121, o_13_122, o_13_123, o_13_124, o_13_125, o_13_126, o_13_127, o_13_128, o_13_129, o_13_130, o_13_131, o_13_132, o_13_133, o_13_134, o_13_135, o_13_136, o_13_137, o_13_138, o_13_139, o_13_140, o_13_141, o_13_142, o_13_143, o_13_144, o_13_145, o_13_146, o_13_147, o_13_148, o_13_149, o_13_150, o_13_151, o_13_152, o_13_153, o_13_154, o_13_155, o_13_156, o_13_157, o_13_158, o_13_159, o_13_160, o_13_161, o_13_162, o_13_163, o_13_164, o_13_165, o_13_166, o_13_167, o_13_168, o_13_169, o_13_170, o_13_171, o_13_172, o_13_173, o_13_174, o_13_175, o_13_176, o_13_177, o_13_178, o_13_179, o_13_180, o_13_181, o_13_182, o_13_183, o_13_184, o_13_185, o_13_186, o_13_187, o_13_188, o_13_189, o_13_190, o_13_191, o_13_192, o_13_193, o_13_194, o_13_195, o_13_196, o_13_197, o_13_198, o_13_199, o_13_200, o_13_201, o_13_202, o_13_203, o_13_204, o_13_205, o_13_206, o_13_207, o_13_208, o_13_209, o_13_210, o_13_211, o_13_212, o_13_213, o_13_214, o_13_215, o_13_216, o_13_217, o_13_218, o_13_219, o_13_220, o_13_221, o_13_222, o_13_223, o_13_224, o_13_225, o_13_226, o_13_227, o_13_228, o_13_229, o_13_230, o_13_231, o_13_232, o_13_233, o_13_234, o_13_235, o_13_236, o_13_237, o_13_238, o_13_239, o_13_240, o_13_241, o_13_242, o_13_243, o_13_244, o_13_245, o_13_246, o_13_247, o_13_248, o_13_249, o_13_250, o_13_251, o_13_252, o_13_253, o_13_254, o_13_255, o_13_256, o_13_257, o_13_258, o_13_259, o_13_260, o_13_261, o_13_262, o_13_263, o_13_264, o_13_265, o_13_266, o_13_267, o_13_268, o_13_269, o_13_270, o_13_271, o_13_272, o_13_273, o_13_274, o_13_275, o_13_276, o_13_277, o_13_278, o_13_279, o_13_280, o_13_281, o_13_282, o_13_283, o_13_284, o_13_285, o_13_286, o_13_287, o_13_288, o_13_289, o_13_290, o_13_291, o_13_292, o_13_293, o_13_294, o_13_295, o_13_296, o_13_297, o_13_298, o_13_299, o_13_300, o_13_301, o_13_302, o_13_303, o_13_304, o_13_305, o_13_306, o_13_307, o_13_308, o_13_309, o_13_310, o_13_311, o_13_312, o_13_313, o_13_314, o_13_315, o_13_316, o_13_317, o_13_318, o_13_319, o_13_320, o_13_321, o_13_322, o_13_323, o_13_324, o_13_325, o_13_326, o_13_327, o_13_328, o_13_329, o_13_330, o_13_331, o_13_332, o_13_333, o_13_334, o_13_335, o_13_336, o_13_337, o_13_338, o_13_339, o_13_340, o_13_341, o_13_342, o_13_343, o_13_344, o_13_345, o_13_346, o_13_347, o_13_348, o_13_349, o_13_350, o_13_351, o_13_352, o_13_353, o_13_354, o_13_355, o_13_356, o_13_357, o_13_358, o_13_359, o_13_360, o_13_361, o_13_362, o_13_363, o_13_364, o_13_365, o_13_366, o_13_367, o_13_368, o_13_369, o_13_370, o_13_371, o_13_372, o_13_373, o_13_374, o_13_375, o_13_376, o_13_377, o_13_378, o_13_379, o_13_380, o_13_381, o_13_382, o_13_383, o_13_384, o_13_385, o_13_386, o_13_387, o_13_388, o_13_389, o_13_390, o_13_391, o_13_392, o_13_393, o_13_394, o_13_395, o_13_396, o_13_397, o_13_398, o_13_399, o_13_400, o_13_401, o_13_402, o_13_403, o_13_404, o_13_405, o_13_406, o_13_407, o_13_408, o_13_409, o_13_410, o_13_411, o_13_412, o_13_413, o_13_414, o_13_415, o_13_416, o_13_417, o_13_418, o_13_419, o_13_420, o_13_421, o_13_422, o_13_423, o_13_424, o_13_425, o_13_426, o_13_427, o_13_428, o_13_429, o_13_430, o_13_431, o_13_432, o_13_433, o_13_434, o_13_435, o_13_436, o_13_437, o_13_438, o_13_439, o_13_440, o_13_441, o_13_442, o_13_443, o_13_444, o_13_445, o_13_446, o_13_447, o_13_448, o_13_449, o_13_450, o_13_451, o_13_452, o_13_453, o_13_454, o_13_455, o_13_456, o_13_457, o_13_458, o_13_459, o_13_460, o_13_461, o_13_462, o_13_463, o_13_464, o_13_465, o_13_466, o_13_467, o_13_468, o_13_469, o_13_470, o_13_471, o_13_472, o_13_473, o_13_474, o_13_475, o_13_476, o_13_477, o_13_478, o_13_479, o_13_480, o_13_481, o_13_482, o_13_483, o_13_484, o_13_485, o_13_486, o_13_487, o_13_488, o_13_489, o_13_490, o_13_491, o_13_492, o_13_493, o_13_494, o_13_495, o_13_496, o_13_497, o_13_498, o_13_499, o_13_500, o_13_501, o_13_502, o_13_503, o_13_504, o_13_505, o_13_506, o_13_507, o_13_508, o_13_509, o_13_510, o_13_511;

  kernel_13 kernel_nulla( i_13_0, i_13_1, i_13_2, i_13_3, i_13_4, i_13_5, i_13_6, i_13_7, i_13_8, i_13_9, i_13_10, i_13_11, i_13_12, i_13_13, i_13_14, i_13_15, i_13_16, i_13_17, i_13_18, i_13_19, i_13_20, i_13_21, i_13_22, i_13_23, i_13_24, i_13_25, i_13_26, i_13_27, i_13_28, i_13_29, i_13_30, i_13_31, i_13_32, i_13_33, i_13_34, i_13_35, i_13_36, i_13_37, i_13_38, i_13_39, i_13_40, i_13_41, i_13_42, i_13_43, i_13_44, i_13_45, i_13_46, i_13_47, i_13_48, i_13_49, i_13_50, i_13_51, i_13_52, i_13_53, i_13_54, i_13_55, i_13_56, i_13_57, i_13_58, i_13_59, i_13_60, i_13_61, i_13_62, i_13_63, i_13_64, i_13_65, i_13_66, i_13_67, i_13_68, i_13_69, i_13_70, i_13_71, i_13_72, i_13_73, i_13_74, i_13_75, i_13_76, i_13_77, i_13_78, i_13_79, i_13_80, i_13_81, i_13_82, i_13_83, i_13_84, i_13_85, i_13_86, i_13_87, i_13_88, i_13_89, i_13_90, i_13_91, i_13_92, i_13_93, i_13_94, i_13_95, i_13_96, i_13_97, i_13_98, i_13_99, i_13_100, i_13_101, i_13_102, i_13_103, i_13_104, i_13_105, i_13_106, i_13_107, i_13_108, i_13_109, i_13_110, i_13_111, i_13_112, i_13_113, i_13_114, i_13_115, i_13_116, i_13_117, i_13_118, i_13_119, i_13_120, i_13_121, i_13_122, i_13_123, i_13_124, i_13_125, i_13_126, i_13_127, i_13_128, i_13_129, i_13_130, i_13_131, i_13_132, i_13_133, i_13_134, i_13_135, i_13_136, i_13_137, i_13_138, i_13_139, i_13_140, i_13_141, i_13_142, i_13_143, i_13_144, i_13_145, i_13_146, i_13_147, i_13_148, i_13_149, i_13_150, i_13_151, i_13_152, i_13_153, i_13_154, i_13_155, i_13_156, i_13_157, i_13_158, i_13_159, i_13_160, i_13_161, i_13_162, i_13_163, i_13_164, i_13_165, i_13_166, i_13_167, i_13_168, i_13_169, i_13_170, i_13_171, i_13_172, i_13_173, i_13_174, i_13_175, i_13_176, i_13_177, i_13_178, i_13_179, i_13_180, i_13_181, i_13_182, i_13_183, i_13_184, i_13_185, i_13_186, i_13_187, i_13_188, i_13_189, i_13_190, i_13_191, i_13_192, i_13_193, i_13_194, i_13_195, i_13_196, i_13_197, i_13_198, i_13_199, i_13_200, i_13_201, i_13_202, i_13_203, i_13_204, i_13_205, i_13_206, i_13_207, i_13_208, i_13_209, i_13_210, i_13_211, i_13_212, i_13_213, i_13_214, i_13_215, i_13_216, i_13_217, i_13_218, i_13_219, i_13_220, i_13_221, i_13_222, i_13_223, i_13_224, i_13_225, i_13_226, i_13_227, i_13_228, i_13_229, i_13_230, i_13_231, i_13_232, i_13_233, i_13_234, i_13_235, i_13_236, i_13_237, i_13_238, i_13_239, i_13_240, i_13_241, i_13_242, i_13_243, i_13_244, i_13_245, i_13_246, i_13_247, i_13_248, i_13_249, i_13_250, i_13_251, i_13_252, i_13_253, i_13_254, i_13_255, i_13_256, i_13_257, i_13_258, i_13_259, i_13_260, i_13_261, i_13_262, i_13_263, i_13_264, i_13_265, i_13_266, i_13_267, i_13_268, i_13_269, i_13_270, i_13_271, i_13_272, i_13_273, i_13_274, i_13_275, i_13_276, i_13_277, i_13_278, i_13_279, i_13_280, i_13_281, i_13_282, i_13_283, i_13_284, i_13_285, i_13_286, i_13_287, i_13_288, i_13_289, i_13_290, i_13_291, i_13_292, i_13_293, i_13_294, i_13_295, i_13_296, i_13_297, i_13_298, i_13_299, i_13_300, i_13_301, i_13_302, i_13_303, i_13_304, i_13_305, i_13_306, i_13_307, i_13_308, i_13_309, i_13_310, i_13_311, i_13_312, i_13_313, i_13_314, i_13_315, i_13_316, i_13_317, i_13_318, i_13_319, i_13_320, i_13_321, i_13_322, i_13_323, i_13_324, i_13_325, i_13_326, i_13_327, i_13_328, i_13_329, i_13_330, i_13_331, i_13_332, i_13_333, i_13_334, i_13_335, i_13_336, i_13_337, i_13_338, i_13_339, i_13_340, i_13_341, i_13_342, i_13_343, i_13_344, i_13_345, i_13_346, i_13_347, i_13_348, i_13_349, i_13_350, i_13_351, i_13_352, i_13_353, i_13_354, i_13_355, i_13_356, i_13_357, i_13_358, i_13_359, i_13_360, i_13_361, i_13_362, i_13_363, i_13_364, i_13_365, i_13_366, i_13_367, i_13_368, i_13_369, i_13_370, i_13_371, i_13_372, i_13_373, i_13_374, i_13_375, i_13_376, i_13_377, i_13_378, i_13_379, i_13_380, i_13_381, i_13_382, i_13_383, i_13_384, i_13_385, i_13_386, i_13_387, i_13_388, i_13_389, i_13_390, i_13_391, i_13_392, i_13_393, i_13_394, i_13_395, i_13_396, i_13_397, i_13_398, i_13_399, i_13_400, i_13_401, i_13_402, i_13_403, i_13_404, i_13_405, i_13_406, i_13_407, i_13_408, i_13_409, i_13_410, i_13_411, i_13_412, i_13_413, i_13_414, i_13_415, i_13_416, i_13_417, i_13_418, i_13_419, i_13_420, i_13_421, i_13_422, i_13_423, i_13_424, i_13_425, i_13_426, i_13_427, i_13_428, i_13_429, i_13_430, i_13_431, i_13_432, i_13_433, i_13_434, i_13_435, i_13_436, i_13_437, i_13_438, i_13_439, i_13_440, i_13_441, i_13_442, i_13_443, i_13_444, i_13_445, i_13_446, i_13_447, i_13_448, i_13_449, i_13_450, i_13_451, i_13_452, i_13_453, i_13_454, i_13_455, i_13_456, i_13_457, i_13_458, i_13_459, i_13_460, i_13_461, i_13_462, i_13_463, i_13_464, i_13_465, i_13_466, i_13_467, i_13_468, i_13_469, i_13_470, i_13_471, i_13_472, i_13_473, i_13_474, i_13_475, i_13_476, i_13_477, i_13_478, i_13_479, i_13_480, i_13_481, i_13_482, i_13_483, i_13_484, i_13_485, i_13_486, i_13_487, i_13_488, i_13_489, i_13_490, i_13_491, i_13_492, i_13_493, i_13_494, i_13_495, i_13_496, i_13_497, i_13_498, i_13_499, i_13_500, i_13_501, i_13_502, i_13_503, i_13_504, i_13_505, i_13_506, i_13_507, i_13_508, i_13_509, i_13_510, i_13_511, i_13_512, i_13_513, i_13_514, i_13_515, i_13_516, i_13_517, i_13_518, i_13_519, i_13_520, i_13_521, i_13_522, i_13_523, i_13_524, i_13_525, i_13_526, i_13_527, i_13_528, i_13_529, i_13_530, i_13_531, i_13_532, i_13_533, i_13_534, i_13_535, i_13_536, i_13_537, i_13_538, i_13_539, i_13_540, i_13_541, i_13_542, i_13_543, i_13_544, i_13_545, i_13_546, i_13_547, i_13_548, i_13_549, i_13_550, i_13_551, i_13_552, i_13_553, i_13_554, i_13_555, i_13_556, i_13_557, i_13_558, i_13_559, i_13_560, i_13_561, i_13_562, i_13_563, i_13_564, i_13_565, i_13_566, i_13_567, i_13_568, i_13_569, i_13_570, i_13_571, i_13_572, i_13_573, i_13_574, i_13_575, i_13_576, i_13_577, i_13_578, i_13_579, i_13_580, i_13_581, i_13_582, i_13_583, i_13_584, i_13_585, i_13_586, i_13_587, i_13_588, i_13_589, i_13_590, i_13_591, i_13_592, i_13_593, i_13_594, i_13_595, i_13_596, i_13_597, i_13_598, i_13_599, i_13_600, i_13_601, i_13_602, i_13_603, i_13_604, i_13_605, i_13_606, i_13_607, i_13_608, i_13_609, i_13_610, i_13_611, i_13_612, i_13_613, i_13_614, i_13_615, i_13_616, i_13_617, i_13_618, i_13_619, i_13_620, i_13_621, i_13_622, i_13_623, i_13_624, i_13_625, i_13_626, i_13_627, i_13_628, i_13_629, i_13_630, i_13_631, i_13_632, i_13_633, i_13_634, i_13_635, i_13_636, i_13_637, i_13_638, i_13_639, i_13_640, i_13_641, i_13_642, i_13_643, i_13_644, i_13_645, i_13_646, i_13_647, i_13_648, i_13_649, i_13_650, i_13_651, i_13_652, i_13_653, i_13_654, i_13_655, i_13_656, i_13_657, i_13_658, i_13_659, i_13_660, i_13_661, i_13_662, i_13_663, i_13_664, i_13_665, i_13_666, i_13_667, i_13_668, i_13_669, i_13_670, i_13_671, i_13_672, i_13_673, i_13_674, i_13_675, i_13_676, i_13_677, i_13_678, i_13_679, i_13_680, i_13_681, i_13_682, i_13_683, i_13_684, i_13_685, i_13_686, i_13_687, i_13_688, i_13_689, i_13_690, i_13_691, i_13_692, i_13_693, i_13_694, i_13_695, i_13_696, i_13_697, i_13_698, i_13_699, i_13_700, i_13_701, i_13_702, i_13_703, i_13_704, i_13_705, i_13_706, i_13_707, i_13_708, i_13_709, i_13_710, i_13_711, i_13_712, i_13_713, i_13_714, i_13_715, i_13_716, i_13_717, i_13_718, i_13_719, i_13_720, i_13_721, i_13_722, i_13_723, i_13_724, i_13_725, i_13_726, i_13_727, i_13_728, i_13_729, i_13_730, i_13_731, i_13_732, i_13_733, i_13_734, i_13_735, i_13_736, i_13_737, i_13_738, i_13_739, i_13_740, i_13_741, i_13_742, i_13_743, i_13_744, i_13_745, i_13_746, i_13_747, i_13_748, i_13_749, i_13_750, i_13_751, i_13_752, i_13_753, i_13_754, i_13_755, i_13_756, i_13_757, i_13_758, i_13_759, i_13_760, i_13_761, i_13_762, i_13_763, i_13_764, i_13_765, i_13_766, i_13_767, i_13_768, i_13_769, i_13_770, i_13_771, i_13_772, i_13_773, i_13_774, i_13_775, i_13_776, i_13_777, i_13_778, i_13_779, i_13_780, i_13_781, i_13_782, i_13_783, i_13_784, i_13_785, i_13_786, i_13_787, i_13_788, i_13_789, i_13_790, i_13_791, i_13_792, i_13_793, i_13_794, i_13_795, i_13_796, i_13_797, i_13_798, i_13_799, i_13_800, i_13_801, i_13_802, i_13_803, i_13_804, i_13_805, i_13_806, i_13_807, i_13_808, i_13_809, i_13_810, i_13_811, i_13_812, i_13_813, i_13_814, i_13_815, i_13_816, i_13_817, i_13_818, i_13_819, i_13_820, i_13_821, i_13_822, i_13_823, i_13_824, i_13_825, i_13_826, i_13_827, i_13_828, i_13_829, i_13_830, i_13_831, i_13_832, i_13_833, i_13_834, i_13_835, i_13_836, i_13_837, i_13_838, i_13_839, i_13_840, i_13_841, i_13_842, i_13_843, i_13_844, i_13_845, i_13_846, i_13_847, i_13_848, i_13_849, i_13_850, i_13_851, i_13_852, i_13_853, i_13_854, i_13_855, i_13_856, i_13_857, i_13_858, i_13_859, i_13_860, i_13_861, i_13_862, i_13_863, i_13_864, i_13_865, i_13_866, i_13_867, i_13_868, i_13_869, i_13_870, i_13_871, i_13_872, i_13_873, i_13_874, i_13_875, i_13_876, i_13_877, i_13_878, i_13_879, i_13_880, i_13_881, i_13_882, i_13_883, i_13_884, i_13_885, i_13_886, i_13_887, i_13_888, i_13_889, i_13_890, i_13_891, i_13_892, i_13_893, i_13_894, i_13_895, i_13_896, i_13_897, i_13_898, i_13_899, i_13_900, i_13_901, i_13_902, i_13_903, i_13_904, i_13_905, i_13_906, i_13_907, i_13_908, i_13_909, i_13_910, i_13_911, i_13_912, i_13_913, i_13_914, i_13_915, i_13_916, i_13_917, i_13_918, i_13_919, i_13_920, i_13_921, i_13_922, i_13_923, i_13_924, i_13_925, i_13_926, i_13_927, i_13_928, i_13_929, i_13_930, i_13_931, i_13_932, i_13_933, i_13_934, i_13_935, i_13_936, i_13_937, i_13_938, i_13_939, i_13_940, i_13_941, i_13_942, i_13_943, i_13_944, i_13_945, i_13_946, i_13_947, i_13_948, i_13_949, i_13_950, i_13_951, i_13_952, i_13_953, i_13_954, i_13_955, i_13_956, i_13_957, i_13_958, i_13_959, i_13_960, i_13_961, i_13_962, i_13_963, i_13_964, i_13_965, i_13_966, i_13_967, i_13_968, i_13_969, i_13_970, i_13_971, i_13_972, i_13_973, i_13_974, i_13_975, i_13_976, i_13_977, i_13_978, i_13_979, i_13_980, i_13_981, i_13_982, i_13_983, i_13_984, i_13_985, i_13_986, i_13_987, i_13_988, i_13_989, i_13_990, i_13_991, i_13_992, i_13_993, i_13_994, i_13_995, i_13_996, i_13_997, i_13_998, i_13_999, i_13_1000, i_13_1001, i_13_1002, i_13_1003, i_13_1004, i_13_1005, i_13_1006, i_13_1007, i_13_1008, i_13_1009, i_13_1010, i_13_1011, i_13_1012, i_13_1013, i_13_1014, i_13_1015, i_13_1016, i_13_1017, i_13_1018, i_13_1019, i_13_1020, i_13_1021, i_13_1022, i_13_1023, i_13_1024, i_13_1025, i_13_1026, i_13_1027, i_13_1028, i_13_1029, i_13_1030, i_13_1031, i_13_1032, i_13_1033, i_13_1034, i_13_1035, i_13_1036, i_13_1037, i_13_1038, i_13_1039, i_13_1040, i_13_1041, i_13_1042, i_13_1043, i_13_1044, i_13_1045, i_13_1046, i_13_1047, i_13_1048, i_13_1049, i_13_1050, i_13_1051, i_13_1052, i_13_1053, i_13_1054, i_13_1055, i_13_1056, i_13_1057, i_13_1058, i_13_1059, i_13_1060, i_13_1061, i_13_1062, i_13_1063, i_13_1064, i_13_1065, i_13_1066, i_13_1067, i_13_1068, i_13_1069, i_13_1070, i_13_1071, i_13_1072, i_13_1073, i_13_1074, i_13_1075, i_13_1076, i_13_1077, i_13_1078, i_13_1079, i_13_1080, i_13_1081, i_13_1082, i_13_1083, i_13_1084, i_13_1085, i_13_1086, i_13_1087, i_13_1088, i_13_1089, i_13_1090, i_13_1091, i_13_1092, i_13_1093, i_13_1094, i_13_1095, i_13_1096, i_13_1097, i_13_1098, i_13_1099, i_13_1100, i_13_1101, i_13_1102, i_13_1103, i_13_1104, i_13_1105, i_13_1106, i_13_1107, i_13_1108, i_13_1109, i_13_1110, i_13_1111, i_13_1112, i_13_1113, i_13_1114, i_13_1115, i_13_1116, i_13_1117, i_13_1118, i_13_1119, i_13_1120, i_13_1121, i_13_1122, i_13_1123, i_13_1124, i_13_1125, i_13_1126, i_13_1127, i_13_1128, i_13_1129, i_13_1130, i_13_1131, i_13_1132, i_13_1133, i_13_1134, i_13_1135, i_13_1136, i_13_1137, i_13_1138, i_13_1139, i_13_1140, i_13_1141, i_13_1142, i_13_1143, i_13_1144, i_13_1145, i_13_1146, i_13_1147, i_13_1148, i_13_1149, i_13_1150, i_13_1151, i_13_1152, i_13_1153, i_13_1154, i_13_1155, i_13_1156, i_13_1157, i_13_1158, i_13_1159, i_13_1160, i_13_1161, i_13_1162, i_13_1163, i_13_1164, i_13_1165, i_13_1166, i_13_1167, i_13_1168, i_13_1169, i_13_1170, i_13_1171, i_13_1172, i_13_1173, i_13_1174, i_13_1175, i_13_1176, i_13_1177, i_13_1178, i_13_1179, i_13_1180, i_13_1181, i_13_1182, i_13_1183, i_13_1184, i_13_1185, i_13_1186, i_13_1187, i_13_1188, i_13_1189, i_13_1190, i_13_1191, i_13_1192, i_13_1193, i_13_1194, i_13_1195, i_13_1196, i_13_1197, i_13_1198, i_13_1199, i_13_1200, i_13_1201, i_13_1202, i_13_1203, i_13_1204, i_13_1205, i_13_1206, i_13_1207, i_13_1208, i_13_1209, i_13_1210, i_13_1211, i_13_1212, i_13_1213, i_13_1214, i_13_1215, i_13_1216, i_13_1217, i_13_1218, i_13_1219, i_13_1220, i_13_1221, i_13_1222, i_13_1223, i_13_1224, i_13_1225, i_13_1226, i_13_1227, i_13_1228, i_13_1229, i_13_1230, i_13_1231, i_13_1232, i_13_1233, i_13_1234, i_13_1235, i_13_1236, i_13_1237, i_13_1238, i_13_1239, i_13_1240, i_13_1241, i_13_1242, i_13_1243, i_13_1244, i_13_1245, i_13_1246, i_13_1247, i_13_1248, i_13_1249, i_13_1250, i_13_1251, i_13_1252, i_13_1253, i_13_1254, i_13_1255, i_13_1256, i_13_1257, i_13_1258, i_13_1259, i_13_1260, i_13_1261, i_13_1262, i_13_1263, i_13_1264, i_13_1265, i_13_1266, i_13_1267, i_13_1268, i_13_1269, i_13_1270, i_13_1271, i_13_1272, i_13_1273, i_13_1274, i_13_1275, i_13_1276, i_13_1277, i_13_1278, i_13_1279, i_13_1280, i_13_1281, i_13_1282, i_13_1283, i_13_1284, i_13_1285, i_13_1286, i_13_1287, i_13_1288, i_13_1289, i_13_1290, i_13_1291, i_13_1292, i_13_1293, i_13_1294, i_13_1295, i_13_1296, i_13_1297, i_13_1298, i_13_1299, i_13_1300, i_13_1301, i_13_1302, i_13_1303, i_13_1304, i_13_1305, i_13_1306, i_13_1307, i_13_1308, i_13_1309, i_13_1310, i_13_1311, i_13_1312, i_13_1313, i_13_1314, i_13_1315, i_13_1316, i_13_1317, i_13_1318, i_13_1319, i_13_1320, i_13_1321, i_13_1322, i_13_1323, i_13_1324, i_13_1325, i_13_1326, i_13_1327, i_13_1328, i_13_1329, i_13_1330, i_13_1331, i_13_1332, i_13_1333, i_13_1334, i_13_1335, i_13_1336, i_13_1337, i_13_1338, i_13_1339, i_13_1340, i_13_1341, i_13_1342, i_13_1343, i_13_1344, i_13_1345, i_13_1346, i_13_1347, i_13_1348, i_13_1349, i_13_1350, i_13_1351, i_13_1352, i_13_1353, i_13_1354, i_13_1355, i_13_1356, i_13_1357, i_13_1358, i_13_1359, i_13_1360, i_13_1361, i_13_1362, i_13_1363, i_13_1364, i_13_1365, i_13_1366, i_13_1367, i_13_1368, i_13_1369, i_13_1370, i_13_1371, i_13_1372, i_13_1373, i_13_1374, i_13_1375, i_13_1376, i_13_1377, i_13_1378, i_13_1379, i_13_1380, i_13_1381, i_13_1382, i_13_1383, i_13_1384, i_13_1385, i_13_1386, i_13_1387, i_13_1388, i_13_1389, i_13_1390, i_13_1391, i_13_1392, i_13_1393, i_13_1394, i_13_1395, i_13_1396, i_13_1397, i_13_1398, i_13_1399, i_13_1400, i_13_1401, i_13_1402, i_13_1403, i_13_1404, i_13_1405, i_13_1406, i_13_1407, i_13_1408, i_13_1409, i_13_1410, i_13_1411, i_13_1412, i_13_1413, i_13_1414, i_13_1415, i_13_1416, i_13_1417, i_13_1418, i_13_1419, i_13_1420, i_13_1421, i_13_1422, i_13_1423, i_13_1424, i_13_1425, i_13_1426, i_13_1427, i_13_1428, i_13_1429, i_13_1430, i_13_1431, i_13_1432, i_13_1433, i_13_1434, i_13_1435, i_13_1436, i_13_1437, i_13_1438, i_13_1439, i_13_1440, i_13_1441, i_13_1442, i_13_1443, i_13_1444, i_13_1445, i_13_1446, i_13_1447, i_13_1448, i_13_1449, i_13_1450, i_13_1451, i_13_1452, i_13_1453, i_13_1454, i_13_1455, i_13_1456, i_13_1457, i_13_1458, i_13_1459, i_13_1460, i_13_1461, i_13_1462, i_13_1463, i_13_1464, i_13_1465, i_13_1466, i_13_1467, i_13_1468, i_13_1469, i_13_1470, i_13_1471, i_13_1472, i_13_1473, i_13_1474, i_13_1475, i_13_1476, i_13_1477, i_13_1478, i_13_1479, i_13_1480, i_13_1481, i_13_1482, i_13_1483, i_13_1484, i_13_1485, i_13_1486, i_13_1487, i_13_1488, i_13_1489, i_13_1490, i_13_1491, i_13_1492, i_13_1493, i_13_1494, i_13_1495, i_13_1496, i_13_1497, i_13_1498, i_13_1499, i_13_1500, i_13_1501, i_13_1502, i_13_1503, i_13_1504, i_13_1505, i_13_1506, i_13_1507, i_13_1508, i_13_1509, i_13_1510, i_13_1511, i_13_1512, i_13_1513, i_13_1514, i_13_1515, i_13_1516, i_13_1517, i_13_1518, i_13_1519, i_13_1520, i_13_1521, i_13_1522, i_13_1523, i_13_1524, i_13_1525, i_13_1526, i_13_1527, i_13_1528, i_13_1529, i_13_1530, i_13_1531, i_13_1532, i_13_1533, i_13_1534, i_13_1535, i_13_1536, i_13_1537, i_13_1538, i_13_1539, i_13_1540, i_13_1541, i_13_1542, i_13_1543, i_13_1544, i_13_1545, i_13_1546, i_13_1547, i_13_1548, i_13_1549, i_13_1550, i_13_1551, i_13_1552, i_13_1553, i_13_1554, i_13_1555, i_13_1556, i_13_1557, i_13_1558, i_13_1559, i_13_1560, i_13_1561, i_13_1562, i_13_1563, i_13_1564, i_13_1565, i_13_1566, i_13_1567, i_13_1568, i_13_1569, i_13_1570, i_13_1571, i_13_1572, i_13_1573, i_13_1574, i_13_1575, i_13_1576, i_13_1577, i_13_1578, i_13_1579, i_13_1580, i_13_1581, i_13_1582, i_13_1583, i_13_1584, i_13_1585, i_13_1586, i_13_1587, i_13_1588, i_13_1589, i_13_1590, i_13_1591, i_13_1592, i_13_1593, i_13_1594, i_13_1595, i_13_1596, i_13_1597, i_13_1598, i_13_1599, i_13_1600, i_13_1601, i_13_1602, i_13_1603, i_13_1604, i_13_1605, i_13_1606, i_13_1607, i_13_1608, i_13_1609, i_13_1610, i_13_1611, i_13_1612, i_13_1613, i_13_1614, i_13_1615, i_13_1616, i_13_1617, i_13_1618, i_13_1619, i_13_1620, i_13_1621, i_13_1622, i_13_1623, i_13_1624, i_13_1625, i_13_1626, i_13_1627, i_13_1628, i_13_1629, i_13_1630, i_13_1631, i_13_1632, i_13_1633, i_13_1634, i_13_1635, i_13_1636, i_13_1637, i_13_1638, i_13_1639, i_13_1640, i_13_1641, i_13_1642, i_13_1643, i_13_1644, i_13_1645, i_13_1646, i_13_1647, i_13_1648, i_13_1649, i_13_1650, i_13_1651, i_13_1652, i_13_1653, i_13_1654, i_13_1655, i_13_1656, i_13_1657, i_13_1658, i_13_1659, i_13_1660, i_13_1661, i_13_1662, i_13_1663, i_13_1664, i_13_1665, i_13_1666, i_13_1667, i_13_1668, i_13_1669, i_13_1670, i_13_1671, i_13_1672, i_13_1673, i_13_1674, i_13_1675, i_13_1676, i_13_1677, i_13_1678, i_13_1679, i_13_1680, i_13_1681, i_13_1682, i_13_1683, i_13_1684, i_13_1685, i_13_1686, i_13_1687, i_13_1688, i_13_1689, i_13_1690, i_13_1691, i_13_1692, i_13_1693, i_13_1694, i_13_1695, i_13_1696, i_13_1697, i_13_1698, i_13_1699, i_13_1700, i_13_1701, i_13_1702, i_13_1703, i_13_1704, i_13_1705, i_13_1706, i_13_1707, i_13_1708, i_13_1709, i_13_1710, i_13_1711, i_13_1712, i_13_1713, i_13_1714, i_13_1715, i_13_1716, i_13_1717, i_13_1718, i_13_1719, i_13_1720, i_13_1721, i_13_1722, i_13_1723, i_13_1724, i_13_1725, i_13_1726, i_13_1727, i_13_1728, i_13_1729, i_13_1730, i_13_1731, i_13_1732, i_13_1733, i_13_1734, i_13_1735, i_13_1736, i_13_1737, i_13_1738, i_13_1739, i_13_1740, i_13_1741, i_13_1742, i_13_1743, i_13_1744, i_13_1745, i_13_1746, i_13_1747, i_13_1748, i_13_1749, i_13_1750, i_13_1751, i_13_1752, i_13_1753, i_13_1754, i_13_1755, i_13_1756, i_13_1757, i_13_1758, i_13_1759, i_13_1760, i_13_1761, i_13_1762, i_13_1763, i_13_1764, i_13_1765, i_13_1766, i_13_1767, i_13_1768, i_13_1769, i_13_1770, i_13_1771, i_13_1772, i_13_1773, i_13_1774, i_13_1775, i_13_1776, i_13_1777, i_13_1778, i_13_1779, i_13_1780, i_13_1781, i_13_1782, i_13_1783, i_13_1784, i_13_1785, i_13_1786, i_13_1787, i_13_1788, i_13_1789, i_13_1790, i_13_1791, i_13_1792, i_13_1793, i_13_1794, i_13_1795, i_13_1796, i_13_1797, i_13_1798, i_13_1799, i_13_1800, i_13_1801, i_13_1802, i_13_1803, i_13_1804, i_13_1805, i_13_1806, i_13_1807, i_13_1808, i_13_1809, i_13_1810, i_13_1811, i_13_1812, i_13_1813, i_13_1814, i_13_1815, i_13_1816, i_13_1817, i_13_1818, i_13_1819, i_13_1820, i_13_1821, i_13_1822, i_13_1823, i_13_1824, i_13_1825, i_13_1826, i_13_1827, i_13_1828, i_13_1829, i_13_1830, i_13_1831, i_13_1832, i_13_1833, i_13_1834, i_13_1835, i_13_1836, i_13_1837, i_13_1838, i_13_1839, i_13_1840, i_13_1841, i_13_1842, i_13_1843, i_13_1844, i_13_1845, i_13_1846, i_13_1847, i_13_1848, i_13_1849, i_13_1850, i_13_1851, i_13_1852, i_13_1853, i_13_1854, i_13_1855, i_13_1856, i_13_1857, i_13_1858, i_13_1859, i_13_1860, i_13_1861, i_13_1862, i_13_1863, i_13_1864, i_13_1865, i_13_1866, i_13_1867, i_13_1868, i_13_1869, i_13_1870, i_13_1871, i_13_1872, i_13_1873, i_13_1874, i_13_1875, i_13_1876, i_13_1877, i_13_1878, i_13_1879, i_13_1880, i_13_1881, i_13_1882, i_13_1883, i_13_1884, i_13_1885, i_13_1886, i_13_1887, i_13_1888, i_13_1889, i_13_1890, i_13_1891, i_13_1892, i_13_1893, i_13_1894, i_13_1895, i_13_1896, i_13_1897, i_13_1898, i_13_1899, i_13_1900, i_13_1901, i_13_1902, i_13_1903, i_13_1904, i_13_1905, i_13_1906, i_13_1907, i_13_1908, i_13_1909, i_13_1910, i_13_1911, i_13_1912, i_13_1913, i_13_1914, i_13_1915, i_13_1916, i_13_1917, i_13_1918, i_13_1919, i_13_1920, i_13_1921, i_13_1922, i_13_1923, i_13_1924, i_13_1925, i_13_1926, i_13_1927, i_13_1928, i_13_1929, i_13_1930, i_13_1931, i_13_1932, i_13_1933, i_13_1934, i_13_1935, i_13_1936, i_13_1937, i_13_1938, i_13_1939, i_13_1940, i_13_1941, i_13_1942, i_13_1943, i_13_1944, i_13_1945, i_13_1946, i_13_1947, i_13_1948, i_13_1949, i_13_1950, i_13_1951, i_13_1952, i_13_1953, i_13_1954, i_13_1955, i_13_1956, i_13_1957, i_13_1958, i_13_1959, i_13_1960, i_13_1961, i_13_1962, i_13_1963, i_13_1964, i_13_1965, i_13_1966, i_13_1967, i_13_1968, i_13_1969, i_13_1970, i_13_1971, i_13_1972, i_13_1973, i_13_1974, i_13_1975, i_13_1976, i_13_1977, i_13_1978, i_13_1979, i_13_1980, i_13_1981, i_13_1982, i_13_1983, i_13_1984, i_13_1985, i_13_1986, i_13_1987, i_13_1988, i_13_1989, i_13_1990, i_13_1991, i_13_1992, i_13_1993, i_13_1994, i_13_1995, i_13_1996, i_13_1997, i_13_1998, i_13_1999, i_13_2000, i_13_2001, i_13_2002, i_13_2003, i_13_2004, i_13_2005, i_13_2006, i_13_2007, i_13_2008, i_13_2009, i_13_2010, i_13_2011, i_13_2012, i_13_2013, i_13_2014, i_13_2015, i_13_2016, i_13_2017, i_13_2018, i_13_2019, i_13_2020, i_13_2021, i_13_2022, i_13_2023, i_13_2024, i_13_2025, i_13_2026, i_13_2027, i_13_2028, i_13_2029, i_13_2030, i_13_2031, i_13_2032, i_13_2033, i_13_2034, i_13_2035, i_13_2036, i_13_2037, i_13_2038, i_13_2039, i_13_2040, i_13_2041, i_13_2042, i_13_2043, i_13_2044, i_13_2045, i_13_2046, i_13_2047, i_13_2048, i_13_2049, i_13_2050, i_13_2051, i_13_2052, i_13_2053, i_13_2054, i_13_2055, i_13_2056, i_13_2057, i_13_2058, i_13_2059, i_13_2060, i_13_2061, i_13_2062, i_13_2063, i_13_2064, i_13_2065, i_13_2066, i_13_2067, i_13_2068, i_13_2069, i_13_2070, i_13_2071, i_13_2072, i_13_2073, i_13_2074, i_13_2075, i_13_2076, i_13_2077, i_13_2078, i_13_2079, i_13_2080, i_13_2081, i_13_2082, i_13_2083, i_13_2084, i_13_2085, i_13_2086, i_13_2087, i_13_2088, i_13_2089, i_13_2090, i_13_2091, i_13_2092, i_13_2093, i_13_2094, i_13_2095, i_13_2096, i_13_2097, i_13_2098, i_13_2099, i_13_2100, i_13_2101, i_13_2102, i_13_2103, i_13_2104, i_13_2105, i_13_2106, i_13_2107, i_13_2108, i_13_2109, i_13_2110, i_13_2111, i_13_2112, i_13_2113, i_13_2114, i_13_2115, i_13_2116, i_13_2117, i_13_2118, i_13_2119, i_13_2120, i_13_2121, i_13_2122, i_13_2123, i_13_2124, i_13_2125, i_13_2126, i_13_2127, i_13_2128, i_13_2129, i_13_2130, i_13_2131, i_13_2132, i_13_2133, i_13_2134, i_13_2135, i_13_2136, i_13_2137, i_13_2138, i_13_2139, i_13_2140, i_13_2141, i_13_2142, i_13_2143, i_13_2144, i_13_2145, i_13_2146, i_13_2147, i_13_2148, i_13_2149, i_13_2150, i_13_2151, i_13_2152, i_13_2153, i_13_2154, i_13_2155, i_13_2156, i_13_2157, i_13_2158, i_13_2159, i_13_2160, i_13_2161, i_13_2162, i_13_2163, i_13_2164, i_13_2165, i_13_2166, i_13_2167, i_13_2168, i_13_2169, i_13_2170, i_13_2171, i_13_2172, i_13_2173, i_13_2174, i_13_2175, i_13_2176, i_13_2177, i_13_2178, i_13_2179, i_13_2180, i_13_2181, i_13_2182, i_13_2183, i_13_2184, i_13_2185, i_13_2186, i_13_2187, i_13_2188, i_13_2189, i_13_2190, i_13_2191, i_13_2192, i_13_2193, i_13_2194, i_13_2195, i_13_2196, i_13_2197, i_13_2198, i_13_2199, i_13_2200, i_13_2201, i_13_2202, i_13_2203, i_13_2204, i_13_2205, i_13_2206, i_13_2207, i_13_2208, i_13_2209, i_13_2210, i_13_2211, i_13_2212, i_13_2213, i_13_2214, i_13_2215, i_13_2216, i_13_2217, i_13_2218, i_13_2219, i_13_2220, i_13_2221, i_13_2222, i_13_2223, i_13_2224, i_13_2225, i_13_2226, i_13_2227, i_13_2228, i_13_2229, i_13_2230, i_13_2231, i_13_2232, i_13_2233, i_13_2234, i_13_2235, i_13_2236, i_13_2237, i_13_2238, i_13_2239, i_13_2240, i_13_2241, i_13_2242, i_13_2243, i_13_2244, i_13_2245, i_13_2246, i_13_2247, i_13_2248, i_13_2249, i_13_2250, i_13_2251, i_13_2252, i_13_2253, i_13_2254, i_13_2255, i_13_2256, i_13_2257, i_13_2258, i_13_2259, i_13_2260, i_13_2261, i_13_2262, i_13_2263, i_13_2264, i_13_2265, i_13_2266, i_13_2267, i_13_2268, i_13_2269, i_13_2270, i_13_2271, i_13_2272, i_13_2273, i_13_2274, i_13_2275, i_13_2276, i_13_2277, i_13_2278, i_13_2279, i_13_2280, i_13_2281, i_13_2282, i_13_2283, i_13_2284, i_13_2285, i_13_2286, i_13_2287, i_13_2288, i_13_2289, i_13_2290, i_13_2291, i_13_2292, i_13_2293, i_13_2294, i_13_2295, i_13_2296, i_13_2297, i_13_2298, i_13_2299, i_13_2300, i_13_2301, i_13_2302, i_13_2303, i_13_2304, i_13_2305, i_13_2306, i_13_2307, i_13_2308, i_13_2309, i_13_2310, i_13_2311, i_13_2312, i_13_2313, i_13_2314, i_13_2315, i_13_2316, i_13_2317, i_13_2318, i_13_2319, i_13_2320, i_13_2321, i_13_2322, i_13_2323, i_13_2324, i_13_2325, i_13_2326, i_13_2327, i_13_2328, i_13_2329, i_13_2330, i_13_2331, i_13_2332, i_13_2333, i_13_2334, i_13_2335, i_13_2336, i_13_2337, i_13_2338, i_13_2339, i_13_2340, i_13_2341, i_13_2342, i_13_2343, i_13_2344, i_13_2345, i_13_2346, i_13_2347, i_13_2348, i_13_2349, i_13_2350, i_13_2351, i_13_2352, i_13_2353, i_13_2354, i_13_2355, i_13_2356, i_13_2357, i_13_2358, i_13_2359, i_13_2360, i_13_2361, i_13_2362, i_13_2363, i_13_2364, i_13_2365, i_13_2366, i_13_2367, i_13_2368, i_13_2369, i_13_2370, i_13_2371, i_13_2372, i_13_2373, i_13_2374, i_13_2375, i_13_2376, i_13_2377, i_13_2378, i_13_2379, i_13_2380, i_13_2381, i_13_2382, i_13_2383, i_13_2384, i_13_2385, i_13_2386, i_13_2387, i_13_2388, i_13_2389, i_13_2390, i_13_2391, i_13_2392, i_13_2393, i_13_2394, i_13_2395, i_13_2396, i_13_2397, i_13_2398, i_13_2399, i_13_2400, i_13_2401, i_13_2402, i_13_2403, i_13_2404, i_13_2405, i_13_2406, i_13_2407, i_13_2408, i_13_2409, i_13_2410, i_13_2411, i_13_2412, i_13_2413, i_13_2414, i_13_2415, i_13_2416, i_13_2417, i_13_2418, i_13_2419, i_13_2420, i_13_2421, i_13_2422, i_13_2423, i_13_2424, i_13_2425, i_13_2426, i_13_2427, i_13_2428, i_13_2429, i_13_2430, i_13_2431, i_13_2432, i_13_2433, i_13_2434, i_13_2435, i_13_2436, i_13_2437, i_13_2438, i_13_2439, i_13_2440, i_13_2441, i_13_2442, i_13_2443, i_13_2444, i_13_2445, i_13_2446, i_13_2447, i_13_2448, i_13_2449, i_13_2450, i_13_2451, i_13_2452, i_13_2453, i_13_2454, i_13_2455, i_13_2456, i_13_2457, i_13_2458, i_13_2459, i_13_2460, i_13_2461, i_13_2462, i_13_2463, i_13_2464, i_13_2465, i_13_2466, i_13_2467, i_13_2468, i_13_2469, i_13_2470, i_13_2471, i_13_2472, i_13_2473, i_13_2474, i_13_2475, i_13_2476, i_13_2477, i_13_2478, i_13_2479, i_13_2480, i_13_2481, i_13_2482, i_13_2483, i_13_2484, i_13_2485, i_13_2486, i_13_2487, i_13_2488, i_13_2489, i_13_2490, i_13_2491, i_13_2492, i_13_2493, i_13_2494, i_13_2495, i_13_2496, i_13_2497, i_13_2498, i_13_2499, i_13_2500, i_13_2501, i_13_2502, i_13_2503, i_13_2504, i_13_2505, i_13_2506, i_13_2507, i_13_2508, i_13_2509, i_13_2510, i_13_2511, i_13_2512, i_13_2513, i_13_2514, i_13_2515, i_13_2516, i_13_2517, i_13_2518, i_13_2519, i_13_2520, i_13_2521, i_13_2522, i_13_2523, i_13_2524, i_13_2525, i_13_2526, i_13_2527, i_13_2528, i_13_2529, i_13_2530, i_13_2531, i_13_2532, i_13_2533, i_13_2534, i_13_2535, i_13_2536, i_13_2537, i_13_2538, i_13_2539, i_13_2540, i_13_2541, i_13_2542, i_13_2543, i_13_2544, i_13_2545, i_13_2546, i_13_2547, i_13_2548, i_13_2549, i_13_2550, i_13_2551, i_13_2552, i_13_2553, i_13_2554, i_13_2555, i_13_2556, i_13_2557, i_13_2558, i_13_2559, i_13_2560, i_13_2561, i_13_2562, i_13_2563, i_13_2564, i_13_2565, i_13_2566, i_13_2567, i_13_2568, i_13_2569, i_13_2570, i_13_2571, i_13_2572, i_13_2573, i_13_2574, i_13_2575, i_13_2576, i_13_2577, i_13_2578, i_13_2579, i_13_2580, i_13_2581, i_13_2582, i_13_2583, i_13_2584, i_13_2585, i_13_2586, i_13_2587, i_13_2588, i_13_2589, i_13_2590, i_13_2591, i_13_2592, i_13_2593, i_13_2594, i_13_2595, i_13_2596, i_13_2597, i_13_2598, i_13_2599, i_13_2600, i_13_2601, i_13_2602, i_13_2603, i_13_2604, i_13_2605, i_13_2606, i_13_2607, i_13_2608, i_13_2609, i_13_2610, i_13_2611, i_13_2612, i_13_2613, i_13_2614, i_13_2615, i_13_2616, i_13_2617, i_13_2618, i_13_2619, i_13_2620, i_13_2621, i_13_2622, i_13_2623, i_13_2624, i_13_2625, i_13_2626, i_13_2627, i_13_2628, i_13_2629, i_13_2630, i_13_2631, i_13_2632, i_13_2633, i_13_2634, i_13_2635, i_13_2636, i_13_2637, i_13_2638, i_13_2639, i_13_2640, i_13_2641, i_13_2642, i_13_2643, i_13_2644, i_13_2645, i_13_2646, i_13_2647, i_13_2648, i_13_2649, i_13_2650, i_13_2651, i_13_2652, i_13_2653, i_13_2654, i_13_2655, i_13_2656, i_13_2657, i_13_2658, i_13_2659, i_13_2660, i_13_2661, i_13_2662, i_13_2663, i_13_2664, i_13_2665, i_13_2666, i_13_2667, i_13_2668, i_13_2669, i_13_2670, i_13_2671, i_13_2672, i_13_2673, i_13_2674, i_13_2675, i_13_2676, i_13_2677, i_13_2678, i_13_2679, i_13_2680, i_13_2681, i_13_2682, i_13_2683, i_13_2684, i_13_2685, i_13_2686, i_13_2687, i_13_2688, i_13_2689, i_13_2690, i_13_2691, i_13_2692, i_13_2693, i_13_2694, i_13_2695, i_13_2696, i_13_2697, i_13_2698, i_13_2699, i_13_2700, i_13_2701, i_13_2702, i_13_2703, i_13_2704, i_13_2705, i_13_2706, i_13_2707, i_13_2708, i_13_2709, i_13_2710, i_13_2711, i_13_2712, i_13_2713, i_13_2714, i_13_2715, i_13_2716, i_13_2717, i_13_2718, i_13_2719, i_13_2720, i_13_2721, i_13_2722, i_13_2723, i_13_2724, i_13_2725, i_13_2726, i_13_2727, i_13_2728, i_13_2729, i_13_2730, i_13_2731, i_13_2732, i_13_2733, i_13_2734, i_13_2735, i_13_2736, i_13_2737, i_13_2738, i_13_2739, i_13_2740, i_13_2741, i_13_2742, i_13_2743, i_13_2744, i_13_2745, i_13_2746, i_13_2747, i_13_2748, i_13_2749, i_13_2750, i_13_2751, i_13_2752, i_13_2753, i_13_2754, i_13_2755, i_13_2756, i_13_2757, i_13_2758, i_13_2759, i_13_2760, i_13_2761, i_13_2762, i_13_2763, i_13_2764, i_13_2765, i_13_2766, i_13_2767, i_13_2768, i_13_2769, i_13_2770, i_13_2771, i_13_2772, i_13_2773, i_13_2774, i_13_2775, i_13_2776, i_13_2777, i_13_2778, i_13_2779, i_13_2780, i_13_2781, i_13_2782, i_13_2783, i_13_2784, i_13_2785, i_13_2786, i_13_2787, i_13_2788, i_13_2789, i_13_2790, i_13_2791, i_13_2792, i_13_2793, i_13_2794, i_13_2795, i_13_2796, i_13_2797, i_13_2798, i_13_2799, i_13_2800, i_13_2801, i_13_2802, i_13_2803, i_13_2804, i_13_2805, i_13_2806, i_13_2807, i_13_2808, i_13_2809, i_13_2810, i_13_2811, i_13_2812, i_13_2813, i_13_2814, i_13_2815, i_13_2816, i_13_2817, i_13_2818, i_13_2819, i_13_2820, i_13_2821, i_13_2822, i_13_2823, i_13_2824, i_13_2825, i_13_2826, i_13_2827, i_13_2828, i_13_2829, i_13_2830, i_13_2831, i_13_2832, i_13_2833, i_13_2834, i_13_2835, i_13_2836, i_13_2837, i_13_2838, i_13_2839, i_13_2840, i_13_2841, i_13_2842, i_13_2843, i_13_2844, i_13_2845, i_13_2846, i_13_2847, i_13_2848, i_13_2849, i_13_2850, i_13_2851, i_13_2852, i_13_2853, i_13_2854, i_13_2855, i_13_2856, i_13_2857, i_13_2858, i_13_2859, i_13_2860, i_13_2861, i_13_2862, i_13_2863, i_13_2864, i_13_2865, i_13_2866, i_13_2867, i_13_2868, i_13_2869, i_13_2870, i_13_2871, i_13_2872, i_13_2873, i_13_2874, i_13_2875, i_13_2876, i_13_2877, i_13_2878, i_13_2879, i_13_2880, i_13_2881, i_13_2882, i_13_2883, i_13_2884, i_13_2885, i_13_2886, i_13_2887, i_13_2888, i_13_2889, i_13_2890, i_13_2891, i_13_2892, i_13_2893, i_13_2894, i_13_2895, i_13_2896, i_13_2897, i_13_2898, i_13_2899, i_13_2900, i_13_2901, i_13_2902, i_13_2903, i_13_2904, i_13_2905, i_13_2906, i_13_2907, i_13_2908, i_13_2909, i_13_2910, i_13_2911, i_13_2912, i_13_2913, i_13_2914, i_13_2915, i_13_2916, i_13_2917, i_13_2918, i_13_2919, i_13_2920, i_13_2921, i_13_2922, i_13_2923, i_13_2924, i_13_2925, i_13_2926, i_13_2927, i_13_2928, i_13_2929, i_13_2930, i_13_2931, i_13_2932, i_13_2933, i_13_2934, i_13_2935, i_13_2936, i_13_2937, i_13_2938, i_13_2939, i_13_2940, i_13_2941, i_13_2942, i_13_2943, i_13_2944, i_13_2945, i_13_2946, i_13_2947, i_13_2948, i_13_2949, i_13_2950, i_13_2951, i_13_2952, i_13_2953, i_13_2954, i_13_2955, i_13_2956, i_13_2957, i_13_2958, i_13_2959, i_13_2960, i_13_2961, i_13_2962, i_13_2963, i_13_2964, i_13_2965, i_13_2966, i_13_2967, i_13_2968, i_13_2969, i_13_2970, i_13_2971, i_13_2972, i_13_2973, i_13_2974, i_13_2975, i_13_2976, i_13_2977, i_13_2978, i_13_2979, i_13_2980, i_13_2981, i_13_2982, i_13_2983, i_13_2984, i_13_2985, i_13_2986, i_13_2987, i_13_2988, i_13_2989, i_13_2990, i_13_2991, i_13_2992, i_13_2993, i_13_2994, i_13_2995, i_13_2996, i_13_2997, i_13_2998, i_13_2999, i_13_3000, i_13_3001, i_13_3002, i_13_3003, i_13_3004, i_13_3005, i_13_3006, i_13_3007, i_13_3008, i_13_3009, i_13_3010, i_13_3011, i_13_3012, i_13_3013, i_13_3014, i_13_3015, i_13_3016, i_13_3017, i_13_3018, i_13_3019, i_13_3020, i_13_3021, i_13_3022, i_13_3023, i_13_3024, i_13_3025, i_13_3026, i_13_3027, i_13_3028, i_13_3029, i_13_3030, i_13_3031, i_13_3032, i_13_3033, i_13_3034, i_13_3035, i_13_3036, i_13_3037, i_13_3038, i_13_3039, i_13_3040, i_13_3041, i_13_3042, i_13_3043, i_13_3044, i_13_3045, i_13_3046, i_13_3047, i_13_3048, i_13_3049, i_13_3050, i_13_3051, i_13_3052, i_13_3053, i_13_3054, i_13_3055, i_13_3056, i_13_3057, i_13_3058, i_13_3059, i_13_3060, i_13_3061, i_13_3062, i_13_3063, i_13_3064, i_13_3065, i_13_3066, i_13_3067, i_13_3068, i_13_3069, i_13_3070, i_13_3071, i_13_3072, i_13_3073, i_13_3074, i_13_3075, i_13_3076, i_13_3077, i_13_3078, i_13_3079, i_13_3080, i_13_3081, i_13_3082, i_13_3083, i_13_3084, i_13_3085, i_13_3086, i_13_3087, i_13_3088, i_13_3089, i_13_3090, i_13_3091, i_13_3092, i_13_3093, i_13_3094, i_13_3095, i_13_3096, i_13_3097, i_13_3098, i_13_3099, i_13_3100, i_13_3101, i_13_3102, i_13_3103, i_13_3104, i_13_3105, i_13_3106, i_13_3107, i_13_3108, i_13_3109, i_13_3110, i_13_3111, i_13_3112, i_13_3113, i_13_3114, i_13_3115, i_13_3116, i_13_3117, i_13_3118, i_13_3119, i_13_3120, i_13_3121, i_13_3122, i_13_3123, i_13_3124, i_13_3125, i_13_3126, i_13_3127, i_13_3128, i_13_3129, i_13_3130, i_13_3131, i_13_3132, i_13_3133, i_13_3134, i_13_3135, i_13_3136, i_13_3137, i_13_3138, i_13_3139, i_13_3140, i_13_3141, i_13_3142, i_13_3143, i_13_3144, i_13_3145, i_13_3146, i_13_3147, i_13_3148, i_13_3149, i_13_3150, i_13_3151, i_13_3152, i_13_3153, i_13_3154, i_13_3155, i_13_3156, i_13_3157, i_13_3158, i_13_3159, i_13_3160, i_13_3161, i_13_3162, i_13_3163, i_13_3164, i_13_3165, i_13_3166, i_13_3167, i_13_3168, i_13_3169, i_13_3170, i_13_3171, i_13_3172, i_13_3173, i_13_3174, i_13_3175, i_13_3176, i_13_3177, i_13_3178, i_13_3179, i_13_3180, i_13_3181, i_13_3182, i_13_3183, i_13_3184, i_13_3185, i_13_3186, i_13_3187, i_13_3188, i_13_3189, i_13_3190, i_13_3191, i_13_3192, i_13_3193, i_13_3194, i_13_3195, i_13_3196, i_13_3197, i_13_3198, i_13_3199, i_13_3200, i_13_3201, i_13_3202, i_13_3203, i_13_3204, i_13_3205, i_13_3206, i_13_3207, i_13_3208, i_13_3209, i_13_3210, i_13_3211, i_13_3212, i_13_3213, i_13_3214, i_13_3215, i_13_3216, i_13_3217, i_13_3218, i_13_3219, i_13_3220, i_13_3221, i_13_3222, i_13_3223, i_13_3224, i_13_3225, i_13_3226, i_13_3227, i_13_3228, i_13_3229, i_13_3230, i_13_3231, i_13_3232, i_13_3233, i_13_3234, i_13_3235, i_13_3236, i_13_3237, i_13_3238, i_13_3239, i_13_3240, i_13_3241, i_13_3242, i_13_3243, i_13_3244, i_13_3245, i_13_3246, i_13_3247, i_13_3248, i_13_3249, i_13_3250, i_13_3251, i_13_3252, i_13_3253, i_13_3254, i_13_3255, i_13_3256, i_13_3257, i_13_3258, i_13_3259, i_13_3260, i_13_3261, i_13_3262, i_13_3263, i_13_3264, i_13_3265, i_13_3266, i_13_3267, i_13_3268, i_13_3269, i_13_3270, i_13_3271, i_13_3272, i_13_3273, i_13_3274, i_13_3275, i_13_3276, i_13_3277, i_13_3278, i_13_3279, i_13_3280, i_13_3281, i_13_3282, i_13_3283, i_13_3284, i_13_3285, i_13_3286, i_13_3287, i_13_3288, i_13_3289, i_13_3290, i_13_3291, i_13_3292, i_13_3293, i_13_3294, i_13_3295, i_13_3296, i_13_3297, i_13_3298, i_13_3299, i_13_3300, i_13_3301, i_13_3302, i_13_3303, i_13_3304, i_13_3305, i_13_3306, i_13_3307, i_13_3308, i_13_3309, i_13_3310, i_13_3311, i_13_3312, i_13_3313, i_13_3314, i_13_3315, i_13_3316, i_13_3317, i_13_3318, i_13_3319, i_13_3320, i_13_3321, i_13_3322, i_13_3323, i_13_3324, i_13_3325, i_13_3326, i_13_3327, i_13_3328, i_13_3329, i_13_3330, i_13_3331, i_13_3332, i_13_3333, i_13_3334, i_13_3335, i_13_3336, i_13_3337, i_13_3338, i_13_3339, i_13_3340, i_13_3341, i_13_3342, i_13_3343, i_13_3344, i_13_3345, i_13_3346, i_13_3347, i_13_3348, i_13_3349, i_13_3350, i_13_3351, i_13_3352, i_13_3353, i_13_3354, i_13_3355, i_13_3356, i_13_3357, i_13_3358, i_13_3359, i_13_3360, i_13_3361, i_13_3362, i_13_3363, i_13_3364, i_13_3365, i_13_3366, i_13_3367, i_13_3368, i_13_3369, i_13_3370, i_13_3371, i_13_3372, i_13_3373, i_13_3374, i_13_3375, i_13_3376, i_13_3377, i_13_3378, i_13_3379, i_13_3380, i_13_3381, i_13_3382, i_13_3383, i_13_3384, i_13_3385, i_13_3386, i_13_3387, i_13_3388, i_13_3389, i_13_3390, i_13_3391, i_13_3392, i_13_3393, i_13_3394, i_13_3395, i_13_3396, i_13_3397, i_13_3398, i_13_3399, i_13_3400, i_13_3401, i_13_3402, i_13_3403, i_13_3404, i_13_3405, i_13_3406, i_13_3407, i_13_3408, i_13_3409, i_13_3410, i_13_3411, i_13_3412, i_13_3413, i_13_3414, i_13_3415, i_13_3416, i_13_3417, i_13_3418, i_13_3419, i_13_3420, i_13_3421, i_13_3422, i_13_3423, i_13_3424, i_13_3425, i_13_3426, i_13_3427, i_13_3428, i_13_3429, i_13_3430, i_13_3431, i_13_3432, i_13_3433, i_13_3434, i_13_3435, i_13_3436, i_13_3437, i_13_3438, i_13_3439, i_13_3440, i_13_3441, i_13_3442, i_13_3443, i_13_3444, i_13_3445, i_13_3446, i_13_3447, i_13_3448, i_13_3449, i_13_3450, i_13_3451, i_13_3452, i_13_3453, i_13_3454, i_13_3455, i_13_3456, i_13_3457, i_13_3458, i_13_3459, i_13_3460, i_13_3461, i_13_3462, i_13_3463, i_13_3464, i_13_3465, i_13_3466, i_13_3467, i_13_3468, i_13_3469, i_13_3470, i_13_3471, i_13_3472, i_13_3473, i_13_3474, i_13_3475, i_13_3476, i_13_3477, i_13_3478, i_13_3479, i_13_3480, i_13_3481, i_13_3482, i_13_3483, i_13_3484, i_13_3485, i_13_3486, i_13_3487, i_13_3488, i_13_3489, i_13_3490, i_13_3491, i_13_3492, i_13_3493, i_13_3494, i_13_3495, i_13_3496, i_13_3497, i_13_3498, i_13_3499, i_13_3500, i_13_3501, i_13_3502, i_13_3503, i_13_3504, i_13_3505, i_13_3506, i_13_3507, i_13_3508, i_13_3509, i_13_3510, i_13_3511, i_13_3512, i_13_3513, i_13_3514, i_13_3515, i_13_3516, i_13_3517, i_13_3518, i_13_3519, i_13_3520, i_13_3521, i_13_3522, i_13_3523, i_13_3524, i_13_3525, i_13_3526, i_13_3527, i_13_3528, i_13_3529, i_13_3530, i_13_3531, i_13_3532, i_13_3533, i_13_3534, i_13_3535, i_13_3536, i_13_3537, i_13_3538, i_13_3539, i_13_3540, i_13_3541, i_13_3542, i_13_3543, i_13_3544, i_13_3545, i_13_3546, i_13_3547, i_13_3548, i_13_3549, i_13_3550, i_13_3551, i_13_3552, i_13_3553, i_13_3554, i_13_3555, i_13_3556, i_13_3557, i_13_3558, i_13_3559, i_13_3560, i_13_3561, i_13_3562, i_13_3563, i_13_3564, i_13_3565, i_13_3566, i_13_3567, i_13_3568, i_13_3569, i_13_3570, i_13_3571, i_13_3572, i_13_3573, i_13_3574, i_13_3575, i_13_3576, i_13_3577, i_13_3578, i_13_3579, i_13_3580, i_13_3581, i_13_3582, i_13_3583, i_13_3584, i_13_3585, i_13_3586, i_13_3587, i_13_3588, i_13_3589, i_13_3590, i_13_3591, i_13_3592, i_13_3593, i_13_3594, i_13_3595, i_13_3596, i_13_3597, i_13_3598, i_13_3599, i_13_3600, i_13_3601, i_13_3602, i_13_3603, i_13_3604, i_13_3605, i_13_3606, i_13_3607, i_13_3608, i_13_3609, i_13_3610, i_13_3611, i_13_3612, i_13_3613, i_13_3614, i_13_3615, i_13_3616, i_13_3617, i_13_3618, i_13_3619, i_13_3620, i_13_3621, i_13_3622, i_13_3623, i_13_3624, i_13_3625, i_13_3626, i_13_3627, i_13_3628, i_13_3629, i_13_3630, i_13_3631, i_13_3632, i_13_3633, i_13_3634, i_13_3635, i_13_3636, i_13_3637, i_13_3638, i_13_3639, i_13_3640, i_13_3641, i_13_3642, i_13_3643, i_13_3644, i_13_3645, i_13_3646, i_13_3647, i_13_3648, i_13_3649, i_13_3650, i_13_3651, i_13_3652, i_13_3653, i_13_3654, i_13_3655, i_13_3656, i_13_3657, i_13_3658, i_13_3659, i_13_3660, i_13_3661, i_13_3662, i_13_3663, i_13_3664, i_13_3665, i_13_3666, i_13_3667, i_13_3668, i_13_3669, i_13_3670, i_13_3671, i_13_3672, i_13_3673, i_13_3674, i_13_3675, i_13_3676, i_13_3677, i_13_3678, i_13_3679, i_13_3680, i_13_3681, i_13_3682, i_13_3683, i_13_3684, i_13_3685, i_13_3686, i_13_3687, i_13_3688, i_13_3689, i_13_3690, i_13_3691, i_13_3692, i_13_3693, i_13_3694, i_13_3695, i_13_3696, i_13_3697, i_13_3698, i_13_3699, i_13_3700, i_13_3701, i_13_3702, i_13_3703, i_13_3704, i_13_3705, i_13_3706, i_13_3707, i_13_3708, i_13_3709, i_13_3710, i_13_3711, i_13_3712, i_13_3713, i_13_3714, i_13_3715, i_13_3716, i_13_3717, i_13_3718, i_13_3719, i_13_3720, i_13_3721, i_13_3722, i_13_3723, i_13_3724, i_13_3725, i_13_3726, i_13_3727, i_13_3728, i_13_3729, i_13_3730, i_13_3731, i_13_3732, i_13_3733, i_13_3734, i_13_3735, i_13_3736, i_13_3737, i_13_3738, i_13_3739, i_13_3740, i_13_3741, i_13_3742, i_13_3743, i_13_3744, i_13_3745, i_13_3746, i_13_3747, i_13_3748, i_13_3749, i_13_3750, i_13_3751, i_13_3752, i_13_3753, i_13_3754, i_13_3755, i_13_3756, i_13_3757, i_13_3758, i_13_3759, i_13_3760, i_13_3761, i_13_3762, i_13_3763, i_13_3764, i_13_3765, i_13_3766, i_13_3767, i_13_3768, i_13_3769, i_13_3770, i_13_3771, i_13_3772, i_13_3773, i_13_3774, i_13_3775, i_13_3776, i_13_3777, i_13_3778, i_13_3779, i_13_3780, i_13_3781, i_13_3782, i_13_3783, i_13_3784, i_13_3785, i_13_3786, i_13_3787, i_13_3788, i_13_3789, i_13_3790, i_13_3791, i_13_3792, i_13_3793, i_13_3794, i_13_3795, i_13_3796, i_13_3797, i_13_3798, i_13_3799, i_13_3800, i_13_3801, i_13_3802, i_13_3803, i_13_3804, i_13_3805, i_13_3806, i_13_3807, i_13_3808, i_13_3809, i_13_3810, i_13_3811, i_13_3812, i_13_3813, i_13_3814, i_13_3815, i_13_3816, i_13_3817, i_13_3818, i_13_3819, i_13_3820, i_13_3821, i_13_3822, i_13_3823, i_13_3824, i_13_3825, i_13_3826, i_13_3827, i_13_3828, i_13_3829, i_13_3830, i_13_3831, i_13_3832, i_13_3833, i_13_3834, i_13_3835, i_13_3836, i_13_3837, i_13_3838, i_13_3839, i_13_3840, i_13_3841, i_13_3842, i_13_3843, i_13_3844, i_13_3845, i_13_3846, i_13_3847, i_13_3848, i_13_3849, i_13_3850, i_13_3851, i_13_3852, i_13_3853, i_13_3854, i_13_3855, i_13_3856, i_13_3857, i_13_3858, i_13_3859, i_13_3860, i_13_3861, i_13_3862, i_13_3863, i_13_3864, i_13_3865, i_13_3866, i_13_3867, i_13_3868, i_13_3869, i_13_3870, i_13_3871, i_13_3872, i_13_3873, i_13_3874, i_13_3875, i_13_3876, i_13_3877, i_13_3878, i_13_3879, i_13_3880, i_13_3881, i_13_3882, i_13_3883, i_13_3884, i_13_3885, i_13_3886, i_13_3887, i_13_3888, i_13_3889, i_13_3890, i_13_3891, i_13_3892, i_13_3893, i_13_3894, i_13_3895, i_13_3896, i_13_3897, i_13_3898, i_13_3899, i_13_3900, i_13_3901, i_13_3902, i_13_3903, i_13_3904, i_13_3905, i_13_3906, i_13_3907, i_13_3908, i_13_3909, i_13_3910, i_13_3911, i_13_3912, i_13_3913, i_13_3914, i_13_3915, i_13_3916, i_13_3917, i_13_3918, i_13_3919, i_13_3920, i_13_3921, i_13_3922, i_13_3923, i_13_3924, i_13_3925, i_13_3926, i_13_3927, i_13_3928, i_13_3929, i_13_3930, i_13_3931, i_13_3932, i_13_3933, i_13_3934, i_13_3935, i_13_3936, i_13_3937, i_13_3938, i_13_3939, i_13_3940, i_13_3941, i_13_3942, i_13_3943, i_13_3944, i_13_3945, i_13_3946, i_13_3947, i_13_3948, i_13_3949, i_13_3950, i_13_3951, i_13_3952, i_13_3953, i_13_3954, i_13_3955, i_13_3956, i_13_3957, i_13_3958, i_13_3959, i_13_3960, i_13_3961, i_13_3962, i_13_3963, i_13_3964, i_13_3965, i_13_3966, i_13_3967, i_13_3968, i_13_3969, i_13_3970, i_13_3971, i_13_3972, i_13_3973, i_13_3974, i_13_3975, i_13_3976, i_13_3977, i_13_3978, i_13_3979, i_13_3980, i_13_3981, i_13_3982, i_13_3983, i_13_3984, i_13_3985, i_13_3986, i_13_3987, i_13_3988, i_13_3989, i_13_3990, i_13_3991, i_13_3992, i_13_3993, i_13_3994, i_13_3995, i_13_3996, i_13_3997, i_13_3998, i_13_3999, i_13_4000, i_13_4001, i_13_4002, i_13_4003, i_13_4004, i_13_4005, i_13_4006, i_13_4007, i_13_4008, i_13_4009, i_13_4010, i_13_4011, i_13_4012, i_13_4013, i_13_4014, i_13_4015, i_13_4016, i_13_4017, i_13_4018, i_13_4019, i_13_4020, i_13_4021, i_13_4022, i_13_4023, i_13_4024, i_13_4025, i_13_4026, i_13_4027, i_13_4028, i_13_4029, i_13_4030, i_13_4031, i_13_4032, i_13_4033, i_13_4034, i_13_4035, i_13_4036, i_13_4037, i_13_4038, i_13_4039, i_13_4040, i_13_4041, i_13_4042, i_13_4043, i_13_4044, i_13_4045, i_13_4046, i_13_4047, i_13_4048, i_13_4049, i_13_4050, i_13_4051, i_13_4052, i_13_4053, i_13_4054, i_13_4055, i_13_4056, i_13_4057, i_13_4058, i_13_4059, i_13_4060, i_13_4061, i_13_4062, i_13_4063, i_13_4064, i_13_4065, i_13_4066, i_13_4067, i_13_4068, i_13_4069, i_13_4070, i_13_4071, i_13_4072, i_13_4073, i_13_4074, i_13_4075, i_13_4076, i_13_4077, i_13_4078, i_13_4079, i_13_4080, i_13_4081, i_13_4082, i_13_4083, i_13_4084, i_13_4085, i_13_4086, i_13_4087, i_13_4088, i_13_4089, i_13_4090, i_13_4091, i_13_4092, i_13_4093, i_13_4094, i_13_4095, i_13_4096, i_13_4097, i_13_4098, i_13_4099, i_13_4100, i_13_4101, i_13_4102, i_13_4103, i_13_4104, i_13_4105, i_13_4106, i_13_4107, i_13_4108, i_13_4109, i_13_4110, i_13_4111, i_13_4112, i_13_4113, i_13_4114, i_13_4115, i_13_4116, i_13_4117, i_13_4118, i_13_4119, i_13_4120, i_13_4121, i_13_4122, i_13_4123, i_13_4124, i_13_4125, i_13_4126, i_13_4127, i_13_4128, i_13_4129, i_13_4130, i_13_4131, i_13_4132, i_13_4133, i_13_4134, i_13_4135, i_13_4136, i_13_4137, i_13_4138, i_13_4139, i_13_4140, i_13_4141, i_13_4142, i_13_4143, i_13_4144, i_13_4145, i_13_4146, i_13_4147, i_13_4148, i_13_4149, i_13_4150, i_13_4151, i_13_4152, i_13_4153, i_13_4154, i_13_4155, i_13_4156, i_13_4157, i_13_4158, i_13_4159, i_13_4160, i_13_4161, i_13_4162, i_13_4163, i_13_4164, i_13_4165, i_13_4166, i_13_4167, i_13_4168, i_13_4169, i_13_4170, i_13_4171, i_13_4172, i_13_4173, i_13_4174, i_13_4175, i_13_4176, i_13_4177, i_13_4178, i_13_4179, i_13_4180, i_13_4181, i_13_4182, i_13_4183, i_13_4184, i_13_4185, i_13_4186, i_13_4187, i_13_4188, i_13_4189, i_13_4190, i_13_4191, i_13_4192, i_13_4193, i_13_4194, i_13_4195, i_13_4196, i_13_4197, i_13_4198, i_13_4199, i_13_4200, i_13_4201, i_13_4202, i_13_4203, i_13_4204, i_13_4205, i_13_4206, i_13_4207, i_13_4208, i_13_4209, i_13_4210, i_13_4211, i_13_4212, i_13_4213, i_13_4214, i_13_4215, i_13_4216, i_13_4217, i_13_4218, i_13_4219, i_13_4220, i_13_4221, i_13_4222, i_13_4223, i_13_4224, i_13_4225, i_13_4226, i_13_4227, i_13_4228, i_13_4229, i_13_4230, i_13_4231, i_13_4232, i_13_4233, i_13_4234, i_13_4235, i_13_4236, i_13_4237, i_13_4238, i_13_4239, i_13_4240, i_13_4241, i_13_4242, i_13_4243, i_13_4244, i_13_4245, i_13_4246, i_13_4247, i_13_4248, i_13_4249, i_13_4250, i_13_4251, i_13_4252, i_13_4253, i_13_4254, i_13_4255, i_13_4256, i_13_4257, i_13_4258, i_13_4259, i_13_4260, i_13_4261, i_13_4262, i_13_4263, i_13_4264, i_13_4265, i_13_4266, i_13_4267, i_13_4268, i_13_4269, i_13_4270, i_13_4271, i_13_4272, i_13_4273, i_13_4274, i_13_4275, i_13_4276, i_13_4277, i_13_4278, i_13_4279, i_13_4280, i_13_4281, i_13_4282, i_13_4283, i_13_4284, i_13_4285, i_13_4286, i_13_4287, i_13_4288, i_13_4289, i_13_4290, i_13_4291, i_13_4292, i_13_4293, i_13_4294, i_13_4295, i_13_4296, i_13_4297, i_13_4298, i_13_4299, i_13_4300, i_13_4301, i_13_4302, i_13_4303, i_13_4304, i_13_4305, i_13_4306, i_13_4307, i_13_4308, i_13_4309, i_13_4310, i_13_4311, i_13_4312, i_13_4313, i_13_4314, i_13_4315, i_13_4316, i_13_4317, i_13_4318, i_13_4319, i_13_4320, i_13_4321, i_13_4322, i_13_4323, i_13_4324, i_13_4325, i_13_4326, i_13_4327, i_13_4328, i_13_4329, i_13_4330, i_13_4331, i_13_4332, i_13_4333, i_13_4334, i_13_4335, i_13_4336, i_13_4337, i_13_4338, i_13_4339, i_13_4340, i_13_4341, i_13_4342, i_13_4343, i_13_4344, i_13_4345, i_13_4346, i_13_4347, i_13_4348, i_13_4349, i_13_4350, i_13_4351, i_13_4352, i_13_4353, i_13_4354, i_13_4355, i_13_4356, i_13_4357, i_13_4358, i_13_4359, i_13_4360, i_13_4361, i_13_4362, i_13_4363, i_13_4364, i_13_4365, i_13_4366, i_13_4367, i_13_4368, i_13_4369, i_13_4370, i_13_4371, i_13_4372, i_13_4373, i_13_4374, i_13_4375, i_13_4376, i_13_4377, i_13_4378, i_13_4379, i_13_4380, i_13_4381, i_13_4382, i_13_4383, i_13_4384, i_13_4385, i_13_4386, i_13_4387, i_13_4388, i_13_4389, i_13_4390, i_13_4391, i_13_4392, i_13_4393, i_13_4394, i_13_4395, i_13_4396, i_13_4397, i_13_4398, i_13_4399, i_13_4400, i_13_4401, i_13_4402, i_13_4403, i_13_4404, i_13_4405, i_13_4406, i_13_4407, i_13_4408, i_13_4409, i_13_4410, i_13_4411, i_13_4412, i_13_4413, i_13_4414, i_13_4415, i_13_4416, i_13_4417, i_13_4418, i_13_4419, i_13_4420, i_13_4421, i_13_4422, i_13_4423, i_13_4424, i_13_4425, i_13_4426, i_13_4427, i_13_4428, i_13_4429, i_13_4430, i_13_4431, i_13_4432, i_13_4433, i_13_4434, i_13_4435, i_13_4436, i_13_4437, i_13_4438, i_13_4439, i_13_4440, i_13_4441, i_13_4442, i_13_4443, i_13_4444, i_13_4445, i_13_4446, i_13_4447, i_13_4448, i_13_4449, i_13_4450, i_13_4451, i_13_4452, i_13_4453, i_13_4454, i_13_4455, i_13_4456, i_13_4457, i_13_4458, i_13_4459, i_13_4460, i_13_4461, i_13_4462, i_13_4463, i_13_4464, i_13_4465, i_13_4466, i_13_4467, i_13_4468, i_13_4469, i_13_4470, i_13_4471, i_13_4472, i_13_4473, i_13_4474, i_13_4475, i_13_4476, i_13_4477, i_13_4478, i_13_4479, i_13_4480, i_13_4481, i_13_4482, i_13_4483, i_13_4484, i_13_4485, i_13_4486, i_13_4487, i_13_4488, i_13_4489, i_13_4490, i_13_4491, i_13_4492, i_13_4493, i_13_4494, i_13_4495, i_13_4496, i_13_4497, i_13_4498, i_13_4499, i_13_4500, i_13_4501, i_13_4502, i_13_4503, i_13_4504, i_13_4505, i_13_4506, i_13_4507, i_13_4508, i_13_4509, i_13_4510, i_13_4511, i_13_4512, i_13_4513, i_13_4514, i_13_4515, i_13_4516, i_13_4517, i_13_4518, i_13_4519, i_13_4520, i_13_4521, i_13_4522, i_13_4523, i_13_4524, i_13_4525, i_13_4526, i_13_4527, i_13_4528, i_13_4529, i_13_4530, i_13_4531, i_13_4532, i_13_4533, i_13_4534, i_13_4535, i_13_4536, i_13_4537, i_13_4538, i_13_4539, i_13_4540, i_13_4541, i_13_4542, i_13_4543, i_13_4544, i_13_4545, i_13_4546, i_13_4547, i_13_4548, i_13_4549, i_13_4550, i_13_4551, i_13_4552, i_13_4553, i_13_4554, i_13_4555, i_13_4556, i_13_4557, i_13_4558, i_13_4559, i_13_4560, i_13_4561, i_13_4562, i_13_4563, i_13_4564, i_13_4565, i_13_4566, i_13_4567, i_13_4568, i_13_4569, i_13_4570, i_13_4571, i_13_4572, i_13_4573, i_13_4574, i_13_4575, i_13_4576, i_13_4577, i_13_4578, i_13_4579, i_13_4580, i_13_4581, i_13_4582, i_13_4583, i_13_4584, i_13_4585, i_13_4586, i_13_4587, i_13_4588, i_13_4589, i_13_4590, i_13_4591, i_13_4592, i_13_4593, i_13_4594, i_13_4595, i_13_4596, i_13_4597, i_13_4598, i_13_4599, i_13_4600, i_13_4601, i_13_4602, i_13_4603, i_13_4604, i_13_4605, i_13_4606, i_13_4607, o_13_0, o_13_1, o_13_2, o_13_3, o_13_4, o_13_5, o_13_6, o_13_7, o_13_8, o_13_9, o_13_10, o_13_11, o_13_12, o_13_13, o_13_14, o_13_15, o_13_16, o_13_17, o_13_18, o_13_19, o_13_20, o_13_21, o_13_22, o_13_23, o_13_24, o_13_25, o_13_26, o_13_27, o_13_28, o_13_29, o_13_30, o_13_31, o_13_32, o_13_33, o_13_34, o_13_35, o_13_36, o_13_37, o_13_38, o_13_39, o_13_40, o_13_41, o_13_42, o_13_43, o_13_44, o_13_45, o_13_46, o_13_47, o_13_48, o_13_49, o_13_50, o_13_51, o_13_52, o_13_53, o_13_54, o_13_55, o_13_56, o_13_57, o_13_58, o_13_59, o_13_60, o_13_61, o_13_62, o_13_63, o_13_64, o_13_65, o_13_66, o_13_67, o_13_68, o_13_69, o_13_70, o_13_71, o_13_72, o_13_73, o_13_74, o_13_75, o_13_76, o_13_77, o_13_78, o_13_79, o_13_80, o_13_81, o_13_82, o_13_83, o_13_84, o_13_85, o_13_86, o_13_87, o_13_88, o_13_89, o_13_90, o_13_91, o_13_92, o_13_93, o_13_94, o_13_95, o_13_96, o_13_97, o_13_98, o_13_99, o_13_100, o_13_101, o_13_102, o_13_103, o_13_104, o_13_105, o_13_106, o_13_107, o_13_108, o_13_109, o_13_110, o_13_111, o_13_112, o_13_113, o_13_114, o_13_115, o_13_116, o_13_117, o_13_118, o_13_119, o_13_120, o_13_121, o_13_122, o_13_123, o_13_124, o_13_125, o_13_126, o_13_127, o_13_128, o_13_129, o_13_130, o_13_131, o_13_132, o_13_133, o_13_134, o_13_135, o_13_136, o_13_137, o_13_138, o_13_139, o_13_140, o_13_141, o_13_142, o_13_143, o_13_144, o_13_145, o_13_146, o_13_147, o_13_148, o_13_149, o_13_150, o_13_151, o_13_152, o_13_153, o_13_154, o_13_155, o_13_156, o_13_157, o_13_158, o_13_159, o_13_160, o_13_161, o_13_162, o_13_163, o_13_164, o_13_165, o_13_166, o_13_167, o_13_168, o_13_169, o_13_170, o_13_171, o_13_172, o_13_173, o_13_174, o_13_175, o_13_176, o_13_177, o_13_178, o_13_179, o_13_180, o_13_181, o_13_182, o_13_183, o_13_184, o_13_185, o_13_186, o_13_187, o_13_188, o_13_189, o_13_190, o_13_191, o_13_192, o_13_193, o_13_194, o_13_195, o_13_196, o_13_197, o_13_198, o_13_199, o_13_200, o_13_201, o_13_202, o_13_203, o_13_204, o_13_205, o_13_206, o_13_207, o_13_208, o_13_209, o_13_210, o_13_211, o_13_212, o_13_213, o_13_214, o_13_215, o_13_216, o_13_217, o_13_218, o_13_219, o_13_220, o_13_221, o_13_222, o_13_223, o_13_224, o_13_225, o_13_226, o_13_227, o_13_228, o_13_229, o_13_230, o_13_231, o_13_232, o_13_233, o_13_234, o_13_235, o_13_236, o_13_237, o_13_238, o_13_239, o_13_240, o_13_241, o_13_242, o_13_243, o_13_244, o_13_245, o_13_246, o_13_247, o_13_248, o_13_249, o_13_250, o_13_251, o_13_252, o_13_253, o_13_254, o_13_255, o_13_256, o_13_257, o_13_258, o_13_259, o_13_260, o_13_261, o_13_262, o_13_263, o_13_264, o_13_265, o_13_266, o_13_267, o_13_268, o_13_269, o_13_270, o_13_271, o_13_272, o_13_273, o_13_274, o_13_275, o_13_276, o_13_277, o_13_278, o_13_279, o_13_280, o_13_281, o_13_282, o_13_283, o_13_284, o_13_285, o_13_286, o_13_287, o_13_288, o_13_289, o_13_290, o_13_291, o_13_292, o_13_293, o_13_294, o_13_295, o_13_296, o_13_297, o_13_298, o_13_299, o_13_300, o_13_301, o_13_302, o_13_303, o_13_304, o_13_305, o_13_306, o_13_307, o_13_308, o_13_309, o_13_310, o_13_311, o_13_312, o_13_313, o_13_314, o_13_315, o_13_316, o_13_317, o_13_318, o_13_319, o_13_320, o_13_321, o_13_322, o_13_323, o_13_324, o_13_325, o_13_326, o_13_327, o_13_328, o_13_329, o_13_330, o_13_331, o_13_332, o_13_333, o_13_334, o_13_335, o_13_336, o_13_337, o_13_338, o_13_339, o_13_340, o_13_341, o_13_342, o_13_343, o_13_344, o_13_345, o_13_346, o_13_347, o_13_348, o_13_349, o_13_350, o_13_351, o_13_352, o_13_353, o_13_354, o_13_355, o_13_356, o_13_357, o_13_358, o_13_359, o_13_360, o_13_361, o_13_362, o_13_363, o_13_364, o_13_365, o_13_366, o_13_367, o_13_368, o_13_369, o_13_370, o_13_371, o_13_372, o_13_373, o_13_374, o_13_375, o_13_376, o_13_377, o_13_378, o_13_379, o_13_380, o_13_381, o_13_382, o_13_383, o_13_384, o_13_385, o_13_386, o_13_387, o_13_388, o_13_389, o_13_390, o_13_391, o_13_392, o_13_393, o_13_394, o_13_395, o_13_396, o_13_397, o_13_398, o_13_399, o_13_400, o_13_401, o_13_402, o_13_403, o_13_404, o_13_405, o_13_406, o_13_407, o_13_408, o_13_409, o_13_410, o_13_411, o_13_412, o_13_413, o_13_414, o_13_415, o_13_416, o_13_417, o_13_418, o_13_419, o_13_420, o_13_421, o_13_422, o_13_423, o_13_424, o_13_425, o_13_426, o_13_427, o_13_428, o_13_429, o_13_430, o_13_431, o_13_432, o_13_433, o_13_434, o_13_435, o_13_436, o_13_437, o_13_438, o_13_439, o_13_440, o_13_441, o_13_442, o_13_443, o_13_444, o_13_445, o_13_446, o_13_447, o_13_448, o_13_449, o_13_450, o_13_451, o_13_452, o_13_453, o_13_454, o_13_455, o_13_456, o_13_457, o_13_458, o_13_459, o_13_460, o_13_461, o_13_462, o_13_463, o_13_464, o_13_465, o_13_466, o_13_467, o_13_468, o_13_469, o_13_470, o_13_471, o_13_472, o_13_473, o_13_474, o_13_475, o_13_476, o_13_477, o_13_478, o_13_479, o_13_480, o_13_481, o_13_482, o_13_483, o_13_484, o_13_485, o_13_486, o_13_487, o_13_488, o_13_489, o_13_490, o_13_491, o_13_492, o_13_493, o_13_494, o_13_495, o_13_496, o_13_497, o_13_498, o_13_499, o_13_500, o_13_501, o_13_502, o_13_503, o_13_504, o_13_505, o_13_506, o_13_507, o_13_508, o_13_509, o_13_510, o_13_511);

  always @ (posedge ap_clk)
    if (ap_rst)
      begin
        out_reg <= 0;
        i_13_0 <= 0;
        i_13_1 <= 0;
        i_13_2 <= 0;
        i_13_3 <= 0;
        i_13_4 <= 0;
        i_13_5 <= 0;
        i_13_6 <= 0;
        i_13_7 <= 0;
        i_13_8 <= 0;
        i_13_9 <= 0;
        i_13_10 <= 0;
        i_13_11 <= 0;
        i_13_12 <= 0;
        i_13_13 <= 0;
        i_13_14 <= 0;
        i_13_15 <= 0;
        i_13_16 <= 0;
        i_13_17 <= 0;
        i_13_18 <= 0;
        i_13_19 <= 0;
        i_13_20 <= 0;
        i_13_21 <= 0;
        i_13_22 <= 0;
        i_13_23 <= 0;
        i_13_24 <= 0;
        i_13_25 <= 0;
        i_13_26 <= 0;
        i_13_27 <= 0;
        i_13_28 <= 0;
        i_13_29 <= 0;
        i_13_30 <= 0;
        i_13_31 <= 0;
        i_13_32 <= 0;
        i_13_33 <= 0;
        i_13_34 <= 0;
        i_13_35 <= 0;
        i_13_36 <= 0;
        i_13_37 <= 0;
        i_13_38 <= 0;
        i_13_39 <= 0;
        i_13_40 <= 0;
        i_13_41 <= 0;
        i_13_42 <= 0;
        i_13_43 <= 0;
        i_13_44 <= 0;
        i_13_45 <= 0;
        i_13_46 <= 0;
        i_13_47 <= 0;
        i_13_48 <= 0;
        i_13_49 <= 0;
        i_13_50 <= 0;
        i_13_51 <= 0;
        i_13_52 <= 0;
        i_13_53 <= 0;
        i_13_54 <= 0;
        i_13_55 <= 0;
        i_13_56 <= 0;
        i_13_57 <= 0;
        i_13_58 <= 0;
        i_13_59 <= 0;
        i_13_60 <= 0;
        i_13_61 <= 0;
        i_13_62 <= 0;
        i_13_63 <= 0;
        i_13_64 <= 0;
        i_13_65 <= 0;
        i_13_66 <= 0;
        i_13_67 <= 0;
        i_13_68 <= 0;
        i_13_69 <= 0;
        i_13_70 <= 0;
        i_13_71 <= 0;
        i_13_72 <= 0;
        i_13_73 <= 0;
        i_13_74 <= 0;
        i_13_75 <= 0;
        i_13_76 <= 0;
        i_13_77 <= 0;
        i_13_78 <= 0;
        i_13_79 <= 0;
        i_13_80 <= 0;
        i_13_81 <= 0;
        i_13_82 <= 0;
        i_13_83 <= 0;
        i_13_84 <= 0;
        i_13_85 <= 0;
        i_13_86 <= 0;
        i_13_87 <= 0;
        i_13_88 <= 0;
        i_13_89 <= 0;
        i_13_90 <= 0;
        i_13_91 <= 0;
        i_13_92 <= 0;
        i_13_93 <= 0;
        i_13_94 <= 0;
        i_13_95 <= 0;
        i_13_96 <= 0;
        i_13_97 <= 0;
        i_13_98 <= 0;
        i_13_99 <= 0;
        i_13_100 <= 0;
        i_13_101 <= 0;
        i_13_102 <= 0;
        i_13_103 <= 0;
        i_13_104 <= 0;
        i_13_105 <= 0;
        i_13_106 <= 0;
        i_13_107 <= 0;
        i_13_108 <= 0;
        i_13_109 <= 0;
        i_13_110 <= 0;
        i_13_111 <= 0;
        i_13_112 <= 0;
        i_13_113 <= 0;
        i_13_114 <= 0;
        i_13_115 <= 0;
        i_13_116 <= 0;
        i_13_117 <= 0;
        i_13_118 <= 0;
        i_13_119 <= 0;
        i_13_120 <= 0;
        i_13_121 <= 0;
        i_13_122 <= 0;
        i_13_123 <= 0;
        i_13_124 <= 0;
        i_13_125 <= 0;
        i_13_126 <= 0;
        i_13_127 <= 0;
        i_13_128 <= 0;
        i_13_129 <= 0;
        i_13_130 <= 0;
        i_13_131 <= 0;
        i_13_132 <= 0;
        i_13_133 <= 0;
        i_13_134 <= 0;
        i_13_135 <= 0;
        i_13_136 <= 0;
        i_13_137 <= 0;
        i_13_138 <= 0;
        i_13_139 <= 0;
        i_13_140 <= 0;
        i_13_141 <= 0;
        i_13_142 <= 0;
        i_13_143 <= 0;
        i_13_144 <= 0;
        i_13_145 <= 0;
        i_13_146 <= 0;
        i_13_147 <= 0;
        i_13_148 <= 0;
        i_13_149 <= 0;
        i_13_150 <= 0;
        i_13_151 <= 0;
        i_13_152 <= 0;
        i_13_153 <= 0;
        i_13_154 <= 0;
        i_13_155 <= 0;
        i_13_156 <= 0;
        i_13_157 <= 0;
        i_13_158 <= 0;
        i_13_159 <= 0;
        i_13_160 <= 0;
        i_13_161 <= 0;
        i_13_162 <= 0;
        i_13_163 <= 0;
        i_13_164 <= 0;
        i_13_165 <= 0;
        i_13_166 <= 0;
        i_13_167 <= 0;
        i_13_168 <= 0;
        i_13_169 <= 0;
        i_13_170 <= 0;
        i_13_171 <= 0;
        i_13_172 <= 0;
        i_13_173 <= 0;
        i_13_174 <= 0;
        i_13_175 <= 0;
        i_13_176 <= 0;
        i_13_177 <= 0;
        i_13_178 <= 0;
        i_13_179 <= 0;
        i_13_180 <= 0;
        i_13_181 <= 0;
        i_13_182 <= 0;
        i_13_183 <= 0;
        i_13_184 <= 0;
        i_13_185 <= 0;
        i_13_186 <= 0;
        i_13_187 <= 0;
        i_13_188 <= 0;
        i_13_189 <= 0;
        i_13_190 <= 0;
        i_13_191 <= 0;
        i_13_192 <= 0;
        i_13_193 <= 0;
        i_13_194 <= 0;
        i_13_195 <= 0;
        i_13_196 <= 0;
        i_13_197 <= 0;
        i_13_198 <= 0;
        i_13_199 <= 0;
        i_13_200 <= 0;
        i_13_201 <= 0;
        i_13_202 <= 0;
        i_13_203 <= 0;
        i_13_204 <= 0;
        i_13_205 <= 0;
        i_13_206 <= 0;
        i_13_207 <= 0;
        i_13_208 <= 0;
        i_13_209 <= 0;
        i_13_210 <= 0;
        i_13_211 <= 0;
        i_13_212 <= 0;
        i_13_213 <= 0;
        i_13_214 <= 0;
        i_13_215 <= 0;
        i_13_216 <= 0;
        i_13_217 <= 0;
        i_13_218 <= 0;
        i_13_219 <= 0;
        i_13_220 <= 0;
        i_13_221 <= 0;
        i_13_222 <= 0;
        i_13_223 <= 0;
        i_13_224 <= 0;
        i_13_225 <= 0;
        i_13_226 <= 0;
        i_13_227 <= 0;
        i_13_228 <= 0;
        i_13_229 <= 0;
        i_13_230 <= 0;
        i_13_231 <= 0;
        i_13_232 <= 0;
        i_13_233 <= 0;
        i_13_234 <= 0;
        i_13_235 <= 0;
        i_13_236 <= 0;
        i_13_237 <= 0;
        i_13_238 <= 0;
        i_13_239 <= 0;
        i_13_240 <= 0;
        i_13_241 <= 0;
        i_13_242 <= 0;
        i_13_243 <= 0;
        i_13_244 <= 0;
        i_13_245 <= 0;
        i_13_246 <= 0;
        i_13_247 <= 0;
        i_13_248 <= 0;
        i_13_249 <= 0;
        i_13_250 <= 0;
        i_13_251 <= 0;
        i_13_252 <= 0;
        i_13_253 <= 0;
        i_13_254 <= 0;
        i_13_255 <= 0;
        i_13_256 <= 0;
        i_13_257 <= 0;
        i_13_258 <= 0;
        i_13_259 <= 0;
        i_13_260 <= 0;
        i_13_261 <= 0;
        i_13_262 <= 0;
        i_13_263 <= 0;
        i_13_264 <= 0;
        i_13_265 <= 0;
        i_13_266 <= 0;
        i_13_267 <= 0;
        i_13_268 <= 0;
        i_13_269 <= 0;
        i_13_270 <= 0;
        i_13_271 <= 0;
        i_13_272 <= 0;
        i_13_273 <= 0;
        i_13_274 <= 0;
        i_13_275 <= 0;
        i_13_276 <= 0;
        i_13_277 <= 0;
        i_13_278 <= 0;
        i_13_279 <= 0;
        i_13_280 <= 0;
        i_13_281 <= 0;
        i_13_282 <= 0;
        i_13_283 <= 0;
        i_13_284 <= 0;
        i_13_285 <= 0;
        i_13_286 <= 0;
        i_13_287 <= 0;
        i_13_288 <= 0;
        i_13_289 <= 0;
        i_13_290 <= 0;
        i_13_291 <= 0;
        i_13_292 <= 0;
        i_13_293 <= 0;
        i_13_294 <= 0;
        i_13_295 <= 0;
        i_13_296 <= 0;
        i_13_297 <= 0;
        i_13_298 <= 0;
        i_13_299 <= 0;
        i_13_300 <= 0;
        i_13_301 <= 0;
        i_13_302 <= 0;
        i_13_303 <= 0;
        i_13_304 <= 0;
        i_13_305 <= 0;
        i_13_306 <= 0;
        i_13_307 <= 0;
        i_13_308 <= 0;
        i_13_309 <= 0;
        i_13_310 <= 0;
        i_13_311 <= 0;
        i_13_312 <= 0;
        i_13_313 <= 0;
        i_13_314 <= 0;
        i_13_315 <= 0;
        i_13_316 <= 0;
        i_13_317 <= 0;
        i_13_318 <= 0;
        i_13_319 <= 0;
        i_13_320 <= 0;
        i_13_321 <= 0;
        i_13_322 <= 0;
        i_13_323 <= 0;
        i_13_324 <= 0;
        i_13_325 <= 0;
        i_13_326 <= 0;
        i_13_327 <= 0;
        i_13_328 <= 0;
        i_13_329 <= 0;
        i_13_330 <= 0;
        i_13_331 <= 0;
        i_13_332 <= 0;
        i_13_333 <= 0;
        i_13_334 <= 0;
        i_13_335 <= 0;
        i_13_336 <= 0;
        i_13_337 <= 0;
        i_13_338 <= 0;
        i_13_339 <= 0;
        i_13_340 <= 0;
        i_13_341 <= 0;
        i_13_342 <= 0;
        i_13_343 <= 0;
        i_13_344 <= 0;
        i_13_345 <= 0;
        i_13_346 <= 0;
        i_13_347 <= 0;
        i_13_348 <= 0;
        i_13_349 <= 0;
        i_13_350 <= 0;
        i_13_351 <= 0;
        i_13_352 <= 0;
        i_13_353 <= 0;
        i_13_354 <= 0;
        i_13_355 <= 0;
        i_13_356 <= 0;
        i_13_357 <= 0;
        i_13_358 <= 0;
        i_13_359 <= 0;
        i_13_360 <= 0;
        i_13_361 <= 0;
        i_13_362 <= 0;
        i_13_363 <= 0;
        i_13_364 <= 0;
        i_13_365 <= 0;
        i_13_366 <= 0;
        i_13_367 <= 0;
        i_13_368 <= 0;
        i_13_369 <= 0;
        i_13_370 <= 0;
        i_13_371 <= 0;
        i_13_372 <= 0;
        i_13_373 <= 0;
        i_13_374 <= 0;
        i_13_375 <= 0;
        i_13_376 <= 0;
        i_13_377 <= 0;
        i_13_378 <= 0;
        i_13_379 <= 0;
        i_13_380 <= 0;
        i_13_381 <= 0;
        i_13_382 <= 0;
        i_13_383 <= 0;
        i_13_384 <= 0;
        i_13_385 <= 0;
        i_13_386 <= 0;
        i_13_387 <= 0;
        i_13_388 <= 0;
        i_13_389 <= 0;
        i_13_390 <= 0;
        i_13_391 <= 0;
        i_13_392 <= 0;
        i_13_393 <= 0;
        i_13_394 <= 0;
        i_13_395 <= 0;
        i_13_396 <= 0;
        i_13_397 <= 0;
        i_13_398 <= 0;
        i_13_399 <= 0;
        i_13_400 <= 0;
        i_13_401 <= 0;
        i_13_402 <= 0;
        i_13_403 <= 0;
        i_13_404 <= 0;
        i_13_405 <= 0;
        i_13_406 <= 0;
        i_13_407 <= 0;
        i_13_408 <= 0;
        i_13_409 <= 0;
        i_13_410 <= 0;
        i_13_411 <= 0;
        i_13_412 <= 0;
        i_13_413 <= 0;
        i_13_414 <= 0;
        i_13_415 <= 0;
        i_13_416 <= 0;
        i_13_417 <= 0;
        i_13_418 <= 0;
        i_13_419 <= 0;
        i_13_420 <= 0;
        i_13_421 <= 0;
        i_13_422 <= 0;
        i_13_423 <= 0;
        i_13_424 <= 0;
        i_13_425 <= 0;
        i_13_426 <= 0;
        i_13_427 <= 0;
        i_13_428 <= 0;
        i_13_429 <= 0;
        i_13_430 <= 0;
        i_13_431 <= 0;
        i_13_432 <= 0;
        i_13_433 <= 0;
        i_13_434 <= 0;
        i_13_435 <= 0;
        i_13_436 <= 0;
        i_13_437 <= 0;
        i_13_438 <= 0;
        i_13_439 <= 0;
        i_13_440 <= 0;
        i_13_441 <= 0;
        i_13_442 <= 0;
        i_13_443 <= 0;
        i_13_444 <= 0;
        i_13_445 <= 0;
        i_13_446 <= 0;
        i_13_447 <= 0;
        i_13_448 <= 0;
        i_13_449 <= 0;
        i_13_450 <= 0;
        i_13_451 <= 0;
        i_13_452 <= 0;
        i_13_453 <= 0;
        i_13_454 <= 0;
        i_13_455 <= 0;
        i_13_456 <= 0;
        i_13_457 <= 0;
        i_13_458 <= 0;
        i_13_459 <= 0;
        i_13_460 <= 0;
        i_13_461 <= 0;
        i_13_462 <= 0;
        i_13_463 <= 0;
        i_13_464 <= 0;
        i_13_465 <= 0;
        i_13_466 <= 0;
        i_13_467 <= 0;
        i_13_468 <= 0;
        i_13_469 <= 0;
        i_13_470 <= 0;
        i_13_471 <= 0;
        i_13_472 <= 0;
        i_13_473 <= 0;
        i_13_474 <= 0;
        i_13_475 <= 0;
        i_13_476 <= 0;
        i_13_477 <= 0;
        i_13_478 <= 0;
        i_13_479 <= 0;
        i_13_480 <= 0;
        i_13_481 <= 0;
        i_13_482 <= 0;
        i_13_483 <= 0;
        i_13_484 <= 0;
        i_13_485 <= 0;
        i_13_486 <= 0;
        i_13_487 <= 0;
        i_13_488 <= 0;
        i_13_489 <= 0;
        i_13_490 <= 0;
        i_13_491 <= 0;
        i_13_492 <= 0;
        i_13_493 <= 0;
        i_13_494 <= 0;
        i_13_495 <= 0;
        i_13_496 <= 0;
        i_13_497 <= 0;
        i_13_498 <= 0;
        i_13_499 <= 0;
        i_13_500 <= 0;
        i_13_501 <= 0;
        i_13_502 <= 0;
        i_13_503 <= 0;
        i_13_504 <= 0;
        i_13_505 <= 0;
        i_13_506 <= 0;
        i_13_507 <= 0;
        i_13_508 <= 0;
        i_13_509 <= 0;
        i_13_510 <= 0;
        i_13_511 <= 0;
        i_13_512 <= 0;
        i_13_513 <= 0;
        i_13_514 <= 0;
        i_13_515 <= 0;
        i_13_516 <= 0;
        i_13_517 <= 0;
        i_13_518 <= 0;
        i_13_519 <= 0;
        i_13_520 <= 0;
        i_13_521 <= 0;
        i_13_522 <= 0;
        i_13_523 <= 0;
        i_13_524 <= 0;
        i_13_525 <= 0;
        i_13_526 <= 0;
        i_13_527 <= 0;
        i_13_528 <= 0;
        i_13_529 <= 0;
        i_13_530 <= 0;
        i_13_531 <= 0;
        i_13_532 <= 0;
        i_13_533 <= 0;
        i_13_534 <= 0;
        i_13_535 <= 0;
        i_13_536 <= 0;
        i_13_537 <= 0;
        i_13_538 <= 0;
        i_13_539 <= 0;
        i_13_540 <= 0;
        i_13_541 <= 0;
        i_13_542 <= 0;
        i_13_543 <= 0;
        i_13_544 <= 0;
        i_13_545 <= 0;
        i_13_546 <= 0;
        i_13_547 <= 0;
        i_13_548 <= 0;
        i_13_549 <= 0;
        i_13_550 <= 0;
        i_13_551 <= 0;
        i_13_552 <= 0;
        i_13_553 <= 0;
        i_13_554 <= 0;
        i_13_555 <= 0;
        i_13_556 <= 0;
        i_13_557 <= 0;
        i_13_558 <= 0;
        i_13_559 <= 0;
        i_13_560 <= 0;
        i_13_561 <= 0;
        i_13_562 <= 0;
        i_13_563 <= 0;
        i_13_564 <= 0;
        i_13_565 <= 0;
        i_13_566 <= 0;
        i_13_567 <= 0;
        i_13_568 <= 0;
        i_13_569 <= 0;
        i_13_570 <= 0;
        i_13_571 <= 0;
        i_13_572 <= 0;
        i_13_573 <= 0;
        i_13_574 <= 0;
        i_13_575 <= 0;
        i_13_576 <= 0;
        i_13_577 <= 0;
        i_13_578 <= 0;
        i_13_579 <= 0;
        i_13_580 <= 0;
        i_13_581 <= 0;
        i_13_582 <= 0;
        i_13_583 <= 0;
        i_13_584 <= 0;
        i_13_585 <= 0;
        i_13_586 <= 0;
        i_13_587 <= 0;
        i_13_588 <= 0;
        i_13_589 <= 0;
        i_13_590 <= 0;
        i_13_591 <= 0;
        i_13_592 <= 0;
        i_13_593 <= 0;
        i_13_594 <= 0;
        i_13_595 <= 0;
        i_13_596 <= 0;
        i_13_597 <= 0;
        i_13_598 <= 0;
        i_13_599 <= 0;
        i_13_600 <= 0;
        i_13_601 <= 0;
        i_13_602 <= 0;
        i_13_603 <= 0;
        i_13_604 <= 0;
        i_13_605 <= 0;
        i_13_606 <= 0;
        i_13_607 <= 0;
        i_13_608 <= 0;
        i_13_609 <= 0;
        i_13_610 <= 0;
        i_13_611 <= 0;
        i_13_612 <= 0;
        i_13_613 <= 0;
        i_13_614 <= 0;
        i_13_615 <= 0;
        i_13_616 <= 0;
        i_13_617 <= 0;
        i_13_618 <= 0;
        i_13_619 <= 0;
        i_13_620 <= 0;
        i_13_621 <= 0;
        i_13_622 <= 0;
        i_13_623 <= 0;
        i_13_624 <= 0;
        i_13_625 <= 0;
        i_13_626 <= 0;
        i_13_627 <= 0;
        i_13_628 <= 0;
        i_13_629 <= 0;
        i_13_630 <= 0;
        i_13_631 <= 0;
        i_13_632 <= 0;
        i_13_633 <= 0;
        i_13_634 <= 0;
        i_13_635 <= 0;
        i_13_636 <= 0;
        i_13_637 <= 0;
        i_13_638 <= 0;
        i_13_639 <= 0;
        i_13_640 <= 0;
        i_13_641 <= 0;
        i_13_642 <= 0;
        i_13_643 <= 0;
        i_13_644 <= 0;
        i_13_645 <= 0;
        i_13_646 <= 0;
        i_13_647 <= 0;
        i_13_648 <= 0;
        i_13_649 <= 0;
        i_13_650 <= 0;
        i_13_651 <= 0;
        i_13_652 <= 0;
        i_13_653 <= 0;
        i_13_654 <= 0;
        i_13_655 <= 0;
        i_13_656 <= 0;
        i_13_657 <= 0;
        i_13_658 <= 0;
        i_13_659 <= 0;
        i_13_660 <= 0;
        i_13_661 <= 0;
        i_13_662 <= 0;
        i_13_663 <= 0;
        i_13_664 <= 0;
        i_13_665 <= 0;
        i_13_666 <= 0;
        i_13_667 <= 0;
        i_13_668 <= 0;
        i_13_669 <= 0;
        i_13_670 <= 0;
        i_13_671 <= 0;
        i_13_672 <= 0;
        i_13_673 <= 0;
        i_13_674 <= 0;
        i_13_675 <= 0;
        i_13_676 <= 0;
        i_13_677 <= 0;
        i_13_678 <= 0;
        i_13_679 <= 0;
        i_13_680 <= 0;
        i_13_681 <= 0;
        i_13_682 <= 0;
        i_13_683 <= 0;
        i_13_684 <= 0;
        i_13_685 <= 0;
        i_13_686 <= 0;
        i_13_687 <= 0;
        i_13_688 <= 0;
        i_13_689 <= 0;
        i_13_690 <= 0;
        i_13_691 <= 0;
        i_13_692 <= 0;
        i_13_693 <= 0;
        i_13_694 <= 0;
        i_13_695 <= 0;
        i_13_696 <= 0;
        i_13_697 <= 0;
        i_13_698 <= 0;
        i_13_699 <= 0;
        i_13_700 <= 0;
        i_13_701 <= 0;
        i_13_702 <= 0;
        i_13_703 <= 0;
        i_13_704 <= 0;
        i_13_705 <= 0;
        i_13_706 <= 0;
        i_13_707 <= 0;
        i_13_708 <= 0;
        i_13_709 <= 0;
        i_13_710 <= 0;
        i_13_711 <= 0;
        i_13_712 <= 0;
        i_13_713 <= 0;
        i_13_714 <= 0;
        i_13_715 <= 0;
        i_13_716 <= 0;
        i_13_717 <= 0;
        i_13_718 <= 0;
        i_13_719 <= 0;
        i_13_720 <= 0;
        i_13_721 <= 0;
        i_13_722 <= 0;
        i_13_723 <= 0;
        i_13_724 <= 0;
        i_13_725 <= 0;
        i_13_726 <= 0;
        i_13_727 <= 0;
        i_13_728 <= 0;
        i_13_729 <= 0;
        i_13_730 <= 0;
        i_13_731 <= 0;
        i_13_732 <= 0;
        i_13_733 <= 0;
        i_13_734 <= 0;
        i_13_735 <= 0;
        i_13_736 <= 0;
        i_13_737 <= 0;
        i_13_738 <= 0;
        i_13_739 <= 0;
        i_13_740 <= 0;
        i_13_741 <= 0;
        i_13_742 <= 0;
        i_13_743 <= 0;
        i_13_744 <= 0;
        i_13_745 <= 0;
        i_13_746 <= 0;
        i_13_747 <= 0;
        i_13_748 <= 0;
        i_13_749 <= 0;
        i_13_750 <= 0;
        i_13_751 <= 0;
        i_13_752 <= 0;
        i_13_753 <= 0;
        i_13_754 <= 0;
        i_13_755 <= 0;
        i_13_756 <= 0;
        i_13_757 <= 0;
        i_13_758 <= 0;
        i_13_759 <= 0;
        i_13_760 <= 0;
        i_13_761 <= 0;
        i_13_762 <= 0;
        i_13_763 <= 0;
        i_13_764 <= 0;
        i_13_765 <= 0;
        i_13_766 <= 0;
        i_13_767 <= 0;
        i_13_768 <= 0;
        i_13_769 <= 0;
        i_13_770 <= 0;
        i_13_771 <= 0;
        i_13_772 <= 0;
        i_13_773 <= 0;
        i_13_774 <= 0;
        i_13_775 <= 0;
        i_13_776 <= 0;
        i_13_777 <= 0;
        i_13_778 <= 0;
        i_13_779 <= 0;
        i_13_780 <= 0;
        i_13_781 <= 0;
        i_13_782 <= 0;
        i_13_783 <= 0;
        i_13_784 <= 0;
        i_13_785 <= 0;
        i_13_786 <= 0;
        i_13_787 <= 0;
        i_13_788 <= 0;
        i_13_789 <= 0;
        i_13_790 <= 0;
        i_13_791 <= 0;
        i_13_792 <= 0;
        i_13_793 <= 0;
        i_13_794 <= 0;
        i_13_795 <= 0;
        i_13_796 <= 0;
        i_13_797 <= 0;
        i_13_798 <= 0;
        i_13_799 <= 0;
        i_13_800 <= 0;
        i_13_801 <= 0;
        i_13_802 <= 0;
        i_13_803 <= 0;
        i_13_804 <= 0;
        i_13_805 <= 0;
        i_13_806 <= 0;
        i_13_807 <= 0;
        i_13_808 <= 0;
        i_13_809 <= 0;
        i_13_810 <= 0;
        i_13_811 <= 0;
        i_13_812 <= 0;
        i_13_813 <= 0;
        i_13_814 <= 0;
        i_13_815 <= 0;
        i_13_816 <= 0;
        i_13_817 <= 0;
        i_13_818 <= 0;
        i_13_819 <= 0;
        i_13_820 <= 0;
        i_13_821 <= 0;
        i_13_822 <= 0;
        i_13_823 <= 0;
        i_13_824 <= 0;
        i_13_825 <= 0;
        i_13_826 <= 0;
        i_13_827 <= 0;
        i_13_828 <= 0;
        i_13_829 <= 0;
        i_13_830 <= 0;
        i_13_831 <= 0;
        i_13_832 <= 0;
        i_13_833 <= 0;
        i_13_834 <= 0;
        i_13_835 <= 0;
        i_13_836 <= 0;
        i_13_837 <= 0;
        i_13_838 <= 0;
        i_13_839 <= 0;
        i_13_840 <= 0;
        i_13_841 <= 0;
        i_13_842 <= 0;
        i_13_843 <= 0;
        i_13_844 <= 0;
        i_13_845 <= 0;
        i_13_846 <= 0;
        i_13_847 <= 0;
        i_13_848 <= 0;
        i_13_849 <= 0;
        i_13_850 <= 0;
        i_13_851 <= 0;
        i_13_852 <= 0;
        i_13_853 <= 0;
        i_13_854 <= 0;
        i_13_855 <= 0;
        i_13_856 <= 0;
        i_13_857 <= 0;
        i_13_858 <= 0;
        i_13_859 <= 0;
        i_13_860 <= 0;
        i_13_861 <= 0;
        i_13_862 <= 0;
        i_13_863 <= 0;
        i_13_864 <= 0;
        i_13_865 <= 0;
        i_13_866 <= 0;
        i_13_867 <= 0;
        i_13_868 <= 0;
        i_13_869 <= 0;
        i_13_870 <= 0;
        i_13_871 <= 0;
        i_13_872 <= 0;
        i_13_873 <= 0;
        i_13_874 <= 0;
        i_13_875 <= 0;
        i_13_876 <= 0;
        i_13_877 <= 0;
        i_13_878 <= 0;
        i_13_879 <= 0;
        i_13_880 <= 0;
        i_13_881 <= 0;
        i_13_882 <= 0;
        i_13_883 <= 0;
        i_13_884 <= 0;
        i_13_885 <= 0;
        i_13_886 <= 0;
        i_13_887 <= 0;
        i_13_888 <= 0;
        i_13_889 <= 0;
        i_13_890 <= 0;
        i_13_891 <= 0;
        i_13_892 <= 0;
        i_13_893 <= 0;
        i_13_894 <= 0;
        i_13_895 <= 0;
        i_13_896 <= 0;
        i_13_897 <= 0;
        i_13_898 <= 0;
        i_13_899 <= 0;
        i_13_900 <= 0;
        i_13_901 <= 0;
        i_13_902 <= 0;
        i_13_903 <= 0;
        i_13_904 <= 0;
        i_13_905 <= 0;
        i_13_906 <= 0;
        i_13_907 <= 0;
        i_13_908 <= 0;
        i_13_909 <= 0;
        i_13_910 <= 0;
        i_13_911 <= 0;
        i_13_912 <= 0;
        i_13_913 <= 0;
        i_13_914 <= 0;
        i_13_915 <= 0;
        i_13_916 <= 0;
        i_13_917 <= 0;
        i_13_918 <= 0;
        i_13_919 <= 0;
        i_13_920 <= 0;
        i_13_921 <= 0;
        i_13_922 <= 0;
        i_13_923 <= 0;
        i_13_924 <= 0;
        i_13_925 <= 0;
        i_13_926 <= 0;
        i_13_927 <= 0;
        i_13_928 <= 0;
        i_13_929 <= 0;
        i_13_930 <= 0;
        i_13_931 <= 0;
        i_13_932 <= 0;
        i_13_933 <= 0;
        i_13_934 <= 0;
        i_13_935 <= 0;
        i_13_936 <= 0;
        i_13_937 <= 0;
        i_13_938 <= 0;
        i_13_939 <= 0;
        i_13_940 <= 0;
        i_13_941 <= 0;
        i_13_942 <= 0;
        i_13_943 <= 0;
        i_13_944 <= 0;
        i_13_945 <= 0;
        i_13_946 <= 0;
        i_13_947 <= 0;
        i_13_948 <= 0;
        i_13_949 <= 0;
        i_13_950 <= 0;
        i_13_951 <= 0;
        i_13_952 <= 0;
        i_13_953 <= 0;
        i_13_954 <= 0;
        i_13_955 <= 0;
        i_13_956 <= 0;
        i_13_957 <= 0;
        i_13_958 <= 0;
        i_13_959 <= 0;
        i_13_960 <= 0;
        i_13_961 <= 0;
        i_13_962 <= 0;
        i_13_963 <= 0;
        i_13_964 <= 0;
        i_13_965 <= 0;
        i_13_966 <= 0;
        i_13_967 <= 0;
        i_13_968 <= 0;
        i_13_969 <= 0;
        i_13_970 <= 0;
        i_13_971 <= 0;
        i_13_972 <= 0;
        i_13_973 <= 0;
        i_13_974 <= 0;
        i_13_975 <= 0;
        i_13_976 <= 0;
        i_13_977 <= 0;
        i_13_978 <= 0;
        i_13_979 <= 0;
        i_13_980 <= 0;
        i_13_981 <= 0;
        i_13_982 <= 0;
        i_13_983 <= 0;
        i_13_984 <= 0;
        i_13_985 <= 0;
        i_13_986 <= 0;
        i_13_987 <= 0;
        i_13_988 <= 0;
        i_13_989 <= 0;
        i_13_990 <= 0;
        i_13_991 <= 0;
        i_13_992 <= 0;
        i_13_993 <= 0;
        i_13_994 <= 0;
        i_13_995 <= 0;
        i_13_996 <= 0;
        i_13_997 <= 0;
        i_13_998 <= 0;
        i_13_999 <= 0;
        i_13_1000 <= 0;
        i_13_1001 <= 0;
        i_13_1002 <= 0;
        i_13_1003 <= 0;
        i_13_1004 <= 0;
        i_13_1005 <= 0;
        i_13_1006 <= 0;
        i_13_1007 <= 0;
        i_13_1008 <= 0;
        i_13_1009 <= 0;
        i_13_1010 <= 0;
        i_13_1011 <= 0;
        i_13_1012 <= 0;
        i_13_1013 <= 0;
        i_13_1014 <= 0;
        i_13_1015 <= 0;
        i_13_1016 <= 0;
        i_13_1017 <= 0;
        i_13_1018 <= 0;
        i_13_1019 <= 0;
        i_13_1020 <= 0;
        i_13_1021 <= 0;
        i_13_1022 <= 0;
        i_13_1023 <= 0;
        i_13_1024 <= 0;
        i_13_1025 <= 0;
        i_13_1026 <= 0;
        i_13_1027 <= 0;
        i_13_1028 <= 0;
        i_13_1029 <= 0;
        i_13_1030 <= 0;
        i_13_1031 <= 0;
        i_13_1032 <= 0;
        i_13_1033 <= 0;
        i_13_1034 <= 0;
        i_13_1035 <= 0;
        i_13_1036 <= 0;
        i_13_1037 <= 0;
        i_13_1038 <= 0;
        i_13_1039 <= 0;
        i_13_1040 <= 0;
        i_13_1041 <= 0;
        i_13_1042 <= 0;
        i_13_1043 <= 0;
        i_13_1044 <= 0;
        i_13_1045 <= 0;
        i_13_1046 <= 0;
        i_13_1047 <= 0;
        i_13_1048 <= 0;
        i_13_1049 <= 0;
        i_13_1050 <= 0;
        i_13_1051 <= 0;
        i_13_1052 <= 0;
        i_13_1053 <= 0;
        i_13_1054 <= 0;
        i_13_1055 <= 0;
        i_13_1056 <= 0;
        i_13_1057 <= 0;
        i_13_1058 <= 0;
        i_13_1059 <= 0;
        i_13_1060 <= 0;
        i_13_1061 <= 0;
        i_13_1062 <= 0;
        i_13_1063 <= 0;
        i_13_1064 <= 0;
        i_13_1065 <= 0;
        i_13_1066 <= 0;
        i_13_1067 <= 0;
        i_13_1068 <= 0;
        i_13_1069 <= 0;
        i_13_1070 <= 0;
        i_13_1071 <= 0;
        i_13_1072 <= 0;
        i_13_1073 <= 0;
        i_13_1074 <= 0;
        i_13_1075 <= 0;
        i_13_1076 <= 0;
        i_13_1077 <= 0;
        i_13_1078 <= 0;
        i_13_1079 <= 0;
        i_13_1080 <= 0;
        i_13_1081 <= 0;
        i_13_1082 <= 0;
        i_13_1083 <= 0;
        i_13_1084 <= 0;
        i_13_1085 <= 0;
        i_13_1086 <= 0;
        i_13_1087 <= 0;
        i_13_1088 <= 0;
        i_13_1089 <= 0;
        i_13_1090 <= 0;
        i_13_1091 <= 0;
        i_13_1092 <= 0;
        i_13_1093 <= 0;
        i_13_1094 <= 0;
        i_13_1095 <= 0;
        i_13_1096 <= 0;
        i_13_1097 <= 0;
        i_13_1098 <= 0;
        i_13_1099 <= 0;
        i_13_1100 <= 0;
        i_13_1101 <= 0;
        i_13_1102 <= 0;
        i_13_1103 <= 0;
        i_13_1104 <= 0;
        i_13_1105 <= 0;
        i_13_1106 <= 0;
        i_13_1107 <= 0;
        i_13_1108 <= 0;
        i_13_1109 <= 0;
        i_13_1110 <= 0;
        i_13_1111 <= 0;
        i_13_1112 <= 0;
        i_13_1113 <= 0;
        i_13_1114 <= 0;
        i_13_1115 <= 0;
        i_13_1116 <= 0;
        i_13_1117 <= 0;
        i_13_1118 <= 0;
        i_13_1119 <= 0;
        i_13_1120 <= 0;
        i_13_1121 <= 0;
        i_13_1122 <= 0;
        i_13_1123 <= 0;
        i_13_1124 <= 0;
        i_13_1125 <= 0;
        i_13_1126 <= 0;
        i_13_1127 <= 0;
        i_13_1128 <= 0;
        i_13_1129 <= 0;
        i_13_1130 <= 0;
        i_13_1131 <= 0;
        i_13_1132 <= 0;
        i_13_1133 <= 0;
        i_13_1134 <= 0;
        i_13_1135 <= 0;
        i_13_1136 <= 0;
        i_13_1137 <= 0;
        i_13_1138 <= 0;
        i_13_1139 <= 0;
        i_13_1140 <= 0;
        i_13_1141 <= 0;
        i_13_1142 <= 0;
        i_13_1143 <= 0;
        i_13_1144 <= 0;
        i_13_1145 <= 0;
        i_13_1146 <= 0;
        i_13_1147 <= 0;
        i_13_1148 <= 0;
        i_13_1149 <= 0;
        i_13_1150 <= 0;
        i_13_1151 <= 0;
        i_13_1152 <= 0;
        i_13_1153 <= 0;
        i_13_1154 <= 0;
        i_13_1155 <= 0;
        i_13_1156 <= 0;
        i_13_1157 <= 0;
        i_13_1158 <= 0;
        i_13_1159 <= 0;
        i_13_1160 <= 0;
        i_13_1161 <= 0;
        i_13_1162 <= 0;
        i_13_1163 <= 0;
        i_13_1164 <= 0;
        i_13_1165 <= 0;
        i_13_1166 <= 0;
        i_13_1167 <= 0;
        i_13_1168 <= 0;
        i_13_1169 <= 0;
        i_13_1170 <= 0;
        i_13_1171 <= 0;
        i_13_1172 <= 0;
        i_13_1173 <= 0;
        i_13_1174 <= 0;
        i_13_1175 <= 0;
        i_13_1176 <= 0;
        i_13_1177 <= 0;
        i_13_1178 <= 0;
        i_13_1179 <= 0;
        i_13_1180 <= 0;
        i_13_1181 <= 0;
        i_13_1182 <= 0;
        i_13_1183 <= 0;
        i_13_1184 <= 0;
        i_13_1185 <= 0;
        i_13_1186 <= 0;
        i_13_1187 <= 0;
        i_13_1188 <= 0;
        i_13_1189 <= 0;
        i_13_1190 <= 0;
        i_13_1191 <= 0;
        i_13_1192 <= 0;
        i_13_1193 <= 0;
        i_13_1194 <= 0;
        i_13_1195 <= 0;
        i_13_1196 <= 0;
        i_13_1197 <= 0;
        i_13_1198 <= 0;
        i_13_1199 <= 0;
        i_13_1200 <= 0;
        i_13_1201 <= 0;
        i_13_1202 <= 0;
        i_13_1203 <= 0;
        i_13_1204 <= 0;
        i_13_1205 <= 0;
        i_13_1206 <= 0;
        i_13_1207 <= 0;
        i_13_1208 <= 0;
        i_13_1209 <= 0;
        i_13_1210 <= 0;
        i_13_1211 <= 0;
        i_13_1212 <= 0;
        i_13_1213 <= 0;
        i_13_1214 <= 0;
        i_13_1215 <= 0;
        i_13_1216 <= 0;
        i_13_1217 <= 0;
        i_13_1218 <= 0;
        i_13_1219 <= 0;
        i_13_1220 <= 0;
        i_13_1221 <= 0;
        i_13_1222 <= 0;
        i_13_1223 <= 0;
        i_13_1224 <= 0;
        i_13_1225 <= 0;
        i_13_1226 <= 0;
        i_13_1227 <= 0;
        i_13_1228 <= 0;
        i_13_1229 <= 0;
        i_13_1230 <= 0;
        i_13_1231 <= 0;
        i_13_1232 <= 0;
        i_13_1233 <= 0;
        i_13_1234 <= 0;
        i_13_1235 <= 0;
        i_13_1236 <= 0;
        i_13_1237 <= 0;
        i_13_1238 <= 0;
        i_13_1239 <= 0;
        i_13_1240 <= 0;
        i_13_1241 <= 0;
        i_13_1242 <= 0;
        i_13_1243 <= 0;
        i_13_1244 <= 0;
        i_13_1245 <= 0;
        i_13_1246 <= 0;
        i_13_1247 <= 0;
        i_13_1248 <= 0;
        i_13_1249 <= 0;
        i_13_1250 <= 0;
        i_13_1251 <= 0;
        i_13_1252 <= 0;
        i_13_1253 <= 0;
        i_13_1254 <= 0;
        i_13_1255 <= 0;
        i_13_1256 <= 0;
        i_13_1257 <= 0;
        i_13_1258 <= 0;
        i_13_1259 <= 0;
        i_13_1260 <= 0;
        i_13_1261 <= 0;
        i_13_1262 <= 0;
        i_13_1263 <= 0;
        i_13_1264 <= 0;
        i_13_1265 <= 0;
        i_13_1266 <= 0;
        i_13_1267 <= 0;
        i_13_1268 <= 0;
        i_13_1269 <= 0;
        i_13_1270 <= 0;
        i_13_1271 <= 0;
        i_13_1272 <= 0;
        i_13_1273 <= 0;
        i_13_1274 <= 0;
        i_13_1275 <= 0;
        i_13_1276 <= 0;
        i_13_1277 <= 0;
        i_13_1278 <= 0;
        i_13_1279 <= 0;
        i_13_1280 <= 0;
        i_13_1281 <= 0;
        i_13_1282 <= 0;
        i_13_1283 <= 0;
        i_13_1284 <= 0;
        i_13_1285 <= 0;
        i_13_1286 <= 0;
        i_13_1287 <= 0;
        i_13_1288 <= 0;
        i_13_1289 <= 0;
        i_13_1290 <= 0;
        i_13_1291 <= 0;
        i_13_1292 <= 0;
        i_13_1293 <= 0;
        i_13_1294 <= 0;
        i_13_1295 <= 0;
        i_13_1296 <= 0;
        i_13_1297 <= 0;
        i_13_1298 <= 0;
        i_13_1299 <= 0;
        i_13_1300 <= 0;
        i_13_1301 <= 0;
        i_13_1302 <= 0;
        i_13_1303 <= 0;
        i_13_1304 <= 0;
        i_13_1305 <= 0;
        i_13_1306 <= 0;
        i_13_1307 <= 0;
        i_13_1308 <= 0;
        i_13_1309 <= 0;
        i_13_1310 <= 0;
        i_13_1311 <= 0;
        i_13_1312 <= 0;
        i_13_1313 <= 0;
        i_13_1314 <= 0;
        i_13_1315 <= 0;
        i_13_1316 <= 0;
        i_13_1317 <= 0;
        i_13_1318 <= 0;
        i_13_1319 <= 0;
        i_13_1320 <= 0;
        i_13_1321 <= 0;
        i_13_1322 <= 0;
        i_13_1323 <= 0;
        i_13_1324 <= 0;
        i_13_1325 <= 0;
        i_13_1326 <= 0;
        i_13_1327 <= 0;
        i_13_1328 <= 0;
        i_13_1329 <= 0;
        i_13_1330 <= 0;
        i_13_1331 <= 0;
        i_13_1332 <= 0;
        i_13_1333 <= 0;
        i_13_1334 <= 0;
        i_13_1335 <= 0;
        i_13_1336 <= 0;
        i_13_1337 <= 0;
        i_13_1338 <= 0;
        i_13_1339 <= 0;
        i_13_1340 <= 0;
        i_13_1341 <= 0;
        i_13_1342 <= 0;
        i_13_1343 <= 0;
        i_13_1344 <= 0;
        i_13_1345 <= 0;
        i_13_1346 <= 0;
        i_13_1347 <= 0;
        i_13_1348 <= 0;
        i_13_1349 <= 0;
        i_13_1350 <= 0;
        i_13_1351 <= 0;
        i_13_1352 <= 0;
        i_13_1353 <= 0;
        i_13_1354 <= 0;
        i_13_1355 <= 0;
        i_13_1356 <= 0;
        i_13_1357 <= 0;
        i_13_1358 <= 0;
        i_13_1359 <= 0;
        i_13_1360 <= 0;
        i_13_1361 <= 0;
        i_13_1362 <= 0;
        i_13_1363 <= 0;
        i_13_1364 <= 0;
        i_13_1365 <= 0;
        i_13_1366 <= 0;
        i_13_1367 <= 0;
        i_13_1368 <= 0;
        i_13_1369 <= 0;
        i_13_1370 <= 0;
        i_13_1371 <= 0;
        i_13_1372 <= 0;
        i_13_1373 <= 0;
        i_13_1374 <= 0;
        i_13_1375 <= 0;
        i_13_1376 <= 0;
        i_13_1377 <= 0;
        i_13_1378 <= 0;
        i_13_1379 <= 0;
        i_13_1380 <= 0;
        i_13_1381 <= 0;
        i_13_1382 <= 0;
        i_13_1383 <= 0;
        i_13_1384 <= 0;
        i_13_1385 <= 0;
        i_13_1386 <= 0;
        i_13_1387 <= 0;
        i_13_1388 <= 0;
        i_13_1389 <= 0;
        i_13_1390 <= 0;
        i_13_1391 <= 0;
        i_13_1392 <= 0;
        i_13_1393 <= 0;
        i_13_1394 <= 0;
        i_13_1395 <= 0;
        i_13_1396 <= 0;
        i_13_1397 <= 0;
        i_13_1398 <= 0;
        i_13_1399 <= 0;
        i_13_1400 <= 0;
        i_13_1401 <= 0;
        i_13_1402 <= 0;
        i_13_1403 <= 0;
        i_13_1404 <= 0;
        i_13_1405 <= 0;
        i_13_1406 <= 0;
        i_13_1407 <= 0;
        i_13_1408 <= 0;
        i_13_1409 <= 0;
        i_13_1410 <= 0;
        i_13_1411 <= 0;
        i_13_1412 <= 0;
        i_13_1413 <= 0;
        i_13_1414 <= 0;
        i_13_1415 <= 0;
        i_13_1416 <= 0;
        i_13_1417 <= 0;
        i_13_1418 <= 0;
        i_13_1419 <= 0;
        i_13_1420 <= 0;
        i_13_1421 <= 0;
        i_13_1422 <= 0;
        i_13_1423 <= 0;
        i_13_1424 <= 0;
        i_13_1425 <= 0;
        i_13_1426 <= 0;
        i_13_1427 <= 0;
        i_13_1428 <= 0;
        i_13_1429 <= 0;
        i_13_1430 <= 0;
        i_13_1431 <= 0;
        i_13_1432 <= 0;
        i_13_1433 <= 0;
        i_13_1434 <= 0;
        i_13_1435 <= 0;
        i_13_1436 <= 0;
        i_13_1437 <= 0;
        i_13_1438 <= 0;
        i_13_1439 <= 0;
        i_13_1440 <= 0;
        i_13_1441 <= 0;
        i_13_1442 <= 0;
        i_13_1443 <= 0;
        i_13_1444 <= 0;
        i_13_1445 <= 0;
        i_13_1446 <= 0;
        i_13_1447 <= 0;
        i_13_1448 <= 0;
        i_13_1449 <= 0;
        i_13_1450 <= 0;
        i_13_1451 <= 0;
        i_13_1452 <= 0;
        i_13_1453 <= 0;
        i_13_1454 <= 0;
        i_13_1455 <= 0;
        i_13_1456 <= 0;
        i_13_1457 <= 0;
        i_13_1458 <= 0;
        i_13_1459 <= 0;
        i_13_1460 <= 0;
        i_13_1461 <= 0;
        i_13_1462 <= 0;
        i_13_1463 <= 0;
        i_13_1464 <= 0;
        i_13_1465 <= 0;
        i_13_1466 <= 0;
        i_13_1467 <= 0;
        i_13_1468 <= 0;
        i_13_1469 <= 0;
        i_13_1470 <= 0;
        i_13_1471 <= 0;
        i_13_1472 <= 0;
        i_13_1473 <= 0;
        i_13_1474 <= 0;
        i_13_1475 <= 0;
        i_13_1476 <= 0;
        i_13_1477 <= 0;
        i_13_1478 <= 0;
        i_13_1479 <= 0;
        i_13_1480 <= 0;
        i_13_1481 <= 0;
        i_13_1482 <= 0;
        i_13_1483 <= 0;
        i_13_1484 <= 0;
        i_13_1485 <= 0;
        i_13_1486 <= 0;
        i_13_1487 <= 0;
        i_13_1488 <= 0;
        i_13_1489 <= 0;
        i_13_1490 <= 0;
        i_13_1491 <= 0;
        i_13_1492 <= 0;
        i_13_1493 <= 0;
        i_13_1494 <= 0;
        i_13_1495 <= 0;
        i_13_1496 <= 0;
        i_13_1497 <= 0;
        i_13_1498 <= 0;
        i_13_1499 <= 0;
        i_13_1500 <= 0;
        i_13_1501 <= 0;
        i_13_1502 <= 0;
        i_13_1503 <= 0;
        i_13_1504 <= 0;
        i_13_1505 <= 0;
        i_13_1506 <= 0;
        i_13_1507 <= 0;
        i_13_1508 <= 0;
        i_13_1509 <= 0;
        i_13_1510 <= 0;
        i_13_1511 <= 0;
        i_13_1512 <= 0;
        i_13_1513 <= 0;
        i_13_1514 <= 0;
        i_13_1515 <= 0;
        i_13_1516 <= 0;
        i_13_1517 <= 0;
        i_13_1518 <= 0;
        i_13_1519 <= 0;
        i_13_1520 <= 0;
        i_13_1521 <= 0;
        i_13_1522 <= 0;
        i_13_1523 <= 0;
        i_13_1524 <= 0;
        i_13_1525 <= 0;
        i_13_1526 <= 0;
        i_13_1527 <= 0;
        i_13_1528 <= 0;
        i_13_1529 <= 0;
        i_13_1530 <= 0;
        i_13_1531 <= 0;
        i_13_1532 <= 0;
        i_13_1533 <= 0;
        i_13_1534 <= 0;
        i_13_1535 <= 0;
        i_13_1536 <= 0;
        i_13_1537 <= 0;
        i_13_1538 <= 0;
        i_13_1539 <= 0;
        i_13_1540 <= 0;
        i_13_1541 <= 0;
        i_13_1542 <= 0;
        i_13_1543 <= 0;
        i_13_1544 <= 0;
        i_13_1545 <= 0;
        i_13_1546 <= 0;
        i_13_1547 <= 0;
        i_13_1548 <= 0;
        i_13_1549 <= 0;
        i_13_1550 <= 0;
        i_13_1551 <= 0;
        i_13_1552 <= 0;
        i_13_1553 <= 0;
        i_13_1554 <= 0;
        i_13_1555 <= 0;
        i_13_1556 <= 0;
        i_13_1557 <= 0;
        i_13_1558 <= 0;
        i_13_1559 <= 0;
        i_13_1560 <= 0;
        i_13_1561 <= 0;
        i_13_1562 <= 0;
        i_13_1563 <= 0;
        i_13_1564 <= 0;
        i_13_1565 <= 0;
        i_13_1566 <= 0;
        i_13_1567 <= 0;
        i_13_1568 <= 0;
        i_13_1569 <= 0;
        i_13_1570 <= 0;
        i_13_1571 <= 0;
        i_13_1572 <= 0;
        i_13_1573 <= 0;
        i_13_1574 <= 0;
        i_13_1575 <= 0;
        i_13_1576 <= 0;
        i_13_1577 <= 0;
        i_13_1578 <= 0;
        i_13_1579 <= 0;
        i_13_1580 <= 0;
        i_13_1581 <= 0;
        i_13_1582 <= 0;
        i_13_1583 <= 0;
        i_13_1584 <= 0;
        i_13_1585 <= 0;
        i_13_1586 <= 0;
        i_13_1587 <= 0;
        i_13_1588 <= 0;
        i_13_1589 <= 0;
        i_13_1590 <= 0;
        i_13_1591 <= 0;
        i_13_1592 <= 0;
        i_13_1593 <= 0;
        i_13_1594 <= 0;
        i_13_1595 <= 0;
        i_13_1596 <= 0;
        i_13_1597 <= 0;
        i_13_1598 <= 0;
        i_13_1599 <= 0;
        i_13_1600 <= 0;
        i_13_1601 <= 0;
        i_13_1602 <= 0;
        i_13_1603 <= 0;
        i_13_1604 <= 0;
        i_13_1605 <= 0;
        i_13_1606 <= 0;
        i_13_1607 <= 0;
        i_13_1608 <= 0;
        i_13_1609 <= 0;
        i_13_1610 <= 0;
        i_13_1611 <= 0;
        i_13_1612 <= 0;
        i_13_1613 <= 0;
        i_13_1614 <= 0;
        i_13_1615 <= 0;
        i_13_1616 <= 0;
        i_13_1617 <= 0;
        i_13_1618 <= 0;
        i_13_1619 <= 0;
        i_13_1620 <= 0;
        i_13_1621 <= 0;
        i_13_1622 <= 0;
        i_13_1623 <= 0;
        i_13_1624 <= 0;
        i_13_1625 <= 0;
        i_13_1626 <= 0;
        i_13_1627 <= 0;
        i_13_1628 <= 0;
        i_13_1629 <= 0;
        i_13_1630 <= 0;
        i_13_1631 <= 0;
        i_13_1632 <= 0;
        i_13_1633 <= 0;
        i_13_1634 <= 0;
        i_13_1635 <= 0;
        i_13_1636 <= 0;
        i_13_1637 <= 0;
        i_13_1638 <= 0;
        i_13_1639 <= 0;
        i_13_1640 <= 0;
        i_13_1641 <= 0;
        i_13_1642 <= 0;
        i_13_1643 <= 0;
        i_13_1644 <= 0;
        i_13_1645 <= 0;
        i_13_1646 <= 0;
        i_13_1647 <= 0;
        i_13_1648 <= 0;
        i_13_1649 <= 0;
        i_13_1650 <= 0;
        i_13_1651 <= 0;
        i_13_1652 <= 0;
        i_13_1653 <= 0;
        i_13_1654 <= 0;
        i_13_1655 <= 0;
        i_13_1656 <= 0;
        i_13_1657 <= 0;
        i_13_1658 <= 0;
        i_13_1659 <= 0;
        i_13_1660 <= 0;
        i_13_1661 <= 0;
        i_13_1662 <= 0;
        i_13_1663 <= 0;
        i_13_1664 <= 0;
        i_13_1665 <= 0;
        i_13_1666 <= 0;
        i_13_1667 <= 0;
        i_13_1668 <= 0;
        i_13_1669 <= 0;
        i_13_1670 <= 0;
        i_13_1671 <= 0;
        i_13_1672 <= 0;
        i_13_1673 <= 0;
        i_13_1674 <= 0;
        i_13_1675 <= 0;
        i_13_1676 <= 0;
        i_13_1677 <= 0;
        i_13_1678 <= 0;
        i_13_1679 <= 0;
        i_13_1680 <= 0;
        i_13_1681 <= 0;
        i_13_1682 <= 0;
        i_13_1683 <= 0;
        i_13_1684 <= 0;
        i_13_1685 <= 0;
        i_13_1686 <= 0;
        i_13_1687 <= 0;
        i_13_1688 <= 0;
        i_13_1689 <= 0;
        i_13_1690 <= 0;
        i_13_1691 <= 0;
        i_13_1692 <= 0;
        i_13_1693 <= 0;
        i_13_1694 <= 0;
        i_13_1695 <= 0;
        i_13_1696 <= 0;
        i_13_1697 <= 0;
        i_13_1698 <= 0;
        i_13_1699 <= 0;
        i_13_1700 <= 0;
        i_13_1701 <= 0;
        i_13_1702 <= 0;
        i_13_1703 <= 0;
        i_13_1704 <= 0;
        i_13_1705 <= 0;
        i_13_1706 <= 0;
        i_13_1707 <= 0;
        i_13_1708 <= 0;
        i_13_1709 <= 0;
        i_13_1710 <= 0;
        i_13_1711 <= 0;
        i_13_1712 <= 0;
        i_13_1713 <= 0;
        i_13_1714 <= 0;
        i_13_1715 <= 0;
        i_13_1716 <= 0;
        i_13_1717 <= 0;
        i_13_1718 <= 0;
        i_13_1719 <= 0;
        i_13_1720 <= 0;
        i_13_1721 <= 0;
        i_13_1722 <= 0;
        i_13_1723 <= 0;
        i_13_1724 <= 0;
        i_13_1725 <= 0;
        i_13_1726 <= 0;
        i_13_1727 <= 0;
        i_13_1728 <= 0;
        i_13_1729 <= 0;
        i_13_1730 <= 0;
        i_13_1731 <= 0;
        i_13_1732 <= 0;
        i_13_1733 <= 0;
        i_13_1734 <= 0;
        i_13_1735 <= 0;
        i_13_1736 <= 0;
        i_13_1737 <= 0;
        i_13_1738 <= 0;
        i_13_1739 <= 0;
        i_13_1740 <= 0;
        i_13_1741 <= 0;
        i_13_1742 <= 0;
        i_13_1743 <= 0;
        i_13_1744 <= 0;
        i_13_1745 <= 0;
        i_13_1746 <= 0;
        i_13_1747 <= 0;
        i_13_1748 <= 0;
        i_13_1749 <= 0;
        i_13_1750 <= 0;
        i_13_1751 <= 0;
        i_13_1752 <= 0;
        i_13_1753 <= 0;
        i_13_1754 <= 0;
        i_13_1755 <= 0;
        i_13_1756 <= 0;
        i_13_1757 <= 0;
        i_13_1758 <= 0;
        i_13_1759 <= 0;
        i_13_1760 <= 0;
        i_13_1761 <= 0;
        i_13_1762 <= 0;
        i_13_1763 <= 0;
        i_13_1764 <= 0;
        i_13_1765 <= 0;
        i_13_1766 <= 0;
        i_13_1767 <= 0;
        i_13_1768 <= 0;
        i_13_1769 <= 0;
        i_13_1770 <= 0;
        i_13_1771 <= 0;
        i_13_1772 <= 0;
        i_13_1773 <= 0;
        i_13_1774 <= 0;
        i_13_1775 <= 0;
        i_13_1776 <= 0;
        i_13_1777 <= 0;
        i_13_1778 <= 0;
        i_13_1779 <= 0;
        i_13_1780 <= 0;
        i_13_1781 <= 0;
        i_13_1782 <= 0;
        i_13_1783 <= 0;
        i_13_1784 <= 0;
        i_13_1785 <= 0;
        i_13_1786 <= 0;
        i_13_1787 <= 0;
        i_13_1788 <= 0;
        i_13_1789 <= 0;
        i_13_1790 <= 0;
        i_13_1791 <= 0;
        i_13_1792 <= 0;
        i_13_1793 <= 0;
        i_13_1794 <= 0;
        i_13_1795 <= 0;
        i_13_1796 <= 0;
        i_13_1797 <= 0;
        i_13_1798 <= 0;
        i_13_1799 <= 0;
        i_13_1800 <= 0;
        i_13_1801 <= 0;
        i_13_1802 <= 0;
        i_13_1803 <= 0;
        i_13_1804 <= 0;
        i_13_1805 <= 0;
        i_13_1806 <= 0;
        i_13_1807 <= 0;
        i_13_1808 <= 0;
        i_13_1809 <= 0;
        i_13_1810 <= 0;
        i_13_1811 <= 0;
        i_13_1812 <= 0;
        i_13_1813 <= 0;
        i_13_1814 <= 0;
        i_13_1815 <= 0;
        i_13_1816 <= 0;
        i_13_1817 <= 0;
        i_13_1818 <= 0;
        i_13_1819 <= 0;
        i_13_1820 <= 0;
        i_13_1821 <= 0;
        i_13_1822 <= 0;
        i_13_1823 <= 0;
        i_13_1824 <= 0;
        i_13_1825 <= 0;
        i_13_1826 <= 0;
        i_13_1827 <= 0;
        i_13_1828 <= 0;
        i_13_1829 <= 0;
        i_13_1830 <= 0;
        i_13_1831 <= 0;
        i_13_1832 <= 0;
        i_13_1833 <= 0;
        i_13_1834 <= 0;
        i_13_1835 <= 0;
        i_13_1836 <= 0;
        i_13_1837 <= 0;
        i_13_1838 <= 0;
        i_13_1839 <= 0;
        i_13_1840 <= 0;
        i_13_1841 <= 0;
        i_13_1842 <= 0;
        i_13_1843 <= 0;
        i_13_1844 <= 0;
        i_13_1845 <= 0;
        i_13_1846 <= 0;
        i_13_1847 <= 0;
        i_13_1848 <= 0;
        i_13_1849 <= 0;
        i_13_1850 <= 0;
        i_13_1851 <= 0;
        i_13_1852 <= 0;
        i_13_1853 <= 0;
        i_13_1854 <= 0;
        i_13_1855 <= 0;
        i_13_1856 <= 0;
        i_13_1857 <= 0;
        i_13_1858 <= 0;
        i_13_1859 <= 0;
        i_13_1860 <= 0;
        i_13_1861 <= 0;
        i_13_1862 <= 0;
        i_13_1863 <= 0;
        i_13_1864 <= 0;
        i_13_1865 <= 0;
        i_13_1866 <= 0;
        i_13_1867 <= 0;
        i_13_1868 <= 0;
        i_13_1869 <= 0;
        i_13_1870 <= 0;
        i_13_1871 <= 0;
        i_13_1872 <= 0;
        i_13_1873 <= 0;
        i_13_1874 <= 0;
        i_13_1875 <= 0;
        i_13_1876 <= 0;
        i_13_1877 <= 0;
        i_13_1878 <= 0;
        i_13_1879 <= 0;
        i_13_1880 <= 0;
        i_13_1881 <= 0;
        i_13_1882 <= 0;
        i_13_1883 <= 0;
        i_13_1884 <= 0;
        i_13_1885 <= 0;
        i_13_1886 <= 0;
        i_13_1887 <= 0;
        i_13_1888 <= 0;
        i_13_1889 <= 0;
        i_13_1890 <= 0;
        i_13_1891 <= 0;
        i_13_1892 <= 0;
        i_13_1893 <= 0;
        i_13_1894 <= 0;
        i_13_1895 <= 0;
        i_13_1896 <= 0;
        i_13_1897 <= 0;
        i_13_1898 <= 0;
        i_13_1899 <= 0;
        i_13_1900 <= 0;
        i_13_1901 <= 0;
        i_13_1902 <= 0;
        i_13_1903 <= 0;
        i_13_1904 <= 0;
        i_13_1905 <= 0;
        i_13_1906 <= 0;
        i_13_1907 <= 0;
        i_13_1908 <= 0;
        i_13_1909 <= 0;
        i_13_1910 <= 0;
        i_13_1911 <= 0;
        i_13_1912 <= 0;
        i_13_1913 <= 0;
        i_13_1914 <= 0;
        i_13_1915 <= 0;
        i_13_1916 <= 0;
        i_13_1917 <= 0;
        i_13_1918 <= 0;
        i_13_1919 <= 0;
        i_13_1920 <= 0;
        i_13_1921 <= 0;
        i_13_1922 <= 0;
        i_13_1923 <= 0;
        i_13_1924 <= 0;
        i_13_1925 <= 0;
        i_13_1926 <= 0;
        i_13_1927 <= 0;
        i_13_1928 <= 0;
        i_13_1929 <= 0;
        i_13_1930 <= 0;
        i_13_1931 <= 0;
        i_13_1932 <= 0;
        i_13_1933 <= 0;
        i_13_1934 <= 0;
        i_13_1935 <= 0;
        i_13_1936 <= 0;
        i_13_1937 <= 0;
        i_13_1938 <= 0;
        i_13_1939 <= 0;
        i_13_1940 <= 0;
        i_13_1941 <= 0;
        i_13_1942 <= 0;
        i_13_1943 <= 0;
        i_13_1944 <= 0;
        i_13_1945 <= 0;
        i_13_1946 <= 0;
        i_13_1947 <= 0;
        i_13_1948 <= 0;
        i_13_1949 <= 0;
        i_13_1950 <= 0;
        i_13_1951 <= 0;
        i_13_1952 <= 0;
        i_13_1953 <= 0;
        i_13_1954 <= 0;
        i_13_1955 <= 0;
        i_13_1956 <= 0;
        i_13_1957 <= 0;
        i_13_1958 <= 0;
        i_13_1959 <= 0;
        i_13_1960 <= 0;
        i_13_1961 <= 0;
        i_13_1962 <= 0;
        i_13_1963 <= 0;
        i_13_1964 <= 0;
        i_13_1965 <= 0;
        i_13_1966 <= 0;
        i_13_1967 <= 0;
        i_13_1968 <= 0;
        i_13_1969 <= 0;
        i_13_1970 <= 0;
        i_13_1971 <= 0;
        i_13_1972 <= 0;
        i_13_1973 <= 0;
        i_13_1974 <= 0;
        i_13_1975 <= 0;
        i_13_1976 <= 0;
        i_13_1977 <= 0;
        i_13_1978 <= 0;
        i_13_1979 <= 0;
        i_13_1980 <= 0;
        i_13_1981 <= 0;
        i_13_1982 <= 0;
        i_13_1983 <= 0;
        i_13_1984 <= 0;
        i_13_1985 <= 0;
        i_13_1986 <= 0;
        i_13_1987 <= 0;
        i_13_1988 <= 0;
        i_13_1989 <= 0;
        i_13_1990 <= 0;
        i_13_1991 <= 0;
        i_13_1992 <= 0;
        i_13_1993 <= 0;
        i_13_1994 <= 0;
        i_13_1995 <= 0;
        i_13_1996 <= 0;
        i_13_1997 <= 0;
        i_13_1998 <= 0;
        i_13_1999 <= 0;
        i_13_2000 <= 0;
        i_13_2001 <= 0;
        i_13_2002 <= 0;
        i_13_2003 <= 0;
        i_13_2004 <= 0;
        i_13_2005 <= 0;
        i_13_2006 <= 0;
        i_13_2007 <= 0;
        i_13_2008 <= 0;
        i_13_2009 <= 0;
        i_13_2010 <= 0;
        i_13_2011 <= 0;
        i_13_2012 <= 0;
        i_13_2013 <= 0;
        i_13_2014 <= 0;
        i_13_2015 <= 0;
        i_13_2016 <= 0;
        i_13_2017 <= 0;
        i_13_2018 <= 0;
        i_13_2019 <= 0;
        i_13_2020 <= 0;
        i_13_2021 <= 0;
        i_13_2022 <= 0;
        i_13_2023 <= 0;
        i_13_2024 <= 0;
        i_13_2025 <= 0;
        i_13_2026 <= 0;
        i_13_2027 <= 0;
        i_13_2028 <= 0;
        i_13_2029 <= 0;
        i_13_2030 <= 0;
        i_13_2031 <= 0;
        i_13_2032 <= 0;
        i_13_2033 <= 0;
        i_13_2034 <= 0;
        i_13_2035 <= 0;
        i_13_2036 <= 0;
        i_13_2037 <= 0;
        i_13_2038 <= 0;
        i_13_2039 <= 0;
        i_13_2040 <= 0;
        i_13_2041 <= 0;
        i_13_2042 <= 0;
        i_13_2043 <= 0;
        i_13_2044 <= 0;
        i_13_2045 <= 0;
        i_13_2046 <= 0;
        i_13_2047 <= 0;
        i_13_2048 <= 0;
        i_13_2049 <= 0;
        i_13_2050 <= 0;
        i_13_2051 <= 0;
        i_13_2052 <= 0;
        i_13_2053 <= 0;
        i_13_2054 <= 0;
        i_13_2055 <= 0;
        i_13_2056 <= 0;
        i_13_2057 <= 0;
        i_13_2058 <= 0;
        i_13_2059 <= 0;
        i_13_2060 <= 0;
        i_13_2061 <= 0;
        i_13_2062 <= 0;
        i_13_2063 <= 0;
        i_13_2064 <= 0;
        i_13_2065 <= 0;
        i_13_2066 <= 0;
        i_13_2067 <= 0;
        i_13_2068 <= 0;
        i_13_2069 <= 0;
        i_13_2070 <= 0;
        i_13_2071 <= 0;
        i_13_2072 <= 0;
        i_13_2073 <= 0;
        i_13_2074 <= 0;
        i_13_2075 <= 0;
        i_13_2076 <= 0;
        i_13_2077 <= 0;
        i_13_2078 <= 0;
        i_13_2079 <= 0;
        i_13_2080 <= 0;
        i_13_2081 <= 0;
        i_13_2082 <= 0;
        i_13_2083 <= 0;
        i_13_2084 <= 0;
        i_13_2085 <= 0;
        i_13_2086 <= 0;
        i_13_2087 <= 0;
        i_13_2088 <= 0;
        i_13_2089 <= 0;
        i_13_2090 <= 0;
        i_13_2091 <= 0;
        i_13_2092 <= 0;
        i_13_2093 <= 0;
        i_13_2094 <= 0;
        i_13_2095 <= 0;
        i_13_2096 <= 0;
        i_13_2097 <= 0;
        i_13_2098 <= 0;
        i_13_2099 <= 0;
        i_13_2100 <= 0;
        i_13_2101 <= 0;
        i_13_2102 <= 0;
        i_13_2103 <= 0;
        i_13_2104 <= 0;
        i_13_2105 <= 0;
        i_13_2106 <= 0;
        i_13_2107 <= 0;
        i_13_2108 <= 0;
        i_13_2109 <= 0;
        i_13_2110 <= 0;
        i_13_2111 <= 0;
        i_13_2112 <= 0;
        i_13_2113 <= 0;
        i_13_2114 <= 0;
        i_13_2115 <= 0;
        i_13_2116 <= 0;
        i_13_2117 <= 0;
        i_13_2118 <= 0;
        i_13_2119 <= 0;
        i_13_2120 <= 0;
        i_13_2121 <= 0;
        i_13_2122 <= 0;
        i_13_2123 <= 0;
        i_13_2124 <= 0;
        i_13_2125 <= 0;
        i_13_2126 <= 0;
        i_13_2127 <= 0;
        i_13_2128 <= 0;
        i_13_2129 <= 0;
        i_13_2130 <= 0;
        i_13_2131 <= 0;
        i_13_2132 <= 0;
        i_13_2133 <= 0;
        i_13_2134 <= 0;
        i_13_2135 <= 0;
        i_13_2136 <= 0;
        i_13_2137 <= 0;
        i_13_2138 <= 0;
        i_13_2139 <= 0;
        i_13_2140 <= 0;
        i_13_2141 <= 0;
        i_13_2142 <= 0;
        i_13_2143 <= 0;
        i_13_2144 <= 0;
        i_13_2145 <= 0;
        i_13_2146 <= 0;
        i_13_2147 <= 0;
        i_13_2148 <= 0;
        i_13_2149 <= 0;
        i_13_2150 <= 0;
        i_13_2151 <= 0;
        i_13_2152 <= 0;
        i_13_2153 <= 0;
        i_13_2154 <= 0;
        i_13_2155 <= 0;
        i_13_2156 <= 0;
        i_13_2157 <= 0;
        i_13_2158 <= 0;
        i_13_2159 <= 0;
        i_13_2160 <= 0;
        i_13_2161 <= 0;
        i_13_2162 <= 0;
        i_13_2163 <= 0;
        i_13_2164 <= 0;
        i_13_2165 <= 0;
        i_13_2166 <= 0;
        i_13_2167 <= 0;
        i_13_2168 <= 0;
        i_13_2169 <= 0;
        i_13_2170 <= 0;
        i_13_2171 <= 0;
        i_13_2172 <= 0;
        i_13_2173 <= 0;
        i_13_2174 <= 0;
        i_13_2175 <= 0;
        i_13_2176 <= 0;
        i_13_2177 <= 0;
        i_13_2178 <= 0;
        i_13_2179 <= 0;
        i_13_2180 <= 0;
        i_13_2181 <= 0;
        i_13_2182 <= 0;
        i_13_2183 <= 0;
        i_13_2184 <= 0;
        i_13_2185 <= 0;
        i_13_2186 <= 0;
        i_13_2187 <= 0;
        i_13_2188 <= 0;
        i_13_2189 <= 0;
        i_13_2190 <= 0;
        i_13_2191 <= 0;
        i_13_2192 <= 0;
        i_13_2193 <= 0;
        i_13_2194 <= 0;
        i_13_2195 <= 0;
        i_13_2196 <= 0;
        i_13_2197 <= 0;
        i_13_2198 <= 0;
        i_13_2199 <= 0;
        i_13_2200 <= 0;
        i_13_2201 <= 0;
        i_13_2202 <= 0;
        i_13_2203 <= 0;
        i_13_2204 <= 0;
        i_13_2205 <= 0;
        i_13_2206 <= 0;
        i_13_2207 <= 0;
        i_13_2208 <= 0;
        i_13_2209 <= 0;
        i_13_2210 <= 0;
        i_13_2211 <= 0;
        i_13_2212 <= 0;
        i_13_2213 <= 0;
        i_13_2214 <= 0;
        i_13_2215 <= 0;
        i_13_2216 <= 0;
        i_13_2217 <= 0;
        i_13_2218 <= 0;
        i_13_2219 <= 0;
        i_13_2220 <= 0;
        i_13_2221 <= 0;
        i_13_2222 <= 0;
        i_13_2223 <= 0;
        i_13_2224 <= 0;
        i_13_2225 <= 0;
        i_13_2226 <= 0;
        i_13_2227 <= 0;
        i_13_2228 <= 0;
        i_13_2229 <= 0;
        i_13_2230 <= 0;
        i_13_2231 <= 0;
        i_13_2232 <= 0;
        i_13_2233 <= 0;
        i_13_2234 <= 0;
        i_13_2235 <= 0;
        i_13_2236 <= 0;
        i_13_2237 <= 0;
        i_13_2238 <= 0;
        i_13_2239 <= 0;
        i_13_2240 <= 0;
        i_13_2241 <= 0;
        i_13_2242 <= 0;
        i_13_2243 <= 0;
        i_13_2244 <= 0;
        i_13_2245 <= 0;
        i_13_2246 <= 0;
        i_13_2247 <= 0;
        i_13_2248 <= 0;
        i_13_2249 <= 0;
        i_13_2250 <= 0;
        i_13_2251 <= 0;
        i_13_2252 <= 0;
        i_13_2253 <= 0;
        i_13_2254 <= 0;
        i_13_2255 <= 0;
        i_13_2256 <= 0;
        i_13_2257 <= 0;
        i_13_2258 <= 0;
        i_13_2259 <= 0;
        i_13_2260 <= 0;
        i_13_2261 <= 0;
        i_13_2262 <= 0;
        i_13_2263 <= 0;
        i_13_2264 <= 0;
        i_13_2265 <= 0;
        i_13_2266 <= 0;
        i_13_2267 <= 0;
        i_13_2268 <= 0;
        i_13_2269 <= 0;
        i_13_2270 <= 0;
        i_13_2271 <= 0;
        i_13_2272 <= 0;
        i_13_2273 <= 0;
        i_13_2274 <= 0;
        i_13_2275 <= 0;
        i_13_2276 <= 0;
        i_13_2277 <= 0;
        i_13_2278 <= 0;
        i_13_2279 <= 0;
        i_13_2280 <= 0;
        i_13_2281 <= 0;
        i_13_2282 <= 0;
        i_13_2283 <= 0;
        i_13_2284 <= 0;
        i_13_2285 <= 0;
        i_13_2286 <= 0;
        i_13_2287 <= 0;
        i_13_2288 <= 0;
        i_13_2289 <= 0;
        i_13_2290 <= 0;
        i_13_2291 <= 0;
        i_13_2292 <= 0;
        i_13_2293 <= 0;
        i_13_2294 <= 0;
        i_13_2295 <= 0;
        i_13_2296 <= 0;
        i_13_2297 <= 0;
        i_13_2298 <= 0;
        i_13_2299 <= 0;
        i_13_2300 <= 0;
        i_13_2301 <= 0;
        i_13_2302 <= 0;
        i_13_2303 <= 0;
        i_13_2304 <= 0;
        i_13_2305 <= 0;
        i_13_2306 <= 0;
        i_13_2307 <= 0;
        i_13_2308 <= 0;
        i_13_2309 <= 0;
        i_13_2310 <= 0;
        i_13_2311 <= 0;
        i_13_2312 <= 0;
        i_13_2313 <= 0;
        i_13_2314 <= 0;
        i_13_2315 <= 0;
        i_13_2316 <= 0;
        i_13_2317 <= 0;
        i_13_2318 <= 0;
        i_13_2319 <= 0;
        i_13_2320 <= 0;
        i_13_2321 <= 0;
        i_13_2322 <= 0;
        i_13_2323 <= 0;
        i_13_2324 <= 0;
        i_13_2325 <= 0;
        i_13_2326 <= 0;
        i_13_2327 <= 0;
        i_13_2328 <= 0;
        i_13_2329 <= 0;
        i_13_2330 <= 0;
        i_13_2331 <= 0;
        i_13_2332 <= 0;
        i_13_2333 <= 0;
        i_13_2334 <= 0;
        i_13_2335 <= 0;
        i_13_2336 <= 0;
        i_13_2337 <= 0;
        i_13_2338 <= 0;
        i_13_2339 <= 0;
        i_13_2340 <= 0;
        i_13_2341 <= 0;
        i_13_2342 <= 0;
        i_13_2343 <= 0;
        i_13_2344 <= 0;
        i_13_2345 <= 0;
        i_13_2346 <= 0;
        i_13_2347 <= 0;
        i_13_2348 <= 0;
        i_13_2349 <= 0;
        i_13_2350 <= 0;
        i_13_2351 <= 0;
        i_13_2352 <= 0;
        i_13_2353 <= 0;
        i_13_2354 <= 0;
        i_13_2355 <= 0;
        i_13_2356 <= 0;
        i_13_2357 <= 0;
        i_13_2358 <= 0;
        i_13_2359 <= 0;
        i_13_2360 <= 0;
        i_13_2361 <= 0;
        i_13_2362 <= 0;
        i_13_2363 <= 0;
        i_13_2364 <= 0;
        i_13_2365 <= 0;
        i_13_2366 <= 0;
        i_13_2367 <= 0;
        i_13_2368 <= 0;
        i_13_2369 <= 0;
        i_13_2370 <= 0;
        i_13_2371 <= 0;
        i_13_2372 <= 0;
        i_13_2373 <= 0;
        i_13_2374 <= 0;
        i_13_2375 <= 0;
        i_13_2376 <= 0;
        i_13_2377 <= 0;
        i_13_2378 <= 0;
        i_13_2379 <= 0;
        i_13_2380 <= 0;
        i_13_2381 <= 0;
        i_13_2382 <= 0;
        i_13_2383 <= 0;
        i_13_2384 <= 0;
        i_13_2385 <= 0;
        i_13_2386 <= 0;
        i_13_2387 <= 0;
        i_13_2388 <= 0;
        i_13_2389 <= 0;
        i_13_2390 <= 0;
        i_13_2391 <= 0;
        i_13_2392 <= 0;
        i_13_2393 <= 0;
        i_13_2394 <= 0;
        i_13_2395 <= 0;
        i_13_2396 <= 0;
        i_13_2397 <= 0;
        i_13_2398 <= 0;
        i_13_2399 <= 0;
        i_13_2400 <= 0;
        i_13_2401 <= 0;
        i_13_2402 <= 0;
        i_13_2403 <= 0;
        i_13_2404 <= 0;
        i_13_2405 <= 0;
        i_13_2406 <= 0;
        i_13_2407 <= 0;
        i_13_2408 <= 0;
        i_13_2409 <= 0;
        i_13_2410 <= 0;
        i_13_2411 <= 0;
        i_13_2412 <= 0;
        i_13_2413 <= 0;
        i_13_2414 <= 0;
        i_13_2415 <= 0;
        i_13_2416 <= 0;
        i_13_2417 <= 0;
        i_13_2418 <= 0;
        i_13_2419 <= 0;
        i_13_2420 <= 0;
        i_13_2421 <= 0;
        i_13_2422 <= 0;
        i_13_2423 <= 0;
        i_13_2424 <= 0;
        i_13_2425 <= 0;
        i_13_2426 <= 0;
        i_13_2427 <= 0;
        i_13_2428 <= 0;
        i_13_2429 <= 0;
        i_13_2430 <= 0;
        i_13_2431 <= 0;
        i_13_2432 <= 0;
        i_13_2433 <= 0;
        i_13_2434 <= 0;
        i_13_2435 <= 0;
        i_13_2436 <= 0;
        i_13_2437 <= 0;
        i_13_2438 <= 0;
        i_13_2439 <= 0;
        i_13_2440 <= 0;
        i_13_2441 <= 0;
        i_13_2442 <= 0;
        i_13_2443 <= 0;
        i_13_2444 <= 0;
        i_13_2445 <= 0;
        i_13_2446 <= 0;
        i_13_2447 <= 0;
        i_13_2448 <= 0;
        i_13_2449 <= 0;
        i_13_2450 <= 0;
        i_13_2451 <= 0;
        i_13_2452 <= 0;
        i_13_2453 <= 0;
        i_13_2454 <= 0;
        i_13_2455 <= 0;
        i_13_2456 <= 0;
        i_13_2457 <= 0;
        i_13_2458 <= 0;
        i_13_2459 <= 0;
        i_13_2460 <= 0;
        i_13_2461 <= 0;
        i_13_2462 <= 0;
        i_13_2463 <= 0;
        i_13_2464 <= 0;
        i_13_2465 <= 0;
        i_13_2466 <= 0;
        i_13_2467 <= 0;
        i_13_2468 <= 0;
        i_13_2469 <= 0;
        i_13_2470 <= 0;
        i_13_2471 <= 0;
        i_13_2472 <= 0;
        i_13_2473 <= 0;
        i_13_2474 <= 0;
        i_13_2475 <= 0;
        i_13_2476 <= 0;
        i_13_2477 <= 0;
        i_13_2478 <= 0;
        i_13_2479 <= 0;
        i_13_2480 <= 0;
        i_13_2481 <= 0;
        i_13_2482 <= 0;
        i_13_2483 <= 0;
        i_13_2484 <= 0;
        i_13_2485 <= 0;
        i_13_2486 <= 0;
        i_13_2487 <= 0;
        i_13_2488 <= 0;
        i_13_2489 <= 0;
        i_13_2490 <= 0;
        i_13_2491 <= 0;
        i_13_2492 <= 0;
        i_13_2493 <= 0;
        i_13_2494 <= 0;
        i_13_2495 <= 0;
        i_13_2496 <= 0;
        i_13_2497 <= 0;
        i_13_2498 <= 0;
        i_13_2499 <= 0;
        i_13_2500 <= 0;
        i_13_2501 <= 0;
        i_13_2502 <= 0;
        i_13_2503 <= 0;
        i_13_2504 <= 0;
        i_13_2505 <= 0;
        i_13_2506 <= 0;
        i_13_2507 <= 0;
        i_13_2508 <= 0;
        i_13_2509 <= 0;
        i_13_2510 <= 0;
        i_13_2511 <= 0;
        i_13_2512 <= 0;
        i_13_2513 <= 0;
        i_13_2514 <= 0;
        i_13_2515 <= 0;
        i_13_2516 <= 0;
        i_13_2517 <= 0;
        i_13_2518 <= 0;
        i_13_2519 <= 0;
        i_13_2520 <= 0;
        i_13_2521 <= 0;
        i_13_2522 <= 0;
        i_13_2523 <= 0;
        i_13_2524 <= 0;
        i_13_2525 <= 0;
        i_13_2526 <= 0;
        i_13_2527 <= 0;
        i_13_2528 <= 0;
        i_13_2529 <= 0;
        i_13_2530 <= 0;
        i_13_2531 <= 0;
        i_13_2532 <= 0;
        i_13_2533 <= 0;
        i_13_2534 <= 0;
        i_13_2535 <= 0;
        i_13_2536 <= 0;
        i_13_2537 <= 0;
        i_13_2538 <= 0;
        i_13_2539 <= 0;
        i_13_2540 <= 0;
        i_13_2541 <= 0;
        i_13_2542 <= 0;
        i_13_2543 <= 0;
        i_13_2544 <= 0;
        i_13_2545 <= 0;
        i_13_2546 <= 0;
        i_13_2547 <= 0;
        i_13_2548 <= 0;
        i_13_2549 <= 0;
        i_13_2550 <= 0;
        i_13_2551 <= 0;
        i_13_2552 <= 0;
        i_13_2553 <= 0;
        i_13_2554 <= 0;
        i_13_2555 <= 0;
        i_13_2556 <= 0;
        i_13_2557 <= 0;
        i_13_2558 <= 0;
        i_13_2559 <= 0;
        i_13_2560 <= 0;
        i_13_2561 <= 0;
        i_13_2562 <= 0;
        i_13_2563 <= 0;
        i_13_2564 <= 0;
        i_13_2565 <= 0;
        i_13_2566 <= 0;
        i_13_2567 <= 0;
        i_13_2568 <= 0;
        i_13_2569 <= 0;
        i_13_2570 <= 0;
        i_13_2571 <= 0;
        i_13_2572 <= 0;
        i_13_2573 <= 0;
        i_13_2574 <= 0;
        i_13_2575 <= 0;
        i_13_2576 <= 0;
        i_13_2577 <= 0;
        i_13_2578 <= 0;
        i_13_2579 <= 0;
        i_13_2580 <= 0;
        i_13_2581 <= 0;
        i_13_2582 <= 0;
        i_13_2583 <= 0;
        i_13_2584 <= 0;
        i_13_2585 <= 0;
        i_13_2586 <= 0;
        i_13_2587 <= 0;
        i_13_2588 <= 0;
        i_13_2589 <= 0;
        i_13_2590 <= 0;
        i_13_2591 <= 0;
        i_13_2592 <= 0;
        i_13_2593 <= 0;
        i_13_2594 <= 0;
        i_13_2595 <= 0;
        i_13_2596 <= 0;
        i_13_2597 <= 0;
        i_13_2598 <= 0;
        i_13_2599 <= 0;
        i_13_2600 <= 0;
        i_13_2601 <= 0;
        i_13_2602 <= 0;
        i_13_2603 <= 0;
        i_13_2604 <= 0;
        i_13_2605 <= 0;
        i_13_2606 <= 0;
        i_13_2607 <= 0;
        i_13_2608 <= 0;
        i_13_2609 <= 0;
        i_13_2610 <= 0;
        i_13_2611 <= 0;
        i_13_2612 <= 0;
        i_13_2613 <= 0;
        i_13_2614 <= 0;
        i_13_2615 <= 0;
        i_13_2616 <= 0;
        i_13_2617 <= 0;
        i_13_2618 <= 0;
        i_13_2619 <= 0;
        i_13_2620 <= 0;
        i_13_2621 <= 0;
        i_13_2622 <= 0;
        i_13_2623 <= 0;
        i_13_2624 <= 0;
        i_13_2625 <= 0;
        i_13_2626 <= 0;
        i_13_2627 <= 0;
        i_13_2628 <= 0;
        i_13_2629 <= 0;
        i_13_2630 <= 0;
        i_13_2631 <= 0;
        i_13_2632 <= 0;
        i_13_2633 <= 0;
        i_13_2634 <= 0;
        i_13_2635 <= 0;
        i_13_2636 <= 0;
        i_13_2637 <= 0;
        i_13_2638 <= 0;
        i_13_2639 <= 0;
        i_13_2640 <= 0;
        i_13_2641 <= 0;
        i_13_2642 <= 0;
        i_13_2643 <= 0;
        i_13_2644 <= 0;
        i_13_2645 <= 0;
        i_13_2646 <= 0;
        i_13_2647 <= 0;
        i_13_2648 <= 0;
        i_13_2649 <= 0;
        i_13_2650 <= 0;
        i_13_2651 <= 0;
        i_13_2652 <= 0;
        i_13_2653 <= 0;
        i_13_2654 <= 0;
        i_13_2655 <= 0;
        i_13_2656 <= 0;
        i_13_2657 <= 0;
        i_13_2658 <= 0;
        i_13_2659 <= 0;
        i_13_2660 <= 0;
        i_13_2661 <= 0;
        i_13_2662 <= 0;
        i_13_2663 <= 0;
        i_13_2664 <= 0;
        i_13_2665 <= 0;
        i_13_2666 <= 0;
        i_13_2667 <= 0;
        i_13_2668 <= 0;
        i_13_2669 <= 0;
        i_13_2670 <= 0;
        i_13_2671 <= 0;
        i_13_2672 <= 0;
        i_13_2673 <= 0;
        i_13_2674 <= 0;
        i_13_2675 <= 0;
        i_13_2676 <= 0;
        i_13_2677 <= 0;
        i_13_2678 <= 0;
        i_13_2679 <= 0;
        i_13_2680 <= 0;
        i_13_2681 <= 0;
        i_13_2682 <= 0;
        i_13_2683 <= 0;
        i_13_2684 <= 0;
        i_13_2685 <= 0;
        i_13_2686 <= 0;
        i_13_2687 <= 0;
        i_13_2688 <= 0;
        i_13_2689 <= 0;
        i_13_2690 <= 0;
        i_13_2691 <= 0;
        i_13_2692 <= 0;
        i_13_2693 <= 0;
        i_13_2694 <= 0;
        i_13_2695 <= 0;
        i_13_2696 <= 0;
        i_13_2697 <= 0;
        i_13_2698 <= 0;
        i_13_2699 <= 0;
        i_13_2700 <= 0;
        i_13_2701 <= 0;
        i_13_2702 <= 0;
        i_13_2703 <= 0;
        i_13_2704 <= 0;
        i_13_2705 <= 0;
        i_13_2706 <= 0;
        i_13_2707 <= 0;
        i_13_2708 <= 0;
        i_13_2709 <= 0;
        i_13_2710 <= 0;
        i_13_2711 <= 0;
        i_13_2712 <= 0;
        i_13_2713 <= 0;
        i_13_2714 <= 0;
        i_13_2715 <= 0;
        i_13_2716 <= 0;
        i_13_2717 <= 0;
        i_13_2718 <= 0;
        i_13_2719 <= 0;
        i_13_2720 <= 0;
        i_13_2721 <= 0;
        i_13_2722 <= 0;
        i_13_2723 <= 0;
        i_13_2724 <= 0;
        i_13_2725 <= 0;
        i_13_2726 <= 0;
        i_13_2727 <= 0;
        i_13_2728 <= 0;
        i_13_2729 <= 0;
        i_13_2730 <= 0;
        i_13_2731 <= 0;
        i_13_2732 <= 0;
        i_13_2733 <= 0;
        i_13_2734 <= 0;
        i_13_2735 <= 0;
        i_13_2736 <= 0;
        i_13_2737 <= 0;
        i_13_2738 <= 0;
        i_13_2739 <= 0;
        i_13_2740 <= 0;
        i_13_2741 <= 0;
        i_13_2742 <= 0;
        i_13_2743 <= 0;
        i_13_2744 <= 0;
        i_13_2745 <= 0;
        i_13_2746 <= 0;
        i_13_2747 <= 0;
        i_13_2748 <= 0;
        i_13_2749 <= 0;
        i_13_2750 <= 0;
        i_13_2751 <= 0;
        i_13_2752 <= 0;
        i_13_2753 <= 0;
        i_13_2754 <= 0;
        i_13_2755 <= 0;
        i_13_2756 <= 0;
        i_13_2757 <= 0;
        i_13_2758 <= 0;
        i_13_2759 <= 0;
        i_13_2760 <= 0;
        i_13_2761 <= 0;
        i_13_2762 <= 0;
        i_13_2763 <= 0;
        i_13_2764 <= 0;
        i_13_2765 <= 0;
        i_13_2766 <= 0;
        i_13_2767 <= 0;
        i_13_2768 <= 0;
        i_13_2769 <= 0;
        i_13_2770 <= 0;
        i_13_2771 <= 0;
        i_13_2772 <= 0;
        i_13_2773 <= 0;
        i_13_2774 <= 0;
        i_13_2775 <= 0;
        i_13_2776 <= 0;
        i_13_2777 <= 0;
        i_13_2778 <= 0;
        i_13_2779 <= 0;
        i_13_2780 <= 0;
        i_13_2781 <= 0;
        i_13_2782 <= 0;
        i_13_2783 <= 0;
        i_13_2784 <= 0;
        i_13_2785 <= 0;
        i_13_2786 <= 0;
        i_13_2787 <= 0;
        i_13_2788 <= 0;
        i_13_2789 <= 0;
        i_13_2790 <= 0;
        i_13_2791 <= 0;
        i_13_2792 <= 0;
        i_13_2793 <= 0;
        i_13_2794 <= 0;
        i_13_2795 <= 0;
        i_13_2796 <= 0;
        i_13_2797 <= 0;
        i_13_2798 <= 0;
        i_13_2799 <= 0;
        i_13_2800 <= 0;
        i_13_2801 <= 0;
        i_13_2802 <= 0;
        i_13_2803 <= 0;
        i_13_2804 <= 0;
        i_13_2805 <= 0;
        i_13_2806 <= 0;
        i_13_2807 <= 0;
        i_13_2808 <= 0;
        i_13_2809 <= 0;
        i_13_2810 <= 0;
        i_13_2811 <= 0;
        i_13_2812 <= 0;
        i_13_2813 <= 0;
        i_13_2814 <= 0;
        i_13_2815 <= 0;
        i_13_2816 <= 0;
        i_13_2817 <= 0;
        i_13_2818 <= 0;
        i_13_2819 <= 0;
        i_13_2820 <= 0;
        i_13_2821 <= 0;
        i_13_2822 <= 0;
        i_13_2823 <= 0;
        i_13_2824 <= 0;
        i_13_2825 <= 0;
        i_13_2826 <= 0;
        i_13_2827 <= 0;
        i_13_2828 <= 0;
        i_13_2829 <= 0;
        i_13_2830 <= 0;
        i_13_2831 <= 0;
        i_13_2832 <= 0;
        i_13_2833 <= 0;
        i_13_2834 <= 0;
        i_13_2835 <= 0;
        i_13_2836 <= 0;
        i_13_2837 <= 0;
        i_13_2838 <= 0;
        i_13_2839 <= 0;
        i_13_2840 <= 0;
        i_13_2841 <= 0;
        i_13_2842 <= 0;
        i_13_2843 <= 0;
        i_13_2844 <= 0;
        i_13_2845 <= 0;
        i_13_2846 <= 0;
        i_13_2847 <= 0;
        i_13_2848 <= 0;
        i_13_2849 <= 0;
        i_13_2850 <= 0;
        i_13_2851 <= 0;
        i_13_2852 <= 0;
        i_13_2853 <= 0;
        i_13_2854 <= 0;
        i_13_2855 <= 0;
        i_13_2856 <= 0;
        i_13_2857 <= 0;
        i_13_2858 <= 0;
        i_13_2859 <= 0;
        i_13_2860 <= 0;
        i_13_2861 <= 0;
        i_13_2862 <= 0;
        i_13_2863 <= 0;
        i_13_2864 <= 0;
        i_13_2865 <= 0;
        i_13_2866 <= 0;
        i_13_2867 <= 0;
        i_13_2868 <= 0;
        i_13_2869 <= 0;
        i_13_2870 <= 0;
        i_13_2871 <= 0;
        i_13_2872 <= 0;
        i_13_2873 <= 0;
        i_13_2874 <= 0;
        i_13_2875 <= 0;
        i_13_2876 <= 0;
        i_13_2877 <= 0;
        i_13_2878 <= 0;
        i_13_2879 <= 0;
        i_13_2880 <= 0;
        i_13_2881 <= 0;
        i_13_2882 <= 0;
        i_13_2883 <= 0;
        i_13_2884 <= 0;
        i_13_2885 <= 0;
        i_13_2886 <= 0;
        i_13_2887 <= 0;
        i_13_2888 <= 0;
        i_13_2889 <= 0;
        i_13_2890 <= 0;
        i_13_2891 <= 0;
        i_13_2892 <= 0;
        i_13_2893 <= 0;
        i_13_2894 <= 0;
        i_13_2895 <= 0;
        i_13_2896 <= 0;
        i_13_2897 <= 0;
        i_13_2898 <= 0;
        i_13_2899 <= 0;
        i_13_2900 <= 0;
        i_13_2901 <= 0;
        i_13_2902 <= 0;
        i_13_2903 <= 0;
        i_13_2904 <= 0;
        i_13_2905 <= 0;
        i_13_2906 <= 0;
        i_13_2907 <= 0;
        i_13_2908 <= 0;
        i_13_2909 <= 0;
        i_13_2910 <= 0;
        i_13_2911 <= 0;
        i_13_2912 <= 0;
        i_13_2913 <= 0;
        i_13_2914 <= 0;
        i_13_2915 <= 0;
        i_13_2916 <= 0;
        i_13_2917 <= 0;
        i_13_2918 <= 0;
        i_13_2919 <= 0;
        i_13_2920 <= 0;
        i_13_2921 <= 0;
        i_13_2922 <= 0;
        i_13_2923 <= 0;
        i_13_2924 <= 0;
        i_13_2925 <= 0;
        i_13_2926 <= 0;
        i_13_2927 <= 0;
        i_13_2928 <= 0;
        i_13_2929 <= 0;
        i_13_2930 <= 0;
        i_13_2931 <= 0;
        i_13_2932 <= 0;
        i_13_2933 <= 0;
        i_13_2934 <= 0;
        i_13_2935 <= 0;
        i_13_2936 <= 0;
        i_13_2937 <= 0;
        i_13_2938 <= 0;
        i_13_2939 <= 0;
        i_13_2940 <= 0;
        i_13_2941 <= 0;
        i_13_2942 <= 0;
        i_13_2943 <= 0;
        i_13_2944 <= 0;
        i_13_2945 <= 0;
        i_13_2946 <= 0;
        i_13_2947 <= 0;
        i_13_2948 <= 0;
        i_13_2949 <= 0;
        i_13_2950 <= 0;
        i_13_2951 <= 0;
        i_13_2952 <= 0;
        i_13_2953 <= 0;
        i_13_2954 <= 0;
        i_13_2955 <= 0;
        i_13_2956 <= 0;
        i_13_2957 <= 0;
        i_13_2958 <= 0;
        i_13_2959 <= 0;
        i_13_2960 <= 0;
        i_13_2961 <= 0;
        i_13_2962 <= 0;
        i_13_2963 <= 0;
        i_13_2964 <= 0;
        i_13_2965 <= 0;
        i_13_2966 <= 0;
        i_13_2967 <= 0;
        i_13_2968 <= 0;
        i_13_2969 <= 0;
        i_13_2970 <= 0;
        i_13_2971 <= 0;
        i_13_2972 <= 0;
        i_13_2973 <= 0;
        i_13_2974 <= 0;
        i_13_2975 <= 0;
        i_13_2976 <= 0;
        i_13_2977 <= 0;
        i_13_2978 <= 0;
        i_13_2979 <= 0;
        i_13_2980 <= 0;
        i_13_2981 <= 0;
        i_13_2982 <= 0;
        i_13_2983 <= 0;
        i_13_2984 <= 0;
        i_13_2985 <= 0;
        i_13_2986 <= 0;
        i_13_2987 <= 0;
        i_13_2988 <= 0;
        i_13_2989 <= 0;
        i_13_2990 <= 0;
        i_13_2991 <= 0;
        i_13_2992 <= 0;
        i_13_2993 <= 0;
        i_13_2994 <= 0;
        i_13_2995 <= 0;
        i_13_2996 <= 0;
        i_13_2997 <= 0;
        i_13_2998 <= 0;
        i_13_2999 <= 0;
        i_13_3000 <= 0;
        i_13_3001 <= 0;
        i_13_3002 <= 0;
        i_13_3003 <= 0;
        i_13_3004 <= 0;
        i_13_3005 <= 0;
        i_13_3006 <= 0;
        i_13_3007 <= 0;
        i_13_3008 <= 0;
        i_13_3009 <= 0;
        i_13_3010 <= 0;
        i_13_3011 <= 0;
        i_13_3012 <= 0;
        i_13_3013 <= 0;
        i_13_3014 <= 0;
        i_13_3015 <= 0;
        i_13_3016 <= 0;
        i_13_3017 <= 0;
        i_13_3018 <= 0;
        i_13_3019 <= 0;
        i_13_3020 <= 0;
        i_13_3021 <= 0;
        i_13_3022 <= 0;
        i_13_3023 <= 0;
        i_13_3024 <= 0;
        i_13_3025 <= 0;
        i_13_3026 <= 0;
        i_13_3027 <= 0;
        i_13_3028 <= 0;
        i_13_3029 <= 0;
        i_13_3030 <= 0;
        i_13_3031 <= 0;
        i_13_3032 <= 0;
        i_13_3033 <= 0;
        i_13_3034 <= 0;
        i_13_3035 <= 0;
        i_13_3036 <= 0;
        i_13_3037 <= 0;
        i_13_3038 <= 0;
        i_13_3039 <= 0;
        i_13_3040 <= 0;
        i_13_3041 <= 0;
        i_13_3042 <= 0;
        i_13_3043 <= 0;
        i_13_3044 <= 0;
        i_13_3045 <= 0;
        i_13_3046 <= 0;
        i_13_3047 <= 0;
        i_13_3048 <= 0;
        i_13_3049 <= 0;
        i_13_3050 <= 0;
        i_13_3051 <= 0;
        i_13_3052 <= 0;
        i_13_3053 <= 0;
        i_13_3054 <= 0;
        i_13_3055 <= 0;
        i_13_3056 <= 0;
        i_13_3057 <= 0;
        i_13_3058 <= 0;
        i_13_3059 <= 0;
        i_13_3060 <= 0;
        i_13_3061 <= 0;
        i_13_3062 <= 0;
        i_13_3063 <= 0;
        i_13_3064 <= 0;
        i_13_3065 <= 0;
        i_13_3066 <= 0;
        i_13_3067 <= 0;
        i_13_3068 <= 0;
        i_13_3069 <= 0;
        i_13_3070 <= 0;
        i_13_3071 <= 0;
        i_13_3072 <= 0;
        i_13_3073 <= 0;
        i_13_3074 <= 0;
        i_13_3075 <= 0;
        i_13_3076 <= 0;
        i_13_3077 <= 0;
        i_13_3078 <= 0;
        i_13_3079 <= 0;
        i_13_3080 <= 0;
        i_13_3081 <= 0;
        i_13_3082 <= 0;
        i_13_3083 <= 0;
        i_13_3084 <= 0;
        i_13_3085 <= 0;
        i_13_3086 <= 0;
        i_13_3087 <= 0;
        i_13_3088 <= 0;
        i_13_3089 <= 0;
        i_13_3090 <= 0;
        i_13_3091 <= 0;
        i_13_3092 <= 0;
        i_13_3093 <= 0;
        i_13_3094 <= 0;
        i_13_3095 <= 0;
        i_13_3096 <= 0;
        i_13_3097 <= 0;
        i_13_3098 <= 0;
        i_13_3099 <= 0;
        i_13_3100 <= 0;
        i_13_3101 <= 0;
        i_13_3102 <= 0;
        i_13_3103 <= 0;
        i_13_3104 <= 0;
        i_13_3105 <= 0;
        i_13_3106 <= 0;
        i_13_3107 <= 0;
        i_13_3108 <= 0;
        i_13_3109 <= 0;
        i_13_3110 <= 0;
        i_13_3111 <= 0;
        i_13_3112 <= 0;
        i_13_3113 <= 0;
        i_13_3114 <= 0;
        i_13_3115 <= 0;
        i_13_3116 <= 0;
        i_13_3117 <= 0;
        i_13_3118 <= 0;
        i_13_3119 <= 0;
        i_13_3120 <= 0;
        i_13_3121 <= 0;
        i_13_3122 <= 0;
        i_13_3123 <= 0;
        i_13_3124 <= 0;
        i_13_3125 <= 0;
        i_13_3126 <= 0;
        i_13_3127 <= 0;
        i_13_3128 <= 0;
        i_13_3129 <= 0;
        i_13_3130 <= 0;
        i_13_3131 <= 0;
        i_13_3132 <= 0;
        i_13_3133 <= 0;
        i_13_3134 <= 0;
        i_13_3135 <= 0;
        i_13_3136 <= 0;
        i_13_3137 <= 0;
        i_13_3138 <= 0;
        i_13_3139 <= 0;
        i_13_3140 <= 0;
        i_13_3141 <= 0;
        i_13_3142 <= 0;
        i_13_3143 <= 0;
        i_13_3144 <= 0;
        i_13_3145 <= 0;
        i_13_3146 <= 0;
        i_13_3147 <= 0;
        i_13_3148 <= 0;
        i_13_3149 <= 0;
        i_13_3150 <= 0;
        i_13_3151 <= 0;
        i_13_3152 <= 0;
        i_13_3153 <= 0;
        i_13_3154 <= 0;
        i_13_3155 <= 0;
        i_13_3156 <= 0;
        i_13_3157 <= 0;
        i_13_3158 <= 0;
        i_13_3159 <= 0;
        i_13_3160 <= 0;
        i_13_3161 <= 0;
        i_13_3162 <= 0;
        i_13_3163 <= 0;
        i_13_3164 <= 0;
        i_13_3165 <= 0;
        i_13_3166 <= 0;
        i_13_3167 <= 0;
        i_13_3168 <= 0;
        i_13_3169 <= 0;
        i_13_3170 <= 0;
        i_13_3171 <= 0;
        i_13_3172 <= 0;
        i_13_3173 <= 0;
        i_13_3174 <= 0;
        i_13_3175 <= 0;
        i_13_3176 <= 0;
        i_13_3177 <= 0;
        i_13_3178 <= 0;
        i_13_3179 <= 0;
        i_13_3180 <= 0;
        i_13_3181 <= 0;
        i_13_3182 <= 0;
        i_13_3183 <= 0;
        i_13_3184 <= 0;
        i_13_3185 <= 0;
        i_13_3186 <= 0;
        i_13_3187 <= 0;
        i_13_3188 <= 0;
        i_13_3189 <= 0;
        i_13_3190 <= 0;
        i_13_3191 <= 0;
        i_13_3192 <= 0;
        i_13_3193 <= 0;
        i_13_3194 <= 0;
        i_13_3195 <= 0;
        i_13_3196 <= 0;
        i_13_3197 <= 0;
        i_13_3198 <= 0;
        i_13_3199 <= 0;
        i_13_3200 <= 0;
        i_13_3201 <= 0;
        i_13_3202 <= 0;
        i_13_3203 <= 0;
        i_13_3204 <= 0;
        i_13_3205 <= 0;
        i_13_3206 <= 0;
        i_13_3207 <= 0;
        i_13_3208 <= 0;
        i_13_3209 <= 0;
        i_13_3210 <= 0;
        i_13_3211 <= 0;
        i_13_3212 <= 0;
        i_13_3213 <= 0;
        i_13_3214 <= 0;
        i_13_3215 <= 0;
        i_13_3216 <= 0;
        i_13_3217 <= 0;
        i_13_3218 <= 0;
        i_13_3219 <= 0;
        i_13_3220 <= 0;
        i_13_3221 <= 0;
        i_13_3222 <= 0;
        i_13_3223 <= 0;
        i_13_3224 <= 0;
        i_13_3225 <= 0;
        i_13_3226 <= 0;
        i_13_3227 <= 0;
        i_13_3228 <= 0;
        i_13_3229 <= 0;
        i_13_3230 <= 0;
        i_13_3231 <= 0;
        i_13_3232 <= 0;
        i_13_3233 <= 0;
        i_13_3234 <= 0;
        i_13_3235 <= 0;
        i_13_3236 <= 0;
        i_13_3237 <= 0;
        i_13_3238 <= 0;
        i_13_3239 <= 0;
        i_13_3240 <= 0;
        i_13_3241 <= 0;
        i_13_3242 <= 0;
        i_13_3243 <= 0;
        i_13_3244 <= 0;
        i_13_3245 <= 0;
        i_13_3246 <= 0;
        i_13_3247 <= 0;
        i_13_3248 <= 0;
        i_13_3249 <= 0;
        i_13_3250 <= 0;
        i_13_3251 <= 0;
        i_13_3252 <= 0;
        i_13_3253 <= 0;
        i_13_3254 <= 0;
        i_13_3255 <= 0;
        i_13_3256 <= 0;
        i_13_3257 <= 0;
        i_13_3258 <= 0;
        i_13_3259 <= 0;
        i_13_3260 <= 0;
        i_13_3261 <= 0;
        i_13_3262 <= 0;
        i_13_3263 <= 0;
        i_13_3264 <= 0;
        i_13_3265 <= 0;
        i_13_3266 <= 0;
        i_13_3267 <= 0;
        i_13_3268 <= 0;
        i_13_3269 <= 0;
        i_13_3270 <= 0;
        i_13_3271 <= 0;
        i_13_3272 <= 0;
        i_13_3273 <= 0;
        i_13_3274 <= 0;
        i_13_3275 <= 0;
        i_13_3276 <= 0;
        i_13_3277 <= 0;
        i_13_3278 <= 0;
        i_13_3279 <= 0;
        i_13_3280 <= 0;
        i_13_3281 <= 0;
        i_13_3282 <= 0;
        i_13_3283 <= 0;
        i_13_3284 <= 0;
        i_13_3285 <= 0;
        i_13_3286 <= 0;
        i_13_3287 <= 0;
        i_13_3288 <= 0;
        i_13_3289 <= 0;
        i_13_3290 <= 0;
        i_13_3291 <= 0;
        i_13_3292 <= 0;
        i_13_3293 <= 0;
        i_13_3294 <= 0;
        i_13_3295 <= 0;
        i_13_3296 <= 0;
        i_13_3297 <= 0;
        i_13_3298 <= 0;
        i_13_3299 <= 0;
        i_13_3300 <= 0;
        i_13_3301 <= 0;
        i_13_3302 <= 0;
        i_13_3303 <= 0;
        i_13_3304 <= 0;
        i_13_3305 <= 0;
        i_13_3306 <= 0;
        i_13_3307 <= 0;
        i_13_3308 <= 0;
        i_13_3309 <= 0;
        i_13_3310 <= 0;
        i_13_3311 <= 0;
        i_13_3312 <= 0;
        i_13_3313 <= 0;
        i_13_3314 <= 0;
        i_13_3315 <= 0;
        i_13_3316 <= 0;
        i_13_3317 <= 0;
        i_13_3318 <= 0;
        i_13_3319 <= 0;
        i_13_3320 <= 0;
        i_13_3321 <= 0;
        i_13_3322 <= 0;
        i_13_3323 <= 0;
        i_13_3324 <= 0;
        i_13_3325 <= 0;
        i_13_3326 <= 0;
        i_13_3327 <= 0;
        i_13_3328 <= 0;
        i_13_3329 <= 0;
        i_13_3330 <= 0;
        i_13_3331 <= 0;
        i_13_3332 <= 0;
        i_13_3333 <= 0;
        i_13_3334 <= 0;
        i_13_3335 <= 0;
        i_13_3336 <= 0;
        i_13_3337 <= 0;
        i_13_3338 <= 0;
        i_13_3339 <= 0;
        i_13_3340 <= 0;
        i_13_3341 <= 0;
        i_13_3342 <= 0;
        i_13_3343 <= 0;
        i_13_3344 <= 0;
        i_13_3345 <= 0;
        i_13_3346 <= 0;
        i_13_3347 <= 0;
        i_13_3348 <= 0;
        i_13_3349 <= 0;
        i_13_3350 <= 0;
        i_13_3351 <= 0;
        i_13_3352 <= 0;
        i_13_3353 <= 0;
        i_13_3354 <= 0;
        i_13_3355 <= 0;
        i_13_3356 <= 0;
        i_13_3357 <= 0;
        i_13_3358 <= 0;
        i_13_3359 <= 0;
        i_13_3360 <= 0;
        i_13_3361 <= 0;
        i_13_3362 <= 0;
        i_13_3363 <= 0;
        i_13_3364 <= 0;
        i_13_3365 <= 0;
        i_13_3366 <= 0;
        i_13_3367 <= 0;
        i_13_3368 <= 0;
        i_13_3369 <= 0;
        i_13_3370 <= 0;
        i_13_3371 <= 0;
        i_13_3372 <= 0;
        i_13_3373 <= 0;
        i_13_3374 <= 0;
        i_13_3375 <= 0;
        i_13_3376 <= 0;
        i_13_3377 <= 0;
        i_13_3378 <= 0;
        i_13_3379 <= 0;
        i_13_3380 <= 0;
        i_13_3381 <= 0;
        i_13_3382 <= 0;
        i_13_3383 <= 0;
        i_13_3384 <= 0;
        i_13_3385 <= 0;
        i_13_3386 <= 0;
        i_13_3387 <= 0;
        i_13_3388 <= 0;
        i_13_3389 <= 0;
        i_13_3390 <= 0;
        i_13_3391 <= 0;
        i_13_3392 <= 0;
        i_13_3393 <= 0;
        i_13_3394 <= 0;
        i_13_3395 <= 0;
        i_13_3396 <= 0;
        i_13_3397 <= 0;
        i_13_3398 <= 0;
        i_13_3399 <= 0;
        i_13_3400 <= 0;
        i_13_3401 <= 0;
        i_13_3402 <= 0;
        i_13_3403 <= 0;
        i_13_3404 <= 0;
        i_13_3405 <= 0;
        i_13_3406 <= 0;
        i_13_3407 <= 0;
        i_13_3408 <= 0;
        i_13_3409 <= 0;
        i_13_3410 <= 0;
        i_13_3411 <= 0;
        i_13_3412 <= 0;
        i_13_3413 <= 0;
        i_13_3414 <= 0;
        i_13_3415 <= 0;
        i_13_3416 <= 0;
        i_13_3417 <= 0;
        i_13_3418 <= 0;
        i_13_3419 <= 0;
        i_13_3420 <= 0;
        i_13_3421 <= 0;
        i_13_3422 <= 0;
        i_13_3423 <= 0;
        i_13_3424 <= 0;
        i_13_3425 <= 0;
        i_13_3426 <= 0;
        i_13_3427 <= 0;
        i_13_3428 <= 0;
        i_13_3429 <= 0;
        i_13_3430 <= 0;
        i_13_3431 <= 0;
        i_13_3432 <= 0;
        i_13_3433 <= 0;
        i_13_3434 <= 0;
        i_13_3435 <= 0;
        i_13_3436 <= 0;
        i_13_3437 <= 0;
        i_13_3438 <= 0;
        i_13_3439 <= 0;
        i_13_3440 <= 0;
        i_13_3441 <= 0;
        i_13_3442 <= 0;
        i_13_3443 <= 0;
        i_13_3444 <= 0;
        i_13_3445 <= 0;
        i_13_3446 <= 0;
        i_13_3447 <= 0;
        i_13_3448 <= 0;
        i_13_3449 <= 0;
        i_13_3450 <= 0;
        i_13_3451 <= 0;
        i_13_3452 <= 0;
        i_13_3453 <= 0;
        i_13_3454 <= 0;
        i_13_3455 <= 0;
        i_13_3456 <= 0;
        i_13_3457 <= 0;
        i_13_3458 <= 0;
        i_13_3459 <= 0;
        i_13_3460 <= 0;
        i_13_3461 <= 0;
        i_13_3462 <= 0;
        i_13_3463 <= 0;
        i_13_3464 <= 0;
        i_13_3465 <= 0;
        i_13_3466 <= 0;
        i_13_3467 <= 0;
        i_13_3468 <= 0;
        i_13_3469 <= 0;
        i_13_3470 <= 0;
        i_13_3471 <= 0;
        i_13_3472 <= 0;
        i_13_3473 <= 0;
        i_13_3474 <= 0;
        i_13_3475 <= 0;
        i_13_3476 <= 0;
        i_13_3477 <= 0;
        i_13_3478 <= 0;
        i_13_3479 <= 0;
        i_13_3480 <= 0;
        i_13_3481 <= 0;
        i_13_3482 <= 0;
        i_13_3483 <= 0;
        i_13_3484 <= 0;
        i_13_3485 <= 0;
        i_13_3486 <= 0;
        i_13_3487 <= 0;
        i_13_3488 <= 0;
        i_13_3489 <= 0;
        i_13_3490 <= 0;
        i_13_3491 <= 0;
        i_13_3492 <= 0;
        i_13_3493 <= 0;
        i_13_3494 <= 0;
        i_13_3495 <= 0;
        i_13_3496 <= 0;
        i_13_3497 <= 0;
        i_13_3498 <= 0;
        i_13_3499 <= 0;
        i_13_3500 <= 0;
        i_13_3501 <= 0;
        i_13_3502 <= 0;
        i_13_3503 <= 0;
        i_13_3504 <= 0;
        i_13_3505 <= 0;
        i_13_3506 <= 0;
        i_13_3507 <= 0;
        i_13_3508 <= 0;
        i_13_3509 <= 0;
        i_13_3510 <= 0;
        i_13_3511 <= 0;
        i_13_3512 <= 0;
        i_13_3513 <= 0;
        i_13_3514 <= 0;
        i_13_3515 <= 0;
        i_13_3516 <= 0;
        i_13_3517 <= 0;
        i_13_3518 <= 0;
        i_13_3519 <= 0;
        i_13_3520 <= 0;
        i_13_3521 <= 0;
        i_13_3522 <= 0;
        i_13_3523 <= 0;
        i_13_3524 <= 0;
        i_13_3525 <= 0;
        i_13_3526 <= 0;
        i_13_3527 <= 0;
        i_13_3528 <= 0;
        i_13_3529 <= 0;
        i_13_3530 <= 0;
        i_13_3531 <= 0;
        i_13_3532 <= 0;
        i_13_3533 <= 0;
        i_13_3534 <= 0;
        i_13_3535 <= 0;
        i_13_3536 <= 0;
        i_13_3537 <= 0;
        i_13_3538 <= 0;
        i_13_3539 <= 0;
        i_13_3540 <= 0;
        i_13_3541 <= 0;
        i_13_3542 <= 0;
        i_13_3543 <= 0;
        i_13_3544 <= 0;
        i_13_3545 <= 0;
        i_13_3546 <= 0;
        i_13_3547 <= 0;
        i_13_3548 <= 0;
        i_13_3549 <= 0;
        i_13_3550 <= 0;
        i_13_3551 <= 0;
        i_13_3552 <= 0;
        i_13_3553 <= 0;
        i_13_3554 <= 0;
        i_13_3555 <= 0;
        i_13_3556 <= 0;
        i_13_3557 <= 0;
        i_13_3558 <= 0;
        i_13_3559 <= 0;
        i_13_3560 <= 0;
        i_13_3561 <= 0;
        i_13_3562 <= 0;
        i_13_3563 <= 0;
        i_13_3564 <= 0;
        i_13_3565 <= 0;
        i_13_3566 <= 0;
        i_13_3567 <= 0;
        i_13_3568 <= 0;
        i_13_3569 <= 0;
        i_13_3570 <= 0;
        i_13_3571 <= 0;
        i_13_3572 <= 0;
        i_13_3573 <= 0;
        i_13_3574 <= 0;
        i_13_3575 <= 0;
        i_13_3576 <= 0;
        i_13_3577 <= 0;
        i_13_3578 <= 0;
        i_13_3579 <= 0;
        i_13_3580 <= 0;
        i_13_3581 <= 0;
        i_13_3582 <= 0;
        i_13_3583 <= 0;
        i_13_3584 <= 0;
        i_13_3585 <= 0;
        i_13_3586 <= 0;
        i_13_3587 <= 0;
        i_13_3588 <= 0;
        i_13_3589 <= 0;
        i_13_3590 <= 0;
        i_13_3591 <= 0;
        i_13_3592 <= 0;
        i_13_3593 <= 0;
        i_13_3594 <= 0;
        i_13_3595 <= 0;
        i_13_3596 <= 0;
        i_13_3597 <= 0;
        i_13_3598 <= 0;
        i_13_3599 <= 0;
        i_13_3600 <= 0;
        i_13_3601 <= 0;
        i_13_3602 <= 0;
        i_13_3603 <= 0;
        i_13_3604 <= 0;
        i_13_3605 <= 0;
        i_13_3606 <= 0;
        i_13_3607 <= 0;
        i_13_3608 <= 0;
        i_13_3609 <= 0;
        i_13_3610 <= 0;
        i_13_3611 <= 0;
        i_13_3612 <= 0;
        i_13_3613 <= 0;
        i_13_3614 <= 0;
        i_13_3615 <= 0;
        i_13_3616 <= 0;
        i_13_3617 <= 0;
        i_13_3618 <= 0;
        i_13_3619 <= 0;
        i_13_3620 <= 0;
        i_13_3621 <= 0;
        i_13_3622 <= 0;
        i_13_3623 <= 0;
        i_13_3624 <= 0;
        i_13_3625 <= 0;
        i_13_3626 <= 0;
        i_13_3627 <= 0;
        i_13_3628 <= 0;
        i_13_3629 <= 0;
        i_13_3630 <= 0;
        i_13_3631 <= 0;
        i_13_3632 <= 0;
        i_13_3633 <= 0;
        i_13_3634 <= 0;
        i_13_3635 <= 0;
        i_13_3636 <= 0;
        i_13_3637 <= 0;
        i_13_3638 <= 0;
        i_13_3639 <= 0;
        i_13_3640 <= 0;
        i_13_3641 <= 0;
        i_13_3642 <= 0;
        i_13_3643 <= 0;
        i_13_3644 <= 0;
        i_13_3645 <= 0;
        i_13_3646 <= 0;
        i_13_3647 <= 0;
        i_13_3648 <= 0;
        i_13_3649 <= 0;
        i_13_3650 <= 0;
        i_13_3651 <= 0;
        i_13_3652 <= 0;
        i_13_3653 <= 0;
        i_13_3654 <= 0;
        i_13_3655 <= 0;
        i_13_3656 <= 0;
        i_13_3657 <= 0;
        i_13_3658 <= 0;
        i_13_3659 <= 0;
        i_13_3660 <= 0;
        i_13_3661 <= 0;
        i_13_3662 <= 0;
        i_13_3663 <= 0;
        i_13_3664 <= 0;
        i_13_3665 <= 0;
        i_13_3666 <= 0;
        i_13_3667 <= 0;
        i_13_3668 <= 0;
        i_13_3669 <= 0;
        i_13_3670 <= 0;
        i_13_3671 <= 0;
        i_13_3672 <= 0;
        i_13_3673 <= 0;
        i_13_3674 <= 0;
        i_13_3675 <= 0;
        i_13_3676 <= 0;
        i_13_3677 <= 0;
        i_13_3678 <= 0;
        i_13_3679 <= 0;
        i_13_3680 <= 0;
        i_13_3681 <= 0;
        i_13_3682 <= 0;
        i_13_3683 <= 0;
        i_13_3684 <= 0;
        i_13_3685 <= 0;
        i_13_3686 <= 0;
        i_13_3687 <= 0;
        i_13_3688 <= 0;
        i_13_3689 <= 0;
        i_13_3690 <= 0;
        i_13_3691 <= 0;
        i_13_3692 <= 0;
        i_13_3693 <= 0;
        i_13_3694 <= 0;
        i_13_3695 <= 0;
        i_13_3696 <= 0;
        i_13_3697 <= 0;
        i_13_3698 <= 0;
        i_13_3699 <= 0;
        i_13_3700 <= 0;
        i_13_3701 <= 0;
        i_13_3702 <= 0;
        i_13_3703 <= 0;
        i_13_3704 <= 0;
        i_13_3705 <= 0;
        i_13_3706 <= 0;
        i_13_3707 <= 0;
        i_13_3708 <= 0;
        i_13_3709 <= 0;
        i_13_3710 <= 0;
        i_13_3711 <= 0;
        i_13_3712 <= 0;
        i_13_3713 <= 0;
        i_13_3714 <= 0;
        i_13_3715 <= 0;
        i_13_3716 <= 0;
        i_13_3717 <= 0;
        i_13_3718 <= 0;
        i_13_3719 <= 0;
        i_13_3720 <= 0;
        i_13_3721 <= 0;
        i_13_3722 <= 0;
        i_13_3723 <= 0;
        i_13_3724 <= 0;
        i_13_3725 <= 0;
        i_13_3726 <= 0;
        i_13_3727 <= 0;
        i_13_3728 <= 0;
        i_13_3729 <= 0;
        i_13_3730 <= 0;
        i_13_3731 <= 0;
        i_13_3732 <= 0;
        i_13_3733 <= 0;
        i_13_3734 <= 0;
        i_13_3735 <= 0;
        i_13_3736 <= 0;
        i_13_3737 <= 0;
        i_13_3738 <= 0;
        i_13_3739 <= 0;
        i_13_3740 <= 0;
        i_13_3741 <= 0;
        i_13_3742 <= 0;
        i_13_3743 <= 0;
        i_13_3744 <= 0;
        i_13_3745 <= 0;
        i_13_3746 <= 0;
        i_13_3747 <= 0;
        i_13_3748 <= 0;
        i_13_3749 <= 0;
        i_13_3750 <= 0;
        i_13_3751 <= 0;
        i_13_3752 <= 0;
        i_13_3753 <= 0;
        i_13_3754 <= 0;
        i_13_3755 <= 0;
        i_13_3756 <= 0;
        i_13_3757 <= 0;
        i_13_3758 <= 0;
        i_13_3759 <= 0;
        i_13_3760 <= 0;
        i_13_3761 <= 0;
        i_13_3762 <= 0;
        i_13_3763 <= 0;
        i_13_3764 <= 0;
        i_13_3765 <= 0;
        i_13_3766 <= 0;
        i_13_3767 <= 0;
        i_13_3768 <= 0;
        i_13_3769 <= 0;
        i_13_3770 <= 0;
        i_13_3771 <= 0;
        i_13_3772 <= 0;
        i_13_3773 <= 0;
        i_13_3774 <= 0;
        i_13_3775 <= 0;
        i_13_3776 <= 0;
        i_13_3777 <= 0;
        i_13_3778 <= 0;
        i_13_3779 <= 0;
        i_13_3780 <= 0;
        i_13_3781 <= 0;
        i_13_3782 <= 0;
        i_13_3783 <= 0;
        i_13_3784 <= 0;
        i_13_3785 <= 0;
        i_13_3786 <= 0;
        i_13_3787 <= 0;
        i_13_3788 <= 0;
        i_13_3789 <= 0;
        i_13_3790 <= 0;
        i_13_3791 <= 0;
        i_13_3792 <= 0;
        i_13_3793 <= 0;
        i_13_3794 <= 0;
        i_13_3795 <= 0;
        i_13_3796 <= 0;
        i_13_3797 <= 0;
        i_13_3798 <= 0;
        i_13_3799 <= 0;
        i_13_3800 <= 0;
        i_13_3801 <= 0;
        i_13_3802 <= 0;
        i_13_3803 <= 0;
        i_13_3804 <= 0;
        i_13_3805 <= 0;
        i_13_3806 <= 0;
        i_13_3807 <= 0;
        i_13_3808 <= 0;
        i_13_3809 <= 0;
        i_13_3810 <= 0;
        i_13_3811 <= 0;
        i_13_3812 <= 0;
        i_13_3813 <= 0;
        i_13_3814 <= 0;
        i_13_3815 <= 0;
        i_13_3816 <= 0;
        i_13_3817 <= 0;
        i_13_3818 <= 0;
        i_13_3819 <= 0;
        i_13_3820 <= 0;
        i_13_3821 <= 0;
        i_13_3822 <= 0;
        i_13_3823 <= 0;
        i_13_3824 <= 0;
        i_13_3825 <= 0;
        i_13_3826 <= 0;
        i_13_3827 <= 0;
        i_13_3828 <= 0;
        i_13_3829 <= 0;
        i_13_3830 <= 0;
        i_13_3831 <= 0;
        i_13_3832 <= 0;
        i_13_3833 <= 0;
        i_13_3834 <= 0;
        i_13_3835 <= 0;
        i_13_3836 <= 0;
        i_13_3837 <= 0;
        i_13_3838 <= 0;
        i_13_3839 <= 0;
        i_13_3840 <= 0;
        i_13_3841 <= 0;
        i_13_3842 <= 0;
        i_13_3843 <= 0;
        i_13_3844 <= 0;
        i_13_3845 <= 0;
        i_13_3846 <= 0;
        i_13_3847 <= 0;
        i_13_3848 <= 0;
        i_13_3849 <= 0;
        i_13_3850 <= 0;
        i_13_3851 <= 0;
        i_13_3852 <= 0;
        i_13_3853 <= 0;
        i_13_3854 <= 0;
        i_13_3855 <= 0;
        i_13_3856 <= 0;
        i_13_3857 <= 0;
        i_13_3858 <= 0;
        i_13_3859 <= 0;
        i_13_3860 <= 0;
        i_13_3861 <= 0;
        i_13_3862 <= 0;
        i_13_3863 <= 0;
        i_13_3864 <= 0;
        i_13_3865 <= 0;
        i_13_3866 <= 0;
        i_13_3867 <= 0;
        i_13_3868 <= 0;
        i_13_3869 <= 0;
        i_13_3870 <= 0;
        i_13_3871 <= 0;
        i_13_3872 <= 0;
        i_13_3873 <= 0;
        i_13_3874 <= 0;
        i_13_3875 <= 0;
        i_13_3876 <= 0;
        i_13_3877 <= 0;
        i_13_3878 <= 0;
        i_13_3879 <= 0;
        i_13_3880 <= 0;
        i_13_3881 <= 0;
        i_13_3882 <= 0;
        i_13_3883 <= 0;
        i_13_3884 <= 0;
        i_13_3885 <= 0;
        i_13_3886 <= 0;
        i_13_3887 <= 0;
        i_13_3888 <= 0;
        i_13_3889 <= 0;
        i_13_3890 <= 0;
        i_13_3891 <= 0;
        i_13_3892 <= 0;
        i_13_3893 <= 0;
        i_13_3894 <= 0;
        i_13_3895 <= 0;
        i_13_3896 <= 0;
        i_13_3897 <= 0;
        i_13_3898 <= 0;
        i_13_3899 <= 0;
        i_13_3900 <= 0;
        i_13_3901 <= 0;
        i_13_3902 <= 0;
        i_13_3903 <= 0;
        i_13_3904 <= 0;
        i_13_3905 <= 0;
        i_13_3906 <= 0;
        i_13_3907 <= 0;
        i_13_3908 <= 0;
        i_13_3909 <= 0;
        i_13_3910 <= 0;
        i_13_3911 <= 0;
        i_13_3912 <= 0;
        i_13_3913 <= 0;
        i_13_3914 <= 0;
        i_13_3915 <= 0;
        i_13_3916 <= 0;
        i_13_3917 <= 0;
        i_13_3918 <= 0;
        i_13_3919 <= 0;
        i_13_3920 <= 0;
        i_13_3921 <= 0;
        i_13_3922 <= 0;
        i_13_3923 <= 0;
        i_13_3924 <= 0;
        i_13_3925 <= 0;
        i_13_3926 <= 0;
        i_13_3927 <= 0;
        i_13_3928 <= 0;
        i_13_3929 <= 0;
        i_13_3930 <= 0;
        i_13_3931 <= 0;
        i_13_3932 <= 0;
        i_13_3933 <= 0;
        i_13_3934 <= 0;
        i_13_3935 <= 0;
        i_13_3936 <= 0;
        i_13_3937 <= 0;
        i_13_3938 <= 0;
        i_13_3939 <= 0;
        i_13_3940 <= 0;
        i_13_3941 <= 0;
        i_13_3942 <= 0;
        i_13_3943 <= 0;
        i_13_3944 <= 0;
        i_13_3945 <= 0;
        i_13_3946 <= 0;
        i_13_3947 <= 0;
        i_13_3948 <= 0;
        i_13_3949 <= 0;
        i_13_3950 <= 0;
        i_13_3951 <= 0;
        i_13_3952 <= 0;
        i_13_3953 <= 0;
        i_13_3954 <= 0;
        i_13_3955 <= 0;
        i_13_3956 <= 0;
        i_13_3957 <= 0;
        i_13_3958 <= 0;
        i_13_3959 <= 0;
        i_13_3960 <= 0;
        i_13_3961 <= 0;
        i_13_3962 <= 0;
        i_13_3963 <= 0;
        i_13_3964 <= 0;
        i_13_3965 <= 0;
        i_13_3966 <= 0;
        i_13_3967 <= 0;
        i_13_3968 <= 0;
        i_13_3969 <= 0;
        i_13_3970 <= 0;
        i_13_3971 <= 0;
        i_13_3972 <= 0;
        i_13_3973 <= 0;
        i_13_3974 <= 0;
        i_13_3975 <= 0;
        i_13_3976 <= 0;
        i_13_3977 <= 0;
        i_13_3978 <= 0;
        i_13_3979 <= 0;
        i_13_3980 <= 0;
        i_13_3981 <= 0;
        i_13_3982 <= 0;
        i_13_3983 <= 0;
        i_13_3984 <= 0;
        i_13_3985 <= 0;
        i_13_3986 <= 0;
        i_13_3987 <= 0;
        i_13_3988 <= 0;
        i_13_3989 <= 0;
        i_13_3990 <= 0;
        i_13_3991 <= 0;
        i_13_3992 <= 0;
        i_13_3993 <= 0;
        i_13_3994 <= 0;
        i_13_3995 <= 0;
        i_13_3996 <= 0;
        i_13_3997 <= 0;
        i_13_3998 <= 0;
        i_13_3999 <= 0;
        i_13_4000 <= 0;
        i_13_4001 <= 0;
        i_13_4002 <= 0;
        i_13_4003 <= 0;
        i_13_4004 <= 0;
        i_13_4005 <= 0;
        i_13_4006 <= 0;
        i_13_4007 <= 0;
        i_13_4008 <= 0;
        i_13_4009 <= 0;
        i_13_4010 <= 0;
        i_13_4011 <= 0;
        i_13_4012 <= 0;
        i_13_4013 <= 0;
        i_13_4014 <= 0;
        i_13_4015 <= 0;
        i_13_4016 <= 0;
        i_13_4017 <= 0;
        i_13_4018 <= 0;
        i_13_4019 <= 0;
        i_13_4020 <= 0;
        i_13_4021 <= 0;
        i_13_4022 <= 0;
        i_13_4023 <= 0;
        i_13_4024 <= 0;
        i_13_4025 <= 0;
        i_13_4026 <= 0;
        i_13_4027 <= 0;
        i_13_4028 <= 0;
        i_13_4029 <= 0;
        i_13_4030 <= 0;
        i_13_4031 <= 0;
        i_13_4032 <= 0;
        i_13_4033 <= 0;
        i_13_4034 <= 0;
        i_13_4035 <= 0;
        i_13_4036 <= 0;
        i_13_4037 <= 0;
        i_13_4038 <= 0;
        i_13_4039 <= 0;
        i_13_4040 <= 0;
        i_13_4041 <= 0;
        i_13_4042 <= 0;
        i_13_4043 <= 0;
        i_13_4044 <= 0;
        i_13_4045 <= 0;
        i_13_4046 <= 0;
        i_13_4047 <= 0;
        i_13_4048 <= 0;
        i_13_4049 <= 0;
        i_13_4050 <= 0;
        i_13_4051 <= 0;
        i_13_4052 <= 0;
        i_13_4053 <= 0;
        i_13_4054 <= 0;
        i_13_4055 <= 0;
        i_13_4056 <= 0;
        i_13_4057 <= 0;
        i_13_4058 <= 0;
        i_13_4059 <= 0;
        i_13_4060 <= 0;
        i_13_4061 <= 0;
        i_13_4062 <= 0;
        i_13_4063 <= 0;
        i_13_4064 <= 0;
        i_13_4065 <= 0;
        i_13_4066 <= 0;
        i_13_4067 <= 0;
        i_13_4068 <= 0;
        i_13_4069 <= 0;
        i_13_4070 <= 0;
        i_13_4071 <= 0;
        i_13_4072 <= 0;
        i_13_4073 <= 0;
        i_13_4074 <= 0;
        i_13_4075 <= 0;
        i_13_4076 <= 0;
        i_13_4077 <= 0;
        i_13_4078 <= 0;
        i_13_4079 <= 0;
        i_13_4080 <= 0;
        i_13_4081 <= 0;
        i_13_4082 <= 0;
        i_13_4083 <= 0;
        i_13_4084 <= 0;
        i_13_4085 <= 0;
        i_13_4086 <= 0;
        i_13_4087 <= 0;
        i_13_4088 <= 0;
        i_13_4089 <= 0;
        i_13_4090 <= 0;
        i_13_4091 <= 0;
        i_13_4092 <= 0;
        i_13_4093 <= 0;
        i_13_4094 <= 0;
        i_13_4095 <= 0;
        i_13_4096 <= 0;
        i_13_4097 <= 0;
        i_13_4098 <= 0;
        i_13_4099 <= 0;
        i_13_4100 <= 0;
        i_13_4101 <= 0;
        i_13_4102 <= 0;
        i_13_4103 <= 0;
        i_13_4104 <= 0;
        i_13_4105 <= 0;
        i_13_4106 <= 0;
        i_13_4107 <= 0;
        i_13_4108 <= 0;
        i_13_4109 <= 0;
        i_13_4110 <= 0;
        i_13_4111 <= 0;
        i_13_4112 <= 0;
        i_13_4113 <= 0;
        i_13_4114 <= 0;
        i_13_4115 <= 0;
        i_13_4116 <= 0;
        i_13_4117 <= 0;
        i_13_4118 <= 0;
        i_13_4119 <= 0;
        i_13_4120 <= 0;
        i_13_4121 <= 0;
        i_13_4122 <= 0;
        i_13_4123 <= 0;
        i_13_4124 <= 0;
        i_13_4125 <= 0;
        i_13_4126 <= 0;
        i_13_4127 <= 0;
        i_13_4128 <= 0;
        i_13_4129 <= 0;
        i_13_4130 <= 0;
        i_13_4131 <= 0;
        i_13_4132 <= 0;
        i_13_4133 <= 0;
        i_13_4134 <= 0;
        i_13_4135 <= 0;
        i_13_4136 <= 0;
        i_13_4137 <= 0;
        i_13_4138 <= 0;
        i_13_4139 <= 0;
        i_13_4140 <= 0;
        i_13_4141 <= 0;
        i_13_4142 <= 0;
        i_13_4143 <= 0;
        i_13_4144 <= 0;
        i_13_4145 <= 0;
        i_13_4146 <= 0;
        i_13_4147 <= 0;
        i_13_4148 <= 0;
        i_13_4149 <= 0;
        i_13_4150 <= 0;
        i_13_4151 <= 0;
        i_13_4152 <= 0;
        i_13_4153 <= 0;
        i_13_4154 <= 0;
        i_13_4155 <= 0;
        i_13_4156 <= 0;
        i_13_4157 <= 0;
        i_13_4158 <= 0;
        i_13_4159 <= 0;
        i_13_4160 <= 0;
        i_13_4161 <= 0;
        i_13_4162 <= 0;
        i_13_4163 <= 0;
        i_13_4164 <= 0;
        i_13_4165 <= 0;
        i_13_4166 <= 0;
        i_13_4167 <= 0;
        i_13_4168 <= 0;
        i_13_4169 <= 0;
        i_13_4170 <= 0;
        i_13_4171 <= 0;
        i_13_4172 <= 0;
        i_13_4173 <= 0;
        i_13_4174 <= 0;
        i_13_4175 <= 0;
        i_13_4176 <= 0;
        i_13_4177 <= 0;
        i_13_4178 <= 0;
        i_13_4179 <= 0;
        i_13_4180 <= 0;
        i_13_4181 <= 0;
        i_13_4182 <= 0;
        i_13_4183 <= 0;
        i_13_4184 <= 0;
        i_13_4185 <= 0;
        i_13_4186 <= 0;
        i_13_4187 <= 0;
        i_13_4188 <= 0;
        i_13_4189 <= 0;
        i_13_4190 <= 0;
        i_13_4191 <= 0;
        i_13_4192 <= 0;
        i_13_4193 <= 0;
        i_13_4194 <= 0;
        i_13_4195 <= 0;
        i_13_4196 <= 0;
        i_13_4197 <= 0;
        i_13_4198 <= 0;
        i_13_4199 <= 0;
        i_13_4200 <= 0;
        i_13_4201 <= 0;
        i_13_4202 <= 0;
        i_13_4203 <= 0;
        i_13_4204 <= 0;
        i_13_4205 <= 0;
        i_13_4206 <= 0;
        i_13_4207 <= 0;
        i_13_4208 <= 0;
        i_13_4209 <= 0;
        i_13_4210 <= 0;
        i_13_4211 <= 0;
        i_13_4212 <= 0;
        i_13_4213 <= 0;
        i_13_4214 <= 0;
        i_13_4215 <= 0;
        i_13_4216 <= 0;
        i_13_4217 <= 0;
        i_13_4218 <= 0;
        i_13_4219 <= 0;
        i_13_4220 <= 0;
        i_13_4221 <= 0;
        i_13_4222 <= 0;
        i_13_4223 <= 0;
        i_13_4224 <= 0;
        i_13_4225 <= 0;
        i_13_4226 <= 0;
        i_13_4227 <= 0;
        i_13_4228 <= 0;
        i_13_4229 <= 0;
        i_13_4230 <= 0;
        i_13_4231 <= 0;
        i_13_4232 <= 0;
        i_13_4233 <= 0;
        i_13_4234 <= 0;
        i_13_4235 <= 0;
        i_13_4236 <= 0;
        i_13_4237 <= 0;
        i_13_4238 <= 0;
        i_13_4239 <= 0;
        i_13_4240 <= 0;
        i_13_4241 <= 0;
        i_13_4242 <= 0;
        i_13_4243 <= 0;
        i_13_4244 <= 0;
        i_13_4245 <= 0;
        i_13_4246 <= 0;
        i_13_4247 <= 0;
        i_13_4248 <= 0;
        i_13_4249 <= 0;
        i_13_4250 <= 0;
        i_13_4251 <= 0;
        i_13_4252 <= 0;
        i_13_4253 <= 0;
        i_13_4254 <= 0;
        i_13_4255 <= 0;
        i_13_4256 <= 0;
        i_13_4257 <= 0;
        i_13_4258 <= 0;
        i_13_4259 <= 0;
        i_13_4260 <= 0;
        i_13_4261 <= 0;
        i_13_4262 <= 0;
        i_13_4263 <= 0;
        i_13_4264 <= 0;
        i_13_4265 <= 0;
        i_13_4266 <= 0;
        i_13_4267 <= 0;
        i_13_4268 <= 0;
        i_13_4269 <= 0;
        i_13_4270 <= 0;
        i_13_4271 <= 0;
        i_13_4272 <= 0;
        i_13_4273 <= 0;
        i_13_4274 <= 0;
        i_13_4275 <= 0;
        i_13_4276 <= 0;
        i_13_4277 <= 0;
        i_13_4278 <= 0;
        i_13_4279 <= 0;
        i_13_4280 <= 0;
        i_13_4281 <= 0;
        i_13_4282 <= 0;
        i_13_4283 <= 0;
        i_13_4284 <= 0;
        i_13_4285 <= 0;
        i_13_4286 <= 0;
        i_13_4287 <= 0;
        i_13_4288 <= 0;
        i_13_4289 <= 0;
        i_13_4290 <= 0;
        i_13_4291 <= 0;
        i_13_4292 <= 0;
        i_13_4293 <= 0;
        i_13_4294 <= 0;
        i_13_4295 <= 0;
        i_13_4296 <= 0;
        i_13_4297 <= 0;
        i_13_4298 <= 0;
        i_13_4299 <= 0;
        i_13_4300 <= 0;
        i_13_4301 <= 0;
        i_13_4302 <= 0;
        i_13_4303 <= 0;
        i_13_4304 <= 0;
        i_13_4305 <= 0;
        i_13_4306 <= 0;
        i_13_4307 <= 0;
        i_13_4308 <= 0;
        i_13_4309 <= 0;
        i_13_4310 <= 0;
        i_13_4311 <= 0;
        i_13_4312 <= 0;
        i_13_4313 <= 0;
        i_13_4314 <= 0;
        i_13_4315 <= 0;
        i_13_4316 <= 0;
        i_13_4317 <= 0;
        i_13_4318 <= 0;
        i_13_4319 <= 0;
        i_13_4320 <= 0;
        i_13_4321 <= 0;
        i_13_4322 <= 0;
        i_13_4323 <= 0;
        i_13_4324 <= 0;
        i_13_4325 <= 0;
        i_13_4326 <= 0;
        i_13_4327 <= 0;
        i_13_4328 <= 0;
        i_13_4329 <= 0;
        i_13_4330 <= 0;
        i_13_4331 <= 0;
        i_13_4332 <= 0;
        i_13_4333 <= 0;
        i_13_4334 <= 0;
        i_13_4335 <= 0;
        i_13_4336 <= 0;
        i_13_4337 <= 0;
        i_13_4338 <= 0;
        i_13_4339 <= 0;
        i_13_4340 <= 0;
        i_13_4341 <= 0;
        i_13_4342 <= 0;
        i_13_4343 <= 0;
        i_13_4344 <= 0;
        i_13_4345 <= 0;
        i_13_4346 <= 0;
        i_13_4347 <= 0;
        i_13_4348 <= 0;
        i_13_4349 <= 0;
        i_13_4350 <= 0;
        i_13_4351 <= 0;
        i_13_4352 <= 0;
        i_13_4353 <= 0;
        i_13_4354 <= 0;
        i_13_4355 <= 0;
        i_13_4356 <= 0;
        i_13_4357 <= 0;
        i_13_4358 <= 0;
        i_13_4359 <= 0;
        i_13_4360 <= 0;
        i_13_4361 <= 0;
        i_13_4362 <= 0;
        i_13_4363 <= 0;
        i_13_4364 <= 0;
        i_13_4365 <= 0;
        i_13_4366 <= 0;
        i_13_4367 <= 0;
        i_13_4368 <= 0;
        i_13_4369 <= 0;
        i_13_4370 <= 0;
        i_13_4371 <= 0;
        i_13_4372 <= 0;
        i_13_4373 <= 0;
        i_13_4374 <= 0;
        i_13_4375 <= 0;
        i_13_4376 <= 0;
        i_13_4377 <= 0;
        i_13_4378 <= 0;
        i_13_4379 <= 0;
        i_13_4380 <= 0;
        i_13_4381 <= 0;
        i_13_4382 <= 0;
        i_13_4383 <= 0;
        i_13_4384 <= 0;
        i_13_4385 <= 0;
        i_13_4386 <= 0;
        i_13_4387 <= 0;
        i_13_4388 <= 0;
        i_13_4389 <= 0;
        i_13_4390 <= 0;
        i_13_4391 <= 0;
        i_13_4392 <= 0;
        i_13_4393 <= 0;
        i_13_4394 <= 0;
        i_13_4395 <= 0;
        i_13_4396 <= 0;
        i_13_4397 <= 0;
        i_13_4398 <= 0;
        i_13_4399 <= 0;
        i_13_4400 <= 0;
        i_13_4401 <= 0;
        i_13_4402 <= 0;
        i_13_4403 <= 0;
        i_13_4404 <= 0;
        i_13_4405 <= 0;
        i_13_4406 <= 0;
        i_13_4407 <= 0;
        i_13_4408 <= 0;
        i_13_4409 <= 0;
        i_13_4410 <= 0;
        i_13_4411 <= 0;
        i_13_4412 <= 0;
        i_13_4413 <= 0;
        i_13_4414 <= 0;
        i_13_4415 <= 0;
        i_13_4416 <= 0;
        i_13_4417 <= 0;
        i_13_4418 <= 0;
        i_13_4419 <= 0;
        i_13_4420 <= 0;
        i_13_4421 <= 0;
        i_13_4422 <= 0;
        i_13_4423 <= 0;
        i_13_4424 <= 0;
        i_13_4425 <= 0;
        i_13_4426 <= 0;
        i_13_4427 <= 0;
        i_13_4428 <= 0;
        i_13_4429 <= 0;
        i_13_4430 <= 0;
        i_13_4431 <= 0;
        i_13_4432 <= 0;
        i_13_4433 <= 0;
        i_13_4434 <= 0;
        i_13_4435 <= 0;
        i_13_4436 <= 0;
        i_13_4437 <= 0;
        i_13_4438 <= 0;
        i_13_4439 <= 0;
        i_13_4440 <= 0;
        i_13_4441 <= 0;
        i_13_4442 <= 0;
        i_13_4443 <= 0;
        i_13_4444 <= 0;
        i_13_4445 <= 0;
        i_13_4446 <= 0;
        i_13_4447 <= 0;
        i_13_4448 <= 0;
        i_13_4449 <= 0;
        i_13_4450 <= 0;
        i_13_4451 <= 0;
        i_13_4452 <= 0;
        i_13_4453 <= 0;
        i_13_4454 <= 0;
        i_13_4455 <= 0;
        i_13_4456 <= 0;
        i_13_4457 <= 0;
        i_13_4458 <= 0;
        i_13_4459 <= 0;
        i_13_4460 <= 0;
        i_13_4461 <= 0;
        i_13_4462 <= 0;
        i_13_4463 <= 0;
        i_13_4464 <= 0;
        i_13_4465 <= 0;
        i_13_4466 <= 0;
        i_13_4467 <= 0;
        i_13_4468 <= 0;
        i_13_4469 <= 0;
        i_13_4470 <= 0;
        i_13_4471 <= 0;
        i_13_4472 <= 0;
        i_13_4473 <= 0;
        i_13_4474 <= 0;
        i_13_4475 <= 0;
        i_13_4476 <= 0;
        i_13_4477 <= 0;
        i_13_4478 <= 0;
        i_13_4479 <= 0;
        i_13_4480 <= 0;
        i_13_4481 <= 0;
        i_13_4482 <= 0;
        i_13_4483 <= 0;
        i_13_4484 <= 0;
        i_13_4485 <= 0;
        i_13_4486 <= 0;
        i_13_4487 <= 0;
        i_13_4488 <= 0;
        i_13_4489 <= 0;
        i_13_4490 <= 0;
        i_13_4491 <= 0;
        i_13_4492 <= 0;
        i_13_4493 <= 0;
        i_13_4494 <= 0;
        i_13_4495 <= 0;
        i_13_4496 <= 0;
        i_13_4497 <= 0;
        i_13_4498 <= 0;
        i_13_4499 <= 0;
        i_13_4500 <= 0;
        i_13_4501 <= 0;
        i_13_4502 <= 0;
        i_13_4503 <= 0;
        i_13_4504 <= 0;
        i_13_4505 <= 0;
        i_13_4506 <= 0;
        i_13_4507 <= 0;
        i_13_4508 <= 0;
        i_13_4509 <= 0;
        i_13_4510 <= 0;
        i_13_4511 <= 0;
        i_13_4512 <= 0;
        i_13_4513 <= 0;
        i_13_4514 <= 0;
        i_13_4515 <= 0;
        i_13_4516 <= 0;
        i_13_4517 <= 0;
        i_13_4518 <= 0;
        i_13_4519 <= 0;
        i_13_4520 <= 0;
        i_13_4521 <= 0;
        i_13_4522 <= 0;
        i_13_4523 <= 0;
        i_13_4524 <= 0;
        i_13_4525 <= 0;
        i_13_4526 <= 0;
        i_13_4527 <= 0;
        i_13_4528 <= 0;
        i_13_4529 <= 0;
        i_13_4530 <= 0;
        i_13_4531 <= 0;
        i_13_4532 <= 0;
        i_13_4533 <= 0;
        i_13_4534 <= 0;
        i_13_4535 <= 0;
        i_13_4536 <= 0;
        i_13_4537 <= 0;
        i_13_4538 <= 0;
        i_13_4539 <= 0;
        i_13_4540 <= 0;
        i_13_4541 <= 0;
        i_13_4542 <= 0;
        i_13_4543 <= 0;
        i_13_4544 <= 0;
        i_13_4545 <= 0;
        i_13_4546 <= 0;
        i_13_4547 <= 0;
        i_13_4548 <= 0;
        i_13_4549 <= 0;
        i_13_4550 <= 0;
        i_13_4551 <= 0;
        i_13_4552 <= 0;
        i_13_4553 <= 0;
        i_13_4554 <= 0;
        i_13_4555 <= 0;
        i_13_4556 <= 0;
        i_13_4557 <= 0;
        i_13_4558 <= 0;
        i_13_4559 <= 0;
        i_13_4560 <= 0;
        i_13_4561 <= 0;
        i_13_4562 <= 0;
        i_13_4563 <= 0;
        i_13_4564 <= 0;
        i_13_4565 <= 0;
        i_13_4566 <= 0;
        i_13_4567 <= 0;
        i_13_4568 <= 0;
        i_13_4569 <= 0;
        i_13_4570 <= 0;
        i_13_4571 <= 0;
        i_13_4572 <= 0;
        i_13_4573 <= 0;
        i_13_4574 <= 0;
        i_13_4575 <= 0;
        i_13_4576 <= 0;
        i_13_4577 <= 0;
        i_13_4578 <= 0;
        i_13_4579 <= 0;
        i_13_4580 <= 0;
        i_13_4581 <= 0;
        i_13_4582 <= 0;
        i_13_4583 <= 0;
        i_13_4584 <= 0;
        i_13_4585 <= 0;
        i_13_4586 <= 0;
        i_13_4587 <= 0;
        i_13_4588 <= 0;
        i_13_4589 <= 0;
        i_13_4590 <= 0;
        i_13_4591 <= 0;
        i_13_4592 <= 0;
        i_13_4593 <= 0;
        i_13_4594 <= 0;
        i_13_4595 <= 0;
        i_13_4596 <= 0;
        i_13_4597 <= 0;
        i_13_4598 <= 0;
        i_13_4599 <= 0;
        i_13_4600 <= 0;
        i_13_4601 <= 0;
        i_13_4602 <= 0;
        i_13_4603 <= 0;
        i_13_4604 <= 0;
        i_13_4605 <= 0;
        i_13_4606 <= 0;
        i_13_4607 <= 0;
        dly1 <= 0;
        dly2 <= 0;
      end
    else if (ce)
      begin
        out_reg <= { o_13_511, o_13_510, o_13_509, o_13_508, o_13_507, o_13_506, o_13_505, o_13_504, o_13_503, o_13_502, o_13_501, o_13_500, o_13_499, o_13_498, o_13_497, o_13_496, o_13_495, o_13_494, o_13_493, o_13_492, o_13_491, o_13_490, o_13_489, o_13_488, o_13_487, o_13_486, o_13_485, o_13_484, o_13_483, o_13_482, o_13_481, o_13_480, o_13_479, o_13_478, o_13_477, o_13_476, o_13_475, o_13_474, o_13_473, o_13_472, o_13_471, o_13_470, o_13_469, o_13_468, o_13_467, o_13_466, o_13_465, o_13_464, o_13_463, o_13_462, o_13_461, o_13_460, o_13_459, o_13_458, o_13_457, o_13_456, o_13_455, o_13_454, o_13_453, o_13_452, o_13_451, o_13_450, o_13_449, o_13_448, o_13_447, o_13_446, o_13_445, o_13_444, o_13_443, o_13_442, o_13_441, o_13_440, o_13_439, o_13_438, o_13_437, o_13_436, o_13_435, o_13_434, o_13_433, o_13_432, o_13_431, o_13_430, o_13_429, o_13_428, o_13_427, o_13_426, o_13_425, o_13_424, o_13_423, o_13_422, o_13_421, o_13_420, o_13_419, o_13_418, o_13_417, o_13_416, o_13_415, o_13_414, o_13_413, o_13_412, o_13_411, o_13_410, o_13_409, o_13_408, o_13_407, o_13_406, o_13_405, o_13_404, o_13_403, o_13_402, o_13_401, o_13_400, o_13_399, o_13_398, o_13_397, o_13_396, o_13_395, o_13_394, o_13_393, o_13_392, o_13_391, o_13_390, o_13_389, o_13_388, o_13_387, o_13_386, o_13_385, o_13_384, o_13_383, o_13_382, o_13_381, o_13_380, o_13_379, o_13_378, o_13_377, o_13_376, o_13_375, o_13_374, o_13_373, o_13_372, o_13_371, o_13_370, o_13_369, o_13_368, o_13_367, o_13_366, o_13_365, o_13_364, o_13_363, o_13_362, o_13_361, o_13_360, o_13_359, o_13_358, o_13_357, o_13_356, o_13_355, o_13_354, o_13_353, o_13_352, o_13_351, o_13_350, o_13_349, o_13_348, o_13_347, o_13_346, o_13_345, o_13_344, o_13_343, o_13_342, o_13_341, o_13_340, o_13_339, o_13_338, o_13_337, o_13_336, o_13_335, o_13_334, o_13_333, o_13_332, o_13_331, o_13_330, o_13_329, o_13_328, o_13_327, o_13_326, o_13_325, o_13_324, o_13_323, o_13_322, o_13_321, o_13_320, o_13_319, o_13_318, o_13_317, o_13_316, o_13_315, o_13_314, o_13_313, o_13_312, o_13_311, o_13_310, o_13_309, o_13_308, o_13_307, o_13_306, o_13_305, o_13_304, o_13_303, o_13_302, o_13_301, o_13_300, o_13_299, o_13_298, o_13_297, o_13_296, o_13_295, o_13_294, o_13_293, o_13_292, o_13_291, o_13_290, o_13_289, o_13_288, o_13_287, o_13_286, o_13_285, o_13_284, o_13_283, o_13_282, o_13_281, o_13_280, o_13_279, o_13_278, o_13_277, o_13_276, o_13_275, o_13_274, o_13_273, o_13_272, o_13_271, o_13_270, o_13_269, o_13_268, o_13_267, o_13_266, o_13_265, o_13_264, o_13_263, o_13_262, o_13_261, o_13_260, o_13_259, o_13_258, o_13_257, o_13_256, o_13_255, o_13_254, o_13_253, o_13_252, o_13_251, o_13_250, o_13_249, o_13_248, o_13_247, o_13_246, o_13_245, o_13_244, o_13_243, o_13_242, o_13_241, o_13_240, o_13_239, o_13_238, o_13_237, o_13_236, o_13_235, o_13_234, o_13_233, o_13_232, o_13_231, o_13_230, o_13_229, o_13_228, o_13_227, o_13_226, o_13_225, o_13_224, o_13_223, o_13_222, o_13_221, o_13_220, o_13_219, o_13_218, o_13_217, o_13_216, o_13_215, o_13_214, o_13_213, o_13_212, o_13_211, o_13_210, o_13_209, o_13_208, o_13_207, o_13_206, o_13_205, o_13_204, o_13_203, o_13_202, o_13_201, o_13_200, o_13_199, o_13_198, o_13_197, o_13_196, o_13_195, o_13_194, o_13_193, o_13_192, o_13_191, o_13_190, o_13_189, o_13_188, o_13_187, o_13_186, o_13_185, o_13_184, o_13_183, o_13_182, o_13_181, o_13_180, o_13_179, o_13_178, o_13_177, o_13_176, o_13_175, o_13_174, o_13_173, o_13_172, o_13_171, o_13_170, o_13_169, o_13_168, o_13_167, o_13_166, o_13_165, o_13_164, o_13_163, o_13_162, o_13_161, o_13_160, o_13_159, o_13_158, o_13_157, o_13_156, o_13_155, o_13_154, o_13_153, o_13_152, o_13_151, o_13_150, o_13_149, o_13_148, o_13_147, o_13_146, o_13_145, o_13_144, o_13_143, o_13_142, o_13_141, o_13_140, o_13_139, o_13_138, o_13_137, o_13_136, o_13_135, o_13_134, o_13_133, o_13_132, o_13_131, o_13_130, o_13_129, o_13_128, o_13_127, o_13_126, o_13_125, o_13_124, o_13_123, o_13_122, o_13_121, o_13_120, o_13_119, o_13_118, o_13_117, o_13_116, o_13_115, o_13_114, o_13_113, o_13_112, o_13_111, o_13_110, o_13_109, o_13_108, o_13_107, o_13_106, o_13_105, o_13_104, o_13_103, o_13_102, o_13_101, o_13_100, o_13_99, o_13_98, o_13_97, o_13_96, o_13_95, o_13_94, o_13_93, o_13_92, o_13_91, o_13_90, o_13_89, o_13_88, o_13_87, o_13_86, o_13_85, o_13_84, o_13_83, o_13_82, o_13_81, o_13_80, o_13_79, o_13_78, o_13_77, o_13_76, o_13_75, o_13_74, o_13_73, o_13_72, o_13_71, o_13_70, o_13_69, o_13_68, o_13_67, o_13_66, o_13_65, o_13_64, o_13_63, o_13_62, o_13_61, o_13_60, o_13_59, o_13_58, o_13_57, o_13_56, o_13_55, o_13_54, o_13_53, o_13_52, o_13_51, o_13_50, o_13_49, o_13_48, o_13_47, o_13_46, o_13_45, o_13_44, o_13_43, o_13_42, o_13_41, o_13_40, o_13_39, o_13_38, o_13_37, o_13_36, o_13_35, o_13_34, o_13_33, o_13_32, o_13_31, o_13_30, o_13_29, o_13_28, o_13_27, o_13_26, o_13_25, o_13_24, o_13_23, o_13_22, o_13_21, o_13_20, o_13_19, o_13_18, o_13_17, o_13_16, o_13_15, o_13_14, o_13_13, o_13_12, o_13_11, o_13_10, o_13_9, o_13_8, o_13_7, o_13_6, o_13_5, o_13_4, o_13_3, o_13_2, o_13_1, o_13_0};
        i_13_0 <= in_reg[0];
        i_13_1 <= in_reg[512];
        i_13_2 <= in_reg[1024];
        i_13_3 <= in_reg[1536];
        i_13_4 <= in_reg[2048];
        i_13_5 <= in_reg[2560];
        i_13_6 <= in_reg[3072];
        i_13_7 <= in_reg[3584];
        i_13_8 <= in_reg[4096];
        i_13_9 <= in_reg[1];
        i_13_10 <= in_reg[513];
        i_13_11 <= in_reg[1025];
        i_13_12 <= in_reg[1537];
        i_13_13 <= in_reg[2049];
        i_13_14 <= in_reg[2561];
        i_13_15 <= in_reg[3073];
        i_13_16 <= in_reg[3585];
        i_13_17 <= in_reg[4097];
        i_13_18 <= in_reg[2];
        i_13_19 <= in_reg[514];
        i_13_20 <= in_reg[1026];
        i_13_21 <= in_reg[1538];
        i_13_22 <= in_reg[2050];
        i_13_23 <= in_reg[2562];
        i_13_24 <= in_reg[3074];
        i_13_25 <= in_reg[3586];
        i_13_26 <= in_reg[4098];
        i_13_27 <= in_reg[3];
        i_13_28 <= in_reg[515];
        i_13_29 <= in_reg[1027];
        i_13_30 <= in_reg[1539];
        i_13_31 <= in_reg[2051];
        i_13_32 <= in_reg[2563];
        i_13_33 <= in_reg[3075];
        i_13_34 <= in_reg[3587];
        i_13_35 <= in_reg[4099];
        i_13_36 <= in_reg[4];
        i_13_37 <= in_reg[516];
        i_13_38 <= in_reg[1028];
        i_13_39 <= in_reg[1540];
        i_13_40 <= in_reg[2052];
        i_13_41 <= in_reg[2564];
        i_13_42 <= in_reg[3076];
        i_13_43 <= in_reg[3588];
        i_13_44 <= in_reg[4100];
        i_13_45 <= in_reg[5];
        i_13_46 <= in_reg[517];
        i_13_47 <= in_reg[1029];
        i_13_48 <= in_reg[1541];
        i_13_49 <= in_reg[2053];
        i_13_50 <= in_reg[2565];
        i_13_51 <= in_reg[3077];
        i_13_52 <= in_reg[3589];
        i_13_53 <= in_reg[4101];
        i_13_54 <= in_reg[6];
        i_13_55 <= in_reg[518];
        i_13_56 <= in_reg[1030];
        i_13_57 <= in_reg[1542];
        i_13_58 <= in_reg[2054];
        i_13_59 <= in_reg[2566];
        i_13_60 <= in_reg[3078];
        i_13_61 <= in_reg[3590];
        i_13_62 <= in_reg[4102];
        i_13_63 <= in_reg[7];
        i_13_64 <= in_reg[519];
        i_13_65 <= in_reg[1031];
        i_13_66 <= in_reg[1543];
        i_13_67 <= in_reg[2055];
        i_13_68 <= in_reg[2567];
        i_13_69 <= in_reg[3079];
        i_13_70 <= in_reg[3591];
        i_13_71 <= in_reg[4103];
        i_13_72 <= in_reg[8];
        i_13_73 <= in_reg[520];
        i_13_74 <= in_reg[1032];
        i_13_75 <= in_reg[1544];
        i_13_76 <= in_reg[2056];
        i_13_77 <= in_reg[2568];
        i_13_78 <= in_reg[3080];
        i_13_79 <= in_reg[3592];
        i_13_80 <= in_reg[4104];
        i_13_81 <= in_reg[9];
        i_13_82 <= in_reg[521];
        i_13_83 <= in_reg[1033];
        i_13_84 <= in_reg[1545];
        i_13_85 <= in_reg[2057];
        i_13_86 <= in_reg[2569];
        i_13_87 <= in_reg[3081];
        i_13_88 <= in_reg[3593];
        i_13_89 <= in_reg[4105];
        i_13_90 <= in_reg[10];
        i_13_91 <= in_reg[522];
        i_13_92 <= in_reg[1034];
        i_13_93 <= in_reg[1546];
        i_13_94 <= in_reg[2058];
        i_13_95 <= in_reg[2570];
        i_13_96 <= in_reg[3082];
        i_13_97 <= in_reg[3594];
        i_13_98 <= in_reg[4106];
        i_13_99 <= in_reg[11];
        i_13_100 <= in_reg[523];
        i_13_101 <= in_reg[1035];
        i_13_102 <= in_reg[1547];
        i_13_103 <= in_reg[2059];
        i_13_104 <= in_reg[2571];
        i_13_105 <= in_reg[3083];
        i_13_106 <= in_reg[3595];
        i_13_107 <= in_reg[4107];
        i_13_108 <= in_reg[12];
        i_13_109 <= in_reg[524];
        i_13_110 <= in_reg[1036];
        i_13_111 <= in_reg[1548];
        i_13_112 <= in_reg[2060];
        i_13_113 <= in_reg[2572];
        i_13_114 <= in_reg[3084];
        i_13_115 <= in_reg[3596];
        i_13_116 <= in_reg[4108];
        i_13_117 <= in_reg[13];
        i_13_118 <= in_reg[525];
        i_13_119 <= in_reg[1037];
        i_13_120 <= in_reg[1549];
        i_13_121 <= in_reg[2061];
        i_13_122 <= in_reg[2573];
        i_13_123 <= in_reg[3085];
        i_13_124 <= in_reg[3597];
        i_13_125 <= in_reg[4109];
        i_13_126 <= in_reg[14];
        i_13_127 <= in_reg[526];
        i_13_128 <= in_reg[1038];
        i_13_129 <= in_reg[1550];
        i_13_130 <= in_reg[2062];
        i_13_131 <= in_reg[2574];
        i_13_132 <= in_reg[3086];
        i_13_133 <= in_reg[3598];
        i_13_134 <= in_reg[4110];
        i_13_135 <= in_reg[15];
        i_13_136 <= in_reg[527];
        i_13_137 <= in_reg[1039];
        i_13_138 <= in_reg[1551];
        i_13_139 <= in_reg[2063];
        i_13_140 <= in_reg[2575];
        i_13_141 <= in_reg[3087];
        i_13_142 <= in_reg[3599];
        i_13_143 <= in_reg[4111];
        i_13_144 <= in_reg[16];
        i_13_145 <= in_reg[528];
        i_13_146 <= in_reg[1040];
        i_13_147 <= in_reg[1552];
        i_13_148 <= in_reg[2064];
        i_13_149 <= in_reg[2576];
        i_13_150 <= in_reg[3088];
        i_13_151 <= in_reg[3600];
        i_13_152 <= in_reg[4112];
        i_13_153 <= in_reg[17];
        i_13_154 <= in_reg[529];
        i_13_155 <= in_reg[1041];
        i_13_156 <= in_reg[1553];
        i_13_157 <= in_reg[2065];
        i_13_158 <= in_reg[2577];
        i_13_159 <= in_reg[3089];
        i_13_160 <= in_reg[3601];
        i_13_161 <= in_reg[4113];
        i_13_162 <= in_reg[18];
        i_13_163 <= in_reg[530];
        i_13_164 <= in_reg[1042];
        i_13_165 <= in_reg[1554];
        i_13_166 <= in_reg[2066];
        i_13_167 <= in_reg[2578];
        i_13_168 <= in_reg[3090];
        i_13_169 <= in_reg[3602];
        i_13_170 <= in_reg[4114];
        i_13_171 <= in_reg[19];
        i_13_172 <= in_reg[531];
        i_13_173 <= in_reg[1043];
        i_13_174 <= in_reg[1555];
        i_13_175 <= in_reg[2067];
        i_13_176 <= in_reg[2579];
        i_13_177 <= in_reg[3091];
        i_13_178 <= in_reg[3603];
        i_13_179 <= in_reg[4115];
        i_13_180 <= in_reg[20];
        i_13_181 <= in_reg[532];
        i_13_182 <= in_reg[1044];
        i_13_183 <= in_reg[1556];
        i_13_184 <= in_reg[2068];
        i_13_185 <= in_reg[2580];
        i_13_186 <= in_reg[3092];
        i_13_187 <= in_reg[3604];
        i_13_188 <= in_reg[4116];
        i_13_189 <= in_reg[21];
        i_13_190 <= in_reg[533];
        i_13_191 <= in_reg[1045];
        i_13_192 <= in_reg[1557];
        i_13_193 <= in_reg[2069];
        i_13_194 <= in_reg[2581];
        i_13_195 <= in_reg[3093];
        i_13_196 <= in_reg[3605];
        i_13_197 <= in_reg[4117];
        i_13_198 <= in_reg[22];
        i_13_199 <= in_reg[534];
        i_13_200 <= in_reg[1046];
        i_13_201 <= in_reg[1558];
        i_13_202 <= in_reg[2070];
        i_13_203 <= in_reg[2582];
        i_13_204 <= in_reg[3094];
        i_13_205 <= in_reg[3606];
        i_13_206 <= in_reg[4118];
        i_13_207 <= in_reg[23];
        i_13_208 <= in_reg[535];
        i_13_209 <= in_reg[1047];
        i_13_210 <= in_reg[1559];
        i_13_211 <= in_reg[2071];
        i_13_212 <= in_reg[2583];
        i_13_213 <= in_reg[3095];
        i_13_214 <= in_reg[3607];
        i_13_215 <= in_reg[4119];
        i_13_216 <= in_reg[24];
        i_13_217 <= in_reg[536];
        i_13_218 <= in_reg[1048];
        i_13_219 <= in_reg[1560];
        i_13_220 <= in_reg[2072];
        i_13_221 <= in_reg[2584];
        i_13_222 <= in_reg[3096];
        i_13_223 <= in_reg[3608];
        i_13_224 <= in_reg[4120];
        i_13_225 <= in_reg[25];
        i_13_226 <= in_reg[537];
        i_13_227 <= in_reg[1049];
        i_13_228 <= in_reg[1561];
        i_13_229 <= in_reg[2073];
        i_13_230 <= in_reg[2585];
        i_13_231 <= in_reg[3097];
        i_13_232 <= in_reg[3609];
        i_13_233 <= in_reg[4121];
        i_13_234 <= in_reg[26];
        i_13_235 <= in_reg[538];
        i_13_236 <= in_reg[1050];
        i_13_237 <= in_reg[1562];
        i_13_238 <= in_reg[2074];
        i_13_239 <= in_reg[2586];
        i_13_240 <= in_reg[3098];
        i_13_241 <= in_reg[3610];
        i_13_242 <= in_reg[4122];
        i_13_243 <= in_reg[27];
        i_13_244 <= in_reg[539];
        i_13_245 <= in_reg[1051];
        i_13_246 <= in_reg[1563];
        i_13_247 <= in_reg[2075];
        i_13_248 <= in_reg[2587];
        i_13_249 <= in_reg[3099];
        i_13_250 <= in_reg[3611];
        i_13_251 <= in_reg[4123];
        i_13_252 <= in_reg[28];
        i_13_253 <= in_reg[540];
        i_13_254 <= in_reg[1052];
        i_13_255 <= in_reg[1564];
        i_13_256 <= in_reg[2076];
        i_13_257 <= in_reg[2588];
        i_13_258 <= in_reg[3100];
        i_13_259 <= in_reg[3612];
        i_13_260 <= in_reg[4124];
        i_13_261 <= in_reg[29];
        i_13_262 <= in_reg[541];
        i_13_263 <= in_reg[1053];
        i_13_264 <= in_reg[1565];
        i_13_265 <= in_reg[2077];
        i_13_266 <= in_reg[2589];
        i_13_267 <= in_reg[3101];
        i_13_268 <= in_reg[3613];
        i_13_269 <= in_reg[4125];
        i_13_270 <= in_reg[30];
        i_13_271 <= in_reg[542];
        i_13_272 <= in_reg[1054];
        i_13_273 <= in_reg[1566];
        i_13_274 <= in_reg[2078];
        i_13_275 <= in_reg[2590];
        i_13_276 <= in_reg[3102];
        i_13_277 <= in_reg[3614];
        i_13_278 <= in_reg[4126];
        i_13_279 <= in_reg[31];
        i_13_280 <= in_reg[543];
        i_13_281 <= in_reg[1055];
        i_13_282 <= in_reg[1567];
        i_13_283 <= in_reg[2079];
        i_13_284 <= in_reg[2591];
        i_13_285 <= in_reg[3103];
        i_13_286 <= in_reg[3615];
        i_13_287 <= in_reg[4127];
        i_13_288 <= in_reg[32];
        i_13_289 <= in_reg[544];
        i_13_290 <= in_reg[1056];
        i_13_291 <= in_reg[1568];
        i_13_292 <= in_reg[2080];
        i_13_293 <= in_reg[2592];
        i_13_294 <= in_reg[3104];
        i_13_295 <= in_reg[3616];
        i_13_296 <= in_reg[4128];
        i_13_297 <= in_reg[33];
        i_13_298 <= in_reg[545];
        i_13_299 <= in_reg[1057];
        i_13_300 <= in_reg[1569];
        i_13_301 <= in_reg[2081];
        i_13_302 <= in_reg[2593];
        i_13_303 <= in_reg[3105];
        i_13_304 <= in_reg[3617];
        i_13_305 <= in_reg[4129];
        i_13_306 <= in_reg[34];
        i_13_307 <= in_reg[546];
        i_13_308 <= in_reg[1058];
        i_13_309 <= in_reg[1570];
        i_13_310 <= in_reg[2082];
        i_13_311 <= in_reg[2594];
        i_13_312 <= in_reg[3106];
        i_13_313 <= in_reg[3618];
        i_13_314 <= in_reg[4130];
        i_13_315 <= in_reg[35];
        i_13_316 <= in_reg[547];
        i_13_317 <= in_reg[1059];
        i_13_318 <= in_reg[1571];
        i_13_319 <= in_reg[2083];
        i_13_320 <= in_reg[2595];
        i_13_321 <= in_reg[3107];
        i_13_322 <= in_reg[3619];
        i_13_323 <= in_reg[4131];
        i_13_324 <= in_reg[36];
        i_13_325 <= in_reg[548];
        i_13_326 <= in_reg[1060];
        i_13_327 <= in_reg[1572];
        i_13_328 <= in_reg[2084];
        i_13_329 <= in_reg[2596];
        i_13_330 <= in_reg[3108];
        i_13_331 <= in_reg[3620];
        i_13_332 <= in_reg[4132];
        i_13_333 <= in_reg[37];
        i_13_334 <= in_reg[549];
        i_13_335 <= in_reg[1061];
        i_13_336 <= in_reg[1573];
        i_13_337 <= in_reg[2085];
        i_13_338 <= in_reg[2597];
        i_13_339 <= in_reg[3109];
        i_13_340 <= in_reg[3621];
        i_13_341 <= in_reg[4133];
        i_13_342 <= in_reg[38];
        i_13_343 <= in_reg[550];
        i_13_344 <= in_reg[1062];
        i_13_345 <= in_reg[1574];
        i_13_346 <= in_reg[2086];
        i_13_347 <= in_reg[2598];
        i_13_348 <= in_reg[3110];
        i_13_349 <= in_reg[3622];
        i_13_350 <= in_reg[4134];
        i_13_351 <= in_reg[39];
        i_13_352 <= in_reg[551];
        i_13_353 <= in_reg[1063];
        i_13_354 <= in_reg[1575];
        i_13_355 <= in_reg[2087];
        i_13_356 <= in_reg[2599];
        i_13_357 <= in_reg[3111];
        i_13_358 <= in_reg[3623];
        i_13_359 <= in_reg[4135];
        i_13_360 <= in_reg[40];
        i_13_361 <= in_reg[552];
        i_13_362 <= in_reg[1064];
        i_13_363 <= in_reg[1576];
        i_13_364 <= in_reg[2088];
        i_13_365 <= in_reg[2600];
        i_13_366 <= in_reg[3112];
        i_13_367 <= in_reg[3624];
        i_13_368 <= in_reg[4136];
        i_13_369 <= in_reg[41];
        i_13_370 <= in_reg[553];
        i_13_371 <= in_reg[1065];
        i_13_372 <= in_reg[1577];
        i_13_373 <= in_reg[2089];
        i_13_374 <= in_reg[2601];
        i_13_375 <= in_reg[3113];
        i_13_376 <= in_reg[3625];
        i_13_377 <= in_reg[4137];
        i_13_378 <= in_reg[42];
        i_13_379 <= in_reg[554];
        i_13_380 <= in_reg[1066];
        i_13_381 <= in_reg[1578];
        i_13_382 <= in_reg[2090];
        i_13_383 <= in_reg[2602];
        i_13_384 <= in_reg[3114];
        i_13_385 <= in_reg[3626];
        i_13_386 <= in_reg[4138];
        i_13_387 <= in_reg[43];
        i_13_388 <= in_reg[555];
        i_13_389 <= in_reg[1067];
        i_13_390 <= in_reg[1579];
        i_13_391 <= in_reg[2091];
        i_13_392 <= in_reg[2603];
        i_13_393 <= in_reg[3115];
        i_13_394 <= in_reg[3627];
        i_13_395 <= in_reg[4139];
        i_13_396 <= in_reg[44];
        i_13_397 <= in_reg[556];
        i_13_398 <= in_reg[1068];
        i_13_399 <= in_reg[1580];
        i_13_400 <= in_reg[2092];
        i_13_401 <= in_reg[2604];
        i_13_402 <= in_reg[3116];
        i_13_403 <= in_reg[3628];
        i_13_404 <= in_reg[4140];
        i_13_405 <= in_reg[45];
        i_13_406 <= in_reg[557];
        i_13_407 <= in_reg[1069];
        i_13_408 <= in_reg[1581];
        i_13_409 <= in_reg[2093];
        i_13_410 <= in_reg[2605];
        i_13_411 <= in_reg[3117];
        i_13_412 <= in_reg[3629];
        i_13_413 <= in_reg[4141];
        i_13_414 <= in_reg[46];
        i_13_415 <= in_reg[558];
        i_13_416 <= in_reg[1070];
        i_13_417 <= in_reg[1582];
        i_13_418 <= in_reg[2094];
        i_13_419 <= in_reg[2606];
        i_13_420 <= in_reg[3118];
        i_13_421 <= in_reg[3630];
        i_13_422 <= in_reg[4142];
        i_13_423 <= in_reg[47];
        i_13_424 <= in_reg[559];
        i_13_425 <= in_reg[1071];
        i_13_426 <= in_reg[1583];
        i_13_427 <= in_reg[2095];
        i_13_428 <= in_reg[2607];
        i_13_429 <= in_reg[3119];
        i_13_430 <= in_reg[3631];
        i_13_431 <= in_reg[4143];
        i_13_432 <= in_reg[48];
        i_13_433 <= in_reg[560];
        i_13_434 <= in_reg[1072];
        i_13_435 <= in_reg[1584];
        i_13_436 <= in_reg[2096];
        i_13_437 <= in_reg[2608];
        i_13_438 <= in_reg[3120];
        i_13_439 <= in_reg[3632];
        i_13_440 <= in_reg[4144];
        i_13_441 <= in_reg[49];
        i_13_442 <= in_reg[561];
        i_13_443 <= in_reg[1073];
        i_13_444 <= in_reg[1585];
        i_13_445 <= in_reg[2097];
        i_13_446 <= in_reg[2609];
        i_13_447 <= in_reg[3121];
        i_13_448 <= in_reg[3633];
        i_13_449 <= in_reg[4145];
        i_13_450 <= in_reg[50];
        i_13_451 <= in_reg[562];
        i_13_452 <= in_reg[1074];
        i_13_453 <= in_reg[1586];
        i_13_454 <= in_reg[2098];
        i_13_455 <= in_reg[2610];
        i_13_456 <= in_reg[3122];
        i_13_457 <= in_reg[3634];
        i_13_458 <= in_reg[4146];
        i_13_459 <= in_reg[51];
        i_13_460 <= in_reg[563];
        i_13_461 <= in_reg[1075];
        i_13_462 <= in_reg[1587];
        i_13_463 <= in_reg[2099];
        i_13_464 <= in_reg[2611];
        i_13_465 <= in_reg[3123];
        i_13_466 <= in_reg[3635];
        i_13_467 <= in_reg[4147];
        i_13_468 <= in_reg[52];
        i_13_469 <= in_reg[564];
        i_13_470 <= in_reg[1076];
        i_13_471 <= in_reg[1588];
        i_13_472 <= in_reg[2100];
        i_13_473 <= in_reg[2612];
        i_13_474 <= in_reg[3124];
        i_13_475 <= in_reg[3636];
        i_13_476 <= in_reg[4148];
        i_13_477 <= in_reg[53];
        i_13_478 <= in_reg[565];
        i_13_479 <= in_reg[1077];
        i_13_480 <= in_reg[1589];
        i_13_481 <= in_reg[2101];
        i_13_482 <= in_reg[2613];
        i_13_483 <= in_reg[3125];
        i_13_484 <= in_reg[3637];
        i_13_485 <= in_reg[4149];
        i_13_486 <= in_reg[54];
        i_13_487 <= in_reg[566];
        i_13_488 <= in_reg[1078];
        i_13_489 <= in_reg[1590];
        i_13_490 <= in_reg[2102];
        i_13_491 <= in_reg[2614];
        i_13_492 <= in_reg[3126];
        i_13_493 <= in_reg[3638];
        i_13_494 <= in_reg[4150];
        i_13_495 <= in_reg[55];
        i_13_496 <= in_reg[567];
        i_13_497 <= in_reg[1079];
        i_13_498 <= in_reg[1591];
        i_13_499 <= in_reg[2103];
        i_13_500 <= in_reg[2615];
        i_13_501 <= in_reg[3127];
        i_13_502 <= in_reg[3639];
        i_13_503 <= in_reg[4151];
        i_13_504 <= in_reg[56];
        i_13_505 <= in_reg[568];
        i_13_506 <= in_reg[1080];
        i_13_507 <= in_reg[1592];
        i_13_508 <= in_reg[2104];
        i_13_509 <= in_reg[2616];
        i_13_510 <= in_reg[3128];
        i_13_511 <= in_reg[3640];
        i_13_512 <= in_reg[4152];
        i_13_513 <= in_reg[57];
        i_13_514 <= in_reg[569];
        i_13_515 <= in_reg[1081];
        i_13_516 <= in_reg[1593];
        i_13_517 <= in_reg[2105];
        i_13_518 <= in_reg[2617];
        i_13_519 <= in_reg[3129];
        i_13_520 <= in_reg[3641];
        i_13_521 <= in_reg[4153];
        i_13_522 <= in_reg[58];
        i_13_523 <= in_reg[570];
        i_13_524 <= in_reg[1082];
        i_13_525 <= in_reg[1594];
        i_13_526 <= in_reg[2106];
        i_13_527 <= in_reg[2618];
        i_13_528 <= in_reg[3130];
        i_13_529 <= in_reg[3642];
        i_13_530 <= in_reg[4154];
        i_13_531 <= in_reg[59];
        i_13_532 <= in_reg[571];
        i_13_533 <= in_reg[1083];
        i_13_534 <= in_reg[1595];
        i_13_535 <= in_reg[2107];
        i_13_536 <= in_reg[2619];
        i_13_537 <= in_reg[3131];
        i_13_538 <= in_reg[3643];
        i_13_539 <= in_reg[4155];
        i_13_540 <= in_reg[60];
        i_13_541 <= in_reg[572];
        i_13_542 <= in_reg[1084];
        i_13_543 <= in_reg[1596];
        i_13_544 <= in_reg[2108];
        i_13_545 <= in_reg[2620];
        i_13_546 <= in_reg[3132];
        i_13_547 <= in_reg[3644];
        i_13_548 <= in_reg[4156];
        i_13_549 <= in_reg[61];
        i_13_550 <= in_reg[573];
        i_13_551 <= in_reg[1085];
        i_13_552 <= in_reg[1597];
        i_13_553 <= in_reg[2109];
        i_13_554 <= in_reg[2621];
        i_13_555 <= in_reg[3133];
        i_13_556 <= in_reg[3645];
        i_13_557 <= in_reg[4157];
        i_13_558 <= in_reg[62];
        i_13_559 <= in_reg[574];
        i_13_560 <= in_reg[1086];
        i_13_561 <= in_reg[1598];
        i_13_562 <= in_reg[2110];
        i_13_563 <= in_reg[2622];
        i_13_564 <= in_reg[3134];
        i_13_565 <= in_reg[3646];
        i_13_566 <= in_reg[4158];
        i_13_567 <= in_reg[63];
        i_13_568 <= in_reg[575];
        i_13_569 <= in_reg[1087];
        i_13_570 <= in_reg[1599];
        i_13_571 <= in_reg[2111];
        i_13_572 <= in_reg[2623];
        i_13_573 <= in_reg[3135];
        i_13_574 <= in_reg[3647];
        i_13_575 <= in_reg[4159];
        i_13_576 <= in_reg[64];
        i_13_577 <= in_reg[576];
        i_13_578 <= in_reg[1088];
        i_13_579 <= in_reg[1600];
        i_13_580 <= in_reg[2112];
        i_13_581 <= in_reg[2624];
        i_13_582 <= in_reg[3136];
        i_13_583 <= in_reg[3648];
        i_13_584 <= in_reg[4160];
        i_13_585 <= in_reg[65];
        i_13_586 <= in_reg[577];
        i_13_587 <= in_reg[1089];
        i_13_588 <= in_reg[1601];
        i_13_589 <= in_reg[2113];
        i_13_590 <= in_reg[2625];
        i_13_591 <= in_reg[3137];
        i_13_592 <= in_reg[3649];
        i_13_593 <= in_reg[4161];
        i_13_594 <= in_reg[66];
        i_13_595 <= in_reg[578];
        i_13_596 <= in_reg[1090];
        i_13_597 <= in_reg[1602];
        i_13_598 <= in_reg[2114];
        i_13_599 <= in_reg[2626];
        i_13_600 <= in_reg[3138];
        i_13_601 <= in_reg[3650];
        i_13_602 <= in_reg[4162];
        i_13_603 <= in_reg[67];
        i_13_604 <= in_reg[579];
        i_13_605 <= in_reg[1091];
        i_13_606 <= in_reg[1603];
        i_13_607 <= in_reg[2115];
        i_13_608 <= in_reg[2627];
        i_13_609 <= in_reg[3139];
        i_13_610 <= in_reg[3651];
        i_13_611 <= in_reg[4163];
        i_13_612 <= in_reg[68];
        i_13_613 <= in_reg[580];
        i_13_614 <= in_reg[1092];
        i_13_615 <= in_reg[1604];
        i_13_616 <= in_reg[2116];
        i_13_617 <= in_reg[2628];
        i_13_618 <= in_reg[3140];
        i_13_619 <= in_reg[3652];
        i_13_620 <= in_reg[4164];
        i_13_621 <= in_reg[69];
        i_13_622 <= in_reg[581];
        i_13_623 <= in_reg[1093];
        i_13_624 <= in_reg[1605];
        i_13_625 <= in_reg[2117];
        i_13_626 <= in_reg[2629];
        i_13_627 <= in_reg[3141];
        i_13_628 <= in_reg[3653];
        i_13_629 <= in_reg[4165];
        i_13_630 <= in_reg[70];
        i_13_631 <= in_reg[582];
        i_13_632 <= in_reg[1094];
        i_13_633 <= in_reg[1606];
        i_13_634 <= in_reg[2118];
        i_13_635 <= in_reg[2630];
        i_13_636 <= in_reg[3142];
        i_13_637 <= in_reg[3654];
        i_13_638 <= in_reg[4166];
        i_13_639 <= in_reg[71];
        i_13_640 <= in_reg[583];
        i_13_641 <= in_reg[1095];
        i_13_642 <= in_reg[1607];
        i_13_643 <= in_reg[2119];
        i_13_644 <= in_reg[2631];
        i_13_645 <= in_reg[3143];
        i_13_646 <= in_reg[3655];
        i_13_647 <= in_reg[4167];
        i_13_648 <= in_reg[72];
        i_13_649 <= in_reg[584];
        i_13_650 <= in_reg[1096];
        i_13_651 <= in_reg[1608];
        i_13_652 <= in_reg[2120];
        i_13_653 <= in_reg[2632];
        i_13_654 <= in_reg[3144];
        i_13_655 <= in_reg[3656];
        i_13_656 <= in_reg[4168];
        i_13_657 <= in_reg[73];
        i_13_658 <= in_reg[585];
        i_13_659 <= in_reg[1097];
        i_13_660 <= in_reg[1609];
        i_13_661 <= in_reg[2121];
        i_13_662 <= in_reg[2633];
        i_13_663 <= in_reg[3145];
        i_13_664 <= in_reg[3657];
        i_13_665 <= in_reg[4169];
        i_13_666 <= in_reg[74];
        i_13_667 <= in_reg[586];
        i_13_668 <= in_reg[1098];
        i_13_669 <= in_reg[1610];
        i_13_670 <= in_reg[2122];
        i_13_671 <= in_reg[2634];
        i_13_672 <= in_reg[3146];
        i_13_673 <= in_reg[3658];
        i_13_674 <= in_reg[4170];
        i_13_675 <= in_reg[75];
        i_13_676 <= in_reg[587];
        i_13_677 <= in_reg[1099];
        i_13_678 <= in_reg[1611];
        i_13_679 <= in_reg[2123];
        i_13_680 <= in_reg[2635];
        i_13_681 <= in_reg[3147];
        i_13_682 <= in_reg[3659];
        i_13_683 <= in_reg[4171];
        i_13_684 <= in_reg[76];
        i_13_685 <= in_reg[588];
        i_13_686 <= in_reg[1100];
        i_13_687 <= in_reg[1612];
        i_13_688 <= in_reg[2124];
        i_13_689 <= in_reg[2636];
        i_13_690 <= in_reg[3148];
        i_13_691 <= in_reg[3660];
        i_13_692 <= in_reg[4172];
        i_13_693 <= in_reg[77];
        i_13_694 <= in_reg[589];
        i_13_695 <= in_reg[1101];
        i_13_696 <= in_reg[1613];
        i_13_697 <= in_reg[2125];
        i_13_698 <= in_reg[2637];
        i_13_699 <= in_reg[3149];
        i_13_700 <= in_reg[3661];
        i_13_701 <= in_reg[4173];
        i_13_702 <= in_reg[78];
        i_13_703 <= in_reg[590];
        i_13_704 <= in_reg[1102];
        i_13_705 <= in_reg[1614];
        i_13_706 <= in_reg[2126];
        i_13_707 <= in_reg[2638];
        i_13_708 <= in_reg[3150];
        i_13_709 <= in_reg[3662];
        i_13_710 <= in_reg[4174];
        i_13_711 <= in_reg[79];
        i_13_712 <= in_reg[591];
        i_13_713 <= in_reg[1103];
        i_13_714 <= in_reg[1615];
        i_13_715 <= in_reg[2127];
        i_13_716 <= in_reg[2639];
        i_13_717 <= in_reg[3151];
        i_13_718 <= in_reg[3663];
        i_13_719 <= in_reg[4175];
        i_13_720 <= in_reg[80];
        i_13_721 <= in_reg[592];
        i_13_722 <= in_reg[1104];
        i_13_723 <= in_reg[1616];
        i_13_724 <= in_reg[2128];
        i_13_725 <= in_reg[2640];
        i_13_726 <= in_reg[3152];
        i_13_727 <= in_reg[3664];
        i_13_728 <= in_reg[4176];
        i_13_729 <= in_reg[81];
        i_13_730 <= in_reg[593];
        i_13_731 <= in_reg[1105];
        i_13_732 <= in_reg[1617];
        i_13_733 <= in_reg[2129];
        i_13_734 <= in_reg[2641];
        i_13_735 <= in_reg[3153];
        i_13_736 <= in_reg[3665];
        i_13_737 <= in_reg[4177];
        i_13_738 <= in_reg[82];
        i_13_739 <= in_reg[594];
        i_13_740 <= in_reg[1106];
        i_13_741 <= in_reg[1618];
        i_13_742 <= in_reg[2130];
        i_13_743 <= in_reg[2642];
        i_13_744 <= in_reg[3154];
        i_13_745 <= in_reg[3666];
        i_13_746 <= in_reg[4178];
        i_13_747 <= in_reg[83];
        i_13_748 <= in_reg[595];
        i_13_749 <= in_reg[1107];
        i_13_750 <= in_reg[1619];
        i_13_751 <= in_reg[2131];
        i_13_752 <= in_reg[2643];
        i_13_753 <= in_reg[3155];
        i_13_754 <= in_reg[3667];
        i_13_755 <= in_reg[4179];
        i_13_756 <= in_reg[84];
        i_13_757 <= in_reg[596];
        i_13_758 <= in_reg[1108];
        i_13_759 <= in_reg[1620];
        i_13_760 <= in_reg[2132];
        i_13_761 <= in_reg[2644];
        i_13_762 <= in_reg[3156];
        i_13_763 <= in_reg[3668];
        i_13_764 <= in_reg[4180];
        i_13_765 <= in_reg[85];
        i_13_766 <= in_reg[597];
        i_13_767 <= in_reg[1109];
        i_13_768 <= in_reg[1621];
        i_13_769 <= in_reg[2133];
        i_13_770 <= in_reg[2645];
        i_13_771 <= in_reg[3157];
        i_13_772 <= in_reg[3669];
        i_13_773 <= in_reg[4181];
        i_13_774 <= in_reg[86];
        i_13_775 <= in_reg[598];
        i_13_776 <= in_reg[1110];
        i_13_777 <= in_reg[1622];
        i_13_778 <= in_reg[2134];
        i_13_779 <= in_reg[2646];
        i_13_780 <= in_reg[3158];
        i_13_781 <= in_reg[3670];
        i_13_782 <= in_reg[4182];
        i_13_783 <= in_reg[87];
        i_13_784 <= in_reg[599];
        i_13_785 <= in_reg[1111];
        i_13_786 <= in_reg[1623];
        i_13_787 <= in_reg[2135];
        i_13_788 <= in_reg[2647];
        i_13_789 <= in_reg[3159];
        i_13_790 <= in_reg[3671];
        i_13_791 <= in_reg[4183];
        i_13_792 <= in_reg[88];
        i_13_793 <= in_reg[600];
        i_13_794 <= in_reg[1112];
        i_13_795 <= in_reg[1624];
        i_13_796 <= in_reg[2136];
        i_13_797 <= in_reg[2648];
        i_13_798 <= in_reg[3160];
        i_13_799 <= in_reg[3672];
        i_13_800 <= in_reg[4184];
        i_13_801 <= in_reg[89];
        i_13_802 <= in_reg[601];
        i_13_803 <= in_reg[1113];
        i_13_804 <= in_reg[1625];
        i_13_805 <= in_reg[2137];
        i_13_806 <= in_reg[2649];
        i_13_807 <= in_reg[3161];
        i_13_808 <= in_reg[3673];
        i_13_809 <= in_reg[4185];
        i_13_810 <= in_reg[90];
        i_13_811 <= in_reg[602];
        i_13_812 <= in_reg[1114];
        i_13_813 <= in_reg[1626];
        i_13_814 <= in_reg[2138];
        i_13_815 <= in_reg[2650];
        i_13_816 <= in_reg[3162];
        i_13_817 <= in_reg[3674];
        i_13_818 <= in_reg[4186];
        i_13_819 <= in_reg[91];
        i_13_820 <= in_reg[603];
        i_13_821 <= in_reg[1115];
        i_13_822 <= in_reg[1627];
        i_13_823 <= in_reg[2139];
        i_13_824 <= in_reg[2651];
        i_13_825 <= in_reg[3163];
        i_13_826 <= in_reg[3675];
        i_13_827 <= in_reg[4187];
        i_13_828 <= in_reg[92];
        i_13_829 <= in_reg[604];
        i_13_830 <= in_reg[1116];
        i_13_831 <= in_reg[1628];
        i_13_832 <= in_reg[2140];
        i_13_833 <= in_reg[2652];
        i_13_834 <= in_reg[3164];
        i_13_835 <= in_reg[3676];
        i_13_836 <= in_reg[4188];
        i_13_837 <= in_reg[93];
        i_13_838 <= in_reg[605];
        i_13_839 <= in_reg[1117];
        i_13_840 <= in_reg[1629];
        i_13_841 <= in_reg[2141];
        i_13_842 <= in_reg[2653];
        i_13_843 <= in_reg[3165];
        i_13_844 <= in_reg[3677];
        i_13_845 <= in_reg[4189];
        i_13_846 <= in_reg[94];
        i_13_847 <= in_reg[606];
        i_13_848 <= in_reg[1118];
        i_13_849 <= in_reg[1630];
        i_13_850 <= in_reg[2142];
        i_13_851 <= in_reg[2654];
        i_13_852 <= in_reg[3166];
        i_13_853 <= in_reg[3678];
        i_13_854 <= in_reg[4190];
        i_13_855 <= in_reg[95];
        i_13_856 <= in_reg[607];
        i_13_857 <= in_reg[1119];
        i_13_858 <= in_reg[1631];
        i_13_859 <= in_reg[2143];
        i_13_860 <= in_reg[2655];
        i_13_861 <= in_reg[3167];
        i_13_862 <= in_reg[3679];
        i_13_863 <= in_reg[4191];
        i_13_864 <= in_reg[96];
        i_13_865 <= in_reg[608];
        i_13_866 <= in_reg[1120];
        i_13_867 <= in_reg[1632];
        i_13_868 <= in_reg[2144];
        i_13_869 <= in_reg[2656];
        i_13_870 <= in_reg[3168];
        i_13_871 <= in_reg[3680];
        i_13_872 <= in_reg[4192];
        i_13_873 <= in_reg[97];
        i_13_874 <= in_reg[609];
        i_13_875 <= in_reg[1121];
        i_13_876 <= in_reg[1633];
        i_13_877 <= in_reg[2145];
        i_13_878 <= in_reg[2657];
        i_13_879 <= in_reg[3169];
        i_13_880 <= in_reg[3681];
        i_13_881 <= in_reg[4193];
        i_13_882 <= in_reg[98];
        i_13_883 <= in_reg[610];
        i_13_884 <= in_reg[1122];
        i_13_885 <= in_reg[1634];
        i_13_886 <= in_reg[2146];
        i_13_887 <= in_reg[2658];
        i_13_888 <= in_reg[3170];
        i_13_889 <= in_reg[3682];
        i_13_890 <= in_reg[4194];
        i_13_891 <= in_reg[99];
        i_13_892 <= in_reg[611];
        i_13_893 <= in_reg[1123];
        i_13_894 <= in_reg[1635];
        i_13_895 <= in_reg[2147];
        i_13_896 <= in_reg[2659];
        i_13_897 <= in_reg[3171];
        i_13_898 <= in_reg[3683];
        i_13_899 <= in_reg[4195];
        i_13_900 <= in_reg[100];
        i_13_901 <= in_reg[612];
        i_13_902 <= in_reg[1124];
        i_13_903 <= in_reg[1636];
        i_13_904 <= in_reg[2148];
        i_13_905 <= in_reg[2660];
        i_13_906 <= in_reg[3172];
        i_13_907 <= in_reg[3684];
        i_13_908 <= in_reg[4196];
        i_13_909 <= in_reg[101];
        i_13_910 <= in_reg[613];
        i_13_911 <= in_reg[1125];
        i_13_912 <= in_reg[1637];
        i_13_913 <= in_reg[2149];
        i_13_914 <= in_reg[2661];
        i_13_915 <= in_reg[3173];
        i_13_916 <= in_reg[3685];
        i_13_917 <= in_reg[4197];
        i_13_918 <= in_reg[102];
        i_13_919 <= in_reg[614];
        i_13_920 <= in_reg[1126];
        i_13_921 <= in_reg[1638];
        i_13_922 <= in_reg[2150];
        i_13_923 <= in_reg[2662];
        i_13_924 <= in_reg[3174];
        i_13_925 <= in_reg[3686];
        i_13_926 <= in_reg[4198];
        i_13_927 <= in_reg[103];
        i_13_928 <= in_reg[615];
        i_13_929 <= in_reg[1127];
        i_13_930 <= in_reg[1639];
        i_13_931 <= in_reg[2151];
        i_13_932 <= in_reg[2663];
        i_13_933 <= in_reg[3175];
        i_13_934 <= in_reg[3687];
        i_13_935 <= in_reg[4199];
        i_13_936 <= in_reg[104];
        i_13_937 <= in_reg[616];
        i_13_938 <= in_reg[1128];
        i_13_939 <= in_reg[1640];
        i_13_940 <= in_reg[2152];
        i_13_941 <= in_reg[2664];
        i_13_942 <= in_reg[3176];
        i_13_943 <= in_reg[3688];
        i_13_944 <= in_reg[4200];
        i_13_945 <= in_reg[105];
        i_13_946 <= in_reg[617];
        i_13_947 <= in_reg[1129];
        i_13_948 <= in_reg[1641];
        i_13_949 <= in_reg[2153];
        i_13_950 <= in_reg[2665];
        i_13_951 <= in_reg[3177];
        i_13_952 <= in_reg[3689];
        i_13_953 <= in_reg[4201];
        i_13_954 <= in_reg[106];
        i_13_955 <= in_reg[618];
        i_13_956 <= in_reg[1130];
        i_13_957 <= in_reg[1642];
        i_13_958 <= in_reg[2154];
        i_13_959 <= in_reg[2666];
        i_13_960 <= in_reg[3178];
        i_13_961 <= in_reg[3690];
        i_13_962 <= in_reg[4202];
        i_13_963 <= in_reg[107];
        i_13_964 <= in_reg[619];
        i_13_965 <= in_reg[1131];
        i_13_966 <= in_reg[1643];
        i_13_967 <= in_reg[2155];
        i_13_968 <= in_reg[2667];
        i_13_969 <= in_reg[3179];
        i_13_970 <= in_reg[3691];
        i_13_971 <= in_reg[4203];
        i_13_972 <= in_reg[108];
        i_13_973 <= in_reg[620];
        i_13_974 <= in_reg[1132];
        i_13_975 <= in_reg[1644];
        i_13_976 <= in_reg[2156];
        i_13_977 <= in_reg[2668];
        i_13_978 <= in_reg[3180];
        i_13_979 <= in_reg[3692];
        i_13_980 <= in_reg[4204];
        i_13_981 <= in_reg[109];
        i_13_982 <= in_reg[621];
        i_13_983 <= in_reg[1133];
        i_13_984 <= in_reg[1645];
        i_13_985 <= in_reg[2157];
        i_13_986 <= in_reg[2669];
        i_13_987 <= in_reg[3181];
        i_13_988 <= in_reg[3693];
        i_13_989 <= in_reg[4205];
        i_13_990 <= in_reg[110];
        i_13_991 <= in_reg[622];
        i_13_992 <= in_reg[1134];
        i_13_993 <= in_reg[1646];
        i_13_994 <= in_reg[2158];
        i_13_995 <= in_reg[2670];
        i_13_996 <= in_reg[3182];
        i_13_997 <= in_reg[3694];
        i_13_998 <= in_reg[4206];
        i_13_999 <= in_reg[111];
        i_13_1000 <= in_reg[623];
        i_13_1001 <= in_reg[1135];
        i_13_1002 <= in_reg[1647];
        i_13_1003 <= in_reg[2159];
        i_13_1004 <= in_reg[2671];
        i_13_1005 <= in_reg[3183];
        i_13_1006 <= in_reg[3695];
        i_13_1007 <= in_reg[4207];
        i_13_1008 <= in_reg[112];
        i_13_1009 <= in_reg[624];
        i_13_1010 <= in_reg[1136];
        i_13_1011 <= in_reg[1648];
        i_13_1012 <= in_reg[2160];
        i_13_1013 <= in_reg[2672];
        i_13_1014 <= in_reg[3184];
        i_13_1015 <= in_reg[3696];
        i_13_1016 <= in_reg[4208];
        i_13_1017 <= in_reg[113];
        i_13_1018 <= in_reg[625];
        i_13_1019 <= in_reg[1137];
        i_13_1020 <= in_reg[1649];
        i_13_1021 <= in_reg[2161];
        i_13_1022 <= in_reg[2673];
        i_13_1023 <= in_reg[3185];
        i_13_1024 <= in_reg[3697];
        i_13_1025 <= in_reg[4209];
        i_13_1026 <= in_reg[114];
        i_13_1027 <= in_reg[626];
        i_13_1028 <= in_reg[1138];
        i_13_1029 <= in_reg[1650];
        i_13_1030 <= in_reg[2162];
        i_13_1031 <= in_reg[2674];
        i_13_1032 <= in_reg[3186];
        i_13_1033 <= in_reg[3698];
        i_13_1034 <= in_reg[4210];
        i_13_1035 <= in_reg[115];
        i_13_1036 <= in_reg[627];
        i_13_1037 <= in_reg[1139];
        i_13_1038 <= in_reg[1651];
        i_13_1039 <= in_reg[2163];
        i_13_1040 <= in_reg[2675];
        i_13_1041 <= in_reg[3187];
        i_13_1042 <= in_reg[3699];
        i_13_1043 <= in_reg[4211];
        i_13_1044 <= in_reg[116];
        i_13_1045 <= in_reg[628];
        i_13_1046 <= in_reg[1140];
        i_13_1047 <= in_reg[1652];
        i_13_1048 <= in_reg[2164];
        i_13_1049 <= in_reg[2676];
        i_13_1050 <= in_reg[3188];
        i_13_1051 <= in_reg[3700];
        i_13_1052 <= in_reg[4212];
        i_13_1053 <= in_reg[117];
        i_13_1054 <= in_reg[629];
        i_13_1055 <= in_reg[1141];
        i_13_1056 <= in_reg[1653];
        i_13_1057 <= in_reg[2165];
        i_13_1058 <= in_reg[2677];
        i_13_1059 <= in_reg[3189];
        i_13_1060 <= in_reg[3701];
        i_13_1061 <= in_reg[4213];
        i_13_1062 <= in_reg[118];
        i_13_1063 <= in_reg[630];
        i_13_1064 <= in_reg[1142];
        i_13_1065 <= in_reg[1654];
        i_13_1066 <= in_reg[2166];
        i_13_1067 <= in_reg[2678];
        i_13_1068 <= in_reg[3190];
        i_13_1069 <= in_reg[3702];
        i_13_1070 <= in_reg[4214];
        i_13_1071 <= in_reg[119];
        i_13_1072 <= in_reg[631];
        i_13_1073 <= in_reg[1143];
        i_13_1074 <= in_reg[1655];
        i_13_1075 <= in_reg[2167];
        i_13_1076 <= in_reg[2679];
        i_13_1077 <= in_reg[3191];
        i_13_1078 <= in_reg[3703];
        i_13_1079 <= in_reg[4215];
        i_13_1080 <= in_reg[120];
        i_13_1081 <= in_reg[632];
        i_13_1082 <= in_reg[1144];
        i_13_1083 <= in_reg[1656];
        i_13_1084 <= in_reg[2168];
        i_13_1085 <= in_reg[2680];
        i_13_1086 <= in_reg[3192];
        i_13_1087 <= in_reg[3704];
        i_13_1088 <= in_reg[4216];
        i_13_1089 <= in_reg[121];
        i_13_1090 <= in_reg[633];
        i_13_1091 <= in_reg[1145];
        i_13_1092 <= in_reg[1657];
        i_13_1093 <= in_reg[2169];
        i_13_1094 <= in_reg[2681];
        i_13_1095 <= in_reg[3193];
        i_13_1096 <= in_reg[3705];
        i_13_1097 <= in_reg[4217];
        i_13_1098 <= in_reg[122];
        i_13_1099 <= in_reg[634];
        i_13_1100 <= in_reg[1146];
        i_13_1101 <= in_reg[1658];
        i_13_1102 <= in_reg[2170];
        i_13_1103 <= in_reg[2682];
        i_13_1104 <= in_reg[3194];
        i_13_1105 <= in_reg[3706];
        i_13_1106 <= in_reg[4218];
        i_13_1107 <= in_reg[123];
        i_13_1108 <= in_reg[635];
        i_13_1109 <= in_reg[1147];
        i_13_1110 <= in_reg[1659];
        i_13_1111 <= in_reg[2171];
        i_13_1112 <= in_reg[2683];
        i_13_1113 <= in_reg[3195];
        i_13_1114 <= in_reg[3707];
        i_13_1115 <= in_reg[4219];
        i_13_1116 <= in_reg[124];
        i_13_1117 <= in_reg[636];
        i_13_1118 <= in_reg[1148];
        i_13_1119 <= in_reg[1660];
        i_13_1120 <= in_reg[2172];
        i_13_1121 <= in_reg[2684];
        i_13_1122 <= in_reg[3196];
        i_13_1123 <= in_reg[3708];
        i_13_1124 <= in_reg[4220];
        i_13_1125 <= in_reg[125];
        i_13_1126 <= in_reg[637];
        i_13_1127 <= in_reg[1149];
        i_13_1128 <= in_reg[1661];
        i_13_1129 <= in_reg[2173];
        i_13_1130 <= in_reg[2685];
        i_13_1131 <= in_reg[3197];
        i_13_1132 <= in_reg[3709];
        i_13_1133 <= in_reg[4221];
        i_13_1134 <= in_reg[126];
        i_13_1135 <= in_reg[638];
        i_13_1136 <= in_reg[1150];
        i_13_1137 <= in_reg[1662];
        i_13_1138 <= in_reg[2174];
        i_13_1139 <= in_reg[2686];
        i_13_1140 <= in_reg[3198];
        i_13_1141 <= in_reg[3710];
        i_13_1142 <= in_reg[4222];
        i_13_1143 <= in_reg[127];
        i_13_1144 <= in_reg[639];
        i_13_1145 <= in_reg[1151];
        i_13_1146 <= in_reg[1663];
        i_13_1147 <= in_reg[2175];
        i_13_1148 <= in_reg[2687];
        i_13_1149 <= in_reg[3199];
        i_13_1150 <= in_reg[3711];
        i_13_1151 <= in_reg[4223];
        i_13_1152 <= in_reg[128];
        i_13_1153 <= in_reg[640];
        i_13_1154 <= in_reg[1152];
        i_13_1155 <= in_reg[1664];
        i_13_1156 <= in_reg[2176];
        i_13_1157 <= in_reg[2688];
        i_13_1158 <= in_reg[3200];
        i_13_1159 <= in_reg[3712];
        i_13_1160 <= in_reg[4224];
        i_13_1161 <= in_reg[129];
        i_13_1162 <= in_reg[641];
        i_13_1163 <= in_reg[1153];
        i_13_1164 <= in_reg[1665];
        i_13_1165 <= in_reg[2177];
        i_13_1166 <= in_reg[2689];
        i_13_1167 <= in_reg[3201];
        i_13_1168 <= in_reg[3713];
        i_13_1169 <= in_reg[4225];
        i_13_1170 <= in_reg[130];
        i_13_1171 <= in_reg[642];
        i_13_1172 <= in_reg[1154];
        i_13_1173 <= in_reg[1666];
        i_13_1174 <= in_reg[2178];
        i_13_1175 <= in_reg[2690];
        i_13_1176 <= in_reg[3202];
        i_13_1177 <= in_reg[3714];
        i_13_1178 <= in_reg[4226];
        i_13_1179 <= in_reg[131];
        i_13_1180 <= in_reg[643];
        i_13_1181 <= in_reg[1155];
        i_13_1182 <= in_reg[1667];
        i_13_1183 <= in_reg[2179];
        i_13_1184 <= in_reg[2691];
        i_13_1185 <= in_reg[3203];
        i_13_1186 <= in_reg[3715];
        i_13_1187 <= in_reg[4227];
        i_13_1188 <= in_reg[132];
        i_13_1189 <= in_reg[644];
        i_13_1190 <= in_reg[1156];
        i_13_1191 <= in_reg[1668];
        i_13_1192 <= in_reg[2180];
        i_13_1193 <= in_reg[2692];
        i_13_1194 <= in_reg[3204];
        i_13_1195 <= in_reg[3716];
        i_13_1196 <= in_reg[4228];
        i_13_1197 <= in_reg[133];
        i_13_1198 <= in_reg[645];
        i_13_1199 <= in_reg[1157];
        i_13_1200 <= in_reg[1669];
        i_13_1201 <= in_reg[2181];
        i_13_1202 <= in_reg[2693];
        i_13_1203 <= in_reg[3205];
        i_13_1204 <= in_reg[3717];
        i_13_1205 <= in_reg[4229];
        i_13_1206 <= in_reg[134];
        i_13_1207 <= in_reg[646];
        i_13_1208 <= in_reg[1158];
        i_13_1209 <= in_reg[1670];
        i_13_1210 <= in_reg[2182];
        i_13_1211 <= in_reg[2694];
        i_13_1212 <= in_reg[3206];
        i_13_1213 <= in_reg[3718];
        i_13_1214 <= in_reg[4230];
        i_13_1215 <= in_reg[135];
        i_13_1216 <= in_reg[647];
        i_13_1217 <= in_reg[1159];
        i_13_1218 <= in_reg[1671];
        i_13_1219 <= in_reg[2183];
        i_13_1220 <= in_reg[2695];
        i_13_1221 <= in_reg[3207];
        i_13_1222 <= in_reg[3719];
        i_13_1223 <= in_reg[4231];
        i_13_1224 <= in_reg[136];
        i_13_1225 <= in_reg[648];
        i_13_1226 <= in_reg[1160];
        i_13_1227 <= in_reg[1672];
        i_13_1228 <= in_reg[2184];
        i_13_1229 <= in_reg[2696];
        i_13_1230 <= in_reg[3208];
        i_13_1231 <= in_reg[3720];
        i_13_1232 <= in_reg[4232];
        i_13_1233 <= in_reg[137];
        i_13_1234 <= in_reg[649];
        i_13_1235 <= in_reg[1161];
        i_13_1236 <= in_reg[1673];
        i_13_1237 <= in_reg[2185];
        i_13_1238 <= in_reg[2697];
        i_13_1239 <= in_reg[3209];
        i_13_1240 <= in_reg[3721];
        i_13_1241 <= in_reg[4233];
        i_13_1242 <= in_reg[138];
        i_13_1243 <= in_reg[650];
        i_13_1244 <= in_reg[1162];
        i_13_1245 <= in_reg[1674];
        i_13_1246 <= in_reg[2186];
        i_13_1247 <= in_reg[2698];
        i_13_1248 <= in_reg[3210];
        i_13_1249 <= in_reg[3722];
        i_13_1250 <= in_reg[4234];
        i_13_1251 <= in_reg[139];
        i_13_1252 <= in_reg[651];
        i_13_1253 <= in_reg[1163];
        i_13_1254 <= in_reg[1675];
        i_13_1255 <= in_reg[2187];
        i_13_1256 <= in_reg[2699];
        i_13_1257 <= in_reg[3211];
        i_13_1258 <= in_reg[3723];
        i_13_1259 <= in_reg[4235];
        i_13_1260 <= in_reg[140];
        i_13_1261 <= in_reg[652];
        i_13_1262 <= in_reg[1164];
        i_13_1263 <= in_reg[1676];
        i_13_1264 <= in_reg[2188];
        i_13_1265 <= in_reg[2700];
        i_13_1266 <= in_reg[3212];
        i_13_1267 <= in_reg[3724];
        i_13_1268 <= in_reg[4236];
        i_13_1269 <= in_reg[141];
        i_13_1270 <= in_reg[653];
        i_13_1271 <= in_reg[1165];
        i_13_1272 <= in_reg[1677];
        i_13_1273 <= in_reg[2189];
        i_13_1274 <= in_reg[2701];
        i_13_1275 <= in_reg[3213];
        i_13_1276 <= in_reg[3725];
        i_13_1277 <= in_reg[4237];
        i_13_1278 <= in_reg[142];
        i_13_1279 <= in_reg[654];
        i_13_1280 <= in_reg[1166];
        i_13_1281 <= in_reg[1678];
        i_13_1282 <= in_reg[2190];
        i_13_1283 <= in_reg[2702];
        i_13_1284 <= in_reg[3214];
        i_13_1285 <= in_reg[3726];
        i_13_1286 <= in_reg[4238];
        i_13_1287 <= in_reg[143];
        i_13_1288 <= in_reg[655];
        i_13_1289 <= in_reg[1167];
        i_13_1290 <= in_reg[1679];
        i_13_1291 <= in_reg[2191];
        i_13_1292 <= in_reg[2703];
        i_13_1293 <= in_reg[3215];
        i_13_1294 <= in_reg[3727];
        i_13_1295 <= in_reg[4239];
        i_13_1296 <= in_reg[144];
        i_13_1297 <= in_reg[656];
        i_13_1298 <= in_reg[1168];
        i_13_1299 <= in_reg[1680];
        i_13_1300 <= in_reg[2192];
        i_13_1301 <= in_reg[2704];
        i_13_1302 <= in_reg[3216];
        i_13_1303 <= in_reg[3728];
        i_13_1304 <= in_reg[4240];
        i_13_1305 <= in_reg[145];
        i_13_1306 <= in_reg[657];
        i_13_1307 <= in_reg[1169];
        i_13_1308 <= in_reg[1681];
        i_13_1309 <= in_reg[2193];
        i_13_1310 <= in_reg[2705];
        i_13_1311 <= in_reg[3217];
        i_13_1312 <= in_reg[3729];
        i_13_1313 <= in_reg[4241];
        i_13_1314 <= in_reg[146];
        i_13_1315 <= in_reg[658];
        i_13_1316 <= in_reg[1170];
        i_13_1317 <= in_reg[1682];
        i_13_1318 <= in_reg[2194];
        i_13_1319 <= in_reg[2706];
        i_13_1320 <= in_reg[3218];
        i_13_1321 <= in_reg[3730];
        i_13_1322 <= in_reg[4242];
        i_13_1323 <= in_reg[147];
        i_13_1324 <= in_reg[659];
        i_13_1325 <= in_reg[1171];
        i_13_1326 <= in_reg[1683];
        i_13_1327 <= in_reg[2195];
        i_13_1328 <= in_reg[2707];
        i_13_1329 <= in_reg[3219];
        i_13_1330 <= in_reg[3731];
        i_13_1331 <= in_reg[4243];
        i_13_1332 <= in_reg[148];
        i_13_1333 <= in_reg[660];
        i_13_1334 <= in_reg[1172];
        i_13_1335 <= in_reg[1684];
        i_13_1336 <= in_reg[2196];
        i_13_1337 <= in_reg[2708];
        i_13_1338 <= in_reg[3220];
        i_13_1339 <= in_reg[3732];
        i_13_1340 <= in_reg[4244];
        i_13_1341 <= in_reg[149];
        i_13_1342 <= in_reg[661];
        i_13_1343 <= in_reg[1173];
        i_13_1344 <= in_reg[1685];
        i_13_1345 <= in_reg[2197];
        i_13_1346 <= in_reg[2709];
        i_13_1347 <= in_reg[3221];
        i_13_1348 <= in_reg[3733];
        i_13_1349 <= in_reg[4245];
        i_13_1350 <= in_reg[150];
        i_13_1351 <= in_reg[662];
        i_13_1352 <= in_reg[1174];
        i_13_1353 <= in_reg[1686];
        i_13_1354 <= in_reg[2198];
        i_13_1355 <= in_reg[2710];
        i_13_1356 <= in_reg[3222];
        i_13_1357 <= in_reg[3734];
        i_13_1358 <= in_reg[4246];
        i_13_1359 <= in_reg[151];
        i_13_1360 <= in_reg[663];
        i_13_1361 <= in_reg[1175];
        i_13_1362 <= in_reg[1687];
        i_13_1363 <= in_reg[2199];
        i_13_1364 <= in_reg[2711];
        i_13_1365 <= in_reg[3223];
        i_13_1366 <= in_reg[3735];
        i_13_1367 <= in_reg[4247];
        i_13_1368 <= in_reg[152];
        i_13_1369 <= in_reg[664];
        i_13_1370 <= in_reg[1176];
        i_13_1371 <= in_reg[1688];
        i_13_1372 <= in_reg[2200];
        i_13_1373 <= in_reg[2712];
        i_13_1374 <= in_reg[3224];
        i_13_1375 <= in_reg[3736];
        i_13_1376 <= in_reg[4248];
        i_13_1377 <= in_reg[153];
        i_13_1378 <= in_reg[665];
        i_13_1379 <= in_reg[1177];
        i_13_1380 <= in_reg[1689];
        i_13_1381 <= in_reg[2201];
        i_13_1382 <= in_reg[2713];
        i_13_1383 <= in_reg[3225];
        i_13_1384 <= in_reg[3737];
        i_13_1385 <= in_reg[4249];
        i_13_1386 <= in_reg[154];
        i_13_1387 <= in_reg[666];
        i_13_1388 <= in_reg[1178];
        i_13_1389 <= in_reg[1690];
        i_13_1390 <= in_reg[2202];
        i_13_1391 <= in_reg[2714];
        i_13_1392 <= in_reg[3226];
        i_13_1393 <= in_reg[3738];
        i_13_1394 <= in_reg[4250];
        i_13_1395 <= in_reg[155];
        i_13_1396 <= in_reg[667];
        i_13_1397 <= in_reg[1179];
        i_13_1398 <= in_reg[1691];
        i_13_1399 <= in_reg[2203];
        i_13_1400 <= in_reg[2715];
        i_13_1401 <= in_reg[3227];
        i_13_1402 <= in_reg[3739];
        i_13_1403 <= in_reg[4251];
        i_13_1404 <= in_reg[156];
        i_13_1405 <= in_reg[668];
        i_13_1406 <= in_reg[1180];
        i_13_1407 <= in_reg[1692];
        i_13_1408 <= in_reg[2204];
        i_13_1409 <= in_reg[2716];
        i_13_1410 <= in_reg[3228];
        i_13_1411 <= in_reg[3740];
        i_13_1412 <= in_reg[4252];
        i_13_1413 <= in_reg[157];
        i_13_1414 <= in_reg[669];
        i_13_1415 <= in_reg[1181];
        i_13_1416 <= in_reg[1693];
        i_13_1417 <= in_reg[2205];
        i_13_1418 <= in_reg[2717];
        i_13_1419 <= in_reg[3229];
        i_13_1420 <= in_reg[3741];
        i_13_1421 <= in_reg[4253];
        i_13_1422 <= in_reg[158];
        i_13_1423 <= in_reg[670];
        i_13_1424 <= in_reg[1182];
        i_13_1425 <= in_reg[1694];
        i_13_1426 <= in_reg[2206];
        i_13_1427 <= in_reg[2718];
        i_13_1428 <= in_reg[3230];
        i_13_1429 <= in_reg[3742];
        i_13_1430 <= in_reg[4254];
        i_13_1431 <= in_reg[159];
        i_13_1432 <= in_reg[671];
        i_13_1433 <= in_reg[1183];
        i_13_1434 <= in_reg[1695];
        i_13_1435 <= in_reg[2207];
        i_13_1436 <= in_reg[2719];
        i_13_1437 <= in_reg[3231];
        i_13_1438 <= in_reg[3743];
        i_13_1439 <= in_reg[4255];
        i_13_1440 <= in_reg[160];
        i_13_1441 <= in_reg[672];
        i_13_1442 <= in_reg[1184];
        i_13_1443 <= in_reg[1696];
        i_13_1444 <= in_reg[2208];
        i_13_1445 <= in_reg[2720];
        i_13_1446 <= in_reg[3232];
        i_13_1447 <= in_reg[3744];
        i_13_1448 <= in_reg[4256];
        i_13_1449 <= in_reg[161];
        i_13_1450 <= in_reg[673];
        i_13_1451 <= in_reg[1185];
        i_13_1452 <= in_reg[1697];
        i_13_1453 <= in_reg[2209];
        i_13_1454 <= in_reg[2721];
        i_13_1455 <= in_reg[3233];
        i_13_1456 <= in_reg[3745];
        i_13_1457 <= in_reg[4257];
        i_13_1458 <= in_reg[162];
        i_13_1459 <= in_reg[674];
        i_13_1460 <= in_reg[1186];
        i_13_1461 <= in_reg[1698];
        i_13_1462 <= in_reg[2210];
        i_13_1463 <= in_reg[2722];
        i_13_1464 <= in_reg[3234];
        i_13_1465 <= in_reg[3746];
        i_13_1466 <= in_reg[4258];
        i_13_1467 <= in_reg[163];
        i_13_1468 <= in_reg[675];
        i_13_1469 <= in_reg[1187];
        i_13_1470 <= in_reg[1699];
        i_13_1471 <= in_reg[2211];
        i_13_1472 <= in_reg[2723];
        i_13_1473 <= in_reg[3235];
        i_13_1474 <= in_reg[3747];
        i_13_1475 <= in_reg[4259];
        i_13_1476 <= in_reg[164];
        i_13_1477 <= in_reg[676];
        i_13_1478 <= in_reg[1188];
        i_13_1479 <= in_reg[1700];
        i_13_1480 <= in_reg[2212];
        i_13_1481 <= in_reg[2724];
        i_13_1482 <= in_reg[3236];
        i_13_1483 <= in_reg[3748];
        i_13_1484 <= in_reg[4260];
        i_13_1485 <= in_reg[165];
        i_13_1486 <= in_reg[677];
        i_13_1487 <= in_reg[1189];
        i_13_1488 <= in_reg[1701];
        i_13_1489 <= in_reg[2213];
        i_13_1490 <= in_reg[2725];
        i_13_1491 <= in_reg[3237];
        i_13_1492 <= in_reg[3749];
        i_13_1493 <= in_reg[4261];
        i_13_1494 <= in_reg[166];
        i_13_1495 <= in_reg[678];
        i_13_1496 <= in_reg[1190];
        i_13_1497 <= in_reg[1702];
        i_13_1498 <= in_reg[2214];
        i_13_1499 <= in_reg[2726];
        i_13_1500 <= in_reg[3238];
        i_13_1501 <= in_reg[3750];
        i_13_1502 <= in_reg[4262];
        i_13_1503 <= in_reg[167];
        i_13_1504 <= in_reg[679];
        i_13_1505 <= in_reg[1191];
        i_13_1506 <= in_reg[1703];
        i_13_1507 <= in_reg[2215];
        i_13_1508 <= in_reg[2727];
        i_13_1509 <= in_reg[3239];
        i_13_1510 <= in_reg[3751];
        i_13_1511 <= in_reg[4263];
        i_13_1512 <= in_reg[168];
        i_13_1513 <= in_reg[680];
        i_13_1514 <= in_reg[1192];
        i_13_1515 <= in_reg[1704];
        i_13_1516 <= in_reg[2216];
        i_13_1517 <= in_reg[2728];
        i_13_1518 <= in_reg[3240];
        i_13_1519 <= in_reg[3752];
        i_13_1520 <= in_reg[4264];
        i_13_1521 <= in_reg[169];
        i_13_1522 <= in_reg[681];
        i_13_1523 <= in_reg[1193];
        i_13_1524 <= in_reg[1705];
        i_13_1525 <= in_reg[2217];
        i_13_1526 <= in_reg[2729];
        i_13_1527 <= in_reg[3241];
        i_13_1528 <= in_reg[3753];
        i_13_1529 <= in_reg[4265];
        i_13_1530 <= in_reg[170];
        i_13_1531 <= in_reg[682];
        i_13_1532 <= in_reg[1194];
        i_13_1533 <= in_reg[1706];
        i_13_1534 <= in_reg[2218];
        i_13_1535 <= in_reg[2730];
        i_13_1536 <= in_reg[3242];
        i_13_1537 <= in_reg[3754];
        i_13_1538 <= in_reg[4266];
        i_13_1539 <= in_reg[171];
        i_13_1540 <= in_reg[683];
        i_13_1541 <= in_reg[1195];
        i_13_1542 <= in_reg[1707];
        i_13_1543 <= in_reg[2219];
        i_13_1544 <= in_reg[2731];
        i_13_1545 <= in_reg[3243];
        i_13_1546 <= in_reg[3755];
        i_13_1547 <= in_reg[4267];
        i_13_1548 <= in_reg[172];
        i_13_1549 <= in_reg[684];
        i_13_1550 <= in_reg[1196];
        i_13_1551 <= in_reg[1708];
        i_13_1552 <= in_reg[2220];
        i_13_1553 <= in_reg[2732];
        i_13_1554 <= in_reg[3244];
        i_13_1555 <= in_reg[3756];
        i_13_1556 <= in_reg[4268];
        i_13_1557 <= in_reg[173];
        i_13_1558 <= in_reg[685];
        i_13_1559 <= in_reg[1197];
        i_13_1560 <= in_reg[1709];
        i_13_1561 <= in_reg[2221];
        i_13_1562 <= in_reg[2733];
        i_13_1563 <= in_reg[3245];
        i_13_1564 <= in_reg[3757];
        i_13_1565 <= in_reg[4269];
        i_13_1566 <= in_reg[174];
        i_13_1567 <= in_reg[686];
        i_13_1568 <= in_reg[1198];
        i_13_1569 <= in_reg[1710];
        i_13_1570 <= in_reg[2222];
        i_13_1571 <= in_reg[2734];
        i_13_1572 <= in_reg[3246];
        i_13_1573 <= in_reg[3758];
        i_13_1574 <= in_reg[4270];
        i_13_1575 <= in_reg[175];
        i_13_1576 <= in_reg[687];
        i_13_1577 <= in_reg[1199];
        i_13_1578 <= in_reg[1711];
        i_13_1579 <= in_reg[2223];
        i_13_1580 <= in_reg[2735];
        i_13_1581 <= in_reg[3247];
        i_13_1582 <= in_reg[3759];
        i_13_1583 <= in_reg[4271];
        i_13_1584 <= in_reg[176];
        i_13_1585 <= in_reg[688];
        i_13_1586 <= in_reg[1200];
        i_13_1587 <= in_reg[1712];
        i_13_1588 <= in_reg[2224];
        i_13_1589 <= in_reg[2736];
        i_13_1590 <= in_reg[3248];
        i_13_1591 <= in_reg[3760];
        i_13_1592 <= in_reg[4272];
        i_13_1593 <= in_reg[177];
        i_13_1594 <= in_reg[689];
        i_13_1595 <= in_reg[1201];
        i_13_1596 <= in_reg[1713];
        i_13_1597 <= in_reg[2225];
        i_13_1598 <= in_reg[2737];
        i_13_1599 <= in_reg[3249];
        i_13_1600 <= in_reg[3761];
        i_13_1601 <= in_reg[4273];
        i_13_1602 <= in_reg[178];
        i_13_1603 <= in_reg[690];
        i_13_1604 <= in_reg[1202];
        i_13_1605 <= in_reg[1714];
        i_13_1606 <= in_reg[2226];
        i_13_1607 <= in_reg[2738];
        i_13_1608 <= in_reg[3250];
        i_13_1609 <= in_reg[3762];
        i_13_1610 <= in_reg[4274];
        i_13_1611 <= in_reg[179];
        i_13_1612 <= in_reg[691];
        i_13_1613 <= in_reg[1203];
        i_13_1614 <= in_reg[1715];
        i_13_1615 <= in_reg[2227];
        i_13_1616 <= in_reg[2739];
        i_13_1617 <= in_reg[3251];
        i_13_1618 <= in_reg[3763];
        i_13_1619 <= in_reg[4275];
        i_13_1620 <= in_reg[180];
        i_13_1621 <= in_reg[692];
        i_13_1622 <= in_reg[1204];
        i_13_1623 <= in_reg[1716];
        i_13_1624 <= in_reg[2228];
        i_13_1625 <= in_reg[2740];
        i_13_1626 <= in_reg[3252];
        i_13_1627 <= in_reg[3764];
        i_13_1628 <= in_reg[4276];
        i_13_1629 <= in_reg[181];
        i_13_1630 <= in_reg[693];
        i_13_1631 <= in_reg[1205];
        i_13_1632 <= in_reg[1717];
        i_13_1633 <= in_reg[2229];
        i_13_1634 <= in_reg[2741];
        i_13_1635 <= in_reg[3253];
        i_13_1636 <= in_reg[3765];
        i_13_1637 <= in_reg[4277];
        i_13_1638 <= in_reg[182];
        i_13_1639 <= in_reg[694];
        i_13_1640 <= in_reg[1206];
        i_13_1641 <= in_reg[1718];
        i_13_1642 <= in_reg[2230];
        i_13_1643 <= in_reg[2742];
        i_13_1644 <= in_reg[3254];
        i_13_1645 <= in_reg[3766];
        i_13_1646 <= in_reg[4278];
        i_13_1647 <= in_reg[183];
        i_13_1648 <= in_reg[695];
        i_13_1649 <= in_reg[1207];
        i_13_1650 <= in_reg[1719];
        i_13_1651 <= in_reg[2231];
        i_13_1652 <= in_reg[2743];
        i_13_1653 <= in_reg[3255];
        i_13_1654 <= in_reg[3767];
        i_13_1655 <= in_reg[4279];
        i_13_1656 <= in_reg[184];
        i_13_1657 <= in_reg[696];
        i_13_1658 <= in_reg[1208];
        i_13_1659 <= in_reg[1720];
        i_13_1660 <= in_reg[2232];
        i_13_1661 <= in_reg[2744];
        i_13_1662 <= in_reg[3256];
        i_13_1663 <= in_reg[3768];
        i_13_1664 <= in_reg[4280];
        i_13_1665 <= in_reg[185];
        i_13_1666 <= in_reg[697];
        i_13_1667 <= in_reg[1209];
        i_13_1668 <= in_reg[1721];
        i_13_1669 <= in_reg[2233];
        i_13_1670 <= in_reg[2745];
        i_13_1671 <= in_reg[3257];
        i_13_1672 <= in_reg[3769];
        i_13_1673 <= in_reg[4281];
        i_13_1674 <= in_reg[186];
        i_13_1675 <= in_reg[698];
        i_13_1676 <= in_reg[1210];
        i_13_1677 <= in_reg[1722];
        i_13_1678 <= in_reg[2234];
        i_13_1679 <= in_reg[2746];
        i_13_1680 <= in_reg[3258];
        i_13_1681 <= in_reg[3770];
        i_13_1682 <= in_reg[4282];
        i_13_1683 <= in_reg[187];
        i_13_1684 <= in_reg[699];
        i_13_1685 <= in_reg[1211];
        i_13_1686 <= in_reg[1723];
        i_13_1687 <= in_reg[2235];
        i_13_1688 <= in_reg[2747];
        i_13_1689 <= in_reg[3259];
        i_13_1690 <= in_reg[3771];
        i_13_1691 <= in_reg[4283];
        i_13_1692 <= in_reg[188];
        i_13_1693 <= in_reg[700];
        i_13_1694 <= in_reg[1212];
        i_13_1695 <= in_reg[1724];
        i_13_1696 <= in_reg[2236];
        i_13_1697 <= in_reg[2748];
        i_13_1698 <= in_reg[3260];
        i_13_1699 <= in_reg[3772];
        i_13_1700 <= in_reg[4284];
        i_13_1701 <= in_reg[189];
        i_13_1702 <= in_reg[701];
        i_13_1703 <= in_reg[1213];
        i_13_1704 <= in_reg[1725];
        i_13_1705 <= in_reg[2237];
        i_13_1706 <= in_reg[2749];
        i_13_1707 <= in_reg[3261];
        i_13_1708 <= in_reg[3773];
        i_13_1709 <= in_reg[4285];
        i_13_1710 <= in_reg[190];
        i_13_1711 <= in_reg[702];
        i_13_1712 <= in_reg[1214];
        i_13_1713 <= in_reg[1726];
        i_13_1714 <= in_reg[2238];
        i_13_1715 <= in_reg[2750];
        i_13_1716 <= in_reg[3262];
        i_13_1717 <= in_reg[3774];
        i_13_1718 <= in_reg[4286];
        i_13_1719 <= in_reg[191];
        i_13_1720 <= in_reg[703];
        i_13_1721 <= in_reg[1215];
        i_13_1722 <= in_reg[1727];
        i_13_1723 <= in_reg[2239];
        i_13_1724 <= in_reg[2751];
        i_13_1725 <= in_reg[3263];
        i_13_1726 <= in_reg[3775];
        i_13_1727 <= in_reg[4287];
        i_13_1728 <= in_reg[192];
        i_13_1729 <= in_reg[704];
        i_13_1730 <= in_reg[1216];
        i_13_1731 <= in_reg[1728];
        i_13_1732 <= in_reg[2240];
        i_13_1733 <= in_reg[2752];
        i_13_1734 <= in_reg[3264];
        i_13_1735 <= in_reg[3776];
        i_13_1736 <= in_reg[4288];
        i_13_1737 <= in_reg[193];
        i_13_1738 <= in_reg[705];
        i_13_1739 <= in_reg[1217];
        i_13_1740 <= in_reg[1729];
        i_13_1741 <= in_reg[2241];
        i_13_1742 <= in_reg[2753];
        i_13_1743 <= in_reg[3265];
        i_13_1744 <= in_reg[3777];
        i_13_1745 <= in_reg[4289];
        i_13_1746 <= in_reg[194];
        i_13_1747 <= in_reg[706];
        i_13_1748 <= in_reg[1218];
        i_13_1749 <= in_reg[1730];
        i_13_1750 <= in_reg[2242];
        i_13_1751 <= in_reg[2754];
        i_13_1752 <= in_reg[3266];
        i_13_1753 <= in_reg[3778];
        i_13_1754 <= in_reg[4290];
        i_13_1755 <= in_reg[195];
        i_13_1756 <= in_reg[707];
        i_13_1757 <= in_reg[1219];
        i_13_1758 <= in_reg[1731];
        i_13_1759 <= in_reg[2243];
        i_13_1760 <= in_reg[2755];
        i_13_1761 <= in_reg[3267];
        i_13_1762 <= in_reg[3779];
        i_13_1763 <= in_reg[4291];
        i_13_1764 <= in_reg[196];
        i_13_1765 <= in_reg[708];
        i_13_1766 <= in_reg[1220];
        i_13_1767 <= in_reg[1732];
        i_13_1768 <= in_reg[2244];
        i_13_1769 <= in_reg[2756];
        i_13_1770 <= in_reg[3268];
        i_13_1771 <= in_reg[3780];
        i_13_1772 <= in_reg[4292];
        i_13_1773 <= in_reg[197];
        i_13_1774 <= in_reg[709];
        i_13_1775 <= in_reg[1221];
        i_13_1776 <= in_reg[1733];
        i_13_1777 <= in_reg[2245];
        i_13_1778 <= in_reg[2757];
        i_13_1779 <= in_reg[3269];
        i_13_1780 <= in_reg[3781];
        i_13_1781 <= in_reg[4293];
        i_13_1782 <= in_reg[198];
        i_13_1783 <= in_reg[710];
        i_13_1784 <= in_reg[1222];
        i_13_1785 <= in_reg[1734];
        i_13_1786 <= in_reg[2246];
        i_13_1787 <= in_reg[2758];
        i_13_1788 <= in_reg[3270];
        i_13_1789 <= in_reg[3782];
        i_13_1790 <= in_reg[4294];
        i_13_1791 <= in_reg[199];
        i_13_1792 <= in_reg[711];
        i_13_1793 <= in_reg[1223];
        i_13_1794 <= in_reg[1735];
        i_13_1795 <= in_reg[2247];
        i_13_1796 <= in_reg[2759];
        i_13_1797 <= in_reg[3271];
        i_13_1798 <= in_reg[3783];
        i_13_1799 <= in_reg[4295];
        i_13_1800 <= in_reg[200];
        i_13_1801 <= in_reg[712];
        i_13_1802 <= in_reg[1224];
        i_13_1803 <= in_reg[1736];
        i_13_1804 <= in_reg[2248];
        i_13_1805 <= in_reg[2760];
        i_13_1806 <= in_reg[3272];
        i_13_1807 <= in_reg[3784];
        i_13_1808 <= in_reg[4296];
        i_13_1809 <= in_reg[201];
        i_13_1810 <= in_reg[713];
        i_13_1811 <= in_reg[1225];
        i_13_1812 <= in_reg[1737];
        i_13_1813 <= in_reg[2249];
        i_13_1814 <= in_reg[2761];
        i_13_1815 <= in_reg[3273];
        i_13_1816 <= in_reg[3785];
        i_13_1817 <= in_reg[4297];
        i_13_1818 <= in_reg[202];
        i_13_1819 <= in_reg[714];
        i_13_1820 <= in_reg[1226];
        i_13_1821 <= in_reg[1738];
        i_13_1822 <= in_reg[2250];
        i_13_1823 <= in_reg[2762];
        i_13_1824 <= in_reg[3274];
        i_13_1825 <= in_reg[3786];
        i_13_1826 <= in_reg[4298];
        i_13_1827 <= in_reg[203];
        i_13_1828 <= in_reg[715];
        i_13_1829 <= in_reg[1227];
        i_13_1830 <= in_reg[1739];
        i_13_1831 <= in_reg[2251];
        i_13_1832 <= in_reg[2763];
        i_13_1833 <= in_reg[3275];
        i_13_1834 <= in_reg[3787];
        i_13_1835 <= in_reg[4299];
        i_13_1836 <= in_reg[204];
        i_13_1837 <= in_reg[716];
        i_13_1838 <= in_reg[1228];
        i_13_1839 <= in_reg[1740];
        i_13_1840 <= in_reg[2252];
        i_13_1841 <= in_reg[2764];
        i_13_1842 <= in_reg[3276];
        i_13_1843 <= in_reg[3788];
        i_13_1844 <= in_reg[4300];
        i_13_1845 <= in_reg[205];
        i_13_1846 <= in_reg[717];
        i_13_1847 <= in_reg[1229];
        i_13_1848 <= in_reg[1741];
        i_13_1849 <= in_reg[2253];
        i_13_1850 <= in_reg[2765];
        i_13_1851 <= in_reg[3277];
        i_13_1852 <= in_reg[3789];
        i_13_1853 <= in_reg[4301];
        i_13_1854 <= in_reg[206];
        i_13_1855 <= in_reg[718];
        i_13_1856 <= in_reg[1230];
        i_13_1857 <= in_reg[1742];
        i_13_1858 <= in_reg[2254];
        i_13_1859 <= in_reg[2766];
        i_13_1860 <= in_reg[3278];
        i_13_1861 <= in_reg[3790];
        i_13_1862 <= in_reg[4302];
        i_13_1863 <= in_reg[207];
        i_13_1864 <= in_reg[719];
        i_13_1865 <= in_reg[1231];
        i_13_1866 <= in_reg[1743];
        i_13_1867 <= in_reg[2255];
        i_13_1868 <= in_reg[2767];
        i_13_1869 <= in_reg[3279];
        i_13_1870 <= in_reg[3791];
        i_13_1871 <= in_reg[4303];
        i_13_1872 <= in_reg[208];
        i_13_1873 <= in_reg[720];
        i_13_1874 <= in_reg[1232];
        i_13_1875 <= in_reg[1744];
        i_13_1876 <= in_reg[2256];
        i_13_1877 <= in_reg[2768];
        i_13_1878 <= in_reg[3280];
        i_13_1879 <= in_reg[3792];
        i_13_1880 <= in_reg[4304];
        i_13_1881 <= in_reg[209];
        i_13_1882 <= in_reg[721];
        i_13_1883 <= in_reg[1233];
        i_13_1884 <= in_reg[1745];
        i_13_1885 <= in_reg[2257];
        i_13_1886 <= in_reg[2769];
        i_13_1887 <= in_reg[3281];
        i_13_1888 <= in_reg[3793];
        i_13_1889 <= in_reg[4305];
        i_13_1890 <= in_reg[210];
        i_13_1891 <= in_reg[722];
        i_13_1892 <= in_reg[1234];
        i_13_1893 <= in_reg[1746];
        i_13_1894 <= in_reg[2258];
        i_13_1895 <= in_reg[2770];
        i_13_1896 <= in_reg[3282];
        i_13_1897 <= in_reg[3794];
        i_13_1898 <= in_reg[4306];
        i_13_1899 <= in_reg[211];
        i_13_1900 <= in_reg[723];
        i_13_1901 <= in_reg[1235];
        i_13_1902 <= in_reg[1747];
        i_13_1903 <= in_reg[2259];
        i_13_1904 <= in_reg[2771];
        i_13_1905 <= in_reg[3283];
        i_13_1906 <= in_reg[3795];
        i_13_1907 <= in_reg[4307];
        i_13_1908 <= in_reg[212];
        i_13_1909 <= in_reg[724];
        i_13_1910 <= in_reg[1236];
        i_13_1911 <= in_reg[1748];
        i_13_1912 <= in_reg[2260];
        i_13_1913 <= in_reg[2772];
        i_13_1914 <= in_reg[3284];
        i_13_1915 <= in_reg[3796];
        i_13_1916 <= in_reg[4308];
        i_13_1917 <= in_reg[213];
        i_13_1918 <= in_reg[725];
        i_13_1919 <= in_reg[1237];
        i_13_1920 <= in_reg[1749];
        i_13_1921 <= in_reg[2261];
        i_13_1922 <= in_reg[2773];
        i_13_1923 <= in_reg[3285];
        i_13_1924 <= in_reg[3797];
        i_13_1925 <= in_reg[4309];
        i_13_1926 <= in_reg[214];
        i_13_1927 <= in_reg[726];
        i_13_1928 <= in_reg[1238];
        i_13_1929 <= in_reg[1750];
        i_13_1930 <= in_reg[2262];
        i_13_1931 <= in_reg[2774];
        i_13_1932 <= in_reg[3286];
        i_13_1933 <= in_reg[3798];
        i_13_1934 <= in_reg[4310];
        i_13_1935 <= in_reg[215];
        i_13_1936 <= in_reg[727];
        i_13_1937 <= in_reg[1239];
        i_13_1938 <= in_reg[1751];
        i_13_1939 <= in_reg[2263];
        i_13_1940 <= in_reg[2775];
        i_13_1941 <= in_reg[3287];
        i_13_1942 <= in_reg[3799];
        i_13_1943 <= in_reg[4311];
        i_13_1944 <= in_reg[216];
        i_13_1945 <= in_reg[728];
        i_13_1946 <= in_reg[1240];
        i_13_1947 <= in_reg[1752];
        i_13_1948 <= in_reg[2264];
        i_13_1949 <= in_reg[2776];
        i_13_1950 <= in_reg[3288];
        i_13_1951 <= in_reg[3800];
        i_13_1952 <= in_reg[4312];
        i_13_1953 <= in_reg[217];
        i_13_1954 <= in_reg[729];
        i_13_1955 <= in_reg[1241];
        i_13_1956 <= in_reg[1753];
        i_13_1957 <= in_reg[2265];
        i_13_1958 <= in_reg[2777];
        i_13_1959 <= in_reg[3289];
        i_13_1960 <= in_reg[3801];
        i_13_1961 <= in_reg[4313];
        i_13_1962 <= in_reg[218];
        i_13_1963 <= in_reg[730];
        i_13_1964 <= in_reg[1242];
        i_13_1965 <= in_reg[1754];
        i_13_1966 <= in_reg[2266];
        i_13_1967 <= in_reg[2778];
        i_13_1968 <= in_reg[3290];
        i_13_1969 <= in_reg[3802];
        i_13_1970 <= in_reg[4314];
        i_13_1971 <= in_reg[219];
        i_13_1972 <= in_reg[731];
        i_13_1973 <= in_reg[1243];
        i_13_1974 <= in_reg[1755];
        i_13_1975 <= in_reg[2267];
        i_13_1976 <= in_reg[2779];
        i_13_1977 <= in_reg[3291];
        i_13_1978 <= in_reg[3803];
        i_13_1979 <= in_reg[4315];
        i_13_1980 <= in_reg[220];
        i_13_1981 <= in_reg[732];
        i_13_1982 <= in_reg[1244];
        i_13_1983 <= in_reg[1756];
        i_13_1984 <= in_reg[2268];
        i_13_1985 <= in_reg[2780];
        i_13_1986 <= in_reg[3292];
        i_13_1987 <= in_reg[3804];
        i_13_1988 <= in_reg[4316];
        i_13_1989 <= in_reg[221];
        i_13_1990 <= in_reg[733];
        i_13_1991 <= in_reg[1245];
        i_13_1992 <= in_reg[1757];
        i_13_1993 <= in_reg[2269];
        i_13_1994 <= in_reg[2781];
        i_13_1995 <= in_reg[3293];
        i_13_1996 <= in_reg[3805];
        i_13_1997 <= in_reg[4317];
        i_13_1998 <= in_reg[222];
        i_13_1999 <= in_reg[734];
        i_13_2000 <= in_reg[1246];
        i_13_2001 <= in_reg[1758];
        i_13_2002 <= in_reg[2270];
        i_13_2003 <= in_reg[2782];
        i_13_2004 <= in_reg[3294];
        i_13_2005 <= in_reg[3806];
        i_13_2006 <= in_reg[4318];
        i_13_2007 <= in_reg[223];
        i_13_2008 <= in_reg[735];
        i_13_2009 <= in_reg[1247];
        i_13_2010 <= in_reg[1759];
        i_13_2011 <= in_reg[2271];
        i_13_2012 <= in_reg[2783];
        i_13_2013 <= in_reg[3295];
        i_13_2014 <= in_reg[3807];
        i_13_2015 <= in_reg[4319];
        i_13_2016 <= in_reg[224];
        i_13_2017 <= in_reg[736];
        i_13_2018 <= in_reg[1248];
        i_13_2019 <= in_reg[1760];
        i_13_2020 <= in_reg[2272];
        i_13_2021 <= in_reg[2784];
        i_13_2022 <= in_reg[3296];
        i_13_2023 <= in_reg[3808];
        i_13_2024 <= in_reg[4320];
        i_13_2025 <= in_reg[225];
        i_13_2026 <= in_reg[737];
        i_13_2027 <= in_reg[1249];
        i_13_2028 <= in_reg[1761];
        i_13_2029 <= in_reg[2273];
        i_13_2030 <= in_reg[2785];
        i_13_2031 <= in_reg[3297];
        i_13_2032 <= in_reg[3809];
        i_13_2033 <= in_reg[4321];
        i_13_2034 <= in_reg[226];
        i_13_2035 <= in_reg[738];
        i_13_2036 <= in_reg[1250];
        i_13_2037 <= in_reg[1762];
        i_13_2038 <= in_reg[2274];
        i_13_2039 <= in_reg[2786];
        i_13_2040 <= in_reg[3298];
        i_13_2041 <= in_reg[3810];
        i_13_2042 <= in_reg[4322];
        i_13_2043 <= in_reg[227];
        i_13_2044 <= in_reg[739];
        i_13_2045 <= in_reg[1251];
        i_13_2046 <= in_reg[1763];
        i_13_2047 <= in_reg[2275];
        i_13_2048 <= in_reg[2787];
        i_13_2049 <= in_reg[3299];
        i_13_2050 <= in_reg[3811];
        i_13_2051 <= in_reg[4323];
        i_13_2052 <= in_reg[228];
        i_13_2053 <= in_reg[740];
        i_13_2054 <= in_reg[1252];
        i_13_2055 <= in_reg[1764];
        i_13_2056 <= in_reg[2276];
        i_13_2057 <= in_reg[2788];
        i_13_2058 <= in_reg[3300];
        i_13_2059 <= in_reg[3812];
        i_13_2060 <= in_reg[4324];
        i_13_2061 <= in_reg[229];
        i_13_2062 <= in_reg[741];
        i_13_2063 <= in_reg[1253];
        i_13_2064 <= in_reg[1765];
        i_13_2065 <= in_reg[2277];
        i_13_2066 <= in_reg[2789];
        i_13_2067 <= in_reg[3301];
        i_13_2068 <= in_reg[3813];
        i_13_2069 <= in_reg[4325];
        i_13_2070 <= in_reg[230];
        i_13_2071 <= in_reg[742];
        i_13_2072 <= in_reg[1254];
        i_13_2073 <= in_reg[1766];
        i_13_2074 <= in_reg[2278];
        i_13_2075 <= in_reg[2790];
        i_13_2076 <= in_reg[3302];
        i_13_2077 <= in_reg[3814];
        i_13_2078 <= in_reg[4326];
        i_13_2079 <= in_reg[231];
        i_13_2080 <= in_reg[743];
        i_13_2081 <= in_reg[1255];
        i_13_2082 <= in_reg[1767];
        i_13_2083 <= in_reg[2279];
        i_13_2084 <= in_reg[2791];
        i_13_2085 <= in_reg[3303];
        i_13_2086 <= in_reg[3815];
        i_13_2087 <= in_reg[4327];
        i_13_2088 <= in_reg[232];
        i_13_2089 <= in_reg[744];
        i_13_2090 <= in_reg[1256];
        i_13_2091 <= in_reg[1768];
        i_13_2092 <= in_reg[2280];
        i_13_2093 <= in_reg[2792];
        i_13_2094 <= in_reg[3304];
        i_13_2095 <= in_reg[3816];
        i_13_2096 <= in_reg[4328];
        i_13_2097 <= in_reg[233];
        i_13_2098 <= in_reg[745];
        i_13_2099 <= in_reg[1257];
        i_13_2100 <= in_reg[1769];
        i_13_2101 <= in_reg[2281];
        i_13_2102 <= in_reg[2793];
        i_13_2103 <= in_reg[3305];
        i_13_2104 <= in_reg[3817];
        i_13_2105 <= in_reg[4329];
        i_13_2106 <= in_reg[234];
        i_13_2107 <= in_reg[746];
        i_13_2108 <= in_reg[1258];
        i_13_2109 <= in_reg[1770];
        i_13_2110 <= in_reg[2282];
        i_13_2111 <= in_reg[2794];
        i_13_2112 <= in_reg[3306];
        i_13_2113 <= in_reg[3818];
        i_13_2114 <= in_reg[4330];
        i_13_2115 <= in_reg[235];
        i_13_2116 <= in_reg[747];
        i_13_2117 <= in_reg[1259];
        i_13_2118 <= in_reg[1771];
        i_13_2119 <= in_reg[2283];
        i_13_2120 <= in_reg[2795];
        i_13_2121 <= in_reg[3307];
        i_13_2122 <= in_reg[3819];
        i_13_2123 <= in_reg[4331];
        i_13_2124 <= in_reg[236];
        i_13_2125 <= in_reg[748];
        i_13_2126 <= in_reg[1260];
        i_13_2127 <= in_reg[1772];
        i_13_2128 <= in_reg[2284];
        i_13_2129 <= in_reg[2796];
        i_13_2130 <= in_reg[3308];
        i_13_2131 <= in_reg[3820];
        i_13_2132 <= in_reg[4332];
        i_13_2133 <= in_reg[237];
        i_13_2134 <= in_reg[749];
        i_13_2135 <= in_reg[1261];
        i_13_2136 <= in_reg[1773];
        i_13_2137 <= in_reg[2285];
        i_13_2138 <= in_reg[2797];
        i_13_2139 <= in_reg[3309];
        i_13_2140 <= in_reg[3821];
        i_13_2141 <= in_reg[4333];
        i_13_2142 <= in_reg[238];
        i_13_2143 <= in_reg[750];
        i_13_2144 <= in_reg[1262];
        i_13_2145 <= in_reg[1774];
        i_13_2146 <= in_reg[2286];
        i_13_2147 <= in_reg[2798];
        i_13_2148 <= in_reg[3310];
        i_13_2149 <= in_reg[3822];
        i_13_2150 <= in_reg[4334];
        i_13_2151 <= in_reg[239];
        i_13_2152 <= in_reg[751];
        i_13_2153 <= in_reg[1263];
        i_13_2154 <= in_reg[1775];
        i_13_2155 <= in_reg[2287];
        i_13_2156 <= in_reg[2799];
        i_13_2157 <= in_reg[3311];
        i_13_2158 <= in_reg[3823];
        i_13_2159 <= in_reg[4335];
        i_13_2160 <= in_reg[240];
        i_13_2161 <= in_reg[752];
        i_13_2162 <= in_reg[1264];
        i_13_2163 <= in_reg[1776];
        i_13_2164 <= in_reg[2288];
        i_13_2165 <= in_reg[2800];
        i_13_2166 <= in_reg[3312];
        i_13_2167 <= in_reg[3824];
        i_13_2168 <= in_reg[4336];
        i_13_2169 <= in_reg[241];
        i_13_2170 <= in_reg[753];
        i_13_2171 <= in_reg[1265];
        i_13_2172 <= in_reg[1777];
        i_13_2173 <= in_reg[2289];
        i_13_2174 <= in_reg[2801];
        i_13_2175 <= in_reg[3313];
        i_13_2176 <= in_reg[3825];
        i_13_2177 <= in_reg[4337];
        i_13_2178 <= in_reg[242];
        i_13_2179 <= in_reg[754];
        i_13_2180 <= in_reg[1266];
        i_13_2181 <= in_reg[1778];
        i_13_2182 <= in_reg[2290];
        i_13_2183 <= in_reg[2802];
        i_13_2184 <= in_reg[3314];
        i_13_2185 <= in_reg[3826];
        i_13_2186 <= in_reg[4338];
        i_13_2187 <= in_reg[243];
        i_13_2188 <= in_reg[755];
        i_13_2189 <= in_reg[1267];
        i_13_2190 <= in_reg[1779];
        i_13_2191 <= in_reg[2291];
        i_13_2192 <= in_reg[2803];
        i_13_2193 <= in_reg[3315];
        i_13_2194 <= in_reg[3827];
        i_13_2195 <= in_reg[4339];
        i_13_2196 <= in_reg[244];
        i_13_2197 <= in_reg[756];
        i_13_2198 <= in_reg[1268];
        i_13_2199 <= in_reg[1780];
        i_13_2200 <= in_reg[2292];
        i_13_2201 <= in_reg[2804];
        i_13_2202 <= in_reg[3316];
        i_13_2203 <= in_reg[3828];
        i_13_2204 <= in_reg[4340];
        i_13_2205 <= in_reg[245];
        i_13_2206 <= in_reg[757];
        i_13_2207 <= in_reg[1269];
        i_13_2208 <= in_reg[1781];
        i_13_2209 <= in_reg[2293];
        i_13_2210 <= in_reg[2805];
        i_13_2211 <= in_reg[3317];
        i_13_2212 <= in_reg[3829];
        i_13_2213 <= in_reg[4341];
        i_13_2214 <= in_reg[246];
        i_13_2215 <= in_reg[758];
        i_13_2216 <= in_reg[1270];
        i_13_2217 <= in_reg[1782];
        i_13_2218 <= in_reg[2294];
        i_13_2219 <= in_reg[2806];
        i_13_2220 <= in_reg[3318];
        i_13_2221 <= in_reg[3830];
        i_13_2222 <= in_reg[4342];
        i_13_2223 <= in_reg[247];
        i_13_2224 <= in_reg[759];
        i_13_2225 <= in_reg[1271];
        i_13_2226 <= in_reg[1783];
        i_13_2227 <= in_reg[2295];
        i_13_2228 <= in_reg[2807];
        i_13_2229 <= in_reg[3319];
        i_13_2230 <= in_reg[3831];
        i_13_2231 <= in_reg[4343];
        i_13_2232 <= in_reg[248];
        i_13_2233 <= in_reg[760];
        i_13_2234 <= in_reg[1272];
        i_13_2235 <= in_reg[1784];
        i_13_2236 <= in_reg[2296];
        i_13_2237 <= in_reg[2808];
        i_13_2238 <= in_reg[3320];
        i_13_2239 <= in_reg[3832];
        i_13_2240 <= in_reg[4344];
        i_13_2241 <= in_reg[249];
        i_13_2242 <= in_reg[761];
        i_13_2243 <= in_reg[1273];
        i_13_2244 <= in_reg[1785];
        i_13_2245 <= in_reg[2297];
        i_13_2246 <= in_reg[2809];
        i_13_2247 <= in_reg[3321];
        i_13_2248 <= in_reg[3833];
        i_13_2249 <= in_reg[4345];
        i_13_2250 <= in_reg[250];
        i_13_2251 <= in_reg[762];
        i_13_2252 <= in_reg[1274];
        i_13_2253 <= in_reg[1786];
        i_13_2254 <= in_reg[2298];
        i_13_2255 <= in_reg[2810];
        i_13_2256 <= in_reg[3322];
        i_13_2257 <= in_reg[3834];
        i_13_2258 <= in_reg[4346];
        i_13_2259 <= in_reg[251];
        i_13_2260 <= in_reg[763];
        i_13_2261 <= in_reg[1275];
        i_13_2262 <= in_reg[1787];
        i_13_2263 <= in_reg[2299];
        i_13_2264 <= in_reg[2811];
        i_13_2265 <= in_reg[3323];
        i_13_2266 <= in_reg[3835];
        i_13_2267 <= in_reg[4347];
        i_13_2268 <= in_reg[252];
        i_13_2269 <= in_reg[764];
        i_13_2270 <= in_reg[1276];
        i_13_2271 <= in_reg[1788];
        i_13_2272 <= in_reg[2300];
        i_13_2273 <= in_reg[2812];
        i_13_2274 <= in_reg[3324];
        i_13_2275 <= in_reg[3836];
        i_13_2276 <= in_reg[4348];
        i_13_2277 <= in_reg[253];
        i_13_2278 <= in_reg[765];
        i_13_2279 <= in_reg[1277];
        i_13_2280 <= in_reg[1789];
        i_13_2281 <= in_reg[2301];
        i_13_2282 <= in_reg[2813];
        i_13_2283 <= in_reg[3325];
        i_13_2284 <= in_reg[3837];
        i_13_2285 <= in_reg[4349];
        i_13_2286 <= in_reg[254];
        i_13_2287 <= in_reg[766];
        i_13_2288 <= in_reg[1278];
        i_13_2289 <= in_reg[1790];
        i_13_2290 <= in_reg[2302];
        i_13_2291 <= in_reg[2814];
        i_13_2292 <= in_reg[3326];
        i_13_2293 <= in_reg[3838];
        i_13_2294 <= in_reg[4350];
        i_13_2295 <= in_reg[255];
        i_13_2296 <= in_reg[767];
        i_13_2297 <= in_reg[1279];
        i_13_2298 <= in_reg[1791];
        i_13_2299 <= in_reg[2303];
        i_13_2300 <= in_reg[2815];
        i_13_2301 <= in_reg[3327];
        i_13_2302 <= in_reg[3839];
        i_13_2303 <= in_reg[4351];
        i_13_2304 <= in_reg[256];
        i_13_2305 <= in_reg[768];
        i_13_2306 <= in_reg[1280];
        i_13_2307 <= in_reg[1792];
        i_13_2308 <= in_reg[2304];
        i_13_2309 <= in_reg[2816];
        i_13_2310 <= in_reg[3328];
        i_13_2311 <= in_reg[3840];
        i_13_2312 <= in_reg[4352];
        i_13_2313 <= in_reg[257];
        i_13_2314 <= in_reg[769];
        i_13_2315 <= in_reg[1281];
        i_13_2316 <= in_reg[1793];
        i_13_2317 <= in_reg[2305];
        i_13_2318 <= in_reg[2817];
        i_13_2319 <= in_reg[3329];
        i_13_2320 <= in_reg[3841];
        i_13_2321 <= in_reg[4353];
        i_13_2322 <= in_reg[258];
        i_13_2323 <= in_reg[770];
        i_13_2324 <= in_reg[1282];
        i_13_2325 <= in_reg[1794];
        i_13_2326 <= in_reg[2306];
        i_13_2327 <= in_reg[2818];
        i_13_2328 <= in_reg[3330];
        i_13_2329 <= in_reg[3842];
        i_13_2330 <= in_reg[4354];
        i_13_2331 <= in_reg[259];
        i_13_2332 <= in_reg[771];
        i_13_2333 <= in_reg[1283];
        i_13_2334 <= in_reg[1795];
        i_13_2335 <= in_reg[2307];
        i_13_2336 <= in_reg[2819];
        i_13_2337 <= in_reg[3331];
        i_13_2338 <= in_reg[3843];
        i_13_2339 <= in_reg[4355];
        i_13_2340 <= in_reg[260];
        i_13_2341 <= in_reg[772];
        i_13_2342 <= in_reg[1284];
        i_13_2343 <= in_reg[1796];
        i_13_2344 <= in_reg[2308];
        i_13_2345 <= in_reg[2820];
        i_13_2346 <= in_reg[3332];
        i_13_2347 <= in_reg[3844];
        i_13_2348 <= in_reg[4356];
        i_13_2349 <= in_reg[261];
        i_13_2350 <= in_reg[773];
        i_13_2351 <= in_reg[1285];
        i_13_2352 <= in_reg[1797];
        i_13_2353 <= in_reg[2309];
        i_13_2354 <= in_reg[2821];
        i_13_2355 <= in_reg[3333];
        i_13_2356 <= in_reg[3845];
        i_13_2357 <= in_reg[4357];
        i_13_2358 <= in_reg[262];
        i_13_2359 <= in_reg[774];
        i_13_2360 <= in_reg[1286];
        i_13_2361 <= in_reg[1798];
        i_13_2362 <= in_reg[2310];
        i_13_2363 <= in_reg[2822];
        i_13_2364 <= in_reg[3334];
        i_13_2365 <= in_reg[3846];
        i_13_2366 <= in_reg[4358];
        i_13_2367 <= in_reg[263];
        i_13_2368 <= in_reg[775];
        i_13_2369 <= in_reg[1287];
        i_13_2370 <= in_reg[1799];
        i_13_2371 <= in_reg[2311];
        i_13_2372 <= in_reg[2823];
        i_13_2373 <= in_reg[3335];
        i_13_2374 <= in_reg[3847];
        i_13_2375 <= in_reg[4359];
        i_13_2376 <= in_reg[264];
        i_13_2377 <= in_reg[776];
        i_13_2378 <= in_reg[1288];
        i_13_2379 <= in_reg[1800];
        i_13_2380 <= in_reg[2312];
        i_13_2381 <= in_reg[2824];
        i_13_2382 <= in_reg[3336];
        i_13_2383 <= in_reg[3848];
        i_13_2384 <= in_reg[4360];
        i_13_2385 <= in_reg[265];
        i_13_2386 <= in_reg[777];
        i_13_2387 <= in_reg[1289];
        i_13_2388 <= in_reg[1801];
        i_13_2389 <= in_reg[2313];
        i_13_2390 <= in_reg[2825];
        i_13_2391 <= in_reg[3337];
        i_13_2392 <= in_reg[3849];
        i_13_2393 <= in_reg[4361];
        i_13_2394 <= in_reg[266];
        i_13_2395 <= in_reg[778];
        i_13_2396 <= in_reg[1290];
        i_13_2397 <= in_reg[1802];
        i_13_2398 <= in_reg[2314];
        i_13_2399 <= in_reg[2826];
        i_13_2400 <= in_reg[3338];
        i_13_2401 <= in_reg[3850];
        i_13_2402 <= in_reg[4362];
        i_13_2403 <= in_reg[267];
        i_13_2404 <= in_reg[779];
        i_13_2405 <= in_reg[1291];
        i_13_2406 <= in_reg[1803];
        i_13_2407 <= in_reg[2315];
        i_13_2408 <= in_reg[2827];
        i_13_2409 <= in_reg[3339];
        i_13_2410 <= in_reg[3851];
        i_13_2411 <= in_reg[4363];
        i_13_2412 <= in_reg[268];
        i_13_2413 <= in_reg[780];
        i_13_2414 <= in_reg[1292];
        i_13_2415 <= in_reg[1804];
        i_13_2416 <= in_reg[2316];
        i_13_2417 <= in_reg[2828];
        i_13_2418 <= in_reg[3340];
        i_13_2419 <= in_reg[3852];
        i_13_2420 <= in_reg[4364];
        i_13_2421 <= in_reg[269];
        i_13_2422 <= in_reg[781];
        i_13_2423 <= in_reg[1293];
        i_13_2424 <= in_reg[1805];
        i_13_2425 <= in_reg[2317];
        i_13_2426 <= in_reg[2829];
        i_13_2427 <= in_reg[3341];
        i_13_2428 <= in_reg[3853];
        i_13_2429 <= in_reg[4365];
        i_13_2430 <= in_reg[270];
        i_13_2431 <= in_reg[782];
        i_13_2432 <= in_reg[1294];
        i_13_2433 <= in_reg[1806];
        i_13_2434 <= in_reg[2318];
        i_13_2435 <= in_reg[2830];
        i_13_2436 <= in_reg[3342];
        i_13_2437 <= in_reg[3854];
        i_13_2438 <= in_reg[4366];
        i_13_2439 <= in_reg[271];
        i_13_2440 <= in_reg[783];
        i_13_2441 <= in_reg[1295];
        i_13_2442 <= in_reg[1807];
        i_13_2443 <= in_reg[2319];
        i_13_2444 <= in_reg[2831];
        i_13_2445 <= in_reg[3343];
        i_13_2446 <= in_reg[3855];
        i_13_2447 <= in_reg[4367];
        i_13_2448 <= in_reg[272];
        i_13_2449 <= in_reg[784];
        i_13_2450 <= in_reg[1296];
        i_13_2451 <= in_reg[1808];
        i_13_2452 <= in_reg[2320];
        i_13_2453 <= in_reg[2832];
        i_13_2454 <= in_reg[3344];
        i_13_2455 <= in_reg[3856];
        i_13_2456 <= in_reg[4368];
        i_13_2457 <= in_reg[273];
        i_13_2458 <= in_reg[785];
        i_13_2459 <= in_reg[1297];
        i_13_2460 <= in_reg[1809];
        i_13_2461 <= in_reg[2321];
        i_13_2462 <= in_reg[2833];
        i_13_2463 <= in_reg[3345];
        i_13_2464 <= in_reg[3857];
        i_13_2465 <= in_reg[4369];
        i_13_2466 <= in_reg[274];
        i_13_2467 <= in_reg[786];
        i_13_2468 <= in_reg[1298];
        i_13_2469 <= in_reg[1810];
        i_13_2470 <= in_reg[2322];
        i_13_2471 <= in_reg[2834];
        i_13_2472 <= in_reg[3346];
        i_13_2473 <= in_reg[3858];
        i_13_2474 <= in_reg[4370];
        i_13_2475 <= in_reg[275];
        i_13_2476 <= in_reg[787];
        i_13_2477 <= in_reg[1299];
        i_13_2478 <= in_reg[1811];
        i_13_2479 <= in_reg[2323];
        i_13_2480 <= in_reg[2835];
        i_13_2481 <= in_reg[3347];
        i_13_2482 <= in_reg[3859];
        i_13_2483 <= in_reg[4371];
        i_13_2484 <= in_reg[276];
        i_13_2485 <= in_reg[788];
        i_13_2486 <= in_reg[1300];
        i_13_2487 <= in_reg[1812];
        i_13_2488 <= in_reg[2324];
        i_13_2489 <= in_reg[2836];
        i_13_2490 <= in_reg[3348];
        i_13_2491 <= in_reg[3860];
        i_13_2492 <= in_reg[4372];
        i_13_2493 <= in_reg[277];
        i_13_2494 <= in_reg[789];
        i_13_2495 <= in_reg[1301];
        i_13_2496 <= in_reg[1813];
        i_13_2497 <= in_reg[2325];
        i_13_2498 <= in_reg[2837];
        i_13_2499 <= in_reg[3349];
        i_13_2500 <= in_reg[3861];
        i_13_2501 <= in_reg[4373];
        i_13_2502 <= in_reg[278];
        i_13_2503 <= in_reg[790];
        i_13_2504 <= in_reg[1302];
        i_13_2505 <= in_reg[1814];
        i_13_2506 <= in_reg[2326];
        i_13_2507 <= in_reg[2838];
        i_13_2508 <= in_reg[3350];
        i_13_2509 <= in_reg[3862];
        i_13_2510 <= in_reg[4374];
        i_13_2511 <= in_reg[279];
        i_13_2512 <= in_reg[791];
        i_13_2513 <= in_reg[1303];
        i_13_2514 <= in_reg[1815];
        i_13_2515 <= in_reg[2327];
        i_13_2516 <= in_reg[2839];
        i_13_2517 <= in_reg[3351];
        i_13_2518 <= in_reg[3863];
        i_13_2519 <= in_reg[4375];
        i_13_2520 <= in_reg[280];
        i_13_2521 <= in_reg[792];
        i_13_2522 <= in_reg[1304];
        i_13_2523 <= in_reg[1816];
        i_13_2524 <= in_reg[2328];
        i_13_2525 <= in_reg[2840];
        i_13_2526 <= in_reg[3352];
        i_13_2527 <= in_reg[3864];
        i_13_2528 <= in_reg[4376];
        i_13_2529 <= in_reg[281];
        i_13_2530 <= in_reg[793];
        i_13_2531 <= in_reg[1305];
        i_13_2532 <= in_reg[1817];
        i_13_2533 <= in_reg[2329];
        i_13_2534 <= in_reg[2841];
        i_13_2535 <= in_reg[3353];
        i_13_2536 <= in_reg[3865];
        i_13_2537 <= in_reg[4377];
        i_13_2538 <= in_reg[282];
        i_13_2539 <= in_reg[794];
        i_13_2540 <= in_reg[1306];
        i_13_2541 <= in_reg[1818];
        i_13_2542 <= in_reg[2330];
        i_13_2543 <= in_reg[2842];
        i_13_2544 <= in_reg[3354];
        i_13_2545 <= in_reg[3866];
        i_13_2546 <= in_reg[4378];
        i_13_2547 <= in_reg[283];
        i_13_2548 <= in_reg[795];
        i_13_2549 <= in_reg[1307];
        i_13_2550 <= in_reg[1819];
        i_13_2551 <= in_reg[2331];
        i_13_2552 <= in_reg[2843];
        i_13_2553 <= in_reg[3355];
        i_13_2554 <= in_reg[3867];
        i_13_2555 <= in_reg[4379];
        i_13_2556 <= in_reg[284];
        i_13_2557 <= in_reg[796];
        i_13_2558 <= in_reg[1308];
        i_13_2559 <= in_reg[1820];
        i_13_2560 <= in_reg[2332];
        i_13_2561 <= in_reg[2844];
        i_13_2562 <= in_reg[3356];
        i_13_2563 <= in_reg[3868];
        i_13_2564 <= in_reg[4380];
        i_13_2565 <= in_reg[285];
        i_13_2566 <= in_reg[797];
        i_13_2567 <= in_reg[1309];
        i_13_2568 <= in_reg[1821];
        i_13_2569 <= in_reg[2333];
        i_13_2570 <= in_reg[2845];
        i_13_2571 <= in_reg[3357];
        i_13_2572 <= in_reg[3869];
        i_13_2573 <= in_reg[4381];
        i_13_2574 <= in_reg[286];
        i_13_2575 <= in_reg[798];
        i_13_2576 <= in_reg[1310];
        i_13_2577 <= in_reg[1822];
        i_13_2578 <= in_reg[2334];
        i_13_2579 <= in_reg[2846];
        i_13_2580 <= in_reg[3358];
        i_13_2581 <= in_reg[3870];
        i_13_2582 <= in_reg[4382];
        i_13_2583 <= in_reg[287];
        i_13_2584 <= in_reg[799];
        i_13_2585 <= in_reg[1311];
        i_13_2586 <= in_reg[1823];
        i_13_2587 <= in_reg[2335];
        i_13_2588 <= in_reg[2847];
        i_13_2589 <= in_reg[3359];
        i_13_2590 <= in_reg[3871];
        i_13_2591 <= in_reg[4383];
        i_13_2592 <= in_reg[288];
        i_13_2593 <= in_reg[800];
        i_13_2594 <= in_reg[1312];
        i_13_2595 <= in_reg[1824];
        i_13_2596 <= in_reg[2336];
        i_13_2597 <= in_reg[2848];
        i_13_2598 <= in_reg[3360];
        i_13_2599 <= in_reg[3872];
        i_13_2600 <= in_reg[4384];
        i_13_2601 <= in_reg[289];
        i_13_2602 <= in_reg[801];
        i_13_2603 <= in_reg[1313];
        i_13_2604 <= in_reg[1825];
        i_13_2605 <= in_reg[2337];
        i_13_2606 <= in_reg[2849];
        i_13_2607 <= in_reg[3361];
        i_13_2608 <= in_reg[3873];
        i_13_2609 <= in_reg[4385];
        i_13_2610 <= in_reg[290];
        i_13_2611 <= in_reg[802];
        i_13_2612 <= in_reg[1314];
        i_13_2613 <= in_reg[1826];
        i_13_2614 <= in_reg[2338];
        i_13_2615 <= in_reg[2850];
        i_13_2616 <= in_reg[3362];
        i_13_2617 <= in_reg[3874];
        i_13_2618 <= in_reg[4386];
        i_13_2619 <= in_reg[291];
        i_13_2620 <= in_reg[803];
        i_13_2621 <= in_reg[1315];
        i_13_2622 <= in_reg[1827];
        i_13_2623 <= in_reg[2339];
        i_13_2624 <= in_reg[2851];
        i_13_2625 <= in_reg[3363];
        i_13_2626 <= in_reg[3875];
        i_13_2627 <= in_reg[4387];
        i_13_2628 <= in_reg[292];
        i_13_2629 <= in_reg[804];
        i_13_2630 <= in_reg[1316];
        i_13_2631 <= in_reg[1828];
        i_13_2632 <= in_reg[2340];
        i_13_2633 <= in_reg[2852];
        i_13_2634 <= in_reg[3364];
        i_13_2635 <= in_reg[3876];
        i_13_2636 <= in_reg[4388];
        i_13_2637 <= in_reg[293];
        i_13_2638 <= in_reg[805];
        i_13_2639 <= in_reg[1317];
        i_13_2640 <= in_reg[1829];
        i_13_2641 <= in_reg[2341];
        i_13_2642 <= in_reg[2853];
        i_13_2643 <= in_reg[3365];
        i_13_2644 <= in_reg[3877];
        i_13_2645 <= in_reg[4389];
        i_13_2646 <= in_reg[294];
        i_13_2647 <= in_reg[806];
        i_13_2648 <= in_reg[1318];
        i_13_2649 <= in_reg[1830];
        i_13_2650 <= in_reg[2342];
        i_13_2651 <= in_reg[2854];
        i_13_2652 <= in_reg[3366];
        i_13_2653 <= in_reg[3878];
        i_13_2654 <= in_reg[4390];
        i_13_2655 <= in_reg[295];
        i_13_2656 <= in_reg[807];
        i_13_2657 <= in_reg[1319];
        i_13_2658 <= in_reg[1831];
        i_13_2659 <= in_reg[2343];
        i_13_2660 <= in_reg[2855];
        i_13_2661 <= in_reg[3367];
        i_13_2662 <= in_reg[3879];
        i_13_2663 <= in_reg[4391];
        i_13_2664 <= in_reg[296];
        i_13_2665 <= in_reg[808];
        i_13_2666 <= in_reg[1320];
        i_13_2667 <= in_reg[1832];
        i_13_2668 <= in_reg[2344];
        i_13_2669 <= in_reg[2856];
        i_13_2670 <= in_reg[3368];
        i_13_2671 <= in_reg[3880];
        i_13_2672 <= in_reg[4392];
        i_13_2673 <= in_reg[297];
        i_13_2674 <= in_reg[809];
        i_13_2675 <= in_reg[1321];
        i_13_2676 <= in_reg[1833];
        i_13_2677 <= in_reg[2345];
        i_13_2678 <= in_reg[2857];
        i_13_2679 <= in_reg[3369];
        i_13_2680 <= in_reg[3881];
        i_13_2681 <= in_reg[4393];
        i_13_2682 <= in_reg[298];
        i_13_2683 <= in_reg[810];
        i_13_2684 <= in_reg[1322];
        i_13_2685 <= in_reg[1834];
        i_13_2686 <= in_reg[2346];
        i_13_2687 <= in_reg[2858];
        i_13_2688 <= in_reg[3370];
        i_13_2689 <= in_reg[3882];
        i_13_2690 <= in_reg[4394];
        i_13_2691 <= in_reg[299];
        i_13_2692 <= in_reg[811];
        i_13_2693 <= in_reg[1323];
        i_13_2694 <= in_reg[1835];
        i_13_2695 <= in_reg[2347];
        i_13_2696 <= in_reg[2859];
        i_13_2697 <= in_reg[3371];
        i_13_2698 <= in_reg[3883];
        i_13_2699 <= in_reg[4395];
        i_13_2700 <= in_reg[300];
        i_13_2701 <= in_reg[812];
        i_13_2702 <= in_reg[1324];
        i_13_2703 <= in_reg[1836];
        i_13_2704 <= in_reg[2348];
        i_13_2705 <= in_reg[2860];
        i_13_2706 <= in_reg[3372];
        i_13_2707 <= in_reg[3884];
        i_13_2708 <= in_reg[4396];
        i_13_2709 <= in_reg[301];
        i_13_2710 <= in_reg[813];
        i_13_2711 <= in_reg[1325];
        i_13_2712 <= in_reg[1837];
        i_13_2713 <= in_reg[2349];
        i_13_2714 <= in_reg[2861];
        i_13_2715 <= in_reg[3373];
        i_13_2716 <= in_reg[3885];
        i_13_2717 <= in_reg[4397];
        i_13_2718 <= in_reg[302];
        i_13_2719 <= in_reg[814];
        i_13_2720 <= in_reg[1326];
        i_13_2721 <= in_reg[1838];
        i_13_2722 <= in_reg[2350];
        i_13_2723 <= in_reg[2862];
        i_13_2724 <= in_reg[3374];
        i_13_2725 <= in_reg[3886];
        i_13_2726 <= in_reg[4398];
        i_13_2727 <= in_reg[303];
        i_13_2728 <= in_reg[815];
        i_13_2729 <= in_reg[1327];
        i_13_2730 <= in_reg[1839];
        i_13_2731 <= in_reg[2351];
        i_13_2732 <= in_reg[2863];
        i_13_2733 <= in_reg[3375];
        i_13_2734 <= in_reg[3887];
        i_13_2735 <= in_reg[4399];
        i_13_2736 <= in_reg[304];
        i_13_2737 <= in_reg[816];
        i_13_2738 <= in_reg[1328];
        i_13_2739 <= in_reg[1840];
        i_13_2740 <= in_reg[2352];
        i_13_2741 <= in_reg[2864];
        i_13_2742 <= in_reg[3376];
        i_13_2743 <= in_reg[3888];
        i_13_2744 <= in_reg[4400];
        i_13_2745 <= in_reg[305];
        i_13_2746 <= in_reg[817];
        i_13_2747 <= in_reg[1329];
        i_13_2748 <= in_reg[1841];
        i_13_2749 <= in_reg[2353];
        i_13_2750 <= in_reg[2865];
        i_13_2751 <= in_reg[3377];
        i_13_2752 <= in_reg[3889];
        i_13_2753 <= in_reg[4401];
        i_13_2754 <= in_reg[306];
        i_13_2755 <= in_reg[818];
        i_13_2756 <= in_reg[1330];
        i_13_2757 <= in_reg[1842];
        i_13_2758 <= in_reg[2354];
        i_13_2759 <= in_reg[2866];
        i_13_2760 <= in_reg[3378];
        i_13_2761 <= in_reg[3890];
        i_13_2762 <= in_reg[4402];
        i_13_2763 <= in_reg[307];
        i_13_2764 <= in_reg[819];
        i_13_2765 <= in_reg[1331];
        i_13_2766 <= in_reg[1843];
        i_13_2767 <= in_reg[2355];
        i_13_2768 <= in_reg[2867];
        i_13_2769 <= in_reg[3379];
        i_13_2770 <= in_reg[3891];
        i_13_2771 <= in_reg[4403];
        i_13_2772 <= in_reg[308];
        i_13_2773 <= in_reg[820];
        i_13_2774 <= in_reg[1332];
        i_13_2775 <= in_reg[1844];
        i_13_2776 <= in_reg[2356];
        i_13_2777 <= in_reg[2868];
        i_13_2778 <= in_reg[3380];
        i_13_2779 <= in_reg[3892];
        i_13_2780 <= in_reg[4404];
        i_13_2781 <= in_reg[309];
        i_13_2782 <= in_reg[821];
        i_13_2783 <= in_reg[1333];
        i_13_2784 <= in_reg[1845];
        i_13_2785 <= in_reg[2357];
        i_13_2786 <= in_reg[2869];
        i_13_2787 <= in_reg[3381];
        i_13_2788 <= in_reg[3893];
        i_13_2789 <= in_reg[4405];
        i_13_2790 <= in_reg[310];
        i_13_2791 <= in_reg[822];
        i_13_2792 <= in_reg[1334];
        i_13_2793 <= in_reg[1846];
        i_13_2794 <= in_reg[2358];
        i_13_2795 <= in_reg[2870];
        i_13_2796 <= in_reg[3382];
        i_13_2797 <= in_reg[3894];
        i_13_2798 <= in_reg[4406];
        i_13_2799 <= in_reg[311];
        i_13_2800 <= in_reg[823];
        i_13_2801 <= in_reg[1335];
        i_13_2802 <= in_reg[1847];
        i_13_2803 <= in_reg[2359];
        i_13_2804 <= in_reg[2871];
        i_13_2805 <= in_reg[3383];
        i_13_2806 <= in_reg[3895];
        i_13_2807 <= in_reg[4407];
        i_13_2808 <= in_reg[312];
        i_13_2809 <= in_reg[824];
        i_13_2810 <= in_reg[1336];
        i_13_2811 <= in_reg[1848];
        i_13_2812 <= in_reg[2360];
        i_13_2813 <= in_reg[2872];
        i_13_2814 <= in_reg[3384];
        i_13_2815 <= in_reg[3896];
        i_13_2816 <= in_reg[4408];
        i_13_2817 <= in_reg[313];
        i_13_2818 <= in_reg[825];
        i_13_2819 <= in_reg[1337];
        i_13_2820 <= in_reg[1849];
        i_13_2821 <= in_reg[2361];
        i_13_2822 <= in_reg[2873];
        i_13_2823 <= in_reg[3385];
        i_13_2824 <= in_reg[3897];
        i_13_2825 <= in_reg[4409];
        i_13_2826 <= in_reg[314];
        i_13_2827 <= in_reg[826];
        i_13_2828 <= in_reg[1338];
        i_13_2829 <= in_reg[1850];
        i_13_2830 <= in_reg[2362];
        i_13_2831 <= in_reg[2874];
        i_13_2832 <= in_reg[3386];
        i_13_2833 <= in_reg[3898];
        i_13_2834 <= in_reg[4410];
        i_13_2835 <= in_reg[315];
        i_13_2836 <= in_reg[827];
        i_13_2837 <= in_reg[1339];
        i_13_2838 <= in_reg[1851];
        i_13_2839 <= in_reg[2363];
        i_13_2840 <= in_reg[2875];
        i_13_2841 <= in_reg[3387];
        i_13_2842 <= in_reg[3899];
        i_13_2843 <= in_reg[4411];
        i_13_2844 <= in_reg[316];
        i_13_2845 <= in_reg[828];
        i_13_2846 <= in_reg[1340];
        i_13_2847 <= in_reg[1852];
        i_13_2848 <= in_reg[2364];
        i_13_2849 <= in_reg[2876];
        i_13_2850 <= in_reg[3388];
        i_13_2851 <= in_reg[3900];
        i_13_2852 <= in_reg[4412];
        i_13_2853 <= in_reg[317];
        i_13_2854 <= in_reg[829];
        i_13_2855 <= in_reg[1341];
        i_13_2856 <= in_reg[1853];
        i_13_2857 <= in_reg[2365];
        i_13_2858 <= in_reg[2877];
        i_13_2859 <= in_reg[3389];
        i_13_2860 <= in_reg[3901];
        i_13_2861 <= in_reg[4413];
        i_13_2862 <= in_reg[318];
        i_13_2863 <= in_reg[830];
        i_13_2864 <= in_reg[1342];
        i_13_2865 <= in_reg[1854];
        i_13_2866 <= in_reg[2366];
        i_13_2867 <= in_reg[2878];
        i_13_2868 <= in_reg[3390];
        i_13_2869 <= in_reg[3902];
        i_13_2870 <= in_reg[4414];
        i_13_2871 <= in_reg[319];
        i_13_2872 <= in_reg[831];
        i_13_2873 <= in_reg[1343];
        i_13_2874 <= in_reg[1855];
        i_13_2875 <= in_reg[2367];
        i_13_2876 <= in_reg[2879];
        i_13_2877 <= in_reg[3391];
        i_13_2878 <= in_reg[3903];
        i_13_2879 <= in_reg[4415];
        i_13_2880 <= in_reg[320];
        i_13_2881 <= in_reg[832];
        i_13_2882 <= in_reg[1344];
        i_13_2883 <= in_reg[1856];
        i_13_2884 <= in_reg[2368];
        i_13_2885 <= in_reg[2880];
        i_13_2886 <= in_reg[3392];
        i_13_2887 <= in_reg[3904];
        i_13_2888 <= in_reg[4416];
        i_13_2889 <= in_reg[321];
        i_13_2890 <= in_reg[833];
        i_13_2891 <= in_reg[1345];
        i_13_2892 <= in_reg[1857];
        i_13_2893 <= in_reg[2369];
        i_13_2894 <= in_reg[2881];
        i_13_2895 <= in_reg[3393];
        i_13_2896 <= in_reg[3905];
        i_13_2897 <= in_reg[4417];
        i_13_2898 <= in_reg[322];
        i_13_2899 <= in_reg[834];
        i_13_2900 <= in_reg[1346];
        i_13_2901 <= in_reg[1858];
        i_13_2902 <= in_reg[2370];
        i_13_2903 <= in_reg[2882];
        i_13_2904 <= in_reg[3394];
        i_13_2905 <= in_reg[3906];
        i_13_2906 <= in_reg[4418];
        i_13_2907 <= in_reg[323];
        i_13_2908 <= in_reg[835];
        i_13_2909 <= in_reg[1347];
        i_13_2910 <= in_reg[1859];
        i_13_2911 <= in_reg[2371];
        i_13_2912 <= in_reg[2883];
        i_13_2913 <= in_reg[3395];
        i_13_2914 <= in_reg[3907];
        i_13_2915 <= in_reg[4419];
        i_13_2916 <= in_reg[324];
        i_13_2917 <= in_reg[836];
        i_13_2918 <= in_reg[1348];
        i_13_2919 <= in_reg[1860];
        i_13_2920 <= in_reg[2372];
        i_13_2921 <= in_reg[2884];
        i_13_2922 <= in_reg[3396];
        i_13_2923 <= in_reg[3908];
        i_13_2924 <= in_reg[4420];
        i_13_2925 <= in_reg[325];
        i_13_2926 <= in_reg[837];
        i_13_2927 <= in_reg[1349];
        i_13_2928 <= in_reg[1861];
        i_13_2929 <= in_reg[2373];
        i_13_2930 <= in_reg[2885];
        i_13_2931 <= in_reg[3397];
        i_13_2932 <= in_reg[3909];
        i_13_2933 <= in_reg[4421];
        i_13_2934 <= in_reg[326];
        i_13_2935 <= in_reg[838];
        i_13_2936 <= in_reg[1350];
        i_13_2937 <= in_reg[1862];
        i_13_2938 <= in_reg[2374];
        i_13_2939 <= in_reg[2886];
        i_13_2940 <= in_reg[3398];
        i_13_2941 <= in_reg[3910];
        i_13_2942 <= in_reg[4422];
        i_13_2943 <= in_reg[327];
        i_13_2944 <= in_reg[839];
        i_13_2945 <= in_reg[1351];
        i_13_2946 <= in_reg[1863];
        i_13_2947 <= in_reg[2375];
        i_13_2948 <= in_reg[2887];
        i_13_2949 <= in_reg[3399];
        i_13_2950 <= in_reg[3911];
        i_13_2951 <= in_reg[4423];
        i_13_2952 <= in_reg[328];
        i_13_2953 <= in_reg[840];
        i_13_2954 <= in_reg[1352];
        i_13_2955 <= in_reg[1864];
        i_13_2956 <= in_reg[2376];
        i_13_2957 <= in_reg[2888];
        i_13_2958 <= in_reg[3400];
        i_13_2959 <= in_reg[3912];
        i_13_2960 <= in_reg[4424];
        i_13_2961 <= in_reg[329];
        i_13_2962 <= in_reg[841];
        i_13_2963 <= in_reg[1353];
        i_13_2964 <= in_reg[1865];
        i_13_2965 <= in_reg[2377];
        i_13_2966 <= in_reg[2889];
        i_13_2967 <= in_reg[3401];
        i_13_2968 <= in_reg[3913];
        i_13_2969 <= in_reg[4425];
        i_13_2970 <= in_reg[330];
        i_13_2971 <= in_reg[842];
        i_13_2972 <= in_reg[1354];
        i_13_2973 <= in_reg[1866];
        i_13_2974 <= in_reg[2378];
        i_13_2975 <= in_reg[2890];
        i_13_2976 <= in_reg[3402];
        i_13_2977 <= in_reg[3914];
        i_13_2978 <= in_reg[4426];
        i_13_2979 <= in_reg[331];
        i_13_2980 <= in_reg[843];
        i_13_2981 <= in_reg[1355];
        i_13_2982 <= in_reg[1867];
        i_13_2983 <= in_reg[2379];
        i_13_2984 <= in_reg[2891];
        i_13_2985 <= in_reg[3403];
        i_13_2986 <= in_reg[3915];
        i_13_2987 <= in_reg[4427];
        i_13_2988 <= in_reg[332];
        i_13_2989 <= in_reg[844];
        i_13_2990 <= in_reg[1356];
        i_13_2991 <= in_reg[1868];
        i_13_2992 <= in_reg[2380];
        i_13_2993 <= in_reg[2892];
        i_13_2994 <= in_reg[3404];
        i_13_2995 <= in_reg[3916];
        i_13_2996 <= in_reg[4428];
        i_13_2997 <= in_reg[333];
        i_13_2998 <= in_reg[845];
        i_13_2999 <= in_reg[1357];
        i_13_3000 <= in_reg[1869];
        i_13_3001 <= in_reg[2381];
        i_13_3002 <= in_reg[2893];
        i_13_3003 <= in_reg[3405];
        i_13_3004 <= in_reg[3917];
        i_13_3005 <= in_reg[4429];
        i_13_3006 <= in_reg[334];
        i_13_3007 <= in_reg[846];
        i_13_3008 <= in_reg[1358];
        i_13_3009 <= in_reg[1870];
        i_13_3010 <= in_reg[2382];
        i_13_3011 <= in_reg[2894];
        i_13_3012 <= in_reg[3406];
        i_13_3013 <= in_reg[3918];
        i_13_3014 <= in_reg[4430];
        i_13_3015 <= in_reg[335];
        i_13_3016 <= in_reg[847];
        i_13_3017 <= in_reg[1359];
        i_13_3018 <= in_reg[1871];
        i_13_3019 <= in_reg[2383];
        i_13_3020 <= in_reg[2895];
        i_13_3021 <= in_reg[3407];
        i_13_3022 <= in_reg[3919];
        i_13_3023 <= in_reg[4431];
        i_13_3024 <= in_reg[336];
        i_13_3025 <= in_reg[848];
        i_13_3026 <= in_reg[1360];
        i_13_3027 <= in_reg[1872];
        i_13_3028 <= in_reg[2384];
        i_13_3029 <= in_reg[2896];
        i_13_3030 <= in_reg[3408];
        i_13_3031 <= in_reg[3920];
        i_13_3032 <= in_reg[4432];
        i_13_3033 <= in_reg[337];
        i_13_3034 <= in_reg[849];
        i_13_3035 <= in_reg[1361];
        i_13_3036 <= in_reg[1873];
        i_13_3037 <= in_reg[2385];
        i_13_3038 <= in_reg[2897];
        i_13_3039 <= in_reg[3409];
        i_13_3040 <= in_reg[3921];
        i_13_3041 <= in_reg[4433];
        i_13_3042 <= in_reg[338];
        i_13_3043 <= in_reg[850];
        i_13_3044 <= in_reg[1362];
        i_13_3045 <= in_reg[1874];
        i_13_3046 <= in_reg[2386];
        i_13_3047 <= in_reg[2898];
        i_13_3048 <= in_reg[3410];
        i_13_3049 <= in_reg[3922];
        i_13_3050 <= in_reg[4434];
        i_13_3051 <= in_reg[339];
        i_13_3052 <= in_reg[851];
        i_13_3053 <= in_reg[1363];
        i_13_3054 <= in_reg[1875];
        i_13_3055 <= in_reg[2387];
        i_13_3056 <= in_reg[2899];
        i_13_3057 <= in_reg[3411];
        i_13_3058 <= in_reg[3923];
        i_13_3059 <= in_reg[4435];
        i_13_3060 <= in_reg[340];
        i_13_3061 <= in_reg[852];
        i_13_3062 <= in_reg[1364];
        i_13_3063 <= in_reg[1876];
        i_13_3064 <= in_reg[2388];
        i_13_3065 <= in_reg[2900];
        i_13_3066 <= in_reg[3412];
        i_13_3067 <= in_reg[3924];
        i_13_3068 <= in_reg[4436];
        i_13_3069 <= in_reg[341];
        i_13_3070 <= in_reg[853];
        i_13_3071 <= in_reg[1365];
        i_13_3072 <= in_reg[1877];
        i_13_3073 <= in_reg[2389];
        i_13_3074 <= in_reg[2901];
        i_13_3075 <= in_reg[3413];
        i_13_3076 <= in_reg[3925];
        i_13_3077 <= in_reg[4437];
        i_13_3078 <= in_reg[342];
        i_13_3079 <= in_reg[854];
        i_13_3080 <= in_reg[1366];
        i_13_3081 <= in_reg[1878];
        i_13_3082 <= in_reg[2390];
        i_13_3083 <= in_reg[2902];
        i_13_3084 <= in_reg[3414];
        i_13_3085 <= in_reg[3926];
        i_13_3086 <= in_reg[4438];
        i_13_3087 <= in_reg[343];
        i_13_3088 <= in_reg[855];
        i_13_3089 <= in_reg[1367];
        i_13_3090 <= in_reg[1879];
        i_13_3091 <= in_reg[2391];
        i_13_3092 <= in_reg[2903];
        i_13_3093 <= in_reg[3415];
        i_13_3094 <= in_reg[3927];
        i_13_3095 <= in_reg[4439];
        i_13_3096 <= in_reg[344];
        i_13_3097 <= in_reg[856];
        i_13_3098 <= in_reg[1368];
        i_13_3099 <= in_reg[1880];
        i_13_3100 <= in_reg[2392];
        i_13_3101 <= in_reg[2904];
        i_13_3102 <= in_reg[3416];
        i_13_3103 <= in_reg[3928];
        i_13_3104 <= in_reg[4440];
        i_13_3105 <= in_reg[345];
        i_13_3106 <= in_reg[857];
        i_13_3107 <= in_reg[1369];
        i_13_3108 <= in_reg[1881];
        i_13_3109 <= in_reg[2393];
        i_13_3110 <= in_reg[2905];
        i_13_3111 <= in_reg[3417];
        i_13_3112 <= in_reg[3929];
        i_13_3113 <= in_reg[4441];
        i_13_3114 <= in_reg[346];
        i_13_3115 <= in_reg[858];
        i_13_3116 <= in_reg[1370];
        i_13_3117 <= in_reg[1882];
        i_13_3118 <= in_reg[2394];
        i_13_3119 <= in_reg[2906];
        i_13_3120 <= in_reg[3418];
        i_13_3121 <= in_reg[3930];
        i_13_3122 <= in_reg[4442];
        i_13_3123 <= in_reg[347];
        i_13_3124 <= in_reg[859];
        i_13_3125 <= in_reg[1371];
        i_13_3126 <= in_reg[1883];
        i_13_3127 <= in_reg[2395];
        i_13_3128 <= in_reg[2907];
        i_13_3129 <= in_reg[3419];
        i_13_3130 <= in_reg[3931];
        i_13_3131 <= in_reg[4443];
        i_13_3132 <= in_reg[348];
        i_13_3133 <= in_reg[860];
        i_13_3134 <= in_reg[1372];
        i_13_3135 <= in_reg[1884];
        i_13_3136 <= in_reg[2396];
        i_13_3137 <= in_reg[2908];
        i_13_3138 <= in_reg[3420];
        i_13_3139 <= in_reg[3932];
        i_13_3140 <= in_reg[4444];
        i_13_3141 <= in_reg[349];
        i_13_3142 <= in_reg[861];
        i_13_3143 <= in_reg[1373];
        i_13_3144 <= in_reg[1885];
        i_13_3145 <= in_reg[2397];
        i_13_3146 <= in_reg[2909];
        i_13_3147 <= in_reg[3421];
        i_13_3148 <= in_reg[3933];
        i_13_3149 <= in_reg[4445];
        i_13_3150 <= in_reg[350];
        i_13_3151 <= in_reg[862];
        i_13_3152 <= in_reg[1374];
        i_13_3153 <= in_reg[1886];
        i_13_3154 <= in_reg[2398];
        i_13_3155 <= in_reg[2910];
        i_13_3156 <= in_reg[3422];
        i_13_3157 <= in_reg[3934];
        i_13_3158 <= in_reg[4446];
        i_13_3159 <= in_reg[351];
        i_13_3160 <= in_reg[863];
        i_13_3161 <= in_reg[1375];
        i_13_3162 <= in_reg[1887];
        i_13_3163 <= in_reg[2399];
        i_13_3164 <= in_reg[2911];
        i_13_3165 <= in_reg[3423];
        i_13_3166 <= in_reg[3935];
        i_13_3167 <= in_reg[4447];
        i_13_3168 <= in_reg[352];
        i_13_3169 <= in_reg[864];
        i_13_3170 <= in_reg[1376];
        i_13_3171 <= in_reg[1888];
        i_13_3172 <= in_reg[2400];
        i_13_3173 <= in_reg[2912];
        i_13_3174 <= in_reg[3424];
        i_13_3175 <= in_reg[3936];
        i_13_3176 <= in_reg[4448];
        i_13_3177 <= in_reg[353];
        i_13_3178 <= in_reg[865];
        i_13_3179 <= in_reg[1377];
        i_13_3180 <= in_reg[1889];
        i_13_3181 <= in_reg[2401];
        i_13_3182 <= in_reg[2913];
        i_13_3183 <= in_reg[3425];
        i_13_3184 <= in_reg[3937];
        i_13_3185 <= in_reg[4449];
        i_13_3186 <= in_reg[354];
        i_13_3187 <= in_reg[866];
        i_13_3188 <= in_reg[1378];
        i_13_3189 <= in_reg[1890];
        i_13_3190 <= in_reg[2402];
        i_13_3191 <= in_reg[2914];
        i_13_3192 <= in_reg[3426];
        i_13_3193 <= in_reg[3938];
        i_13_3194 <= in_reg[4450];
        i_13_3195 <= in_reg[355];
        i_13_3196 <= in_reg[867];
        i_13_3197 <= in_reg[1379];
        i_13_3198 <= in_reg[1891];
        i_13_3199 <= in_reg[2403];
        i_13_3200 <= in_reg[2915];
        i_13_3201 <= in_reg[3427];
        i_13_3202 <= in_reg[3939];
        i_13_3203 <= in_reg[4451];
        i_13_3204 <= in_reg[356];
        i_13_3205 <= in_reg[868];
        i_13_3206 <= in_reg[1380];
        i_13_3207 <= in_reg[1892];
        i_13_3208 <= in_reg[2404];
        i_13_3209 <= in_reg[2916];
        i_13_3210 <= in_reg[3428];
        i_13_3211 <= in_reg[3940];
        i_13_3212 <= in_reg[4452];
        i_13_3213 <= in_reg[357];
        i_13_3214 <= in_reg[869];
        i_13_3215 <= in_reg[1381];
        i_13_3216 <= in_reg[1893];
        i_13_3217 <= in_reg[2405];
        i_13_3218 <= in_reg[2917];
        i_13_3219 <= in_reg[3429];
        i_13_3220 <= in_reg[3941];
        i_13_3221 <= in_reg[4453];
        i_13_3222 <= in_reg[358];
        i_13_3223 <= in_reg[870];
        i_13_3224 <= in_reg[1382];
        i_13_3225 <= in_reg[1894];
        i_13_3226 <= in_reg[2406];
        i_13_3227 <= in_reg[2918];
        i_13_3228 <= in_reg[3430];
        i_13_3229 <= in_reg[3942];
        i_13_3230 <= in_reg[4454];
        i_13_3231 <= in_reg[359];
        i_13_3232 <= in_reg[871];
        i_13_3233 <= in_reg[1383];
        i_13_3234 <= in_reg[1895];
        i_13_3235 <= in_reg[2407];
        i_13_3236 <= in_reg[2919];
        i_13_3237 <= in_reg[3431];
        i_13_3238 <= in_reg[3943];
        i_13_3239 <= in_reg[4455];
        i_13_3240 <= in_reg[360];
        i_13_3241 <= in_reg[872];
        i_13_3242 <= in_reg[1384];
        i_13_3243 <= in_reg[1896];
        i_13_3244 <= in_reg[2408];
        i_13_3245 <= in_reg[2920];
        i_13_3246 <= in_reg[3432];
        i_13_3247 <= in_reg[3944];
        i_13_3248 <= in_reg[4456];
        i_13_3249 <= in_reg[361];
        i_13_3250 <= in_reg[873];
        i_13_3251 <= in_reg[1385];
        i_13_3252 <= in_reg[1897];
        i_13_3253 <= in_reg[2409];
        i_13_3254 <= in_reg[2921];
        i_13_3255 <= in_reg[3433];
        i_13_3256 <= in_reg[3945];
        i_13_3257 <= in_reg[4457];
        i_13_3258 <= in_reg[362];
        i_13_3259 <= in_reg[874];
        i_13_3260 <= in_reg[1386];
        i_13_3261 <= in_reg[1898];
        i_13_3262 <= in_reg[2410];
        i_13_3263 <= in_reg[2922];
        i_13_3264 <= in_reg[3434];
        i_13_3265 <= in_reg[3946];
        i_13_3266 <= in_reg[4458];
        i_13_3267 <= in_reg[363];
        i_13_3268 <= in_reg[875];
        i_13_3269 <= in_reg[1387];
        i_13_3270 <= in_reg[1899];
        i_13_3271 <= in_reg[2411];
        i_13_3272 <= in_reg[2923];
        i_13_3273 <= in_reg[3435];
        i_13_3274 <= in_reg[3947];
        i_13_3275 <= in_reg[4459];
        i_13_3276 <= in_reg[364];
        i_13_3277 <= in_reg[876];
        i_13_3278 <= in_reg[1388];
        i_13_3279 <= in_reg[1900];
        i_13_3280 <= in_reg[2412];
        i_13_3281 <= in_reg[2924];
        i_13_3282 <= in_reg[3436];
        i_13_3283 <= in_reg[3948];
        i_13_3284 <= in_reg[4460];
        i_13_3285 <= in_reg[365];
        i_13_3286 <= in_reg[877];
        i_13_3287 <= in_reg[1389];
        i_13_3288 <= in_reg[1901];
        i_13_3289 <= in_reg[2413];
        i_13_3290 <= in_reg[2925];
        i_13_3291 <= in_reg[3437];
        i_13_3292 <= in_reg[3949];
        i_13_3293 <= in_reg[4461];
        i_13_3294 <= in_reg[366];
        i_13_3295 <= in_reg[878];
        i_13_3296 <= in_reg[1390];
        i_13_3297 <= in_reg[1902];
        i_13_3298 <= in_reg[2414];
        i_13_3299 <= in_reg[2926];
        i_13_3300 <= in_reg[3438];
        i_13_3301 <= in_reg[3950];
        i_13_3302 <= in_reg[4462];
        i_13_3303 <= in_reg[367];
        i_13_3304 <= in_reg[879];
        i_13_3305 <= in_reg[1391];
        i_13_3306 <= in_reg[1903];
        i_13_3307 <= in_reg[2415];
        i_13_3308 <= in_reg[2927];
        i_13_3309 <= in_reg[3439];
        i_13_3310 <= in_reg[3951];
        i_13_3311 <= in_reg[4463];
        i_13_3312 <= in_reg[368];
        i_13_3313 <= in_reg[880];
        i_13_3314 <= in_reg[1392];
        i_13_3315 <= in_reg[1904];
        i_13_3316 <= in_reg[2416];
        i_13_3317 <= in_reg[2928];
        i_13_3318 <= in_reg[3440];
        i_13_3319 <= in_reg[3952];
        i_13_3320 <= in_reg[4464];
        i_13_3321 <= in_reg[369];
        i_13_3322 <= in_reg[881];
        i_13_3323 <= in_reg[1393];
        i_13_3324 <= in_reg[1905];
        i_13_3325 <= in_reg[2417];
        i_13_3326 <= in_reg[2929];
        i_13_3327 <= in_reg[3441];
        i_13_3328 <= in_reg[3953];
        i_13_3329 <= in_reg[4465];
        i_13_3330 <= in_reg[370];
        i_13_3331 <= in_reg[882];
        i_13_3332 <= in_reg[1394];
        i_13_3333 <= in_reg[1906];
        i_13_3334 <= in_reg[2418];
        i_13_3335 <= in_reg[2930];
        i_13_3336 <= in_reg[3442];
        i_13_3337 <= in_reg[3954];
        i_13_3338 <= in_reg[4466];
        i_13_3339 <= in_reg[371];
        i_13_3340 <= in_reg[883];
        i_13_3341 <= in_reg[1395];
        i_13_3342 <= in_reg[1907];
        i_13_3343 <= in_reg[2419];
        i_13_3344 <= in_reg[2931];
        i_13_3345 <= in_reg[3443];
        i_13_3346 <= in_reg[3955];
        i_13_3347 <= in_reg[4467];
        i_13_3348 <= in_reg[372];
        i_13_3349 <= in_reg[884];
        i_13_3350 <= in_reg[1396];
        i_13_3351 <= in_reg[1908];
        i_13_3352 <= in_reg[2420];
        i_13_3353 <= in_reg[2932];
        i_13_3354 <= in_reg[3444];
        i_13_3355 <= in_reg[3956];
        i_13_3356 <= in_reg[4468];
        i_13_3357 <= in_reg[373];
        i_13_3358 <= in_reg[885];
        i_13_3359 <= in_reg[1397];
        i_13_3360 <= in_reg[1909];
        i_13_3361 <= in_reg[2421];
        i_13_3362 <= in_reg[2933];
        i_13_3363 <= in_reg[3445];
        i_13_3364 <= in_reg[3957];
        i_13_3365 <= in_reg[4469];
        i_13_3366 <= in_reg[374];
        i_13_3367 <= in_reg[886];
        i_13_3368 <= in_reg[1398];
        i_13_3369 <= in_reg[1910];
        i_13_3370 <= in_reg[2422];
        i_13_3371 <= in_reg[2934];
        i_13_3372 <= in_reg[3446];
        i_13_3373 <= in_reg[3958];
        i_13_3374 <= in_reg[4470];
        i_13_3375 <= in_reg[375];
        i_13_3376 <= in_reg[887];
        i_13_3377 <= in_reg[1399];
        i_13_3378 <= in_reg[1911];
        i_13_3379 <= in_reg[2423];
        i_13_3380 <= in_reg[2935];
        i_13_3381 <= in_reg[3447];
        i_13_3382 <= in_reg[3959];
        i_13_3383 <= in_reg[4471];
        i_13_3384 <= in_reg[376];
        i_13_3385 <= in_reg[888];
        i_13_3386 <= in_reg[1400];
        i_13_3387 <= in_reg[1912];
        i_13_3388 <= in_reg[2424];
        i_13_3389 <= in_reg[2936];
        i_13_3390 <= in_reg[3448];
        i_13_3391 <= in_reg[3960];
        i_13_3392 <= in_reg[4472];
        i_13_3393 <= in_reg[377];
        i_13_3394 <= in_reg[889];
        i_13_3395 <= in_reg[1401];
        i_13_3396 <= in_reg[1913];
        i_13_3397 <= in_reg[2425];
        i_13_3398 <= in_reg[2937];
        i_13_3399 <= in_reg[3449];
        i_13_3400 <= in_reg[3961];
        i_13_3401 <= in_reg[4473];
        i_13_3402 <= in_reg[378];
        i_13_3403 <= in_reg[890];
        i_13_3404 <= in_reg[1402];
        i_13_3405 <= in_reg[1914];
        i_13_3406 <= in_reg[2426];
        i_13_3407 <= in_reg[2938];
        i_13_3408 <= in_reg[3450];
        i_13_3409 <= in_reg[3962];
        i_13_3410 <= in_reg[4474];
        i_13_3411 <= in_reg[379];
        i_13_3412 <= in_reg[891];
        i_13_3413 <= in_reg[1403];
        i_13_3414 <= in_reg[1915];
        i_13_3415 <= in_reg[2427];
        i_13_3416 <= in_reg[2939];
        i_13_3417 <= in_reg[3451];
        i_13_3418 <= in_reg[3963];
        i_13_3419 <= in_reg[4475];
        i_13_3420 <= in_reg[380];
        i_13_3421 <= in_reg[892];
        i_13_3422 <= in_reg[1404];
        i_13_3423 <= in_reg[1916];
        i_13_3424 <= in_reg[2428];
        i_13_3425 <= in_reg[2940];
        i_13_3426 <= in_reg[3452];
        i_13_3427 <= in_reg[3964];
        i_13_3428 <= in_reg[4476];
        i_13_3429 <= in_reg[381];
        i_13_3430 <= in_reg[893];
        i_13_3431 <= in_reg[1405];
        i_13_3432 <= in_reg[1917];
        i_13_3433 <= in_reg[2429];
        i_13_3434 <= in_reg[2941];
        i_13_3435 <= in_reg[3453];
        i_13_3436 <= in_reg[3965];
        i_13_3437 <= in_reg[4477];
        i_13_3438 <= in_reg[382];
        i_13_3439 <= in_reg[894];
        i_13_3440 <= in_reg[1406];
        i_13_3441 <= in_reg[1918];
        i_13_3442 <= in_reg[2430];
        i_13_3443 <= in_reg[2942];
        i_13_3444 <= in_reg[3454];
        i_13_3445 <= in_reg[3966];
        i_13_3446 <= in_reg[4478];
        i_13_3447 <= in_reg[383];
        i_13_3448 <= in_reg[895];
        i_13_3449 <= in_reg[1407];
        i_13_3450 <= in_reg[1919];
        i_13_3451 <= in_reg[2431];
        i_13_3452 <= in_reg[2943];
        i_13_3453 <= in_reg[3455];
        i_13_3454 <= in_reg[3967];
        i_13_3455 <= in_reg[4479];
        i_13_3456 <= in_reg[384];
        i_13_3457 <= in_reg[896];
        i_13_3458 <= in_reg[1408];
        i_13_3459 <= in_reg[1920];
        i_13_3460 <= in_reg[2432];
        i_13_3461 <= in_reg[2944];
        i_13_3462 <= in_reg[3456];
        i_13_3463 <= in_reg[3968];
        i_13_3464 <= in_reg[4480];
        i_13_3465 <= in_reg[385];
        i_13_3466 <= in_reg[897];
        i_13_3467 <= in_reg[1409];
        i_13_3468 <= in_reg[1921];
        i_13_3469 <= in_reg[2433];
        i_13_3470 <= in_reg[2945];
        i_13_3471 <= in_reg[3457];
        i_13_3472 <= in_reg[3969];
        i_13_3473 <= in_reg[4481];
        i_13_3474 <= in_reg[386];
        i_13_3475 <= in_reg[898];
        i_13_3476 <= in_reg[1410];
        i_13_3477 <= in_reg[1922];
        i_13_3478 <= in_reg[2434];
        i_13_3479 <= in_reg[2946];
        i_13_3480 <= in_reg[3458];
        i_13_3481 <= in_reg[3970];
        i_13_3482 <= in_reg[4482];
        i_13_3483 <= in_reg[387];
        i_13_3484 <= in_reg[899];
        i_13_3485 <= in_reg[1411];
        i_13_3486 <= in_reg[1923];
        i_13_3487 <= in_reg[2435];
        i_13_3488 <= in_reg[2947];
        i_13_3489 <= in_reg[3459];
        i_13_3490 <= in_reg[3971];
        i_13_3491 <= in_reg[4483];
        i_13_3492 <= in_reg[388];
        i_13_3493 <= in_reg[900];
        i_13_3494 <= in_reg[1412];
        i_13_3495 <= in_reg[1924];
        i_13_3496 <= in_reg[2436];
        i_13_3497 <= in_reg[2948];
        i_13_3498 <= in_reg[3460];
        i_13_3499 <= in_reg[3972];
        i_13_3500 <= in_reg[4484];
        i_13_3501 <= in_reg[389];
        i_13_3502 <= in_reg[901];
        i_13_3503 <= in_reg[1413];
        i_13_3504 <= in_reg[1925];
        i_13_3505 <= in_reg[2437];
        i_13_3506 <= in_reg[2949];
        i_13_3507 <= in_reg[3461];
        i_13_3508 <= in_reg[3973];
        i_13_3509 <= in_reg[4485];
        i_13_3510 <= in_reg[390];
        i_13_3511 <= in_reg[902];
        i_13_3512 <= in_reg[1414];
        i_13_3513 <= in_reg[1926];
        i_13_3514 <= in_reg[2438];
        i_13_3515 <= in_reg[2950];
        i_13_3516 <= in_reg[3462];
        i_13_3517 <= in_reg[3974];
        i_13_3518 <= in_reg[4486];
        i_13_3519 <= in_reg[391];
        i_13_3520 <= in_reg[903];
        i_13_3521 <= in_reg[1415];
        i_13_3522 <= in_reg[1927];
        i_13_3523 <= in_reg[2439];
        i_13_3524 <= in_reg[2951];
        i_13_3525 <= in_reg[3463];
        i_13_3526 <= in_reg[3975];
        i_13_3527 <= in_reg[4487];
        i_13_3528 <= in_reg[392];
        i_13_3529 <= in_reg[904];
        i_13_3530 <= in_reg[1416];
        i_13_3531 <= in_reg[1928];
        i_13_3532 <= in_reg[2440];
        i_13_3533 <= in_reg[2952];
        i_13_3534 <= in_reg[3464];
        i_13_3535 <= in_reg[3976];
        i_13_3536 <= in_reg[4488];
        i_13_3537 <= in_reg[393];
        i_13_3538 <= in_reg[905];
        i_13_3539 <= in_reg[1417];
        i_13_3540 <= in_reg[1929];
        i_13_3541 <= in_reg[2441];
        i_13_3542 <= in_reg[2953];
        i_13_3543 <= in_reg[3465];
        i_13_3544 <= in_reg[3977];
        i_13_3545 <= in_reg[4489];
        i_13_3546 <= in_reg[394];
        i_13_3547 <= in_reg[906];
        i_13_3548 <= in_reg[1418];
        i_13_3549 <= in_reg[1930];
        i_13_3550 <= in_reg[2442];
        i_13_3551 <= in_reg[2954];
        i_13_3552 <= in_reg[3466];
        i_13_3553 <= in_reg[3978];
        i_13_3554 <= in_reg[4490];
        i_13_3555 <= in_reg[395];
        i_13_3556 <= in_reg[907];
        i_13_3557 <= in_reg[1419];
        i_13_3558 <= in_reg[1931];
        i_13_3559 <= in_reg[2443];
        i_13_3560 <= in_reg[2955];
        i_13_3561 <= in_reg[3467];
        i_13_3562 <= in_reg[3979];
        i_13_3563 <= in_reg[4491];
        i_13_3564 <= in_reg[396];
        i_13_3565 <= in_reg[908];
        i_13_3566 <= in_reg[1420];
        i_13_3567 <= in_reg[1932];
        i_13_3568 <= in_reg[2444];
        i_13_3569 <= in_reg[2956];
        i_13_3570 <= in_reg[3468];
        i_13_3571 <= in_reg[3980];
        i_13_3572 <= in_reg[4492];
        i_13_3573 <= in_reg[397];
        i_13_3574 <= in_reg[909];
        i_13_3575 <= in_reg[1421];
        i_13_3576 <= in_reg[1933];
        i_13_3577 <= in_reg[2445];
        i_13_3578 <= in_reg[2957];
        i_13_3579 <= in_reg[3469];
        i_13_3580 <= in_reg[3981];
        i_13_3581 <= in_reg[4493];
        i_13_3582 <= in_reg[398];
        i_13_3583 <= in_reg[910];
        i_13_3584 <= in_reg[1422];
        i_13_3585 <= in_reg[1934];
        i_13_3586 <= in_reg[2446];
        i_13_3587 <= in_reg[2958];
        i_13_3588 <= in_reg[3470];
        i_13_3589 <= in_reg[3982];
        i_13_3590 <= in_reg[4494];
        i_13_3591 <= in_reg[399];
        i_13_3592 <= in_reg[911];
        i_13_3593 <= in_reg[1423];
        i_13_3594 <= in_reg[1935];
        i_13_3595 <= in_reg[2447];
        i_13_3596 <= in_reg[2959];
        i_13_3597 <= in_reg[3471];
        i_13_3598 <= in_reg[3983];
        i_13_3599 <= in_reg[4495];
        i_13_3600 <= in_reg[400];
        i_13_3601 <= in_reg[912];
        i_13_3602 <= in_reg[1424];
        i_13_3603 <= in_reg[1936];
        i_13_3604 <= in_reg[2448];
        i_13_3605 <= in_reg[2960];
        i_13_3606 <= in_reg[3472];
        i_13_3607 <= in_reg[3984];
        i_13_3608 <= in_reg[4496];
        i_13_3609 <= in_reg[401];
        i_13_3610 <= in_reg[913];
        i_13_3611 <= in_reg[1425];
        i_13_3612 <= in_reg[1937];
        i_13_3613 <= in_reg[2449];
        i_13_3614 <= in_reg[2961];
        i_13_3615 <= in_reg[3473];
        i_13_3616 <= in_reg[3985];
        i_13_3617 <= in_reg[4497];
        i_13_3618 <= in_reg[402];
        i_13_3619 <= in_reg[914];
        i_13_3620 <= in_reg[1426];
        i_13_3621 <= in_reg[1938];
        i_13_3622 <= in_reg[2450];
        i_13_3623 <= in_reg[2962];
        i_13_3624 <= in_reg[3474];
        i_13_3625 <= in_reg[3986];
        i_13_3626 <= in_reg[4498];
        i_13_3627 <= in_reg[403];
        i_13_3628 <= in_reg[915];
        i_13_3629 <= in_reg[1427];
        i_13_3630 <= in_reg[1939];
        i_13_3631 <= in_reg[2451];
        i_13_3632 <= in_reg[2963];
        i_13_3633 <= in_reg[3475];
        i_13_3634 <= in_reg[3987];
        i_13_3635 <= in_reg[4499];
        i_13_3636 <= in_reg[404];
        i_13_3637 <= in_reg[916];
        i_13_3638 <= in_reg[1428];
        i_13_3639 <= in_reg[1940];
        i_13_3640 <= in_reg[2452];
        i_13_3641 <= in_reg[2964];
        i_13_3642 <= in_reg[3476];
        i_13_3643 <= in_reg[3988];
        i_13_3644 <= in_reg[4500];
        i_13_3645 <= in_reg[405];
        i_13_3646 <= in_reg[917];
        i_13_3647 <= in_reg[1429];
        i_13_3648 <= in_reg[1941];
        i_13_3649 <= in_reg[2453];
        i_13_3650 <= in_reg[2965];
        i_13_3651 <= in_reg[3477];
        i_13_3652 <= in_reg[3989];
        i_13_3653 <= in_reg[4501];
        i_13_3654 <= in_reg[406];
        i_13_3655 <= in_reg[918];
        i_13_3656 <= in_reg[1430];
        i_13_3657 <= in_reg[1942];
        i_13_3658 <= in_reg[2454];
        i_13_3659 <= in_reg[2966];
        i_13_3660 <= in_reg[3478];
        i_13_3661 <= in_reg[3990];
        i_13_3662 <= in_reg[4502];
        i_13_3663 <= in_reg[407];
        i_13_3664 <= in_reg[919];
        i_13_3665 <= in_reg[1431];
        i_13_3666 <= in_reg[1943];
        i_13_3667 <= in_reg[2455];
        i_13_3668 <= in_reg[2967];
        i_13_3669 <= in_reg[3479];
        i_13_3670 <= in_reg[3991];
        i_13_3671 <= in_reg[4503];
        i_13_3672 <= in_reg[408];
        i_13_3673 <= in_reg[920];
        i_13_3674 <= in_reg[1432];
        i_13_3675 <= in_reg[1944];
        i_13_3676 <= in_reg[2456];
        i_13_3677 <= in_reg[2968];
        i_13_3678 <= in_reg[3480];
        i_13_3679 <= in_reg[3992];
        i_13_3680 <= in_reg[4504];
        i_13_3681 <= in_reg[409];
        i_13_3682 <= in_reg[921];
        i_13_3683 <= in_reg[1433];
        i_13_3684 <= in_reg[1945];
        i_13_3685 <= in_reg[2457];
        i_13_3686 <= in_reg[2969];
        i_13_3687 <= in_reg[3481];
        i_13_3688 <= in_reg[3993];
        i_13_3689 <= in_reg[4505];
        i_13_3690 <= in_reg[410];
        i_13_3691 <= in_reg[922];
        i_13_3692 <= in_reg[1434];
        i_13_3693 <= in_reg[1946];
        i_13_3694 <= in_reg[2458];
        i_13_3695 <= in_reg[2970];
        i_13_3696 <= in_reg[3482];
        i_13_3697 <= in_reg[3994];
        i_13_3698 <= in_reg[4506];
        i_13_3699 <= in_reg[411];
        i_13_3700 <= in_reg[923];
        i_13_3701 <= in_reg[1435];
        i_13_3702 <= in_reg[1947];
        i_13_3703 <= in_reg[2459];
        i_13_3704 <= in_reg[2971];
        i_13_3705 <= in_reg[3483];
        i_13_3706 <= in_reg[3995];
        i_13_3707 <= in_reg[4507];
        i_13_3708 <= in_reg[412];
        i_13_3709 <= in_reg[924];
        i_13_3710 <= in_reg[1436];
        i_13_3711 <= in_reg[1948];
        i_13_3712 <= in_reg[2460];
        i_13_3713 <= in_reg[2972];
        i_13_3714 <= in_reg[3484];
        i_13_3715 <= in_reg[3996];
        i_13_3716 <= in_reg[4508];
        i_13_3717 <= in_reg[413];
        i_13_3718 <= in_reg[925];
        i_13_3719 <= in_reg[1437];
        i_13_3720 <= in_reg[1949];
        i_13_3721 <= in_reg[2461];
        i_13_3722 <= in_reg[2973];
        i_13_3723 <= in_reg[3485];
        i_13_3724 <= in_reg[3997];
        i_13_3725 <= in_reg[4509];
        i_13_3726 <= in_reg[414];
        i_13_3727 <= in_reg[926];
        i_13_3728 <= in_reg[1438];
        i_13_3729 <= in_reg[1950];
        i_13_3730 <= in_reg[2462];
        i_13_3731 <= in_reg[2974];
        i_13_3732 <= in_reg[3486];
        i_13_3733 <= in_reg[3998];
        i_13_3734 <= in_reg[4510];
        i_13_3735 <= in_reg[415];
        i_13_3736 <= in_reg[927];
        i_13_3737 <= in_reg[1439];
        i_13_3738 <= in_reg[1951];
        i_13_3739 <= in_reg[2463];
        i_13_3740 <= in_reg[2975];
        i_13_3741 <= in_reg[3487];
        i_13_3742 <= in_reg[3999];
        i_13_3743 <= in_reg[4511];
        i_13_3744 <= in_reg[416];
        i_13_3745 <= in_reg[928];
        i_13_3746 <= in_reg[1440];
        i_13_3747 <= in_reg[1952];
        i_13_3748 <= in_reg[2464];
        i_13_3749 <= in_reg[2976];
        i_13_3750 <= in_reg[3488];
        i_13_3751 <= in_reg[4000];
        i_13_3752 <= in_reg[4512];
        i_13_3753 <= in_reg[417];
        i_13_3754 <= in_reg[929];
        i_13_3755 <= in_reg[1441];
        i_13_3756 <= in_reg[1953];
        i_13_3757 <= in_reg[2465];
        i_13_3758 <= in_reg[2977];
        i_13_3759 <= in_reg[3489];
        i_13_3760 <= in_reg[4001];
        i_13_3761 <= in_reg[4513];
        i_13_3762 <= in_reg[418];
        i_13_3763 <= in_reg[930];
        i_13_3764 <= in_reg[1442];
        i_13_3765 <= in_reg[1954];
        i_13_3766 <= in_reg[2466];
        i_13_3767 <= in_reg[2978];
        i_13_3768 <= in_reg[3490];
        i_13_3769 <= in_reg[4002];
        i_13_3770 <= in_reg[4514];
        i_13_3771 <= in_reg[419];
        i_13_3772 <= in_reg[931];
        i_13_3773 <= in_reg[1443];
        i_13_3774 <= in_reg[1955];
        i_13_3775 <= in_reg[2467];
        i_13_3776 <= in_reg[2979];
        i_13_3777 <= in_reg[3491];
        i_13_3778 <= in_reg[4003];
        i_13_3779 <= in_reg[4515];
        i_13_3780 <= in_reg[420];
        i_13_3781 <= in_reg[932];
        i_13_3782 <= in_reg[1444];
        i_13_3783 <= in_reg[1956];
        i_13_3784 <= in_reg[2468];
        i_13_3785 <= in_reg[2980];
        i_13_3786 <= in_reg[3492];
        i_13_3787 <= in_reg[4004];
        i_13_3788 <= in_reg[4516];
        i_13_3789 <= in_reg[421];
        i_13_3790 <= in_reg[933];
        i_13_3791 <= in_reg[1445];
        i_13_3792 <= in_reg[1957];
        i_13_3793 <= in_reg[2469];
        i_13_3794 <= in_reg[2981];
        i_13_3795 <= in_reg[3493];
        i_13_3796 <= in_reg[4005];
        i_13_3797 <= in_reg[4517];
        i_13_3798 <= in_reg[422];
        i_13_3799 <= in_reg[934];
        i_13_3800 <= in_reg[1446];
        i_13_3801 <= in_reg[1958];
        i_13_3802 <= in_reg[2470];
        i_13_3803 <= in_reg[2982];
        i_13_3804 <= in_reg[3494];
        i_13_3805 <= in_reg[4006];
        i_13_3806 <= in_reg[4518];
        i_13_3807 <= in_reg[423];
        i_13_3808 <= in_reg[935];
        i_13_3809 <= in_reg[1447];
        i_13_3810 <= in_reg[1959];
        i_13_3811 <= in_reg[2471];
        i_13_3812 <= in_reg[2983];
        i_13_3813 <= in_reg[3495];
        i_13_3814 <= in_reg[4007];
        i_13_3815 <= in_reg[4519];
        i_13_3816 <= in_reg[424];
        i_13_3817 <= in_reg[936];
        i_13_3818 <= in_reg[1448];
        i_13_3819 <= in_reg[1960];
        i_13_3820 <= in_reg[2472];
        i_13_3821 <= in_reg[2984];
        i_13_3822 <= in_reg[3496];
        i_13_3823 <= in_reg[4008];
        i_13_3824 <= in_reg[4520];
        i_13_3825 <= in_reg[425];
        i_13_3826 <= in_reg[937];
        i_13_3827 <= in_reg[1449];
        i_13_3828 <= in_reg[1961];
        i_13_3829 <= in_reg[2473];
        i_13_3830 <= in_reg[2985];
        i_13_3831 <= in_reg[3497];
        i_13_3832 <= in_reg[4009];
        i_13_3833 <= in_reg[4521];
        i_13_3834 <= in_reg[426];
        i_13_3835 <= in_reg[938];
        i_13_3836 <= in_reg[1450];
        i_13_3837 <= in_reg[1962];
        i_13_3838 <= in_reg[2474];
        i_13_3839 <= in_reg[2986];
        i_13_3840 <= in_reg[3498];
        i_13_3841 <= in_reg[4010];
        i_13_3842 <= in_reg[4522];
        i_13_3843 <= in_reg[427];
        i_13_3844 <= in_reg[939];
        i_13_3845 <= in_reg[1451];
        i_13_3846 <= in_reg[1963];
        i_13_3847 <= in_reg[2475];
        i_13_3848 <= in_reg[2987];
        i_13_3849 <= in_reg[3499];
        i_13_3850 <= in_reg[4011];
        i_13_3851 <= in_reg[4523];
        i_13_3852 <= in_reg[428];
        i_13_3853 <= in_reg[940];
        i_13_3854 <= in_reg[1452];
        i_13_3855 <= in_reg[1964];
        i_13_3856 <= in_reg[2476];
        i_13_3857 <= in_reg[2988];
        i_13_3858 <= in_reg[3500];
        i_13_3859 <= in_reg[4012];
        i_13_3860 <= in_reg[4524];
        i_13_3861 <= in_reg[429];
        i_13_3862 <= in_reg[941];
        i_13_3863 <= in_reg[1453];
        i_13_3864 <= in_reg[1965];
        i_13_3865 <= in_reg[2477];
        i_13_3866 <= in_reg[2989];
        i_13_3867 <= in_reg[3501];
        i_13_3868 <= in_reg[4013];
        i_13_3869 <= in_reg[4525];
        i_13_3870 <= in_reg[430];
        i_13_3871 <= in_reg[942];
        i_13_3872 <= in_reg[1454];
        i_13_3873 <= in_reg[1966];
        i_13_3874 <= in_reg[2478];
        i_13_3875 <= in_reg[2990];
        i_13_3876 <= in_reg[3502];
        i_13_3877 <= in_reg[4014];
        i_13_3878 <= in_reg[4526];
        i_13_3879 <= in_reg[431];
        i_13_3880 <= in_reg[943];
        i_13_3881 <= in_reg[1455];
        i_13_3882 <= in_reg[1967];
        i_13_3883 <= in_reg[2479];
        i_13_3884 <= in_reg[2991];
        i_13_3885 <= in_reg[3503];
        i_13_3886 <= in_reg[4015];
        i_13_3887 <= in_reg[4527];
        i_13_3888 <= in_reg[432];
        i_13_3889 <= in_reg[944];
        i_13_3890 <= in_reg[1456];
        i_13_3891 <= in_reg[1968];
        i_13_3892 <= in_reg[2480];
        i_13_3893 <= in_reg[2992];
        i_13_3894 <= in_reg[3504];
        i_13_3895 <= in_reg[4016];
        i_13_3896 <= in_reg[4528];
        i_13_3897 <= in_reg[433];
        i_13_3898 <= in_reg[945];
        i_13_3899 <= in_reg[1457];
        i_13_3900 <= in_reg[1969];
        i_13_3901 <= in_reg[2481];
        i_13_3902 <= in_reg[2993];
        i_13_3903 <= in_reg[3505];
        i_13_3904 <= in_reg[4017];
        i_13_3905 <= in_reg[4529];
        i_13_3906 <= in_reg[434];
        i_13_3907 <= in_reg[946];
        i_13_3908 <= in_reg[1458];
        i_13_3909 <= in_reg[1970];
        i_13_3910 <= in_reg[2482];
        i_13_3911 <= in_reg[2994];
        i_13_3912 <= in_reg[3506];
        i_13_3913 <= in_reg[4018];
        i_13_3914 <= in_reg[4530];
        i_13_3915 <= in_reg[435];
        i_13_3916 <= in_reg[947];
        i_13_3917 <= in_reg[1459];
        i_13_3918 <= in_reg[1971];
        i_13_3919 <= in_reg[2483];
        i_13_3920 <= in_reg[2995];
        i_13_3921 <= in_reg[3507];
        i_13_3922 <= in_reg[4019];
        i_13_3923 <= in_reg[4531];
        i_13_3924 <= in_reg[436];
        i_13_3925 <= in_reg[948];
        i_13_3926 <= in_reg[1460];
        i_13_3927 <= in_reg[1972];
        i_13_3928 <= in_reg[2484];
        i_13_3929 <= in_reg[2996];
        i_13_3930 <= in_reg[3508];
        i_13_3931 <= in_reg[4020];
        i_13_3932 <= in_reg[4532];
        i_13_3933 <= in_reg[437];
        i_13_3934 <= in_reg[949];
        i_13_3935 <= in_reg[1461];
        i_13_3936 <= in_reg[1973];
        i_13_3937 <= in_reg[2485];
        i_13_3938 <= in_reg[2997];
        i_13_3939 <= in_reg[3509];
        i_13_3940 <= in_reg[4021];
        i_13_3941 <= in_reg[4533];
        i_13_3942 <= in_reg[438];
        i_13_3943 <= in_reg[950];
        i_13_3944 <= in_reg[1462];
        i_13_3945 <= in_reg[1974];
        i_13_3946 <= in_reg[2486];
        i_13_3947 <= in_reg[2998];
        i_13_3948 <= in_reg[3510];
        i_13_3949 <= in_reg[4022];
        i_13_3950 <= in_reg[4534];
        i_13_3951 <= in_reg[439];
        i_13_3952 <= in_reg[951];
        i_13_3953 <= in_reg[1463];
        i_13_3954 <= in_reg[1975];
        i_13_3955 <= in_reg[2487];
        i_13_3956 <= in_reg[2999];
        i_13_3957 <= in_reg[3511];
        i_13_3958 <= in_reg[4023];
        i_13_3959 <= in_reg[4535];
        i_13_3960 <= in_reg[440];
        i_13_3961 <= in_reg[952];
        i_13_3962 <= in_reg[1464];
        i_13_3963 <= in_reg[1976];
        i_13_3964 <= in_reg[2488];
        i_13_3965 <= in_reg[3000];
        i_13_3966 <= in_reg[3512];
        i_13_3967 <= in_reg[4024];
        i_13_3968 <= in_reg[4536];
        i_13_3969 <= in_reg[441];
        i_13_3970 <= in_reg[953];
        i_13_3971 <= in_reg[1465];
        i_13_3972 <= in_reg[1977];
        i_13_3973 <= in_reg[2489];
        i_13_3974 <= in_reg[3001];
        i_13_3975 <= in_reg[3513];
        i_13_3976 <= in_reg[4025];
        i_13_3977 <= in_reg[4537];
        i_13_3978 <= in_reg[442];
        i_13_3979 <= in_reg[954];
        i_13_3980 <= in_reg[1466];
        i_13_3981 <= in_reg[1978];
        i_13_3982 <= in_reg[2490];
        i_13_3983 <= in_reg[3002];
        i_13_3984 <= in_reg[3514];
        i_13_3985 <= in_reg[4026];
        i_13_3986 <= in_reg[4538];
        i_13_3987 <= in_reg[443];
        i_13_3988 <= in_reg[955];
        i_13_3989 <= in_reg[1467];
        i_13_3990 <= in_reg[1979];
        i_13_3991 <= in_reg[2491];
        i_13_3992 <= in_reg[3003];
        i_13_3993 <= in_reg[3515];
        i_13_3994 <= in_reg[4027];
        i_13_3995 <= in_reg[4539];
        i_13_3996 <= in_reg[444];
        i_13_3997 <= in_reg[956];
        i_13_3998 <= in_reg[1468];
        i_13_3999 <= in_reg[1980];
        i_13_4000 <= in_reg[2492];
        i_13_4001 <= in_reg[3004];
        i_13_4002 <= in_reg[3516];
        i_13_4003 <= in_reg[4028];
        i_13_4004 <= in_reg[4540];
        i_13_4005 <= in_reg[445];
        i_13_4006 <= in_reg[957];
        i_13_4007 <= in_reg[1469];
        i_13_4008 <= in_reg[1981];
        i_13_4009 <= in_reg[2493];
        i_13_4010 <= in_reg[3005];
        i_13_4011 <= in_reg[3517];
        i_13_4012 <= in_reg[4029];
        i_13_4013 <= in_reg[4541];
        i_13_4014 <= in_reg[446];
        i_13_4015 <= in_reg[958];
        i_13_4016 <= in_reg[1470];
        i_13_4017 <= in_reg[1982];
        i_13_4018 <= in_reg[2494];
        i_13_4019 <= in_reg[3006];
        i_13_4020 <= in_reg[3518];
        i_13_4021 <= in_reg[4030];
        i_13_4022 <= in_reg[4542];
        i_13_4023 <= in_reg[447];
        i_13_4024 <= in_reg[959];
        i_13_4025 <= in_reg[1471];
        i_13_4026 <= in_reg[1983];
        i_13_4027 <= in_reg[2495];
        i_13_4028 <= in_reg[3007];
        i_13_4029 <= in_reg[3519];
        i_13_4030 <= in_reg[4031];
        i_13_4031 <= in_reg[4543];
        i_13_4032 <= in_reg[448];
        i_13_4033 <= in_reg[960];
        i_13_4034 <= in_reg[1472];
        i_13_4035 <= in_reg[1984];
        i_13_4036 <= in_reg[2496];
        i_13_4037 <= in_reg[3008];
        i_13_4038 <= in_reg[3520];
        i_13_4039 <= in_reg[4032];
        i_13_4040 <= in_reg[4544];
        i_13_4041 <= in_reg[449];
        i_13_4042 <= in_reg[961];
        i_13_4043 <= in_reg[1473];
        i_13_4044 <= in_reg[1985];
        i_13_4045 <= in_reg[2497];
        i_13_4046 <= in_reg[3009];
        i_13_4047 <= in_reg[3521];
        i_13_4048 <= in_reg[4033];
        i_13_4049 <= in_reg[4545];
        i_13_4050 <= in_reg[450];
        i_13_4051 <= in_reg[962];
        i_13_4052 <= in_reg[1474];
        i_13_4053 <= in_reg[1986];
        i_13_4054 <= in_reg[2498];
        i_13_4055 <= in_reg[3010];
        i_13_4056 <= in_reg[3522];
        i_13_4057 <= in_reg[4034];
        i_13_4058 <= in_reg[4546];
        i_13_4059 <= in_reg[451];
        i_13_4060 <= in_reg[963];
        i_13_4061 <= in_reg[1475];
        i_13_4062 <= in_reg[1987];
        i_13_4063 <= in_reg[2499];
        i_13_4064 <= in_reg[3011];
        i_13_4065 <= in_reg[3523];
        i_13_4066 <= in_reg[4035];
        i_13_4067 <= in_reg[4547];
        i_13_4068 <= in_reg[452];
        i_13_4069 <= in_reg[964];
        i_13_4070 <= in_reg[1476];
        i_13_4071 <= in_reg[1988];
        i_13_4072 <= in_reg[2500];
        i_13_4073 <= in_reg[3012];
        i_13_4074 <= in_reg[3524];
        i_13_4075 <= in_reg[4036];
        i_13_4076 <= in_reg[4548];
        i_13_4077 <= in_reg[453];
        i_13_4078 <= in_reg[965];
        i_13_4079 <= in_reg[1477];
        i_13_4080 <= in_reg[1989];
        i_13_4081 <= in_reg[2501];
        i_13_4082 <= in_reg[3013];
        i_13_4083 <= in_reg[3525];
        i_13_4084 <= in_reg[4037];
        i_13_4085 <= in_reg[4549];
        i_13_4086 <= in_reg[454];
        i_13_4087 <= in_reg[966];
        i_13_4088 <= in_reg[1478];
        i_13_4089 <= in_reg[1990];
        i_13_4090 <= in_reg[2502];
        i_13_4091 <= in_reg[3014];
        i_13_4092 <= in_reg[3526];
        i_13_4093 <= in_reg[4038];
        i_13_4094 <= in_reg[4550];
        i_13_4095 <= in_reg[455];
        i_13_4096 <= in_reg[967];
        i_13_4097 <= in_reg[1479];
        i_13_4098 <= in_reg[1991];
        i_13_4099 <= in_reg[2503];
        i_13_4100 <= in_reg[3015];
        i_13_4101 <= in_reg[3527];
        i_13_4102 <= in_reg[4039];
        i_13_4103 <= in_reg[4551];
        i_13_4104 <= in_reg[456];
        i_13_4105 <= in_reg[968];
        i_13_4106 <= in_reg[1480];
        i_13_4107 <= in_reg[1992];
        i_13_4108 <= in_reg[2504];
        i_13_4109 <= in_reg[3016];
        i_13_4110 <= in_reg[3528];
        i_13_4111 <= in_reg[4040];
        i_13_4112 <= in_reg[4552];
        i_13_4113 <= in_reg[457];
        i_13_4114 <= in_reg[969];
        i_13_4115 <= in_reg[1481];
        i_13_4116 <= in_reg[1993];
        i_13_4117 <= in_reg[2505];
        i_13_4118 <= in_reg[3017];
        i_13_4119 <= in_reg[3529];
        i_13_4120 <= in_reg[4041];
        i_13_4121 <= in_reg[4553];
        i_13_4122 <= in_reg[458];
        i_13_4123 <= in_reg[970];
        i_13_4124 <= in_reg[1482];
        i_13_4125 <= in_reg[1994];
        i_13_4126 <= in_reg[2506];
        i_13_4127 <= in_reg[3018];
        i_13_4128 <= in_reg[3530];
        i_13_4129 <= in_reg[4042];
        i_13_4130 <= in_reg[4554];
        i_13_4131 <= in_reg[459];
        i_13_4132 <= in_reg[971];
        i_13_4133 <= in_reg[1483];
        i_13_4134 <= in_reg[1995];
        i_13_4135 <= in_reg[2507];
        i_13_4136 <= in_reg[3019];
        i_13_4137 <= in_reg[3531];
        i_13_4138 <= in_reg[4043];
        i_13_4139 <= in_reg[4555];
        i_13_4140 <= in_reg[460];
        i_13_4141 <= in_reg[972];
        i_13_4142 <= in_reg[1484];
        i_13_4143 <= in_reg[1996];
        i_13_4144 <= in_reg[2508];
        i_13_4145 <= in_reg[3020];
        i_13_4146 <= in_reg[3532];
        i_13_4147 <= in_reg[4044];
        i_13_4148 <= in_reg[4556];
        i_13_4149 <= in_reg[461];
        i_13_4150 <= in_reg[973];
        i_13_4151 <= in_reg[1485];
        i_13_4152 <= in_reg[1997];
        i_13_4153 <= in_reg[2509];
        i_13_4154 <= in_reg[3021];
        i_13_4155 <= in_reg[3533];
        i_13_4156 <= in_reg[4045];
        i_13_4157 <= in_reg[4557];
        i_13_4158 <= in_reg[462];
        i_13_4159 <= in_reg[974];
        i_13_4160 <= in_reg[1486];
        i_13_4161 <= in_reg[1998];
        i_13_4162 <= in_reg[2510];
        i_13_4163 <= in_reg[3022];
        i_13_4164 <= in_reg[3534];
        i_13_4165 <= in_reg[4046];
        i_13_4166 <= in_reg[4558];
        i_13_4167 <= in_reg[463];
        i_13_4168 <= in_reg[975];
        i_13_4169 <= in_reg[1487];
        i_13_4170 <= in_reg[1999];
        i_13_4171 <= in_reg[2511];
        i_13_4172 <= in_reg[3023];
        i_13_4173 <= in_reg[3535];
        i_13_4174 <= in_reg[4047];
        i_13_4175 <= in_reg[4559];
        i_13_4176 <= in_reg[464];
        i_13_4177 <= in_reg[976];
        i_13_4178 <= in_reg[1488];
        i_13_4179 <= in_reg[2000];
        i_13_4180 <= in_reg[2512];
        i_13_4181 <= in_reg[3024];
        i_13_4182 <= in_reg[3536];
        i_13_4183 <= in_reg[4048];
        i_13_4184 <= in_reg[4560];
        i_13_4185 <= in_reg[465];
        i_13_4186 <= in_reg[977];
        i_13_4187 <= in_reg[1489];
        i_13_4188 <= in_reg[2001];
        i_13_4189 <= in_reg[2513];
        i_13_4190 <= in_reg[3025];
        i_13_4191 <= in_reg[3537];
        i_13_4192 <= in_reg[4049];
        i_13_4193 <= in_reg[4561];
        i_13_4194 <= in_reg[466];
        i_13_4195 <= in_reg[978];
        i_13_4196 <= in_reg[1490];
        i_13_4197 <= in_reg[2002];
        i_13_4198 <= in_reg[2514];
        i_13_4199 <= in_reg[3026];
        i_13_4200 <= in_reg[3538];
        i_13_4201 <= in_reg[4050];
        i_13_4202 <= in_reg[4562];
        i_13_4203 <= in_reg[467];
        i_13_4204 <= in_reg[979];
        i_13_4205 <= in_reg[1491];
        i_13_4206 <= in_reg[2003];
        i_13_4207 <= in_reg[2515];
        i_13_4208 <= in_reg[3027];
        i_13_4209 <= in_reg[3539];
        i_13_4210 <= in_reg[4051];
        i_13_4211 <= in_reg[4563];
        i_13_4212 <= in_reg[468];
        i_13_4213 <= in_reg[980];
        i_13_4214 <= in_reg[1492];
        i_13_4215 <= in_reg[2004];
        i_13_4216 <= in_reg[2516];
        i_13_4217 <= in_reg[3028];
        i_13_4218 <= in_reg[3540];
        i_13_4219 <= in_reg[4052];
        i_13_4220 <= in_reg[4564];
        i_13_4221 <= in_reg[469];
        i_13_4222 <= in_reg[981];
        i_13_4223 <= in_reg[1493];
        i_13_4224 <= in_reg[2005];
        i_13_4225 <= in_reg[2517];
        i_13_4226 <= in_reg[3029];
        i_13_4227 <= in_reg[3541];
        i_13_4228 <= in_reg[4053];
        i_13_4229 <= in_reg[4565];
        i_13_4230 <= in_reg[470];
        i_13_4231 <= in_reg[982];
        i_13_4232 <= in_reg[1494];
        i_13_4233 <= in_reg[2006];
        i_13_4234 <= in_reg[2518];
        i_13_4235 <= in_reg[3030];
        i_13_4236 <= in_reg[3542];
        i_13_4237 <= in_reg[4054];
        i_13_4238 <= in_reg[4566];
        i_13_4239 <= in_reg[471];
        i_13_4240 <= in_reg[983];
        i_13_4241 <= in_reg[1495];
        i_13_4242 <= in_reg[2007];
        i_13_4243 <= in_reg[2519];
        i_13_4244 <= in_reg[3031];
        i_13_4245 <= in_reg[3543];
        i_13_4246 <= in_reg[4055];
        i_13_4247 <= in_reg[4567];
        i_13_4248 <= in_reg[472];
        i_13_4249 <= in_reg[984];
        i_13_4250 <= in_reg[1496];
        i_13_4251 <= in_reg[2008];
        i_13_4252 <= in_reg[2520];
        i_13_4253 <= in_reg[3032];
        i_13_4254 <= in_reg[3544];
        i_13_4255 <= in_reg[4056];
        i_13_4256 <= in_reg[4568];
        i_13_4257 <= in_reg[473];
        i_13_4258 <= in_reg[985];
        i_13_4259 <= in_reg[1497];
        i_13_4260 <= in_reg[2009];
        i_13_4261 <= in_reg[2521];
        i_13_4262 <= in_reg[3033];
        i_13_4263 <= in_reg[3545];
        i_13_4264 <= in_reg[4057];
        i_13_4265 <= in_reg[4569];
        i_13_4266 <= in_reg[474];
        i_13_4267 <= in_reg[986];
        i_13_4268 <= in_reg[1498];
        i_13_4269 <= in_reg[2010];
        i_13_4270 <= in_reg[2522];
        i_13_4271 <= in_reg[3034];
        i_13_4272 <= in_reg[3546];
        i_13_4273 <= in_reg[4058];
        i_13_4274 <= in_reg[4570];
        i_13_4275 <= in_reg[475];
        i_13_4276 <= in_reg[987];
        i_13_4277 <= in_reg[1499];
        i_13_4278 <= in_reg[2011];
        i_13_4279 <= in_reg[2523];
        i_13_4280 <= in_reg[3035];
        i_13_4281 <= in_reg[3547];
        i_13_4282 <= in_reg[4059];
        i_13_4283 <= in_reg[4571];
        i_13_4284 <= in_reg[476];
        i_13_4285 <= in_reg[988];
        i_13_4286 <= in_reg[1500];
        i_13_4287 <= in_reg[2012];
        i_13_4288 <= in_reg[2524];
        i_13_4289 <= in_reg[3036];
        i_13_4290 <= in_reg[3548];
        i_13_4291 <= in_reg[4060];
        i_13_4292 <= in_reg[4572];
        i_13_4293 <= in_reg[477];
        i_13_4294 <= in_reg[989];
        i_13_4295 <= in_reg[1501];
        i_13_4296 <= in_reg[2013];
        i_13_4297 <= in_reg[2525];
        i_13_4298 <= in_reg[3037];
        i_13_4299 <= in_reg[3549];
        i_13_4300 <= in_reg[4061];
        i_13_4301 <= in_reg[4573];
        i_13_4302 <= in_reg[478];
        i_13_4303 <= in_reg[990];
        i_13_4304 <= in_reg[1502];
        i_13_4305 <= in_reg[2014];
        i_13_4306 <= in_reg[2526];
        i_13_4307 <= in_reg[3038];
        i_13_4308 <= in_reg[3550];
        i_13_4309 <= in_reg[4062];
        i_13_4310 <= in_reg[4574];
        i_13_4311 <= in_reg[479];
        i_13_4312 <= in_reg[991];
        i_13_4313 <= in_reg[1503];
        i_13_4314 <= in_reg[2015];
        i_13_4315 <= in_reg[2527];
        i_13_4316 <= in_reg[3039];
        i_13_4317 <= in_reg[3551];
        i_13_4318 <= in_reg[4063];
        i_13_4319 <= in_reg[4575];
        i_13_4320 <= in_reg[480];
        i_13_4321 <= in_reg[992];
        i_13_4322 <= in_reg[1504];
        i_13_4323 <= in_reg[2016];
        i_13_4324 <= in_reg[2528];
        i_13_4325 <= in_reg[3040];
        i_13_4326 <= in_reg[3552];
        i_13_4327 <= in_reg[4064];
        i_13_4328 <= in_reg[4576];
        i_13_4329 <= in_reg[481];
        i_13_4330 <= in_reg[993];
        i_13_4331 <= in_reg[1505];
        i_13_4332 <= in_reg[2017];
        i_13_4333 <= in_reg[2529];
        i_13_4334 <= in_reg[3041];
        i_13_4335 <= in_reg[3553];
        i_13_4336 <= in_reg[4065];
        i_13_4337 <= in_reg[4577];
        i_13_4338 <= in_reg[482];
        i_13_4339 <= in_reg[994];
        i_13_4340 <= in_reg[1506];
        i_13_4341 <= in_reg[2018];
        i_13_4342 <= in_reg[2530];
        i_13_4343 <= in_reg[3042];
        i_13_4344 <= in_reg[3554];
        i_13_4345 <= in_reg[4066];
        i_13_4346 <= in_reg[4578];
        i_13_4347 <= in_reg[483];
        i_13_4348 <= in_reg[995];
        i_13_4349 <= in_reg[1507];
        i_13_4350 <= in_reg[2019];
        i_13_4351 <= in_reg[2531];
        i_13_4352 <= in_reg[3043];
        i_13_4353 <= in_reg[3555];
        i_13_4354 <= in_reg[4067];
        i_13_4355 <= in_reg[4579];
        i_13_4356 <= in_reg[484];
        i_13_4357 <= in_reg[996];
        i_13_4358 <= in_reg[1508];
        i_13_4359 <= in_reg[2020];
        i_13_4360 <= in_reg[2532];
        i_13_4361 <= in_reg[3044];
        i_13_4362 <= in_reg[3556];
        i_13_4363 <= in_reg[4068];
        i_13_4364 <= in_reg[4580];
        i_13_4365 <= in_reg[485];
        i_13_4366 <= in_reg[997];
        i_13_4367 <= in_reg[1509];
        i_13_4368 <= in_reg[2021];
        i_13_4369 <= in_reg[2533];
        i_13_4370 <= in_reg[3045];
        i_13_4371 <= in_reg[3557];
        i_13_4372 <= in_reg[4069];
        i_13_4373 <= in_reg[4581];
        i_13_4374 <= in_reg[486];
        i_13_4375 <= in_reg[998];
        i_13_4376 <= in_reg[1510];
        i_13_4377 <= in_reg[2022];
        i_13_4378 <= in_reg[2534];
        i_13_4379 <= in_reg[3046];
        i_13_4380 <= in_reg[3558];
        i_13_4381 <= in_reg[4070];
        i_13_4382 <= in_reg[4582];
        i_13_4383 <= in_reg[487];
        i_13_4384 <= in_reg[999];
        i_13_4385 <= in_reg[1511];
        i_13_4386 <= in_reg[2023];
        i_13_4387 <= in_reg[2535];
        i_13_4388 <= in_reg[3047];
        i_13_4389 <= in_reg[3559];
        i_13_4390 <= in_reg[4071];
        i_13_4391 <= in_reg[4583];
        i_13_4392 <= in_reg[488];
        i_13_4393 <= in_reg[1000];
        i_13_4394 <= in_reg[1512];
        i_13_4395 <= in_reg[2024];
        i_13_4396 <= in_reg[2536];
        i_13_4397 <= in_reg[3048];
        i_13_4398 <= in_reg[3560];
        i_13_4399 <= in_reg[4072];
        i_13_4400 <= in_reg[4584];
        i_13_4401 <= in_reg[489];
        i_13_4402 <= in_reg[1001];
        i_13_4403 <= in_reg[1513];
        i_13_4404 <= in_reg[2025];
        i_13_4405 <= in_reg[2537];
        i_13_4406 <= in_reg[3049];
        i_13_4407 <= in_reg[3561];
        i_13_4408 <= in_reg[4073];
        i_13_4409 <= in_reg[4585];
        i_13_4410 <= in_reg[490];
        i_13_4411 <= in_reg[1002];
        i_13_4412 <= in_reg[1514];
        i_13_4413 <= in_reg[2026];
        i_13_4414 <= in_reg[2538];
        i_13_4415 <= in_reg[3050];
        i_13_4416 <= in_reg[3562];
        i_13_4417 <= in_reg[4074];
        i_13_4418 <= in_reg[4586];
        i_13_4419 <= in_reg[491];
        i_13_4420 <= in_reg[1003];
        i_13_4421 <= in_reg[1515];
        i_13_4422 <= in_reg[2027];
        i_13_4423 <= in_reg[2539];
        i_13_4424 <= in_reg[3051];
        i_13_4425 <= in_reg[3563];
        i_13_4426 <= in_reg[4075];
        i_13_4427 <= in_reg[4587];
        i_13_4428 <= in_reg[492];
        i_13_4429 <= in_reg[1004];
        i_13_4430 <= in_reg[1516];
        i_13_4431 <= in_reg[2028];
        i_13_4432 <= in_reg[2540];
        i_13_4433 <= in_reg[3052];
        i_13_4434 <= in_reg[3564];
        i_13_4435 <= in_reg[4076];
        i_13_4436 <= in_reg[4588];
        i_13_4437 <= in_reg[493];
        i_13_4438 <= in_reg[1005];
        i_13_4439 <= in_reg[1517];
        i_13_4440 <= in_reg[2029];
        i_13_4441 <= in_reg[2541];
        i_13_4442 <= in_reg[3053];
        i_13_4443 <= in_reg[3565];
        i_13_4444 <= in_reg[4077];
        i_13_4445 <= in_reg[4589];
        i_13_4446 <= in_reg[494];
        i_13_4447 <= in_reg[1006];
        i_13_4448 <= in_reg[1518];
        i_13_4449 <= in_reg[2030];
        i_13_4450 <= in_reg[2542];
        i_13_4451 <= in_reg[3054];
        i_13_4452 <= in_reg[3566];
        i_13_4453 <= in_reg[4078];
        i_13_4454 <= in_reg[4590];
        i_13_4455 <= in_reg[495];
        i_13_4456 <= in_reg[1007];
        i_13_4457 <= in_reg[1519];
        i_13_4458 <= in_reg[2031];
        i_13_4459 <= in_reg[2543];
        i_13_4460 <= in_reg[3055];
        i_13_4461 <= in_reg[3567];
        i_13_4462 <= in_reg[4079];
        i_13_4463 <= in_reg[4591];
        i_13_4464 <= in_reg[496];
        i_13_4465 <= in_reg[1008];
        i_13_4466 <= in_reg[1520];
        i_13_4467 <= in_reg[2032];
        i_13_4468 <= in_reg[2544];
        i_13_4469 <= in_reg[3056];
        i_13_4470 <= in_reg[3568];
        i_13_4471 <= in_reg[4080];
        i_13_4472 <= in_reg[4592];
        i_13_4473 <= in_reg[497];
        i_13_4474 <= in_reg[1009];
        i_13_4475 <= in_reg[1521];
        i_13_4476 <= in_reg[2033];
        i_13_4477 <= in_reg[2545];
        i_13_4478 <= in_reg[3057];
        i_13_4479 <= in_reg[3569];
        i_13_4480 <= in_reg[4081];
        i_13_4481 <= in_reg[4593];
        i_13_4482 <= in_reg[498];
        i_13_4483 <= in_reg[1010];
        i_13_4484 <= in_reg[1522];
        i_13_4485 <= in_reg[2034];
        i_13_4486 <= in_reg[2546];
        i_13_4487 <= in_reg[3058];
        i_13_4488 <= in_reg[3570];
        i_13_4489 <= in_reg[4082];
        i_13_4490 <= in_reg[4594];
        i_13_4491 <= in_reg[499];
        i_13_4492 <= in_reg[1011];
        i_13_4493 <= in_reg[1523];
        i_13_4494 <= in_reg[2035];
        i_13_4495 <= in_reg[2547];
        i_13_4496 <= in_reg[3059];
        i_13_4497 <= in_reg[3571];
        i_13_4498 <= in_reg[4083];
        i_13_4499 <= in_reg[4595];
        i_13_4500 <= in_reg[500];
        i_13_4501 <= in_reg[1012];
        i_13_4502 <= in_reg[1524];
        i_13_4503 <= in_reg[2036];
        i_13_4504 <= in_reg[2548];
        i_13_4505 <= in_reg[3060];
        i_13_4506 <= in_reg[3572];
        i_13_4507 <= in_reg[4084];
        i_13_4508 <= in_reg[4596];
        i_13_4509 <= in_reg[501];
        i_13_4510 <= in_reg[1013];
        i_13_4511 <= in_reg[1525];
        i_13_4512 <= in_reg[2037];
        i_13_4513 <= in_reg[2549];
        i_13_4514 <= in_reg[3061];
        i_13_4515 <= in_reg[3573];
        i_13_4516 <= in_reg[4085];
        i_13_4517 <= in_reg[4597];
        i_13_4518 <= in_reg[502];
        i_13_4519 <= in_reg[1014];
        i_13_4520 <= in_reg[1526];
        i_13_4521 <= in_reg[2038];
        i_13_4522 <= in_reg[2550];
        i_13_4523 <= in_reg[3062];
        i_13_4524 <= in_reg[3574];
        i_13_4525 <= in_reg[4086];
        i_13_4526 <= in_reg[4598];
        i_13_4527 <= in_reg[503];
        i_13_4528 <= in_reg[1015];
        i_13_4529 <= in_reg[1527];
        i_13_4530 <= in_reg[2039];
        i_13_4531 <= in_reg[2551];
        i_13_4532 <= in_reg[3063];
        i_13_4533 <= in_reg[3575];
        i_13_4534 <= in_reg[4087];
        i_13_4535 <= in_reg[4599];
        i_13_4536 <= in_reg[504];
        i_13_4537 <= in_reg[1016];
        i_13_4538 <= in_reg[1528];
        i_13_4539 <= in_reg[2040];
        i_13_4540 <= in_reg[2552];
        i_13_4541 <= in_reg[3064];
        i_13_4542 <= in_reg[3576];
        i_13_4543 <= in_reg[4088];
        i_13_4544 <= in_reg[4600];
        i_13_4545 <= in_reg[505];
        i_13_4546 <= in_reg[1017];
        i_13_4547 <= in_reg[1529];
        i_13_4548 <= in_reg[2041];
        i_13_4549 <= in_reg[2553];
        i_13_4550 <= in_reg[3065];
        i_13_4551 <= in_reg[3577];
        i_13_4552 <= in_reg[4089];
        i_13_4553 <= in_reg[4601];
        i_13_4554 <= in_reg[506];
        i_13_4555 <= in_reg[1018];
        i_13_4556 <= in_reg[1530];
        i_13_4557 <= in_reg[2042];
        i_13_4558 <= in_reg[2554];
        i_13_4559 <= in_reg[3066];
        i_13_4560 <= in_reg[3578];
        i_13_4561 <= in_reg[4090];
        i_13_4562 <= in_reg[4602];
        i_13_4563 <= in_reg[507];
        i_13_4564 <= in_reg[1019];
        i_13_4565 <= in_reg[1531];
        i_13_4566 <= in_reg[2043];
        i_13_4567 <= in_reg[2555];
        i_13_4568 <= in_reg[3067];
        i_13_4569 <= in_reg[3579];
        i_13_4570 <= in_reg[4091];
        i_13_4571 <= in_reg[4603];
        i_13_4572 <= in_reg[508];
        i_13_4573 <= in_reg[1020];
        i_13_4574 <= in_reg[1532];
        i_13_4575 <= in_reg[2044];
        i_13_4576 <= in_reg[2556];
        i_13_4577 <= in_reg[3068];
        i_13_4578 <= in_reg[3580];
        i_13_4579 <= in_reg[4092];
        i_13_4580 <= in_reg[4604];
        i_13_4581 <= in_reg[509];
        i_13_4582 <= in_reg[1021];
        i_13_4583 <= in_reg[1533];
        i_13_4584 <= in_reg[2045];
        i_13_4585 <= in_reg[2557];
        i_13_4586 <= in_reg[3069];
        i_13_4587 <= in_reg[3581];
        i_13_4588 <= in_reg[4093];
        i_13_4589 <= in_reg[4605];
        i_13_4590 <= in_reg[510];
        i_13_4591 <= in_reg[1022];
        i_13_4592 <= in_reg[1534];
        i_13_4593 <= in_reg[2046];
        i_13_4594 <= in_reg[2558];
        i_13_4595 <= in_reg[3070];
        i_13_4596 <= in_reg[3582];
        i_13_4597 <= in_reg[4094];
        i_13_4598 <= in_reg[4606];
        i_13_4599 <= in_reg[511];
        i_13_4600 <= in_reg[1023];
        i_13_4601 <= in_reg[1535];
        i_13_4602 <= in_reg[2047];
        i_13_4603 <= in_reg[2559];
        i_13_4604 <= in_reg[3071];
        i_13_4605 <= in_reg[3583];
        i_13_4606 <= in_reg[4095];
        i_13_4607 <= in_reg[4607];
        dly1 <= ap_start;
        dly2 <= dly1;
      end

  assign out_reg_ap_vld = dly2;
  assign ap_ready = dly2;
  assign ap_done = dly2;
  assign ap_idle = ~ap_start;

endmodule
