// Benchmark "kernel_8_0" written by ABC on Sun Jul 19 10:03:02 2020

module kernel_8_0 ( 
    i_8_0_85_0, i_8_0_86_0, i_8_0_136_0, i_8_0_154_0, i_8_0_155_0,
    i_8_0_157_0, i_8_0_181_0, i_8_0_216_0, i_8_0_218_0, i_8_0_220_0,
    i_8_0_221_0, i_8_0_239_0, i_8_0_265_0, i_8_0_330_0, i_8_0_349_0,
    i_8_0_350_0, i_8_0_365_0, i_8_0_377_0, i_8_0_482_0, i_8_0_499_0,
    i_8_0_500_0, i_8_0_526_0, i_8_0_528_0, i_8_0_552_0, i_8_0_614_0,
    i_8_0_676_0, i_8_0_708_0, i_8_0_716_0, i_8_0_719_0, i_8_0_758_0,
    i_8_0_789_0, i_8_0_813_0, i_8_0_824_0, i_8_0_893_0, i_8_0_918_0,
    i_8_0_919_0, i_8_0_940_0, i_8_0_941_0, i_8_0_946_0, i_8_0_985_0,
    i_8_0_1026_0, i_8_0_1029_0, i_8_0_1030_0, i_8_0_1113_0, i_8_0_1114_0,
    i_8_0_1128_0, i_8_0_1134_0, i_8_0_1154_0, i_8_0_1157_0, i_8_0_1264_0,
    i_8_0_1305_0, i_8_0_1306_0, i_8_0_1307_0, i_8_0_1342_0, i_8_0_1343_0,
    i_8_0_1345_0, i_8_0_1346_0, i_8_0_1405_0, i_8_0_1410_0, i_8_0_1434_0,
    i_8_0_1437_0, i_8_0_1468_0, i_8_0_1474_0, i_8_0_1491_0, i_8_0_1508_0,
    i_8_0_1541_0, i_8_0_1547_0, i_8_0_1549_0, i_8_0_1550_0, i_8_0_1562_0,
    i_8_0_1633_0, i_8_0_1647_0, i_8_0_1649_0, i_8_0_1676_0, i_8_0_1678_0,
    i_8_0_1683_0, i_8_0_1702_0, i_8_0_1747_0, i_8_0_1749_0, i_8_0_1751_0,
    i_8_0_1786_0, i_8_0_1790_0, i_8_0_1805_0, i_8_0_1821_0, i_8_0_1825_0,
    i_8_0_1865_0, i_8_0_1868_0, i_8_0_1889_0, i_8_0_1949_0, i_8_0_1988_0,
    i_8_0_2043_0, i_8_0_2048_0, i_8_0_2216_0, i_8_0_2227_0, i_8_0_2243_0,
    i_8_0_2271_0, i_8_0_2273_0, i_8_0_2275_0, i_8_0_2290_0, i_8_0_2291_0,
    o_8_0_0_0  );
  input  i_8_0_85_0, i_8_0_86_0, i_8_0_136_0, i_8_0_154_0, i_8_0_155_0,
    i_8_0_157_0, i_8_0_181_0, i_8_0_216_0, i_8_0_218_0, i_8_0_220_0,
    i_8_0_221_0, i_8_0_239_0, i_8_0_265_0, i_8_0_330_0, i_8_0_349_0,
    i_8_0_350_0, i_8_0_365_0, i_8_0_377_0, i_8_0_482_0, i_8_0_499_0,
    i_8_0_500_0, i_8_0_526_0, i_8_0_528_0, i_8_0_552_0, i_8_0_614_0,
    i_8_0_676_0, i_8_0_708_0, i_8_0_716_0, i_8_0_719_0, i_8_0_758_0,
    i_8_0_789_0, i_8_0_813_0, i_8_0_824_0, i_8_0_893_0, i_8_0_918_0,
    i_8_0_919_0, i_8_0_940_0, i_8_0_941_0, i_8_0_946_0, i_8_0_985_0,
    i_8_0_1026_0, i_8_0_1029_0, i_8_0_1030_0, i_8_0_1113_0, i_8_0_1114_0,
    i_8_0_1128_0, i_8_0_1134_0, i_8_0_1154_0, i_8_0_1157_0, i_8_0_1264_0,
    i_8_0_1305_0, i_8_0_1306_0, i_8_0_1307_0, i_8_0_1342_0, i_8_0_1343_0,
    i_8_0_1345_0, i_8_0_1346_0, i_8_0_1405_0, i_8_0_1410_0, i_8_0_1434_0,
    i_8_0_1437_0, i_8_0_1468_0, i_8_0_1474_0, i_8_0_1491_0, i_8_0_1508_0,
    i_8_0_1541_0, i_8_0_1547_0, i_8_0_1549_0, i_8_0_1550_0, i_8_0_1562_0,
    i_8_0_1633_0, i_8_0_1647_0, i_8_0_1649_0, i_8_0_1676_0, i_8_0_1678_0,
    i_8_0_1683_0, i_8_0_1702_0, i_8_0_1747_0, i_8_0_1749_0, i_8_0_1751_0,
    i_8_0_1786_0, i_8_0_1790_0, i_8_0_1805_0, i_8_0_1821_0, i_8_0_1825_0,
    i_8_0_1865_0, i_8_0_1868_0, i_8_0_1889_0, i_8_0_1949_0, i_8_0_1988_0,
    i_8_0_2043_0, i_8_0_2048_0, i_8_0_2216_0, i_8_0_2227_0, i_8_0_2243_0,
    i_8_0_2271_0, i_8_0_2273_0, i_8_0_2275_0, i_8_0_2290_0, i_8_0_2291_0;
  output o_8_0_0_0;
  assign o_8_0_0_0 = 0;
endmodule



// Benchmark "kernel_8_1" written by ABC on Sun Jul 19 10:03:03 2020

module kernel_8_1 ( 
    i_8_1_32_0, i_8_1_34_0, i_8_1_42_0, i_8_1_53_0, i_8_1_67_0, i_8_1_80_0,
    i_8_1_226_0, i_8_1_233_0, i_8_1_280_0, i_8_1_329_0, i_8_1_364_0,
    i_8_1_386_0, i_8_1_389_0, i_8_1_400_0, i_8_1_415_0, i_8_1_416_0,
    i_8_1_493_0, i_8_1_506_0, i_8_1_529_0, i_8_1_579_0, i_8_1_592_0,
    i_8_1_607_0, i_8_1_635_0, i_8_1_637_0, i_8_1_662_0, i_8_1_669_0,
    i_8_1_673_0, i_8_1_679_0, i_8_1_680_0, i_8_1_700_0, i_8_1_738_0,
    i_8_1_825_0, i_8_1_826_0, i_8_1_837_0, i_8_1_841_0, i_8_1_843_0,
    i_8_1_844_0, i_8_1_856_0, i_8_1_861_0, i_8_1_868_0, i_8_1_968_0,
    i_8_1_1012_0, i_8_1_1056_0, i_8_1_1071_0, i_8_1_1102_0, i_8_1_1105_0,
    i_8_1_1144_0, i_8_1_1189_0, i_8_1_1199_0, i_8_1_1240_0, i_8_1_1243_0,
    i_8_1_1263_0, i_8_1_1283_0, i_8_1_1300_0, i_8_1_1301_0, i_8_1_1316_0,
    i_8_1_1320_0, i_8_1_1363_0, i_8_1_1400_0, i_8_1_1439_0, i_8_1_1440_0,
    i_8_1_1445_0, i_8_1_1460_0, i_8_1_1464_0, i_8_1_1479_0, i_8_1_1480_0,
    i_8_1_1483_0, i_8_1_1505_0, i_8_1_1524_0, i_8_1_1542_0, i_8_1_1545_0,
    i_8_1_1571_0, i_8_1_1573_0, i_8_1_1633_0, i_8_1_1659_0, i_8_1_1687_0,
    i_8_1_1696_0, i_8_1_1767_0, i_8_1_1781_0, i_8_1_1782_0, i_8_1_1785_0,
    i_8_1_1793_0, i_8_1_1804_0, i_8_1_1858_0, i_8_1_1885_0, i_8_1_1929_0,
    i_8_1_1960_0, i_8_1_1984_0, i_8_1_1993_0, i_8_1_1996_0, i_8_1_2038_0,
    i_8_1_2047_0, i_8_1_2058_0, i_8_1_2110_0, i_8_1_2137_0, i_8_1_2143_0,
    i_8_1_2146_0, i_8_1_2155_0, i_8_1_2156_0, i_8_1_2248_0,
    o_8_1_0_0  );
  input  i_8_1_32_0, i_8_1_34_0, i_8_1_42_0, i_8_1_53_0, i_8_1_67_0,
    i_8_1_80_0, i_8_1_226_0, i_8_1_233_0, i_8_1_280_0, i_8_1_329_0,
    i_8_1_364_0, i_8_1_386_0, i_8_1_389_0, i_8_1_400_0, i_8_1_415_0,
    i_8_1_416_0, i_8_1_493_0, i_8_1_506_0, i_8_1_529_0, i_8_1_579_0,
    i_8_1_592_0, i_8_1_607_0, i_8_1_635_0, i_8_1_637_0, i_8_1_662_0,
    i_8_1_669_0, i_8_1_673_0, i_8_1_679_0, i_8_1_680_0, i_8_1_700_0,
    i_8_1_738_0, i_8_1_825_0, i_8_1_826_0, i_8_1_837_0, i_8_1_841_0,
    i_8_1_843_0, i_8_1_844_0, i_8_1_856_0, i_8_1_861_0, i_8_1_868_0,
    i_8_1_968_0, i_8_1_1012_0, i_8_1_1056_0, i_8_1_1071_0, i_8_1_1102_0,
    i_8_1_1105_0, i_8_1_1144_0, i_8_1_1189_0, i_8_1_1199_0, i_8_1_1240_0,
    i_8_1_1243_0, i_8_1_1263_0, i_8_1_1283_0, i_8_1_1300_0, i_8_1_1301_0,
    i_8_1_1316_0, i_8_1_1320_0, i_8_1_1363_0, i_8_1_1400_0, i_8_1_1439_0,
    i_8_1_1440_0, i_8_1_1445_0, i_8_1_1460_0, i_8_1_1464_0, i_8_1_1479_0,
    i_8_1_1480_0, i_8_1_1483_0, i_8_1_1505_0, i_8_1_1524_0, i_8_1_1542_0,
    i_8_1_1545_0, i_8_1_1571_0, i_8_1_1573_0, i_8_1_1633_0, i_8_1_1659_0,
    i_8_1_1687_0, i_8_1_1696_0, i_8_1_1767_0, i_8_1_1781_0, i_8_1_1782_0,
    i_8_1_1785_0, i_8_1_1793_0, i_8_1_1804_0, i_8_1_1858_0, i_8_1_1885_0,
    i_8_1_1929_0, i_8_1_1960_0, i_8_1_1984_0, i_8_1_1993_0, i_8_1_1996_0,
    i_8_1_2038_0, i_8_1_2047_0, i_8_1_2058_0, i_8_1_2110_0, i_8_1_2137_0,
    i_8_1_2143_0, i_8_1_2146_0, i_8_1_2155_0, i_8_1_2156_0, i_8_1_2248_0;
  output o_8_1_0_0;
  assign o_8_1_0_0 = 0;
endmodule



// Benchmark "kernel_8_2" written by ABC on Sun Jul 19 10:03:04 2020

module kernel_8_2 ( 
    i_8_2_2_0, i_8_2_11_0, i_8_2_40_0, i_8_2_55_0, i_8_2_73_0, i_8_2_101_0,
    i_8_2_135_0, i_8_2_181_0, i_8_2_192_0, i_8_2_195_0, i_8_2_225_0,
    i_8_2_228_0, i_8_2_306_0, i_8_2_315_0, i_8_2_321_0, i_8_2_361_0,
    i_8_2_368_0, i_8_2_388_0, i_8_2_493_0, i_8_2_504_0, i_8_2_508_0,
    i_8_2_509_0, i_8_2_534_0, i_8_2_550_0, i_8_2_568_0, i_8_2_577_0,
    i_8_2_622_0, i_8_2_640_0, i_8_2_675_0, i_8_2_697_0, i_8_2_704_0,
    i_8_2_747_0, i_8_2_865_0, i_8_2_866_0, i_8_2_873_0, i_8_2_874_0,
    i_8_2_949_0, i_8_2_950_0, i_8_2_977_0, i_8_2_978_0, i_8_2_1009_0,
    i_8_2_1066_0, i_8_2_1074_0, i_8_2_1099_0, i_8_2_1127_0, i_8_2_1203_0,
    i_8_2_1228_0, i_8_2_1243_0, i_8_2_1263_0, i_8_2_1266_0, i_8_2_1268_0,
    i_8_2_1282_0, i_8_2_1301_0, i_8_2_1328_0, i_8_2_1360_0, i_8_2_1403_0,
    i_8_2_1433_0, i_8_2_1477_0, i_8_2_1479_0, i_8_2_1488_0, i_8_2_1513_0,
    i_8_2_1515_0, i_8_2_1545_0, i_8_2_1567_0, i_8_2_1577_0, i_8_2_1580_0,
    i_8_2_1595_0, i_8_2_1598_0, i_8_2_1632_0, i_8_2_1634_0, i_8_2_1651_0,
    i_8_2_1674_0, i_8_2_1701_0, i_8_2_1702_0, i_8_2_1747_0, i_8_2_1753_0,
    i_8_2_1756_0, i_8_2_1757_0, i_8_2_1773_0, i_8_2_1787_0, i_8_2_1790_0,
    i_8_2_1809_0, i_8_2_1810_0, i_8_2_1824_0, i_8_2_1837_0, i_8_2_1946_0,
    i_8_2_1949_0, i_8_2_1953_0, i_8_2_1954_0, i_8_2_1995_0, i_8_2_2038_0,
    i_8_2_2070_0, i_8_2_2097_0, i_8_2_2098_0, i_8_2_2142_0, i_8_2_2172_0,
    i_8_2_2227_0, i_8_2_2281_0, i_8_2_2288_0, i_8_2_2292_0,
    o_8_2_0_0  );
  input  i_8_2_2_0, i_8_2_11_0, i_8_2_40_0, i_8_2_55_0, i_8_2_73_0,
    i_8_2_101_0, i_8_2_135_0, i_8_2_181_0, i_8_2_192_0, i_8_2_195_0,
    i_8_2_225_0, i_8_2_228_0, i_8_2_306_0, i_8_2_315_0, i_8_2_321_0,
    i_8_2_361_0, i_8_2_368_0, i_8_2_388_0, i_8_2_493_0, i_8_2_504_0,
    i_8_2_508_0, i_8_2_509_0, i_8_2_534_0, i_8_2_550_0, i_8_2_568_0,
    i_8_2_577_0, i_8_2_622_0, i_8_2_640_0, i_8_2_675_0, i_8_2_697_0,
    i_8_2_704_0, i_8_2_747_0, i_8_2_865_0, i_8_2_866_0, i_8_2_873_0,
    i_8_2_874_0, i_8_2_949_0, i_8_2_950_0, i_8_2_977_0, i_8_2_978_0,
    i_8_2_1009_0, i_8_2_1066_0, i_8_2_1074_0, i_8_2_1099_0, i_8_2_1127_0,
    i_8_2_1203_0, i_8_2_1228_0, i_8_2_1243_0, i_8_2_1263_0, i_8_2_1266_0,
    i_8_2_1268_0, i_8_2_1282_0, i_8_2_1301_0, i_8_2_1328_0, i_8_2_1360_0,
    i_8_2_1403_0, i_8_2_1433_0, i_8_2_1477_0, i_8_2_1479_0, i_8_2_1488_0,
    i_8_2_1513_0, i_8_2_1515_0, i_8_2_1545_0, i_8_2_1567_0, i_8_2_1577_0,
    i_8_2_1580_0, i_8_2_1595_0, i_8_2_1598_0, i_8_2_1632_0, i_8_2_1634_0,
    i_8_2_1651_0, i_8_2_1674_0, i_8_2_1701_0, i_8_2_1702_0, i_8_2_1747_0,
    i_8_2_1753_0, i_8_2_1756_0, i_8_2_1757_0, i_8_2_1773_0, i_8_2_1787_0,
    i_8_2_1790_0, i_8_2_1809_0, i_8_2_1810_0, i_8_2_1824_0, i_8_2_1837_0,
    i_8_2_1946_0, i_8_2_1949_0, i_8_2_1953_0, i_8_2_1954_0, i_8_2_1995_0,
    i_8_2_2038_0, i_8_2_2070_0, i_8_2_2097_0, i_8_2_2098_0, i_8_2_2142_0,
    i_8_2_2172_0, i_8_2_2227_0, i_8_2_2281_0, i_8_2_2288_0, i_8_2_2292_0;
  output o_8_2_0_0;
  assign o_8_2_0_0 = 0;
endmodule



// Benchmark "kernel_8_3" written by ABC on Sun Jul 19 10:03:05 2020

module kernel_8_3 ( 
    i_8_3_72_0, i_8_3_103_0, i_8_3_126_0, i_8_3_147_0, i_8_3_202_0,
    i_8_3_208_0, i_8_3_262_0, i_8_3_273_0, i_8_3_275_0, i_8_3_318_0,
    i_8_3_378_0, i_8_3_383_0, i_8_3_397_0, i_8_3_420_0, i_8_3_441_0,
    i_8_3_476_0, i_8_3_492_0, i_8_3_507_0, i_8_3_514_0, i_8_3_577_0,
    i_8_3_580_0, i_8_3_630_0, i_8_3_665_0, i_8_3_668_0, i_8_3_679_0,
    i_8_3_702_0, i_8_3_800_0, i_8_3_838_0, i_8_3_841_0, i_8_3_847_0,
    i_8_3_910_0, i_8_3_926_0, i_8_3_948_0, i_8_3_955_0, i_8_3_966_0,
    i_8_3_1083_0, i_8_3_1111_0, i_8_3_1128_0, i_8_3_1153_0, i_8_3_1198_0,
    i_8_3_1224_0, i_8_3_1225_0, i_8_3_1269_0, i_8_3_1270_0, i_8_3_1281_0,
    i_8_3_1297_0, i_8_3_1335_0, i_8_3_1350_0, i_8_3_1385_0, i_8_3_1386_0,
    i_8_3_1387_0, i_8_3_1388_0, i_8_3_1405_0, i_8_3_1410_0, i_8_3_1461_0,
    i_8_3_1470_0, i_8_3_1478_0, i_8_3_1485_0, i_8_3_1494_0, i_8_3_1495_0,
    i_8_3_1521_0, i_8_3_1536_0, i_8_3_1537_0, i_8_3_1549_0, i_8_3_1650_0,
    i_8_3_1652_0, i_8_3_1675_0, i_8_3_1678_0, i_8_3_1686_0, i_8_3_1693_0,
    i_8_3_1701_0, i_8_3_1746_0, i_8_3_1747_0, i_8_3_1791_0, i_8_3_1803_0,
    i_8_3_1820_0, i_8_3_1821_0, i_8_3_1826_0, i_8_3_1841_0, i_8_3_1864_0,
    i_8_3_1926_0, i_8_3_1962_0, i_8_3_1992_0, i_8_3_2011_0, i_8_3_2044_0,
    i_8_3_2046_0, i_8_3_2136_0, i_8_3_2143_0, i_8_3_2149_0, i_8_3_2169_0,
    i_8_3_2170_0, i_8_3_2178_0, i_8_3_2226_0, i_8_3_2232_0, i_8_3_2234_0,
    i_8_3_2253_0, i_8_3_2256_0, i_8_3_2280_0, i_8_3_2295_0, i_8_3_2296_0,
    o_8_3_0_0  );
  input  i_8_3_72_0, i_8_3_103_0, i_8_3_126_0, i_8_3_147_0, i_8_3_202_0,
    i_8_3_208_0, i_8_3_262_0, i_8_3_273_0, i_8_3_275_0, i_8_3_318_0,
    i_8_3_378_0, i_8_3_383_0, i_8_3_397_0, i_8_3_420_0, i_8_3_441_0,
    i_8_3_476_0, i_8_3_492_0, i_8_3_507_0, i_8_3_514_0, i_8_3_577_0,
    i_8_3_580_0, i_8_3_630_0, i_8_3_665_0, i_8_3_668_0, i_8_3_679_0,
    i_8_3_702_0, i_8_3_800_0, i_8_3_838_0, i_8_3_841_0, i_8_3_847_0,
    i_8_3_910_0, i_8_3_926_0, i_8_3_948_0, i_8_3_955_0, i_8_3_966_0,
    i_8_3_1083_0, i_8_3_1111_0, i_8_3_1128_0, i_8_3_1153_0, i_8_3_1198_0,
    i_8_3_1224_0, i_8_3_1225_0, i_8_3_1269_0, i_8_3_1270_0, i_8_3_1281_0,
    i_8_3_1297_0, i_8_3_1335_0, i_8_3_1350_0, i_8_3_1385_0, i_8_3_1386_0,
    i_8_3_1387_0, i_8_3_1388_0, i_8_3_1405_0, i_8_3_1410_0, i_8_3_1461_0,
    i_8_3_1470_0, i_8_3_1478_0, i_8_3_1485_0, i_8_3_1494_0, i_8_3_1495_0,
    i_8_3_1521_0, i_8_3_1536_0, i_8_3_1537_0, i_8_3_1549_0, i_8_3_1650_0,
    i_8_3_1652_0, i_8_3_1675_0, i_8_3_1678_0, i_8_3_1686_0, i_8_3_1693_0,
    i_8_3_1701_0, i_8_3_1746_0, i_8_3_1747_0, i_8_3_1791_0, i_8_3_1803_0,
    i_8_3_1820_0, i_8_3_1821_0, i_8_3_1826_0, i_8_3_1841_0, i_8_3_1864_0,
    i_8_3_1926_0, i_8_3_1962_0, i_8_3_1992_0, i_8_3_2011_0, i_8_3_2044_0,
    i_8_3_2046_0, i_8_3_2136_0, i_8_3_2143_0, i_8_3_2149_0, i_8_3_2169_0,
    i_8_3_2170_0, i_8_3_2178_0, i_8_3_2226_0, i_8_3_2232_0, i_8_3_2234_0,
    i_8_3_2253_0, i_8_3_2256_0, i_8_3_2280_0, i_8_3_2295_0, i_8_3_2296_0;
  output o_8_3_0_0;
  assign o_8_3_0_0 = 0;
endmodule



// Benchmark "kernel_8_4" written by ABC on Sun Jul 19 10:03:07 2020

module kernel_8_4 ( 
    i_8_4_28_0, i_8_4_47_0, i_8_4_49_0, i_8_4_108_0, i_8_4_109_0,
    i_8_4_111_0, i_8_4_180_0, i_8_4_181_0, i_8_4_182_0, i_8_4_185_0,
    i_8_4_191_0, i_8_4_220_0, i_8_4_221_0, i_8_4_237_0, i_8_4_238_0,
    i_8_4_256_0, i_8_4_263_0, i_8_4_300_0, i_8_4_343_0, i_8_4_345_0,
    i_8_4_362_0, i_8_4_364_0, i_8_4_378_0, i_8_4_379_0, i_8_4_387_0,
    i_8_4_388_0, i_8_4_477_0, i_8_4_478_0, i_8_4_550_0, i_8_4_596_0,
    i_8_4_599_0, i_8_4_615_0, i_8_4_631_0, i_8_4_665_0, i_8_4_685_0,
    i_8_4_704_0, i_8_4_707_0, i_8_4_758_0, i_8_4_759_0, i_8_4_884_0,
    i_8_4_919_0, i_8_4_937_0, i_8_4_938_0, i_8_4_991_0, i_8_4_1089_0,
    i_8_4_1110_0, i_8_4_1117_0, i_8_4_1179_0, i_8_4_1180_0, i_8_4_1181_0,
    i_8_4_1189_0, i_8_4_1283_0, i_8_4_1288_0, i_8_4_1314_0, i_8_4_1334_0,
    i_8_4_1407_0, i_8_4_1409_0, i_8_4_1434_0, i_8_4_1435_0, i_8_4_1455_0,
    i_8_4_1467_0, i_8_4_1468_0, i_8_4_1476_0, i_8_4_1487_0, i_8_4_1506_0,
    i_8_4_1507_0, i_8_4_1542_0, i_8_4_1549_0, i_8_4_1554_0, i_8_4_1561_0,
    i_8_4_1631_0, i_8_4_1648_0, i_8_4_1651_0, i_8_4_1674_0, i_8_4_1675_0,
    i_8_4_1720_0, i_8_4_1724_0, i_8_4_1729_0, i_8_4_1739_0, i_8_4_1760_0,
    i_8_4_1778_0, i_8_4_1818_0, i_8_4_1819_0, i_8_4_1821_0, i_8_4_1827_0,
    i_8_4_1831_0, i_8_4_1857_0, i_8_4_1858_0, i_8_4_1864_0, i_8_4_1901_0,
    i_8_4_1948_0, i_8_4_1993_0, i_8_4_1996_0, i_8_4_2044_0, i_8_4_2143_0,
    i_8_4_2219_0, i_8_4_2245_0, i_8_4_2246_0, i_8_4_2281_0, i_8_4_2297_0,
    o_8_4_0_0  );
  input  i_8_4_28_0, i_8_4_47_0, i_8_4_49_0, i_8_4_108_0, i_8_4_109_0,
    i_8_4_111_0, i_8_4_180_0, i_8_4_181_0, i_8_4_182_0, i_8_4_185_0,
    i_8_4_191_0, i_8_4_220_0, i_8_4_221_0, i_8_4_237_0, i_8_4_238_0,
    i_8_4_256_0, i_8_4_263_0, i_8_4_300_0, i_8_4_343_0, i_8_4_345_0,
    i_8_4_362_0, i_8_4_364_0, i_8_4_378_0, i_8_4_379_0, i_8_4_387_0,
    i_8_4_388_0, i_8_4_477_0, i_8_4_478_0, i_8_4_550_0, i_8_4_596_0,
    i_8_4_599_0, i_8_4_615_0, i_8_4_631_0, i_8_4_665_0, i_8_4_685_0,
    i_8_4_704_0, i_8_4_707_0, i_8_4_758_0, i_8_4_759_0, i_8_4_884_0,
    i_8_4_919_0, i_8_4_937_0, i_8_4_938_0, i_8_4_991_0, i_8_4_1089_0,
    i_8_4_1110_0, i_8_4_1117_0, i_8_4_1179_0, i_8_4_1180_0, i_8_4_1181_0,
    i_8_4_1189_0, i_8_4_1283_0, i_8_4_1288_0, i_8_4_1314_0, i_8_4_1334_0,
    i_8_4_1407_0, i_8_4_1409_0, i_8_4_1434_0, i_8_4_1435_0, i_8_4_1455_0,
    i_8_4_1467_0, i_8_4_1468_0, i_8_4_1476_0, i_8_4_1487_0, i_8_4_1506_0,
    i_8_4_1507_0, i_8_4_1542_0, i_8_4_1549_0, i_8_4_1554_0, i_8_4_1561_0,
    i_8_4_1631_0, i_8_4_1648_0, i_8_4_1651_0, i_8_4_1674_0, i_8_4_1675_0,
    i_8_4_1720_0, i_8_4_1724_0, i_8_4_1729_0, i_8_4_1739_0, i_8_4_1760_0,
    i_8_4_1778_0, i_8_4_1818_0, i_8_4_1819_0, i_8_4_1821_0, i_8_4_1827_0,
    i_8_4_1831_0, i_8_4_1857_0, i_8_4_1858_0, i_8_4_1864_0, i_8_4_1901_0,
    i_8_4_1948_0, i_8_4_1993_0, i_8_4_1996_0, i_8_4_2044_0, i_8_4_2143_0,
    i_8_4_2219_0, i_8_4_2245_0, i_8_4_2246_0, i_8_4_2281_0, i_8_4_2297_0;
  output o_8_4_0_0;
  assign o_8_4_0_0 = ~((i_8_4_49_0 & ((i_8_4_665_0 & i_8_4_1409_0 & ~i_8_4_1434_0) | (~i_8_4_1110_0 & ~i_8_4_1554_0 & ~i_8_4_1720_0 & ~i_8_4_1760_0 & ~i_8_4_1858_0))) | (~i_8_4_49_0 & ((~i_8_4_237_0 & i_8_4_300_0 & ~i_8_4_685_0 & ~i_8_4_759_0 & ~i_8_4_1435_0 & ~i_8_4_1857_0) | (~i_8_4_477_0 & ~i_8_4_1288_0 & ~i_8_4_1760_0 & i_8_4_1819_0 & ~i_8_4_1948_0))) | (~i_8_4_1179_0 & ((~i_8_4_191_0 & ~i_8_4_1476_0 & ((~i_8_4_28_0 & i_8_4_345_0 & ~i_8_4_631_0 & ~i_8_4_1181_0 & i_8_4_1467_0) | (i_8_4_181_0 & ~i_8_4_938_0 & ~i_8_4_1554_0 & ~i_8_4_2044_0 & ~i_8_4_2281_0))) | (~i_8_4_1181_0 & ((i_8_4_47_0 & ~i_8_4_108_0 & ~i_8_4_1487_0) | (~i_8_4_550_0 & ~i_8_4_631_0 & i_8_4_685_0 & ~i_8_4_1110_0 & ~i_8_4_1674_0 & ~i_8_4_1858_0 & ~i_8_4_1901_0))) | (~i_8_4_1674_0 & ((i_8_4_109_0 & ~i_8_4_237_0 & ~i_8_4_345_0 & ~i_8_4_1334_0 & ~i_8_4_1435_0 & i_8_4_1858_0 & ~i_8_4_1993_0 & ~i_8_4_2219_0) | (~i_8_4_238_0 & i_8_4_379_0 & ~i_8_4_1675_0 & ~i_8_4_2297_0))) | (~i_8_4_111_0 & ~i_8_4_1434_0 & i_8_4_1821_0))) | (~i_8_4_28_0 & ((i_8_4_185_0 & ~i_8_4_1407_0) | (~i_8_4_47_0 & ~i_8_4_111_0 & ~i_8_4_238_0 & i_8_4_599_0 & ~i_8_4_884_0 & ~i_8_4_1857_0))) | (i_8_4_221_0 & ((i_8_4_362_0 & ~i_8_4_937_0 & ~i_8_4_938_0 & ~i_8_4_1554_0) | (~i_8_4_256_0 & ~i_8_4_685_0 & ~i_8_4_1180_0 & ~i_8_4_1181_0 & ~i_8_4_1542_0 & ~i_8_4_1857_0))) | (i_8_4_238_0 & ((~i_8_4_237_0 & i_8_4_300_0 & ~i_8_4_615_0 & ~i_8_4_685_0 & i_8_4_1435_0 & ~i_8_4_1760_0) | (i_8_4_1821_0 & i_8_4_1996_0))) | (i_8_4_345_0 & ((~i_8_4_221_0 & ~i_8_4_256_0 & ~i_8_4_478_0 & ~i_8_4_615_0 & ~i_8_4_1675_0) | (~i_8_4_387_0 & i_8_4_1821_0))) | (~i_8_4_256_0 & ((i_8_4_220_0 & ~i_8_4_237_0 & ~i_8_4_263_0 & ~i_8_4_685_0 & ~i_8_4_1110_0 & ~i_8_4_1739_0) | (i_8_4_378_0 & i_8_4_1993_0))) | (i_8_4_220_0 & ((~i_8_4_1181_0 & ~i_8_4_1314_0 & ~i_8_4_1760_0 & ~i_8_4_1827_0 & i_8_4_1948_0 & ~i_8_4_2044_0) | (~i_8_4_300_0 & ~i_8_4_1110_0 & ~i_8_4_1180_0 & ~i_8_4_1334_0 & ~i_8_4_1455_0 & ~i_8_4_1468_0 & ~i_8_4_1648_0 & ~i_8_4_2219_0))) | (~i_8_4_1334_0 & ((~i_8_4_263_0 & ((~i_8_4_345_0 & i_8_4_388_0 & ~i_8_4_665_0 & ~i_8_4_937_0 & ~i_8_4_1720_0 & i_8_4_1778_0) | (~i_8_4_108_0 & i_8_4_364_0 & ~i_8_4_685_0 & ~i_8_4_759_0 & ~i_8_4_1996_0 & ~i_8_4_2245_0))) | (~i_8_4_1434_0 & ((~i_8_4_1435_0 & i_8_4_1996_0) | (~i_8_4_237_0 & ~i_8_4_238_0 & ~i_8_4_665_0 & ~i_8_4_685_0 & ~i_8_4_1554_0 & ~i_8_4_1827_0 & ~i_8_4_1858_0 & ~i_8_4_2219_0 & ~i_8_4_2245_0))))) | (~i_8_4_665_0 & ((~i_8_4_938_0 & ~i_8_4_991_0 & ~i_8_4_1288_0 & ~i_8_4_1407_0 & ~i_8_4_1455_0 & ~i_8_4_1821_0 & ~i_8_4_1831_0 & i_8_4_1948_0) | (~i_8_4_108_0 & ~i_8_4_237_0 & ~i_8_4_238_0 & ~i_8_4_758_0 & ~i_8_4_1434_0 & ~i_8_4_1651_0 & ~i_8_4_1858_0 & ~i_8_4_2245_0))) | (~i_8_4_758_0 & ((~i_8_4_108_0 & ~i_8_4_2297_0 & ((i_8_4_379_0 & ~i_8_4_387_0 & ~i_8_4_615_0 & ~i_8_4_1110_0) | (~i_8_4_220_0 & ~i_8_4_300_0 & ~i_8_4_477_0 & ~i_8_4_1549_0 & i_8_4_1778_0))) | (~i_8_4_759_0 & ((~i_8_4_1089_0 & i_8_4_1409_0 & ~i_8_4_1435_0 & ~i_8_4_1455_0 & ~i_8_4_1554_0 & ~i_8_4_1724_0) | (~i_8_4_477_0 & ~i_8_4_938_0 & ~i_8_4_1110_0 & i_8_4_1283_0 & ~i_8_4_1651_0 & ~i_8_4_1821_0 & ~i_8_4_1831_0))))) | (~i_8_4_615_0 & ((~i_8_4_1407_0 & ~i_8_4_1435_0 & ~i_8_4_1831_0 & ~i_8_4_1996_0 & i_8_4_2245_0) | (~i_8_4_378_0 & ~i_8_4_1089_0 & i_8_4_1407_0 & ~i_8_4_1651_0 & ~i_8_4_2245_0))) | (~i_8_4_685_0 & ((i_8_4_1434_0 & i_8_4_1435_0 & ~i_8_4_1476_0 & ~i_8_4_1831_0 & i_8_4_2143_0) | (~i_8_4_220_0 & ~i_8_4_238_0 & ~i_8_4_1675_0 & i_8_4_1993_0 & ~i_8_4_2246_0))) | (~i_8_4_220_0 & ~i_8_4_1651_0 & ((~i_8_4_237_0 & i_8_4_665_0 & ~i_8_4_1409_0 & ~i_8_4_1554_0 & ~i_8_4_1760_0 & ~i_8_4_1858_0) | (i_8_4_2245_0 & i_8_4_2246_0 & ~i_8_4_2281_0))) | (~i_8_4_1434_0 & ((~i_8_4_237_0 & ((~i_8_4_238_0 & ~i_8_4_478_0 & ~i_8_4_937_0 & ~i_8_4_1283_0 & ~i_8_4_1435_0 & ~i_8_4_1739_0 & ~i_8_4_1827_0 & ~i_8_4_1831_0) | (~i_8_4_1110_0 & i_8_4_1651_0 & ~i_8_4_2245_0 & ~i_8_4_2297_0))) | (~i_8_4_300_0 & i_8_4_707_0 & ~i_8_4_1739_0))) | (i_8_4_1821_0 & ((~i_8_4_300_0 & ~i_8_4_478_0 & ((~i_8_4_477_0 & ~i_8_4_1110_0 & ~i_8_4_1407_0) | (i_8_4_1407_0 & ~i_8_4_1455_0))) | (i_8_4_111_0 & ~i_8_4_991_0 & ~i_8_4_1110_0) | (~i_8_4_111_0 & ~i_8_4_238_0 & ~i_8_4_477_0 & ~i_8_4_1857_0))) | (~i_8_4_991_0 & ((i_8_4_478_0 & i_8_4_1561_0 & ~i_8_4_1948_0 & ~i_8_4_2219_0) | (i_8_4_364_0 & ~i_8_4_759_0 & ~i_8_4_1561_0 & ~i_8_4_2044_0 & i_8_4_2245_0))) | (~i_8_4_1729_0 & ((~i_8_4_477_0 & i_8_4_1818_0 & ~i_8_4_1858_0) | (~i_8_4_109_0 & i_8_4_1858_0 & i_8_4_2143_0))) | (i_8_4_1818_0 & ((i_8_4_387_0 & i_8_4_1549_0) | (~i_8_4_759_0 & ~i_8_4_1549_0 & ~i_8_4_1561_0 & i_8_4_1858_0))) | (~i_8_4_759_0 & ((i_8_4_1542_0 & ~i_8_4_1858_0) | (i_8_4_237_0 & ~i_8_4_300_0 & ~i_8_4_345_0 & i_8_4_1554_0 & i_8_4_1651_0 & ~i_8_4_1675_0 & ~i_8_4_2219_0) | (i_8_4_1506_0 & i_8_4_1996_0 & ~i_8_4_2297_0))) | (i_8_4_1314_0 & i_8_4_2219_0 & i_8_4_2281_0));
endmodule



// Benchmark "kernel_8_5" written by ABC on Sun Jul 19 10:03:07 2020

module kernel_8_5 ( 
    i_8_5_3_0, i_8_5_66_0, i_8_5_67_0, i_8_5_79_0, i_8_5_84_0, i_8_5_85_0,
    i_8_5_190_0, i_8_5_193_0, i_8_5_210_0, i_8_5_223_0, i_8_5_238_0,
    i_8_5_361_0, i_8_5_364_0, i_8_5_414_0, i_8_5_481_0, i_8_5_498_0,
    i_8_5_516_0, i_8_5_517_0, i_8_5_525_0, i_8_5_582_0, i_8_5_603_0,
    i_8_5_612_0, i_8_5_615_0, i_8_5_624_0, i_8_5_625_0, i_8_5_636_0,
    i_8_5_672_0, i_8_5_705_0, i_8_5_708_0, i_8_5_760_0, i_8_5_789_0,
    i_8_5_795_0, i_8_5_814_0, i_8_5_835_0, i_8_5_843_0, i_8_5_844_0,
    i_8_5_858_0, i_8_5_937_0, i_8_5_959_0, i_8_5_999_0, i_8_5_1002_0,
    i_8_5_1057_0, i_8_5_1059_0, i_8_5_1074_0, i_8_5_1114_0, i_8_5_1141_0,
    i_8_5_1168_0, i_8_5_1182_0, i_8_5_1183_0, i_8_5_1192_0, i_8_5_1219_0,
    i_8_5_1227_0, i_8_5_1236_0, i_8_5_1237_0, i_8_5_1239_0, i_8_5_1249_0,
    i_8_5_1275_0, i_8_5_1286_0, i_8_5_1300_0, i_8_5_1345_0, i_8_5_1348_0,
    i_8_5_1382_0, i_8_5_1407_0, i_8_5_1410_0, i_8_5_1497_0, i_8_5_1530_0,
    i_8_5_1533_0, i_8_5_1633_0, i_8_5_1650_0, i_8_5_1668_0, i_8_5_1689_0,
    i_8_5_1704_0, i_8_5_1741_0, i_8_5_1764_0, i_8_5_1818_0, i_8_5_1821_0,
    i_8_5_1839_0, i_8_5_1848_0, i_8_5_1857_0, i_8_5_1884_0, i_8_5_1885_0,
    i_8_5_1888_0, i_8_5_1896_0, i_8_5_2011_0, i_8_5_2037_0, i_8_5_2044_0,
    i_8_5_2047_0, i_8_5_2065_0, i_8_5_2104_0, i_8_5_2118_0, i_8_5_2119_0,
    i_8_5_2122_0, i_8_5_2146_0, i_8_5_2169_0, i_8_5_2174_0, i_8_5_2211_0,
    i_8_5_2214_0, i_8_5_2257_0, i_8_5_2290_0, i_8_5_2299_0,
    o_8_5_0_0  );
  input  i_8_5_3_0, i_8_5_66_0, i_8_5_67_0, i_8_5_79_0, i_8_5_84_0,
    i_8_5_85_0, i_8_5_190_0, i_8_5_193_0, i_8_5_210_0, i_8_5_223_0,
    i_8_5_238_0, i_8_5_361_0, i_8_5_364_0, i_8_5_414_0, i_8_5_481_0,
    i_8_5_498_0, i_8_5_516_0, i_8_5_517_0, i_8_5_525_0, i_8_5_582_0,
    i_8_5_603_0, i_8_5_612_0, i_8_5_615_0, i_8_5_624_0, i_8_5_625_0,
    i_8_5_636_0, i_8_5_672_0, i_8_5_705_0, i_8_5_708_0, i_8_5_760_0,
    i_8_5_789_0, i_8_5_795_0, i_8_5_814_0, i_8_5_835_0, i_8_5_843_0,
    i_8_5_844_0, i_8_5_858_0, i_8_5_937_0, i_8_5_959_0, i_8_5_999_0,
    i_8_5_1002_0, i_8_5_1057_0, i_8_5_1059_0, i_8_5_1074_0, i_8_5_1114_0,
    i_8_5_1141_0, i_8_5_1168_0, i_8_5_1182_0, i_8_5_1183_0, i_8_5_1192_0,
    i_8_5_1219_0, i_8_5_1227_0, i_8_5_1236_0, i_8_5_1237_0, i_8_5_1239_0,
    i_8_5_1249_0, i_8_5_1275_0, i_8_5_1286_0, i_8_5_1300_0, i_8_5_1345_0,
    i_8_5_1348_0, i_8_5_1382_0, i_8_5_1407_0, i_8_5_1410_0, i_8_5_1497_0,
    i_8_5_1530_0, i_8_5_1533_0, i_8_5_1633_0, i_8_5_1650_0, i_8_5_1668_0,
    i_8_5_1689_0, i_8_5_1704_0, i_8_5_1741_0, i_8_5_1764_0, i_8_5_1818_0,
    i_8_5_1821_0, i_8_5_1839_0, i_8_5_1848_0, i_8_5_1857_0, i_8_5_1884_0,
    i_8_5_1885_0, i_8_5_1888_0, i_8_5_1896_0, i_8_5_2011_0, i_8_5_2037_0,
    i_8_5_2044_0, i_8_5_2047_0, i_8_5_2065_0, i_8_5_2104_0, i_8_5_2118_0,
    i_8_5_2119_0, i_8_5_2122_0, i_8_5_2146_0, i_8_5_2169_0, i_8_5_2174_0,
    i_8_5_2211_0, i_8_5_2214_0, i_8_5_2257_0, i_8_5_2290_0, i_8_5_2299_0;
  output o_8_5_0_0;
  assign o_8_5_0_0 = 0;
endmodule



// Benchmark "kernel_8_6" written by ABC on Sun Jul 19 10:03:09 2020

module kernel_8_6 ( 
    i_8_6_12_0, i_8_6_37_0, i_8_6_40_0, i_8_6_50_0, i_8_6_57_0, i_8_6_64_0,
    i_8_6_68_0, i_8_6_256_0, i_8_6_262_0, i_8_6_305_0, i_8_6_319_0,
    i_8_6_381_0, i_8_6_382_0, i_8_6_391_0, i_8_6_435_0, i_8_6_453_0,
    i_8_6_454_0, i_8_6_460_0, i_8_6_486_0, i_8_6_490_0, i_8_6_504_0,
    i_8_6_622_0, i_8_6_662_0, i_8_6_665_0, i_8_6_684_0, i_8_6_693_0,
    i_8_6_695_0, i_8_6_698_0, i_8_6_708_0, i_8_6_748_0, i_8_6_844_0,
    i_8_6_874_0, i_8_6_875_0, i_8_6_877_0, i_8_6_895_0, i_8_6_990_0,
    i_8_6_993_0, i_8_6_1034_0, i_8_6_1051_0, i_8_6_1054_0, i_8_6_1071_0,
    i_8_6_1114_0, i_8_6_1136_0, i_8_6_1198_0, i_8_6_1201_0, i_8_6_1225_0,
    i_8_6_1236_0, i_8_6_1237_0, i_8_6_1264_0, i_8_6_1265_0, i_8_6_1276_0,
    i_8_6_1282_0, i_8_6_1296_0, i_8_6_1328_0, i_8_6_1335_0, i_8_6_1354_0,
    i_8_6_1381_0, i_8_6_1383_0, i_8_6_1399_0, i_8_6_1404_0, i_8_6_1438_0,
    i_8_6_1461_0, i_8_6_1462_0, i_8_6_1486_0, i_8_6_1515_0, i_8_6_1530_0,
    i_8_6_1550_0, i_8_6_1623_0, i_8_6_1631_0, i_8_6_1632_0, i_8_6_1702_0,
    i_8_6_1746_0, i_8_6_1748_0, i_8_6_1754_0, i_8_6_1776_0, i_8_6_1791_0,
    i_8_6_1795_0, i_8_6_1812_0, i_8_6_1822_0, i_8_6_1836_0, i_8_6_1882_0,
    i_8_6_1903_0, i_8_6_1909_0, i_8_6_1911_0, i_8_6_1913_0, i_8_6_1936_0,
    i_8_6_1980_0, i_8_6_1992_0, i_8_6_1994_0, i_8_6_2038_0, i_8_6_2043_0,
    i_8_6_2044_0, i_8_6_2048_0, i_8_6_2055_0, i_8_6_2070_0, i_8_6_2106_0,
    i_8_6_2110_0, i_8_6_2142_0, i_8_6_2144_0, i_8_6_2296_0,
    o_8_6_0_0  );
  input  i_8_6_12_0, i_8_6_37_0, i_8_6_40_0, i_8_6_50_0, i_8_6_57_0,
    i_8_6_64_0, i_8_6_68_0, i_8_6_256_0, i_8_6_262_0, i_8_6_305_0,
    i_8_6_319_0, i_8_6_381_0, i_8_6_382_0, i_8_6_391_0, i_8_6_435_0,
    i_8_6_453_0, i_8_6_454_0, i_8_6_460_0, i_8_6_486_0, i_8_6_490_0,
    i_8_6_504_0, i_8_6_622_0, i_8_6_662_0, i_8_6_665_0, i_8_6_684_0,
    i_8_6_693_0, i_8_6_695_0, i_8_6_698_0, i_8_6_708_0, i_8_6_748_0,
    i_8_6_844_0, i_8_6_874_0, i_8_6_875_0, i_8_6_877_0, i_8_6_895_0,
    i_8_6_990_0, i_8_6_993_0, i_8_6_1034_0, i_8_6_1051_0, i_8_6_1054_0,
    i_8_6_1071_0, i_8_6_1114_0, i_8_6_1136_0, i_8_6_1198_0, i_8_6_1201_0,
    i_8_6_1225_0, i_8_6_1236_0, i_8_6_1237_0, i_8_6_1264_0, i_8_6_1265_0,
    i_8_6_1276_0, i_8_6_1282_0, i_8_6_1296_0, i_8_6_1328_0, i_8_6_1335_0,
    i_8_6_1354_0, i_8_6_1381_0, i_8_6_1383_0, i_8_6_1399_0, i_8_6_1404_0,
    i_8_6_1438_0, i_8_6_1461_0, i_8_6_1462_0, i_8_6_1486_0, i_8_6_1515_0,
    i_8_6_1530_0, i_8_6_1550_0, i_8_6_1623_0, i_8_6_1631_0, i_8_6_1632_0,
    i_8_6_1702_0, i_8_6_1746_0, i_8_6_1748_0, i_8_6_1754_0, i_8_6_1776_0,
    i_8_6_1791_0, i_8_6_1795_0, i_8_6_1812_0, i_8_6_1822_0, i_8_6_1836_0,
    i_8_6_1882_0, i_8_6_1903_0, i_8_6_1909_0, i_8_6_1911_0, i_8_6_1913_0,
    i_8_6_1936_0, i_8_6_1980_0, i_8_6_1992_0, i_8_6_1994_0, i_8_6_2038_0,
    i_8_6_2043_0, i_8_6_2044_0, i_8_6_2048_0, i_8_6_2055_0, i_8_6_2070_0,
    i_8_6_2106_0, i_8_6_2110_0, i_8_6_2142_0, i_8_6_2144_0, i_8_6_2296_0;
  output o_8_6_0_0;
  assign o_8_6_0_0 = ~((~i_8_6_460_0 & ((~i_8_6_12_0 & ((~i_8_6_40_0 & ~i_8_6_391_0 & ~i_8_6_1702_0 & ~i_8_6_1911_0 & ~i_8_6_2043_0) | (~i_8_6_504_0 & ~i_8_6_1034_0 & ~i_8_6_1201_0 & ~i_8_6_1383_0 & ~i_8_6_1461_0 & ~i_8_6_2044_0 & ~i_8_6_2048_0))) | (~i_8_6_40_0 & ~i_8_6_504_0 & ((~i_8_6_262_0 & ~i_8_6_1201_0 & ~i_8_6_1225_0 & ~i_8_6_1748_0 & ~i_8_6_1909_0 & ~i_8_6_1911_0) | (~i_8_6_319_0 & ~i_8_6_665_0 & i_8_6_1265_0 & ~i_8_6_1461_0 & ~i_8_6_2142_0))) | (~i_8_6_1911_0 & ((~i_8_6_37_0 & ~i_8_6_708_0 & ~i_8_6_748_0 & ~i_8_6_895_0 & ~i_8_6_1791_0 & ~i_8_6_1795_0 & ~i_8_6_1913_0) | (~i_8_6_1054_0 & ~i_8_6_1530_0 & ~i_8_6_1702_0 & ~i_8_6_1746_0 & ~i_8_6_1776_0 & ~i_8_6_1936_0 & ~i_8_6_2048_0))))) | (~i_8_6_68_0 & ((~i_8_6_40_0 & ((~i_8_6_256_0 & ~i_8_6_262_0 & ~i_8_6_504_0 & ~i_8_6_1383_0 & ~i_8_6_1702_0 & ~i_8_6_1812_0 & ~i_8_6_1909_0) | (~i_8_6_844_0 & ~i_8_6_1198_0 & ~i_8_6_1296_0 & i_8_6_1994_0 & ~i_8_6_2106_0))) | (~i_8_6_391_0 & ~i_8_6_1335_0 & ~i_8_6_1354_0 & ~i_8_6_1632_0 & ~i_8_6_1702_0 & ~i_8_6_1795_0 & ~i_8_6_2296_0))) | (~i_8_6_57_0 & ~i_8_6_708_0 & ((~i_8_6_381_0 & ~i_8_6_1071_0 & ~i_8_6_1201_0 & ~i_8_6_1383_0 & ~i_8_6_1791_0 & ~i_8_6_1882_0) | (~i_8_6_435_0 & ~i_8_6_1530_0 & ~i_8_6_1550_0 & ~i_8_6_1836_0 & ~i_8_6_1994_0 & ~i_8_6_2044_0))) | (~i_8_6_1992_0 & ((~i_8_6_64_0 & ~i_8_6_1461_0 & ((~i_8_6_37_0 & ~i_8_6_1237_0 & ~i_8_6_1631_0 & ~i_8_6_1909_0 & ~i_8_6_1911_0) | (~i_8_6_319_0 & ~i_8_6_1071_0 & ~i_8_6_1276_0 & ~i_8_6_1913_0 & ~i_8_6_2043_0 & ~i_8_6_2070_0 & ~i_8_6_2296_0))) | (~i_8_6_50_0 & i_8_6_1114_0 & ~i_8_6_1264_0 & ~i_8_6_1265_0 & ~i_8_6_1354_0))) | (~i_8_6_319_0 & ~i_8_6_2038_0 & ((~i_8_6_622_0 & ~i_8_6_1265_0 & ~i_8_6_1354_0 & ~i_8_6_1486_0 & ~i_8_6_1530_0 & ~i_8_6_1911_0) | (~i_8_6_381_0 & ~i_8_6_1237_0 & ~i_8_6_1264_0 & ~i_8_6_1791_0 & ~i_8_6_2043_0 & ~i_8_6_2044_0))) | (~i_8_6_1795_0 & ((~i_8_6_1909_0 & ((~i_8_6_435_0 & i_8_6_993_0 & ~i_8_6_1201_0 & ~i_8_6_1882_0) | (~i_8_6_1198_0 & ~i_8_6_1404_0 & ~i_8_6_1462_0 & ~i_8_6_1515_0 & ~i_8_6_1748_0 & ~i_8_6_1791_0 & ~i_8_6_2142_0))) | (~i_8_6_391_0 & ~i_8_6_748_0 & ~i_8_6_1276_0 & ~i_8_6_1399_0 & ~i_8_6_1776_0 & ~i_8_6_2043_0))) | (i_8_6_50_0 & i_8_6_1903_0 & ~i_8_6_2296_0));
endmodule



// Benchmark "kernel_8_7" written by ABC on Sun Jul 19 10:03:10 2020

module kernel_8_7 ( 
    i_8_7_12_0, i_8_7_13_0, i_8_7_46_0, i_8_7_52_0, i_8_7_78_0,
    i_8_7_139_0, i_8_7_159_0, i_8_7_211_0, i_8_7_237_0, i_8_7_262_0,
    i_8_7_264_0, i_8_7_265_0, i_8_7_285_0, i_8_7_322_0, i_8_7_328_0,
    i_8_7_336_0, i_8_7_337_0, i_8_7_381_0, i_8_7_384_0, i_8_7_400_0,
    i_8_7_417_0, i_8_7_420_0, i_8_7_421_0, i_8_7_471_0, i_8_7_510_0,
    i_8_7_556_0, i_8_7_573_0, i_8_7_574_0, i_8_7_580_0, i_8_7_660_0,
    i_8_7_687_0, i_8_7_688_0, i_8_7_697_0, i_8_7_753_0, i_8_7_807_0,
    i_8_7_822_0, i_8_7_894_0, i_8_7_895_0, i_8_7_898_0, i_8_7_919_0,
    i_8_7_966_0, i_8_7_975_0, i_8_7_976_0, i_8_7_1011_0, i_8_7_1012_0,
    i_8_7_1039_0, i_8_7_1041_0, i_8_7_1110_0, i_8_7_1113_0, i_8_7_1114_0,
    i_8_7_1239_0, i_8_7_1249_0, i_8_7_1260_0, i_8_7_1263_0, i_8_7_1267_0,
    i_8_7_1272_0, i_8_7_1273_0, i_8_7_1275_0, i_8_7_1282_0, i_8_7_1302_0,
    i_8_7_1303_0, i_8_7_1314_0, i_8_7_1315_0, i_8_7_1335_0, i_8_7_1338_0,
    i_8_7_1425_0, i_8_7_1426_0, i_8_7_1434_0, i_8_7_1437_0, i_8_7_1467_0,
    i_8_7_1510_0, i_8_7_1524_0, i_8_7_1525_0, i_8_7_1527_0, i_8_7_1528_0,
    i_8_7_1551_0, i_8_7_1554_0, i_8_7_1560_0, i_8_7_1572_0, i_8_7_1632_0,
    i_8_7_1668_0, i_8_7_1669_0, i_8_7_1722_0, i_8_7_1723_0, i_8_7_1726_0,
    i_8_7_1749_0, i_8_7_1768_0, i_8_7_1783_0, i_8_7_1797_0, i_8_7_1900_0,
    i_8_7_1939_0, i_8_7_1959_0, i_8_7_1969_0, i_8_7_1993_0, i_8_7_2154_0,
    i_8_7_2176_0, i_8_7_2229_0, i_8_7_2246_0, i_8_7_2249_0, i_8_7_2294_0,
    o_8_7_0_0  );
  input  i_8_7_12_0, i_8_7_13_0, i_8_7_46_0, i_8_7_52_0, i_8_7_78_0,
    i_8_7_139_0, i_8_7_159_0, i_8_7_211_0, i_8_7_237_0, i_8_7_262_0,
    i_8_7_264_0, i_8_7_265_0, i_8_7_285_0, i_8_7_322_0, i_8_7_328_0,
    i_8_7_336_0, i_8_7_337_0, i_8_7_381_0, i_8_7_384_0, i_8_7_400_0,
    i_8_7_417_0, i_8_7_420_0, i_8_7_421_0, i_8_7_471_0, i_8_7_510_0,
    i_8_7_556_0, i_8_7_573_0, i_8_7_574_0, i_8_7_580_0, i_8_7_660_0,
    i_8_7_687_0, i_8_7_688_0, i_8_7_697_0, i_8_7_753_0, i_8_7_807_0,
    i_8_7_822_0, i_8_7_894_0, i_8_7_895_0, i_8_7_898_0, i_8_7_919_0,
    i_8_7_966_0, i_8_7_975_0, i_8_7_976_0, i_8_7_1011_0, i_8_7_1012_0,
    i_8_7_1039_0, i_8_7_1041_0, i_8_7_1110_0, i_8_7_1113_0, i_8_7_1114_0,
    i_8_7_1239_0, i_8_7_1249_0, i_8_7_1260_0, i_8_7_1263_0, i_8_7_1267_0,
    i_8_7_1272_0, i_8_7_1273_0, i_8_7_1275_0, i_8_7_1282_0, i_8_7_1302_0,
    i_8_7_1303_0, i_8_7_1314_0, i_8_7_1315_0, i_8_7_1335_0, i_8_7_1338_0,
    i_8_7_1425_0, i_8_7_1426_0, i_8_7_1434_0, i_8_7_1437_0, i_8_7_1467_0,
    i_8_7_1510_0, i_8_7_1524_0, i_8_7_1525_0, i_8_7_1527_0, i_8_7_1528_0,
    i_8_7_1551_0, i_8_7_1554_0, i_8_7_1560_0, i_8_7_1572_0, i_8_7_1632_0,
    i_8_7_1668_0, i_8_7_1669_0, i_8_7_1722_0, i_8_7_1723_0, i_8_7_1726_0,
    i_8_7_1749_0, i_8_7_1768_0, i_8_7_1783_0, i_8_7_1797_0, i_8_7_1900_0,
    i_8_7_1939_0, i_8_7_1959_0, i_8_7_1969_0, i_8_7_1993_0, i_8_7_2154_0,
    i_8_7_2176_0, i_8_7_2229_0, i_8_7_2246_0, i_8_7_2249_0, i_8_7_2294_0;
  output o_8_7_0_0;
  assign o_8_7_0_0 = ~((~i_8_7_574_0 & ((~i_8_7_13_0 & ((~i_8_7_159_0 & ~i_8_7_919_0 & ~i_8_7_1425_0 & i_8_7_1434_0 & ~i_8_7_1669_0 & ~i_8_7_1783_0 & ~i_8_7_1797_0) | (~i_8_7_52_0 & ~i_8_7_237_0 & ~i_8_7_556_0 & ~i_8_7_580_0 & ~i_8_7_975_0 & ~i_8_7_1338_0 & ~i_8_7_1527_0 & ~i_8_7_2294_0))) | (~i_8_7_265_0 & ~i_8_7_322_0 & ~i_8_7_336_0 & ~i_8_7_337_0 & ~i_8_7_400_0 & ~i_8_7_807_0 & ~i_8_7_1012_0 & ~i_8_7_1282_0 & ~i_8_7_1572_0) | (~i_8_7_139_0 & ~i_8_7_328_0 & ~i_8_7_822_0 & ~i_8_7_898_0 & ~i_8_7_1338_0 & ~i_8_7_1528_0 & ~i_8_7_1668_0 & ~i_8_7_1783_0 & ~i_8_7_1900_0))) | (~i_8_7_46_0 & ((~i_8_7_421_0 & ~i_8_7_895_0 & i_8_7_1510_0 & ~i_8_7_1797_0) | (~i_8_7_265_0 & ~i_8_7_580_0 & i_8_7_753_0 & ~i_8_7_975_0 & i_8_7_1554_0 & ~i_8_7_1572_0 & ~i_8_7_1669_0 & ~i_8_7_2249_0))) | (~i_8_7_1524_0 & ((~i_8_7_211_0 & ((~i_8_7_322_0 & ~i_8_7_400_0 & ~i_8_7_660_0 & ~i_8_7_822_0 & ~i_8_7_1426_0 & ~i_8_7_1437_0 & ~i_8_7_1722_0) | (~i_8_7_894_0 & ~i_8_7_1110_0 & ~i_8_7_1113_0 & ~i_8_7_1314_0 & ~i_8_7_1527_0 & ~i_8_7_1669_0 & ~i_8_7_1939_0 & ~i_8_7_1959_0))) | (~i_8_7_262_0 & ~i_8_7_400_0 & ((~i_8_7_337_0 & ~i_8_7_421_0 & ~i_8_7_573_0 & ~i_8_7_1528_0 & ~i_8_7_1783_0) | (~i_8_7_159_0 & ~i_8_7_898_0 & ~i_8_7_1426_0 & ~i_8_7_1525_0 & ~i_8_7_1669_0 & ~i_8_7_1797_0 & ~i_8_7_2229_0 & ~i_8_7_2246_0))) | (~i_8_7_52_0 & ~i_8_7_264_0 & ~i_8_7_976_0 & ~i_8_7_1260_0 & ~i_8_7_1273_0 & ~i_8_7_1510_0 & ~i_8_7_1525_0 & ~i_8_7_1528_0 & i_8_7_1993_0))) | (~i_8_7_265_0 & ((~i_8_7_400_0 & ~i_8_7_660_0 & ~i_8_7_822_0 & ~i_8_7_895_0 & ~i_8_7_1041_0 & ~i_8_7_1669_0 & ~i_8_7_1768_0 & ~i_8_7_1900_0 & ~i_8_7_1993_0) | (~i_8_7_285_0 & ~i_8_7_322_0 & ~i_8_7_556_0 & i_8_7_1282_0 & ~i_8_7_1632_0 & ~i_8_7_1797_0 & ~i_8_7_2249_0))) | (~i_8_7_894_0 & ((~i_8_7_264_0 & ~i_8_7_895_0 & ~i_8_7_976_0 & ~i_8_7_1425_0 & ~i_8_7_1426_0 & ~i_8_7_1527_0 & ~i_8_7_1528_0 & ~i_8_7_1722_0 & ~i_8_7_1939_0) | (~i_8_7_381_0 & ~i_8_7_510_0 & ~i_8_7_898_0 & ~i_8_7_975_0 & ~i_8_7_1302_0 & ~i_8_7_1723_0 & ~i_8_7_1749_0 & ~i_8_7_1797_0 & ~i_8_7_1959_0))) | (~i_8_7_895_0 & ((~i_8_7_976_0 & ((~i_8_7_12_0 & ~i_8_7_556_0 & ~i_8_7_753_0 & ~i_8_7_898_0 & ~i_8_7_1011_0) | (~i_8_7_322_0 & i_8_7_1272_0 & ~i_8_7_1315_0 & ~i_8_7_1726_0))) | (~i_8_7_285_0 & ~i_8_7_417_0 & ~i_8_7_573_0 & ~i_8_7_1039_0 & ~i_8_7_1551_0 & ~i_8_7_1668_0 & ~i_8_7_1723_0))));
endmodule



// Benchmark "kernel_8_8" written by ABC on Sun Jul 19 10:03:10 2020

module kernel_8_8 ( 
    i_8_8_31_0, i_8_8_40_0, i_8_8_54_0, i_8_8_57_0, i_8_8_88_0,
    i_8_8_111_0, i_8_8_112_0, i_8_8_153_0, i_8_8_165_0, i_8_8_226_0,
    i_8_8_241_0, i_8_8_333_0, i_8_8_335_0, i_8_8_348_0, i_8_8_372_0,
    i_8_8_375_0, i_8_8_376_0, i_8_8_450_0, i_8_8_454_0, i_8_8_469_0,
    i_8_8_523_0, i_8_8_525_0, i_8_8_529_0, i_8_8_530_0, i_8_8_540_0,
    i_8_8_543_0, i_8_8_551_0, i_8_8_556_0, i_8_8_570_0, i_8_8_571_0,
    i_8_8_613_0, i_8_8_616_0, i_8_8_687_0, i_8_8_688_0, i_8_8_705_0,
    i_8_8_706_0, i_8_8_775_0, i_8_8_777_0, i_8_8_786_0, i_8_8_800_0,
    i_8_8_810_0, i_8_8_814_0, i_8_8_844_0, i_8_8_850_0, i_8_8_858_0,
    i_8_8_916_0, i_8_8_1056_0, i_8_8_1113_0, i_8_8_1114_0, i_8_8_1115_0,
    i_8_8_1124_0, i_8_8_1160_0, i_8_8_1182_0, i_8_8_1240_0, i_8_8_1267_0,
    i_8_8_1291_0, i_8_8_1292_0, i_8_8_1299_0, i_8_8_1308_0, i_8_8_1317_0,
    i_8_8_1323_0, i_8_8_1407_0, i_8_8_1490_0, i_8_8_1588_0, i_8_8_1596_0,
    i_8_8_1630_0, i_8_8_1651_0, i_8_8_1653_0, i_8_8_1654_0, i_8_8_1671_0,
    i_8_8_1696_0, i_8_8_1719_0, i_8_8_1722_0, i_8_8_1737_0, i_8_8_1741_0,
    i_8_8_1745_0, i_8_8_1749_0, i_8_8_1790_0, i_8_8_1840_0, i_8_8_1847_0,
    i_8_8_1856_0, i_8_8_1857_0, i_8_8_1884_0, i_8_8_1888_0, i_8_8_1946_0,
    i_8_8_1993_0, i_8_8_1997_0, i_8_8_2020_0, i_8_8_2022_0, i_8_8_2023_0,
    i_8_8_2037_0, i_8_8_2043_0, i_8_8_2044_0, i_8_8_2047_0, i_8_8_2050_0,
    i_8_8_2092_0, i_8_8_2123_0, i_8_8_2172_0, i_8_8_2233_0, i_8_8_2299_0,
    o_8_8_0_0  );
  input  i_8_8_31_0, i_8_8_40_0, i_8_8_54_0, i_8_8_57_0, i_8_8_88_0,
    i_8_8_111_0, i_8_8_112_0, i_8_8_153_0, i_8_8_165_0, i_8_8_226_0,
    i_8_8_241_0, i_8_8_333_0, i_8_8_335_0, i_8_8_348_0, i_8_8_372_0,
    i_8_8_375_0, i_8_8_376_0, i_8_8_450_0, i_8_8_454_0, i_8_8_469_0,
    i_8_8_523_0, i_8_8_525_0, i_8_8_529_0, i_8_8_530_0, i_8_8_540_0,
    i_8_8_543_0, i_8_8_551_0, i_8_8_556_0, i_8_8_570_0, i_8_8_571_0,
    i_8_8_613_0, i_8_8_616_0, i_8_8_687_0, i_8_8_688_0, i_8_8_705_0,
    i_8_8_706_0, i_8_8_775_0, i_8_8_777_0, i_8_8_786_0, i_8_8_800_0,
    i_8_8_810_0, i_8_8_814_0, i_8_8_844_0, i_8_8_850_0, i_8_8_858_0,
    i_8_8_916_0, i_8_8_1056_0, i_8_8_1113_0, i_8_8_1114_0, i_8_8_1115_0,
    i_8_8_1124_0, i_8_8_1160_0, i_8_8_1182_0, i_8_8_1240_0, i_8_8_1267_0,
    i_8_8_1291_0, i_8_8_1292_0, i_8_8_1299_0, i_8_8_1308_0, i_8_8_1317_0,
    i_8_8_1323_0, i_8_8_1407_0, i_8_8_1490_0, i_8_8_1588_0, i_8_8_1596_0,
    i_8_8_1630_0, i_8_8_1651_0, i_8_8_1653_0, i_8_8_1654_0, i_8_8_1671_0,
    i_8_8_1696_0, i_8_8_1719_0, i_8_8_1722_0, i_8_8_1737_0, i_8_8_1741_0,
    i_8_8_1745_0, i_8_8_1749_0, i_8_8_1790_0, i_8_8_1840_0, i_8_8_1847_0,
    i_8_8_1856_0, i_8_8_1857_0, i_8_8_1884_0, i_8_8_1888_0, i_8_8_1946_0,
    i_8_8_1993_0, i_8_8_1997_0, i_8_8_2020_0, i_8_8_2022_0, i_8_8_2023_0,
    i_8_8_2037_0, i_8_8_2043_0, i_8_8_2044_0, i_8_8_2047_0, i_8_8_2050_0,
    i_8_8_2092_0, i_8_8_2123_0, i_8_8_2172_0, i_8_8_2233_0, i_8_8_2299_0;
  output o_8_8_0_0;
  assign o_8_8_0_0 = 0;
endmodule



// Benchmark "kernel_8_9" written by ABC on Sun Jul 19 10:03:11 2020

module kernel_8_9 ( 
    i_8_9_46_0, i_8_9_58_0, i_8_9_59_0, i_8_9_85_0, i_8_9_87_0, i_8_9_88_0,
    i_8_9_106_0, i_8_9_140_0, i_8_9_142_0, i_8_9_143_0, i_8_9_187_0,
    i_8_9_188_0, i_8_9_252_0, i_8_9_256_0, i_8_9_259_0, i_8_9_303_0,
    i_8_9_304_0, i_8_9_311_0, i_8_9_331_0, i_8_9_346_0, i_8_9_378_0,
    i_8_9_401_0, i_8_9_422_0, i_8_9_445_0, i_8_9_478_0, i_8_9_479_0,
    i_8_9_480_0, i_8_9_482_0, i_8_9_484_0, i_8_9_490_0, i_8_9_501_0,
    i_8_9_528_0, i_8_9_530_0, i_8_9_548_0, i_8_9_579_0, i_8_9_609_0,
    i_8_9_678_0, i_8_9_705_0, i_8_9_714_0, i_8_9_715_0, i_8_9_781_0,
    i_8_9_850_0, i_8_9_922_0, i_8_9_937_0, i_8_9_952_0, i_8_9_955_0,
    i_8_9_994_0, i_8_9_995_0, i_8_9_1030_0, i_8_9_1031_0, i_8_9_1075_0,
    i_8_9_1079_0, i_8_9_1112_0, i_8_9_1127_0, i_8_9_1243_0, i_8_9_1265_0,
    i_8_9_1270_0, i_8_9_1271_0, i_8_9_1274_0, i_8_9_1283_0, i_8_9_1306_0,
    i_8_9_1307_0, i_8_9_1390_0, i_8_9_1479_0, i_8_9_1492_0, i_8_9_1503_0,
    i_8_9_1521_0, i_8_9_1543_0, i_8_9_1544_0, i_8_9_1550_0, i_8_9_1574_0,
    i_8_9_1579_0, i_8_9_1653_0, i_8_9_1669_0, i_8_9_1684_0, i_8_9_1707_0,
    i_8_9_1716_0, i_8_9_1746_0, i_8_9_1750_0, i_8_9_1774_0, i_8_9_1779_0,
    i_8_9_1780_0, i_8_9_1804_0, i_8_9_1821_0, i_8_9_1894_0, i_8_9_1917_0,
    i_8_9_1920_0, i_8_9_2129_0, i_8_9_2130_0, i_8_9_2131_0, i_8_9_2143_0,
    i_8_9_2148_0, i_8_9_2214_0, i_8_9_2215_0, i_8_9_2218_0, i_8_9_2229_0,
    i_8_9_2235_0, i_8_9_2242_0, i_8_9_2281_0, i_8_9_2282_0,
    o_8_9_0_0  );
  input  i_8_9_46_0, i_8_9_58_0, i_8_9_59_0, i_8_9_85_0, i_8_9_87_0,
    i_8_9_88_0, i_8_9_106_0, i_8_9_140_0, i_8_9_142_0, i_8_9_143_0,
    i_8_9_187_0, i_8_9_188_0, i_8_9_252_0, i_8_9_256_0, i_8_9_259_0,
    i_8_9_303_0, i_8_9_304_0, i_8_9_311_0, i_8_9_331_0, i_8_9_346_0,
    i_8_9_378_0, i_8_9_401_0, i_8_9_422_0, i_8_9_445_0, i_8_9_478_0,
    i_8_9_479_0, i_8_9_480_0, i_8_9_482_0, i_8_9_484_0, i_8_9_490_0,
    i_8_9_501_0, i_8_9_528_0, i_8_9_530_0, i_8_9_548_0, i_8_9_579_0,
    i_8_9_609_0, i_8_9_678_0, i_8_9_705_0, i_8_9_714_0, i_8_9_715_0,
    i_8_9_781_0, i_8_9_850_0, i_8_9_922_0, i_8_9_937_0, i_8_9_952_0,
    i_8_9_955_0, i_8_9_994_0, i_8_9_995_0, i_8_9_1030_0, i_8_9_1031_0,
    i_8_9_1075_0, i_8_9_1079_0, i_8_9_1112_0, i_8_9_1127_0, i_8_9_1243_0,
    i_8_9_1265_0, i_8_9_1270_0, i_8_9_1271_0, i_8_9_1274_0, i_8_9_1283_0,
    i_8_9_1306_0, i_8_9_1307_0, i_8_9_1390_0, i_8_9_1479_0, i_8_9_1492_0,
    i_8_9_1503_0, i_8_9_1521_0, i_8_9_1543_0, i_8_9_1544_0, i_8_9_1550_0,
    i_8_9_1574_0, i_8_9_1579_0, i_8_9_1653_0, i_8_9_1669_0, i_8_9_1684_0,
    i_8_9_1707_0, i_8_9_1716_0, i_8_9_1746_0, i_8_9_1750_0, i_8_9_1774_0,
    i_8_9_1779_0, i_8_9_1780_0, i_8_9_1804_0, i_8_9_1821_0, i_8_9_1894_0,
    i_8_9_1917_0, i_8_9_1920_0, i_8_9_2129_0, i_8_9_2130_0, i_8_9_2131_0,
    i_8_9_2143_0, i_8_9_2148_0, i_8_9_2214_0, i_8_9_2215_0, i_8_9_2218_0,
    i_8_9_2229_0, i_8_9_2235_0, i_8_9_2242_0, i_8_9_2281_0, i_8_9_2282_0;
  output o_8_9_0_0;
  assign o_8_9_0_0 = 0;
endmodule



// Benchmark "kernel_8_10" written by ABC on Sun Jul 19 10:03:13 2020

module kernel_8_10 ( 
    i_8_10_3_0, i_8_10_22_0, i_8_10_40_0, i_8_10_94_0, i_8_10_193_0,
    i_8_10_201_0, i_8_10_246_0, i_8_10_256_0, i_8_10_277_0, i_8_10_283_0,
    i_8_10_352_0, i_8_10_355_0, i_8_10_356_0, i_8_10_358_0, i_8_10_367_0,
    i_8_10_426_0, i_8_10_457_0, i_8_10_516_0, i_8_10_517_0, i_8_10_527_0,
    i_8_10_528_0, i_8_10_556_0, i_8_10_594_0, i_8_10_612_0, i_8_10_613_0,
    i_8_10_616_0, i_8_10_622_0, i_8_10_632_0, i_8_10_633_0, i_8_10_666_0,
    i_8_10_698_0, i_8_10_704_0, i_8_10_705_0, i_8_10_782_0, i_8_10_814_0,
    i_8_10_832_0, i_8_10_838_0, i_8_10_877_0, i_8_10_912_0, i_8_10_958_0,
    i_8_10_995_0, i_8_10_1128_0, i_8_10_1174_0, i_8_10_1192_0,
    i_8_10_1201_0, i_8_10_1228_0, i_8_10_1263_0, i_8_10_1284_0,
    i_8_10_1299_0, i_8_10_1305_0, i_8_10_1306_0, i_8_10_1307_0,
    i_8_10_1315_0, i_8_10_1354_0, i_8_10_1390_0, i_8_10_1467_0,
    i_8_10_1473_0, i_8_10_1497_0, i_8_10_1524_0, i_8_10_1525_0,
    i_8_10_1534_0, i_8_10_1570_0, i_8_10_1624_0, i_8_10_1635_0,
    i_8_10_1648_0, i_8_10_1678_0, i_8_10_1686_0, i_8_10_1696_0,
    i_8_10_1714_0, i_8_10_1746_0, i_8_10_1747_0, i_8_10_1752_0,
    i_8_10_1776_0, i_8_10_1791_0, i_8_10_1795_0, i_8_10_1801_0,
    i_8_10_1806_0, i_8_10_1818_0, i_8_10_1822_0, i_8_10_1848_0,
    i_8_10_1849_0, i_8_10_1876_0, i_8_10_1906_0, i_8_10_1918_0,
    i_8_10_1976_0, i_8_10_2014_0, i_8_10_2046_0, i_8_10_2047_0,
    i_8_10_2064_0, i_8_10_2065_0, i_8_10_2066_0, i_8_10_2091_0,
    i_8_10_2092_0, i_8_10_2119_0, i_8_10_2122_0, i_8_10_2155_0,
    i_8_10_2215_0, i_8_10_2216_0, i_8_10_2256_0, i_8_10_2291_0,
    o_8_10_0_0  );
  input  i_8_10_3_0, i_8_10_22_0, i_8_10_40_0, i_8_10_94_0, i_8_10_193_0,
    i_8_10_201_0, i_8_10_246_0, i_8_10_256_0, i_8_10_277_0, i_8_10_283_0,
    i_8_10_352_0, i_8_10_355_0, i_8_10_356_0, i_8_10_358_0, i_8_10_367_0,
    i_8_10_426_0, i_8_10_457_0, i_8_10_516_0, i_8_10_517_0, i_8_10_527_0,
    i_8_10_528_0, i_8_10_556_0, i_8_10_594_0, i_8_10_612_0, i_8_10_613_0,
    i_8_10_616_0, i_8_10_622_0, i_8_10_632_0, i_8_10_633_0, i_8_10_666_0,
    i_8_10_698_0, i_8_10_704_0, i_8_10_705_0, i_8_10_782_0, i_8_10_814_0,
    i_8_10_832_0, i_8_10_838_0, i_8_10_877_0, i_8_10_912_0, i_8_10_958_0,
    i_8_10_995_0, i_8_10_1128_0, i_8_10_1174_0, i_8_10_1192_0,
    i_8_10_1201_0, i_8_10_1228_0, i_8_10_1263_0, i_8_10_1284_0,
    i_8_10_1299_0, i_8_10_1305_0, i_8_10_1306_0, i_8_10_1307_0,
    i_8_10_1315_0, i_8_10_1354_0, i_8_10_1390_0, i_8_10_1467_0,
    i_8_10_1473_0, i_8_10_1497_0, i_8_10_1524_0, i_8_10_1525_0,
    i_8_10_1534_0, i_8_10_1570_0, i_8_10_1624_0, i_8_10_1635_0,
    i_8_10_1648_0, i_8_10_1678_0, i_8_10_1686_0, i_8_10_1696_0,
    i_8_10_1714_0, i_8_10_1746_0, i_8_10_1747_0, i_8_10_1752_0,
    i_8_10_1776_0, i_8_10_1791_0, i_8_10_1795_0, i_8_10_1801_0,
    i_8_10_1806_0, i_8_10_1818_0, i_8_10_1822_0, i_8_10_1848_0,
    i_8_10_1849_0, i_8_10_1876_0, i_8_10_1906_0, i_8_10_1918_0,
    i_8_10_1976_0, i_8_10_2014_0, i_8_10_2046_0, i_8_10_2047_0,
    i_8_10_2064_0, i_8_10_2065_0, i_8_10_2066_0, i_8_10_2091_0,
    i_8_10_2092_0, i_8_10_2119_0, i_8_10_2122_0, i_8_10_2155_0,
    i_8_10_2215_0, i_8_10_2216_0, i_8_10_2256_0, i_8_10_2291_0;
  output o_8_10_0_0;
  assign o_8_10_0_0 = ~((~i_8_10_356_0 & ((~i_8_10_201_0 & ((~i_8_10_3_0 & ~i_8_10_246_0 & ~i_8_10_352_0 & ~i_8_10_832_0 & ~i_8_10_1849_0 & ~i_8_10_2066_0 & ~i_8_10_2256_0) | (~i_8_10_516_0 & ~i_8_10_616_0 & ~i_8_10_1128_0 & ~i_8_10_1534_0 & i_8_10_1648_0 & ~i_8_10_1776_0 & ~i_8_10_2119_0 & ~i_8_10_2291_0))) | (~i_8_10_1305_0 & ((~i_8_10_283_0 & ~i_8_10_832_0 & ~i_8_10_958_0 & ~i_8_10_1201_0 & ~i_8_10_1686_0 & ~i_8_10_1848_0 & ~i_8_10_1876_0 & ~i_8_10_2064_0) | (~i_8_10_516_0 & ~i_8_10_632_0 & ~i_8_10_633_0 & ~i_8_10_1228_0 & ~i_8_10_1849_0 & i_8_10_2092_0))) | (~i_8_10_2091_0 & ((i_8_10_1284_0 & ~i_8_10_1635_0 & ~i_8_10_1795_0 & ~i_8_10_2014_0) | (~i_8_10_1263_0 & ~i_8_10_1534_0 & ~i_8_10_1791_0 & ~i_8_10_1876_0 & ~i_8_10_2065_0))))) | (~i_8_10_527_0 & ((~i_8_10_40_0 & i_8_10_1648_0 & ((~i_8_10_355_0 & ~i_8_10_516_0 & ~i_8_10_594_0 & ~i_8_10_1174_0 & ~i_8_10_1201_0 & ~i_8_10_1525_0 & i_8_10_1818_0) | (~i_8_10_457_0 & ~i_8_10_1696_0 & i_8_10_1822_0 & ~i_8_10_1848_0 & ~i_8_10_1849_0 & ~i_8_10_2119_0))) | (~i_8_10_528_0 & ~i_8_10_1307_0 & ((~i_8_10_246_0 & ~i_8_10_352_0 & ~i_8_10_367_0 & ~i_8_10_516_0 & ~i_8_10_632_0 & ~i_8_10_704_0 & ~i_8_10_1467_0 & ~i_8_10_1648_0) | (~i_8_10_517_0 & ~i_8_10_832_0 & ~i_8_10_2065_0 & ~i_8_10_2215_0))))) | (~i_8_10_1497_0 & ((~i_8_10_352_0 & ((~i_8_10_22_0 & i_8_10_528_0 & ~i_8_10_1876_0) | (~i_8_10_358_0 & ~i_8_10_516_0 & ~i_8_10_517_0 & i_8_10_527_0 & ~i_8_10_612_0 & ~i_8_10_613_0 & ~i_8_10_2122_0 & ~i_8_10_2215_0))) | (~i_8_10_613_0 & i_8_10_838_0 & ~i_8_10_1201_0 & ~i_8_10_1534_0) | (i_8_10_256_0 & ~i_8_10_517_0 & ~i_8_10_704_0 & ~i_8_10_1776_0) | (~i_8_10_516_0 & i_8_10_1534_0 & i_8_10_1678_0 & ~i_8_10_1714_0 & ~i_8_10_1795_0 & ~i_8_10_1806_0 & ~i_8_10_2064_0 & ~i_8_10_2065_0) | (~i_8_10_40_0 & ~i_8_10_612_0 & i_8_10_877_0 & ~i_8_10_1299_0 & ~i_8_10_1746_0 & ~i_8_10_2092_0))) | (~i_8_10_516_0 & ((i_8_10_1524_0 & ~i_8_10_1648_0) | (~i_8_10_355_0 & ~i_8_10_1467_0 & i_8_10_1624_0 & ~i_8_10_2047_0))) | (~i_8_10_355_0 & ((~i_8_10_612_0 & ~i_8_10_632_0 & ~i_8_10_1174_0 & ~i_8_10_1776_0 & ~i_8_10_2065_0 & ~i_8_10_2215_0) | (~i_8_10_256_0 & ~i_8_10_698_0 & i_8_10_1746_0 & ~i_8_10_1806_0 & ~i_8_10_1849_0 & ~i_8_10_2092_0 & ~i_8_10_2291_0))) | (~i_8_10_517_0 & ((~i_8_10_426_0 & i_8_10_613_0 & i_8_10_622_0 & ~i_8_10_705_0 & ~i_8_10_1648_0) | (i_8_10_612_0 & ~i_8_10_838_0 & ~i_8_10_1174_0 & i_8_10_1801_0 & ~i_8_10_2066_0))) | (~i_8_10_2047_0 & ((i_8_10_94_0 & i_8_10_556_0) | (~i_8_10_1849_0 & ~i_8_10_2064_0 & ~i_8_10_2065_0 & ~i_8_10_2066_0))) | (~i_8_10_632_0 & ~i_8_10_633_0 & ~i_8_10_1263_0 & ~i_8_10_1299_0 & ~i_8_10_1307_0 & i_8_10_1678_0 & i_8_10_2091_0 & ~i_8_10_2122_0));
endmodule



// Benchmark "kernel_8_11" written by ABC on Sun Jul 19 10:03:13 2020

module kernel_8_11 ( 
    i_8_11_64_0, i_8_11_79_0, i_8_11_111_0, i_8_11_141_0, i_8_11_197_0,
    i_8_11_231_0, i_8_11_262_0, i_8_11_265_0, i_8_11_311_0, i_8_11_326_0,
    i_8_11_329_0, i_8_11_364_0, i_8_11_367_0, i_8_11_379_0, i_8_11_392_0,
    i_8_11_401_0, i_8_11_419_0, i_8_11_424_0, i_8_11_439_0, i_8_11_475_0,
    i_8_11_486_0, i_8_11_499_0, i_8_11_509_0, i_8_11_525_0, i_8_11_528_0,
    i_8_11_529_0, i_8_11_557_0, i_8_11_571_0, i_8_11_616_0, i_8_11_625_0,
    i_8_11_631_0, i_8_11_635_0, i_8_11_656_0, i_8_11_659_0, i_8_11_661_0,
    i_8_11_673_0, i_8_11_700_0, i_8_11_703_0, i_8_11_718_0, i_8_11_724_0,
    i_8_11_725_0, i_8_11_734_0, i_8_11_754_0, i_8_11_771_0, i_8_11_824_0,
    i_8_11_835_0, i_8_11_837_0, i_8_11_838_0, i_8_11_840_0, i_8_11_841_0,
    i_8_11_968_0, i_8_11_1012_0, i_8_11_1110_0, i_8_11_1191_0,
    i_8_11_1229_0, i_8_11_1231_0, i_8_11_1246_0, i_8_11_1267_0,
    i_8_11_1301_0, i_8_11_1354_0, i_8_11_1355_0, i_8_11_1399_0,
    i_8_11_1411_0, i_8_11_1462_0, i_8_11_1471_0, i_8_11_1547_0,
    i_8_11_1571_0, i_8_11_1625_0, i_8_11_1647_0, i_8_11_1653_0,
    i_8_11_1655_0, i_8_11_1679_0, i_8_11_1696_0, i_8_11_1699_0,
    i_8_11_1747_0, i_8_11_1748_0, i_8_11_1750_0, i_8_11_1754_0,
    i_8_11_1769_0, i_8_11_1773_0, i_8_11_1795_0, i_8_11_1798_0,
    i_8_11_1819_0, i_8_11_1840_0, i_8_11_1849_0, i_8_11_1858_0,
    i_8_11_1912_0, i_8_11_1913_0, i_8_11_1952_0, i_8_11_1981_0,
    i_8_11_2011_0, i_8_11_2012_0, i_8_11_2048_0, i_8_11_2074_0,
    i_8_11_2095_0, i_8_11_2119_0, i_8_11_2136_0, i_8_11_2191_0,
    i_8_11_2257_0, i_8_11_2298_0,
    o_8_11_0_0  );
  input  i_8_11_64_0, i_8_11_79_0, i_8_11_111_0, i_8_11_141_0,
    i_8_11_197_0, i_8_11_231_0, i_8_11_262_0, i_8_11_265_0, i_8_11_311_0,
    i_8_11_326_0, i_8_11_329_0, i_8_11_364_0, i_8_11_367_0, i_8_11_379_0,
    i_8_11_392_0, i_8_11_401_0, i_8_11_419_0, i_8_11_424_0, i_8_11_439_0,
    i_8_11_475_0, i_8_11_486_0, i_8_11_499_0, i_8_11_509_0, i_8_11_525_0,
    i_8_11_528_0, i_8_11_529_0, i_8_11_557_0, i_8_11_571_0, i_8_11_616_0,
    i_8_11_625_0, i_8_11_631_0, i_8_11_635_0, i_8_11_656_0, i_8_11_659_0,
    i_8_11_661_0, i_8_11_673_0, i_8_11_700_0, i_8_11_703_0, i_8_11_718_0,
    i_8_11_724_0, i_8_11_725_0, i_8_11_734_0, i_8_11_754_0, i_8_11_771_0,
    i_8_11_824_0, i_8_11_835_0, i_8_11_837_0, i_8_11_838_0, i_8_11_840_0,
    i_8_11_841_0, i_8_11_968_0, i_8_11_1012_0, i_8_11_1110_0,
    i_8_11_1191_0, i_8_11_1229_0, i_8_11_1231_0, i_8_11_1246_0,
    i_8_11_1267_0, i_8_11_1301_0, i_8_11_1354_0, i_8_11_1355_0,
    i_8_11_1399_0, i_8_11_1411_0, i_8_11_1462_0, i_8_11_1471_0,
    i_8_11_1547_0, i_8_11_1571_0, i_8_11_1625_0, i_8_11_1647_0,
    i_8_11_1653_0, i_8_11_1655_0, i_8_11_1679_0, i_8_11_1696_0,
    i_8_11_1699_0, i_8_11_1747_0, i_8_11_1748_0, i_8_11_1750_0,
    i_8_11_1754_0, i_8_11_1769_0, i_8_11_1773_0, i_8_11_1795_0,
    i_8_11_1798_0, i_8_11_1819_0, i_8_11_1840_0, i_8_11_1849_0,
    i_8_11_1858_0, i_8_11_1912_0, i_8_11_1913_0, i_8_11_1952_0,
    i_8_11_1981_0, i_8_11_2011_0, i_8_11_2012_0, i_8_11_2048_0,
    i_8_11_2074_0, i_8_11_2095_0, i_8_11_2119_0, i_8_11_2136_0,
    i_8_11_2191_0, i_8_11_2257_0, i_8_11_2298_0;
  output o_8_11_0_0;
  assign o_8_11_0_0 = 0;
endmodule



// Benchmark "kernel_8_12" written by ABC on Sun Jul 19 10:03:14 2020

module kernel_8_12 ( 
    i_8_12_13_0, i_8_12_92_0, i_8_12_94_0, i_8_12_121_0, i_8_12_138_0,
    i_8_12_139_0, i_8_12_183_0, i_8_12_192_0, i_8_12_193_0, i_8_12_209_0,
    i_8_12_221_0, i_8_12_278_0, i_8_12_284_0, i_8_12_318_0, i_8_12_325_0,
    i_8_12_326_0, i_8_12_350_0, i_8_12_363_0, i_8_12_390_0, i_8_12_471_0,
    i_8_12_472_0, i_8_12_473_0, i_8_12_478_0, i_8_12_480_0, i_8_12_481_0,
    i_8_12_505_0, i_8_12_523_0, i_8_12_554_0, i_8_12_569_0, i_8_12_632_0,
    i_8_12_656_0, i_8_12_694_0, i_8_12_696_0, i_8_12_697_0, i_8_12_712_0,
    i_8_12_731_0, i_8_12_749_0, i_8_12_750_0, i_8_12_863_0, i_8_12_877_0,
    i_8_12_883_0, i_8_12_893_0, i_8_12_959_0, i_8_12_962_0, i_8_12_964_0,
    i_8_12_967_0, i_8_12_991_0, i_8_12_995_0, i_8_12_1027_0, i_8_12_1094_0,
    i_8_12_1120_0, i_8_12_1144_0, i_8_12_1201_0, i_8_12_1202_0,
    i_8_12_1234_0, i_8_12_1286_0, i_8_12_1309_0, i_8_12_1315_0,
    i_8_12_1316_0, i_8_12_1328_0, i_8_12_1342_0, i_8_12_1372_0,
    i_8_12_1382_0, i_8_12_1413_0, i_8_12_1432_0, i_8_12_1434_0,
    i_8_12_1442_0, i_8_12_1621_0, i_8_12_1625_0, i_8_12_1651_0,
    i_8_12_1665_0, i_8_12_1666_0, i_8_12_1696_0, i_8_12_1699_0,
    i_8_12_1705_0, i_8_12_1712_0, i_8_12_1749_0, i_8_12_1751_0,
    i_8_12_1805_0, i_8_12_1818_0, i_8_12_1857_0, i_8_12_1874_0,
    i_8_12_1981_0, i_8_12_1982_0, i_8_12_2008_0, i_8_12_2009_0,
    i_8_12_2025_0, i_8_12_2053_0, i_8_12_2083_0, i_8_12_2084_0,
    i_8_12_2090_0, i_8_12_2122_0, i_8_12_2123_0, i_8_12_2143_0,
    i_8_12_2170_0, i_8_12_2189_0, i_8_12_2227_0, i_8_12_2284_0,
    i_8_12_2285_0, i_8_12_2299_0,
    o_8_12_0_0  );
  input  i_8_12_13_0, i_8_12_92_0, i_8_12_94_0, i_8_12_121_0,
    i_8_12_138_0, i_8_12_139_0, i_8_12_183_0, i_8_12_192_0, i_8_12_193_0,
    i_8_12_209_0, i_8_12_221_0, i_8_12_278_0, i_8_12_284_0, i_8_12_318_0,
    i_8_12_325_0, i_8_12_326_0, i_8_12_350_0, i_8_12_363_0, i_8_12_390_0,
    i_8_12_471_0, i_8_12_472_0, i_8_12_473_0, i_8_12_478_0, i_8_12_480_0,
    i_8_12_481_0, i_8_12_505_0, i_8_12_523_0, i_8_12_554_0, i_8_12_569_0,
    i_8_12_632_0, i_8_12_656_0, i_8_12_694_0, i_8_12_696_0, i_8_12_697_0,
    i_8_12_712_0, i_8_12_731_0, i_8_12_749_0, i_8_12_750_0, i_8_12_863_0,
    i_8_12_877_0, i_8_12_883_0, i_8_12_893_0, i_8_12_959_0, i_8_12_962_0,
    i_8_12_964_0, i_8_12_967_0, i_8_12_991_0, i_8_12_995_0, i_8_12_1027_0,
    i_8_12_1094_0, i_8_12_1120_0, i_8_12_1144_0, i_8_12_1201_0,
    i_8_12_1202_0, i_8_12_1234_0, i_8_12_1286_0, i_8_12_1309_0,
    i_8_12_1315_0, i_8_12_1316_0, i_8_12_1328_0, i_8_12_1342_0,
    i_8_12_1372_0, i_8_12_1382_0, i_8_12_1413_0, i_8_12_1432_0,
    i_8_12_1434_0, i_8_12_1442_0, i_8_12_1621_0, i_8_12_1625_0,
    i_8_12_1651_0, i_8_12_1665_0, i_8_12_1666_0, i_8_12_1696_0,
    i_8_12_1699_0, i_8_12_1705_0, i_8_12_1712_0, i_8_12_1749_0,
    i_8_12_1751_0, i_8_12_1805_0, i_8_12_1818_0, i_8_12_1857_0,
    i_8_12_1874_0, i_8_12_1981_0, i_8_12_1982_0, i_8_12_2008_0,
    i_8_12_2009_0, i_8_12_2025_0, i_8_12_2053_0, i_8_12_2083_0,
    i_8_12_2084_0, i_8_12_2090_0, i_8_12_2122_0, i_8_12_2123_0,
    i_8_12_2143_0, i_8_12_2170_0, i_8_12_2189_0, i_8_12_2227_0,
    i_8_12_2284_0, i_8_12_2285_0, i_8_12_2299_0;
  output o_8_12_0_0;
  assign o_8_12_0_0 = 0;
endmodule



// Benchmark "kernel_8_13" written by ABC on Sun Jul 19 10:03:15 2020

module kernel_8_13 ( 
    i_8_13_4_0, i_8_13_28_0, i_8_13_33_0, i_8_13_47_0, i_8_13_58_0,
    i_8_13_59_0, i_8_13_71_0, i_8_13_166_0, i_8_13_170_0, i_8_13_190_0,
    i_8_13_227_0, i_8_13_256_0, i_8_13_257_0, i_8_13_281_0, i_8_13_293_0,
    i_8_13_320_0, i_8_13_326_0, i_8_13_328_0, i_8_13_364_0, i_8_13_379_0,
    i_8_13_380_0, i_8_13_421_0, i_8_13_424_0, i_8_13_444_0, i_8_13_453_0,
    i_8_13_593_0, i_8_13_603_0, i_8_13_660_0, i_8_13_693_0, i_8_13_703_0,
    i_8_13_704_0, i_8_13_705_0, i_8_13_706_0, i_8_13_708_0, i_8_13_778_0,
    i_8_13_784_0, i_8_13_787_0, i_8_13_826_0, i_8_13_832_0, i_8_13_833_0,
    i_8_13_838_0, i_8_13_842_0, i_8_13_844_0, i_8_13_873_0, i_8_13_877_0,
    i_8_13_886_0, i_8_13_890_0, i_8_13_928_0, i_8_13_932_0, i_8_13_977_0,
    i_8_13_1083_0, i_8_13_1108_0, i_8_13_1115_0, i_8_13_1174_0,
    i_8_13_1180_0, i_8_13_1183_0, i_8_13_1234_0, i_8_13_1236_0,
    i_8_13_1271_0, i_8_13_1282_0, i_8_13_1286_0, i_8_13_1327_0,
    i_8_13_1352_0, i_8_13_1360_0, i_8_13_1435_0, i_8_13_1442_0,
    i_8_13_1472_0, i_8_13_1474_0, i_8_13_1498_0, i_8_13_1533_0,
    i_8_13_1597_0, i_8_13_1603_0, i_8_13_1607_0, i_8_13_1634_0,
    i_8_13_1673_0, i_8_13_1706_0, i_8_13_1746_0, i_8_13_1748_0,
    i_8_13_1764_0, i_8_13_1769_0, i_8_13_1789_0, i_8_13_1807_0,
    i_8_13_1813_0, i_8_13_1824_0, i_8_13_1881_0, i_8_13_1907_0,
    i_8_13_1965_0, i_8_13_1967_0, i_8_13_1984_0, i_8_13_1987_0,
    i_8_13_1989_0, i_8_13_2038_0, i_8_13_2052_0, i_8_13_2056_0,
    i_8_13_2060_0, i_8_13_2143_0, i_8_13_2150_0, i_8_13_2224_0,
    i_8_13_2263_0, i_8_13_2264_0,
    o_8_13_0_0  );
  input  i_8_13_4_0, i_8_13_28_0, i_8_13_33_0, i_8_13_47_0, i_8_13_58_0,
    i_8_13_59_0, i_8_13_71_0, i_8_13_166_0, i_8_13_170_0, i_8_13_190_0,
    i_8_13_227_0, i_8_13_256_0, i_8_13_257_0, i_8_13_281_0, i_8_13_293_0,
    i_8_13_320_0, i_8_13_326_0, i_8_13_328_0, i_8_13_364_0, i_8_13_379_0,
    i_8_13_380_0, i_8_13_421_0, i_8_13_424_0, i_8_13_444_0, i_8_13_453_0,
    i_8_13_593_0, i_8_13_603_0, i_8_13_660_0, i_8_13_693_0, i_8_13_703_0,
    i_8_13_704_0, i_8_13_705_0, i_8_13_706_0, i_8_13_708_0, i_8_13_778_0,
    i_8_13_784_0, i_8_13_787_0, i_8_13_826_0, i_8_13_832_0, i_8_13_833_0,
    i_8_13_838_0, i_8_13_842_0, i_8_13_844_0, i_8_13_873_0, i_8_13_877_0,
    i_8_13_886_0, i_8_13_890_0, i_8_13_928_0, i_8_13_932_0, i_8_13_977_0,
    i_8_13_1083_0, i_8_13_1108_0, i_8_13_1115_0, i_8_13_1174_0,
    i_8_13_1180_0, i_8_13_1183_0, i_8_13_1234_0, i_8_13_1236_0,
    i_8_13_1271_0, i_8_13_1282_0, i_8_13_1286_0, i_8_13_1327_0,
    i_8_13_1352_0, i_8_13_1360_0, i_8_13_1435_0, i_8_13_1442_0,
    i_8_13_1472_0, i_8_13_1474_0, i_8_13_1498_0, i_8_13_1533_0,
    i_8_13_1597_0, i_8_13_1603_0, i_8_13_1607_0, i_8_13_1634_0,
    i_8_13_1673_0, i_8_13_1706_0, i_8_13_1746_0, i_8_13_1748_0,
    i_8_13_1764_0, i_8_13_1769_0, i_8_13_1789_0, i_8_13_1807_0,
    i_8_13_1813_0, i_8_13_1824_0, i_8_13_1881_0, i_8_13_1907_0,
    i_8_13_1965_0, i_8_13_1967_0, i_8_13_1984_0, i_8_13_1987_0,
    i_8_13_1989_0, i_8_13_2038_0, i_8_13_2052_0, i_8_13_2056_0,
    i_8_13_2060_0, i_8_13_2143_0, i_8_13_2150_0, i_8_13_2224_0,
    i_8_13_2263_0, i_8_13_2264_0;
  output o_8_13_0_0;
  assign o_8_13_0_0 = 0;
endmodule



// Benchmark "kernel_8_14" written by ABC on Sun Jul 19 10:03:16 2020

module kernel_8_14 ( 
    i_8_14_25_0, i_8_14_41_0, i_8_14_170_0, i_8_14_174_0, i_8_14_178_0,
    i_8_14_228_0, i_8_14_230_0, i_8_14_231_0, i_8_14_233_0, i_8_14_248_0,
    i_8_14_273_0, i_8_14_277_0, i_8_14_278_0, i_8_14_355_0, i_8_14_356_0,
    i_8_14_359_0, i_8_14_363_0, i_8_14_364_0, i_8_14_385_0, i_8_14_391_0,
    i_8_14_476_0, i_8_14_484_0, i_8_14_499_0, i_8_14_516_0, i_8_14_518_0,
    i_8_14_592_0, i_8_14_597_0, i_8_14_607_0, i_8_14_608_0, i_8_14_611_0,
    i_8_14_626_0, i_8_14_634_0, i_8_14_772_0, i_8_14_799_0, i_8_14_825_0,
    i_8_14_830_0, i_8_14_841_0, i_8_14_879_0, i_8_14_889_0, i_8_14_925_0,
    i_8_14_935_0, i_8_14_955_0, i_8_14_958_0, i_8_14_959_0, i_8_14_994_0,
    i_8_14_996_0, i_8_14_1039_0, i_8_14_1075_0, i_8_14_1076_0,
    i_8_14_1087_0, i_8_14_1178_0, i_8_14_1192_0, i_8_14_1228_0,
    i_8_14_1232_0, i_8_14_1241_0, i_8_14_1258_0, i_8_14_1273_0,
    i_8_14_1274_0, i_8_14_1277_0, i_8_14_1285_0, i_8_14_1385_0,
    i_8_14_1387_0, i_8_14_1391_0, i_8_14_1408_0, i_8_14_1412_0,
    i_8_14_1497_0, i_8_14_1525_0, i_8_14_1528_0, i_8_14_1546_0,
    i_8_14_1552_0, i_8_14_1645_0, i_8_14_1647_0, i_8_14_1650_0,
    i_8_14_1659_0, i_8_14_1680_0, i_8_14_1681_0, i_8_14_1726_0,
    i_8_14_1767_0, i_8_14_1768_0, i_8_14_1771_0, i_8_14_1800_0,
    i_8_14_1807_0, i_8_14_1849_0, i_8_14_1866_0, i_8_14_1870_0,
    i_8_14_1906_0, i_8_14_1919_0, i_8_14_1940_0, i_8_14_1967_0,
    i_8_14_1996_0, i_8_14_2040_0, i_8_14_2041_0, i_8_14_2066_0,
    i_8_14_2075_0, i_8_14_2146_0, i_8_14_2150_0, i_8_14_2159_0,
    i_8_14_2212_0, i_8_14_2219_0, i_8_14_2249_0,
    o_8_14_0_0  );
  input  i_8_14_25_0, i_8_14_41_0, i_8_14_170_0, i_8_14_174_0,
    i_8_14_178_0, i_8_14_228_0, i_8_14_230_0, i_8_14_231_0, i_8_14_233_0,
    i_8_14_248_0, i_8_14_273_0, i_8_14_277_0, i_8_14_278_0, i_8_14_355_0,
    i_8_14_356_0, i_8_14_359_0, i_8_14_363_0, i_8_14_364_0, i_8_14_385_0,
    i_8_14_391_0, i_8_14_476_0, i_8_14_484_0, i_8_14_499_0, i_8_14_516_0,
    i_8_14_518_0, i_8_14_592_0, i_8_14_597_0, i_8_14_607_0, i_8_14_608_0,
    i_8_14_611_0, i_8_14_626_0, i_8_14_634_0, i_8_14_772_0, i_8_14_799_0,
    i_8_14_825_0, i_8_14_830_0, i_8_14_841_0, i_8_14_879_0, i_8_14_889_0,
    i_8_14_925_0, i_8_14_935_0, i_8_14_955_0, i_8_14_958_0, i_8_14_959_0,
    i_8_14_994_0, i_8_14_996_0, i_8_14_1039_0, i_8_14_1075_0,
    i_8_14_1076_0, i_8_14_1087_0, i_8_14_1178_0, i_8_14_1192_0,
    i_8_14_1228_0, i_8_14_1232_0, i_8_14_1241_0, i_8_14_1258_0,
    i_8_14_1273_0, i_8_14_1274_0, i_8_14_1277_0, i_8_14_1285_0,
    i_8_14_1385_0, i_8_14_1387_0, i_8_14_1391_0, i_8_14_1408_0,
    i_8_14_1412_0, i_8_14_1497_0, i_8_14_1525_0, i_8_14_1528_0,
    i_8_14_1546_0, i_8_14_1552_0, i_8_14_1645_0, i_8_14_1647_0,
    i_8_14_1650_0, i_8_14_1659_0, i_8_14_1680_0, i_8_14_1681_0,
    i_8_14_1726_0, i_8_14_1767_0, i_8_14_1768_0, i_8_14_1771_0,
    i_8_14_1800_0, i_8_14_1807_0, i_8_14_1849_0, i_8_14_1866_0,
    i_8_14_1870_0, i_8_14_1906_0, i_8_14_1919_0, i_8_14_1940_0,
    i_8_14_1967_0, i_8_14_1996_0, i_8_14_2040_0, i_8_14_2041_0,
    i_8_14_2066_0, i_8_14_2075_0, i_8_14_2146_0, i_8_14_2150_0,
    i_8_14_2159_0, i_8_14_2212_0, i_8_14_2219_0, i_8_14_2249_0;
  output o_8_14_0_0;
  assign o_8_14_0_0 = ~((~i_8_14_230_0 & ((~i_8_14_273_0 & ~i_8_14_385_0 & ~i_8_14_597_0 & ~i_8_14_955_0 & ~i_8_14_1241_0 & ~i_8_14_1385_0 & ~i_8_14_1387_0 & ~i_8_14_1408_0 & i_8_14_1552_0) | (~i_8_14_25_0 & ~i_8_14_41_0 & ~i_8_14_174_0 & ~i_8_14_476_0 & ~i_8_14_799_0 & ~i_8_14_830_0 & ~i_8_14_1232_0 & ~i_8_14_1258_0 & ~i_8_14_1273_0 & ~i_8_14_1647_0 & ~i_8_14_2159_0))) | (~i_8_14_25_0 & ((~i_8_14_592_0 & i_8_14_626_0 & ~i_8_14_955_0 & ~i_8_14_1277_0 & ~i_8_14_1546_0 & i_8_14_1552_0) | (~i_8_14_41_0 & ~i_8_14_174_0 & ~i_8_14_356_0 & ~i_8_14_359_0 & ~i_8_14_364_0 & ~i_8_14_597_0 & ~i_8_14_772_0 & ~i_8_14_1385_0 & ~i_8_14_1552_0 & ~i_8_14_1906_0 & ~i_8_14_2146_0))) | (~i_8_14_178_0 & ((~i_8_14_174_0 & ~i_8_14_355_0 & ((~i_8_14_959_0 & ~i_8_14_1076_0 & ~i_8_14_1178_0 & ~i_8_14_1258_0 & ~i_8_14_1277_0 & ~i_8_14_1391_0 & ~i_8_14_1849_0 & ~i_8_14_1940_0) | (~i_8_14_170_0 & ~i_8_14_248_0 & ~i_8_14_359_0 & ~i_8_14_499_0 & ~i_8_14_830_0 & ~i_8_14_1232_0 & ~i_8_14_1546_0 & ~i_8_14_1647_0 & ~i_8_14_1870_0 & ~i_8_14_2041_0))) | (~i_8_14_248_0 & ((~i_8_14_499_0 & ~i_8_14_516_0 & ~i_8_14_925_0 & ~i_8_14_935_0 & i_8_14_1039_0 & ~i_8_14_1228_0) | (~i_8_14_356_0 & ~i_8_14_889_0 & ~i_8_14_958_0 & ~i_8_14_1232_0 & ~i_8_14_1241_0 & ~i_8_14_1285_0 & ~i_8_14_1497_0 & ~i_8_14_1919_0 & ~i_8_14_2066_0 & ~i_8_14_2249_0))) | (~i_8_14_518_0 & ~i_8_14_1387_0 & ((~i_8_14_359_0 & i_8_14_608_0 & ~i_8_14_1076_0 & ~i_8_14_1232_0 & ~i_8_14_1391_0) | (~i_8_14_799_0 & ~i_8_14_825_0 & ~i_8_14_935_0 & ~i_8_14_959_0 & ~i_8_14_1075_0 & ~i_8_14_1412_0 & ~i_8_14_1497_0 & ~i_8_14_1866_0 & ~i_8_14_1996_0))) | (~i_8_14_41_0 & ~i_8_14_273_0 & ~i_8_14_278_0 & ~i_8_14_385_0 & ~i_8_14_959_0 & ~i_8_14_1391_0 & ~i_8_14_1849_0 & ~i_8_14_2146_0))) | (~i_8_14_278_0 & ~i_8_14_958_0 & ~i_8_14_1178_0 & ((~i_8_14_248_0 & ~i_8_14_772_0 & ~i_8_14_955_0 & ~i_8_14_1192_0 & ~i_8_14_1274_0 & ~i_8_14_1800_0 & ~i_8_14_1849_0 & ~i_8_14_1906_0 & ~i_8_14_2040_0) | (~i_8_14_41_0 & ~i_8_14_170_0 & ~i_8_14_356_0 & ~i_8_14_499_0 & ~i_8_14_607_0 & ~i_8_14_608_0 & ~i_8_14_799_0 & ~i_8_14_1258_0 & ~i_8_14_1659_0 & ~i_8_14_2075_0 & ~i_8_14_2159_0))) | (~i_8_14_41_0 & ~i_8_14_2066_0 & ((~i_8_14_1087_0 & ~i_8_14_1232_0 & ~i_8_14_1273_0 & ~i_8_14_1385_0 & ~i_8_14_1807_0 & ~i_8_14_2041_0 & i_8_14_2146_0) | (~i_8_14_170_0 & ~i_8_14_516_0 & ~i_8_14_1075_0 & ~i_8_14_1241_0 & ~i_8_14_1391_0 & ~i_8_14_1412_0 & ~i_8_14_1645_0 & ~i_8_14_2146_0))) | (~i_8_14_2159_0 & ((~i_8_14_355_0 & ~i_8_14_799_0 & ((i_8_14_607_0 & ~i_8_14_994_0 & ~i_8_14_1075_0 & ~i_8_14_2041_0) | (~i_8_14_356_0 & ~i_8_14_364_0 & ~i_8_14_516_0 & ~i_8_14_592_0 & ~i_8_14_1391_0 & ~i_8_14_1866_0 & ~i_8_14_1870_0 & ~i_8_14_1940_0 & ~i_8_14_2219_0))) | (~i_8_14_170_0 & ~i_8_14_273_0 & ~i_8_14_499_0 & ~i_8_14_955_0 & i_8_14_1768_0 & ~i_8_14_2041_0))) | (i_8_14_889_0 & ~i_8_14_935_0 & i_8_14_994_0 & ~i_8_14_1866_0) | (~i_8_14_476_0 & i_8_14_484_0 & ~i_8_14_955_0 & ~i_8_14_1228_0 & ~i_8_14_1277_0 & ~i_8_14_1385_0 & i_8_14_1681_0) | (~i_8_14_597_0 & i_8_14_825_0 & i_8_14_1767_0 & ~i_8_14_1996_0 & i_8_14_2066_0) | (~i_8_14_356_0 & ~i_8_14_385_0 & ~i_8_14_634_0 & ~i_8_14_841_0 & ~i_8_14_1258_0 & ~i_8_14_1768_0 & ~i_8_14_1849_0 & ~i_8_14_1870_0 & ~i_8_14_2146_0 & ~i_8_14_2150_0));
endmodule



// Benchmark "kernel_8_15" written by ABC on Sun Jul 19 10:03:17 2020

module kernel_8_15 ( 
    i_8_15_5_0, i_8_15_19_0, i_8_15_76_0, i_8_15_83_0, i_8_15_112_0,
    i_8_15_140_0, i_8_15_148_0, i_8_15_150_0, i_8_15_169_0, i_8_15_173_0,
    i_8_15_192_0, i_8_15_193_0, i_8_15_226_0, i_8_15_239_0, i_8_15_245_0,
    i_8_15_274_0, i_8_15_275_0, i_8_15_325_0, i_8_15_335_0, i_8_15_341_0,
    i_8_15_353_0, i_8_15_361_0, i_8_15_364_0, i_8_15_365_0, i_8_15_442_0,
    i_8_15_515_0, i_8_15_581_0, i_8_15_587_0, i_8_15_596_0, i_8_15_652_0,
    i_8_15_667_0, i_8_15_668_0, i_8_15_680_0, i_8_15_703_0, i_8_15_704_0,
    i_8_15_707_0, i_8_15_730_0, i_8_15_733_0, i_8_15_751_0, i_8_15_756_0,
    i_8_15_830_0, i_8_15_910_0, i_8_15_911_0, i_8_15_968_0, i_8_15_1111_0,
    i_8_15_1129_0, i_8_15_1171_0, i_8_15_1297_0, i_8_15_1355_0,
    i_8_15_1483_0, i_8_15_1495_0, i_8_15_1521_0, i_8_15_1522_0,
    i_8_15_1531_0, i_8_15_1549_0, i_8_15_1594_0, i_8_15_1634_0,
    i_8_15_1651_0, i_8_15_1652_0, i_8_15_1682_0, i_8_15_1694_0,
    i_8_15_1705_0, i_8_15_1748_0, i_8_15_1765_0, i_8_15_1766_0,
    i_8_15_1774_0, i_8_15_1777_0, i_8_15_1805_0, i_8_15_1818_0,
    i_8_15_1819_0, i_8_15_1821_0, i_8_15_1822_0, i_8_15_1826_0,
    i_8_15_1857_0, i_8_15_1864_0, i_8_15_1874_0, i_8_15_1881_0,
    i_8_15_1892_0, i_8_15_1946_0, i_8_15_1967_0, i_8_15_1991_0,
    i_8_15_1994_0, i_8_15_1995_0, i_8_15_1996_0, i_8_15_2008_0,
    i_8_15_2009_0, i_8_15_2011_0, i_8_15_2062_0, i_8_15_2063_0,
    i_8_15_2074_0, i_8_15_2146_0, i_8_15_2147_0, i_8_15_2215_0,
    i_8_15_2227_0, i_8_15_2255_0, i_8_15_2256_0, i_8_15_2258_0,
    i_8_15_2269_0, i_8_15_2294_0, i_8_15_2300_0,
    o_8_15_0_0  );
  input  i_8_15_5_0, i_8_15_19_0, i_8_15_76_0, i_8_15_83_0, i_8_15_112_0,
    i_8_15_140_0, i_8_15_148_0, i_8_15_150_0, i_8_15_169_0, i_8_15_173_0,
    i_8_15_192_0, i_8_15_193_0, i_8_15_226_0, i_8_15_239_0, i_8_15_245_0,
    i_8_15_274_0, i_8_15_275_0, i_8_15_325_0, i_8_15_335_0, i_8_15_341_0,
    i_8_15_353_0, i_8_15_361_0, i_8_15_364_0, i_8_15_365_0, i_8_15_442_0,
    i_8_15_515_0, i_8_15_581_0, i_8_15_587_0, i_8_15_596_0, i_8_15_652_0,
    i_8_15_667_0, i_8_15_668_0, i_8_15_680_0, i_8_15_703_0, i_8_15_704_0,
    i_8_15_707_0, i_8_15_730_0, i_8_15_733_0, i_8_15_751_0, i_8_15_756_0,
    i_8_15_830_0, i_8_15_910_0, i_8_15_911_0, i_8_15_968_0, i_8_15_1111_0,
    i_8_15_1129_0, i_8_15_1171_0, i_8_15_1297_0, i_8_15_1355_0,
    i_8_15_1483_0, i_8_15_1495_0, i_8_15_1521_0, i_8_15_1522_0,
    i_8_15_1531_0, i_8_15_1549_0, i_8_15_1594_0, i_8_15_1634_0,
    i_8_15_1651_0, i_8_15_1652_0, i_8_15_1682_0, i_8_15_1694_0,
    i_8_15_1705_0, i_8_15_1748_0, i_8_15_1765_0, i_8_15_1766_0,
    i_8_15_1774_0, i_8_15_1777_0, i_8_15_1805_0, i_8_15_1818_0,
    i_8_15_1819_0, i_8_15_1821_0, i_8_15_1822_0, i_8_15_1826_0,
    i_8_15_1857_0, i_8_15_1864_0, i_8_15_1874_0, i_8_15_1881_0,
    i_8_15_1892_0, i_8_15_1946_0, i_8_15_1967_0, i_8_15_1991_0,
    i_8_15_1994_0, i_8_15_1995_0, i_8_15_1996_0, i_8_15_2008_0,
    i_8_15_2009_0, i_8_15_2011_0, i_8_15_2062_0, i_8_15_2063_0,
    i_8_15_2074_0, i_8_15_2146_0, i_8_15_2147_0, i_8_15_2215_0,
    i_8_15_2227_0, i_8_15_2255_0, i_8_15_2256_0, i_8_15_2258_0,
    i_8_15_2269_0, i_8_15_2294_0, i_8_15_2300_0;
  output o_8_15_0_0;
  assign o_8_15_0_0 = 0;
endmodule



// Benchmark "kernel_8_16" written by ABC on Sun Jul 19 10:03:18 2020

module kernel_8_16 ( 
    i_8_16_4_0, i_8_16_8_0, i_8_16_19_0, i_8_16_41_0, i_8_16_76_0,
    i_8_16_138_0, i_8_16_176_0, i_8_16_184_0, i_8_16_248_0, i_8_16_275_0,
    i_8_16_277_0, i_8_16_356_0, i_8_16_364_0, i_8_16_365_0, i_8_16_382_0,
    i_8_16_422_0, i_8_16_463_0, i_8_16_464_0, i_8_16_493_0, i_8_16_497_0,
    i_8_16_500_0, i_8_16_517_0, i_8_16_518_0, i_8_16_527_0, i_8_16_555_0,
    i_8_16_571_0, i_8_16_593_0, i_8_16_596_0, i_8_16_598_0, i_8_16_608_0,
    i_8_16_658_0, i_8_16_661_0, i_8_16_705_0, i_8_16_732_0, i_8_16_733_0,
    i_8_16_734_0, i_8_16_754_0, i_8_16_832_0, i_8_16_833_0, i_8_16_840_0,
    i_8_16_894_0, i_8_16_914_0, i_8_16_959_0, i_8_16_965_0, i_8_16_990_0,
    i_8_16_994_0, i_8_16_1073_0, i_8_16_1084_0, i_8_16_1175_0,
    i_8_16_1264_0, i_8_16_1298_0, i_8_16_1308_0, i_8_16_1331_0,
    i_8_16_1354_0, i_8_16_1358_0, i_8_16_1391_0, i_8_16_1466_0,
    i_8_16_1481_0, i_8_16_1484_0, i_8_16_1498_0, i_8_16_1499_0,
    i_8_16_1517_0, i_8_16_1534_0, i_8_16_1535_0, i_8_16_1597_0,
    i_8_16_1598_0, i_8_16_1654_0, i_8_16_1655_0, i_8_16_1660_0,
    i_8_16_1666_0, i_8_16_1678_0, i_8_16_1679_0, i_8_16_1695_0,
    i_8_16_1698_0, i_8_16_1777_0, i_8_16_1795_0, i_8_16_1812_0,
    i_8_16_1824_0, i_8_16_1826_0, i_8_16_1843_0, i_8_16_1849_0,
    i_8_16_1867_0, i_8_16_1876_0, i_8_16_1885_0, i_8_16_1894_0,
    i_8_16_1918_0, i_8_16_1951_0, i_8_16_1967_0, i_8_16_1995_0,
    i_8_16_2011_0, i_8_16_2039_0, i_8_16_2048_0, i_8_16_2172_0,
    i_8_16_2215_0, i_8_16_2227_0, i_8_16_2230_0, i_8_16_2234_0,
    i_8_16_2245_0, i_8_16_2284_0, i_8_16_2294_0,
    o_8_16_0_0  );
  input  i_8_16_4_0, i_8_16_8_0, i_8_16_19_0, i_8_16_41_0, i_8_16_76_0,
    i_8_16_138_0, i_8_16_176_0, i_8_16_184_0, i_8_16_248_0, i_8_16_275_0,
    i_8_16_277_0, i_8_16_356_0, i_8_16_364_0, i_8_16_365_0, i_8_16_382_0,
    i_8_16_422_0, i_8_16_463_0, i_8_16_464_0, i_8_16_493_0, i_8_16_497_0,
    i_8_16_500_0, i_8_16_517_0, i_8_16_518_0, i_8_16_527_0, i_8_16_555_0,
    i_8_16_571_0, i_8_16_593_0, i_8_16_596_0, i_8_16_598_0, i_8_16_608_0,
    i_8_16_658_0, i_8_16_661_0, i_8_16_705_0, i_8_16_732_0, i_8_16_733_0,
    i_8_16_734_0, i_8_16_754_0, i_8_16_832_0, i_8_16_833_0, i_8_16_840_0,
    i_8_16_894_0, i_8_16_914_0, i_8_16_959_0, i_8_16_965_0, i_8_16_990_0,
    i_8_16_994_0, i_8_16_1073_0, i_8_16_1084_0, i_8_16_1175_0,
    i_8_16_1264_0, i_8_16_1298_0, i_8_16_1308_0, i_8_16_1331_0,
    i_8_16_1354_0, i_8_16_1358_0, i_8_16_1391_0, i_8_16_1466_0,
    i_8_16_1481_0, i_8_16_1484_0, i_8_16_1498_0, i_8_16_1499_0,
    i_8_16_1517_0, i_8_16_1534_0, i_8_16_1535_0, i_8_16_1597_0,
    i_8_16_1598_0, i_8_16_1654_0, i_8_16_1655_0, i_8_16_1660_0,
    i_8_16_1666_0, i_8_16_1678_0, i_8_16_1679_0, i_8_16_1695_0,
    i_8_16_1698_0, i_8_16_1777_0, i_8_16_1795_0, i_8_16_1812_0,
    i_8_16_1824_0, i_8_16_1826_0, i_8_16_1843_0, i_8_16_1849_0,
    i_8_16_1867_0, i_8_16_1876_0, i_8_16_1885_0, i_8_16_1894_0,
    i_8_16_1918_0, i_8_16_1951_0, i_8_16_1967_0, i_8_16_1995_0,
    i_8_16_2011_0, i_8_16_2039_0, i_8_16_2048_0, i_8_16_2172_0,
    i_8_16_2215_0, i_8_16_2227_0, i_8_16_2230_0, i_8_16_2234_0,
    i_8_16_2245_0, i_8_16_2284_0, i_8_16_2294_0;
  output o_8_16_0_0;
  assign o_8_16_0_0 = 0;
endmodule



// Benchmark "kernel_8_17" written by ABC on Sun Jul 19 10:03:19 2020

module kernel_8_17 ( 
    i_8_17_27_0, i_8_17_28_0, i_8_17_34_0, i_8_17_51_0, i_8_17_82_0,
    i_8_17_85_0, i_8_17_93_0, i_8_17_156_0, i_8_17_199_0, i_8_17_233_0,
    i_8_17_243_0, i_8_17_252_0, i_8_17_255_0, i_8_17_288_0, i_8_17_297_0,
    i_8_17_324_0, i_8_17_342_0, i_8_17_345_0, i_8_17_371_0, i_8_17_378_0,
    i_8_17_435_0, i_8_17_436_0, i_8_17_450_0, i_8_17_471_0, i_8_17_530_0,
    i_8_17_551_0, i_8_17_562_0, i_8_17_565_0, i_8_17_585_0, i_8_17_586_0,
    i_8_17_615_0, i_8_17_621_0, i_8_17_624_0, i_8_17_633_0, i_8_17_637_0,
    i_8_17_657_0, i_8_17_665_0, i_8_17_666_0, i_8_17_669_0, i_8_17_694_0,
    i_8_17_700_0, i_8_17_715_0, i_8_17_810_0, i_8_17_972_0, i_8_17_973_0,
    i_8_17_975_0, i_8_17_990_0, i_8_17_1011_0, i_8_17_1188_0,
    i_8_17_1215_0, i_8_17_1216_0, i_8_17_1219_0, i_8_17_1224_0,
    i_8_17_1233_0, i_8_17_1247_0, i_8_17_1263_0, i_8_17_1278_0,
    i_8_17_1279_0, i_8_17_1284_0, i_8_17_1326_0, i_8_17_1345_0,
    i_8_17_1375_0, i_8_17_1434_0, i_8_17_1443_0, i_8_17_1503_0,
    i_8_17_1539_0, i_8_17_1584_0, i_8_17_1585_0, i_8_17_1587_0,
    i_8_17_1593_0, i_8_17_1594_0, i_8_17_1633_0, i_8_17_1665_0,
    i_8_17_1680_0, i_8_17_1701_0, i_8_17_1710_0, i_8_17_1751_0,
    i_8_17_1758_0, i_8_17_1799_0, i_8_17_1831_0, i_8_17_1845_0,
    i_8_17_1848_0, i_8_17_1854_0, i_8_17_1890_0, i_8_17_1899_0,
    i_8_17_1963_0, i_8_17_2043_0, i_8_17_2046_0, i_8_17_2092_0,
    i_8_17_2106_0, i_8_17_2110_0, i_8_17_2124_0, i_8_17_2126_0,
    i_8_17_2178_0, i_8_17_2179_0, i_8_17_2187_0, i_8_17_2259_0,
    i_8_17_2260_0, i_8_17_2269_0, i_8_17_2277_0,
    o_8_17_0_0  );
  input  i_8_17_27_0, i_8_17_28_0, i_8_17_34_0, i_8_17_51_0, i_8_17_82_0,
    i_8_17_85_0, i_8_17_93_0, i_8_17_156_0, i_8_17_199_0, i_8_17_233_0,
    i_8_17_243_0, i_8_17_252_0, i_8_17_255_0, i_8_17_288_0, i_8_17_297_0,
    i_8_17_324_0, i_8_17_342_0, i_8_17_345_0, i_8_17_371_0, i_8_17_378_0,
    i_8_17_435_0, i_8_17_436_0, i_8_17_450_0, i_8_17_471_0, i_8_17_530_0,
    i_8_17_551_0, i_8_17_562_0, i_8_17_565_0, i_8_17_585_0, i_8_17_586_0,
    i_8_17_615_0, i_8_17_621_0, i_8_17_624_0, i_8_17_633_0, i_8_17_637_0,
    i_8_17_657_0, i_8_17_665_0, i_8_17_666_0, i_8_17_669_0, i_8_17_694_0,
    i_8_17_700_0, i_8_17_715_0, i_8_17_810_0, i_8_17_972_0, i_8_17_973_0,
    i_8_17_975_0, i_8_17_990_0, i_8_17_1011_0, i_8_17_1188_0,
    i_8_17_1215_0, i_8_17_1216_0, i_8_17_1219_0, i_8_17_1224_0,
    i_8_17_1233_0, i_8_17_1247_0, i_8_17_1263_0, i_8_17_1278_0,
    i_8_17_1279_0, i_8_17_1284_0, i_8_17_1326_0, i_8_17_1345_0,
    i_8_17_1375_0, i_8_17_1434_0, i_8_17_1443_0, i_8_17_1503_0,
    i_8_17_1539_0, i_8_17_1584_0, i_8_17_1585_0, i_8_17_1587_0,
    i_8_17_1593_0, i_8_17_1594_0, i_8_17_1633_0, i_8_17_1665_0,
    i_8_17_1680_0, i_8_17_1701_0, i_8_17_1710_0, i_8_17_1751_0,
    i_8_17_1758_0, i_8_17_1799_0, i_8_17_1831_0, i_8_17_1845_0,
    i_8_17_1848_0, i_8_17_1854_0, i_8_17_1890_0, i_8_17_1899_0,
    i_8_17_1963_0, i_8_17_2043_0, i_8_17_2046_0, i_8_17_2092_0,
    i_8_17_2106_0, i_8_17_2110_0, i_8_17_2124_0, i_8_17_2126_0,
    i_8_17_2178_0, i_8_17_2179_0, i_8_17_2187_0, i_8_17_2259_0,
    i_8_17_2260_0, i_8_17_2269_0, i_8_17_2277_0;
  output o_8_17_0_0;
  assign o_8_17_0_0 = 0;
endmodule



// Benchmark "kernel_8_18" written by ABC on Sun Jul 19 10:03:20 2020

module kernel_8_18 ( 
    i_8_18_12_0, i_8_18_13_0, i_8_18_14_0, i_8_18_31_0, i_8_18_41_0,
    i_8_18_67_0, i_8_18_88_0, i_8_18_114_0, i_8_18_122_0, i_8_18_136_0,
    i_8_18_150_0, i_8_18_175_0, i_8_18_178_0, i_8_18_193_0, i_8_18_202_0,
    i_8_18_211_0, i_8_18_274_0, i_8_18_276_0, i_8_18_277_0, i_8_18_292_0,
    i_8_18_354_0, i_8_18_362_0, i_8_18_401_0, i_8_18_410_0, i_8_18_421_0,
    i_8_18_427_0, i_8_18_507_0, i_8_18_534_0, i_8_18_535_0, i_8_18_544_0,
    i_8_18_553_0, i_8_18_571_0, i_8_18_574_0, i_8_18_616_0, i_8_18_633_0,
    i_8_18_634_0, i_8_18_653_0, i_8_18_660_0, i_8_18_662_0, i_8_18_676_0,
    i_8_18_680_0, i_8_18_697_0, i_8_18_700_0, i_8_18_703_0, i_8_18_707_0,
    i_8_18_729_0, i_8_18_732_0, i_8_18_804_0, i_8_18_826_0, i_8_18_864_0,
    i_8_18_866_0, i_8_18_867_0, i_8_18_868_0, i_8_18_973_0, i_8_18_976_0,
    i_8_18_1031_0, i_8_18_1084_0, i_8_18_1102_0, i_8_18_1108_0,
    i_8_18_1153_0, i_8_18_1155_0, i_8_18_1174_0, i_8_18_1243_0,
    i_8_18_1245_0, i_8_18_1278_0, i_8_18_1299_0, i_8_18_1301_0,
    i_8_18_1314_0, i_8_18_1315_0, i_8_18_1336_0, i_8_18_1372_0,
    i_8_18_1387_0, i_8_18_1398_0, i_8_18_1405_0, i_8_18_1423_0,
    i_8_18_1440_0, i_8_18_1477_0, i_8_18_1525_0, i_8_18_1549_0,
    i_8_18_1576_0, i_8_18_1606_0, i_8_18_1642_0, i_8_18_1665_0,
    i_8_18_1683_0, i_8_18_1689_0, i_8_18_1791_0, i_8_18_1805_0,
    i_8_18_1822_0, i_8_18_1826_0, i_8_18_1884_0, i_8_18_1938_0,
    i_8_18_1995_0, i_8_18_2119_0, i_8_18_2147_0, i_8_18_2148_0,
    i_8_18_2173_0, i_8_18_2181_0, i_8_18_2188_0, i_8_18_2244_0,
    i_8_18_2272_0,
    o_8_18_0_0  );
  input  i_8_18_12_0, i_8_18_13_0, i_8_18_14_0, i_8_18_31_0, i_8_18_41_0,
    i_8_18_67_0, i_8_18_88_0, i_8_18_114_0, i_8_18_122_0, i_8_18_136_0,
    i_8_18_150_0, i_8_18_175_0, i_8_18_178_0, i_8_18_193_0, i_8_18_202_0,
    i_8_18_211_0, i_8_18_274_0, i_8_18_276_0, i_8_18_277_0, i_8_18_292_0,
    i_8_18_354_0, i_8_18_362_0, i_8_18_401_0, i_8_18_410_0, i_8_18_421_0,
    i_8_18_427_0, i_8_18_507_0, i_8_18_534_0, i_8_18_535_0, i_8_18_544_0,
    i_8_18_553_0, i_8_18_571_0, i_8_18_574_0, i_8_18_616_0, i_8_18_633_0,
    i_8_18_634_0, i_8_18_653_0, i_8_18_660_0, i_8_18_662_0, i_8_18_676_0,
    i_8_18_680_0, i_8_18_697_0, i_8_18_700_0, i_8_18_703_0, i_8_18_707_0,
    i_8_18_729_0, i_8_18_732_0, i_8_18_804_0, i_8_18_826_0, i_8_18_864_0,
    i_8_18_866_0, i_8_18_867_0, i_8_18_868_0, i_8_18_973_0, i_8_18_976_0,
    i_8_18_1031_0, i_8_18_1084_0, i_8_18_1102_0, i_8_18_1108_0,
    i_8_18_1153_0, i_8_18_1155_0, i_8_18_1174_0, i_8_18_1243_0,
    i_8_18_1245_0, i_8_18_1278_0, i_8_18_1299_0, i_8_18_1301_0,
    i_8_18_1314_0, i_8_18_1315_0, i_8_18_1336_0, i_8_18_1372_0,
    i_8_18_1387_0, i_8_18_1398_0, i_8_18_1405_0, i_8_18_1423_0,
    i_8_18_1440_0, i_8_18_1477_0, i_8_18_1525_0, i_8_18_1549_0,
    i_8_18_1576_0, i_8_18_1606_0, i_8_18_1642_0, i_8_18_1665_0,
    i_8_18_1683_0, i_8_18_1689_0, i_8_18_1791_0, i_8_18_1805_0,
    i_8_18_1822_0, i_8_18_1826_0, i_8_18_1884_0, i_8_18_1938_0,
    i_8_18_1995_0, i_8_18_2119_0, i_8_18_2147_0, i_8_18_2148_0,
    i_8_18_2173_0, i_8_18_2181_0, i_8_18_2188_0, i_8_18_2244_0,
    i_8_18_2272_0;
  output o_8_18_0_0;
  assign o_8_18_0_0 = 0;
endmodule



// Benchmark "kernel_8_19" written by ABC on Sun Jul 19 10:03:20 2020

module kernel_8_19 ( 
    i_8_19_52_0, i_8_19_57_0, i_8_19_58_0, i_8_19_59_0, i_8_19_87_0,
    i_8_19_88_0, i_8_19_142_0, i_8_19_143_0, i_8_19_166_0, i_8_19_168_0,
    i_8_19_169_0, i_8_19_229_0, i_8_19_230_0, i_8_19_233_0, i_8_19_257_0,
    i_8_19_258_0, i_8_19_260_0, i_8_19_328_0, i_8_19_329_0, i_8_19_369_0,
    i_8_19_370_0, i_8_19_377_0, i_8_19_379_0, i_8_19_421_0, i_8_19_437_0,
    i_8_19_483_0, i_8_19_485_0, i_8_19_502_0, i_8_19_508_0, i_8_19_522_0,
    i_8_19_529_0, i_8_19_530_0, i_8_19_552_0, i_8_19_553_0, i_8_19_556_0,
    i_8_19_557_0, i_8_19_596_0, i_8_19_633_0, i_8_19_634_0, i_8_19_635_0,
    i_8_19_689_0, i_8_19_691_0, i_8_19_692_0, i_8_19_735_0, i_8_19_736_0,
    i_8_19_752_0, i_8_19_762_0, i_8_19_768_0, i_8_19_815_0, i_8_19_850_0,
    i_8_19_868_0, i_8_19_993_0, i_8_19_994_0, i_8_19_1050_0, i_8_19_1051_0,
    i_8_19_1052_0, i_8_19_1057_0, i_8_19_1073_0, i_8_19_1110_0,
    i_8_19_1112_0, i_8_19_1119_0, i_8_19_1120_0, i_8_19_1188_0,
    i_8_19_1189_0, i_8_19_1292_0, i_8_19_1305_0, i_8_19_1306_0,
    i_8_19_1307_0, i_8_19_1315_0, i_8_19_1317_0, i_8_19_1327_0,
    i_8_19_1407_0, i_8_19_1437_0, i_8_19_1438_0, i_8_19_1506_0,
    i_8_19_1516_0, i_8_19_1560_0, i_8_19_1574_0, i_8_19_1631_0,
    i_8_19_1632_0, i_8_19_1633_0, i_8_19_1680_0, i_8_19_1684_0,
    i_8_19_1723_0, i_8_19_1749_0, i_8_19_1750_0, i_8_19_1754_0,
    i_8_19_1823_0, i_8_19_1861_0, i_8_19_1919_0, i_8_19_1958_0,
    i_8_19_1959_0, i_8_19_1960_0, i_8_19_1992_0, i_8_19_2003_0,
    i_8_19_2005_0, i_8_19_2032_0, i_8_19_2057_0, i_8_19_2093_0,
    i_8_19_2096_0,
    o_8_19_0_0  );
  input  i_8_19_52_0, i_8_19_57_0, i_8_19_58_0, i_8_19_59_0, i_8_19_87_0,
    i_8_19_88_0, i_8_19_142_0, i_8_19_143_0, i_8_19_166_0, i_8_19_168_0,
    i_8_19_169_0, i_8_19_229_0, i_8_19_230_0, i_8_19_233_0, i_8_19_257_0,
    i_8_19_258_0, i_8_19_260_0, i_8_19_328_0, i_8_19_329_0, i_8_19_369_0,
    i_8_19_370_0, i_8_19_377_0, i_8_19_379_0, i_8_19_421_0, i_8_19_437_0,
    i_8_19_483_0, i_8_19_485_0, i_8_19_502_0, i_8_19_508_0, i_8_19_522_0,
    i_8_19_529_0, i_8_19_530_0, i_8_19_552_0, i_8_19_553_0, i_8_19_556_0,
    i_8_19_557_0, i_8_19_596_0, i_8_19_633_0, i_8_19_634_0, i_8_19_635_0,
    i_8_19_689_0, i_8_19_691_0, i_8_19_692_0, i_8_19_735_0, i_8_19_736_0,
    i_8_19_752_0, i_8_19_762_0, i_8_19_768_0, i_8_19_815_0, i_8_19_850_0,
    i_8_19_868_0, i_8_19_993_0, i_8_19_994_0, i_8_19_1050_0, i_8_19_1051_0,
    i_8_19_1052_0, i_8_19_1057_0, i_8_19_1073_0, i_8_19_1110_0,
    i_8_19_1112_0, i_8_19_1119_0, i_8_19_1120_0, i_8_19_1188_0,
    i_8_19_1189_0, i_8_19_1292_0, i_8_19_1305_0, i_8_19_1306_0,
    i_8_19_1307_0, i_8_19_1315_0, i_8_19_1317_0, i_8_19_1327_0,
    i_8_19_1407_0, i_8_19_1437_0, i_8_19_1438_0, i_8_19_1506_0,
    i_8_19_1516_0, i_8_19_1560_0, i_8_19_1574_0, i_8_19_1631_0,
    i_8_19_1632_0, i_8_19_1633_0, i_8_19_1680_0, i_8_19_1684_0,
    i_8_19_1723_0, i_8_19_1749_0, i_8_19_1750_0, i_8_19_1754_0,
    i_8_19_1823_0, i_8_19_1861_0, i_8_19_1919_0, i_8_19_1958_0,
    i_8_19_1959_0, i_8_19_1960_0, i_8_19_1992_0, i_8_19_2003_0,
    i_8_19_2005_0, i_8_19_2032_0, i_8_19_2057_0, i_8_19_2093_0,
    i_8_19_2096_0;
  output o_8_19_0_0;
  assign o_8_19_0_0 = 0;
endmodule



// Benchmark "kernel_8_20" written by ABC on Sun Jul 19 10:03:21 2020

module kernel_8_20 ( 
    i_8_20_16_0, i_8_20_37_0, i_8_20_79_0, i_8_20_80_0, i_8_20_147_0,
    i_8_20_158_0, i_8_20_197_0, i_8_20_226_0, i_8_20_229_0, i_8_20_230_0,
    i_8_20_233_0, i_8_20_310_0, i_8_20_364_0, i_8_20_404_0, i_8_20_418_0,
    i_8_20_430_0, i_8_20_456_0, i_8_20_471_0, i_8_20_579_0, i_8_20_583_0,
    i_8_20_598_0, i_8_20_611_0, i_8_20_638_0, i_8_20_645_0, i_8_20_652_0,
    i_8_20_656_0, i_8_20_662_0, i_8_20_670_0, i_8_20_700_0, i_8_20_702_0,
    i_8_20_780_0, i_8_20_825_0, i_8_20_843_0, i_8_20_861_0, i_8_20_862_0,
    i_8_20_881_0, i_8_20_899_0, i_8_20_967_0, i_8_20_1015_0, i_8_20_1043_0,
    i_8_20_1089_0, i_8_20_1112_0, i_8_20_1129_0, i_8_20_1131_0,
    i_8_20_1187_0, i_8_20_1228_0, i_8_20_1263_0, i_8_20_1285_0,
    i_8_20_1299_0, i_8_20_1303_0, i_8_20_1310_0, i_8_20_1339_0,
    i_8_20_1340_0, i_8_20_1353_0, i_8_20_1384_0, i_8_20_1403_0,
    i_8_20_1426_0, i_8_20_1439_0, i_8_20_1474_0, i_8_20_1488_0,
    i_8_20_1489_0, i_8_20_1520_0, i_8_20_1545_0, i_8_20_1551_0,
    i_8_20_1552_0, i_8_20_1624_0, i_8_20_1628_0, i_8_20_1642_0,
    i_8_20_1653_0, i_8_20_1681_0, i_8_20_1706_0, i_8_20_1752_0,
    i_8_20_1771_0, i_8_20_1789_0, i_8_20_1806_0, i_8_20_1807_0,
    i_8_20_1812_0, i_8_20_1831_0, i_8_20_1843_0, i_8_20_1844_0,
    i_8_20_1854_0, i_8_20_1870_0, i_8_20_1875_0, i_8_20_1921_0,
    i_8_20_1943_0, i_8_20_1974_0, i_8_20_1978_0, i_8_20_1987_0,
    i_8_20_1993_0, i_8_20_2041_0, i_8_20_2091_0, i_8_20_2092_0,
    i_8_20_2110_0, i_8_20_2141_0, i_8_20_2215_0, i_8_20_2229_0,
    i_8_20_2238_0, i_8_20_2253_0, i_8_20_2265_0, i_8_20_2301_0,
    o_8_20_0_0  );
  input  i_8_20_16_0, i_8_20_37_0, i_8_20_79_0, i_8_20_80_0,
    i_8_20_147_0, i_8_20_158_0, i_8_20_197_0, i_8_20_226_0, i_8_20_229_0,
    i_8_20_230_0, i_8_20_233_0, i_8_20_310_0, i_8_20_364_0, i_8_20_404_0,
    i_8_20_418_0, i_8_20_430_0, i_8_20_456_0, i_8_20_471_0, i_8_20_579_0,
    i_8_20_583_0, i_8_20_598_0, i_8_20_611_0, i_8_20_638_0, i_8_20_645_0,
    i_8_20_652_0, i_8_20_656_0, i_8_20_662_0, i_8_20_670_0, i_8_20_700_0,
    i_8_20_702_0, i_8_20_780_0, i_8_20_825_0, i_8_20_843_0, i_8_20_861_0,
    i_8_20_862_0, i_8_20_881_0, i_8_20_899_0, i_8_20_967_0, i_8_20_1015_0,
    i_8_20_1043_0, i_8_20_1089_0, i_8_20_1112_0, i_8_20_1129_0,
    i_8_20_1131_0, i_8_20_1187_0, i_8_20_1228_0, i_8_20_1263_0,
    i_8_20_1285_0, i_8_20_1299_0, i_8_20_1303_0, i_8_20_1310_0,
    i_8_20_1339_0, i_8_20_1340_0, i_8_20_1353_0, i_8_20_1384_0,
    i_8_20_1403_0, i_8_20_1426_0, i_8_20_1439_0, i_8_20_1474_0,
    i_8_20_1488_0, i_8_20_1489_0, i_8_20_1520_0, i_8_20_1545_0,
    i_8_20_1551_0, i_8_20_1552_0, i_8_20_1624_0, i_8_20_1628_0,
    i_8_20_1642_0, i_8_20_1653_0, i_8_20_1681_0, i_8_20_1706_0,
    i_8_20_1752_0, i_8_20_1771_0, i_8_20_1789_0, i_8_20_1806_0,
    i_8_20_1807_0, i_8_20_1812_0, i_8_20_1831_0, i_8_20_1843_0,
    i_8_20_1844_0, i_8_20_1854_0, i_8_20_1870_0, i_8_20_1875_0,
    i_8_20_1921_0, i_8_20_1943_0, i_8_20_1974_0, i_8_20_1978_0,
    i_8_20_1987_0, i_8_20_1993_0, i_8_20_2041_0, i_8_20_2091_0,
    i_8_20_2092_0, i_8_20_2110_0, i_8_20_2141_0, i_8_20_2215_0,
    i_8_20_2229_0, i_8_20_2238_0, i_8_20_2253_0, i_8_20_2265_0,
    i_8_20_2301_0;
  output o_8_20_0_0;
  assign o_8_20_0_0 = 0;
endmodule



// Benchmark "kernel_8_21" written by ABC on Sun Jul 19 10:03:23 2020

module kernel_8_21 ( 
    i_8_21_28_0, i_8_21_29_0, i_8_21_60_0, i_8_21_138_0, i_8_21_139_0,
    i_8_21_158_0, i_8_21_159_0, i_8_21_166_0, i_8_21_193_0, i_8_21_229_0,
    i_8_21_230_0, i_8_21_232_0, i_8_21_363_0, i_8_21_364_0, i_8_21_365_0,
    i_8_21_366_0, i_8_21_368_0, i_8_21_381_0, i_8_21_484_0, i_8_21_510_0,
    i_8_21_528_0, i_8_21_657_0, i_8_21_661_0, i_8_21_687_0, i_8_21_688_0,
    i_8_21_690_0, i_8_21_691_0, i_8_21_692_0, i_8_21_695_0, i_8_21_707_0,
    i_8_21_709_0, i_8_21_762_0, i_8_21_763_0, i_8_21_764_0, i_8_21_822_0,
    i_8_21_827_0, i_8_21_844_0, i_8_21_845_0, i_8_21_868_0, i_8_21_994_0,
    i_8_21_1013_0, i_8_21_1026_0, i_8_21_1030_0, i_8_21_1033_0,
    i_8_21_1034_0, i_8_21_1051_0, i_8_21_1056_0, i_8_21_1059_0,
    i_8_21_1090_0, i_8_21_1115_0, i_8_21_1159_0, i_8_21_1160_0,
    i_8_21_1184_0, i_8_21_1255_0, i_8_21_1265_0, i_8_21_1296_0,
    i_8_21_1305_0, i_8_21_1306_0, i_8_21_1308_0, i_8_21_1310_0,
    i_8_21_1325_0, i_8_21_1344_0, i_8_21_1404_0, i_8_21_1556_0,
    i_8_21_1572_0, i_8_21_1634_0, i_8_21_1672_0, i_8_21_1674_0,
    i_8_21_1723_0, i_8_21_1741_0, i_8_21_1742_0, i_8_21_1743_0,
    i_8_21_1744_0, i_8_21_1745_0, i_8_21_1801_0, i_8_21_1805_0,
    i_8_21_1806_0, i_8_21_1808_0, i_8_21_1821_0, i_8_21_1822_0,
    i_8_21_1824_0, i_8_21_1825_0, i_8_21_1832_0, i_8_21_1834_0,
    i_8_21_1854_0, i_8_21_1918_0, i_8_21_2076_0, i_8_21_2119_0,
    i_8_21_2215_0, i_8_21_2216_0, i_8_21_2217_0, i_8_21_2224_0,
    i_8_21_2226_0, i_8_21_2233_0, i_8_21_2234_0, i_8_21_2271_0,
    i_8_21_2274_0, i_8_21_2275_0, i_8_21_2289_0, i_8_21_2290_0,
    o_8_21_0_0  );
  input  i_8_21_28_0, i_8_21_29_0, i_8_21_60_0, i_8_21_138_0,
    i_8_21_139_0, i_8_21_158_0, i_8_21_159_0, i_8_21_166_0, i_8_21_193_0,
    i_8_21_229_0, i_8_21_230_0, i_8_21_232_0, i_8_21_363_0, i_8_21_364_0,
    i_8_21_365_0, i_8_21_366_0, i_8_21_368_0, i_8_21_381_0, i_8_21_484_0,
    i_8_21_510_0, i_8_21_528_0, i_8_21_657_0, i_8_21_661_0, i_8_21_687_0,
    i_8_21_688_0, i_8_21_690_0, i_8_21_691_0, i_8_21_692_0, i_8_21_695_0,
    i_8_21_707_0, i_8_21_709_0, i_8_21_762_0, i_8_21_763_0, i_8_21_764_0,
    i_8_21_822_0, i_8_21_827_0, i_8_21_844_0, i_8_21_845_0, i_8_21_868_0,
    i_8_21_994_0, i_8_21_1013_0, i_8_21_1026_0, i_8_21_1030_0,
    i_8_21_1033_0, i_8_21_1034_0, i_8_21_1051_0, i_8_21_1056_0,
    i_8_21_1059_0, i_8_21_1090_0, i_8_21_1115_0, i_8_21_1159_0,
    i_8_21_1160_0, i_8_21_1184_0, i_8_21_1255_0, i_8_21_1265_0,
    i_8_21_1296_0, i_8_21_1305_0, i_8_21_1306_0, i_8_21_1308_0,
    i_8_21_1310_0, i_8_21_1325_0, i_8_21_1344_0, i_8_21_1404_0,
    i_8_21_1556_0, i_8_21_1572_0, i_8_21_1634_0, i_8_21_1672_0,
    i_8_21_1674_0, i_8_21_1723_0, i_8_21_1741_0, i_8_21_1742_0,
    i_8_21_1743_0, i_8_21_1744_0, i_8_21_1745_0, i_8_21_1801_0,
    i_8_21_1805_0, i_8_21_1806_0, i_8_21_1808_0, i_8_21_1821_0,
    i_8_21_1822_0, i_8_21_1824_0, i_8_21_1825_0, i_8_21_1832_0,
    i_8_21_1834_0, i_8_21_1854_0, i_8_21_1918_0, i_8_21_2076_0,
    i_8_21_2119_0, i_8_21_2215_0, i_8_21_2216_0, i_8_21_2217_0,
    i_8_21_2224_0, i_8_21_2226_0, i_8_21_2233_0, i_8_21_2234_0,
    i_8_21_2271_0, i_8_21_2274_0, i_8_21_2275_0, i_8_21_2289_0,
    i_8_21_2290_0;
  output o_8_21_0_0;
  assign o_8_21_0_0 = ~((~i_8_21_166_0 & ((~i_8_21_484_0 & i_8_21_690_0 & ~i_8_21_822_0 & ~i_8_21_1026_0 & ~i_8_21_1308_0 & ~i_8_21_1741_0 & ~i_8_21_1832_0 & ~i_8_21_2076_0 & ~i_8_21_2119_0 & ~i_8_21_2224_0 & ~i_8_21_2233_0) | (~i_8_21_29_0 & ~i_8_21_60_0 & ~i_8_21_158_0 & ~i_8_21_687_0 & ~i_8_21_688_0 & i_8_21_1090_0 & ~i_8_21_1184_0 & ~i_8_21_1310_0 & ~i_8_21_1742_0 & ~i_8_21_1805_0 & ~i_8_21_2234_0))) | (~i_8_21_158_0 & ((i_8_21_29_0 & ~i_8_21_138_0 & ~i_8_21_139_0 & i_8_21_695_0 & ~i_8_21_1090_0 & ~i_8_21_1805_0 & ~i_8_21_1821_0) | (~i_8_21_60_0 & ~i_8_21_232_0 & i_8_21_364_0 & ~i_8_21_1265_0 & ~i_8_21_1723_0 & ~i_8_21_2217_0 & ~i_8_21_2290_0))) | (~i_8_21_1743_0 & ((~i_8_21_2234_0 & ((~i_8_21_138_0 & ~i_8_21_484_0 & ~i_8_21_1741_0 & ((~i_8_21_29_0 & ~i_8_21_139_0 & ~i_8_21_193_0 & ~i_8_21_691_0 & ~i_8_21_695_0 & ~i_8_21_844_0 & ~i_8_21_1296_0 & ~i_8_21_1832_0 & i_8_21_1918_0) | (~i_8_21_510_0 & ~i_8_21_764_0 & ~i_8_21_1265_0 & ~i_8_21_1306_0 & ~i_8_21_1918_0 & ~i_8_21_2216_0))) | (i_8_21_661_0 & ~i_8_21_688_0 & ~i_8_21_1184_0 & ~i_8_21_1296_0 & ~i_8_21_2076_0 & ~i_8_21_2215_0))) | (~i_8_21_139_0 & ((~i_8_21_229_0 & ~i_8_21_1030_0 & i_8_21_1404_0 & ~i_8_21_1723_0 & i_8_21_1918_0) | (i_8_21_1034_0 & ~i_8_21_1745_0 & ~i_8_21_1832_0 & ~i_8_21_2119_0 & ~i_8_21_2290_0))) | (~i_8_21_1745_0 & ((~i_8_21_230_0 & ~i_8_21_845_0 & ~i_8_21_1059_0 & ~i_8_21_1184_0 & ~i_8_21_1325_0 & i_8_21_1801_0 & ~i_8_21_1854_0) | (~i_8_21_60_0 & ~i_8_21_510_0 & i_8_21_763_0 & ~i_8_21_1310_0 & ~i_8_21_1404_0 & ~i_8_21_1634_0 & ~i_8_21_1806_0 & ~i_8_21_2216_0))) | (~i_8_21_687_0 & ~i_8_21_764_0 & ~i_8_21_1090_0 & ~i_8_21_1296_0 & ~i_8_21_1742_0 & i_8_21_1801_0 & ~i_8_21_2076_0) | (~i_8_21_762_0 & ~i_8_21_763_0 & i_8_21_1824_0 & i_8_21_2215_0))) | (~i_8_21_1310_0 & ((~i_8_21_510_0 & ((i_8_21_365_0 & ~i_8_21_688_0 & ~i_8_21_763_0 & ~i_8_21_1634_0 & ~i_8_21_1723_0 & ~i_8_21_1744_0) | (~i_8_21_690_0 & i_8_21_1115_0 & ~i_8_21_1344_0 & i_8_21_1805_0))) | (~i_8_21_229_0 & ~i_8_21_690_0 & ~i_8_21_762_0 & ~i_8_21_1159_0 & ~i_8_21_1325_0 & ~i_8_21_1745_0 & i_8_21_1822_0))) | (~i_8_21_2216_0 & ((~i_8_21_1325_0 & ((~i_8_21_1306_0 & ((~i_8_21_29_0 & ~i_8_21_690_0 & ~i_8_21_1296_0 & ((~i_8_21_60_0 & ((~i_8_21_661_0 & ~i_8_21_687_0 & ~i_8_21_764_0 & ~i_8_21_1051_0 & ~i_8_21_1184_0 & ~i_8_21_1744_0 & ~i_8_21_1918_0) | (~i_8_21_139_0 & ~i_8_21_691_0 & ~i_8_21_692_0 & ~i_8_21_707_0 & ~i_8_21_1059_0 & ~i_8_21_1090_0 & ~i_8_21_1745_0 & ~i_8_21_2234_0))) | (~i_8_21_139_0 & ~i_8_21_229_0 & ~i_8_21_364_0 & ~i_8_21_366_0 & ~i_8_21_661_0 & ~i_8_21_687_0 & ~i_8_21_762_0 & ~i_8_21_764_0 & ~i_8_21_1059_0 & ~i_8_21_1832_0 & ~i_8_21_2215_0 & ~i_8_21_2233_0))) | (~i_8_21_687_0 & i_8_21_1090_0 & ~i_8_21_1742_0 & ~i_8_21_2217_0))) | (~i_8_21_28_0 & ~i_8_21_688_0 & ~i_8_21_691_0 & ~i_8_21_1305_0 & ~i_8_21_1742_0 & i_8_21_1918_0 & ~i_8_21_2233_0 & ~i_8_21_2234_0))) | (~i_8_21_1741_0 & ((~i_8_21_691_0 & i_8_21_845_0) | (i_8_21_695_0 & i_8_21_1805_0))) | (~i_8_21_60_0 & i_8_21_707_0 & ~i_8_21_1115_0 & ~i_8_21_1305_0 & ~i_8_21_1742_0 & i_8_21_1822_0))) | (~i_8_21_688_0 & ((~i_8_21_29_0 & ((~i_8_21_139_0 & i_8_21_1030_0 & ~i_8_21_1742_0 & ~i_8_21_1745_0) | (~i_8_21_1059_0 & ~i_8_21_1265_0 & i_8_21_1821_0))) | (~i_8_21_691_0 & ((~i_8_21_139_0 & ~i_8_21_695_0 & ~i_8_21_764_0 & ~i_8_21_1184_0 & i_8_21_1265_0 & ~i_8_21_1325_0 & ~i_8_21_2215_0) | (i_8_21_845_0 & ~i_8_21_1801_0 & ~i_8_21_2233_0))) | (i_8_21_707_0 & ~i_8_21_1296_0 & ~i_8_21_1305_0 & i_8_21_1634_0 & ~i_8_21_1742_0))) | (~i_8_21_229_0 & ((~i_8_21_29_0 & i_8_21_707_0 & ~i_8_21_1090_0 & ~i_8_21_1742_0 & ~i_8_21_1745_0 & ~i_8_21_1296_0 & ~i_8_21_1741_0) | (~i_8_21_692_0 & ~i_8_21_1744_0 & i_8_21_1808_0))) | (~i_8_21_687_0 & (i_8_21_2271_0 | (i_8_21_1824_0 & ~i_8_21_2217_0))) | (~i_8_21_690_0 & ((~i_8_21_692_0 & i_8_21_827_0 & ~i_8_21_1306_0) | (~i_8_21_1265_0 & ~i_8_21_1745_0 & i_8_21_1806_0 & ~i_8_21_1918_0 & ~i_8_21_2119_0 & ~i_8_21_2233_0))) | (~i_8_21_764_0 & ((i_8_21_1013_0 & ~i_8_21_1308_0 & ~i_8_21_1741_0) | (~i_8_21_365_0 & ~i_8_21_692_0 & ~i_8_21_994_0 & ~i_8_21_1059_0 & ~i_8_21_1184_0 & i_8_21_1556_0 & ~i_8_21_2215_0))) | (~i_8_21_1306_0 & ((~i_8_21_762_0 & ~i_8_21_1674_0 & i_8_21_1825_0 & ~i_8_21_2119_0) | (~i_8_21_230_0 & ~i_8_21_691_0 & i_8_21_1344_0 & ~i_8_21_1742_0 & ~i_8_21_2217_0))) | (~i_8_21_1742_0 & ((i_8_21_692_0 & ~i_8_21_1741_0 & i_8_21_1832_0 & ~i_8_21_1918_0) | (i_8_21_1854_0 & i_8_21_2234_0))) | (i_8_21_363_0 & ~i_8_21_763_0 & ~i_8_21_844_0 & ~i_8_21_1051_0 & ~i_8_21_1723_0) | (i_8_21_709_0 & i_8_21_1808_0) | (i_8_21_1743_0 & i_8_21_1806_0 & i_8_21_1918_0) | (~i_8_21_232_0 & ~i_8_21_1059_0 & i_8_21_1296_0 & i_8_21_1674_0 & ~i_8_21_1854_0 & ~i_8_21_2233_0));
endmodule



// Benchmark "kernel_8_22" written by ABC on Sun Jul 19 10:03:24 2020

module kernel_8_22 ( 
    i_8_22_9_0, i_8_22_49_0, i_8_22_118_0, i_8_22_126_0, i_8_22_300_0,
    i_8_22_360_0, i_8_22_361_0, i_8_22_382_0, i_8_22_390_0, i_8_22_391_0,
    i_8_22_399_0, i_8_22_400_0, i_8_22_417_0, i_8_22_426_0, i_8_22_453_0,
    i_8_22_504_0, i_8_22_505_0, i_8_22_558_0, i_8_22_559_0, i_8_22_561_0,
    i_8_22_568_0, i_8_22_639_0, i_8_22_640_0, i_8_22_660_0, i_8_22_661_0,
    i_8_22_676_0, i_8_22_679_0, i_8_22_696_0, i_8_22_697_0, i_8_22_702_0,
    i_8_22_766_0, i_8_22_783_0, i_8_22_784_0, i_8_22_847_0, i_8_22_891_0,
    i_8_22_892_0, i_8_22_969_0, i_8_22_999_0, i_8_22_1036_0, i_8_22_1045_0,
    i_8_22_1054_0, i_8_22_1102_0, i_8_22_1111_0, i_8_22_1130_0,
    i_8_22_1152_0, i_8_22_1179_0, i_8_22_1198_0, i_8_22_1234_0,
    i_8_22_1236_0, i_8_22_1263_0, i_8_22_1281_0, i_8_22_1295_0,
    i_8_22_1299_0, i_8_22_1339_0, i_8_22_1359_0, i_8_22_1360_0,
    i_8_22_1362_0, i_8_22_1363_0, i_8_22_1381_0, i_8_22_1399_0,
    i_8_22_1422_0, i_8_22_1423_0, i_8_22_1432_0, i_8_22_1440_0,
    i_8_22_1448_0, i_8_22_1450_0, i_8_22_1484_0, i_8_22_1486_0,
    i_8_22_1512_0, i_8_22_1513_0, i_8_22_1515_0, i_8_22_1521_0,
    i_8_22_1524_0, i_8_22_1551_0, i_8_22_1569_0, i_8_22_1639_0,
    i_8_22_1651_0, i_8_22_1656_0, i_8_22_1677_0, i_8_22_1678_0,
    i_8_22_1686_0, i_8_22_1746_0, i_8_22_1750_0, i_8_22_1767_0,
    i_8_22_1822_0, i_8_22_1839_0, i_8_22_1840_0, i_8_22_1845_0,
    i_8_22_1881_0, i_8_22_1974_0, i_8_22_1981_0, i_8_22_1992_0,
    i_8_22_2145_0, i_8_22_2147_0, i_8_22_2152_0, i_8_22_2190_0,
    i_8_22_2191_0, i_8_22_2224_0, i_8_22_2244_0, i_8_22_2245_0,
    o_8_22_0_0  );
  input  i_8_22_9_0, i_8_22_49_0, i_8_22_118_0, i_8_22_126_0,
    i_8_22_300_0, i_8_22_360_0, i_8_22_361_0, i_8_22_382_0, i_8_22_390_0,
    i_8_22_391_0, i_8_22_399_0, i_8_22_400_0, i_8_22_417_0, i_8_22_426_0,
    i_8_22_453_0, i_8_22_504_0, i_8_22_505_0, i_8_22_558_0, i_8_22_559_0,
    i_8_22_561_0, i_8_22_568_0, i_8_22_639_0, i_8_22_640_0, i_8_22_660_0,
    i_8_22_661_0, i_8_22_676_0, i_8_22_679_0, i_8_22_696_0, i_8_22_697_0,
    i_8_22_702_0, i_8_22_766_0, i_8_22_783_0, i_8_22_784_0, i_8_22_847_0,
    i_8_22_891_0, i_8_22_892_0, i_8_22_969_0, i_8_22_999_0, i_8_22_1036_0,
    i_8_22_1045_0, i_8_22_1054_0, i_8_22_1102_0, i_8_22_1111_0,
    i_8_22_1130_0, i_8_22_1152_0, i_8_22_1179_0, i_8_22_1198_0,
    i_8_22_1234_0, i_8_22_1236_0, i_8_22_1263_0, i_8_22_1281_0,
    i_8_22_1295_0, i_8_22_1299_0, i_8_22_1339_0, i_8_22_1359_0,
    i_8_22_1360_0, i_8_22_1362_0, i_8_22_1363_0, i_8_22_1381_0,
    i_8_22_1399_0, i_8_22_1422_0, i_8_22_1423_0, i_8_22_1432_0,
    i_8_22_1440_0, i_8_22_1448_0, i_8_22_1450_0, i_8_22_1484_0,
    i_8_22_1486_0, i_8_22_1512_0, i_8_22_1513_0, i_8_22_1515_0,
    i_8_22_1521_0, i_8_22_1524_0, i_8_22_1551_0, i_8_22_1569_0,
    i_8_22_1639_0, i_8_22_1651_0, i_8_22_1656_0, i_8_22_1677_0,
    i_8_22_1678_0, i_8_22_1686_0, i_8_22_1746_0, i_8_22_1750_0,
    i_8_22_1767_0, i_8_22_1822_0, i_8_22_1839_0, i_8_22_1840_0,
    i_8_22_1845_0, i_8_22_1881_0, i_8_22_1974_0, i_8_22_1981_0,
    i_8_22_1992_0, i_8_22_2145_0, i_8_22_2147_0, i_8_22_2152_0,
    i_8_22_2190_0, i_8_22_2191_0, i_8_22_2224_0, i_8_22_2244_0,
    i_8_22_2245_0;
  output o_8_22_0_0;
  assign o_8_22_0_0 = 0;
endmodule



// Benchmark "kernel_8_23" written by ABC on Sun Jul 19 10:03:25 2020

module kernel_8_23 ( 
    i_8_23_22_0, i_8_23_37_0, i_8_23_40_0, i_8_23_52_0, i_8_23_75_0,
    i_8_23_82_0, i_8_23_85_0, i_8_23_94_0, i_8_23_123_0, i_8_23_126_0,
    i_8_23_165_0, i_8_23_175_0, i_8_23_214_0, i_8_23_255_0, i_8_23_288_0,
    i_8_23_346_0, i_8_23_355_0, i_8_23_364_0, i_8_23_373_0, i_8_23_382_0,
    i_8_23_383_0, i_8_23_400_0, i_8_23_427_0, i_8_23_453_0, i_8_23_484_0,
    i_8_23_500_0, i_8_23_551_0, i_8_23_555_0, i_8_23_586_0, i_8_23_587_0,
    i_8_23_589_0, i_8_23_595_0, i_8_23_598_0, i_8_23_606_0, i_8_23_607_0,
    i_8_23_662_0, i_8_23_679_0, i_8_23_696_0, i_8_23_702_0, i_8_23_709_0,
    i_8_23_786_0, i_8_23_799_0, i_8_23_868_0, i_8_23_880_0, i_8_23_955_0,
    i_8_23_975_0, i_8_23_1020_0, i_8_23_1069_0, i_8_23_1071_0,
    i_8_23_1072_0, i_8_23_1090_0, i_8_23_1119_0, i_8_23_1123_0,
    i_8_23_1221_0, i_8_23_1227_0, i_8_23_1267_0, i_8_23_1272_0,
    i_8_23_1291_0, i_8_23_1298_0, i_8_23_1305_0, i_8_23_1308_0,
    i_8_23_1324_0, i_8_23_1327_0, i_8_23_1365_0, i_8_23_1470_0,
    i_8_23_1542_0, i_8_23_1606_0, i_8_23_1614_0, i_8_23_1626_0,
    i_8_23_1686_0, i_8_23_1749_0, i_8_23_1794_0, i_8_23_1821_0,
    i_8_23_1822_0, i_8_23_1824_0, i_8_23_1825_0, i_8_23_1830_0,
    i_8_23_1849_0, i_8_23_1855_0, i_8_23_1935_0, i_8_23_1938_0,
    i_8_23_1944_0, i_8_23_1993_0, i_8_23_1996_0, i_8_23_2002_0,
    i_8_23_2075_0, i_8_23_2103_0, i_8_23_2137_0, i_8_23_2142_0,
    i_8_23_2182_0, i_8_23_2212_0, i_8_23_2226_0, i_8_23_2227_0,
    i_8_23_2232_0, i_8_23_2235_0, i_8_23_2236_0, i_8_23_2245_0,
    i_8_23_2263_0, i_8_23_2280_0, i_8_23_2281_0,
    o_8_23_0_0  );
  input  i_8_23_22_0, i_8_23_37_0, i_8_23_40_0, i_8_23_52_0, i_8_23_75_0,
    i_8_23_82_0, i_8_23_85_0, i_8_23_94_0, i_8_23_123_0, i_8_23_126_0,
    i_8_23_165_0, i_8_23_175_0, i_8_23_214_0, i_8_23_255_0, i_8_23_288_0,
    i_8_23_346_0, i_8_23_355_0, i_8_23_364_0, i_8_23_373_0, i_8_23_382_0,
    i_8_23_383_0, i_8_23_400_0, i_8_23_427_0, i_8_23_453_0, i_8_23_484_0,
    i_8_23_500_0, i_8_23_551_0, i_8_23_555_0, i_8_23_586_0, i_8_23_587_0,
    i_8_23_589_0, i_8_23_595_0, i_8_23_598_0, i_8_23_606_0, i_8_23_607_0,
    i_8_23_662_0, i_8_23_679_0, i_8_23_696_0, i_8_23_702_0, i_8_23_709_0,
    i_8_23_786_0, i_8_23_799_0, i_8_23_868_0, i_8_23_880_0, i_8_23_955_0,
    i_8_23_975_0, i_8_23_1020_0, i_8_23_1069_0, i_8_23_1071_0,
    i_8_23_1072_0, i_8_23_1090_0, i_8_23_1119_0, i_8_23_1123_0,
    i_8_23_1221_0, i_8_23_1227_0, i_8_23_1267_0, i_8_23_1272_0,
    i_8_23_1291_0, i_8_23_1298_0, i_8_23_1305_0, i_8_23_1308_0,
    i_8_23_1324_0, i_8_23_1327_0, i_8_23_1365_0, i_8_23_1470_0,
    i_8_23_1542_0, i_8_23_1606_0, i_8_23_1614_0, i_8_23_1626_0,
    i_8_23_1686_0, i_8_23_1749_0, i_8_23_1794_0, i_8_23_1821_0,
    i_8_23_1822_0, i_8_23_1824_0, i_8_23_1825_0, i_8_23_1830_0,
    i_8_23_1849_0, i_8_23_1855_0, i_8_23_1935_0, i_8_23_1938_0,
    i_8_23_1944_0, i_8_23_1993_0, i_8_23_1996_0, i_8_23_2002_0,
    i_8_23_2075_0, i_8_23_2103_0, i_8_23_2137_0, i_8_23_2142_0,
    i_8_23_2182_0, i_8_23_2212_0, i_8_23_2226_0, i_8_23_2227_0,
    i_8_23_2232_0, i_8_23_2235_0, i_8_23_2236_0, i_8_23_2245_0,
    i_8_23_2263_0, i_8_23_2280_0, i_8_23_2281_0;
  output o_8_23_0_0;
  assign o_8_23_0_0 = 0;
endmodule



// Benchmark "kernel_8_24" written by ABC on Sun Jul 19 10:03:25 2020

module kernel_8_24 ( 
    i_8_24_34_0, i_8_24_69_0, i_8_24_78_0, i_8_24_79_0, i_8_24_115_0,
    i_8_24_133_0, i_8_24_169_0, i_8_24_250_0, i_8_24_312_0, i_8_24_337_0,
    i_8_24_380_0, i_8_24_384_0, i_8_24_475_0, i_8_24_500_0, i_8_24_501_0,
    i_8_24_511_0, i_8_24_519_0, i_8_24_525_0, i_8_24_528_0, i_8_24_539_0,
    i_8_24_553_0, i_8_24_555_0, i_8_24_574_0, i_8_24_583_0, i_8_24_600_0,
    i_8_24_628_0, i_8_24_637_0, i_8_24_664_0, i_8_24_673_0, i_8_24_733_0,
    i_8_24_750_0, i_8_24_834_0, i_8_24_843_0, i_8_24_916_0, i_8_24_1033_0,
    i_8_24_1087_0, i_8_24_1111_0, i_8_24_1177_0, i_8_24_1183_0,
    i_8_24_1245_0, i_8_24_1258_0, i_8_24_1273_0, i_8_24_1285_0,
    i_8_24_1291_0, i_8_24_1302_0, i_8_24_1303_0, i_8_24_1304_0,
    i_8_24_1365_0, i_8_24_1401_0, i_8_24_1407_0, i_8_24_1416_0,
    i_8_24_1438_0, i_8_24_1470_0, i_8_24_1489_0, i_8_24_1492_0,
    i_8_24_1501_0, i_8_24_1528_0, i_8_24_1536_0, i_8_24_1537_0,
    i_8_24_1544_0, i_8_24_1552_0, i_8_24_1608_0, i_8_24_1614_0,
    i_8_24_1653_0, i_8_24_1663_0, i_8_24_1672_0, i_8_24_1696_0,
    i_8_24_1702_0, i_8_24_1752_0, i_8_24_1762_0, i_8_24_1781_0,
    i_8_24_1794_0, i_8_24_1798_0, i_8_24_1816_0, i_8_24_1821_0,
    i_8_24_1851_0, i_8_24_1879_0, i_8_24_1884_0, i_8_24_1887_0,
    i_8_24_1898_0, i_8_24_1915_0, i_8_24_1951_0, i_8_24_1968_0,
    i_8_24_1970_0, i_8_24_2013_0, i_8_24_2041_0, i_8_24_2050_0,
    i_8_24_2064_0, i_8_24_2122_0, i_8_24_2153_0, i_8_24_2176_0,
    i_8_24_2186_0, i_8_24_2216_0, i_8_24_2218_0, i_8_24_2219_0,
    i_8_24_2228_0, i_8_24_2229_0, i_8_24_2247_0, i_8_24_2248_0,
    i_8_24_2257_0,
    o_8_24_0_0  );
  input  i_8_24_34_0, i_8_24_69_0, i_8_24_78_0, i_8_24_79_0,
    i_8_24_115_0, i_8_24_133_0, i_8_24_169_0, i_8_24_250_0, i_8_24_312_0,
    i_8_24_337_0, i_8_24_380_0, i_8_24_384_0, i_8_24_475_0, i_8_24_500_0,
    i_8_24_501_0, i_8_24_511_0, i_8_24_519_0, i_8_24_525_0, i_8_24_528_0,
    i_8_24_539_0, i_8_24_553_0, i_8_24_555_0, i_8_24_574_0, i_8_24_583_0,
    i_8_24_600_0, i_8_24_628_0, i_8_24_637_0, i_8_24_664_0, i_8_24_673_0,
    i_8_24_733_0, i_8_24_750_0, i_8_24_834_0, i_8_24_843_0, i_8_24_916_0,
    i_8_24_1033_0, i_8_24_1087_0, i_8_24_1111_0, i_8_24_1177_0,
    i_8_24_1183_0, i_8_24_1245_0, i_8_24_1258_0, i_8_24_1273_0,
    i_8_24_1285_0, i_8_24_1291_0, i_8_24_1302_0, i_8_24_1303_0,
    i_8_24_1304_0, i_8_24_1365_0, i_8_24_1401_0, i_8_24_1407_0,
    i_8_24_1416_0, i_8_24_1438_0, i_8_24_1470_0, i_8_24_1489_0,
    i_8_24_1492_0, i_8_24_1501_0, i_8_24_1528_0, i_8_24_1536_0,
    i_8_24_1537_0, i_8_24_1544_0, i_8_24_1552_0, i_8_24_1608_0,
    i_8_24_1614_0, i_8_24_1653_0, i_8_24_1663_0, i_8_24_1672_0,
    i_8_24_1696_0, i_8_24_1702_0, i_8_24_1752_0, i_8_24_1762_0,
    i_8_24_1781_0, i_8_24_1794_0, i_8_24_1798_0, i_8_24_1816_0,
    i_8_24_1821_0, i_8_24_1851_0, i_8_24_1879_0, i_8_24_1884_0,
    i_8_24_1887_0, i_8_24_1898_0, i_8_24_1915_0, i_8_24_1951_0,
    i_8_24_1968_0, i_8_24_1970_0, i_8_24_2013_0, i_8_24_2041_0,
    i_8_24_2050_0, i_8_24_2064_0, i_8_24_2122_0, i_8_24_2153_0,
    i_8_24_2176_0, i_8_24_2186_0, i_8_24_2216_0, i_8_24_2218_0,
    i_8_24_2219_0, i_8_24_2228_0, i_8_24_2229_0, i_8_24_2247_0,
    i_8_24_2248_0, i_8_24_2257_0;
  output o_8_24_0_0;
  assign o_8_24_0_0 = 0;
endmodule



// Benchmark "kernel_8_25" written by ABC on Sun Jul 19 10:03:26 2020

module kernel_8_25 ( 
    i_8_25_20_0, i_8_25_27_0, i_8_25_44_0, i_8_25_48_0, i_8_25_54_0,
    i_8_25_87_0, i_8_25_108_0, i_8_25_115_0, i_8_25_220_0, i_8_25_304_0,
    i_8_25_325_0, i_8_25_345_0, i_8_25_355_0, i_8_25_365_0, i_8_25_489_0,
    i_8_25_491_0, i_8_25_553_0, i_8_25_571_0, i_8_25_606_0, i_8_25_607_0,
    i_8_25_613_0, i_8_25_617_0, i_8_25_643_0, i_8_25_651_0, i_8_25_655_0,
    i_8_25_675_0, i_8_25_694_0, i_8_25_698_0, i_8_25_701_0, i_8_25_782_0,
    i_8_25_791_0, i_8_25_802_0, i_8_25_876_0, i_8_25_882_0, i_8_25_993_0,
    i_8_25_1038_0, i_8_25_1040_0, i_8_25_1054_0, i_8_25_1071_0,
    i_8_25_1074_0, i_8_25_1093_0, i_8_25_1094_0, i_8_25_1098_0,
    i_8_25_1102_0, i_8_25_1125_0, i_8_25_1131_0, i_8_25_1137_0,
    i_8_25_1142_0, i_8_25_1146_0, i_8_25_1147_0, i_8_25_1164_0,
    i_8_25_1224_0, i_8_25_1237_0, i_8_25_1254_0, i_8_25_1313_0,
    i_8_25_1318_0, i_8_25_1322_0, i_8_25_1330_0, i_8_25_1351_0,
    i_8_25_1362_0, i_8_25_1422_0, i_8_25_1482_0, i_8_25_1526_0,
    i_8_25_1549_0, i_8_25_1600_0, i_8_25_1607_0, i_8_25_1621_0,
    i_8_25_1654_0, i_8_25_1677_0, i_8_25_1704_0, i_8_25_1737_0,
    i_8_25_1738_0, i_8_25_1739_0, i_8_25_1741_0, i_8_25_1770_0,
    i_8_25_1790_0, i_8_25_1804_0, i_8_25_1806_0, i_8_25_1808_0,
    i_8_25_1809_0, i_8_25_1821_0, i_8_25_1822_0, i_8_25_1949_0,
    i_8_25_1958_0, i_8_25_1966_0, i_8_25_1983_0, i_8_25_1995_0,
    i_8_25_2055_0, i_8_25_2058_0, i_8_25_2076_0, i_8_25_2097_0,
    i_8_25_2101_0, i_8_25_2104_0, i_8_25_2124_0, i_8_25_2154_0,
    i_8_25_2163_0, i_8_25_2173_0, i_8_25_2190_0, i_8_25_2191_0,
    i_8_25_2233_0,
    o_8_25_0_0  );
  input  i_8_25_20_0, i_8_25_27_0, i_8_25_44_0, i_8_25_48_0, i_8_25_54_0,
    i_8_25_87_0, i_8_25_108_0, i_8_25_115_0, i_8_25_220_0, i_8_25_304_0,
    i_8_25_325_0, i_8_25_345_0, i_8_25_355_0, i_8_25_365_0, i_8_25_489_0,
    i_8_25_491_0, i_8_25_553_0, i_8_25_571_0, i_8_25_606_0, i_8_25_607_0,
    i_8_25_613_0, i_8_25_617_0, i_8_25_643_0, i_8_25_651_0, i_8_25_655_0,
    i_8_25_675_0, i_8_25_694_0, i_8_25_698_0, i_8_25_701_0, i_8_25_782_0,
    i_8_25_791_0, i_8_25_802_0, i_8_25_876_0, i_8_25_882_0, i_8_25_993_0,
    i_8_25_1038_0, i_8_25_1040_0, i_8_25_1054_0, i_8_25_1071_0,
    i_8_25_1074_0, i_8_25_1093_0, i_8_25_1094_0, i_8_25_1098_0,
    i_8_25_1102_0, i_8_25_1125_0, i_8_25_1131_0, i_8_25_1137_0,
    i_8_25_1142_0, i_8_25_1146_0, i_8_25_1147_0, i_8_25_1164_0,
    i_8_25_1224_0, i_8_25_1237_0, i_8_25_1254_0, i_8_25_1313_0,
    i_8_25_1318_0, i_8_25_1322_0, i_8_25_1330_0, i_8_25_1351_0,
    i_8_25_1362_0, i_8_25_1422_0, i_8_25_1482_0, i_8_25_1526_0,
    i_8_25_1549_0, i_8_25_1600_0, i_8_25_1607_0, i_8_25_1621_0,
    i_8_25_1654_0, i_8_25_1677_0, i_8_25_1704_0, i_8_25_1737_0,
    i_8_25_1738_0, i_8_25_1739_0, i_8_25_1741_0, i_8_25_1770_0,
    i_8_25_1790_0, i_8_25_1804_0, i_8_25_1806_0, i_8_25_1808_0,
    i_8_25_1809_0, i_8_25_1821_0, i_8_25_1822_0, i_8_25_1949_0,
    i_8_25_1958_0, i_8_25_1966_0, i_8_25_1983_0, i_8_25_1995_0,
    i_8_25_2055_0, i_8_25_2058_0, i_8_25_2076_0, i_8_25_2097_0,
    i_8_25_2101_0, i_8_25_2104_0, i_8_25_2124_0, i_8_25_2154_0,
    i_8_25_2163_0, i_8_25_2173_0, i_8_25_2190_0, i_8_25_2191_0,
    i_8_25_2233_0;
  output o_8_25_0_0;
  assign o_8_25_0_0 = 0;
endmodule



// Benchmark "kernel_8_26" written by ABC on Sun Jul 19 10:03:27 2020

module kernel_8_26 ( 
    i_8_26_19_0, i_8_26_32_0, i_8_26_33_0, i_8_26_138_0, i_8_26_153_0,
    i_8_26_157_0, i_8_26_184_0, i_8_26_193_0, i_8_26_373_0, i_8_26_379_0,
    i_8_26_387_0, i_8_26_388_0, i_8_26_436_0, i_8_26_441_0, i_8_26_442_0,
    i_8_26_479_0, i_8_26_495_0, i_8_26_496_0, i_8_26_507_0, i_8_26_508_0,
    i_8_26_525_0, i_8_26_526_0, i_8_26_536_0, i_8_26_551_0, i_8_26_554_0,
    i_8_26_586_0, i_8_26_604_0, i_8_26_613_0, i_8_26_660_0, i_8_26_662_0,
    i_8_26_666_0, i_8_26_678_0, i_8_26_760_0, i_8_26_761_0, i_8_26_769_0,
    i_8_26_819_0, i_8_26_822_0, i_8_26_823_0, i_8_26_824_0, i_8_26_864_0,
    i_8_26_865_0, i_8_26_918_0, i_8_26_922_0, i_8_26_981_0, i_8_26_982_0,
    i_8_26_983_0, i_8_26_1008_0, i_8_26_1030_0, i_8_26_1108_0,
    i_8_26_1112_0, i_8_26_1129_0, i_8_26_1130_0, i_8_26_1153_0,
    i_8_26_1233_0, i_8_26_1236_0, i_8_26_1242_0, i_8_26_1243_0,
    i_8_26_1245_0, i_8_26_1246_0, i_8_26_1252_0, i_8_26_1263_0,
    i_8_26_1264_0, i_8_26_1278_0, i_8_26_1279_0, i_8_26_1323_0,
    i_8_26_1341_0, i_8_26_1400_0, i_8_26_1435_0, i_8_26_1503_0,
    i_8_26_1506_0, i_8_26_1513_0, i_8_26_1530_0, i_8_26_1531_0,
    i_8_26_1550_0, i_8_26_1561_0, i_8_26_1576_0, i_8_26_1594_0,
    i_8_26_1611_0, i_8_26_1614_0, i_8_26_1647_0, i_8_26_1667_0,
    i_8_26_1755_0, i_8_26_1756_0, i_8_26_1777_0, i_8_26_1785_0,
    i_8_26_1800_0, i_8_26_1837_0, i_8_26_1848_0, i_8_26_1890_0,
    i_8_26_1943_0, i_8_26_1999_0, i_8_26_2037_0, i_8_26_2043_0,
    i_8_26_2106_0, i_8_26_2107_0, i_8_26_2178_0, i_8_26_2223_0,
    i_8_26_2236_0, i_8_26_2237_0, i_8_26_2245_0,
    o_8_26_0_0  );
  input  i_8_26_19_0, i_8_26_32_0, i_8_26_33_0, i_8_26_138_0,
    i_8_26_153_0, i_8_26_157_0, i_8_26_184_0, i_8_26_193_0, i_8_26_373_0,
    i_8_26_379_0, i_8_26_387_0, i_8_26_388_0, i_8_26_436_0, i_8_26_441_0,
    i_8_26_442_0, i_8_26_479_0, i_8_26_495_0, i_8_26_496_0, i_8_26_507_0,
    i_8_26_508_0, i_8_26_525_0, i_8_26_526_0, i_8_26_536_0, i_8_26_551_0,
    i_8_26_554_0, i_8_26_586_0, i_8_26_604_0, i_8_26_613_0, i_8_26_660_0,
    i_8_26_662_0, i_8_26_666_0, i_8_26_678_0, i_8_26_760_0, i_8_26_761_0,
    i_8_26_769_0, i_8_26_819_0, i_8_26_822_0, i_8_26_823_0, i_8_26_824_0,
    i_8_26_864_0, i_8_26_865_0, i_8_26_918_0, i_8_26_922_0, i_8_26_981_0,
    i_8_26_982_0, i_8_26_983_0, i_8_26_1008_0, i_8_26_1030_0,
    i_8_26_1108_0, i_8_26_1112_0, i_8_26_1129_0, i_8_26_1130_0,
    i_8_26_1153_0, i_8_26_1233_0, i_8_26_1236_0, i_8_26_1242_0,
    i_8_26_1243_0, i_8_26_1245_0, i_8_26_1246_0, i_8_26_1252_0,
    i_8_26_1263_0, i_8_26_1264_0, i_8_26_1278_0, i_8_26_1279_0,
    i_8_26_1323_0, i_8_26_1341_0, i_8_26_1400_0, i_8_26_1435_0,
    i_8_26_1503_0, i_8_26_1506_0, i_8_26_1513_0, i_8_26_1530_0,
    i_8_26_1531_0, i_8_26_1550_0, i_8_26_1561_0, i_8_26_1576_0,
    i_8_26_1594_0, i_8_26_1611_0, i_8_26_1614_0, i_8_26_1647_0,
    i_8_26_1667_0, i_8_26_1755_0, i_8_26_1756_0, i_8_26_1777_0,
    i_8_26_1785_0, i_8_26_1800_0, i_8_26_1837_0, i_8_26_1848_0,
    i_8_26_1890_0, i_8_26_1943_0, i_8_26_1999_0, i_8_26_2037_0,
    i_8_26_2043_0, i_8_26_2106_0, i_8_26_2107_0, i_8_26_2178_0,
    i_8_26_2223_0, i_8_26_2236_0, i_8_26_2237_0, i_8_26_2245_0;
  output o_8_26_0_0;
  assign o_8_26_0_0 = 0;
endmodule



// Benchmark "kernel_8_27" written by ABC on Sun Jul 19 10:03:28 2020

module kernel_8_27 ( 
    i_8_27_4_0, i_8_27_5_0, i_8_27_25_0, i_8_27_35_0, i_8_27_44_0,
    i_8_27_77_0, i_8_27_87_0, i_8_27_148_0, i_8_27_211_0, i_8_27_230_0,
    i_8_27_244_0, i_8_27_247_0, i_8_27_248_0, i_8_27_274_0, i_8_27_275_0,
    i_8_27_323_0, i_8_27_363_0, i_8_27_368_0, i_8_27_385_0, i_8_27_421_0,
    i_8_27_422_0, i_8_27_431_0, i_8_27_527_0, i_8_27_528_0, i_8_27_530_0,
    i_8_27_565_0, i_8_27_571_0, i_8_27_572_0, i_8_27_575_0, i_8_27_582_0,
    i_8_27_583_0, i_8_27_586_0, i_8_27_644_0, i_8_27_652_0, i_8_27_655_0,
    i_8_27_670_0, i_8_27_671_0, i_8_27_681_0, i_8_27_682_0, i_8_27_696_0,
    i_8_27_703_0, i_8_27_706_0, i_8_27_733_0, i_8_27_734_0, i_8_27_760_0,
    i_8_27_781_0, i_8_27_844_0, i_8_27_850_0, i_8_27_859_0, i_8_27_889_0,
    i_8_27_943_0, i_8_27_956_0, i_8_27_991_0, i_8_27_992_0, i_8_27_1105_0,
    i_8_27_1111_0, i_8_27_1129_0, i_8_27_1132_0, i_8_27_1172_0,
    i_8_27_1321_0, i_8_27_1329_0, i_8_27_1330_0, i_8_27_1354_0,
    i_8_27_1355_0, i_8_27_1358_0, i_8_27_1382_0, i_8_27_1399_0,
    i_8_27_1400_0, i_8_27_1465_0, i_8_27_1468_0, i_8_27_1480_0,
    i_8_27_1481_0, i_8_27_1518_0, i_8_27_1531_0, i_8_27_1535_0,
    i_8_27_1541_0, i_8_27_1598_0, i_8_27_1699_0, i_8_27_1703_0,
    i_8_27_1705_0, i_8_27_1753_0, i_8_27_1754_0, i_8_27_1772_0,
    i_8_27_1795_0, i_8_27_1796_0, i_8_27_1804_0, i_8_27_1807_0,
    i_8_27_1813_0, i_8_27_1843_0, i_8_27_1928_0, i_8_27_1960_0,
    i_8_27_2042_0, i_8_27_2065_0, i_8_27_2066_0, i_8_27_2194_0,
    i_8_27_2216_0, i_8_27_2244_0, i_8_27_2254_0, i_8_27_2255_0,
    i_8_27_2256_0,
    o_8_27_0_0  );
  input  i_8_27_4_0, i_8_27_5_0, i_8_27_25_0, i_8_27_35_0, i_8_27_44_0,
    i_8_27_77_0, i_8_27_87_0, i_8_27_148_0, i_8_27_211_0, i_8_27_230_0,
    i_8_27_244_0, i_8_27_247_0, i_8_27_248_0, i_8_27_274_0, i_8_27_275_0,
    i_8_27_323_0, i_8_27_363_0, i_8_27_368_0, i_8_27_385_0, i_8_27_421_0,
    i_8_27_422_0, i_8_27_431_0, i_8_27_527_0, i_8_27_528_0, i_8_27_530_0,
    i_8_27_565_0, i_8_27_571_0, i_8_27_572_0, i_8_27_575_0, i_8_27_582_0,
    i_8_27_583_0, i_8_27_586_0, i_8_27_644_0, i_8_27_652_0, i_8_27_655_0,
    i_8_27_670_0, i_8_27_671_0, i_8_27_681_0, i_8_27_682_0, i_8_27_696_0,
    i_8_27_703_0, i_8_27_706_0, i_8_27_733_0, i_8_27_734_0, i_8_27_760_0,
    i_8_27_781_0, i_8_27_844_0, i_8_27_850_0, i_8_27_859_0, i_8_27_889_0,
    i_8_27_943_0, i_8_27_956_0, i_8_27_991_0, i_8_27_992_0, i_8_27_1105_0,
    i_8_27_1111_0, i_8_27_1129_0, i_8_27_1132_0, i_8_27_1172_0,
    i_8_27_1321_0, i_8_27_1329_0, i_8_27_1330_0, i_8_27_1354_0,
    i_8_27_1355_0, i_8_27_1358_0, i_8_27_1382_0, i_8_27_1399_0,
    i_8_27_1400_0, i_8_27_1465_0, i_8_27_1468_0, i_8_27_1480_0,
    i_8_27_1481_0, i_8_27_1518_0, i_8_27_1531_0, i_8_27_1535_0,
    i_8_27_1541_0, i_8_27_1598_0, i_8_27_1699_0, i_8_27_1703_0,
    i_8_27_1705_0, i_8_27_1753_0, i_8_27_1754_0, i_8_27_1772_0,
    i_8_27_1795_0, i_8_27_1796_0, i_8_27_1804_0, i_8_27_1807_0,
    i_8_27_1813_0, i_8_27_1843_0, i_8_27_1928_0, i_8_27_1960_0,
    i_8_27_2042_0, i_8_27_2065_0, i_8_27_2066_0, i_8_27_2194_0,
    i_8_27_2216_0, i_8_27_2244_0, i_8_27_2254_0, i_8_27_2255_0,
    i_8_27_2256_0;
  output o_8_27_0_0;
  assign o_8_27_0_0 = 0;
endmodule



// Benchmark "kernel_8_28" written by ABC on Sun Jul 19 10:03:28 2020

module kernel_8_28 ( 
    i_8_28_1_0, i_8_28_19_0, i_8_28_20_0, i_8_28_85_0, i_8_28_118_0,
    i_8_28_136_0, i_8_28_143_0, i_8_28_144_0, i_8_28_190_0, i_8_28_202_0,
    i_8_28_352_0, i_8_28_381_0, i_8_28_382_0, i_8_28_391_0, i_8_28_414_0,
    i_8_28_442_0, i_8_28_469_0, i_8_28_514_0, i_8_28_522_0, i_8_28_523_0,
    i_8_28_524_0, i_8_28_525_0, i_8_28_567_0, i_8_28_577_0, i_8_28_595_0,
    i_8_28_596_0, i_8_28_607_0, i_8_28_610_0, i_8_28_631_0, i_8_28_634_0,
    i_8_28_637_0, i_8_28_658_0, i_8_28_667_0, i_8_28_702_0, i_8_28_703_0,
    i_8_28_712_0, i_8_28_748_0, i_8_28_751_0, i_8_28_829_0, i_8_28_838_0,
    i_8_28_844_0, i_8_28_859_0, i_8_28_881_0, i_8_28_910_0, i_8_28_929_0,
    i_8_28_955_0, i_8_28_964_0, i_8_28_967_0, i_8_28_968_0, i_8_28_997_0,
    i_8_28_1179_0, i_8_28_1198_0, i_8_28_1234_0, i_8_28_1252_0,
    i_8_28_1282_0, i_8_28_1354_0, i_8_28_1387_0, i_8_28_1396_0,
    i_8_28_1467_0, i_8_28_1468_0, i_8_28_1486_0, i_8_28_1495_0,
    i_8_28_1507_0, i_8_28_1531_0, i_8_28_1533_0, i_8_28_1536_0,
    i_8_28_1594_0, i_8_28_1629_0, i_8_28_1639_0, i_8_28_1647_0,
    i_8_28_1657_0, i_8_28_1702_0, i_8_28_1703_0, i_8_28_1747_0,
    i_8_28_1757_0, i_8_28_1774_0, i_8_28_1775_0, i_8_28_1791_0,
    i_8_28_1792_0, i_8_28_1801_0, i_8_28_1802_0, i_8_28_1818_0,
    i_8_28_1819_0, i_8_28_1822_0, i_8_28_1846_0, i_8_28_1864_0,
    i_8_28_1873_0, i_8_28_1900_0, i_8_28_1910_0, i_8_28_1963_0,
    i_8_28_2008_0, i_8_28_2044_0, i_8_28_2062_0, i_8_28_2089_0,
    i_8_28_2116_0, i_8_28_2133_0, i_8_28_2134_0, i_8_28_2173_0,
    i_8_28_2227_0, i_8_28_2284_0,
    o_8_28_0_0  );
  input  i_8_28_1_0, i_8_28_19_0, i_8_28_20_0, i_8_28_85_0, i_8_28_118_0,
    i_8_28_136_0, i_8_28_143_0, i_8_28_144_0, i_8_28_190_0, i_8_28_202_0,
    i_8_28_352_0, i_8_28_381_0, i_8_28_382_0, i_8_28_391_0, i_8_28_414_0,
    i_8_28_442_0, i_8_28_469_0, i_8_28_514_0, i_8_28_522_0, i_8_28_523_0,
    i_8_28_524_0, i_8_28_525_0, i_8_28_567_0, i_8_28_577_0, i_8_28_595_0,
    i_8_28_596_0, i_8_28_607_0, i_8_28_610_0, i_8_28_631_0, i_8_28_634_0,
    i_8_28_637_0, i_8_28_658_0, i_8_28_667_0, i_8_28_702_0, i_8_28_703_0,
    i_8_28_712_0, i_8_28_748_0, i_8_28_751_0, i_8_28_829_0, i_8_28_838_0,
    i_8_28_844_0, i_8_28_859_0, i_8_28_881_0, i_8_28_910_0, i_8_28_929_0,
    i_8_28_955_0, i_8_28_964_0, i_8_28_967_0, i_8_28_968_0, i_8_28_997_0,
    i_8_28_1179_0, i_8_28_1198_0, i_8_28_1234_0, i_8_28_1252_0,
    i_8_28_1282_0, i_8_28_1354_0, i_8_28_1387_0, i_8_28_1396_0,
    i_8_28_1467_0, i_8_28_1468_0, i_8_28_1486_0, i_8_28_1495_0,
    i_8_28_1507_0, i_8_28_1531_0, i_8_28_1533_0, i_8_28_1536_0,
    i_8_28_1594_0, i_8_28_1629_0, i_8_28_1639_0, i_8_28_1647_0,
    i_8_28_1657_0, i_8_28_1702_0, i_8_28_1703_0, i_8_28_1747_0,
    i_8_28_1757_0, i_8_28_1774_0, i_8_28_1775_0, i_8_28_1791_0,
    i_8_28_1792_0, i_8_28_1801_0, i_8_28_1802_0, i_8_28_1818_0,
    i_8_28_1819_0, i_8_28_1822_0, i_8_28_1846_0, i_8_28_1864_0,
    i_8_28_1873_0, i_8_28_1900_0, i_8_28_1910_0, i_8_28_1963_0,
    i_8_28_2008_0, i_8_28_2044_0, i_8_28_2062_0, i_8_28_2089_0,
    i_8_28_2116_0, i_8_28_2133_0, i_8_28_2134_0, i_8_28_2173_0,
    i_8_28_2227_0, i_8_28_2284_0;
  output o_8_28_0_0;
  assign o_8_28_0_0 = 0;
endmodule



// Benchmark "kernel_8_29" written by ABC on Sun Jul 19 10:03:30 2020

module kernel_8_29 ( 
    i_8_29_58_0, i_8_29_77_0, i_8_29_80_0, i_8_29_104_0, i_8_29_107_0,
    i_8_29_116_0, i_8_29_140_0, i_8_29_182_0, i_8_29_185_0, i_8_29_188_0,
    i_8_29_197_0, i_8_29_247_0, i_8_29_366_0, i_8_29_367_0, i_8_29_389_0,
    i_8_29_391_0, i_8_29_394_0, i_8_29_400_0, i_8_29_401_0, i_8_29_428_0,
    i_8_29_431_0, i_8_29_451_0, i_8_29_453_0, i_8_29_490_0, i_8_29_575_0,
    i_8_29_584_0, i_8_29_594_0, i_8_29_604_0, i_8_29_608_0, i_8_29_610_0,
    i_8_29_638_0, i_8_29_814_0, i_8_29_853_0, i_8_29_856_0, i_8_29_860_0,
    i_8_29_879_0, i_8_29_962_0, i_8_29_1012_0, i_8_29_1013_0,
    i_8_29_1015_0, i_8_29_1016_0, i_8_29_1029_0, i_8_29_1040_0,
    i_8_29_1105_0, i_8_29_1106_0, i_8_29_1129_0, i_8_29_1130_0,
    i_8_29_1142_0, i_8_29_1157_0, i_8_29_1160_0, i_8_29_1228_0,
    i_8_29_1322_0, i_8_29_1328_0, i_8_29_1331_0, i_8_29_1350_0,
    i_8_29_1407_0, i_8_29_1465_0, i_8_29_1493_0, i_8_29_1507_0,
    i_8_29_1510_0, i_8_29_1519_0, i_8_29_1538_0, i_8_29_1550_0,
    i_8_29_1553_0, i_8_29_1658_0, i_8_29_1688_0, i_8_29_1690_0,
    i_8_29_1697_0, i_8_29_1784_0, i_8_29_1817_0, i_8_29_1822_0,
    i_8_29_1838_0, i_8_29_1840_0, i_8_29_1844_0, i_8_29_1850_0,
    i_8_29_1860_0, i_8_29_1882_0, i_8_29_1885_0, i_8_29_1894_0,
    i_8_29_1895_0, i_8_29_1946_0, i_8_29_1966_0, i_8_29_2017_0,
    i_8_29_2038_0, i_8_29_2041_0, i_8_29_2072_0, i_8_29_2116_0,
    i_8_29_2119_0, i_8_29_2120_0, i_8_29_2126_0, i_8_29_2150_0,
    i_8_29_2154_0, i_8_29_2172_0, i_8_29_2177_0, i_8_29_2231_0,
    i_8_29_2263_0, i_8_29_2264_0, i_8_29_2266_0, i_8_29_2273_0,
    i_8_29_2276_0,
    o_8_29_0_0  );
  input  i_8_29_58_0, i_8_29_77_0, i_8_29_80_0, i_8_29_104_0,
    i_8_29_107_0, i_8_29_116_0, i_8_29_140_0, i_8_29_182_0, i_8_29_185_0,
    i_8_29_188_0, i_8_29_197_0, i_8_29_247_0, i_8_29_366_0, i_8_29_367_0,
    i_8_29_389_0, i_8_29_391_0, i_8_29_394_0, i_8_29_400_0, i_8_29_401_0,
    i_8_29_428_0, i_8_29_431_0, i_8_29_451_0, i_8_29_453_0, i_8_29_490_0,
    i_8_29_575_0, i_8_29_584_0, i_8_29_594_0, i_8_29_604_0, i_8_29_608_0,
    i_8_29_610_0, i_8_29_638_0, i_8_29_814_0, i_8_29_853_0, i_8_29_856_0,
    i_8_29_860_0, i_8_29_879_0, i_8_29_962_0, i_8_29_1012_0, i_8_29_1013_0,
    i_8_29_1015_0, i_8_29_1016_0, i_8_29_1029_0, i_8_29_1040_0,
    i_8_29_1105_0, i_8_29_1106_0, i_8_29_1129_0, i_8_29_1130_0,
    i_8_29_1142_0, i_8_29_1157_0, i_8_29_1160_0, i_8_29_1228_0,
    i_8_29_1322_0, i_8_29_1328_0, i_8_29_1331_0, i_8_29_1350_0,
    i_8_29_1407_0, i_8_29_1465_0, i_8_29_1493_0, i_8_29_1507_0,
    i_8_29_1510_0, i_8_29_1519_0, i_8_29_1538_0, i_8_29_1550_0,
    i_8_29_1553_0, i_8_29_1658_0, i_8_29_1688_0, i_8_29_1690_0,
    i_8_29_1697_0, i_8_29_1784_0, i_8_29_1817_0, i_8_29_1822_0,
    i_8_29_1838_0, i_8_29_1840_0, i_8_29_1844_0, i_8_29_1850_0,
    i_8_29_1860_0, i_8_29_1882_0, i_8_29_1885_0, i_8_29_1894_0,
    i_8_29_1895_0, i_8_29_1946_0, i_8_29_1966_0, i_8_29_2017_0,
    i_8_29_2038_0, i_8_29_2041_0, i_8_29_2072_0, i_8_29_2116_0,
    i_8_29_2119_0, i_8_29_2120_0, i_8_29_2126_0, i_8_29_2150_0,
    i_8_29_2154_0, i_8_29_2172_0, i_8_29_2177_0, i_8_29_2231_0,
    i_8_29_2263_0, i_8_29_2264_0, i_8_29_2266_0, i_8_29_2273_0,
    i_8_29_2276_0;
  output o_8_29_0_0;
  assign o_8_29_0_0 = ~((~i_8_29_2126_0 & ((~i_8_29_1040_0 & ((~i_8_29_879_0 & ((~i_8_29_80_0 & ~i_8_29_1894_0 & ((~i_8_29_431_0 & ~i_8_29_490_0 & ~i_8_29_584_0 & ~i_8_29_1510_0 & ~i_8_29_1697_0 & ~i_8_29_2072_0) | (~i_8_29_608_0 & ~i_8_29_1130_0 & ~i_8_29_1322_0 & ~i_8_29_1407_0 & ~i_8_29_1519_0 & ~i_8_29_1688_0 & ~i_8_29_1822_0 & ~i_8_29_1838_0 & ~i_8_29_2273_0))) | (~i_8_29_490_0 & ~i_8_29_584_0 & ~i_8_29_610_0 & ~i_8_29_1016_0 & ~i_8_29_1838_0 & ~i_8_29_2116_0 & ~i_8_29_2120_0 & ~i_8_29_2231_0 & i_8_29_2273_0))) | (~i_8_29_182_0 & ~i_8_29_1015_0 & ~i_8_29_1016_0 & i_8_29_1840_0 & i_8_29_2172_0 & ~i_8_29_2266_0))) | (~i_8_29_182_0 & ((~i_8_29_185_0 & ((i_8_29_107_0 & ~i_8_29_575_0 & ~i_8_29_1507_0 & ~i_8_29_1510_0 & ~i_8_29_1658_0 & ~i_8_29_1840_0) | (~i_8_29_188_0 & ~i_8_29_391_0 & ~i_8_29_401_0 & ~i_8_29_1160_0 & ~i_8_29_1465_0 & ~i_8_29_1688_0 & ~i_8_29_1690_0 & ~i_8_29_1838_0 & ~i_8_29_1894_0 & ~i_8_29_1946_0 & ~i_8_29_2116_0))) | (~i_8_29_188_0 & ~i_8_29_394_0 & i_8_29_490_0 & ~i_8_29_608_0 & ~i_8_29_1129_0 & ~i_8_29_1130_0 & ~i_8_29_1328_0 & ~i_8_29_1407_0 & ~i_8_29_1507_0 & ~i_8_29_1688_0 & ~i_8_29_1838_0) | (~i_8_29_428_0 & ~i_8_29_490_0 & ~i_8_29_610_0 & ~i_8_29_1013_0 & ~i_8_29_1160_0 & ~i_8_29_1322_0 & ~i_8_29_1331_0 & ~i_8_29_1538_0 & ~i_8_29_1822_0 & ~i_8_29_1894_0 & ~i_8_29_2072_0))) | (~i_8_29_584_0 & ((i_8_29_428_0 & ~i_8_29_575_0 & ~i_8_29_608_0 & ~i_8_29_1331_0 & ~i_8_29_1507_0 & ~i_8_29_1688_0 & ~i_8_29_1697_0 & ~i_8_29_1838_0 & ~i_8_29_2041_0) | (i_8_29_1228_0 & ~i_8_29_1690_0 & i_8_29_2116_0 & ~i_8_29_2154_0))) | (i_8_29_58_0 & ~i_8_29_116_0 & ~i_8_29_604_0 & ~i_8_29_1012_0 & ~i_8_29_1013_0 & ~i_8_29_1015_0 & ~i_8_29_1350_0 & ~i_8_29_1465_0 & ~i_8_29_1946_0 & ~i_8_29_2017_0 & ~i_8_29_2273_0))) | (~i_8_29_1013_0 & ((i_8_29_140_0 & ((~i_8_29_247_0 & ~i_8_29_584_0 & ~i_8_29_1350_0 & ~i_8_29_1493_0 & ~i_8_29_1519_0 & i_8_29_1885_0 & ~i_8_29_2154_0) | (~i_8_29_401_0 & ~i_8_29_1105_0 & ~i_8_29_1130_0 & ~i_8_29_1157_0 & ~i_8_29_1507_0 & ~i_8_29_1510_0 & ~i_8_29_1840_0 & ~i_8_29_1894_0 & ~i_8_29_1895_0 & ~i_8_29_2017_0 & ~i_8_29_2231_0))) | (~i_8_29_182_0 & ((~i_8_29_185_0 & ~i_8_29_1331_0 & ~i_8_29_1465_0 & ((~i_8_29_188_0 & ~i_8_29_389_0 & ~i_8_29_610_0 & ~i_8_29_1012_0 & ~i_8_29_1105_0 & ~i_8_29_1130_0 & ~i_8_29_1322_0 & ~i_8_29_1328_0 & ~i_8_29_1350_0 & ~i_8_29_1885_0) | (~i_8_29_400_0 & ~i_8_29_490_0 & ~i_8_29_1157_0 & ~i_8_29_1507_0 & ~i_8_29_1690_0 & ~i_8_29_1838_0 & ~i_8_29_1894_0))) | (~i_8_29_140_0 & ~i_8_29_1040_0 & ~i_8_29_1160_0 & ~i_8_29_1322_0 & ~i_8_29_1510_0 & ~i_8_29_1553_0 & ~i_8_29_1697_0 & ~i_8_29_1822_0 & ~i_8_29_1860_0))) | (i_8_29_1966_0 & ~i_8_29_2273_0 & ((i_8_29_860_0 & i_8_29_1040_0) | (~i_8_29_391_0 & ~i_8_29_610_0 & i_8_29_1840_0 & ~i_8_29_1895_0 & ~i_8_29_2231_0))) | (~i_8_29_428_0 & ~i_8_29_1157_0 & ~i_8_29_1507_0 & i_8_29_1882_0 & ~i_8_29_2017_0 & i_8_29_2116_0 & ~i_8_29_2150_0))) | (~i_8_29_182_0 & ((~i_8_29_116_0 & ~i_8_29_1012_0 & ((~i_8_29_451_0 & ~i_8_29_584_0 & ~i_8_29_1322_0 & ~i_8_29_1331_0 & ~i_8_29_1407_0 & ~i_8_29_1519_0 & ~i_8_29_1538_0 & ~i_8_29_1658_0 & ~i_8_29_1688_0 & ~i_8_29_1840_0 & ~i_8_29_1946_0 & ~i_8_29_2038_0 & ~i_8_29_2116_0) | (~i_8_29_140_0 & ~i_8_29_389_0 & ~i_8_29_1016_0 & ~i_8_29_1350_0 & ~i_8_29_1465_0 & ~i_8_29_1895_0 & i_8_29_1966_0 & ~i_8_29_2017_0 & ~i_8_29_2231_0))) | (~i_8_29_1658_0 & ((~i_8_29_185_0 & ~i_8_29_1844_0 & ~i_8_29_2017_0 & ((i_8_29_490_0 & ~i_8_29_575_0 & ~i_8_29_879_0 & ~i_8_29_1015_0 & ~i_8_29_1040_0 & ~i_8_29_1157_0 & ~i_8_29_1465_0 & ~i_8_29_1507_0 & ~i_8_29_1553_0) | (~i_8_29_389_0 & ~i_8_29_394_0 & ~i_8_29_431_0 & ~i_8_29_853_0 & ~i_8_29_1322_0 & ~i_8_29_1328_0 & ~i_8_29_1550_0 & ~i_8_29_1690_0 & ~i_8_29_1817_0 & ~i_8_29_1838_0 & ~i_8_29_1885_0 & ~i_8_29_1946_0))) | (i_8_29_77_0 & ~i_8_29_1106_0 & ~i_8_29_1322_0 & ~i_8_29_1688_0 & ~i_8_29_1690_0 & ~i_8_29_1838_0 & ~i_8_29_1882_0 & ~i_8_29_1885_0 & ~i_8_29_1895_0 & ~i_8_29_2177_0))) | (~i_8_29_1519_0 & ((~i_8_29_188_0 & ((~i_8_29_400_0 & ~i_8_29_1160_0 & ~i_8_29_1894_0 & ~i_8_29_2072_0 & ~i_8_29_2150_0 & i_8_29_2154_0) | (~i_8_29_1510_0 & ~i_8_29_1553_0 & ~i_8_29_1105_0 & ~i_8_29_1322_0 & ~i_8_29_1688_0 & ~i_8_29_1690_0 & ~i_8_29_1838_0 & ~i_8_29_1840_0 & ~i_8_29_2273_0))) | (i_8_29_366_0 & ~i_8_29_394_0 & ~i_8_29_401_0 & i_8_29_1822_0 & ~i_8_29_1850_0 & i_8_29_1860_0 & ~i_8_29_2041_0))) | (~i_8_29_197_0 & i_8_29_389_0 & ~i_8_29_401_0 & ~i_8_29_962_0 & ~i_8_29_1040_0 & ~i_8_29_1157_0 & ~i_8_29_2276_0))) | (~i_8_29_1838_0 & ((~i_8_29_116_0 & ((i_8_29_366_0 & ~i_8_29_431_0 & ~i_8_29_604_0 & ~i_8_29_1519_0 & ~i_8_29_1688_0 & ~i_8_29_1690_0 & ~i_8_29_1784_0 & ~i_8_29_2017_0) | (~i_8_29_1465_0 & ~i_8_29_1697_0 & ~i_8_29_1894_0 & ~i_8_29_2072_0 & i_8_29_2172_0 & ~i_8_29_2177_0))) | (~i_8_29_185_0 & ~i_8_29_584_0 & ~i_8_29_1016_0 & ~i_8_29_1105_0 & ~i_8_29_1129_0 & ~i_8_29_1331_0 & ~i_8_29_1407_0 & ~i_8_29_1465_0 & ~i_8_29_1519_0 & ~i_8_29_1553_0 & ~i_8_29_1860_0 & ~i_8_29_1946_0 & ~i_8_29_2072_0) | (i_8_29_247_0 & ~i_8_29_394_0 & ~i_8_29_1012_0 & ~i_8_29_1322_0 & ~i_8_29_2273_0))) | (~i_8_29_140_0 & ((~i_8_29_400_0 & ~i_8_29_1106_0 & ~i_8_29_1322_0 & ~i_8_29_1331_0 & ~i_8_29_1519_0 & i_8_29_1817_0) | (~i_8_29_389_0 & ~i_8_29_879_0 & ~i_8_29_1040_0 & ~i_8_29_1105_0 & ~i_8_29_1465_0 & ~i_8_29_1510_0 & ~i_8_29_1688_0 & i_8_29_1885_0 & i_8_29_2041_0))) | (~i_8_29_1322_0 & ((~i_8_29_389_0 & ((~i_8_29_1012_0 & i_8_29_1350_0 & ~i_8_29_1519_0 & ~i_8_29_1895_0 & i_8_29_1946_0 & ~i_8_29_2072_0) | (~i_8_29_185_0 & ~i_8_29_594_0 & ~i_8_29_1129_0 & ~i_8_29_1658_0 & i_8_29_1850_0 & ~i_8_29_1860_0 & ~i_8_29_2116_0))) | (~i_8_29_1129_0 & ~i_8_29_2072_0 & ((~i_8_29_197_0 & ~i_8_29_604_0 & ~i_8_29_1130_0 & ~i_8_29_1142_0 & ~i_8_29_1493_0 & ~i_8_29_1658_0 & ~i_8_29_1895_0 & i_8_29_2041_0) | (~i_8_29_366_0 & ~i_8_29_391_0 & i_8_29_879_0 & ~i_8_29_1553_0 & ~i_8_29_1844_0 & ~i_8_29_2273_0))))) | (~i_8_29_185_0 & ((~i_8_29_1040_0 & i_8_29_1130_0 & ~i_8_29_1822_0 & i_8_29_2038_0 & ~i_8_29_2072_0) | (~i_8_29_107_0 & i_8_29_367_0 & ~i_8_29_391_0 & ~i_8_29_394_0 & ~i_8_29_1130_0 & ~i_8_29_1465_0 & ~i_8_29_1510_0 & ~i_8_29_1538_0 & ~i_8_29_1553_0 & ~i_8_29_1840_0 & ~i_8_29_1946_0 & ~i_8_29_2177_0))) | (~i_8_29_1328_0 & i_8_29_1550_0 & i_8_29_1553_0 & ~i_8_29_1850_0 & ~i_8_29_1895_0 & i_8_29_2038_0) | (~i_8_29_77_0 & ~i_8_29_394_0 & ~i_8_29_575_0 & ~i_8_29_1882_0 & ~i_8_29_1894_0 & ~i_8_29_2116_0 & i_8_29_2119_0));
endmodule



// Benchmark "kernel_8_30" written by ABC on Sun Jul 19 10:03:32 2020

module kernel_8_30 ( 
    i_8_30_32_0, i_8_30_49_0, i_8_30_50_0, i_8_30_87_0, i_8_30_95_0,
    i_8_30_116_0, i_8_30_143_0, i_8_30_167_0, i_8_30_176_0, i_8_30_220_0,
    i_8_30_227_0, i_8_30_304_0, i_8_30_347_0, i_8_30_361_0, i_8_30_378_0,
    i_8_30_383_0, i_8_30_385_0, i_8_30_416_0, i_8_30_425_0, i_8_30_490_0,
    i_8_30_525_0, i_8_30_527_0, i_8_30_550_0, i_8_30_553_0, i_8_30_581_0,
    i_8_30_614_0, i_8_30_653_0, i_8_30_656_0, i_8_30_671_0, i_8_30_677_0,
    i_8_30_687_0, i_8_30_689_0, i_8_30_695_0, i_8_30_749_0, i_8_30_794_0,
    i_8_30_796_0, i_8_30_797_0, i_8_30_806_0, i_8_30_830_0, i_8_30_838_0,
    i_8_30_932_0, i_8_30_956_0, i_8_30_991_0, i_8_30_994_0, i_8_30_1058_0,
    i_8_30_1101_0, i_8_30_1126_0, i_8_30_1127_0, i_8_30_1130_0,
    i_8_30_1175_0, i_8_30_1235_0, i_8_30_1256_0, i_8_30_1271_0,
    i_8_30_1277_0, i_8_30_1283_0, i_8_30_1285_0, i_8_30_1323_0,
    i_8_30_1340_0, i_8_30_1358_0, i_8_30_1382_0, i_8_30_1442_0,
    i_8_30_1453_0, i_8_30_1454_0, i_8_30_1471_0, i_8_30_1481_0,
    i_8_30_1489_0, i_8_30_1490_0, i_8_30_1536_0, i_8_30_1544_0,
    i_8_30_1552_0, i_8_30_1625_0, i_8_30_1639_0, i_8_30_1677_0,
    i_8_30_1697_0, i_8_30_1721_0, i_8_30_1741_0, i_8_30_1774_0,
    i_8_30_1775_0, i_8_30_1801_0, i_8_30_1823_0, i_8_30_1856_0,
    i_8_30_1868_0, i_8_30_1886_0, i_8_30_1889_0, i_8_30_1892_0,
    i_8_30_1943_0, i_8_30_1966_0, i_8_30_1991_0, i_8_30_2039_0,
    i_8_30_2050_0, i_8_30_2143_0, i_8_30_2146_0, i_8_30_2171_0,
    i_8_30_2192_0, i_8_30_2210_0, i_8_30_2215_0, i_8_30_2237_0,
    i_8_30_2261_0, i_8_30_2282_0, i_8_30_2291_0,
    o_8_30_0_0  );
  input  i_8_30_32_0, i_8_30_49_0, i_8_30_50_0, i_8_30_87_0, i_8_30_95_0,
    i_8_30_116_0, i_8_30_143_0, i_8_30_167_0, i_8_30_176_0, i_8_30_220_0,
    i_8_30_227_0, i_8_30_304_0, i_8_30_347_0, i_8_30_361_0, i_8_30_378_0,
    i_8_30_383_0, i_8_30_385_0, i_8_30_416_0, i_8_30_425_0, i_8_30_490_0,
    i_8_30_525_0, i_8_30_527_0, i_8_30_550_0, i_8_30_553_0, i_8_30_581_0,
    i_8_30_614_0, i_8_30_653_0, i_8_30_656_0, i_8_30_671_0, i_8_30_677_0,
    i_8_30_687_0, i_8_30_689_0, i_8_30_695_0, i_8_30_749_0, i_8_30_794_0,
    i_8_30_796_0, i_8_30_797_0, i_8_30_806_0, i_8_30_830_0, i_8_30_838_0,
    i_8_30_932_0, i_8_30_956_0, i_8_30_991_0, i_8_30_994_0, i_8_30_1058_0,
    i_8_30_1101_0, i_8_30_1126_0, i_8_30_1127_0, i_8_30_1130_0,
    i_8_30_1175_0, i_8_30_1235_0, i_8_30_1256_0, i_8_30_1271_0,
    i_8_30_1277_0, i_8_30_1283_0, i_8_30_1285_0, i_8_30_1323_0,
    i_8_30_1340_0, i_8_30_1358_0, i_8_30_1382_0, i_8_30_1442_0,
    i_8_30_1453_0, i_8_30_1454_0, i_8_30_1471_0, i_8_30_1481_0,
    i_8_30_1489_0, i_8_30_1490_0, i_8_30_1536_0, i_8_30_1544_0,
    i_8_30_1552_0, i_8_30_1625_0, i_8_30_1639_0, i_8_30_1677_0,
    i_8_30_1697_0, i_8_30_1721_0, i_8_30_1741_0, i_8_30_1774_0,
    i_8_30_1775_0, i_8_30_1801_0, i_8_30_1823_0, i_8_30_1856_0,
    i_8_30_1868_0, i_8_30_1886_0, i_8_30_1889_0, i_8_30_1892_0,
    i_8_30_1943_0, i_8_30_1966_0, i_8_30_1991_0, i_8_30_2039_0,
    i_8_30_2050_0, i_8_30_2143_0, i_8_30_2146_0, i_8_30_2171_0,
    i_8_30_2192_0, i_8_30_2210_0, i_8_30_2215_0, i_8_30_2237_0,
    i_8_30_2261_0, i_8_30_2282_0, i_8_30_2291_0;
  output o_8_30_0_0;
  assign o_8_30_0_0 = ~((~i_8_30_794_0 & ((~i_8_30_32_0 & ((~i_8_30_383_0 & ~i_8_30_677_0 & ~i_8_30_1175_0 & ~i_8_30_1256_0 & ~i_8_30_1856_0 & ~i_8_30_2146_0 & ~i_8_30_2210_0) | (~i_8_30_87_0 & i_8_30_304_0 & ~i_8_30_689_0 & ~i_8_30_994_0 & ~i_8_30_1471_0 & ~i_8_30_1625_0 & ~i_8_30_2237_0 & ~i_8_30_2282_0))) | (~i_8_30_1256_0 & ((~i_8_30_1453_0 & ((~i_8_30_50_0 & ((~i_8_30_383_0 & ~i_8_30_689_0) | (~i_8_30_830_0 & ~i_8_30_932_0 & ~i_8_30_1130_0 & ~i_8_30_1868_0 & ~i_8_30_1943_0 & ~i_8_30_2192_0))) | (~i_8_30_830_0 & ~i_8_30_932_0 & ~i_8_30_1277_0 & ~i_8_30_1856_0 & ~i_8_30_1868_0 & ~i_8_30_2192_0 & ~i_8_30_2291_0))) | (~i_8_30_167_0 & i_8_30_1058_0 & ~i_8_30_2261_0))))) | (~i_8_30_385_0 & ((~i_8_30_143_0 & ~i_8_30_689_0 & ~i_8_30_1271_0 & i_8_30_1358_0 & ~i_8_30_1382_0 & ~i_8_30_1544_0 & ~i_8_30_2215_0) | (~i_8_30_49_0 & ~i_8_30_347_0 & ~i_8_30_656_0 & ~i_8_30_806_0 & ~i_8_30_932_0 & ~i_8_30_956_0 & ~i_8_30_1058_0 & ~i_8_30_1625_0 & ~i_8_30_2192_0 & ~i_8_30_2282_0))) | (~i_8_30_581_0 & ((i_8_30_383_0 & ~i_8_30_671_0 & ~i_8_30_695_0 & ~i_8_30_1256_0 & ~i_8_30_1552_0 & ~i_8_30_2039_0) | (~i_8_30_830_0 & ~i_8_30_994_0 & ~i_8_30_1454_0 & ~i_8_30_1868_0 & i_8_30_2146_0 & ~i_8_30_2282_0))) | (~i_8_30_2192_0 & ((~i_8_30_614_0 & ~i_8_30_1889_0 & ((~i_8_30_1058_0 & i_8_30_1283_0 & ~i_8_30_1442_0 & ~i_8_30_1454_0 & ~i_8_30_1856_0 & ~i_8_30_1868_0 & ~i_8_30_2039_0) | (i_8_30_347_0 & ~i_8_30_838_0 & ~i_8_30_1552_0 & ~i_8_30_1625_0 & ~i_8_30_2237_0))) | (~i_8_30_176_0 & i_8_30_385_0 & ~i_8_30_677_0 & ~i_8_30_932_0 & ~i_8_30_1058_0 & ~i_8_30_1442_0 & ~i_8_30_1453_0 & ~i_8_30_2210_0) | (~i_8_30_167_0 & ~i_8_30_361_0 & i_8_30_838_0 & ~i_8_30_1454_0 & ~i_8_30_2215_0 & ~i_8_30_2261_0 & ~i_8_30_2282_0))) | (~i_8_30_167_0 & ((~i_8_30_796_0 & i_8_30_1490_0 & i_8_30_1552_0 & i_8_30_1801_0) | (~i_8_30_304_0 & ~i_8_30_687_0 & ~i_8_30_689_0 & ~i_8_30_1235_0 & ~i_8_30_1283_0 & ~i_8_30_2291_0))) | (~i_8_30_671_0 & ((~i_8_30_116_0 & ~i_8_30_490_0 & ~i_8_30_797_0 & ~i_8_30_932_0 & ~i_8_30_1175_0 & ~i_8_30_1625_0) | (~i_8_30_95_0 & ~i_8_30_1382_0 & ~i_8_30_1697_0 & i_8_30_1801_0 & ~i_8_30_2210_0 & ~i_8_30_2215_0))) | (~i_8_30_116_0 & ((~i_8_30_50_0 & ~i_8_30_838_0 & ~i_8_30_1235_0 & ~i_8_30_1489_0 & ~i_8_30_1544_0 & ~i_8_30_1625_0 & ~i_8_30_1966_0 & ~i_8_30_2050_0) | (i_8_30_220_0 & ~i_8_30_656_0 & ~i_8_30_806_0 & ~i_8_30_1130_0 & ~i_8_30_2210_0 & ~i_8_30_2261_0))) | (~i_8_30_1256_0 & (i_8_30_1774_0 | (~i_8_30_797_0 & ~i_8_30_1283_0 & ~i_8_30_1544_0 & ~i_8_30_2261_0))) | (i_8_30_677_0 & i_8_30_1126_0) | (~i_8_30_677_0 & ~i_8_30_1271_0 & i_8_30_1677_0 & ~i_8_30_1697_0 & ~i_8_30_1774_0 & ~i_8_30_2261_0) | (~i_8_30_796_0 & ~i_8_30_1175_0 & ~i_8_30_1235_0 & i_8_30_1489_0 & ~i_8_30_1856_0));
endmodule



// Benchmark "kernel_8_31" written by ABC on Sun Jul 19 10:03:33 2020

module kernel_8_31 ( 
    i_8_31_10_0, i_8_31_37_0, i_8_31_73_0, i_8_31_114_0, i_8_31_169_0,
    i_8_31_172_0, i_8_31_363_0, i_8_31_364_0, i_8_31_373_0, i_8_31_442_0,
    i_8_31_454_0, i_8_31_471_0, i_8_31_486_0, i_8_31_487_0, i_8_31_493_0,
    i_8_31_507_0, i_8_31_522_0, i_8_31_526_0, i_8_31_535_0, i_8_31_555_0,
    i_8_31_580_0, i_8_31_616_0, i_8_31_656_0, i_8_31_664_0, i_8_31_669_0,
    i_8_31_684_0, i_8_31_694_0, i_8_31_696_0, i_8_31_697_0, i_8_31_704_0,
    i_8_31_766_0, i_8_31_837_0, i_8_31_840_0, i_8_31_841_0, i_8_31_847_0,
    i_8_31_913_0, i_8_31_948_0, i_8_31_949_0, i_8_31_955_0, i_8_31_956_0,
    i_8_31_1102_0, i_8_31_1103_0, i_8_31_1108_0, i_8_31_1110_0,
    i_8_31_1127_0, i_8_31_1129_0, i_8_31_1130_0, i_8_31_1224_0,
    i_8_31_1225_0, i_8_31_1227_0, i_8_31_1228_0, i_8_31_1281_0,
    i_8_31_1286_0, i_8_31_1305_0, i_8_31_1352_0, i_8_31_1357_0,
    i_8_31_1369_0, i_8_31_1390_0, i_8_31_1399_0, i_8_31_1456_0,
    i_8_31_1480_0, i_8_31_1489_0, i_8_31_1497_0, i_8_31_1516_0,
    i_8_31_1533_0, i_8_31_1549_0, i_8_31_1558_0, i_8_31_1673_0,
    i_8_31_1685_0, i_8_31_1704_0, i_8_31_1784_0, i_8_31_1794_0,
    i_8_31_1803_0, i_8_31_1805_0, i_8_31_1822_0, i_8_31_1824_0,
    i_8_31_1864_0, i_8_31_1885_0, i_8_31_1912_0, i_8_31_1917_0,
    i_8_31_1939_0, i_8_31_1957_0, i_8_31_1990_0, i_8_31_1993_0,
    i_8_31_2006_0, i_8_31_2021_0, i_8_31_2048_0, i_8_31_2133_0,
    i_8_31_2134_0, i_8_31_2143_0, i_8_31_2146_0, i_8_31_2147_0,
    i_8_31_2148_0, i_8_31_2165_0, i_8_31_2215_0, i_8_31_2232_0,
    i_8_31_2236_0, i_8_31_2242_0, i_8_31_2296_0, i_8_31_2299_0,
    o_8_31_0_0  );
  input  i_8_31_10_0, i_8_31_37_0, i_8_31_73_0, i_8_31_114_0,
    i_8_31_169_0, i_8_31_172_0, i_8_31_363_0, i_8_31_364_0, i_8_31_373_0,
    i_8_31_442_0, i_8_31_454_0, i_8_31_471_0, i_8_31_486_0, i_8_31_487_0,
    i_8_31_493_0, i_8_31_507_0, i_8_31_522_0, i_8_31_526_0, i_8_31_535_0,
    i_8_31_555_0, i_8_31_580_0, i_8_31_616_0, i_8_31_656_0, i_8_31_664_0,
    i_8_31_669_0, i_8_31_684_0, i_8_31_694_0, i_8_31_696_0, i_8_31_697_0,
    i_8_31_704_0, i_8_31_766_0, i_8_31_837_0, i_8_31_840_0, i_8_31_841_0,
    i_8_31_847_0, i_8_31_913_0, i_8_31_948_0, i_8_31_949_0, i_8_31_955_0,
    i_8_31_956_0, i_8_31_1102_0, i_8_31_1103_0, i_8_31_1108_0,
    i_8_31_1110_0, i_8_31_1127_0, i_8_31_1129_0, i_8_31_1130_0,
    i_8_31_1224_0, i_8_31_1225_0, i_8_31_1227_0, i_8_31_1228_0,
    i_8_31_1281_0, i_8_31_1286_0, i_8_31_1305_0, i_8_31_1352_0,
    i_8_31_1357_0, i_8_31_1369_0, i_8_31_1390_0, i_8_31_1399_0,
    i_8_31_1456_0, i_8_31_1480_0, i_8_31_1489_0, i_8_31_1497_0,
    i_8_31_1516_0, i_8_31_1533_0, i_8_31_1549_0, i_8_31_1558_0,
    i_8_31_1673_0, i_8_31_1685_0, i_8_31_1704_0, i_8_31_1784_0,
    i_8_31_1794_0, i_8_31_1803_0, i_8_31_1805_0, i_8_31_1822_0,
    i_8_31_1824_0, i_8_31_1864_0, i_8_31_1885_0, i_8_31_1912_0,
    i_8_31_1917_0, i_8_31_1939_0, i_8_31_1957_0, i_8_31_1990_0,
    i_8_31_1993_0, i_8_31_2006_0, i_8_31_2021_0, i_8_31_2048_0,
    i_8_31_2133_0, i_8_31_2134_0, i_8_31_2143_0, i_8_31_2146_0,
    i_8_31_2147_0, i_8_31_2148_0, i_8_31_2165_0, i_8_31_2215_0,
    i_8_31_2232_0, i_8_31_2236_0, i_8_31_2242_0, i_8_31_2296_0,
    i_8_31_2299_0;
  output o_8_31_0_0;
  assign o_8_31_0_0 = 0;
endmodule



// Benchmark "kernel_8_32" written by ABC on Sun Jul 19 10:03:34 2020

module kernel_8_32 ( 
    i_8_32_22_0, i_8_32_39_0, i_8_32_196_0, i_8_32_232_0, i_8_32_300_0,
    i_8_32_303_0, i_8_32_304_0, i_8_32_330_0, i_8_32_360_0, i_8_32_364_0,
    i_8_32_365_0, i_8_32_367_0, i_8_32_368_0, i_8_32_420_0, i_8_32_421_0,
    i_8_32_448_0, i_8_32_457_0, i_8_32_510_0, i_8_32_511_0, i_8_32_520_0,
    i_8_32_525_0, i_8_32_528_0, i_8_32_605_0, i_8_32_606_0, i_8_32_658_0,
    i_8_32_660_0, i_8_32_700_0, i_8_32_751_0, i_8_32_762_0, i_8_32_781_0,
    i_8_32_782_0, i_8_32_795_0, i_8_32_823_0, i_8_32_835_0, i_8_32_842_0,
    i_8_32_843_0, i_8_32_852_0, i_8_32_996_0, i_8_32_997_0, i_8_32_1028_0,
    i_8_32_1050_0, i_8_32_1158_0, i_8_32_1159_0, i_8_32_1192_0,
    i_8_32_1249_0, i_8_32_1274_0, i_8_32_1282_0, i_8_32_1305_0,
    i_8_32_1308_0, i_8_32_1330_0, i_8_32_1382_0, i_8_32_1389_0,
    i_8_32_1391_0, i_8_32_1393_0, i_8_32_1432_0, i_8_32_1437_0,
    i_8_32_1438_0, i_8_32_1439_0, i_8_32_1545_0, i_8_32_1546_0,
    i_8_32_1554_0, i_8_32_1596_0, i_8_32_1635_0, i_8_32_1643_0,
    i_8_32_1679_0, i_8_32_1699_0, i_8_32_1700_0, i_8_32_1708_0,
    i_8_32_1764_0, i_8_32_1784_0, i_8_32_1818_0, i_8_32_1820_0,
    i_8_32_1840_0, i_8_32_1858_0, i_8_32_1875_0, i_8_32_1876_0,
    i_8_32_1879_0, i_8_32_1880_0, i_8_32_1887_0, i_8_32_2013_0,
    i_8_32_2014_0, i_8_32_2075_0, i_8_32_2077_0, i_8_32_2091_0,
    i_8_32_2092_0, i_8_32_2093_0, i_8_32_2095_0, i_8_32_2096_0,
    i_8_32_2122_0, i_8_32_2147_0, i_8_32_2154_0, i_8_32_2214_0,
    i_8_32_2215_0, i_8_32_2216_0, i_8_32_2218_0, i_8_32_2235_0,
    i_8_32_2236_0, i_8_32_2239_0, i_8_32_2244_0, i_8_32_2293_0,
    o_8_32_0_0  );
  input  i_8_32_22_0, i_8_32_39_0, i_8_32_196_0, i_8_32_232_0,
    i_8_32_300_0, i_8_32_303_0, i_8_32_304_0, i_8_32_330_0, i_8_32_360_0,
    i_8_32_364_0, i_8_32_365_0, i_8_32_367_0, i_8_32_368_0, i_8_32_420_0,
    i_8_32_421_0, i_8_32_448_0, i_8_32_457_0, i_8_32_510_0, i_8_32_511_0,
    i_8_32_520_0, i_8_32_525_0, i_8_32_528_0, i_8_32_605_0, i_8_32_606_0,
    i_8_32_658_0, i_8_32_660_0, i_8_32_700_0, i_8_32_751_0, i_8_32_762_0,
    i_8_32_781_0, i_8_32_782_0, i_8_32_795_0, i_8_32_823_0, i_8_32_835_0,
    i_8_32_842_0, i_8_32_843_0, i_8_32_852_0, i_8_32_996_0, i_8_32_997_0,
    i_8_32_1028_0, i_8_32_1050_0, i_8_32_1158_0, i_8_32_1159_0,
    i_8_32_1192_0, i_8_32_1249_0, i_8_32_1274_0, i_8_32_1282_0,
    i_8_32_1305_0, i_8_32_1308_0, i_8_32_1330_0, i_8_32_1382_0,
    i_8_32_1389_0, i_8_32_1391_0, i_8_32_1393_0, i_8_32_1432_0,
    i_8_32_1437_0, i_8_32_1438_0, i_8_32_1439_0, i_8_32_1545_0,
    i_8_32_1546_0, i_8_32_1554_0, i_8_32_1596_0, i_8_32_1635_0,
    i_8_32_1643_0, i_8_32_1679_0, i_8_32_1699_0, i_8_32_1700_0,
    i_8_32_1708_0, i_8_32_1764_0, i_8_32_1784_0, i_8_32_1818_0,
    i_8_32_1820_0, i_8_32_1840_0, i_8_32_1858_0, i_8_32_1875_0,
    i_8_32_1876_0, i_8_32_1879_0, i_8_32_1880_0, i_8_32_1887_0,
    i_8_32_2013_0, i_8_32_2014_0, i_8_32_2075_0, i_8_32_2077_0,
    i_8_32_2091_0, i_8_32_2092_0, i_8_32_2093_0, i_8_32_2095_0,
    i_8_32_2096_0, i_8_32_2122_0, i_8_32_2147_0, i_8_32_2154_0,
    i_8_32_2214_0, i_8_32_2215_0, i_8_32_2216_0, i_8_32_2218_0,
    i_8_32_2235_0, i_8_32_2236_0, i_8_32_2239_0, i_8_32_2244_0,
    i_8_32_2293_0;
  output o_8_32_0_0;
  assign o_8_32_0_0 = ~((~i_8_32_996_0 & ((i_8_32_365_0 & ~i_8_32_2215_0 & ((~i_8_32_421_0 & ~i_8_32_1159_0 & ~i_8_32_1875_0 & ~i_8_32_2014_0 & ~i_8_32_2095_0 & ~i_8_32_2218_0) | (~i_8_32_448_0 & ~i_8_32_511_0 & ~i_8_32_782_0 & ~i_8_32_1554_0 & ~i_8_32_2077_0 & ~i_8_32_2239_0))) | (~i_8_32_1876_0 & ((~i_8_32_520_0 & ~i_8_32_1393_0 & ((i_8_32_762_0 & ~i_8_32_852_0 & ~i_8_32_1432_0 & ~i_8_32_2214_0) | (~i_8_32_457_0 & ~i_8_32_525_0 & ~i_8_32_1308_0 & ~i_8_32_1382_0 & ~i_8_32_1546_0 & ~i_8_32_1708_0 & ~i_8_32_1820_0 & ~i_8_32_1880_0 & ~i_8_32_2096_0 & ~i_8_32_2216_0))) | (i_8_32_367_0 & ~i_8_32_525_0 & ~i_8_32_997_0 & ~i_8_32_1820_0 & ~i_8_32_1879_0 & ~i_8_32_1880_0 & ~i_8_32_2239_0))))) | (~i_8_32_2014_0 & ((~i_8_32_1880_0 & ((~i_8_32_420_0 & ((~i_8_32_196_0 & ~i_8_32_232_0 & ~i_8_32_421_0 & ~i_8_32_1192_0 & ~i_8_32_1282_0 & ~i_8_32_1330_0 & ~i_8_32_1391_0 & ~i_8_32_1784_0 & ~i_8_32_1820_0 & ~i_8_32_2013_0 & ~i_8_32_2092_0) | (~i_8_32_22_0 & i_8_32_700_0 & ~i_8_32_1050_0 & ~i_8_32_1274_0 & ~i_8_32_2239_0))) | (~i_8_32_421_0 & ~i_8_32_525_0 & ~i_8_32_528_0 & ~i_8_32_1274_0 & ~i_8_32_1820_0 & ~i_8_32_1876_0 & i_8_32_2092_0 & ~i_8_32_2239_0) | (~i_8_32_1393_0 & ~i_8_32_1596_0 & i_8_32_1679_0 & ~i_8_32_1879_0 & ~i_8_32_1887_0 & ~i_8_32_2236_0))) | (~i_8_32_2013_0 & ((~i_8_32_762_0 & ((~i_8_32_510_0 & ~i_8_32_511_0 & ~i_8_32_1546_0 & ~i_8_32_1784_0 & i_8_32_1818_0) | (~i_8_32_528_0 & i_8_32_606_0 & ~i_8_32_1840_0 & ~i_8_32_1875_0 & ~i_8_32_2077_0))) | (i_8_32_510_0 & ~i_8_32_520_0 & i_8_32_852_0 & ~i_8_32_1545_0 & ~i_8_32_1875_0 & ~i_8_32_1879_0 & ~i_8_32_2236_0))) | (i_8_32_700_0 & ~i_8_32_1635_0 & ~i_8_32_2091_0 & ~i_8_32_2096_0 & ~i_8_32_2122_0 & ~i_8_32_2147_0 & ~i_8_32_2235_0))) | (~i_8_32_520_0 & ((~i_8_32_22_0 & ~i_8_32_1389_0 & ~i_8_32_1545_0 & ((~i_8_32_420_0 & ~i_8_32_421_0 & ~i_8_32_510_0 & ~i_8_32_751_0 & ~i_8_32_762_0 & ~i_8_32_1391_0 & ~i_8_32_1700_0 & ~i_8_32_1708_0 & ~i_8_32_1879_0 & ~i_8_32_1880_0 & ~i_8_32_2091_0 & ~i_8_32_2154_0) | (i_8_32_525_0 & ~i_8_32_528_0 & ~i_8_32_1784_0 & ~i_8_32_1875_0 & ~i_8_32_2096_0 & ~i_8_32_2215_0))) | (~i_8_32_232_0 & i_8_32_511_0 & ~i_8_32_835_0 & ~i_8_32_852_0 & ~i_8_32_1050_0 & ~i_8_32_1393_0 & ~i_8_32_1643_0 & ~i_8_32_1879_0 & ~i_8_32_2013_0 & ~i_8_32_2214_0 & ~i_8_32_2236_0 & ~i_8_32_2239_0))) | (~i_8_32_1391_0 & ((~i_8_32_196_0 & ~i_8_32_1546_0 & ((~i_8_32_368_0 & ~i_8_32_420_0 & ~i_8_32_1389_0 & ~i_8_32_1545_0 & ~i_8_32_1708_0 & ~i_8_32_1875_0 & ~i_8_32_2095_0 & ~i_8_32_2096_0 & ~i_8_32_2122_0 & i_8_32_2218_0) | (i_8_32_367_0 & ~i_8_32_448_0 & ~i_8_32_457_0 & ~i_8_32_2013_0 & i_8_32_2092_0 & ~i_8_32_2214_0 & ~i_8_32_2239_0))) | (~i_8_32_1880_0 & ((~i_8_32_421_0 & ~i_8_32_835_0 & i_8_32_1439_0 & ~i_8_32_2013_0) | (~i_8_32_511_0 & ~i_8_32_1274_0 & ~i_8_32_1308_0 & ~i_8_32_1596_0 & ~i_8_32_1820_0 & ~i_8_32_1875_0 & ~i_8_32_2091_0 & ~i_8_32_2095_0 & ~i_8_32_2096_0 & ~i_8_32_2122_0 & ~i_8_32_2293_0))) | (~i_8_32_232_0 & ~i_8_32_367_0 & ~i_8_32_420_0 & ~i_8_32_782_0 & ~i_8_32_1393_0 & ~i_8_32_1635_0 & ~i_8_32_2013_0 & ~i_8_32_2092_0 & ~i_8_32_2093_0 & ~i_8_32_2218_0 & ~i_8_32_2235_0 & ~i_8_32_2239_0))) | (~i_8_32_2236_0 & ((~i_8_32_420_0 & ((i_8_32_303_0 & ~i_8_32_852_0 & ~i_8_32_1393_0 & ~i_8_32_1880_0 & ~i_8_32_1887_0) | (~i_8_32_232_0 & ~i_8_32_510_0 & ~i_8_32_1192_0 & i_8_32_1437_0 & ~i_8_32_1643_0 & ~i_8_32_1708_0 & ~i_8_32_2013_0))) | (~i_8_32_1700_0 & i_8_32_1820_0 & ~i_8_32_1876_0 & ~i_8_32_2092_0 & ~i_8_32_2239_0))) | (~i_8_32_232_0 & ((i_8_32_368_0 & i_8_32_842_0 & ~i_8_32_997_0 & ~i_8_32_1876_0 & ~i_8_32_2095_0) | (~i_8_32_330_0 & ~i_8_32_510_0 & ~i_8_32_511_0 & ~i_8_32_852_0 & ~i_8_32_1028_0 & ~i_8_32_1875_0 & ~i_8_32_2122_0 & i_8_32_2293_0))) | (~i_8_32_751_0 & ((~i_8_32_510_0 & ~i_8_32_1050_0 & ~i_8_32_1282_0 & ~i_8_32_1546_0 & ~i_8_32_1596_0 & ~i_8_32_1643_0 & ~i_8_32_1764_0 & ~i_8_32_1875_0 & ~i_8_32_1879_0 & ~i_8_32_2092_0 & ~i_8_32_2096_0) | (~i_8_32_605_0 & ~i_8_32_762_0 & i_8_32_842_0 & ~i_8_32_1382_0 & ~i_8_32_1820_0 & ~i_8_32_2013_0 & ~i_8_32_2147_0 & ~i_8_32_2216_0 & ~i_8_32_2218_0))) | (~i_8_32_852_0 & ((~i_8_32_762_0 & ~i_8_32_1635_0 & ~i_8_32_1708_0 & ~i_8_32_1764_0 & ~i_8_32_1875_0 & ~i_8_32_1879_0 & ~i_8_32_2122_0 & i_8_32_2154_0 & ~i_8_32_2214_0) | (i_8_32_364_0 & ~i_8_32_843_0 & ~i_8_32_1818_0 & ~i_8_32_1876_0 & ~i_8_32_1880_0 & ~i_8_32_2235_0 & ~i_8_32_2244_0))) | (i_8_32_781_0 & i_8_32_1439_0 & ~i_8_32_1879_0 & ~i_8_32_2093_0 & ~i_8_32_2235_0) | (~i_8_32_1305_0 & ~i_8_32_1596_0 & ~i_8_32_1643_0 & ~i_8_32_2013_0 & ~i_8_32_2092_0 & ~i_8_32_2095_0 & ~i_8_32_2096_0 & ~i_8_32_2215_0 & ~i_8_32_2218_0) | (i_8_32_1159_0 & i_8_32_2122_0 & i_8_32_2293_0));
endmodule



// Benchmark "kernel_8_33" written by ABC on Sun Jul 19 10:03:36 2020

module kernel_8_33 ( 
    i_8_33_30_0, i_8_33_33_0, i_8_33_34_0, i_8_33_48_0, i_8_33_49_0,
    i_8_33_53_0, i_8_33_76_0, i_8_33_164_0, i_8_33_174_0, i_8_33_193_0,
    i_8_33_227_0, i_8_33_258_0, i_8_33_305_0, i_8_33_345_0, i_8_33_348_0,
    i_8_33_366_0, i_8_33_385_0, i_8_33_453_0, i_8_33_479_0, i_8_33_510_0,
    i_8_33_552_0, i_8_33_585_0, i_8_33_634_0, i_8_33_651_0, i_8_33_652_0,
    i_8_33_653_0, i_8_33_718_0, i_8_33_719_0, i_8_33_770_0, i_8_33_773_0,
    i_8_33_778_0, i_8_33_796_0, i_8_33_797_0, i_8_33_805_0, i_8_33_862_0,
    i_8_33_885_0, i_8_33_890_0, i_8_33_921_0, i_8_33_923_0, i_8_33_930_0,
    i_8_33_935_0, i_8_33_992_0, i_8_33_1091_0, i_8_33_1102_0,
    i_8_33_1159_0, i_8_33_1170_0, i_8_33_1258_0, i_8_33_1259_0,
    i_8_33_1263_0, i_8_33_1265_0, i_8_33_1274_0, i_8_33_1301_0,
    i_8_33_1302_0, i_8_33_1305_0, i_8_33_1330_0, i_8_33_1331_0,
    i_8_33_1355_0, i_8_33_1399_0, i_8_33_1408_0, i_8_33_1470_0,
    i_8_33_1471_0, i_8_33_1473_0, i_8_33_1489_0, i_8_33_1490_0,
    i_8_33_1549_0, i_8_33_1562_0, i_8_33_1587_0, i_8_33_1678_0,
    i_8_33_1700_0, i_8_33_1733_0, i_8_33_1753_0, i_8_33_1773_0,
    i_8_33_1774_0, i_8_33_1776_0, i_8_33_1778_0, i_8_33_1788_0,
    i_8_33_1805_0, i_8_33_1864_0, i_8_33_1939_0, i_8_33_1993_0,
    i_8_33_2017_0, i_8_33_2031_0, i_8_33_2048_0, i_8_33_2111_0,
    i_8_33_2172_0, i_8_33_2174_0, i_8_33_2175_0, i_8_33_2176_0,
    i_8_33_2177_0, i_8_33_2194_0, i_8_33_2200_0, i_8_33_2206_0,
    i_8_33_2244_0, i_8_33_2245_0, i_8_33_2246_0, i_8_33_2249_0,
    i_8_33_2264_0, i_8_33_2276_0, i_8_33_2291_0, i_8_33_2292_0,
    o_8_33_0_0  );
  input  i_8_33_30_0, i_8_33_33_0, i_8_33_34_0, i_8_33_48_0, i_8_33_49_0,
    i_8_33_53_0, i_8_33_76_0, i_8_33_164_0, i_8_33_174_0, i_8_33_193_0,
    i_8_33_227_0, i_8_33_258_0, i_8_33_305_0, i_8_33_345_0, i_8_33_348_0,
    i_8_33_366_0, i_8_33_385_0, i_8_33_453_0, i_8_33_479_0, i_8_33_510_0,
    i_8_33_552_0, i_8_33_585_0, i_8_33_634_0, i_8_33_651_0, i_8_33_652_0,
    i_8_33_653_0, i_8_33_718_0, i_8_33_719_0, i_8_33_770_0, i_8_33_773_0,
    i_8_33_778_0, i_8_33_796_0, i_8_33_797_0, i_8_33_805_0, i_8_33_862_0,
    i_8_33_885_0, i_8_33_890_0, i_8_33_921_0, i_8_33_923_0, i_8_33_930_0,
    i_8_33_935_0, i_8_33_992_0, i_8_33_1091_0, i_8_33_1102_0,
    i_8_33_1159_0, i_8_33_1170_0, i_8_33_1258_0, i_8_33_1259_0,
    i_8_33_1263_0, i_8_33_1265_0, i_8_33_1274_0, i_8_33_1301_0,
    i_8_33_1302_0, i_8_33_1305_0, i_8_33_1330_0, i_8_33_1331_0,
    i_8_33_1355_0, i_8_33_1399_0, i_8_33_1408_0, i_8_33_1470_0,
    i_8_33_1471_0, i_8_33_1473_0, i_8_33_1489_0, i_8_33_1490_0,
    i_8_33_1549_0, i_8_33_1562_0, i_8_33_1587_0, i_8_33_1678_0,
    i_8_33_1700_0, i_8_33_1733_0, i_8_33_1753_0, i_8_33_1773_0,
    i_8_33_1774_0, i_8_33_1776_0, i_8_33_1778_0, i_8_33_1788_0,
    i_8_33_1805_0, i_8_33_1864_0, i_8_33_1939_0, i_8_33_1993_0,
    i_8_33_2017_0, i_8_33_2031_0, i_8_33_2048_0, i_8_33_2111_0,
    i_8_33_2172_0, i_8_33_2174_0, i_8_33_2175_0, i_8_33_2176_0,
    i_8_33_2177_0, i_8_33_2194_0, i_8_33_2200_0, i_8_33_2206_0,
    i_8_33_2244_0, i_8_33_2245_0, i_8_33_2246_0, i_8_33_2249_0,
    i_8_33_2264_0, i_8_33_2276_0, i_8_33_2291_0, i_8_33_2292_0;
  output o_8_33_0_0;
  assign o_8_33_0_0 = ~((~i_8_33_770_0 & ((~i_8_33_773_0 & ((~i_8_33_34_0 & ((~i_8_33_49_0 & i_8_33_1355_0 & ~i_8_33_2031_0 & i_8_33_2174_0 & ~i_8_33_2194_0) | (~i_8_33_164_0 & ~i_8_33_890_0 & ~i_8_33_921_0 & ~i_8_33_1170_0 & ~i_8_33_1258_0 & ~i_8_33_1259_0 & i_8_33_1265_0 & ~i_8_33_1331_0 & ~i_8_33_1549_0 & ~i_8_33_1864_0 & ~i_8_33_2200_0 & ~i_8_33_2206_0 & ~i_8_33_2264_0 & ~i_8_33_2291_0))) | (~i_8_33_453_0 & ~i_8_33_797_0 & ((~i_8_33_1170_0 & ~i_8_33_1258_0 & ~i_8_33_479_0 & ~i_8_33_719_0 & ~i_8_33_1259_0 & ~i_8_33_1274_0 & ~i_8_33_2031_0 & ~i_8_33_2194_0 & i_8_33_2246_0) | (~i_8_33_796_0 & ~i_8_33_923_0 & ~i_8_33_992_0 & ~i_8_33_1159_0 & ~i_8_33_1470_0 & ~i_8_33_1549_0 & i_8_33_1778_0 & ~i_8_33_1939_0 & ~i_8_33_1993_0 & ~i_8_33_2200_0 & ~i_8_33_2291_0 & ~i_8_33_2292_0))) | (~i_8_33_49_0 & i_8_33_193_0 & ~i_8_33_510_0 & ~i_8_33_805_0 & ~i_8_33_1259_0 & ~i_8_33_1302_0 & ~i_8_33_1408_0 & ~i_8_33_2017_0 & ~i_8_33_2177_0))) | (~i_8_33_53_0 & ((~i_8_33_48_0 & ~i_8_33_1259_0 & ((~i_8_33_164_0 & ~i_8_33_258_0 & ~i_8_33_348_0 & ~i_8_33_453_0 & ~i_8_33_1159_0 & ~i_8_33_1473_0 & i_8_33_2172_0 & ~i_8_33_2206_0) | (~i_8_33_49_0 & ~i_8_33_345_0 & ~i_8_33_796_0 & ~i_8_33_1091_0 & ~i_8_33_1471_0 & ~i_8_33_1549_0 & ~i_8_33_2111_0 & i_8_33_2177_0 & ~i_8_33_2264_0))) | (~i_8_33_1258_0 & i_8_33_1490_0 & ~i_8_33_1753_0 & i_8_33_2174_0 & ~i_8_33_2291_0))) | (~i_8_33_164_0 & ((~i_8_33_76_0 & ~i_8_33_227_0 & ~i_8_33_1091_0 & ~i_8_33_1305_0 & i_8_33_1678_0 & ~i_8_33_1733_0 & i_8_33_1778_0 & ~i_8_33_1805_0 & ~i_8_33_2017_0 & ~i_8_33_2172_0 & ~i_8_33_2264_0) | (i_8_33_193_0 & ~i_8_33_935_0 & i_8_33_2245_0 & ~i_8_33_2292_0))) | (~i_8_33_1091_0 & ((~i_8_33_345_0 & ((~i_8_33_923_0 & ~i_8_33_992_0 & ~i_8_33_366_0 & ~i_8_33_718_0 & ~i_8_33_1274_0 & ~i_8_33_1470_0 & i_8_33_1490_0 & ~i_8_33_1562_0) | (~i_8_33_719_0 & ~i_8_33_921_0 & ~i_8_33_1102_0 & i_8_33_1263_0 & i_8_33_1678_0 & ~i_8_33_2031_0))) | (~i_8_33_348_0 & ~i_8_33_479_0 & ~i_8_33_921_0 & i_8_33_1263_0 & ~i_8_33_1473_0 & ~i_8_33_1700_0 & ~i_8_33_1939_0 & ~i_8_33_2017_0 & ~i_8_33_2031_0 & ~i_8_33_2292_0))) | (~i_8_33_510_0 & ((i_8_33_653_0 & ~i_8_33_935_0 & ~i_8_33_1473_0 & ~i_8_33_2017_0 & ~i_8_33_2175_0 & i_8_33_2249_0) | (~i_8_33_1259_0 & i_8_33_1301_0 & ~i_8_33_1408_0 & i_8_33_1778_0 & ~i_8_33_2249_0))) | (~i_8_33_1753_0 & ((~i_8_33_385_0 & i_8_33_634_0 & ~i_8_33_1864_0 & ~i_8_33_2200_0 & i_8_33_2264_0) | (~i_8_33_718_0 & ~i_8_33_992_0 & ~i_8_33_1159_0 & i_8_33_1301_0 & ~i_8_33_1330_0 & ~i_8_33_1331_0 & ~i_8_33_1355_0 & ~i_8_33_1490_0 & ~i_8_33_1678_0 & ~i_8_33_1993_0 & ~i_8_33_2291_0))) | (i_8_33_651_0 & ~i_8_33_921_0 & i_8_33_1263_0 & ~i_8_33_1408_0 & ~i_8_33_1587_0) | (~i_8_33_348_0 & ~i_8_33_552_0 & ~i_8_33_1471_0 & i_8_33_1489_0 & i_8_33_1678_0 & ~i_8_33_2291_0))) | (~i_8_33_453_0 & ((~i_8_33_49_0 & ~i_8_33_385_0 & ((~i_8_33_1473_0 & i_8_33_1587_0 & ~i_8_33_1733_0 & ~i_8_33_1753_0 & ~i_8_33_1774_0 & ~i_8_33_1776_0) | (~i_8_33_718_0 & ~i_8_33_1170_0 & i_8_33_1774_0 & ~i_8_33_1788_0 & ~i_8_33_1993_0 & ~i_8_33_2017_0 & ~i_8_33_2291_0))) | (~i_8_33_76_0 & ~i_8_33_921_0 & ((~i_8_33_53_0 & i_8_33_193_0 & ~i_8_33_348_0 & ~i_8_33_773_0 & ~i_8_33_1159_0 & ~i_8_33_1263_0 & ~i_8_33_1471_0 & ~i_8_33_1549_0 & ~i_8_33_1805_0) | (~i_8_33_805_0 & i_8_33_885_0 & ~i_8_33_1170_0 & ~i_8_33_1470_0 & ~i_8_33_2017_0 & ~i_8_33_2249_0))) | (~i_8_33_1778_0 & ((~i_8_33_48_0 & ~i_8_33_348_0 & i_8_33_552_0 & ~i_8_33_773_0 & ~i_8_33_1678_0 & i_8_33_1788_0) | (~i_8_33_719_0 & ~i_8_33_796_0 & ~i_8_33_1301_0 & ~i_8_33_1355_0 & ~i_8_33_1753_0 & ~i_8_33_1774_0 & ~i_8_33_1788_0 & i_8_33_1993_0 & ~i_8_33_2174_0 & ~i_8_33_2264_0 & ~i_8_33_2291_0))) | (i_8_33_193_0 & ~i_8_33_1159_0 & i_8_33_1302_0 & ~i_8_33_2249_0) | (~i_8_33_1788_0 & i_8_33_1993_0 & i_8_33_652_0 & ~i_8_33_1330_0 & ~i_8_33_2017_0 & ~i_8_33_2194_0 & ~i_8_33_2206_0 & ~i_8_33_2292_0))) | (~i_8_33_164_0 & ((~i_8_33_48_0 & ~i_8_33_227_0 & ~i_8_33_345_0 & ~i_8_33_719_0 & i_8_33_1549_0 & ~i_8_33_1678_0 & i_8_33_1778_0 & ~i_8_33_1805_0 & ~i_8_33_2111_0 & ~i_8_33_2177_0 & ~i_8_33_2291_0) | (i_8_33_48_0 & i_8_33_49_0 & ~i_8_33_305_0 & ~i_8_33_366_0 & ~i_8_33_921_0 & ~i_8_33_1170_0 & ~i_8_33_1265_0 & ~i_8_33_1301_0 & ~i_8_33_1305_0 & ~i_8_33_1355_0 & ~i_8_33_2206_0 & ~i_8_33_2292_0 & ~i_8_33_1399_0 & ~i_8_33_1788_0))) | (~i_8_33_2292_0 & ((~i_8_33_193_0 & ((~i_8_33_258_0 & ~i_8_33_552_0 & ~i_8_33_719_0 & ~i_8_33_1159_0 & ~i_8_33_1259_0 & ~i_8_33_1330_0 & i_8_33_1399_0 & ~i_8_33_1549_0 & ~i_8_33_1587_0 & ~i_8_33_1678_0) | (~i_8_33_30_0 & ~i_8_33_48_0 & ~i_8_33_385_0 & i_8_33_552_0 & ~i_8_33_773_0 & ~i_8_33_1258_0 & ~i_8_33_1301_0 & ~i_8_33_1305_0 & ~i_8_33_1331_0 & ~i_8_33_1470_0 & ~i_8_33_1473_0 & ~i_8_33_2031_0 & ~i_8_33_2175_0))) | (~i_8_33_48_0 & ~i_8_33_2031_0 & ((i_8_33_33_0 & ~i_8_33_1159_0 & ~i_8_33_1263_0 & ~i_8_33_1587_0) | (~i_8_33_348_0 & ~i_8_33_1102_0 & ~i_8_33_1753_0 & ~i_8_33_1939_0 & i_8_33_2244_0))) | (~i_8_33_719_0 & ((~i_8_33_653_0 & i_8_33_778_0 & ~i_8_33_797_0 & ~i_8_33_1330_0 & ~i_8_33_1331_0 & ~i_8_33_1471_0 & ~i_8_33_1562_0 & ~i_8_33_1753_0 & ~i_8_33_1788_0 & ~i_8_33_1864_0 & ~i_8_33_2111_0) | (i_8_33_653_0 & ~i_8_33_1274_0 & i_8_33_1778_0 & ~i_8_33_2276_0 & ~i_8_33_2291_0))) | (~i_8_33_2194_0 & ((~i_8_33_1549_0 & ((~i_8_33_53_0 & ~i_8_33_258_0 & ~i_8_33_479_0 & ~i_8_33_796_0 & ~i_8_33_805_0 & ~i_8_33_1305_0 & i_8_33_1489_0 & ~i_8_33_1805_0 & ~i_8_33_2200_0 & ~i_8_33_2245_0) | (~i_8_33_885_0 & ~i_8_33_921_0 & ~i_8_33_935_0 & ~i_8_33_1331_0 & ~i_8_33_1774_0 & i_8_33_1805_0 & ~i_8_33_1939_0 & ~i_8_33_2048_0 & i_8_33_2176_0 & ~i_8_33_2264_0))) | (i_8_33_652_0 & ~i_8_33_992_0 & ~i_8_33_1473_0 & ~i_8_33_2206_0 & i_8_33_2244_0))) | (i_8_33_348_0 & ~i_8_33_1159_0 & i_8_33_1773_0 & ~i_8_33_1993_0))) | (~i_8_33_258_0 & ((~i_8_33_53_0 & ~i_8_33_718_0 & ~i_8_33_773_0 & i_8_33_778_0 & ~i_8_33_805_0 & ~i_8_33_1274_0 & ~i_8_33_1331_0 & ~i_8_33_1470_0 & i_8_33_1489_0) | (i_8_33_585_0 & ~i_8_33_930_0 & ~i_8_33_1587_0 & i_8_33_1774_0 & i_8_33_1993_0))) | (~i_8_33_1473_0 & ((~i_8_33_348_0 & ~i_8_33_1788_0 & ((i_8_33_651_0 & ~i_8_33_718_0 & ~i_8_33_2017_0 & ~i_8_33_2206_0 & ~i_8_33_2245_0) | (i_8_33_193_0 & ~i_8_33_653_0 & ~i_8_33_921_0 & ~i_8_33_1159_0 & ~i_8_33_1259_0 & ~i_8_33_1274_0 & ~i_8_33_1331_0 & ~i_8_33_1549_0 & ~i_8_33_2031_0 & ~i_8_33_2276_0))) | (~i_8_33_1408_0 & ~i_8_33_2291_0 & ((~i_8_33_48_0 & ~i_8_33_305_0 & i_8_33_348_0 & ~i_8_33_1258_0 & ~i_8_33_1263_0 & ~i_8_33_1753_0 & ~i_8_33_1776_0) | (~i_8_33_53_0 & ~i_8_33_479_0 & ~i_8_33_796_0 & ~i_8_33_1159_0 & ~i_8_33_1259_0 & ~i_8_33_885_0 & ~i_8_33_930_0 & ~i_8_33_1471_0 & ~i_8_33_1562_0 & ~i_8_33_1587_0 & i_8_33_1993_0 & ~i_8_33_2172_0 & ~i_8_33_2206_0 & ~i_8_33_2264_0))))) | (~i_8_33_49_0 & ((~i_8_33_366_0 & ((~i_8_33_1102_0 & ~i_8_33_1170_0 & ~i_8_33_1263_0 & ~i_8_33_1753_0 & ~i_8_33_1774_0 & i_8_33_1776_0 & ~i_8_33_1864_0) | (~i_8_33_552_0 & i_8_33_585_0 & ~i_8_33_634_0 & ~i_8_33_718_0 & ~i_8_33_1490_0 & ~i_8_33_1562_0 & ~i_8_33_2017_0 & ~i_8_33_2175_0))) | (~i_8_33_385_0 & ((~i_8_33_305_0 & ~i_8_33_1159_0 & ~i_8_33_1170_0 & i_8_33_1549_0 & i_8_33_1776_0 & ~i_8_33_2017_0 & ~i_8_33_2111_0) | (~i_8_33_53_0 & ~i_8_33_719_0 & ~i_8_33_773_0 & ~i_8_33_1331_0 & i_8_33_1355_0 & ~i_8_33_1549_0 & ~i_8_33_1864_0 & ~i_8_33_2177_0 & ~i_8_33_2264_0 & ~i_8_33_2291_0))) | (~i_8_33_53_0 & ~i_8_33_305_0 & ((~i_8_33_1091_0 & ~i_8_33_1470_0 & i_8_33_1549_0 & ~i_8_33_1700_0 & i_8_33_1774_0 & ~i_8_33_2017_0 & ~i_8_33_2111_0 & ~i_8_33_2206_0) | (~i_8_33_510_0 & i_8_33_1265_0 & ~i_8_33_1408_0 & ~i_8_33_1778_0 & ~i_8_33_2291_0))))) | (~i_8_33_510_0 & ((~i_8_33_48_0 & ~i_8_33_305_0 & i_8_33_385_0 & ~i_8_33_652_0 & ~i_8_33_718_0 & ~i_8_33_773_0 & ~i_8_33_1330_0 & ~i_8_33_1331_0 & ~i_8_33_1753_0 & ~i_8_33_1788_0 & ~i_8_33_2176_0) | (~i_8_33_385_0 & ~i_8_33_1091_0 & i_8_33_1355_0 & ~i_8_33_1993_0 & i_8_33_2177_0 & ~i_8_33_2194_0 & ~i_8_33_2276_0))) | (~i_8_33_48_0 & ~i_8_33_1330_0 & ((~i_8_33_718_0 & i_8_33_885_0 & i_8_33_2172_0 & ~i_8_33_2249_0) | (~i_8_33_719_0 & i_8_33_890_0 & ~i_8_33_1274_0 & ~i_8_33_1331_0 & ~i_8_33_1753_0 & ~i_8_33_2031_0 & ~i_8_33_2264_0))) | (~i_8_33_385_0 & ((~i_8_33_1258_0 & ((~i_8_33_885_0 & i_8_33_1302_0 & i_8_33_1399_0 & ~i_8_33_2031_0 & i_8_33_2175_0) | (~i_8_33_890_0 & ~i_8_33_1355_0 & ~i_8_33_1408_0 & ~i_8_33_1700_0 & ~i_8_33_1753_0 & i_8_33_2249_0))) | (i_8_33_76_0 & ~i_8_33_345_0 & ~i_8_33_773_0 & ~i_8_33_1259_0 & i_8_33_1265_0 & ~i_8_33_1678_0 & ~i_8_33_1776_0 & ~i_8_33_2194_0 & ~i_8_33_2249_0))) | (~i_8_33_1549_0 & ((~i_8_33_719_0 & i_8_33_1265_0 & ~i_8_33_1331_0 & ~i_8_33_2017_0 & i_8_33_2174_0) | (i_8_33_651_0 & ~i_8_33_718_0 & ~i_8_33_1091_0 & ~i_8_33_2031_0 & ~i_8_33_2111_0 & i_8_33_2175_0))) | (i_8_33_479_0 & ~i_8_33_1562_0 & ~i_8_33_1805_0 & i_8_33_2048_0) | (~i_8_33_479_0 & ~i_8_33_805_0 & ~i_8_33_923_0 & i_8_33_992_0 & i_8_33_1733_0 & ~i_8_33_2246_0 & ~i_8_33_2291_0));
endmodule



// Benchmark "kernel_8_34" written by ABC on Sun Jul 19 10:03:38 2020

module kernel_8_34 ( 
    i_8_34_40_0, i_8_34_51_0, i_8_34_57_0, i_8_34_79_0, i_8_34_143_0,
    i_8_34_174_0, i_8_34_220_0, i_8_34_225_0, i_8_34_252_0, i_8_34_265_0,
    i_8_34_364_0, i_8_34_365_0, i_8_34_367_0, i_8_34_369_0, i_8_34_453_0,
    i_8_34_492_0, i_8_34_499_0, i_8_34_589_0, i_8_34_590_0, i_8_34_591_0,
    i_8_34_595_0, i_8_34_597_0, i_8_34_598_0, i_8_34_634_0, i_8_34_635_0,
    i_8_34_651_0, i_8_34_659_0, i_8_34_660_0, i_8_34_675_0, i_8_34_679_0,
    i_8_34_680_0, i_8_34_693_0, i_8_34_705_0, i_8_34_706_0, i_8_34_729_0,
    i_8_34_779_0, i_8_34_819_0, i_8_34_820_0, i_8_34_855_0, i_8_34_866_0,
    i_8_34_882_0, i_8_34_885_0, i_8_34_937_0, i_8_34_968_0, i_8_34_969_0,
    i_8_34_971_0, i_8_34_1035_0, i_8_34_1039_0, i_8_34_1137_0,
    i_8_34_1147_0, i_8_34_1164_0, i_8_34_1165_0, i_8_34_1182_0,
    i_8_34_1220_0, i_8_34_1227_0, i_8_34_1260_0, i_8_34_1262_0,
    i_8_34_1297_0, i_8_34_1318_0, i_8_34_1369_0, i_8_34_1389_0,
    i_8_34_1479_0, i_8_34_1507_0, i_8_34_1524_0, i_8_34_1545_0,
    i_8_34_1546_0, i_8_34_1547_0, i_8_34_1564_0, i_8_34_1607_0,
    i_8_34_1610_0, i_8_34_1614_0, i_8_34_1675_0, i_8_34_1677_0,
    i_8_34_1703_0, i_8_34_1714_0, i_8_34_1762_0, i_8_34_1807_0,
    i_8_34_1850_0, i_8_34_1885_0, i_8_34_1927_0, i_8_34_1981_0,
    i_8_34_1984_0, i_8_34_2004_0, i_8_34_2052_0, i_8_34_2056_0,
    i_8_34_2091_0, i_8_34_2100_0, i_8_34_2101_0, i_8_34_2133_0,
    i_8_34_2135_0, i_8_34_2155_0, i_8_34_2163_0, i_8_34_2173_0,
    i_8_34_2176_0, i_8_34_2214_0, i_8_34_2224_0, i_8_34_2227_0,
    i_8_34_2241_0, i_8_34_2244_0, i_8_34_2262_0,
    o_8_34_0_0  );
  input  i_8_34_40_0, i_8_34_51_0, i_8_34_57_0, i_8_34_79_0,
    i_8_34_143_0, i_8_34_174_0, i_8_34_220_0, i_8_34_225_0, i_8_34_252_0,
    i_8_34_265_0, i_8_34_364_0, i_8_34_365_0, i_8_34_367_0, i_8_34_369_0,
    i_8_34_453_0, i_8_34_492_0, i_8_34_499_0, i_8_34_589_0, i_8_34_590_0,
    i_8_34_591_0, i_8_34_595_0, i_8_34_597_0, i_8_34_598_0, i_8_34_634_0,
    i_8_34_635_0, i_8_34_651_0, i_8_34_659_0, i_8_34_660_0, i_8_34_675_0,
    i_8_34_679_0, i_8_34_680_0, i_8_34_693_0, i_8_34_705_0, i_8_34_706_0,
    i_8_34_729_0, i_8_34_779_0, i_8_34_819_0, i_8_34_820_0, i_8_34_855_0,
    i_8_34_866_0, i_8_34_882_0, i_8_34_885_0, i_8_34_937_0, i_8_34_968_0,
    i_8_34_969_0, i_8_34_971_0, i_8_34_1035_0, i_8_34_1039_0,
    i_8_34_1137_0, i_8_34_1147_0, i_8_34_1164_0, i_8_34_1165_0,
    i_8_34_1182_0, i_8_34_1220_0, i_8_34_1227_0, i_8_34_1260_0,
    i_8_34_1262_0, i_8_34_1297_0, i_8_34_1318_0, i_8_34_1369_0,
    i_8_34_1389_0, i_8_34_1479_0, i_8_34_1507_0, i_8_34_1524_0,
    i_8_34_1545_0, i_8_34_1546_0, i_8_34_1547_0, i_8_34_1564_0,
    i_8_34_1607_0, i_8_34_1610_0, i_8_34_1614_0, i_8_34_1675_0,
    i_8_34_1677_0, i_8_34_1703_0, i_8_34_1714_0, i_8_34_1762_0,
    i_8_34_1807_0, i_8_34_1850_0, i_8_34_1885_0, i_8_34_1927_0,
    i_8_34_1981_0, i_8_34_1984_0, i_8_34_2004_0, i_8_34_2052_0,
    i_8_34_2056_0, i_8_34_2091_0, i_8_34_2100_0, i_8_34_2101_0,
    i_8_34_2133_0, i_8_34_2135_0, i_8_34_2155_0, i_8_34_2163_0,
    i_8_34_2173_0, i_8_34_2176_0, i_8_34_2214_0, i_8_34_2224_0,
    i_8_34_2227_0, i_8_34_2241_0, i_8_34_2244_0, i_8_34_2262_0;
  output o_8_34_0_0;
  assign o_8_34_0_0 = 0;
endmodule



// Benchmark "kernel_8_35" written by ABC on Sun Jul 19 10:03:39 2020

module kernel_8_35 ( 
    i_8_35_25_0, i_8_35_28_0, i_8_35_31_0, i_8_35_83_0, i_8_35_203_0,
    i_8_35_299_0, i_8_35_352_0, i_8_35_371_0, i_8_35_418_0, i_8_35_440_0,
    i_8_35_443_0, i_8_35_469_0, i_8_35_478_0, i_8_35_481_0, i_8_35_482_0,
    i_8_35_484_0, i_8_35_496_0, i_8_35_587_0, i_8_35_667_0, i_8_35_671_0,
    i_8_35_793_0, i_8_35_815_0, i_8_35_918_0, i_8_35_919_0, i_8_35_1003_0,
    i_8_35_1008_0, i_8_35_1013_0, i_8_35_1027_0, i_8_35_1108_0,
    i_8_35_1109_0, i_8_35_1125_0, i_8_35_1126_0, i_8_35_1127_0,
    i_8_35_1135_0, i_8_35_1139_0, i_8_35_1157_0, i_8_35_1217_0,
    i_8_35_1234_0, i_8_35_1256_0, i_8_35_1325_0, i_8_35_1346_0,
    i_8_35_1348_0, i_8_35_1435_0, i_8_35_1437_0, i_8_35_1468_0,
    i_8_35_1506_0, i_8_35_1521_0, i_8_35_1548_0, i_8_35_1556_0,
    i_8_35_1582_0, i_8_35_1603_0, i_8_35_1612_0, i_8_35_1640_0,
    i_8_35_1668_0, i_8_35_1669_0, i_8_35_1674_0, i_8_35_1675_0,
    i_8_35_1703_0, i_8_35_1704_0, i_8_35_1705_0, i_8_35_1714_0,
    i_8_35_1715_0, i_8_35_1717_0, i_8_35_1720_0, i_8_35_1746_0,
    i_8_35_1748_0, i_8_35_1749_0, i_8_35_1750_0, i_8_35_1751_0,
    i_8_35_1752_0, i_8_35_1776_0, i_8_35_1785_0, i_8_35_1791_0,
    i_8_35_1801_0, i_8_35_1808_0, i_8_35_1809_0, i_8_35_1812_0,
    i_8_35_1813_0, i_8_35_1838_0, i_8_35_1849_0, i_8_35_1859_0,
    i_8_35_1882_0, i_8_35_1918_0, i_8_35_1947_0, i_8_35_1951_0,
    i_8_35_1964_0, i_8_35_1986_0, i_8_35_1996_0, i_8_35_2000_0,
    i_8_35_2044_0, i_8_35_2107_0, i_8_35_2111_0, i_8_35_2125_0,
    i_8_35_2128_0, i_8_35_2143_0, i_8_35_2180_0, i_8_35_2188_0,
    i_8_35_2189_0, i_8_35_2245_0, i_8_35_2289_0,
    o_8_35_0_0  );
  input  i_8_35_25_0, i_8_35_28_0, i_8_35_31_0, i_8_35_83_0,
    i_8_35_203_0, i_8_35_299_0, i_8_35_352_0, i_8_35_371_0, i_8_35_418_0,
    i_8_35_440_0, i_8_35_443_0, i_8_35_469_0, i_8_35_478_0, i_8_35_481_0,
    i_8_35_482_0, i_8_35_484_0, i_8_35_496_0, i_8_35_587_0, i_8_35_667_0,
    i_8_35_671_0, i_8_35_793_0, i_8_35_815_0, i_8_35_918_0, i_8_35_919_0,
    i_8_35_1003_0, i_8_35_1008_0, i_8_35_1013_0, i_8_35_1027_0,
    i_8_35_1108_0, i_8_35_1109_0, i_8_35_1125_0, i_8_35_1126_0,
    i_8_35_1127_0, i_8_35_1135_0, i_8_35_1139_0, i_8_35_1157_0,
    i_8_35_1217_0, i_8_35_1234_0, i_8_35_1256_0, i_8_35_1325_0,
    i_8_35_1346_0, i_8_35_1348_0, i_8_35_1435_0, i_8_35_1437_0,
    i_8_35_1468_0, i_8_35_1506_0, i_8_35_1521_0, i_8_35_1548_0,
    i_8_35_1556_0, i_8_35_1582_0, i_8_35_1603_0, i_8_35_1612_0,
    i_8_35_1640_0, i_8_35_1668_0, i_8_35_1669_0, i_8_35_1674_0,
    i_8_35_1675_0, i_8_35_1703_0, i_8_35_1704_0, i_8_35_1705_0,
    i_8_35_1714_0, i_8_35_1715_0, i_8_35_1717_0, i_8_35_1720_0,
    i_8_35_1746_0, i_8_35_1748_0, i_8_35_1749_0, i_8_35_1750_0,
    i_8_35_1751_0, i_8_35_1752_0, i_8_35_1776_0, i_8_35_1785_0,
    i_8_35_1791_0, i_8_35_1801_0, i_8_35_1808_0, i_8_35_1809_0,
    i_8_35_1812_0, i_8_35_1813_0, i_8_35_1838_0, i_8_35_1849_0,
    i_8_35_1859_0, i_8_35_1882_0, i_8_35_1918_0, i_8_35_1947_0,
    i_8_35_1951_0, i_8_35_1964_0, i_8_35_1986_0, i_8_35_1996_0,
    i_8_35_2000_0, i_8_35_2044_0, i_8_35_2107_0, i_8_35_2111_0,
    i_8_35_2125_0, i_8_35_2128_0, i_8_35_2143_0, i_8_35_2180_0,
    i_8_35_2188_0, i_8_35_2189_0, i_8_35_2245_0, i_8_35_2289_0;
  output o_8_35_0_0;
  assign o_8_35_0_0 = 0;
endmodule



// Benchmark "kernel_8_36" written by ABC on Sun Jul 19 10:03:39 2020

module kernel_8_36 ( 
    i_8_36_31_0, i_8_36_33_0, i_8_36_35_0, i_8_36_43_0, i_8_36_49_0,
    i_8_36_54_0, i_8_36_57_0, i_8_36_73_0, i_8_36_93_0, i_8_36_94_0,
    i_8_36_101_0, i_8_36_183_0, i_8_36_228_0, i_8_36_230_0, i_8_36_238_0,
    i_8_36_300_0, i_8_36_334_0, i_8_36_345_0, i_8_36_360_0, i_8_36_368_0,
    i_8_36_380_0, i_8_36_417_0, i_8_36_472_0, i_8_36_489_0, i_8_36_503_0,
    i_8_36_508_0, i_8_36_527_0, i_8_36_528_0, i_8_36_571_0, i_8_36_599_0,
    i_8_36_617_0, i_8_36_634_0, i_8_36_670_0, i_8_36_686_0, i_8_36_689_0,
    i_8_36_710_0, i_8_36_733_0, i_8_36_760_0, i_8_36_764_0, i_8_36_775_0,
    i_8_36_780_0, i_8_36_781_0, i_8_36_805_0, i_8_36_809_0, i_8_36_826_0,
    i_8_36_841_0, i_8_36_859_0, i_8_36_877_0, i_8_36_883_0, i_8_36_904_0,
    i_8_36_939_0, i_8_36_940_0, i_8_36_941_0, i_8_36_990_0, i_8_36_1075_0,
    i_8_36_1144_0, i_8_36_1160_0, i_8_36_1169_0, i_8_36_1228_0,
    i_8_36_1229_0, i_8_36_1236_0, i_8_36_1294_0, i_8_36_1300_0,
    i_8_36_1312_0, i_8_36_1331_0, i_8_36_1399_0, i_8_36_1467_0,
    i_8_36_1492_0, i_8_36_1506_0, i_8_36_1539_0, i_8_36_1585_0,
    i_8_36_1625_0, i_8_36_1632_0, i_8_36_1655_0, i_8_36_1678_0,
    i_8_36_1681_0, i_8_36_1682_0, i_8_36_1696_0, i_8_36_1697_0,
    i_8_36_1723_0, i_8_36_1741_0, i_8_36_1750_0, i_8_36_1753_0,
    i_8_36_1784_0, i_8_36_1813_0, i_8_36_1835_0, i_8_36_1903_0,
    i_8_36_1986_0, i_8_36_2058_0, i_8_36_2059_0, i_8_36_2098_0,
    i_8_36_2119_0, i_8_36_2137_0, i_8_36_2171_0, i_8_36_2173_0,
    i_8_36_2176_0, i_8_36_2191_0, i_8_36_2276_0, i_8_36_2296_0,
    i_8_36_2299_0,
    o_8_36_0_0  );
  input  i_8_36_31_0, i_8_36_33_0, i_8_36_35_0, i_8_36_43_0, i_8_36_49_0,
    i_8_36_54_0, i_8_36_57_0, i_8_36_73_0, i_8_36_93_0, i_8_36_94_0,
    i_8_36_101_0, i_8_36_183_0, i_8_36_228_0, i_8_36_230_0, i_8_36_238_0,
    i_8_36_300_0, i_8_36_334_0, i_8_36_345_0, i_8_36_360_0, i_8_36_368_0,
    i_8_36_380_0, i_8_36_417_0, i_8_36_472_0, i_8_36_489_0, i_8_36_503_0,
    i_8_36_508_0, i_8_36_527_0, i_8_36_528_0, i_8_36_571_0, i_8_36_599_0,
    i_8_36_617_0, i_8_36_634_0, i_8_36_670_0, i_8_36_686_0, i_8_36_689_0,
    i_8_36_710_0, i_8_36_733_0, i_8_36_760_0, i_8_36_764_0, i_8_36_775_0,
    i_8_36_780_0, i_8_36_781_0, i_8_36_805_0, i_8_36_809_0, i_8_36_826_0,
    i_8_36_841_0, i_8_36_859_0, i_8_36_877_0, i_8_36_883_0, i_8_36_904_0,
    i_8_36_939_0, i_8_36_940_0, i_8_36_941_0, i_8_36_990_0, i_8_36_1075_0,
    i_8_36_1144_0, i_8_36_1160_0, i_8_36_1169_0, i_8_36_1228_0,
    i_8_36_1229_0, i_8_36_1236_0, i_8_36_1294_0, i_8_36_1300_0,
    i_8_36_1312_0, i_8_36_1331_0, i_8_36_1399_0, i_8_36_1467_0,
    i_8_36_1492_0, i_8_36_1506_0, i_8_36_1539_0, i_8_36_1585_0,
    i_8_36_1625_0, i_8_36_1632_0, i_8_36_1655_0, i_8_36_1678_0,
    i_8_36_1681_0, i_8_36_1682_0, i_8_36_1696_0, i_8_36_1697_0,
    i_8_36_1723_0, i_8_36_1741_0, i_8_36_1750_0, i_8_36_1753_0,
    i_8_36_1784_0, i_8_36_1813_0, i_8_36_1835_0, i_8_36_1903_0,
    i_8_36_1986_0, i_8_36_2058_0, i_8_36_2059_0, i_8_36_2098_0,
    i_8_36_2119_0, i_8_36_2137_0, i_8_36_2171_0, i_8_36_2173_0,
    i_8_36_2176_0, i_8_36_2191_0, i_8_36_2276_0, i_8_36_2296_0,
    i_8_36_2299_0;
  output o_8_36_0_0;
  assign o_8_36_0_0 = 0;
endmodule



// Benchmark "kernel_8_37" written by ABC on Sun Jul 19 10:03:41 2020

module kernel_8_37 ( 
    i_8_37_42_0, i_8_37_70_0, i_8_37_78_0, i_8_37_87_0, i_8_37_94_0,
    i_8_37_102_0, i_8_37_283_0, i_8_37_286_0, i_8_37_303_0, i_8_37_310_0,
    i_8_37_322_0, i_8_37_365_0, i_8_37_394_0, i_8_37_400_0, i_8_37_403_0,
    i_8_37_420_0, i_8_37_421_0, i_8_37_444_0, i_8_37_511_0, i_8_37_529_0,
    i_8_37_552_0, i_8_37_571_0, i_8_37_573_0, i_8_37_633_0, i_8_37_637_0,
    i_8_37_642_0, i_8_37_643_0, i_8_37_652_0, i_8_37_662_0, i_8_37_706_0,
    i_8_37_760_0, i_8_37_814_0, i_8_37_825_0, i_8_37_861_0, i_8_37_871_0,
    i_8_37_895_0, i_8_37_970_0, i_8_37_992_0, i_8_37_1071_0, i_8_37_1086_0,
    i_8_37_1104_0, i_8_37_1131_0, i_8_37_1156_0, i_8_37_1236_0,
    i_8_37_1262_0, i_8_37_1291_0, i_8_37_1318_0, i_8_37_1330_0,
    i_8_37_1338_0, i_8_37_1345_0, i_8_37_1365_0, i_8_37_1366_0,
    i_8_37_1393_0, i_8_37_1402_0, i_8_37_1407_0, i_8_37_1411_0,
    i_8_37_1425_0, i_8_37_1438_0, i_8_37_1464_0, i_8_37_1465_0,
    i_8_37_1471_0, i_8_37_1473_0, i_8_37_1479_0, i_8_37_1482_0,
    i_8_37_1483_0, i_8_37_1486_0, i_8_37_1515_0, i_8_37_1516_0,
    i_8_37_1518_0, i_8_37_1524_0, i_8_37_1527_0, i_8_37_1528_0,
    i_8_37_1536_0, i_8_37_1554_0, i_8_37_1635_0, i_8_37_1660_0,
    i_8_37_1669_0, i_8_37_1671_0, i_8_37_1676_0, i_8_37_1681_0,
    i_8_37_1690_0, i_8_37_1696_0, i_8_37_1704_0, i_8_37_1705_0,
    i_8_37_1707_0, i_8_37_1708_0, i_8_37_1779_0, i_8_37_1794_0,
    i_8_37_1823_0, i_8_37_1839_0, i_8_37_1840_0, i_8_37_1843_0,
    i_8_37_1914_0, i_8_37_1938_0, i_8_37_1977_0, i_8_37_2146_0,
    i_8_37_2149_0, i_8_37_2206_0, i_8_37_2223_0, i_8_37_2294_0,
    o_8_37_0_0  );
  input  i_8_37_42_0, i_8_37_70_0, i_8_37_78_0, i_8_37_87_0, i_8_37_94_0,
    i_8_37_102_0, i_8_37_283_0, i_8_37_286_0, i_8_37_303_0, i_8_37_310_0,
    i_8_37_322_0, i_8_37_365_0, i_8_37_394_0, i_8_37_400_0, i_8_37_403_0,
    i_8_37_420_0, i_8_37_421_0, i_8_37_444_0, i_8_37_511_0, i_8_37_529_0,
    i_8_37_552_0, i_8_37_571_0, i_8_37_573_0, i_8_37_633_0, i_8_37_637_0,
    i_8_37_642_0, i_8_37_643_0, i_8_37_652_0, i_8_37_662_0, i_8_37_706_0,
    i_8_37_760_0, i_8_37_814_0, i_8_37_825_0, i_8_37_861_0, i_8_37_871_0,
    i_8_37_895_0, i_8_37_970_0, i_8_37_992_0, i_8_37_1071_0, i_8_37_1086_0,
    i_8_37_1104_0, i_8_37_1131_0, i_8_37_1156_0, i_8_37_1236_0,
    i_8_37_1262_0, i_8_37_1291_0, i_8_37_1318_0, i_8_37_1330_0,
    i_8_37_1338_0, i_8_37_1345_0, i_8_37_1365_0, i_8_37_1366_0,
    i_8_37_1393_0, i_8_37_1402_0, i_8_37_1407_0, i_8_37_1411_0,
    i_8_37_1425_0, i_8_37_1438_0, i_8_37_1464_0, i_8_37_1465_0,
    i_8_37_1471_0, i_8_37_1473_0, i_8_37_1479_0, i_8_37_1482_0,
    i_8_37_1483_0, i_8_37_1486_0, i_8_37_1515_0, i_8_37_1516_0,
    i_8_37_1518_0, i_8_37_1524_0, i_8_37_1527_0, i_8_37_1528_0,
    i_8_37_1536_0, i_8_37_1554_0, i_8_37_1635_0, i_8_37_1660_0,
    i_8_37_1669_0, i_8_37_1671_0, i_8_37_1676_0, i_8_37_1681_0,
    i_8_37_1690_0, i_8_37_1696_0, i_8_37_1704_0, i_8_37_1705_0,
    i_8_37_1707_0, i_8_37_1708_0, i_8_37_1779_0, i_8_37_1794_0,
    i_8_37_1823_0, i_8_37_1839_0, i_8_37_1840_0, i_8_37_1843_0,
    i_8_37_1914_0, i_8_37_1938_0, i_8_37_1977_0, i_8_37_2146_0,
    i_8_37_2149_0, i_8_37_2206_0, i_8_37_2223_0, i_8_37_2294_0;
  output o_8_37_0_0;
  assign o_8_37_0_0 = 0;
endmodule



// Benchmark "kernel_8_38" written by ABC on Sun Jul 19 10:03:41 2020

module kernel_8_38 ( 
    i_8_38_25_0, i_8_38_170_0, i_8_38_247_0, i_8_38_293_0, i_8_38_296_0,
    i_8_38_319_0, i_8_38_329_0, i_8_38_334_0, i_8_38_341_0, i_8_38_361_0,
    i_8_38_363_0, i_8_38_366_0, i_8_38_367_0, i_8_38_383_0, i_8_38_454_0,
    i_8_38_480_0, i_8_38_535_0, i_8_38_553_0, i_8_38_562_0, i_8_38_580_0,
    i_8_38_592_0, i_8_38_604_0, i_8_38_608_0, i_8_38_621_0, i_8_38_628_0,
    i_8_38_631_0, i_8_38_634_0, i_8_38_662_0, i_8_38_693_0, i_8_38_696_0,
    i_8_38_698_0, i_8_38_703_0, i_8_38_705_0, i_8_38_714_0, i_8_38_718_0,
    i_8_38_719_0, i_8_38_783_0, i_8_38_809_0, i_8_38_840_0, i_8_38_843_0,
    i_8_38_871_0, i_8_38_880_0, i_8_38_954_0, i_8_38_957_0, i_8_38_966_0,
    i_8_38_969_0, i_8_38_1015_0, i_8_38_1051_0, i_8_38_1075_0,
    i_8_38_1076_0, i_8_38_1115_0, i_8_38_1226_0, i_8_38_1228_0,
    i_8_38_1231_0, i_8_38_1240_0, i_8_38_1273_0, i_8_38_1285_0,
    i_8_38_1286_0, i_8_38_1321_0, i_8_38_1330_0, i_8_38_1372_0,
    i_8_38_1445_0, i_8_38_1456_0, i_8_38_1470_0, i_8_38_1518_0,
    i_8_38_1542_0, i_8_38_1552_0, i_8_38_1553_0, i_8_38_1560_0,
    i_8_38_1561_0, i_8_38_1563_0, i_8_38_1571_0, i_8_38_1591_0,
    i_8_38_1624_0, i_8_38_1632_0, i_8_38_1668_0, i_8_38_1680_0,
    i_8_38_1704_0, i_8_38_1708_0, i_8_38_1733_0, i_8_38_1808_0,
    i_8_38_1809_0, i_8_38_1825_0, i_8_38_1835_0, i_8_38_1854_0,
    i_8_38_1862_0, i_8_38_1870_0, i_8_38_1885_0, i_8_38_1912_0,
    i_8_38_1966_0, i_8_38_1992_0, i_8_38_1996_0, i_8_38_2132_0,
    i_8_38_2134_0, i_8_38_2147_0, i_8_38_2217_0, i_8_38_2244_0,
    i_8_38_2245_0, i_8_38_2248_0, i_8_38_2281_0,
    o_8_38_0_0  );
  input  i_8_38_25_0, i_8_38_170_0, i_8_38_247_0, i_8_38_293_0,
    i_8_38_296_0, i_8_38_319_0, i_8_38_329_0, i_8_38_334_0, i_8_38_341_0,
    i_8_38_361_0, i_8_38_363_0, i_8_38_366_0, i_8_38_367_0, i_8_38_383_0,
    i_8_38_454_0, i_8_38_480_0, i_8_38_535_0, i_8_38_553_0, i_8_38_562_0,
    i_8_38_580_0, i_8_38_592_0, i_8_38_604_0, i_8_38_608_0, i_8_38_621_0,
    i_8_38_628_0, i_8_38_631_0, i_8_38_634_0, i_8_38_662_0, i_8_38_693_0,
    i_8_38_696_0, i_8_38_698_0, i_8_38_703_0, i_8_38_705_0, i_8_38_714_0,
    i_8_38_718_0, i_8_38_719_0, i_8_38_783_0, i_8_38_809_0, i_8_38_840_0,
    i_8_38_843_0, i_8_38_871_0, i_8_38_880_0, i_8_38_954_0, i_8_38_957_0,
    i_8_38_966_0, i_8_38_969_0, i_8_38_1015_0, i_8_38_1051_0,
    i_8_38_1075_0, i_8_38_1076_0, i_8_38_1115_0, i_8_38_1226_0,
    i_8_38_1228_0, i_8_38_1231_0, i_8_38_1240_0, i_8_38_1273_0,
    i_8_38_1285_0, i_8_38_1286_0, i_8_38_1321_0, i_8_38_1330_0,
    i_8_38_1372_0, i_8_38_1445_0, i_8_38_1456_0, i_8_38_1470_0,
    i_8_38_1518_0, i_8_38_1542_0, i_8_38_1552_0, i_8_38_1553_0,
    i_8_38_1560_0, i_8_38_1561_0, i_8_38_1563_0, i_8_38_1571_0,
    i_8_38_1591_0, i_8_38_1624_0, i_8_38_1632_0, i_8_38_1668_0,
    i_8_38_1680_0, i_8_38_1704_0, i_8_38_1708_0, i_8_38_1733_0,
    i_8_38_1808_0, i_8_38_1809_0, i_8_38_1825_0, i_8_38_1835_0,
    i_8_38_1854_0, i_8_38_1862_0, i_8_38_1870_0, i_8_38_1885_0,
    i_8_38_1912_0, i_8_38_1966_0, i_8_38_1992_0, i_8_38_1996_0,
    i_8_38_2132_0, i_8_38_2134_0, i_8_38_2147_0, i_8_38_2217_0,
    i_8_38_2244_0, i_8_38_2245_0, i_8_38_2248_0, i_8_38_2281_0;
  output o_8_38_0_0;
  assign o_8_38_0_0 = 0;
endmodule



// Benchmark "kernel_8_39" written by ABC on Sun Jul 19 10:03:42 2020

module kernel_8_39 ( 
    i_8_39_63_0, i_8_39_64_0, i_8_39_117_0, i_8_39_138_0, i_8_39_147_0,
    i_8_39_192_0, i_8_39_237_0, i_8_39_262_0, i_8_39_273_0, i_8_39_319_0,
    i_8_39_352_0, i_8_39_360_0, i_8_39_364_0, i_8_39_365_0, i_8_39_369_0,
    i_8_39_417_0, i_8_39_450_0, i_8_39_451_0, i_8_39_457_0, i_8_39_460_0,
    i_8_39_489_0, i_8_39_531_0, i_8_39_549_0, i_8_39_585_0, i_8_39_603_0,
    i_8_39_606_0, i_8_39_607_0, i_8_39_651_0, i_8_39_661_0, i_8_39_675_0,
    i_8_39_694_0, i_8_39_700_0, i_8_39_703_0, i_8_39_704_0, i_8_39_729_0,
    i_8_39_751_0, i_8_39_810_0, i_8_39_814_0, i_8_39_828_0, i_8_39_829_0,
    i_8_39_849_0, i_8_39_876_0, i_8_39_981_0, i_8_39_1063_0, i_8_39_1080_0,
    i_8_39_1101_0, i_8_39_1102_0, i_8_39_1114_0, i_8_39_1138_0,
    i_8_39_1162_0, i_8_39_1200_0, i_8_39_1260_0, i_8_39_1278_0,
    i_8_39_1296_0, i_8_39_1306_0, i_8_39_1324_0, i_8_39_1355_0,
    i_8_39_1377_0, i_8_39_1378_0, i_8_39_1386_0, i_8_39_1395_0,
    i_8_39_1396_0, i_8_39_1408_0, i_8_39_1452_0, i_8_39_1468_0,
    i_8_39_1486_0, i_8_39_1488_0, i_8_39_1503_0, i_8_39_1540_0,
    i_8_39_1548_0, i_8_39_1562_0, i_8_39_1624_0, i_8_39_1647_0,
    i_8_39_1650_0, i_8_39_1668_0, i_8_39_1674_0, i_8_39_1681_0,
    i_8_39_1702_0, i_8_39_1758_0, i_8_39_1764_0, i_8_39_1792_0,
    i_8_39_1801_0, i_8_39_1821_0, i_8_39_1824_0, i_8_39_1828_0,
    i_8_39_1857_0, i_8_39_1873_0, i_8_39_1885_0, i_8_39_1908_0,
    i_8_39_1944_0, i_8_39_1962_0, i_8_39_1972_0, i_8_39_1995_0,
    i_8_39_2007_0, i_8_39_2008_0, i_8_39_2089_0, i_8_39_2134_0,
    i_8_39_2148_0, i_8_39_2241_0, i_8_39_2295_0,
    o_8_39_0_0  );
  input  i_8_39_63_0, i_8_39_64_0, i_8_39_117_0, i_8_39_138_0,
    i_8_39_147_0, i_8_39_192_0, i_8_39_237_0, i_8_39_262_0, i_8_39_273_0,
    i_8_39_319_0, i_8_39_352_0, i_8_39_360_0, i_8_39_364_0, i_8_39_365_0,
    i_8_39_369_0, i_8_39_417_0, i_8_39_450_0, i_8_39_451_0, i_8_39_457_0,
    i_8_39_460_0, i_8_39_489_0, i_8_39_531_0, i_8_39_549_0, i_8_39_585_0,
    i_8_39_603_0, i_8_39_606_0, i_8_39_607_0, i_8_39_651_0, i_8_39_661_0,
    i_8_39_675_0, i_8_39_694_0, i_8_39_700_0, i_8_39_703_0, i_8_39_704_0,
    i_8_39_729_0, i_8_39_751_0, i_8_39_810_0, i_8_39_814_0, i_8_39_828_0,
    i_8_39_829_0, i_8_39_849_0, i_8_39_876_0, i_8_39_981_0, i_8_39_1063_0,
    i_8_39_1080_0, i_8_39_1101_0, i_8_39_1102_0, i_8_39_1114_0,
    i_8_39_1138_0, i_8_39_1162_0, i_8_39_1200_0, i_8_39_1260_0,
    i_8_39_1278_0, i_8_39_1296_0, i_8_39_1306_0, i_8_39_1324_0,
    i_8_39_1355_0, i_8_39_1377_0, i_8_39_1378_0, i_8_39_1386_0,
    i_8_39_1395_0, i_8_39_1396_0, i_8_39_1408_0, i_8_39_1452_0,
    i_8_39_1468_0, i_8_39_1486_0, i_8_39_1488_0, i_8_39_1503_0,
    i_8_39_1540_0, i_8_39_1548_0, i_8_39_1562_0, i_8_39_1624_0,
    i_8_39_1647_0, i_8_39_1650_0, i_8_39_1668_0, i_8_39_1674_0,
    i_8_39_1681_0, i_8_39_1702_0, i_8_39_1758_0, i_8_39_1764_0,
    i_8_39_1792_0, i_8_39_1801_0, i_8_39_1821_0, i_8_39_1824_0,
    i_8_39_1828_0, i_8_39_1857_0, i_8_39_1873_0, i_8_39_1885_0,
    i_8_39_1908_0, i_8_39_1944_0, i_8_39_1962_0, i_8_39_1972_0,
    i_8_39_1995_0, i_8_39_2007_0, i_8_39_2008_0, i_8_39_2089_0,
    i_8_39_2134_0, i_8_39_2148_0, i_8_39_2241_0, i_8_39_2295_0;
  output o_8_39_0_0;
  assign o_8_39_0_0 = 0;
endmodule



// Benchmark "kernel_8_40" written by ABC on Sun Jul 19 10:03:43 2020

module kernel_8_40 ( 
    i_8_40_8_0, i_8_40_39_0, i_8_40_66_0, i_8_40_89_0, i_8_40_168_0,
    i_8_40_169_0, i_8_40_175_0, i_8_40_183_0, i_8_40_187_0, i_8_40_191_0,
    i_8_40_324_0, i_8_40_425_0, i_8_40_450_0, i_8_40_456_0, i_8_40_489_0,
    i_8_40_524_0, i_8_40_528_0, i_8_40_529_0, i_8_40_530_0, i_8_40_552_0,
    i_8_40_553_0, i_8_40_589_0, i_8_40_601_0, i_8_40_615_0, i_8_40_636_0,
    i_8_40_685_0, i_8_40_690_0, i_8_40_691_0, i_8_40_699_0, i_8_40_700_0,
    i_8_40_705_0, i_8_40_707_0, i_8_40_737_0, i_8_40_763_0, i_8_40_798_0,
    i_8_40_837_0, i_8_40_838_0, i_8_40_843_0, i_8_40_881_0, i_8_40_892_0,
    i_8_40_957_0, i_8_40_966_0, i_8_40_995_0, i_8_40_1029_0, i_8_40_1030_0,
    i_8_40_1044_0, i_8_40_1076_0, i_8_40_1078_0, i_8_40_1096_0,
    i_8_40_1114_0, i_8_40_1205_0, i_8_40_1213_0, i_8_40_1230_0,
    i_8_40_1239_0, i_8_40_1273_0, i_8_40_1276_0, i_8_40_1284_0,
    i_8_40_1285_0, i_8_40_1340_0, i_8_40_1353_0, i_8_40_1362_0,
    i_8_40_1426_0, i_8_40_1446_0, i_8_40_1447_0, i_8_40_1452_0,
    i_8_40_1471_0, i_8_40_1490_0, i_8_40_1570_0, i_8_40_1605_0,
    i_8_40_1681_0, i_8_40_1689_0, i_8_40_1723_0, i_8_40_1751_0,
    i_8_40_1762_0, i_8_40_1773_0, i_8_40_1776_0, i_8_40_1777_0,
    i_8_40_1815_0, i_8_40_1852_0, i_8_40_1862_0, i_8_40_1903_0,
    i_8_40_1904_0, i_8_40_1941_0, i_8_40_1996_0, i_8_40_2005_0,
    i_8_40_2074_0, i_8_40_2113_0, i_8_40_2140_0, i_8_40_2145_0,
    i_8_40_2150_0, i_8_40_2174_0, i_8_40_2175_0, i_8_40_2185_0,
    i_8_40_2212_0, i_8_40_2226_0, i_8_40_2233_0, i_8_40_2234_0,
    i_8_40_2265_0, i_8_40_2267_0, i_8_40_2289_0,
    o_8_40_0_0  );
  input  i_8_40_8_0, i_8_40_39_0, i_8_40_66_0, i_8_40_89_0, i_8_40_168_0,
    i_8_40_169_0, i_8_40_175_0, i_8_40_183_0, i_8_40_187_0, i_8_40_191_0,
    i_8_40_324_0, i_8_40_425_0, i_8_40_450_0, i_8_40_456_0, i_8_40_489_0,
    i_8_40_524_0, i_8_40_528_0, i_8_40_529_0, i_8_40_530_0, i_8_40_552_0,
    i_8_40_553_0, i_8_40_589_0, i_8_40_601_0, i_8_40_615_0, i_8_40_636_0,
    i_8_40_685_0, i_8_40_690_0, i_8_40_691_0, i_8_40_699_0, i_8_40_700_0,
    i_8_40_705_0, i_8_40_707_0, i_8_40_737_0, i_8_40_763_0, i_8_40_798_0,
    i_8_40_837_0, i_8_40_838_0, i_8_40_843_0, i_8_40_881_0, i_8_40_892_0,
    i_8_40_957_0, i_8_40_966_0, i_8_40_995_0, i_8_40_1029_0, i_8_40_1030_0,
    i_8_40_1044_0, i_8_40_1076_0, i_8_40_1078_0, i_8_40_1096_0,
    i_8_40_1114_0, i_8_40_1205_0, i_8_40_1213_0, i_8_40_1230_0,
    i_8_40_1239_0, i_8_40_1273_0, i_8_40_1276_0, i_8_40_1284_0,
    i_8_40_1285_0, i_8_40_1340_0, i_8_40_1353_0, i_8_40_1362_0,
    i_8_40_1426_0, i_8_40_1446_0, i_8_40_1447_0, i_8_40_1452_0,
    i_8_40_1471_0, i_8_40_1490_0, i_8_40_1570_0, i_8_40_1605_0,
    i_8_40_1681_0, i_8_40_1689_0, i_8_40_1723_0, i_8_40_1751_0,
    i_8_40_1762_0, i_8_40_1773_0, i_8_40_1776_0, i_8_40_1777_0,
    i_8_40_1815_0, i_8_40_1852_0, i_8_40_1862_0, i_8_40_1903_0,
    i_8_40_1904_0, i_8_40_1941_0, i_8_40_1996_0, i_8_40_2005_0,
    i_8_40_2074_0, i_8_40_2113_0, i_8_40_2140_0, i_8_40_2145_0,
    i_8_40_2150_0, i_8_40_2174_0, i_8_40_2175_0, i_8_40_2185_0,
    i_8_40_2212_0, i_8_40_2226_0, i_8_40_2233_0, i_8_40_2234_0,
    i_8_40_2265_0, i_8_40_2267_0, i_8_40_2289_0;
  output o_8_40_0_0;
  assign o_8_40_0_0 = 0;
endmodule



// Benchmark "kernel_8_41" written by ABC on Sun Jul 19 10:03:44 2020

module kernel_8_41 ( 
    i_8_41_13_0, i_8_41_23_0, i_8_41_35_0, i_8_41_85_0, i_8_41_118_0,
    i_8_41_121_0, i_8_41_122_0, i_8_41_139_0, i_8_41_148_0, i_8_41_189_0,
    i_8_41_328_0, i_8_41_348_0, i_8_41_362_0, i_8_41_450_0, i_8_41_483_0,
    i_8_41_484_0, i_8_41_499_0, i_8_41_538_0, i_8_41_552_0, i_8_41_556_0,
    i_8_41_589_0, i_8_41_607_0, i_8_41_636_0, i_8_41_662_0, i_8_41_679_0,
    i_8_41_682_0, i_8_41_686_0, i_8_41_694_0, i_8_41_697_0, i_8_41_699_0,
    i_8_41_733_0, i_8_41_755_0, i_8_41_781_0, i_8_41_785_0, i_8_41_797_0,
    i_8_41_823_0, i_8_41_839_0, i_8_41_843_0, i_8_41_958_0, i_8_41_968_0,
    i_8_41_973_0, i_8_41_977_0, i_8_41_1027_0, i_8_41_1030_0,
    i_8_41_1036_0, i_8_41_1057_0, i_8_41_1087_0, i_8_41_1111_0,
    i_8_41_1113_0, i_8_41_1127_0, i_8_41_1133_0, i_8_41_1157_0,
    i_8_41_1183_0, i_8_41_1230_0, i_8_41_1251_0, i_8_41_1255_0,
    i_8_41_1300_0, i_8_41_1337_0, i_8_41_1355_0, i_8_41_1552_0,
    i_8_41_1564_0, i_8_41_1588_0, i_8_41_1610_0, i_8_41_1612_0,
    i_8_41_1622_0, i_8_41_1624_0, i_8_41_1627_0, i_8_41_1628_0,
    i_8_41_1639_0, i_8_41_1669_0, i_8_41_1684_0, i_8_41_1694_0,
    i_8_41_1748_0, i_8_41_1750_0, i_8_41_1759_0, i_8_41_1768_0,
    i_8_41_1769_0, i_8_41_1777_0, i_8_41_1778_0, i_8_41_1791_0,
    i_8_41_1802_0, i_8_41_1805_0, i_8_41_1816_0, i_8_41_1858_0,
    i_8_41_1926_0, i_8_41_1939_0, i_8_41_1996_0, i_8_41_2011_0,
    i_8_41_2134_0, i_8_41_2138_0, i_8_41_2149_0, i_8_41_2150_0,
    i_8_41_2173_0, i_8_41_2229_0, i_8_41_2230_0, i_8_41_2232_0,
    i_8_41_2245_0, i_8_41_2246_0, i_8_41_2247_0, i_8_41_2263_0,
    o_8_41_0_0  );
  input  i_8_41_13_0, i_8_41_23_0, i_8_41_35_0, i_8_41_85_0,
    i_8_41_118_0, i_8_41_121_0, i_8_41_122_0, i_8_41_139_0, i_8_41_148_0,
    i_8_41_189_0, i_8_41_328_0, i_8_41_348_0, i_8_41_362_0, i_8_41_450_0,
    i_8_41_483_0, i_8_41_484_0, i_8_41_499_0, i_8_41_538_0, i_8_41_552_0,
    i_8_41_556_0, i_8_41_589_0, i_8_41_607_0, i_8_41_636_0, i_8_41_662_0,
    i_8_41_679_0, i_8_41_682_0, i_8_41_686_0, i_8_41_694_0, i_8_41_697_0,
    i_8_41_699_0, i_8_41_733_0, i_8_41_755_0, i_8_41_781_0, i_8_41_785_0,
    i_8_41_797_0, i_8_41_823_0, i_8_41_839_0, i_8_41_843_0, i_8_41_958_0,
    i_8_41_968_0, i_8_41_973_0, i_8_41_977_0, i_8_41_1027_0, i_8_41_1030_0,
    i_8_41_1036_0, i_8_41_1057_0, i_8_41_1087_0, i_8_41_1111_0,
    i_8_41_1113_0, i_8_41_1127_0, i_8_41_1133_0, i_8_41_1157_0,
    i_8_41_1183_0, i_8_41_1230_0, i_8_41_1251_0, i_8_41_1255_0,
    i_8_41_1300_0, i_8_41_1337_0, i_8_41_1355_0, i_8_41_1552_0,
    i_8_41_1564_0, i_8_41_1588_0, i_8_41_1610_0, i_8_41_1612_0,
    i_8_41_1622_0, i_8_41_1624_0, i_8_41_1627_0, i_8_41_1628_0,
    i_8_41_1639_0, i_8_41_1669_0, i_8_41_1684_0, i_8_41_1694_0,
    i_8_41_1748_0, i_8_41_1750_0, i_8_41_1759_0, i_8_41_1768_0,
    i_8_41_1769_0, i_8_41_1777_0, i_8_41_1778_0, i_8_41_1791_0,
    i_8_41_1802_0, i_8_41_1805_0, i_8_41_1816_0, i_8_41_1858_0,
    i_8_41_1926_0, i_8_41_1939_0, i_8_41_1996_0, i_8_41_2011_0,
    i_8_41_2134_0, i_8_41_2138_0, i_8_41_2149_0, i_8_41_2150_0,
    i_8_41_2173_0, i_8_41_2229_0, i_8_41_2230_0, i_8_41_2232_0,
    i_8_41_2245_0, i_8_41_2246_0, i_8_41_2247_0, i_8_41_2263_0;
  output o_8_41_0_0;
  assign o_8_41_0_0 = 0;
endmodule



// Benchmark "kernel_8_42" written by ABC on Sun Jul 19 10:03:45 2020

module kernel_8_42 ( 
    i_8_42_0_0, i_8_42_66_0, i_8_42_72_0, i_8_42_106_0, i_8_42_135_0,
    i_8_42_144_0, i_8_42_199_0, i_8_42_220_0, i_8_42_240_0, i_8_42_244_0,
    i_8_42_309_0, i_8_42_397_0, i_8_42_399_0, i_8_42_400_0, i_8_42_418_0,
    i_8_42_427_0, i_8_42_498_0, i_8_42_507_0, i_8_42_513_0, i_8_42_553_0,
    i_8_42_554_0, i_8_42_570_0, i_8_42_588_0, i_8_42_601_0, i_8_42_603_0,
    i_8_42_614_0, i_8_42_617_0, i_8_42_651_0, i_8_42_655_0, i_8_42_706_0,
    i_8_42_714_0, i_8_42_730_0, i_8_42_747_0, i_8_42_831_0, i_8_42_837_0,
    i_8_42_840_0, i_8_42_891_0, i_8_42_958_0, i_8_42_973_0, i_8_42_1108_0,
    i_8_42_1152_0, i_8_42_1170_0, i_8_42_1197_0, i_8_42_1200_0,
    i_8_42_1224_0, i_8_42_1236_0, i_8_42_1266_0, i_8_42_1294_0,
    i_8_42_1350_0, i_8_42_1353_0, i_8_42_1359_0, i_8_42_1363_0,
    i_8_42_1390_0, i_8_42_1399_0, i_8_42_1422_0, i_8_42_1431_0,
    i_8_42_1440_0, i_8_42_1461_0, i_8_42_1462_0, i_8_42_1467_0,
    i_8_42_1476_0, i_8_42_1494_0, i_8_42_1556_0, i_8_42_1632_0,
    i_8_42_1635_0, i_8_42_1692_0, i_8_42_1693_0, i_8_42_1722_0,
    i_8_42_1748_0, i_8_42_1749_0, i_8_42_1750_0, i_8_42_1751_0,
    i_8_42_1764_0, i_8_42_1782_0, i_8_42_1792_0, i_8_42_1805_0,
    i_8_42_1815_0, i_8_42_1822_0, i_8_42_1836_0, i_8_42_1840_0,
    i_8_42_1866_0, i_8_42_1881_0, i_8_42_1885_0, i_8_42_1917_0,
    i_8_42_1926_0, i_8_42_1947_0, i_8_42_1950_0, i_8_42_1974_0,
    i_8_42_1980_0, i_8_42_2007_0, i_8_42_2043_0, i_8_42_2044_0,
    i_8_42_2062_0, i_8_42_2116_0, i_8_42_2142_0, i_8_42_2143_0,
    i_8_42_2145_0, i_8_42_2146_0, i_8_42_2149_0, i_8_42_2248_0,
    o_8_42_0_0  );
  input  i_8_42_0_0, i_8_42_66_0, i_8_42_72_0, i_8_42_106_0,
    i_8_42_135_0, i_8_42_144_0, i_8_42_199_0, i_8_42_220_0, i_8_42_240_0,
    i_8_42_244_0, i_8_42_309_0, i_8_42_397_0, i_8_42_399_0, i_8_42_400_0,
    i_8_42_418_0, i_8_42_427_0, i_8_42_498_0, i_8_42_507_0, i_8_42_513_0,
    i_8_42_553_0, i_8_42_554_0, i_8_42_570_0, i_8_42_588_0, i_8_42_601_0,
    i_8_42_603_0, i_8_42_614_0, i_8_42_617_0, i_8_42_651_0, i_8_42_655_0,
    i_8_42_706_0, i_8_42_714_0, i_8_42_730_0, i_8_42_747_0, i_8_42_831_0,
    i_8_42_837_0, i_8_42_840_0, i_8_42_891_0, i_8_42_958_0, i_8_42_973_0,
    i_8_42_1108_0, i_8_42_1152_0, i_8_42_1170_0, i_8_42_1197_0,
    i_8_42_1200_0, i_8_42_1224_0, i_8_42_1236_0, i_8_42_1266_0,
    i_8_42_1294_0, i_8_42_1350_0, i_8_42_1353_0, i_8_42_1359_0,
    i_8_42_1363_0, i_8_42_1390_0, i_8_42_1399_0, i_8_42_1422_0,
    i_8_42_1431_0, i_8_42_1440_0, i_8_42_1461_0, i_8_42_1462_0,
    i_8_42_1467_0, i_8_42_1476_0, i_8_42_1494_0, i_8_42_1556_0,
    i_8_42_1632_0, i_8_42_1635_0, i_8_42_1692_0, i_8_42_1693_0,
    i_8_42_1722_0, i_8_42_1748_0, i_8_42_1749_0, i_8_42_1750_0,
    i_8_42_1751_0, i_8_42_1764_0, i_8_42_1782_0, i_8_42_1792_0,
    i_8_42_1805_0, i_8_42_1815_0, i_8_42_1822_0, i_8_42_1836_0,
    i_8_42_1840_0, i_8_42_1866_0, i_8_42_1881_0, i_8_42_1885_0,
    i_8_42_1917_0, i_8_42_1926_0, i_8_42_1947_0, i_8_42_1950_0,
    i_8_42_1974_0, i_8_42_1980_0, i_8_42_2007_0, i_8_42_2043_0,
    i_8_42_2044_0, i_8_42_2062_0, i_8_42_2116_0, i_8_42_2142_0,
    i_8_42_2143_0, i_8_42_2145_0, i_8_42_2146_0, i_8_42_2149_0,
    i_8_42_2248_0;
  output o_8_42_0_0;
  assign o_8_42_0_0 = 0;
endmodule



// Benchmark "kernel_8_43" written by ABC on Sun Jul 19 10:03:46 2020

module kernel_8_43 ( 
    i_8_43_3_0, i_8_43_30_0, i_8_43_31_0, i_8_43_34_0, i_8_43_42_0,
    i_8_43_94_0, i_8_43_99_0, i_8_43_100_0, i_8_43_117_0, i_8_43_120_0,
    i_8_43_126_0, i_8_43_220_0, i_8_43_274_0, i_8_43_279_0, i_8_43_288_0,
    i_8_43_309_0, i_8_43_315_0, i_8_43_345_0, i_8_43_348_0, i_8_43_356_0,
    i_8_43_378_0, i_8_43_381_0, i_8_43_384_0, i_8_43_402_0, i_8_43_427_0,
    i_8_43_432_0, i_8_43_433_0, i_8_43_435_0, i_8_43_442_0, i_8_43_517_0,
    i_8_43_527_0, i_8_43_530_0, i_8_43_547_0, i_8_43_660_0, i_8_43_665_0,
    i_8_43_723_0, i_8_43_774_0, i_8_43_814_0, i_8_43_819_0, i_8_43_841_0,
    i_8_43_861_0, i_8_43_894_0, i_8_43_913_0, i_8_43_967_0, i_8_43_972_0,
    i_8_43_981_0, i_8_43_999_0, i_8_43_1102_0, i_8_43_1200_0,
    i_8_43_1206_0, i_8_43_1251_0, i_8_43_1263_0, i_8_43_1266_0,
    i_8_43_1284_0, i_8_43_1372_0, i_8_43_1410_0, i_8_43_1434_0,
    i_8_43_1445_0, i_8_43_1453_0, i_8_43_1456_0, i_8_43_1491_0,
    i_8_43_1510_0, i_8_43_1539_0, i_8_43_1555_0, i_8_43_1565_0,
    i_8_43_1566_0, i_8_43_1584_0, i_8_43_1609_0, i_8_43_1611_0,
    i_8_43_1623_0, i_8_43_1627_0, i_8_43_1684_0, i_8_43_1755_0,
    i_8_43_1759_0, i_8_43_1776_0, i_8_43_1866_0, i_8_43_1873_0,
    i_8_43_1899_0, i_8_43_1902_0, i_8_43_1905_0, i_8_43_1936_0,
    i_8_43_1942_0, i_8_43_1975_0, i_8_43_1976_0, i_8_43_2001_0,
    i_8_43_2025_0, i_8_43_2062_0, i_8_43_2065_0, i_8_43_2080_0,
    i_8_43_2083_0, i_8_43_2115_0, i_8_43_2142_0, i_8_43_2143_0,
    i_8_43_2149_0, i_8_43_2169_0, i_8_43_2173_0, i_8_43_2187_0,
    i_8_43_2205_0, i_8_43_2209_0, i_8_43_2257_0,
    o_8_43_0_0  );
  input  i_8_43_3_0, i_8_43_30_0, i_8_43_31_0, i_8_43_34_0, i_8_43_42_0,
    i_8_43_94_0, i_8_43_99_0, i_8_43_100_0, i_8_43_117_0, i_8_43_120_0,
    i_8_43_126_0, i_8_43_220_0, i_8_43_274_0, i_8_43_279_0, i_8_43_288_0,
    i_8_43_309_0, i_8_43_315_0, i_8_43_345_0, i_8_43_348_0, i_8_43_356_0,
    i_8_43_378_0, i_8_43_381_0, i_8_43_384_0, i_8_43_402_0, i_8_43_427_0,
    i_8_43_432_0, i_8_43_433_0, i_8_43_435_0, i_8_43_442_0, i_8_43_517_0,
    i_8_43_527_0, i_8_43_530_0, i_8_43_547_0, i_8_43_660_0, i_8_43_665_0,
    i_8_43_723_0, i_8_43_774_0, i_8_43_814_0, i_8_43_819_0, i_8_43_841_0,
    i_8_43_861_0, i_8_43_894_0, i_8_43_913_0, i_8_43_967_0, i_8_43_972_0,
    i_8_43_981_0, i_8_43_999_0, i_8_43_1102_0, i_8_43_1200_0,
    i_8_43_1206_0, i_8_43_1251_0, i_8_43_1263_0, i_8_43_1266_0,
    i_8_43_1284_0, i_8_43_1372_0, i_8_43_1410_0, i_8_43_1434_0,
    i_8_43_1445_0, i_8_43_1453_0, i_8_43_1456_0, i_8_43_1491_0,
    i_8_43_1510_0, i_8_43_1539_0, i_8_43_1555_0, i_8_43_1565_0,
    i_8_43_1566_0, i_8_43_1584_0, i_8_43_1609_0, i_8_43_1611_0,
    i_8_43_1623_0, i_8_43_1627_0, i_8_43_1684_0, i_8_43_1755_0,
    i_8_43_1759_0, i_8_43_1776_0, i_8_43_1866_0, i_8_43_1873_0,
    i_8_43_1899_0, i_8_43_1902_0, i_8_43_1905_0, i_8_43_1936_0,
    i_8_43_1942_0, i_8_43_1975_0, i_8_43_1976_0, i_8_43_2001_0,
    i_8_43_2025_0, i_8_43_2062_0, i_8_43_2065_0, i_8_43_2080_0,
    i_8_43_2083_0, i_8_43_2115_0, i_8_43_2142_0, i_8_43_2143_0,
    i_8_43_2149_0, i_8_43_2169_0, i_8_43_2173_0, i_8_43_2187_0,
    i_8_43_2205_0, i_8_43_2209_0, i_8_43_2257_0;
  output o_8_43_0_0;
  assign o_8_43_0_0 = 0;
endmodule



// Benchmark "kernel_8_44" written by ABC on Sun Jul 19 10:03:47 2020

module kernel_8_44 ( 
    i_8_44_11_0, i_8_44_23_0, i_8_44_28_0, i_8_44_95_0, i_8_44_97_0,
    i_8_44_157_0, i_8_44_158_0, i_8_44_202_0, i_8_44_203_0, i_8_44_209_0,
    i_8_44_223_0, i_8_44_244_0, i_8_44_245_0, i_8_44_248_0, i_8_44_266_0,
    i_8_44_326_0, i_8_44_348_0, i_8_44_355_0, i_8_44_364_0, i_8_44_380_0,
    i_8_44_437_0, i_8_44_452_0, i_8_44_483_0, i_8_44_484_0, i_8_44_498_0,
    i_8_44_508_0, i_8_44_526_0, i_8_44_536_0, i_8_44_551_0, i_8_44_554_0,
    i_8_44_556_0, i_8_44_557_0, i_8_44_587_0, i_8_44_626_0, i_8_44_628_0,
    i_8_44_657_0, i_8_44_779_0, i_8_44_793_0, i_8_44_827_0, i_8_44_841_0,
    i_8_44_851_0, i_8_44_877_0, i_8_44_878_0, i_8_44_896_0, i_8_44_992_0,
    i_8_44_996_0, i_8_44_1012_0, i_8_44_1061_0, i_8_44_1066_0,
    i_8_44_1067_0, i_8_44_1084_0, i_8_44_1112_0, i_8_44_1115_0,
    i_8_44_1133_0, i_8_44_1148_0, i_8_44_1175_0, i_8_44_1246_0,
    i_8_44_1247_0, i_8_44_1261_0, i_8_44_1328_0, i_8_44_1346_0,
    i_8_44_1350_0, i_8_44_1417_0, i_8_44_1418_0, i_8_44_1451_0,
    i_8_44_1523_0, i_8_44_1525_0, i_8_44_1526_0, i_8_44_1550_0,
    i_8_44_1579_0, i_8_44_1613_0, i_8_44_1654_0, i_8_44_1667_0,
    i_8_44_1679_0, i_8_44_1681_0, i_8_44_1682_0, i_8_44_1729_0,
    i_8_44_1730_0, i_8_44_1733_0, i_8_44_1739_0, i_8_44_1747_0,
    i_8_44_1750_0, i_8_44_1753_0, i_8_44_1777_0, i_8_44_1778_0,
    i_8_44_1802_0, i_8_44_1808_0, i_8_44_1856_0, i_8_44_1867_0,
    i_8_44_1903_0, i_8_44_1904_0, i_8_44_1959_0, i_8_44_1990_0,
    i_8_44_1996_0, i_8_44_2011_0, i_8_44_2012_0, i_8_44_2077_0,
    i_8_44_2078_0, i_8_44_2153_0, i_8_44_2288_0,
    o_8_44_0_0  );
  input  i_8_44_11_0, i_8_44_23_0, i_8_44_28_0, i_8_44_95_0, i_8_44_97_0,
    i_8_44_157_0, i_8_44_158_0, i_8_44_202_0, i_8_44_203_0, i_8_44_209_0,
    i_8_44_223_0, i_8_44_244_0, i_8_44_245_0, i_8_44_248_0, i_8_44_266_0,
    i_8_44_326_0, i_8_44_348_0, i_8_44_355_0, i_8_44_364_0, i_8_44_380_0,
    i_8_44_437_0, i_8_44_452_0, i_8_44_483_0, i_8_44_484_0, i_8_44_498_0,
    i_8_44_508_0, i_8_44_526_0, i_8_44_536_0, i_8_44_551_0, i_8_44_554_0,
    i_8_44_556_0, i_8_44_557_0, i_8_44_587_0, i_8_44_626_0, i_8_44_628_0,
    i_8_44_657_0, i_8_44_779_0, i_8_44_793_0, i_8_44_827_0, i_8_44_841_0,
    i_8_44_851_0, i_8_44_877_0, i_8_44_878_0, i_8_44_896_0, i_8_44_992_0,
    i_8_44_996_0, i_8_44_1012_0, i_8_44_1061_0, i_8_44_1066_0,
    i_8_44_1067_0, i_8_44_1084_0, i_8_44_1112_0, i_8_44_1115_0,
    i_8_44_1133_0, i_8_44_1148_0, i_8_44_1175_0, i_8_44_1246_0,
    i_8_44_1247_0, i_8_44_1261_0, i_8_44_1328_0, i_8_44_1346_0,
    i_8_44_1350_0, i_8_44_1417_0, i_8_44_1418_0, i_8_44_1451_0,
    i_8_44_1523_0, i_8_44_1525_0, i_8_44_1526_0, i_8_44_1550_0,
    i_8_44_1579_0, i_8_44_1613_0, i_8_44_1654_0, i_8_44_1667_0,
    i_8_44_1679_0, i_8_44_1681_0, i_8_44_1682_0, i_8_44_1729_0,
    i_8_44_1730_0, i_8_44_1733_0, i_8_44_1739_0, i_8_44_1747_0,
    i_8_44_1750_0, i_8_44_1753_0, i_8_44_1777_0, i_8_44_1778_0,
    i_8_44_1802_0, i_8_44_1808_0, i_8_44_1856_0, i_8_44_1867_0,
    i_8_44_1903_0, i_8_44_1904_0, i_8_44_1959_0, i_8_44_1990_0,
    i_8_44_1996_0, i_8_44_2011_0, i_8_44_2012_0, i_8_44_2077_0,
    i_8_44_2078_0, i_8_44_2153_0, i_8_44_2288_0;
  output o_8_44_0_0;
  assign o_8_44_0_0 = 0;
endmodule



// Benchmark "kernel_8_45" written by ABC on Sun Jul 19 10:03:48 2020

module kernel_8_45 ( 
    i_8_45_41_0, i_8_45_44_0, i_8_45_77_0, i_8_45_112_0, i_8_45_114_0,
    i_8_45_115_0, i_8_45_116_0, i_8_45_141_0, i_8_45_182_0, i_8_45_317_0,
    i_8_45_319_0, i_8_45_320_0, i_8_45_322_0, i_8_45_381_0, i_8_45_382_0,
    i_8_45_392_0, i_8_45_398_0, i_8_45_489_0, i_8_45_537_0, i_8_45_547_0,
    i_8_45_553_0, i_8_45_556_0, i_8_45_568_0, i_8_45_571_0, i_8_45_580_0,
    i_8_45_589_0, i_8_45_598_0, i_8_45_612_0, i_8_45_634_0, i_8_45_640_0,
    i_8_45_652_0, i_8_45_655_0, i_8_45_657_0, i_8_45_670_0, i_8_45_680_0,
    i_8_45_716_0, i_8_45_732_0, i_8_45_859_0, i_8_45_860_0, i_8_45_895_0,
    i_8_45_966_0, i_8_45_970_0, i_8_45_975_0, i_8_45_1102_0, i_8_45_1111_0,
    i_8_45_1187_0, i_8_45_1192_0, i_8_45_1193_0, i_8_45_1201_0,
    i_8_45_1225_0, i_8_45_1228_0, i_8_45_1243_0, i_8_45_1296_0,
    i_8_45_1316_0, i_8_45_1326_0, i_8_45_1327_0, i_8_45_1363_0,
    i_8_45_1384_0, i_8_45_1407_0, i_8_45_1423_0, i_8_45_1427_0,
    i_8_45_1435_0, i_8_45_1462_0, i_8_45_1463_0, i_8_45_1467_0,
    i_8_45_1469_0, i_8_45_1477_0, i_8_45_1481_0, i_8_45_1516_0,
    i_8_45_1546_0, i_8_45_1573_0, i_8_45_1625_0, i_8_45_1630_0,
    i_8_45_1633_0, i_8_45_1694_0, i_8_45_1697_0, i_8_45_1750_0,
    i_8_45_1765_0, i_8_45_1768_0, i_8_45_1771_0, i_8_45_1776_0,
    i_8_45_1783_0, i_8_45_1840_0, i_8_45_1885_0, i_8_45_1894_0,
    i_8_45_1906_0, i_8_45_1912_0, i_8_45_1918_0, i_8_45_1949_0,
    i_8_45_1957_0, i_8_45_1972_0, i_8_45_1975_0, i_8_45_1979_0,
    i_8_45_1984_0, i_8_45_2041_0, i_8_45_2069_0, i_8_45_2095_0,
    i_8_45_2135_0, i_8_45_2192_0, i_8_45_2226_0,
    o_8_45_0_0  );
  input  i_8_45_41_0, i_8_45_44_0, i_8_45_77_0, i_8_45_112_0,
    i_8_45_114_0, i_8_45_115_0, i_8_45_116_0, i_8_45_141_0, i_8_45_182_0,
    i_8_45_317_0, i_8_45_319_0, i_8_45_320_0, i_8_45_322_0, i_8_45_381_0,
    i_8_45_382_0, i_8_45_392_0, i_8_45_398_0, i_8_45_489_0, i_8_45_537_0,
    i_8_45_547_0, i_8_45_553_0, i_8_45_556_0, i_8_45_568_0, i_8_45_571_0,
    i_8_45_580_0, i_8_45_589_0, i_8_45_598_0, i_8_45_612_0, i_8_45_634_0,
    i_8_45_640_0, i_8_45_652_0, i_8_45_655_0, i_8_45_657_0, i_8_45_670_0,
    i_8_45_680_0, i_8_45_716_0, i_8_45_732_0, i_8_45_859_0, i_8_45_860_0,
    i_8_45_895_0, i_8_45_966_0, i_8_45_970_0, i_8_45_975_0, i_8_45_1102_0,
    i_8_45_1111_0, i_8_45_1187_0, i_8_45_1192_0, i_8_45_1193_0,
    i_8_45_1201_0, i_8_45_1225_0, i_8_45_1228_0, i_8_45_1243_0,
    i_8_45_1296_0, i_8_45_1316_0, i_8_45_1326_0, i_8_45_1327_0,
    i_8_45_1363_0, i_8_45_1384_0, i_8_45_1407_0, i_8_45_1423_0,
    i_8_45_1427_0, i_8_45_1435_0, i_8_45_1462_0, i_8_45_1463_0,
    i_8_45_1467_0, i_8_45_1469_0, i_8_45_1477_0, i_8_45_1481_0,
    i_8_45_1516_0, i_8_45_1546_0, i_8_45_1573_0, i_8_45_1625_0,
    i_8_45_1630_0, i_8_45_1633_0, i_8_45_1694_0, i_8_45_1697_0,
    i_8_45_1750_0, i_8_45_1765_0, i_8_45_1768_0, i_8_45_1771_0,
    i_8_45_1776_0, i_8_45_1783_0, i_8_45_1840_0, i_8_45_1885_0,
    i_8_45_1894_0, i_8_45_1906_0, i_8_45_1912_0, i_8_45_1918_0,
    i_8_45_1949_0, i_8_45_1957_0, i_8_45_1972_0, i_8_45_1975_0,
    i_8_45_1979_0, i_8_45_1984_0, i_8_45_2041_0, i_8_45_2069_0,
    i_8_45_2095_0, i_8_45_2135_0, i_8_45_2192_0, i_8_45_2226_0;
  output o_8_45_0_0;
  assign o_8_45_0_0 = 0;
endmodule



// Benchmark "kernel_8_46" written by ABC on Sun Jul 19 10:03:49 2020

module kernel_8_46 ( 
    i_8_46_77_0, i_8_46_107_0, i_8_46_250_0, i_8_46_259_0, i_8_46_284_0,
    i_8_46_296_0, i_8_46_322_0, i_8_46_323_0, i_8_46_368_0, i_8_46_431_0,
    i_8_46_457_0, i_8_46_490_0, i_8_46_494_0, i_8_46_530_0, i_8_46_587_0,
    i_8_46_593_0, i_8_46_599_0, i_8_46_628_0, i_8_46_643_0, i_8_46_653_0,
    i_8_46_661_0, i_8_46_673_0, i_8_46_681_0, i_8_46_691_0, i_8_46_697_0,
    i_8_46_698_0, i_8_46_707_0, i_8_46_719_0, i_8_46_728_0, i_8_46_736_0,
    i_8_46_763_0, i_8_46_775_0, i_8_46_809_0, i_8_46_815_0, i_8_46_817_0,
    i_8_46_838_0, i_8_46_842_0, i_8_46_845_0, i_8_46_881_0, i_8_46_970_0,
    i_8_46_971_0, i_8_46_1031_0, i_8_46_1033_0, i_8_46_1078_0,
    i_8_46_1205_0, i_8_46_1227_0, i_8_46_1228_0, i_8_46_1232_0,
    i_8_46_1238_0, i_8_46_1239_0, i_8_46_1240_0, i_8_46_1265_0,
    i_8_46_1268_0, i_8_46_1321_0, i_8_46_1350_0, i_8_46_1358_0,
    i_8_46_1363_0, i_8_46_1391_0, i_8_46_1407_0, i_8_46_1408_0,
    i_8_46_1432_0, i_8_46_1436_0, i_8_46_1475_0, i_8_46_1492_0,
    i_8_46_1519_0, i_8_46_1520_0, i_8_46_1527_0, i_8_46_1528_0,
    i_8_46_1570_0, i_8_46_1574_0, i_8_46_1591_0, i_8_46_1592_0,
    i_8_46_1625_0, i_8_46_1642_0, i_8_46_1706_0, i_8_46_1744_0,
    i_8_46_1754_0, i_8_46_1768_0, i_8_46_1771_0, i_8_46_1813_0,
    i_8_46_1822_0, i_8_46_1823_0, i_8_46_1826_0, i_8_46_1858_0,
    i_8_46_1859_0, i_8_46_1880_0, i_8_46_1885_0, i_8_46_1889_0,
    i_8_46_1982_0, i_8_46_1994_0, i_8_46_2029_0, i_8_46_2032_0,
    i_8_46_2077_0, i_8_46_2132_0, i_8_46_2149_0, i_8_46_2156_0,
    i_8_46_2195_0, i_8_46_2224_0, i_8_46_2285_0, i_8_46_2290_0,
    o_8_46_0_0  );
  input  i_8_46_77_0, i_8_46_107_0, i_8_46_250_0, i_8_46_259_0,
    i_8_46_284_0, i_8_46_296_0, i_8_46_322_0, i_8_46_323_0, i_8_46_368_0,
    i_8_46_431_0, i_8_46_457_0, i_8_46_490_0, i_8_46_494_0, i_8_46_530_0,
    i_8_46_587_0, i_8_46_593_0, i_8_46_599_0, i_8_46_628_0, i_8_46_643_0,
    i_8_46_653_0, i_8_46_661_0, i_8_46_673_0, i_8_46_681_0, i_8_46_691_0,
    i_8_46_697_0, i_8_46_698_0, i_8_46_707_0, i_8_46_719_0, i_8_46_728_0,
    i_8_46_736_0, i_8_46_763_0, i_8_46_775_0, i_8_46_809_0, i_8_46_815_0,
    i_8_46_817_0, i_8_46_838_0, i_8_46_842_0, i_8_46_845_0, i_8_46_881_0,
    i_8_46_970_0, i_8_46_971_0, i_8_46_1031_0, i_8_46_1033_0,
    i_8_46_1078_0, i_8_46_1205_0, i_8_46_1227_0, i_8_46_1228_0,
    i_8_46_1232_0, i_8_46_1238_0, i_8_46_1239_0, i_8_46_1240_0,
    i_8_46_1265_0, i_8_46_1268_0, i_8_46_1321_0, i_8_46_1350_0,
    i_8_46_1358_0, i_8_46_1363_0, i_8_46_1391_0, i_8_46_1407_0,
    i_8_46_1408_0, i_8_46_1432_0, i_8_46_1436_0, i_8_46_1475_0,
    i_8_46_1492_0, i_8_46_1519_0, i_8_46_1520_0, i_8_46_1527_0,
    i_8_46_1528_0, i_8_46_1570_0, i_8_46_1574_0, i_8_46_1591_0,
    i_8_46_1592_0, i_8_46_1625_0, i_8_46_1642_0, i_8_46_1706_0,
    i_8_46_1744_0, i_8_46_1754_0, i_8_46_1768_0, i_8_46_1771_0,
    i_8_46_1813_0, i_8_46_1822_0, i_8_46_1823_0, i_8_46_1826_0,
    i_8_46_1858_0, i_8_46_1859_0, i_8_46_1880_0, i_8_46_1885_0,
    i_8_46_1889_0, i_8_46_1982_0, i_8_46_1994_0, i_8_46_2029_0,
    i_8_46_2032_0, i_8_46_2077_0, i_8_46_2132_0, i_8_46_2149_0,
    i_8_46_2156_0, i_8_46_2195_0, i_8_46_2224_0, i_8_46_2285_0,
    i_8_46_2290_0;
  output o_8_46_0_0;
  assign o_8_46_0_0 = 0;
endmodule



// Benchmark "kernel_8_47" written by ABC on Sun Jul 19 10:03:50 2020

module kernel_8_47 ( 
    i_8_47_7_0, i_8_47_24_0, i_8_47_70_0, i_8_47_79_0, i_8_47_88_0,
    i_8_47_129_0, i_8_47_151_0, i_8_47_195_0, i_8_47_212_0, i_8_47_214_0,
    i_8_47_247_0, i_8_47_250_0, i_8_47_277_0, i_8_47_313_0, i_8_47_358_0,
    i_8_47_376_0, i_8_47_396_0, i_8_47_450_0, i_8_47_467_0, i_8_47_503_0,
    i_8_47_528_0, i_8_47_529_0, i_8_47_570_0, i_8_47_597_0, i_8_47_602_0,
    i_8_47_609_0, i_8_47_615_0, i_8_47_636_0, i_8_47_654_0, i_8_47_655_0,
    i_8_47_672_0, i_8_47_681_0, i_8_47_695_0, i_8_47_700_0, i_8_47_708_0,
    i_8_47_709_0, i_8_47_735_0, i_8_47_751_0, i_8_47_754_0, i_8_47_762_0,
    i_8_47_772_0, i_8_47_835_0, i_8_47_862_0, i_8_47_1060_0, i_8_47_1061_0,
    i_8_47_1069_0, i_8_47_1137_0, i_8_47_1155_0, i_8_47_1177_0,
    i_8_47_1227_0, i_8_47_1257_0, i_8_47_1266_0, i_8_47_1267_0,
    i_8_47_1300_0, i_8_47_1303_0, i_8_47_1357_0, i_8_47_1384_0,
    i_8_47_1393_0, i_8_47_1410_0, i_8_47_1455_0, i_8_47_1496_0,
    i_8_47_1498_0, i_8_47_1501_0, i_8_47_1534_0, i_8_47_1551_0,
    i_8_47_1552_0, i_8_47_1599_0, i_8_47_1645_0, i_8_47_1648_0,
    i_8_47_1653_0, i_8_47_1654_0, i_8_47_1662_0, i_8_47_1690_0,
    i_8_47_1735_0, i_8_47_1750_0, i_8_47_1813_0, i_8_47_1851_0,
    i_8_47_1852_0, i_8_47_1870_0, i_8_47_1914_0, i_8_47_1915_0,
    i_8_47_1920_0, i_8_47_1921_0, i_8_47_1968_0, i_8_47_1969_0,
    i_8_47_1996_0, i_8_47_2013_0, i_8_47_2014_0, i_8_47_2068_0,
    i_8_47_2095_0, i_8_47_2112_0, i_8_47_2122_0, i_8_47_2172_0,
    i_8_47_2175_0, i_8_47_2184_0, i_8_47_2185_0, i_8_47_2217_0,
    i_8_47_2218_0, i_8_47_2272_0, i_8_47_2292_0,
    o_8_47_0_0  );
  input  i_8_47_7_0, i_8_47_24_0, i_8_47_70_0, i_8_47_79_0, i_8_47_88_0,
    i_8_47_129_0, i_8_47_151_0, i_8_47_195_0, i_8_47_212_0, i_8_47_214_0,
    i_8_47_247_0, i_8_47_250_0, i_8_47_277_0, i_8_47_313_0, i_8_47_358_0,
    i_8_47_376_0, i_8_47_396_0, i_8_47_450_0, i_8_47_467_0, i_8_47_503_0,
    i_8_47_528_0, i_8_47_529_0, i_8_47_570_0, i_8_47_597_0, i_8_47_602_0,
    i_8_47_609_0, i_8_47_615_0, i_8_47_636_0, i_8_47_654_0, i_8_47_655_0,
    i_8_47_672_0, i_8_47_681_0, i_8_47_695_0, i_8_47_700_0, i_8_47_708_0,
    i_8_47_709_0, i_8_47_735_0, i_8_47_751_0, i_8_47_754_0, i_8_47_762_0,
    i_8_47_772_0, i_8_47_835_0, i_8_47_862_0, i_8_47_1060_0, i_8_47_1061_0,
    i_8_47_1069_0, i_8_47_1137_0, i_8_47_1155_0, i_8_47_1177_0,
    i_8_47_1227_0, i_8_47_1257_0, i_8_47_1266_0, i_8_47_1267_0,
    i_8_47_1300_0, i_8_47_1303_0, i_8_47_1357_0, i_8_47_1384_0,
    i_8_47_1393_0, i_8_47_1410_0, i_8_47_1455_0, i_8_47_1496_0,
    i_8_47_1498_0, i_8_47_1501_0, i_8_47_1534_0, i_8_47_1551_0,
    i_8_47_1552_0, i_8_47_1599_0, i_8_47_1645_0, i_8_47_1648_0,
    i_8_47_1653_0, i_8_47_1654_0, i_8_47_1662_0, i_8_47_1690_0,
    i_8_47_1735_0, i_8_47_1750_0, i_8_47_1813_0, i_8_47_1851_0,
    i_8_47_1852_0, i_8_47_1870_0, i_8_47_1914_0, i_8_47_1915_0,
    i_8_47_1920_0, i_8_47_1921_0, i_8_47_1968_0, i_8_47_1969_0,
    i_8_47_1996_0, i_8_47_2013_0, i_8_47_2014_0, i_8_47_2068_0,
    i_8_47_2095_0, i_8_47_2112_0, i_8_47_2122_0, i_8_47_2172_0,
    i_8_47_2175_0, i_8_47_2184_0, i_8_47_2185_0, i_8_47_2217_0,
    i_8_47_2218_0, i_8_47_2272_0, i_8_47_2292_0;
  output o_8_47_0_0;
  assign o_8_47_0_0 = 0;
endmodule



// Benchmark "kernel_8_48" written by ABC on Sun Jul 19 10:03:51 2020

module kernel_8_48 ( 
    i_8_48_22_0, i_8_48_82_0, i_8_48_104_0, i_8_48_263_0, i_8_48_292_0,
    i_8_48_302_0, i_8_48_303_0, i_8_48_346_0, i_8_48_347_0, i_8_48_377_0,
    i_8_48_418_0, i_8_48_463_0, i_8_48_464_0, i_8_48_476_0, i_8_48_482_0,
    i_8_48_500_0, i_8_48_503_0, i_8_48_547_0, i_8_48_554_0, i_8_48_556_0,
    i_8_48_557_0, i_8_48_589_0, i_8_48_593_0, i_8_48_597_0, i_8_48_599_0,
    i_8_48_625_0, i_8_48_674_0, i_8_48_716_0, i_8_48_796_0, i_8_48_827_0,
    i_8_48_892_0, i_8_48_895_0, i_8_48_1030_0, i_8_48_1114_0,
    i_8_48_1115_0, i_8_48_1121_0, i_8_48_1129_0, i_8_48_1130_0,
    i_8_48_1258_0, i_8_48_1271_0, i_8_48_1274_0, i_8_48_1283_0,
    i_8_48_1286_0, i_8_48_1307_0, i_8_48_1314_0, i_8_48_1323_0,
    i_8_48_1347_0, i_8_48_1350_0, i_8_48_1432_0, i_8_48_1453_0,
    i_8_48_1454_0, i_8_48_1470_0, i_8_48_1471_0, i_8_48_1472_0,
    i_8_48_1535_0, i_8_48_1587_0, i_8_48_1597_0, i_8_48_1604_0,
    i_8_48_1681_0, i_8_48_1706_0, i_8_48_1711_0, i_8_48_1714_0,
    i_8_48_1749_0, i_8_48_1763_0, i_8_48_1787_0, i_8_48_1790_0,
    i_8_48_1802_0, i_8_48_1807_0, i_8_48_1841_0, i_8_48_1854_0,
    i_8_48_1855_0, i_8_48_1867_0, i_8_48_1871_0, i_8_48_1895_0,
    i_8_48_1918_0, i_8_48_1919_0, i_8_48_1927_0, i_8_48_1948_0,
    i_8_48_1970_0, i_8_48_2033_0, i_8_48_2050_0, i_8_48_2051_0,
    i_8_48_2110_0, i_8_48_2111_0, i_8_48_2129_0, i_8_48_2134_0,
    i_8_48_2140_0, i_8_48_2183_0, i_8_48_2191_0, i_8_48_2192_0,
    i_8_48_2214_0, i_8_48_2215_0, i_8_48_2216_0, i_8_48_2230_0,
    i_8_48_2234_0, i_8_48_2247_0, i_8_48_2261_0, i_8_48_2273_0,
    i_8_48_2276_0, i_8_48_2290_0,
    o_8_48_0_0  );
  input  i_8_48_22_0, i_8_48_82_0, i_8_48_104_0, i_8_48_263_0,
    i_8_48_292_0, i_8_48_302_0, i_8_48_303_0, i_8_48_346_0, i_8_48_347_0,
    i_8_48_377_0, i_8_48_418_0, i_8_48_463_0, i_8_48_464_0, i_8_48_476_0,
    i_8_48_482_0, i_8_48_500_0, i_8_48_503_0, i_8_48_547_0, i_8_48_554_0,
    i_8_48_556_0, i_8_48_557_0, i_8_48_589_0, i_8_48_593_0, i_8_48_597_0,
    i_8_48_599_0, i_8_48_625_0, i_8_48_674_0, i_8_48_716_0, i_8_48_796_0,
    i_8_48_827_0, i_8_48_892_0, i_8_48_895_0, i_8_48_1030_0, i_8_48_1114_0,
    i_8_48_1115_0, i_8_48_1121_0, i_8_48_1129_0, i_8_48_1130_0,
    i_8_48_1258_0, i_8_48_1271_0, i_8_48_1274_0, i_8_48_1283_0,
    i_8_48_1286_0, i_8_48_1307_0, i_8_48_1314_0, i_8_48_1323_0,
    i_8_48_1347_0, i_8_48_1350_0, i_8_48_1432_0, i_8_48_1453_0,
    i_8_48_1454_0, i_8_48_1470_0, i_8_48_1471_0, i_8_48_1472_0,
    i_8_48_1535_0, i_8_48_1587_0, i_8_48_1597_0, i_8_48_1604_0,
    i_8_48_1681_0, i_8_48_1706_0, i_8_48_1711_0, i_8_48_1714_0,
    i_8_48_1749_0, i_8_48_1763_0, i_8_48_1787_0, i_8_48_1790_0,
    i_8_48_1802_0, i_8_48_1807_0, i_8_48_1841_0, i_8_48_1854_0,
    i_8_48_1855_0, i_8_48_1867_0, i_8_48_1871_0, i_8_48_1895_0,
    i_8_48_1918_0, i_8_48_1919_0, i_8_48_1927_0, i_8_48_1948_0,
    i_8_48_1970_0, i_8_48_2033_0, i_8_48_2050_0, i_8_48_2051_0,
    i_8_48_2110_0, i_8_48_2111_0, i_8_48_2129_0, i_8_48_2134_0,
    i_8_48_2140_0, i_8_48_2183_0, i_8_48_2191_0, i_8_48_2192_0,
    i_8_48_2214_0, i_8_48_2215_0, i_8_48_2216_0, i_8_48_2230_0,
    i_8_48_2234_0, i_8_48_2247_0, i_8_48_2261_0, i_8_48_2273_0,
    i_8_48_2276_0, i_8_48_2290_0;
  output o_8_48_0_0;
  assign o_8_48_0_0 = 0;
endmodule



// Benchmark "kernel_8_49" written by ABC on Sun Jul 19 10:03:52 2020

module kernel_8_49 ( 
    i_8_49_22_0, i_8_49_39_0, i_8_49_53_0, i_8_49_126_0, i_8_49_147_0,
    i_8_49_318_0, i_8_49_319_0, i_8_49_320_0, i_8_49_321_0, i_8_49_322_0,
    i_8_49_323_0, i_8_49_336_0, i_8_49_342_0, i_8_49_396_0, i_8_49_397_0,
    i_8_49_424_0, i_8_49_425_0, i_8_49_427_0, i_8_49_439_0, i_8_49_547_0,
    i_8_49_552_0, i_8_49_561_0, i_8_49_571_0, i_8_49_580_0, i_8_49_588_0,
    i_8_49_589_0, i_8_49_596_0, i_8_49_603_0, i_8_49_604_0, i_8_49_610_0,
    i_8_49_611_0, i_8_49_658_0, i_8_49_676_0, i_8_49_695_0, i_8_49_750_0,
    i_8_49_766_0, i_8_49_777_0, i_8_49_841_0, i_8_49_865_0, i_8_49_875_0,
    i_8_49_894_0, i_8_49_969_0, i_8_49_976_0, i_8_49_1022_0, i_8_49_1100_0,
    i_8_49_1102_0, i_8_49_1103_0, i_8_49_1110_0, i_8_49_1180_0,
    i_8_49_1236_0, i_8_49_1237_0, i_8_49_1243_0, i_8_49_1264_0,
    i_8_49_1286_0, i_8_49_1327_0, i_8_49_1357_0, i_8_49_1362_0,
    i_8_49_1363_0, i_8_49_1380_0, i_8_49_1381_0, i_8_49_1399_0,
    i_8_49_1431_0, i_8_49_1432_0, i_8_49_1461_0, i_8_49_1463_0,
    i_8_49_1477_0, i_8_49_1514_0, i_8_49_1526_0, i_8_49_1536_0,
    i_8_49_1573_0, i_8_49_1605_0, i_8_49_1606_0, i_8_49_1626_0,
    i_8_49_1632_0, i_8_49_1681_0, i_8_49_1707_0, i_8_49_1735_0,
    i_8_49_1749_0, i_8_49_1750_0, i_8_49_1760_0, i_8_49_1766_0,
    i_8_49_1767_0, i_8_49_1781_0, i_8_49_1866_0, i_8_49_1884_0,
    i_8_49_1929_0, i_8_49_1930_0, i_8_49_1937_0, i_8_49_1957_0,
    i_8_49_1974_0, i_8_49_1975_0, i_8_49_1996_0, i_8_49_2091_0,
    i_8_49_2119_0, i_8_49_2143_0, i_8_49_2191_0, i_8_49_2244_0,
    i_8_49_2245_0, i_8_49_2246_0, i_8_49_2271_0,
    o_8_49_0_0  );
  input  i_8_49_22_0, i_8_49_39_0, i_8_49_53_0, i_8_49_126_0,
    i_8_49_147_0, i_8_49_318_0, i_8_49_319_0, i_8_49_320_0, i_8_49_321_0,
    i_8_49_322_0, i_8_49_323_0, i_8_49_336_0, i_8_49_342_0, i_8_49_396_0,
    i_8_49_397_0, i_8_49_424_0, i_8_49_425_0, i_8_49_427_0, i_8_49_439_0,
    i_8_49_547_0, i_8_49_552_0, i_8_49_561_0, i_8_49_571_0, i_8_49_580_0,
    i_8_49_588_0, i_8_49_589_0, i_8_49_596_0, i_8_49_603_0, i_8_49_604_0,
    i_8_49_610_0, i_8_49_611_0, i_8_49_658_0, i_8_49_676_0, i_8_49_695_0,
    i_8_49_750_0, i_8_49_766_0, i_8_49_777_0, i_8_49_841_0, i_8_49_865_0,
    i_8_49_875_0, i_8_49_894_0, i_8_49_969_0, i_8_49_976_0, i_8_49_1022_0,
    i_8_49_1100_0, i_8_49_1102_0, i_8_49_1103_0, i_8_49_1110_0,
    i_8_49_1180_0, i_8_49_1236_0, i_8_49_1237_0, i_8_49_1243_0,
    i_8_49_1264_0, i_8_49_1286_0, i_8_49_1327_0, i_8_49_1357_0,
    i_8_49_1362_0, i_8_49_1363_0, i_8_49_1380_0, i_8_49_1381_0,
    i_8_49_1399_0, i_8_49_1431_0, i_8_49_1432_0, i_8_49_1461_0,
    i_8_49_1463_0, i_8_49_1477_0, i_8_49_1514_0, i_8_49_1526_0,
    i_8_49_1536_0, i_8_49_1573_0, i_8_49_1605_0, i_8_49_1606_0,
    i_8_49_1626_0, i_8_49_1632_0, i_8_49_1681_0, i_8_49_1707_0,
    i_8_49_1735_0, i_8_49_1749_0, i_8_49_1750_0, i_8_49_1760_0,
    i_8_49_1766_0, i_8_49_1767_0, i_8_49_1781_0, i_8_49_1866_0,
    i_8_49_1884_0, i_8_49_1929_0, i_8_49_1930_0, i_8_49_1937_0,
    i_8_49_1957_0, i_8_49_1974_0, i_8_49_1975_0, i_8_49_1996_0,
    i_8_49_2091_0, i_8_49_2119_0, i_8_49_2143_0, i_8_49_2191_0,
    i_8_49_2244_0, i_8_49_2245_0, i_8_49_2246_0, i_8_49_2271_0;
  output o_8_49_0_0;
  assign o_8_49_0_0 = 0;
endmodule



// Benchmark "kernel_8_50" written by ABC on Sun Jul 19 10:03:53 2020

module kernel_8_50 ( 
    i_8_50_14_0, i_8_50_18_0, i_8_50_85_0, i_8_50_93_0, i_8_50_117_0,
    i_8_50_151_0, i_8_50_192_0, i_8_50_193_0, i_8_50_258_0, i_8_50_259_0,
    i_8_50_273_0, i_8_50_325_0, i_8_50_360_0, i_8_50_363_0, i_8_50_364_0,
    i_8_50_423_0, i_8_50_426_0, i_8_50_427_0, i_8_50_447_0, i_8_50_468_0,
    i_8_50_526_0, i_8_50_529_0, i_8_50_554_0, i_8_50_567_0, i_8_50_568_0,
    i_8_50_615_0, i_8_50_622_0, i_8_50_630_0, i_8_50_652_0, i_8_50_684_0,
    i_8_50_694_0, i_8_50_699_0, i_8_50_707_0, i_8_50_832_0, i_8_50_837_0,
    i_8_50_865_0, i_8_50_873_0, i_8_50_874_0, i_8_50_876_0, i_8_50_882_0,
    i_8_50_981_0, i_8_50_1023_0, i_8_50_1030_0, i_8_50_1036_0,
    i_8_50_1051_0, i_8_50_1089_0, i_8_50_1092_0, i_8_50_1102_0,
    i_8_50_1137_0, i_8_50_1138_0, i_8_50_1147_0, i_8_50_1237_0,
    i_8_50_1267_0, i_8_50_1314_0, i_8_50_1332_0, i_8_50_1349_0,
    i_8_50_1407_0, i_8_50_1455_0, i_8_50_1486_0, i_8_50_1597_0,
    i_8_50_1602_0, i_8_50_1605_0, i_8_50_1620_0, i_8_50_1638_0,
    i_8_50_1650_0, i_8_50_1696_0, i_8_50_1702_0, i_8_50_1765_0,
    i_8_50_1768_0, i_8_50_1774_0, i_8_50_1804_0, i_8_50_1807_0,
    i_8_50_1810_0, i_8_50_1818_0, i_8_50_1821_0, i_8_50_1857_0,
    i_8_50_1881_0, i_8_50_1882_0, i_8_50_1884_0, i_8_50_1893_0,
    i_8_50_1929_0, i_8_50_1938_0, i_8_50_2007_0, i_8_50_2044_0,
    i_8_50_2055_0, i_8_50_2066_0, i_8_50_2070_0, i_8_50_2079_0,
    i_8_50_2092_0, i_8_50_2097_0, i_8_50_2114_0, i_8_50_2124_0,
    i_8_50_2144_0, i_8_50_2146_0, i_8_50_2147_0, i_8_50_2152_0,
    i_8_50_2170_0, i_8_50_2241_0, i_8_50_2246_0, i_8_50_2294_0,
    o_8_50_0_0  );
  input  i_8_50_14_0, i_8_50_18_0, i_8_50_85_0, i_8_50_93_0,
    i_8_50_117_0, i_8_50_151_0, i_8_50_192_0, i_8_50_193_0, i_8_50_258_0,
    i_8_50_259_0, i_8_50_273_0, i_8_50_325_0, i_8_50_360_0, i_8_50_363_0,
    i_8_50_364_0, i_8_50_423_0, i_8_50_426_0, i_8_50_427_0, i_8_50_447_0,
    i_8_50_468_0, i_8_50_526_0, i_8_50_529_0, i_8_50_554_0, i_8_50_567_0,
    i_8_50_568_0, i_8_50_615_0, i_8_50_622_0, i_8_50_630_0, i_8_50_652_0,
    i_8_50_684_0, i_8_50_694_0, i_8_50_699_0, i_8_50_707_0, i_8_50_832_0,
    i_8_50_837_0, i_8_50_865_0, i_8_50_873_0, i_8_50_874_0, i_8_50_876_0,
    i_8_50_882_0, i_8_50_981_0, i_8_50_1023_0, i_8_50_1030_0,
    i_8_50_1036_0, i_8_50_1051_0, i_8_50_1089_0, i_8_50_1092_0,
    i_8_50_1102_0, i_8_50_1137_0, i_8_50_1138_0, i_8_50_1147_0,
    i_8_50_1237_0, i_8_50_1267_0, i_8_50_1314_0, i_8_50_1332_0,
    i_8_50_1349_0, i_8_50_1407_0, i_8_50_1455_0, i_8_50_1486_0,
    i_8_50_1597_0, i_8_50_1602_0, i_8_50_1605_0, i_8_50_1620_0,
    i_8_50_1638_0, i_8_50_1650_0, i_8_50_1696_0, i_8_50_1702_0,
    i_8_50_1765_0, i_8_50_1768_0, i_8_50_1774_0, i_8_50_1804_0,
    i_8_50_1807_0, i_8_50_1810_0, i_8_50_1818_0, i_8_50_1821_0,
    i_8_50_1857_0, i_8_50_1881_0, i_8_50_1882_0, i_8_50_1884_0,
    i_8_50_1893_0, i_8_50_1929_0, i_8_50_1938_0, i_8_50_2007_0,
    i_8_50_2044_0, i_8_50_2055_0, i_8_50_2066_0, i_8_50_2070_0,
    i_8_50_2079_0, i_8_50_2092_0, i_8_50_2097_0, i_8_50_2114_0,
    i_8_50_2124_0, i_8_50_2144_0, i_8_50_2146_0, i_8_50_2147_0,
    i_8_50_2152_0, i_8_50_2170_0, i_8_50_2241_0, i_8_50_2246_0,
    i_8_50_2294_0;
  output o_8_50_0_0;
  assign o_8_50_0_0 = 0;
endmodule



// Benchmark "kernel_8_51" written by ABC on Sun Jul 19 10:03:54 2020

module kernel_8_51 ( 
    i_8_51_26_0, i_8_51_69_0, i_8_51_88_0, i_8_51_176_0, i_8_51_193_0,
    i_8_51_197_0, i_8_51_204_0, i_8_51_205_0, i_8_51_206_0, i_8_51_214_0,
    i_8_51_215_0, i_8_51_278_0, i_8_51_345_0, i_8_51_358_0, i_8_51_359_0,
    i_8_51_364_0, i_8_51_367_0, i_8_51_377_0, i_8_51_379_0, i_8_51_383_0,
    i_8_51_384_0, i_8_51_398_0, i_8_51_449_0, i_8_51_458_0, i_8_51_475_0,
    i_8_51_500_0, i_8_51_503_0, i_8_51_520_0, i_8_51_521_0, i_8_51_530_0,
    i_8_51_575_0, i_8_51_592_0, i_8_51_593_0, i_8_51_619_0, i_8_51_634_0,
    i_8_51_673_0, i_8_51_674_0, i_8_51_692_0, i_8_51_719_0, i_8_51_772_0,
    i_8_51_773_0, i_8_51_818_0, i_8_51_826_0, i_8_51_833_0, i_8_51_881_0,
    i_8_51_890_0, i_8_51_959_0, i_8_51_995_0, i_8_51_1035_0, i_8_51_1043_0,
    i_8_51_1079_0, i_8_51_1087_0, i_8_51_1196_0, i_8_51_1232_0,
    i_8_51_1261_0, i_8_51_1264_0, i_8_51_1285_0, i_8_51_1294_0,
    i_8_51_1300_0, i_8_51_1304_0, i_8_51_1312_0, i_8_51_1353_0,
    i_8_51_1410_0, i_8_51_1439_0, i_8_51_1473_0, i_8_51_1501_0,
    i_8_51_1504_0, i_8_51_1544_0, i_8_51_1565_0, i_8_51_1646_0,
    i_8_51_1672_0, i_8_51_1673_0, i_8_51_1691_0, i_8_51_1699_0,
    i_8_51_1700_0, i_8_51_1717_0, i_8_51_1718_0, i_8_51_1722_0,
    i_8_51_1735_0, i_8_51_1771_0, i_8_51_1772_0, i_8_51_1789_0,
    i_8_51_1807_0, i_8_51_1816_0, i_8_51_1844_0, i_8_51_1853_0,
    i_8_51_1880_0, i_8_51_1886_0, i_8_51_1887_0, i_8_51_1948_0,
    i_8_51_2014_0, i_8_51_2015_0, i_8_51_2074_0, i_8_51_2152_0,
    i_8_51_2186_0, i_8_51_2194_0, i_8_51_2195_0, i_8_51_2218_0,
    i_8_51_2249_0, i_8_51_2267_0,
    o_8_51_0_0  );
  input  i_8_51_26_0, i_8_51_69_0, i_8_51_88_0, i_8_51_176_0,
    i_8_51_193_0, i_8_51_197_0, i_8_51_204_0, i_8_51_205_0, i_8_51_206_0,
    i_8_51_214_0, i_8_51_215_0, i_8_51_278_0, i_8_51_345_0, i_8_51_358_0,
    i_8_51_359_0, i_8_51_364_0, i_8_51_367_0, i_8_51_377_0, i_8_51_379_0,
    i_8_51_383_0, i_8_51_384_0, i_8_51_398_0, i_8_51_449_0, i_8_51_458_0,
    i_8_51_475_0, i_8_51_500_0, i_8_51_503_0, i_8_51_520_0, i_8_51_521_0,
    i_8_51_530_0, i_8_51_575_0, i_8_51_592_0, i_8_51_593_0, i_8_51_619_0,
    i_8_51_634_0, i_8_51_673_0, i_8_51_674_0, i_8_51_692_0, i_8_51_719_0,
    i_8_51_772_0, i_8_51_773_0, i_8_51_818_0, i_8_51_826_0, i_8_51_833_0,
    i_8_51_881_0, i_8_51_890_0, i_8_51_959_0, i_8_51_995_0, i_8_51_1035_0,
    i_8_51_1043_0, i_8_51_1079_0, i_8_51_1087_0, i_8_51_1196_0,
    i_8_51_1232_0, i_8_51_1261_0, i_8_51_1264_0, i_8_51_1285_0,
    i_8_51_1294_0, i_8_51_1300_0, i_8_51_1304_0, i_8_51_1312_0,
    i_8_51_1353_0, i_8_51_1410_0, i_8_51_1439_0, i_8_51_1473_0,
    i_8_51_1501_0, i_8_51_1504_0, i_8_51_1544_0, i_8_51_1565_0,
    i_8_51_1646_0, i_8_51_1672_0, i_8_51_1673_0, i_8_51_1691_0,
    i_8_51_1699_0, i_8_51_1700_0, i_8_51_1717_0, i_8_51_1718_0,
    i_8_51_1722_0, i_8_51_1735_0, i_8_51_1771_0, i_8_51_1772_0,
    i_8_51_1789_0, i_8_51_1807_0, i_8_51_1816_0, i_8_51_1844_0,
    i_8_51_1853_0, i_8_51_1880_0, i_8_51_1886_0, i_8_51_1887_0,
    i_8_51_1948_0, i_8_51_2014_0, i_8_51_2015_0, i_8_51_2074_0,
    i_8_51_2152_0, i_8_51_2186_0, i_8_51_2194_0, i_8_51_2195_0,
    i_8_51_2218_0, i_8_51_2249_0, i_8_51_2267_0;
  output o_8_51_0_0;
  assign o_8_51_0_0 = ~((~i_8_51_26_0 & ((~i_8_51_206_0 & ~i_8_51_692_0 & ~i_8_51_1087_0 & ~i_8_51_1691_0 & ~i_8_51_1735_0) | (~i_8_51_176_0 & ~i_8_51_278_0 & ~i_8_51_345_0 & ~i_8_51_359_0 & ~i_8_51_772_0 & ~i_8_51_818_0 & ~i_8_51_1717_0 & ~i_8_51_2186_0))) | (~i_8_51_214_0 & ((~i_8_51_197_0 & ~i_8_51_359_0 & i_8_51_719_0 & ~i_8_51_1294_0 & ~i_8_51_1300_0 & ~i_8_51_1844_0) | (~i_8_51_204_0 & ~i_8_51_1673_0 & i_8_51_2249_0))) | (~i_8_51_204_0 & ((~i_8_51_206_0 & ~i_8_51_503_0 & ~i_8_51_1232_0 & ~i_8_51_1816_0) | (~i_8_51_176_0 & ~i_8_51_383_0 & ~i_8_51_384_0 & ~i_8_51_673_0 & ~i_8_51_674_0 & i_8_51_995_0 & ~i_8_51_1264_0 & ~i_8_51_1501_0 & ~i_8_51_1948_0))) | (~i_8_51_215_0 & ((~i_8_51_358_0 & ~i_8_51_449_0 & ~i_8_51_818_0 & ~i_8_51_1087_0 & ~i_8_51_1261_0 & ~i_8_51_1646_0) | (~i_8_51_379_0 & ~i_8_51_1501_0 & ~i_8_51_1853_0 & ~i_8_51_2015_0))) | (~i_8_51_278_0 & ((~i_8_51_205_0 & ~i_8_51_449_0 & ~i_8_51_1087_0 & ~i_8_51_1886_0) | (~i_8_51_521_0 & ~i_8_51_818_0 & ~i_8_51_1261_0 & ~i_8_51_1700_0 & ~i_8_51_1735_0 & ~i_8_51_2267_0))) | (~i_8_51_377_0 & ~i_8_51_1880_0 & ((i_8_51_383_0 & ~i_8_51_1035_0 & ~i_8_51_1294_0 & ~i_8_51_1646_0) | (~i_8_51_818_0 & ~i_8_51_1312_0 & ~i_8_51_1691_0 & i_8_51_2014_0 & ~i_8_51_2218_0))) | (~i_8_51_2014_0 & ((~i_8_51_359_0 & ~i_8_51_449_0 & ~i_8_51_773_0 & ~i_8_51_1079_0) | (i_8_51_206_0 & ~i_8_51_1565_0 & ~i_8_51_1673_0 & ~i_8_51_1718_0 & i_8_51_2218_0))) | (i_8_51_449_0 & ~i_8_51_503_0 & ~i_8_51_692_0 & ~i_8_51_1501_0 & ~i_8_51_1504_0 & i_8_51_1807_0 & ~i_8_51_2152_0 & ~i_8_51_2186_0));
endmodule



// Benchmark "kernel_8_52" written by ABC on Sun Jul 19 10:03:55 2020

module kernel_8_52 ( 
    i_8_52_3_0, i_8_52_17_0, i_8_52_20_0, i_8_52_21_0, i_8_52_29_0,
    i_8_52_31_0, i_8_52_37_0, i_8_52_53_0, i_8_52_87_0, i_8_52_88_0,
    i_8_52_104_0, i_8_52_263_0, i_8_52_290_0, i_8_52_307_0, i_8_52_316_0,
    i_8_52_335_0, i_8_52_348_0, i_8_52_363_0, i_8_52_379_0, i_8_52_380_0,
    i_8_52_402_0, i_8_52_417_0, i_8_52_483_0, i_8_52_489_0, i_8_52_528_0,
    i_8_52_529_0, i_8_52_586_0, i_8_52_587_0, i_8_52_605_0, i_8_52_621_0,
    i_8_52_634_0, i_8_52_649_0, i_8_52_660_0, i_8_52_675_0, i_8_52_693_0,
    i_8_52_703_0, i_8_52_721_0, i_8_52_730_0, i_8_52_791_0, i_8_52_824_0,
    i_8_52_841_0, i_8_52_843_0, i_8_52_874_0, i_8_52_888_0, i_8_52_918_0,
    i_8_52_923_0, i_8_52_950_0, i_8_52_968_0, i_8_52_974_0, i_8_52_1078_0,
    i_8_52_1120_0, i_8_52_1180_0, i_8_52_1222_0, i_8_52_1264_0,
    i_8_52_1276_0, i_8_52_1284_0, i_8_52_1290_0, i_8_52_1324_0,
    i_8_52_1334_0, i_8_52_1440_0, i_8_52_1469_0, i_8_52_1474_0,
    i_8_52_1504_0, i_8_52_1585_0, i_8_52_1680_0, i_8_52_1682_0,
    i_8_52_1698_0, i_8_52_1743_0, i_8_52_1745_0, i_8_52_1748_0,
    i_8_52_1752_0, i_8_52_1760_0, i_8_52_1764_0, i_8_52_1768_0,
    i_8_52_1773_0, i_8_52_1796_0, i_8_52_1817_0, i_8_52_1820_0,
    i_8_52_1854_0, i_8_52_1861_0, i_8_52_1901_0, i_8_52_1904_0,
    i_8_52_1981_0, i_8_52_1993_0, i_8_52_1999_0, i_8_52_2026_0,
    i_8_52_2071_0, i_8_52_2105_0, i_8_52_2117_0, i_8_52_2130_0,
    i_8_52_2139_0, i_8_52_2140_0, i_8_52_2141_0, i_8_52_2143_0,
    i_8_52_2187_0, i_8_52_2188_0, i_8_52_2234_0, i_8_52_2243_0,
    i_8_52_2287_0, i_8_52_2301_0,
    o_8_52_0_0  );
  input  i_8_52_3_0, i_8_52_17_0, i_8_52_20_0, i_8_52_21_0, i_8_52_29_0,
    i_8_52_31_0, i_8_52_37_0, i_8_52_53_0, i_8_52_87_0, i_8_52_88_0,
    i_8_52_104_0, i_8_52_263_0, i_8_52_290_0, i_8_52_307_0, i_8_52_316_0,
    i_8_52_335_0, i_8_52_348_0, i_8_52_363_0, i_8_52_379_0, i_8_52_380_0,
    i_8_52_402_0, i_8_52_417_0, i_8_52_483_0, i_8_52_489_0, i_8_52_528_0,
    i_8_52_529_0, i_8_52_586_0, i_8_52_587_0, i_8_52_605_0, i_8_52_621_0,
    i_8_52_634_0, i_8_52_649_0, i_8_52_660_0, i_8_52_675_0, i_8_52_693_0,
    i_8_52_703_0, i_8_52_721_0, i_8_52_730_0, i_8_52_791_0, i_8_52_824_0,
    i_8_52_841_0, i_8_52_843_0, i_8_52_874_0, i_8_52_888_0, i_8_52_918_0,
    i_8_52_923_0, i_8_52_950_0, i_8_52_968_0, i_8_52_974_0, i_8_52_1078_0,
    i_8_52_1120_0, i_8_52_1180_0, i_8_52_1222_0, i_8_52_1264_0,
    i_8_52_1276_0, i_8_52_1284_0, i_8_52_1290_0, i_8_52_1324_0,
    i_8_52_1334_0, i_8_52_1440_0, i_8_52_1469_0, i_8_52_1474_0,
    i_8_52_1504_0, i_8_52_1585_0, i_8_52_1680_0, i_8_52_1682_0,
    i_8_52_1698_0, i_8_52_1743_0, i_8_52_1745_0, i_8_52_1748_0,
    i_8_52_1752_0, i_8_52_1760_0, i_8_52_1764_0, i_8_52_1768_0,
    i_8_52_1773_0, i_8_52_1796_0, i_8_52_1817_0, i_8_52_1820_0,
    i_8_52_1854_0, i_8_52_1861_0, i_8_52_1901_0, i_8_52_1904_0,
    i_8_52_1981_0, i_8_52_1993_0, i_8_52_1999_0, i_8_52_2026_0,
    i_8_52_2071_0, i_8_52_2105_0, i_8_52_2117_0, i_8_52_2130_0,
    i_8_52_2139_0, i_8_52_2140_0, i_8_52_2141_0, i_8_52_2143_0,
    i_8_52_2187_0, i_8_52_2188_0, i_8_52_2234_0, i_8_52_2243_0,
    i_8_52_2287_0, i_8_52_2301_0;
  output o_8_52_0_0;
  assign o_8_52_0_0 = 0;
endmodule



// Benchmark "kernel_8_53" written by ABC on Sun Jul 19 10:03:56 2020

module kernel_8_53 ( 
    i_8_53_32_0, i_8_53_37_0, i_8_53_41_0, i_8_53_43_0, i_8_53_51_0,
    i_8_53_57_0, i_8_53_64_0, i_8_53_67_0, i_8_53_120_0, i_8_53_160_0,
    i_8_53_172_0, i_8_53_205_0, i_8_53_228_0, i_8_53_229_0, i_8_53_230_0,
    i_8_53_325_0, i_8_53_326_0, i_8_53_329_0, i_8_53_334_0, i_8_53_352_0,
    i_8_53_392_0, i_8_53_400_0, i_8_53_401_0, i_8_53_417_0, i_8_53_462_0,
    i_8_53_502_0, i_8_53_552_0, i_8_53_555_0, i_8_53_556_0, i_8_53_557_0,
    i_8_53_697_0, i_8_53_698_0, i_8_53_699_0, i_8_53_700_0, i_8_53_701_0,
    i_8_53_748_0, i_8_53_838_0, i_8_53_839_0, i_8_53_850_0, i_8_53_883_0,
    i_8_53_885_0, i_8_53_886_0, i_8_53_889_0, i_8_53_995_0, i_8_53_1012_0,
    i_8_53_1128_0, i_8_53_1129_0, i_8_53_1131_0, i_8_53_1133_0,
    i_8_53_1156_0, i_8_53_1158_0, i_8_53_1202_0, i_8_53_1203_0,
    i_8_53_1205_0, i_8_53_1236_0, i_8_53_1322_0, i_8_53_1328_0,
    i_8_53_1331_0, i_8_53_1381_0, i_8_53_1427_0, i_8_53_1489_0,
    i_8_53_1551_0, i_8_53_1552_0, i_8_53_1555_0, i_8_53_1682_0,
    i_8_53_1705_0, i_8_53_1709_0, i_8_53_1726_0, i_8_53_1732_0,
    i_8_53_1749_0, i_8_53_1751_0, i_8_53_1753_0, i_8_53_1797_0,
    i_8_53_1806_0, i_8_53_1807_0, i_8_53_1841_0, i_8_53_1912_0,
    i_8_53_1913_0, i_8_53_1914_0, i_8_53_1915_0, i_8_53_1916_0,
    i_8_53_1936_0, i_8_53_1939_0, i_8_53_1982_0, i_8_53_1983_0,
    i_8_53_1985_0, i_8_53_1992_0, i_8_53_1999_0, i_8_53_2017_0,
    i_8_53_2055_0, i_8_53_2057_0, i_8_53_2058_0, i_8_53_2059_0,
    i_8_53_2144_0, i_8_53_2146_0, i_8_53_2147_0, i_8_53_2154_0,
    i_8_53_2159_0, i_8_53_2177_0, i_8_53_2272_0,
    o_8_53_0_0  );
  input  i_8_53_32_0, i_8_53_37_0, i_8_53_41_0, i_8_53_43_0, i_8_53_51_0,
    i_8_53_57_0, i_8_53_64_0, i_8_53_67_0, i_8_53_120_0, i_8_53_160_0,
    i_8_53_172_0, i_8_53_205_0, i_8_53_228_0, i_8_53_229_0, i_8_53_230_0,
    i_8_53_325_0, i_8_53_326_0, i_8_53_329_0, i_8_53_334_0, i_8_53_352_0,
    i_8_53_392_0, i_8_53_400_0, i_8_53_401_0, i_8_53_417_0, i_8_53_462_0,
    i_8_53_502_0, i_8_53_552_0, i_8_53_555_0, i_8_53_556_0, i_8_53_557_0,
    i_8_53_697_0, i_8_53_698_0, i_8_53_699_0, i_8_53_700_0, i_8_53_701_0,
    i_8_53_748_0, i_8_53_838_0, i_8_53_839_0, i_8_53_850_0, i_8_53_883_0,
    i_8_53_885_0, i_8_53_886_0, i_8_53_889_0, i_8_53_995_0, i_8_53_1012_0,
    i_8_53_1128_0, i_8_53_1129_0, i_8_53_1131_0, i_8_53_1133_0,
    i_8_53_1156_0, i_8_53_1158_0, i_8_53_1202_0, i_8_53_1203_0,
    i_8_53_1205_0, i_8_53_1236_0, i_8_53_1322_0, i_8_53_1328_0,
    i_8_53_1331_0, i_8_53_1381_0, i_8_53_1427_0, i_8_53_1489_0,
    i_8_53_1551_0, i_8_53_1552_0, i_8_53_1555_0, i_8_53_1682_0,
    i_8_53_1705_0, i_8_53_1709_0, i_8_53_1726_0, i_8_53_1732_0,
    i_8_53_1749_0, i_8_53_1751_0, i_8_53_1753_0, i_8_53_1797_0,
    i_8_53_1806_0, i_8_53_1807_0, i_8_53_1841_0, i_8_53_1912_0,
    i_8_53_1913_0, i_8_53_1914_0, i_8_53_1915_0, i_8_53_1916_0,
    i_8_53_1936_0, i_8_53_1939_0, i_8_53_1982_0, i_8_53_1983_0,
    i_8_53_1985_0, i_8_53_1992_0, i_8_53_1999_0, i_8_53_2017_0,
    i_8_53_2055_0, i_8_53_2057_0, i_8_53_2058_0, i_8_53_2059_0,
    i_8_53_2144_0, i_8_53_2146_0, i_8_53_2147_0, i_8_53_2154_0,
    i_8_53_2159_0, i_8_53_2177_0, i_8_53_2272_0;
  output o_8_53_0_0;
  assign o_8_53_0_0 = ~((~i_8_53_352_0 & ((~i_8_53_1916_0 & ((~i_8_53_334_0 & ((~i_8_53_32_0 & ((~i_8_53_67_0 & ~i_8_53_172_0 & ~i_8_53_462_0 & ~i_8_53_699_0 & ~i_8_53_995_0 & ~i_8_53_1131_0 & ~i_8_53_1205_0 & ~i_8_53_1331_0 & ~i_8_53_1551_0 & ~i_8_53_1552_0 & ~i_8_53_1705_0 & ~i_8_53_1806_0 & ~i_8_53_1841_0 & ~i_8_53_2059_0 & ~i_8_53_2154_0) | (~i_8_53_43_0 & ~i_8_53_57_0 & ~i_8_53_64_0 & ~i_8_53_160_0 & ~i_8_53_502_0 & i_8_53_995_0 & ~i_8_53_1158_0 & ~i_8_53_1381_0 & ~i_8_53_1709_0 & ~i_8_53_1913_0 & ~i_8_53_2272_0))) | (~i_8_53_41_0 & ~i_8_53_43_0 & ~i_8_53_64_0 & ~i_8_53_230_0 & ~i_8_53_502_0 & ~i_8_53_1555_0 & ~i_8_53_1682_0 & ~i_8_53_1749_0 & ~i_8_53_1807_0 & ~i_8_53_1841_0 & ~i_8_53_1914_0 & ~i_8_53_1983_0 & ~i_8_53_2272_0))) | (~i_8_53_502_0 & ((~i_8_53_41_0 & ~i_8_53_1381_0 & ((~i_8_53_37_0 & ~i_8_53_64_0 & ~i_8_53_400_0 & ~i_8_53_462_0 & ~i_8_53_552_0 & ~i_8_53_557_0 & ~i_8_53_1158_0 & ~i_8_53_1202_0 & ~i_8_53_1322_0 & ~i_8_53_1331_0 & ~i_8_53_1841_0 & ~i_8_53_1912_0 & ~i_8_53_1914_0 & ~i_8_53_1915_0 & ~i_8_53_1936_0 & ~i_8_53_1999_0 & ~i_8_53_2017_0) | (~i_8_53_172_0 & ~i_8_53_401_0 & ~i_8_53_556_0 & ~i_8_53_1156_0 & ~i_8_53_1705_0 & ~i_8_53_1709_0 & ~i_8_53_1806_0 & i_8_53_2159_0 & ~i_8_53_2272_0))) | (~i_8_53_64_0 & ~i_8_53_67_0 & ~i_8_53_392_0 & ~i_8_53_838_0 & ~i_8_53_1156_0 & ~i_8_53_1158_0 & ~i_8_53_1236_0 & ~i_8_53_1328_0 & ~i_8_53_1427_0 & ~i_8_53_1709_0 & ~i_8_53_1749_0 & ~i_8_53_1753_0 & ~i_8_53_1841_0 & ~i_8_53_2017_0 & ~i_8_53_2146_0 & ~i_8_53_2177_0))) | (~i_8_53_41_0 & ~i_8_53_325_0 & ~i_8_53_552_0 & ~i_8_53_555_0 & ~i_8_53_557_0 & ~i_8_53_839_0 & ~i_8_53_1129_0 & ~i_8_53_1489_0 & ~i_8_53_1555_0 & ~i_8_53_1705_0 & ~i_8_53_1749_0 & ~i_8_53_1913_0 & ~i_8_53_1936_0 & ~i_8_53_1992_0 & ~i_8_53_2017_0 & ~i_8_53_2057_0 & ~i_8_53_2159_0 & ~i_8_53_2272_0))) | (~i_8_53_160_0 & ((i_8_53_885_0 & ~i_8_53_1128_0 & ~i_8_53_1555_0 & ~i_8_53_1936_0) | (i_8_53_229_0 & i_8_53_230_0 & ~i_8_53_839_0 & ~i_8_53_1129_0 & ~i_8_53_1203_0 & ~i_8_53_2147_0))) | (~i_8_53_205_0 & ~i_8_53_556_0 & ((~i_8_53_41_0 & ~i_8_53_172_0 & i_8_53_325_0 & ~i_8_53_400_0 & ~i_8_53_462_0 & ~i_8_53_850_0 & ~i_8_53_1131_0 & ~i_8_53_1381_0 & ~i_8_53_1749_0 & ~i_8_53_1913_0) | (~i_8_53_37_0 & ~i_8_53_64_0 & ~i_8_53_67_0 & ~i_8_53_417_0 & ~i_8_53_1156_0 & ~i_8_53_1202_0 & ~i_8_53_1203_0 & ~i_8_53_1205_0 & ~i_8_53_1427_0 & ~i_8_53_1705_0 & i_8_53_2057_0 & ~i_8_53_2177_0 & ~i_8_53_2272_0))) | (~i_8_53_172_0 & ((~i_8_53_555_0 & ~i_8_53_701_0 & ~i_8_53_1129_0 & ~i_8_53_1156_0 & i_8_53_1236_0 & ~i_8_53_1551_0 & i_8_53_1552_0 & ~i_8_53_1705_0 & ~i_8_53_2057_0 & ~i_8_53_2147_0) | (~i_8_53_37_0 & ~i_8_53_334_0 & ~i_8_53_1128_0 & ~i_8_53_1133_0 & ~i_8_53_1158_0 & ~i_8_53_1202_0 & ~i_8_53_1328_0 & ~i_8_53_1749_0 & ~i_8_53_1751_0 & ~i_8_53_1806_0 & ~i_8_53_1807_0 & ~i_8_53_1913_0 & ~i_8_53_1915_0 & ~i_8_53_1982_0 & ~i_8_53_2159_0))) | (~i_8_53_37_0 & ~i_8_53_1129_0 & ~i_8_53_1203_0 & ((~i_8_53_57_0 & ~i_8_53_228_0 & ~i_8_53_462_0 & ~i_8_53_502_0 & ~i_8_53_839_0 & ~i_8_53_1236_0 & i_8_53_1749_0 & i_8_53_1753_0 & ~i_8_53_1914_0 & ~i_8_53_2017_0) | (~i_8_53_400_0 & ~i_8_53_1133_0 & ~i_8_53_1322_0 & ~i_8_53_1705_0 & ~i_8_53_1806_0 & ~i_8_53_1936_0 & ~i_8_53_1985_0 & i_8_53_2055_0))))) | (~i_8_53_555_0 & ((~i_8_53_334_0 & ((~i_8_53_41_0 & ~i_8_53_1205_0 & ((~i_8_53_57_0 & ~i_8_53_160_0 & i_8_53_229_0 & ~i_8_53_400_0 & ~i_8_53_838_0 & ~i_8_53_1913_0 & ~i_8_53_1914_0) | (~i_8_53_43_0 & ~i_8_53_417_0 & ~i_8_53_557_0 & ~i_8_53_700_0 & ~i_8_53_1158_0 & ~i_8_53_1203_0 & ~i_8_53_1381_0 & ~i_8_53_1489_0 & ~i_8_53_1705_0 & ~i_8_53_1709_0 & ~i_8_53_1749_0 & ~i_8_53_1841_0 & ~i_8_53_1916_0 & ~i_8_53_1983_0 & ~i_8_53_2144_0))) | (~i_8_53_64_0 & ~i_8_53_1381_0 & i_8_53_1551_0 & ~i_8_53_1555_0 & ~i_8_53_1751_0 & i_8_53_1992_0 & ~i_8_53_2055_0 & ~i_8_53_2147_0))) | (~i_8_53_1133_0 & ((~i_8_53_43_0 & ~i_8_53_1012_0 & ~i_8_53_2144_0 & ((~i_8_53_400_0 & ~i_8_53_462_0 & ~i_8_53_556_0 & ~i_8_53_1328_0 & ~i_8_53_1732_0 & ~i_8_53_1797_0 & ~i_8_53_1999_0 & i_8_53_2154_0) | (~i_8_53_160_0 & ~i_8_53_417_0 & ~i_8_53_557_0 & ~i_8_53_697_0 & ~i_8_53_700_0 & ~i_8_53_838_0 & ~i_8_53_839_0 & ~i_8_53_995_0 & ~i_8_53_1322_0 & ~i_8_53_1331_0 & ~i_8_53_1156_0 & ~i_8_53_1158_0 & ~i_8_53_1916_0 & ~i_8_53_1936_0 & ~i_8_53_1985_0 & ~i_8_53_2146_0 & ~i_8_53_2272_0))) | (~i_8_53_64_0 & ~i_8_53_67_0 & ~i_8_53_172_0 & i_8_53_700_0 & ~i_8_53_1128_0 & ~i_8_53_1129_0 & ~i_8_53_1156_0 & ~i_8_53_1705_0 & ~i_8_53_1751_0 & ~i_8_53_1841_0 & ~i_8_53_1914_0 & ~i_8_53_1916_0 & ~i_8_53_2057_0 & ~i_8_53_2058_0))))) | (~i_8_53_64_0 & ((~i_8_53_67_0 & ((~i_8_53_43_0 & ~i_8_53_392_0 & ~i_8_53_1551_0 & ~i_8_53_2055_0 & ((~i_8_53_172_0 & ~i_8_53_334_0 & ~i_8_53_400_0 & ~i_8_53_401_0 & ~i_8_53_502_0 & ~i_8_53_557_0 & ~i_8_53_1427_0 & ~i_8_53_1489_0 & ~i_8_53_1555_0 & ~i_8_53_1732_0 & ~i_8_53_1916_0) | (~i_8_53_32_0 & ~i_8_53_37_0 & i_8_53_700_0 & ~i_8_53_995_0 & ~i_8_53_1331_0 & ~i_8_53_1709_0 & ~i_8_53_1726_0 & ~i_8_53_1806_0 & ~i_8_53_1913_0 & ~i_8_53_1999_0))) | (i_8_53_120_0 & ~i_8_53_1709_0 & ~i_8_53_1797_0 & ~i_8_53_1915_0 & i_8_53_1992_0))) | (~i_8_53_1131_0 & ~i_8_53_2017_0 & ((~i_8_53_839_0 & ~i_8_53_1133_0 & ~i_8_53_1203_0 & ~i_8_53_1489_0 & ~i_8_53_1912_0 & ~i_8_53_1913_0 & ~i_8_53_1914_0 & ~i_8_53_1916_0 & i_8_53_2058_0) | (~i_8_53_41_0 & i_8_53_57_0 & ~i_8_53_552_0 & ~i_8_53_1128_0 & ~i_8_53_1129_0 & ~i_8_53_1202_0 & ~i_8_53_1915_0 & ~i_8_53_2159_0))) | (i_8_53_326_0 & ~i_8_53_995_0 & ~i_8_53_1427_0 & ~i_8_53_1489_0 & ~i_8_53_1555_0 & ~i_8_53_1841_0 & ~i_8_53_1939_0))) | (~i_8_53_2017_0 & ((~i_8_53_172_0 & ~i_8_53_1331_0 & ((i_8_53_230_0 & ~i_8_53_502_0 & ~i_8_53_748_0 & ~i_8_53_1128_0 & ~i_8_53_1202_0 & ~i_8_53_1381_0 & ~i_8_53_1797_0 & ~i_8_53_1916_0 & ~i_8_53_1992_0 & ~i_8_53_2154_0) | (~i_8_53_41_0 & ~i_8_53_120_0 & ~i_8_53_334_0 & ~i_8_53_392_0 & ~i_8_53_556_0 & ~i_8_53_557_0 & ~i_8_53_839_0 & ~i_8_53_1158_0 & ~i_8_53_1328_0 & ~i_8_53_1489_0 & i_8_53_1552_0 & ~i_8_53_1807_0 & ~i_8_53_1999_0 & ~i_8_53_2057_0 & ~i_8_53_2059_0 & ~i_8_53_2272_0))) | (~i_8_53_1236_0 & ((~i_8_53_1156_0 & ((i_8_53_838_0 & ~i_8_53_1128_0 & i_8_53_1983_0 & ~i_8_53_2147_0) | (~i_8_53_401_0 & ~i_8_53_502_0 & ~i_8_53_67_0 & ~i_8_53_334_0 & ~i_8_53_850_0 & ~i_8_53_1131_0 & ~i_8_53_557_0 & ~i_8_53_838_0 & ~i_8_53_1205_0 & ~i_8_53_1427_0 & ~i_8_53_1709_0 & ~i_8_53_1751_0 & ~i_8_53_1753_0 & ~i_8_53_1914_0 & ~i_8_53_1936_0 & ~i_8_53_2059_0 & ~i_8_53_2177_0))) | (~i_8_53_1322_0 & ~i_8_53_1381_0 & i_8_53_1552_0 & ~i_8_53_1753_0 & ~i_8_53_1841_0 & ~i_8_53_1912_0 & ~i_8_53_1936_0 & ~i_8_53_1983_0 & i_8_53_1985_0))))) | (~i_8_53_37_0 & ((~i_8_53_41_0 & ~i_8_53_1131_0 & ((~i_8_53_172_0 & ~i_8_53_552_0 & ~i_8_53_557_0 & ~i_8_53_1205_0 & ~i_8_53_1328_0 & i_8_53_1555_0 & ~i_8_53_1705_0 & ~i_8_53_1709_0 & ~i_8_53_1751_0 & ~i_8_53_1806_0 & ~i_8_53_1807_0) | (i_8_53_699_0 & ~i_8_53_1133_0 & ~i_8_53_1158_0 & ~i_8_53_1914_0 & ~i_8_53_1915_0 & i_8_53_2055_0 & ~i_8_53_2272_0))) | (~i_8_53_462_0 & ~i_8_53_1202_0 & ~i_8_53_1328_0 & ~i_8_53_1427_0 & ~i_8_53_1705_0 & ~i_8_53_1912_0 & ~i_8_53_1913_0 & ~i_8_53_1916_0 & i_8_53_1985_0 & ~i_8_53_2144_0 & ~i_8_53_2154_0))) | (~i_8_53_1427_0 & ~i_8_53_1916_0 & ((~i_8_53_172_0 & ~i_8_53_400_0 & i_8_53_698_0 & ~i_8_53_748_0 & ~i_8_53_839_0 & ~i_8_53_1012_0 & ~i_8_53_1131_0 & ~i_8_53_1331_0 & ~i_8_53_1705_0 & ~i_8_53_1751_0 & ~i_8_53_1999_0) | (i_8_53_228_0 & i_8_53_229_0 & ~i_8_53_462_0 & ~i_8_53_1797_0 & ~i_8_53_1915_0 & ~i_8_53_1985_0 & ~i_8_53_2144_0))) | (i_8_53_329_0 & ~i_8_53_417_0 & ~i_8_53_556_0 & ~i_8_53_1322_0 & ~i_8_53_1705_0 & ~i_8_53_1709_0 & ~i_8_53_1913_0 & ~i_8_53_1999_0 & i_8_53_2057_0) | (~i_8_53_838_0 & ~i_8_53_1128_0 & i_8_53_1551_0 & i_8_53_1555_0 & ~i_8_53_1682_0 & ~i_8_53_1726_0 & ~i_8_53_1749_0 & ~i_8_53_1807_0 & ~i_8_53_2147_0 & ~i_8_53_2154_0) | (i_8_53_325_0 & i_8_53_995_0 & i_8_53_2154_0 & ~i_8_53_2272_0));
endmodule



// Benchmark "kernel_8_54" written by ABC on Sun Jul 19 10:03:57 2020

module kernel_8_54 ( 
    i_8_54_31_0, i_8_54_32_0, i_8_54_52_0, i_8_54_55_0, i_8_54_79_0,
    i_8_54_97_0, i_8_54_104_0, i_8_54_208_0, i_8_54_212_0, i_8_54_258_0,
    i_8_54_262_0, i_8_54_283_0, i_8_54_292_0, i_8_54_301_0, i_8_54_363_0,
    i_8_54_382_0, i_8_54_384_0, i_8_54_427_0, i_8_54_454_0, i_8_54_456_0,
    i_8_54_492_0, i_8_54_624_0, i_8_54_625_0, i_8_54_628_0, i_8_54_636_0,
    i_8_54_669_0, i_8_54_670_0, i_8_54_679_0, i_8_54_682_0, i_8_54_696_0,
    i_8_54_698_0, i_8_54_701_0, i_8_54_719_0, i_8_54_727_0, i_8_54_733_0,
    i_8_54_738_0, i_8_54_781_0, i_8_54_784_0, i_8_54_786_0, i_8_54_792_0,
    i_8_54_800_0, i_8_54_827_0, i_8_54_840_0, i_8_54_853_0, i_8_54_880_0,
    i_8_54_915_0, i_8_54_958_0, i_8_54_1029_0, i_8_54_1059_0,
    i_8_54_1108_0, i_8_54_1114_0, i_8_54_1138_0, i_8_54_1229_0,
    i_8_54_1249_0, i_8_54_1282_0, i_8_54_1285_0, i_8_54_1335_0,
    i_8_54_1354_0, i_8_54_1355_0, i_8_54_1381_0, i_8_54_1438_0,
    i_8_54_1444_0, i_8_54_1454_0, i_8_54_1542_0, i_8_54_1543_0,
    i_8_54_1565_0, i_8_54_1588_0, i_8_54_1591_0, i_8_54_1606_0,
    i_8_54_1683_0, i_8_54_1684_0, i_8_54_1700_0, i_8_54_1706_0,
    i_8_54_1732_0, i_8_54_1736_0, i_8_54_1762_0, i_8_54_1771_0,
    i_8_54_1794_0, i_8_54_1805_0, i_8_54_1808_0, i_8_54_1822_0,
    i_8_54_1823_0, i_8_54_1825_0, i_8_54_1858_0, i_8_54_1860_0,
    i_8_54_1867_0, i_8_54_1885_0, i_8_54_1912_0, i_8_54_1966_0,
    i_8_54_1983_0, i_8_54_1997_0, i_8_54_2147_0, i_8_54_2190_0,
    i_8_54_2193_0, i_8_54_2200_0, i_8_54_2215_0, i_8_54_2229_0,
    i_8_54_2247_0, i_8_54_2263_0, i_8_54_2284_0,
    o_8_54_0_0  );
  input  i_8_54_31_0, i_8_54_32_0, i_8_54_52_0, i_8_54_55_0, i_8_54_79_0,
    i_8_54_97_0, i_8_54_104_0, i_8_54_208_0, i_8_54_212_0, i_8_54_258_0,
    i_8_54_262_0, i_8_54_283_0, i_8_54_292_0, i_8_54_301_0, i_8_54_363_0,
    i_8_54_382_0, i_8_54_384_0, i_8_54_427_0, i_8_54_454_0, i_8_54_456_0,
    i_8_54_492_0, i_8_54_624_0, i_8_54_625_0, i_8_54_628_0, i_8_54_636_0,
    i_8_54_669_0, i_8_54_670_0, i_8_54_679_0, i_8_54_682_0, i_8_54_696_0,
    i_8_54_698_0, i_8_54_701_0, i_8_54_719_0, i_8_54_727_0, i_8_54_733_0,
    i_8_54_738_0, i_8_54_781_0, i_8_54_784_0, i_8_54_786_0, i_8_54_792_0,
    i_8_54_800_0, i_8_54_827_0, i_8_54_840_0, i_8_54_853_0, i_8_54_880_0,
    i_8_54_915_0, i_8_54_958_0, i_8_54_1029_0, i_8_54_1059_0,
    i_8_54_1108_0, i_8_54_1114_0, i_8_54_1138_0, i_8_54_1229_0,
    i_8_54_1249_0, i_8_54_1282_0, i_8_54_1285_0, i_8_54_1335_0,
    i_8_54_1354_0, i_8_54_1355_0, i_8_54_1381_0, i_8_54_1438_0,
    i_8_54_1444_0, i_8_54_1454_0, i_8_54_1542_0, i_8_54_1543_0,
    i_8_54_1565_0, i_8_54_1588_0, i_8_54_1591_0, i_8_54_1606_0,
    i_8_54_1683_0, i_8_54_1684_0, i_8_54_1700_0, i_8_54_1706_0,
    i_8_54_1732_0, i_8_54_1736_0, i_8_54_1762_0, i_8_54_1771_0,
    i_8_54_1794_0, i_8_54_1805_0, i_8_54_1808_0, i_8_54_1822_0,
    i_8_54_1823_0, i_8_54_1825_0, i_8_54_1858_0, i_8_54_1860_0,
    i_8_54_1867_0, i_8_54_1885_0, i_8_54_1912_0, i_8_54_1966_0,
    i_8_54_1983_0, i_8_54_1997_0, i_8_54_2147_0, i_8_54_2190_0,
    i_8_54_2193_0, i_8_54_2200_0, i_8_54_2215_0, i_8_54_2229_0,
    i_8_54_2247_0, i_8_54_2263_0, i_8_54_2284_0;
  output o_8_54_0_0;
  assign o_8_54_0_0 = 0;
endmodule



// Benchmark "kernel_8_55" written by ABC on Sun Jul 19 10:03:58 2020

module kernel_8_55 ( 
    i_8_55_6_0, i_8_55_23_0, i_8_55_30_0, i_8_55_41_0, i_8_55_65_0,
    i_8_55_68_0, i_8_55_85_0, i_8_55_86_0, i_8_55_137_0, i_8_55_142_0,
    i_8_55_145_0, i_8_55_175_0, i_8_55_176_0, i_8_55_199_0, i_8_55_205_0,
    i_8_55_247_0, i_8_55_282_0, i_8_55_335_0, i_8_55_355_0, i_8_55_356_0,
    i_8_55_364_0, i_8_55_368_0, i_8_55_437_0, i_8_55_440_0, i_8_55_444_0,
    i_8_55_445_0, i_8_55_497_0, i_8_55_517_0, i_8_55_527_0, i_8_55_550_0,
    i_8_55_588_0, i_8_55_597_0, i_8_55_615_0, i_8_55_661_0, i_8_55_682_0,
    i_8_55_699_0, i_8_55_707_0, i_8_55_710_0, i_8_55_713_0, i_8_55_715_0,
    i_8_55_727_0, i_8_55_728_0, i_8_55_770_0, i_8_55_914_0, i_8_55_958_0,
    i_8_55_971_0, i_8_55_992_0, i_8_55_1084_0, i_8_55_1127_0,
    i_8_55_1134_0, i_8_55_1229_0, i_8_55_1236_0, i_8_55_1267_0,
    i_8_55_1282_0, i_8_55_1305_0, i_8_55_1351_0, i_8_55_1363_0,
    i_8_55_1391_0, i_8_55_1407_0, i_8_55_1425_0, i_8_55_1437_0,
    i_8_55_1438_0, i_8_55_1447_0, i_8_55_1484_0, i_8_55_1487_0,
    i_8_55_1490_0, i_8_55_1525_0, i_8_55_1549_0, i_8_55_1598_0,
    i_8_55_1629_0, i_8_55_1642_0, i_8_55_1646_0, i_8_55_1654_0,
    i_8_55_1687_0, i_8_55_1700_0, i_8_55_1706_0, i_8_55_1745_0,
    i_8_55_1779_0, i_8_55_1781_0, i_8_55_1794_0, i_8_55_1813_0,
    i_8_55_1819_0, i_8_55_1820_0, i_8_55_1823_0, i_8_55_1837_0,
    i_8_55_1850_0, i_8_55_1873_0, i_8_55_1884_0, i_8_55_1916_0,
    i_8_55_1980_0, i_8_55_2004_0, i_8_55_2044_0, i_8_55_2046_0,
    i_8_55_2066_0, i_8_55_2090_0, i_8_55_2098_0, i_8_55_2147_0,
    i_8_55_2183_0, i_8_55_2238_0, i_8_55_2289_0,
    o_8_55_0_0  );
  input  i_8_55_6_0, i_8_55_23_0, i_8_55_30_0, i_8_55_41_0, i_8_55_65_0,
    i_8_55_68_0, i_8_55_85_0, i_8_55_86_0, i_8_55_137_0, i_8_55_142_0,
    i_8_55_145_0, i_8_55_175_0, i_8_55_176_0, i_8_55_199_0, i_8_55_205_0,
    i_8_55_247_0, i_8_55_282_0, i_8_55_335_0, i_8_55_355_0, i_8_55_356_0,
    i_8_55_364_0, i_8_55_368_0, i_8_55_437_0, i_8_55_440_0, i_8_55_444_0,
    i_8_55_445_0, i_8_55_497_0, i_8_55_517_0, i_8_55_527_0, i_8_55_550_0,
    i_8_55_588_0, i_8_55_597_0, i_8_55_615_0, i_8_55_661_0, i_8_55_682_0,
    i_8_55_699_0, i_8_55_707_0, i_8_55_710_0, i_8_55_713_0, i_8_55_715_0,
    i_8_55_727_0, i_8_55_728_0, i_8_55_770_0, i_8_55_914_0, i_8_55_958_0,
    i_8_55_971_0, i_8_55_992_0, i_8_55_1084_0, i_8_55_1127_0,
    i_8_55_1134_0, i_8_55_1229_0, i_8_55_1236_0, i_8_55_1267_0,
    i_8_55_1282_0, i_8_55_1305_0, i_8_55_1351_0, i_8_55_1363_0,
    i_8_55_1391_0, i_8_55_1407_0, i_8_55_1425_0, i_8_55_1437_0,
    i_8_55_1438_0, i_8_55_1447_0, i_8_55_1484_0, i_8_55_1487_0,
    i_8_55_1490_0, i_8_55_1525_0, i_8_55_1549_0, i_8_55_1598_0,
    i_8_55_1629_0, i_8_55_1642_0, i_8_55_1646_0, i_8_55_1654_0,
    i_8_55_1687_0, i_8_55_1700_0, i_8_55_1706_0, i_8_55_1745_0,
    i_8_55_1779_0, i_8_55_1781_0, i_8_55_1794_0, i_8_55_1813_0,
    i_8_55_1819_0, i_8_55_1820_0, i_8_55_1823_0, i_8_55_1837_0,
    i_8_55_1850_0, i_8_55_1873_0, i_8_55_1884_0, i_8_55_1916_0,
    i_8_55_1980_0, i_8_55_2004_0, i_8_55_2044_0, i_8_55_2046_0,
    i_8_55_2066_0, i_8_55_2090_0, i_8_55_2098_0, i_8_55_2147_0,
    i_8_55_2183_0, i_8_55_2238_0, i_8_55_2289_0;
  output o_8_55_0_0;
  assign o_8_55_0_0 = 0;
endmodule



// Benchmark "kernel_8_56" written by ABC on Sun Jul 19 10:03:59 2020

module kernel_8_56 ( 
    i_8_56_20_0, i_8_56_65_0, i_8_56_76_0, i_8_56_77_0, i_8_56_94_0,
    i_8_56_112_0, i_8_56_245_0, i_8_56_353_0, i_8_56_388_0, i_8_56_389_0,
    i_8_56_443_0, i_8_56_461_0, i_8_56_481_0, i_8_56_486_0, i_8_56_497_0,
    i_8_56_515_0, i_8_56_524_0, i_8_56_529_0, i_8_56_549_0, i_8_56_550_0,
    i_8_56_595_0, i_8_56_605_0, i_8_56_631_0, i_8_56_632_0, i_8_56_633_0,
    i_8_56_658_0, i_8_56_716_0, i_8_56_812_0, i_8_56_830_0, i_8_56_841_0,
    i_8_56_843_0, i_8_56_873_0, i_8_56_875_0, i_8_56_877_0, i_8_56_883_0,
    i_8_56_926_0, i_8_56_965_0, i_8_56_967_0, i_8_56_1040_0, i_8_56_1073_0,
    i_8_56_1127_0, i_8_56_1143_0, i_8_56_1144_0, i_8_56_1153_0,
    i_8_56_1171_0, i_8_56_1198_0, i_8_56_1199_0, i_8_56_1269_0,
    i_8_56_1283_0, i_8_56_1298_0, i_8_56_1315_0, i_8_56_1351_0,
    i_8_56_1382_0, i_8_56_1396_0, i_8_56_1397_0, i_8_56_1424_0,
    i_8_56_1431_0, i_8_56_1433_0, i_8_56_1451_0, i_8_56_1468_0,
    i_8_56_1495_0, i_8_56_1513_0, i_8_56_1514_0, i_8_56_1523_0,
    i_8_56_1532_0, i_8_56_1621_0, i_8_56_1649_0, i_8_56_1657_0,
    i_8_56_1658_0, i_8_56_1681_0, i_8_56_1702_0, i_8_56_1703_0,
    i_8_56_1730_0, i_8_56_1747_0, i_8_56_1773_0, i_8_56_1791_0,
    i_8_56_1792_0, i_8_56_1793_0, i_8_56_1823_0, i_8_56_1824_0,
    i_8_56_1864_0, i_8_56_1882_0, i_8_56_1909_0, i_8_56_1910_0,
    i_8_56_1936_0, i_8_56_1981_0, i_8_56_2044_0, i_8_56_2052_0,
    i_8_56_2053_0, i_8_56_2099_0, i_8_56_2117_0, i_8_56_2134_0,
    i_8_56_2143_0, i_8_56_2169_0, i_8_56_2171_0, i_8_56_2224_0,
    i_8_56_2234_0, i_8_56_2243_0, i_8_56_2254_0, i_8_56_2283_0,
    o_8_56_0_0  );
  input  i_8_56_20_0, i_8_56_65_0, i_8_56_76_0, i_8_56_77_0, i_8_56_94_0,
    i_8_56_112_0, i_8_56_245_0, i_8_56_353_0, i_8_56_388_0, i_8_56_389_0,
    i_8_56_443_0, i_8_56_461_0, i_8_56_481_0, i_8_56_486_0, i_8_56_497_0,
    i_8_56_515_0, i_8_56_524_0, i_8_56_529_0, i_8_56_549_0, i_8_56_550_0,
    i_8_56_595_0, i_8_56_605_0, i_8_56_631_0, i_8_56_632_0, i_8_56_633_0,
    i_8_56_658_0, i_8_56_716_0, i_8_56_812_0, i_8_56_830_0, i_8_56_841_0,
    i_8_56_843_0, i_8_56_873_0, i_8_56_875_0, i_8_56_877_0, i_8_56_883_0,
    i_8_56_926_0, i_8_56_965_0, i_8_56_967_0, i_8_56_1040_0, i_8_56_1073_0,
    i_8_56_1127_0, i_8_56_1143_0, i_8_56_1144_0, i_8_56_1153_0,
    i_8_56_1171_0, i_8_56_1198_0, i_8_56_1199_0, i_8_56_1269_0,
    i_8_56_1283_0, i_8_56_1298_0, i_8_56_1315_0, i_8_56_1351_0,
    i_8_56_1382_0, i_8_56_1396_0, i_8_56_1397_0, i_8_56_1424_0,
    i_8_56_1431_0, i_8_56_1433_0, i_8_56_1451_0, i_8_56_1468_0,
    i_8_56_1495_0, i_8_56_1513_0, i_8_56_1514_0, i_8_56_1523_0,
    i_8_56_1532_0, i_8_56_1621_0, i_8_56_1649_0, i_8_56_1657_0,
    i_8_56_1658_0, i_8_56_1681_0, i_8_56_1702_0, i_8_56_1703_0,
    i_8_56_1730_0, i_8_56_1747_0, i_8_56_1773_0, i_8_56_1791_0,
    i_8_56_1792_0, i_8_56_1793_0, i_8_56_1823_0, i_8_56_1824_0,
    i_8_56_1864_0, i_8_56_1882_0, i_8_56_1909_0, i_8_56_1910_0,
    i_8_56_1936_0, i_8_56_1981_0, i_8_56_2044_0, i_8_56_2052_0,
    i_8_56_2053_0, i_8_56_2099_0, i_8_56_2117_0, i_8_56_2134_0,
    i_8_56_2143_0, i_8_56_2169_0, i_8_56_2171_0, i_8_56_2224_0,
    i_8_56_2234_0, i_8_56_2243_0, i_8_56_2254_0, i_8_56_2283_0;
  output o_8_56_0_0;
  assign o_8_56_0_0 = 0;
endmodule



// Benchmark "kernel_8_57" written by ABC on Sun Jul 19 10:04:00 2020

module kernel_8_57 ( 
    i_8_57_156_0, i_8_57_258_0, i_8_57_348_0, i_8_57_372_0, i_8_57_380_0,
    i_8_57_441_0, i_8_57_458_0, i_8_57_462_0, i_8_57_463_0, i_8_57_468_0,
    i_8_57_474_0, i_8_57_475_0, i_8_57_480_0, i_8_57_503_0, i_8_57_552_0,
    i_8_57_585_0, i_8_57_607_0, i_8_57_639_0, i_8_57_642_0, i_8_57_669_0,
    i_8_57_719_0, i_8_57_720_0, i_8_57_778_0, i_8_57_793_0, i_8_57_811_0,
    i_8_57_831_0, i_8_57_837_0, i_8_57_838_0, i_8_57_841_0, i_8_57_870_0,
    i_8_57_950_0, i_8_57_973_0, i_8_57_1011_0, i_8_57_1014_0,
    i_8_57_1066_0, i_8_57_1071_0, i_8_57_1072_0, i_8_57_1074_0,
    i_8_57_1075_0, i_8_57_1083_0, i_8_57_1084_0, i_8_57_1129_0,
    i_8_57_1134_0, i_8_57_1218_0, i_8_57_1225_0, i_8_57_1236_0,
    i_8_57_1237_0, i_8_57_1249_0, i_8_57_1252_0, i_8_57_1254_0,
    i_8_57_1255_0, i_8_57_1261_0, i_8_57_1263_0, i_8_57_1272_0,
    i_8_57_1283_0, i_8_57_1285_0, i_8_57_1288_0, i_8_57_1305_0,
    i_8_57_1306_0, i_8_57_1307_0, i_8_57_1378_0, i_8_57_1419_0,
    i_8_57_1452_0, i_8_57_1467_0, i_8_57_1519_0, i_8_57_1535_0,
    i_8_57_1542_0, i_8_57_1584_0, i_8_57_1587_0, i_8_57_1593_0,
    i_8_57_1596_0, i_8_57_1605_0, i_8_57_1606_0, i_8_57_1611_0,
    i_8_57_1624_0, i_8_57_1641_0, i_8_57_1659_0, i_8_57_1680_0,
    i_8_57_1704_0, i_8_57_1705_0, i_8_57_1718_0, i_8_57_1720_0,
    i_8_57_1747_0, i_8_57_1764_0, i_8_57_1767_0, i_8_57_1783_0,
    i_8_57_1803_0, i_8_57_1804_0, i_8_57_1805_0, i_8_57_1815_0,
    i_8_57_1828_0, i_8_57_1864_0, i_8_57_1981_0, i_8_57_2037_0,
    i_8_57_2124_0, i_8_57_2143_0, i_8_57_2146_0, i_8_57_2154_0,
    i_8_57_2272_0, i_8_57_2274_0,
    o_8_57_0_0  );
  input  i_8_57_156_0, i_8_57_258_0, i_8_57_348_0, i_8_57_372_0,
    i_8_57_380_0, i_8_57_441_0, i_8_57_458_0, i_8_57_462_0, i_8_57_463_0,
    i_8_57_468_0, i_8_57_474_0, i_8_57_475_0, i_8_57_480_0, i_8_57_503_0,
    i_8_57_552_0, i_8_57_585_0, i_8_57_607_0, i_8_57_639_0, i_8_57_642_0,
    i_8_57_669_0, i_8_57_719_0, i_8_57_720_0, i_8_57_778_0, i_8_57_793_0,
    i_8_57_811_0, i_8_57_831_0, i_8_57_837_0, i_8_57_838_0, i_8_57_841_0,
    i_8_57_870_0, i_8_57_950_0, i_8_57_973_0, i_8_57_1011_0, i_8_57_1014_0,
    i_8_57_1066_0, i_8_57_1071_0, i_8_57_1072_0, i_8_57_1074_0,
    i_8_57_1075_0, i_8_57_1083_0, i_8_57_1084_0, i_8_57_1129_0,
    i_8_57_1134_0, i_8_57_1218_0, i_8_57_1225_0, i_8_57_1236_0,
    i_8_57_1237_0, i_8_57_1249_0, i_8_57_1252_0, i_8_57_1254_0,
    i_8_57_1255_0, i_8_57_1261_0, i_8_57_1263_0, i_8_57_1272_0,
    i_8_57_1283_0, i_8_57_1285_0, i_8_57_1288_0, i_8_57_1305_0,
    i_8_57_1306_0, i_8_57_1307_0, i_8_57_1378_0, i_8_57_1419_0,
    i_8_57_1452_0, i_8_57_1467_0, i_8_57_1519_0, i_8_57_1535_0,
    i_8_57_1542_0, i_8_57_1584_0, i_8_57_1587_0, i_8_57_1593_0,
    i_8_57_1596_0, i_8_57_1605_0, i_8_57_1606_0, i_8_57_1611_0,
    i_8_57_1624_0, i_8_57_1641_0, i_8_57_1659_0, i_8_57_1680_0,
    i_8_57_1704_0, i_8_57_1705_0, i_8_57_1718_0, i_8_57_1720_0,
    i_8_57_1747_0, i_8_57_1764_0, i_8_57_1767_0, i_8_57_1783_0,
    i_8_57_1803_0, i_8_57_1804_0, i_8_57_1805_0, i_8_57_1815_0,
    i_8_57_1828_0, i_8_57_1864_0, i_8_57_1981_0, i_8_57_2037_0,
    i_8_57_2124_0, i_8_57_2143_0, i_8_57_2146_0, i_8_57_2154_0,
    i_8_57_2272_0, i_8_57_2274_0;
  output o_8_57_0_0;
  assign o_8_57_0_0 = 0;
endmodule



// Benchmark "kernel_8_58" written by ABC on Sun Jul 19 10:04:00 2020

module kernel_8_58 ( 
    i_8_58_54_0, i_8_58_86_0, i_8_58_89_0, i_8_58_97_0, i_8_58_111_0,
    i_8_58_254_0, i_8_58_257_0, i_8_58_259_0, i_8_58_266_0, i_8_58_279_0,
    i_8_58_328_0, i_8_58_334_0, i_8_58_344_0, i_8_58_390_0, i_8_58_449_0,
    i_8_58_454_0, i_8_58_455_0, i_8_58_489_0, i_8_58_500_0, i_8_58_511_0,
    i_8_58_525_0, i_8_58_527_0, i_8_58_530_0, i_8_58_628_0, i_8_58_662_0,
    i_8_58_666_0, i_8_58_670_0, i_8_58_674_0, i_8_58_683_0, i_8_58_716_0,
    i_8_58_725_0, i_8_58_742_0, i_8_58_759_0, i_8_58_789_0, i_8_58_791_0,
    i_8_58_796_0, i_8_58_815_0, i_8_58_834_0, i_8_58_842_0, i_8_58_856_0,
    i_8_58_874_0, i_8_58_881_0, i_8_58_952_0, i_8_58_953_0, i_8_58_1030_0,
    i_8_58_1114_0, i_8_58_1120_0, i_8_58_1132_0, i_8_58_1138_0,
    i_8_58_1159_0, i_8_58_1160_0, i_8_58_1200_0, i_8_58_1236_0,
    i_8_58_1237_0, i_8_58_1238_0, i_8_58_1262_0, i_8_58_1283_0,
    i_8_58_1294_0, i_8_58_1321_0, i_8_58_1347_0, i_8_58_1406_0,
    i_8_58_1473_0, i_8_58_1527_0, i_8_58_1528_0, i_8_58_1536_0,
    i_8_58_1548_0, i_8_58_1588_0, i_8_58_1589_0, i_8_58_1634_0,
    i_8_58_1676_0, i_8_58_1700_0, i_8_58_1707_0, i_8_58_1717_0,
    i_8_58_1727_0, i_8_58_1729_0, i_8_58_1732_0, i_8_58_1751_0,
    i_8_58_1796_0, i_8_58_1807_0, i_8_58_1808_0, i_8_58_1814_0,
    i_8_58_1858_0, i_8_58_1859_0, i_8_58_1903_0, i_8_58_1904_0,
    i_8_58_1918_0, i_8_58_1921_0, i_8_58_1930_0, i_8_58_1976_0,
    i_8_58_1984_0, i_8_58_2011_0, i_8_58_2012_0, i_8_58_2028_0,
    i_8_58_2029_0, i_8_58_2032_0, i_8_58_2151_0, i_8_58_2174_0,
    i_8_58_2215_0, i_8_58_2216_0, i_8_58_2292_0,
    o_8_58_0_0  );
  input  i_8_58_54_0, i_8_58_86_0, i_8_58_89_0, i_8_58_97_0,
    i_8_58_111_0, i_8_58_254_0, i_8_58_257_0, i_8_58_259_0, i_8_58_266_0,
    i_8_58_279_0, i_8_58_328_0, i_8_58_334_0, i_8_58_344_0, i_8_58_390_0,
    i_8_58_449_0, i_8_58_454_0, i_8_58_455_0, i_8_58_489_0, i_8_58_500_0,
    i_8_58_511_0, i_8_58_525_0, i_8_58_527_0, i_8_58_530_0, i_8_58_628_0,
    i_8_58_662_0, i_8_58_666_0, i_8_58_670_0, i_8_58_674_0, i_8_58_683_0,
    i_8_58_716_0, i_8_58_725_0, i_8_58_742_0, i_8_58_759_0, i_8_58_789_0,
    i_8_58_791_0, i_8_58_796_0, i_8_58_815_0, i_8_58_834_0, i_8_58_842_0,
    i_8_58_856_0, i_8_58_874_0, i_8_58_881_0, i_8_58_952_0, i_8_58_953_0,
    i_8_58_1030_0, i_8_58_1114_0, i_8_58_1120_0, i_8_58_1132_0,
    i_8_58_1138_0, i_8_58_1159_0, i_8_58_1160_0, i_8_58_1200_0,
    i_8_58_1236_0, i_8_58_1237_0, i_8_58_1238_0, i_8_58_1262_0,
    i_8_58_1283_0, i_8_58_1294_0, i_8_58_1321_0, i_8_58_1347_0,
    i_8_58_1406_0, i_8_58_1473_0, i_8_58_1527_0, i_8_58_1528_0,
    i_8_58_1536_0, i_8_58_1548_0, i_8_58_1588_0, i_8_58_1589_0,
    i_8_58_1634_0, i_8_58_1676_0, i_8_58_1700_0, i_8_58_1707_0,
    i_8_58_1717_0, i_8_58_1727_0, i_8_58_1729_0, i_8_58_1732_0,
    i_8_58_1751_0, i_8_58_1796_0, i_8_58_1807_0, i_8_58_1808_0,
    i_8_58_1814_0, i_8_58_1858_0, i_8_58_1859_0, i_8_58_1903_0,
    i_8_58_1904_0, i_8_58_1918_0, i_8_58_1921_0, i_8_58_1930_0,
    i_8_58_1976_0, i_8_58_1984_0, i_8_58_2011_0, i_8_58_2012_0,
    i_8_58_2028_0, i_8_58_2029_0, i_8_58_2032_0, i_8_58_2151_0,
    i_8_58_2174_0, i_8_58_2215_0, i_8_58_2216_0, i_8_58_2292_0;
  output o_8_58_0_0;
  assign o_8_58_0_0 = 0;
endmodule



// Benchmark "kernel_8_59" written by ABC on Sun Jul 19 10:04:01 2020

module kernel_8_59 ( 
    i_8_59_20_0, i_8_59_29_0, i_8_59_30_0, i_8_59_47_0, i_8_59_50_0,
    i_8_59_56_0, i_8_59_74_0, i_8_59_77_0, i_8_59_112_0, i_8_59_113_0,
    i_8_59_137_0, i_8_59_165_0, i_8_59_229_0, i_8_59_253_0, i_8_59_254_0,
    i_8_59_256_0, i_8_59_262_0, i_8_59_376_0, i_8_59_420_0, i_8_59_442_0,
    i_8_59_451_0, i_8_59_452_0, i_8_59_454_0, i_8_59_455_0, i_8_59_590_0,
    i_8_59_596_0, i_8_59_644_0, i_8_59_665_0, i_8_59_677_0, i_8_59_694_0,
    i_8_59_695_0, i_8_59_707_0, i_8_59_776_0, i_8_59_784_0, i_8_59_796_0,
    i_8_59_823_0, i_8_59_875_0, i_8_59_878_0, i_8_59_965_0, i_8_59_991_0,
    i_8_59_994_0, i_8_59_1038_0, i_8_59_1111_0, i_8_59_1120_0,
    i_8_59_1139_0, i_8_59_1163_0, i_8_59_1202_0, i_8_59_1226_0,
    i_8_59_1253_0, i_8_59_1255_0, i_8_59_1260_0, i_8_59_1289_0,
    i_8_59_1318_0, i_8_59_1334_0, i_8_59_1342_0, i_8_59_1379_0,
    i_8_59_1400_0, i_8_59_1487_0, i_8_59_1538_0, i_8_59_1546_0,
    i_8_59_1552_0, i_8_59_1559_0, i_8_59_1631_0, i_8_59_1637_0,
    i_8_59_1666_0, i_8_59_1675_0, i_8_59_1679_0, i_8_59_1681_0,
    i_8_59_1682_0, i_8_59_1687_0, i_8_59_1697_0, i_8_59_1701_0,
    i_8_59_1755_0, i_8_59_1757_0, i_8_59_1770_0, i_8_59_1772_0,
    i_8_59_1784_0, i_8_59_1789_0, i_8_59_1840_0, i_8_59_1882_0,
    i_8_59_1885_0, i_8_59_1904_0, i_8_59_1910_0, i_8_59_1918_0,
    i_8_59_1960_0, i_8_59_1984_0, i_8_59_1990_0, i_8_59_1994_0,
    i_8_59_1995_0, i_8_59_2033_0, i_8_59_2075_0, i_8_59_2099_0,
    i_8_59_2108_0, i_8_59_2136_0, i_8_59_2146_0, i_8_59_2156_0,
    i_8_59_2224_0, i_8_59_2233_0, i_8_59_2241_0, i_8_59_2260_0,
    o_8_59_0_0  );
  input  i_8_59_20_0, i_8_59_29_0, i_8_59_30_0, i_8_59_47_0, i_8_59_50_0,
    i_8_59_56_0, i_8_59_74_0, i_8_59_77_0, i_8_59_112_0, i_8_59_113_0,
    i_8_59_137_0, i_8_59_165_0, i_8_59_229_0, i_8_59_253_0, i_8_59_254_0,
    i_8_59_256_0, i_8_59_262_0, i_8_59_376_0, i_8_59_420_0, i_8_59_442_0,
    i_8_59_451_0, i_8_59_452_0, i_8_59_454_0, i_8_59_455_0, i_8_59_590_0,
    i_8_59_596_0, i_8_59_644_0, i_8_59_665_0, i_8_59_677_0, i_8_59_694_0,
    i_8_59_695_0, i_8_59_707_0, i_8_59_776_0, i_8_59_784_0, i_8_59_796_0,
    i_8_59_823_0, i_8_59_875_0, i_8_59_878_0, i_8_59_965_0, i_8_59_991_0,
    i_8_59_994_0, i_8_59_1038_0, i_8_59_1111_0, i_8_59_1120_0,
    i_8_59_1139_0, i_8_59_1163_0, i_8_59_1202_0, i_8_59_1226_0,
    i_8_59_1253_0, i_8_59_1255_0, i_8_59_1260_0, i_8_59_1289_0,
    i_8_59_1318_0, i_8_59_1334_0, i_8_59_1342_0, i_8_59_1379_0,
    i_8_59_1400_0, i_8_59_1487_0, i_8_59_1538_0, i_8_59_1546_0,
    i_8_59_1552_0, i_8_59_1559_0, i_8_59_1631_0, i_8_59_1637_0,
    i_8_59_1666_0, i_8_59_1675_0, i_8_59_1679_0, i_8_59_1681_0,
    i_8_59_1682_0, i_8_59_1687_0, i_8_59_1697_0, i_8_59_1701_0,
    i_8_59_1755_0, i_8_59_1757_0, i_8_59_1770_0, i_8_59_1772_0,
    i_8_59_1784_0, i_8_59_1789_0, i_8_59_1840_0, i_8_59_1882_0,
    i_8_59_1885_0, i_8_59_1904_0, i_8_59_1910_0, i_8_59_1918_0,
    i_8_59_1960_0, i_8_59_1984_0, i_8_59_1990_0, i_8_59_1994_0,
    i_8_59_1995_0, i_8_59_2033_0, i_8_59_2075_0, i_8_59_2099_0,
    i_8_59_2108_0, i_8_59_2136_0, i_8_59_2146_0, i_8_59_2156_0,
    i_8_59_2224_0, i_8_59_2233_0, i_8_59_2241_0, i_8_59_2260_0;
  output o_8_59_0_0;
  assign o_8_59_0_0 = 0;
endmodule



// Benchmark "kernel_8_60" written by ABC on Sun Jul 19 10:04:02 2020

module kernel_8_60 ( 
    i_8_60_25_0, i_8_60_41_0, i_8_60_44_0, i_8_60_88_0, i_8_60_116_0,
    i_8_60_248_0, i_8_60_283_0, i_8_60_363_0, i_8_60_365_0, i_8_60_389_0,
    i_8_60_400_0, i_8_60_419_0, i_8_60_422_0, i_8_60_430_0, i_8_60_472_0,
    i_8_60_473_0, i_8_60_493_0, i_8_60_508_0, i_8_60_517_0, i_8_60_527_0,
    i_8_60_574_0, i_8_60_575_0, i_8_60_580_0, i_8_60_581_0, i_8_60_592_0,
    i_8_60_593_0, i_8_60_604_0, i_8_60_608_0, i_8_60_661_0, i_8_60_679_0,
    i_8_60_680_0, i_8_60_693_0, i_8_60_697_0, i_8_60_751_0, i_8_60_752_0,
    i_8_60_781_0, i_8_60_824_0, i_8_60_833_0, i_8_60_839_0, i_8_60_841_0,
    i_8_60_848_0, i_8_60_881_0, i_8_60_882_0, i_8_60_886_0, i_8_60_895_0,
    i_8_60_955_0, i_8_60_1036_0, i_8_60_1040_0, i_8_60_1103_0,
    i_8_60_1111_0, i_8_60_1129_0, i_8_60_1184_0, i_8_60_1238_0,
    i_8_60_1241_0, i_8_60_1318_0, i_8_60_1325_0, i_8_60_1330_0,
    i_8_60_1337_0, i_8_60_1353_0, i_8_60_1358_0, i_8_60_1363_0,
    i_8_60_1364_0, i_8_60_1427_0, i_8_60_1436_0, i_8_60_1444_0,
    i_8_60_1480_0, i_8_60_1481_0, i_8_60_1490_0, i_8_60_1532_0,
    i_8_60_1552_0, i_8_60_1633_0, i_8_60_1651_0, i_8_60_1664_0,
    i_8_60_1682_0, i_8_60_1694_0, i_8_60_1697_0, i_8_60_1706_0,
    i_8_60_1733_0, i_8_60_1751_0, i_8_60_1772_0, i_8_60_1774_0,
    i_8_60_1775_0, i_8_60_1781_0, i_8_60_1784_0, i_8_60_1787_0,
    i_8_60_1790_0, i_8_60_1810_0, i_8_60_1855_0, i_8_60_1858_0,
    i_8_60_1859_0, i_8_60_1867_0, i_8_60_1877_0, i_8_60_1913_0,
    i_8_60_1975_0, i_8_60_1978_0, i_8_60_1997_0, i_8_60_2137_0,
    i_8_60_2150_0, i_8_60_2177_0, i_8_60_2249_0,
    o_8_60_0_0  );
  input  i_8_60_25_0, i_8_60_41_0, i_8_60_44_0, i_8_60_88_0,
    i_8_60_116_0, i_8_60_248_0, i_8_60_283_0, i_8_60_363_0, i_8_60_365_0,
    i_8_60_389_0, i_8_60_400_0, i_8_60_419_0, i_8_60_422_0, i_8_60_430_0,
    i_8_60_472_0, i_8_60_473_0, i_8_60_493_0, i_8_60_508_0, i_8_60_517_0,
    i_8_60_527_0, i_8_60_574_0, i_8_60_575_0, i_8_60_580_0, i_8_60_581_0,
    i_8_60_592_0, i_8_60_593_0, i_8_60_604_0, i_8_60_608_0, i_8_60_661_0,
    i_8_60_679_0, i_8_60_680_0, i_8_60_693_0, i_8_60_697_0, i_8_60_751_0,
    i_8_60_752_0, i_8_60_781_0, i_8_60_824_0, i_8_60_833_0, i_8_60_839_0,
    i_8_60_841_0, i_8_60_848_0, i_8_60_881_0, i_8_60_882_0, i_8_60_886_0,
    i_8_60_895_0, i_8_60_955_0, i_8_60_1036_0, i_8_60_1040_0,
    i_8_60_1103_0, i_8_60_1111_0, i_8_60_1129_0, i_8_60_1184_0,
    i_8_60_1238_0, i_8_60_1241_0, i_8_60_1318_0, i_8_60_1325_0,
    i_8_60_1330_0, i_8_60_1337_0, i_8_60_1353_0, i_8_60_1358_0,
    i_8_60_1363_0, i_8_60_1364_0, i_8_60_1427_0, i_8_60_1436_0,
    i_8_60_1444_0, i_8_60_1480_0, i_8_60_1481_0, i_8_60_1490_0,
    i_8_60_1532_0, i_8_60_1552_0, i_8_60_1633_0, i_8_60_1651_0,
    i_8_60_1664_0, i_8_60_1682_0, i_8_60_1694_0, i_8_60_1697_0,
    i_8_60_1706_0, i_8_60_1733_0, i_8_60_1751_0, i_8_60_1772_0,
    i_8_60_1774_0, i_8_60_1775_0, i_8_60_1781_0, i_8_60_1784_0,
    i_8_60_1787_0, i_8_60_1790_0, i_8_60_1810_0, i_8_60_1855_0,
    i_8_60_1858_0, i_8_60_1859_0, i_8_60_1867_0, i_8_60_1877_0,
    i_8_60_1913_0, i_8_60_1975_0, i_8_60_1978_0, i_8_60_1997_0,
    i_8_60_2137_0, i_8_60_2150_0, i_8_60_2177_0, i_8_60_2249_0;
  output o_8_60_0_0;
  assign o_8_60_0_0 = 0;
endmodule



// Benchmark "kernel_8_61" written by ABC on Sun Jul 19 10:04:03 2020

module kernel_8_61 ( 
    i_8_61_11_0, i_8_61_19_0, i_8_61_21_0, i_8_61_22_0, i_8_61_102_0,
    i_8_61_219_0, i_8_61_224_0, i_8_61_265_0, i_8_61_306_0, i_8_61_391_0,
    i_8_61_398_0, i_8_61_404_0, i_8_61_429_0, i_8_61_437_0, i_8_61_464_0,
    i_8_61_487_0, i_8_61_488_0, i_8_61_530_0, i_8_61_538_0, i_8_61_565_0,
    i_8_61_583_0, i_8_61_590_0, i_8_61_601_0, i_8_61_610_0, i_8_61_646_0,
    i_8_61_657_0, i_8_61_661_0, i_8_61_664_0, i_8_61_696_0, i_8_61_709_0,
    i_8_61_749_0, i_8_61_754_0, i_8_61_781_0, i_8_61_783_0, i_8_61_797_0,
    i_8_61_799_0, i_8_61_842_0, i_8_61_858_0, i_8_61_869_0, i_8_61_894_0,
    i_8_61_994_0, i_8_61_1035_0, i_8_61_1065_0, i_8_61_1067_0,
    i_8_61_1137_0, i_8_61_1138_0, i_8_61_1139_0, i_8_61_1189_0,
    i_8_61_1190_0, i_8_61_1202_0, i_8_61_1249_0, i_8_61_1266_0,
    i_8_61_1292_0, i_8_61_1294_0, i_8_61_1298_0, i_8_61_1317_0,
    i_8_61_1363_0, i_8_61_1373_0, i_8_61_1425_0, i_8_61_1443_0,
    i_8_61_1444_0, i_8_61_1446_0, i_8_61_1508_0, i_8_61_1550_0,
    i_8_61_1605_0, i_8_61_1606_0, i_8_61_1607_0, i_8_61_1746_0,
    i_8_61_1747_0, i_8_61_1748_0, i_8_61_1752_0, i_8_61_1759_0,
    i_8_61_1771_0, i_8_61_1773_0, i_8_61_1778_0, i_8_61_1816_0,
    i_8_61_1823_0, i_8_61_1825_0, i_8_61_1831_0, i_8_61_1835_0,
    i_8_61_1841_0, i_8_61_1888_0, i_8_61_1907_0, i_8_61_1951_0,
    i_8_61_1963_0, i_8_61_1966_0, i_8_61_1972_0, i_8_61_1993_0,
    i_8_61_1995_0, i_8_61_2032_0, i_8_61_2043_0, i_8_61_2052_0,
    i_8_61_2053_0, i_8_61_2110_0, i_8_61_2166_0, i_8_61_2169_0,
    i_8_61_2225_0, i_8_61_2237_0, i_8_61_2244_0, i_8_61_2293_0,
    o_8_61_0_0  );
  input  i_8_61_11_0, i_8_61_19_0, i_8_61_21_0, i_8_61_22_0,
    i_8_61_102_0, i_8_61_219_0, i_8_61_224_0, i_8_61_265_0, i_8_61_306_0,
    i_8_61_391_0, i_8_61_398_0, i_8_61_404_0, i_8_61_429_0, i_8_61_437_0,
    i_8_61_464_0, i_8_61_487_0, i_8_61_488_0, i_8_61_530_0, i_8_61_538_0,
    i_8_61_565_0, i_8_61_583_0, i_8_61_590_0, i_8_61_601_0, i_8_61_610_0,
    i_8_61_646_0, i_8_61_657_0, i_8_61_661_0, i_8_61_664_0, i_8_61_696_0,
    i_8_61_709_0, i_8_61_749_0, i_8_61_754_0, i_8_61_781_0, i_8_61_783_0,
    i_8_61_797_0, i_8_61_799_0, i_8_61_842_0, i_8_61_858_0, i_8_61_869_0,
    i_8_61_894_0, i_8_61_994_0, i_8_61_1035_0, i_8_61_1065_0,
    i_8_61_1067_0, i_8_61_1137_0, i_8_61_1138_0, i_8_61_1139_0,
    i_8_61_1189_0, i_8_61_1190_0, i_8_61_1202_0, i_8_61_1249_0,
    i_8_61_1266_0, i_8_61_1292_0, i_8_61_1294_0, i_8_61_1298_0,
    i_8_61_1317_0, i_8_61_1363_0, i_8_61_1373_0, i_8_61_1425_0,
    i_8_61_1443_0, i_8_61_1444_0, i_8_61_1446_0, i_8_61_1508_0,
    i_8_61_1550_0, i_8_61_1605_0, i_8_61_1606_0, i_8_61_1607_0,
    i_8_61_1746_0, i_8_61_1747_0, i_8_61_1748_0, i_8_61_1752_0,
    i_8_61_1759_0, i_8_61_1771_0, i_8_61_1773_0, i_8_61_1778_0,
    i_8_61_1816_0, i_8_61_1823_0, i_8_61_1825_0, i_8_61_1831_0,
    i_8_61_1835_0, i_8_61_1841_0, i_8_61_1888_0, i_8_61_1907_0,
    i_8_61_1951_0, i_8_61_1963_0, i_8_61_1966_0, i_8_61_1972_0,
    i_8_61_1993_0, i_8_61_1995_0, i_8_61_2032_0, i_8_61_2043_0,
    i_8_61_2052_0, i_8_61_2053_0, i_8_61_2110_0, i_8_61_2166_0,
    i_8_61_2169_0, i_8_61_2225_0, i_8_61_2237_0, i_8_61_2244_0,
    i_8_61_2293_0;
  output o_8_61_0_0;
  assign o_8_61_0_0 = 0;
endmodule



// Benchmark "kernel_8_62" written by ABC on Sun Jul 19 10:04:05 2020

module kernel_8_62 ( 
    i_8_62_35_0, i_8_62_61_0, i_8_62_96_0, i_8_62_97_0, i_8_62_258_0,
    i_8_62_325_0, i_8_62_328_0, i_8_62_331_0, i_8_62_367_0, i_8_62_372_0,
    i_8_62_381_0, i_8_62_382_0, i_8_62_458_0, i_8_62_465_0, i_8_62_467_0,
    i_8_62_487_0, i_8_62_504_0, i_8_62_525_0, i_8_62_552_0, i_8_62_586_0,
    i_8_62_590_0, i_8_62_610_0, i_8_62_630_0, i_8_62_632_0, i_8_62_633_0,
    i_8_62_637_0, i_8_62_661_0, i_8_62_664_0, i_8_62_693_0, i_8_62_694_0,
    i_8_62_698_0, i_8_62_762_0, i_8_62_763_0, i_8_62_768_0, i_8_62_790_0,
    i_8_62_855_0, i_8_62_876_0, i_8_62_877_0, i_8_62_879_0, i_8_62_995_0,
    i_8_62_998_0, i_8_62_1137_0, i_8_62_1195_0, i_8_62_1236_0,
    i_8_62_1237_0, i_8_62_1239_0, i_8_62_1240_0, i_8_62_1261_0,
    i_8_62_1264_0, i_8_62_1285_0, i_8_62_1296_0, i_8_62_1297_0,
    i_8_62_1299_0, i_8_62_1333_0, i_8_62_1369_0, i_8_62_1396_0,
    i_8_62_1399_0, i_8_62_1410_0, i_8_62_1489_0, i_8_62_1535_0,
    i_8_62_1536_0, i_8_62_1538_0, i_8_62_1591_0, i_8_62_1599_0,
    i_8_62_1600_0, i_8_62_1602_0, i_8_62_1605_0, i_8_62_1629_0,
    i_8_62_1630_0, i_8_62_1704_0, i_8_62_1722_0, i_8_62_1744_0,
    i_8_62_1746_0, i_8_62_1791_0, i_8_62_1792_0, i_8_62_1795_0,
    i_8_62_1842_0, i_8_62_1843_0, i_8_62_1854_0, i_8_62_1855_0,
    i_8_62_1900_0, i_8_62_1903_0, i_8_62_1915_0, i_8_62_1947_0,
    i_8_62_1951_0, i_8_62_1969_0, i_8_62_2004_0, i_8_62_2047_0,
    i_8_62_2146_0, i_8_62_2154_0, i_8_62_2155_0, i_8_62_2156_0,
    i_8_62_2194_0, i_8_62_2218_0, i_8_62_2233_0, i_8_62_2246_0,
    i_8_62_2263_0, i_8_62_2264_0, i_8_62_2298_0, i_8_62_2299_0,
    o_8_62_0_0  );
  input  i_8_62_35_0, i_8_62_61_0, i_8_62_96_0, i_8_62_97_0,
    i_8_62_258_0, i_8_62_325_0, i_8_62_328_0, i_8_62_331_0, i_8_62_367_0,
    i_8_62_372_0, i_8_62_381_0, i_8_62_382_0, i_8_62_458_0, i_8_62_465_0,
    i_8_62_467_0, i_8_62_487_0, i_8_62_504_0, i_8_62_525_0, i_8_62_552_0,
    i_8_62_586_0, i_8_62_590_0, i_8_62_610_0, i_8_62_630_0, i_8_62_632_0,
    i_8_62_633_0, i_8_62_637_0, i_8_62_661_0, i_8_62_664_0, i_8_62_693_0,
    i_8_62_694_0, i_8_62_698_0, i_8_62_762_0, i_8_62_763_0, i_8_62_768_0,
    i_8_62_790_0, i_8_62_855_0, i_8_62_876_0, i_8_62_877_0, i_8_62_879_0,
    i_8_62_995_0, i_8_62_998_0, i_8_62_1137_0, i_8_62_1195_0,
    i_8_62_1236_0, i_8_62_1237_0, i_8_62_1239_0, i_8_62_1240_0,
    i_8_62_1261_0, i_8_62_1264_0, i_8_62_1285_0, i_8_62_1296_0,
    i_8_62_1297_0, i_8_62_1299_0, i_8_62_1333_0, i_8_62_1369_0,
    i_8_62_1396_0, i_8_62_1399_0, i_8_62_1410_0, i_8_62_1489_0,
    i_8_62_1535_0, i_8_62_1536_0, i_8_62_1538_0, i_8_62_1591_0,
    i_8_62_1599_0, i_8_62_1600_0, i_8_62_1602_0, i_8_62_1605_0,
    i_8_62_1629_0, i_8_62_1630_0, i_8_62_1704_0, i_8_62_1722_0,
    i_8_62_1744_0, i_8_62_1746_0, i_8_62_1791_0, i_8_62_1792_0,
    i_8_62_1795_0, i_8_62_1842_0, i_8_62_1843_0, i_8_62_1854_0,
    i_8_62_1855_0, i_8_62_1900_0, i_8_62_1903_0, i_8_62_1915_0,
    i_8_62_1947_0, i_8_62_1951_0, i_8_62_1969_0, i_8_62_2004_0,
    i_8_62_2047_0, i_8_62_2146_0, i_8_62_2154_0, i_8_62_2155_0,
    i_8_62_2156_0, i_8_62_2194_0, i_8_62_2218_0, i_8_62_2233_0,
    i_8_62_2246_0, i_8_62_2263_0, i_8_62_2264_0, i_8_62_2298_0,
    i_8_62_2299_0;
  output o_8_62_0_0;
  assign o_8_62_0_0 = ~((~i_8_62_1296_0 & ((~i_8_62_1630_0 & ((~i_8_62_61_0 & ((~i_8_62_331_0 & i_8_62_879_0 & ~i_8_62_998_0 & ~i_8_62_1236_0 & ~i_8_62_1239_0 & ~i_8_62_1299_0 & ~i_8_62_1591_0 & ~i_8_62_1602_0 & ~i_8_62_1795_0 & ~i_8_62_2047_0) | (~i_8_62_467_0 & ~i_8_62_552_0 & ~i_8_62_661_0 & ~i_8_62_1240_0 & ~i_8_62_1297_0 & ~i_8_62_1704_0 & ~i_8_62_1843_0 & ~i_8_62_1915_0 & ~i_8_62_1969_0 & ~i_8_62_2218_0))) | (i_8_62_367_0 & ~i_8_62_465_0 & ~i_8_62_467_0 & ~i_8_62_762_0 & ~i_8_62_995_0 & ~i_8_62_1722_0 & ~i_8_62_1947_0 & ~i_8_62_2194_0 & ~i_8_62_2246_0 & ~i_8_62_2298_0))) | (~i_8_62_1333_0 & ((~i_8_62_467_0 & ((~i_8_62_637_0 & ~i_8_62_1236_0 & ~i_8_62_1237_0 & ~i_8_62_1239_0 & ~i_8_62_1264_0 & ~i_8_62_1396_0 & ~i_8_62_1599_0 & ~i_8_62_1744_0 & ~i_8_62_1947_0 & ~i_8_62_1951_0) | (~i_8_62_465_0 & ~i_8_62_610_0 & ~i_8_62_1240_0 & ~i_8_62_1600_0 & ~i_8_62_1602_0 & ~i_8_62_1704_0 & ~i_8_62_1792_0 & ~i_8_62_1842_0 & ~i_8_62_2047_0 & ~i_8_62_2299_0))) | (~i_8_62_1951_0 & ~i_8_62_2298_0 & ((~i_8_62_458_0 & ~i_8_62_693_0 & ~i_8_62_1239_0 & ~i_8_62_1285_0 & i_8_62_1630_0 & ~i_8_62_1969_0) | (i_8_62_525_0 & ~i_8_62_637_0 & ~i_8_62_1264_0 & ~i_8_62_1297_0 & ~i_8_62_1629_0 & ~i_8_62_1915_0 & i_8_62_1947_0 & ~i_8_62_2047_0 & ~i_8_62_2146_0))))) | (~i_8_62_465_0 & ~i_8_62_632_0 & ~i_8_62_1396_0 & ~i_8_62_1536_0 & ~i_8_62_1791_0 & ((~i_8_62_504_0 & ~i_8_62_1195_0 & ~i_8_62_1261_0 & ~i_8_62_1299_0 & ~i_8_62_1591_0 & ~i_8_62_1843_0 & ~i_8_62_2047_0) | (~i_8_62_372_0 & ~i_8_62_610_0 & ~i_8_62_633_0 & ~i_8_62_1410_0 & ~i_8_62_1599_0 & ~i_8_62_1704_0 & ~i_8_62_1722_0 & ~i_8_62_1854_0 & ~i_8_62_1969_0 & ~i_8_62_2298_0))) | (~i_8_62_1746_0 & ((~i_8_62_637_0 & ~i_8_62_876_0 & ~i_8_62_1239_0 & ~i_8_62_1297_0 & ~i_8_62_1410_0 & ~i_8_62_1538_0 & ~i_8_62_1599_0 & ~i_8_62_1792_0 & ~i_8_62_1915_0 & ~i_8_62_2218_0) | (~i_8_62_768_0 & ~i_8_62_1285_0 & i_8_62_1903_0 & ~i_8_62_2298_0))))) | (~i_8_62_2194_0 & ((i_8_62_328_0 & ((i_8_62_661_0 & ~i_8_62_1236_0 & ~i_8_62_1602_0 & ~i_8_62_1722_0 & ~i_8_62_1792_0 & ~i_8_62_1915_0) | (~i_8_62_698_0 & i_8_62_768_0 & ~i_8_62_1333_0 & ~i_8_62_1410_0 & ~i_8_62_1951_0))) | (~i_8_62_465_0 & ((i_8_62_610_0 & i_8_62_877_0 & i_8_62_1285_0 & ~i_8_62_1410_0 & ~i_8_62_1535_0 & ~i_8_62_1599_0 & ~i_8_62_1903_0 & ~i_8_62_2298_0) | (~i_8_62_35_0 & ~i_8_62_637_0 & ~i_8_62_1239_0 & ~i_8_62_1261_0 & ~i_8_62_1285_0 & ~i_8_62_1297_0 & ~i_8_62_1299_0 & ~i_8_62_1536_0 & ~i_8_62_1602_0 & ~i_8_62_1915_0 & ~i_8_62_2146_0 & ~i_8_62_2246_0 & ~i_8_62_2299_0))) | (~i_8_62_328_0 & ~i_8_62_633_0 & i_8_62_664_0 & ~i_8_62_763_0 & ~i_8_62_855_0 & ~i_8_62_1261_0 & ~i_8_62_1410_0 & ~i_8_62_1489_0 & ~i_8_62_1704_0 & ~i_8_62_1744_0 & ~i_8_62_1791_0 & ~i_8_62_2246_0))) | (~i_8_62_610_0 & ((~i_8_62_372_0 & ((~i_8_62_1239_0 & ~i_8_62_1264_0 & i_8_62_458_0 & ~i_8_62_698_0) | (~i_8_62_694_0 & i_8_62_877_0 & ~i_8_62_1399_0 & ~i_8_62_1410_0 & ~i_8_62_1536_0 & ~i_8_62_1602_0 & ~i_8_62_1629_0 & ~i_8_62_1791_0))) | (i_8_62_381_0 & ~i_8_62_487_0 & ~i_8_62_586_0 & ~i_8_62_998_0 & ~i_8_62_1261_0 & ~i_8_62_1600_0 & ~i_8_62_1792_0 & ~i_8_62_1951_0 & ~i_8_62_2218_0 & ~i_8_62_2233_0))) | (~i_8_62_504_0 & ((~i_8_62_762_0 & ((~i_8_62_1915_0 & ((~i_8_62_465_0 & ((~i_8_62_552_0 & ~i_8_62_632_0 & ~i_8_62_1297_0 & i_8_62_1410_0 & ~i_8_62_1591_0 & ~i_8_62_1599_0 & ~i_8_62_1722_0 & ~i_8_62_1746_0 & ~i_8_62_1795_0) | (i_8_62_661_0 & i_8_62_877_0 & ~i_8_62_1369_0 & ~i_8_62_1538_0 & ~i_8_62_1704_0 & ~i_8_62_1792_0 & ~i_8_62_2298_0))) | (~i_8_62_586_0 & ~i_8_62_630_0 & ~i_8_62_1396_0 & ~i_8_62_1489_0 & ~i_8_62_1538_0 & ~i_8_62_1600_0 & ~i_8_62_1842_0 & ~i_8_62_1969_0 & ~i_8_62_2246_0))) | (~i_8_62_35_0 & ~i_8_62_552_0 & ~i_8_62_586_0 & ~i_8_62_632_0 & ~i_8_62_763_0 & ~i_8_62_1261_0 & ~i_8_62_1333_0 & ~i_8_62_1795_0 & ~i_8_62_1947_0 & ~i_8_62_2154_0 & ~i_8_62_2298_0 & ~i_8_62_2299_0))) | (~i_8_62_1237_0 & ((~i_8_62_552_0 & ~i_8_62_630_0 & ((~i_8_62_458_0 & ~i_8_62_1240_0 & ~i_8_62_1261_0 & ~i_8_62_1264_0 & ~i_8_62_1600_0 & ~i_8_62_1842_0 & ~i_8_62_1951_0) | (~i_8_62_586_0 & i_8_62_664_0 & ~i_8_62_1410_0 & ~i_8_62_2298_0))) | (~i_8_62_328_0 & ~i_8_62_855_0 & i_8_62_1264_0 & ~i_8_62_1536_0 & ~i_8_62_1599_0 & ~i_8_62_1630_0 & ~i_8_62_1843_0 & ~i_8_62_1969_0 & ~i_8_62_2263_0))))) | (~i_8_62_1951_0 & ((~i_8_62_35_0 & ((~i_8_62_1237_0 & ~i_8_62_1240_0 & ~i_8_62_1399_0 & ~i_8_62_1536_0 & i_8_62_1591_0) | (i_8_62_367_0 & ~i_8_62_382_0 & ~i_8_62_467_0 & ~i_8_62_487_0 & ~i_8_62_693_0 & ~i_8_62_763_0 & ~i_8_62_1195_0 & ~i_8_62_1297_0 & ~i_8_62_1600_0 & ~i_8_62_1744_0 & ~i_8_62_1746_0))) | (~i_8_62_633_0 & i_8_62_698_0 & ~i_8_62_768_0 & ~i_8_62_855_0 & ~i_8_62_1297_0 & ~i_8_62_1591_0 & ~i_8_62_1600_0 & ~i_8_62_1795_0) | (~i_8_62_1792_0 & ~i_8_62_1842_0 & ~i_8_62_1900_0 & i_8_62_1947_0 & ~i_8_62_2146_0 & i_8_62_2155_0 & ~i_8_62_2156_0 & ~i_8_62_2218_0 & ~i_8_62_2233_0 & ~i_8_62_2298_0))) | (~i_8_62_465_0 & ((i_8_62_61_0 & ~i_8_62_467_0 & i_8_62_763_0 & ~i_8_62_1297_0 & ~i_8_62_1396_0 & ~i_8_62_1599_0 & ~i_8_62_1600_0 & ~i_8_62_1722_0) | (i_8_62_487_0 & ~i_8_62_630_0 & ~i_8_62_633_0 & ~i_8_62_855_0 & ~i_8_62_1237_0 & ~i_8_62_1240_0 & ~i_8_62_1369_0 & ~i_8_62_2155_0 & ~i_8_62_2298_0))) | (~i_8_62_2218_0 & ((~i_8_62_467_0 & ((~i_8_62_525_0 & ~i_8_62_552_0 & ~i_8_62_633_0 & ~i_8_62_876_0 & ~i_8_62_1261_0 & ~i_8_62_1297_0 & ~i_8_62_1399_0 & ~i_8_62_1744_0 & ~i_8_62_1915_0) | (~i_8_62_328_0 & i_8_62_664_0 & ~i_8_62_693_0 & ~i_8_62_855_0 & ~i_8_62_1536_0 & ~i_8_62_1842_0 & ~i_8_62_2246_0))) | (~i_8_62_633_0 & i_8_62_698_0 & ~i_8_62_1299_0 & ~i_8_62_1630_0 & ~i_8_62_2047_0 & i_8_62_2156_0))) | (~i_8_62_328_0 & ~i_8_62_998_0 & ~i_8_62_1591_0 & ((i_8_62_381_0 & i_8_62_382_0 & ~i_8_62_633_0 & ~i_8_62_763_0 & ~i_8_62_1261_0 & ~i_8_62_1842_0 & ~i_8_62_1915_0 & ~i_8_62_2156_0) | (~i_8_62_325_0 & ~i_8_62_525_0 & ~i_8_62_552_0 & ~i_8_62_762_0 & ~i_8_62_1237_0 & ~i_8_62_1297_0 & ~i_8_62_1333_0 & ~i_8_62_1410_0 & ~i_8_62_1599_0 & ~i_8_62_1744_0 & ~i_8_62_1792_0 & ~i_8_62_1843_0 & ~i_8_62_2047_0 & ~i_8_62_2246_0))) | (i_8_62_487_0 & ((~i_8_62_586_0 & i_8_62_876_0 & ~i_8_62_1630_0) | (~i_8_62_525_0 & ~i_8_62_1746_0 & i_8_62_1903_0))) | (~i_8_62_2233_0 & ((i_8_62_1137_0 & ~i_8_62_1264_0 & ~i_8_62_1297_0 & ~i_8_62_1399_0 & ~i_8_62_1792_0 & ~i_8_62_1842_0 & ~i_8_62_1410_0 & ~i_8_62_1538_0) | (~i_8_62_258_0 & i_8_62_325_0 & i_8_62_694_0 & ~i_8_62_1299_0 & ~i_8_62_1535_0 & ~i_8_62_1629_0 & ~i_8_62_2156_0 & ~i_8_62_2298_0))) | (~i_8_62_630_0 & i_8_62_633_0 & ~i_8_62_637_0 & ~i_8_62_1396_0 & ~i_8_62_1605_0 & i_8_62_1947_0 & ~i_8_62_2298_0));
endmodule



// Benchmark "kernel_8_63" written by ABC on Sun Jul 19 10:04:06 2020

module kernel_8_63 ( 
    i_8_63_26_0, i_8_63_77_0, i_8_63_89_0, i_8_63_160_0, i_8_63_161_0,
    i_8_63_224_0, i_8_63_259_0, i_8_63_286_0, i_8_63_296_0, i_8_63_312_0,
    i_8_63_337_0, i_8_63_349_0, i_8_63_367_0, i_8_63_404_0, i_8_63_422_0,
    i_8_63_457_0, i_8_63_485_0, i_8_63_525_0, i_8_63_526_0, i_8_63_556_0,
    i_8_63_606_0, i_8_63_628_0, i_8_63_636_0, i_8_63_682_0, i_8_63_694_0,
    i_8_63_696_0, i_8_63_718_0, i_8_63_763_0, i_8_63_818_0, i_8_63_843_0,
    i_8_63_844_0, i_8_63_872_0, i_8_63_898_0, i_8_63_926_0, i_8_63_951_0,
    i_8_63_952_0, i_8_63_953_0, i_8_63_958_0, i_8_63_980_0, i_8_63_1016_0,
    i_8_63_1033_0, i_8_63_1086_0, i_8_63_1106_0, i_8_63_1114_0,
    i_8_63_1151_0, i_8_63_1222_0, i_8_63_1223_0, i_8_63_1273_0,
    i_8_63_1274_0, i_8_63_1282_0, i_8_63_1286_0, i_8_63_1314_0,
    i_8_63_1324_0, i_8_63_1328_0, i_8_63_1393_0, i_8_63_1404_0,
    i_8_63_1411_0, i_8_63_1437_0, i_8_63_1447_0, i_8_63_1457_0,
    i_8_63_1471_0, i_8_63_1484_0, i_8_63_1524_0, i_8_63_1528_0,
    i_8_63_1534_0, i_8_63_1537_0, i_8_63_1546_0, i_8_63_1547_0,
    i_8_63_1574_0, i_8_63_1582_0, i_8_63_1591_0, i_8_63_1628_0,
    i_8_63_1636_0, i_8_63_1655_0, i_8_63_1658_0, i_8_63_1672_0,
    i_8_63_1690_0, i_8_63_1750_0, i_8_63_1753_0, i_8_63_1807_0,
    i_8_63_1815_0, i_8_63_1823_0, i_8_63_1825_0, i_8_63_1834_0,
    i_8_63_1840_0, i_8_63_1861_0, i_8_63_1870_0, i_8_63_1880_0,
    i_8_63_1888_0, i_8_63_1903_0, i_8_63_1905_0, i_8_63_1906_0,
    i_8_63_1907_0, i_8_63_1975_0, i_8_63_1986_0, i_8_63_2005_0,
    i_8_63_2049_0, i_8_63_2051_0, i_8_63_2060_0, i_8_63_2274_0,
    o_8_63_0_0  );
  input  i_8_63_26_0, i_8_63_77_0, i_8_63_89_0, i_8_63_160_0,
    i_8_63_161_0, i_8_63_224_0, i_8_63_259_0, i_8_63_286_0, i_8_63_296_0,
    i_8_63_312_0, i_8_63_337_0, i_8_63_349_0, i_8_63_367_0, i_8_63_404_0,
    i_8_63_422_0, i_8_63_457_0, i_8_63_485_0, i_8_63_525_0, i_8_63_526_0,
    i_8_63_556_0, i_8_63_606_0, i_8_63_628_0, i_8_63_636_0, i_8_63_682_0,
    i_8_63_694_0, i_8_63_696_0, i_8_63_718_0, i_8_63_763_0, i_8_63_818_0,
    i_8_63_843_0, i_8_63_844_0, i_8_63_872_0, i_8_63_898_0, i_8_63_926_0,
    i_8_63_951_0, i_8_63_952_0, i_8_63_953_0, i_8_63_958_0, i_8_63_980_0,
    i_8_63_1016_0, i_8_63_1033_0, i_8_63_1086_0, i_8_63_1106_0,
    i_8_63_1114_0, i_8_63_1151_0, i_8_63_1222_0, i_8_63_1223_0,
    i_8_63_1273_0, i_8_63_1274_0, i_8_63_1282_0, i_8_63_1286_0,
    i_8_63_1314_0, i_8_63_1324_0, i_8_63_1328_0, i_8_63_1393_0,
    i_8_63_1404_0, i_8_63_1411_0, i_8_63_1437_0, i_8_63_1447_0,
    i_8_63_1457_0, i_8_63_1471_0, i_8_63_1484_0, i_8_63_1524_0,
    i_8_63_1528_0, i_8_63_1534_0, i_8_63_1537_0, i_8_63_1546_0,
    i_8_63_1547_0, i_8_63_1574_0, i_8_63_1582_0, i_8_63_1591_0,
    i_8_63_1628_0, i_8_63_1636_0, i_8_63_1655_0, i_8_63_1658_0,
    i_8_63_1672_0, i_8_63_1690_0, i_8_63_1750_0, i_8_63_1753_0,
    i_8_63_1807_0, i_8_63_1815_0, i_8_63_1823_0, i_8_63_1825_0,
    i_8_63_1834_0, i_8_63_1840_0, i_8_63_1861_0, i_8_63_1870_0,
    i_8_63_1880_0, i_8_63_1888_0, i_8_63_1903_0, i_8_63_1905_0,
    i_8_63_1906_0, i_8_63_1907_0, i_8_63_1975_0, i_8_63_1986_0,
    i_8_63_2005_0, i_8_63_2049_0, i_8_63_2051_0, i_8_63_2060_0,
    i_8_63_2274_0;
  output o_8_63_0_0;
  assign o_8_63_0_0 = 0;
endmodule



// Benchmark "kernel_8_64" written by ABC on Sun Jul 19 10:04:07 2020

module kernel_8_64 ( 
    i_8_64_12_0, i_8_64_13_0, i_8_64_62_0, i_8_64_75_0, i_8_64_89_0,
    i_8_64_129_0, i_8_64_130_0, i_8_64_193_0, i_8_64_223_0, i_8_64_363_0,
    i_8_64_365_0, i_8_64_366_0, i_8_64_390_0, i_8_64_426_0, i_8_64_499_0,
    i_8_64_522_0, i_8_64_526_0, i_8_64_528_0, i_8_64_530_0, i_8_64_591_0,
    i_8_64_593_0, i_8_64_604_0, i_8_64_609_0, i_8_64_610_0, i_8_64_627_0,
    i_8_64_637_0, i_8_64_654_0, i_8_64_660_0, i_8_64_661_0, i_8_64_665_0,
    i_8_64_678_0, i_8_64_681_0, i_8_64_705_0, i_8_64_708_0, i_8_64_718_0,
    i_8_64_815_0, i_8_64_834_0, i_8_64_835_0, i_8_64_894_0, i_8_64_1032_0,
    i_8_64_1033_0, i_8_64_1078_0, i_8_64_1266_0, i_8_64_1272_0,
    i_8_64_1274_0, i_8_64_1302_0, i_8_64_1308_0, i_8_64_1338_0,
    i_8_64_1339_0, i_8_64_1340_0, i_8_64_1398_0, i_8_64_1403_0,
    i_8_64_1434_0, i_8_64_1439_0, i_8_64_1449_0, i_8_64_1461_0,
    i_8_64_1464_0, i_8_64_1507_0, i_8_64_1547_0, i_8_64_1599_0,
    i_8_64_1601_0, i_8_64_1625_0, i_8_64_1627_0, i_8_64_1636_0,
    i_8_64_1637_0, i_8_64_1641_0, i_8_64_1643_0, i_8_64_1662_0,
    i_8_64_1731_0, i_8_64_1734_0, i_8_64_1749_0, i_8_64_1779_0,
    i_8_64_1780_0, i_8_64_1787_0, i_8_64_1788_0, i_8_64_1789_0,
    i_8_64_1790_0, i_8_64_1804_0, i_8_64_1851_0, i_8_64_1853_0,
    i_8_64_1857_0, i_8_64_1860_0, i_8_64_1861_0, i_8_64_1866_0,
    i_8_64_1867_0, i_8_64_1869_0, i_8_64_1879_0, i_8_64_1905_0,
    i_8_64_1906_0, i_8_64_1907_0, i_8_64_1951_0, i_8_64_1952_0,
    i_8_64_2032_0, i_8_64_2040_0, i_8_64_2092_0, i_8_64_2093_0,
    i_8_64_2158_0, i_8_64_2215_0, i_8_64_2242_0, i_8_64_2249_0,
    o_8_64_0_0  );
  input  i_8_64_12_0, i_8_64_13_0, i_8_64_62_0, i_8_64_75_0, i_8_64_89_0,
    i_8_64_129_0, i_8_64_130_0, i_8_64_193_0, i_8_64_223_0, i_8_64_363_0,
    i_8_64_365_0, i_8_64_366_0, i_8_64_390_0, i_8_64_426_0, i_8_64_499_0,
    i_8_64_522_0, i_8_64_526_0, i_8_64_528_0, i_8_64_530_0, i_8_64_591_0,
    i_8_64_593_0, i_8_64_604_0, i_8_64_609_0, i_8_64_610_0, i_8_64_627_0,
    i_8_64_637_0, i_8_64_654_0, i_8_64_660_0, i_8_64_661_0, i_8_64_665_0,
    i_8_64_678_0, i_8_64_681_0, i_8_64_705_0, i_8_64_708_0, i_8_64_718_0,
    i_8_64_815_0, i_8_64_834_0, i_8_64_835_0, i_8_64_894_0, i_8_64_1032_0,
    i_8_64_1033_0, i_8_64_1078_0, i_8_64_1266_0, i_8_64_1272_0,
    i_8_64_1274_0, i_8_64_1302_0, i_8_64_1308_0, i_8_64_1338_0,
    i_8_64_1339_0, i_8_64_1340_0, i_8_64_1398_0, i_8_64_1403_0,
    i_8_64_1434_0, i_8_64_1439_0, i_8_64_1449_0, i_8_64_1461_0,
    i_8_64_1464_0, i_8_64_1507_0, i_8_64_1547_0, i_8_64_1599_0,
    i_8_64_1601_0, i_8_64_1625_0, i_8_64_1627_0, i_8_64_1636_0,
    i_8_64_1637_0, i_8_64_1641_0, i_8_64_1643_0, i_8_64_1662_0,
    i_8_64_1731_0, i_8_64_1734_0, i_8_64_1749_0, i_8_64_1779_0,
    i_8_64_1780_0, i_8_64_1787_0, i_8_64_1788_0, i_8_64_1789_0,
    i_8_64_1790_0, i_8_64_1804_0, i_8_64_1851_0, i_8_64_1853_0,
    i_8_64_1857_0, i_8_64_1860_0, i_8_64_1861_0, i_8_64_1866_0,
    i_8_64_1867_0, i_8_64_1869_0, i_8_64_1879_0, i_8_64_1905_0,
    i_8_64_1906_0, i_8_64_1907_0, i_8_64_1951_0, i_8_64_1952_0,
    i_8_64_2032_0, i_8_64_2040_0, i_8_64_2092_0, i_8_64_2093_0,
    i_8_64_2158_0, i_8_64_2215_0, i_8_64_2242_0, i_8_64_2249_0;
  output o_8_64_0_0;
  assign o_8_64_0_0 = ~((i_8_64_129_0 & ((~i_8_64_1398_0 & ~i_8_64_1779_0 & ~i_8_64_1780_0 & ~i_8_64_1787_0 & ~i_8_64_1804_0 & ~i_8_64_1952_0) | (~i_8_64_530_0 & ~i_8_64_593_0 & ~i_8_64_678_0 & ~i_8_64_1449_0 & ~i_8_64_1636_0 & ~i_8_64_1637_0 & ~i_8_64_1788_0 & ~i_8_64_2032_0))) | (i_8_64_130_0 & ((~i_8_64_593_0 & ~i_8_64_894_0 & ~i_8_64_1340_0 & ~i_8_64_1780_0) | (i_8_64_365_0 & ~i_8_64_610_0 & i_8_64_1340_0 & i_8_64_1439_0 & ~i_8_64_1636_0 & i_8_64_1952_0 & ~i_8_64_2032_0 & ~i_8_64_2092_0 & ~i_8_64_2242_0))) | (~i_8_64_1338_0 & ((~i_8_64_130_0 & ((~i_8_64_609_0 & ~i_8_64_894_0 & ~i_8_64_1339_0 & i_8_64_1398_0 & ~i_8_64_1599_0 & i_8_64_1749_0 & ~i_8_64_1860_0 & ~i_8_64_1861_0 & ~i_8_64_1866_0) | (~i_8_64_223_0 & ~i_8_64_363_0 & ~i_8_64_366_0 & ~i_8_64_390_0 & ~i_8_64_1403_0 & ~i_8_64_1439_0 & ~i_8_64_1449_0 & ~i_8_64_1627_0 & ~i_8_64_1787_0 & ~i_8_64_2032_0))) | (~i_8_64_678_0 & ((~i_8_64_12_0 & ~i_8_64_62_0 & ~i_8_64_654_0 & ~i_8_64_708_0 & ~i_8_64_894_0 & ~i_8_64_1266_0 & ~i_8_64_1308_0 & ~i_8_64_1547_0 & ~i_8_64_1601_0 & ~i_8_64_1787_0 & ~i_8_64_1790_0) | (i_8_64_499_0 & ~i_8_64_1302_0 & ~i_8_64_1339_0 & ~i_8_64_1340_0 & ~i_8_64_1857_0))) | (~i_8_64_1403_0 & ((~i_8_64_75_0 & ~i_8_64_426_0 & ~i_8_64_661_0 & ~i_8_64_1339_0 & ~i_8_64_1398_0 & ~i_8_64_1439_0 & ~i_8_64_1787_0) | (~i_8_64_1636_0 & i_8_64_1853_0 & ~i_8_64_1869_0))) | (~i_8_64_1789_0 & ((~i_8_64_1434_0 & ~i_8_64_1547_0 & ~i_8_64_2158_0 & i_8_64_2215_0) | (~i_8_64_13_0 & ~i_8_64_193_0 & ~i_8_64_593_0 & ~i_8_64_681_0 & ~i_8_64_894_0 & ~i_8_64_1749_0 & ~i_8_64_2032_0 & ~i_8_64_2249_0))) | (~i_8_64_591_0 & ~i_8_64_604_0 & ~i_8_64_610_0 & ~i_8_64_1274_0 & i_8_64_1731_0))) | (~i_8_64_75_0 & ((~i_8_64_62_0 & ~i_8_64_591_0 & ~i_8_64_604_0 & ~i_8_64_678_0 & ~i_8_64_705_0 & ~i_8_64_1643_0 & ~i_8_64_1779_0 & ~i_8_64_1787_0 & ~i_8_64_1790_0 & ~i_8_64_1952_0) | (~i_8_64_627_0 & ~i_8_64_654_0 & ~i_8_64_665_0 & ~i_8_64_1434_0 & ~i_8_64_1461_0 & ~i_8_64_1749_0 & ~i_8_64_1780_0 & ~i_8_64_1789_0 & ~i_8_64_1853_0 & ~i_8_64_2040_0 & ~i_8_64_2249_0))) | (~i_8_64_223_0 & ((~i_8_64_604_0 & ~i_8_64_610_0 & ~i_8_64_708_0 & ~i_8_64_1302_0 & ~i_8_64_1787_0 & ~i_8_64_1790_0 & ~i_8_64_1340_0 & ~i_8_64_1749_0) | (~i_8_64_593_0 & i_8_64_1434_0 & ~i_8_64_1449_0 & ~i_8_64_1780_0 & ~i_8_64_1853_0 & i_8_64_2158_0))) | (~i_8_64_363_0 & ((i_8_64_530_0 & i_8_64_1601_0) | (i_8_64_526_0 & ~i_8_64_604_0 & ~i_8_64_661_0 & ~i_8_64_1340_0 & ~i_8_64_1599_0 & ~i_8_64_1734_0 & i_8_64_1749_0))) | (~i_8_64_499_0 & ((~i_8_64_660_0 & i_8_64_1731_0 & ~i_8_64_1749_0 & ~i_8_64_1804_0 & ~i_8_64_2158_0) | (~i_8_64_62_0 & i_8_64_526_0 & ~i_8_64_530_0 & ~i_8_64_591_0 & ~i_8_64_1403_0 & ~i_8_64_1449_0 & ~i_8_64_1637_0 & ~i_8_64_2249_0))) | (~i_8_64_681_0 & ((~i_8_64_62_0 & ~i_8_64_637_0 & ~i_8_64_2249_0 & ((~i_8_64_604_0 & ~i_8_64_610_0 & ~i_8_64_1266_0 & ~i_8_64_1302_0 & i_8_64_1780_0) | (~i_8_64_13_0 & ~i_8_64_1339_0 & ~i_8_64_1340_0 & ~i_8_64_1636_0 & i_8_64_1789_0 & ~i_8_64_1951_0 & ~i_8_64_2158_0 & ~i_8_64_2242_0))) | (~i_8_64_1403_0 & ((~i_8_64_604_0 & ~i_8_64_1339_0 & ~i_8_64_1434_0 & i_8_64_1547_0) | (~i_8_64_365_0 & ~i_8_64_661_0 & ~i_8_64_678_0 & ~i_8_64_1461_0 & ~i_8_64_1734_0 & ~i_8_64_1879_0 & i_8_64_2215_0))) | (~i_8_64_12_0 & i_8_64_528_0 & i_8_64_834_0) | (i_8_64_593_0 & ~i_8_64_665_0 & ~i_8_64_1274_0 & ~i_8_64_1627_0 & ~i_8_64_1804_0 & i_8_64_1860_0 & ~i_8_64_1907_0) | (i_8_64_193_0 & ~i_8_64_708_0 & ~i_8_64_1637_0 & i_8_64_1804_0 & ~i_8_64_1952_0))) | (~i_8_64_390_0 & ((~i_8_64_13_0 & ((~i_8_64_366_0 & ~i_8_64_1439_0 & i_8_64_1507_0 & ~i_8_64_1780_0) | (~i_8_64_193_0 & ~i_8_64_609_0 & ~i_8_64_637_0 & i_8_64_678_0 & i_8_64_705_0 & ~i_8_64_1787_0 & ~i_8_64_1951_0 & ~i_8_64_2158_0 & ~i_8_64_2215_0))) | (~i_8_64_604_0 & ~i_8_64_1643_0 & ((~i_8_64_678_0 & ~i_8_64_1340_0 & ~i_8_64_1449_0 & i_8_64_1857_0 & ~i_8_64_2158_0) | (i_8_64_522_0 & ~i_8_64_591_0 & ~i_8_64_660_0 & ~i_8_64_1308_0 & ~i_8_64_2249_0))))) | (~i_8_64_522_0 & ((~i_8_64_654_0 & ~i_8_64_894_0 & ~i_8_64_1547_0 & i_8_64_1641_0 & i_8_64_1780_0 & ~i_8_64_1952_0) | (i_8_64_661_0 & ~i_8_64_678_0 & ~i_8_64_1398_0 & ~i_8_64_1779_0 & ~i_8_64_1787_0 & ~i_8_64_1788_0 & ~i_8_64_2158_0 & ~i_8_64_2249_0))) | (~i_8_64_661_0 & ((~i_8_64_12_0 & ~i_8_64_593_0 & ~i_8_64_678_0 & ~i_8_64_894_0 & ~i_8_64_1266_0 & ~i_8_64_1779_0 & ~i_8_64_1780_0 & ~i_8_64_1787_0 & ~i_8_64_1789_0) | (~i_8_64_1339_0 & ~i_8_64_1398_0 & i_8_64_609_0 & ~i_8_64_1274_0 & ~i_8_64_1636_0 & ~i_8_64_1637_0 & ~i_8_64_1749_0 & ~i_8_64_2249_0))) | (~i_8_64_12_0 & ~i_8_64_678_0 & ((i_8_64_89_0 & ~i_8_64_1340_0) | (i_8_64_426_0 & i_8_64_526_0 & ~i_8_64_609_0 & ~i_8_64_1790_0 & i_8_64_1804_0))) | (~i_8_64_665_0 & ((~i_8_64_426_0 & i_8_64_530_0 & ~i_8_64_1032_0 & ~i_8_64_1398_0 & ~i_8_64_1403_0) | (~i_8_64_1339_0 & ~i_8_64_1340_0 & ~i_8_64_1788_0 & ~i_8_64_1951_0 & i_8_64_2249_0))) | (~i_8_64_1461_0 & ((~i_8_64_637_0 & ~i_8_64_1308_0 & i_8_64_1804_0 & i_8_64_1857_0) | (i_8_64_604_0 & ~i_8_64_660_0 & ~i_8_64_894_0 & ~i_8_64_1636_0 & ~i_8_64_1749_0 & ~i_8_64_1867_0 & ~i_8_64_1907_0 & i_8_64_2242_0 & ~i_8_64_2249_0))) | (~i_8_64_1749_0 & i_8_64_1851_0 & ~i_8_64_1951_0 & ~i_8_64_1952_0) | (i_8_64_1907_0 & ~i_8_64_2032_0 & i_8_64_2215_0));
endmodule



// Benchmark "kernel_8_65" written by ABC on Sun Jul 19 10:04:08 2020

module kernel_8_65 ( 
    i_8_65_43_0, i_8_65_53_0, i_8_65_76_0, i_8_65_127_0, i_8_65_145_0,
    i_8_65_196_0, i_8_65_210_0, i_8_65_284_0, i_8_65_301_0, i_8_65_319_0,
    i_8_65_325_0, i_8_65_328_0, i_8_65_347_0, i_8_65_361_0, i_8_65_384_0,
    i_8_65_390_0, i_8_65_453_0, i_8_65_454_0, i_8_65_508_0, i_8_65_526_0,
    i_8_65_562_0, i_8_65_583_0, i_8_65_599_0, i_8_65_608_0, i_8_65_611_0,
    i_8_65_643_0, i_8_65_656_0, i_8_65_658_0, i_8_65_664_0, i_8_65_695_0,
    i_8_65_697_0, i_8_65_709_0, i_8_65_710_0, i_8_65_775_0, i_8_65_792_0,
    i_8_65_839_0, i_8_65_840_0, i_8_65_895_0, i_8_65_926_0, i_8_65_967_0,
    i_8_65_968_0, i_8_65_1015_0, i_8_65_1074_0, i_8_65_1103_0,
    i_8_65_1106_0, i_8_65_1107_0, i_8_65_1115_0, i_8_65_1126_0,
    i_8_65_1183_0, i_8_65_1204_0, i_8_65_1231_0, i_8_65_1240_0,
    i_8_65_1263_0, i_8_65_1264_0, i_8_65_1267_0, i_8_65_1268_0,
    i_8_65_1286_0, i_8_65_1299_0, i_8_65_1339_0, i_8_65_1365_0,
    i_8_65_1410_0, i_8_65_1436_0, i_8_65_1444_0, i_8_65_1474_0,
    i_8_65_1490_0, i_8_65_1525_0, i_8_65_1546_0, i_8_65_1572_0,
    i_8_65_1603_0, i_8_65_1607_0, i_8_65_1609_0, i_8_65_1669_0,
    i_8_65_1690_0, i_8_65_1749_0, i_8_65_1751_0, i_8_65_1780_0,
    i_8_65_1786_0, i_8_65_1787_0, i_8_65_1806_0, i_8_65_1825_0,
    i_8_65_1886_0, i_8_65_1915_0, i_8_65_1930_0, i_8_65_1948_0,
    i_8_65_1949_0, i_8_65_1950_0, i_8_65_1992_0, i_8_65_1994_0,
    i_8_65_1995_0, i_8_65_2112_0, i_8_65_2142_0, i_8_65_2144_0,
    i_8_65_2147_0, i_8_65_2148_0, i_8_65_2150_0, i_8_65_2212_0,
    i_8_65_2260_0, i_8_65_2272_0, i_8_65_2290_0, i_8_65_2294_0,
    o_8_65_0_0  );
  input  i_8_65_43_0, i_8_65_53_0, i_8_65_76_0, i_8_65_127_0,
    i_8_65_145_0, i_8_65_196_0, i_8_65_210_0, i_8_65_284_0, i_8_65_301_0,
    i_8_65_319_0, i_8_65_325_0, i_8_65_328_0, i_8_65_347_0, i_8_65_361_0,
    i_8_65_384_0, i_8_65_390_0, i_8_65_453_0, i_8_65_454_0, i_8_65_508_0,
    i_8_65_526_0, i_8_65_562_0, i_8_65_583_0, i_8_65_599_0, i_8_65_608_0,
    i_8_65_611_0, i_8_65_643_0, i_8_65_656_0, i_8_65_658_0, i_8_65_664_0,
    i_8_65_695_0, i_8_65_697_0, i_8_65_709_0, i_8_65_710_0, i_8_65_775_0,
    i_8_65_792_0, i_8_65_839_0, i_8_65_840_0, i_8_65_895_0, i_8_65_926_0,
    i_8_65_967_0, i_8_65_968_0, i_8_65_1015_0, i_8_65_1074_0,
    i_8_65_1103_0, i_8_65_1106_0, i_8_65_1107_0, i_8_65_1115_0,
    i_8_65_1126_0, i_8_65_1183_0, i_8_65_1204_0, i_8_65_1231_0,
    i_8_65_1240_0, i_8_65_1263_0, i_8_65_1264_0, i_8_65_1267_0,
    i_8_65_1268_0, i_8_65_1286_0, i_8_65_1299_0, i_8_65_1339_0,
    i_8_65_1365_0, i_8_65_1410_0, i_8_65_1436_0, i_8_65_1444_0,
    i_8_65_1474_0, i_8_65_1490_0, i_8_65_1525_0, i_8_65_1546_0,
    i_8_65_1572_0, i_8_65_1603_0, i_8_65_1607_0, i_8_65_1609_0,
    i_8_65_1669_0, i_8_65_1690_0, i_8_65_1749_0, i_8_65_1751_0,
    i_8_65_1780_0, i_8_65_1786_0, i_8_65_1787_0, i_8_65_1806_0,
    i_8_65_1825_0, i_8_65_1886_0, i_8_65_1915_0, i_8_65_1930_0,
    i_8_65_1948_0, i_8_65_1949_0, i_8_65_1950_0, i_8_65_1992_0,
    i_8_65_1994_0, i_8_65_1995_0, i_8_65_2112_0, i_8_65_2142_0,
    i_8_65_2144_0, i_8_65_2147_0, i_8_65_2148_0, i_8_65_2150_0,
    i_8_65_2212_0, i_8_65_2260_0, i_8_65_2272_0, i_8_65_2290_0,
    i_8_65_2294_0;
  output o_8_65_0_0;
  assign o_8_65_0_0 = 0;
endmodule



// Benchmark "kernel_8_66" written by ABC on Sun Jul 19 10:04:10 2020

module kernel_8_66 ( 
    i_8_66_27_0, i_8_66_30_0, i_8_66_78_0, i_8_66_79_0, i_8_66_114_0,
    i_8_66_165_0, i_8_66_166_0, i_8_66_192_0, i_8_66_193_0, i_8_66_211_0,
    i_8_66_224_0, i_8_66_234_0, i_8_66_237_0, i_8_66_238_0, i_8_66_240_0,
    i_8_66_241_0, i_8_66_301_0, i_8_66_302_0, i_8_66_337_0, i_8_66_338_0,
    i_8_66_346_0, i_8_66_384_0, i_8_66_462_0, i_8_66_476_0, i_8_66_489_0,
    i_8_66_510_0, i_8_66_525_0, i_8_66_591_0, i_8_66_592_0, i_8_66_593_0,
    i_8_66_600_0, i_8_66_602_0, i_8_66_604_0, i_8_66_616_0, i_8_66_617_0,
    i_8_66_658_0, i_8_66_701_0, i_8_66_710_0, i_8_66_717_0, i_8_66_720_0,
    i_8_66_747_0, i_8_66_774_0, i_8_66_787_0, i_8_66_804_0, i_8_66_825_0,
    i_8_66_850_0, i_8_66_864_0, i_8_66_996_0, i_8_66_1047_0, i_8_66_1056_0,
    i_8_66_1120_0, i_8_66_1128_0, i_8_66_1260_0, i_8_66_1279_0,
    i_8_66_1284_0, i_8_66_1292_0, i_8_66_1306_0, i_8_66_1410_0,
    i_8_66_1412_0, i_8_66_1437_0, i_8_66_1438_0, i_8_66_1527_0,
    i_8_66_1528_0, i_8_66_1572_0, i_8_66_1611_0, i_8_66_1624_0,
    i_8_66_1625_0, i_8_66_1632_0, i_8_66_1633_0, i_8_66_1634_0,
    i_8_66_1635_0, i_8_66_1637_0, i_8_66_1653_0, i_8_66_1654_0,
    i_8_66_1655_0, i_8_66_1672_0, i_8_66_1699_0, i_8_66_1754_0,
    i_8_66_1782_0, i_8_66_1824_0, i_8_66_1832_0, i_8_66_1854_0,
    i_8_66_1857_0, i_8_66_1947_0, i_8_66_1983_0, i_8_66_1984_0,
    i_8_66_1992_0, i_8_66_1993_0, i_8_66_1994_0, i_8_66_1997_0,
    i_8_66_2031_0, i_8_66_2040_0, i_8_66_2076_0, i_8_66_2077_0,
    i_8_66_2088_0, i_8_66_2154_0, i_8_66_2212_0, i_8_66_2214_0,
    i_8_66_2259_0, i_8_66_2262_0,
    o_8_66_0_0  );
  input  i_8_66_27_0, i_8_66_30_0, i_8_66_78_0, i_8_66_79_0,
    i_8_66_114_0, i_8_66_165_0, i_8_66_166_0, i_8_66_192_0, i_8_66_193_0,
    i_8_66_211_0, i_8_66_224_0, i_8_66_234_0, i_8_66_237_0, i_8_66_238_0,
    i_8_66_240_0, i_8_66_241_0, i_8_66_301_0, i_8_66_302_0, i_8_66_337_0,
    i_8_66_338_0, i_8_66_346_0, i_8_66_384_0, i_8_66_462_0, i_8_66_476_0,
    i_8_66_489_0, i_8_66_510_0, i_8_66_525_0, i_8_66_591_0, i_8_66_592_0,
    i_8_66_593_0, i_8_66_600_0, i_8_66_602_0, i_8_66_604_0, i_8_66_616_0,
    i_8_66_617_0, i_8_66_658_0, i_8_66_701_0, i_8_66_710_0, i_8_66_717_0,
    i_8_66_720_0, i_8_66_747_0, i_8_66_774_0, i_8_66_787_0, i_8_66_804_0,
    i_8_66_825_0, i_8_66_850_0, i_8_66_864_0, i_8_66_996_0, i_8_66_1047_0,
    i_8_66_1056_0, i_8_66_1120_0, i_8_66_1128_0, i_8_66_1260_0,
    i_8_66_1279_0, i_8_66_1284_0, i_8_66_1292_0, i_8_66_1306_0,
    i_8_66_1410_0, i_8_66_1412_0, i_8_66_1437_0, i_8_66_1438_0,
    i_8_66_1527_0, i_8_66_1528_0, i_8_66_1572_0, i_8_66_1611_0,
    i_8_66_1624_0, i_8_66_1625_0, i_8_66_1632_0, i_8_66_1633_0,
    i_8_66_1634_0, i_8_66_1635_0, i_8_66_1637_0, i_8_66_1653_0,
    i_8_66_1654_0, i_8_66_1655_0, i_8_66_1672_0, i_8_66_1699_0,
    i_8_66_1754_0, i_8_66_1782_0, i_8_66_1824_0, i_8_66_1832_0,
    i_8_66_1854_0, i_8_66_1857_0, i_8_66_1947_0, i_8_66_1983_0,
    i_8_66_1984_0, i_8_66_1992_0, i_8_66_1993_0, i_8_66_1994_0,
    i_8_66_1997_0, i_8_66_2031_0, i_8_66_2040_0, i_8_66_2076_0,
    i_8_66_2077_0, i_8_66_2088_0, i_8_66_2154_0, i_8_66_2212_0,
    i_8_66_2214_0, i_8_66_2259_0, i_8_66_2262_0;
  output o_8_66_0_0;
  assign o_8_66_0_0 = ~((i_8_66_78_0 & ((~i_8_66_114_0 & ~i_8_66_710_0 & ~i_8_66_804_0 & ~i_8_66_825_0 & ~i_8_66_2076_0) | (~i_8_66_237_0 & ~i_8_66_604_0 & ~i_8_66_1611_0 & ~i_8_66_2040_0 & ~i_8_66_2077_0))) | (~i_8_66_1292_0 & ((~i_8_66_27_0 & ((~i_8_66_30_0 & ~i_8_66_1527_0 & ~i_8_66_2262_0 & ((~i_8_66_165_0 & ~i_8_66_489_0 & i_8_66_1284_0 & i_8_66_1438_0 & ~i_8_66_1654_0 & ~i_8_66_1655_0 & ~i_8_66_1824_0 & ~i_8_66_1854_0) | (i_8_66_193_0 & ~i_8_66_240_0 & ~i_8_66_384_0 & ~i_8_66_710_0 & ~i_8_66_720_0 & ~i_8_66_864_0 & ~i_8_66_1260_0 & ~i_8_66_1624_0 & ~i_8_66_2077_0))) | (~i_8_66_238_0 & ~i_8_66_864_0 & i_8_66_1120_0 & ~i_8_66_1279_0 & ~i_8_66_1654_0 & ~i_8_66_1672_0 & ~i_8_66_2259_0))) | (i_8_66_302_0 & ((~i_8_66_337_0 & i_8_66_338_0 & ~i_8_66_617_0 & ~i_8_66_1047_0) | (~i_8_66_238_0 & ~i_8_66_1056_0 & ~i_8_66_1437_0 & ~i_8_66_1625_0 & ~i_8_66_1832_0 & ~i_8_66_1984_0 & ~i_8_66_1993_0))) | (~i_8_66_804_0 & ((i_8_66_224_0 & ~i_8_66_234_0 & ~i_8_66_241_0 & ~i_8_66_701_0 & ~i_8_66_864_0 & ~i_8_66_1412_0 & ~i_8_66_1528_0) | (i_8_66_489_0 & i_8_66_591_0 & ~i_8_66_720_0 & ~i_8_66_1306_0 & ~i_8_66_1438_0 & ~i_8_66_1994_0))) | (~i_8_66_996_0 & ~i_8_66_1625_0 & ~i_8_66_2259_0 & ((~i_8_66_240_0 & ~i_8_66_476_0 & ~i_8_66_617_0 & i_8_66_710_0 & ~i_8_66_1437_0) | (~i_8_66_237_0 & ~i_8_66_864_0 & i_8_66_1128_0 & ~i_8_66_1857_0))) | (i_8_66_338_0 & i_8_66_476_0 & i_8_66_1412_0 & ~i_8_66_1984_0 & i_8_66_1994_0) | (i_8_66_193_0 & ~i_8_66_717_0 & ~i_8_66_774_0 & ~i_8_66_1120_0 & ~i_8_66_1412_0 & ~i_8_66_1611_0 & ~i_8_66_1633_0 & ~i_8_66_1854_0 & ~i_8_66_1983_0 & ~i_8_66_1997_0 & ~i_8_66_2040_0 & ~i_8_66_2076_0))) | (~i_8_66_30_0 & ((~i_8_66_489_0 & i_8_66_850_0 & i_8_66_864_0 & ~i_8_66_1056_0 & ~i_8_66_1306_0) | (~i_8_66_114_0 & ~i_8_66_774_0 & ~i_8_66_1047_0 & ~i_8_66_1260_0 & ~i_8_66_1624_0 & ~i_8_66_1625_0 & ~i_8_66_1632_0 & ~i_8_66_1653_0 & ~i_8_66_1654_0 & i_8_66_1947_0 & ~i_8_66_1983_0 & ~i_8_66_1984_0))) | (~i_8_66_338_0 & ((~i_8_66_27_0 & ~i_8_66_211_0 & ~i_8_66_525_0 & ~i_8_66_1279_0 & ((~i_8_66_114_0 & ~i_8_66_384_0 & i_8_66_616_0 & ~i_8_66_617_0 & ~i_8_66_864_0 & ~i_8_66_1672_0 & ~i_8_66_1832_0 & ~i_8_66_1983_0 & ~i_8_66_2040_0 & ~i_8_66_2088_0) | (~i_8_66_237_0 & ~i_8_66_240_0 & ~i_8_66_1047_0 & ~i_8_66_1611_0 & ~i_8_66_1625_0 & i_8_66_1983_0 & ~i_8_66_2076_0 & ~i_8_66_2214_0))) | (~i_8_66_617_0 & ((~i_8_66_701_0 & ~i_8_66_1260_0 & ((~i_8_66_1625_0 & ((~i_8_66_234_0 & ~i_8_66_1047_0 & ((~i_8_66_238_0 & ~i_8_66_774_0 & i_8_66_1279_0 & ~i_8_66_1854_0) | (~i_8_66_658_0 & ~i_8_66_864_0 & ~i_8_66_1284_0 & ~i_8_66_1437_0 & ~i_8_66_1655_0 & ~i_8_66_1947_0 & ~i_8_66_1984_0 & ~i_8_66_2076_0 & ~i_8_66_2077_0 & ~i_8_66_2154_0 & ~i_8_66_2259_0))) | (~i_8_66_241_0 & ~i_8_66_337_0 & ~i_8_66_658_0 & ~i_8_66_774_0 & ~i_8_66_996_0 & ~i_8_66_1056_0 & ~i_8_66_1437_0 & ~i_8_66_1984_0 & ~i_8_66_2076_0 & ~i_8_66_2212_0 & ~i_8_66_2214_0))) | (~i_8_66_114_0 & ~i_8_66_337_0 & ~i_8_66_616_0 & ~i_8_66_658_0 & ~i_8_66_850_0 & ~i_8_66_864_0 & ~i_8_66_1284_0 & ~i_8_66_1412_0 & ~i_8_66_1528_0 & ~i_8_66_1624_0 & ~i_8_66_1782_0 & ~i_8_66_1857_0 & ~i_8_66_1994_0 & ~i_8_66_2076_0 & ~i_8_66_2259_0))) | (~i_8_66_238_0 & ~i_8_66_337_0 & ~i_8_66_864_0 & ~i_8_66_996_0 & ~i_8_66_1527_0 & ~i_8_66_1611_0 & ~i_8_66_1782_0 & ~i_8_66_1983_0 & i_8_66_1993_0 & ~i_8_66_2212_0 & ~i_8_66_2214_0))) | (~i_8_66_234_0 & ~i_8_66_616_0 & ((~i_8_66_241_0 & i_8_66_301_0 & ~i_8_66_774_0 & ~i_8_66_804_0 & ~i_8_66_1653_0) | (~i_8_66_237_0 & ~i_8_66_346_0 & ~i_8_66_591_0 & ~i_8_66_658_0 & ~i_8_66_701_0 & ~i_8_66_864_0 & ~i_8_66_996_0 & ~i_8_66_1056_0 & ~i_8_66_1260_0 & ~i_8_66_1410_0 & ~i_8_66_1528_0 & ~i_8_66_1625_0 & ~i_8_66_1654_0 & ~i_8_66_1832_0 & ~i_8_66_1854_0 & ~i_8_66_1947_0 & ~i_8_66_1984_0 & ~i_8_66_1994_0))) | (~i_8_66_489_0 & ~i_8_66_1857_0 & ((~i_8_66_166_0 & i_8_66_476_0 & ~i_8_66_1637_0 & ~i_8_66_1984_0 & i_8_66_1997_0 & ~i_8_66_2077_0) | (~i_8_66_193_0 & i_8_66_462_0 & ~i_8_66_787_0 & ~i_8_66_1854_0 & ~i_8_66_2214_0 & ~i_8_66_2259_0))) | (~i_8_66_774_0 & ~i_8_66_1284_0 & ~i_8_66_1654_0 & ~i_8_66_1655_0 & ~i_8_66_1854_0 & i_8_66_1997_0))) | (~i_8_66_234_0 & ((~i_8_66_2040_0 & ((~i_8_66_165_0 & ((~i_8_66_27_0 & ~i_8_66_701_0 & ~i_8_66_804_0 & ~i_8_66_1410_0 & i_8_66_1632_0 & ~i_8_66_1699_0 & ~i_8_66_2212_0) | (~i_8_66_166_0 & ~i_8_66_193_0 & ~i_8_66_241_0 & i_8_66_489_0 & ~i_8_66_616_0 & ~i_8_66_774_0 & ~i_8_66_1824_0 & ~i_8_66_1857_0 & ~i_8_66_1992_0 & ~i_8_66_2214_0))) | (i_8_66_346_0 & i_8_66_604_0 & ~i_8_66_774_0 & ~i_8_66_1625_0 & ~i_8_66_2259_0))) | (~i_8_66_238_0 & ~i_8_66_616_0 & i_8_66_747_0 & i_8_66_774_0 & ~i_8_66_1056_0 & ~i_8_66_1632_0 & ~i_8_66_1699_0 & ~i_8_66_1854_0))) | (~i_8_66_240_0 & ((i_8_66_591_0 & i_8_66_600_0 & ~i_8_66_1832_0) | (~i_8_66_384_0 & i_8_66_489_0 & ~i_8_66_720_0 & ~i_8_66_1260_0 & ~i_8_66_1279_0 & ~i_8_66_1527_0 & i_8_66_2088_0))) | (~i_8_66_27_0 & ((~i_8_66_237_0 & ((~i_8_66_1832_0 & ((~i_8_66_241_0 & ~i_8_66_337_0 & ~i_8_66_864_0 & ((i_8_66_301_0 & ~i_8_66_476_0 & ~i_8_66_774_0 & ~i_8_66_1572_0 & ~i_8_66_1611_0 & ~i_8_66_1653_0) | (~i_8_66_211_0 & i_8_66_604_0 & ~i_8_66_1528_0 & ~i_8_66_1624_0 & ~i_8_66_1947_0 & ~i_8_66_1983_0 & ~i_8_66_2077_0 & ~i_8_66_2259_0))) | (i_8_66_462_0 & i_8_66_1947_0 & ~i_8_66_2214_0))) | (i_8_66_301_0 & i_8_66_302_0 & ~i_8_66_1056_0 & ~i_8_66_1306_0 & ~i_8_66_1412_0 & ~i_8_66_1625_0 & ~i_8_66_2262_0))) | (~i_8_66_1260_0 & ((i_8_66_224_0 & ~i_8_66_462_0 & ~i_8_66_804_0 & ~i_8_66_1410_0 & i_8_66_1633_0 & ~i_8_66_1654_0) | (~i_8_66_617_0 & ~i_8_66_701_0 & ~i_8_66_720_0 & ~i_8_66_1056_0 & ~i_8_66_1527_0 & ~i_8_66_1572_0 & ~i_8_66_1634_0 & ~i_8_66_1635_0 & ~i_8_66_1854_0 & ~i_8_66_1984_0 & ~i_8_66_1992_0 & i_8_66_2154_0 & ~i_8_66_2262_0))))) | (~i_8_66_211_0 & ((i_8_66_79_0 & i_8_66_224_0 & ~i_8_66_1056_0 & ~i_8_66_1528_0 & ~i_8_66_1625_0 & ~i_8_66_1854_0) | (~i_8_66_774_0 & ~i_8_66_996_0 & ~i_8_66_1120_0 & i_8_66_1279_0 & i_8_66_1993_0 & i_8_66_1994_0))) | (i_8_66_224_0 & ((~i_8_66_476_0 & i_8_66_701_0 & ~i_8_66_1284_0 & ~i_8_66_1306_0 & ~i_8_66_1528_0 & ~i_8_66_1654_0 & ~i_8_66_1832_0) | (~i_8_66_238_0 & ~i_8_66_1625_0 & ~i_8_66_1672_0 & ~i_8_66_2077_0))) | (~i_8_66_1625_0 & ((~i_8_66_237_0 & ((~i_8_66_238_0 & ~i_8_66_774_0 & ~i_8_66_1410_0 & ~i_8_66_1637_0 & ~i_8_66_1983_0 & i_8_66_2088_0) | (~i_8_66_337_0 & ~i_8_66_1611_0 & ~i_8_66_1857_0 & ~i_8_66_2076_0 & i_8_66_2154_0))) | (~i_8_66_1306_0 & ((~i_8_66_238_0 & i_8_66_592_0 & i_8_66_710_0 & ~i_8_66_996_0) | (i_8_66_510_0 & i_8_66_1635_0 & ~i_8_66_1782_0) | (~i_8_66_337_0 & ~i_8_66_616_0 & ~i_8_66_1279_0 & ~i_8_66_1284_0 & ~i_8_66_1857_0 & i_8_66_1994_0) | (~i_8_66_1624_0 & i_8_66_1637_0 & i_8_66_1997_0 & ~i_8_66_2076_0))) | (i_8_66_593_0 & ~i_8_66_617_0 & ~i_8_66_1832_0 & ~i_8_66_2154_0 & ~i_8_66_2259_0 & ~i_8_66_1854_0 & ~i_8_66_1984_0))) | (~i_8_66_238_0 & ((~i_8_66_616_0 & ~i_8_66_710_0 & ~i_8_66_864_0 & ~i_8_66_1260_0 & ~i_8_66_1279_0 & ~i_8_66_1284_0 & ~i_8_66_1306_0 & ~i_8_66_1410_0 & i_8_66_1438_0 & ~i_8_66_1672_0 & ~i_8_66_1832_0) | (~i_8_66_166_0 & i_8_66_592_0 & i_8_66_593_0 & ~i_8_66_1854_0 & i_8_66_1997_0))) | (~i_8_66_616_0 & ((i_8_66_462_0 & ((i_8_66_1047_0 & ~i_8_66_1611_0 & i_8_66_1782_0 & ~i_8_66_1992_0 & ~i_8_66_1994_0) | (~i_8_66_525_0 & ~i_8_66_617_0 & ~i_8_66_747_0 & ~i_8_66_804_0 & i_8_66_1279_0 & i_8_66_1983_0 & ~i_8_66_2259_0))) | (~i_8_66_864_0 & ~i_8_66_1284_0 & ~i_8_66_462_0 & ~i_8_66_489_0 & ~i_8_66_1653_0 & ~i_8_66_1857_0 & ~i_8_66_1983_0 & ~i_8_66_1984_0 & i_8_66_2214_0))) | (~i_8_66_604_0 & i_8_66_1997_0 & ((~i_8_66_241_0 & ~i_8_66_346_0 & i_8_66_850_0 & ~i_8_66_1260_0 & ~i_8_66_1624_0) | (~i_8_66_193_0 & ~i_8_66_476_0 & ~i_8_66_602_0 & ~i_8_66_658_0 & ~i_8_66_1284_0 & ~i_8_66_1306_0 & i_8_66_1624_0 & ~i_8_66_1653_0))) | (~i_8_66_617_0 & ~i_8_66_1624_0 & ((~i_8_66_337_0 & i_8_66_701_0 & ~i_8_66_1412_0 & ~i_8_66_1438_0 & i_8_66_1625_0) | (~i_8_66_804_0 & ~i_8_66_1527_0 & ~i_8_66_1611_0 & ~i_8_66_1634_0 & ~i_8_66_1854_0 & i_8_66_1992_0 & i_8_66_1993_0 & ~i_8_66_2040_0 & ~i_8_66_2262_0))) | (~i_8_66_720_0 & ~i_8_66_2077_0 & ((~i_8_66_804_0 & i_8_66_850_0 & ~i_8_66_1983_0 & i_8_66_1992_0) | (i_8_66_600_0 & ~i_8_66_1284_0 & ~i_8_66_1410_0 & ~i_8_66_1984_0 & ~i_8_66_2259_0))) | (i_8_66_1993_0 & ((~i_8_66_658_0 & i_8_66_747_0 & ~i_8_66_1260_0 & ~i_8_66_1655_0) | (~i_8_66_1654_0 & ~i_8_66_1854_0 & i_8_66_1992_0 & i_8_66_2154_0))) | (~i_8_66_774_0 & i_8_66_1633_0 & ~i_8_66_1634_0 & ~i_8_66_1984_0 & i_8_66_1994_0));
endmodule



// Benchmark "kernel_8_67" written by ABC on Sun Jul 19 10:04:11 2020

module kernel_8_67 ( 
    i_8_67_3_0, i_8_67_26_0, i_8_67_31_0, i_8_67_64_0, i_8_67_75_0,
    i_8_67_84_0, i_8_67_111_0, i_8_67_114_0, i_8_67_138_0, i_8_67_229_0,
    i_8_67_300_0, i_8_67_301_0, i_8_67_304_0, i_8_67_318_0, i_8_67_352_0,
    i_8_67_399_0, i_8_67_416_0, i_8_67_420_0, i_8_67_437_0, i_8_67_469_0,
    i_8_67_470_0, i_8_67_553_0, i_8_67_567_0, i_8_67_570_0, i_8_67_579_0,
    i_8_67_591_0, i_8_67_598_0, i_8_67_607_0, i_8_67_624_0, i_8_67_633_0,
    i_8_67_667_0, i_8_67_676_0, i_8_67_699_0, i_8_67_705_0, i_8_67_729_0,
    i_8_67_811_0, i_8_67_832_0, i_8_67_838_0, i_8_67_839_0, i_8_67_840_0,
    i_8_67_955_0, i_8_67_956_0, i_8_67_959_0, i_8_67_1101_0, i_8_67_1107_0,
    i_8_67_1152_0, i_8_67_1225_0, i_8_67_1228_0, i_8_67_1234_0,
    i_8_67_1296_0, i_8_67_1298_0, i_8_67_1318_0, i_8_67_1326_0,
    i_8_67_1335_0, i_8_67_1344_0, i_8_67_1353_0, i_8_67_1397_0,
    i_8_67_1399_0, i_8_67_1431_0, i_8_67_1432_0, i_8_67_1434_0,
    i_8_67_1440_0, i_8_67_1483_0, i_8_67_1487_0, i_8_67_1492_0,
    i_8_67_1495_0, i_8_67_1521_0, i_8_67_1624_0, i_8_67_1635_0,
    i_8_67_1642_0, i_8_67_1647_0, i_8_67_1686_0, i_8_67_1696_0,
    i_8_67_1705_0, i_8_67_1768_0, i_8_67_1779_0, i_8_67_1786_0,
    i_8_67_1804_0, i_8_67_1806_0, i_8_67_1807_0, i_8_67_1813_0,
    i_8_67_1827_0, i_8_67_1836_0, i_8_67_1848_0, i_8_67_1911_0,
    i_8_67_1915_0, i_8_67_1917_0, i_8_67_2038_0, i_8_67_2045_0,
    i_8_67_2056_0, i_8_67_2065_0, i_8_67_2073_0, i_8_67_2074_0,
    i_8_67_2090_0, i_8_67_2119_0, i_8_67_2120_0, i_8_67_2190_0,
    i_8_67_2244_0, i_8_67_2272_0, i_8_67_2297_0,
    o_8_67_0_0  );
  input  i_8_67_3_0, i_8_67_26_0, i_8_67_31_0, i_8_67_64_0, i_8_67_75_0,
    i_8_67_84_0, i_8_67_111_0, i_8_67_114_0, i_8_67_138_0, i_8_67_229_0,
    i_8_67_300_0, i_8_67_301_0, i_8_67_304_0, i_8_67_318_0, i_8_67_352_0,
    i_8_67_399_0, i_8_67_416_0, i_8_67_420_0, i_8_67_437_0, i_8_67_469_0,
    i_8_67_470_0, i_8_67_553_0, i_8_67_567_0, i_8_67_570_0, i_8_67_579_0,
    i_8_67_591_0, i_8_67_598_0, i_8_67_607_0, i_8_67_624_0, i_8_67_633_0,
    i_8_67_667_0, i_8_67_676_0, i_8_67_699_0, i_8_67_705_0, i_8_67_729_0,
    i_8_67_811_0, i_8_67_832_0, i_8_67_838_0, i_8_67_839_0, i_8_67_840_0,
    i_8_67_955_0, i_8_67_956_0, i_8_67_959_0, i_8_67_1101_0, i_8_67_1107_0,
    i_8_67_1152_0, i_8_67_1225_0, i_8_67_1228_0, i_8_67_1234_0,
    i_8_67_1296_0, i_8_67_1298_0, i_8_67_1318_0, i_8_67_1326_0,
    i_8_67_1335_0, i_8_67_1344_0, i_8_67_1353_0, i_8_67_1397_0,
    i_8_67_1399_0, i_8_67_1431_0, i_8_67_1432_0, i_8_67_1434_0,
    i_8_67_1440_0, i_8_67_1483_0, i_8_67_1487_0, i_8_67_1492_0,
    i_8_67_1495_0, i_8_67_1521_0, i_8_67_1624_0, i_8_67_1635_0,
    i_8_67_1642_0, i_8_67_1647_0, i_8_67_1686_0, i_8_67_1696_0,
    i_8_67_1705_0, i_8_67_1768_0, i_8_67_1779_0, i_8_67_1786_0,
    i_8_67_1804_0, i_8_67_1806_0, i_8_67_1807_0, i_8_67_1813_0,
    i_8_67_1827_0, i_8_67_1836_0, i_8_67_1848_0, i_8_67_1911_0,
    i_8_67_1915_0, i_8_67_1917_0, i_8_67_2038_0, i_8_67_2045_0,
    i_8_67_2056_0, i_8_67_2065_0, i_8_67_2073_0, i_8_67_2074_0,
    i_8_67_2090_0, i_8_67_2119_0, i_8_67_2120_0, i_8_67_2190_0,
    i_8_67_2244_0, i_8_67_2272_0, i_8_67_2297_0;
  output o_8_67_0_0;
  assign o_8_67_0_0 = 0;
endmodule



// Benchmark "kernel_8_68" written by ABC on Sun Jul 19 10:04:11 2020

module kernel_8_68 ( 
    i_8_68_29_0, i_8_68_49_0, i_8_68_52_0, i_8_68_95_0, i_8_68_131_0,
    i_8_68_173_0, i_8_68_328_0, i_8_68_337_0, i_8_68_364_0, i_8_68_371_0,
    i_8_68_373_0, i_8_68_434_0, i_8_68_445_0, i_8_68_454_0, i_8_68_475_0,
    i_8_68_510_0, i_8_68_527_0, i_8_68_528_0, i_8_68_596_0, i_8_68_630_0,
    i_8_68_667_0, i_8_68_717_0, i_8_68_753_0, i_8_68_760_0, i_8_68_777_0,
    i_8_68_780_0, i_8_68_826_0, i_8_68_827_0, i_8_68_840_0, i_8_68_841_0,
    i_8_68_842_0, i_8_68_843_0, i_8_68_844_0, i_8_68_886_0, i_8_68_901_0,
    i_8_68_943_0, i_8_68_977_0, i_8_68_1031_0, i_8_68_1046_0,
    i_8_68_1103_0, i_8_68_1248_0, i_8_68_1249_0, i_8_68_1259_0,
    i_8_68_1300_0, i_8_68_1401_0, i_8_68_1427_0, i_8_68_1434_0,
    i_8_68_1435_0, i_8_68_1438_0, i_8_68_1439_0, i_8_68_1450_0,
    i_8_68_1451_0, i_8_68_1471_0, i_8_68_1533_0, i_8_68_1534_0,
    i_8_68_1535_0, i_8_68_1543_0, i_8_68_1544_0, i_8_68_1547_0,
    i_8_68_1573_0, i_8_68_1606_0, i_8_68_1626_0, i_8_68_1627_0,
    i_8_68_1628_0, i_8_68_1634_0, i_8_68_1637_0, i_8_68_1648_0,
    i_8_68_1678_0, i_8_68_1679_0, i_8_68_1681_0, i_8_68_1682_0,
    i_8_68_1701_0, i_8_68_1705_0, i_8_68_1723_0, i_8_68_1748_0,
    i_8_68_1753_0, i_8_68_1758_0, i_8_68_1759_0, i_8_68_1760_0,
    i_8_68_1761_0, i_8_68_1762_0, i_8_68_1763_0, i_8_68_1767_0,
    i_8_68_1774_0, i_8_68_1777_0, i_8_68_1857_0, i_8_68_1877_0,
    i_8_68_1929_0, i_8_68_1940_0, i_8_68_1966_0, i_8_68_1980_0,
    i_8_68_1993_0, i_8_68_2003_0, i_8_68_2109_0, i_8_68_2110_0,
    i_8_68_2119_0, i_8_68_2150_0, i_8_68_2214_0, i_8_68_2215_0,
    i_8_68_2216_0,
    o_8_68_0_0  );
  input  i_8_68_29_0, i_8_68_49_0, i_8_68_52_0, i_8_68_95_0,
    i_8_68_131_0, i_8_68_173_0, i_8_68_328_0, i_8_68_337_0, i_8_68_364_0,
    i_8_68_371_0, i_8_68_373_0, i_8_68_434_0, i_8_68_445_0, i_8_68_454_0,
    i_8_68_475_0, i_8_68_510_0, i_8_68_527_0, i_8_68_528_0, i_8_68_596_0,
    i_8_68_630_0, i_8_68_667_0, i_8_68_717_0, i_8_68_753_0, i_8_68_760_0,
    i_8_68_777_0, i_8_68_780_0, i_8_68_826_0, i_8_68_827_0, i_8_68_840_0,
    i_8_68_841_0, i_8_68_842_0, i_8_68_843_0, i_8_68_844_0, i_8_68_886_0,
    i_8_68_901_0, i_8_68_943_0, i_8_68_977_0, i_8_68_1031_0, i_8_68_1046_0,
    i_8_68_1103_0, i_8_68_1248_0, i_8_68_1249_0, i_8_68_1259_0,
    i_8_68_1300_0, i_8_68_1401_0, i_8_68_1427_0, i_8_68_1434_0,
    i_8_68_1435_0, i_8_68_1438_0, i_8_68_1439_0, i_8_68_1450_0,
    i_8_68_1451_0, i_8_68_1471_0, i_8_68_1533_0, i_8_68_1534_0,
    i_8_68_1535_0, i_8_68_1543_0, i_8_68_1544_0, i_8_68_1547_0,
    i_8_68_1573_0, i_8_68_1606_0, i_8_68_1626_0, i_8_68_1627_0,
    i_8_68_1628_0, i_8_68_1634_0, i_8_68_1637_0, i_8_68_1648_0,
    i_8_68_1678_0, i_8_68_1679_0, i_8_68_1681_0, i_8_68_1682_0,
    i_8_68_1701_0, i_8_68_1705_0, i_8_68_1723_0, i_8_68_1748_0,
    i_8_68_1753_0, i_8_68_1758_0, i_8_68_1759_0, i_8_68_1760_0,
    i_8_68_1761_0, i_8_68_1762_0, i_8_68_1763_0, i_8_68_1767_0,
    i_8_68_1774_0, i_8_68_1777_0, i_8_68_1857_0, i_8_68_1877_0,
    i_8_68_1929_0, i_8_68_1940_0, i_8_68_1966_0, i_8_68_1980_0,
    i_8_68_1993_0, i_8_68_2003_0, i_8_68_2109_0, i_8_68_2110_0,
    i_8_68_2119_0, i_8_68_2150_0, i_8_68_2214_0, i_8_68_2215_0,
    i_8_68_2216_0;
  output o_8_68_0_0;
  assign o_8_68_0_0 = 0;
endmodule



// Benchmark "kernel_8_69" written by ABC on Sun Jul 19 10:04:13 2020

module kernel_8_69 ( 
    i_8_69_3_0, i_8_69_6_0, i_8_69_7_0, i_8_69_98_0, i_8_69_115_0,
    i_8_69_203_0, i_8_69_205_0, i_8_69_206_0, i_8_69_226_0, i_8_69_227_0,
    i_8_69_228_0, i_8_69_229_0, i_8_69_230_0, i_8_69_231_0, i_8_69_232_0,
    i_8_69_233_0, i_8_69_248_0, i_8_69_325_0, i_8_69_356_0, i_8_69_357_0,
    i_8_69_383_0, i_8_69_497_0, i_8_69_499_0, i_8_69_501_0, i_8_69_502_0,
    i_8_69_571_0, i_8_69_572_0, i_8_69_574_0, i_8_69_605_0, i_8_69_606_0,
    i_8_69_609_0, i_8_69_610_0, i_8_69_611_0, i_8_69_671_0, i_8_69_672_0,
    i_8_69_714_0, i_8_69_716_0, i_8_69_717_0, i_8_69_812_0, i_8_69_822_0,
    i_8_69_838_0, i_8_69_883_0, i_8_69_884_0, i_8_69_888_0, i_8_69_889_0,
    i_8_69_890_0, i_8_69_930_0, i_8_69_932_0, i_8_69_934_0, i_8_69_958_0,
    i_8_69_966_0, i_8_69_990_0, i_8_69_1047_0, i_8_69_1049_0,
    i_8_69_1175_0, i_8_69_1236_0, i_8_69_1256_0, i_8_69_1258_0,
    i_8_69_1272_0, i_8_69_1279_0, i_8_69_1300_0, i_8_69_1336_0,
    i_8_69_1446_0, i_8_69_1491_0, i_8_69_1642_0, i_8_69_1648_0,
    i_8_69_1720_0, i_8_69_1721_0, i_8_69_1724_0, i_8_69_1747_0,
    i_8_69_1768_0, i_8_69_1769_0, i_8_69_1789_0, i_8_69_1805_0,
    i_8_69_1807_0, i_8_69_1818_0, i_8_69_1849_0, i_8_69_1850_0,
    i_8_69_1858_0, i_8_69_1865_0, i_8_69_1866_0, i_8_69_1868_0,
    i_8_69_1871_0, i_8_69_1980_0, i_8_69_1982_0, i_8_69_1983_0,
    i_8_69_1995_0, i_8_69_2074_0, i_8_69_2104_0, i_8_69_2142_0,
    i_8_69_2143_0, i_8_69_2145_0, i_8_69_2153_0, i_8_69_2176_0,
    i_8_69_2245_0, i_8_69_2246_0, i_8_69_2275_0, i_8_69_2289_0,
    i_8_69_2290_0, i_8_69_2291_0,
    o_8_69_0_0  );
  input  i_8_69_3_0, i_8_69_6_0, i_8_69_7_0, i_8_69_98_0, i_8_69_115_0,
    i_8_69_203_0, i_8_69_205_0, i_8_69_206_0, i_8_69_226_0, i_8_69_227_0,
    i_8_69_228_0, i_8_69_229_0, i_8_69_230_0, i_8_69_231_0, i_8_69_232_0,
    i_8_69_233_0, i_8_69_248_0, i_8_69_325_0, i_8_69_356_0, i_8_69_357_0,
    i_8_69_383_0, i_8_69_497_0, i_8_69_499_0, i_8_69_501_0, i_8_69_502_0,
    i_8_69_571_0, i_8_69_572_0, i_8_69_574_0, i_8_69_605_0, i_8_69_606_0,
    i_8_69_609_0, i_8_69_610_0, i_8_69_611_0, i_8_69_671_0, i_8_69_672_0,
    i_8_69_714_0, i_8_69_716_0, i_8_69_717_0, i_8_69_812_0, i_8_69_822_0,
    i_8_69_838_0, i_8_69_883_0, i_8_69_884_0, i_8_69_888_0, i_8_69_889_0,
    i_8_69_890_0, i_8_69_930_0, i_8_69_932_0, i_8_69_934_0, i_8_69_958_0,
    i_8_69_966_0, i_8_69_990_0, i_8_69_1047_0, i_8_69_1049_0,
    i_8_69_1175_0, i_8_69_1236_0, i_8_69_1256_0, i_8_69_1258_0,
    i_8_69_1272_0, i_8_69_1279_0, i_8_69_1300_0, i_8_69_1336_0,
    i_8_69_1446_0, i_8_69_1491_0, i_8_69_1642_0, i_8_69_1648_0,
    i_8_69_1720_0, i_8_69_1721_0, i_8_69_1724_0, i_8_69_1747_0,
    i_8_69_1768_0, i_8_69_1769_0, i_8_69_1789_0, i_8_69_1805_0,
    i_8_69_1807_0, i_8_69_1818_0, i_8_69_1849_0, i_8_69_1850_0,
    i_8_69_1858_0, i_8_69_1865_0, i_8_69_1866_0, i_8_69_1868_0,
    i_8_69_1871_0, i_8_69_1980_0, i_8_69_1982_0, i_8_69_1983_0,
    i_8_69_1995_0, i_8_69_2074_0, i_8_69_2104_0, i_8_69_2142_0,
    i_8_69_2143_0, i_8_69_2145_0, i_8_69_2153_0, i_8_69_2176_0,
    i_8_69_2245_0, i_8_69_2246_0, i_8_69_2275_0, i_8_69_2289_0,
    i_8_69_2290_0, i_8_69_2291_0;
  output o_8_69_0_0;
  assign o_8_69_0_0 = ~((~i_8_69_1769_0 & ((~i_8_69_205_0 & ((~i_8_69_228_0 & ~i_8_69_325_0 & ~i_8_69_609_0 & ~i_8_69_610_0 & ~i_8_69_990_0 & ~i_8_69_1272_0 & ~i_8_69_1336_0 & ~i_8_69_1648_0 & ~i_8_69_1724_0 & i_8_69_1789_0 & ~i_8_69_1980_0) | (~i_8_69_226_0 & ~i_8_69_229_0 & ~i_8_69_232_0 & ~i_8_69_233_0 & ~i_8_69_356_0 & i_8_69_671_0 & ~i_8_69_883_0 & ~i_8_69_1049_0 & ~i_8_69_1300_0 & ~i_8_69_1995_0 & ~i_8_69_2246_0))) | (~i_8_69_325_0 & ((~i_8_69_231_0 & ~i_8_69_610_0 & ~i_8_69_611_0 & ~i_8_69_990_0 & ~i_8_69_1768_0 & ((~i_8_69_233_0 & ~i_8_69_572_0 & ~i_8_69_605_0 & ~i_8_69_812_0 & ~i_8_69_888_0 & ~i_8_69_1047_0 & ~i_8_69_1279_0 & ~i_8_69_1789_0 & ~i_8_69_1980_0 & ~i_8_69_2153_0 & ~i_8_69_2176_0) | (~i_8_69_232_0 & ~i_8_69_248_0 & ~i_8_69_606_0 & ~i_8_69_609_0 & ~i_8_69_883_0 & ~i_8_69_1720_0 & ~i_8_69_1721_0 & ~i_8_69_1724_0 & ~i_8_69_1747_0 & ~i_8_69_1807_0 & ~i_8_69_1865_0 & ~i_8_69_1982_0 & ~i_8_69_2104_0 & ~i_8_69_2245_0))) | (~i_8_69_356_0 & ~i_8_69_574_0 & ~i_8_69_671_0 & ~i_8_69_884_0 & i_8_69_1279_0 & ~i_8_69_1648_0 & ~i_8_69_1724_0 & ~i_8_69_1789_0 & ~i_8_69_1858_0 & ~i_8_69_2143_0 & i_8_69_2153_0))) | (~i_8_69_574_0 & ((i_8_69_501_0 & ~i_8_69_571_0 & ~i_8_69_610_0 & ~i_8_69_890_0 & ~i_8_69_1300_0) | (~i_8_69_572_0 & ~i_8_69_609_0 & i_8_69_671_0 & ~i_8_69_1336_0 & ~i_8_69_1865_0 & ~i_8_69_1982_0 & ~i_8_69_2104_0 & ~i_8_69_2153_0))) | (~i_8_69_889_0 & ~i_8_69_890_0 & ~i_8_69_1336_0 & ~i_8_69_1446_0 & ~i_8_69_1768_0 & i_8_69_1805_0 & i_8_69_1807_0) | (~i_8_69_230_0 & ~i_8_69_497_0 & ~i_8_69_1047_0 & ~i_8_69_1721_0 & ~i_8_69_1747_0 & ~i_8_69_1805_0 & ~i_8_69_1858_0 & ~i_8_69_1866_0 & ~i_8_69_1983_0 & i_8_69_2143_0 & ~i_8_69_2153_0 & ~i_8_69_2245_0 & ~i_8_69_2290_0))) | (~i_8_69_889_0 & ((~i_8_69_230_0 & ((~i_8_69_231_0 & ~i_8_69_572_0 & i_8_69_1256_0 & ~i_8_69_1300_0 & ~i_8_69_1336_0 & ~i_8_69_1642_0 & ~i_8_69_2153_0) | (~i_8_69_115_0 & ~i_8_69_229_0 & ~i_8_69_716_0 & ~i_8_69_966_0 & ~i_8_69_1279_0 & ~i_8_69_1491_0 & ~i_8_69_1720_0 & ~i_8_69_1818_0 & ~i_8_69_1995_0 & i_8_69_2290_0))) | (~i_8_69_884_0 & ((~i_8_69_1789_0 & ((~i_8_69_115_0 & ~i_8_69_890_0 & ~i_8_69_1047_0 & ((~i_8_69_248_0 & ~i_8_69_574_0 & ~i_8_69_610_0 & ~i_8_69_611_0 & i_8_69_671_0 & ~i_8_69_1721_0) | (~i_8_69_572_0 & ~i_8_69_605_0 & ~i_8_69_1724_0 & i_8_69_1805_0 & ~i_8_69_1980_0 & ~i_8_69_2104_0))) | (~i_8_69_325_0 & ~i_8_69_2074_0 & i_8_69_2142_0 & i_8_69_2290_0))) | (~i_8_69_2153_0 & ((~i_8_69_574_0 & ~i_8_69_611_0 & i_8_69_716_0 & ~i_8_69_1279_0 & ~i_8_69_1642_0 & ~i_8_69_1724_0 & ~i_8_69_1768_0) | (~i_8_69_497_0 & i_8_69_930_0 & ~i_8_69_1747_0 & ~i_8_69_1865_0 & ~i_8_69_2104_0))))) | (~i_8_69_888_0 & ((~i_8_69_229_0 & ~i_8_69_1336_0 & ~i_8_69_2246_0 & ((~i_8_69_383_0 & ~i_8_69_497_0 & ~i_8_69_609_0 & ~i_8_69_611_0 & ~i_8_69_671_0 & ~i_8_69_883_0 & ~i_8_69_890_0 & ~i_8_69_966_0 & ~i_8_69_1175_0 & ~i_8_69_1279_0 & ~i_8_69_1300_0 & ~i_8_69_1721_0 & ~i_8_69_1724_0 & ~i_8_69_1768_0 & ~i_8_69_1871_0 & ~i_8_69_1980_0 & ~i_8_69_1982_0 & ~i_8_69_1983_0) | (i_8_69_714_0 & ~i_8_69_716_0 & ~i_8_69_958_0 & ~i_8_69_1491_0 & ~i_8_69_1747_0 & ~i_8_69_2074_0 & ~i_8_69_2104_0))) | (~i_8_69_571_0 & ~i_8_69_990_0 & ~i_8_69_2104_0 & ((~i_8_69_610_0 & ~i_8_69_883_0 & i_8_69_966_0 & ~i_8_69_1049_0 & ~i_8_69_1279_0 & ~i_8_69_1648_0 & i_8_69_2145_0) | (~i_8_69_231_0 & ~i_8_69_233_0 & i_8_69_497_0 & ~i_8_69_966_0 & i_8_69_1747_0 & ~i_8_69_1768_0 & ~i_8_69_1980_0 & ~i_8_69_1982_0 & ~i_8_69_2176_0))))) | (~i_8_69_571_0 & ~i_8_69_574_0 & ((~i_8_69_233_0 & ~i_8_69_883_0 & ~i_8_69_890_0 & ~i_8_69_990_0 & ~i_8_69_1721_0 & i_8_69_1850_0 & ~i_8_69_1983_0) | (~i_8_69_605_0 & ~i_8_69_606_0 & ~i_8_69_611_0 & ~i_8_69_717_0 & ~i_8_69_1049_0 & ~i_8_69_1336_0 & ~i_8_69_1724_0 & ~i_8_69_1818_0 & i_8_69_2275_0 & ~i_8_69_2290_0))) | (~i_8_69_572_0 & ((i_8_69_356_0 & ~i_8_69_605_0 & ~i_8_69_1818_0 & ~i_8_69_1865_0 & ~i_8_69_1980_0 & ~i_8_69_1982_0) | (~i_8_69_231_0 & ~i_8_69_611_0 & ~i_8_69_838_0 & ~i_8_69_890_0 & ~i_8_69_1049_0 & ~i_8_69_1648_0 & ~i_8_69_1747_0 & i_8_69_1805_0 & ~i_8_69_2074_0))) | (~i_8_69_606_0 & ~i_8_69_610_0 & ~i_8_69_671_0 & ~i_8_69_714_0 & ~i_8_69_838_0 & ~i_8_69_1047_0 & i_8_69_1491_0 & i_8_69_1995_0) | (i_8_69_1446_0 & ~i_8_69_1491_0 & ~i_8_69_1789_0 & ~i_8_69_1983_0 & ~i_8_69_1995_0) | (~i_8_69_232_0 & ~i_8_69_966_0 & ~i_8_69_990_0 & ~i_8_69_1805_0 & i_8_69_2104_0 & i_8_69_2145_0 & ~i_8_69_2246_0))) | (~i_8_69_1720_0 & ((~i_8_69_1768_0 & ((~i_8_69_115_0 & ~i_8_69_714_0 & ~i_8_69_2153_0 & ((~i_8_69_227_0 & ~i_8_69_233_0 & ~i_8_69_888_0 & ~i_8_69_1336_0 & i_8_69_1491_0 & ~i_8_69_1980_0) | (~i_8_69_226_0 & ~i_8_69_231_0 & ~i_8_69_232_0 & ~i_8_69_574_0 & ~i_8_69_606_0 & ~i_8_69_610_0 & ~i_8_69_611_0 & ~i_8_69_1049_0 & ~i_8_69_1648_0 & ~i_8_69_1789_0 & ~i_8_69_1818_0 & ~i_8_69_1865_0 & ~i_8_69_2143_0 & ~i_8_69_2246_0))) | (~i_8_69_230_0 & i_8_69_383_0 & ~i_8_69_609_0 & ~i_8_69_610_0 & ~i_8_69_890_0 & ~i_8_69_1983_0 & ~i_8_69_2104_0 & ~i_8_69_2246_0))) | (~i_8_69_227_0 & ((~i_8_69_572_0 & ~i_8_69_672_0 & i_8_69_958_0 & ~i_8_69_1279_0 & ~i_8_69_1642_0 & ~i_8_69_1721_0 & ~i_8_69_1805_0 & ~i_8_69_1865_0 & ~i_8_69_1980_0 & ~i_8_69_2104_0) | (~i_8_69_231_0 & ~i_8_69_606_0 & ~i_8_69_610_0 & i_8_69_838_0 & ~i_8_69_883_0 & i_8_69_1236_0 & ~i_8_69_1982_0 & i_8_69_2145_0))) | (~i_8_69_231_0 & ~i_8_69_1049_0 & ((~i_8_69_98_0 & ~i_8_69_232_0 & ~i_8_69_572_0 & ~i_8_69_605_0 & ~i_8_69_606_0 & ~i_8_69_611_0 & ~i_8_69_822_0 & ~i_8_69_883_0 & i_8_69_1648_0 & ~i_8_69_1721_0 & ~i_8_69_1866_0 & ~i_8_69_2145_0) | (~i_8_69_325_0 & i_8_69_1849_0 & ~i_8_69_1980_0 & ~i_8_69_2246_0))) | (~i_8_69_229_0 & ~i_8_69_611_0 & ~i_8_69_883_0 & ~i_8_69_884_0 & ~i_8_69_888_0 & i_8_69_1236_0 & ~i_8_69_1300_0 & ~i_8_69_1983_0 & i_8_69_2142_0) | (~i_8_69_228_0 & ~i_8_69_605_0 & ~i_8_69_990_0 & ~i_8_69_1272_0 & ~i_8_69_1721_0 & i_8_69_1849_0 & ~i_8_69_2074_0 & ~i_8_69_2289_0 & ~i_8_69_2291_0))) | (~i_8_69_609_0 & ((~i_8_69_227_0 & ~i_8_69_1300_0 & ((~i_8_69_226_0 & ~i_8_69_228_0 & ~i_8_69_231_0 & ~i_8_69_325_0 & ~i_8_69_605_0 & ~i_8_69_610_0 & ~i_8_69_611_0 & ~i_8_69_883_0 & ~i_8_69_884_0 & ~i_8_69_890_0 & ~i_8_69_990_0 & ~i_8_69_1049_0 & ~i_8_69_1236_0 & ~i_8_69_1336_0 & ~i_8_69_1818_0 & ~i_8_69_2104_0) | (~i_8_69_229_0 & ~i_8_69_1648_0 & i_8_69_1868_0 & ~i_8_69_1980_0 & ~i_8_69_2176_0))) | (~i_8_69_1049_0 & ~i_8_69_1995_0 & ((~i_8_69_966_0 & ~i_8_69_990_0 & ~i_8_69_610_0 & ~i_8_69_838_0 & i_8_69_1047_0 & ~i_8_69_1642_0 & ~i_8_69_1648_0 & ~i_8_69_1747_0) | (~i_8_69_1336_0 & ~i_8_69_1724_0 & i_8_69_115_0 & ~i_8_69_890_0 & ~i_8_69_2104_0 & ~i_8_69_2153_0 & ~i_8_69_2176_0 & ~i_8_69_2245_0 & ~i_8_69_2290_0))))) | (~i_8_69_883_0 & ((~i_8_69_966_0 & ((~i_8_69_228_0 & ~i_8_69_572_0 & ~i_8_69_932_0 & ~i_8_69_1047_0 & ~i_8_69_2104_0 & ((~i_8_69_231_0 & ~i_8_69_499_0 & ~i_8_69_822_0 & ~i_8_69_838_0 & ~i_8_69_1721_0 & ~i_8_69_1807_0 & i_8_69_1858_0 & ~i_8_69_1982_0 & ~i_8_69_2176_0 & ~i_8_69_2246_0) | (~i_8_69_233_0 & ~i_8_69_714_0 & ~i_8_69_717_0 & ~i_8_69_884_0 & ~i_8_69_888_0 & ~i_8_69_890_0 & ~i_8_69_958_0 & ~i_8_69_1049_0 & ~i_8_69_1272_0 & ~i_8_69_1279_0 & ~i_8_69_1336_0 & ~i_8_69_1446_0 & ~i_8_69_1648_0 & ~i_8_69_1805_0 & ~i_8_69_1858_0 & ~i_8_69_2142_0 & ~i_8_69_2289_0))) | (~i_8_69_838_0 & ((~i_8_69_229_0 & ~i_8_69_232_0 & ~i_8_69_574_0 & ~i_8_69_605_0 & ~i_8_69_672_0 & i_8_69_714_0 & ~i_8_69_1336_0 & ~i_8_69_1995_0 & ~i_8_69_2145_0) | (~i_8_69_714_0 & i_8_69_1336_0 & i_8_69_2289_0))))) | (~i_8_69_884_0 & ~i_8_69_1980_0 & ((~i_8_69_206_0 & i_8_69_499_0 & ~i_8_69_572_0 & ~i_8_69_610_0 & ~i_8_69_888_0 & ~i_8_69_990_0 & ~i_8_69_1724_0) | (~i_8_69_232_0 & ~i_8_69_605_0 & ~i_8_69_606_0 & ~i_8_69_611_0 & ~i_8_69_1491_0 & ~i_8_69_1789_0 & ~i_8_69_2074_0 & ~i_8_69_2104_0 & i_8_69_2142_0 & ~i_8_69_2153_0))))) | (~i_8_69_229_0 & ((~i_8_69_232_0 & ~i_8_69_325_0 & i_8_69_717_0 & i_8_69_2275_0) | (~i_8_69_226_0 & ~i_8_69_571_0 & ~i_8_69_572_0 & ~i_8_69_812_0 & ~i_8_69_888_0 & ~i_8_69_605_0 & ~i_8_69_611_0 & ~i_8_69_1256_0 & ~i_8_69_1491_0 & ~i_8_69_1724_0 & ~i_8_69_1982_0 & ~i_8_69_2074_0 & ~i_8_69_2245_0 & i_8_69_2291_0))) | (~i_8_69_605_0 & ((~i_8_69_226_0 & ~i_8_69_325_0 & ~i_8_69_884_0 & ((~i_8_69_890_0 & ~i_8_69_1047_0 & ~i_8_69_1300_0 & ~i_8_69_1805_0 & i_8_69_1982_0 & ~i_8_69_2104_0 & ~i_8_69_2176_0) | (~i_8_69_611_0 & i_8_69_958_0 & ~i_8_69_1995_0 & i_8_69_2143_0 & ~i_8_69_2246_0 & ~i_8_69_2291_0))) | (~i_8_69_838_0 & ~i_8_69_890_0 & ~i_8_69_233_0 & ~i_8_69_610_0 & ~i_8_69_1336_0 & ~i_8_69_1747_0 & ~i_8_69_1768_0 & ~i_8_69_1980_0 & i_8_69_2145_0))) | (i_8_69_502_0 & ((~i_8_69_230_0 & ~i_8_69_231_0 & ~i_8_69_233_0 & ~i_8_69_932_0 & ~i_8_69_1049_0 & ~i_8_69_1768_0 & ~i_8_69_1980_0 & ~i_8_69_1983_0) | (~i_8_69_610_0 & ~i_8_69_717_0 & ~i_8_69_990_0 & ~i_8_69_1491_0 & ~i_8_69_1648_0 & ~i_8_69_1747_0 & ~i_8_69_1789_0 & ~i_8_69_2246_0))) | (~i_8_69_990_0 & ((i_8_69_714_0 & ~i_8_69_822_0 & ~i_8_69_1049_0 & ~i_8_69_1648_0 & i_8_69_1747_0 & ~i_8_69_1789_0 & ~i_8_69_1850_0) | (i_8_69_606_0 & ~i_8_69_610_0 & ~i_8_69_671_0 & i_8_69_1047_0 & ~i_8_69_1300_0 & ~i_8_69_1642_0 & i_8_69_1983_0 & i_8_69_2142_0 & ~i_8_69_2153_0))) | (i_8_69_1789_0 & ~i_8_69_2176_0 & ((~i_8_69_1724_0 & i_8_69_1769_0 & i_8_69_1805_0 & ~i_8_69_2104_0 & ~i_8_69_2153_0 & ~i_8_69_1858_0 & ~i_8_69_1995_0) | (~i_8_69_502_0 & i_8_69_609_0 & ~i_8_69_672_0 & ~i_8_69_1047_0 & ~i_8_69_1049_0 & ~i_8_69_1336_0 & ~i_8_69_1768_0 & ~i_8_69_1980_0 & ~i_8_69_1983_0 & ~i_8_69_2245_0))) | (i_8_69_206_0 & ~i_8_69_232_0 & ~i_8_69_890_0 & ~i_8_69_2074_0 & ~i_8_69_2246_0));
endmodule



// Benchmark "kernel_8_70" written by ABC on Sun Jul 19 10:04:14 2020

module kernel_8_70 ( 
    i_8_70_21_0, i_8_70_28_0, i_8_70_31_0, i_8_70_46_0, i_8_70_101_0,
    i_8_70_119_0, i_8_70_136_0, i_8_70_230_0, i_8_70_232_0, i_8_70_298_0,
    i_8_70_302_0, i_8_70_316_0, i_8_70_326_0, i_8_70_374_0, i_8_70_388_0,
    i_8_70_423_0, i_8_70_468_0, i_8_70_489_0, i_8_70_490_0, i_8_70_521_0,
    i_8_70_551_0, i_8_70_556_0, i_8_70_608_0, i_8_70_616_0, i_8_70_622_0,
    i_8_70_623_0, i_8_70_634_0, i_8_70_637_0, i_8_70_649_0, i_8_70_677_0,
    i_8_70_684_0, i_8_70_692_0, i_8_70_702_0, i_8_70_704_0, i_8_70_830_0,
    i_8_70_839_0, i_8_70_958_0, i_8_70_974_0, i_8_70_982_0, i_8_70_983_0,
    i_8_70_992_0, i_8_70_1000_0, i_8_70_1001_0, i_8_70_1037_0,
    i_8_70_1046_0, i_8_70_1089_0, i_8_70_1216_0, i_8_70_1262_0,
    i_8_70_1271_0, i_8_70_1309_0, i_8_70_1345_0, i_8_70_1370_0,
    i_8_70_1388_0, i_8_70_1423_0, i_8_70_1424_0, i_8_70_1433_0,
    i_8_70_1460_0, i_8_70_1462_0, i_8_70_1463_0, i_8_70_1478_0,
    i_8_70_1493_0, i_8_70_1495_0, i_8_70_1514_0, i_8_70_1522_0,
    i_8_70_1536_0, i_8_70_1550_0, i_8_70_1586_0, i_8_70_1600_0,
    i_8_70_1671_0, i_8_70_1674_0, i_8_70_1678_0, i_8_70_1711_0,
    i_8_70_1714_0, i_8_70_1721_0, i_8_70_1724_0, i_8_70_1746_0,
    i_8_70_1747_0, i_8_70_1784_0, i_8_70_1805_0, i_8_70_1808_0,
    i_8_70_1821_0, i_8_70_1823_0, i_8_70_1854_0, i_8_70_1891_0,
    i_8_70_1901_0, i_8_70_2008_0, i_8_70_2038_0, i_8_70_2039_0,
    i_8_70_2054_0, i_8_70_2065_0, i_8_70_2075_0, i_8_70_2098_0,
    i_8_70_2120_0, i_8_70_2143_0, i_8_70_2149_0, i_8_70_2215_0,
    i_8_70_2225_0, i_8_70_2230_0, i_8_70_2243_0, i_8_70_2260_0,
    o_8_70_0_0  );
  input  i_8_70_21_0, i_8_70_28_0, i_8_70_31_0, i_8_70_46_0,
    i_8_70_101_0, i_8_70_119_0, i_8_70_136_0, i_8_70_230_0, i_8_70_232_0,
    i_8_70_298_0, i_8_70_302_0, i_8_70_316_0, i_8_70_326_0, i_8_70_374_0,
    i_8_70_388_0, i_8_70_423_0, i_8_70_468_0, i_8_70_489_0, i_8_70_490_0,
    i_8_70_521_0, i_8_70_551_0, i_8_70_556_0, i_8_70_608_0, i_8_70_616_0,
    i_8_70_622_0, i_8_70_623_0, i_8_70_634_0, i_8_70_637_0, i_8_70_649_0,
    i_8_70_677_0, i_8_70_684_0, i_8_70_692_0, i_8_70_702_0, i_8_70_704_0,
    i_8_70_830_0, i_8_70_839_0, i_8_70_958_0, i_8_70_974_0, i_8_70_982_0,
    i_8_70_983_0, i_8_70_992_0, i_8_70_1000_0, i_8_70_1001_0,
    i_8_70_1037_0, i_8_70_1046_0, i_8_70_1089_0, i_8_70_1216_0,
    i_8_70_1262_0, i_8_70_1271_0, i_8_70_1309_0, i_8_70_1345_0,
    i_8_70_1370_0, i_8_70_1388_0, i_8_70_1423_0, i_8_70_1424_0,
    i_8_70_1433_0, i_8_70_1460_0, i_8_70_1462_0, i_8_70_1463_0,
    i_8_70_1478_0, i_8_70_1493_0, i_8_70_1495_0, i_8_70_1514_0,
    i_8_70_1522_0, i_8_70_1536_0, i_8_70_1550_0, i_8_70_1586_0,
    i_8_70_1600_0, i_8_70_1671_0, i_8_70_1674_0, i_8_70_1678_0,
    i_8_70_1711_0, i_8_70_1714_0, i_8_70_1721_0, i_8_70_1724_0,
    i_8_70_1746_0, i_8_70_1747_0, i_8_70_1784_0, i_8_70_1805_0,
    i_8_70_1808_0, i_8_70_1821_0, i_8_70_1823_0, i_8_70_1854_0,
    i_8_70_1891_0, i_8_70_1901_0, i_8_70_2008_0, i_8_70_2038_0,
    i_8_70_2039_0, i_8_70_2054_0, i_8_70_2065_0, i_8_70_2075_0,
    i_8_70_2098_0, i_8_70_2120_0, i_8_70_2143_0, i_8_70_2149_0,
    i_8_70_2215_0, i_8_70_2225_0, i_8_70_2230_0, i_8_70_2243_0,
    i_8_70_2260_0;
  output o_8_70_0_0;
  assign o_8_70_0_0 = 0;
endmodule



// Benchmark "kernel_8_71" written by ABC on Sun Jul 19 10:04:15 2020

module kernel_8_71 ( 
    i_8_71_22_0, i_8_71_29_0, i_8_71_80_0, i_8_71_112_0, i_8_71_139_0,
    i_8_71_148_0, i_8_71_221_0, i_8_71_224_0, i_8_71_256_0, i_8_71_296_0,
    i_8_71_304_0, i_8_71_305_0, i_8_71_329_0, i_8_71_377_0, i_8_71_414_0,
    i_8_71_457_0, i_8_71_485_0, i_8_71_486_0, i_8_71_549_0, i_8_71_550_0,
    i_8_71_551_0, i_8_71_554_0, i_8_71_578_0, i_8_71_585_0, i_8_71_586_0,
    i_8_71_587_0, i_8_71_590_0, i_8_71_596_0, i_8_71_605_0, i_8_71_612_0,
    i_8_71_638_0, i_8_71_662_0, i_8_71_675_0, i_8_71_676_0, i_8_71_677_0,
    i_8_71_699_0, i_8_71_716_0, i_8_71_719_0, i_8_71_784_0, i_8_71_790_0,
    i_8_71_821_0, i_8_71_822_0, i_8_71_838_0, i_8_71_839_0, i_8_71_851_0,
    i_8_71_864_0, i_8_71_865_0, i_8_71_946_0, i_8_71_983_0, i_8_71_1045_0,
    i_8_71_1046_0, i_8_71_1100_0, i_8_71_1130_0, i_8_71_1201_0,
    i_8_71_1233_0, i_8_71_1243_0, i_8_71_1267_0, i_8_71_1305_0,
    i_8_71_1308_0, i_8_71_1316_0, i_8_71_1355_0, i_8_71_1404_0,
    i_8_71_1405_0, i_8_71_1438_0, i_8_71_1453_0, i_8_71_1458_0,
    i_8_71_1477_0, i_8_71_1478_0, i_8_71_1486_0, i_8_71_1510_0,
    i_8_71_1550_0, i_8_71_1557_0, i_8_71_1558_0, i_8_71_1559_0,
    i_8_71_1603_0, i_8_71_1620_0, i_8_71_1647_0, i_8_71_1650_0,
    i_8_71_1669_0, i_8_71_1671_0, i_8_71_1694_0, i_8_71_1712_0,
    i_8_71_1730_0, i_8_71_1746_0, i_8_71_1757_0, i_8_71_1780_0,
    i_8_71_1792_0, i_8_71_1881_0, i_8_71_1882_0, i_8_71_1883_0,
    i_8_71_1944_0, i_8_71_1946_0, i_8_71_1965_0, i_8_71_1989_0,
    i_8_71_1990_0, i_8_71_2093_0, i_8_71_2135_0, i_8_71_2144_0,
    i_8_71_2268_0, i_8_71_2296_0,
    o_8_71_0_0  );
  input  i_8_71_22_0, i_8_71_29_0, i_8_71_80_0, i_8_71_112_0,
    i_8_71_139_0, i_8_71_148_0, i_8_71_221_0, i_8_71_224_0, i_8_71_256_0,
    i_8_71_296_0, i_8_71_304_0, i_8_71_305_0, i_8_71_329_0, i_8_71_377_0,
    i_8_71_414_0, i_8_71_457_0, i_8_71_485_0, i_8_71_486_0, i_8_71_549_0,
    i_8_71_550_0, i_8_71_551_0, i_8_71_554_0, i_8_71_578_0, i_8_71_585_0,
    i_8_71_586_0, i_8_71_587_0, i_8_71_590_0, i_8_71_596_0, i_8_71_605_0,
    i_8_71_612_0, i_8_71_638_0, i_8_71_662_0, i_8_71_675_0, i_8_71_676_0,
    i_8_71_677_0, i_8_71_699_0, i_8_71_716_0, i_8_71_719_0, i_8_71_784_0,
    i_8_71_790_0, i_8_71_821_0, i_8_71_822_0, i_8_71_838_0, i_8_71_839_0,
    i_8_71_851_0, i_8_71_864_0, i_8_71_865_0, i_8_71_946_0, i_8_71_983_0,
    i_8_71_1045_0, i_8_71_1046_0, i_8_71_1100_0, i_8_71_1130_0,
    i_8_71_1201_0, i_8_71_1233_0, i_8_71_1243_0, i_8_71_1267_0,
    i_8_71_1305_0, i_8_71_1308_0, i_8_71_1316_0, i_8_71_1355_0,
    i_8_71_1404_0, i_8_71_1405_0, i_8_71_1438_0, i_8_71_1453_0,
    i_8_71_1458_0, i_8_71_1477_0, i_8_71_1478_0, i_8_71_1486_0,
    i_8_71_1510_0, i_8_71_1550_0, i_8_71_1557_0, i_8_71_1558_0,
    i_8_71_1559_0, i_8_71_1603_0, i_8_71_1620_0, i_8_71_1647_0,
    i_8_71_1650_0, i_8_71_1669_0, i_8_71_1671_0, i_8_71_1694_0,
    i_8_71_1712_0, i_8_71_1730_0, i_8_71_1746_0, i_8_71_1757_0,
    i_8_71_1780_0, i_8_71_1792_0, i_8_71_1881_0, i_8_71_1882_0,
    i_8_71_1883_0, i_8_71_1944_0, i_8_71_1946_0, i_8_71_1965_0,
    i_8_71_1989_0, i_8_71_1990_0, i_8_71_2093_0, i_8_71_2135_0,
    i_8_71_2144_0, i_8_71_2268_0, i_8_71_2296_0;
  output o_8_71_0_0;
  assign o_8_71_0_0 = 0;
endmodule



// Benchmark "kernel_8_72" written by ABC on Sun Jul 19 10:04:16 2020

module kernel_8_72 ( 
    i_8_72_19_0, i_8_72_49_0, i_8_72_52_0, i_8_72_53_0, i_8_72_66_0,
    i_8_72_74_0, i_8_72_87_0, i_8_72_103_0, i_8_72_107_0, i_8_72_223_0,
    i_8_72_243_0, i_8_72_284_0, i_8_72_288_0, i_8_72_289_0, i_8_72_325_0,
    i_8_72_367_0, i_8_72_418_0, i_8_72_427_0, i_8_72_436_0, i_8_72_491_0,
    i_8_72_523_0, i_8_72_525_0, i_8_72_526_0, i_8_72_528_0, i_8_72_530_0,
    i_8_72_598_0, i_8_72_604_0, i_8_72_608_0, i_8_72_630_0, i_8_72_631_0,
    i_8_72_643_0, i_8_72_657_0, i_8_72_683_0, i_8_72_690_0, i_8_72_693_0,
    i_8_72_694_0, i_8_72_696_0, i_8_72_698_0, i_8_72_702_0, i_8_72_703_0,
    i_8_72_706_0, i_8_72_709_0, i_8_72_710_0, i_8_72_720_0, i_8_72_721_0,
    i_8_72_723_0, i_8_72_724_0, i_8_72_725_0, i_8_72_734_0, i_8_72_763_0,
    i_8_72_778_0, i_8_72_801_0, i_8_72_805_0, i_8_72_806_0, i_8_72_829_0,
    i_8_72_838_0, i_8_72_877_0, i_8_72_967_0, i_8_72_969_0, i_8_72_970_0,
    i_8_72_976_0, i_8_72_1026_0, i_8_72_1112_0, i_8_72_1183_0,
    i_8_72_1261_0, i_8_72_1262_0, i_8_72_1264_0, i_8_72_1282_0,
    i_8_72_1299_0, i_8_72_1317_0, i_8_72_1327_0, i_8_72_1352_0,
    i_8_72_1362_0, i_8_72_1400_0, i_8_72_1407_0, i_8_72_1408_0,
    i_8_72_1435_0, i_8_72_1445_0, i_8_72_1486_0, i_8_72_1544_0,
    i_8_72_1588_0, i_8_72_1622_0, i_8_72_1750_0, i_8_72_1776_0,
    i_8_72_1777_0, i_8_72_1855_0, i_8_72_1882_0, i_8_72_1885_0,
    i_8_72_1904_0, i_8_72_1964_0, i_8_72_1984_0, i_8_72_2025_0,
    i_8_72_2028_0, i_8_72_2038_0, i_8_72_2115_0, i_8_72_2116_0,
    i_8_72_2151_0, i_8_72_2191_0, i_8_72_2228_0, i_8_72_2241_0,
    o_8_72_0_0  );
  input  i_8_72_19_0, i_8_72_49_0, i_8_72_52_0, i_8_72_53_0, i_8_72_66_0,
    i_8_72_74_0, i_8_72_87_0, i_8_72_103_0, i_8_72_107_0, i_8_72_223_0,
    i_8_72_243_0, i_8_72_284_0, i_8_72_288_0, i_8_72_289_0, i_8_72_325_0,
    i_8_72_367_0, i_8_72_418_0, i_8_72_427_0, i_8_72_436_0, i_8_72_491_0,
    i_8_72_523_0, i_8_72_525_0, i_8_72_526_0, i_8_72_528_0, i_8_72_530_0,
    i_8_72_598_0, i_8_72_604_0, i_8_72_608_0, i_8_72_630_0, i_8_72_631_0,
    i_8_72_643_0, i_8_72_657_0, i_8_72_683_0, i_8_72_690_0, i_8_72_693_0,
    i_8_72_694_0, i_8_72_696_0, i_8_72_698_0, i_8_72_702_0, i_8_72_703_0,
    i_8_72_706_0, i_8_72_709_0, i_8_72_710_0, i_8_72_720_0, i_8_72_721_0,
    i_8_72_723_0, i_8_72_724_0, i_8_72_725_0, i_8_72_734_0, i_8_72_763_0,
    i_8_72_778_0, i_8_72_801_0, i_8_72_805_0, i_8_72_806_0, i_8_72_829_0,
    i_8_72_838_0, i_8_72_877_0, i_8_72_967_0, i_8_72_969_0, i_8_72_970_0,
    i_8_72_976_0, i_8_72_1026_0, i_8_72_1112_0, i_8_72_1183_0,
    i_8_72_1261_0, i_8_72_1262_0, i_8_72_1264_0, i_8_72_1282_0,
    i_8_72_1299_0, i_8_72_1317_0, i_8_72_1327_0, i_8_72_1352_0,
    i_8_72_1362_0, i_8_72_1400_0, i_8_72_1407_0, i_8_72_1408_0,
    i_8_72_1435_0, i_8_72_1445_0, i_8_72_1486_0, i_8_72_1544_0,
    i_8_72_1588_0, i_8_72_1622_0, i_8_72_1750_0, i_8_72_1776_0,
    i_8_72_1777_0, i_8_72_1855_0, i_8_72_1882_0, i_8_72_1885_0,
    i_8_72_1904_0, i_8_72_1964_0, i_8_72_1984_0, i_8_72_2025_0,
    i_8_72_2028_0, i_8_72_2038_0, i_8_72_2115_0, i_8_72_2116_0,
    i_8_72_2151_0, i_8_72_2191_0, i_8_72_2228_0, i_8_72_2241_0;
  output o_8_72_0_0;
  assign o_8_72_0_0 = ~((~i_8_72_107_0 & ((~i_8_72_87_0 & ~i_8_72_243_0 & ~i_8_72_418_0 & ~i_8_72_720_0 & ~i_8_72_721_0 & ~i_8_72_725_0 & ~i_8_72_778_0 & ~i_8_72_1026_0 & ~i_8_72_1262_0) | (~i_8_72_52_0 & ~i_8_72_723_0 & i_8_72_1435_0 & ~i_8_72_1445_0 & ~i_8_72_2116_0 & ~i_8_72_2151_0))) | (~i_8_72_806_0 & ((~i_8_72_52_0 & ((i_8_72_427_0 & ~i_8_72_721_0) | (~i_8_72_284_0 & ~i_8_72_725_0 & ~i_8_72_801_0 & ~i_8_72_1435_0 & ~i_8_72_1588_0 & ~i_8_72_1855_0))) | (~i_8_72_694_0 & ~i_8_72_967_0 & ~i_8_72_1282_0) | (~i_8_72_53_0 & ~i_8_72_74_0 & ~i_8_72_243_0 & ~i_8_72_436_0 & ~i_8_72_631_0 & ~i_8_72_1352_0) | (~i_8_72_491_0 & ~i_8_72_1904_0 & ~i_8_72_2025_0 & ~i_8_72_2028_0 & ~i_8_72_2115_0 & ~i_8_72_2116_0))) | (~i_8_72_724_0 & ((~i_8_72_53_0 & ((i_8_72_703_0 & ~i_8_72_720_0) | (~i_8_72_657_0 & ~i_8_72_694_0 & ~i_8_72_698_0 & ~i_8_72_721_0))) | (i_8_72_53_0 & ~i_8_72_526_0 & ~i_8_72_734_0 & ~i_8_72_778_0 & ~i_8_72_829_0 & ~i_8_72_1544_0 & ~i_8_72_2025_0 & ~i_8_72_2038_0))) | (~i_8_72_725_0 & ((~i_8_72_720_0 & ((~i_8_72_838_0 & ~i_8_72_970_0 & ~i_8_72_1544_0 & ~i_8_72_2025_0) | (~i_8_72_608_0 & ~i_8_72_657_0 & ~i_8_72_709_0 & ~i_8_72_710_0 & ~i_8_72_734_0 & ~i_8_72_1445_0 & ~i_8_72_1588_0 & ~i_8_72_2116_0 & ~i_8_72_2151_0))) | (~i_8_72_103_0 & ~i_8_72_1622_0 & i_8_72_2228_0))) | (i_8_72_525_0 & ~i_8_72_696_0) | (~i_8_72_683_0 & ~i_8_72_877_0 & i_8_72_1882_0) | (i_8_72_523_0 & i_8_72_1282_0 & i_8_72_1984_0));
endmodule



// Benchmark "kernel_8_73" written by ABC on Sun Jul 19 10:04:17 2020

module kernel_8_73 ( 
    i_8_73_32_0, i_8_73_33_0, i_8_73_48_0, i_8_73_52_0, i_8_73_58_0,
    i_8_73_61_0, i_8_73_85_0, i_8_73_120_0, i_8_73_141_0, i_8_73_170_0,
    i_8_73_183_0, i_8_73_222_0, i_8_73_223_0, i_8_73_259_0, i_8_73_295_0,
    i_8_73_301_0, i_8_73_312_0, i_8_73_328_0, i_8_73_373_0, i_8_73_391_0,
    i_8_73_440_0, i_8_73_480_0, i_8_73_481_0, i_8_73_483_0, i_8_73_500_0,
    i_8_73_502_0, i_8_73_507_0, i_8_73_527_0, i_8_73_530_0, i_8_73_556_0,
    i_8_73_594_0, i_8_73_607_0, i_8_73_687_0, i_8_73_690_0, i_8_73_759_0,
    i_8_73_786_0, i_8_73_787_0, i_8_73_789_0, i_8_73_800_0, i_8_73_844_0,
    i_8_73_849_0, i_8_73_862_0, i_8_73_868_0, i_8_73_876_0, i_8_73_947_0,
    i_8_73_994_0, i_8_73_1050_0, i_8_73_1060_0, i_8_73_1075_0,
    i_8_73_1120_0, i_8_73_1218_0, i_8_73_1219_0, i_8_73_1221_0,
    i_8_73_1222_0, i_8_73_1282_0, i_8_73_1305_0, i_8_73_1306_0,
    i_8_73_1307_0, i_8_73_1308_0, i_8_73_1314_0, i_8_73_1330_0,
    i_8_73_1345_0, i_8_73_1387_0, i_8_73_1390_0, i_8_73_1410_0,
    i_8_73_1471_0, i_8_73_1506_0, i_8_73_1509_0, i_8_73_1545_0,
    i_8_73_1547_0, i_8_73_1551_0, i_8_73_1555_0, i_8_73_1560_0,
    i_8_73_1570_0, i_8_73_1654_0, i_8_73_1677_0, i_8_73_1683_0,
    i_8_73_1707_0, i_8_73_1722_0, i_8_73_1726_0, i_8_73_1738_0,
    i_8_73_1740_0, i_8_73_1749_0, i_8_73_1750_0, i_8_73_1752_0,
    i_8_73_1753_0, i_8_73_1761_0, i_8_73_1788_0, i_8_73_1791_0,
    i_8_73_1804_0, i_8_73_1879_0, i_8_73_1906_0, i_8_73_2028_0,
    i_8_73_2046_0, i_8_73_2092_0, i_8_73_2145_0, i_8_73_2172_0,
    i_8_73_2215_0, i_8_73_2216_0, i_8_73_2285_0,
    o_8_73_0_0  );
  input  i_8_73_32_0, i_8_73_33_0, i_8_73_48_0, i_8_73_52_0, i_8_73_58_0,
    i_8_73_61_0, i_8_73_85_0, i_8_73_120_0, i_8_73_141_0, i_8_73_170_0,
    i_8_73_183_0, i_8_73_222_0, i_8_73_223_0, i_8_73_259_0, i_8_73_295_0,
    i_8_73_301_0, i_8_73_312_0, i_8_73_328_0, i_8_73_373_0, i_8_73_391_0,
    i_8_73_440_0, i_8_73_480_0, i_8_73_481_0, i_8_73_483_0, i_8_73_500_0,
    i_8_73_502_0, i_8_73_507_0, i_8_73_527_0, i_8_73_530_0, i_8_73_556_0,
    i_8_73_594_0, i_8_73_607_0, i_8_73_687_0, i_8_73_690_0, i_8_73_759_0,
    i_8_73_786_0, i_8_73_787_0, i_8_73_789_0, i_8_73_800_0, i_8_73_844_0,
    i_8_73_849_0, i_8_73_862_0, i_8_73_868_0, i_8_73_876_0, i_8_73_947_0,
    i_8_73_994_0, i_8_73_1050_0, i_8_73_1060_0, i_8_73_1075_0,
    i_8_73_1120_0, i_8_73_1218_0, i_8_73_1219_0, i_8_73_1221_0,
    i_8_73_1222_0, i_8_73_1282_0, i_8_73_1305_0, i_8_73_1306_0,
    i_8_73_1307_0, i_8_73_1308_0, i_8_73_1314_0, i_8_73_1330_0,
    i_8_73_1345_0, i_8_73_1387_0, i_8_73_1390_0, i_8_73_1410_0,
    i_8_73_1471_0, i_8_73_1506_0, i_8_73_1509_0, i_8_73_1545_0,
    i_8_73_1547_0, i_8_73_1551_0, i_8_73_1555_0, i_8_73_1560_0,
    i_8_73_1570_0, i_8_73_1654_0, i_8_73_1677_0, i_8_73_1683_0,
    i_8_73_1707_0, i_8_73_1722_0, i_8_73_1726_0, i_8_73_1738_0,
    i_8_73_1740_0, i_8_73_1749_0, i_8_73_1750_0, i_8_73_1752_0,
    i_8_73_1753_0, i_8_73_1761_0, i_8_73_1788_0, i_8_73_1791_0,
    i_8_73_1804_0, i_8_73_1879_0, i_8_73_1906_0, i_8_73_2028_0,
    i_8_73_2046_0, i_8_73_2092_0, i_8_73_2145_0, i_8_73_2172_0,
    i_8_73_2215_0, i_8_73_2216_0, i_8_73_2285_0;
  output o_8_73_0_0;
  assign o_8_73_0_0 = 0;
endmodule



// Benchmark "kernel_8_74" written by ABC on Sun Jul 19 10:04:18 2020

module kernel_8_74 ( 
    i_8_74_82_0, i_8_74_136_0, i_8_74_139_0, i_8_74_157_0, i_8_74_208_0,
    i_8_74_255_0, i_8_74_289_0, i_8_74_297_0, i_8_74_339_0, i_8_74_343_0,
    i_8_74_387_0, i_8_74_388_0, i_8_74_392_0, i_8_74_445_0, i_8_74_450_0,
    i_8_74_451_0, i_8_74_460_0, i_8_74_507_0, i_8_74_508_0, i_8_74_529_0,
    i_8_74_540_0, i_8_74_549_0, i_8_74_595_0, i_8_74_598_0, i_8_74_603_0,
    i_8_74_604_0, i_8_74_610_0, i_8_74_621_0, i_8_74_669_0, i_8_74_679_0,
    i_8_74_711_0, i_8_74_712_0, i_8_74_716_0, i_8_74_735_0, i_8_74_748_0,
    i_8_74_760_0, i_8_74_765_0, i_8_74_766_0, i_8_74_770_0, i_8_74_793_0,
    i_8_74_814_0, i_8_74_828_0, i_8_74_844_0, i_8_74_877_0, i_8_74_907_0,
    i_8_74_939_0, i_8_74_946_0, i_8_74_994_0, i_8_74_1011_0, i_8_74_1012_0,
    i_8_74_1026_0, i_8_74_1071_0, i_8_74_1074_0, i_8_74_1081_0,
    i_8_74_1099_0, i_8_74_1108_0, i_8_74_1137_0, i_8_74_1251_0,
    i_8_74_1267_0, i_8_74_1323_0, i_8_74_1324_0, i_8_74_1344_0,
    i_8_74_1367_0, i_8_74_1441_0, i_8_74_1480_0, i_8_74_1503_0,
    i_8_74_1524_0, i_8_74_1548_0, i_8_74_1549_0, i_8_74_1552_0,
    i_8_74_1594_0, i_8_74_1597_0, i_8_74_1602_0, i_8_74_1605_0,
    i_8_74_1606_0, i_8_74_1611_0, i_8_74_1642_0, i_8_74_1648_0,
    i_8_74_1675_0, i_8_74_1681_0, i_8_74_1695_0, i_8_74_1701_0,
    i_8_74_1720_0, i_8_74_1730_0, i_8_74_1749_0, i_8_74_1776_0,
    i_8_74_1778_0, i_8_74_1779_0, i_8_74_1812_0, i_8_74_1819_0,
    i_8_74_1821_0, i_8_74_1890_0, i_8_74_1891_0, i_8_74_1947_0,
    i_8_74_1963_0, i_8_74_1994_0, i_8_74_2070_0, i_8_74_2140_0,
    i_8_74_2150_0, i_8_74_2214_0,
    o_8_74_0_0  );
  input  i_8_74_82_0, i_8_74_136_0, i_8_74_139_0, i_8_74_157_0,
    i_8_74_208_0, i_8_74_255_0, i_8_74_289_0, i_8_74_297_0, i_8_74_339_0,
    i_8_74_343_0, i_8_74_387_0, i_8_74_388_0, i_8_74_392_0, i_8_74_445_0,
    i_8_74_450_0, i_8_74_451_0, i_8_74_460_0, i_8_74_507_0, i_8_74_508_0,
    i_8_74_529_0, i_8_74_540_0, i_8_74_549_0, i_8_74_595_0, i_8_74_598_0,
    i_8_74_603_0, i_8_74_604_0, i_8_74_610_0, i_8_74_621_0, i_8_74_669_0,
    i_8_74_679_0, i_8_74_711_0, i_8_74_712_0, i_8_74_716_0, i_8_74_735_0,
    i_8_74_748_0, i_8_74_760_0, i_8_74_765_0, i_8_74_766_0, i_8_74_770_0,
    i_8_74_793_0, i_8_74_814_0, i_8_74_828_0, i_8_74_844_0, i_8_74_877_0,
    i_8_74_907_0, i_8_74_939_0, i_8_74_946_0, i_8_74_994_0, i_8_74_1011_0,
    i_8_74_1012_0, i_8_74_1026_0, i_8_74_1071_0, i_8_74_1074_0,
    i_8_74_1081_0, i_8_74_1099_0, i_8_74_1108_0, i_8_74_1137_0,
    i_8_74_1251_0, i_8_74_1267_0, i_8_74_1323_0, i_8_74_1324_0,
    i_8_74_1344_0, i_8_74_1367_0, i_8_74_1441_0, i_8_74_1480_0,
    i_8_74_1503_0, i_8_74_1524_0, i_8_74_1548_0, i_8_74_1549_0,
    i_8_74_1552_0, i_8_74_1594_0, i_8_74_1597_0, i_8_74_1602_0,
    i_8_74_1605_0, i_8_74_1606_0, i_8_74_1611_0, i_8_74_1642_0,
    i_8_74_1648_0, i_8_74_1675_0, i_8_74_1681_0, i_8_74_1695_0,
    i_8_74_1701_0, i_8_74_1720_0, i_8_74_1730_0, i_8_74_1749_0,
    i_8_74_1776_0, i_8_74_1778_0, i_8_74_1779_0, i_8_74_1812_0,
    i_8_74_1819_0, i_8_74_1821_0, i_8_74_1890_0, i_8_74_1891_0,
    i_8_74_1947_0, i_8_74_1963_0, i_8_74_1994_0, i_8_74_2070_0,
    i_8_74_2140_0, i_8_74_2150_0, i_8_74_2214_0;
  output o_8_74_0_0;
  assign o_8_74_0_0 = 0;
endmodule



// Benchmark "kernel_8_75" written by ABC on Sun Jul 19 10:04:19 2020

module kernel_8_75 ( 
    i_8_75_33_0, i_8_75_35_0, i_8_75_40_0, i_8_75_42_0, i_8_75_78_0,
    i_8_75_105_0, i_8_75_142_0, i_8_75_150_0, i_8_75_172_0, i_8_75_184_0,
    i_8_75_190_0, i_8_75_193_0, i_8_75_223_0, i_8_75_313_0, i_8_75_321_0,
    i_8_75_330_0, i_8_75_364_0, i_8_75_417_0, i_8_75_420_0, i_8_75_453_0,
    i_8_75_507_0, i_8_75_510_0, i_8_75_524_0, i_8_75_528_0, i_8_75_537_0,
    i_8_75_555_0, i_8_75_571_0, i_8_75_601_0, i_8_75_607_0, i_8_75_664_0,
    i_8_75_665_0, i_8_75_687_0, i_8_75_696_0, i_8_75_701_0, i_8_75_753_0,
    i_8_75_799_0, i_8_75_837_0, i_8_75_840_0, i_8_75_844_0, i_8_75_845_0,
    i_8_75_877_0, i_8_75_897_0, i_8_75_945_0, i_8_75_946_0, i_8_75_951_0,
    i_8_75_952_0, i_8_75_978_0, i_8_75_993_0, i_8_75_1014_0, i_8_75_1015_0,
    i_8_75_1120_0, i_8_75_1129_0, i_8_75_1158_0, i_8_75_1239_0,
    i_8_75_1257_0, i_8_75_1330_0, i_8_75_1339_0, i_8_75_1425_0,
    i_8_75_1464_0, i_8_75_1469_0, i_8_75_1482_0, i_8_75_1515_0,
    i_8_75_1527_0, i_8_75_1528_0, i_8_75_1536_0, i_8_75_1549_0,
    i_8_75_1555_0, i_8_75_1560_0, i_8_75_1572_0, i_8_75_1617_0,
    i_8_75_1647_0, i_8_75_1653_0, i_8_75_1662_0, i_8_75_1686_0,
    i_8_75_1689_0, i_8_75_1752_0, i_8_75_1807_0, i_8_75_1822_0,
    i_8_75_1861_0, i_8_75_1884_0, i_8_75_1887_0, i_8_75_1894_0,
    i_8_75_1914_0, i_8_75_1933_0, i_8_75_1951_0, i_8_75_1983_0,
    i_8_75_1995_0, i_8_75_1996_0, i_8_75_2050_0, i_8_75_2095_0,
    i_8_75_2104_0, i_8_75_2116_0, i_8_75_2128_0, i_8_75_2139_0,
    i_8_75_2152_0, i_8_75_2153_0, i_8_75_2183_0, i_8_75_2190_0,
    i_8_75_2226_0, i_8_75_2248_0,
    o_8_75_0_0  );
  input  i_8_75_33_0, i_8_75_35_0, i_8_75_40_0, i_8_75_42_0, i_8_75_78_0,
    i_8_75_105_0, i_8_75_142_0, i_8_75_150_0, i_8_75_172_0, i_8_75_184_0,
    i_8_75_190_0, i_8_75_193_0, i_8_75_223_0, i_8_75_313_0, i_8_75_321_0,
    i_8_75_330_0, i_8_75_364_0, i_8_75_417_0, i_8_75_420_0, i_8_75_453_0,
    i_8_75_507_0, i_8_75_510_0, i_8_75_524_0, i_8_75_528_0, i_8_75_537_0,
    i_8_75_555_0, i_8_75_571_0, i_8_75_601_0, i_8_75_607_0, i_8_75_664_0,
    i_8_75_665_0, i_8_75_687_0, i_8_75_696_0, i_8_75_701_0, i_8_75_753_0,
    i_8_75_799_0, i_8_75_837_0, i_8_75_840_0, i_8_75_844_0, i_8_75_845_0,
    i_8_75_877_0, i_8_75_897_0, i_8_75_945_0, i_8_75_946_0, i_8_75_951_0,
    i_8_75_952_0, i_8_75_978_0, i_8_75_993_0, i_8_75_1014_0, i_8_75_1015_0,
    i_8_75_1120_0, i_8_75_1129_0, i_8_75_1158_0, i_8_75_1239_0,
    i_8_75_1257_0, i_8_75_1330_0, i_8_75_1339_0, i_8_75_1425_0,
    i_8_75_1464_0, i_8_75_1469_0, i_8_75_1482_0, i_8_75_1515_0,
    i_8_75_1527_0, i_8_75_1528_0, i_8_75_1536_0, i_8_75_1549_0,
    i_8_75_1555_0, i_8_75_1560_0, i_8_75_1572_0, i_8_75_1617_0,
    i_8_75_1647_0, i_8_75_1653_0, i_8_75_1662_0, i_8_75_1686_0,
    i_8_75_1689_0, i_8_75_1752_0, i_8_75_1807_0, i_8_75_1822_0,
    i_8_75_1861_0, i_8_75_1884_0, i_8_75_1887_0, i_8_75_1894_0,
    i_8_75_1914_0, i_8_75_1933_0, i_8_75_1951_0, i_8_75_1983_0,
    i_8_75_1995_0, i_8_75_1996_0, i_8_75_2050_0, i_8_75_2095_0,
    i_8_75_2104_0, i_8_75_2116_0, i_8_75_2128_0, i_8_75_2139_0,
    i_8_75_2152_0, i_8_75_2153_0, i_8_75_2183_0, i_8_75_2190_0,
    i_8_75_2226_0, i_8_75_2248_0;
  output o_8_75_0_0;
  assign o_8_75_0_0 = 0;
endmodule



// Benchmark "kernel_8_76" written by ABC on Sun Jul 19 10:04:20 2020

module kernel_8_76 ( 
    i_8_76_1_0, i_8_76_77_0, i_8_76_115_0, i_8_76_318_0, i_8_76_319_0,
    i_8_76_362_0, i_8_76_368_0, i_8_76_398_0, i_8_76_464_0, i_8_76_505_0,
    i_8_76_526_0, i_8_76_571_0, i_8_76_575_0, i_8_76_578_0, i_8_76_580_0,
    i_8_76_581_0, i_8_76_587_0, i_8_76_589_0, i_8_76_595_0, i_8_76_607_0,
    i_8_76_610_0, i_8_76_634_0, i_8_76_636_0, i_8_76_637_0, i_8_76_692_0,
    i_8_76_707_0, i_8_76_784_0, i_8_76_840_0, i_8_76_844_0, i_8_76_883_0,
    i_8_76_892_0, i_8_76_967_0, i_8_76_995_0, i_8_76_1036_0, i_8_76_1037_0,
    i_8_76_1072_0, i_8_76_1103_0, i_8_76_1111_0, i_8_76_1127_0,
    i_8_76_1262_0, i_8_76_1264_0, i_8_76_1271_0, i_8_76_1298_0,
    i_8_76_1300_0, i_8_76_1315_0, i_8_76_1328_0, i_8_76_1334_0,
    i_8_76_1336_0, i_8_76_1337_0, i_8_76_1363_0, i_8_76_1400_0,
    i_8_76_1440_0, i_8_76_1441_0, i_8_76_1462_0, i_8_76_1471_0,
    i_8_76_1515_0, i_8_76_1524_0, i_8_76_1526_0, i_8_76_1544_0,
    i_8_76_1553_0, i_8_76_1558_0, i_8_76_1595_0, i_8_76_1603_0,
    i_8_76_1655_0, i_8_76_1684_0, i_8_76_1697_0, i_8_76_1700_0,
    i_8_76_1703_0, i_8_76_1706_0, i_8_76_1747_0, i_8_76_1748_0,
    i_8_76_1795_0, i_8_76_1819_0, i_8_76_1825_0, i_8_76_1867_0,
    i_8_76_1869_0, i_8_76_1871_0, i_8_76_1885_0, i_8_76_1888_0,
    i_8_76_1912_0, i_8_76_1913_0, i_8_76_1927_0, i_8_76_1950_0,
    i_8_76_2045_0, i_8_76_2122_0, i_8_76_2150_0, i_8_76_2154_0,
    i_8_76_2155_0, i_8_76_2157_0, i_8_76_2176_0, i_8_76_2190_0,
    i_8_76_2191_0, i_8_76_2218_0, i_8_76_2223_0, i_8_76_2224_0,
    i_8_76_2225_0, i_8_76_2243_0, i_8_76_2245_0, i_8_76_2286_0,
    i_8_76_2297_0,
    o_8_76_0_0  );
  input  i_8_76_1_0, i_8_76_77_0, i_8_76_115_0, i_8_76_318_0,
    i_8_76_319_0, i_8_76_362_0, i_8_76_368_0, i_8_76_398_0, i_8_76_464_0,
    i_8_76_505_0, i_8_76_526_0, i_8_76_571_0, i_8_76_575_0, i_8_76_578_0,
    i_8_76_580_0, i_8_76_581_0, i_8_76_587_0, i_8_76_589_0, i_8_76_595_0,
    i_8_76_607_0, i_8_76_610_0, i_8_76_634_0, i_8_76_636_0, i_8_76_637_0,
    i_8_76_692_0, i_8_76_707_0, i_8_76_784_0, i_8_76_840_0, i_8_76_844_0,
    i_8_76_883_0, i_8_76_892_0, i_8_76_967_0, i_8_76_995_0, i_8_76_1036_0,
    i_8_76_1037_0, i_8_76_1072_0, i_8_76_1103_0, i_8_76_1111_0,
    i_8_76_1127_0, i_8_76_1262_0, i_8_76_1264_0, i_8_76_1271_0,
    i_8_76_1298_0, i_8_76_1300_0, i_8_76_1315_0, i_8_76_1328_0,
    i_8_76_1334_0, i_8_76_1336_0, i_8_76_1337_0, i_8_76_1363_0,
    i_8_76_1400_0, i_8_76_1440_0, i_8_76_1441_0, i_8_76_1462_0,
    i_8_76_1471_0, i_8_76_1515_0, i_8_76_1524_0, i_8_76_1526_0,
    i_8_76_1544_0, i_8_76_1553_0, i_8_76_1558_0, i_8_76_1595_0,
    i_8_76_1603_0, i_8_76_1655_0, i_8_76_1684_0, i_8_76_1697_0,
    i_8_76_1700_0, i_8_76_1703_0, i_8_76_1706_0, i_8_76_1747_0,
    i_8_76_1748_0, i_8_76_1795_0, i_8_76_1819_0, i_8_76_1825_0,
    i_8_76_1867_0, i_8_76_1869_0, i_8_76_1871_0, i_8_76_1885_0,
    i_8_76_1888_0, i_8_76_1912_0, i_8_76_1913_0, i_8_76_1927_0,
    i_8_76_1950_0, i_8_76_2045_0, i_8_76_2122_0, i_8_76_2150_0,
    i_8_76_2154_0, i_8_76_2155_0, i_8_76_2157_0, i_8_76_2176_0,
    i_8_76_2190_0, i_8_76_2191_0, i_8_76_2218_0, i_8_76_2223_0,
    i_8_76_2224_0, i_8_76_2225_0, i_8_76_2243_0, i_8_76_2245_0,
    i_8_76_2286_0, i_8_76_2297_0;
  output o_8_76_0_0;
  assign o_8_76_0_0 = 0;
endmodule



// Benchmark "kernel_8_77" written by ABC on Sun Jul 19 10:04:20 2020

module kernel_8_77 ( 
    i_8_77_12_0, i_8_77_27_0, i_8_77_28_0, i_8_77_33_0, i_8_77_34_0,
    i_8_77_40_0, i_8_77_58_0, i_8_77_102_0, i_8_77_165_0, i_8_77_166_0,
    i_8_77_183_0, i_8_77_186_0, i_8_77_231_0, i_8_77_298_0, i_8_77_304_0,
    i_8_77_310_0, i_8_77_336_0, i_8_77_337_0, i_8_77_365_0, i_8_77_368_0,
    i_8_77_379_0, i_8_77_380_0, i_8_77_418_0, i_8_77_424_0, i_8_77_426_0,
    i_8_77_444_0, i_8_77_454_0, i_8_77_467_0, i_8_77_480_0, i_8_77_483_0,
    i_8_77_507_0, i_8_77_508_0, i_8_77_529_0, i_8_77_543_0, i_8_77_544_0,
    i_8_77_556_0, i_8_77_580_0, i_8_77_588_0, i_8_77_615_0, i_8_77_675_0,
    i_8_77_678_0, i_8_77_679_0, i_8_77_687_0, i_8_77_694_0, i_8_77_702_0,
    i_8_77_705_0, i_8_77_729_0, i_8_77_763_0, i_8_77_781_0, i_8_77_817_0,
    i_8_77_849_0, i_8_77_885_0, i_8_77_886_0, i_8_77_921_0, i_8_77_959_0,
    i_8_77_967_0, i_8_77_1054_0, i_8_77_1059_0, i_8_77_1103_0,
    i_8_77_1108_0, i_8_77_1192_0, i_8_77_1267_0, i_8_77_1284_0,
    i_8_77_1285_0, i_8_77_1290_0, i_8_77_1299_0, i_8_77_1326_0,
    i_8_77_1333_0, i_8_77_1354_0, i_8_77_1389_0, i_8_77_1395_0,
    i_8_77_1432_0, i_8_77_1468_0, i_8_77_1641_0, i_8_77_1649_0,
    i_8_77_1653_0, i_8_77_1690_0, i_8_77_1731_0, i_8_77_1740_0,
    i_8_77_1741_0, i_8_77_1769_0, i_8_77_1824_0, i_8_77_1825_0,
    i_8_77_1828_0, i_8_77_1831_0, i_8_77_1837_0, i_8_77_1884_0,
    i_8_77_1948_0, i_8_77_1983_0, i_8_77_1984_0, i_8_77_2002_0,
    i_8_77_2040_0, i_8_77_2047_0, i_8_77_2134_0, i_8_77_2146_0,
    i_8_77_2172_0, i_8_77_2214_0, i_8_77_2215_0, i_8_77_2248_0,
    i_8_77_2299_0,
    o_8_77_0_0  );
  input  i_8_77_12_0, i_8_77_27_0, i_8_77_28_0, i_8_77_33_0, i_8_77_34_0,
    i_8_77_40_0, i_8_77_58_0, i_8_77_102_0, i_8_77_165_0, i_8_77_166_0,
    i_8_77_183_0, i_8_77_186_0, i_8_77_231_0, i_8_77_298_0, i_8_77_304_0,
    i_8_77_310_0, i_8_77_336_0, i_8_77_337_0, i_8_77_365_0, i_8_77_368_0,
    i_8_77_379_0, i_8_77_380_0, i_8_77_418_0, i_8_77_424_0, i_8_77_426_0,
    i_8_77_444_0, i_8_77_454_0, i_8_77_467_0, i_8_77_480_0, i_8_77_483_0,
    i_8_77_507_0, i_8_77_508_0, i_8_77_529_0, i_8_77_543_0, i_8_77_544_0,
    i_8_77_556_0, i_8_77_580_0, i_8_77_588_0, i_8_77_615_0, i_8_77_675_0,
    i_8_77_678_0, i_8_77_679_0, i_8_77_687_0, i_8_77_694_0, i_8_77_702_0,
    i_8_77_705_0, i_8_77_729_0, i_8_77_763_0, i_8_77_781_0, i_8_77_817_0,
    i_8_77_849_0, i_8_77_885_0, i_8_77_886_0, i_8_77_921_0, i_8_77_959_0,
    i_8_77_967_0, i_8_77_1054_0, i_8_77_1059_0, i_8_77_1103_0,
    i_8_77_1108_0, i_8_77_1192_0, i_8_77_1267_0, i_8_77_1284_0,
    i_8_77_1285_0, i_8_77_1290_0, i_8_77_1299_0, i_8_77_1326_0,
    i_8_77_1333_0, i_8_77_1354_0, i_8_77_1389_0, i_8_77_1395_0,
    i_8_77_1432_0, i_8_77_1468_0, i_8_77_1641_0, i_8_77_1649_0,
    i_8_77_1653_0, i_8_77_1690_0, i_8_77_1731_0, i_8_77_1740_0,
    i_8_77_1741_0, i_8_77_1769_0, i_8_77_1824_0, i_8_77_1825_0,
    i_8_77_1828_0, i_8_77_1831_0, i_8_77_1837_0, i_8_77_1884_0,
    i_8_77_1948_0, i_8_77_1983_0, i_8_77_1984_0, i_8_77_2002_0,
    i_8_77_2040_0, i_8_77_2047_0, i_8_77_2134_0, i_8_77_2146_0,
    i_8_77_2172_0, i_8_77_2214_0, i_8_77_2215_0, i_8_77_2248_0,
    i_8_77_2299_0;
  output o_8_77_0_0;
  assign o_8_77_0_0 = 0;
endmodule



// Benchmark "kernel_8_78" written by ABC on Sun Jul 19 10:04:21 2020

module kernel_8_78 ( 
    i_8_78_1_0, i_8_78_4_0, i_8_78_74_0, i_8_78_81_0, i_8_78_82_0,
    i_8_78_243_0, i_8_78_244_0, i_8_78_249_0, i_8_78_270_0, i_8_78_370_0,
    i_8_78_371_0, i_8_78_391_0, i_8_78_421_0, i_8_78_423_0, i_8_78_504_0,
    i_8_78_505_0, i_8_78_514_0, i_8_78_550_0, i_8_78_553_0, i_8_78_568_0,
    i_8_78_575_0, i_8_78_622_0, i_8_78_636_0, i_8_78_638_0, i_8_78_649_0,
    i_8_78_658_0, i_8_78_664_0, i_8_78_704_0, i_8_78_729_0, i_8_78_730_0,
    i_8_78_799_0, i_8_78_843_0, i_8_78_844_0, i_8_78_856_0, i_8_78_895_0,
    i_8_78_896_0, i_8_78_954_0, i_8_78_970_0, i_8_78_1005_0, i_8_78_1035_0,
    i_8_78_1071_0, i_8_78_1080_0, i_8_78_1098_0, i_8_78_1108_0,
    i_8_78_1156_0, i_8_78_1239_0, i_8_78_1260_0, i_8_78_1282_0,
    i_8_78_1297_0, i_8_78_1298_0, i_8_78_1318_0, i_8_78_1353_0,
    i_8_78_1359_0, i_8_78_1363_0, i_8_78_1396_0, i_8_78_1407_0,
    i_8_78_1426_0, i_8_78_1435_0, i_8_78_1469_0, i_8_78_1474_0,
    i_8_78_1481_0, i_8_78_1489_0, i_8_78_1494_0, i_8_78_1495_0,
    i_8_78_1516_0, i_8_78_1530_0, i_8_78_1531_0, i_8_78_1543_0,
    i_8_78_1552_0, i_8_78_1553_0, i_8_78_1555_0, i_8_78_1639_0,
    i_8_78_1651_0, i_8_78_1657_0, i_8_78_1672_0, i_8_78_1707_0,
    i_8_78_1746_0, i_8_78_1749_0, i_8_78_1750_0, i_8_78_1774_0,
    i_8_78_1780_0, i_8_78_1792_0, i_8_78_1819_0, i_8_78_1823_0,
    i_8_78_1846_0, i_8_78_1873_0, i_8_78_1877_0, i_8_78_1881_0,
    i_8_78_1888_0, i_8_78_1945_0, i_8_78_1948_0, i_8_78_2035_0,
    i_8_78_2044_0, i_8_78_2062_0, i_8_78_2074_0, i_8_78_2092_0,
    i_8_78_2122_0, i_8_78_2172_0, i_8_78_2173_0, i_8_78_2296_0,
    o_8_78_0_0  );
  input  i_8_78_1_0, i_8_78_4_0, i_8_78_74_0, i_8_78_81_0, i_8_78_82_0,
    i_8_78_243_0, i_8_78_244_0, i_8_78_249_0, i_8_78_270_0, i_8_78_370_0,
    i_8_78_371_0, i_8_78_391_0, i_8_78_421_0, i_8_78_423_0, i_8_78_504_0,
    i_8_78_505_0, i_8_78_514_0, i_8_78_550_0, i_8_78_553_0, i_8_78_568_0,
    i_8_78_575_0, i_8_78_622_0, i_8_78_636_0, i_8_78_638_0, i_8_78_649_0,
    i_8_78_658_0, i_8_78_664_0, i_8_78_704_0, i_8_78_729_0, i_8_78_730_0,
    i_8_78_799_0, i_8_78_843_0, i_8_78_844_0, i_8_78_856_0, i_8_78_895_0,
    i_8_78_896_0, i_8_78_954_0, i_8_78_970_0, i_8_78_1005_0, i_8_78_1035_0,
    i_8_78_1071_0, i_8_78_1080_0, i_8_78_1098_0, i_8_78_1108_0,
    i_8_78_1156_0, i_8_78_1239_0, i_8_78_1260_0, i_8_78_1282_0,
    i_8_78_1297_0, i_8_78_1298_0, i_8_78_1318_0, i_8_78_1353_0,
    i_8_78_1359_0, i_8_78_1363_0, i_8_78_1396_0, i_8_78_1407_0,
    i_8_78_1426_0, i_8_78_1435_0, i_8_78_1469_0, i_8_78_1474_0,
    i_8_78_1481_0, i_8_78_1489_0, i_8_78_1494_0, i_8_78_1495_0,
    i_8_78_1516_0, i_8_78_1530_0, i_8_78_1531_0, i_8_78_1543_0,
    i_8_78_1552_0, i_8_78_1553_0, i_8_78_1555_0, i_8_78_1639_0,
    i_8_78_1651_0, i_8_78_1657_0, i_8_78_1672_0, i_8_78_1707_0,
    i_8_78_1746_0, i_8_78_1749_0, i_8_78_1750_0, i_8_78_1774_0,
    i_8_78_1780_0, i_8_78_1792_0, i_8_78_1819_0, i_8_78_1823_0,
    i_8_78_1846_0, i_8_78_1873_0, i_8_78_1877_0, i_8_78_1881_0,
    i_8_78_1888_0, i_8_78_1945_0, i_8_78_1948_0, i_8_78_2035_0,
    i_8_78_2044_0, i_8_78_2062_0, i_8_78_2074_0, i_8_78_2092_0,
    i_8_78_2122_0, i_8_78_2172_0, i_8_78_2173_0, i_8_78_2296_0;
  output o_8_78_0_0;
  assign o_8_78_0_0 = 0;
endmodule



// Benchmark "kernel_8_79" written by ABC on Sun Jul 19 10:04:22 2020

module kernel_8_79 ( 
    i_8_79_67_0, i_8_79_79_0, i_8_79_88_0, i_8_79_106_0, i_8_79_138_0,
    i_8_79_143_0, i_8_79_150_0, i_8_79_178_0, i_8_79_265_0, i_8_79_301_0,
    i_8_79_381_0, i_8_79_391_0, i_8_79_421_0, i_8_79_422_0, i_8_79_427_0,
    i_8_79_538_0, i_8_79_553_0, i_8_79_573_0, i_8_79_598_0, i_8_79_599_0,
    i_8_79_655_0, i_8_79_706_0, i_8_79_707_0, i_8_79_735_0, i_8_79_744_0,
    i_8_79_763_0, i_8_79_816_0, i_8_79_817_0, i_8_79_834_0, i_8_79_835_0,
    i_8_79_838_0, i_8_79_841_0, i_8_79_842_0, i_8_79_853_0, i_8_79_876_0,
    i_8_79_891_0, i_8_79_892_0, i_8_79_916_0, i_8_79_951_0, i_8_79_1087_0,
    i_8_79_1126_0, i_8_79_1127_0, i_8_79_1131_0, i_8_79_1135_0,
    i_8_79_1141_0, i_8_79_1178_0, i_8_79_1201_0, i_8_79_1267_0,
    i_8_79_1305_0, i_8_79_1306_0, i_8_79_1308_0, i_8_79_1338_0,
    i_8_79_1403_0, i_8_79_1410_0, i_8_79_1475_0, i_8_79_1481_0,
    i_8_79_1489_0, i_8_79_1492_0, i_8_79_1543_0, i_8_79_1544_0,
    i_8_79_1552_0, i_8_79_1601_0, i_8_79_1609_0, i_8_79_1645_0,
    i_8_79_1649_0, i_8_79_1651_0, i_8_79_1655_0, i_8_79_1690_0,
    i_8_79_1704_0, i_8_79_1709_0, i_8_79_1723_0, i_8_79_1750_0,
    i_8_79_1780_0, i_8_79_1814_0, i_8_79_1816_0, i_8_79_1824_0,
    i_8_79_1843_0, i_8_79_1855_0, i_8_79_1869_0, i_8_79_1885_0,
    i_8_79_1889_0, i_8_79_1912_0, i_8_79_1921_0, i_8_79_1957_0,
    i_8_79_1969_0, i_8_79_1976_0, i_8_79_1996_0, i_8_79_2023_0,
    i_8_79_2096_0, i_8_79_2119_0, i_8_79_2122_0, i_8_79_2141_0,
    i_8_79_2146_0, i_8_79_2150_0, i_8_79_2217_0, i_8_79_2218_0,
    i_8_79_2226_0, i_8_79_2227_0, i_8_79_2245_0, i_8_79_2299_0,
    o_8_79_0_0  );
  input  i_8_79_67_0, i_8_79_79_0, i_8_79_88_0, i_8_79_106_0,
    i_8_79_138_0, i_8_79_143_0, i_8_79_150_0, i_8_79_178_0, i_8_79_265_0,
    i_8_79_301_0, i_8_79_381_0, i_8_79_391_0, i_8_79_421_0, i_8_79_422_0,
    i_8_79_427_0, i_8_79_538_0, i_8_79_553_0, i_8_79_573_0, i_8_79_598_0,
    i_8_79_599_0, i_8_79_655_0, i_8_79_706_0, i_8_79_707_0, i_8_79_735_0,
    i_8_79_744_0, i_8_79_763_0, i_8_79_816_0, i_8_79_817_0, i_8_79_834_0,
    i_8_79_835_0, i_8_79_838_0, i_8_79_841_0, i_8_79_842_0, i_8_79_853_0,
    i_8_79_876_0, i_8_79_891_0, i_8_79_892_0, i_8_79_916_0, i_8_79_951_0,
    i_8_79_1087_0, i_8_79_1126_0, i_8_79_1127_0, i_8_79_1131_0,
    i_8_79_1135_0, i_8_79_1141_0, i_8_79_1178_0, i_8_79_1201_0,
    i_8_79_1267_0, i_8_79_1305_0, i_8_79_1306_0, i_8_79_1308_0,
    i_8_79_1338_0, i_8_79_1403_0, i_8_79_1410_0, i_8_79_1475_0,
    i_8_79_1481_0, i_8_79_1489_0, i_8_79_1492_0, i_8_79_1543_0,
    i_8_79_1544_0, i_8_79_1552_0, i_8_79_1601_0, i_8_79_1609_0,
    i_8_79_1645_0, i_8_79_1649_0, i_8_79_1651_0, i_8_79_1655_0,
    i_8_79_1690_0, i_8_79_1704_0, i_8_79_1709_0, i_8_79_1723_0,
    i_8_79_1750_0, i_8_79_1780_0, i_8_79_1814_0, i_8_79_1816_0,
    i_8_79_1824_0, i_8_79_1843_0, i_8_79_1855_0, i_8_79_1869_0,
    i_8_79_1885_0, i_8_79_1889_0, i_8_79_1912_0, i_8_79_1921_0,
    i_8_79_1957_0, i_8_79_1969_0, i_8_79_1976_0, i_8_79_1996_0,
    i_8_79_2023_0, i_8_79_2096_0, i_8_79_2119_0, i_8_79_2122_0,
    i_8_79_2141_0, i_8_79_2146_0, i_8_79_2150_0, i_8_79_2217_0,
    i_8_79_2218_0, i_8_79_2226_0, i_8_79_2227_0, i_8_79_2245_0,
    i_8_79_2299_0;
  output o_8_79_0_0;
  assign o_8_79_0_0 = 0;
endmodule



// Benchmark "kernel_8_80" written by ABC on Sun Jul 19 10:04:23 2020

module kernel_8_80 ( 
    i_8_80_38_0, i_8_80_41_0, i_8_80_50_0, i_8_80_57_0, i_8_80_60_0,
    i_8_80_62_0, i_8_80_95_0, i_8_80_166_0, i_8_80_239_0, i_8_80_260_0,
    i_8_80_300_0, i_8_80_319_0, i_8_80_335_0, i_8_80_338_0, i_8_80_365_0,
    i_8_80_382_0, i_8_80_421_0, i_8_80_425_0, i_8_80_427_0, i_8_80_437_0,
    i_8_80_490_0, i_8_80_493_0, i_8_80_496_0, i_8_80_497_0, i_8_80_552_0,
    i_8_80_554_0, i_8_80_555_0, i_8_80_556_0, i_8_80_584_0, i_8_80_604_0,
    i_8_80_613_0, i_8_80_653_0, i_8_80_658_0, i_8_80_676_0, i_8_80_700_0,
    i_8_80_751_0, i_8_80_755_0, i_8_80_761_0, i_8_80_799_0, i_8_80_800_0,
    i_8_80_803_0, i_8_80_932_0, i_8_80_968_0, i_8_80_1066_0, i_8_80_1073_0,
    i_8_80_1091_0, i_8_80_1156_0, i_8_80_1189_0, i_8_80_1264_0,
    i_8_80_1274_0, i_8_80_1282_0, i_8_80_1283_0, i_8_80_1285_0,
    i_8_80_1289_0, i_8_80_1292_0, i_8_80_1328_0, i_8_80_1355_0,
    i_8_80_1356_0, i_8_80_1382_0, i_8_80_1393_0, i_8_80_1409_0,
    i_8_80_1466_0, i_8_80_1472_0, i_8_80_1481_0, i_8_80_1552_0,
    i_8_80_1555_0, i_8_80_1562_0, i_8_80_1622_0, i_8_80_1625_0,
    i_8_80_1634_0, i_8_80_1651_0, i_8_80_1652_0, i_8_80_1655_0,
    i_8_80_1660_0, i_8_80_1669_0, i_8_80_1688_0, i_8_80_1706_0,
    i_8_80_1777_0, i_8_80_1781_0, i_8_80_1819_0, i_8_80_1828_0,
    i_8_80_1832_0, i_8_80_1867_0, i_8_80_1904_0, i_8_80_1939_0,
    i_8_80_1940_0, i_8_80_1943_0, i_8_80_1993_0, i_8_80_2005_0,
    i_8_80_2026_0, i_8_80_2107_0, i_8_80_2146_0, i_8_80_2153_0,
    i_8_80_2155_0, i_8_80_2156_0, i_8_80_2165_0, i_8_80_2179_0,
    i_8_80_2210_0, i_8_80_2225_0, i_8_80_2227_0,
    o_8_80_0_0  );
  input  i_8_80_38_0, i_8_80_41_0, i_8_80_50_0, i_8_80_57_0, i_8_80_60_0,
    i_8_80_62_0, i_8_80_95_0, i_8_80_166_0, i_8_80_239_0, i_8_80_260_0,
    i_8_80_300_0, i_8_80_319_0, i_8_80_335_0, i_8_80_338_0, i_8_80_365_0,
    i_8_80_382_0, i_8_80_421_0, i_8_80_425_0, i_8_80_427_0, i_8_80_437_0,
    i_8_80_490_0, i_8_80_493_0, i_8_80_496_0, i_8_80_497_0, i_8_80_552_0,
    i_8_80_554_0, i_8_80_555_0, i_8_80_556_0, i_8_80_584_0, i_8_80_604_0,
    i_8_80_613_0, i_8_80_653_0, i_8_80_658_0, i_8_80_676_0, i_8_80_700_0,
    i_8_80_751_0, i_8_80_755_0, i_8_80_761_0, i_8_80_799_0, i_8_80_800_0,
    i_8_80_803_0, i_8_80_932_0, i_8_80_968_0, i_8_80_1066_0, i_8_80_1073_0,
    i_8_80_1091_0, i_8_80_1156_0, i_8_80_1189_0, i_8_80_1264_0,
    i_8_80_1274_0, i_8_80_1282_0, i_8_80_1283_0, i_8_80_1285_0,
    i_8_80_1289_0, i_8_80_1292_0, i_8_80_1328_0, i_8_80_1355_0,
    i_8_80_1356_0, i_8_80_1382_0, i_8_80_1393_0, i_8_80_1409_0,
    i_8_80_1466_0, i_8_80_1472_0, i_8_80_1481_0, i_8_80_1552_0,
    i_8_80_1555_0, i_8_80_1562_0, i_8_80_1622_0, i_8_80_1625_0,
    i_8_80_1634_0, i_8_80_1651_0, i_8_80_1652_0, i_8_80_1655_0,
    i_8_80_1660_0, i_8_80_1669_0, i_8_80_1688_0, i_8_80_1706_0,
    i_8_80_1777_0, i_8_80_1781_0, i_8_80_1819_0, i_8_80_1828_0,
    i_8_80_1832_0, i_8_80_1867_0, i_8_80_1904_0, i_8_80_1939_0,
    i_8_80_1940_0, i_8_80_1943_0, i_8_80_1993_0, i_8_80_2005_0,
    i_8_80_2026_0, i_8_80_2107_0, i_8_80_2146_0, i_8_80_2153_0,
    i_8_80_2155_0, i_8_80_2156_0, i_8_80_2165_0, i_8_80_2179_0,
    i_8_80_2210_0, i_8_80_2225_0, i_8_80_2227_0;
  output o_8_80_0_0;
  assign o_8_80_0_0 = 0;
endmodule



// Benchmark "kernel_8_81" written by ABC on Sun Jul 19 10:04:25 2020

module kernel_8_81 ( 
    i_8_81_45_0, i_8_81_108_0, i_8_81_111_0, i_8_81_120_0, i_8_81_156_0,
    i_8_81_160_0, i_8_81_229_0, i_8_81_230_0, i_8_81_291_0, i_8_81_330_0,
    i_8_81_345_0, i_8_81_381_0, i_8_81_391_0, i_8_81_433_0, i_8_81_434_0,
    i_8_81_437_0, i_8_81_483_0, i_8_81_485_0, i_8_81_486_0, i_8_81_489_0,
    i_8_81_493_0, i_8_81_502_0, i_8_81_588_0, i_8_81_593_0, i_8_81_606_0,
    i_8_81_621_0, i_8_81_624_0, i_8_81_627_0, i_8_81_669_0, i_8_81_670_0,
    i_8_81_687_0, i_8_81_694_0, i_8_81_703_0, i_8_81_705_0, i_8_81_706_0,
    i_8_81_707_0, i_8_81_714_0, i_8_81_716_0, i_8_81_718_0, i_8_81_723_0,
    i_8_81_724_0, i_8_81_774_0, i_8_81_780_0, i_8_81_781_0, i_8_81_807_0,
    i_8_81_822_0, i_8_81_823_0, i_8_81_825_0, i_8_81_826_0, i_8_81_827_0,
    i_8_81_848_0, i_8_81_873_0, i_8_81_875_0, i_8_81_973_0, i_8_81_991_0,
    i_8_81_1015_0, i_8_81_1027_0, i_8_81_1029_0, i_8_81_1030_0,
    i_8_81_1059_0, i_8_81_1233_0, i_8_81_1254_0, i_8_81_1270_0,
    i_8_81_1288_0, i_8_81_1300_0, i_8_81_1318_0, i_8_81_1346_0,
    i_8_81_1356_0, i_8_81_1398_0, i_8_81_1399_0, i_8_81_1426_0,
    i_8_81_1437_0, i_8_81_1443_0, i_8_81_1587_0, i_8_81_1625_0,
    i_8_81_1645_0, i_8_81_1649_0, i_8_81_1652_0, i_8_81_1773_0,
    i_8_81_1803_0, i_8_81_1823_0, i_8_81_1824_0, i_8_81_1825_0,
    i_8_81_1854_0, i_8_81_1858_0, i_8_81_1864_0, i_8_81_1882_0,
    i_8_81_1884_0, i_8_81_1885_0, i_8_81_1951_0, i_8_81_1968_0,
    i_8_81_2026_0, i_8_81_2029_0, i_8_81_2073_0, i_8_81_2091_0,
    i_8_81_2122_0, i_8_81_2172_0, i_8_81_2242_0, i_8_81_2273_0,
    i_8_81_2290_0,
    o_8_81_0_0  );
  input  i_8_81_45_0, i_8_81_108_0, i_8_81_111_0, i_8_81_120_0,
    i_8_81_156_0, i_8_81_160_0, i_8_81_229_0, i_8_81_230_0, i_8_81_291_0,
    i_8_81_330_0, i_8_81_345_0, i_8_81_381_0, i_8_81_391_0, i_8_81_433_0,
    i_8_81_434_0, i_8_81_437_0, i_8_81_483_0, i_8_81_485_0, i_8_81_486_0,
    i_8_81_489_0, i_8_81_493_0, i_8_81_502_0, i_8_81_588_0, i_8_81_593_0,
    i_8_81_606_0, i_8_81_621_0, i_8_81_624_0, i_8_81_627_0, i_8_81_669_0,
    i_8_81_670_0, i_8_81_687_0, i_8_81_694_0, i_8_81_703_0, i_8_81_705_0,
    i_8_81_706_0, i_8_81_707_0, i_8_81_714_0, i_8_81_716_0, i_8_81_718_0,
    i_8_81_723_0, i_8_81_724_0, i_8_81_774_0, i_8_81_780_0, i_8_81_781_0,
    i_8_81_807_0, i_8_81_822_0, i_8_81_823_0, i_8_81_825_0, i_8_81_826_0,
    i_8_81_827_0, i_8_81_848_0, i_8_81_873_0, i_8_81_875_0, i_8_81_973_0,
    i_8_81_991_0, i_8_81_1015_0, i_8_81_1027_0, i_8_81_1029_0,
    i_8_81_1030_0, i_8_81_1059_0, i_8_81_1233_0, i_8_81_1254_0,
    i_8_81_1270_0, i_8_81_1288_0, i_8_81_1300_0, i_8_81_1318_0,
    i_8_81_1346_0, i_8_81_1356_0, i_8_81_1398_0, i_8_81_1399_0,
    i_8_81_1426_0, i_8_81_1437_0, i_8_81_1443_0, i_8_81_1587_0,
    i_8_81_1625_0, i_8_81_1645_0, i_8_81_1649_0, i_8_81_1652_0,
    i_8_81_1773_0, i_8_81_1803_0, i_8_81_1823_0, i_8_81_1824_0,
    i_8_81_1825_0, i_8_81_1854_0, i_8_81_1858_0, i_8_81_1864_0,
    i_8_81_1882_0, i_8_81_1884_0, i_8_81_1885_0, i_8_81_1951_0,
    i_8_81_1968_0, i_8_81_2026_0, i_8_81_2029_0, i_8_81_2073_0,
    i_8_81_2091_0, i_8_81_2122_0, i_8_81_2172_0, i_8_81_2242_0,
    i_8_81_2273_0, i_8_81_2290_0;
  output o_8_81_0_0;
  assign o_8_81_0_0 = ~((~i_8_81_120_0 & ((~i_8_81_433_0 & i_8_81_588_0 & ~i_8_81_669_0 & ~i_8_81_1027_0 & ~i_8_81_1346_0 & ~i_8_81_1882_0 & ~i_8_81_1951_0 & ~i_8_81_2026_0 & ~i_8_81_2242_0) | (~i_8_81_502_0 & ~i_8_81_724_0 & ~i_8_81_1587_0 & ~i_8_81_1645_0 & i_8_81_1823_0 & ~i_8_81_1858_0 & ~i_8_81_2122_0 & ~i_8_81_2290_0))) | (~i_8_81_434_0 & ((~i_8_81_502_0 & ((~i_8_81_160_0 & ((~i_8_81_483_0 & ~i_8_81_669_0 & ~i_8_81_716_0 & ~i_8_81_718_0 & ~i_8_81_807_0 & ~i_8_81_1027_0 & ~i_8_81_1029_0 & ~i_8_81_1854_0) | (~i_8_81_1426_0 & i_8_81_1645_0 & ~i_8_81_2242_0))) | (~i_8_81_621_0 & i_8_81_687_0 & ~i_8_81_822_0 & ~i_8_81_1443_0 & ~i_8_81_1587_0) | (~i_8_81_45_0 & ~i_8_81_823_0 & i_8_81_848_0 & ~i_8_81_973_0 & ~i_8_81_1858_0))) | (~i_8_81_483_0 & ((~i_8_81_156_0 & ((~i_8_81_291_0 & ~i_8_81_437_0 & ~i_8_81_827_0 & ~i_8_81_1270_0 & ~i_8_81_1587_0 & ~i_8_81_1882_0 & i_8_81_2091_0) | (~i_8_81_486_0 & ~i_8_81_624_0 & ~i_8_81_716_0 & ~i_8_81_807_0 & ~i_8_81_1015_0 & ~i_8_81_1346_0 & ~i_8_81_1437_0 & ~i_8_81_1443_0 & ~i_8_81_1625_0 & ~i_8_81_1854_0 & ~i_8_81_2122_0))) | (~i_8_81_291_0 & ~i_8_81_485_0 & ~i_8_81_489_0 & i_8_81_502_0 & ~i_8_81_1027_0))) | (~i_8_81_111_0 & ~i_8_81_156_0 & i_8_81_705_0 & ~i_8_81_822_0 & ~i_8_81_1443_0) | (~i_8_81_381_0 & i_8_81_694_0 & ~i_8_81_714_0 & ~i_8_81_827_0 & i_8_81_1649_0))) | (~i_8_81_826_0 & ((~i_8_81_45_0 & ~i_8_81_669_0 & ((i_8_81_330_0 & ~i_8_81_433_0 & ~i_8_81_485_0 & ~i_8_81_621_0 & ~i_8_81_1029_0 & ~i_8_81_1587_0 & ~i_8_81_1625_0 & ~i_8_81_1882_0 & ~i_8_81_2172_0) | (~i_8_81_502_0 & ~i_8_81_588_0 & ~i_8_81_624_0 & ~i_8_81_718_0 & ~i_8_81_781_0 & ~i_8_81_1027_0 & ~i_8_81_1346_0 & ~i_8_81_2242_0))) | (~i_8_81_716_0 & ((~i_8_81_160_0 & ~i_8_81_723_0 & ((~i_8_81_391_0 & ~i_8_81_621_0 & ~i_8_81_670_0 & ~i_8_81_694_0 & ~i_8_81_827_0 & ~i_8_81_1015_0 & ~i_8_81_1027_0 & ~i_8_81_1864_0 & ~i_8_81_2026_0) | (~i_8_81_156_0 & ~i_8_81_483_0 & ~i_8_81_486_0 & ~i_8_81_774_0 & ~i_8_81_875_0 & ~i_8_81_991_0 & ~i_8_81_1030_0 & ~i_8_81_2122_0 & ~i_8_81_2242_0))) | (~i_8_81_391_0 & ~i_8_81_433_0 & ~i_8_81_437_0 & ~i_8_81_621_0 & ~i_8_81_714_0 & ~i_8_81_780_0 & ~i_8_81_825_0 & ~i_8_81_827_0 & ~i_8_81_1426_0 & ~i_8_81_1858_0))) | (~i_8_81_489_0 & ~i_8_81_502_0 & ~i_8_81_723_0 & ~i_8_81_774_0 & ~i_8_81_807_0 & ~i_8_81_823_0 & ~i_8_81_827_0 & ~i_8_81_973_0 & ~i_8_81_1027_0 & ~i_8_81_1030_0 & ~i_8_81_1858_0 & ~i_8_81_2122_0 & ~i_8_81_2273_0))) | (~i_8_81_156_0 & ((~i_8_81_391_0 & ~i_8_81_437_0 & i_8_81_493_0 & ~i_8_81_807_0 & ~i_8_81_1015_0 & ~i_8_81_1254_0 & ~i_8_81_1346_0 & ~i_8_81_1426_0 & ~i_8_81_1587_0) | (i_8_81_483_0 & ~i_8_81_489_0 & ~i_8_81_502_0 & ~i_8_81_716_0 & ~i_8_81_1029_0 & ~i_8_81_1233_0 & ~i_8_81_1649_0 & ~i_8_81_2029_0))) | (~i_8_81_1027_0 & ((~i_8_81_345_0 & ~i_8_81_716_0 & ((~i_8_81_624_0 & ~i_8_81_718_0 & ~i_8_81_807_0 & ~i_8_81_848_0 & i_8_81_1346_0) | (i_8_81_588_0 & ~i_8_81_714_0 & ~i_8_81_780_0 & ~i_8_81_823_0 & ~i_8_81_2026_0))) | (~i_8_81_437_0 & ~i_8_81_1029_0 & ~i_8_81_2273_0 & ((~i_8_81_160_0 & ~i_8_81_483_0 & ~i_8_81_670_0 & ~i_8_81_694_0 & ~i_8_81_718_0 & ~i_8_81_827_0 & ~i_8_81_1854_0) | (~i_8_81_485_0 & ~i_8_81_621_0 & ~i_8_81_627_0 & ~i_8_81_780_0 & ~i_8_81_825_0 & ~i_8_81_1030_0 & ~i_8_81_2026_0 & ~i_8_81_2122_0))))) | (~i_8_81_160_0 & ~i_8_81_714_0 & ((~i_8_81_493_0 & ~i_8_81_502_0 & ~i_8_81_1399_0 & i_8_81_1951_0) | (~i_8_81_108_0 & ~i_8_81_588_0 & ~i_8_81_823_0 & ~i_8_81_875_0 & ~i_8_81_991_0 & i_8_81_1030_0 & ~i_8_81_1587_0 & ~i_8_81_2273_0))) | (~i_8_81_483_0 & ((~i_8_81_621_0 & i_8_81_705_0 & ~i_8_81_1346_0) | (~i_8_81_433_0 & ~i_8_81_670_0 & ~i_8_81_875_0 & i_8_81_1773_0 & ~i_8_81_1854_0 & ~i_8_81_2026_0))) | (~i_8_81_485_0 & ~i_8_81_606_0 & ((~i_8_81_345_0 & ~i_8_81_822_0 & ~i_8_81_827_0 & i_8_81_1399_0 & ~i_8_81_1443_0) | (~i_8_81_381_0 & ~i_8_81_391_0 & ~i_8_81_502_0 & ~i_8_81_624_0 & ~i_8_81_848_0 & ~i_8_81_1300_0 & ~i_8_81_1346_0 & ~i_8_81_1437_0 & ~i_8_81_1858_0 & ~i_8_81_2026_0 & ~i_8_81_2029_0 & ~i_8_81_2273_0 & ~i_8_81_2290_0))) | (~i_8_81_627_0 & ((~i_8_81_973_0 & i_8_81_1399_0 & i_8_81_1587_0) | (i_8_81_493_0 & ~i_8_81_502_0 & ~i_8_81_1030_0 & ~i_8_81_1233_0 & ~i_8_81_1587_0 & ~i_8_81_1858_0))) | (~i_8_81_718_0 & ~i_8_81_823_0 & ~i_8_81_1346_0 & ((~i_8_81_621_0 & ~i_8_81_825_0 & ~i_8_81_848_0 & ~i_8_81_1015_0 & ~i_8_81_1029_0 & ~i_8_81_1233_0 & ~i_8_81_1356_0 & ~i_8_81_1587_0 & ~i_8_81_1649_0 & ~i_8_81_1854_0 & ~i_8_81_2122_0) | (~i_8_81_716_0 & ~i_8_81_723_0 & ~i_8_81_822_0 & i_8_81_1858_0 & ~i_8_81_1864_0 & ~i_8_81_2026_0 & ~i_8_81_2290_0))) | (i_8_81_1858_0 & ((i_8_81_1854_0 & i_8_81_1882_0 & i_8_81_2091_0) | (i_8_81_45_0 & i_8_81_345_0 & ~i_8_81_822_0 & i_8_81_2242_0))) | (~i_8_81_670_0 & i_8_81_706_0 & ~i_8_81_707_0 & ~i_8_81_973_0 & ~i_8_81_1426_0 & ~i_8_81_1587_0 & ~i_8_81_1825_0) | (i_8_81_707_0 & i_8_81_1652_0 & ~i_8_81_2026_0));
endmodule



// Benchmark "kernel_8_82" written by ABC on Sun Jul 19 10:04:26 2020

module kernel_8_82 ( 
    i_8_82_18_0, i_8_82_31_0, i_8_82_89_0, i_8_82_93_0, i_8_82_200_0,
    i_8_82_211_0, i_8_82_230_0, i_8_82_301_0, i_8_82_343_0, i_8_82_374_0,
    i_8_82_378_0, i_8_82_379_0, i_8_82_440_0, i_8_82_453_0, i_8_82_454_0,
    i_8_82_462_0, i_8_82_476_0, i_8_82_551_0, i_8_82_557_0, i_8_82_568_0,
    i_8_82_572_0, i_8_82_588_0, i_8_82_596_0, i_8_82_601_0, i_8_82_611_0,
    i_8_82_615_0, i_8_82_616_0, i_8_82_621_0, i_8_82_633_0, i_8_82_660_0,
    i_8_82_672_0, i_8_82_693_0, i_8_82_732_0, i_8_82_772_0, i_8_82_779_0,
    i_8_82_795_0, i_8_82_796_0, i_8_82_811_0, i_8_82_846_0, i_8_82_847_0,
    i_8_82_850_0, i_8_82_855_0, i_8_82_856_0, i_8_82_946_0, i_8_82_980_0,
    i_8_82_1012_0, i_8_82_1027_0, i_8_82_1065_0, i_8_82_1088_0,
    i_8_82_1125_0, i_8_82_1128_0, i_8_82_1137_0, i_8_82_1183_0,
    i_8_82_1191_0, i_8_82_1255_0, i_8_82_1256_0, i_8_82_1281_0,
    i_8_82_1307_0, i_8_82_1309_0, i_8_82_1391_0, i_8_82_1437_0,
    i_8_82_1439_0, i_8_82_1450_0, i_8_82_1488_0, i_8_82_1489_0,
    i_8_82_1525_0, i_8_82_1528_0, i_8_82_1538_0, i_8_82_1541_0,
    i_8_82_1587_0, i_8_82_1588_0, i_8_82_1614_0, i_8_82_1624_0,
    i_8_82_1630_0, i_8_82_1632_0, i_8_82_1669_0, i_8_82_1702_0,
    i_8_82_1724_0, i_8_82_1728_0, i_8_82_1741_0, i_8_82_1742_0,
    i_8_82_1795_0, i_8_82_1808_0, i_8_82_1818_0, i_8_82_1839_0,
    i_8_82_1845_0, i_8_82_1858_0, i_8_82_1870_0, i_8_82_1884_0,
    i_8_82_1903_0, i_8_82_1906_0, i_8_82_1966_0, i_8_82_1995_0,
    i_8_82_2048_0, i_8_82_2151_0, i_8_82_2188_0, i_8_82_2216_0,
    i_8_82_2217_0, i_8_82_2291_0, i_8_82_2299_0,
    o_8_82_0_0  );
  input  i_8_82_18_0, i_8_82_31_0, i_8_82_89_0, i_8_82_93_0,
    i_8_82_200_0, i_8_82_211_0, i_8_82_230_0, i_8_82_301_0, i_8_82_343_0,
    i_8_82_374_0, i_8_82_378_0, i_8_82_379_0, i_8_82_440_0, i_8_82_453_0,
    i_8_82_454_0, i_8_82_462_0, i_8_82_476_0, i_8_82_551_0, i_8_82_557_0,
    i_8_82_568_0, i_8_82_572_0, i_8_82_588_0, i_8_82_596_0, i_8_82_601_0,
    i_8_82_611_0, i_8_82_615_0, i_8_82_616_0, i_8_82_621_0, i_8_82_633_0,
    i_8_82_660_0, i_8_82_672_0, i_8_82_693_0, i_8_82_732_0, i_8_82_772_0,
    i_8_82_779_0, i_8_82_795_0, i_8_82_796_0, i_8_82_811_0, i_8_82_846_0,
    i_8_82_847_0, i_8_82_850_0, i_8_82_855_0, i_8_82_856_0, i_8_82_946_0,
    i_8_82_980_0, i_8_82_1012_0, i_8_82_1027_0, i_8_82_1065_0,
    i_8_82_1088_0, i_8_82_1125_0, i_8_82_1128_0, i_8_82_1137_0,
    i_8_82_1183_0, i_8_82_1191_0, i_8_82_1255_0, i_8_82_1256_0,
    i_8_82_1281_0, i_8_82_1307_0, i_8_82_1309_0, i_8_82_1391_0,
    i_8_82_1437_0, i_8_82_1439_0, i_8_82_1450_0, i_8_82_1488_0,
    i_8_82_1489_0, i_8_82_1525_0, i_8_82_1528_0, i_8_82_1538_0,
    i_8_82_1541_0, i_8_82_1587_0, i_8_82_1588_0, i_8_82_1614_0,
    i_8_82_1624_0, i_8_82_1630_0, i_8_82_1632_0, i_8_82_1669_0,
    i_8_82_1702_0, i_8_82_1724_0, i_8_82_1728_0, i_8_82_1741_0,
    i_8_82_1742_0, i_8_82_1795_0, i_8_82_1808_0, i_8_82_1818_0,
    i_8_82_1839_0, i_8_82_1845_0, i_8_82_1858_0, i_8_82_1870_0,
    i_8_82_1884_0, i_8_82_1903_0, i_8_82_1906_0, i_8_82_1966_0,
    i_8_82_1995_0, i_8_82_2048_0, i_8_82_2151_0, i_8_82_2188_0,
    i_8_82_2216_0, i_8_82_2217_0, i_8_82_2291_0, i_8_82_2299_0;
  output o_8_82_0_0;
  assign o_8_82_0_0 = 0;
endmodule



// Benchmark "kernel_8_83" written by ABC on Sun Jul 19 10:04:26 2020

module kernel_8_83 ( 
    i_8_83_25_0, i_8_83_26_0, i_8_83_41_0, i_8_83_44_0, i_8_83_86_0,
    i_8_83_107_0, i_8_83_176_0, i_8_83_191_0, i_8_83_214_0, i_8_83_215_0,
    i_8_83_314_0, i_8_83_331_0, i_8_83_347_0, i_8_83_377_0, i_8_83_430_0,
    i_8_83_440_0, i_8_83_457_0, i_8_83_469_0, i_8_83_470_0, i_8_83_493_0,
    i_8_83_499_0, i_8_83_500_0, i_8_83_502_0, i_8_83_611_0, i_8_83_629_0,
    i_8_83_637_0, i_8_83_661_0, i_8_83_664_0, i_8_83_665_0, i_8_83_733_0,
    i_8_83_764_0, i_8_83_772_0, i_8_83_773_0, i_8_83_799_0, i_8_83_985_0,
    i_8_83_995_0, i_8_83_1012_0, i_8_83_1015_0, i_8_83_1024_0,
    i_8_83_1033_0, i_8_83_1060_0, i_8_83_1097_0, i_8_83_1132_0,
    i_8_83_1160_0, i_8_83_1175_0, i_8_83_1187_0, i_8_83_1258_0,
    i_8_83_1268_0, i_8_83_1310_0, i_8_83_1313_0, i_8_83_1348_0,
    i_8_83_1350_0, i_8_83_1358_0, i_8_83_1411_0, i_8_83_1412_0,
    i_8_83_1592_0, i_8_83_1596_0, i_8_83_1609_0, i_8_83_1636_0,
    i_8_83_1649_0, i_8_83_1655_0, i_8_83_1675_0, i_8_83_1691_0,
    i_8_83_1736_0, i_8_83_1753_0, i_8_83_1754_0, i_8_83_1858_0,
    i_8_83_1870_0, i_8_83_1871_0, i_8_83_1889_0, i_8_83_1897_0,
    i_8_83_1907_0, i_8_83_1917_0, i_8_83_1919_0, i_8_83_1922_0,
    i_8_83_1990_0, i_8_83_1995_0, i_8_83_2002_0, i_8_83_2005_0,
    i_8_83_2006_0, i_8_83_2023_0, i_8_83_2122_0, i_8_83_2123_0,
    i_8_83_2132_0, i_8_83_2158_0, i_8_83_2159_0, i_8_83_2164_0,
    i_8_83_2174_0, i_8_83_2176_0, i_8_83_2186_0, i_8_83_2195_0,
    i_8_83_2203_0, i_8_83_2215_0, i_8_83_2216_0, i_8_83_2218_0,
    i_8_83_2263_0, i_8_83_2276_0, i_8_83_2281_0, i_8_83_2284_0,
    i_8_83_2294_0,
    o_8_83_0_0  );
  input  i_8_83_25_0, i_8_83_26_0, i_8_83_41_0, i_8_83_44_0, i_8_83_86_0,
    i_8_83_107_0, i_8_83_176_0, i_8_83_191_0, i_8_83_214_0, i_8_83_215_0,
    i_8_83_314_0, i_8_83_331_0, i_8_83_347_0, i_8_83_377_0, i_8_83_430_0,
    i_8_83_440_0, i_8_83_457_0, i_8_83_469_0, i_8_83_470_0, i_8_83_493_0,
    i_8_83_499_0, i_8_83_500_0, i_8_83_502_0, i_8_83_611_0, i_8_83_629_0,
    i_8_83_637_0, i_8_83_661_0, i_8_83_664_0, i_8_83_665_0, i_8_83_733_0,
    i_8_83_764_0, i_8_83_772_0, i_8_83_773_0, i_8_83_799_0, i_8_83_985_0,
    i_8_83_995_0, i_8_83_1012_0, i_8_83_1015_0, i_8_83_1024_0,
    i_8_83_1033_0, i_8_83_1060_0, i_8_83_1097_0, i_8_83_1132_0,
    i_8_83_1160_0, i_8_83_1175_0, i_8_83_1187_0, i_8_83_1258_0,
    i_8_83_1268_0, i_8_83_1310_0, i_8_83_1313_0, i_8_83_1348_0,
    i_8_83_1350_0, i_8_83_1358_0, i_8_83_1411_0, i_8_83_1412_0,
    i_8_83_1592_0, i_8_83_1596_0, i_8_83_1609_0, i_8_83_1636_0,
    i_8_83_1649_0, i_8_83_1655_0, i_8_83_1675_0, i_8_83_1691_0,
    i_8_83_1736_0, i_8_83_1753_0, i_8_83_1754_0, i_8_83_1858_0,
    i_8_83_1870_0, i_8_83_1871_0, i_8_83_1889_0, i_8_83_1897_0,
    i_8_83_1907_0, i_8_83_1917_0, i_8_83_1919_0, i_8_83_1922_0,
    i_8_83_1990_0, i_8_83_1995_0, i_8_83_2002_0, i_8_83_2005_0,
    i_8_83_2006_0, i_8_83_2023_0, i_8_83_2122_0, i_8_83_2123_0,
    i_8_83_2132_0, i_8_83_2158_0, i_8_83_2159_0, i_8_83_2164_0,
    i_8_83_2174_0, i_8_83_2176_0, i_8_83_2186_0, i_8_83_2195_0,
    i_8_83_2203_0, i_8_83_2215_0, i_8_83_2216_0, i_8_83_2218_0,
    i_8_83_2263_0, i_8_83_2276_0, i_8_83_2281_0, i_8_83_2284_0,
    i_8_83_2294_0;
  output o_8_83_0_0;
  assign o_8_83_0_0 = 0;
endmodule



// Benchmark "kernel_8_84" written by ABC on Sun Jul 19 10:04:27 2020

module kernel_8_84 ( 
    i_8_84_30_0, i_8_84_87_0, i_8_84_103_0, i_8_84_224_0, i_8_84_255_0,
    i_8_84_259_0, i_8_84_296_0, i_8_84_301_0, i_8_84_305_0, i_8_84_327_0,
    i_8_84_328_0, i_8_84_336_0, i_8_84_364_0, i_8_84_386_0, i_8_84_420_0,
    i_8_84_422_0, i_8_84_440_0, i_8_84_447_0, i_8_84_448_0, i_8_84_454_0,
    i_8_84_476_0, i_8_84_483_0, i_8_84_485_0, i_8_84_495_0, i_8_84_555_0,
    i_8_84_557_0, i_8_84_592_0, i_8_84_593_0, i_8_84_603_0, i_8_84_616_0,
    i_8_84_619_0, i_8_84_628_0, i_8_84_649_0, i_8_84_663_0, i_8_84_664_0,
    i_8_84_682_0, i_8_84_763_0, i_8_84_764_0, i_8_84_817_0, i_8_84_850_0,
    i_8_84_853_0, i_8_84_880_0, i_8_84_881_0, i_8_84_951_0, i_8_84_952_0,
    i_8_84_986_0, i_8_84_1032_0, i_8_84_1059_0, i_8_84_1071_0,
    i_8_84_1075_0, i_8_84_1114_0, i_8_84_1124_0, i_8_84_1307_0,
    i_8_84_1308_0, i_8_84_1311_0, i_8_84_1329_0, i_8_84_1330_0,
    i_8_84_1341_0, i_8_84_1349_0, i_8_84_1431_0, i_8_84_1432_0,
    i_8_84_1533_0, i_8_84_1537_0, i_8_84_1591_0, i_8_84_1600_0,
    i_8_84_1633_0, i_8_84_1637_0, i_8_84_1654_0, i_8_84_1671_0,
    i_8_84_1680_0, i_8_84_1723_0, i_8_84_1734_0, i_8_84_1743_0,
    i_8_84_1744_0, i_8_84_1749_0, i_8_84_1751_0, i_8_84_1786_0,
    i_8_84_1787_0, i_8_84_1790_0, i_8_84_1807_0, i_8_84_1837_0,
    i_8_84_1839_0, i_8_84_1844_0, i_8_84_1864_0, i_8_84_1867_0,
    i_8_84_1894_0, i_8_84_1951_0, i_8_84_1962_0, i_8_84_1965_0,
    i_8_84_1978_0, i_8_84_2013_0, i_8_84_2112_0, i_8_84_2131_0,
    i_8_84_2132_0, i_8_84_2146_0, i_8_84_2152_0, i_8_84_2194_0,
    i_8_84_2231_0, i_8_84_2239_0, i_8_84_2240_0,
    o_8_84_0_0  );
  input  i_8_84_30_0, i_8_84_87_0, i_8_84_103_0, i_8_84_224_0,
    i_8_84_255_0, i_8_84_259_0, i_8_84_296_0, i_8_84_301_0, i_8_84_305_0,
    i_8_84_327_0, i_8_84_328_0, i_8_84_336_0, i_8_84_364_0, i_8_84_386_0,
    i_8_84_420_0, i_8_84_422_0, i_8_84_440_0, i_8_84_447_0, i_8_84_448_0,
    i_8_84_454_0, i_8_84_476_0, i_8_84_483_0, i_8_84_485_0, i_8_84_495_0,
    i_8_84_555_0, i_8_84_557_0, i_8_84_592_0, i_8_84_593_0, i_8_84_603_0,
    i_8_84_616_0, i_8_84_619_0, i_8_84_628_0, i_8_84_649_0, i_8_84_663_0,
    i_8_84_664_0, i_8_84_682_0, i_8_84_763_0, i_8_84_764_0, i_8_84_817_0,
    i_8_84_850_0, i_8_84_853_0, i_8_84_880_0, i_8_84_881_0, i_8_84_951_0,
    i_8_84_952_0, i_8_84_986_0, i_8_84_1032_0, i_8_84_1059_0,
    i_8_84_1071_0, i_8_84_1075_0, i_8_84_1114_0, i_8_84_1124_0,
    i_8_84_1307_0, i_8_84_1308_0, i_8_84_1311_0, i_8_84_1329_0,
    i_8_84_1330_0, i_8_84_1341_0, i_8_84_1349_0, i_8_84_1431_0,
    i_8_84_1432_0, i_8_84_1533_0, i_8_84_1537_0, i_8_84_1591_0,
    i_8_84_1600_0, i_8_84_1633_0, i_8_84_1637_0, i_8_84_1654_0,
    i_8_84_1671_0, i_8_84_1680_0, i_8_84_1723_0, i_8_84_1734_0,
    i_8_84_1743_0, i_8_84_1744_0, i_8_84_1749_0, i_8_84_1751_0,
    i_8_84_1786_0, i_8_84_1787_0, i_8_84_1790_0, i_8_84_1807_0,
    i_8_84_1837_0, i_8_84_1839_0, i_8_84_1844_0, i_8_84_1864_0,
    i_8_84_1867_0, i_8_84_1894_0, i_8_84_1951_0, i_8_84_1962_0,
    i_8_84_1965_0, i_8_84_1978_0, i_8_84_2013_0, i_8_84_2112_0,
    i_8_84_2131_0, i_8_84_2132_0, i_8_84_2146_0, i_8_84_2152_0,
    i_8_84_2194_0, i_8_84_2231_0, i_8_84_2239_0, i_8_84_2240_0;
  output o_8_84_0_0;
  assign o_8_84_0_0 = 0;
endmodule



// Benchmark "kernel_8_85" written by ABC on Sun Jul 19 10:04:28 2020

module kernel_8_85 ( 
    i_8_85_14_0, i_8_85_24_0, i_8_85_26_0, i_8_85_76_0, i_8_85_78_0,
    i_8_85_86_0, i_8_85_121_0, i_8_85_140_0, i_8_85_187_0, i_8_85_189_0,
    i_8_85_196_0, i_8_85_229_0, i_8_85_238_0, i_8_85_295_0, i_8_85_303_0,
    i_8_85_327_0, i_8_85_348_0, i_8_85_383_0, i_8_85_385_0, i_8_85_386_0,
    i_8_85_401_0, i_8_85_420_0, i_8_85_447_0, i_8_85_465_0, i_8_85_525_0,
    i_8_85_528_0, i_8_85_574_0, i_8_85_609_0, i_8_85_610_0, i_8_85_611_0,
    i_8_85_638_0, i_8_85_661_0, i_8_85_798_0, i_8_85_872_0, i_8_85_877_0,
    i_8_85_956_0, i_8_85_970_0, i_8_85_1006_0, i_8_85_1034_0,
    i_8_85_1102_0, i_8_85_1120_0, i_8_85_1123_0, i_8_85_1132_0,
    i_8_85_1159_0, i_8_85_1188_0, i_8_85_1192_0, i_8_85_1194_0,
    i_8_85_1197_0, i_8_85_1221_0, i_8_85_1237_0, i_8_85_1266_0,
    i_8_85_1285_0, i_8_85_1328_0, i_8_85_1330_0, i_8_85_1398_0,
    i_8_85_1422_0, i_8_85_1455_0, i_8_85_1456_0, i_8_85_1468_0,
    i_8_85_1469_0, i_8_85_1475_0, i_8_85_1493_0, i_8_85_1504_0,
    i_8_85_1509_0, i_8_85_1510_0, i_8_85_1542_0, i_8_85_1545_0,
    i_8_85_1546_0, i_8_85_1590_0, i_8_85_1600_0, i_8_85_1617_0,
    i_8_85_1618_0, i_8_85_1639_0, i_8_85_1640_0, i_8_85_1711_0,
    i_8_85_1750_0, i_8_85_1751_0, i_8_85_1816_0, i_8_85_1842_0,
    i_8_85_1843_0, i_8_85_1876_0, i_8_85_1877_0, i_8_85_1888_0,
    i_8_85_1894_0, i_8_85_1896_0, i_8_85_1905_0, i_8_85_1949_0,
    i_8_85_1988_0, i_8_85_1995_0, i_8_85_2041_0, i_8_85_2057_0,
    i_8_85_2112_0, i_8_85_2130_0, i_8_85_2135_0, i_8_85_2149_0,
    i_8_85_2156_0, i_8_85_2185_0, i_8_85_2193_0, i_8_85_2267_0,
    i_8_85_2274_0,
    o_8_85_0_0  );
  input  i_8_85_14_0, i_8_85_24_0, i_8_85_26_0, i_8_85_76_0, i_8_85_78_0,
    i_8_85_86_0, i_8_85_121_0, i_8_85_140_0, i_8_85_187_0, i_8_85_189_0,
    i_8_85_196_0, i_8_85_229_0, i_8_85_238_0, i_8_85_295_0, i_8_85_303_0,
    i_8_85_327_0, i_8_85_348_0, i_8_85_383_0, i_8_85_385_0, i_8_85_386_0,
    i_8_85_401_0, i_8_85_420_0, i_8_85_447_0, i_8_85_465_0, i_8_85_525_0,
    i_8_85_528_0, i_8_85_574_0, i_8_85_609_0, i_8_85_610_0, i_8_85_611_0,
    i_8_85_638_0, i_8_85_661_0, i_8_85_798_0, i_8_85_872_0, i_8_85_877_0,
    i_8_85_956_0, i_8_85_970_0, i_8_85_1006_0, i_8_85_1034_0,
    i_8_85_1102_0, i_8_85_1120_0, i_8_85_1123_0, i_8_85_1132_0,
    i_8_85_1159_0, i_8_85_1188_0, i_8_85_1192_0, i_8_85_1194_0,
    i_8_85_1197_0, i_8_85_1221_0, i_8_85_1237_0, i_8_85_1266_0,
    i_8_85_1285_0, i_8_85_1328_0, i_8_85_1330_0, i_8_85_1398_0,
    i_8_85_1422_0, i_8_85_1455_0, i_8_85_1456_0, i_8_85_1468_0,
    i_8_85_1469_0, i_8_85_1475_0, i_8_85_1493_0, i_8_85_1504_0,
    i_8_85_1509_0, i_8_85_1510_0, i_8_85_1542_0, i_8_85_1545_0,
    i_8_85_1546_0, i_8_85_1590_0, i_8_85_1600_0, i_8_85_1617_0,
    i_8_85_1618_0, i_8_85_1639_0, i_8_85_1640_0, i_8_85_1711_0,
    i_8_85_1750_0, i_8_85_1751_0, i_8_85_1816_0, i_8_85_1842_0,
    i_8_85_1843_0, i_8_85_1876_0, i_8_85_1877_0, i_8_85_1888_0,
    i_8_85_1894_0, i_8_85_1896_0, i_8_85_1905_0, i_8_85_1949_0,
    i_8_85_1988_0, i_8_85_1995_0, i_8_85_2041_0, i_8_85_2057_0,
    i_8_85_2112_0, i_8_85_2130_0, i_8_85_2135_0, i_8_85_2149_0,
    i_8_85_2156_0, i_8_85_2185_0, i_8_85_2193_0, i_8_85_2267_0,
    i_8_85_2274_0;
  output o_8_85_0_0;
  assign o_8_85_0_0 = ~((~i_8_85_295_0 & ((~i_8_85_420_0 & i_8_85_528_0 & ~i_8_85_1123_0 & ~i_8_85_1455_0 & ~i_8_85_1545_0) | (~i_8_85_196_0 & ~i_8_85_447_0 & ~i_8_85_638_0 & ~i_8_85_1102_0 & ~i_8_85_1398_0 & ~i_8_85_1843_0))) | (~i_8_85_574_0 & ((~i_8_85_609_0 & ~i_8_85_798_0) | (~i_8_85_1188_0 & ~i_8_85_1192_0 & ~i_8_85_1546_0 & i_8_85_1843_0 & ~i_8_85_1905_0 & ~i_8_85_1949_0 & ~i_8_85_2193_0))) | (~i_8_85_1132_0 & ((~i_8_85_798_0 & ~i_8_85_1600_0 & ~i_8_85_1896_0) | (~i_8_85_610_0 & ~i_8_85_1188_0 & ~i_8_85_1237_0 & ~i_8_85_1590_0 & ~i_8_85_2185_0))) | (~i_8_85_24_0 & ((~i_8_85_1842_0 & ((~i_8_85_1504_0 & i_8_85_1510_0 & i_8_85_1546_0 & ~i_8_85_1905_0) | (~i_8_85_348_0 & ~i_8_85_2193_0))) | (~i_8_85_121_0 & ~i_8_85_420_0 & ~i_8_85_447_0 & ~i_8_85_528_0 & ~i_8_85_638_0))) | (~i_8_85_1888_0 & ((~i_8_85_1542_0 & i_8_85_1590_0 & ~i_8_85_1876_0 & ~i_8_85_1988_0 & ~i_8_85_2112_0) | (~i_8_85_1546_0 & ~i_8_85_1600_0 & ~i_8_85_1640_0 & ~i_8_85_2135_0 & ~i_8_85_2274_0))) | (~i_8_85_1542_0 & ((~i_8_85_76_0 & ~i_8_85_609_0 & ~i_8_85_1034_0 & ~i_8_85_1188_0) | (~i_8_85_189_0 & ~i_8_85_611_0 & ~i_8_85_956_0 & ~i_8_85_1123_0 & ~i_8_85_1456_0 & ~i_8_85_2112_0))) | i_8_85_1618_0 | (~i_8_85_26_0 & i_8_85_420_0 & ~i_8_85_661_0 & ~i_8_85_1843_0) | (i_8_85_78_0 & ~i_8_85_187_0 & ~i_8_85_1102_0 & ~i_8_85_1455_0 & ~i_8_85_1711_0 & ~i_8_85_2057_0));
endmodule



// Benchmark "kernel_8_86" written by ABC on Sun Jul 19 10:04:29 2020

module kernel_8_86 ( 
    i_8_86_7_0, i_8_86_40_0, i_8_86_64_0, i_8_86_76_0, i_8_86_79_0,
    i_8_86_139_0, i_8_86_150_0, i_8_86_151_0, i_8_86_190_0, i_8_86_214_0,
    i_8_86_230_0, i_8_86_304_0, i_8_86_322_0, i_8_86_364_0, i_8_86_376_0,
    i_8_86_394_0, i_8_86_395_0, i_8_86_400_0, i_8_86_401_0, i_8_86_420_0,
    i_8_86_421_0, i_8_86_422_0, i_8_86_446_0, i_8_86_479_0, i_8_86_482_0,
    i_8_86_483_0, i_8_86_485_0, i_8_86_490_0, i_8_86_526_0, i_8_86_530_0,
    i_8_86_570_0, i_8_86_574_0, i_8_86_592_0, i_8_86_593_0, i_8_86_594_0,
    i_8_86_596_0, i_8_86_602_0, i_8_86_611_0, i_8_86_639_0, i_8_86_642_0,
    i_8_86_705_0, i_8_86_715_0, i_8_86_728_0, i_8_86_751_0, i_8_86_762_0,
    i_8_86_814_0, i_8_86_827_0, i_8_86_843_0, i_8_86_844_0, i_8_86_845_0,
    i_8_86_859_0, i_8_86_886_0, i_8_86_895_0, i_8_86_899_0, i_8_86_925_0,
    i_8_86_1012_0, i_8_86_1027_0, i_8_86_1076_0, i_8_86_1101_0,
    i_8_86_1120_0, i_8_86_1229_0, i_8_86_1240_0, i_8_86_1271_0,
    i_8_86_1305_0, i_8_86_1308_0, i_8_86_1326_0, i_8_86_1328_0,
    i_8_86_1331_0, i_8_86_1335_0, i_8_86_1357_0, i_8_86_1416_0,
    i_8_86_1436_0, i_8_86_1437_0, i_8_86_1455_0, i_8_86_1465_0,
    i_8_86_1472_0, i_8_86_1480_0, i_8_86_1483_0, i_8_86_1547_0,
    i_8_86_1551_0, i_8_86_1573_0, i_8_86_1634_0, i_8_86_1636_0,
    i_8_86_1645_0, i_8_86_1654_0, i_8_86_1687_0, i_8_86_1707_0,
    i_8_86_1708_0, i_8_86_1723_0, i_8_86_1751_0, i_8_86_1754_0,
    i_8_86_1772_0, i_8_86_1808_0, i_8_86_1858_0, i_8_86_1912_0,
    i_8_86_1966_0, i_8_86_1996_0, i_8_86_2051_0, i_8_86_2152_0,
    i_8_86_2214_0,
    o_8_86_0_0  );
  input  i_8_86_7_0, i_8_86_40_0, i_8_86_64_0, i_8_86_76_0, i_8_86_79_0,
    i_8_86_139_0, i_8_86_150_0, i_8_86_151_0, i_8_86_190_0, i_8_86_214_0,
    i_8_86_230_0, i_8_86_304_0, i_8_86_322_0, i_8_86_364_0, i_8_86_376_0,
    i_8_86_394_0, i_8_86_395_0, i_8_86_400_0, i_8_86_401_0, i_8_86_420_0,
    i_8_86_421_0, i_8_86_422_0, i_8_86_446_0, i_8_86_479_0, i_8_86_482_0,
    i_8_86_483_0, i_8_86_485_0, i_8_86_490_0, i_8_86_526_0, i_8_86_530_0,
    i_8_86_570_0, i_8_86_574_0, i_8_86_592_0, i_8_86_593_0, i_8_86_594_0,
    i_8_86_596_0, i_8_86_602_0, i_8_86_611_0, i_8_86_639_0, i_8_86_642_0,
    i_8_86_705_0, i_8_86_715_0, i_8_86_728_0, i_8_86_751_0, i_8_86_762_0,
    i_8_86_814_0, i_8_86_827_0, i_8_86_843_0, i_8_86_844_0, i_8_86_845_0,
    i_8_86_859_0, i_8_86_886_0, i_8_86_895_0, i_8_86_899_0, i_8_86_925_0,
    i_8_86_1012_0, i_8_86_1027_0, i_8_86_1076_0, i_8_86_1101_0,
    i_8_86_1120_0, i_8_86_1229_0, i_8_86_1240_0, i_8_86_1271_0,
    i_8_86_1305_0, i_8_86_1308_0, i_8_86_1326_0, i_8_86_1328_0,
    i_8_86_1331_0, i_8_86_1335_0, i_8_86_1357_0, i_8_86_1416_0,
    i_8_86_1436_0, i_8_86_1437_0, i_8_86_1455_0, i_8_86_1465_0,
    i_8_86_1472_0, i_8_86_1480_0, i_8_86_1483_0, i_8_86_1547_0,
    i_8_86_1551_0, i_8_86_1573_0, i_8_86_1634_0, i_8_86_1636_0,
    i_8_86_1645_0, i_8_86_1654_0, i_8_86_1687_0, i_8_86_1707_0,
    i_8_86_1708_0, i_8_86_1723_0, i_8_86_1751_0, i_8_86_1754_0,
    i_8_86_1772_0, i_8_86_1808_0, i_8_86_1858_0, i_8_86_1912_0,
    i_8_86_1966_0, i_8_86_1996_0, i_8_86_2051_0, i_8_86_2152_0,
    i_8_86_2214_0;
  output o_8_86_0_0;
  assign o_8_86_0_0 = 0;
endmodule



// Benchmark "kernel_8_87" written by ABC on Sun Jul 19 10:04:30 2020

module kernel_8_87 ( 
    i_8_87_19_0, i_8_87_22_0, i_8_87_23_0, i_8_87_41_0, i_8_87_73_0,
    i_8_87_74_0, i_8_87_84_0, i_8_87_103_0, i_8_87_167_0, i_8_87_198_0,
    i_8_87_199_0, i_8_87_271_0, i_8_87_272_0, i_8_87_352_0, i_8_87_371_0,
    i_8_87_382_0, i_8_87_388_0, i_8_87_452_0, i_8_87_526_0, i_8_87_532_0,
    i_8_87_549_0, i_8_87_553_0, i_8_87_594_0, i_8_87_630_0, i_8_87_631_0,
    i_8_87_653_0, i_8_87_657_0, i_8_87_685_0, i_8_87_694_0, i_8_87_695_0,
    i_8_87_747_0, i_8_87_819_0, i_8_87_829_0, i_8_87_838_0, i_8_87_860_0,
    i_8_87_875_0, i_8_87_910_0, i_8_87_914_0, i_8_87_919_0, i_8_87_1029_0,
    i_8_87_1110_0, i_8_87_1111_0, i_8_87_1156_0, i_8_87_1198_0,
    i_8_87_1225_0, i_8_87_1233_0, i_8_87_1234_0, i_8_87_1268_0,
    i_8_87_1296_0, i_8_87_1297_0, i_8_87_1315_0, i_8_87_1318_0,
    i_8_87_1332_0, i_8_87_1354_0, i_8_87_1387_0, i_8_87_1390_0,
    i_8_87_1435_0, i_8_87_1458_0, i_8_87_1471_0, i_8_87_1477_0,
    i_8_87_1486_0, i_8_87_1530_0, i_8_87_1534_0, i_8_87_1540_0,
    i_8_87_1547_0, i_8_87_1548_0, i_8_87_1594_0, i_8_87_1595_0,
    i_8_87_1630_0, i_8_87_1631_0, i_8_87_1633_0, i_8_87_1639_0,
    i_8_87_1649_0, i_8_87_1657_0, i_8_87_1773_0, i_8_87_1782_0,
    i_8_87_1784_0, i_8_87_1791_0, i_8_87_1793_0, i_8_87_1818_0,
    i_8_87_1865_0, i_8_87_1873_0, i_8_87_1886_0, i_8_87_1909_0,
    i_8_87_1918_0, i_8_87_1944_0, i_8_87_1947_0, i_8_87_1964_0,
    i_8_87_1972_0, i_8_87_1980_0, i_8_87_2007_0, i_8_87_2063_0,
    i_8_87_2093_0, i_8_87_2107_0, i_8_87_2147_0, i_8_87_2157_0,
    i_8_87_2223_0, i_8_87_2233_0, i_8_87_2243_0, i_8_87_2287_0,
    o_8_87_0_0  );
  input  i_8_87_19_0, i_8_87_22_0, i_8_87_23_0, i_8_87_41_0, i_8_87_73_0,
    i_8_87_74_0, i_8_87_84_0, i_8_87_103_0, i_8_87_167_0, i_8_87_198_0,
    i_8_87_199_0, i_8_87_271_0, i_8_87_272_0, i_8_87_352_0, i_8_87_371_0,
    i_8_87_382_0, i_8_87_388_0, i_8_87_452_0, i_8_87_526_0, i_8_87_532_0,
    i_8_87_549_0, i_8_87_553_0, i_8_87_594_0, i_8_87_630_0, i_8_87_631_0,
    i_8_87_653_0, i_8_87_657_0, i_8_87_685_0, i_8_87_694_0, i_8_87_695_0,
    i_8_87_747_0, i_8_87_819_0, i_8_87_829_0, i_8_87_838_0, i_8_87_860_0,
    i_8_87_875_0, i_8_87_910_0, i_8_87_914_0, i_8_87_919_0, i_8_87_1029_0,
    i_8_87_1110_0, i_8_87_1111_0, i_8_87_1156_0, i_8_87_1198_0,
    i_8_87_1225_0, i_8_87_1233_0, i_8_87_1234_0, i_8_87_1268_0,
    i_8_87_1296_0, i_8_87_1297_0, i_8_87_1315_0, i_8_87_1318_0,
    i_8_87_1332_0, i_8_87_1354_0, i_8_87_1387_0, i_8_87_1390_0,
    i_8_87_1435_0, i_8_87_1458_0, i_8_87_1471_0, i_8_87_1477_0,
    i_8_87_1486_0, i_8_87_1530_0, i_8_87_1534_0, i_8_87_1540_0,
    i_8_87_1547_0, i_8_87_1548_0, i_8_87_1594_0, i_8_87_1595_0,
    i_8_87_1630_0, i_8_87_1631_0, i_8_87_1633_0, i_8_87_1639_0,
    i_8_87_1649_0, i_8_87_1657_0, i_8_87_1773_0, i_8_87_1782_0,
    i_8_87_1784_0, i_8_87_1791_0, i_8_87_1793_0, i_8_87_1818_0,
    i_8_87_1865_0, i_8_87_1873_0, i_8_87_1886_0, i_8_87_1909_0,
    i_8_87_1918_0, i_8_87_1944_0, i_8_87_1947_0, i_8_87_1964_0,
    i_8_87_1972_0, i_8_87_1980_0, i_8_87_2007_0, i_8_87_2063_0,
    i_8_87_2093_0, i_8_87_2107_0, i_8_87_2147_0, i_8_87_2157_0,
    i_8_87_2223_0, i_8_87_2233_0, i_8_87_2243_0, i_8_87_2287_0;
  output o_8_87_0_0;
  assign o_8_87_0_0 = 0;
endmodule



// Benchmark "kernel_8_88" written by ABC on Sun Jul 19 10:04:31 2020

module kernel_8_88 ( 
    i_8_88_93_0, i_8_88_94_0, i_8_88_107_0, i_8_88_143_0, i_8_88_197_0,
    i_8_88_223_0, i_8_88_266_0, i_8_88_283_0, i_8_88_284_0, i_8_88_288_0,
    i_8_88_296_0, i_8_88_299_0, i_8_88_305_0, i_8_88_319_0, i_8_88_322_0,
    i_8_88_328_0, i_8_88_368_0, i_8_88_382_0, i_8_88_404_0, i_8_88_431_0,
    i_8_88_437_0, i_8_88_489_0, i_8_88_492_0, i_8_88_553_0, i_8_88_557_0,
    i_8_88_593_0, i_8_88_599_0, i_8_88_628_0, i_8_88_637_0, i_8_88_643_0,
    i_8_88_656_0, i_8_88_661_0, i_8_88_664_0, i_8_88_724_0, i_8_88_727_0,
    i_8_88_781_0, i_8_88_782_0, i_8_88_790_0, i_8_88_791_0, i_8_88_824_0,
    i_8_88_827_0, i_8_88_840_0, i_8_88_843_0, i_8_88_845_0, i_8_88_930_0,
    i_8_88_931_0, i_8_88_953_0, i_8_88_976_0, i_8_88_991_0, i_8_88_1056_0,
    i_8_88_1075_0, i_8_88_1155_0, i_8_88_1157_0, i_8_88_1214_0,
    i_8_88_1240_0, i_8_88_1273_0, i_8_88_1283_0, i_8_88_1324_0,
    i_8_88_1345_0, i_8_88_1354_0, i_8_88_1366_0, i_8_88_1375_0,
    i_8_88_1390_0, i_8_88_1391_0, i_8_88_1454_0, i_8_88_1483_0,
    i_8_88_1490_0, i_8_88_1592_0, i_8_88_1647_0, i_8_88_1681_0,
    i_8_88_1751_0, i_8_88_1771_0, i_8_88_1789_0, i_8_88_1803_0,
    i_8_88_1806_0, i_8_88_1810_0, i_8_88_1837_0, i_8_88_1853_0,
    i_8_88_1859_0, i_8_88_1893_0, i_8_88_1903_0, i_8_88_1907_0,
    i_8_88_1949_0, i_8_88_1950_0, i_8_88_1994_0, i_8_88_1995_0,
    i_8_88_2046_0, i_8_88_2120_0, i_8_88_2129_0, i_8_88_2132_0,
    i_8_88_2150_0, i_8_88_2174_0, i_8_88_2177_0, i_8_88_2194_0,
    i_8_88_2195_0, i_8_88_2227_0, i_8_88_2248_0, i_8_88_2249_0,
    i_8_88_2282_0, i_8_88_2287_0,
    o_8_88_0_0  );
  input  i_8_88_93_0, i_8_88_94_0, i_8_88_107_0, i_8_88_143_0,
    i_8_88_197_0, i_8_88_223_0, i_8_88_266_0, i_8_88_283_0, i_8_88_284_0,
    i_8_88_288_0, i_8_88_296_0, i_8_88_299_0, i_8_88_305_0, i_8_88_319_0,
    i_8_88_322_0, i_8_88_328_0, i_8_88_368_0, i_8_88_382_0, i_8_88_404_0,
    i_8_88_431_0, i_8_88_437_0, i_8_88_489_0, i_8_88_492_0, i_8_88_553_0,
    i_8_88_557_0, i_8_88_593_0, i_8_88_599_0, i_8_88_628_0, i_8_88_637_0,
    i_8_88_643_0, i_8_88_656_0, i_8_88_661_0, i_8_88_664_0, i_8_88_724_0,
    i_8_88_727_0, i_8_88_781_0, i_8_88_782_0, i_8_88_790_0, i_8_88_791_0,
    i_8_88_824_0, i_8_88_827_0, i_8_88_840_0, i_8_88_843_0, i_8_88_845_0,
    i_8_88_930_0, i_8_88_931_0, i_8_88_953_0, i_8_88_976_0, i_8_88_991_0,
    i_8_88_1056_0, i_8_88_1075_0, i_8_88_1155_0, i_8_88_1157_0,
    i_8_88_1214_0, i_8_88_1240_0, i_8_88_1273_0, i_8_88_1283_0,
    i_8_88_1324_0, i_8_88_1345_0, i_8_88_1354_0, i_8_88_1366_0,
    i_8_88_1375_0, i_8_88_1390_0, i_8_88_1391_0, i_8_88_1454_0,
    i_8_88_1483_0, i_8_88_1490_0, i_8_88_1592_0, i_8_88_1647_0,
    i_8_88_1681_0, i_8_88_1751_0, i_8_88_1771_0, i_8_88_1789_0,
    i_8_88_1803_0, i_8_88_1806_0, i_8_88_1810_0, i_8_88_1837_0,
    i_8_88_1853_0, i_8_88_1859_0, i_8_88_1893_0, i_8_88_1903_0,
    i_8_88_1907_0, i_8_88_1949_0, i_8_88_1950_0, i_8_88_1994_0,
    i_8_88_1995_0, i_8_88_2046_0, i_8_88_2120_0, i_8_88_2129_0,
    i_8_88_2132_0, i_8_88_2150_0, i_8_88_2174_0, i_8_88_2177_0,
    i_8_88_2194_0, i_8_88_2195_0, i_8_88_2227_0, i_8_88_2248_0,
    i_8_88_2249_0, i_8_88_2282_0, i_8_88_2287_0;
  output o_8_88_0_0;
  assign o_8_88_0_0 = 0;
endmodule



// Benchmark "kernel_8_89" written by ABC on Sun Jul 19 10:04:32 2020

module kernel_8_89 ( 
    i_8_89_23_0, i_8_89_34_0, i_8_89_35_0, i_8_89_96_0, i_8_89_106_0,
    i_8_89_141_0, i_8_89_142_0, i_8_89_160_0, i_8_89_161_0, i_8_89_187_0,
    i_8_89_201_0, i_8_89_204_0, i_8_89_206_0, i_8_89_220_0, i_8_89_257_0,
    i_8_89_289_0, i_8_89_302_0, i_8_89_305_0, i_8_89_328_0, i_8_89_345_0,
    i_8_89_346_0, i_8_89_367_0, i_8_89_373_0, i_8_89_440_0, i_8_89_458_0,
    i_8_89_463_0, i_8_89_610_0, i_8_89_615_0, i_8_89_617_0, i_8_89_628_0,
    i_8_89_697_0, i_8_89_782_0, i_8_89_984_0, i_8_89_985_0, i_8_89_991_0,
    i_8_89_992_0, i_8_89_993_0, i_8_89_994_0, i_8_89_1014_0, i_8_89_1087_0,
    i_8_89_1112_0, i_8_89_1114_0, i_8_89_1135_0, i_8_89_1136_0,
    i_8_89_1138_0, i_8_89_1189_0, i_8_89_1192_0, i_8_89_1270_0,
    i_8_89_1271_0, i_8_89_1273_0, i_8_89_1306_0, i_8_89_1344_0,
    i_8_89_1397_0, i_8_89_1417_0, i_8_89_1434_0, i_8_89_1436_0,
    i_8_89_1438_0, i_8_89_1511_0, i_8_89_1537_0, i_8_89_1541_0,
    i_8_89_1542_0, i_8_89_1544_0, i_8_89_1564_0, i_8_89_1578_0,
    i_8_89_1612_0, i_8_89_1616_0, i_8_89_1629_0, i_8_89_1631_0,
    i_8_89_1714_0, i_8_89_1715_0, i_8_89_1723_0, i_8_89_1726_0,
    i_8_89_1727_0, i_8_89_1736_0, i_8_89_1801_0, i_8_89_1804_0,
    i_8_89_1807_0, i_8_89_1810_0, i_8_89_1812_0, i_8_89_1831_0,
    i_8_89_1838_0, i_8_89_1840_0, i_8_89_1841_0, i_8_89_1858_0,
    i_8_89_1922_0, i_8_89_2002_0, i_8_89_2015_0, i_8_89_2049_0,
    i_8_89_2050_0, i_8_89_2051_0, i_8_89_2134_0, i_8_89_2150_0,
    i_8_89_2182_0, i_8_89_2215_0, i_8_89_2230_0, i_8_89_2260_0,
    i_8_89_2261_0, i_8_89_2264_0, i_8_89_2272_0, i_8_89_2282_0,
    o_8_89_0_0  );
  input  i_8_89_23_0, i_8_89_34_0, i_8_89_35_0, i_8_89_96_0,
    i_8_89_106_0, i_8_89_141_0, i_8_89_142_0, i_8_89_160_0, i_8_89_161_0,
    i_8_89_187_0, i_8_89_201_0, i_8_89_204_0, i_8_89_206_0, i_8_89_220_0,
    i_8_89_257_0, i_8_89_289_0, i_8_89_302_0, i_8_89_305_0, i_8_89_328_0,
    i_8_89_345_0, i_8_89_346_0, i_8_89_367_0, i_8_89_373_0, i_8_89_440_0,
    i_8_89_458_0, i_8_89_463_0, i_8_89_610_0, i_8_89_615_0, i_8_89_617_0,
    i_8_89_628_0, i_8_89_697_0, i_8_89_782_0, i_8_89_984_0, i_8_89_985_0,
    i_8_89_991_0, i_8_89_992_0, i_8_89_993_0, i_8_89_994_0, i_8_89_1014_0,
    i_8_89_1087_0, i_8_89_1112_0, i_8_89_1114_0, i_8_89_1135_0,
    i_8_89_1136_0, i_8_89_1138_0, i_8_89_1189_0, i_8_89_1192_0,
    i_8_89_1270_0, i_8_89_1271_0, i_8_89_1273_0, i_8_89_1306_0,
    i_8_89_1344_0, i_8_89_1397_0, i_8_89_1417_0, i_8_89_1434_0,
    i_8_89_1436_0, i_8_89_1438_0, i_8_89_1511_0, i_8_89_1537_0,
    i_8_89_1541_0, i_8_89_1542_0, i_8_89_1544_0, i_8_89_1564_0,
    i_8_89_1578_0, i_8_89_1612_0, i_8_89_1616_0, i_8_89_1629_0,
    i_8_89_1631_0, i_8_89_1714_0, i_8_89_1715_0, i_8_89_1723_0,
    i_8_89_1726_0, i_8_89_1727_0, i_8_89_1736_0, i_8_89_1801_0,
    i_8_89_1804_0, i_8_89_1807_0, i_8_89_1810_0, i_8_89_1812_0,
    i_8_89_1831_0, i_8_89_1838_0, i_8_89_1840_0, i_8_89_1841_0,
    i_8_89_1858_0, i_8_89_1922_0, i_8_89_2002_0, i_8_89_2015_0,
    i_8_89_2049_0, i_8_89_2050_0, i_8_89_2051_0, i_8_89_2134_0,
    i_8_89_2150_0, i_8_89_2182_0, i_8_89_2215_0, i_8_89_2230_0,
    i_8_89_2260_0, i_8_89_2261_0, i_8_89_2264_0, i_8_89_2272_0,
    i_8_89_2282_0;
  output o_8_89_0_0;
  assign o_8_89_0_0 = ~((~i_8_89_201_0 & ((~i_8_89_206_0 & i_8_89_610_0 & ~i_8_89_984_0 & ~i_8_89_1397_0 & ~i_8_89_1631_0 & ~i_8_89_1812_0) | (~i_8_89_34_0 & ~i_8_89_96_0 & ~i_8_89_160_0 & ~i_8_89_1714_0 & ~i_8_89_2050_0 & ~i_8_89_2051_0 & ~i_8_89_2134_0))) | (~i_8_89_96_0 & ((~i_8_89_204_0 & ~i_8_89_991_0 & ~i_8_89_994_0 & ~i_8_89_1135_0 & ~i_8_89_1138_0 & ~i_8_89_1736_0) | (~i_8_89_141_0 & ~i_8_89_161_0 & ~i_8_89_373_0 & i_8_89_610_0 & ~i_8_89_985_0 & ~i_8_89_1629_0 & ~i_8_89_1726_0 & i_8_89_1922_0))) | (~i_8_89_141_0 & ((~i_8_89_204_0 & i_8_89_220_0 & ~i_8_89_1135_0 & ~i_8_89_1629_0 & ~i_8_89_1715_0 & ~i_8_89_1727_0 & ~i_8_89_2049_0 & ~i_8_89_2050_0) | (~i_8_89_35_0 & ~i_8_89_440_0 & ~i_8_89_615_0 & ~i_8_89_782_0 & ~i_8_89_984_0 & ~i_8_89_1397_0 & ~i_8_89_2002_0 & ~i_8_89_2015_0 & ~i_8_89_2051_0 & ~i_8_89_2230_0))) | (~i_8_89_160_0 & ((~i_8_89_142_0 & ~i_8_89_992_0 & i_8_89_1138_0 & ~i_8_89_1306_0 & ~i_8_89_1511_0 & ~i_8_89_1715_0 & ~i_8_89_2015_0 & ~i_8_89_2215_0 & ~i_8_89_2230_0) | (~i_8_89_34_0 & ~i_8_89_161_0 & ~i_8_89_1135_0 & i_8_89_2230_0 & ~i_8_89_2260_0 & ~i_8_89_2261_0))) | (~i_8_89_34_0 & ((i_8_89_346_0 & ~i_8_89_782_0 & ~i_8_89_1087_0 & ~i_8_89_1397_0) | (~i_8_89_991_0 & ~i_8_89_1014_0 & ~i_8_89_1629_0 & ~i_8_89_1715_0 & i_8_89_2182_0))) | (~i_8_89_142_0 & ((i_8_89_345_0 & ~i_8_89_985_0 & ~i_8_89_1714_0) | (~i_8_89_35_0 & ~i_8_89_204_0 & ~i_8_89_328_0 & ~i_8_89_1616_0 & ~i_8_89_1629_0 & ~i_8_89_2049_0 & ~i_8_89_2260_0 & ~i_8_89_2264_0))) | (~i_8_89_1344_0 & ((~i_8_89_35_0 & ~i_8_89_1616_0 & ~i_8_89_2261_0 & ((~i_8_89_220_0 & ~i_8_89_628_0 & ~i_8_89_2015_0) | (~i_8_89_1087_0 & ~i_8_89_1438_0 & ~i_8_89_1714_0 & ~i_8_89_1812_0 & ~i_8_89_2260_0))) | (i_8_89_697_0 & ~i_8_89_984_0 & ~i_8_89_992_0 & ~i_8_89_993_0 & ~i_8_89_1564_0 & ~i_8_89_1631_0 & ~i_8_89_2051_0))) | (~i_8_89_204_0 & ~i_8_89_2264_0 & ((~i_8_89_302_0 & ~i_8_89_458_0 & ~i_8_89_628_0 & ~i_8_89_1136_0 & ~i_8_89_1138_0 & ~i_8_89_1612_0 & ~i_8_89_1715_0 & ~i_8_89_2002_0) | (~i_8_89_257_0 & ~i_8_89_697_0 & ~i_8_89_984_0 & ~i_8_89_993_0 & ~i_8_89_1397_0 & ~i_8_89_1723_0 & ~i_8_89_1727_0 & ~i_8_89_2230_0 & ~i_8_89_2261_0))) | (~i_8_89_1436_0 & ~i_8_89_2230_0 & ((~i_8_89_187_0 & ~i_8_89_782_0 & ~i_8_89_984_0 & ~i_8_89_991_0 & ~i_8_89_1136_0 & ~i_8_89_1564_0 & ~i_8_89_2049_0) | (~i_8_89_161_0 & ~i_8_89_302_0 & ~i_8_89_458_0 & i_8_89_1544_0 & ~i_8_89_2215_0))) | (i_8_89_463_0 & i_8_89_1840_0 & ~i_8_89_1922_0) | (~i_8_89_440_0 & ~i_8_89_1014_0 & ~i_8_89_1715_0 & ~i_8_89_1727_0 & ~i_8_89_1810_0 & ~i_8_89_2049_0 & ~i_8_89_2260_0));
endmodule



// Benchmark "kernel_8_90" written by ABC on Sun Jul 19 10:04:33 2020

module kernel_8_90 ( 
    i_8_90_11_0, i_8_90_40_0, i_8_90_48_0, i_8_90_57_0, i_8_90_88_0,
    i_8_90_115_0, i_8_90_120_0, i_8_90_127_0, i_8_90_138_0, i_8_90_146_0,
    i_8_90_165_0, i_8_90_191_0, i_8_90_203_0, i_8_90_226_0, i_8_90_228_0,
    i_8_90_236_0, i_8_90_283_0, i_8_90_285_0, i_8_90_295_0, i_8_90_321_0,
    i_8_90_328_0, i_8_90_331_0, i_8_90_336_0, i_8_90_363_0, i_8_90_373_0,
    i_8_90_383_0, i_8_90_386_0, i_8_90_398_0, i_8_90_403_0, i_8_90_420_0,
    i_8_90_453_0, i_8_90_526_0, i_8_90_555_0, i_8_90_571_0, i_8_90_609_0,
    i_8_90_627_0, i_8_90_654_0, i_8_90_662_0, i_8_90_665_0, i_8_90_696_0,
    i_8_90_700_0, i_8_90_739_0, i_8_90_771_0, i_8_90_779_0, i_8_90_788_0,
    i_8_90_794_0, i_8_90_857_0, i_8_90_917_0, i_8_90_966_0, i_8_90_1059_0,
    i_8_90_1068_0, i_8_90_1118_0, i_8_90_1138_0, i_8_90_1235_0,
    i_8_90_1238_0, i_8_90_1253_0, i_8_90_1300_0, i_8_90_1319_0,
    i_8_90_1324_0, i_8_90_1353_0, i_8_90_1357_0, i_8_90_1408_0,
    i_8_90_1451_0, i_8_90_1455_0, i_8_90_1473_0, i_8_90_1534_0,
    i_8_90_1545_0, i_8_90_1547_0, i_8_90_1605_0, i_8_90_1606_0,
    i_8_90_1617_0, i_8_90_1623_0, i_8_90_1635_0, i_8_90_1649_0,
    i_8_90_1669_0, i_8_90_1708_0, i_8_90_1731_0, i_8_90_1732_0,
    i_8_90_1739_0, i_8_90_1770_0, i_8_90_1784_0, i_8_90_1830_0,
    i_8_90_1867_0, i_8_90_1886_0, i_8_90_1969_0, i_8_90_1983_0,
    i_8_90_2118_0, i_8_90_2127_0, i_8_90_2145_0, i_8_90_2149_0,
    i_8_90_2208_0, i_8_90_2211_0, i_8_90_2212_0, i_8_90_2218_0,
    i_8_90_2229_0, i_8_90_2238_0, i_8_90_2244_0, i_8_90_2245_0,
    i_8_90_2247_0, i_8_90_2248_0,
    o_8_90_0_0  );
  input  i_8_90_11_0, i_8_90_40_0, i_8_90_48_0, i_8_90_57_0, i_8_90_88_0,
    i_8_90_115_0, i_8_90_120_0, i_8_90_127_0, i_8_90_138_0, i_8_90_146_0,
    i_8_90_165_0, i_8_90_191_0, i_8_90_203_0, i_8_90_226_0, i_8_90_228_0,
    i_8_90_236_0, i_8_90_283_0, i_8_90_285_0, i_8_90_295_0, i_8_90_321_0,
    i_8_90_328_0, i_8_90_331_0, i_8_90_336_0, i_8_90_363_0, i_8_90_373_0,
    i_8_90_383_0, i_8_90_386_0, i_8_90_398_0, i_8_90_403_0, i_8_90_420_0,
    i_8_90_453_0, i_8_90_526_0, i_8_90_555_0, i_8_90_571_0, i_8_90_609_0,
    i_8_90_627_0, i_8_90_654_0, i_8_90_662_0, i_8_90_665_0, i_8_90_696_0,
    i_8_90_700_0, i_8_90_739_0, i_8_90_771_0, i_8_90_779_0, i_8_90_788_0,
    i_8_90_794_0, i_8_90_857_0, i_8_90_917_0, i_8_90_966_0, i_8_90_1059_0,
    i_8_90_1068_0, i_8_90_1118_0, i_8_90_1138_0, i_8_90_1235_0,
    i_8_90_1238_0, i_8_90_1253_0, i_8_90_1300_0, i_8_90_1319_0,
    i_8_90_1324_0, i_8_90_1353_0, i_8_90_1357_0, i_8_90_1408_0,
    i_8_90_1451_0, i_8_90_1455_0, i_8_90_1473_0, i_8_90_1534_0,
    i_8_90_1545_0, i_8_90_1547_0, i_8_90_1605_0, i_8_90_1606_0,
    i_8_90_1617_0, i_8_90_1623_0, i_8_90_1635_0, i_8_90_1649_0,
    i_8_90_1669_0, i_8_90_1708_0, i_8_90_1731_0, i_8_90_1732_0,
    i_8_90_1739_0, i_8_90_1770_0, i_8_90_1784_0, i_8_90_1830_0,
    i_8_90_1867_0, i_8_90_1886_0, i_8_90_1969_0, i_8_90_1983_0,
    i_8_90_2118_0, i_8_90_2127_0, i_8_90_2145_0, i_8_90_2149_0,
    i_8_90_2208_0, i_8_90_2211_0, i_8_90_2212_0, i_8_90_2218_0,
    i_8_90_2229_0, i_8_90_2238_0, i_8_90_2244_0, i_8_90_2245_0,
    i_8_90_2247_0, i_8_90_2248_0;
  output o_8_90_0_0;
  assign o_8_90_0_0 = 0;
endmodule



// Benchmark "kernel_8_91" written by ABC on Sun Jul 19 10:04:34 2020

module kernel_8_91 ( 
    i_8_91_22_0, i_8_91_25_0, i_8_91_28_0, i_8_91_63_0, i_8_91_67_0,
    i_8_91_80_0, i_8_91_144_0, i_8_91_172_0, i_8_91_303_0, i_8_91_318_0,
    i_8_91_351_0, i_8_91_352_0, i_8_91_360_0, i_8_91_364_0, i_8_91_379_0,
    i_8_91_401_0, i_8_91_421_0, i_8_91_441_0, i_8_91_513_0, i_8_91_514_0,
    i_8_91_522_0, i_8_91_557_0, i_8_91_571_0, i_8_91_631_0, i_8_91_644_0,
    i_8_91_657_0, i_8_91_666_0, i_8_91_667_0, i_8_91_676_0, i_8_91_697_0,
    i_8_91_702_0, i_8_91_703_0, i_8_91_766_0, i_8_91_824_0, i_8_91_846_0,
    i_8_91_880_0, i_8_91_949_0, i_8_91_955_0, i_8_91_956_0, i_8_91_1047_0,
    i_8_91_1057_0, i_8_91_1107_0, i_8_91_1115_0, i_8_91_1170_0,
    i_8_91_1180_0, i_8_91_1201_0, i_8_91_1228_0, i_8_91_1231_0,
    i_8_91_1269_0, i_8_91_1270_0, i_8_91_1296_0, i_8_91_1351_0,
    i_8_91_1353_0, i_8_91_1355_0, i_8_91_1386_0, i_8_91_1396_0,
    i_8_91_1404_0, i_8_91_1408_0, i_8_91_1434_0, i_8_91_1462_0,
    i_8_91_1463_0, i_8_91_1467_0, i_8_91_1494_0, i_8_91_1497_0,
    i_8_91_1535_0, i_8_91_1562_0, i_8_91_1631_0, i_8_91_1632_0,
    i_8_91_1634_0, i_8_91_1656_0, i_8_91_1701_0, i_8_91_1702_0,
    i_8_91_1746_0, i_8_91_1767_0, i_8_91_1768_0, i_8_91_1769_0,
    i_8_91_1780_0, i_8_91_1791_0, i_8_91_1794_0, i_8_91_1809_0,
    i_8_91_1822_0, i_8_91_1831_0, i_8_91_1845_0, i_8_91_1849_0,
    i_8_91_1863_0, i_8_91_1867_0, i_8_91_1872_0, i_8_91_1901_0,
    i_8_91_1944_0, i_8_91_1993_0, i_8_91_2034_0, i_8_91_2043_0,
    i_8_91_2065_0, i_8_91_2089_0, i_8_91_2135_0, i_8_91_2142_0,
    i_8_91_2147_0, i_8_91_2223_0, i_8_91_2226_0, i_8_91_2274_0,
    o_8_91_0_0  );
  input  i_8_91_22_0, i_8_91_25_0, i_8_91_28_0, i_8_91_63_0, i_8_91_67_0,
    i_8_91_80_0, i_8_91_144_0, i_8_91_172_0, i_8_91_303_0, i_8_91_318_0,
    i_8_91_351_0, i_8_91_352_0, i_8_91_360_0, i_8_91_364_0, i_8_91_379_0,
    i_8_91_401_0, i_8_91_421_0, i_8_91_441_0, i_8_91_513_0, i_8_91_514_0,
    i_8_91_522_0, i_8_91_557_0, i_8_91_571_0, i_8_91_631_0, i_8_91_644_0,
    i_8_91_657_0, i_8_91_666_0, i_8_91_667_0, i_8_91_676_0, i_8_91_697_0,
    i_8_91_702_0, i_8_91_703_0, i_8_91_766_0, i_8_91_824_0, i_8_91_846_0,
    i_8_91_880_0, i_8_91_949_0, i_8_91_955_0, i_8_91_956_0, i_8_91_1047_0,
    i_8_91_1057_0, i_8_91_1107_0, i_8_91_1115_0, i_8_91_1170_0,
    i_8_91_1180_0, i_8_91_1201_0, i_8_91_1228_0, i_8_91_1231_0,
    i_8_91_1269_0, i_8_91_1270_0, i_8_91_1296_0, i_8_91_1351_0,
    i_8_91_1353_0, i_8_91_1355_0, i_8_91_1386_0, i_8_91_1396_0,
    i_8_91_1404_0, i_8_91_1408_0, i_8_91_1434_0, i_8_91_1462_0,
    i_8_91_1463_0, i_8_91_1467_0, i_8_91_1494_0, i_8_91_1497_0,
    i_8_91_1535_0, i_8_91_1562_0, i_8_91_1631_0, i_8_91_1632_0,
    i_8_91_1634_0, i_8_91_1656_0, i_8_91_1701_0, i_8_91_1702_0,
    i_8_91_1746_0, i_8_91_1767_0, i_8_91_1768_0, i_8_91_1769_0,
    i_8_91_1780_0, i_8_91_1791_0, i_8_91_1794_0, i_8_91_1809_0,
    i_8_91_1822_0, i_8_91_1831_0, i_8_91_1845_0, i_8_91_1849_0,
    i_8_91_1863_0, i_8_91_1867_0, i_8_91_1872_0, i_8_91_1901_0,
    i_8_91_1944_0, i_8_91_1993_0, i_8_91_2034_0, i_8_91_2043_0,
    i_8_91_2065_0, i_8_91_2089_0, i_8_91_2135_0, i_8_91_2142_0,
    i_8_91_2147_0, i_8_91_2223_0, i_8_91_2226_0, i_8_91_2274_0;
  output o_8_91_0_0;
  assign o_8_91_0_0 = 0;
endmodule



// Benchmark "kernel_8_92" written by ABC on Sun Jul 19 10:04:35 2020

module kernel_8_92 ( 
    i_8_92_77_0, i_8_92_80_0, i_8_92_119_0, i_8_92_163_0, i_8_92_220_0,
    i_8_92_314_0, i_8_92_363_0, i_8_92_364_0, i_8_92_366_0, i_8_92_367_0,
    i_8_92_370_0, i_8_92_381_0, i_8_92_484_0, i_8_92_487_0, i_8_92_489_0,
    i_8_92_490_0, i_8_92_492_0, i_8_92_493_0, i_8_92_494_0, i_8_92_507_0,
    i_8_92_509_0, i_8_92_523_0, i_8_92_524_0, i_8_92_527_0, i_8_92_554_0,
    i_8_92_556_0, i_8_92_597_0, i_8_92_604_0, i_8_92_637_0, i_8_92_638_0,
    i_8_92_691_0, i_8_92_693_0, i_8_92_694_0, i_8_92_695_0, i_8_92_698_0,
    i_8_92_699_0, i_8_92_760_0, i_8_92_827_0, i_8_92_838_0, i_8_92_841_0,
    i_8_92_843_0, i_8_92_851_0, i_8_92_880_0, i_8_92_964_0, i_8_92_1027_0,
    i_8_92_1072_0, i_8_92_1110_0, i_8_92_1113_0, i_8_92_1255_0,
    i_8_92_1263_0, i_8_92_1265_0, i_8_92_1296_0, i_8_92_1301_0,
    i_8_92_1339_0, i_8_92_1355_0, i_8_92_1369_0, i_8_92_1370_0,
    i_8_92_1372_0, i_8_92_1373_0, i_8_92_1398_0, i_8_92_1399_0,
    i_8_92_1400_0, i_8_92_1437_0, i_8_92_1438_0, i_8_92_1439_0,
    i_8_92_1455_0, i_8_92_1468_0, i_8_92_1535_0, i_8_92_1620_0,
    i_8_92_1621_0, i_8_92_1623_0, i_8_92_1624_0, i_8_92_1625_0,
    i_8_92_1628_0, i_8_92_1629_0, i_8_92_1632_0, i_8_92_1634_0,
    i_8_92_1672_0, i_8_92_1693_0, i_8_92_1733_0, i_8_92_1746_0,
    i_8_92_1747_0, i_8_92_1748_0, i_8_92_1749_0, i_8_92_1752_0,
    i_8_92_1753_0, i_8_92_1763_0, i_8_92_1825_0, i_8_92_1826_0,
    i_8_92_1854_0, i_8_92_1861_0, i_8_92_1888_0, i_8_92_1900_0,
    i_8_92_1904_0, i_8_92_1945_0, i_8_92_1996_0, i_8_92_2171_0,
    i_8_92_2241_0, i_8_92_2246_0, i_8_92_2276_0,
    o_8_92_0_0  );
  input  i_8_92_77_0, i_8_92_80_0, i_8_92_119_0, i_8_92_163_0,
    i_8_92_220_0, i_8_92_314_0, i_8_92_363_0, i_8_92_364_0, i_8_92_366_0,
    i_8_92_367_0, i_8_92_370_0, i_8_92_381_0, i_8_92_484_0, i_8_92_487_0,
    i_8_92_489_0, i_8_92_490_0, i_8_92_492_0, i_8_92_493_0, i_8_92_494_0,
    i_8_92_507_0, i_8_92_509_0, i_8_92_523_0, i_8_92_524_0, i_8_92_527_0,
    i_8_92_554_0, i_8_92_556_0, i_8_92_597_0, i_8_92_604_0, i_8_92_637_0,
    i_8_92_638_0, i_8_92_691_0, i_8_92_693_0, i_8_92_694_0, i_8_92_695_0,
    i_8_92_698_0, i_8_92_699_0, i_8_92_760_0, i_8_92_827_0, i_8_92_838_0,
    i_8_92_841_0, i_8_92_843_0, i_8_92_851_0, i_8_92_880_0, i_8_92_964_0,
    i_8_92_1027_0, i_8_92_1072_0, i_8_92_1110_0, i_8_92_1113_0,
    i_8_92_1255_0, i_8_92_1263_0, i_8_92_1265_0, i_8_92_1296_0,
    i_8_92_1301_0, i_8_92_1339_0, i_8_92_1355_0, i_8_92_1369_0,
    i_8_92_1370_0, i_8_92_1372_0, i_8_92_1373_0, i_8_92_1398_0,
    i_8_92_1399_0, i_8_92_1400_0, i_8_92_1437_0, i_8_92_1438_0,
    i_8_92_1439_0, i_8_92_1455_0, i_8_92_1468_0, i_8_92_1535_0,
    i_8_92_1620_0, i_8_92_1621_0, i_8_92_1623_0, i_8_92_1624_0,
    i_8_92_1625_0, i_8_92_1628_0, i_8_92_1629_0, i_8_92_1632_0,
    i_8_92_1634_0, i_8_92_1672_0, i_8_92_1693_0, i_8_92_1733_0,
    i_8_92_1746_0, i_8_92_1747_0, i_8_92_1748_0, i_8_92_1749_0,
    i_8_92_1752_0, i_8_92_1753_0, i_8_92_1763_0, i_8_92_1825_0,
    i_8_92_1826_0, i_8_92_1854_0, i_8_92_1861_0, i_8_92_1888_0,
    i_8_92_1900_0, i_8_92_1904_0, i_8_92_1945_0, i_8_92_1996_0,
    i_8_92_2171_0, i_8_92_2241_0, i_8_92_2246_0, i_8_92_2276_0;
  output o_8_92_0_0;
  assign o_8_92_0_0 = ~((~i_8_92_1693_0 & ((~i_8_92_1370_0 & ((~i_8_92_119_0 & ~i_8_92_1900_0 & ((~i_8_92_80_0 & ~i_8_92_492_0 & ~i_8_92_693_0 & ~i_8_92_695_0 & ~i_8_92_843_0 & ~i_8_92_880_0 & ~i_8_92_1027_0 & ~i_8_92_1296_0 & ~i_8_92_1399_0 & ~i_8_92_1620_0 & ~i_8_92_1628_0 & ~i_8_92_1733_0 & ~i_8_92_1945_0) | (~i_8_92_367_0 & ~i_8_92_381_0 & ~i_8_92_489_0 & ~i_8_92_698_0 & ~i_8_92_838_0 & ~i_8_92_1263_0 & ~i_8_92_1369_0 & ~i_8_92_1455_0 & ~i_8_92_1623_0 & ~i_8_92_1625_0 & ~i_8_92_1904_0 & ~i_8_92_2246_0 & ~i_8_92_2276_0))) | (~i_8_92_364_0 & ~i_8_92_366_0 & ~i_8_92_487_0 & ~i_8_92_492_0 & ~i_8_92_694_0 & ~i_8_92_698_0 & ~i_8_92_964_0 & ~i_8_92_1263_0 & ~i_8_92_1535_0 & ~i_8_92_1628_0))) | (i_8_92_77_0 & ~i_8_92_163_0 & ~i_8_92_1369_0 & ~i_8_92_1621_0 & i_8_92_1748_0) | (~i_8_92_366_0 & i_8_92_507_0 & ~i_8_92_1672_0 & ~i_8_92_1854_0 & ~i_8_92_1900_0) | (i_8_92_1265_0 & i_8_92_1535_0 & ~i_8_92_1620_0 & i_8_92_2241_0))) | (~i_8_92_119_0 & ((~i_8_92_1370_0 & ((~i_8_92_314_0 & ((i_8_92_509_0 & ~i_8_92_1373_0 & ~i_8_92_1621_0) | (i_8_92_523_0 & ~i_8_92_637_0 & ~i_8_92_838_0 & ~i_8_92_1027_0 & ~i_8_92_1255_0 & ~i_8_92_1369_0 & ~i_8_92_1372_0 & ~i_8_92_1455_0 & ~i_8_92_1468_0 & ~i_8_92_1825_0 & ~i_8_92_1854_0))) | (~i_8_92_487_0 & ~i_8_92_493_0 & ~i_8_92_698_0 & ~i_8_92_843_0 & ~i_8_92_1027_0 & ~i_8_92_1263_0 & ~i_8_92_1623_0 & ~i_8_92_1628_0 & ~i_8_92_1854_0))) | (~i_8_92_364_0 & ~i_8_92_487_0 & ~i_8_92_490_0 & ~i_8_92_492_0 & i_8_92_1263_0 & ~i_8_92_1369_0 & ~i_8_92_1468_0 & ~i_8_92_1733_0 & ~i_8_92_1888_0) | (i_8_92_509_0 & ~i_8_92_691_0 & i_8_92_1301_0 & ~i_8_92_1900_0 & ~i_8_92_2241_0))) | (~i_8_92_490_0 & ((~i_8_92_693_0 & ~i_8_92_1296_0 & ~i_8_92_1620_0 & ~i_8_92_1624_0 & ~i_8_92_1625_0 & i_8_92_1747_0) | (~i_8_92_163_0 & ~i_8_92_314_0 & ~i_8_92_523_0 & ~i_8_92_527_0 & ~i_8_92_1370_0 & ~i_8_92_1373_0 & i_8_92_2171_0))) | (~i_8_92_163_0 & ((~i_8_92_487_0 & ~i_8_92_494_0 & ~i_8_92_841_0 & i_8_92_1265_0 & ~i_8_92_1370_0 & ~i_8_92_1625_0) | (i_8_92_523_0 & ~i_8_92_698_0 & ~i_8_92_1296_0 & i_8_92_1438_0 & ~i_8_92_1825_0))) | (~i_8_92_487_0 & ((~i_8_92_367_0 & ~i_8_92_843_0 & ~i_8_92_880_0 & ~i_8_92_1373_0 & i_8_92_1439_0 & i_8_92_1628_0) | (i_8_92_1110_0 & i_8_92_1746_0))) | (~i_8_92_1623_0 & ((~i_8_92_367_0 & ((i_8_92_489_0 & i_8_92_493_0 & ~i_8_92_699_0 & ~i_8_92_1854_0) | (~i_8_92_489_0 & ~i_8_92_1455_0 & ~i_8_92_1621_0 & ~i_8_92_1625_0 & i_8_92_1753_0 & ~i_8_92_1904_0))) | (~i_8_92_694_0 & ~i_8_92_1628_0 & ((~i_8_92_843_0 & i_8_92_851_0 & ~i_8_92_1400_0 & ~i_8_92_1904_0) | (i_8_92_80_0 & ~i_8_92_364_0 & ~i_8_92_527_0 & ~i_8_92_2171_0))) | (i_8_92_366_0 & ~i_8_92_1620_0 & ~i_8_92_1624_0 & i_8_92_1632_0) | (i_8_92_638_0 & ~i_8_92_880_0 & ~i_8_92_1621_0 & ~i_8_92_1749_0 & i_8_92_1888_0))) | (i_8_92_80_0 & ((~i_8_92_493_0 & ~i_8_92_693_0 & ~i_8_92_1369_0 & ~i_8_92_1455_0 & ~i_8_92_1625_0) | (i_8_92_220_0 & ~i_8_92_1621_0 & i_8_92_1825_0))) | (~i_8_92_694_0 & ((~i_8_92_693_0 & ((~i_8_92_494_0 & ((~i_8_92_314_0 & ~i_8_92_492_0 & i_8_92_880_0 & ~i_8_92_1398_0 & ~i_8_92_1621_0 & ~i_8_92_1625_0 & ~i_8_92_1672_0 & ~i_8_92_1888_0 & ~i_8_92_1900_0) | (~i_8_92_493_0 & ~i_8_92_695_0 & ~i_8_92_698_0 & ~i_8_92_699_0 & ~i_8_92_964_0 & ~i_8_92_1296_0 & ~i_8_92_1372_0 & ~i_8_92_1373_0 & ~i_8_92_1854_0 & ~i_8_92_1996_0))) | (~i_8_92_381_0 & ~i_8_92_699_0 & ~i_8_92_964_0 & ~i_8_92_1372_0 & i_8_92_1753_0 & ~i_8_92_1904_0))) | (~i_8_92_1255_0 & ~i_8_92_1373_0 & ~i_8_92_1624_0 & ~i_8_92_1747_0 & i_8_92_1749_0))) | (~i_8_92_314_0 & ((~i_8_92_492_0 & ~i_8_92_1255_0 & i_8_92_1399_0 & ~i_8_92_1854_0 & ~i_8_92_1900_0 & ~i_8_92_1624_0 & ~i_8_92_1625_0) | (~i_8_92_364_0 & i_8_92_527_0 & ~i_8_92_843_0 & ~i_8_92_964_0 & ~i_8_92_1370_0 & ~i_8_92_1888_0 & ~i_8_92_1996_0 & ~i_8_92_2241_0 & ~i_8_92_2276_0))) | (~i_8_92_364_0 & ((~i_8_92_363_0 & i_8_92_1398_0 & ~i_8_92_1861_0) | (~i_8_92_1263_0 & i_8_92_1746_0 & ~i_8_92_1900_0))) | (~i_8_92_1624_0 & ((~i_8_92_363_0 & ((~i_8_92_851_0 & i_8_92_1265_0 & i_8_92_1355_0 & ~i_8_92_1620_0 & ~i_8_92_1861_0) | (i_8_92_490_0 & ~i_8_92_698_0 & i_8_92_1438_0 & i_8_92_1825_0 & ~i_8_92_2276_0))) | (~i_8_92_493_0 & ~i_8_92_1369_0 & ~i_8_92_1370_0 & ~i_8_92_1621_0 & i_8_92_1629_0 & ~i_8_92_1904_0))) | (~i_8_92_492_0 & ((i_8_92_1632_0 & ~i_8_92_1854_0) | (~i_8_92_381_0 & ~i_8_92_493_0 & ~i_8_92_554_0 & ~i_8_92_597_0 & ~i_8_92_1072_0 & i_8_92_1110_0 & ~i_8_92_1263_0 & ~i_8_92_1265_0 & ~i_8_92_1399_0 & ~i_8_92_1439_0 & ~i_8_92_1455_0 & ~i_8_92_1900_0))) | (~i_8_92_1372_0 & ((~i_8_92_381_0 & ((~i_8_92_493_0 & ~i_8_92_698_0 & ~i_8_92_1296_0 & ~i_8_92_1370_0 & i_8_92_1747_0 & ~i_8_92_1854_0) | (~i_8_92_841_0 & ~i_8_92_1255_0 & ~i_8_92_1301_0 & ~i_8_92_1369_0 & ~i_8_92_1620_0 & ~i_8_92_1733_0 & i_8_92_1748_0 & ~i_8_92_1900_0))) | (~i_8_92_695_0 & ~i_8_92_838_0 & ~i_8_92_1370_0 & ~i_8_92_1620_0 & ~i_8_92_1628_0 & ~i_8_92_1854_0 & i_8_92_1945_0) | (i_8_92_1113_0 & ~i_8_92_1369_0 & i_8_92_1437_0 & ~i_8_92_2276_0))) | (~i_8_92_1370_0 & ((~i_8_92_1255_0 & ((i_8_92_484_0 & ~i_8_92_841_0 & ~i_8_92_843_0 & ~i_8_92_1826_0) | (~i_8_92_484_0 & ~i_8_92_523_0 & ~i_8_92_1027_0 & i_8_92_1355_0 & i_8_92_1439_0 & ~i_8_92_1455_0 & ~i_8_92_1634_0 & i_8_92_1861_0))) | (i_8_92_556_0 & i_8_92_827_0 & ~i_8_92_1369_0 & ~i_8_92_1535_0))) | (~i_8_92_1620_0 & ((~i_8_92_1027_0 & ((~i_8_92_880_0 & i_8_92_1110_0 & ~i_8_92_1369_0 & ~i_8_92_1438_0 & ~i_8_92_1455_0 & ~i_8_92_1861_0) | (i_8_92_699_0 & i_8_92_1437_0 & i_8_92_1753_0 & ~i_8_92_1825_0 & i_8_92_1888_0))) | (i_8_92_370_0 & ~i_8_92_698_0 & i_8_92_1263_0 & ~i_8_92_1854_0))));
endmodule



// Benchmark "kernel_8_93" written by ABC on Sun Jul 19 10:04:37 2020

module kernel_8_93 ( 
    i_8_93_22_0, i_8_93_23_0, i_8_93_31_0, i_8_93_70_0, i_8_93_140_0,
    i_8_93_188_0, i_8_93_202_0, i_8_93_223_0, i_8_93_224_0, i_8_93_275_0,
    i_8_93_292_0, i_8_93_293_0, i_8_93_301_0, i_8_93_345_0, i_8_93_346_0,
    i_8_93_364_0, i_8_93_374_0, i_8_93_377_0, i_8_93_379_0, i_8_93_390_0,
    i_8_93_451_0, i_8_93_484_0, i_8_93_507_0, i_8_93_555_0, i_8_93_556_0,
    i_8_93_577_0, i_8_93_589_0, i_8_93_599_0, i_8_93_634_0, i_8_93_636_0,
    i_8_93_672_0, i_8_93_711_0, i_8_93_715_0, i_8_93_716_0, i_8_93_772_0,
    i_8_93_786_0, i_8_93_826_0, i_8_93_839_0, i_8_93_840_0, i_8_93_872_0,
    i_8_93_881_0, i_8_93_985_0, i_8_93_994_0, i_8_93_1029_0, i_8_93_1119_0,
    i_8_93_1120_0, i_8_93_1121_0, i_8_93_1124_0, i_8_93_1186_0,
    i_8_93_1192_0, i_8_93_1219_0, i_8_93_1220_0, i_8_93_1236_0,
    i_8_93_1256_0, i_8_93_1271_0, i_8_93_1274_0, i_8_93_1283_0,
    i_8_93_1299_0, i_8_93_1305_0, i_8_93_1306_0, i_8_93_1314_0,
    i_8_93_1328_0, i_8_93_1329_0, i_8_93_1331_0, i_8_93_1410_0,
    i_8_93_1467_0, i_8_93_1470_0, i_8_93_1478_0, i_8_93_1497_0,
    i_8_93_1506_0, i_8_93_1507_0, i_8_93_1508_0, i_8_93_1542_0,
    i_8_93_1573_0, i_8_93_1615_0, i_8_93_1653_0, i_8_93_1654_0,
    i_8_93_1669_0, i_8_93_1742_0, i_8_93_1752_0, i_8_93_1763_0,
    i_8_93_1788_0, i_8_93_1789_0, i_8_93_1790_0, i_8_93_1832_0,
    i_8_93_1857_0, i_8_93_1858_0, i_8_93_1859_0, i_8_93_1885_0,
    i_8_93_1985_0, i_8_93_2047_0, i_8_93_2137_0, i_8_93_2153_0,
    i_8_93_2214_0, i_8_93_2215_0, i_8_93_2216_0, i_8_93_2226_0,
    i_8_93_2249_0, i_8_93_2261_0, i_8_93_2273_0,
    o_8_93_0_0  );
  input  i_8_93_22_0, i_8_93_23_0, i_8_93_31_0, i_8_93_70_0,
    i_8_93_140_0, i_8_93_188_0, i_8_93_202_0, i_8_93_223_0, i_8_93_224_0,
    i_8_93_275_0, i_8_93_292_0, i_8_93_293_0, i_8_93_301_0, i_8_93_345_0,
    i_8_93_346_0, i_8_93_364_0, i_8_93_374_0, i_8_93_377_0, i_8_93_379_0,
    i_8_93_390_0, i_8_93_451_0, i_8_93_484_0, i_8_93_507_0, i_8_93_555_0,
    i_8_93_556_0, i_8_93_577_0, i_8_93_589_0, i_8_93_599_0, i_8_93_634_0,
    i_8_93_636_0, i_8_93_672_0, i_8_93_711_0, i_8_93_715_0, i_8_93_716_0,
    i_8_93_772_0, i_8_93_786_0, i_8_93_826_0, i_8_93_839_0, i_8_93_840_0,
    i_8_93_872_0, i_8_93_881_0, i_8_93_985_0, i_8_93_994_0, i_8_93_1029_0,
    i_8_93_1119_0, i_8_93_1120_0, i_8_93_1121_0, i_8_93_1124_0,
    i_8_93_1186_0, i_8_93_1192_0, i_8_93_1219_0, i_8_93_1220_0,
    i_8_93_1236_0, i_8_93_1256_0, i_8_93_1271_0, i_8_93_1274_0,
    i_8_93_1283_0, i_8_93_1299_0, i_8_93_1305_0, i_8_93_1306_0,
    i_8_93_1314_0, i_8_93_1328_0, i_8_93_1329_0, i_8_93_1331_0,
    i_8_93_1410_0, i_8_93_1467_0, i_8_93_1470_0, i_8_93_1478_0,
    i_8_93_1497_0, i_8_93_1506_0, i_8_93_1507_0, i_8_93_1508_0,
    i_8_93_1542_0, i_8_93_1573_0, i_8_93_1615_0, i_8_93_1653_0,
    i_8_93_1654_0, i_8_93_1669_0, i_8_93_1742_0, i_8_93_1752_0,
    i_8_93_1763_0, i_8_93_1788_0, i_8_93_1789_0, i_8_93_1790_0,
    i_8_93_1832_0, i_8_93_1857_0, i_8_93_1858_0, i_8_93_1859_0,
    i_8_93_1885_0, i_8_93_1985_0, i_8_93_2047_0, i_8_93_2137_0,
    i_8_93_2153_0, i_8_93_2214_0, i_8_93_2215_0, i_8_93_2216_0,
    i_8_93_2226_0, i_8_93_2249_0, i_8_93_2261_0, i_8_93_2273_0;
  output o_8_93_0_0;
  assign o_8_93_0_0 = ~((~i_8_93_1314_0 & ((~i_8_93_22_0 & ((~i_8_93_1192_0 & ~i_8_93_1885_0 & i_8_93_2137_0) | (~i_8_93_188_0 & ~i_8_93_292_0 & ~i_8_93_507_0 & ~i_8_93_672_0 & ~i_8_93_1274_0 & ~i_8_93_1763_0 & ~i_8_93_2216_0))) | (~i_8_93_484_0 & ~i_8_93_786_0 & ~i_8_93_1029_0 & ~i_8_93_1271_0 & ~i_8_93_1573_0 & ~i_8_93_2216_0) | (~i_8_93_377_0 & ~i_8_93_826_0 & ~i_8_93_1120_0 & ~i_8_93_1331_0 & ~i_8_93_1615_0 & ~i_8_93_1752_0 & ~i_8_93_1788_0 & ~i_8_93_2153_0))) | (~i_8_93_1119_0 & ((~i_8_93_223_0 & ((~i_8_93_188_0 & ~i_8_93_292_0 & ~i_8_93_881_0 & ~i_8_93_1506_0) | (~i_8_93_1186_0 & ~i_8_93_1274_0 & ~i_8_93_1542_0 & ~i_8_93_1742_0))) | (~i_8_93_224_0 & ~i_8_93_772_0 & ~i_8_93_872_0 & ~i_8_93_1121_0 & ~i_8_93_1124_0 & ~i_8_93_1467_0 & ~i_8_93_1573_0))) | (~i_8_93_188_0 & ((i_8_93_634_0 & ~i_8_93_1331_0 & ~i_8_93_1467_0) | (~i_8_93_293_0 & ~i_8_93_484_0 & ~i_8_93_786_0 & ~i_8_93_1120_0 & ~i_8_93_1507_0))) | (~i_8_93_301_0 & ((~i_8_93_484_0 & ~i_8_93_1271_0 & ~i_8_93_1331_0 & ~i_8_93_1470_0) | (~i_8_93_556_0 & ~i_8_93_589_0 & ~i_8_93_716_0 & ~i_8_93_994_0 & ~i_8_93_2261_0))) | (~i_8_93_374_0 & ((~i_8_93_377_0 & i_8_93_556_0 & ~i_8_93_1271_0 & ~i_8_93_1542_0 & ~i_8_93_1654_0) | (~i_8_93_672_0 & ~i_8_93_1478_0 & ~i_8_93_1507_0 & ~i_8_93_1788_0))) | (~i_8_93_1124_0 & ((~i_8_93_70_0 & ~i_8_93_1274_0 & ~i_8_93_1283_0 & ~i_8_93_1305_0 & ~i_8_93_1328_0 & ~i_8_93_1329_0 & ~i_8_93_1573_0 & ~i_8_93_1763_0 & ~i_8_93_1832_0) | (~i_8_93_292_0 & i_8_93_1859_0))) | (~i_8_93_293_0 & i_8_93_556_0 & i_8_93_634_0 & ~i_8_93_1832_0) | (i_8_93_301_0 & i_8_93_451_0 & ~i_8_93_484_0 & ~i_8_93_994_0 & ~i_8_93_1305_0) | (~i_8_93_716_0 & ~i_8_93_1121_0 & ~i_8_93_1274_0 & ~i_8_93_1506_0 & ~i_8_93_2214_0) | (~i_8_93_599_0 & ~i_8_93_715_0 & ~i_8_93_1742_0 & ~i_8_93_1790_0 & ~i_8_93_2215_0) | (i_8_93_1985_0 & i_8_93_2249_0));
endmodule



// Benchmark "kernel_8_94" written by ABC on Sun Jul 19 10:04:38 2020

module kernel_8_94 ( 
    i_8_94_13_0, i_8_94_43_0, i_8_94_115_0, i_8_94_139_0, i_8_94_143_0,
    i_8_94_152_0, i_8_94_153_0, i_8_94_201_0, i_8_94_226_0, i_8_94_233_0,
    i_8_94_356_0, i_8_94_382_0, i_8_94_392_0, i_8_94_455_0, i_8_94_458_0,
    i_8_94_522_0, i_8_94_526_0, i_8_94_572_0, i_8_94_591_0, i_8_94_592_0,
    i_8_94_595_0, i_8_94_596_0, i_8_94_635_0, i_8_94_652_0, i_8_94_656_0,
    i_8_94_659_0, i_8_94_661_0, i_8_94_671_0, i_8_94_688_0, i_8_94_706_0,
    i_8_94_733_0, i_8_94_759_0, i_8_94_760_0, i_8_94_838_0, i_8_94_860_0,
    i_8_94_923_0, i_8_94_959_0, i_8_94_1013_0, i_8_94_1032_0,
    i_8_94_1115_0, i_8_94_1156_0, i_8_94_1174_0, i_8_94_1188_0,
    i_8_94_1229_0, i_8_94_1232_0, i_8_94_1267_0, i_8_94_1268_0,
    i_8_94_1271_0, i_8_94_1297_0, i_8_94_1300_0, i_8_94_1305_0,
    i_8_94_1306_0, i_8_94_1307_0, i_8_94_1309_0, i_8_94_1331_0,
    i_8_94_1385_0, i_8_94_1390_0, i_8_94_1400_0, i_8_94_1438_0,
    i_8_94_1469_0, i_8_94_1470_0, i_8_94_1471_0, i_8_94_1478_0,
    i_8_94_1498_0, i_8_94_1531_0, i_8_94_1534_0, i_8_94_1535_0,
    i_8_94_1544_0, i_8_94_1645_0, i_8_94_1651_0, i_8_94_1679_0,
    i_8_94_1697_0, i_8_94_1706_0, i_8_94_1778_0, i_8_94_1798_0,
    i_8_94_1806_0, i_8_94_1807_0, i_8_94_1822_0, i_8_94_1823_0,
    i_8_94_1826_0, i_8_94_1868_0, i_8_94_1874_0, i_8_94_1883_0,
    i_8_94_1884_0, i_8_94_1886_0, i_8_94_1916_0, i_8_94_1960_0,
    i_8_94_1975_0, i_8_94_1992_0, i_8_94_2030_0, i_8_94_2041_0,
    i_8_94_2066_0, i_8_94_2120_0, i_8_94_2155_0, i_8_94_2173_0,
    i_8_94_2216_0, i_8_94_2230_0, i_8_94_2243_0, i_8_94_2248_0,
    i_8_94_2296_0,
    o_8_94_0_0  );
  input  i_8_94_13_0, i_8_94_43_0, i_8_94_115_0, i_8_94_139_0,
    i_8_94_143_0, i_8_94_152_0, i_8_94_153_0, i_8_94_201_0, i_8_94_226_0,
    i_8_94_233_0, i_8_94_356_0, i_8_94_382_0, i_8_94_392_0, i_8_94_455_0,
    i_8_94_458_0, i_8_94_522_0, i_8_94_526_0, i_8_94_572_0, i_8_94_591_0,
    i_8_94_592_0, i_8_94_595_0, i_8_94_596_0, i_8_94_635_0, i_8_94_652_0,
    i_8_94_656_0, i_8_94_659_0, i_8_94_661_0, i_8_94_671_0, i_8_94_688_0,
    i_8_94_706_0, i_8_94_733_0, i_8_94_759_0, i_8_94_760_0, i_8_94_838_0,
    i_8_94_860_0, i_8_94_923_0, i_8_94_959_0, i_8_94_1013_0, i_8_94_1032_0,
    i_8_94_1115_0, i_8_94_1156_0, i_8_94_1174_0, i_8_94_1188_0,
    i_8_94_1229_0, i_8_94_1232_0, i_8_94_1267_0, i_8_94_1268_0,
    i_8_94_1271_0, i_8_94_1297_0, i_8_94_1300_0, i_8_94_1305_0,
    i_8_94_1306_0, i_8_94_1307_0, i_8_94_1309_0, i_8_94_1331_0,
    i_8_94_1385_0, i_8_94_1390_0, i_8_94_1400_0, i_8_94_1438_0,
    i_8_94_1469_0, i_8_94_1470_0, i_8_94_1471_0, i_8_94_1478_0,
    i_8_94_1498_0, i_8_94_1531_0, i_8_94_1534_0, i_8_94_1535_0,
    i_8_94_1544_0, i_8_94_1645_0, i_8_94_1651_0, i_8_94_1679_0,
    i_8_94_1697_0, i_8_94_1706_0, i_8_94_1778_0, i_8_94_1798_0,
    i_8_94_1806_0, i_8_94_1807_0, i_8_94_1822_0, i_8_94_1823_0,
    i_8_94_1826_0, i_8_94_1868_0, i_8_94_1874_0, i_8_94_1883_0,
    i_8_94_1884_0, i_8_94_1886_0, i_8_94_1916_0, i_8_94_1960_0,
    i_8_94_1975_0, i_8_94_1992_0, i_8_94_2030_0, i_8_94_2041_0,
    i_8_94_2066_0, i_8_94_2120_0, i_8_94_2155_0, i_8_94_2173_0,
    i_8_94_2216_0, i_8_94_2230_0, i_8_94_2243_0, i_8_94_2248_0,
    i_8_94_2296_0;
  output o_8_94_0_0;
  assign o_8_94_0_0 = 0;
endmodule



// Benchmark "kernel_8_95" written by ABC on Sun Jul 19 10:04:39 2020

module kernel_8_95 ( 
    i_8_95_3_0, i_8_95_7_0, i_8_95_22_0, i_8_95_124_0, i_8_95_170_0,
    i_8_95_200_0, i_8_95_250_0, i_8_95_287_0, i_8_95_292_0, i_8_95_293_0,
    i_8_95_328_0, i_8_95_329_0, i_8_95_330_0, i_8_95_366_0, i_8_95_383_0,
    i_8_95_385_0, i_8_95_440_0, i_8_95_456_0, i_8_95_493_0, i_8_95_529_0,
    i_8_95_554_0, i_8_95_584_0, i_8_95_626_0, i_8_95_635_0, i_8_95_642_0,
    i_8_95_673_0, i_8_95_674_0, i_8_95_680_0, i_8_95_695_0, i_8_95_700_0,
    i_8_95_701_0, i_8_95_703_0, i_8_95_704_0, i_8_95_763_0, i_8_95_809_0,
    i_8_95_827_0, i_8_95_833_0, i_8_95_836_0, i_8_95_844_0, i_8_95_852_0,
    i_8_95_854_0, i_8_95_958_0, i_8_95_968_0, i_8_95_971_0, i_8_95_986_0,
    i_8_95_989_0, i_8_95_1154_0, i_8_95_1194_0, i_8_95_1227_0,
    i_8_95_1258_0, i_8_95_1259_0, i_8_95_1267_0, i_8_95_1270_0,
    i_8_95_1286_0, i_8_95_1299_0, i_8_95_1323_0, i_8_95_1350_0,
    i_8_95_1358_0, i_8_95_1436_0, i_8_95_1442_0, i_8_95_1468_0,
    i_8_95_1489_0, i_8_95_1493_0, i_8_95_1520_0, i_8_95_1538_0,
    i_8_95_1547_0, i_8_95_1574_0, i_8_95_1585_0, i_8_95_1588_0,
    i_8_95_1591_0, i_8_95_1650_0, i_8_95_1652_0, i_8_95_1675_0,
    i_8_95_1705_0, i_8_95_1724_0, i_8_95_1750_0, i_8_95_1769_0,
    i_8_95_1777_0, i_8_95_1781_0, i_8_95_1817_0, i_8_95_1820_0,
    i_8_95_1824_0, i_8_95_1834_0, i_8_95_1843_0, i_8_95_1860_0,
    i_8_95_1885_0, i_8_95_1892_0, i_8_95_1896_0, i_8_95_2032_0,
    i_8_95_2041_0, i_8_95_2042_0, i_8_95_2089_0, i_8_95_2146_0,
    i_8_95_2149_0, i_8_95_2155_0, i_8_95_2187_0, i_8_95_2191_0,
    i_8_95_2192_0, i_8_95_2244_0, i_8_95_2275_0,
    o_8_95_0_0  );
  input  i_8_95_3_0, i_8_95_7_0, i_8_95_22_0, i_8_95_124_0, i_8_95_170_0,
    i_8_95_200_0, i_8_95_250_0, i_8_95_287_0, i_8_95_292_0, i_8_95_293_0,
    i_8_95_328_0, i_8_95_329_0, i_8_95_330_0, i_8_95_366_0, i_8_95_383_0,
    i_8_95_385_0, i_8_95_440_0, i_8_95_456_0, i_8_95_493_0, i_8_95_529_0,
    i_8_95_554_0, i_8_95_584_0, i_8_95_626_0, i_8_95_635_0, i_8_95_642_0,
    i_8_95_673_0, i_8_95_674_0, i_8_95_680_0, i_8_95_695_0, i_8_95_700_0,
    i_8_95_701_0, i_8_95_703_0, i_8_95_704_0, i_8_95_763_0, i_8_95_809_0,
    i_8_95_827_0, i_8_95_833_0, i_8_95_836_0, i_8_95_844_0, i_8_95_852_0,
    i_8_95_854_0, i_8_95_958_0, i_8_95_968_0, i_8_95_971_0, i_8_95_986_0,
    i_8_95_989_0, i_8_95_1154_0, i_8_95_1194_0, i_8_95_1227_0,
    i_8_95_1258_0, i_8_95_1259_0, i_8_95_1267_0, i_8_95_1270_0,
    i_8_95_1286_0, i_8_95_1299_0, i_8_95_1323_0, i_8_95_1350_0,
    i_8_95_1358_0, i_8_95_1436_0, i_8_95_1442_0, i_8_95_1468_0,
    i_8_95_1489_0, i_8_95_1493_0, i_8_95_1520_0, i_8_95_1538_0,
    i_8_95_1547_0, i_8_95_1574_0, i_8_95_1585_0, i_8_95_1588_0,
    i_8_95_1591_0, i_8_95_1650_0, i_8_95_1652_0, i_8_95_1675_0,
    i_8_95_1705_0, i_8_95_1724_0, i_8_95_1750_0, i_8_95_1769_0,
    i_8_95_1777_0, i_8_95_1781_0, i_8_95_1817_0, i_8_95_1820_0,
    i_8_95_1824_0, i_8_95_1834_0, i_8_95_1843_0, i_8_95_1860_0,
    i_8_95_1885_0, i_8_95_1892_0, i_8_95_1896_0, i_8_95_2032_0,
    i_8_95_2041_0, i_8_95_2042_0, i_8_95_2089_0, i_8_95_2146_0,
    i_8_95_2149_0, i_8_95_2155_0, i_8_95_2187_0, i_8_95_2191_0,
    i_8_95_2192_0, i_8_95_2244_0, i_8_95_2275_0;
  output o_8_95_0_0;
  assign o_8_95_0_0 = ~((~i_8_95_22_0 & ((~i_8_95_809_0 & ~i_8_95_1270_0 & i_8_95_1358_0 & ~i_8_95_1520_0 & ~i_8_95_1574_0 & ~i_8_95_1591_0 & ~i_8_95_1834_0) | (~i_8_95_385_0 & ~i_8_95_584_0 & ~i_8_95_1259_0 & ~i_8_95_2042_0))) | (~i_8_95_293_0 & ((~i_8_95_170_0 & ~i_8_95_440_0 & ~i_8_95_680_0 & ~i_8_95_1259_0) | (~i_8_95_366_0 & ~i_8_95_701_0 & ~i_8_95_2041_0 & ~i_8_95_2146_0))) | (~i_8_95_170_0 & ((~i_8_95_836_0 & ~i_8_95_1258_0 & ~i_8_95_1259_0 & ~i_8_95_1270_0 & ~i_8_95_1323_0 & ~i_8_95_1442_0 & ~i_8_95_1591_0) | (i_8_95_968_0 & ~i_8_95_1267_0 & i_8_95_1817_0))) | (~i_8_95_2032_0 & ((~i_8_95_440_0 & ~i_8_95_2192_0 & ((~i_8_95_680_0 & ~i_8_95_971_0 & ~i_8_95_1436_0 & ~i_8_95_1820_0) | (~i_8_95_827_0 & ~i_8_95_1781_0 & ~i_8_95_1824_0))) | (~i_8_95_330_0 & i_8_95_635_0 & ~i_8_95_1258_0 & ~i_8_95_1442_0 & ~i_8_95_1574_0 & ~i_8_95_2155_0 & ~i_8_95_2191_0))) | (~i_8_95_809_0 & ((~i_8_95_200_0 & ~i_8_95_383_0 & ~i_8_95_844_0 & i_8_95_2149_0) | (~i_8_95_836_0 & ~i_8_95_1358_0 & ~i_8_95_2149_0))) | (~i_8_95_1817_0 & ((~i_8_95_329_0 & ~i_8_95_827_0) | (~i_8_95_7_0 & i_8_95_329_0 & ~i_8_95_833_0 & ~i_8_95_1259_0 & ~i_8_95_2042_0))));
endmodule



// Benchmark "kernel_8_96" written by ABC on Sun Jul 19 10:04:40 2020

module kernel_8_96 ( 
    i_8_96_23_0, i_8_96_35_0, i_8_96_53_0, i_8_96_57_0, i_8_96_62_0,
    i_8_96_74_0, i_8_96_98_0, i_8_96_141_0, i_8_96_158_0, i_8_96_187_0,
    i_8_96_223_0, i_8_96_260_0, i_8_96_304_0, i_8_96_305_0, i_8_96_311_0,
    i_8_96_348_0, i_8_96_349_0, i_8_96_421_0, i_8_96_422_0, i_8_96_524_0,
    i_8_96_527_0, i_8_96_530_0, i_8_96_590_0, i_8_96_602_0, i_8_96_610_0,
    i_8_96_625_0, i_8_96_631_0, i_8_96_632_0, i_8_96_634_0, i_8_96_635_0,
    i_8_96_659_0, i_8_96_662_0, i_8_96_663_0, i_8_96_690_0, i_8_96_691_0,
    i_8_96_715_0, i_8_96_770_0, i_8_96_789_0, i_8_96_814_0, i_8_96_817_0,
    i_8_96_839_0, i_8_96_853_0, i_8_96_854_0, i_8_96_876_0, i_8_96_880_0,
    i_8_96_964_0, i_8_96_994_0, i_8_96_1016_0, i_8_96_1018_0,
    i_8_96_1032_0, i_8_96_1034_0, i_8_96_1052_0, i_8_96_1076_0,
    i_8_96_1129_0, i_8_96_1193_0, i_8_96_1264_0, i_8_96_1277_0,
    i_8_96_1299_0, i_8_96_1305_0, i_8_96_1327_0, i_8_96_1328_0,
    i_8_96_1331_0, i_8_96_1344_0, i_8_96_1346_0, i_8_96_1397_0,
    i_8_96_1411_0, i_8_96_1434_0, i_8_96_1438_0, i_8_96_1506_0,
    i_8_96_1507_0, i_8_96_1545_0, i_8_96_1546_0, i_8_96_1565_0,
    i_8_96_1574_0, i_8_96_1603_0, i_8_96_1624_0, i_8_96_1648_0,
    i_8_96_1654_0, i_8_96_1720_0, i_8_96_1723_0, i_8_96_1736_0,
    i_8_96_1742_0, i_8_96_1806_0, i_8_96_1808_0, i_8_96_1844_0,
    i_8_96_1888_0, i_8_96_1905_0, i_8_96_1906_0, i_8_96_1919_0,
    i_8_96_2017_0, i_8_96_2032_0, i_8_96_2072_0, i_8_96_2093_0,
    i_8_96_2134_0, i_8_96_2157_0, i_8_96_2165_0, i_8_96_2216_0,
    i_8_96_2239_0, i_8_96_2291_0, i_8_96_2292_0,
    o_8_96_0_0  );
  input  i_8_96_23_0, i_8_96_35_0, i_8_96_53_0, i_8_96_57_0, i_8_96_62_0,
    i_8_96_74_0, i_8_96_98_0, i_8_96_141_0, i_8_96_158_0, i_8_96_187_0,
    i_8_96_223_0, i_8_96_260_0, i_8_96_304_0, i_8_96_305_0, i_8_96_311_0,
    i_8_96_348_0, i_8_96_349_0, i_8_96_421_0, i_8_96_422_0, i_8_96_524_0,
    i_8_96_527_0, i_8_96_530_0, i_8_96_590_0, i_8_96_602_0, i_8_96_610_0,
    i_8_96_625_0, i_8_96_631_0, i_8_96_632_0, i_8_96_634_0, i_8_96_635_0,
    i_8_96_659_0, i_8_96_662_0, i_8_96_663_0, i_8_96_690_0, i_8_96_691_0,
    i_8_96_715_0, i_8_96_770_0, i_8_96_789_0, i_8_96_814_0, i_8_96_817_0,
    i_8_96_839_0, i_8_96_853_0, i_8_96_854_0, i_8_96_876_0, i_8_96_880_0,
    i_8_96_964_0, i_8_96_994_0, i_8_96_1016_0, i_8_96_1018_0,
    i_8_96_1032_0, i_8_96_1034_0, i_8_96_1052_0, i_8_96_1076_0,
    i_8_96_1129_0, i_8_96_1193_0, i_8_96_1264_0, i_8_96_1277_0,
    i_8_96_1299_0, i_8_96_1305_0, i_8_96_1327_0, i_8_96_1328_0,
    i_8_96_1331_0, i_8_96_1344_0, i_8_96_1346_0, i_8_96_1397_0,
    i_8_96_1411_0, i_8_96_1434_0, i_8_96_1438_0, i_8_96_1506_0,
    i_8_96_1507_0, i_8_96_1545_0, i_8_96_1546_0, i_8_96_1565_0,
    i_8_96_1574_0, i_8_96_1603_0, i_8_96_1624_0, i_8_96_1648_0,
    i_8_96_1654_0, i_8_96_1720_0, i_8_96_1723_0, i_8_96_1736_0,
    i_8_96_1742_0, i_8_96_1806_0, i_8_96_1808_0, i_8_96_1844_0,
    i_8_96_1888_0, i_8_96_1905_0, i_8_96_1906_0, i_8_96_1919_0,
    i_8_96_2017_0, i_8_96_2032_0, i_8_96_2072_0, i_8_96_2093_0,
    i_8_96_2134_0, i_8_96_2157_0, i_8_96_2165_0, i_8_96_2216_0,
    i_8_96_2239_0, i_8_96_2291_0, i_8_96_2292_0;
  output o_8_96_0_0;
  assign o_8_96_0_0 = 0;
endmodule



// Benchmark "kernel_8_97" written by ABC on Sun Jul 19 10:04:41 2020

module kernel_8_97 ( 
    i_8_97_60_0, i_8_97_61_0, i_8_97_69_0, i_8_97_70_0, i_8_97_115_0,
    i_8_97_132_0, i_8_97_171_0, i_8_97_186_0, i_8_97_189_0, i_8_97_190_0,
    i_8_97_213_0, i_8_97_214_0, i_8_97_295_0, i_8_97_296_0, i_8_97_303_0,
    i_8_97_304_0, i_8_97_339_0, i_8_97_378_0, i_8_97_382_0, i_8_97_420_0,
    i_8_97_456_0, i_8_97_469_0, i_8_97_492_0, i_8_97_582_0, i_8_97_591_0,
    i_8_97_606_0, i_8_97_619_0, i_8_97_633_0, i_8_97_637_0, i_8_97_658_0,
    i_8_97_665_0, i_8_97_753_0, i_8_97_898_0, i_8_97_924_0, i_8_97_1015_0,
    i_8_97_1073_0, i_8_97_1102_0, i_8_97_1105_0, i_8_97_1131_0,
    i_8_97_1141_0, i_8_97_1156_0, i_8_97_1176_0, i_8_97_1263_0,
    i_8_97_1267_0, i_8_97_1284_0, i_8_97_1286_0, i_8_97_1288_0,
    i_8_97_1304_0, i_8_97_1308_0, i_8_97_1332_0, i_8_97_1353_0,
    i_8_97_1356_0, i_8_97_1383_0, i_8_97_1402_0, i_8_97_1410_0,
    i_8_97_1482_0, i_8_97_1484_0, i_8_97_1528_0, i_8_97_1555_0,
    i_8_97_1591_0, i_8_97_1645_0, i_8_97_1671_0, i_8_97_1672_0,
    i_8_97_1673_0, i_8_97_1677_0, i_8_97_1681_0, i_8_97_1689_0,
    i_8_97_1707_0, i_8_97_1713_0, i_8_97_1714_0, i_8_97_1731_0,
    i_8_97_1732_0, i_8_97_1734_0, i_8_97_1746_0, i_8_97_1754_0,
    i_8_97_1762_0, i_8_97_1773_0, i_8_97_1779_0, i_8_97_1821_0,
    i_8_97_1843_0, i_8_97_1857_0, i_8_97_1860_0, i_8_97_1887_0,
    i_8_97_1888_0, i_8_97_1895_0, i_8_97_1942_0, i_8_97_1966_0,
    i_8_97_1986_0, i_8_97_1996_0, i_8_97_1997_0, i_8_97_2004_0,
    i_8_97_2014_0, i_8_97_2076_0, i_8_97_2149_0, i_8_97_2151_0,
    i_8_97_2173_0, i_8_97_2242_0, i_8_97_2250_0, i_8_97_2275_0,
    i_8_97_2292_0,
    o_8_97_0_0  );
  input  i_8_97_60_0, i_8_97_61_0, i_8_97_69_0, i_8_97_70_0,
    i_8_97_115_0, i_8_97_132_0, i_8_97_171_0, i_8_97_186_0, i_8_97_189_0,
    i_8_97_190_0, i_8_97_213_0, i_8_97_214_0, i_8_97_295_0, i_8_97_296_0,
    i_8_97_303_0, i_8_97_304_0, i_8_97_339_0, i_8_97_378_0, i_8_97_382_0,
    i_8_97_420_0, i_8_97_456_0, i_8_97_469_0, i_8_97_492_0, i_8_97_582_0,
    i_8_97_591_0, i_8_97_606_0, i_8_97_619_0, i_8_97_633_0, i_8_97_637_0,
    i_8_97_658_0, i_8_97_665_0, i_8_97_753_0, i_8_97_898_0, i_8_97_924_0,
    i_8_97_1015_0, i_8_97_1073_0, i_8_97_1102_0, i_8_97_1105_0,
    i_8_97_1131_0, i_8_97_1141_0, i_8_97_1156_0, i_8_97_1176_0,
    i_8_97_1263_0, i_8_97_1267_0, i_8_97_1284_0, i_8_97_1286_0,
    i_8_97_1288_0, i_8_97_1304_0, i_8_97_1308_0, i_8_97_1332_0,
    i_8_97_1353_0, i_8_97_1356_0, i_8_97_1383_0, i_8_97_1402_0,
    i_8_97_1410_0, i_8_97_1482_0, i_8_97_1484_0, i_8_97_1528_0,
    i_8_97_1555_0, i_8_97_1591_0, i_8_97_1645_0, i_8_97_1671_0,
    i_8_97_1672_0, i_8_97_1673_0, i_8_97_1677_0, i_8_97_1681_0,
    i_8_97_1689_0, i_8_97_1707_0, i_8_97_1713_0, i_8_97_1714_0,
    i_8_97_1731_0, i_8_97_1732_0, i_8_97_1734_0, i_8_97_1746_0,
    i_8_97_1754_0, i_8_97_1762_0, i_8_97_1773_0, i_8_97_1779_0,
    i_8_97_1821_0, i_8_97_1843_0, i_8_97_1857_0, i_8_97_1860_0,
    i_8_97_1887_0, i_8_97_1888_0, i_8_97_1895_0, i_8_97_1942_0,
    i_8_97_1966_0, i_8_97_1986_0, i_8_97_1996_0, i_8_97_1997_0,
    i_8_97_2004_0, i_8_97_2014_0, i_8_97_2076_0, i_8_97_2149_0,
    i_8_97_2151_0, i_8_97_2173_0, i_8_97_2242_0, i_8_97_2250_0,
    i_8_97_2275_0, i_8_97_2292_0;
  output o_8_97_0_0;
  assign o_8_97_0_0 = ~((~i_8_97_1528_0 & ((~i_8_97_60_0 & ((~i_8_97_115_0 & ~i_8_97_637_0 & ~i_8_97_1105_0 & ~i_8_97_1308_0 & ~i_8_97_1383_0 & ~i_8_97_1410_0 & ~i_8_97_1484_0 & ~i_8_97_1707_0 & i_8_97_1860_0) | (~i_8_97_132_0 & ~i_8_97_214_0 & ~i_8_97_606_0 & ~i_8_97_1482_0 & i_8_97_1966_0 & ~i_8_97_2242_0))) | (~i_8_97_189_0 & ((~i_8_97_132_0 & ~i_8_97_213_0 & i_8_97_606_0 & i_8_97_1966_0) | (~i_8_97_186_0 & ~i_8_97_214_0 & ~i_8_97_898_0 & ~i_8_97_1105_0 & ~i_8_97_1482_0 & ~i_8_97_1671_0 & ~i_8_97_1689_0 & ~i_8_97_1887_0 & ~i_8_97_1942_0 & ~i_8_97_2014_0))) | (~i_8_97_69_0 & ~i_8_97_190_0 & ~i_8_97_382_0 & ~i_8_97_665_0 & ~i_8_97_1073_0 & ~i_8_97_1671_0 & ~i_8_97_1681_0 & ~i_8_97_1731_0 & ~i_8_97_1857_0 & ~i_8_97_2004_0 & ~i_8_97_2076_0 & ~i_8_97_2242_0) | (i_8_97_1267_0 & ~i_8_97_1286_0 & ~i_8_97_1308_0 & i_8_97_1353_0 & ~i_8_97_1673_0 & ~i_8_97_2014_0 & i_8_97_2149_0 & ~i_8_97_2292_0))) | (i_8_97_115_0 & ((~i_8_97_69_0 & ~i_8_97_189_0 & ~i_8_97_214_0 & ~i_8_97_420_0 & ~i_8_97_1383_0 & ~i_8_97_1671_0 & ~i_8_97_1672_0 & ~i_8_97_1673_0 & ~i_8_97_1754_0) | (~i_8_97_186_0 & ~i_8_97_1102_0 & ~i_8_97_1105_0 & ~i_8_97_1176_0 & ~i_8_97_1402_0 & ~i_8_97_1410_0 & ~i_8_97_1591_0 & ~i_8_97_1689_0 & ~i_8_97_1843_0 & ~i_8_97_1997_0 & ~i_8_97_2014_0 & ~i_8_97_2292_0))) | (~i_8_97_69_0 & ((~i_8_97_132_0 & ~i_8_97_190_0 & ~i_8_97_469_0 & ~i_8_97_1105_0 & ~i_8_97_1672_0 & ~i_8_97_1707_0 & ~i_8_97_1843_0 & ~i_8_97_2004_0 & ~i_8_97_2014_0) | (~i_8_97_70_0 & ~i_8_97_214_0 & i_8_97_456_0 & ~i_8_97_1015_0 & ~i_8_97_1131_0 & ~i_8_97_1176_0 & ~i_8_97_2076_0 & ~i_8_97_2151_0))) | (~i_8_97_1887_0 & ((~i_8_97_171_0 & ((~i_8_97_115_0 & ~i_8_97_213_0 & ~i_8_97_924_0 & ~i_8_97_1482_0 & ~i_8_97_1484_0 & ~i_8_97_1714_0 & ~i_8_97_1731_0 & ~i_8_97_1888_0) | (~i_8_97_189_0 & ~i_8_97_214_0 & ~i_8_97_296_0 & ~i_8_97_753_0 & ~i_8_97_1015_0 & ~i_8_97_1156_0 & ~i_8_97_1677_0 & ~i_8_97_1681_0 & ~i_8_97_1689_0 & ~i_8_97_1762_0 & ~i_8_97_1860_0 & ~i_8_97_2076_0 & ~i_8_97_2250_0))) | (~i_8_97_378_0 & ((~i_8_97_214_0 & ~i_8_97_898_0 & ~i_8_97_924_0 & ~i_8_97_1176_0 & ~i_8_97_1482_0 & ~i_8_97_1484_0 & ~i_8_97_1645_0 & ~i_8_97_1673_0) | (~i_8_97_70_0 & ~i_8_97_456_0 & ~i_8_97_492_0 & ~i_8_97_1131_0 & ~i_8_97_1681_0 & ~i_8_97_1714_0 & ~i_8_97_1732_0 & ~i_8_97_1860_0 & ~i_8_97_1966_0 & ~i_8_97_2275_0))) | (~i_8_97_1707_0 & ((~i_8_97_1105_0 & i_8_97_1156_0 & ~i_8_97_1402_0 & ~i_8_97_2004_0) | (i_8_97_469_0 & ~i_8_97_1102_0 & ~i_8_97_1895_0 & i_8_97_1996_0 & ~i_8_97_2014_0 & i_8_97_2149_0))))) | (~i_8_97_70_0 & ((i_8_97_382_0 & i_8_97_658_0 & ~i_8_97_1304_0 & ~i_8_97_1402_0 & ~i_8_97_1888_0) | (~i_8_97_132_0 & ~i_8_97_213_0 & ~i_8_97_420_0 & ~i_8_97_582_0 & ~i_8_97_1645_0 & ~i_8_97_1673_0 & ~i_8_97_2275_0))) | (~i_8_97_213_0 & ~i_8_97_1673_0 & ((~i_8_97_924_0 & ~i_8_97_1015_0 & ~i_8_97_1141_0 & ~i_8_97_1482_0 & ~i_8_97_1555_0 & ~i_8_97_1713_0 & ~i_8_97_1779_0 & ~i_8_97_1942_0) | (~i_8_97_189_0 & ~i_8_97_214_0 & ~i_8_97_1105_0 & ~i_8_97_1383_0 & ~i_8_97_1410_0 & ~i_8_97_1672_0 & ~i_8_97_1689_0 & ~i_8_97_1707_0 & ~i_8_97_1857_0 & ~i_8_97_2151_0))) | (~i_8_97_753_0 & ((~i_8_97_214_0 & ~i_8_97_420_0 & i_8_97_637_0 & ~i_8_97_898_0 & ~i_8_97_1102_0 & i_8_97_1681_0 & ~i_8_97_2076_0) | (i_8_97_469_0 & ~i_8_97_665_0 & ~i_8_97_1383_0 & ~i_8_97_2014_0 & i_8_97_2149_0 & ~i_8_97_1843_0 & ~i_8_97_1997_0) | (i_8_97_304_0 & ~i_8_97_1308_0 & ~i_8_97_1888_0 & ~i_8_97_1942_0 & ~i_8_97_2004_0 & ~i_8_97_2151_0))) | (i_8_97_2014_0 & ~i_8_97_2173_0 & i_8_97_2242_0 & ~i_8_97_2275_0));
endmodule



// Benchmark "kernel_8_98" written by ABC on Sun Jul 19 10:04:42 2020

module kernel_8_98 ( 
    i_8_98_12_0, i_8_98_52_0, i_8_98_70_0, i_8_98_115_0, i_8_98_139_0,
    i_8_98_141_0, i_8_98_228_0, i_8_98_230_0, i_8_98_231_0, i_8_98_314_0,
    i_8_98_319_0, i_8_98_334_0, i_8_98_342_0, i_8_98_345_0, i_8_98_363_0,
    i_8_98_366_0, i_8_98_384_0, i_8_98_400_0, i_8_98_420_0, i_8_98_430_0,
    i_8_98_504_0, i_8_98_525_0, i_8_98_538_0, i_8_98_553_0, i_8_98_557_0,
    i_8_98_570_0, i_8_98_571_0, i_8_98_581_0, i_8_98_583_0, i_8_98_588_0,
    i_8_98_600_0, i_8_98_601_0, i_8_98_603_0, i_8_98_628_0, i_8_98_634_0,
    i_8_98_651_0, i_8_98_657_0, i_8_98_696_0, i_8_98_700_0, i_8_98_704_0,
    i_8_98_732_0, i_8_98_777_0, i_8_98_781_0, i_8_98_819_0, i_8_98_831_0,
    i_8_98_840_0, i_8_98_842_0, i_8_98_843_0, i_8_98_875_0, i_8_98_877_0,
    i_8_98_879_0, i_8_98_895_0, i_8_98_947_0, i_8_98_993_0, i_8_98_1003_0,
    i_8_98_1105_0, i_8_98_1109_0, i_8_98_1115_0, i_8_98_1124_0,
    i_8_98_1156_0, i_8_98_1267_0, i_8_98_1282_0, i_8_98_1284_0,
    i_8_98_1315_0, i_8_98_1317_0, i_8_98_1320_0, i_8_98_1347_0,
    i_8_98_1354_0, i_8_98_1358_0, i_8_98_1366_0, i_8_98_1423_0,
    i_8_98_1426_0, i_8_98_1453_0, i_8_98_1462_0, i_8_98_1490_0,
    i_8_98_1509_0, i_8_98_1519_0, i_8_98_1524_0, i_8_98_1551_0,
    i_8_98_1633_0, i_8_98_1635_0, i_8_98_1680_0, i_8_98_1686_0,
    i_8_98_1690_0, i_8_98_1695_0, i_8_98_1699_0, i_8_98_1700_0,
    i_8_98_1703_0, i_8_98_1723_0, i_8_98_1770_0, i_8_98_1780_0,
    i_8_98_1884_0, i_8_98_1911_0, i_8_98_1956_0, i_8_98_1995_0,
    i_8_98_2132_0, i_8_98_2137_0, i_8_98_2151_0, i_8_98_2240_0,
    i_8_98_2275_0,
    o_8_98_0_0  );
  input  i_8_98_12_0, i_8_98_52_0, i_8_98_70_0, i_8_98_115_0,
    i_8_98_139_0, i_8_98_141_0, i_8_98_228_0, i_8_98_230_0, i_8_98_231_0,
    i_8_98_314_0, i_8_98_319_0, i_8_98_334_0, i_8_98_342_0, i_8_98_345_0,
    i_8_98_363_0, i_8_98_366_0, i_8_98_384_0, i_8_98_400_0, i_8_98_420_0,
    i_8_98_430_0, i_8_98_504_0, i_8_98_525_0, i_8_98_538_0, i_8_98_553_0,
    i_8_98_557_0, i_8_98_570_0, i_8_98_571_0, i_8_98_581_0, i_8_98_583_0,
    i_8_98_588_0, i_8_98_600_0, i_8_98_601_0, i_8_98_603_0, i_8_98_628_0,
    i_8_98_634_0, i_8_98_651_0, i_8_98_657_0, i_8_98_696_0, i_8_98_700_0,
    i_8_98_704_0, i_8_98_732_0, i_8_98_777_0, i_8_98_781_0, i_8_98_819_0,
    i_8_98_831_0, i_8_98_840_0, i_8_98_842_0, i_8_98_843_0, i_8_98_875_0,
    i_8_98_877_0, i_8_98_879_0, i_8_98_895_0, i_8_98_947_0, i_8_98_993_0,
    i_8_98_1003_0, i_8_98_1105_0, i_8_98_1109_0, i_8_98_1115_0,
    i_8_98_1124_0, i_8_98_1156_0, i_8_98_1267_0, i_8_98_1282_0,
    i_8_98_1284_0, i_8_98_1315_0, i_8_98_1317_0, i_8_98_1320_0,
    i_8_98_1347_0, i_8_98_1354_0, i_8_98_1358_0, i_8_98_1366_0,
    i_8_98_1423_0, i_8_98_1426_0, i_8_98_1453_0, i_8_98_1462_0,
    i_8_98_1490_0, i_8_98_1509_0, i_8_98_1519_0, i_8_98_1524_0,
    i_8_98_1551_0, i_8_98_1633_0, i_8_98_1635_0, i_8_98_1680_0,
    i_8_98_1686_0, i_8_98_1690_0, i_8_98_1695_0, i_8_98_1699_0,
    i_8_98_1700_0, i_8_98_1703_0, i_8_98_1723_0, i_8_98_1770_0,
    i_8_98_1780_0, i_8_98_1884_0, i_8_98_1911_0, i_8_98_1956_0,
    i_8_98_1995_0, i_8_98_2132_0, i_8_98_2137_0, i_8_98_2151_0,
    i_8_98_2240_0, i_8_98_2275_0;
  output o_8_98_0_0;
  assign o_8_98_0_0 = 0;
endmodule



// Benchmark "kernel_8_99" written by ABC on Sun Jul 19 10:04:43 2020

module kernel_8_99 ( 
    i_8_99_13_0, i_8_99_34_0, i_8_99_35_0, i_8_99_57_0, i_8_99_67_0,
    i_8_99_97_0, i_8_99_127_0, i_8_99_129_0, i_8_99_255_0, i_8_99_299_0,
    i_8_99_310_0, i_8_99_344_0, i_8_99_364_0, i_8_99_365_0, i_8_99_422_0,
    i_8_99_423_0, i_8_99_480_0, i_8_99_483_0, i_8_99_517_0, i_8_99_523_0,
    i_8_99_528_0, i_8_99_530_0, i_8_99_545_0, i_8_99_571_0, i_8_99_580_0,
    i_8_99_607_0, i_8_99_608_0, i_8_99_631_0, i_8_99_649_0, i_8_99_679_0,
    i_8_99_680_0, i_8_99_705_0, i_8_99_707_0, i_8_99_799_0, i_8_99_826_0,
    i_8_99_839_0, i_8_99_857_0, i_8_99_866_0, i_8_99_964_0, i_8_99_993_0,
    i_8_99_994_0, i_8_99_1013_0, i_8_99_1050_0, i_8_99_1065_0,
    i_8_99_1110_0, i_8_99_1111_0, i_8_99_1153_0, i_8_99_1202_0,
    i_8_99_1237_0, i_8_99_1246_0, i_8_99_1267_0, i_8_99_1270_0,
    i_8_99_1305_0, i_8_99_1306_0, i_8_99_1307_0, i_8_99_1318_0,
    i_8_99_1324_0, i_8_99_1399_0, i_8_99_1423_0, i_8_99_1424_0,
    i_8_99_1437_0, i_8_99_1471_0, i_8_99_1472_0, i_8_99_1486_0,
    i_8_99_1525_0, i_8_99_1573_0, i_8_99_1574_0, i_8_99_1624_0,
    i_8_99_1630_0, i_8_99_1632_0, i_8_99_1673_0, i_8_99_1687_0,
    i_8_99_1705_0, i_8_99_1707_0, i_8_99_1743_0, i_8_99_1768_0,
    i_8_99_1784_0, i_8_99_1793_0, i_8_99_1795_0, i_8_99_1819_0,
    i_8_99_1820_0, i_8_99_1935_0, i_8_99_1937_0, i_8_99_1975_0,
    i_8_99_1995_0, i_8_99_2089_0, i_8_99_2090_0, i_8_99_2101_0,
    i_8_99_2104_0, i_8_99_2129_0, i_8_99_2145_0, i_8_99_2149_0,
    i_8_99_2156_0, i_8_99_2214_0, i_8_99_2216_0, i_8_99_2224_0,
    i_8_99_2225_0, i_8_99_2233_0, i_8_99_2245_0, i_8_99_2248_0,
    o_8_99_0_0  );
  input  i_8_99_13_0, i_8_99_34_0, i_8_99_35_0, i_8_99_57_0, i_8_99_67_0,
    i_8_99_97_0, i_8_99_127_0, i_8_99_129_0, i_8_99_255_0, i_8_99_299_0,
    i_8_99_310_0, i_8_99_344_0, i_8_99_364_0, i_8_99_365_0, i_8_99_422_0,
    i_8_99_423_0, i_8_99_480_0, i_8_99_483_0, i_8_99_517_0, i_8_99_523_0,
    i_8_99_528_0, i_8_99_530_0, i_8_99_545_0, i_8_99_571_0, i_8_99_580_0,
    i_8_99_607_0, i_8_99_608_0, i_8_99_631_0, i_8_99_649_0, i_8_99_679_0,
    i_8_99_680_0, i_8_99_705_0, i_8_99_707_0, i_8_99_799_0, i_8_99_826_0,
    i_8_99_839_0, i_8_99_857_0, i_8_99_866_0, i_8_99_964_0, i_8_99_993_0,
    i_8_99_994_0, i_8_99_1013_0, i_8_99_1050_0, i_8_99_1065_0,
    i_8_99_1110_0, i_8_99_1111_0, i_8_99_1153_0, i_8_99_1202_0,
    i_8_99_1237_0, i_8_99_1246_0, i_8_99_1267_0, i_8_99_1270_0,
    i_8_99_1305_0, i_8_99_1306_0, i_8_99_1307_0, i_8_99_1318_0,
    i_8_99_1324_0, i_8_99_1399_0, i_8_99_1423_0, i_8_99_1424_0,
    i_8_99_1437_0, i_8_99_1471_0, i_8_99_1472_0, i_8_99_1486_0,
    i_8_99_1525_0, i_8_99_1573_0, i_8_99_1574_0, i_8_99_1624_0,
    i_8_99_1630_0, i_8_99_1632_0, i_8_99_1673_0, i_8_99_1687_0,
    i_8_99_1705_0, i_8_99_1707_0, i_8_99_1743_0, i_8_99_1768_0,
    i_8_99_1784_0, i_8_99_1793_0, i_8_99_1795_0, i_8_99_1819_0,
    i_8_99_1820_0, i_8_99_1935_0, i_8_99_1937_0, i_8_99_1975_0,
    i_8_99_1995_0, i_8_99_2089_0, i_8_99_2090_0, i_8_99_2101_0,
    i_8_99_2104_0, i_8_99_2129_0, i_8_99_2145_0, i_8_99_2149_0,
    i_8_99_2156_0, i_8_99_2214_0, i_8_99_2216_0, i_8_99_2224_0,
    i_8_99_2225_0, i_8_99_2233_0, i_8_99_2245_0, i_8_99_2248_0;
  output o_8_99_0_0;
  assign o_8_99_0_0 = 0;
endmodule



// Benchmark "kernel_8_100" written by ABC on Sun Jul 19 10:04:44 2020

module kernel_8_100 ( 
    i_8_100_48_0, i_8_100_50_0, i_8_100_111_0, i_8_100_165_0,
    i_8_100_187_0, i_8_100_226_0, i_8_100_231_0, i_8_100_256_0,
    i_8_100_367_0, i_8_100_373_0, i_8_100_391_0, i_8_100_415_0,
    i_8_100_433_0, i_8_100_444_0, i_8_100_481_0, i_8_100_490_0,
    i_8_100_493_0, i_8_100_504_0, i_8_100_507_0, i_8_100_549_0,
    i_8_100_552_0, i_8_100_553_0, i_8_100_554_0, i_8_100_599_0,
    i_8_100_602_0, i_8_100_630_0, i_8_100_659_0, i_8_100_692_0,
    i_8_100_715_0, i_8_100_778_0, i_8_100_781_0, i_8_100_782_0,
    i_8_100_786_0, i_8_100_804_0, i_8_100_816_0, i_8_100_841_0,
    i_8_100_850_0, i_8_100_931_0, i_8_100_1047_0, i_8_100_1050_0,
    i_8_100_1051_0, i_8_100_1104_0, i_8_100_1110_0, i_8_100_1111_0,
    i_8_100_1120_0, i_8_100_1140_0, i_8_100_1162_0, i_8_100_1185_0,
    i_8_100_1236_0, i_8_100_1265_0, i_8_100_1270_0, i_8_100_1281_0,
    i_8_100_1282_0, i_8_100_1283_0, i_8_100_1285_0, i_8_100_1286_0,
    i_8_100_1306_0, i_8_100_1307_0, i_8_100_1327_0, i_8_100_1331_0,
    i_8_100_1390_0, i_8_100_1396_0, i_8_100_1404_0, i_8_100_1405_0,
    i_8_100_1407_0, i_8_100_1438_0, i_8_100_1506_0, i_8_100_1509_0,
    i_8_100_1536_0, i_8_100_1561_0, i_8_100_1590_0, i_8_100_1641_0,
    i_8_100_1649_0, i_8_100_1650_0, i_8_100_1719_0, i_8_100_1722_0,
    i_8_100_1724_0, i_8_100_1741_0, i_8_100_1846_0, i_8_100_1856_0,
    i_8_100_1857_0, i_8_100_1858_0, i_8_100_1866_0, i_8_100_1873_0,
    i_8_100_1884_0, i_8_100_1903_0, i_8_100_1904_0, i_8_100_1956_0,
    i_8_100_1958_0, i_8_100_2010_0, i_8_100_2016_0, i_8_100_2127_0,
    i_8_100_2140_0, i_8_100_2173_0, i_8_100_2214_0, i_8_100_2215_0,
    i_8_100_2216_0, i_8_100_2236_0, i_8_100_2261_0, i_8_100_2299_0,
    o_8_100_0_0  );
  input  i_8_100_48_0, i_8_100_50_0, i_8_100_111_0, i_8_100_165_0,
    i_8_100_187_0, i_8_100_226_0, i_8_100_231_0, i_8_100_256_0,
    i_8_100_367_0, i_8_100_373_0, i_8_100_391_0, i_8_100_415_0,
    i_8_100_433_0, i_8_100_444_0, i_8_100_481_0, i_8_100_490_0,
    i_8_100_493_0, i_8_100_504_0, i_8_100_507_0, i_8_100_549_0,
    i_8_100_552_0, i_8_100_553_0, i_8_100_554_0, i_8_100_599_0,
    i_8_100_602_0, i_8_100_630_0, i_8_100_659_0, i_8_100_692_0,
    i_8_100_715_0, i_8_100_778_0, i_8_100_781_0, i_8_100_782_0,
    i_8_100_786_0, i_8_100_804_0, i_8_100_816_0, i_8_100_841_0,
    i_8_100_850_0, i_8_100_931_0, i_8_100_1047_0, i_8_100_1050_0,
    i_8_100_1051_0, i_8_100_1104_0, i_8_100_1110_0, i_8_100_1111_0,
    i_8_100_1120_0, i_8_100_1140_0, i_8_100_1162_0, i_8_100_1185_0,
    i_8_100_1236_0, i_8_100_1265_0, i_8_100_1270_0, i_8_100_1281_0,
    i_8_100_1282_0, i_8_100_1283_0, i_8_100_1285_0, i_8_100_1286_0,
    i_8_100_1306_0, i_8_100_1307_0, i_8_100_1327_0, i_8_100_1331_0,
    i_8_100_1390_0, i_8_100_1396_0, i_8_100_1404_0, i_8_100_1405_0,
    i_8_100_1407_0, i_8_100_1438_0, i_8_100_1506_0, i_8_100_1509_0,
    i_8_100_1536_0, i_8_100_1561_0, i_8_100_1590_0, i_8_100_1641_0,
    i_8_100_1649_0, i_8_100_1650_0, i_8_100_1719_0, i_8_100_1722_0,
    i_8_100_1724_0, i_8_100_1741_0, i_8_100_1846_0, i_8_100_1856_0,
    i_8_100_1857_0, i_8_100_1858_0, i_8_100_1866_0, i_8_100_1873_0,
    i_8_100_1884_0, i_8_100_1903_0, i_8_100_1904_0, i_8_100_1956_0,
    i_8_100_1958_0, i_8_100_2010_0, i_8_100_2016_0, i_8_100_2127_0,
    i_8_100_2140_0, i_8_100_2173_0, i_8_100_2214_0, i_8_100_2215_0,
    i_8_100_2216_0, i_8_100_2236_0, i_8_100_2261_0, i_8_100_2299_0;
  output o_8_100_0_0;
  assign o_8_100_0_0 = ~((~i_8_100_48_0 & ((i_8_100_481_0 & i_8_100_778_0 & i_8_100_1110_0) | (i_8_100_1396_0 & i_8_100_1719_0 & ~i_8_100_1903_0 & ~i_8_100_2215_0))) | (~i_8_100_50_0 & ((~i_8_100_187_0 & ~i_8_100_481_0 & ~i_8_100_1047_0 & ~i_8_100_1265_0 & ~i_8_100_1270_0 & ~i_8_100_1390_0 & ~i_8_100_1438_0 & ~i_8_100_1956_0 & ~i_8_100_2140_0) | (~i_8_100_444_0 & ~i_8_100_507_0 & ~i_8_100_630_0 & ~i_8_100_778_0 & ~i_8_100_931_0 & ~i_8_100_1404_0 & ~i_8_100_1561_0 & ~i_8_100_2215_0))) | (~i_8_100_226_0 & ((~i_8_100_187_0 & i_8_100_367_0 & ~i_8_100_804_0 & ~i_8_100_1162_0) | (~i_8_100_850_0 & i_8_100_1281_0))) | (~i_8_100_256_0 & ((i_8_100_490_0 & ~i_8_100_554_0 & ~i_8_100_786_0 & ~i_8_100_1396_0 & ~i_8_100_1722_0) | (~i_8_100_187_0 & i_8_100_549_0 & ~i_8_100_1104_0 & ~i_8_100_1561_0 & ~i_8_100_1903_0 & ~i_8_100_1904_0 & ~i_8_100_2173_0))) | (~i_8_100_187_0 & ~i_8_100_1506_0 & ((~i_8_100_373_0 & ~i_8_100_415_0 & ~i_8_100_444_0 & ~i_8_100_1307_0 & ~i_8_100_1396_0 & ~i_8_100_1561_0 & ~i_8_100_1956_0) | (~i_8_100_433_0 & ~i_8_100_504_0 & ~i_8_100_786_0 & ~i_8_100_1390_0 & ~i_8_100_1866_0 & ~i_8_100_1873_0 & ~i_8_100_1904_0 & ~i_8_100_2215_0))) | (~i_8_100_433_0 & ((~i_8_100_507_0 & ~i_8_100_692_0 & i_8_100_1282_0) | (i_8_100_481_0 & ~i_8_100_490_0 & ~i_8_100_786_0 & ~i_8_100_816_0 & ~i_8_100_1307_0 & ~i_8_100_1390_0 & ~i_8_100_1438_0 & ~i_8_100_1641_0 & ~i_8_100_1866_0))) | (~i_8_100_786_0 & ((~i_8_100_444_0 & ((~i_8_100_549_0 & ~i_8_100_602_0 & ~i_8_100_630_0 & ~i_8_100_1306_0 & ~i_8_100_1719_0 & ~i_8_100_1724_0 & ~i_8_100_1866_0 & ~i_8_100_1873_0 & ~i_8_100_2016_0 & ~i_8_100_2140_0) | (i_8_100_490_0 & ~i_8_100_1140_0 & ~i_8_100_1509_0 & ~i_8_100_1741_0 & ~i_8_100_2010_0 & ~i_8_100_2173_0))) | (i_8_100_1110_0 & i_8_100_1111_0 & ~i_8_100_1120_0 & ~i_8_100_1306_0 & ~i_8_100_1307_0 & ~i_8_100_1858_0) | (~i_8_100_481_0 & ~i_8_100_816_0 & ~i_8_100_1331_0 & ~i_8_100_1509_0 & ~i_8_100_1649_0 & ~i_8_100_1741_0 & ~i_8_100_1873_0 & ~i_8_100_1956_0 & ~i_8_100_2214_0))) | (~i_8_100_504_0 & ((i_8_100_778_0 & ~i_8_100_1390_0) | (~i_8_100_630_0 & ~i_8_100_1561_0 & ~i_8_100_1724_0 & i_8_100_2127_0))) | (~i_8_100_1120_0 & ((~i_8_100_507_0 & ~i_8_100_1270_0 & i_8_100_1438_0 & ~i_8_100_1956_0) | (~i_8_100_850_0 & i_8_100_1327_0 & ~i_8_100_1438_0 & ~i_8_100_2214_0))) | (~i_8_100_2236_0 & ((~i_8_100_493_0 & i_8_100_786_0 & i_8_100_841_0 & ~i_8_100_1306_0) | (i_8_100_554_0 & ~i_8_100_1404_0))) | (~i_8_100_165_0 & i_8_100_444_0 & ~i_8_100_481_0 & ~i_8_100_1846_0 & i_8_100_1884_0 & ~i_8_100_1956_0) | (~i_8_100_1047_0 & ~i_8_100_1050_0 & ~i_8_100_1140_0 & i_8_100_1285_0 & ~i_8_100_1958_0) | (i_8_100_493_0 & i_8_100_1649_0 & ~i_8_100_1866_0 & ~i_8_100_2140_0) | (i_8_100_391_0 & i_8_100_549_0 & ~i_8_100_1561_0 & i_8_100_2173_0) | (i_8_100_782_0 & i_8_100_2261_0) | (~i_8_100_415_0 & i_8_100_1282_0 & ~i_8_100_1719_0 & ~i_8_100_1724_0 & ~i_8_100_1873_0 & ~i_8_100_2299_0));
endmodule



// Benchmark "kernel_8_101" written by ABC on Sun Jul 19 10:04:46 2020

module kernel_8_101 ( 
    i_8_101_1_0, i_8_101_5_0, i_8_101_53_0, i_8_101_65_0, i_8_101_75_0,
    i_8_101_167_0, i_8_101_185_0, i_8_101_200_0, i_8_101_217_0,
    i_8_101_221_0, i_8_101_226_0, i_8_101_227_0, i_8_101_262_0,
    i_8_101_266_0, i_8_101_343_0, i_8_101_360_0, i_8_101_363_0,
    i_8_101_364_0, i_8_101_398_0, i_8_101_424_0, i_8_101_425_0,
    i_8_101_452_0, i_8_101_454_0, i_8_101_490_0, i_8_101_493_0,
    i_8_101_505_0, i_8_101_525_0, i_8_101_581_0, i_8_101_584_0,
    i_8_101_587_0, i_8_101_608_0, i_8_101_611_0, i_8_101_624_0,
    i_8_101_640_0, i_8_101_696_0, i_8_101_724_0, i_8_101_730_0,
    i_8_101_731_0, i_8_101_803_0, i_8_101_806_0, i_8_101_809_0,
    i_8_101_873_0, i_8_101_883_0, i_8_101_935_0, i_8_101_956_0,
    i_8_101_963_0, i_8_101_968_0, i_8_101_980_0, i_8_101_992_0,
    i_8_101_995_0, i_8_101_1073_0, i_8_101_1075_0, i_8_101_1076_0,
    i_8_101_1114_0, i_8_101_1127_0, i_8_101_1171_0, i_8_101_1229_0,
    i_8_101_1234_0, i_8_101_1238_0, i_8_101_1259_0, i_8_101_1274_0,
    i_8_101_1289_0, i_8_101_1298_0, i_8_101_1325_0, i_8_101_1355_0,
    i_8_101_1382_0, i_8_101_1385_0, i_8_101_1391_0, i_8_101_1441_0,
    i_8_101_1487_0, i_8_101_1492_0, i_8_101_1628_0, i_8_101_1636_0,
    i_8_101_1691_0, i_8_101_1703_0, i_8_101_1752_0, i_8_101_1759_0,
    i_8_101_1778_0, i_8_101_1792_0, i_8_101_1793_0, i_8_101_1823_0,
    i_8_101_1847_0, i_8_101_1850_0, i_8_101_1882_0, i_8_101_1909_0,
    i_8_101_1910_0, i_8_101_1980_0, i_8_101_1981_0, i_8_101_1982_0,
    i_8_101_1994_0, i_8_101_2018_0, i_8_101_2078_0, i_8_101_2099_0,
    i_8_101_2139_0, i_8_101_2140_0, i_8_101_2144_0, i_8_101_2147_0,
    i_8_101_2172_0, i_8_101_2213_0, i_8_101_2297_0,
    o_8_101_0_0  );
  input  i_8_101_1_0, i_8_101_5_0, i_8_101_53_0, i_8_101_65_0,
    i_8_101_75_0, i_8_101_167_0, i_8_101_185_0, i_8_101_200_0,
    i_8_101_217_0, i_8_101_221_0, i_8_101_226_0, i_8_101_227_0,
    i_8_101_262_0, i_8_101_266_0, i_8_101_343_0, i_8_101_360_0,
    i_8_101_363_0, i_8_101_364_0, i_8_101_398_0, i_8_101_424_0,
    i_8_101_425_0, i_8_101_452_0, i_8_101_454_0, i_8_101_490_0,
    i_8_101_493_0, i_8_101_505_0, i_8_101_525_0, i_8_101_581_0,
    i_8_101_584_0, i_8_101_587_0, i_8_101_608_0, i_8_101_611_0,
    i_8_101_624_0, i_8_101_640_0, i_8_101_696_0, i_8_101_724_0,
    i_8_101_730_0, i_8_101_731_0, i_8_101_803_0, i_8_101_806_0,
    i_8_101_809_0, i_8_101_873_0, i_8_101_883_0, i_8_101_935_0,
    i_8_101_956_0, i_8_101_963_0, i_8_101_968_0, i_8_101_980_0,
    i_8_101_992_0, i_8_101_995_0, i_8_101_1073_0, i_8_101_1075_0,
    i_8_101_1076_0, i_8_101_1114_0, i_8_101_1127_0, i_8_101_1171_0,
    i_8_101_1229_0, i_8_101_1234_0, i_8_101_1238_0, i_8_101_1259_0,
    i_8_101_1274_0, i_8_101_1289_0, i_8_101_1298_0, i_8_101_1325_0,
    i_8_101_1355_0, i_8_101_1382_0, i_8_101_1385_0, i_8_101_1391_0,
    i_8_101_1441_0, i_8_101_1487_0, i_8_101_1492_0, i_8_101_1628_0,
    i_8_101_1636_0, i_8_101_1691_0, i_8_101_1703_0, i_8_101_1752_0,
    i_8_101_1759_0, i_8_101_1778_0, i_8_101_1792_0, i_8_101_1793_0,
    i_8_101_1823_0, i_8_101_1847_0, i_8_101_1850_0, i_8_101_1882_0,
    i_8_101_1909_0, i_8_101_1910_0, i_8_101_1980_0, i_8_101_1981_0,
    i_8_101_1982_0, i_8_101_1994_0, i_8_101_2018_0, i_8_101_2078_0,
    i_8_101_2099_0, i_8_101_2139_0, i_8_101_2140_0, i_8_101_2144_0,
    i_8_101_2147_0, i_8_101_2172_0, i_8_101_2213_0, i_8_101_2297_0;
  output o_8_101_0_0;
  assign o_8_101_0_0 = ~((i_8_101_227_0 & ((~i_8_101_167_0 & ~i_8_101_505_0 & ~i_8_101_1259_0 & ~i_8_101_1289_0 & ~i_8_101_1298_0) | (~i_8_101_1_0 & ~i_8_101_53_0 & ~i_8_101_266_0 & ~i_8_101_724_0 & ~i_8_101_1274_0 & ~i_8_101_1385_0 & ~i_8_101_1793_0 & ~i_8_101_2018_0))) | (~i_8_101_806_0 & ((~i_8_101_5_0 & ~i_8_101_611_0 & ((~i_8_101_1_0 & ~i_8_101_167_0 & ~i_8_101_360_0 & ~i_8_101_505_0 & ~i_8_101_803_0 & ~i_8_101_980_0 & ~i_8_101_995_0 & ~i_8_101_1075_0 & ~i_8_101_1298_0 & ~i_8_101_1325_0 & ~i_8_101_1703_0) | (~i_8_101_363_0 & ~i_8_101_452_0 & ~i_8_101_490_0 & ~i_8_101_731_0 & ~i_8_101_1259_0 & ~i_8_101_1289_0 & ~i_8_101_1441_0 & ~i_8_101_1981_0))) | (~i_8_101_731_0 & ((~i_8_101_1_0 & ~i_8_101_935_0 & ((~i_8_101_581_0 & ~i_8_101_724_0 & ~i_8_101_883_0 & ~i_8_101_1114_0 & ~i_8_101_1229_0 & ~i_8_101_1441_0 & ~i_8_101_1909_0 & i_8_101_2147_0) | (~i_8_101_227_0 & ~i_8_101_584_0 & ~i_8_101_640_0 & ~i_8_101_803_0 & ~i_8_101_1075_0 & ~i_8_101_1487_0 & ~i_8_101_1703_0 & ~i_8_101_2213_0))) | (~i_8_101_167_0 & ~i_8_101_581_0 & ~i_8_101_584_0 & ~i_8_101_724_0 & ~i_8_101_963_0 & ~i_8_101_1171_0 & ~i_8_101_1910_0 & ~i_8_101_2147_0))))) | (~i_8_101_1_0 & ((~i_8_101_65_0 & ~i_8_101_730_0 & ~i_8_101_731_0 & ~i_8_101_803_0 & ~i_8_101_935_0 & ~i_8_101_968_0 & ~i_8_101_1382_0 & ~i_8_101_1628_0 & ~i_8_101_1909_0) | (~i_8_101_200_0 & ~i_8_101_640_0 & ~i_8_101_1229_0 & ~i_8_101_1259_0 & ~i_8_101_1298_0 & ~i_8_101_1847_0 & ~i_8_101_2147_0))) | (~i_8_101_1910_0 & ((~i_8_101_1850_0 & ((~i_8_101_5_0 & ~i_8_101_640_0 & ~i_8_101_1793_0 & ~i_8_101_1909_0 & ((~i_8_101_65_0 & ~i_8_101_185_0 & ~i_8_101_452_0 & ~i_8_101_956_0 & ~i_8_101_1171_0 & ~i_8_101_1628_0) | (~i_8_101_398_0 & ~i_8_101_584_0 & ~i_8_101_611_0 & ~i_8_101_935_0 & ~i_8_101_980_0 & ~i_8_101_1382_0 & ~i_8_101_1703_0 & ~i_8_101_1847_0))) | (~i_8_101_53_0 & ~i_8_101_185_0 & ~i_8_101_490_0 & ~i_8_101_505_0 & ~i_8_101_611_0 & ~i_8_101_803_0 & ~i_8_101_968_0 & ~i_8_101_1691_0))) | (~i_8_101_1847_0 & ((~i_8_101_53_0 & ~i_8_101_185_0 & ~i_8_101_425_0 & ~i_8_101_452_0 & ~i_8_101_587_0 & ~i_8_101_1234_0 & ~i_8_101_1259_0 & ~i_8_101_2213_0) | (~i_8_101_65_0 & ~i_8_101_266_0 & ~i_8_101_493_0 & i_8_101_611_0 & ~i_8_101_1385_0 & i_8_101_2147_0 & ~i_8_101_2297_0))) | (i_8_101_424_0 & ~i_8_101_581_0 & ~i_8_101_731_0 & ~i_8_101_968_0 & ~i_8_101_995_0 & ~i_8_101_1274_0 & ~i_8_101_1325_0))) | (~i_8_101_53_0 & ((i_8_101_364_0 & i_8_101_424_0 & ~i_8_101_696_0 & ~i_8_101_730_0 & ~i_8_101_1289_0 & ~i_8_101_1325_0 & ~i_8_101_1636_0) | (~i_8_101_5_0 & ~i_8_101_581_0 & ~i_8_101_809_0 & ~i_8_101_956_0 & ~i_8_101_1487_0 & ~i_8_101_1628_0 & ~i_8_101_1847_0 & ~i_8_101_1909_0 & ~i_8_101_2078_0))) | (~i_8_101_803_0 & ((~i_8_101_262_0 & ~i_8_101_398_0 & i_8_101_608_0 & ~i_8_101_956_0 & ~i_8_101_1171_0 & ~i_8_101_1385_0 & ~i_8_101_1703_0 & ~i_8_101_1759_0 & ~i_8_101_1793_0) | (i_8_101_452_0 & i_8_101_525_0 & ~i_8_101_1847_0))) | (~i_8_101_1274_0 & ((~i_8_101_1259_0 & ~i_8_101_1382_0 & i_8_101_1385_0 & ~i_8_101_1703_0 & i_8_101_1823_0) | (~i_8_101_424_0 & ~i_8_101_581_0 & ~i_8_101_935_0 & ~i_8_101_1076_0 & ~i_8_101_1850_0 & ~i_8_101_2144_0 & ~i_8_101_2297_0))));
endmodule



// Benchmark "kernel_8_102" written by ABC on Sun Jul 19 10:04:47 2020

module kernel_8_102 ( 
    i_8_102_28_0, i_8_102_32_0, i_8_102_35_0, i_8_102_89_0, i_8_102_157_0,
    i_8_102_169_0, i_8_102_224_0, i_8_102_283_0, i_8_102_292_0,
    i_8_102_355_0, i_8_102_437_0, i_8_102_455_0, i_8_102_480_0,
    i_8_102_529_0, i_8_102_544_0, i_8_102_552_0, i_8_102_557_0,
    i_8_102_609_0, i_8_102_617_0, i_8_102_658_0, i_8_102_659_0,
    i_8_102_663_0, i_8_102_665_0, i_8_102_703_0, i_8_102_718_0,
    i_8_102_769_0, i_8_102_772_0, i_8_102_850_0, i_8_102_881_0,
    i_8_102_890_0, i_8_102_896_0, i_8_102_951_0, i_8_102_955_0,
    i_8_102_973_0, i_8_102_977_0, i_8_102_1013_0, i_8_102_1032_0,
    i_8_102_1048_0, i_8_102_1050_0, i_8_102_1066_0, i_8_102_1075_0,
    i_8_102_1084_0, i_8_102_1135_0, i_8_102_1137_0, i_8_102_1154_0,
    i_8_102_1157_0, i_8_102_1223_0, i_8_102_1246_0, i_8_102_1247_0,
    i_8_102_1249_0, i_8_102_1256_0, i_8_102_1258_0, i_8_102_1259_0,
    i_8_102_1265_0, i_8_102_1282_0, i_8_102_1283_0, i_8_102_1285_0,
    i_8_102_1297_0, i_8_102_1346_0, i_8_102_1350_0, i_8_102_1367_0,
    i_8_102_1436_0, i_8_102_1449_0, i_8_102_1453_0, i_8_102_1467_0,
    i_8_102_1468_0, i_8_102_1471_0, i_8_102_1482_0, i_8_102_1501_0,
    i_8_102_1502_0, i_8_102_1532_0, i_8_102_1549_0, i_8_102_1577_0,
    i_8_102_1580_0, i_8_102_1613_0, i_8_102_1679_0, i_8_102_1718_0,
    i_8_102_1731_0, i_8_102_1760_0, i_8_102_1771_0, i_8_102_1772_0,
    i_8_102_1776_0, i_8_102_1787_0, i_8_102_1855_0, i_8_102_1856_0,
    i_8_102_1928_0, i_8_102_1931_0, i_8_102_1948_0, i_8_102_1951_0,
    i_8_102_1960_0, i_8_102_2000_0, i_8_102_2030_0, i_8_102_2084_0,
    i_8_102_2143_0, i_8_102_2171_0, i_8_102_2179_0, i_8_102_2214_0,
    i_8_102_2263_0, i_8_102_2264_0, i_8_102_2290_0,
    o_8_102_0_0  );
  input  i_8_102_28_0, i_8_102_32_0, i_8_102_35_0, i_8_102_89_0,
    i_8_102_157_0, i_8_102_169_0, i_8_102_224_0, i_8_102_283_0,
    i_8_102_292_0, i_8_102_355_0, i_8_102_437_0, i_8_102_455_0,
    i_8_102_480_0, i_8_102_529_0, i_8_102_544_0, i_8_102_552_0,
    i_8_102_557_0, i_8_102_609_0, i_8_102_617_0, i_8_102_658_0,
    i_8_102_659_0, i_8_102_663_0, i_8_102_665_0, i_8_102_703_0,
    i_8_102_718_0, i_8_102_769_0, i_8_102_772_0, i_8_102_850_0,
    i_8_102_881_0, i_8_102_890_0, i_8_102_896_0, i_8_102_951_0,
    i_8_102_955_0, i_8_102_973_0, i_8_102_977_0, i_8_102_1013_0,
    i_8_102_1032_0, i_8_102_1048_0, i_8_102_1050_0, i_8_102_1066_0,
    i_8_102_1075_0, i_8_102_1084_0, i_8_102_1135_0, i_8_102_1137_0,
    i_8_102_1154_0, i_8_102_1157_0, i_8_102_1223_0, i_8_102_1246_0,
    i_8_102_1247_0, i_8_102_1249_0, i_8_102_1256_0, i_8_102_1258_0,
    i_8_102_1259_0, i_8_102_1265_0, i_8_102_1282_0, i_8_102_1283_0,
    i_8_102_1285_0, i_8_102_1297_0, i_8_102_1346_0, i_8_102_1350_0,
    i_8_102_1367_0, i_8_102_1436_0, i_8_102_1449_0, i_8_102_1453_0,
    i_8_102_1467_0, i_8_102_1468_0, i_8_102_1471_0, i_8_102_1482_0,
    i_8_102_1501_0, i_8_102_1502_0, i_8_102_1532_0, i_8_102_1549_0,
    i_8_102_1577_0, i_8_102_1580_0, i_8_102_1613_0, i_8_102_1679_0,
    i_8_102_1718_0, i_8_102_1731_0, i_8_102_1760_0, i_8_102_1771_0,
    i_8_102_1772_0, i_8_102_1776_0, i_8_102_1787_0, i_8_102_1855_0,
    i_8_102_1856_0, i_8_102_1928_0, i_8_102_1931_0, i_8_102_1948_0,
    i_8_102_1951_0, i_8_102_1960_0, i_8_102_2000_0, i_8_102_2030_0,
    i_8_102_2084_0, i_8_102_2143_0, i_8_102_2171_0, i_8_102_2179_0,
    i_8_102_2214_0, i_8_102_2263_0, i_8_102_2264_0, i_8_102_2290_0;
  output o_8_102_0_0;
  assign o_8_102_0_0 = 0;
endmodule



// Benchmark "kernel_8_103" written by ABC on Sun Jul 19 10:04:47 2020

module kernel_8_103 ( 
    i_8_103_23_0, i_8_103_26_0, i_8_103_33_0, i_8_103_34_0, i_8_103_35_0,
    i_8_103_61_0, i_8_103_73_0, i_8_103_87_0, i_8_103_114_0, i_8_103_168_0,
    i_8_103_189_0, i_8_103_190_0, i_8_103_223_0, i_8_103_240_0,
    i_8_103_241_0, i_8_103_340_0, i_8_103_375_0, i_8_103_437_0,
    i_8_103_469_0, i_8_103_470_0, i_8_103_483_0, i_8_103_484_0,
    i_8_103_525_0, i_8_103_527_0, i_8_103_574_0, i_8_103_575_0,
    i_8_103_602_0, i_8_103_619_0, i_8_103_636_0, i_8_103_637_0,
    i_8_103_679_0, i_8_103_690_0, i_8_103_691_0, i_8_103_763_0,
    i_8_103_781_0, i_8_103_826_0, i_8_103_861_0, i_8_103_889_0,
    i_8_103_934_0, i_8_103_943_0, i_8_103_944_0, i_8_103_970_0,
    i_8_103_994_0, i_8_103_995_0, i_8_103_1059_0, i_8_103_1060_0,
    i_8_103_1074_0, i_8_103_1111_0, i_8_103_1114_0, i_8_103_1185_0,
    i_8_103_1191_0, i_8_103_1260_0, i_8_103_1284_0, i_8_103_1285_0,
    i_8_103_1295_0, i_8_103_1303_0, i_8_103_1304_0, i_8_103_1305_0,
    i_8_103_1306_0, i_8_103_1339_0, i_8_103_1439_0, i_8_103_1492_0,
    i_8_103_1536_0, i_8_103_1564_0, i_8_103_1575_0, i_8_103_1576_0,
    i_8_103_1591_0, i_8_103_1647_0, i_8_103_1650_0, i_8_103_1653_0,
    i_8_103_1681_0, i_8_103_1699_0, i_8_103_1700_0, i_8_103_1723_0,
    i_8_103_1742_0, i_8_103_1743_0, i_8_103_1744_0, i_8_103_1745_0,
    i_8_103_1753_0, i_8_103_1762_0, i_8_103_1763_0, i_8_103_1780_0,
    i_8_103_1781_0, i_8_103_1834_0, i_8_103_1844_0, i_8_103_1885_0,
    i_8_103_1887_0, i_8_103_1889_0, i_8_103_2050_0, i_8_103_2059_0,
    i_8_103_2060_0, i_8_103_2074_0, i_8_103_2076_0, i_8_103_2123_0,
    i_8_103_2176_0, i_8_103_2218_0, i_8_103_2219_0, i_8_103_2220_0,
    i_8_103_2247_0, i_8_103_2302_0,
    o_8_103_0_0  );
  input  i_8_103_23_0, i_8_103_26_0, i_8_103_33_0, i_8_103_34_0,
    i_8_103_35_0, i_8_103_61_0, i_8_103_73_0, i_8_103_87_0, i_8_103_114_0,
    i_8_103_168_0, i_8_103_189_0, i_8_103_190_0, i_8_103_223_0,
    i_8_103_240_0, i_8_103_241_0, i_8_103_340_0, i_8_103_375_0,
    i_8_103_437_0, i_8_103_469_0, i_8_103_470_0, i_8_103_483_0,
    i_8_103_484_0, i_8_103_525_0, i_8_103_527_0, i_8_103_574_0,
    i_8_103_575_0, i_8_103_602_0, i_8_103_619_0, i_8_103_636_0,
    i_8_103_637_0, i_8_103_679_0, i_8_103_690_0, i_8_103_691_0,
    i_8_103_763_0, i_8_103_781_0, i_8_103_826_0, i_8_103_861_0,
    i_8_103_889_0, i_8_103_934_0, i_8_103_943_0, i_8_103_944_0,
    i_8_103_970_0, i_8_103_994_0, i_8_103_995_0, i_8_103_1059_0,
    i_8_103_1060_0, i_8_103_1074_0, i_8_103_1111_0, i_8_103_1114_0,
    i_8_103_1185_0, i_8_103_1191_0, i_8_103_1260_0, i_8_103_1284_0,
    i_8_103_1285_0, i_8_103_1295_0, i_8_103_1303_0, i_8_103_1304_0,
    i_8_103_1305_0, i_8_103_1306_0, i_8_103_1339_0, i_8_103_1439_0,
    i_8_103_1492_0, i_8_103_1536_0, i_8_103_1564_0, i_8_103_1575_0,
    i_8_103_1576_0, i_8_103_1591_0, i_8_103_1647_0, i_8_103_1650_0,
    i_8_103_1653_0, i_8_103_1681_0, i_8_103_1699_0, i_8_103_1700_0,
    i_8_103_1723_0, i_8_103_1742_0, i_8_103_1743_0, i_8_103_1744_0,
    i_8_103_1745_0, i_8_103_1753_0, i_8_103_1762_0, i_8_103_1763_0,
    i_8_103_1780_0, i_8_103_1781_0, i_8_103_1834_0, i_8_103_1844_0,
    i_8_103_1885_0, i_8_103_1887_0, i_8_103_1889_0, i_8_103_2050_0,
    i_8_103_2059_0, i_8_103_2060_0, i_8_103_2074_0, i_8_103_2076_0,
    i_8_103_2123_0, i_8_103_2176_0, i_8_103_2218_0, i_8_103_2219_0,
    i_8_103_2220_0, i_8_103_2247_0, i_8_103_2302_0;
  output o_8_103_0_0;
  assign o_8_103_0_0 = 0;
endmodule



// Benchmark "kernel_8_104" written by ABC on Sun Jul 19 10:04:48 2020

module kernel_8_104 ( 
    i_8_104_12_0, i_8_104_63_0, i_8_104_72_0, i_8_104_73_0, i_8_104_84_0,
    i_8_104_181_0, i_8_104_298_0, i_8_104_301_0, i_8_104_318_0,
    i_8_104_319_0, i_8_104_334_0, i_8_104_343_0, i_8_104_361_0,
    i_8_104_387_0, i_8_104_418_0, i_8_104_469_0, i_8_104_492_0,
    i_8_104_504_0, i_8_104_505_0, i_8_104_523_0, i_8_104_540_0,
    i_8_104_558_0, i_8_104_577_0, i_8_104_579_0, i_8_104_588_0,
    i_8_104_603_0, i_8_104_630_0, i_8_104_640_0, i_8_104_651_0,
    i_8_104_652_0, i_8_104_657_0, i_8_104_660_0, i_8_104_678_0,
    i_8_104_687_0, i_8_104_707_0, i_8_104_757_0, i_8_104_819_0,
    i_8_104_823_0, i_8_104_839_0, i_8_104_842_0, i_8_104_856_0,
    i_8_104_882_0, i_8_104_886_0, i_8_104_941_0, i_8_104_954_0,
    i_8_104_969_0, i_8_104_1012_0, i_8_104_1026_0, i_8_104_1056_0,
    i_8_104_1071_0, i_8_104_1135_0, i_8_104_1153_0, i_8_104_1170_0,
    i_8_104_1197_0, i_8_104_1215_0, i_8_104_1225_0, i_8_104_1238_0,
    i_8_104_1261_0, i_8_104_1294_0, i_8_104_1381_0, i_8_104_1395_0,
    i_8_104_1398_0, i_8_104_1423_0, i_8_104_1479_0, i_8_104_1487_0,
    i_8_104_1506_0, i_8_104_1507_0, i_8_104_1512_0, i_8_104_1557_0,
    i_8_104_1570_0, i_8_104_1630_0, i_8_104_1654_0, i_8_104_1668_0,
    i_8_104_1671_0, i_8_104_1681_0, i_8_104_1728_0, i_8_104_1747_0,
    i_8_104_1794_0, i_8_104_1824_0, i_8_104_1825_0, i_8_104_1866_0,
    i_8_104_1918_0, i_8_104_1948_0, i_8_104_1962_0, i_8_104_1963_0,
    i_8_104_1989_0, i_8_104_1992_0, i_8_104_1997_0, i_8_104_2103_0,
    i_8_104_2106_0, i_8_104_2107_0, i_8_104_2115_0, i_8_104_2145_0,
    i_8_104_2149_0, i_8_104_2151_0, i_8_104_2152_0, i_8_104_2162_0,
    i_8_104_2190_0, i_8_104_2232_0, i_8_104_2245_0,
    o_8_104_0_0  );
  input  i_8_104_12_0, i_8_104_63_0, i_8_104_72_0, i_8_104_73_0,
    i_8_104_84_0, i_8_104_181_0, i_8_104_298_0, i_8_104_301_0,
    i_8_104_318_0, i_8_104_319_0, i_8_104_334_0, i_8_104_343_0,
    i_8_104_361_0, i_8_104_387_0, i_8_104_418_0, i_8_104_469_0,
    i_8_104_492_0, i_8_104_504_0, i_8_104_505_0, i_8_104_523_0,
    i_8_104_540_0, i_8_104_558_0, i_8_104_577_0, i_8_104_579_0,
    i_8_104_588_0, i_8_104_603_0, i_8_104_630_0, i_8_104_640_0,
    i_8_104_651_0, i_8_104_652_0, i_8_104_657_0, i_8_104_660_0,
    i_8_104_678_0, i_8_104_687_0, i_8_104_707_0, i_8_104_757_0,
    i_8_104_819_0, i_8_104_823_0, i_8_104_839_0, i_8_104_842_0,
    i_8_104_856_0, i_8_104_882_0, i_8_104_886_0, i_8_104_941_0,
    i_8_104_954_0, i_8_104_969_0, i_8_104_1012_0, i_8_104_1026_0,
    i_8_104_1056_0, i_8_104_1071_0, i_8_104_1135_0, i_8_104_1153_0,
    i_8_104_1170_0, i_8_104_1197_0, i_8_104_1215_0, i_8_104_1225_0,
    i_8_104_1238_0, i_8_104_1261_0, i_8_104_1294_0, i_8_104_1381_0,
    i_8_104_1395_0, i_8_104_1398_0, i_8_104_1423_0, i_8_104_1479_0,
    i_8_104_1487_0, i_8_104_1506_0, i_8_104_1507_0, i_8_104_1512_0,
    i_8_104_1557_0, i_8_104_1570_0, i_8_104_1630_0, i_8_104_1654_0,
    i_8_104_1668_0, i_8_104_1671_0, i_8_104_1681_0, i_8_104_1728_0,
    i_8_104_1747_0, i_8_104_1794_0, i_8_104_1824_0, i_8_104_1825_0,
    i_8_104_1866_0, i_8_104_1918_0, i_8_104_1948_0, i_8_104_1962_0,
    i_8_104_1963_0, i_8_104_1989_0, i_8_104_1992_0, i_8_104_1997_0,
    i_8_104_2103_0, i_8_104_2106_0, i_8_104_2107_0, i_8_104_2115_0,
    i_8_104_2145_0, i_8_104_2149_0, i_8_104_2151_0, i_8_104_2152_0,
    i_8_104_2162_0, i_8_104_2190_0, i_8_104_2232_0, i_8_104_2245_0;
  output o_8_104_0_0;
  assign o_8_104_0_0 = 0;
endmodule



// Benchmark "kernel_8_105" written by ABC on Sun Jul 19 10:04:49 2020

module kernel_8_105 ( 
    i_8_105_32_0, i_8_105_33_0, i_8_105_141_0, i_8_105_142_0,
    i_8_105_146_0, i_8_105_189_0, i_8_105_196_0, i_8_105_318_0,
    i_8_105_358_0, i_8_105_393_0, i_8_105_399_0, i_8_105_421_0,
    i_8_105_462_0, i_8_105_502_0, i_8_105_516_0, i_8_105_524_0,
    i_8_105_594_0, i_8_105_597_0, i_8_105_604_0, i_8_105_624_0,
    i_8_105_679_0, i_8_105_702_0, i_8_105_782_0, i_8_105_789_0,
    i_8_105_811_0, i_8_105_834_0, i_8_105_867_0, i_8_105_941_0,
    i_8_105_970_0, i_8_105_993_0, i_8_105_1012_0, i_8_105_1014_0,
    i_8_105_1075_0, i_8_105_1108_0, i_8_105_1110_0, i_8_105_1128_0,
    i_8_105_1137_0, i_8_105_1167_0, i_8_105_1172_0, i_8_105_1230_0,
    i_8_105_1246_0, i_8_105_1272_0, i_8_105_1278_0, i_8_105_1300_0,
    i_8_105_1301_0, i_8_105_1306_0, i_8_105_1318_0, i_8_105_1326_0,
    i_8_105_1331_0, i_8_105_1337_0, i_8_105_1338_0, i_8_105_1355_0,
    i_8_105_1356_0, i_8_105_1411_0, i_8_105_1426_0, i_8_105_1437_0,
    i_8_105_1467_0, i_8_105_1480_0, i_8_105_1534_0, i_8_105_1546_0,
    i_8_105_1552_0, i_8_105_1596_0, i_8_105_1597_0, i_8_105_1642_0,
    i_8_105_1644_0, i_8_105_1645_0, i_8_105_1650_0, i_8_105_1672_0,
    i_8_105_1707_0, i_8_105_1721_0, i_8_105_1749_0, i_8_105_1785_0,
    i_8_105_1795_0, i_8_105_1800_0, i_8_105_1843_0, i_8_105_1852_0,
    i_8_105_1854_0, i_8_105_1858_0, i_8_105_1875_0, i_8_105_1885_0,
    i_8_105_1947_0, i_8_105_1974_0, i_8_105_1975_0, i_8_105_1986_0,
    i_8_105_2047_0, i_8_105_2064_0, i_8_105_2091_0, i_8_105_2094_0,
    i_8_105_2104_0, i_8_105_2119_0, i_8_105_2123_0, i_8_105_2143_0,
    i_8_105_2148_0, i_8_105_2150_0, i_8_105_2155_0, i_8_105_2169_0,
    i_8_105_2214_0, i_8_105_2216_0, i_8_105_2226_0, i_8_105_2244_0,
    o_8_105_0_0  );
  input  i_8_105_32_0, i_8_105_33_0, i_8_105_141_0, i_8_105_142_0,
    i_8_105_146_0, i_8_105_189_0, i_8_105_196_0, i_8_105_318_0,
    i_8_105_358_0, i_8_105_393_0, i_8_105_399_0, i_8_105_421_0,
    i_8_105_462_0, i_8_105_502_0, i_8_105_516_0, i_8_105_524_0,
    i_8_105_594_0, i_8_105_597_0, i_8_105_604_0, i_8_105_624_0,
    i_8_105_679_0, i_8_105_702_0, i_8_105_782_0, i_8_105_789_0,
    i_8_105_811_0, i_8_105_834_0, i_8_105_867_0, i_8_105_941_0,
    i_8_105_970_0, i_8_105_993_0, i_8_105_1012_0, i_8_105_1014_0,
    i_8_105_1075_0, i_8_105_1108_0, i_8_105_1110_0, i_8_105_1128_0,
    i_8_105_1137_0, i_8_105_1167_0, i_8_105_1172_0, i_8_105_1230_0,
    i_8_105_1246_0, i_8_105_1272_0, i_8_105_1278_0, i_8_105_1300_0,
    i_8_105_1301_0, i_8_105_1306_0, i_8_105_1318_0, i_8_105_1326_0,
    i_8_105_1331_0, i_8_105_1337_0, i_8_105_1338_0, i_8_105_1355_0,
    i_8_105_1356_0, i_8_105_1411_0, i_8_105_1426_0, i_8_105_1437_0,
    i_8_105_1467_0, i_8_105_1480_0, i_8_105_1534_0, i_8_105_1546_0,
    i_8_105_1552_0, i_8_105_1596_0, i_8_105_1597_0, i_8_105_1642_0,
    i_8_105_1644_0, i_8_105_1645_0, i_8_105_1650_0, i_8_105_1672_0,
    i_8_105_1707_0, i_8_105_1721_0, i_8_105_1749_0, i_8_105_1785_0,
    i_8_105_1795_0, i_8_105_1800_0, i_8_105_1843_0, i_8_105_1852_0,
    i_8_105_1854_0, i_8_105_1858_0, i_8_105_1875_0, i_8_105_1885_0,
    i_8_105_1947_0, i_8_105_1974_0, i_8_105_1975_0, i_8_105_1986_0,
    i_8_105_2047_0, i_8_105_2064_0, i_8_105_2091_0, i_8_105_2094_0,
    i_8_105_2104_0, i_8_105_2119_0, i_8_105_2123_0, i_8_105_2143_0,
    i_8_105_2148_0, i_8_105_2150_0, i_8_105_2155_0, i_8_105_2169_0,
    i_8_105_2214_0, i_8_105_2216_0, i_8_105_2226_0, i_8_105_2244_0;
  output o_8_105_0_0;
  assign o_8_105_0_0 = 0;
endmodule



// Benchmark "kernel_8_106" written by ABC on Sun Jul 19 10:04:50 2020

module kernel_8_106 ( 
    i_8_106_34_0, i_8_106_71_0, i_8_106_80_0, i_8_106_88_0, i_8_106_107_0,
    i_8_106_115_0, i_8_106_194_0, i_8_106_228_0, i_8_106_241_0,
    i_8_106_242_0, i_8_106_278_0, i_8_106_304_0, i_8_106_379_0,
    i_8_106_381_0, i_8_106_385_0, i_8_106_424_0, i_8_106_484_0,
    i_8_106_489_0, i_8_106_490_0, i_8_106_492_0, i_8_106_523_0,
    i_8_106_529_0, i_8_106_610_0, i_8_106_634_0, i_8_106_637_0,
    i_8_106_658_0, i_8_106_682_0, i_8_106_694_0, i_8_106_706_0,
    i_8_106_715_0, i_8_106_717_0, i_8_106_723_0, i_8_106_735_0,
    i_8_106_738_0, i_8_106_798_0, i_8_106_799_0, i_8_106_817_0,
    i_8_106_853_0, i_8_106_880_0, i_8_106_994_0, i_8_106_1047_0,
    i_8_106_1048_0, i_8_106_1057_0, i_8_106_1066_0, i_8_106_1084_0,
    i_8_106_1105_0, i_8_106_1114_0, i_8_106_1116_0, i_8_106_1117_0,
    i_8_106_1147_0, i_8_106_1171_0, i_8_106_1225_0, i_8_106_1228_0,
    i_8_106_1235_0, i_8_106_1236_0, i_8_106_1278_0, i_8_106_1285_0,
    i_8_106_1288_0, i_8_106_1333_0, i_8_106_1354_0, i_8_106_1357_0,
    i_8_106_1438_0, i_8_106_1545_0, i_8_106_1552_0, i_8_106_1564_0,
    i_8_106_1605_0, i_8_106_1609_0, i_8_106_1615_0, i_8_106_1627_0,
    i_8_106_1646_0, i_8_106_1648_0, i_8_106_1663_0, i_8_106_1696_0,
    i_8_106_1753_0, i_8_106_1763_0, i_8_106_1771_0, i_8_106_1774_0,
    i_8_106_1785_0, i_8_106_1786_0, i_8_106_1821_0, i_8_106_1825_0,
    i_8_106_1843_0, i_8_106_1849_0, i_8_106_1855_0, i_8_106_1860_0,
    i_8_106_1887_0, i_8_106_1903_0, i_8_106_1914_0, i_8_106_1915_0,
    i_8_106_1986_0, i_8_106_1987_0, i_8_106_1988_0, i_8_106_1996_0,
    i_8_106_2041_0, i_8_106_2121_0, i_8_106_2122_0, i_8_106_2149_0,
    i_8_106_2157_0, i_8_106_2242_0, i_8_106_2292_0,
    o_8_106_0_0  );
  input  i_8_106_34_0, i_8_106_71_0, i_8_106_80_0, i_8_106_88_0,
    i_8_106_107_0, i_8_106_115_0, i_8_106_194_0, i_8_106_228_0,
    i_8_106_241_0, i_8_106_242_0, i_8_106_278_0, i_8_106_304_0,
    i_8_106_379_0, i_8_106_381_0, i_8_106_385_0, i_8_106_424_0,
    i_8_106_484_0, i_8_106_489_0, i_8_106_490_0, i_8_106_492_0,
    i_8_106_523_0, i_8_106_529_0, i_8_106_610_0, i_8_106_634_0,
    i_8_106_637_0, i_8_106_658_0, i_8_106_682_0, i_8_106_694_0,
    i_8_106_706_0, i_8_106_715_0, i_8_106_717_0, i_8_106_723_0,
    i_8_106_735_0, i_8_106_738_0, i_8_106_798_0, i_8_106_799_0,
    i_8_106_817_0, i_8_106_853_0, i_8_106_880_0, i_8_106_994_0,
    i_8_106_1047_0, i_8_106_1048_0, i_8_106_1057_0, i_8_106_1066_0,
    i_8_106_1084_0, i_8_106_1105_0, i_8_106_1114_0, i_8_106_1116_0,
    i_8_106_1117_0, i_8_106_1147_0, i_8_106_1171_0, i_8_106_1225_0,
    i_8_106_1228_0, i_8_106_1235_0, i_8_106_1236_0, i_8_106_1278_0,
    i_8_106_1285_0, i_8_106_1288_0, i_8_106_1333_0, i_8_106_1354_0,
    i_8_106_1357_0, i_8_106_1438_0, i_8_106_1545_0, i_8_106_1552_0,
    i_8_106_1564_0, i_8_106_1605_0, i_8_106_1609_0, i_8_106_1615_0,
    i_8_106_1627_0, i_8_106_1646_0, i_8_106_1648_0, i_8_106_1663_0,
    i_8_106_1696_0, i_8_106_1753_0, i_8_106_1763_0, i_8_106_1771_0,
    i_8_106_1774_0, i_8_106_1785_0, i_8_106_1786_0, i_8_106_1821_0,
    i_8_106_1825_0, i_8_106_1843_0, i_8_106_1849_0, i_8_106_1855_0,
    i_8_106_1860_0, i_8_106_1887_0, i_8_106_1903_0, i_8_106_1914_0,
    i_8_106_1915_0, i_8_106_1986_0, i_8_106_1987_0, i_8_106_1988_0,
    i_8_106_1996_0, i_8_106_2041_0, i_8_106_2121_0, i_8_106_2122_0,
    i_8_106_2149_0, i_8_106_2157_0, i_8_106_2242_0, i_8_106_2292_0;
  output o_8_106_0_0;
  assign o_8_106_0_0 = 0;
endmodule



// Benchmark "kernel_8_107" written by ABC on Sun Jul 19 10:04:51 2020

module kernel_8_107 ( 
    i_8_107_31_0, i_8_107_50_0, i_8_107_86_0, i_8_107_167_0, i_8_107_230_0,
    i_8_107_233_0, i_8_107_234_0, i_8_107_326_0, i_8_107_335_0,
    i_8_107_338_0, i_8_107_365_0, i_8_107_368_0, i_8_107_380_0,
    i_8_107_386_0, i_8_107_400_0, i_8_107_419_0, i_8_107_424_0,
    i_8_107_425_0, i_8_107_428_0, i_8_107_440_0, i_8_107_449_0,
    i_8_107_451_0, i_8_107_452_0, i_8_107_494_0, i_8_107_499_0,
    i_8_107_500_0, i_8_107_581_0, i_8_107_613_0, i_8_107_614_0,
    i_8_107_617_0, i_8_107_655_0, i_8_107_694_0, i_8_107_698_0,
    i_8_107_706_0, i_8_107_707_0, i_8_107_733_0, i_8_107_767_0,
    i_8_107_770_0, i_8_107_796_0, i_8_107_797_0, i_8_107_839_0,
    i_8_107_842_0, i_8_107_845_0, i_8_107_878_0, i_8_107_932_0,
    i_8_107_956_0, i_8_107_968_0, i_8_107_1019_0, i_8_107_1022_0,
    i_8_107_1058_0, i_8_107_1097_0, i_8_107_1106_0, i_8_107_1157_0,
    i_8_107_1229_0, i_8_107_1235_0, i_8_107_1238_0, i_8_107_1253_0,
    i_8_107_1256_0, i_8_107_1264_0, i_8_107_1283_0, i_8_107_1292_0,
    i_8_107_1310_0, i_8_107_1404_0, i_8_107_1547_0, i_8_107_1588_0,
    i_8_107_1607_0, i_8_107_1628_0, i_8_107_1652_0, i_8_107_1673_0,
    i_8_107_1681_0, i_8_107_1706_0, i_8_107_1733_0, i_8_107_1763_0,
    i_8_107_1777_0, i_8_107_1819_0, i_8_107_1823_0, i_8_107_1825_0,
    i_8_107_1826_0, i_8_107_1858_0, i_8_107_1889_0, i_8_107_1940_0,
    i_8_107_1996_0, i_8_107_2003_0, i_8_107_2072_0, i_8_107_2108_0,
    i_8_107_2111_0, i_8_107_2134_0, i_8_107_2147_0, i_8_107_2149_0,
    i_8_107_2153_0, i_8_107_2156_0, i_8_107_2173_0, i_8_107_2180_0,
    i_8_107_2192_0, i_8_107_2200_0, i_8_107_2201_0, i_8_107_2225_0,
    i_8_107_2244_0, i_8_107_2273_0, i_8_107_2294_0,
    o_8_107_0_0  );
  input  i_8_107_31_0, i_8_107_50_0, i_8_107_86_0, i_8_107_167_0,
    i_8_107_230_0, i_8_107_233_0, i_8_107_234_0, i_8_107_326_0,
    i_8_107_335_0, i_8_107_338_0, i_8_107_365_0, i_8_107_368_0,
    i_8_107_380_0, i_8_107_386_0, i_8_107_400_0, i_8_107_419_0,
    i_8_107_424_0, i_8_107_425_0, i_8_107_428_0, i_8_107_440_0,
    i_8_107_449_0, i_8_107_451_0, i_8_107_452_0, i_8_107_494_0,
    i_8_107_499_0, i_8_107_500_0, i_8_107_581_0, i_8_107_613_0,
    i_8_107_614_0, i_8_107_617_0, i_8_107_655_0, i_8_107_694_0,
    i_8_107_698_0, i_8_107_706_0, i_8_107_707_0, i_8_107_733_0,
    i_8_107_767_0, i_8_107_770_0, i_8_107_796_0, i_8_107_797_0,
    i_8_107_839_0, i_8_107_842_0, i_8_107_845_0, i_8_107_878_0,
    i_8_107_932_0, i_8_107_956_0, i_8_107_968_0, i_8_107_1019_0,
    i_8_107_1022_0, i_8_107_1058_0, i_8_107_1097_0, i_8_107_1106_0,
    i_8_107_1157_0, i_8_107_1229_0, i_8_107_1235_0, i_8_107_1238_0,
    i_8_107_1253_0, i_8_107_1256_0, i_8_107_1264_0, i_8_107_1283_0,
    i_8_107_1292_0, i_8_107_1310_0, i_8_107_1404_0, i_8_107_1547_0,
    i_8_107_1588_0, i_8_107_1607_0, i_8_107_1628_0, i_8_107_1652_0,
    i_8_107_1673_0, i_8_107_1681_0, i_8_107_1706_0, i_8_107_1733_0,
    i_8_107_1763_0, i_8_107_1777_0, i_8_107_1819_0, i_8_107_1823_0,
    i_8_107_1825_0, i_8_107_1826_0, i_8_107_1858_0, i_8_107_1889_0,
    i_8_107_1940_0, i_8_107_1996_0, i_8_107_2003_0, i_8_107_2072_0,
    i_8_107_2108_0, i_8_107_2111_0, i_8_107_2134_0, i_8_107_2147_0,
    i_8_107_2149_0, i_8_107_2153_0, i_8_107_2156_0, i_8_107_2173_0,
    i_8_107_2180_0, i_8_107_2192_0, i_8_107_2200_0, i_8_107_2201_0,
    i_8_107_2225_0, i_8_107_2244_0, i_8_107_2273_0, i_8_107_2294_0;
  output o_8_107_0_0;
  assign o_8_107_0_0 = 0;
endmodule



// Benchmark "kernel_8_108" written by ABC on Sun Jul 19 10:04:52 2020

module kernel_8_108 ( 
    i_8_108_138_0, i_8_108_163_0, i_8_108_175_0, i_8_108_211_0,
    i_8_108_241_0, i_8_108_262_0, i_8_108_306_0, i_8_108_309_0,
    i_8_108_349_0, i_8_108_363_0, i_8_108_390_0, i_8_108_444_0,
    i_8_108_462_0, i_8_108_492_0, i_8_108_493_0, i_8_108_499_0,
    i_8_108_501_0, i_8_108_504_0, i_8_108_505_0, i_8_108_524_0,
    i_8_108_525_0, i_8_108_528_0, i_8_108_586_0, i_8_108_643_0,
    i_8_108_697_0, i_8_108_701_0, i_8_108_707_0, i_8_108_709_0,
    i_8_108_714_0, i_8_108_750_0, i_8_108_751_0, i_8_108_780_0,
    i_8_108_813_0, i_8_108_842_0, i_8_108_880_0, i_8_108_895_0,
    i_8_108_964_0, i_8_108_996_0, i_8_108_1013_0, i_8_108_1035_0,
    i_8_108_1040_0, i_8_108_1047_0, i_8_108_1071_0, i_8_108_1074_0,
    i_8_108_1084_0, i_8_108_1110_0, i_8_108_1113_0, i_8_108_1132_0,
    i_8_108_1157_0, i_8_108_1267_0, i_8_108_1303_0, i_8_108_1317_0,
    i_8_108_1326_0, i_8_108_1383_0, i_8_108_1401_0, i_8_108_1409_0,
    i_8_108_1422_0, i_8_108_1423_0, i_8_108_1443_0, i_8_108_1462_0,
    i_8_108_1465_0, i_8_108_1506_0, i_8_108_1507_0, i_8_108_1519_0,
    i_8_108_1533_0, i_8_108_1547_0, i_8_108_1548_0, i_8_108_1552_0,
    i_8_108_1553_0, i_8_108_1603_0, i_8_108_1623_0, i_8_108_1638_0,
    i_8_108_1672_0, i_8_108_1674_0, i_8_108_1683_0, i_8_108_1693_0,
    i_8_108_1701_0, i_8_108_1773_0, i_8_108_1775_0, i_8_108_1783_0,
    i_8_108_1832_0, i_8_108_1839_0, i_8_108_1840_0, i_8_108_1881_0,
    i_8_108_1882_0, i_8_108_1883_0, i_8_108_1885_0, i_8_108_1886_0,
    i_8_108_1888_0, i_8_108_1894_0, i_8_108_1900_0, i_8_108_1957_0,
    i_8_108_1984_0, i_8_108_2075_0, i_8_108_2088_0, i_8_108_2109_0,
    i_8_108_2148_0, i_8_108_2156_0, i_8_108_2173_0, i_8_108_2197_0,
    o_8_108_0_0  );
  input  i_8_108_138_0, i_8_108_163_0, i_8_108_175_0, i_8_108_211_0,
    i_8_108_241_0, i_8_108_262_0, i_8_108_306_0, i_8_108_309_0,
    i_8_108_349_0, i_8_108_363_0, i_8_108_390_0, i_8_108_444_0,
    i_8_108_462_0, i_8_108_492_0, i_8_108_493_0, i_8_108_499_0,
    i_8_108_501_0, i_8_108_504_0, i_8_108_505_0, i_8_108_524_0,
    i_8_108_525_0, i_8_108_528_0, i_8_108_586_0, i_8_108_643_0,
    i_8_108_697_0, i_8_108_701_0, i_8_108_707_0, i_8_108_709_0,
    i_8_108_714_0, i_8_108_750_0, i_8_108_751_0, i_8_108_780_0,
    i_8_108_813_0, i_8_108_842_0, i_8_108_880_0, i_8_108_895_0,
    i_8_108_964_0, i_8_108_996_0, i_8_108_1013_0, i_8_108_1035_0,
    i_8_108_1040_0, i_8_108_1047_0, i_8_108_1071_0, i_8_108_1074_0,
    i_8_108_1084_0, i_8_108_1110_0, i_8_108_1113_0, i_8_108_1132_0,
    i_8_108_1157_0, i_8_108_1267_0, i_8_108_1303_0, i_8_108_1317_0,
    i_8_108_1326_0, i_8_108_1383_0, i_8_108_1401_0, i_8_108_1409_0,
    i_8_108_1422_0, i_8_108_1423_0, i_8_108_1443_0, i_8_108_1462_0,
    i_8_108_1465_0, i_8_108_1506_0, i_8_108_1507_0, i_8_108_1519_0,
    i_8_108_1533_0, i_8_108_1547_0, i_8_108_1548_0, i_8_108_1552_0,
    i_8_108_1553_0, i_8_108_1603_0, i_8_108_1623_0, i_8_108_1638_0,
    i_8_108_1672_0, i_8_108_1674_0, i_8_108_1683_0, i_8_108_1693_0,
    i_8_108_1701_0, i_8_108_1773_0, i_8_108_1775_0, i_8_108_1783_0,
    i_8_108_1832_0, i_8_108_1839_0, i_8_108_1840_0, i_8_108_1881_0,
    i_8_108_1882_0, i_8_108_1883_0, i_8_108_1885_0, i_8_108_1886_0,
    i_8_108_1888_0, i_8_108_1894_0, i_8_108_1900_0, i_8_108_1957_0,
    i_8_108_1984_0, i_8_108_2075_0, i_8_108_2088_0, i_8_108_2109_0,
    i_8_108_2148_0, i_8_108_2156_0, i_8_108_2173_0, i_8_108_2197_0;
  output o_8_108_0_0;
  assign o_8_108_0_0 = 0;
endmodule



// Benchmark "kernel_8_109" written by ABC on Sun Jul 19 10:04:54 2020

module kernel_8_109 ( 
    i_8_109_51_0, i_8_109_77_0, i_8_109_194_0, i_8_109_220_0,
    i_8_109_221_0, i_8_109_223_0, i_8_109_224_0, i_8_109_225_0,
    i_8_109_234_0, i_8_109_235_0, i_8_109_236_0, i_8_109_237_0,
    i_8_109_239_0, i_8_109_273_0, i_8_109_303_0, i_8_109_325_0,
    i_8_109_326_0, i_8_109_329_0, i_8_109_334_0, i_8_109_336_0,
    i_8_109_337_0, i_8_109_338_0, i_8_109_365_0, i_8_109_391_0,
    i_8_109_414_0, i_8_109_415_0, i_8_109_418_0, i_8_109_419_0,
    i_8_109_596_0, i_8_109_613_0, i_8_109_614_0, i_8_109_648_0,
    i_8_109_649_0, i_8_109_650_0, i_8_109_651_0, i_8_109_652_0,
    i_8_109_715_0, i_8_109_748_0, i_8_109_749_0, i_8_109_764_0,
    i_8_109_838_0, i_8_109_848_0, i_8_109_970_0, i_8_109_1032_0,
    i_8_109_1048_0, i_8_109_1050_0, i_8_109_1278_0, i_8_109_1287_0,
    i_8_109_1290_0, i_8_109_1291_0, i_8_109_1292_0, i_8_109_1303_0,
    i_8_109_1353_0, i_8_109_1355_0, i_8_109_1439_0, i_8_109_1545_0,
    i_8_109_1546_0, i_8_109_1547_0, i_8_109_1630_0, i_8_109_1631_0,
    i_8_109_1635_0, i_8_109_1675_0, i_8_109_1746_0, i_8_109_1759_0,
    i_8_109_1764_0, i_8_109_1767_0, i_8_109_1769_0, i_8_109_1773_0,
    i_8_109_1774_0, i_8_109_1775_0, i_8_109_1778_0, i_8_109_1808_0,
    i_8_109_1818_0, i_8_109_1819_0, i_8_109_1820_0, i_8_109_1827_0,
    i_8_109_1828_0, i_8_109_1829_0, i_8_109_1830_0, i_8_109_1831_0,
    i_8_109_1859_0, i_8_109_1883_0, i_8_109_1924_0, i_8_109_1949_0,
    i_8_109_1990_0, i_8_109_1992_0, i_8_109_1993_0, i_8_109_1994_0,
    i_8_109_2016_0, i_8_109_2017_0, i_8_109_2019_0, i_8_109_2028_0,
    i_8_109_2088_0, i_8_109_2133_0, i_8_109_2134_0, i_8_109_2152_0,
    i_8_109_2208_0, i_8_109_2209_0, i_8_109_2223_0, i_8_109_2290_0,
    o_8_109_0_0  );
  input  i_8_109_51_0, i_8_109_77_0, i_8_109_194_0, i_8_109_220_0,
    i_8_109_221_0, i_8_109_223_0, i_8_109_224_0, i_8_109_225_0,
    i_8_109_234_0, i_8_109_235_0, i_8_109_236_0, i_8_109_237_0,
    i_8_109_239_0, i_8_109_273_0, i_8_109_303_0, i_8_109_325_0,
    i_8_109_326_0, i_8_109_329_0, i_8_109_334_0, i_8_109_336_0,
    i_8_109_337_0, i_8_109_338_0, i_8_109_365_0, i_8_109_391_0,
    i_8_109_414_0, i_8_109_415_0, i_8_109_418_0, i_8_109_419_0,
    i_8_109_596_0, i_8_109_613_0, i_8_109_614_0, i_8_109_648_0,
    i_8_109_649_0, i_8_109_650_0, i_8_109_651_0, i_8_109_652_0,
    i_8_109_715_0, i_8_109_748_0, i_8_109_749_0, i_8_109_764_0,
    i_8_109_838_0, i_8_109_848_0, i_8_109_970_0, i_8_109_1032_0,
    i_8_109_1048_0, i_8_109_1050_0, i_8_109_1278_0, i_8_109_1287_0,
    i_8_109_1290_0, i_8_109_1291_0, i_8_109_1292_0, i_8_109_1303_0,
    i_8_109_1353_0, i_8_109_1355_0, i_8_109_1439_0, i_8_109_1545_0,
    i_8_109_1546_0, i_8_109_1547_0, i_8_109_1630_0, i_8_109_1631_0,
    i_8_109_1635_0, i_8_109_1675_0, i_8_109_1746_0, i_8_109_1759_0,
    i_8_109_1764_0, i_8_109_1767_0, i_8_109_1769_0, i_8_109_1773_0,
    i_8_109_1774_0, i_8_109_1775_0, i_8_109_1778_0, i_8_109_1808_0,
    i_8_109_1818_0, i_8_109_1819_0, i_8_109_1820_0, i_8_109_1827_0,
    i_8_109_1828_0, i_8_109_1829_0, i_8_109_1830_0, i_8_109_1831_0,
    i_8_109_1859_0, i_8_109_1883_0, i_8_109_1924_0, i_8_109_1949_0,
    i_8_109_1990_0, i_8_109_1992_0, i_8_109_1993_0, i_8_109_1994_0,
    i_8_109_2016_0, i_8_109_2017_0, i_8_109_2019_0, i_8_109_2028_0,
    i_8_109_2088_0, i_8_109_2133_0, i_8_109_2134_0, i_8_109_2152_0,
    i_8_109_2208_0, i_8_109_2209_0, i_8_109_2223_0, i_8_109_2290_0;
  output o_8_109_0_0;
  assign o_8_109_0_0 = ~((~i_8_109_1547_0 & ((~i_8_109_414_0 & ((~i_8_109_220_0 & ~i_8_109_2088_0 & ((~i_8_109_365_0 & ~i_8_109_391_0 & ~i_8_109_418_0 & ~i_8_109_419_0 & ~i_8_109_652_0 & ~i_8_109_970_0 & ~i_8_109_1355_0 & ~i_8_109_1545_0 & ~i_8_109_1746_0 & ~i_8_109_1775_0 & ~i_8_109_1990_0 & ~i_8_109_1992_0) | (~i_8_109_223_0 & ~i_8_109_224_0 & ~i_8_109_225_0 & ~i_8_109_325_0 & ~i_8_109_326_0 & ~i_8_109_649_0 & ~i_8_109_1032_0 & ~i_8_109_1546_0 & ~i_8_109_1767_0 & ~i_8_109_1769_0 & ~i_8_109_1818_0 & ~i_8_109_1994_0 & ~i_8_109_2223_0))) | (~i_8_109_224_0 & ~i_8_109_329_0 & ~i_8_109_418_0 & ~i_8_109_419_0 & ~i_8_109_649_0 & ~i_8_109_652_0 & ~i_8_109_715_0 & ~i_8_109_749_0 & ~i_8_109_848_0 & ~i_8_109_1353_0 & ~i_8_109_1546_0 & ~i_8_109_1630_0 & ~i_8_109_1820_0 & ~i_8_109_1992_0 & ~i_8_109_1993_0))) | (~i_8_109_418_0 & ((~i_8_109_649_0 & ((~i_8_109_224_0 & ~i_8_109_652_0 & ~i_8_109_1355_0 & ((~i_8_109_223_0 & i_8_109_239_0 & ~i_8_109_1287_0 & ~i_8_109_1775_0) | (~i_8_109_221_0 & ~i_8_109_225_0 & ~i_8_109_303_0 & ~i_8_109_325_0 & ~i_8_109_596_0 & ~i_8_109_648_0 & ~i_8_109_749_0 & ~i_8_109_1050_0 & ~i_8_109_1546_0 & ~i_8_109_1773_0 & ~i_8_109_1949_0 & ~i_8_109_1993_0))) | (~i_8_109_273_0 & ~i_8_109_325_0 & ~i_8_109_419_0 & ~i_8_109_651_0 & ~i_8_109_970_0 & i_8_109_1759_0 & ~i_8_109_1924_0 & ~i_8_109_1990_0))) | (~i_8_109_77_0 & ~i_8_109_273_0 & ~i_8_109_326_0 & ~i_8_109_648_0 & ~i_8_109_970_0 & ~i_8_109_1355_0 & ~i_8_109_1630_0 & ~i_8_109_1773_0 & i_8_109_1808_0) | (~i_8_109_325_0 & ~i_8_109_329_0 & ~i_8_109_596_0 & ~i_8_109_749_0 & ~i_8_109_1278_0 & ~i_8_109_1353_0 & i_8_109_1439_0 & ~i_8_109_1759_0 & ~i_8_109_1775_0 & ~i_8_109_2152_0))) | (~i_8_109_748_0 & ((~i_8_109_1994_0 & ((i_8_109_337_0 & ~i_8_109_419_0 & ~i_8_109_764_0 & ~i_8_109_838_0 & ~i_8_109_1032_0 & i_8_109_1831_0 & ~i_8_109_2152_0) | (~i_8_109_51_0 & ~i_8_109_239_0 & i_8_109_336_0 & ~i_8_109_1546_0 & ~i_8_109_1630_0 & ~i_8_109_1769_0 & ~i_8_109_1992_0 & ~i_8_109_2223_0))) | (i_8_109_223_0 & ~i_8_109_273_0 & i_8_109_1032_0 & ~i_8_109_1048_0 & ~i_8_109_1545_0 & ~i_8_109_1675_0 & ~i_8_109_1774_0 & ~i_8_109_1949_0 & ~i_8_109_2134_0))))) | (~i_8_109_1764_0 & ((~i_8_109_223_0 & ((~i_8_109_224_0 & ~i_8_109_325_0 & ~i_8_109_391_0 & ~i_8_109_648_0 & ~i_8_109_650_0 & ~i_8_109_1050_0 & i_8_109_1278_0 & ~i_8_109_1631_0 & ~i_8_109_1808_0 & ~i_8_109_2088_0 & ~i_8_109_2133_0) | (~i_8_109_77_0 & ~i_8_109_651_0 & i_8_109_1545_0 & i_8_109_2152_0))) | (i_8_109_236_0 & ((~i_8_109_225_0 & ~i_8_109_239_0 & ~i_8_109_326_0 & ~i_8_109_419_0 & ~i_8_109_648_0 & ~i_8_109_650_0 & ~i_8_109_749_0 & ~i_8_109_1303_0 & ~i_8_109_1545_0) | (i_8_109_334_0 & ~i_8_109_418_0 & ~i_8_109_1032_0 & ~i_8_109_1769_0 & ~i_8_109_1773_0 & i_8_109_1775_0))) | (~i_8_109_419_0 & ~i_8_109_749_0 & ~i_8_109_848_0 & ~i_8_109_1291_0 & i_8_109_1303_0 & ~i_8_109_1769_0 & ~i_8_109_1819_0 & ~i_8_109_1990_0 & ~i_8_109_1993_0 & ~i_8_109_2028_0 & ~i_8_109_2223_0))) | (~i_8_109_1767_0 & ((~i_8_109_224_0 & ((~i_8_109_1994_0 & ((~i_8_109_329_0 & ((~i_8_109_51_0 & ~i_8_109_418_0 & ~i_8_109_1819_0 & ~i_8_109_1990_0 & ~i_8_109_2088_0 & ((~i_8_109_415_0 & ~i_8_109_419_0 & ~i_8_109_614_0 & ~i_8_109_1303_0 & ~i_8_109_1353_0 & ~i_8_109_1859_0 & ~i_8_109_1949_0 & ~i_8_109_1992_0 & ~i_8_109_2028_0) | (~i_8_109_303_0 & ~i_8_109_596_0 & ~i_8_109_648_0 & ~i_8_109_748_0 & ~i_8_109_848_0 & ~i_8_109_1355_0 & ~i_8_109_1545_0 & ~i_8_109_1635_0 & ~i_8_109_1769_0 & ~i_8_109_1820_0 & ~i_8_109_1993_0 & ~i_8_109_2223_0))) | (~i_8_109_77_0 & ~i_8_109_223_0 & ~i_8_109_391_0 & ~i_8_109_414_0 & ~i_8_109_596_0 & ~i_8_109_650_0 & ~i_8_109_651_0 & ~i_8_109_1546_0 & ~i_8_109_1630_0 & ~i_8_109_1635_0 & ~i_8_109_1746_0 & ~i_8_109_1759_0 & ~i_8_109_1775_0 & ~i_8_109_2028_0))) | (~i_8_109_194_0 & ~i_8_109_273_0 & ~i_8_109_414_0 & ~i_8_109_418_0 & ~i_8_109_650_0 & ~i_8_109_764_0 & ~i_8_109_970_0 & ~i_8_109_1630_0 & ~i_8_109_1775_0 & ~i_8_109_1808_0 & ~i_8_109_1818_0 & ~i_8_109_1820_0 & ~i_8_109_1992_0 & ~i_8_109_1993_0 & ~i_8_109_2028_0 & ~i_8_109_2133_0 & ~i_8_109_2134_0))) | (~i_8_109_419_0 & ~i_8_109_838_0 & ~i_8_109_1546_0 & ~i_8_109_1746_0 & ~i_8_109_1774_0 & ~i_8_109_1775_0 & ~i_8_109_1992_0 & ~i_8_109_2133_0 & i_8_109_2290_0))) | (i_8_109_338_0 & ((i_8_109_329_0 & ~i_8_109_749_0 & ~i_8_109_1353_0 & ~i_8_109_1546_0 & ~i_8_109_1631_0 & ~i_8_109_1635_0 & ~i_8_109_1808_0) | (~i_8_109_325_0 & ~i_8_109_648_0 & ~i_8_109_764_0 & ~i_8_109_1032_0 & ~i_8_109_1355_0 & ~i_8_109_1769_0 & ~i_8_109_1990_0 & ~i_8_109_1994_0))) | (~i_8_109_848_0 & ((~i_8_109_325_0 & ~i_8_109_391_0 & ~i_8_109_1032_0 & ((~i_8_109_329_0 & ~i_8_109_715_0 & ~i_8_109_1050_0 & i_8_109_1303_0 & ~i_8_109_1631_0 & ~i_8_109_1746_0 & ~i_8_109_1949_0) | (i_8_109_51_0 & ~i_8_109_415_0 & ~i_8_109_419_0 & ~i_8_109_748_0 & ~i_8_109_1545_0 & ~i_8_109_1759_0 & ~i_8_109_2017_0 & ~i_8_109_2223_0))) | (~i_8_109_596_0 & ~i_8_109_648_0 & ~i_8_109_77_0 & ~i_8_109_419_0 & ~i_8_109_652_0 & ~i_8_109_749_0 & ~i_8_109_970_0 & ~i_8_109_1050_0 & ~i_8_109_1545_0 & ~i_8_109_1631_0 & ~i_8_109_1769_0 & ~i_8_109_1774_0 & ~i_8_109_1778_0 & ~i_8_109_1808_0 & ~i_8_109_1993_0 & ~i_8_109_2088_0))) | (i_8_109_194_0 & ~i_8_109_419_0 & i_8_109_1355_0 & i_8_109_1759_0 & ~i_8_109_1769_0 & i_8_109_1808_0) | (~i_8_109_748_0 & ~i_8_109_1631_0 & i_8_109_1830_0 & ~i_8_109_1992_0 & ~i_8_109_2028_0 & ~i_8_109_2133_0))) | (~i_8_109_2088_0 & ((~i_8_109_51_0 & ((~i_8_109_338_0 & ~i_8_109_391_0 & i_8_109_1290_0 & ~i_8_109_1439_0 & ~i_8_109_1990_0 & ~i_8_109_2152_0) | (~i_8_109_329_0 & ~i_8_109_415_0 & ~i_8_109_652_0 & ~i_8_109_715_0 & ~i_8_109_749_0 & ~i_8_109_848_0 & ~i_8_109_1746_0 & ~i_8_109_1992_0 & i_8_109_1993_0 & ~i_8_109_1994_0 & ~i_8_109_2290_0))) | (~i_8_109_303_0 & ~i_8_109_325_0 & ~i_8_109_329_0 & i_8_109_338_0 & ~i_8_109_419_0 & ~i_8_109_649_0 & ~i_8_109_748_0 & ~i_8_109_1546_0 & ~i_8_109_1774_0 & ~i_8_109_1819_0 & ~i_8_109_1990_0) | (~i_8_109_221_0 & ~i_8_109_326_0 & ~i_8_109_648_0 & ~i_8_109_650_0 & ~i_8_109_652_0 & ~i_8_109_1032_0 & ~i_8_109_1355_0 & ~i_8_109_1630_0 & ~i_8_109_2028_0 & ~i_8_109_2134_0 & i_8_109_2152_0 & ~i_8_109_2208_0))) | (~i_8_109_1355_0 & ((~i_8_109_194_0 & ~i_8_109_749_0 & ((~i_8_109_225_0 & ~i_8_109_650_0 & ~i_8_109_652_0 & ~i_8_109_1048_0 & ~i_8_109_1546_0 & i_8_109_1635_0 & ~i_8_109_1746_0 & ~i_8_109_1994_0) | (i_8_109_224_0 & ~i_8_109_273_0 & ~i_8_109_1278_0 & ~i_8_109_1545_0 & ~i_8_109_1631_0 & ~i_8_109_1759_0 & ~i_8_109_1769_0 & i_8_109_1808_0 & ~i_8_109_1883_0 & ~i_8_109_1993_0 & ~i_8_109_2152_0))) | (~i_8_109_651_0 & ((~i_8_109_225_0 & ((i_8_109_239_0 & ~i_8_109_329_0 & ~i_8_109_414_0 & ~i_8_109_648_0 & i_8_109_1439_0 & ~i_8_109_1808_0) | (~i_8_109_303_0 & ~i_8_109_419_0 & ~i_8_109_748_0 & ~i_8_109_1769_0 & ~i_8_109_1774_0 & ~i_8_109_848_0 & ~i_8_109_970_0 & ~i_8_109_1775_0 & ~i_8_109_1819_0 & i_8_109_1924_0 & ~i_8_109_1949_0 & ~i_8_109_1990_0 & ~i_8_109_1994_0 & ~i_8_109_2134_0))) | (~i_8_109_596_0 & ~i_8_109_764_0 & ((~i_8_109_336_0 & ~i_8_109_365_0 & ~i_8_109_1774_0 & ~i_8_109_1775_0 & ~i_8_109_1818_0 & ~i_8_109_1924_0 & i_8_109_2152_0) | (i_8_109_235_0 & ~i_8_109_970_0 & ~i_8_109_1808_0 & ~i_8_109_1819_0 & ~i_8_109_1992_0 & ~i_8_109_2028_0 & ~i_8_109_2152_0))))) | (~i_8_109_273_0 & ~i_8_109_303_0 & ~i_8_109_326_0 & ~i_8_109_329_0 & ~i_8_109_414_0 & ~i_8_109_415_0 & ~i_8_109_419_0 & ~i_8_109_648_0 & ~i_8_109_649_0 & ~i_8_109_838_0 & ~i_8_109_1303_0 & ~i_8_109_1353_0 & ~i_8_109_1545_0 & ~i_8_109_1808_0 & ~i_8_109_1993_0 & ~i_8_109_1994_0 & ~i_8_109_2223_0))) | (~i_8_109_326_0 & ~i_8_109_419_0 & ~i_8_109_749_0 & ~i_8_109_1050_0 & ~i_8_109_1545_0 & ~i_8_109_1630_0 & ((i_8_109_336_0 & ~i_8_109_414_0 & ~i_8_109_648_0 & ~i_8_109_650_0 & ~i_8_109_2133_0) | (~i_8_109_194_0 & ~i_8_109_224_0 & ~i_8_109_239_0 & ~i_8_109_303_0 & ~i_8_109_325_0 & ~i_8_109_329_0 & ~i_8_109_365_0 & ~i_8_109_418_0 & ~i_8_109_748_0 & ~i_8_109_1818_0 & ~i_8_109_1949_0 & ~i_8_109_1992_0 & ~i_8_109_2134_0))) | (i_8_109_337_0 & ~i_8_109_596_0 & ~i_8_109_648_0 & ~i_8_109_651_0 & ~i_8_109_652_0 & ~i_8_109_848_0 & i_8_109_1675_0 & ~i_8_109_1769_0 & ~i_8_109_1819_0 & ~i_8_109_1831_0) | (~i_8_109_1818_0 & i_8_109_1819_0 & i_8_109_1859_0 & ~i_8_109_1990_0 & ~i_8_109_2134_0 & i_8_109_2290_0));
endmodule



// Benchmark "kernel_8_110" written by ABC on Sun Jul 19 10:04:55 2020

module kernel_8_110 ( 
    i_8_110_0_0, i_8_110_19_0, i_8_110_20_0, i_8_110_36_0, i_8_110_46_0,
    i_8_110_47_0, i_8_110_100_0, i_8_110_111_0, i_8_110_136_0,
    i_8_110_189_0, i_8_110_347_0, i_8_110_379_0, i_8_110_398_0,
    i_8_110_425_0, i_8_110_487_0, i_8_110_496_0, i_8_110_527_0,
    i_8_110_595_0, i_8_110_607_0, i_8_110_633_0, i_8_110_634_0,
    i_8_110_709_0, i_8_110_766_0, i_8_110_767_0, i_8_110_838_0,
    i_8_110_874_0, i_8_110_879_0, i_8_110_884_0, i_8_110_919_0,
    i_8_110_922_0, i_8_110_966_0, i_8_110_968_0, i_8_110_991_0,
    i_8_110_992_0, i_8_110_1026_0, i_8_110_1036_0, i_8_110_1073_0,
    i_8_110_1135_0, i_8_110_1154_0, i_8_110_1180_0, i_8_110_1225_0,
    i_8_110_1226_0, i_8_110_1252_0, i_8_110_1253_0, i_8_110_1263_0,
    i_8_110_1265_0, i_8_110_1270_0, i_8_110_1279_0, i_8_110_1280_0,
    i_8_110_1399_0, i_8_110_1453_0, i_8_110_1468_0, i_8_110_1478_0,
    i_8_110_1486_0, i_8_110_1487_0, i_8_110_1493_0, i_8_110_1534_0,
    i_8_110_1558_0, i_8_110_1559_0, i_8_110_1603_0, i_8_110_1604_0,
    i_8_110_1634_0, i_8_110_1648_0, i_8_110_1649_0, i_8_110_1681_0,
    i_8_110_1710_0, i_8_110_1719_0, i_8_110_1746_0, i_8_110_1747_0,
    i_8_110_1748_0, i_8_110_1764_0, i_8_110_1768_0, i_8_110_1771_0,
    i_8_110_1779_0, i_8_110_1792_0, i_8_110_1803_0, i_8_110_1832_0,
    i_8_110_1882_0, i_8_110_1884_0, i_8_110_1886_0, i_8_110_1944_0,
    i_8_110_1946_0, i_8_110_1981_0, i_8_110_1991_0, i_8_110_1994_0,
    i_8_110_2008_0, i_8_110_2017_0, i_8_110_2054_0, i_8_110_2090_0,
    i_8_110_2106_0, i_8_110_2107_0, i_8_110_2108_0, i_8_110_2147_0,
    i_8_110_2153_0, i_8_110_2224_0, i_8_110_2242_0, i_8_110_2245_0,
    i_8_110_2270_0, i_8_110_2287_0, i_8_110_2288_0,
    o_8_110_0_0  );
  input  i_8_110_0_0, i_8_110_19_0, i_8_110_20_0, i_8_110_36_0,
    i_8_110_46_0, i_8_110_47_0, i_8_110_100_0, i_8_110_111_0,
    i_8_110_136_0, i_8_110_189_0, i_8_110_347_0, i_8_110_379_0,
    i_8_110_398_0, i_8_110_425_0, i_8_110_487_0, i_8_110_496_0,
    i_8_110_527_0, i_8_110_595_0, i_8_110_607_0, i_8_110_633_0,
    i_8_110_634_0, i_8_110_709_0, i_8_110_766_0, i_8_110_767_0,
    i_8_110_838_0, i_8_110_874_0, i_8_110_879_0, i_8_110_884_0,
    i_8_110_919_0, i_8_110_922_0, i_8_110_966_0, i_8_110_968_0,
    i_8_110_991_0, i_8_110_992_0, i_8_110_1026_0, i_8_110_1036_0,
    i_8_110_1073_0, i_8_110_1135_0, i_8_110_1154_0, i_8_110_1180_0,
    i_8_110_1225_0, i_8_110_1226_0, i_8_110_1252_0, i_8_110_1253_0,
    i_8_110_1263_0, i_8_110_1265_0, i_8_110_1270_0, i_8_110_1279_0,
    i_8_110_1280_0, i_8_110_1399_0, i_8_110_1453_0, i_8_110_1468_0,
    i_8_110_1478_0, i_8_110_1486_0, i_8_110_1487_0, i_8_110_1493_0,
    i_8_110_1534_0, i_8_110_1558_0, i_8_110_1559_0, i_8_110_1603_0,
    i_8_110_1604_0, i_8_110_1634_0, i_8_110_1648_0, i_8_110_1649_0,
    i_8_110_1681_0, i_8_110_1710_0, i_8_110_1719_0, i_8_110_1746_0,
    i_8_110_1747_0, i_8_110_1748_0, i_8_110_1764_0, i_8_110_1768_0,
    i_8_110_1771_0, i_8_110_1779_0, i_8_110_1792_0, i_8_110_1803_0,
    i_8_110_1832_0, i_8_110_1882_0, i_8_110_1884_0, i_8_110_1886_0,
    i_8_110_1944_0, i_8_110_1946_0, i_8_110_1981_0, i_8_110_1991_0,
    i_8_110_1994_0, i_8_110_2008_0, i_8_110_2017_0, i_8_110_2054_0,
    i_8_110_2090_0, i_8_110_2106_0, i_8_110_2107_0, i_8_110_2108_0,
    i_8_110_2147_0, i_8_110_2153_0, i_8_110_2224_0, i_8_110_2242_0,
    i_8_110_2245_0, i_8_110_2270_0, i_8_110_2287_0, i_8_110_2288_0;
  output o_8_110_0_0;
  assign o_8_110_0_0 = ~((~i_8_110_36_0 & ((~i_8_110_379_0 & ~i_8_110_838_0 & ~i_8_110_922_0 & ~i_8_110_966_0 & ~i_8_110_1225_0 & ~i_8_110_1279_0 & ~i_8_110_2108_0) | (~i_8_110_19_0 & ~i_8_110_20_0 & ~i_8_110_398_0 & ~i_8_110_595_0 & ~i_8_110_874_0 & ~i_8_110_1604_0 & ~i_8_110_1944_0 & ~i_8_110_1981_0 & ~i_8_110_2017_0 & ~i_8_110_2287_0))) | (~i_8_110_19_0 & ((~i_8_110_767_0 & ~i_8_110_922_0 & ~i_8_110_1453_0 & ~i_8_110_1468_0 & ~i_8_110_1558_0 & i_8_110_1886_0) | (~i_8_110_47_0 & ~i_8_110_379_0 & ~i_8_110_496_0 & ~i_8_110_1226_0 & ~i_8_110_1710_0 & ~i_8_110_1981_0 & ~i_8_110_2107_0 & ~i_8_110_2147_0 & ~i_8_110_2245_0))) | (~i_8_110_111_0 & ((~i_8_110_767_0 & ((~i_8_110_20_0 & ((~i_8_110_398_0 & ~i_8_110_633_0 & ~i_8_110_966_0 & ~i_8_110_1026_0 & ~i_8_110_1399_0 & ~i_8_110_1648_0 & ~i_8_110_1747_0 & ~i_8_110_1764_0 & ~i_8_110_1946_0 & ~i_8_110_2017_0) | (~i_8_110_766_0 & ~i_8_110_879_0 & ~i_8_110_922_0 & ~i_8_110_1252_0 & ~i_8_110_1604_0 & ~i_8_110_1991_0 & ~i_8_110_2106_0 & ~i_8_110_2107_0 & ~i_8_110_2270_0 & ~i_8_110_2288_0))) | (~i_8_110_1225_0 & ~i_8_110_1468_0 & ~i_8_110_1534_0 & ~i_8_110_1558_0 & ~i_8_110_1559_0 & ~i_8_110_1603_0 & ~i_8_110_1604_0 & ~i_8_110_1944_0 & ~i_8_110_2017_0 & ~i_8_110_2287_0))) | (~i_8_110_46_0 & ~i_8_110_47_0 & ~i_8_110_425_0 & ~i_8_110_874_0 & ~i_8_110_966_0 & ~i_8_110_1225_0 & ~i_8_110_1486_0 & ~i_8_110_1558_0 & ~i_8_110_2106_0 & ~i_8_110_2107_0))) | (~i_8_110_2287_0 & ((~i_8_110_100_0 & ((~i_8_110_379_0 & ~i_8_110_1252_0 & ~i_8_110_1453_0 & ~i_8_110_1603_0 & ~i_8_110_1604_0 & ~i_8_110_2017_0 & ~i_8_110_2108_0) | (~i_8_110_398_0 & ~i_8_110_919_0 & ~i_8_110_1279_0 & ~i_8_110_1280_0 & ~i_8_110_1478_0 & ~i_8_110_2106_0 & ~i_8_110_2224_0))) | (~i_8_110_1558_0 & ((~i_8_110_398_0 & ~i_8_110_425_0 & ~i_8_110_595_0 & ~i_8_110_879_0 & ~i_8_110_1225_0 & ~i_8_110_1604_0 & ~i_8_110_2106_0 & ~i_8_110_2108_0) | (i_8_110_968_0 & ~i_8_110_991_0 & ~i_8_110_1263_0 & ~i_8_110_1603_0 & ~i_8_110_1710_0 & ~i_8_110_2242_0 & ~i_8_110_2270_0))) | (~i_8_110_1746_0 & ((~i_8_110_379_0 & ~i_8_110_1135_0 & ~i_8_110_1280_0 & ~i_8_110_1468_0 & ~i_8_110_1764_0 & ~i_8_110_2106_0) | (~i_8_110_1253_0 & ~i_8_110_1279_0 & i_8_110_2090_0 & i_8_110_2270_0))) | (~i_8_110_46_0 & ~i_8_110_487_0 & ~i_8_110_1886_0 & i_8_110_1981_0 & ~i_8_110_2107_0 & ~i_8_110_2153_0))) | (~i_8_110_46_0 & ((~i_8_110_47_0 & ~i_8_110_922_0 & ~i_8_110_991_0 & ~i_8_110_1453_0 & i_8_110_1648_0 & i_8_110_1747_0 & i_8_110_1882_0) | (~i_8_110_100_0 & ~i_8_110_398_0 & ~i_8_110_766_0 & ~i_8_110_1026_0 & ~i_8_110_1253_0 & ~i_8_110_1681_0 & ~i_8_110_1771_0 & ~i_8_110_1779_0 & ~i_8_110_2106_0 & ~i_8_110_2107_0 & ~i_8_110_2108_0))) | (~i_8_110_595_0 & ~i_8_110_634_0 & ((i_8_110_1135_0 & ~i_8_110_1253_0 & ~i_8_110_1263_0 & ~i_8_110_1468_0 & ~i_8_110_1558_0 & ~i_8_110_1559_0 & ~i_8_110_2224_0) | (i_8_110_111_0 & ~i_8_110_922_0 & i_8_110_966_0 & ~i_8_110_1270_0 & ~i_8_110_1280_0 & ~i_8_110_2017_0 & ~i_8_110_2288_0))) | (~i_8_110_919_0 & ((i_8_110_766_0 & i_8_110_767_0 & ~i_8_110_1225_0 & ~i_8_110_1280_0 & i_8_110_1534_0) | (~i_8_110_487_0 & ~i_8_110_879_0 & ~i_8_110_1252_0 & ~i_8_110_1399_0 & ~i_8_110_1603_0 & ~i_8_110_1604_0 & i_8_110_1746_0 & ~i_8_110_2017_0 & ~i_8_110_2054_0 & ~i_8_110_2107_0 & ~i_8_110_2245_0))) | (~i_8_110_879_0 & ((i_8_110_1036_0 & ~i_8_110_1180_0 & i_8_110_1453_0 & ~i_8_110_1944_0 & ~i_8_110_2242_0) | (i_8_110_1265_0 & ~i_8_110_1558_0 & i_8_110_1748_0 & ~i_8_110_2017_0 & ~i_8_110_2288_0 & i_8_110_1991_0 & i_8_110_1994_0))) | (~i_8_110_1036_0 & ((~i_8_110_1026_0 & ~i_8_110_1253_0 & i_8_110_1486_0 & ~i_8_110_1981_0 & ~i_8_110_2153_0) | (i_8_110_1534_0 & ~i_8_110_1768_0 & i_8_110_1994_0 & ~i_8_110_2054_0 & ~i_8_110_2242_0))) | (~i_8_110_1026_0 & ~i_8_110_1468_0 & ((i_8_110_1263_0 & ~i_8_110_1604_0 & ~i_8_110_1710_0 & i_8_110_1747_0 & ~i_8_110_1946_0 & ~i_8_110_2054_0) | (~i_8_110_922_0 & ~i_8_110_1225_0 & ~i_8_110_1280_0 & ~i_8_110_1558_0 & ~i_8_110_1746_0 & ~i_8_110_1981_0 & ~i_8_110_2017_0 & ~i_8_110_2224_0))) | (~i_8_110_1225_0 & ~i_8_110_1747_0 & ((~i_8_110_874_0 & ~i_8_110_1073_0 & ~i_8_110_1252_0 & ~i_8_110_1253_0 & ~i_8_110_1719_0 & ~i_8_110_1771_0 & ~i_8_110_1946_0 & ~i_8_110_2107_0) | (~i_8_110_100_0 & ~i_8_110_1226_0 & ~i_8_110_1270_0 & ~i_8_110_1558_0 & ~i_8_110_1603_0 & ~i_8_110_1746_0 & ~i_8_110_1944_0 & ~i_8_110_2224_0))) | (i_8_110_379_0 & i_8_110_634_0 & ~i_8_110_1135_0 & ~i_8_110_1226_0 & i_8_110_1263_0 & ~i_8_110_1603_0 & ~i_8_110_1748_0) | (i_8_110_607_0 & i_8_110_1073_0 & i_8_110_1779_0 & i_8_110_2090_0) | (i_8_110_0_0 & ~i_8_110_1252_0 & ~i_8_110_2106_0 & ~i_8_110_2153_0));
endmodule



// Benchmark "kernel_8_111" written by ABC on Sun Jul 19 10:04:56 2020

module kernel_8_111 ( 
    i_8_111_10_0, i_8_111_37_0, i_8_111_49_0, i_8_111_76_0, i_8_111_107_0,
    i_8_111_189_0, i_8_111_223_0, i_8_111_253_0, i_8_111_301_0,
    i_8_111_361_0, i_8_111_363_0, i_8_111_365_0, i_8_111_389_0,
    i_8_111_398_0, i_8_111_426_0, i_8_111_440_0, i_8_111_490_0,
    i_8_111_526_0, i_8_111_532_0, i_8_111_577_0, i_8_111_580_0,
    i_8_111_589_0, i_8_111_590_0, i_8_111_604_0, i_8_111_607_0,
    i_8_111_631_0, i_8_111_632_0, i_8_111_633_0, i_8_111_634_0,
    i_8_111_665_0, i_8_111_671_0, i_8_111_676_0, i_8_111_680_0,
    i_8_111_738_0, i_8_111_740_0, i_8_111_805_0, i_8_111_824_0,
    i_8_111_832_0, i_8_111_837_0, i_8_111_838_0, i_8_111_839_0,
    i_8_111_955_0, i_8_111_965_0, i_8_111_1037_0, i_8_111_1051_0,
    i_8_111_1099_0, i_8_111_1103_0, i_8_111_1127_0, i_8_111_1136_0,
    i_8_111_1152_0, i_8_111_1181_0, i_8_111_1237_0, i_8_111_1238_0,
    i_8_111_1261_0, i_8_111_1262_0, i_8_111_1315_0, i_8_111_1325_0,
    i_8_111_1328_0, i_8_111_1382_0, i_8_111_1398_0, i_8_111_1407_0,
    i_8_111_1414_0, i_8_111_1433_0, i_8_111_1434_0, i_8_111_1442_0,
    i_8_111_1463_0, i_8_111_1470_0, i_8_111_1472_0, i_8_111_1478_0,
    i_8_111_1506_0, i_8_111_1513_0, i_8_111_1550_0, i_8_111_1624_0,
    i_8_111_1629_0, i_8_111_1641_0, i_8_111_1702_0, i_8_111_1724_0,
    i_8_111_1768_0, i_8_111_1784_0, i_8_111_1804_0, i_8_111_1818_0,
    i_8_111_1820_0, i_8_111_1822_0, i_8_111_1837_0, i_8_111_1839_0,
    i_8_111_1903_0, i_8_111_1994_0, i_8_111_2008_0, i_8_111_2009_0,
    i_8_111_2011_0, i_8_111_2038_0, i_8_111_2071_0, i_8_111_2089_0,
    i_8_111_2098_0, i_8_111_2225_0, i_8_111_2227_0, i_8_111_2244_0,
    i_8_111_2245_0, i_8_111_2263_0, i_8_111_2296_0,
    o_8_111_0_0  );
  input  i_8_111_10_0, i_8_111_37_0, i_8_111_49_0, i_8_111_76_0,
    i_8_111_107_0, i_8_111_189_0, i_8_111_223_0, i_8_111_253_0,
    i_8_111_301_0, i_8_111_361_0, i_8_111_363_0, i_8_111_365_0,
    i_8_111_389_0, i_8_111_398_0, i_8_111_426_0, i_8_111_440_0,
    i_8_111_490_0, i_8_111_526_0, i_8_111_532_0, i_8_111_577_0,
    i_8_111_580_0, i_8_111_589_0, i_8_111_590_0, i_8_111_604_0,
    i_8_111_607_0, i_8_111_631_0, i_8_111_632_0, i_8_111_633_0,
    i_8_111_634_0, i_8_111_665_0, i_8_111_671_0, i_8_111_676_0,
    i_8_111_680_0, i_8_111_738_0, i_8_111_740_0, i_8_111_805_0,
    i_8_111_824_0, i_8_111_832_0, i_8_111_837_0, i_8_111_838_0,
    i_8_111_839_0, i_8_111_955_0, i_8_111_965_0, i_8_111_1037_0,
    i_8_111_1051_0, i_8_111_1099_0, i_8_111_1103_0, i_8_111_1127_0,
    i_8_111_1136_0, i_8_111_1152_0, i_8_111_1181_0, i_8_111_1237_0,
    i_8_111_1238_0, i_8_111_1261_0, i_8_111_1262_0, i_8_111_1315_0,
    i_8_111_1325_0, i_8_111_1328_0, i_8_111_1382_0, i_8_111_1398_0,
    i_8_111_1407_0, i_8_111_1414_0, i_8_111_1433_0, i_8_111_1434_0,
    i_8_111_1442_0, i_8_111_1463_0, i_8_111_1470_0, i_8_111_1472_0,
    i_8_111_1478_0, i_8_111_1506_0, i_8_111_1513_0, i_8_111_1550_0,
    i_8_111_1624_0, i_8_111_1629_0, i_8_111_1641_0, i_8_111_1702_0,
    i_8_111_1724_0, i_8_111_1768_0, i_8_111_1784_0, i_8_111_1804_0,
    i_8_111_1818_0, i_8_111_1820_0, i_8_111_1822_0, i_8_111_1837_0,
    i_8_111_1839_0, i_8_111_1903_0, i_8_111_1994_0, i_8_111_2008_0,
    i_8_111_2009_0, i_8_111_2011_0, i_8_111_2038_0, i_8_111_2071_0,
    i_8_111_2089_0, i_8_111_2098_0, i_8_111_2225_0, i_8_111_2227_0,
    i_8_111_2244_0, i_8_111_2245_0, i_8_111_2263_0, i_8_111_2296_0;
  output o_8_111_0_0;
  assign o_8_111_0_0 = 0;
endmodule



// Benchmark "kernel_8_112" written by ABC on Sun Jul 19 10:04:57 2020

module kernel_8_112 ( 
    i_8_112_14_0, i_8_112_45_0, i_8_112_46_0, i_8_112_66_0, i_8_112_82_0,
    i_8_112_136_0, i_8_112_163_0, i_8_112_172_0, i_8_112_193_0,
    i_8_112_207_0, i_8_112_238_0, i_8_112_253_0, i_8_112_255_0,
    i_8_112_307_0, i_8_112_342_0, i_8_112_345_0, i_8_112_375_0,
    i_8_112_423_0, i_8_112_424_0, i_8_112_470_0, i_8_112_481_0,
    i_8_112_495_0, i_8_112_526_0, i_8_112_527_0, i_8_112_544_0,
    i_8_112_549_0, i_8_112_568_0, i_8_112_586_0, i_8_112_603_0,
    i_8_112_613_0, i_8_112_630_0, i_8_112_664_0, i_8_112_676_0,
    i_8_112_765_0, i_8_112_828_0, i_8_112_883_0, i_8_112_918_0,
    i_8_112_927_0, i_8_112_973_0, i_8_112_997_0, i_8_112_998_0,
    i_8_112_1009_0, i_8_112_1017_0, i_8_112_1044_0, i_8_112_1045_0,
    i_8_112_1053_0, i_8_112_1221_0, i_8_112_1228_0, i_8_112_1233_0,
    i_8_112_1269_0, i_8_112_1271_0, i_8_112_1288_0, i_8_112_1296_0,
    i_8_112_1297_0, i_8_112_1306_0, i_8_112_1314_0, i_8_112_1323_0,
    i_8_112_1413_0, i_8_112_1434_0, i_8_112_1435_0, i_8_112_1512_0,
    i_8_112_1524_0, i_8_112_1536_0, i_8_112_1541_0, i_8_112_1558_0,
    i_8_112_1566_0, i_8_112_1611_0, i_8_112_1630_0, i_8_112_1642_0,
    i_8_112_1648_0, i_8_112_1650_0, i_8_112_1680_0, i_8_112_1681_0,
    i_8_112_1682_0, i_8_112_1683_0, i_8_112_1695_0, i_8_112_1707_0,
    i_8_112_1729_0, i_8_112_1763_0, i_8_112_1764_0, i_8_112_1803_0,
    i_8_112_1822_0, i_8_112_1855_0, i_8_112_1884_0, i_8_112_1885_0,
    i_8_112_1886_0, i_8_112_1902_0, i_8_112_1998_0, i_8_112_2106_0,
    i_8_112_2119_0, i_8_112_2142_0, i_8_112_2145_0, i_8_112_2152_0,
    i_8_112_2154_0, i_8_112_2187_0, i_8_112_2196_0, i_8_112_2205_0,
    i_8_112_2259_0, i_8_112_2260_0, i_8_112_2269_0,
    o_8_112_0_0  );
  input  i_8_112_14_0, i_8_112_45_0, i_8_112_46_0, i_8_112_66_0,
    i_8_112_82_0, i_8_112_136_0, i_8_112_163_0, i_8_112_172_0,
    i_8_112_193_0, i_8_112_207_0, i_8_112_238_0, i_8_112_253_0,
    i_8_112_255_0, i_8_112_307_0, i_8_112_342_0, i_8_112_345_0,
    i_8_112_375_0, i_8_112_423_0, i_8_112_424_0, i_8_112_470_0,
    i_8_112_481_0, i_8_112_495_0, i_8_112_526_0, i_8_112_527_0,
    i_8_112_544_0, i_8_112_549_0, i_8_112_568_0, i_8_112_586_0,
    i_8_112_603_0, i_8_112_613_0, i_8_112_630_0, i_8_112_664_0,
    i_8_112_676_0, i_8_112_765_0, i_8_112_828_0, i_8_112_883_0,
    i_8_112_918_0, i_8_112_927_0, i_8_112_973_0, i_8_112_997_0,
    i_8_112_998_0, i_8_112_1009_0, i_8_112_1017_0, i_8_112_1044_0,
    i_8_112_1045_0, i_8_112_1053_0, i_8_112_1221_0, i_8_112_1228_0,
    i_8_112_1233_0, i_8_112_1269_0, i_8_112_1271_0, i_8_112_1288_0,
    i_8_112_1296_0, i_8_112_1297_0, i_8_112_1306_0, i_8_112_1314_0,
    i_8_112_1323_0, i_8_112_1413_0, i_8_112_1434_0, i_8_112_1435_0,
    i_8_112_1512_0, i_8_112_1524_0, i_8_112_1536_0, i_8_112_1541_0,
    i_8_112_1558_0, i_8_112_1566_0, i_8_112_1611_0, i_8_112_1630_0,
    i_8_112_1642_0, i_8_112_1648_0, i_8_112_1650_0, i_8_112_1680_0,
    i_8_112_1681_0, i_8_112_1682_0, i_8_112_1683_0, i_8_112_1695_0,
    i_8_112_1707_0, i_8_112_1729_0, i_8_112_1763_0, i_8_112_1764_0,
    i_8_112_1803_0, i_8_112_1822_0, i_8_112_1855_0, i_8_112_1884_0,
    i_8_112_1885_0, i_8_112_1886_0, i_8_112_1902_0, i_8_112_1998_0,
    i_8_112_2106_0, i_8_112_2119_0, i_8_112_2142_0, i_8_112_2145_0,
    i_8_112_2152_0, i_8_112_2154_0, i_8_112_2187_0, i_8_112_2196_0,
    i_8_112_2205_0, i_8_112_2259_0, i_8_112_2260_0, i_8_112_2269_0;
  output o_8_112_0_0;
  assign o_8_112_0_0 = 0;
endmodule



// Benchmark "kernel_8_113" written by ABC on Sun Jul 19 10:04:58 2020

module kernel_8_113 ( 
    i_8_113_38_0, i_8_113_40_0, i_8_113_43_0, i_8_113_81_0, i_8_113_84_0,
    i_8_113_115_0, i_8_113_148_0, i_8_113_151_0, i_8_113_163_0,
    i_8_113_190_0, i_8_113_194_0, i_8_113_245_0, i_8_113_346_0,
    i_8_113_347_0, i_8_113_352_0, i_8_113_417_0, i_8_113_464_0,
    i_8_113_469_0, i_8_113_470_0, i_8_113_483_0, i_8_113_489_0,
    i_8_113_490_0, i_8_113_522_0, i_8_113_526_0, i_8_113_538_0,
    i_8_113_552_0, i_8_113_555_0, i_8_113_595_0, i_8_113_598_0,
    i_8_113_634_0, i_8_113_648_0, i_8_113_695_0, i_8_113_697_0,
    i_8_113_700_0, i_8_113_702_0, i_8_113_706_0, i_8_113_733_0,
    i_8_113_734_0, i_8_113_770_0, i_8_113_790_0, i_8_113_793_0,
    i_8_113_813_0, i_8_113_833_0, i_8_113_881_0, i_8_113_893_0,
    i_8_113_896_0, i_8_113_926_0, i_8_113_998_0, i_8_113_1154_0,
    i_8_113_1161_0, i_8_113_1171_0, i_8_113_1223_0, i_8_113_1233_0,
    i_8_113_1238_0, i_8_113_1262_0, i_8_113_1288_0, i_8_113_1289_0,
    i_8_113_1292_0, i_8_113_1299_0, i_8_113_1306_0, i_8_113_1309_0,
    i_8_113_1311_0, i_8_113_1312_0, i_8_113_1352_0, i_8_113_1381_0,
    i_8_113_1384_0, i_8_113_1423_0, i_8_113_1442_0, i_8_113_1491_0,
    i_8_113_1498_0, i_8_113_1543_0, i_8_113_1549_0, i_8_113_1562_0,
    i_8_113_1637_0, i_8_113_1648_0, i_8_113_1653_0, i_8_113_1687_0,
    i_8_113_1688_0, i_8_113_1690_0, i_8_113_1701_0, i_8_113_1708_0,
    i_8_113_1748_0, i_8_113_1750_0, i_8_113_1753_0, i_8_113_1803_0,
    i_8_113_1806_0, i_8_113_1832_0, i_8_113_1840_0, i_8_113_1926_0,
    i_8_113_1960_0, i_8_113_1996_0, i_8_113_2038_0, i_8_113_2107_0,
    i_8_113_2203_0, i_8_113_2214_0, i_8_113_2217_0, i_8_113_2227_0,
    i_8_113_2273_0, i_8_113_2286_0, i_8_113_2290_0,
    o_8_113_0_0  );
  input  i_8_113_38_0, i_8_113_40_0, i_8_113_43_0, i_8_113_81_0,
    i_8_113_84_0, i_8_113_115_0, i_8_113_148_0, i_8_113_151_0,
    i_8_113_163_0, i_8_113_190_0, i_8_113_194_0, i_8_113_245_0,
    i_8_113_346_0, i_8_113_347_0, i_8_113_352_0, i_8_113_417_0,
    i_8_113_464_0, i_8_113_469_0, i_8_113_470_0, i_8_113_483_0,
    i_8_113_489_0, i_8_113_490_0, i_8_113_522_0, i_8_113_526_0,
    i_8_113_538_0, i_8_113_552_0, i_8_113_555_0, i_8_113_595_0,
    i_8_113_598_0, i_8_113_634_0, i_8_113_648_0, i_8_113_695_0,
    i_8_113_697_0, i_8_113_700_0, i_8_113_702_0, i_8_113_706_0,
    i_8_113_733_0, i_8_113_734_0, i_8_113_770_0, i_8_113_790_0,
    i_8_113_793_0, i_8_113_813_0, i_8_113_833_0, i_8_113_881_0,
    i_8_113_893_0, i_8_113_896_0, i_8_113_926_0, i_8_113_998_0,
    i_8_113_1154_0, i_8_113_1161_0, i_8_113_1171_0, i_8_113_1223_0,
    i_8_113_1233_0, i_8_113_1238_0, i_8_113_1262_0, i_8_113_1288_0,
    i_8_113_1289_0, i_8_113_1292_0, i_8_113_1299_0, i_8_113_1306_0,
    i_8_113_1309_0, i_8_113_1311_0, i_8_113_1312_0, i_8_113_1352_0,
    i_8_113_1381_0, i_8_113_1384_0, i_8_113_1423_0, i_8_113_1442_0,
    i_8_113_1491_0, i_8_113_1498_0, i_8_113_1543_0, i_8_113_1549_0,
    i_8_113_1562_0, i_8_113_1637_0, i_8_113_1648_0, i_8_113_1653_0,
    i_8_113_1687_0, i_8_113_1688_0, i_8_113_1690_0, i_8_113_1701_0,
    i_8_113_1708_0, i_8_113_1748_0, i_8_113_1750_0, i_8_113_1753_0,
    i_8_113_1803_0, i_8_113_1806_0, i_8_113_1832_0, i_8_113_1840_0,
    i_8_113_1926_0, i_8_113_1960_0, i_8_113_1996_0, i_8_113_2038_0,
    i_8_113_2107_0, i_8_113_2203_0, i_8_113_2214_0, i_8_113_2217_0,
    i_8_113_2227_0, i_8_113_2273_0, i_8_113_2286_0, i_8_113_2290_0;
  output o_8_113_0_0;
  assign o_8_113_0_0 = 0;
endmodule



// Benchmark "kernel_8_114" written by ABC on Sun Jul 19 10:04:58 2020

module kernel_8_114 ( 
    i_8_114_16_0, i_8_114_17_0, i_8_114_43_0, i_8_114_67_0, i_8_114_68_0,
    i_8_114_115_0, i_8_114_143_0, i_8_114_187_0, i_8_114_223_0,
    i_8_114_301_0, i_8_114_322_0, i_8_114_363_0, i_8_114_366_0,
    i_8_114_367_0, i_8_114_368_0, i_8_114_382_0, i_8_114_403_0,
    i_8_114_416_0, i_8_114_430_0, i_8_114_475_0, i_8_114_476_0,
    i_8_114_511_0, i_8_114_529_0, i_8_114_539_0, i_8_114_592_0,
    i_8_114_603_0, i_8_114_606_0, i_8_114_608_0, i_8_114_609_0,
    i_8_114_610_0, i_8_114_611_0, i_8_114_634_0, i_8_114_637_0,
    i_8_114_643_0, i_8_114_655_0, i_8_114_660_0, i_8_114_664_0,
    i_8_114_682_0, i_8_114_840_0, i_8_114_842_0, i_8_114_843_0,
    i_8_114_844_0, i_8_114_845_0, i_8_114_881_0, i_8_114_895_0,
    i_8_114_970_0, i_8_114_977_0, i_8_114_1039_0, i_8_114_1106_0,
    i_8_114_1137_0, i_8_114_1184_0, i_8_114_1201_0, i_8_114_1264_0,
    i_8_114_1267_0, i_8_114_1282_0, i_8_114_1283_0, i_8_114_1285_0,
    i_8_114_1286_0, i_8_114_1301_0, i_8_114_1303_0, i_8_114_1318_0,
    i_8_114_1331_0, i_8_114_1340_0, i_8_114_1351_0, i_8_114_1366_0,
    i_8_114_1403_0, i_8_114_1426_0, i_8_114_1438_0, i_8_114_1465_0,
    i_8_114_1484_0, i_8_114_1493_0, i_8_114_1528_0, i_8_114_1529_0,
    i_8_114_1552_0, i_8_114_1555_0, i_8_114_1574_0, i_8_114_1649_0,
    i_8_114_1689_0, i_8_114_1690_0, i_8_114_1692_0, i_8_114_1697_0,
    i_8_114_1726_0, i_8_114_1771_0, i_8_114_1789_0, i_8_114_1794_0,
    i_8_114_1808_0, i_8_114_1840_0, i_8_114_1874_0, i_8_114_1885_0,
    i_8_114_1979_0, i_8_114_1981_0, i_8_114_2092_0, i_8_114_2096_0,
    i_8_114_2105_0, i_8_114_2173_0, i_8_114_2174_0, i_8_114_2227_0,
    i_8_114_2247_0, i_8_114_2248_0, i_8_114_2300_0,
    o_8_114_0_0  );
  input  i_8_114_16_0, i_8_114_17_0, i_8_114_43_0, i_8_114_67_0,
    i_8_114_68_0, i_8_114_115_0, i_8_114_143_0, i_8_114_187_0,
    i_8_114_223_0, i_8_114_301_0, i_8_114_322_0, i_8_114_363_0,
    i_8_114_366_0, i_8_114_367_0, i_8_114_368_0, i_8_114_382_0,
    i_8_114_403_0, i_8_114_416_0, i_8_114_430_0, i_8_114_475_0,
    i_8_114_476_0, i_8_114_511_0, i_8_114_529_0, i_8_114_539_0,
    i_8_114_592_0, i_8_114_603_0, i_8_114_606_0, i_8_114_608_0,
    i_8_114_609_0, i_8_114_610_0, i_8_114_611_0, i_8_114_634_0,
    i_8_114_637_0, i_8_114_643_0, i_8_114_655_0, i_8_114_660_0,
    i_8_114_664_0, i_8_114_682_0, i_8_114_840_0, i_8_114_842_0,
    i_8_114_843_0, i_8_114_844_0, i_8_114_845_0, i_8_114_881_0,
    i_8_114_895_0, i_8_114_970_0, i_8_114_977_0, i_8_114_1039_0,
    i_8_114_1106_0, i_8_114_1137_0, i_8_114_1184_0, i_8_114_1201_0,
    i_8_114_1264_0, i_8_114_1267_0, i_8_114_1282_0, i_8_114_1283_0,
    i_8_114_1285_0, i_8_114_1286_0, i_8_114_1301_0, i_8_114_1303_0,
    i_8_114_1318_0, i_8_114_1331_0, i_8_114_1340_0, i_8_114_1351_0,
    i_8_114_1366_0, i_8_114_1403_0, i_8_114_1426_0, i_8_114_1438_0,
    i_8_114_1465_0, i_8_114_1484_0, i_8_114_1493_0, i_8_114_1528_0,
    i_8_114_1529_0, i_8_114_1552_0, i_8_114_1555_0, i_8_114_1574_0,
    i_8_114_1649_0, i_8_114_1689_0, i_8_114_1690_0, i_8_114_1692_0,
    i_8_114_1697_0, i_8_114_1726_0, i_8_114_1771_0, i_8_114_1789_0,
    i_8_114_1794_0, i_8_114_1808_0, i_8_114_1840_0, i_8_114_1874_0,
    i_8_114_1885_0, i_8_114_1979_0, i_8_114_1981_0, i_8_114_2092_0,
    i_8_114_2096_0, i_8_114_2105_0, i_8_114_2173_0, i_8_114_2174_0,
    i_8_114_2227_0, i_8_114_2247_0, i_8_114_2248_0, i_8_114_2300_0;
  output o_8_114_0_0;
  assign o_8_114_0_0 = 0;
endmodule



// Benchmark "kernel_8_115" written by ABC on Sun Jul 19 10:05:00 2020

module kernel_8_115 ( 
    i_8_115_49_0, i_8_115_57_0, i_8_115_75_0, i_8_115_77_0, i_8_115_87_0,
    i_8_115_122_0, i_8_115_165_0, i_8_115_166_0, i_8_115_170_0,
    i_8_115_204_0, i_8_115_223_0, i_8_115_229_0, i_8_115_241_0,
    i_8_115_345_0, i_8_115_347_0, i_8_115_377_0, i_8_115_426_0,
    i_8_115_454_0, i_8_115_455_0, i_8_115_458_0, i_8_115_476_0,
    i_8_115_508_0, i_8_115_608_0, i_8_115_615_0, i_8_115_617_0,
    i_8_115_618_0, i_8_115_619_0, i_8_115_633_0, i_8_115_634_0,
    i_8_115_638_0, i_8_115_657_0, i_8_115_658_0, i_8_115_660_0,
    i_8_115_662_0, i_8_115_664_0, i_8_115_695_0, i_8_115_795_0,
    i_8_115_806_0, i_8_115_839_0, i_8_115_851_0, i_8_115_877_0,
    i_8_115_878_0, i_8_115_880_0, i_8_115_896_0, i_8_115_958_0,
    i_8_115_1012_0, i_8_115_1029_0, i_8_115_1030_0, i_8_115_1034_0,
    i_8_115_1037_0, i_8_115_1045_0, i_8_115_1071_0, i_8_115_1072_0,
    i_8_115_1076_0, i_8_115_1130_0, i_8_115_1166_0, i_8_115_1226_0,
    i_8_115_1228_0, i_8_115_1229_0, i_8_115_1240_0, i_8_115_1263_0,
    i_8_115_1264_0, i_8_115_1284_0, i_8_115_1293_0, i_8_115_1296_0,
    i_8_115_1298_0, i_8_115_1300_0, i_8_115_1301_0, i_8_115_1329_0,
    i_8_115_1453_0, i_8_115_1454_0, i_8_115_1455_0, i_8_115_1457_0,
    i_8_115_1506_0, i_8_115_1509_0, i_8_115_1510_0, i_8_115_1542_0,
    i_8_115_1543_0, i_8_115_1544_0, i_8_115_1550_0, i_8_115_1552_0,
    i_8_115_1607_0, i_8_115_1630_0, i_8_115_1806_0, i_8_115_1862_0,
    i_8_115_1893_0, i_8_115_1894_0, i_8_115_1895_0, i_8_115_1898_0,
    i_8_115_1951_0, i_8_115_2041_0, i_8_115_2096_0, i_8_115_2126_0,
    i_8_115_2128_0, i_8_115_2129_0, i_8_115_2143_0, i_8_115_2217_0,
    i_8_115_2218_0, i_8_115_2227_0, i_8_115_2273_0,
    o_8_115_0_0  );
  input  i_8_115_49_0, i_8_115_57_0, i_8_115_75_0, i_8_115_77_0,
    i_8_115_87_0, i_8_115_122_0, i_8_115_165_0, i_8_115_166_0,
    i_8_115_170_0, i_8_115_204_0, i_8_115_223_0, i_8_115_229_0,
    i_8_115_241_0, i_8_115_345_0, i_8_115_347_0, i_8_115_377_0,
    i_8_115_426_0, i_8_115_454_0, i_8_115_455_0, i_8_115_458_0,
    i_8_115_476_0, i_8_115_508_0, i_8_115_608_0, i_8_115_615_0,
    i_8_115_617_0, i_8_115_618_0, i_8_115_619_0, i_8_115_633_0,
    i_8_115_634_0, i_8_115_638_0, i_8_115_657_0, i_8_115_658_0,
    i_8_115_660_0, i_8_115_662_0, i_8_115_664_0, i_8_115_695_0,
    i_8_115_795_0, i_8_115_806_0, i_8_115_839_0, i_8_115_851_0,
    i_8_115_877_0, i_8_115_878_0, i_8_115_880_0, i_8_115_896_0,
    i_8_115_958_0, i_8_115_1012_0, i_8_115_1029_0, i_8_115_1030_0,
    i_8_115_1034_0, i_8_115_1037_0, i_8_115_1045_0, i_8_115_1071_0,
    i_8_115_1072_0, i_8_115_1076_0, i_8_115_1130_0, i_8_115_1166_0,
    i_8_115_1226_0, i_8_115_1228_0, i_8_115_1229_0, i_8_115_1240_0,
    i_8_115_1263_0, i_8_115_1264_0, i_8_115_1284_0, i_8_115_1293_0,
    i_8_115_1296_0, i_8_115_1298_0, i_8_115_1300_0, i_8_115_1301_0,
    i_8_115_1329_0, i_8_115_1453_0, i_8_115_1454_0, i_8_115_1455_0,
    i_8_115_1457_0, i_8_115_1506_0, i_8_115_1509_0, i_8_115_1510_0,
    i_8_115_1542_0, i_8_115_1543_0, i_8_115_1544_0, i_8_115_1550_0,
    i_8_115_1552_0, i_8_115_1607_0, i_8_115_1630_0, i_8_115_1806_0,
    i_8_115_1862_0, i_8_115_1893_0, i_8_115_1894_0, i_8_115_1895_0,
    i_8_115_1898_0, i_8_115_1951_0, i_8_115_2041_0, i_8_115_2096_0,
    i_8_115_2126_0, i_8_115_2128_0, i_8_115_2129_0, i_8_115_2143_0,
    i_8_115_2217_0, i_8_115_2218_0, i_8_115_2227_0, i_8_115_2273_0;
  output o_8_115_0_0;
  assign o_8_115_0_0 = ~((i_8_115_49_0 & ((i_8_115_1284_0 & ~i_8_115_1544_0 & ~i_8_115_1862_0 & ~i_8_115_1893_0 & ~i_8_115_1898_0) | (~i_8_115_229_0 & ~i_8_115_377_0 & ~i_8_115_1029_0 & ~i_8_115_1030_0 & ~i_8_115_1453_0 & ~i_8_115_1457_0 & ~i_8_115_1550_0 & ~i_8_115_1806_0 & ~i_8_115_1895_0 & ~i_8_115_2096_0 & ~i_8_115_2217_0))) | (i_8_115_77_0 & ((~i_8_115_49_0 & ~i_8_115_806_0 & ~i_8_115_1037_0 & ~i_8_115_1045_0 & ~i_8_115_1329_0 & ~i_8_115_1550_0 & ~i_8_115_2218_0) | (~i_8_115_345_0 & ~i_8_115_476_0 & ~i_8_115_695_0 & ~i_8_115_851_0 & ~i_8_115_1510_0 & ~i_8_115_2096_0 & ~i_8_115_2273_0))) | (~i_8_115_204_0 & ((~i_8_115_57_0 & ~i_8_115_241_0 & i_8_115_662_0 & ~i_8_115_851_0 & ~i_8_115_878_0 & ~i_8_115_880_0 & ~i_8_115_1072_0 & ~i_8_115_1607_0 & ~i_8_115_1806_0) | (~i_8_115_377_0 & ~i_8_115_476_0 & ~i_8_115_608_0 & ~i_8_115_618_0 & ~i_8_115_664_0 & ~i_8_115_695_0 & ~i_8_115_1012_0 & ~i_8_115_1029_0 & ~i_8_115_1030_0 & ~i_8_115_1037_0 & ~i_8_115_1045_0 & ~i_8_115_1071_0 & ~i_8_115_1264_0 & ~i_8_115_1296_0 & ~i_8_115_1506_0 & ~i_8_115_1893_0 & ~i_8_115_2217_0 & ~i_8_115_2218_0))) | (i_8_115_455_0 & ((~i_8_115_377_0 & ~i_8_115_795_0 & ~i_8_115_1130_0 & ~i_8_115_1893_0 & ~i_8_115_2128_0) | (~i_8_115_1012_0 & i_8_115_1030_0 & ~i_8_115_1264_0 & i_8_115_2129_0))) | (~i_8_115_508_0 & ((~i_8_115_49_0 & ~i_8_115_638_0 & ~i_8_115_878_0 & ~i_8_115_880_0 & ~i_8_115_1029_0 & ~i_8_115_1166_0 & ~i_8_115_1455_0 & i_8_115_1506_0 & ~i_8_115_1893_0 & ~i_8_115_1951_0) | (~i_8_115_223_0 & ~i_8_115_377_0 & i_8_115_1263_0 & i_8_115_1264_0 & ~i_8_115_1329_0 & ~i_8_115_1454_0 & ~i_8_115_1543_0 & ~i_8_115_1607_0 & ~i_8_115_2126_0))) | (~i_8_115_2126_0 & ((~i_8_115_49_0 & ((~i_8_115_454_0 & i_8_115_660_0 & ~i_8_115_1045_0 & i_8_115_1506_0 & ~i_8_115_1862_0) | (~i_8_115_75_0 & ~i_8_115_170_0 & i_8_115_617_0 & ~i_8_115_1542_0 & ~i_8_115_2129_0 & i_8_115_2273_0))) | (~i_8_115_1029_0 & ((~i_8_115_608_0 & ~i_8_115_1453_0 & ((i_8_115_958_0 & ~i_8_115_1030_0 & ~i_8_115_1166_0 & ~i_8_115_1455_0 & ~i_8_115_1457_0) | (~i_8_115_476_0 & ~i_8_115_1296_0 & ~i_8_115_1543_0 & ~i_8_115_1630_0 & i_8_115_2128_0 & ~i_8_115_2218_0 & ~i_8_115_2273_0))) | (~i_8_115_1895_0 & ((i_8_115_658_0 & ~i_8_115_1455_0 & ~i_8_115_1893_0) | (~i_8_115_223_0 & ~i_8_115_426_0 & ~i_8_115_839_0 & ~i_8_115_877_0 & ~i_8_115_1034_0 & ~i_8_115_1037_0 & ~i_8_115_1166_0 & ~i_8_115_1509_0 & ~i_8_115_1550_0 & ~i_8_115_1898_0 & ~i_8_115_1951_0))))) | (~i_8_115_839_0 & ~i_8_115_896_0 & ~i_8_115_1284_0 & i_8_115_1454_0 & ~i_8_115_1457_0 & i_8_115_1862_0 & ~i_8_115_2096_0) | (~i_8_115_1544_0 & i_8_115_1552_0 & i_8_115_1607_0 & i_8_115_2143_0 & i_8_115_2273_0))) | (~i_8_115_2217_0 & ((~i_8_115_347_0 & ((~i_8_115_426_0 & i_8_115_608_0 & i_8_115_634_0 & ~i_8_115_1130_0 & ~i_8_115_1550_0 & i_8_115_2128_0) | (~i_8_115_57_0 & ~i_8_115_345_0 & ~i_8_115_377_0 & ~i_8_115_880_0 & ~i_8_115_958_0 & ~i_8_115_1037_0 & ~i_8_115_1045_0 & ~i_8_115_1542_0 & ~i_8_115_1862_0 & ~i_8_115_1893_0 & ~i_8_115_1898_0 & ~i_8_115_2096_0 & ~i_8_115_2129_0))) | (~i_8_115_1029_0 & ~i_8_115_1510_0 & ((~i_8_115_229_0 & ~i_8_115_377_0 & ~i_8_115_454_0 & ~i_8_115_1030_0 & i_8_115_1264_0 & ~i_8_115_1454_0 & ~i_8_115_1455_0 & ~i_8_115_1506_0) | (~i_8_115_223_0 & ~i_8_115_476_0 & ~i_8_115_1045_0 & ~i_8_115_1130_0 & ~i_8_115_1166_0 & ~i_8_115_1284_0 & ~i_8_115_1542_0 & i_8_115_1552_0 & ~i_8_115_1893_0 & ~i_8_115_1898_0 & ~i_8_115_2129_0))) | (i_8_115_851_0 & ~i_8_115_1263_0 & ~i_8_115_1453_0 & ~i_8_115_1454_0 & ~i_8_115_1506_0 & ~i_8_115_1552_0 & ~i_8_115_1898_0))) | (~i_8_115_57_0 & ((~i_8_115_878_0 & ~i_8_115_880_0 & ~i_8_115_617_0 & ~i_8_115_658_0 & ~i_8_115_1030_0 & ~i_8_115_1226_0 & ~i_8_115_1506_0 & i_8_115_2143_0) | (i_8_115_87_0 & ~i_8_115_1012_0 & ~i_8_115_1509_0 & ~i_8_115_1510_0 & i_8_115_1806_0 & ~i_8_115_2273_0))) | (~i_8_115_223_0 & ((~i_8_115_345_0 & ~i_8_115_877_0 & ~i_8_115_880_0 & i_8_115_1264_0 & ~i_8_115_1454_0) | (i_8_115_1012_0 & i_8_115_1030_0 & ~i_8_115_1045_0 & ~i_8_115_1453_0 & i_8_115_1552_0))) | (~i_8_115_2096_0 & ((~i_8_115_170_0 & ~i_8_115_1509_0 & ((~i_8_115_1130_0 & i_8_115_1228_0) | (~i_8_115_77_0 & ~i_8_115_345_0 & ~i_8_115_851_0 & ~i_8_115_1012_0 & ~i_8_115_1029_0 & ~i_8_115_1045_0 & ~i_8_115_1510_0 & ~i_8_115_1552_0 & ~i_8_115_1894_0 & ~i_8_115_1898_0 & ~i_8_115_2128_0 & ~i_8_115_2273_0))) | (~i_8_115_1453_0 & ~i_8_115_1543_0 & ((~i_8_115_345_0 & ~i_8_115_476_0 & i_8_115_619_0 & ~i_8_115_1544_0) | (i_8_115_1284_0 & ~i_8_115_1510_0 & ~i_8_115_1542_0 & ~i_8_115_1607_0 & ~i_8_115_1806_0))))) | (~i_8_115_347_0 & ((~i_8_115_426_0 & i_8_115_664_0 & ~i_8_115_877_0 & ~i_8_115_1509_0 & ~i_8_115_1510_0) | (~i_8_115_608_0 & i_8_115_660_0 & ~i_8_115_1045_0 & ~i_8_115_1166_0 & ~i_8_115_1506_0 & ~i_8_115_2128_0))) | (~i_8_115_1898_0 & ((~i_8_115_476_0 & ~i_8_115_1552_0 & ~i_8_115_2227_0 & ((~i_8_115_229_0 & ~i_8_115_454_0 & ~i_8_115_1012_0 & ~i_8_115_1130_0 & ~i_8_115_1166_0 & i_8_115_1240_0 & ~i_8_115_1454_0 & ~i_8_115_1543_0) | (~i_8_115_87_0 & ~i_8_115_122_0 & ~i_8_115_426_0 & ~i_8_115_633_0 & ~i_8_115_658_0 & ~i_8_115_795_0 & i_8_115_877_0 & ~i_8_115_1034_0 & ~i_8_115_1226_0 & ~i_8_115_1298_0 & ~i_8_115_1509_0 & ~i_8_115_1510_0 & ~i_8_115_1607_0 & ~i_8_115_1895_0))) | (~i_8_115_426_0 & ((i_8_115_241_0 & i_8_115_618_0 & ~i_8_115_1228_0 & ~i_8_115_1544_0) | (~i_8_115_880_0 & ~i_8_115_958_0 & ~i_8_115_1329_0 & ~i_8_115_1453_0 & ~i_8_115_1509_0 & ~i_8_115_1895_0 & ~i_8_115_2128_0 & i_8_115_2218_0 & ~i_8_115_2273_0))) | (i_8_115_458_0 & ~i_8_115_634_0 & ~i_8_115_664_0 & ~i_8_115_695_0 & ~i_8_115_795_0 & ~i_8_115_1166_0 & ~i_8_115_1453_0 & ~i_8_115_1509_0 & ~i_8_115_1630_0 & ~i_8_115_1895_0 & i_8_115_2096_0) | (~i_8_115_170_0 & ~i_8_115_877_0 & ~i_8_115_958_0 & ~i_8_115_1130_0 & ~i_8_115_1300_0 & ~i_8_115_1506_0 & ~i_8_115_1607_0 & ~i_8_115_2041_0 & i_8_115_2143_0 & ~i_8_115_2273_0))) | (~i_8_115_229_0 & ((~i_8_115_795_0 & ~i_8_115_1509_0 & ~i_8_115_1552_0 & ~i_8_115_1607_0 & i_8_115_1630_0) | (i_8_115_618_0 & ~i_8_115_1045_0 & i_8_115_1284_0 & ~i_8_115_1806_0))) | (~i_8_115_1607_0 & ((~i_8_115_695_0 & ((i_8_115_633_0 & ~i_8_115_1012_0 & ~i_8_115_1509_0) | (i_8_115_619_0 & ~i_8_115_877_0 & ~i_8_115_958_0 & ~i_8_115_1284_0 & ~i_8_115_1862_0 & ~i_8_115_2273_0))) | (~i_8_115_458_0 & i_8_115_806_0 & ~i_8_115_1542_0))) | (~i_8_115_1029_0 & ~i_8_115_1453_0 & ~i_8_115_1454_0 & ((i_8_115_1298_0 & ~i_8_115_1457_0 & ~i_8_115_2218_0) | (i_8_115_75_0 & ~i_8_115_1030_0 & ~i_8_115_1045_0 & ~i_8_115_1263_0 & ~i_8_115_1455_0 & ~i_8_115_2129_0 & ~i_8_115_2273_0))) | (~i_8_115_1166_0 & ((~i_8_115_1130_0 & i_8_115_1229_0 & ~i_8_115_1542_0 & ~i_8_115_1894_0) | (~i_8_115_634_0 & ~i_8_115_1226_0 & i_8_115_1263_0 & ~i_8_115_1329_0 & ~i_8_115_1506_0 & ~i_8_115_1510_0 & ~i_8_115_1895_0))) | (~i_8_115_1542_0 & ((~i_8_115_166_0 & ~i_8_115_426_0 & ~i_8_115_839_0 & i_8_115_877_0 & i_8_115_1630_0) | (i_8_115_615_0 & ~i_8_115_664_0 & i_8_115_1029_0 & ~i_8_115_1894_0))) | (~i_8_115_455_0 & i_8_115_1045_0 & i_8_115_1076_0 & i_8_115_1264_0) | (~i_8_115_1045_0 & i_8_115_1072_0 & ~i_8_115_1329_0 & ~i_8_115_1543_0));
endmodule



// Benchmark "kernel_8_116" written by ABC on Sun Jul 19 10:05:02 2020

module kernel_8_116 ( 
    i_8_116_160_0, i_8_116_186_0, i_8_116_257_0, i_8_116_293_0,
    i_8_116_331_0, i_8_116_373_0, i_8_116_381_0, i_8_116_394_0,
    i_8_116_430_0, i_8_116_462_0, i_8_116_463_0, i_8_116_464_0,
    i_8_116_528_0, i_8_116_529_0, i_8_116_553_0, i_8_116_556_0,
    i_8_116_592_0, i_8_116_593_0, i_8_116_599_0, i_8_116_607_0,
    i_8_116_608_0, i_8_116_615_0, i_8_116_636_0, i_8_116_653_0,
    i_8_116_661_0, i_8_116_665_0, i_8_116_710_0, i_8_116_760_0,
    i_8_116_780_0, i_8_116_782_0, i_8_116_795_0, i_8_116_817_0,
    i_8_116_827_0, i_8_116_833_0, i_8_116_838_0, i_8_116_955_0,
    i_8_116_998_0, i_8_116_1074_0, i_8_116_1078_0, i_8_116_1114_0,
    i_8_116_1160_0, i_8_116_1191_0, i_8_116_1231_0, i_8_116_1258_0,
    i_8_116_1285_0, i_8_116_1300_0, i_8_116_1318_0, i_8_116_1331_0,
    i_8_116_1382_0, i_8_116_1437_0, i_8_116_1438_0, i_8_116_1439_0,
    i_8_116_1452_0, i_8_116_1453_0, i_8_116_1480_0, i_8_116_1483_0,
    i_8_116_1506_0, i_8_116_1534_0, i_8_116_1535_0, i_8_116_1542_0,
    i_8_116_1547_0, i_8_116_1553_0, i_8_116_1562_0, i_8_116_1588_0,
    i_8_116_1592_0, i_8_116_1605_0, i_8_116_1615_0, i_8_116_1634_0,
    i_8_116_1715_0, i_8_116_1722_0, i_8_116_1762_0, i_8_116_1789_0,
    i_8_116_1799_0, i_8_116_1813_0, i_8_116_1822_0, i_8_116_1830_0,
    i_8_116_1839_0, i_8_116_1841_0, i_8_116_1867_0, i_8_116_1888_0,
    i_8_116_1893_0, i_8_116_1897_0, i_8_116_1898_0, i_8_116_1900_0,
    i_8_116_1922_0, i_8_116_1948_0, i_8_116_1965_0, i_8_116_1966_0,
    i_8_116_1995_0, i_8_116_1996_0, i_8_116_2001_0, i_8_116_2014_0,
    i_8_116_2109_0, i_8_116_2128_0, i_8_116_2163_0, i_8_116_2203_0,
    i_8_116_2216_0, i_8_116_2260_0, i_8_116_2264_0, i_8_116_2274_0,
    o_8_116_0_0  );
  input  i_8_116_160_0, i_8_116_186_0, i_8_116_257_0, i_8_116_293_0,
    i_8_116_331_0, i_8_116_373_0, i_8_116_381_0, i_8_116_394_0,
    i_8_116_430_0, i_8_116_462_0, i_8_116_463_0, i_8_116_464_0,
    i_8_116_528_0, i_8_116_529_0, i_8_116_553_0, i_8_116_556_0,
    i_8_116_592_0, i_8_116_593_0, i_8_116_599_0, i_8_116_607_0,
    i_8_116_608_0, i_8_116_615_0, i_8_116_636_0, i_8_116_653_0,
    i_8_116_661_0, i_8_116_665_0, i_8_116_710_0, i_8_116_760_0,
    i_8_116_780_0, i_8_116_782_0, i_8_116_795_0, i_8_116_817_0,
    i_8_116_827_0, i_8_116_833_0, i_8_116_838_0, i_8_116_955_0,
    i_8_116_998_0, i_8_116_1074_0, i_8_116_1078_0, i_8_116_1114_0,
    i_8_116_1160_0, i_8_116_1191_0, i_8_116_1231_0, i_8_116_1258_0,
    i_8_116_1285_0, i_8_116_1300_0, i_8_116_1318_0, i_8_116_1331_0,
    i_8_116_1382_0, i_8_116_1437_0, i_8_116_1438_0, i_8_116_1439_0,
    i_8_116_1452_0, i_8_116_1453_0, i_8_116_1480_0, i_8_116_1483_0,
    i_8_116_1506_0, i_8_116_1534_0, i_8_116_1535_0, i_8_116_1542_0,
    i_8_116_1547_0, i_8_116_1553_0, i_8_116_1562_0, i_8_116_1588_0,
    i_8_116_1592_0, i_8_116_1605_0, i_8_116_1615_0, i_8_116_1634_0,
    i_8_116_1715_0, i_8_116_1722_0, i_8_116_1762_0, i_8_116_1789_0,
    i_8_116_1799_0, i_8_116_1813_0, i_8_116_1822_0, i_8_116_1830_0,
    i_8_116_1839_0, i_8_116_1841_0, i_8_116_1867_0, i_8_116_1888_0,
    i_8_116_1893_0, i_8_116_1897_0, i_8_116_1898_0, i_8_116_1900_0,
    i_8_116_1922_0, i_8_116_1948_0, i_8_116_1965_0, i_8_116_1966_0,
    i_8_116_1995_0, i_8_116_1996_0, i_8_116_2001_0, i_8_116_2014_0,
    i_8_116_2109_0, i_8_116_2128_0, i_8_116_2163_0, i_8_116_2203_0,
    i_8_116_2216_0, i_8_116_2260_0, i_8_116_2264_0, i_8_116_2274_0;
  output o_8_116_0_0;
  assign o_8_116_0_0 = ~((~i_8_116_160_0 & ((i_8_116_430_0 & ~i_8_116_1588_0 & ~i_8_116_1592_0 & ~i_8_116_1715_0) | (~i_8_116_782_0 & ~i_8_116_795_0 & ~i_8_116_1437_0 & ~i_8_116_1439_0 & ~i_8_116_1762_0))) | (~i_8_116_430_0 & ((~i_8_116_394_0 & ~i_8_116_464_0 & ~i_8_116_556_0 & ~i_8_116_833_0 & ~i_8_116_1300_0 & ~i_8_116_1542_0 & ~i_8_116_1722_0 & ~i_8_116_1799_0 & ~i_8_116_1948_0) | (i_8_116_608_0 & i_8_116_827_0 & ~i_8_116_1535_0 & ~i_8_116_2128_0))) | (~i_8_116_760_0 & ((~i_8_116_394_0 & ((~i_8_116_782_0 & ~i_8_116_1160_0 & ~i_8_116_1191_0 & ~i_8_116_2216_0) | (~i_8_116_1542_0 & ~i_8_116_1588_0 & ~i_8_116_1592_0 & ~i_8_116_1799_0 & ~i_8_116_2274_0))) | (~i_8_116_529_0 & ~i_8_116_608_0 & ~i_8_116_1897_0 & ~i_8_116_1898_0))) | (~i_8_116_463_0 & ((i_8_116_599_0 & ~i_8_116_1535_0 & ~i_8_116_1605_0 & i_8_116_1813_0) | (~i_8_116_782_0 & ~i_8_116_827_0 & ~i_8_116_1258_0 & ~i_8_116_1592_0 & ~i_8_116_1762_0 & ~i_8_116_1965_0))) | (~i_8_116_1258_0 & ((~i_8_116_528_0 & ~i_8_116_608_0 & ~i_8_116_782_0 & ~i_8_116_1078_0 & ~i_8_116_1382_0 & ~i_8_116_1841_0 & ~i_8_116_1897_0 & ~i_8_116_1900_0) | (~i_8_116_331_0 & i_8_116_1300_0 & ~i_8_116_1762_0 & ~i_8_116_2109_0))) | (~i_8_116_1898_0 & ((~i_8_116_608_0 & ((~i_8_116_462_0 & ~i_8_116_553_0 & ~i_8_116_1897_0 & ~i_8_116_1922_0) | (i_8_116_529_0 & ~i_8_116_653_0 & ~i_8_116_710_0 & ~i_8_116_1231_0 & ~i_8_116_1382_0 & ~i_8_116_1715_0 & ~i_8_116_1722_0 & ~i_8_116_1789_0 & ~i_8_116_1841_0 & ~i_8_116_2001_0))) | (i_8_116_553_0 & ~i_8_116_955_0 & i_8_116_1439_0 & ~i_8_116_1452_0 & i_8_116_1534_0 & i_8_116_1588_0 & ~i_8_116_1592_0 & ~i_8_116_1605_0))) | (~i_8_116_1285_0 & ((~i_8_116_1160_0 & ~i_8_116_1191_0 & ~i_8_116_1562_0 & ~i_8_116_1722_0 & ~i_8_116_1893_0 & i_8_116_1966_0) | (~i_8_116_1534_0 & ~i_8_116_1588_0 & ~i_8_116_2128_0))) | (~i_8_116_1592_0 & ((~i_8_116_1506_0 & ~i_8_116_1534_0 & i_8_116_1888_0) | (~i_8_116_464_0 & ~i_8_116_592_0 & i_8_116_1439_0 & ~i_8_116_1605_0 & ~i_8_116_1841_0 & ~i_8_116_1893_0) | (~i_8_116_293_0 & i_8_116_528_0 & ~i_8_116_607_0 & ~i_8_116_665_0 & ~i_8_116_1542_0 & ~i_8_116_1547_0 & ~i_8_116_2128_0))));
endmodule



// Benchmark "kernel_8_117" written by ABC on Sun Jul 19 10:05:04 2020

module kernel_8_117 ( 
    i_8_117_22_0, i_8_117_23_0, i_8_117_109_0, i_8_117_136_0,
    i_8_117_138_0, i_8_117_139_0, i_8_117_140_0, i_8_117_142_0,
    i_8_117_143_0, i_8_117_269_0, i_8_117_324_0, i_8_117_325_0,
    i_8_117_326_0, i_8_117_366_0, i_8_117_385_0, i_8_117_420_0,
    i_8_117_421_0, i_8_117_422_0, i_8_117_446_0, i_8_117_459_0,
    i_8_117_461_0, i_8_117_469_0, i_8_117_472_0, i_8_117_474_0,
    i_8_117_475_0, i_8_117_492_0, i_8_117_496_0, i_8_117_575_0,
    i_8_117_592_0, i_8_117_629_0, i_8_117_657_0, i_8_117_658_0,
    i_8_117_709_0, i_8_117_792_0, i_8_117_795_0, i_8_117_804_0,
    i_8_117_817_0, i_8_117_838_0, i_8_117_877_0, i_8_117_878_0,
    i_8_117_880_0, i_8_117_993_0, i_8_117_1078_0, i_8_117_1111_0,
    i_8_117_1114_0, i_8_117_1159_0, i_8_117_1185_0, i_8_117_1230_0,
    i_8_117_1279_0, i_8_117_1365_0, i_8_117_1393_0, i_8_117_1410_0,
    i_8_117_1426_0, i_8_117_1437_0, i_8_117_1471_0, i_8_117_1480_0,
    i_8_117_1482_0, i_8_117_1524_0, i_8_117_1607_0, i_8_117_1608_0,
    i_8_117_1609_0, i_8_117_1610_0, i_8_117_1652_0, i_8_117_1655_0,
    i_8_117_1677_0, i_8_117_1719_0, i_8_117_1724_0, i_8_117_1725_0,
    i_8_117_1732_0, i_8_117_1736_0, i_8_117_1747_0, i_8_117_1753_0,
    i_8_117_1787_0, i_8_117_1802_0, i_8_117_1805_0, i_8_117_1806_0,
    i_8_117_1856_0, i_8_117_1860_0, i_8_117_1886_0, i_8_117_1901_0,
    i_8_117_1903_0, i_8_117_1904_0, i_8_117_1945_0, i_8_117_1946_0,
    i_8_117_1948_0, i_8_117_1949_0, i_8_117_1951_0, i_8_117_1964_0,
    i_8_117_1967_0, i_8_117_1970_0, i_8_117_1992_0, i_8_117_2031_0,
    i_8_117_2109_0, i_8_117_2112_0, i_8_117_2137_0, i_8_117_2152_0,
    i_8_117_2153_0, i_8_117_2156_0, i_8_117_2158_0, i_8_117_2226_0,
    o_8_117_0_0  );
  input  i_8_117_22_0, i_8_117_23_0, i_8_117_109_0, i_8_117_136_0,
    i_8_117_138_0, i_8_117_139_0, i_8_117_140_0, i_8_117_142_0,
    i_8_117_143_0, i_8_117_269_0, i_8_117_324_0, i_8_117_325_0,
    i_8_117_326_0, i_8_117_366_0, i_8_117_385_0, i_8_117_420_0,
    i_8_117_421_0, i_8_117_422_0, i_8_117_446_0, i_8_117_459_0,
    i_8_117_461_0, i_8_117_469_0, i_8_117_472_0, i_8_117_474_0,
    i_8_117_475_0, i_8_117_492_0, i_8_117_496_0, i_8_117_575_0,
    i_8_117_592_0, i_8_117_629_0, i_8_117_657_0, i_8_117_658_0,
    i_8_117_709_0, i_8_117_792_0, i_8_117_795_0, i_8_117_804_0,
    i_8_117_817_0, i_8_117_838_0, i_8_117_877_0, i_8_117_878_0,
    i_8_117_880_0, i_8_117_993_0, i_8_117_1078_0, i_8_117_1111_0,
    i_8_117_1114_0, i_8_117_1159_0, i_8_117_1185_0, i_8_117_1230_0,
    i_8_117_1279_0, i_8_117_1365_0, i_8_117_1393_0, i_8_117_1410_0,
    i_8_117_1426_0, i_8_117_1437_0, i_8_117_1471_0, i_8_117_1480_0,
    i_8_117_1482_0, i_8_117_1524_0, i_8_117_1607_0, i_8_117_1608_0,
    i_8_117_1609_0, i_8_117_1610_0, i_8_117_1652_0, i_8_117_1655_0,
    i_8_117_1677_0, i_8_117_1719_0, i_8_117_1724_0, i_8_117_1725_0,
    i_8_117_1732_0, i_8_117_1736_0, i_8_117_1747_0, i_8_117_1753_0,
    i_8_117_1787_0, i_8_117_1802_0, i_8_117_1805_0, i_8_117_1806_0,
    i_8_117_1856_0, i_8_117_1860_0, i_8_117_1886_0, i_8_117_1901_0,
    i_8_117_1903_0, i_8_117_1904_0, i_8_117_1945_0, i_8_117_1946_0,
    i_8_117_1948_0, i_8_117_1949_0, i_8_117_1951_0, i_8_117_1964_0,
    i_8_117_1967_0, i_8_117_1970_0, i_8_117_1992_0, i_8_117_2031_0,
    i_8_117_2109_0, i_8_117_2112_0, i_8_117_2137_0, i_8_117_2152_0,
    i_8_117_2153_0, i_8_117_2156_0, i_8_117_2158_0, i_8_117_2226_0;
  output o_8_117_0_0;
  assign o_8_117_0_0 = ~((~i_8_117_138_0 & ((~i_8_117_469_0 & ~i_8_117_1787_0 & i_8_117_1886_0 & ~i_8_117_1948_0 & i_8_117_1970_0 & ~i_8_117_2112_0) | (~i_8_117_496_0 & ~i_8_117_795_0 & ~i_8_117_993_0 & i_8_117_1279_0 & ~i_8_117_1607_0 & ~i_8_117_1652_0 & ~i_8_117_1802_0 & ~i_8_117_1805_0 & ~i_8_117_1951_0 & ~i_8_117_1964_0 & ~i_8_117_2109_0 & i_8_117_2137_0 & ~i_8_117_2158_0))) | (~i_8_117_2112_0 & ((~i_8_117_109_0 & ((~i_8_117_23_0 & ~i_8_117_136_0 & ~i_8_117_366_0 & ~i_8_117_461_0 & ~i_8_117_880_0 & ~i_8_117_1677_0 & ~i_8_117_1886_0 & ~i_8_117_1945_0 & ~i_8_117_1992_0 & ~i_8_117_2109_0 & i_8_117_2156_0 & ~i_8_117_2158_0) | (~i_8_117_657_0 & ~i_8_117_877_0 & ~i_8_117_1230_0 & ~i_8_117_1805_0 & ~i_8_117_1964_0 & ~i_8_117_1967_0 & ~i_8_117_2137_0 & ~i_8_117_2152_0 & ~i_8_117_2156_0 & i_8_117_2158_0 & ~i_8_117_2226_0))) | (i_8_117_139_0 & ((~i_8_117_385_0 & ~i_8_117_475_0 & ~i_8_117_1230_0 & ~i_8_117_1607_0 & ~i_8_117_1652_0 & ~i_8_117_1732_0 & i_8_117_1747_0 & ~i_8_117_1964_0) | (~i_8_117_22_0 & ~i_8_117_469_0 & ~i_8_117_709_0 & ~i_8_117_795_0 & ~i_8_117_1610_0 & ~i_8_117_1747_0 & ~i_8_117_1753_0 & ~i_8_117_1903_0 & ~i_8_117_2109_0))) | (~i_8_117_2109_0 & ((~i_8_117_22_0 & ((i_8_117_421_0 & i_8_117_1393_0 & ~i_8_117_1607_0 & ~i_8_117_1747_0 & ~i_8_117_1787_0) | (i_8_117_136_0 & ~i_8_117_792_0 & ~i_8_117_1471_0 & ~i_8_117_1805_0 & ~i_8_117_1967_0 & ~i_8_117_2153_0))) | (~i_8_117_2153_0 & ((~i_8_117_23_0 & ((~i_8_117_143_0 & ~i_8_117_461_0 & i_8_117_629_0 & i_8_117_709_0 & ~i_8_117_1159_0 & ~i_8_117_1437_0 & ~i_8_117_1967_0) | (~i_8_117_474_0 & ~i_8_117_492_0 & ~i_8_117_795_0 & ~i_8_117_993_0 & i_8_117_1111_0 & ~i_8_117_1230_0 & ~i_8_117_1279_0 & ~i_8_117_1482_0 & ~i_8_117_1607_0 & ~i_8_117_1787_0 & ~i_8_117_1970_0 & ~i_8_117_2152_0))) | (~i_8_117_459_0 & ~i_8_117_1951_0 & ((i_8_117_109_0 & ~i_8_117_795_0 & ~i_8_117_878_0 & ~i_8_117_1111_0 & ~i_8_117_1471_0 & ~i_8_117_1732_0 & ~i_8_117_1856_0) | (~i_8_117_474_0 & ~i_8_117_709_0 & ~i_8_117_993_0 & ~i_8_117_1230_0 & ~i_8_117_1609_0 & ~i_8_117_1610_0 & ~i_8_117_1802_0 & ~i_8_117_1945_0 & ~i_8_117_1964_0 & ~i_8_117_2137_0))))) | (~i_8_117_1607_0 & ~i_8_117_1609_0 & ((~i_8_117_143_0 & i_8_117_658_0 & ~i_8_117_792_0 & i_8_117_838_0 & ~i_8_117_1802_0 & ~i_8_117_1946_0) | (i_8_117_142_0 & ~i_8_117_326_0 & ~i_8_117_1610_0 & i_8_117_1753_0 & ~i_8_117_1806_0 & ~i_8_117_1860_0 & ~i_8_117_2156_0))) | (~i_8_117_139_0 & ~i_8_117_446_0 & ~i_8_117_459_0 & ~i_8_117_474_0 & ~i_8_117_629_0 & ~i_8_117_838_0 & i_8_117_1111_0 & ~i_8_117_1471_0 & ~i_8_117_1608_0 & ~i_8_117_1652_0 & ~i_8_117_1787_0 & ~i_8_117_1805_0 & ~i_8_117_1946_0 & ~i_8_117_1964_0 & ~i_8_117_2152_0))) | (~i_8_117_23_0 & ((i_8_117_492_0 & ~i_8_117_496_0 & ~i_8_117_792_0 & ~i_8_117_878_0 & ~i_8_117_1279_0 & ~i_8_117_1437_0 & ~i_8_117_1609_0 & ~i_8_117_1610_0) | (i_8_117_143_0 & ~i_8_117_385_0 & ~i_8_117_459_0 & ~i_8_117_657_0 & ~i_8_117_1159_0 & ~i_8_117_1607_0 & ~i_8_117_1970_0))) | (~i_8_117_1949_0 & ((i_8_117_109_0 & ((~i_8_117_22_0 & i_8_117_880_0 & ~i_8_117_1652_0 & ~i_8_117_1732_0 & ~i_8_117_1806_0 & ~i_8_117_1945_0) | (~i_8_117_459_0 & ~i_8_117_461_0 & ~i_8_117_496_0 & ~i_8_117_792_0 & ~i_8_117_880_0 & ~i_8_117_1607_0 & ~i_8_117_1736_0 & ~i_8_117_1802_0 & ~i_8_117_1948_0 & ~i_8_117_1951_0))) | (~i_8_117_1607_0 & ((~i_8_117_366_0 & ~i_8_117_459_0 & ~i_8_117_461_0 & ~i_8_117_469_0 & ((~i_8_117_422_0 & ~i_8_117_492_0 & ~i_8_117_657_0 & ~i_8_117_709_0 & ~i_8_117_804_0 & ~i_8_117_878_0 & ~i_8_117_1609_0 & ~i_8_117_1610_0 & ~i_8_117_1945_0) | (~i_8_117_326_0 & ~i_8_117_472_0 & ~i_8_117_792_0 & ~i_8_117_1886_0 & ~i_8_117_1964_0 & ~i_8_117_2152_0 & ~i_8_117_1946_0 & ~i_8_117_1951_0))) | (~i_8_117_325_0 & ~i_8_117_472_0 & ~i_8_117_496_0 & ~i_8_117_657_0 & ~i_8_117_658_0 & ~i_8_117_795_0 & ~i_8_117_1078_0 & ~i_8_117_1410_0 & ~i_8_117_1471_0 & ~i_8_117_1608_0 & ~i_8_117_1787_0 & ~i_8_117_1806_0 & ~i_8_117_1946_0 & ~i_8_117_1948_0 & ~i_8_117_1970_0))))) | (~i_8_117_459_0 & ((i_8_117_469_0 & ~i_8_117_475_0 & ~i_8_117_795_0 & ~i_8_117_878_0 & ~i_8_117_1111_0 & ~i_8_117_1732_0 & ~i_8_117_1860_0 & ~i_8_117_1946_0 & ~i_8_117_1951_0 & ~i_8_117_1992_0 & ~i_8_117_2137_0) | (~i_8_117_140_0 & ~i_8_117_469_0 & ~i_8_117_474_0 & ~i_8_117_1078_0 & ~i_8_117_1159_0 & i_8_117_1480_0 & ~i_8_117_2152_0))) | (~i_8_117_1607_0 & ~i_8_117_1951_0 & ((~i_8_117_472_0 & ~i_8_117_475_0 & ~i_8_117_657_0 & ~i_8_117_993_0 & ~i_8_117_1114_0 & ~i_8_117_1747_0 & ~i_8_117_1945_0 & ~i_8_117_1948_0 & ~i_8_117_1964_0) | (~i_8_117_461_0 & ~i_8_117_474_0 & ~i_8_117_792_0 & ~i_8_117_1608_0 & i_8_117_1677_0 & ~i_8_117_1805_0 & ~i_8_117_1856_0 & ~i_8_117_1860_0 & ~i_8_117_1946_0 & ~i_8_117_2152_0 & ~i_8_117_2153_0))) | (~i_8_117_136_0 & ~i_8_117_420_0 & ~i_8_117_422_0 & ~i_8_117_592_0 & i_8_117_709_0 & ~i_8_117_880_0 & ~i_8_117_1185_0 & ~i_8_117_1610_0 & ~i_8_117_1856_0 & ~i_8_117_1945_0 & ~i_8_117_1948_0 & ~i_8_117_2153_0))) | (~i_8_117_1747_0 & ((~i_8_117_1945_0 & ((i_8_117_109_0 & ((~i_8_117_792_0 & ~i_8_117_1230_0 & i_8_117_1279_0 & ~i_8_117_1753_0 & ~i_8_117_1904_0 & ~i_8_117_1946_0 & ~i_8_117_1948_0 & ~i_8_117_1949_0) | (~i_8_117_136_0 & ~i_8_117_461_0 & ~i_8_117_474_0 & ~i_8_117_592_0 & ~i_8_117_1279_0 & ~i_8_117_1471_0 & ~i_8_117_1482_0 & ~i_8_117_1524_0 & ~i_8_117_1951_0 & ~i_8_117_2158_0))) | (~i_8_117_993_0 & ((~i_8_117_23_0 & ~i_8_117_325_0 & ~i_8_117_1609_0 & i_8_117_1736_0 & ~i_8_117_2137_0) | (~i_8_117_385_0 & ~i_8_117_469_0 & ~i_8_117_475_0 & ~i_8_117_1111_0 & ~i_8_117_1114_0 & ~i_8_117_1608_0 & ~i_8_117_1677_0 & ~i_8_117_1948_0 & ~i_8_117_1967_0 & ~i_8_117_2109_0 & ~i_8_117_2226_0))) | (~i_8_117_1230_0 & i_8_117_1524_0 & ~i_8_117_1736_0 & ~i_8_117_1946_0 & ~i_8_117_1949_0 & ~i_8_117_1964_0))) | (~i_8_117_1949_0 & ((i_8_117_325_0 & ~i_8_117_421_0 & ~i_8_117_469_0 & ~i_8_117_1111_0 & ~i_8_117_1946_0) | (~i_8_117_109_0 & ~i_8_117_139_0 & ~i_8_117_795_0 & ~i_8_117_880_0 & ~i_8_117_1114_0 & ~i_8_117_1608_0 & ~i_8_117_1753_0 & ~i_8_117_1948_0 & ~i_8_117_1964_0 & ~i_8_117_1970_0 & ~i_8_117_1992_0 & ~i_8_117_2153_0))) | (~i_8_117_22_0 & i_8_117_877_0 & i_8_117_1901_0))) | (~i_8_117_472_0 & ((~i_8_117_326_0 & ~i_8_117_1114_0 & ~i_8_117_1967_0 & ((~i_8_117_109_0 & ~i_8_117_420_0 & ~i_8_117_496_0 & ~i_8_117_1279_0 & ~i_8_117_1437_0 & ~i_8_117_1610_0 & ~i_8_117_1802_0 & ~i_8_117_1945_0 & ~i_8_117_1951_0) | (~i_8_117_461_0 & i_8_117_878_0 & ~i_8_117_1805_0 & ~i_8_117_1949_0 & ~i_8_117_2109_0 & ~i_8_117_2137_0 & ~i_8_117_2153_0))) | (~i_8_117_23_0 & ~i_8_117_459_0 & ~i_8_117_475_0 & i_8_117_1114_0 & ~i_8_117_1609_0 & ~i_8_117_1610_0 & i_8_117_1732_0 & ~i_8_117_2109_0) | (i_8_117_143_0 & ~i_8_117_420_0 & ~i_8_117_461_0 & ~i_8_117_474_0 & ~i_8_117_1608_0 & ~i_8_117_1886_0 & ~i_8_117_1949_0) | (~i_8_117_1948_0 & ~i_8_117_1951_0 & i_8_117_1904_0 & ~i_8_117_1946_0))) | (i_8_117_420_0 & ((i_8_117_1903_0 & ~i_8_117_1967_0) | (~i_8_117_1948_0 & ~i_8_117_1949_0 & ~i_8_117_1951_0 & ~i_8_117_2109_0 & ~i_8_117_2152_0 & ~i_8_117_2158_0))) | (~i_8_117_1607_0 & ((~i_8_117_109_0 & ~i_8_117_1608_0 & ((~i_8_117_23_0 & ~i_8_117_474_0 & ~i_8_117_496_0 & ~i_8_117_1159_0 & ~i_8_117_1410_0 & ~i_8_117_1787_0 & ~i_8_117_1802_0 & i_8_117_1886_0 & ~i_8_117_1949_0 & ~i_8_117_1970_0) | (~i_8_117_22_0 & ~i_8_117_385_0 & ~i_8_117_461_0 & ~i_8_117_469_0 & ~i_8_117_817_0 & i_8_117_878_0 & ~i_8_117_1114_0 & ~i_8_117_1856_0 & ~i_8_117_2153_0 & ~i_8_117_2156_0))) | (~i_8_117_461_0 & ~i_8_117_474_0 & ~i_8_117_475_0 & ~i_8_117_1471_0 & i_8_117_1652_0 & ~i_8_117_1860_0 & i_8_117_1992_0))) | (~i_8_117_23_0 & ~i_8_117_1078_0 & ((~i_8_117_459_0 & ~i_8_117_474_0 & ~i_8_117_575_0 & ~i_8_117_1159_0 & ~i_8_117_1393_0 & ~i_8_117_1410_0 & ~i_8_117_1609_0 & ~i_8_117_1610_0 & ~i_8_117_1677_0 & ~i_8_117_1806_0 & i_8_117_1886_0 & ~i_8_117_2156_0) | (~i_8_117_420_0 & ~i_8_117_592_0 & i_8_117_880_0 & ~i_8_117_1111_0 & ~i_8_117_1230_0 & ~i_8_117_1437_0 & ~i_8_117_1903_0 & ~i_8_117_1946_0 & ~i_8_117_1948_0 & ~i_8_117_1967_0 & ~i_8_117_2226_0))) | (~i_8_117_475_0 & ((~i_8_117_492_0 & ~i_8_117_2158_0 & ((~i_8_117_792_0 & ~i_8_117_878_0 & ~i_8_117_1609_0 & i_8_117_1725_0 & ~i_8_117_1805_0) | (~i_8_117_22_0 & ~i_8_117_109_0 & ~i_8_117_385_0 & ~i_8_117_446_0 & ~i_8_117_993_0 & ~i_8_117_1230_0 & ~i_8_117_1279_0 & ~i_8_117_1471_0 & ~i_8_117_1945_0 & ~i_8_117_1951_0 & ~i_8_117_1610_0 & ~i_8_117_1886_0 & ~i_8_117_2152_0 & ~i_8_117_2153_0 & ~i_8_117_1992_0 & ~i_8_117_2109_0))) | (~i_8_117_139_0 & i_8_117_326_0 & i_8_117_658_0 & ~i_8_117_709_0 & i_8_117_878_0 & ~i_8_117_1951_0))) | (~i_8_117_22_0 & ((i_8_117_592_0 & ~i_8_117_880_0 & i_8_117_1655_0 & i_8_117_1787_0 & ~i_8_117_1945_0) | (i_8_117_140_0 & ~i_8_117_496_0 & ~i_8_117_1609_0 & i_8_117_1992_0 & ~i_8_117_2109_0))) | (~i_8_117_385_0 & ((~i_8_117_366_0 & ~i_8_117_592_0 & ~i_8_117_658_0 & i_8_117_838_0 & ~i_8_117_878_0 & ~i_8_117_1471_0 & ~i_8_117_1970_0 & ~i_8_117_2109_0) | (~i_8_117_136_0 & ~i_8_117_496_0 & ~i_8_117_993_0 & i_8_117_1802_0 & i_8_117_1886_0 & ~i_8_117_1946_0 & ~i_8_117_1992_0 & ~i_8_117_2152_0))) | (~i_8_117_709_0 & ((~i_8_117_629_0 & ~i_8_117_792_0 & ~i_8_117_804_0 & i_8_117_838_0 & ~i_8_117_1410_0 & ~i_8_117_1608_0 & ~i_8_117_1725_0 & ~i_8_117_1753_0 & ~i_8_117_1802_0 & ~i_8_117_1946_0 & ~i_8_117_2152_0) | (~i_8_117_469_0 & ~i_8_117_1787_0 & ~i_8_117_1949_0 & i_8_117_2153_0 & i_8_117_2156_0))) | (~i_8_117_1111_0 & ((~i_8_117_474_0 & i_8_117_1437_0 & ~i_8_117_1471_0 & ~i_8_117_1609_0 & ~i_8_117_1806_0 & i_8_117_1860_0 & ~i_8_117_1946_0 & ~i_8_117_2156_0) | (i_8_117_1747_0 & i_8_117_2137_0 & i_8_117_2153_0 & ~i_8_117_2158_0))) | (i_8_117_838_0 & ~i_8_117_1608_0 & i_8_117_1802_0 & i_8_117_1856_0) | (~i_8_117_421_0 & i_8_117_1185_0 & i_8_117_1725_0 & ~i_8_117_2109_0) | (~i_8_117_1949_0 & i_8_117_1967_0 & ~i_8_117_2137_0 & i_8_117_2153_0 & i_8_117_2226_0));
endmodule



// Benchmark "kernel_8_118" written by ABC on Sun Jul 19 10:05:05 2020

module kernel_8_118 ( 
    i_8_118_31_0, i_8_118_84_0, i_8_118_96_0, i_8_118_161_0, i_8_118_192_0,
    i_8_118_224_0, i_8_118_293_0, i_8_118_300_0, i_8_118_301_0,
    i_8_118_368_0, i_8_118_373_0, i_8_118_378_0, i_8_118_379_0,
    i_8_118_381_0, i_8_118_383_0, i_8_118_384_0, i_8_118_386_0,
    i_8_118_394_0, i_8_118_421_0, i_8_118_422_0, i_8_118_446_0,
    i_8_118_456_0, i_8_118_462_0, i_8_118_483_0, i_8_118_493_0,
    i_8_118_494_0, i_8_118_500_0, i_8_118_556_0, i_8_118_588_0,
    i_8_118_593_0, i_8_118_660_0, i_8_118_661_0, i_8_118_673_0,
    i_8_118_715_0, i_8_118_718_0, i_8_118_781_0, i_8_118_783_0,
    i_8_118_795_0, i_8_118_796_0, i_8_118_826_0, i_8_118_827_0,
    i_8_118_842_0, i_8_118_878_0, i_8_118_1012_0, i_8_118_1029_0,
    i_8_118_1077_0, i_8_118_1115_0, i_8_118_1120_0, i_8_118_1156_0,
    i_8_118_1191_0, i_8_118_1228_0, i_8_118_1229_0, i_8_118_1255_0,
    i_8_118_1274_0, i_8_118_1300_0, i_8_118_1331_0, i_8_118_1345_0,
    i_8_118_1346_0, i_8_118_1438_0, i_8_118_1457_0, i_8_118_1471_0,
    i_8_118_1534_0, i_8_118_1535_0, i_8_118_1548_0, i_8_118_1587_0,
    i_8_118_1597_0, i_8_118_1598_0, i_8_118_1606_0, i_8_118_1648_0,
    i_8_118_1649_0, i_8_118_1705_0, i_8_118_1751_0, i_8_118_1763_0,
    i_8_118_1804_0, i_8_118_1807_0, i_8_118_1808_0, i_8_118_1812_0,
    i_8_118_1822_0, i_8_118_1841_0, i_8_118_1844_0, i_8_118_1894_0,
    i_8_118_1903_0, i_8_118_1952_0, i_8_118_1966_0, i_8_118_2110_0,
    i_8_118_2113_0, i_8_118_2127_0, i_8_118_2132_0, i_8_118_2136_0,
    i_8_118_2139_0, i_8_118_2158_0, i_8_118_2172_0, i_8_118_2182_0,
    i_8_118_2190_0, i_8_118_2191_0, i_8_118_2195_0, i_8_118_2216_0,
    i_8_118_2227_0, i_8_118_2273_0, i_8_118_2276_0,
    o_8_118_0_0  );
  input  i_8_118_31_0, i_8_118_84_0, i_8_118_96_0, i_8_118_161_0,
    i_8_118_192_0, i_8_118_224_0, i_8_118_293_0, i_8_118_300_0,
    i_8_118_301_0, i_8_118_368_0, i_8_118_373_0, i_8_118_378_0,
    i_8_118_379_0, i_8_118_381_0, i_8_118_383_0, i_8_118_384_0,
    i_8_118_386_0, i_8_118_394_0, i_8_118_421_0, i_8_118_422_0,
    i_8_118_446_0, i_8_118_456_0, i_8_118_462_0, i_8_118_483_0,
    i_8_118_493_0, i_8_118_494_0, i_8_118_500_0, i_8_118_556_0,
    i_8_118_588_0, i_8_118_593_0, i_8_118_660_0, i_8_118_661_0,
    i_8_118_673_0, i_8_118_715_0, i_8_118_718_0, i_8_118_781_0,
    i_8_118_783_0, i_8_118_795_0, i_8_118_796_0, i_8_118_826_0,
    i_8_118_827_0, i_8_118_842_0, i_8_118_878_0, i_8_118_1012_0,
    i_8_118_1029_0, i_8_118_1077_0, i_8_118_1115_0, i_8_118_1120_0,
    i_8_118_1156_0, i_8_118_1191_0, i_8_118_1228_0, i_8_118_1229_0,
    i_8_118_1255_0, i_8_118_1274_0, i_8_118_1300_0, i_8_118_1331_0,
    i_8_118_1345_0, i_8_118_1346_0, i_8_118_1438_0, i_8_118_1457_0,
    i_8_118_1471_0, i_8_118_1534_0, i_8_118_1535_0, i_8_118_1548_0,
    i_8_118_1587_0, i_8_118_1597_0, i_8_118_1598_0, i_8_118_1606_0,
    i_8_118_1648_0, i_8_118_1649_0, i_8_118_1705_0, i_8_118_1751_0,
    i_8_118_1763_0, i_8_118_1804_0, i_8_118_1807_0, i_8_118_1808_0,
    i_8_118_1812_0, i_8_118_1822_0, i_8_118_1841_0, i_8_118_1844_0,
    i_8_118_1894_0, i_8_118_1903_0, i_8_118_1952_0, i_8_118_1966_0,
    i_8_118_2110_0, i_8_118_2113_0, i_8_118_2127_0, i_8_118_2132_0,
    i_8_118_2136_0, i_8_118_2139_0, i_8_118_2158_0, i_8_118_2172_0,
    i_8_118_2182_0, i_8_118_2190_0, i_8_118_2191_0, i_8_118_2195_0,
    i_8_118_2216_0, i_8_118_2227_0, i_8_118_2273_0, i_8_118_2276_0;
  output o_8_118_0_0;
  assign o_8_118_0_0 = 0;
endmodule



// Benchmark "kernel_8_119" written by ABC on Sun Jul 19 10:05:05 2020

module kernel_8_119 ( 
    i_8_119_50_0, i_8_119_139_0, i_8_119_224_0, i_8_119_225_0,
    i_8_119_230_0, i_8_119_323_0, i_8_119_363_0, i_8_119_365_0,
    i_8_119_385_0, i_8_119_394_0, i_8_119_402_0, i_8_119_403_0,
    i_8_119_489_0, i_8_119_550_0, i_8_119_554_0, i_8_119_569_0,
    i_8_119_604_0, i_8_119_606_0, i_8_119_626_0, i_8_119_632_0,
    i_8_119_638_0, i_8_119_644_0, i_8_119_664_0, i_8_119_665_0,
    i_8_119_675_0, i_8_119_679_0, i_8_119_697_0, i_8_119_700_0,
    i_8_119_781_0, i_8_119_785_0, i_8_119_823_0, i_8_119_833_0,
    i_8_119_839_0, i_8_119_858_0, i_8_119_873_0, i_8_119_876_0,
    i_8_119_893_0, i_8_119_898_0, i_8_119_959_0, i_8_119_968_0,
    i_8_119_992_0, i_8_119_1034_0, i_8_119_1040_0, i_8_119_1073_0,
    i_8_119_1094_0, i_8_119_1134_0, i_8_119_1137_0, i_8_119_1150_0,
    i_8_119_1202_0, i_8_119_1232_0, i_8_119_1264_0, i_8_119_1328_0,
    i_8_119_1340_0, i_8_119_1349_0, i_8_119_1366_0, i_8_119_1367_0,
    i_8_119_1372_0, i_8_119_1404_0, i_8_119_1436_0, i_8_119_1451_0,
    i_8_119_1465_0, i_8_119_1481_0, i_8_119_1490_0, i_8_119_1557_0,
    i_8_119_1558_0, i_8_119_1573_0, i_8_119_1629_0, i_8_119_1633_0,
    i_8_119_1634_0, i_8_119_1700_0, i_8_119_1704_0, i_8_119_1705_0,
    i_8_119_1709_0, i_8_119_1727_0, i_8_119_1733_0, i_8_119_1771_0,
    i_8_119_1772_0, i_8_119_1824_0, i_8_119_1825_0, i_8_119_1826_0,
    i_8_119_1884_0, i_8_119_1886_0, i_8_119_1888_0, i_8_119_1939_0,
    i_8_119_1940_0, i_8_119_1944_0, i_8_119_1960_0, i_8_119_1981_0,
    i_8_119_1997_0, i_8_119_2142_0, i_8_119_2155_0, i_8_119_2157_0,
    i_8_119_2225_0, i_8_119_2226_0, i_8_119_2231_0, i_8_119_2241_0,
    i_8_119_2248_0, i_8_119_2262_0, i_8_119_2282_0, i_8_119_2289_0,
    o_8_119_0_0  );
  input  i_8_119_50_0, i_8_119_139_0, i_8_119_224_0, i_8_119_225_0,
    i_8_119_230_0, i_8_119_323_0, i_8_119_363_0, i_8_119_365_0,
    i_8_119_385_0, i_8_119_394_0, i_8_119_402_0, i_8_119_403_0,
    i_8_119_489_0, i_8_119_550_0, i_8_119_554_0, i_8_119_569_0,
    i_8_119_604_0, i_8_119_606_0, i_8_119_626_0, i_8_119_632_0,
    i_8_119_638_0, i_8_119_644_0, i_8_119_664_0, i_8_119_665_0,
    i_8_119_675_0, i_8_119_679_0, i_8_119_697_0, i_8_119_700_0,
    i_8_119_781_0, i_8_119_785_0, i_8_119_823_0, i_8_119_833_0,
    i_8_119_839_0, i_8_119_858_0, i_8_119_873_0, i_8_119_876_0,
    i_8_119_893_0, i_8_119_898_0, i_8_119_959_0, i_8_119_968_0,
    i_8_119_992_0, i_8_119_1034_0, i_8_119_1040_0, i_8_119_1073_0,
    i_8_119_1094_0, i_8_119_1134_0, i_8_119_1137_0, i_8_119_1150_0,
    i_8_119_1202_0, i_8_119_1232_0, i_8_119_1264_0, i_8_119_1328_0,
    i_8_119_1340_0, i_8_119_1349_0, i_8_119_1366_0, i_8_119_1367_0,
    i_8_119_1372_0, i_8_119_1404_0, i_8_119_1436_0, i_8_119_1451_0,
    i_8_119_1465_0, i_8_119_1481_0, i_8_119_1490_0, i_8_119_1557_0,
    i_8_119_1558_0, i_8_119_1573_0, i_8_119_1629_0, i_8_119_1633_0,
    i_8_119_1634_0, i_8_119_1700_0, i_8_119_1704_0, i_8_119_1705_0,
    i_8_119_1709_0, i_8_119_1727_0, i_8_119_1733_0, i_8_119_1771_0,
    i_8_119_1772_0, i_8_119_1824_0, i_8_119_1825_0, i_8_119_1826_0,
    i_8_119_1884_0, i_8_119_1886_0, i_8_119_1888_0, i_8_119_1939_0,
    i_8_119_1940_0, i_8_119_1944_0, i_8_119_1960_0, i_8_119_1981_0,
    i_8_119_1997_0, i_8_119_2142_0, i_8_119_2155_0, i_8_119_2157_0,
    i_8_119_2225_0, i_8_119_2226_0, i_8_119_2231_0, i_8_119_2241_0,
    i_8_119_2248_0, i_8_119_2262_0, i_8_119_2282_0, i_8_119_2289_0;
  output o_8_119_0_0;
  assign o_8_119_0_0 = 0;
endmodule



// Benchmark "kernel_8_120" written by ABC on Sun Jul 19 10:05:07 2020

module kernel_8_120 ( 
    i_8_120_18_0, i_8_120_19_0, i_8_120_29_0, i_8_120_32_0, i_8_120_83_0,
    i_8_120_95_0, i_8_120_98_0, i_8_120_109_0, i_8_120_112_0,
    i_8_120_116_0, i_8_120_142_0, i_8_120_143_0, i_8_120_163_0,
    i_8_120_164_0, i_8_120_166_0, i_8_120_218_0, i_8_120_221_0,
    i_8_120_239_0, i_8_120_241_0, i_8_120_299_0, i_8_120_331_0,
    i_8_120_344_0, i_8_120_360_0, i_8_120_381_0, i_8_120_479_0,
    i_8_120_481_0, i_8_120_484_0, i_8_120_504_0, i_8_120_526_0,
    i_8_120_591_0, i_8_120_598_0, i_8_120_602_0, i_8_120_605_0,
    i_8_120_614_0, i_8_120_632_0, i_8_120_686_0, i_8_120_701_0,
    i_8_120_702_0, i_8_120_704_0, i_8_120_707_0, i_8_120_713_0,
    i_8_120_737_0, i_8_120_812_0, i_8_120_878_0, i_8_120_921_0,
    i_8_120_938_0, i_8_120_997_0, i_8_120_998_0, i_8_120_1012_0,
    i_8_120_1045_0, i_8_120_1048_0, i_8_120_1058_0, i_8_120_1091_0,
    i_8_120_1107_0, i_8_120_1117_0, i_8_120_1181_0, i_8_120_1235_0,
    i_8_120_1262_0, i_8_120_1265_0, i_8_120_1280_0, i_8_120_1282_0,
    i_8_120_1306_0, i_8_120_1355_0, i_8_120_1412_0, i_8_120_1434_0,
    i_8_120_1462_0, i_8_120_1534_0, i_8_120_1574_0, i_8_120_1586_0,
    i_8_120_1594_0, i_8_120_1679_0, i_8_120_1694_0, i_8_120_1696_0,
    i_8_120_1697_0, i_8_120_1724_0, i_8_120_1729_0, i_8_120_1739_0,
    i_8_120_1751_0, i_8_120_1754_0, i_8_120_1757_0, i_8_120_1804_0,
    i_8_120_1805_0, i_8_120_1814_0, i_8_120_1829_0, i_8_120_1856_0,
    i_8_120_1858_0, i_8_120_1867_0, i_8_120_1993_0, i_8_120_2036_0,
    i_8_120_2038_0, i_8_120_2039_0, i_8_120_2045_0, i_8_120_2047_0,
    i_8_120_2078_0, i_8_120_2096_0, i_8_120_2105_0, i_8_120_2117_0,
    i_8_120_2146_0, i_8_120_2187_0, i_8_120_2246_0,
    o_8_120_0_0  );
  input  i_8_120_18_0, i_8_120_19_0, i_8_120_29_0, i_8_120_32_0,
    i_8_120_83_0, i_8_120_95_0, i_8_120_98_0, i_8_120_109_0, i_8_120_112_0,
    i_8_120_116_0, i_8_120_142_0, i_8_120_143_0, i_8_120_163_0,
    i_8_120_164_0, i_8_120_166_0, i_8_120_218_0, i_8_120_221_0,
    i_8_120_239_0, i_8_120_241_0, i_8_120_299_0, i_8_120_331_0,
    i_8_120_344_0, i_8_120_360_0, i_8_120_381_0, i_8_120_479_0,
    i_8_120_481_0, i_8_120_484_0, i_8_120_504_0, i_8_120_526_0,
    i_8_120_591_0, i_8_120_598_0, i_8_120_602_0, i_8_120_605_0,
    i_8_120_614_0, i_8_120_632_0, i_8_120_686_0, i_8_120_701_0,
    i_8_120_702_0, i_8_120_704_0, i_8_120_707_0, i_8_120_713_0,
    i_8_120_737_0, i_8_120_812_0, i_8_120_878_0, i_8_120_921_0,
    i_8_120_938_0, i_8_120_997_0, i_8_120_998_0, i_8_120_1012_0,
    i_8_120_1045_0, i_8_120_1048_0, i_8_120_1058_0, i_8_120_1091_0,
    i_8_120_1107_0, i_8_120_1117_0, i_8_120_1181_0, i_8_120_1235_0,
    i_8_120_1262_0, i_8_120_1265_0, i_8_120_1280_0, i_8_120_1282_0,
    i_8_120_1306_0, i_8_120_1355_0, i_8_120_1412_0, i_8_120_1434_0,
    i_8_120_1462_0, i_8_120_1534_0, i_8_120_1574_0, i_8_120_1586_0,
    i_8_120_1594_0, i_8_120_1679_0, i_8_120_1694_0, i_8_120_1696_0,
    i_8_120_1697_0, i_8_120_1724_0, i_8_120_1729_0, i_8_120_1739_0,
    i_8_120_1751_0, i_8_120_1754_0, i_8_120_1757_0, i_8_120_1804_0,
    i_8_120_1805_0, i_8_120_1814_0, i_8_120_1829_0, i_8_120_1856_0,
    i_8_120_1858_0, i_8_120_1867_0, i_8_120_1993_0, i_8_120_2036_0,
    i_8_120_2038_0, i_8_120_2039_0, i_8_120_2045_0, i_8_120_2047_0,
    i_8_120_2078_0, i_8_120_2096_0, i_8_120_2105_0, i_8_120_2117_0,
    i_8_120_2146_0, i_8_120_2187_0, i_8_120_2246_0;
  output o_8_120_0_0;
  assign o_8_120_0_0 = ~((~i_8_120_29_0 & ((~i_8_120_164_0 & ~i_8_120_591_0 & ~i_8_120_602_0 & ~i_8_120_632_0 & ~i_8_120_938_0 & ~i_8_120_1181_0) | (~i_8_120_142_0 & i_8_120_239_0 & ~i_8_120_713_0 & ~i_8_120_812_0 & ~i_8_120_2117_0))) | (~i_8_120_32_0 & ((~i_8_120_812_0 & ~i_8_120_998_0 & ~i_8_120_1117_0 & i_8_120_1265_0 & ~i_8_120_1694_0 & ~i_8_120_1858_0) | (i_8_120_299_0 & ~i_8_120_331_0 & ~i_8_120_686_0 & i_8_120_1694_0 & ~i_8_120_2117_0))) | (~i_8_120_83_0 & ((~i_8_120_163_0 & ~i_8_120_164_0 & ~i_8_120_713_0 & ~i_8_120_1574_0 & ~i_8_120_1586_0) | (~i_8_120_112_0 & ~i_8_120_166_0 & ~i_8_120_632_0 & ~i_8_120_1757_0 & ~i_8_120_2039_0))) | (i_8_120_109_0 & ((~i_8_120_19_0 & ~i_8_120_166_0 & ~i_8_120_602_0 & ~i_8_120_713_0 & ~i_8_120_1265_0 & ~i_8_120_1757_0) | (i_8_120_713_0 & ~i_8_120_737_0 & ~i_8_120_2045_0 & i_8_120_2146_0))) | (~i_8_120_299_0 & ((~i_8_120_479_0 & ~i_8_120_591_0 & ~i_8_120_938_0 & ~i_8_120_1181_0 & ~i_8_120_1412_0 & ~i_8_120_1694_0 & ~i_8_120_1856_0) | (~i_8_120_632_0 & i_8_120_1804_0 & ~i_8_120_2246_0))) | (i_8_120_481_0 & ((~i_8_120_1262_0 & ~i_8_120_1355_0 & i_8_120_1679_0 & ~i_8_120_2036_0 & ~i_8_120_2096_0) | (~i_8_120_218_0 & ~i_8_120_1757_0 & ~i_8_120_2039_0 & ~i_8_120_2146_0))) | (~i_8_120_1829_0 & ((~i_8_120_1586_0 & ((~i_8_120_331_0 & ~i_8_120_1181_0 & ~i_8_120_1355_0 & ~i_8_120_1858_0) | (~i_8_120_1739_0 & i_8_120_1867_0))) | (~i_8_120_164_0 & ~i_8_120_239_0 & ~i_8_120_1739_0 & ~i_8_120_2096_0 & ~i_8_120_2117_0))) | (~i_8_120_164_0 & ~i_8_120_2039_0 & ((~i_8_120_98_0 & ~i_8_120_632_0 & ~i_8_120_686_0 & ~i_8_120_1412_0) | (~i_8_120_142_0 & i_8_120_218_0 & ~i_8_120_1754_0 & ~i_8_120_2038_0 & ~i_8_120_2246_0))) | (~i_8_120_632_0 & ((~i_8_120_713_0 & ~i_8_120_1058_0 & ~i_8_120_1235_0 & ~i_8_120_1262_0) | (~i_8_120_1181_0 & ~i_8_120_1574_0 & ~i_8_120_1586_0 & ~i_8_120_1805_0 & ~i_8_120_2105_0 & ~i_8_120_2117_0))) | (i_8_120_98_0 & i_8_120_704_0) | (~i_8_120_166_0 & ~i_8_120_938_0 & ~i_8_120_1045_0 & ~i_8_120_1091_0 & ~i_8_120_1181_0 & ~i_8_120_1265_0 & ~i_8_120_1280_0 & ~i_8_120_1805_0) | (~i_8_120_591_0 & i_8_120_707_0 & ~i_8_120_1117_0 & ~i_8_120_1856_0 & ~i_8_120_2045_0));
endmodule



// Benchmark "kernel_8_121" written by ABC on Sun Jul 19 10:05:08 2020

module kernel_8_121 ( 
    i_8_121_106_0, i_8_121_164_0, i_8_121_166_0, i_8_121_173_0,
    i_8_121_179_0, i_8_121_212_0, i_8_121_253_0, i_8_121_284_0,
    i_8_121_293_0, i_8_121_356_0, i_8_121_365_0, i_8_121_368_0,
    i_8_121_378_0, i_8_121_419_0, i_8_121_430_0, i_8_121_440_0,
    i_8_121_453_0, i_8_121_457_0, i_8_121_473_0, i_8_121_478_0,
    i_8_121_479_0, i_8_121_508_0, i_8_121_535_0, i_8_121_539_0,
    i_8_121_545_0, i_8_121_593_0, i_8_121_599_0, i_8_121_617_0,
    i_8_121_659_0, i_8_121_698_0, i_8_121_742_0, i_8_121_760_0,
    i_8_121_764_0, i_8_121_809_0, i_8_121_827_0, i_8_121_833_0,
    i_8_121_839_0, i_8_121_850_0, i_8_121_868_0, i_8_121_881_0,
    i_8_121_910_0, i_8_121_922_0, i_8_121_940_0, i_8_121_977_0,
    i_8_121_1045_0, i_8_121_1067_0, i_8_121_1075_0, i_8_121_1171_0,
    i_8_121_1208_0, i_8_121_1259_0, i_8_121_1264_0, i_8_121_1282_0,
    i_8_121_1344_0, i_8_121_1401_0, i_8_121_1417_0, i_8_121_1444_0,
    i_8_121_1454_0, i_8_121_1462_0, i_8_121_1508_0, i_8_121_1553_0,
    i_8_121_1574_0, i_8_121_1597_0, i_8_121_1640_0, i_8_121_1648_0,
    i_8_121_1666_0, i_8_121_1680_0, i_8_121_1702_0, i_8_121_1707_0,
    i_8_121_1731_0, i_8_121_1760_0, i_8_121_1779_0, i_8_121_1823_0,
    i_8_121_1826_0, i_8_121_1895_0, i_8_121_1903_0, i_8_121_1907_0,
    i_8_121_1920_0, i_8_121_1931_0, i_8_121_1993_0, i_8_121_1995_0,
    i_8_121_1996_0, i_8_121_2012_0, i_8_121_2117_0, i_8_121_2134_0,
    i_8_121_2137_0, i_8_121_2145_0, i_8_121_2146_0, i_8_121_2153_0,
    i_8_121_2156_0, i_8_121_2182_0, i_8_121_2185_0, i_8_121_2207_0,
    i_8_121_2210_0, i_8_121_2213_0, i_8_121_2215_0, i_8_121_2227_0,
    i_8_121_2245_0, i_8_121_2284_0, i_8_121_2288_0, i_8_121_2293_0,
    o_8_121_0_0  );
  input  i_8_121_106_0, i_8_121_164_0, i_8_121_166_0, i_8_121_173_0,
    i_8_121_179_0, i_8_121_212_0, i_8_121_253_0, i_8_121_284_0,
    i_8_121_293_0, i_8_121_356_0, i_8_121_365_0, i_8_121_368_0,
    i_8_121_378_0, i_8_121_419_0, i_8_121_430_0, i_8_121_440_0,
    i_8_121_453_0, i_8_121_457_0, i_8_121_473_0, i_8_121_478_0,
    i_8_121_479_0, i_8_121_508_0, i_8_121_535_0, i_8_121_539_0,
    i_8_121_545_0, i_8_121_593_0, i_8_121_599_0, i_8_121_617_0,
    i_8_121_659_0, i_8_121_698_0, i_8_121_742_0, i_8_121_760_0,
    i_8_121_764_0, i_8_121_809_0, i_8_121_827_0, i_8_121_833_0,
    i_8_121_839_0, i_8_121_850_0, i_8_121_868_0, i_8_121_881_0,
    i_8_121_910_0, i_8_121_922_0, i_8_121_940_0, i_8_121_977_0,
    i_8_121_1045_0, i_8_121_1067_0, i_8_121_1075_0, i_8_121_1171_0,
    i_8_121_1208_0, i_8_121_1259_0, i_8_121_1264_0, i_8_121_1282_0,
    i_8_121_1344_0, i_8_121_1401_0, i_8_121_1417_0, i_8_121_1444_0,
    i_8_121_1454_0, i_8_121_1462_0, i_8_121_1508_0, i_8_121_1553_0,
    i_8_121_1574_0, i_8_121_1597_0, i_8_121_1640_0, i_8_121_1648_0,
    i_8_121_1666_0, i_8_121_1680_0, i_8_121_1702_0, i_8_121_1707_0,
    i_8_121_1731_0, i_8_121_1760_0, i_8_121_1779_0, i_8_121_1823_0,
    i_8_121_1826_0, i_8_121_1895_0, i_8_121_1903_0, i_8_121_1907_0,
    i_8_121_1920_0, i_8_121_1931_0, i_8_121_1993_0, i_8_121_1995_0,
    i_8_121_1996_0, i_8_121_2012_0, i_8_121_2117_0, i_8_121_2134_0,
    i_8_121_2137_0, i_8_121_2145_0, i_8_121_2146_0, i_8_121_2153_0,
    i_8_121_2156_0, i_8_121_2182_0, i_8_121_2185_0, i_8_121_2207_0,
    i_8_121_2210_0, i_8_121_2213_0, i_8_121_2215_0, i_8_121_2227_0,
    i_8_121_2245_0, i_8_121_2284_0, i_8_121_2288_0, i_8_121_2293_0;
  output o_8_121_0_0;
  assign o_8_121_0_0 = 0;
endmodule



// Benchmark "kernel_8_122" written by ABC on Sun Jul 19 10:05:08 2020

module kernel_8_122 ( 
    i_8_122_57_0, i_8_122_61_0, i_8_122_88_0, i_8_122_96_0, i_8_122_104_0,
    i_8_122_160_0, i_8_122_168_0, i_8_122_169_0, i_8_122_170_0,
    i_8_122_191_0, i_8_122_220_0, i_8_122_232_0, i_8_122_255_0,
    i_8_122_258_0, i_8_122_292_0, i_8_122_303_0, i_8_122_304_0,
    i_8_122_313_0, i_8_122_321_0, i_8_122_328_0, i_8_122_364_0,
    i_8_122_385_0, i_8_122_393_0, i_8_122_417_0, i_8_122_420_0,
    i_8_122_421_0, i_8_122_439_0, i_8_122_440_0, i_8_122_447_0,
    i_8_122_493_0, i_8_122_498_0, i_8_122_522_0, i_8_122_523_0,
    i_8_122_555_0, i_8_122_570_0, i_8_122_597_0, i_8_122_601_0,
    i_8_122_602_0, i_8_122_617_0, i_8_122_624_0, i_8_122_687_0,
    i_8_122_690_0, i_8_122_727_0, i_8_122_786_0, i_8_122_789_0,
    i_8_122_849_0, i_8_122_850_0, i_8_122_856_0, i_8_122_858_0,
    i_8_122_990_0, i_8_122_993_0, i_8_122_996_0, i_8_122_1050_0,
    i_8_122_1071_0, i_8_122_1075_0, i_8_122_1116_0, i_8_122_1122_0,
    i_8_122_1135_0, i_8_122_1188_0, i_8_122_1191_0, i_8_122_1222_0,
    i_8_122_1299_0, i_8_122_1305_0, i_8_122_1306_0, i_8_122_1307_0,
    i_8_122_1314_0, i_8_122_1318_0, i_8_122_1329_0, i_8_122_1346_0,
    i_8_122_1348_0, i_8_122_1470_0, i_8_122_1506_0, i_8_122_1509_0,
    i_8_122_1533_0, i_8_122_1536_0, i_8_122_1545_0, i_8_122_1561_0,
    i_8_122_1564_0, i_8_122_1570_0, i_8_122_1571_0, i_8_122_1574_0,
    i_8_122_1650_0, i_8_122_1651_0, i_8_122_1653_0, i_8_122_1681_0,
    i_8_122_1719_0, i_8_122_1727_0, i_8_122_1747_0, i_8_122_1750_0,
    i_8_122_1753_0, i_8_122_1795_0, i_8_122_1816_0, i_8_122_1956_0,
    i_8_122_1995_0, i_8_122_2031_0, i_8_122_2065_0, i_8_122_2122_0,
    i_8_122_2215_0, i_8_122_2226_0, i_8_122_2275_0,
    o_8_122_0_0  );
  input  i_8_122_57_0, i_8_122_61_0, i_8_122_88_0, i_8_122_96_0,
    i_8_122_104_0, i_8_122_160_0, i_8_122_168_0, i_8_122_169_0,
    i_8_122_170_0, i_8_122_191_0, i_8_122_220_0, i_8_122_232_0,
    i_8_122_255_0, i_8_122_258_0, i_8_122_292_0, i_8_122_303_0,
    i_8_122_304_0, i_8_122_313_0, i_8_122_321_0, i_8_122_328_0,
    i_8_122_364_0, i_8_122_385_0, i_8_122_393_0, i_8_122_417_0,
    i_8_122_420_0, i_8_122_421_0, i_8_122_439_0, i_8_122_440_0,
    i_8_122_447_0, i_8_122_493_0, i_8_122_498_0, i_8_122_522_0,
    i_8_122_523_0, i_8_122_555_0, i_8_122_570_0, i_8_122_597_0,
    i_8_122_601_0, i_8_122_602_0, i_8_122_617_0, i_8_122_624_0,
    i_8_122_687_0, i_8_122_690_0, i_8_122_727_0, i_8_122_786_0,
    i_8_122_789_0, i_8_122_849_0, i_8_122_850_0, i_8_122_856_0,
    i_8_122_858_0, i_8_122_990_0, i_8_122_993_0, i_8_122_996_0,
    i_8_122_1050_0, i_8_122_1071_0, i_8_122_1075_0, i_8_122_1116_0,
    i_8_122_1122_0, i_8_122_1135_0, i_8_122_1188_0, i_8_122_1191_0,
    i_8_122_1222_0, i_8_122_1299_0, i_8_122_1305_0, i_8_122_1306_0,
    i_8_122_1307_0, i_8_122_1314_0, i_8_122_1318_0, i_8_122_1329_0,
    i_8_122_1346_0, i_8_122_1348_0, i_8_122_1470_0, i_8_122_1506_0,
    i_8_122_1509_0, i_8_122_1533_0, i_8_122_1536_0, i_8_122_1545_0,
    i_8_122_1561_0, i_8_122_1564_0, i_8_122_1570_0, i_8_122_1571_0,
    i_8_122_1574_0, i_8_122_1650_0, i_8_122_1651_0, i_8_122_1653_0,
    i_8_122_1681_0, i_8_122_1719_0, i_8_122_1727_0, i_8_122_1747_0,
    i_8_122_1750_0, i_8_122_1753_0, i_8_122_1795_0, i_8_122_1816_0,
    i_8_122_1956_0, i_8_122_1995_0, i_8_122_2031_0, i_8_122_2065_0,
    i_8_122_2122_0, i_8_122_2215_0, i_8_122_2226_0, i_8_122_2275_0;
  output o_8_122_0_0;
  assign o_8_122_0_0 = 0;
endmodule



// Benchmark "kernel_8_123" written by ABC on Sun Jul 19 10:05:10 2020

module kernel_8_123 ( 
    i_8_123_23_0, i_8_123_41_0, i_8_123_72_0, i_8_123_73_0, i_8_123_88_0,
    i_8_123_107_0, i_8_123_118_0, i_8_123_119_0, i_8_123_167_0,
    i_8_123_226_0, i_8_123_258_0, i_8_123_269_0, i_8_123_308_0,
    i_8_123_348_0, i_8_123_349_0, i_8_123_350_0, i_8_123_381_0,
    i_8_123_382_0, i_8_123_440_0, i_8_123_489_0, i_8_123_490_0,
    i_8_123_506_0, i_8_123_585_0, i_8_123_608_0, i_8_123_628_0,
    i_8_123_630_0, i_8_123_631_0, i_8_123_686_0, i_8_123_709_0,
    i_8_123_710_0, i_8_123_727_0, i_8_123_728_0, i_8_123_748_0,
    i_8_123_814_0, i_8_123_826_0, i_8_123_828_0, i_8_123_830_0,
    i_8_123_838_0, i_8_123_873_0, i_8_123_881_0, i_8_123_956_0,
    i_8_123_977_0, i_8_123_980_0, i_8_123_981_0, i_8_123_982_0,
    i_8_123_991_0, i_8_123_1027_0, i_8_123_1028_0, i_8_123_1029_0,
    i_8_123_1030_0, i_8_123_1031_0, i_8_123_1040_0, i_8_123_1058_0,
    i_8_123_1078_0, i_8_123_1161_0, i_8_123_1162_0, i_8_123_1226_0,
    i_8_123_1262_0, i_8_123_1279_0, i_8_123_1281_0, i_8_123_1296_0,
    i_8_123_1297_0, i_8_123_1300_0, i_8_123_1315_0, i_8_123_1319_0,
    i_8_123_1325_0, i_8_123_1327_0, i_8_123_1330_0, i_8_123_1334_0,
    i_8_123_1355_0, i_8_123_1437_0, i_8_123_1449_0, i_8_123_1467_0,
    i_8_123_1470_0, i_8_123_1471_0, i_8_123_1474_0, i_8_123_1705_0,
    i_8_123_1729_0, i_8_123_1746_0, i_8_123_1764_0, i_8_123_1765_0,
    i_8_123_1780_0, i_8_123_1787_0, i_8_123_1813_0, i_8_123_1832_0,
    i_8_123_1862_0, i_8_123_1888_0, i_8_123_1889_0, i_8_123_1949_0,
    i_8_123_1952_0, i_8_123_1965_0, i_8_123_2052_0, i_8_123_2059_0,
    i_8_123_2079_0, i_8_123_2114_0, i_8_123_2126_0, i_8_123_2140_0,
    i_8_123_2158_0, i_8_123_2241_0, i_8_123_2243_0,
    o_8_123_0_0  );
  input  i_8_123_23_0, i_8_123_41_0, i_8_123_72_0, i_8_123_73_0,
    i_8_123_88_0, i_8_123_107_0, i_8_123_118_0, i_8_123_119_0,
    i_8_123_167_0, i_8_123_226_0, i_8_123_258_0, i_8_123_269_0,
    i_8_123_308_0, i_8_123_348_0, i_8_123_349_0, i_8_123_350_0,
    i_8_123_381_0, i_8_123_382_0, i_8_123_440_0, i_8_123_489_0,
    i_8_123_490_0, i_8_123_506_0, i_8_123_585_0, i_8_123_608_0,
    i_8_123_628_0, i_8_123_630_0, i_8_123_631_0, i_8_123_686_0,
    i_8_123_709_0, i_8_123_710_0, i_8_123_727_0, i_8_123_728_0,
    i_8_123_748_0, i_8_123_814_0, i_8_123_826_0, i_8_123_828_0,
    i_8_123_830_0, i_8_123_838_0, i_8_123_873_0, i_8_123_881_0,
    i_8_123_956_0, i_8_123_977_0, i_8_123_980_0, i_8_123_981_0,
    i_8_123_982_0, i_8_123_991_0, i_8_123_1027_0, i_8_123_1028_0,
    i_8_123_1029_0, i_8_123_1030_0, i_8_123_1031_0, i_8_123_1040_0,
    i_8_123_1058_0, i_8_123_1078_0, i_8_123_1161_0, i_8_123_1162_0,
    i_8_123_1226_0, i_8_123_1262_0, i_8_123_1279_0, i_8_123_1281_0,
    i_8_123_1296_0, i_8_123_1297_0, i_8_123_1300_0, i_8_123_1315_0,
    i_8_123_1319_0, i_8_123_1325_0, i_8_123_1327_0, i_8_123_1330_0,
    i_8_123_1334_0, i_8_123_1355_0, i_8_123_1437_0, i_8_123_1449_0,
    i_8_123_1467_0, i_8_123_1470_0, i_8_123_1471_0, i_8_123_1474_0,
    i_8_123_1705_0, i_8_123_1729_0, i_8_123_1746_0, i_8_123_1764_0,
    i_8_123_1765_0, i_8_123_1780_0, i_8_123_1787_0, i_8_123_1813_0,
    i_8_123_1832_0, i_8_123_1862_0, i_8_123_1888_0, i_8_123_1889_0,
    i_8_123_1949_0, i_8_123_1952_0, i_8_123_1965_0, i_8_123_2052_0,
    i_8_123_2059_0, i_8_123_2079_0, i_8_123_2114_0, i_8_123_2126_0,
    i_8_123_2140_0, i_8_123_2158_0, i_8_123_2241_0, i_8_123_2243_0;
  output o_8_123_0_0;
  assign o_8_123_0_0 = ~((~i_8_123_727_0 & ((~i_8_123_88_0 & ((~i_8_123_41_0 & ~i_8_123_118_0 & ~i_8_123_490_0 & ~i_8_123_728_0 & ~i_8_123_748_0 & ~i_8_123_828_0 & ~i_8_123_830_0 & ~i_8_123_956_0 & ~i_8_123_981_0 & ~i_8_123_1813_0 & ~i_8_123_2079_0) | (~i_8_123_107_0 & i_8_123_490_0 & ~i_8_123_814_0 & ~i_8_123_873_0 & ~i_8_123_1029_0 & ~i_8_123_1040_0 & ~i_8_123_1161_0 & ~i_8_123_1729_0 & ~i_8_123_1949_0 & ~i_8_123_2140_0 & ~i_8_123_2158_0))) | (~i_8_123_119_0 & ~i_8_123_2079_0 & ((~i_8_123_269_0 & ~i_8_123_1030_0 & ~i_8_123_1161_0 & ((~i_8_123_107_0 & ~i_8_123_118_0 & ~i_8_123_826_0 & ~i_8_123_830_0 & ~i_8_123_838_0 & ~i_8_123_1813_0) | (~i_8_123_489_0 & ~i_8_123_506_0 & ~i_8_123_728_0 & ~i_8_123_828_0 & ~i_8_123_956_0 & ~i_8_123_991_0 & ~i_8_123_1027_0 & ~i_8_123_1862_0))) | (~i_8_123_381_0 & ~i_8_123_826_0 & ~i_8_123_830_0 & ~i_8_123_873_0 & ~i_8_123_980_0 & ~i_8_123_981_0 & ~i_8_123_1029_0 & ~i_8_123_1031_0 & ~i_8_123_1058_0 & ~i_8_123_1949_0 & ~i_8_123_2052_0 & ~i_8_123_2158_0))) | (~i_8_123_489_0 & ~i_8_123_977_0 & ~i_8_123_981_0 & ~i_8_123_1027_0 & i_8_123_1470_0))) | (~i_8_123_981_0 & ((~i_8_123_308_0 & ((~i_8_123_167_0 & ~i_8_123_490_0 & ((~i_8_123_728_0 & ~i_8_123_826_0 & ~i_8_123_1027_0 & ~i_8_123_1028_0 & ~i_8_123_1029_0 & ~i_8_123_1030_0 & ~i_8_123_1355_0 & ~i_8_123_1437_0 & ~i_8_123_1449_0) | (~i_8_123_119_0 & i_8_123_1028_0 & ~i_8_123_1319_0 & ~i_8_123_1764_0))) | (~i_8_123_107_0 & ~i_8_123_608_0 & ~i_8_123_628_0 & ~i_8_123_748_0 & ~i_8_123_980_0 & ~i_8_123_991_0 & ~i_8_123_1029_0 & ~i_8_123_1030_0 & ~i_8_123_1161_0 & ~i_8_123_1449_0 & ~i_8_123_2059_0))) | (~i_8_123_107_0 & ~i_8_123_980_0 & ((~i_8_123_119_0 & ~i_8_123_628_0 & ~i_8_123_828_0 & ~i_8_123_1226_0 & i_8_123_1813_0) | (~i_8_123_258_0 & ~i_8_123_977_0 & ~i_8_123_1078_0 & ~i_8_123_1355_0 & ~i_8_123_1470_0 & i_8_123_1862_0 & ~i_8_123_2059_0))) | (~i_8_123_728_0 & ((~i_8_123_440_0 & i_8_123_686_0 & ~i_8_123_977_0 & ~i_8_123_1028_0) | (~i_8_123_119_0 & ~i_8_123_748_0 & i_8_123_1279_0 & ~i_8_123_1467_0 & ~i_8_123_1764_0 & ~i_8_123_2114_0))) | (i_8_123_72_0 & i_8_123_838_0 & ~i_8_123_956_0 & ~i_8_123_2052_0) | (~i_8_123_826_0 & ~i_8_123_830_0 & ~i_8_123_977_0 & i_8_123_1787_0 & ~i_8_123_1888_0 & ~i_8_123_2079_0) | (~i_8_123_630_0 & ~i_8_123_982_0 & i_8_123_2059_0 & ~i_8_123_2140_0))) | (~i_8_123_107_0 & ((~i_8_123_258_0 & ~i_8_123_814_0 & ~i_8_123_873_0 & ((~i_8_123_118_0 & ~i_8_123_381_0 & ~i_8_123_628_0 & ~i_8_123_728_0 & ~i_8_123_1162_0 & ~i_8_123_1729_0 & ~i_8_123_1862_0 & ~i_8_123_2079_0) | (~i_8_123_382_0 & ~i_8_123_991_0 & ~i_8_123_1027_0 & ~i_8_123_1746_0 & ~i_8_123_1764_0 & i_8_123_1780_0 & ~i_8_123_2126_0 & ~i_8_123_2241_0))) | (~i_8_123_440_0 & ((~i_8_123_628_0 & ~i_8_123_980_0 & ~i_8_123_1161_0 & i_8_123_1281_0 & ~i_8_123_1729_0) | (~i_8_123_977_0 & ~i_8_123_1027_0 & ~i_8_123_1030_0 & ~i_8_123_1281_0 & i_8_123_1355_0 & ~i_8_123_1765_0 & ~i_8_123_2126_0))) | (~i_8_123_308_0 & ~i_8_123_991_0 & i_8_123_1279_0 & ~i_8_123_1325_0 & ~i_8_123_1330_0 & ~i_8_123_1449_0))) | (~i_8_123_118_0 & ((~i_8_123_873_0 & i_8_123_1467_0) | (~i_8_123_728_0 & ~i_8_123_814_0 & ~i_8_123_991_0 & ~i_8_123_1162_0 & i_8_123_1281_0 & ~i_8_123_1355_0 & ~i_8_123_2079_0 & ~i_8_123_2241_0))) | (~i_8_123_1028_0 & ((~i_8_123_258_0 & ~i_8_123_1449_0 & ((~i_8_123_980_0 & ~i_8_123_982_0 & ~i_8_123_1729_0 & i_8_123_1949_0) | (~i_8_123_119_0 & ~i_8_123_748_0 & ~i_8_123_826_0 & ~i_8_123_828_0 & ~i_8_123_830_0 & ~i_8_123_977_0 & ~i_8_123_991_0 & ~i_8_123_1862_0 & ~i_8_123_2079_0 & ~i_8_123_2140_0 & ~i_8_123_2158_0))) | (~i_8_123_628_0 & i_8_123_710_0 & ~i_8_123_991_0 & ~i_8_123_1031_0 & ~i_8_123_1281_0) | (~i_8_123_828_0 & i_8_123_991_0 & i_8_123_1040_0 & ~i_8_123_1279_0 & ~i_8_123_1355_0 & ~i_8_123_2140_0))) | (~i_8_123_1027_0 & ((i_8_123_73_0 & ~i_8_123_991_0) | (~i_8_123_269_0 & i_8_123_382_0 & ~i_8_123_814_0 & ~i_8_123_977_0 & ~i_8_123_1161_0 & i_8_123_1281_0))) | (~i_8_123_2079_0 & ((~i_8_123_349_0 & ~i_8_123_350_0 & ~i_8_123_1029_0 & i_8_123_1470_0) | (~i_8_123_826_0 & ~i_8_123_1030_0 & ~i_8_123_1162_0 & i_8_123_1226_0 & ~i_8_123_1952_0))) | (i_8_123_608_0 & ~i_8_123_728_0 & ~i_8_123_982_0 & i_8_123_1355_0) | (~i_8_123_226_0 & i_8_123_490_0 & i_8_123_585_0 & ~i_8_123_709_0 & ~i_8_123_1262_0 & ~i_8_123_1746_0 & ~i_8_123_1889_0 & ~i_8_123_2140_0));
endmodule



// Benchmark "kernel_8_124" written by ABC on Sun Jul 19 10:05:11 2020

module kernel_8_124 ( 
    i_8_124_37_0, i_8_124_64_0, i_8_124_72_0, i_8_124_76_0, i_8_124_82_0,
    i_8_124_140_0, i_8_124_144_0, i_8_124_149_0, i_8_124_191_0,
    i_8_124_199_0, i_8_124_244_0, i_8_124_270_0, i_8_124_273_0,
    i_8_124_297_0, i_8_124_348_0, i_8_124_360_0, i_8_124_369_0,
    i_8_124_372_0, i_8_124_397_0, i_8_124_415_0, i_8_124_418_0,
    i_8_124_454_0, i_8_124_489_0, i_8_124_525_0, i_8_124_549_0,
    i_8_124_634_0, i_8_124_637_0, i_8_124_648_0, i_8_124_662_0,
    i_8_124_665_0, i_8_124_676_0, i_8_124_697_0, i_8_124_698_0,
    i_8_124_703_0, i_8_124_705_0, i_8_124_730_0, i_8_124_829_0,
    i_8_124_840_0, i_8_124_841_0, i_8_124_846_0, i_8_124_847_0,
    i_8_124_855_0, i_8_124_873_0, i_8_124_884_0, i_8_124_966_0,
    i_8_124_1027_0, i_8_124_1041_0, i_8_124_1042_0, i_8_124_1111_0,
    i_8_124_1112_0, i_8_124_1170_0, i_8_124_1224_0, i_8_124_1225_0,
    i_8_124_1235_0, i_8_124_1351_0, i_8_124_1387_0, i_8_124_1399_0,
    i_8_124_1458_0, i_8_124_1459_0, i_8_124_1479_0, i_8_124_1496_0,
    i_8_124_1522_0, i_8_124_1543_0, i_8_124_1550_0, i_8_124_1633_0,
    i_8_124_1638_0, i_8_124_1647_0, i_8_124_1648_0, i_8_124_1658_0,
    i_8_124_1682_0, i_8_124_1687_0, i_8_124_1705_0, i_8_124_1749_0,
    i_8_124_1765_0, i_8_124_1800_0, i_8_124_1810_0, i_8_124_1818_0,
    i_8_124_1819_0, i_8_124_1830_0, i_8_124_1845_0, i_8_124_1846_0,
    i_8_124_1864_0, i_8_124_1884_0, i_8_124_1885_0, i_8_124_1945_0,
    i_8_124_1996_0, i_8_124_2035_0, i_8_124_2038_0, i_8_124_2043_0,
    i_8_124_2044_0, i_8_124_2053_0, i_8_124_2125_0, i_8_124_2128_0,
    i_8_124_2141_0, i_8_124_2169_0, i_8_124_2173_0, i_8_124_2182_0,
    i_8_124_2253_0, i_8_124_2254_0, i_8_124_2255_0,
    o_8_124_0_0  );
  input  i_8_124_37_0, i_8_124_64_0, i_8_124_72_0, i_8_124_76_0,
    i_8_124_82_0, i_8_124_140_0, i_8_124_144_0, i_8_124_149_0,
    i_8_124_191_0, i_8_124_199_0, i_8_124_244_0, i_8_124_270_0,
    i_8_124_273_0, i_8_124_297_0, i_8_124_348_0, i_8_124_360_0,
    i_8_124_369_0, i_8_124_372_0, i_8_124_397_0, i_8_124_415_0,
    i_8_124_418_0, i_8_124_454_0, i_8_124_489_0, i_8_124_525_0,
    i_8_124_549_0, i_8_124_634_0, i_8_124_637_0, i_8_124_648_0,
    i_8_124_662_0, i_8_124_665_0, i_8_124_676_0, i_8_124_697_0,
    i_8_124_698_0, i_8_124_703_0, i_8_124_705_0, i_8_124_730_0,
    i_8_124_829_0, i_8_124_840_0, i_8_124_841_0, i_8_124_846_0,
    i_8_124_847_0, i_8_124_855_0, i_8_124_873_0, i_8_124_884_0,
    i_8_124_966_0, i_8_124_1027_0, i_8_124_1041_0, i_8_124_1042_0,
    i_8_124_1111_0, i_8_124_1112_0, i_8_124_1170_0, i_8_124_1224_0,
    i_8_124_1225_0, i_8_124_1235_0, i_8_124_1351_0, i_8_124_1387_0,
    i_8_124_1399_0, i_8_124_1458_0, i_8_124_1459_0, i_8_124_1479_0,
    i_8_124_1496_0, i_8_124_1522_0, i_8_124_1543_0, i_8_124_1550_0,
    i_8_124_1633_0, i_8_124_1638_0, i_8_124_1647_0, i_8_124_1648_0,
    i_8_124_1658_0, i_8_124_1682_0, i_8_124_1687_0, i_8_124_1705_0,
    i_8_124_1749_0, i_8_124_1765_0, i_8_124_1800_0, i_8_124_1810_0,
    i_8_124_1818_0, i_8_124_1819_0, i_8_124_1830_0, i_8_124_1845_0,
    i_8_124_1846_0, i_8_124_1864_0, i_8_124_1884_0, i_8_124_1885_0,
    i_8_124_1945_0, i_8_124_1996_0, i_8_124_2035_0, i_8_124_2038_0,
    i_8_124_2043_0, i_8_124_2044_0, i_8_124_2053_0, i_8_124_2125_0,
    i_8_124_2128_0, i_8_124_2141_0, i_8_124_2169_0, i_8_124_2173_0,
    i_8_124_2182_0, i_8_124_2253_0, i_8_124_2254_0, i_8_124_2255_0;
  output o_8_124_0_0;
  assign o_8_124_0_0 = 0;
endmodule



// Benchmark "kernel_8_125" written by ABC on Sun Jul 19 10:05:12 2020

module kernel_8_125 ( 
    i_8_125_13_0, i_8_125_52_0, i_8_125_103_0, i_8_125_112_0,
    i_8_125_130_0, i_8_125_142_0, i_8_125_165_0, i_8_125_199_0,
    i_8_125_221_0, i_8_125_237_0, i_8_125_254_0, i_8_125_334_0,
    i_8_125_361_0, i_8_125_391_0, i_8_125_424_0, i_8_125_453_0,
    i_8_125_455_0, i_8_125_459_0, i_8_125_475_0, i_8_125_492_0,
    i_8_125_507_0, i_8_125_523_0, i_8_125_544_0, i_8_125_598_0,
    i_8_125_607_0, i_8_125_624_0, i_8_125_654_0, i_8_125_659_0,
    i_8_125_660_0, i_8_125_662_0, i_8_125_685_0, i_8_125_695_0,
    i_8_125_696_0, i_8_125_699_0, i_8_125_704_0, i_8_125_755_0,
    i_8_125_760_0, i_8_125_765_0, i_8_125_786_0, i_8_125_797_0,
    i_8_125_806_0, i_8_125_840_0, i_8_125_841_0, i_8_125_895_0,
    i_8_125_926_0, i_8_125_931_0, i_8_125_940_0, i_8_125_966_0,
    i_8_125_1065_0, i_8_125_1108_0, i_8_125_1155_0, i_8_125_1197_0,
    i_8_125_1219_0, i_8_125_1237_0, i_8_125_1245_0, i_8_125_1258_0,
    i_8_125_1285_0, i_8_125_1290_0, i_8_125_1305_0, i_8_125_1321_0,
    i_8_125_1338_0, i_8_125_1398_0, i_8_125_1419_0, i_8_125_1426_0,
    i_8_125_1431_0, i_8_125_1433_0, i_8_125_1488_0, i_8_125_1527_0,
    i_8_125_1528_0, i_8_125_1650_0, i_8_125_1654_0, i_8_125_1682_0,
    i_8_125_1686_0, i_8_125_1689_0, i_8_125_1705_0, i_8_125_1801_0,
    i_8_125_1803_0, i_8_125_1804_0, i_8_125_1822_0, i_8_125_1825_0,
    i_8_125_1830_0, i_8_125_1831_0, i_8_125_1854_0, i_8_125_1855_0,
    i_8_125_1857_0, i_8_125_1858_0, i_8_125_1885_0, i_8_125_1980_0,
    i_8_125_1996_0, i_8_125_2092_0, i_8_125_2163_0, i_8_125_2203_0,
    i_8_125_2210_0, i_8_125_2224_0, i_8_125_2227_0, i_8_125_2260_0,
    i_8_125_2274_0, i_8_125_2281_0, i_8_125_2283_0, i_8_125_2290_0,
    o_8_125_0_0  );
  input  i_8_125_13_0, i_8_125_52_0, i_8_125_103_0, i_8_125_112_0,
    i_8_125_130_0, i_8_125_142_0, i_8_125_165_0, i_8_125_199_0,
    i_8_125_221_0, i_8_125_237_0, i_8_125_254_0, i_8_125_334_0,
    i_8_125_361_0, i_8_125_391_0, i_8_125_424_0, i_8_125_453_0,
    i_8_125_455_0, i_8_125_459_0, i_8_125_475_0, i_8_125_492_0,
    i_8_125_507_0, i_8_125_523_0, i_8_125_544_0, i_8_125_598_0,
    i_8_125_607_0, i_8_125_624_0, i_8_125_654_0, i_8_125_659_0,
    i_8_125_660_0, i_8_125_662_0, i_8_125_685_0, i_8_125_695_0,
    i_8_125_696_0, i_8_125_699_0, i_8_125_704_0, i_8_125_755_0,
    i_8_125_760_0, i_8_125_765_0, i_8_125_786_0, i_8_125_797_0,
    i_8_125_806_0, i_8_125_840_0, i_8_125_841_0, i_8_125_895_0,
    i_8_125_926_0, i_8_125_931_0, i_8_125_940_0, i_8_125_966_0,
    i_8_125_1065_0, i_8_125_1108_0, i_8_125_1155_0, i_8_125_1197_0,
    i_8_125_1219_0, i_8_125_1237_0, i_8_125_1245_0, i_8_125_1258_0,
    i_8_125_1285_0, i_8_125_1290_0, i_8_125_1305_0, i_8_125_1321_0,
    i_8_125_1338_0, i_8_125_1398_0, i_8_125_1419_0, i_8_125_1426_0,
    i_8_125_1431_0, i_8_125_1433_0, i_8_125_1488_0, i_8_125_1527_0,
    i_8_125_1528_0, i_8_125_1650_0, i_8_125_1654_0, i_8_125_1682_0,
    i_8_125_1686_0, i_8_125_1689_0, i_8_125_1705_0, i_8_125_1801_0,
    i_8_125_1803_0, i_8_125_1804_0, i_8_125_1822_0, i_8_125_1825_0,
    i_8_125_1830_0, i_8_125_1831_0, i_8_125_1854_0, i_8_125_1855_0,
    i_8_125_1857_0, i_8_125_1858_0, i_8_125_1885_0, i_8_125_1980_0,
    i_8_125_1996_0, i_8_125_2092_0, i_8_125_2163_0, i_8_125_2203_0,
    i_8_125_2210_0, i_8_125_2224_0, i_8_125_2227_0, i_8_125_2260_0,
    i_8_125_2274_0, i_8_125_2281_0, i_8_125_2283_0, i_8_125_2290_0;
  output o_8_125_0_0;
  assign o_8_125_0_0 = 0;
endmodule



// Benchmark "kernel_8_126" written by ABC on Sun Jul 19 10:05:12 2020

module kernel_8_126 ( 
    i_8_126_14_0, i_8_126_47_0, i_8_126_53_0, i_8_126_121_0, i_8_126_224_0,
    i_8_126_233_0, i_8_126_247_0, i_8_126_268_0, i_8_126_295_0,
    i_8_126_305_0, i_8_126_346_0, i_8_126_367_0, i_8_126_395_0,
    i_8_126_437_0, i_8_126_455_0, i_8_126_502_0, i_8_126_536_0,
    i_8_126_568_0, i_8_126_608_0, i_8_126_650_0, i_8_126_673_0,
    i_8_126_685_0, i_8_126_716_0, i_8_126_732_0, i_8_126_752_0,
    i_8_126_874_0, i_8_126_877_0, i_8_126_884_0, i_8_126_950_0,
    i_8_126_992_0, i_8_126_1012_0, i_8_126_1039_0, i_8_126_1057_0,
    i_8_126_1114_0, i_8_126_1143_0, i_8_126_1162_0, i_8_126_1222_0,
    i_8_126_1237_0, i_8_126_1262_0, i_8_126_1286_0, i_8_126_1298_0,
    i_8_126_1306_0, i_8_126_1308_0, i_8_126_1311_0, i_8_126_1330_0,
    i_8_126_1331_0, i_8_126_1423_0, i_8_126_1455_0, i_8_126_1456_0,
    i_8_126_1474_0, i_8_126_1483_0, i_8_126_1486_0, i_8_126_1487_0,
    i_8_126_1537_0, i_8_126_1543_0, i_8_126_1546_0, i_8_126_1590_0,
    i_8_126_1600_0, i_8_126_1612_0, i_8_126_1637_0, i_8_126_1651_0,
    i_8_126_1672_0, i_8_126_1723_0, i_8_126_1730_0, i_8_126_1738_0,
    i_8_126_1744_0, i_8_126_1754_0, i_8_126_1761_0, i_8_126_1769_0,
    i_8_126_1772_0, i_8_126_1780_0, i_8_126_1781_0, i_8_126_1798_0,
    i_8_126_1803_0, i_8_126_1822_0, i_8_126_1843_0, i_8_126_1858_0,
    i_8_126_1903_0, i_8_126_1927_0, i_8_126_1978_0, i_8_126_1979_0,
    i_8_126_2003_0, i_8_126_2021_0, i_8_126_2024_0, i_8_126_2045_0,
    i_8_126_2053_0, i_8_126_2069_0, i_8_126_2083_0, i_8_126_2094_0,
    i_8_126_2102_0, i_8_126_2126_0, i_8_126_2130_0, i_8_126_2131_0,
    i_8_126_2149_0, i_8_126_2150_0, i_8_126_2171_0, i_8_126_2172_0,
    i_8_126_2174_0, i_8_126_2273_0, i_8_126_2299_0,
    o_8_126_0_0  );
  input  i_8_126_14_0, i_8_126_47_0, i_8_126_53_0, i_8_126_121_0,
    i_8_126_224_0, i_8_126_233_0, i_8_126_247_0, i_8_126_268_0,
    i_8_126_295_0, i_8_126_305_0, i_8_126_346_0, i_8_126_367_0,
    i_8_126_395_0, i_8_126_437_0, i_8_126_455_0, i_8_126_502_0,
    i_8_126_536_0, i_8_126_568_0, i_8_126_608_0, i_8_126_650_0,
    i_8_126_673_0, i_8_126_685_0, i_8_126_716_0, i_8_126_732_0,
    i_8_126_752_0, i_8_126_874_0, i_8_126_877_0, i_8_126_884_0,
    i_8_126_950_0, i_8_126_992_0, i_8_126_1012_0, i_8_126_1039_0,
    i_8_126_1057_0, i_8_126_1114_0, i_8_126_1143_0, i_8_126_1162_0,
    i_8_126_1222_0, i_8_126_1237_0, i_8_126_1262_0, i_8_126_1286_0,
    i_8_126_1298_0, i_8_126_1306_0, i_8_126_1308_0, i_8_126_1311_0,
    i_8_126_1330_0, i_8_126_1331_0, i_8_126_1423_0, i_8_126_1455_0,
    i_8_126_1456_0, i_8_126_1474_0, i_8_126_1483_0, i_8_126_1486_0,
    i_8_126_1487_0, i_8_126_1537_0, i_8_126_1543_0, i_8_126_1546_0,
    i_8_126_1590_0, i_8_126_1600_0, i_8_126_1612_0, i_8_126_1637_0,
    i_8_126_1651_0, i_8_126_1672_0, i_8_126_1723_0, i_8_126_1730_0,
    i_8_126_1738_0, i_8_126_1744_0, i_8_126_1754_0, i_8_126_1761_0,
    i_8_126_1769_0, i_8_126_1772_0, i_8_126_1780_0, i_8_126_1781_0,
    i_8_126_1798_0, i_8_126_1803_0, i_8_126_1822_0, i_8_126_1843_0,
    i_8_126_1858_0, i_8_126_1903_0, i_8_126_1927_0, i_8_126_1978_0,
    i_8_126_1979_0, i_8_126_2003_0, i_8_126_2021_0, i_8_126_2024_0,
    i_8_126_2045_0, i_8_126_2053_0, i_8_126_2069_0, i_8_126_2083_0,
    i_8_126_2094_0, i_8_126_2102_0, i_8_126_2126_0, i_8_126_2130_0,
    i_8_126_2131_0, i_8_126_2149_0, i_8_126_2150_0, i_8_126_2171_0,
    i_8_126_2172_0, i_8_126_2174_0, i_8_126_2273_0, i_8_126_2299_0;
  output o_8_126_0_0;
  assign o_8_126_0_0 = 0;
endmodule



// Benchmark "kernel_8_127" written by ABC on Sun Jul 19 10:05:13 2020

module kernel_8_127 ( 
    i_8_127_94_0, i_8_127_111_0, i_8_127_124_0, i_8_127_190_0,
    i_8_127_191_0, i_8_127_223_0, i_8_127_231_0, i_8_127_248_0,
    i_8_127_301_0, i_8_127_328_0, i_8_127_346_0, i_8_127_365_0,
    i_8_127_368_0, i_8_127_376_0, i_8_127_420_0, i_8_127_439_0,
    i_8_127_445_0, i_8_127_455_0, i_8_127_471_0, i_8_127_492_0,
    i_8_127_499_0, i_8_127_522_0, i_8_127_523_0, i_8_127_530_0,
    i_8_127_591_0, i_8_127_597_0, i_8_127_634_0, i_8_127_637_0,
    i_8_127_645_0, i_8_127_660_0, i_8_127_673_0, i_8_127_681_0,
    i_8_127_696_0, i_8_127_697_0, i_8_127_770_0, i_8_127_841_0,
    i_8_127_871_0, i_8_127_877_0, i_8_127_879_0, i_8_127_880_0,
    i_8_127_888_0, i_8_127_924_0, i_8_127_958_0, i_8_127_961_0,
    i_8_127_969_0, i_8_127_976_0, i_8_127_993_0, i_8_127_1100_0,
    i_8_127_1105_0, i_8_127_1114_0, i_8_127_1137_0, i_8_127_1149_0,
    i_8_127_1189_0, i_8_127_1191_0, i_8_127_1192_0, i_8_127_1236_0,
    i_8_127_1239_0, i_8_127_1255_0, i_8_127_1266_0, i_8_127_1267_0,
    i_8_127_1281_0, i_8_127_1285_0, i_8_127_1356_0, i_8_127_1390_0,
    i_8_127_1444_0, i_8_127_1527_0, i_8_127_1535_0, i_8_127_1538_0,
    i_8_127_1545_0, i_8_127_1551_0, i_8_127_1596_0, i_8_127_1633_0,
    i_8_127_1634_0, i_8_127_1649_0, i_8_127_1741_0, i_8_127_1767_0,
    i_8_127_1770_0, i_8_127_1771_0, i_8_127_1779_0, i_8_127_1780_0,
    i_8_127_1814_0, i_8_127_1821_0, i_8_127_1840_0, i_8_127_1841_0,
    i_8_127_1859_0, i_8_127_1860_0, i_8_127_1861_0, i_8_127_1904_0,
    i_8_127_1991_0, i_8_127_2112_0, i_8_127_2137_0, i_8_127_2139_0,
    i_8_127_2141_0, i_8_127_2143_0, i_8_127_2146_0, i_8_127_2172_0,
    i_8_127_2215_0, i_8_127_2235_0, i_8_127_2247_0, i_8_127_2248_0,
    o_8_127_0_0  );
  input  i_8_127_94_0, i_8_127_111_0, i_8_127_124_0, i_8_127_190_0,
    i_8_127_191_0, i_8_127_223_0, i_8_127_231_0, i_8_127_248_0,
    i_8_127_301_0, i_8_127_328_0, i_8_127_346_0, i_8_127_365_0,
    i_8_127_368_0, i_8_127_376_0, i_8_127_420_0, i_8_127_439_0,
    i_8_127_445_0, i_8_127_455_0, i_8_127_471_0, i_8_127_492_0,
    i_8_127_499_0, i_8_127_522_0, i_8_127_523_0, i_8_127_530_0,
    i_8_127_591_0, i_8_127_597_0, i_8_127_634_0, i_8_127_637_0,
    i_8_127_645_0, i_8_127_660_0, i_8_127_673_0, i_8_127_681_0,
    i_8_127_696_0, i_8_127_697_0, i_8_127_770_0, i_8_127_841_0,
    i_8_127_871_0, i_8_127_877_0, i_8_127_879_0, i_8_127_880_0,
    i_8_127_888_0, i_8_127_924_0, i_8_127_958_0, i_8_127_961_0,
    i_8_127_969_0, i_8_127_976_0, i_8_127_993_0, i_8_127_1100_0,
    i_8_127_1105_0, i_8_127_1114_0, i_8_127_1137_0, i_8_127_1149_0,
    i_8_127_1189_0, i_8_127_1191_0, i_8_127_1192_0, i_8_127_1236_0,
    i_8_127_1239_0, i_8_127_1255_0, i_8_127_1266_0, i_8_127_1267_0,
    i_8_127_1281_0, i_8_127_1285_0, i_8_127_1356_0, i_8_127_1390_0,
    i_8_127_1444_0, i_8_127_1527_0, i_8_127_1535_0, i_8_127_1538_0,
    i_8_127_1545_0, i_8_127_1551_0, i_8_127_1596_0, i_8_127_1633_0,
    i_8_127_1634_0, i_8_127_1649_0, i_8_127_1741_0, i_8_127_1767_0,
    i_8_127_1770_0, i_8_127_1771_0, i_8_127_1779_0, i_8_127_1780_0,
    i_8_127_1814_0, i_8_127_1821_0, i_8_127_1840_0, i_8_127_1841_0,
    i_8_127_1859_0, i_8_127_1860_0, i_8_127_1861_0, i_8_127_1904_0,
    i_8_127_1991_0, i_8_127_2112_0, i_8_127_2137_0, i_8_127_2139_0,
    i_8_127_2141_0, i_8_127_2143_0, i_8_127_2146_0, i_8_127_2172_0,
    i_8_127_2215_0, i_8_127_2235_0, i_8_127_2247_0, i_8_127_2248_0;
  output o_8_127_0_0;
  assign o_8_127_0_0 = 0;
endmodule



// Benchmark "kernel_8_128" written by ABC on Sun Jul 19 10:05:14 2020

module kernel_8_128 ( 
    i_8_128_64_0, i_8_128_66_0, i_8_128_68_0, i_8_128_74_0, i_8_128_94_0,
    i_8_128_166_0, i_8_128_176_0, i_8_128_186_0, i_8_128_194_0,
    i_8_128_196_0, i_8_128_204_0, i_8_128_227_0, i_8_128_284_0,
    i_8_128_292_0, i_8_128_303_0, i_8_128_312_0, i_8_128_313_0,
    i_8_128_337_0, i_8_128_400_0, i_8_128_421_0, i_8_128_428_0,
    i_8_128_440_0, i_8_128_499_0, i_8_128_524_0, i_8_128_526_0,
    i_8_128_544_0, i_8_128_582_0, i_8_128_595_0, i_8_128_611_0,
    i_8_128_618_0, i_8_128_622_0, i_8_128_634_0, i_8_128_650_0,
    i_8_128_659_0, i_8_128_662_0, i_8_128_676_0, i_8_128_705_0,
    i_8_128_709_0, i_8_128_768_0, i_8_128_778_0, i_8_128_792_0,
    i_8_128_800_0, i_8_128_844_0, i_8_128_880_0, i_8_128_881_0,
    i_8_128_1023_0, i_8_128_1102_0, i_8_128_1104_0, i_8_128_1105_0,
    i_8_128_1123_0, i_8_128_1157_0, i_8_128_1162_0, i_8_128_1163_0,
    i_8_128_1219_0, i_8_128_1267_0, i_8_128_1317_0, i_8_128_1326_0,
    i_8_128_1383_0, i_8_128_1384_0, i_8_128_1427_0, i_8_128_1434_0,
    i_8_128_1437_0, i_8_128_1506_0, i_8_128_1551_0, i_8_128_1554_0,
    i_8_128_1555_0, i_8_128_1558_0, i_8_128_1559_0, i_8_128_1587_0,
    i_8_128_1609_0, i_8_128_1611_0, i_8_128_1681_0, i_8_128_1690_0,
    i_8_128_1743_0, i_8_128_1788_0, i_8_128_1822_0, i_8_128_1823_0,
    i_8_128_1880_0, i_8_128_1894_0, i_8_128_1913_0, i_8_128_1939_0,
    i_8_128_1940_0, i_8_128_1941_0, i_8_128_1942_0, i_8_128_1970_0,
    i_8_128_1974_0, i_8_128_1990_0, i_8_128_1999_0, i_8_128_2005_0,
    i_8_128_2092_0, i_8_128_2141_0, i_8_128_2156_0, i_8_128_2164_0,
    i_8_128_2166_0, i_8_128_2167_0, i_8_128_2183_0, i_8_128_2210_0,
    i_8_128_2216_0, i_8_128_2225_0, i_8_128_2279_0,
    o_8_128_0_0  );
  input  i_8_128_64_0, i_8_128_66_0, i_8_128_68_0, i_8_128_74_0,
    i_8_128_94_0, i_8_128_166_0, i_8_128_176_0, i_8_128_186_0,
    i_8_128_194_0, i_8_128_196_0, i_8_128_204_0, i_8_128_227_0,
    i_8_128_284_0, i_8_128_292_0, i_8_128_303_0, i_8_128_312_0,
    i_8_128_313_0, i_8_128_337_0, i_8_128_400_0, i_8_128_421_0,
    i_8_128_428_0, i_8_128_440_0, i_8_128_499_0, i_8_128_524_0,
    i_8_128_526_0, i_8_128_544_0, i_8_128_582_0, i_8_128_595_0,
    i_8_128_611_0, i_8_128_618_0, i_8_128_622_0, i_8_128_634_0,
    i_8_128_650_0, i_8_128_659_0, i_8_128_662_0, i_8_128_676_0,
    i_8_128_705_0, i_8_128_709_0, i_8_128_768_0, i_8_128_778_0,
    i_8_128_792_0, i_8_128_800_0, i_8_128_844_0, i_8_128_880_0,
    i_8_128_881_0, i_8_128_1023_0, i_8_128_1102_0, i_8_128_1104_0,
    i_8_128_1105_0, i_8_128_1123_0, i_8_128_1157_0, i_8_128_1162_0,
    i_8_128_1163_0, i_8_128_1219_0, i_8_128_1267_0, i_8_128_1317_0,
    i_8_128_1326_0, i_8_128_1383_0, i_8_128_1384_0, i_8_128_1427_0,
    i_8_128_1434_0, i_8_128_1437_0, i_8_128_1506_0, i_8_128_1551_0,
    i_8_128_1554_0, i_8_128_1555_0, i_8_128_1558_0, i_8_128_1559_0,
    i_8_128_1587_0, i_8_128_1609_0, i_8_128_1611_0, i_8_128_1681_0,
    i_8_128_1690_0, i_8_128_1743_0, i_8_128_1788_0, i_8_128_1822_0,
    i_8_128_1823_0, i_8_128_1880_0, i_8_128_1894_0, i_8_128_1913_0,
    i_8_128_1939_0, i_8_128_1940_0, i_8_128_1941_0, i_8_128_1942_0,
    i_8_128_1970_0, i_8_128_1974_0, i_8_128_1990_0, i_8_128_1999_0,
    i_8_128_2005_0, i_8_128_2092_0, i_8_128_2141_0, i_8_128_2156_0,
    i_8_128_2164_0, i_8_128_2166_0, i_8_128_2167_0, i_8_128_2183_0,
    i_8_128_2210_0, i_8_128_2216_0, i_8_128_2225_0, i_8_128_2279_0;
  output o_8_128_0_0;
  assign o_8_128_0_0 = 0;
endmodule



// Benchmark "kernel_8_129" written by ABC on Sun Jul 19 10:05:15 2020

module kernel_8_129 ( 
    i_8_129_22_0, i_8_129_48_0, i_8_129_64_0, i_8_129_72_0, i_8_129_73_0,
    i_8_129_74_0, i_8_129_76_0, i_8_129_90_0, i_8_129_94_0, i_8_129_136_0,
    i_8_129_171_0, i_8_129_194_0, i_8_129_197_0, i_8_129_297_0,
    i_8_129_325_0, i_8_129_505_0, i_8_129_550_0, i_8_129_585_0,
    i_8_129_586_0, i_8_129_588_0, i_8_129_595_0, i_8_129_621_0,
    i_8_129_622_0, i_8_129_624_0, i_8_129_630_0, i_8_129_631_0,
    i_8_129_632_0, i_8_129_652_0, i_8_129_653_0, i_8_129_684_0,
    i_8_129_702_0, i_8_129_703_0, i_8_129_707_0, i_8_129_820_0,
    i_8_129_829_0, i_8_129_969_0, i_8_129_990_0, i_8_129_991_0,
    i_8_129_1003_0, i_8_129_1012_0, i_8_129_1028_0, i_8_129_1029_0,
    i_8_129_1030_0, i_8_129_1031_0, i_8_129_1053_0, i_8_129_1054_0,
    i_8_129_1108_0, i_8_129_1198_0, i_8_129_1225_0, i_8_129_1263_0,
    i_8_129_1264_0, i_8_129_1265_0, i_8_129_1296_0, i_8_129_1297_0,
    i_8_129_1299_0, i_8_129_1351_0, i_8_129_1381_0, i_8_129_1395_0,
    i_8_129_1396_0, i_8_129_1398_0, i_8_129_1399_0, i_8_129_1400_0,
    i_8_129_1431_0, i_8_129_1449_0, i_8_129_1453_0, i_8_129_1454_0,
    i_8_129_1532_0, i_8_129_1621_0, i_8_129_1622_0, i_8_129_1701_0,
    i_8_129_1746_0, i_8_129_1767_0, i_8_129_1773_0, i_8_129_1776_0,
    i_8_129_1791_0, i_8_129_1802_0, i_8_129_1809_0, i_8_129_1818_0,
    i_8_129_1819_0, i_8_129_1821_0, i_8_129_1854_0, i_8_129_1855_0,
    i_8_129_1857_0, i_8_129_1899_0, i_8_129_1900_0, i_8_129_1903_0,
    i_8_129_1908_0, i_8_129_1911_0, i_8_129_1947_0, i_8_129_1948_0,
    i_8_129_1949_0, i_8_129_1963_0, i_8_129_1989_0, i_8_129_1992_0,
    i_8_129_1993_0, i_8_129_2134_0, i_8_129_2143_0, i_8_129_2246_0,
    i_8_129_2289_0, i_8_129_2294_0,
    o_8_129_0_0  );
  input  i_8_129_22_0, i_8_129_48_0, i_8_129_64_0, i_8_129_72_0,
    i_8_129_73_0, i_8_129_74_0, i_8_129_76_0, i_8_129_90_0, i_8_129_94_0,
    i_8_129_136_0, i_8_129_171_0, i_8_129_194_0, i_8_129_197_0,
    i_8_129_297_0, i_8_129_325_0, i_8_129_505_0, i_8_129_550_0,
    i_8_129_585_0, i_8_129_586_0, i_8_129_588_0, i_8_129_595_0,
    i_8_129_621_0, i_8_129_622_0, i_8_129_624_0, i_8_129_630_0,
    i_8_129_631_0, i_8_129_632_0, i_8_129_652_0, i_8_129_653_0,
    i_8_129_684_0, i_8_129_702_0, i_8_129_703_0, i_8_129_707_0,
    i_8_129_820_0, i_8_129_829_0, i_8_129_969_0, i_8_129_990_0,
    i_8_129_991_0, i_8_129_1003_0, i_8_129_1012_0, i_8_129_1028_0,
    i_8_129_1029_0, i_8_129_1030_0, i_8_129_1031_0, i_8_129_1053_0,
    i_8_129_1054_0, i_8_129_1108_0, i_8_129_1198_0, i_8_129_1225_0,
    i_8_129_1263_0, i_8_129_1264_0, i_8_129_1265_0, i_8_129_1296_0,
    i_8_129_1297_0, i_8_129_1299_0, i_8_129_1351_0, i_8_129_1381_0,
    i_8_129_1395_0, i_8_129_1396_0, i_8_129_1398_0, i_8_129_1399_0,
    i_8_129_1400_0, i_8_129_1431_0, i_8_129_1449_0, i_8_129_1453_0,
    i_8_129_1454_0, i_8_129_1532_0, i_8_129_1621_0, i_8_129_1622_0,
    i_8_129_1701_0, i_8_129_1746_0, i_8_129_1767_0, i_8_129_1773_0,
    i_8_129_1776_0, i_8_129_1791_0, i_8_129_1802_0, i_8_129_1809_0,
    i_8_129_1818_0, i_8_129_1819_0, i_8_129_1821_0, i_8_129_1854_0,
    i_8_129_1855_0, i_8_129_1857_0, i_8_129_1899_0, i_8_129_1900_0,
    i_8_129_1903_0, i_8_129_1908_0, i_8_129_1911_0, i_8_129_1947_0,
    i_8_129_1948_0, i_8_129_1949_0, i_8_129_1963_0, i_8_129_1989_0,
    i_8_129_1992_0, i_8_129_1993_0, i_8_129_2134_0, i_8_129_2143_0,
    i_8_129_2246_0, i_8_129_2289_0, i_8_129_2294_0;
  output o_8_129_0_0;
  assign o_8_129_0_0 = ~((~i_8_129_73_0 & ((~i_8_129_76_0 & ~i_8_129_586_0 & ~i_8_129_652_0 & ~i_8_129_702_0 & ~i_8_129_1992_0) | (~i_8_129_632_0 & ~i_8_129_1776_0 & ~i_8_129_1818_0 & ~i_8_129_1949_0 & ~i_8_129_2134_0))) | (~i_8_129_76_0 & ~i_8_129_1791_0 & ((~i_8_129_197_0 & ~i_8_129_505_0 & ~i_8_129_550_0 & ~i_8_129_1264_0 & ~i_8_129_1400_0 & i_8_129_1821_0 & ~i_8_129_1857_0 & i_8_129_1993_0) | (~i_8_129_171_0 & ~i_8_129_1263_0 & ~i_8_129_1399_0 & ~i_8_129_1819_0 & ~i_8_129_2134_0))) | (~i_8_129_586_0 & ((~i_8_129_632_0 & ((~i_8_129_550_0 & ((~i_8_129_1299_0 & ~i_8_129_1396_0 & ~i_8_129_1701_0 & ~i_8_129_1776_0 & ~i_8_129_1908_0 & ~i_8_129_1947_0) | (~i_8_129_585_0 & ~i_8_129_820_0 & ~i_8_129_1398_0 & ~i_8_129_1399_0 & ~i_8_129_1746_0 & ~i_8_129_1949_0))) | (~i_8_129_505_0 & ~i_8_129_702_0 & ~i_8_129_1030_0 & ~i_8_129_1198_0 & ~i_8_129_1225_0 & ~i_8_129_1296_0 & ~i_8_129_1400_0 & ~i_8_129_1949_0 & ~i_8_129_2134_0))) | (~i_8_129_64_0 & ~i_8_129_631_0 & ~i_8_129_1003_0 & ~i_8_129_1029_0 & ~i_8_129_1296_0 & i_8_129_1381_0 & ~i_8_129_1908_0))) | (~i_8_129_1911_0 & ((~i_8_129_64_0 & ((~i_8_129_990_0 & ~i_8_129_1264_0 & ~i_8_129_1395_0 & ~i_8_129_1396_0 & ~i_8_129_1398_0 & ~i_8_129_1400_0 & ~i_8_129_1773_0) | (~i_8_129_325_0 & ~i_8_129_595_0 & ~i_8_129_702_0 & ~i_8_129_1532_0 & ~i_8_129_1947_0 & ~i_8_129_1989_0 & ~i_8_129_1993_0 & ~i_8_129_2246_0))) | (~i_8_129_74_0 & ~i_8_129_1263_0 & ~i_8_129_1297_0 & ~i_8_129_1398_0 & ~i_8_129_1773_0 & ~i_8_129_1821_0) | (~i_8_129_297_0 & ~i_8_129_1030_0 & ~i_8_129_1265_0 & i_8_129_1299_0 & ~i_8_129_1381_0 & ~i_8_129_1908_0 & ~i_8_129_1947_0 & ~i_8_129_1949_0 & i_8_129_1992_0 & i_8_129_1993_0))) | (~i_8_129_585_0 & ((i_8_129_621_0 & ~i_8_129_1400_0) | (~i_8_129_1296_0 & ~i_8_129_1396_0 & ~i_8_129_1819_0 & ~i_8_129_1947_0 & ~i_8_129_1948_0 & ~i_8_129_1949_0))) | (~i_8_129_1400_0 & ((~i_8_129_653_0 & ((i_8_129_707_0 & i_8_129_1396_0 & ~i_8_129_1818_0 & ~i_8_129_1948_0) | (~i_8_129_171_0 & ~i_8_129_505_0 & ~i_8_129_652_0 & ~i_8_129_1296_0 & ~i_8_129_1299_0 & ~i_8_129_1453_0 & ~i_8_129_1903_0 & ~i_8_129_1992_0 & ~i_8_129_1993_0))) | (~i_8_129_702_0 & ~i_8_129_1297_0 & ~i_8_129_1431_0 & ~i_8_129_1821_0 & ~i_8_129_2143_0))) | (~i_8_129_1395_0 & ((~i_8_129_505_0 & ((i_8_129_595_0 & i_8_129_630_0 & ~i_8_129_703_0 & ~i_8_129_707_0 & ~i_8_129_1908_0) | (~i_8_129_22_0 & ~i_8_129_652_0 & ~i_8_129_969_0 & ~i_8_129_1225_0 & ~i_8_129_1396_0 & ~i_8_129_1453_0 & ~i_8_129_1949_0 & ~i_8_129_1989_0))) | (~i_8_129_72_0 & ~i_8_129_1265_0 & ~i_8_129_1297_0 & ~i_8_129_1299_0 & ~i_8_129_1381_0 & ~i_8_129_2246_0))) | (~i_8_129_72_0 & ((~i_8_129_595_0 & i_8_129_1108_0 & ~i_8_129_1396_0 & ~i_8_129_1948_0 & ~i_8_129_1993_0) | (~i_8_129_194_0 & ~i_8_129_703_0 & ~i_8_129_1297_0 & ~i_8_129_1399_0 & ~i_8_129_1773_0 & ~i_8_129_2143_0))) | (~i_8_129_630_0 & ~i_8_129_632_0 & ~i_8_129_652_0 & ~i_8_129_707_0 & ~i_8_129_1297_0 & ~i_8_129_1398_0 & ~i_8_129_1746_0) | (i_8_129_1449_0 & ~i_8_129_1767_0 & ~i_8_129_1776_0 & i_8_129_1993_0) | (~i_8_129_1265_0 & ~i_8_129_1396_0 & i_8_129_1819_0 & ~i_8_129_1821_0 & ~i_8_129_1857_0 & ~i_8_129_1908_0 & ~i_8_129_2246_0));
endmodule



// Benchmark "kernel_8_130" written by ABC on Sun Jul 19 10:05:16 2020

module kernel_8_130 ( 
    i_8_130_22_0, i_8_130_25_0, i_8_130_37_0, i_8_130_54_0, i_8_130_184_0,
    i_8_130_208_0, i_8_130_243_0, i_8_130_247_0, i_8_130_301_0,
    i_8_130_310_0, i_8_130_323_0, i_8_130_346_0, i_8_130_365_0,
    i_8_130_368_0, i_8_130_375_0, i_8_130_376_0, i_8_130_438_0,
    i_8_130_451_0, i_8_130_487_0, i_8_130_490_0, i_8_130_493_0,
    i_8_130_499_0, i_8_130_525_0, i_8_130_529_0, i_8_130_556_0,
    i_8_130_557_0, i_8_130_600_0, i_8_130_637_0, i_8_130_645_0,
    i_8_130_661_0, i_8_130_667_0, i_8_130_673_0, i_8_130_711_0,
    i_8_130_719_0, i_8_130_760_0, i_8_130_773_0, i_8_130_788_0,
    i_8_130_820_0, i_8_130_841_0, i_8_130_869_0, i_8_130_881_0,
    i_8_130_919_0, i_8_130_931_0, i_8_130_941_0, i_8_130_977_0,
    i_8_130_1015_0, i_8_130_1153_0, i_8_130_1171_0, i_8_130_1187_0,
    i_8_130_1204_0, i_8_130_1222_0, i_8_130_1228_0, i_8_130_1238_0,
    i_8_130_1240_0, i_8_130_1255_0, i_8_130_1261_0, i_8_130_1309_0,
    i_8_130_1315_0, i_8_130_1349_0, i_8_130_1388_0, i_8_130_1407_0,
    i_8_130_1408_0, i_8_130_1409_0, i_8_130_1419_0, i_8_130_1438_0,
    i_8_130_1472_0, i_8_130_1501_0, i_8_130_1528_0, i_8_130_1543_0,
    i_8_130_1544_0, i_8_130_1553_0, i_8_130_1600_0, i_8_130_1606_0,
    i_8_130_1705_0, i_8_130_1732_0, i_8_130_1736_0, i_8_130_1787_0,
    i_8_130_1819_0, i_8_130_1824_0, i_8_130_1849_0, i_8_130_1871_0,
    i_8_130_1876_0, i_8_130_1927_0, i_8_130_1992_0, i_8_130_1993_0,
    i_8_130_1996_0, i_8_130_1999_0, i_8_130_2041_0, i_8_130_2124_0,
    i_8_130_2154_0, i_8_130_2155_0, i_8_130_2215_0, i_8_130_2217_0,
    i_8_130_2218_0, i_8_130_2273_0, i_8_130_2278_0, i_8_130_2284_0,
    i_8_130_2286_0, i_8_130_2287_0, i_8_130_2292_0,
    o_8_130_0_0  );
  input  i_8_130_22_0, i_8_130_25_0, i_8_130_37_0, i_8_130_54_0,
    i_8_130_184_0, i_8_130_208_0, i_8_130_243_0, i_8_130_247_0,
    i_8_130_301_0, i_8_130_310_0, i_8_130_323_0, i_8_130_346_0,
    i_8_130_365_0, i_8_130_368_0, i_8_130_375_0, i_8_130_376_0,
    i_8_130_438_0, i_8_130_451_0, i_8_130_487_0, i_8_130_490_0,
    i_8_130_493_0, i_8_130_499_0, i_8_130_525_0, i_8_130_529_0,
    i_8_130_556_0, i_8_130_557_0, i_8_130_600_0, i_8_130_637_0,
    i_8_130_645_0, i_8_130_661_0, i_8_130_667_0, i_8_130_673_0,
    i_8_130_711_0, i_8_130_719_0, i_8_130_760_0, i_8_130_773_0,
    i_8_130_788_0, i_8_130_820_0, i_8_130_841_0, i_8_130_869_0,
    i_8_130_881_0, i_8_130_919_0, i_8_130_931_0, i_8_130_941_0,
    i_8_130_977_0, i_8_130_1015_0, i_8_130_1153_0, i_8_130_1171_0,
    i_8_130_1187_0, i_8_130_1204_0, i_8_130_1222_0, i_8_130_1228_0,
    i_8_130_1238_0, i_8_130_1240_0, i_8_130_1255_0, i_8_130_1261_0,
    i_8_130_1309_0, i_8_130_1315_0, i_8_130_1349_0, i_8_130_1388_0,
    i_8_130_1407_0, i_8_130_1408_0, i_8_130_1409_0, i_8_130_1419_0,
    i_8_130_1438_0, i_8_130_1472_0, i_8_130_1501_0, i_8_130_1528_0,
    i_8_130_1543_0, i_8_130_1544_0, i_8_130_1553_0, i_8_130_1600_0,
    i_8_130_1606_0, i_8_130_1705_0, i_8_130_1732_0, i_8_130_1736_0,
    i_8_130_1787_0, i_8_130_1819_0, i_8_130_1824_0, i_8_130_1849_0,
    i_8_130_1871_0, i_8_130_1876_0, i_8_130_1927_0, i_8_130_1992_0,
    i_8_130_1993_0, i_8_130_1996_0, i_8_130_1999_0, i_8_130_2041_0,
    i_8_130_2124_0, i_8_130_2154_0, i_8_130_2155_0, i_8_130_2215_0,
    i_8_130_2217_0, i_8_130_2218_0, i_8_130_2273_0, i_8_130_2278_0,
    i_8_130_2284_0, i_8_130_2286_0, i_8_130_2287_0, i_8_130_2292_0;
  output o_8_130_0_0;
  assign o_8_130_0_0 = 0;
endmodule



// Benchmark "kernel_8_131" written by ABC on Sun Jul 19 10:05:18 2020

module kernel_8_131 ( 
    i_8_131_73_0, i_8_131_87_0, i_8_131_101_0, i_8_131_181_0,
    i_8_131_182_0, i_8_131_190_0, i_8_131_191_0, i_8_131_232_0,
    i_8_131_243_0, i_8_131_244_0, i_8_131_303_0, i_8_131_304_0,
    i_8_131_339_0, i_8_131_383_0, i_8_131_391_0, i_8_131_396_0,
    i_8_131_397_0, i_8_131_454_0, i_8_131_473_0, i_8_131_490_0,
    i_8_131_594_0, i_8_131_595_0, i_8_131_596_0, i_8_131_628_0,
    i_8_131_629_0, i_8_131_632_0, i_8_131_665_0, i_8_131_716_0,
    i_8_131_719_0, i_8_131_748_0, i_8_131_752_0, i_8_131_757_0,
    i_8_131_850_0, i_8_131_855_0, i_8_131_856_0, i_8_131_858_0,
    i_8_131_969_0, i_8_131_994_0, i_8_131_1033_0, i_8_131_1036_0,
    i_8_131_1047_0, i_8_131_1057_0, i_8_131_1073_0, i_8_131_1078_0,
    i_8_131_1099_0, i_8_131_1100_0, i_8_131_1262_0, i_8_131_1283_0,
    i_8_131_1291_0, i_8_131_1306_0, i_8_131_1307_0, i_8_131_1330_0,
    i_8_131_1354_0, i_8_131_1372_0, i_8_131_1405_0, i_8_131_1439_0,
    i_8_131_1459_0, i_8_131_1470_0, i_8_131_1505_0, i_8_131_1507_0,
    i_8_131_1521_0, i_8_131_1529_0, i_8_131_1538_0, i_8_131_1607_0,
    i_8_131_1647_0, i_8_131_1649_0, i_8_131_1670_0, i_8_131_1675_0,
    i_8_131_1683_0, i_8_131_1736_0, i_8_131_1805_0, i_8_131_1807_0,
    i_8_131_1809_0, i_8_131_1811_0, i_8_131_1837_0, i_8_131_1862_0,
    i_8_131_1882_0, i_8_131_1883_0, i_8_131_1937_0, i_8_131_1964_0,
    i_8_131_1982_0, i_8_131_1993_0, i_8_131_1994_0, i_8_131_2007_0,
    i_8_131_2057_0, i_8_131_2072_0, i_8_131_2106_0, i_8_131_2139_0,
    i_8_131_2140_0, i_8_131_2147_0, i_8_131_2153_0, i_8_131_2155_0,
    i_8_131_2156_0, i_8_131_2161_0, i_8_131_2180_0, i_8_131_2215_0,
    i_8_131_2241_0, i_8_131_2246_0, i_8_131_2267_0, i_8_131_2275_0,
    o_8_131_0_0  );
  input  i_8_131_73_0, i_8_131_87_0, i_8_131_101_0, i_8_131_181_0,
    i_8_131_182_0, i_8_131_190_0, i_8_131_191_0, i_8_131_232_0,
    i_8_131_243_0, i_8_131_244_0, i_8_131_303_0, i_8_131_304_0,
    i_8_131_339_0, i_8_131_383_0, i_8_131_391_0, i_8_131_396_0,
    i_8_131_397_0, i_8_131_454_0, i_8_131_473_0, i_8_131_490_0,
    i_8_131_594_0, i_8_131_595_0, i_8_131_596_0, i_8_131_628_0,
    i_8_131_629_0, i_8_131_632_0, i_8_131_665_0, i_8_131_716_0,
    i_8_131_719_0, i_8_131_748_0, i_8_131_752_0, i_8_131_757_0,
    i_8_131_850_0, i_8_131_855_0, i_8_131_856_0, i_8_131_858_0,
    i_8_131_969_0, i_8_131_994_0, i_8_131_1033_0, i_8_131_1036_0,
    i_8_131_1047_0, i_8_131_1057_0, i_8_131_1073_0, i_8_131_1078_0,
    i_8_131_1099_0, i_8_131_1100_0, i_8_131_1262_0, i_8_131_1283_0,
    i_8_131_1291_0, i_8_131_1306_0, i_8_131_1307_0, i_8_131_1330_0,
    i_8_131_1354_0, i_8_131_1372_0, i_8_131_1405_0, i_8_131_1439_0,
    i_8_131_1459_0, i_8_131_1470_0, i_8_131_1505_0, i_8_131_1507_0,
    i_8_131_1521_0, i_8_131_1529_0, i_8_131_1538_0, i_8_131_1607_0,
    i_8_131_1647_0, i_8_131_1649_0, i_8_131_1670_0, i_8_131_1675_0,
    i_8_131_1683_0, i_8_131_1736_0, i_8_131_1805_0, i_8_131_1807_0,
    i_8_131_1809_0, i_8_131_1811_0, i_8_131_1837_0, i_8_131_1862_0,
    i_8_131_1882_0, i_8_131_1883_0, i_8_131_1937_0, i_8_131_1964_0,
    i_8_131_1982_0, i_8_131_1993_0, i_8_131_1994_0, i_8_131_2007_0,
    i_8_131_2057_0, i_8_131_2072_0, i_8_131_2106_0, i_8_131_2139_0,
    i_8_131_2140_0, i_8_131_2147_0, i_8_131_2153_0, i_8_131_2155_0,
    i_8_131_2156_0, i_8_131_2161_0, i_8_131_2180_0, i_8_131_2215_0,
    i_8_131_2241_0, i_8_131_2246_0, i_8_131_2267_0, i_8_131_2275_0;
  output o_8_131_0_0;
  assign o_8_131_0_0 = ~((i_8_131_391_0 & ((~i_8_131_190_0 & ~i_8_131_303_0 & ~i_8_131_304_0 & ~i_8_131_748_0 & ~i_8_131_1078_0 & ~i_8_131_1538_0 & ~i_8_131_1649_0 & i_8_131_1805_0) | (i_8_131_594_0 & i_8_131_628_0 & i_8_131_1047_0 & ~i_8_131_2139_0))) | (~i_8_131_1100_0 & ((i_8_131_454_0 & ((~i_8_131_190_0 & ~i_8_131_391_0 & ~i_8_131_397_0 & ~i_8_131_629_0 & ~i_8_131_752_0 & ~i_8_131_1459_0 & ~i_8_131_1675_0 & ~i_8_131_1805_0 & ~i_8_131_1883_0 & ~i_8_131_2139_0) | (~i_8_131_719_0 & ~i_8_131_1505_0 & ~i_8_131_1507_0 & ~i_8_131_1647_0 & ~i_8_131_1837_0 & ~i_8_131_1862_0 & ~i_8_131_2215_0 & ~i_8_131_2267_0))) | (~i_8_131_397_0 & ((~i_8_131_87_0 & ~i_8_131_304_0 & ~i_8_131_594_0 & i_8_131_1306_0 & ~i_8_131_1372_0 & ~i_8_131_1521_0 & ~i_8_131_1683_0 & ~i_8_131_1736_0 & ~i_8_131_1837_0 & ~i_8_131_1937_0) | (~i_8_131_101_0 & ~i_8_131_303_0 & ~i_8_131_391_0 & ~i_8_131_396_0 & ~i_8_131_454_0 & ~i_8_131_629_0 & ~i_8_131_719_0 & i_8_131_850_0 & ~i_8_131_1047_0 & ~i_8_131_1529_0 & ~i_8_131_2139_0 & ~i_8_131_2161_0))) | (~i_8_131_182_0 & ((~i_8_131_1683_0 & ((~i_8_131_87_0 & ~i_8_131_628_0 & ~i_8_131_752_0 & ~i_8_131_1033_0 & ((~i_8_131_396_0 & ~i_8_131_454_0 & ~i_8_131_1262_0 & ~i_8_131_1354_0 & ~i_8_131_1521_0 & ~i_8_131_1862_0 & ~i_8_131_1882_0 & ~i_8_131_2140_0 & ~i_8_131_2147_0 & ~i_8_131_2156_0) | (~i_8_131_665_0 & ~i_8_131_969_0 & ~i_8_131_1675_0 & ~i_8_131_1883_0 & ~i_8_131_1993_0 & ~i_8_131_2106_0 & ~i_8_131_2153_0 & ~i_8_131_2241_0 & ~i_8_131_2275_0))) | (i_8_131_473_0 & ~i_8_131_629_0 & ~i_8_131_719_0 & ~i_8_131_850_0 & ~i_8_131_1459_0 & ~i_8_131_1505_0 & ~i_8_131_1507_0 & ~i_8_131_1529_0) | (~i_8_131_181_0 & ~i_8_131_339_0 & ~i_8_131_391_0 & ~i_8_131_2147_0 & ~i_8_131_2153_0 & i_8_131_2215_0 & ~i_8_131_2267_0))) | (~i_8_131_1529_0 & ((~i_8_131_339_0 & ~i_8_131_396_0 & ~i_8_131_490_0 & ~i_8_131_748_0 & ~i_8_131_1283_0 & ~i_8_131_1330_0 & ~i_8_131_1521_0 & ~i_8_131_1538_0 & ~i_8_131_1647_0 & ~i_8_131_1805_0 & ~i_8_131_2007_0 & ~i_8_131_2153_0 & ~i_8_131_2156_0) | (~i_8_131_190_0 & ~i_8_131_191_0 & ~i_8_131_628_0 & ~i_8_131_855_0 & ~i_8_131_1033_0 & ~i_8_131_1099_0 & ~i_8_131_1372_0 & ~i_8_131_1405_0 & ~i_8_131_1439_0 & ~i_8_131_1507_0 & ~i_8_131_1937_0 & ~i_8_131_2241_0))))) | (~i_8_131_1033_0 & ((~i_8_131_190_0 & ~i_8_131_2106_0 & ~i_8_131_2153_0 & ((~i_8_131_473_0 & ~i_8_131_748_0 & ~i_8_131_855_0 & ~i_8_131_1036_0 & ~i_8_131_1439_0 & ~i_8_131_1521_0 & ~i_8_131_1647_0 & ~i_8_131_1670_0 & ~i_8_131_1862_0 & ~i_8_131_2147_0 & ~i_8_131_2180_0) | (~i_8_131_391_0 & ~i_8_131_396_0 & ~i_8_131_629_0 & ~i_8_131_719_0 & ~i_8_131_850_0 & ~i_8_131_969_0 & ~i_8_131_1283_0 & ~i_8_131_1372_0 & ~i_8_131_1470_0 & ~i_8_131_1505_0 & ~i_8_131_1993_0 & ~i_8_131_1994_0 & ~i_8_131_2241_0 & ~i_8_131_2275_0 & ~i_8_131_2007_0 & ~i_8_131_2156_0))) | (~i_8_131_339_0 & ~i_8_131_396_0 & ~i_8_131_752_0 & ~i_8_131_1283_0 & ~i_8_131_1330_0 & ~i_8_131_1078_0 & ~i_8_131_1262_0 & ~i_8_131_1521_0 & ~i_8_131_1647_0 & ~i_8_131_1649_0 & ~i_8_131_1675_0 & ~i_8_131_1805_0 & ~i_8_131_2180_0 & ~i_8_131_2215_0))) | (~i_8_131_396_0 & ~i_8_131_1647_0 & ((~i_8_131_1807_0 & i_8_131_1809_0 & ~i_8_131_1837_0 & ~i_8_131_1882_0 & ~i_8_131_1982_0) | (~i_8_131_628_0 & ~i_8_131_665_0 & i_8_131_1057_0 & ~i_8_131_1521_0 & ~i_8_131_1670_0 & ~i_8_131_1683_0 & ~i_8_131_2072_0 & ~i_8_131_2140_0))) | (i_8_131_595_0 & ~i_8_131_628_0 & ~i_8_131_1099_0 & ~i_8_131_1683_0 & ~i_8_131_1982_0 & ~i_8_131_2007_0 & ~i_8_131_2072_0 & ~i_8_131_2153_0))) | (~i_8_131_629_0 & ((i_8_131_1057_0 & ~i_8_131_1099_0 & ~i_8_131_1683_0 & i_8_131_2007_0 & ~i_8_131_2156_0) | (~i_8_131_182_0 & ~i_8_131_190_0 & ~i_8_131_303_0 & ~i_8_131_304_0 & ~i_8_131_396_0 & ~i_8_131_490_0 & ~i_8_131_719_0 & ~i_8_131_1521_0 & ~i_8_131_1807_0 & ~i_8_131_1837_0 & ~i_8_131_1883_0 & ~i_8_131_1993_0 & ~i_8_131_2057_0 & ~i_8_131_2246_0))) | (~i_8_131_665_0 & ((~i_8_131_190_0 & ~i_8_131_490_0 & ~i_8_131_752_0 & ~i_8_131_1283_0 & i_8_131_1862_0 & ~i_8_131_1883_0 & ~i_8_131_2139_0 & ~i_8_131_2153_0 & ~i_8_131_2267_0) | (~i_8_131_182_0 & ~i_8_131_191_0 & ~i_8_131_748_0 & ~i_8_131_1807_0 & ~i_8_131_1937_0 & i_8_131_2057_0 & ~i_8_131_2275_0))) | (~i_8_131_191_0 & ((~i_8_131_87_0 & ~i_8_131_182_0 & i_8_131_596_0 & ~i_8_131_1372_0 & ~i_8_131_1405_0 & ~i_8_131_1459_0) | (~i_8_131_396_0 & ~i_8_131_490_0 & ~i_8_131_628_0 & ~i_8_131_1439_0 & ~i_8_131_1647_0 & ~i_8_131_1670_0 & ~i_8_131_1837_0 & ~i_8_131_1937_0 & ~i_8_131_1993_0 & ~i_8_131_2180_0 & ~i_8_131_2267_0))) | (~i_8_131_2106_0 & ((~i_8_131_2153_0 & ((~i_8_131_87_0 & ((~i_8_131_181_0 & ~i_8_131_339_0 & ~i_8_131_391_0 & ~i_8_131_396_0 & ~i_8_131_1033_0 & ~i_8_131_1036_0 & i_8_131_1405_0 & ~i_8_131_1507_0 & i_8_131_1882_0 & ~i_8_131_2072_0 & ~i_8_131_2161_0) | (~i_8_131_397_0 & ~i_8_131_490_0 & ~i_8_131_632_0 & ~i_8_131_1078_0 & ~i_8_131_1354_0 & ~i_8_131_1607_0 & ~i_8_131_1647_0 & ~i_8_131_1670_0 & ~i_8_131_1805_0 & ~i_8_131_2140_0 & ~i_8_131_2147_0 & ~i_8_131_2241_0 & ~i_8_131_2275_0 & ~i_8_131_2156_0 & ~i_8_131_2180_0))) | (~i_8_131_181_0 & ~i_8_131_190_0 & ~i_8_131_1033_0 & ~i_8_131_1521_0 & ~i_8_131_1529_0 & ~i_8_131_1649_0 & ~i_8_131_1670_0 & ~i_8_131_1736_0 & ~i_8_131_1837_0 & i_8_131_1993_0 & ~i_8_131_2139_0 & ~i_8_131_2155_0 & ~i_8_131_2215_0 & ~i_8_131_2241_0))) | (~i_8_131_396_0 & ~i_8_131_1807_0 & ((i_8_131_594_0 & i_8_131_628_0 & ~i_8_131_969_0 & ~i_8_131_1047_0 & ~i_8_131_2215_0) | (i_8_131_190_0 & ~i_8_131_490_0 & ~i_8_131_748_0 & ~i_8_131_1099_0 & ~i_8_131_1507_0 & ~i_8_131_1521_0 & ~i_8_131_1649_0 & ~i_8_131_1683_0 & ~i_8_131_2156_0 & ~i_8_131_2246_0))) | (~i_8_131_1937_0 & ((i_8_131_101_0 & ~i_8_131_181_0 & ~i_8_131_1036_0 & ~i_8_131_2072_0 & ~i_8_131_2139_0 & ~i_8_131_2140_0) | (~i_8_131_190_0 & ~i_8_131_232_0 & i_8_131_1047_0 & ~i_8_131_1330_0 & ~i_8_131_1521_0 & ~i_8_131_1647_0 & ~i_8_131_1649_0 & ~i_8_131_1736_0 & ~i_8_131_2246_0))) | (i_8_131_490_0 & ~i_8_131_1047_0 & ~i_8_131_1099_0 & ~i_8_131_1306_0 & i_8_131_2007_0 & i_8_131_2241_0))) | (~i_8_131_397_0 & ((~i_8_131_190_0 & ((~i_8_131_1647_0 & ~i_8_131_1649_0 & i_8_131_595_0 & ~i_8_131_1529_0 & ~i_8_131_1736_0 & ~i_8_131_1982_0 & ~i_8_131_2057_0 & ~i_8_131_2072_0) | (~i_8_131_182_0 & i_8_131_383_0 & ~i_8_131_391_0 & ~i_8_131_719_0 & ~i_8_131_1675_0 & i_8_131_2147_0 & ~i_8_131_2180_0 & ~i_8_131_2241_0))) | (~i_8_131_391_0 & ~i_8_131_1078_0 & i_8_131_1283_0 & ~i_8_131_1505_0 & ~i_8_131_1683_0 & ~i_8_131_1883_0 & i_8_131_1964_0 & ~i_8_131_2007_0 & ~i_8_131_2180_0))) | (i_8_131_383_0 & ((~i_8_131_1073_0 & ~i_8_131_1099_0 & i_8_131_1283_0 & ~i_8_131_1937_0 & i_8_131_1964_0) | (~i_8_131_303_0 & ~i_8_131_391_0 & ~i_8_131_716_0 & ~i_8_131_1330_0 & ~i_8_131_1538_0 & ~i_8_131_1683_0 & ~i_8_131_1982_0 & ~i_8_131_1994_0 & ~i_8_131_2147_0 & ~i_8_131_2153_0))) | (~i_8_131_1647_0 & ((~i_8_131_1538_0 & ((~i_8_131_391_0 & ((~i_8_131_182_0 & ~i_8_131_1805_0 & ~i_8_131_1937_0 & ~i_8_131_2139_0 & ~i_8_131_2241_0 & ((~i_8_131_303_0 & ~i_8_131_1078_0 & ~i_8_131_1262_0 & ~i_8_131_1330_0 & ~i_8_131_1354_0 & ~i_8_131_1372_0 & ~i_8_131_1529_0 & ~i_8_131_1649_0) | (~i_8_131_1033_0 & ~i_8_131_1099_0 & ~i_8_131_1439_0 & ~i_8_131_1505_0 & ~i_8_131_1837_0 & ~i_8_131_1993_0 & ~i_8_131_2267_0))) | (~i_8_131_969_0 & ~i_8_131_1439_0 & i_8_131_1805_0 & ~i_8_131_1811_0 & ~i_8_131_1982_0 & ~i_8_131_2246_0 & ~i_8_131_2267_0))) | (~i_8_131_87_0 & ~i_8_131_748_0 & ~i_8_131_858_0 & ~i_8_131_1033_0 & ~i_8_131_1099_0 & ~i_8_131_1529_0 & ~i_8_131_1670_0 & ~i_8_131_1683_0 & ~i_8_131_1937_0 & i_8_131_2155_0))) | (~i_8_131_303_0 & ~i_8_131_719_0 & ~i_8_131_1405_0 & ~i_8_131_1470_0 & ~i_8_131_1529_0 & ~i_8_131_1649_0 & i_8_131_1807_0 & ~i_8_131_2140_0 & ~i_8_131_2147_0 & ~i_8_131_2153_0) | (~i_8_131_396_0 & i_8_131_1047_0 & ~i_8_131_1078_0 & ~i_8_131_1675_0 & i_8_131_2106_0 & ~i_8_131_2161_0))) | (~i_8_131_1099_0 & ((~i_8_131_87_0 & ~i_8_131_628_0 & ~i_8_131_1670_0 & ((~i_8_131_339_0 & ~i_8_131_396_0 & ~i_8_131_716_0 & ~i_8_131_748_0 & ~i_8_131_1036_0 & i_8_131_1057_0 & ~i_8_131_1078_0 & ~i_8_131_2057_0 & ~i_8_131_2072_0) | (~i_8_131_391_0 & ~i_8_131_719_0 & i_8_131_1033_0 & ~i_8_131_1507_0 & ~i_8_131_1529_0 & ~i_8_131_2246_0))) | (i_8_131_244_0 & i_8_131_716_0 & ~i_8_131_1507_0) | (i_8_131_1036_0 & i_8_131_1047_0 & i_8_131_1675_0 & ~i_8_131_1683_0 & i_8_131_2241_0))) | (~i_8_131_1262_0 & ((~i_8_131_304_0 & ((~i_8_131_339_0 & ~i_8_131_396_0 & ~i_8_131_1036_0 & ~i_8_131_1507_0 & ~i_8_131_1649_0 & i_8_131_1809_0) | (i_8_131_969_0 & ~i_8_131_1047_0 & i_8_131_1078_0 & ~i_8_131_1405_0 & ~i_8_131_1521_0 & ~i_8_131_1529_0 & ~i_8_131_1670_0 & ~i_8_131_1883_0))) | (~i_8_131_339_0 & ~i_8_131_752_0 & ~i_8_131_1047_0 & ~i_8_131_1073_0 & ~i_8_131_1306_0 & ~i_8_131_1683_0 & ~i_8_131_2072_0 & ~i_8_131_2147_0 & i_8_131_2156_0))) | (~i_8_131_304_0 & ~i_8_131_1837_0 & ~i_8_131_1882_0 & ((~i_8_131_1078_0 & ~i_8_131_1354_0 & ~i_8_131_181_0 & ~i_8_131_391_0 & i_8_131_1372_0 & ~i_8_131_1675_0 & ~i_8_131_1736_0 & ~i_8_131_2153_0) | (~i_8_131_1607_0 & ~i_8_131_1670_0 & ~i_8_131_1883_0 & ~i_8_131_2215_0 & ~i_8_131_2241_0 & ~i_8_131_2072_0 & i_8_131_2156_0))) | (~i_8_131_1683_0 & ((i_8_131_73_0 & ~i_8_131_182_0 & ~i_8_131_1033_0 & ~i_8_131_1807_0 & i_8_131_1809_0 & ~i_8_131_1505_0 & ~i_8_131_1538_0) | (~i_8_131_73_0 & ~i_8_131_383_0 & i_8_131_1306_0 & ~i_8_131_1439_0 & ~i_8_131_1521_0 & ~i_8_131_1649_0 & ~i_8_131_2007_0 & ~i_8_131_2153_0))) | (i_8_131_1057_0 & ~i_8_131_1507_0 & i_8_131_1807_0 & ~i_8_131_1993_0 & i_8_131_2139_0 & ~i_8_131_2275_0));
endmodule



// Benchmark "kernel_8_132" written by ABC on Sun Jul 19 10:05:19 2020

module kernel_8_132 ( 
    i_8_132_9_0, i_8_132_12_0, i_8_132_18_0, i_8_132_42_0, i_8_132_69_0,
    i_8_132_78_0, i_8_132_103_0, i_8_132_138_0, i_8_132_151_0,
    i_8_132_166_0, i_8_132_174_0, i_8_132_196_0, i_8_132_229_0,
    i_8_132_283_0, i_8_132_300_0, i_8_132_301_0, i_8_132_318_0,
    i_8_132_337_0, i_8_132_338_0, i_8_132_365_0, i_8_132_367_0,
    i_8_132_397_0, i_8_132_496_0, i_8_132_529_0, i_8_132_537_0,
    i_8_132_544_0, i_8_132_573_0, i_8_132_672_0, i_8_132_703_0,
    i_8_132_704_0, i_8_132_707_0, i_8_132_733_0, i_8_132_773_0,
    i_8_132_806_0, i_8_132_864_0, i_8_132_865_0, i_8_132_866_0,
    i_8_132_937_0, i_8_132_979_0, i_8_132_993_0, i_8_132_1003_0,
    i_8_132_1057_0, i_8_132_1074_0, i_8_132_1104_0, i_8_132_1105_0,
    i_8_132_1151_0, i_8_132_1224_0, i_8_132_1225_0, i_8_132_1228_0,
    i_8_132_1239_0, i_8_132_1258_0, i_8_132_1260_0, i_8_132_1261_0,
    i_8_132_1262_0, i_8_132_1291_0, i_8_132_1292_0, i_8_132_1323_0,
    i_8_132_1333_0, i_8_132_1335_0, i_8_132_1356_0, i_8_132_1384_0,
    i_8_132_1410_0, i_8_132_1412_0, i_8_132_1429_0, i_8_132_1449_0,
    i_8_132_1464_0, i_8_132_1468_0, i_8_132_1471_0, i_8_132_1491_0,
    i_8_132_1515_0, i_8_132_1527_0, i_8_132_1531_0, i_8_132_1562_0,
    i_8_132_1645_0, i_8_132_1653_0, i_8_132_1654_0, i_8_132_1686_0,
    i_8_132_1723_0, i_8_132_1746_0, i_8_132_1751_0, i_8_132_1807_0,
    i_8_132_1823_0, i_8_132_1858_0, i_8_132_1894_0, i_8_132_1907_0,
    i_8_132_1912_0, i_8_132_1956_0, i_8_132_1962_0, i_8_132_1963_0,
    i_8_132_1984_0, i_8_132_1995_0, i_8_132_2106_0, i_8_132_2145_0,
    i_8_132_2151_0, i_8_132_2152_0, i_8_132_2174_0, i_8_132_2200_0,
    i_8_132_2202_0, i_8_132_2245_0, i_8_132_2259_0,
    o_8_132_0_0  );
  input  i_8_132_9_0, i_8_132_12_0, i_8_132_18_0, i_8_132_42_0,
    i_8_132_69_0, i_8_132_78_0, i_8_132_103_0, i_8_132_138_0,
    i_8_132_151_0, i_8_132_166_0, i_8_132_174_0, i_8_132_196_0,
    i_8_132_229_0, i_8_132_283_0, i_8_132_300_0, i_8_132_301_0,
    i_8_132_318_0, i_8_132_337_0, i_8_132_338_0, i_8_132_365_0,
    i_8_132_367_0, i_8_132_397_0, i_8_132_496_0, i_8_132_529_0,
    i_8_132_537_0, i_8_132_544_0, i_8_132_573_0, i_8_132_672_0,
    i_8_132_703_0, i_8_132_704_0, i_8_132_707_0, i_8_132_733_0,
    i_8_132_773_0, i_8_132_806_0, i_8_132_864_0, i_8_132_865_0,
    i_8_132_866_0, i_8_132_937_0, i_8_132_979_0, i_8_132_993_0,
    i_8_132_1003_0, i_8_132_1057_0, i_8_132_1074_0, i_8_132_1104_0,
    i_8_132_1105_0, i_8_132_1151_0, i_8_132_1224_0, i_8_132_1225_0,
    i_8_132_1228_0, i_8_132_1239_0, i_8_132_1258_0, i_8_132_1260_0,
    i_8_132_1261_0, i_8_132_1262_0, i_8_132_1291_0, i_8_132_1292_0,
    i_8_132_1323_0, i_8_132_1333_0, i_8_132_1335_0, i_8_132_1356_0,
    i_8_132_1384_0, i_8_132_1410_0, i_8_132_1412_0, i_8_132_1429_0,
    i_8_132_1449_0, i_8_132_1464_0, i_8_132_1468_0, i_8_132_1471_0,
    i_8_132_1491_0, i_8_132_1515_0, i_8_132_1527_0, i_8_132_1531_0,
    i_8_132_1562_0, i_8_132_1645_0, i_8_132_1653_0, i_8_132_1654_0,
    i_8_132_1686_0, i_8_132_1723_0, i_8_132_1746_0, i_8_132_1751_0,
    i_8_132_1807_0, i_8_132_1823_0, i_8_132_1858_0, i_8_132_1894_0,
    i_8_132_1907_0, i_8_132_1912_0, i_8_132_1956_0, i_8_132_1962_0,
    i_8_132_1963_0, i_8_132_1984_0, i_8_132_1995_0, i_8_132_2106_0,
    i_8_132_2145_0, i_8_132_2151_0, i_8_132_2152_0, i_8_132_2174_0,
    i_8_132_2200_0, i_8_132_2202_0, i_8_132_2245_0, i_8_132_2259_0;
  output o_8_132_0_0;
  assign o_8_132_0_0 = 0;
endmodule



// Benchmark "kernel_8_133" written by ABC on Sun Jul 19 10:05:20 2020

module kernel_8_133 ( 
    i_8_133_13_0, i_8_133_52_0, i_8_133_115_0, i_8_133_139_0,
    i_8_133_151_0, i_8_133_259_0, i_8_133_283_0, i_8_133_301_0,
    i_8_133_304_0, i_8_133_305_0, i_8_133_307_0, i_8_133_367_0,
    i_8_133_382_0, i_8_133_392_0, i_8_133_401_0, i_8_133_420_0,
    i_8_133_421_0, i_8_133_455_0, i_8_133_493_0, i_8_133_508_0,
    i_8_133_509_0, i_8_133_553_0, i_8_133_571_0, i_8_133_580_0,
    i_8_133_583_0, i_8_133_589_0, i_8_133_607_0, i_8_133_610_0,
    i_8_133_631_0, i_8_133_638_0, i_8_133_643_0, i_8_133_644_0,
    i_8_133_661_0, i_8_133_678_0, i_8_133_866_0, i_8_133_895_0,
    i_8_133_967_0, i_8_133_992_0, i_8_133_1012_0, i_8_133_1102_0,
    i_8_133_1103_0, i_8_133_1108_0, i_8_133_1111_0, i_8_133_1130_0,
    i_8_133_1157_0, i_8_133_1183_0, i_8_133_1201_0, i_8_133_1229_0,
    i_8_133_1246_0, i_8_133_1266_0, i_8_133_1267_0, i_8_133_1299_0,
    i_8_133_1301_0, i_8_133_1327_0, i_8_133_1328_0, i_8_133_1336_0,
    i_8_133_1355_0, i_8_133_1357_0, i_8_133_1435_0, i_8_133_1436_0,
    i_8_133_1441_0, i_8_133_1462_0, i_8_133_1463_0, i_8_133_1471_0,
    i_8_133_1477_0, i_8_133_1525_0, i_8_133_1526_0, i_8_133_1538_0,
    i_8_133_1541_0, i_8_133_1542_0, i_8_133_1552_0, i_8_133_1574_0,
    i_8_133_1632_0, i_8_133_1633_0, i_8_133_1642_0, i_8_133_1655_0,
    i_8_133_1678_0, i_8_133_1705_0, i_8_133_1749_0, i_8_133_1750_0,
    i_8_133_1753_0, i_8_133_1767_0, i_8_133_1776_0, i_8_133_1825_0,
    i_8_133_1841_0, i_8_133_1882_0, i_8_133_1894_0, i_8_133_1939_0,
    i_8_133_1940_0, i_8_133_1957_0, i_8_133_1958_0, i_8_133_1967_0,
    i_8_133_1975_0, i_8_133_1992_0, i_8_133_1995_0, i_8_133_1996_0,
    i_8_133_2136_0, i_8_133_2138_0, i_8_133_2210_0, i_8_133_2231_0,
    o_8_133_0_0  );
  input  i_8_133_13_0, i_8_133_52_0, i_8_133_115_0, i_8_133_139_0,
    i_8_133_151_0, i_8_133_259_0, i_8_133_283_0, i_8_133_301_0,
    i_8_133_304_0, i_8_133_305_0, i_8_133_307_0, i_8_133_367_0,
    i_8_133_382_0, i_8_133_392_0, i_8_133_401_0, i_8_133_420_0,
    i_8_133_421_0, i_8_133_455_0, i_8_133_493_0, i_8_133_508_0,
    i_8_133_509_0, i_8_133_553_0, i_8_133_571_0, i_8_133_580_0,
    i_8_133_583_0, i_8_133_589_0, i_8_133_607_0, i_8_133_610_0,
    i_8_133_631_0, i_8_133_638_0, i_8_133_643_0, i_8_133_644_0,
    i_8_133_661_0, i_8_133_678_0, i_8_133_866_0, i_8_133_895_0,
    i_8_133_967_0, i_8_133_992_0, i_8_133_1012_0, i_8_133_1102_0,
    i_8_133_1103_0, i_8_133_1108_0, i_8_133_1111_0, i_8_133_1130_0,
    i_8_133_1157_0, i_8_133_1183_0, i_8_133_1201_0, i_8_133_1229_0,
    i_8_133_1246_0, i_8_133_1266_0, i_8_133_1267_0, i_8_133_1299_0,
    i_8_133_1301_0, i_8_133_1327_0, i_8_133_1328_0, i_8_133_1336_0,
    i_8_133_1355_0, i_8_133_1357_0, i_8_133_1435_0, i_8_133_1436_0,
    i_8_133_1441_0, i_8_133_1462_0, i_8_133_1463_0, i_8_133_1471_0,
    i_8_133_1477_0, i_8_133_1525_0, i_8_133_1526_0, i_8_133_1538_0,
    i_8_133_1541_0, i_8_133_1542_0, i_8_133_1552_0, i_8_133_1574_0,
    i_8_133_1632_0, i_8_133_1633_0, i_8_133_1642_0, i_8_133_1655_0,
    i_8_133_1678_0, i_8_133_1705_0, i_8_133_1749_0, i_8_133_1750_0,
    i_8_133_1753_0, i_8_133_1767_0, i_8_133_1776_0, i_8_133_1825_0,
    i_8_133_1841_0, i_8_133_1882_0, i_8_133_1894_0, i_8_133_1939_0,
    i_8_133_1940_0, i_8_133_1957_0, i_8_133_1958_0, i_8_133_1967_0,
    i_8_133_1975_0, i_8_133_1992_0, i_8_133_1995_0, i_8_133_1996_0,
    i_8_133_2136_0, i_8_133_2138_0, i_8_133_2210_0, i_8_133_2231_0;
  output o_8_133_0_0;
  assign o_8_133_0_0 = 0;
endmodule



// Benchmark "kernel_8_134" written by ABC on Sun Jul 19 10:05:21 2020

module kernel_8_134 ( 
    i_8_134_20_0, i_8_134_31_0, i_8_134_35_0, i_8_134_50_0, i_8_134_55_0,
    i_8_134_103_0, i_8_134_104_0, i_8_134_115_0, i_8_134_142_0,
    i_8_134_167_0, i_8_134_181_0, i_8_134_221_0, i_8_134_232_0,
    i_8_134_233_0, i_8_134_253_0, i_8_134_255_0, i_8_134_289_0,
    i_8_134_292_0, i_8_134_293_0, i_8_134_297_0, i_8_134_306_0,
    i_8_134_343_0, i_8_134_344_0, i_8_134_378_0, i_8_134_386_0,
    i_8_134_414_0, i_8_134_442_0, i_8_134_451_0, i_8_134_476_0,
    i_8_134_479_0, i_8_134_481_0, i_8_134_482_0, i_8_134_484_0,
    i_8_134_497_0, i_8_134_526_0, i_8_134_588_0, i_8_134_589_0,
    i_8_134_595_0, i_8_134_596_0, i_8_134_612_0, i_8_134_689_0,
    i_8_134_706_0, i_8_134_713_0, i_8_134_760_0, i_8_134_761_0,
    i_8_134_766_0, i_8_134_767_0, i_8_134_784_0, i_8_134_787_0,
    i_8_134_797_0, i_8_134_811_0, i_8_134_812_0, i_8_134_838_0,
    i_8_134_847_0, i_8_134_850_0, i_8_134_859_0, i_8_134_929_0,
    i_8_134_992_0, i_8_134_1058_0, i_8_134_1118_0, i_8_134_1183_0,
    i_8_134_1189_0, i_8_134_1216_0, i_8_134_1219_0, i_8_134_1238_0,
    i_8_134_1264_0, i_8_134_1265_0, i_8_134_1269_0, i_8_134_1271_0,
    i_8_134_1282_0, i_8_134_1291_0, i_8_134_1300_0, i_8_134_1306_0,
    i_8_134_1315_0, i_8_134_1318_0, i_8_134_1404_0, i_8_134_1470_0,
    i_8_134_1540_0, i_8_134_1550_0, i_8_134_1557_0, i_8_134_1558_0,
    i_8_134_1560_0, i_8_134_1562_0, i_8_134_1621_0, i_8_134_1633_0,
    i_8_134_1730_0, i_8_134_1739_0, i_8_134_1762_0, i_8_134_1786_0,
    i_8_134_1787_0, i_8_134_1831_0, i_8_134_1873_0, i_8_134_1904_0,
    i_8_134_1949_0, i_8_134_2029_0, i_8_134_2037_0, i_8_134_2089_0,
    i_8_134_2090_0, i_8_134_2093_0, i_8_134_2287_0,
    o_8_134_0_0  );
  input  i_8_134_20_0, i_8_134_31_0, i_8_134_35_0, i_8_134_50_0,
    i_8_134_55_0, i_8_134_103_0, i_8_134_104_0, i_8_134_115_0,
    i_8_134_142_0, i_8_134_167_0, i_8_134_181_0, i_8_134_221_0,
    i_8_134_232_0, i_8_134_233_0, i_8_134_253_0, i_8_134_255_0,
    i_8_134_289_0, i_8_134_292_0, i_8_134_293_0, i_8_134_297_0,
    i_8_134_306_0, i_8_134_343_0, i_8_134_344_0, i_8_134_378_0,
    i_8_134_386_0, i_8_134_414_0, i_8_134_442_0, i_8_134_451_0,
    i_8_134_476_0, i_8_134_479_0, i_8_134_481_0, i_8_134_482_0,
    i_8_134_484_0, i_8_134_497_0, i_8_134_526_0, i_8_134_588_0,
    i_8_134_589_0, i_8_134_595_0, i_8_134_596_0, i_8_134_612_0,
    i_8_134_689_0, i_8_134_706_0, i_8_134_713_0, i_8_134_760_0,
    i_8_134_761_0, i_8_134_766_0, i_8_134_767_0, i_8_134_784_0,
    i_8_134_787_0, i_8_134_797_0, i_8_134_811_0, i_8_134_812_0,
    i_8_134_838_0, i_8_134_847_0, i_8_134_850_0, i_8_134_859_0,
    i_8_134_929_0, i_8_134_992_0, i_8_134_1058_0, i_8_134_1118_0,
    i_8_134_1183_0, i_8_134_1189_0, i_8_134_1216_0, i_8_134_1219_0,
    i_8_134_1238_0, i_8_134_1264_0, i_8_134_1265_0, i_8_134_1269_0,
    i_8_134_1271_0, i_8_134_1282_0, i_8_134_1291_0, i_8_134_1300_0,
    i_8_134_1306_0, i_8_134_1315_0, i_8_134_1318_0, i_8_134_1404_0,
    i_8_134_1470_0, i_8_134_1540_0, i_8_134_1550_0, i_8_134_1557_0,
    i_8_134_1558_0, i_8_134_1560_0, i_8_134_1562_0, i_8_134_1621_0,
    i_8_134_1633_0, i_8_134_1730_0, i_8_134_1739_0, i_8_134_1762_0,
    i_8_134_1786_0, i_8_134_1787_0, i_8_134_1831_0, i_8_134_1873_0,
    i_8_134_1904_0, i_8_134_1949_0, i_8_134_2029_0, i_8_134_2037_0,
    i_8_134_2089_0, i_8_134_2090_0, i_8_134_2093_0, i_8_134_2287_0;
  output o_8_134_0_0;
  assign o_8_134_0_0 = 0;
endmodule



// Benchmark "kernel_8_135" written by ABC on Sun Jul 19 10:05:21 2020

module kernel_8_135 ( 
    i_8_135_32_0, i_8_135_46_0, i_8_135_53_0, i_8_135_56_0, i_8_135_67_0,
    i_8_135_101_0, i_8_135_166_0, i_8_135_257_0, i_8_135_281_0,
    i_8_135_311_0, i_8_135_363_0, i_8_135_371_0, i_8_135_416_0,
    i_8_135_571_0, i_8_135_603_0, i_8_135_606_0, i_8_135_655_0,
    i_8_135_656_0, i_8_135_705_0, i_8_135_768_0, i_8_135_838_0,
    i_8_135_839_0, i_8_135_860_0, i_8_135_866_0, i_8_135_967_0,
    i_8_135_994_0, i_8_135_1056_0, i_8_135_1110_0, i_8_135_1111_0,
    i_8_135_1198_0, i_8_135_1217_0, i_8_135_1220_0, i_8_135_1229_0,
    i_8_135_1234_0, i_8_135_1265_0, i_8_135_1266_0, i_8_135_1267_0,
    i_8_135_1292_0, i_8_135_1318_0, i_8_135_1323_0, i_8_135_1326_0,
    i_8_135_1340_0, i_8_135_1351_0, i_8_135_1360_0, i_8_135_1367_0,
    i_8_135_1400_0, i_8_135_1427_0, i_8_135_1489_0, i_8_135_1504_0,
    i_8_135_1514_0, i_8_135_1522_0, i_8_135_1526_0, i_8_135_1548_0,
    i_8_135_1555_0, i_8_135_1557_0, i_8_135_1622_0, i_8_135_1630_0,
    i_8_135_1651_0, i_8_135_1665_0, i_8_135_1675_0, i_8_135_1684_0,
    i_8_135_1693_0, i_8_135_1703_0, i_8_135_1712_0, i_8_135_1757_0,
    i_8_135_1770_0, i_8_135_1777_0, i_8_135_1814_0, i_8_135_1818_0,
    i_8_135_1819_0, i_8_135_1820_0, i_8_135_1822_0, i_8_135_1825_0,
    i_8_135_1827_0, i_8_135_1856_0, i_8_135_1885_0, i_8_135_1891_0,
    i_8_135_1910_0, i_8_135_1966_0, i_8_135_1973_0, i_8_135_1975_0,
    i_8_135_1996_0, i_8_135_1997_0, i_8_135_2014_0, i_8_135_2097_0,
    i_8_135_2099_0, i_8_135_2128_0, i_8_135_2142_0, i_8_135_2146_0,
    i_8_135_2147_0, i_8_135_2148_0, i_8_135_2153_0, i_8_135_2197_0,
    i_8_135_2225_0, i_8_135_2244_0, i_8_135_2246_0, i_8_135_2258_0,
    i_8_135_2262_0, i_8_135_2272_0, i_8_135_2281_0,
    o_8_135_0_0  );
  input  i_8_135_32_0, i_8_135_46_0, i_8_135_53_0, i_8_135_56_0,
    i_8_135_67_0, i_8_135_101_0, i_8_135_166_0, i_8_135_257_0,
    i_8_135_281_0, i_8_135_311_0, i_8_135_363_0, i_8_135_371_0,
    i_8_135_416_0, i_8_135_571_0, i_8_135_603_0, i_8_135_606_0,
    i_8_135_655_0, i_8_135_656_0, i_8_135_705_0, i_8_135_768_0,
    i_8_135_838_0, i_8_135_839_0, i_8_135_860_0, i_8_135_866_0,
    i_8_135_967_0, i_8_135_994_0, i_8_135_1056_0, i_8_135_1110_0,
    i_8_135_1111_0, i_8_135_1198_0, i_8_135_1217_0, i_8_135_1220_0,
    i_8_135_1229_0, i_8_135_1234_0, i_8_135_1265_0, i_8_135_1266_0,
    i_8_135_1267_0, i_8_135_1292_0, i_8_135_1318_0, i_8_135_1323_0,
    i_8_135_1326_0, i_8_135_1340_0, i_8_135_1351_0, i_8_135_1360_0,
    i_8_135_1367_0, i_8_135_1400_0, i_8_135_1427_0, i_8_135_1489_0,
    i_8_135_1504_0, i_8_135_1514_0, i_8_135_1522_0, i_8_135_1526_0,
    i_8_135_1548_0, i_8_135_1555_0, i_8_135_1557_0, i_8_135_1622_0,
    i_8_135_1630_0, i_8_135_1651_0, i_8_135_1665_0, i_8_135_1675_0,
    i_8_135_1684_0, i_8_135_1693_0, i_8_135_1703_0, i_8_135_1712_0,
    i_8_135_1757_0, i_8_135_1770_0, i_8_135_1777_0, i_8_135_1814_0,
    i_8_135_1818_0, i_8_135_1819_0, i_8_135_1820_0, i_8_135_1822_0,
    i_8_135_1825_0, i_8_135_1827_0, i_8_135_1856_0, i_8_135_1885_0,
    i_8_135_1891_0, i_8_135_1910_0, i_8_135_1966_0, i_8_135_1973_0,
    i_8_135_1975_0, i_8_135_1996_0, i_8_135_1997_0, i_8_135_2014_0,
    i_8_135_2097_0, i_8_135_2099_0, i_8_135_2128_0, i_8_135_2142_0,
    i_8_135_2146_0, i_8_135_2147_0, i_8_135_2148_0, i_8_135_2153_0,
    i_8_135_2197_0, i_8_135_2225_0, i_8_135_2244_0, i_8_135_2246_0,
    i_8_135_2258_0, i_8_135_2262_0, i_8_135_2272_0, i_8_135_2281_0;
  output o_8_135_0_0;
  assign o_8_135_0_0 = 0;
endmodule



// Benchmark "kernel_8_136" written by ABC on Sun Jul 19 10:05:23 2020

module kernel_8_136 ( 
    i_8_136_140_0, i_8_136_147_0, i_8_136_148_0, i_8_136_149_0,
    i_8_136_150_0, i_8_136_151_0, i_8_136_165_0, i_8_136_166_0,
    i_8_136_189_0, i_8_136_192_0, i_8_136_194_0, i_8_136_195_0,
    i_8_136_211_0, i_8_136_214_0, i_8_136_226_0, i_8_136_227_0,
    i_8_136_271_0, i_8_136_303_0, i_8_136_368_0, i_8_136_386_0,
    i_8_136_427_0, i_8_136_453_0, i_8_136_454_0, i_8_136_472_0,
    i_8_136_483_0, i_8_136_484_0, i_8_136_493_0, i_8_136_508_0,
    i_8_136_530_0, i_8_136_582_0, i_8_136_602_0, i_8_136_618_0,
    i_8_136_642_0, i_8_136_657_0, i_8_136_658_0, i_8_136_661_0,
    i_8_136_678_0, i_8_136_701_0, i_8_136_703_0, i_8_136_705_0,
    i_8_136_732_0, i_8_136_750_0, i_8_136_751_0, i_8_136_752_0,
    i_8_136_832_0, i_8_136_833_0, i_8_136_861_0, i_8_136_1003_0,
    i_8_136_1157_0, i_8_136_1160_0, i_8_136_1164_0, i_8_136_1256_0,
    i_8_136_1285_0, i_8_136_1327_0, i_8_136_1335_0, i_8_136_1336_0,
    i_8_136_1355_0, i_8_136_1356_0, i_8_136_1357_0, i_8_136_1399_0,
    i_8_136_1434_0, i_8_136_1436_0, i_8_136_1438_0, i_8_136_1439_0,
    i_8_136_1479_0, i_8_136_1481_0, i_8_136_1488_0, i_8_136_1593_0,
    i_8_136_1596_0, i_8_136_1599_0, i_8_136_1623_0, i_8_136_1644_0,
    i_8_136_1660_0, i_8_136_1662_0, i_8_136_1663_0, i_8_136_1749_0,
    i_8_136_1754_0, i_8_136_1773_0, i_8_136_1776_0, i_8_136_1787_0,
    i_8_136_1824_0, i_8_136_1837_0, i_8_136_1875_0, i_8_136_1886_0,
    i_8_136_1919_0, i_8_136_2003_0, i_8_136_2011_0, i_8_136_2012_0,
    i_8_136_2089_0, i_8_136_2091_0, i_8_136_2095_0, i_8_136_2119_0,
    i_8_136_2154_0, i_8_136_2170_0, i_8_136_2174_0, i_8_136_2177_0,
    i_8_136_2253_0, i_8_136_2256_0, i_8_136_2257_0, i_8_136_2258_0,
    o_8_136_0_0  );
  input  i_8_136_140_0, i_8_136_147_0, i_8_136_148_0, i_8_136_149_0,
    i_8_136_150_0, i_8_136_151_0, i_8_136_165_0, i_8_136_166_0,
    i_8_136_189_0, i_8_136_192_0, i_8_136_194_0, i_8_136_195_0,
    i_8_136_211_0, i_8_136_214_0, i_8_136_226_0, i_8_136_227_0,
    i_8_136_271_0, i_8_136_303_0, i_8_136_368_0, i_8_136_386_0,
    i_8_136_427_0, i_8_136_453_0, i_8_136_454_0, i_8_136_472_0,
    i_8_136_483_0, i_8_136_484_0, i_8_136_493_0, i_8_136_508_0,
    i_8_136_530_0, i_8_136_582_0, i_8_136_602_0, i_8_136_618_0,
    i_8_136_642_0, i_8_136_657_0, i_8_136_658_0, i_8_136_661_0,
    i_8_136_678_0, i_8_136_701_0, i_8_136_703_0, i_8_136_705_0,
    i_8_136_732_0, i_8_136_750_0, i_8_136_751_0, i_8_136_752_0,
    i_8_136_832_0, i_8_136_833_0, i_8_136_861_0, i_8_136_1003_0,
    i_8_136_1157_0, i_8_136_1160_0, i_8_136_1164_0, i_8_136_1256_0,
    i_8_136_1285_0, i_8_136_1327_0, i_8_136_1335_0, i_8_136_1336_0,
    i_8_136_1355_0, i_8_136_1356_0, i_8_136_1357_0, i_8_136_1399_0,
    i_8_136_1434_0, i_8_136_1436_0, i_8_136_1438_0, i_8_136_1439_0,
    i_8_136_1479_0, i_8_136_1481_0, i_8_136_1488_0, i_8_136_1593_0,
    i_8_136_1596_0, i_8_136_1599_0, i_8_136_1623_0, i_8_136_1644_0,
    i_8_136_1660_0, i_8_136_1662_0, i_8_136_1663_0, i_8_136_1749_0,
    i_8_136_1754_0, i_8_136_1773_0, i_8_136_1776_0, i_8_136_1787_0,
    i_8_136_1824_0, i_8_136_1837_0, i_8_136_1875_0, i_8_136_1886_0,
    i_8_136_1919_0, i_8_136_2003_0, i_8_136_2011_0, i_8_136_2012_0,
    i_8_136_2089_0, i_8_136_2091_0, i_8_136_2095_0, i_8_136_2119_0,
    i_8_136_2154_0, i_8_136_2170_0, i_8_136_2174_0, i_8_136_2177_0,
    i_8_136_2253_0, i_8_136_2256_0, i_8_136_2257_0, i_8_136_2258_0;
  output o_8_136_0_0;
  assign o_8_136_0_0 = ~((i_8_136_140_0 & ((~i_8_136_149_0 & ~i_8_136_751_0 & ~i_8_136_1327_0 & ~i_8_136_1356_0 & ~i_8_136_2091_0 & ~i_8_136_2256_0) | (~i_8_136_151_0 & ~i_8_136_832_0 & ~i_8_136_1488_0 & ~i_8_136_2119_0 & ~i_8_136_2174_0 & ~i_8_136_2258_0))) | (~i_8_136_1875_0 & ((~i_8_136_148_0 & ~i_8_136_2011_0 & ((~i_8_136_195_0 & i_8_136_1327_0 & ~i_8_136_1593_0 & ~i_8_136_1644_0 & ~i_8_136_2091_0 & ~i_8_136_2095_0 & ~i_8_136_2177_0 & ~i_8_136_2256_0) | (~i_8_136_149_0 & i_8_136_194_0 & ~i_8_136_271_0 & ~i_8_136_732_0 & ~i_8_136_750_0 & ~i_8_136_1399_0 & ~i_8_136_1623_0 & ~i_8_136_1662_0 & i_8_136_1886_0 & ~i_8_136_2174_0 & ~i_8_136_2257_0))) | (~i_8_136_194_0 & ~i_8_136_227_0 & ((~i_8_136_192_0 & i_8_136_303_0 & ~i_8_136_732_0 & ~i_8_136_2012_0 & ~i_8_136_2091_0 & ~i_8_136_2256_0) | (~i_8_136_195_0 & ~i_8_136_701_0 & ~i_8_136_750_0 & ~i_8_136_752_0 & ~i_8_136_1164_0 & ~i_8_136_1355_0 & ~i_8_136_1593_0 & ~i_8_136_2095_0 & ~i_8_136_2257_0))) | (~i_8_136_1481_0 & ((~i_8_136_147_0 & ~i_8_136_150_0 & i_8_136_658_0 & ~i_8_136_833_0 & ~i_8_136_1773_0) | (~i_8_136_189_0 & i_8_136_453_0 & ~i_8_136_861_0 & ~i_8_136_1593_0 & ~i_8_136_1596_0 & ~i_8_136_1886_0 & ~i_8_136_2095_0 & ~i_8_136_2258_0))) | (~i_8_136_750_0 & ~i_8_136_1003_0 & ~i_8_136_1355_0 & i_8_136_1787_0 & ~i_8_136_2253_0 & ~i_8_136_2257_0))) | (~i_8_136_214_0 & ((~i_8_136_147_0 & ~i_8_136_151_0 & ~i_8_136_189_0 & ~i_8_136_472_0 & ~i_8_136_832_0 & ~i_8_136_833_0 & ~i_8_136_1164_0 & ~i_8_136_1355_0 & ~i_8_136_1356_0 & ~i_8_136_2012_0) | (i_8_136_1285_0 & i_8_136_1355_0 & i_8_136_1357_0 & ~i_8_136_1436_0 & ~i_8_136_2174_0 & ~i_8_136_2177_0 & ~i_8_136_2257_0))) | (~i_8_136_271_0 & ((~i_8_136_151_0 & i_8_136_427_0 & ~i_8_136_751_0 & ~i_8_136_832_0 & ~i_8_136_833_0 & ~i_8_136_1003_0 & ~i_8_136_1660_0 & ~i_8_136_1886_0 & ~i_8_136_2011_0 & ~i_8_136_2256_0) | (~i_8_136_150_0 & ~i_8_136_189_0 & ~i_8_136_192_0 & ~i_8_136_194_0 & ~i_8_136_618_0 & ~i_8_136_703_0 & ~i_8_136_732_0 & ~i_8_136_752_0 & ~i_8_136_1164_0 & ~i_8_136_1481_0 & ~i_8_136_2095_0 & ~i_8_136_2258_0 & ~i_8_136_1662_0 & ~i_8_136_2012_0))) | (~i_8_136_2091_0 & ((~i_8_136_192_0 & ((i_8_136_386_0 & ~i_8_136_703_0 & ~i_8_136_861_0 & ~i_8_136_1164_0 & ~i_8_136_1256_0 & ~i_8_136_1355_0 & ~i_8_136_1660_0 & ~i_8_136_1776_0) | (~i_8_136_147_0 & ~i_8_136_148_0 & ~i_8_136_151_0 & ~i_8_136_166_0 & ~i_8_136_194_0 & ~i_8_136_493_0 & ~i_8_136_751_0 & ~i_8_136_752_0 & ~i_8_136_833_0 & ~i_8_136_1357_0 & ~i_8_136_2089_0))) | (i_8_136_453_0 & i_8_136_454_0 & ~i_8_136_1599_0) | (~i_8_136_149_0 & ~i_8_136_194_0 & ~i_8_136_1660_0 & i_8_136_1754_0 & ~i_8_136_1824_0 & ~i_8_136_2257_0))) | (~i_8_136_148_0 & ((~i_8_136_189_0 & ~i_8_136_701_0 & ~i_8_136_832_0 & ~i_8_136_1003_0 & ~i_8_136_1355_0 & ~i_8_136_1357_0 & ~i_8_136_1662_0 & ~i_8_136_1663_0 & ~i_8_136_1824_0 & ~i_8_136_1886_0 & ~i_8_136_2089_0 & ~i_8_136_2170_0) | (~i_8_136_484_0 & ~i_8_136_703_0 & ~i_8_136_833_0 & ~i_8_136_861_0 & i_8_136_1434_0 & i_8_136_1749_0 & ~i_8_136_2012_0 & ~i_8_136_2253_0))) | (~i_8_136_833_0 & ((~i_8_136_2012_0 & ((~i_8_136_147_0 & ((~i_8_136_508_0 & ~i_8_136_703_0 & ~i_8_136_861_0 & i_8_136_1434_0 & ~i_8_136_1662_0 & ~i_8_136_1919_0 & ~i_8_136_2089_0) | (~i_8_136_149_0 & ~i_8_136_151_0 & ~i_8_136_227_0 & ~i_8_136_701_0 & ~i_8_136_732_0 & ~i_8_136_1356_0 & ~i_8_136_1488_0 & ~i_8_136_1660_0 & ~i_8_136_1663_0 & ~i_8_136_1773_0 & ~i_8_136_1837_0 & ~i_8_136_1886_0 & ~i_8_136_2256_0 & ~i_8_136_2258_0))) | (~i_8_136_151_0 & i_8_136_602_0 & ~i_8_136_1256_0 & ~i_8_136_2003_0 & ~i_8_136_2095_0))) | (~i_8_136_151_0 & ((i_8_136_484_0 & ~i_8_136_1596_0 & ~i_8_136_1599_0 & ~i_8_136_1660_0) | (~i_8_136_192_0 & ~i_8_136_368_0 & ~i_8_136_454_0 & ~i_8_136_661_0 & ~i_8_136_701_0 & ~i_8_136_732_0 & ~i_8_136_1164_0 & ~i_8_136_1623_0 & ~i_8_136_1824_0 & ~i_8_136_1837_0 & ~i_8_136_2089_0 & ~i_8_136_2154_0 & ~i_8_136_2174_0))) | (~i_8_136_149_0 & ~i_8_136_189_0 & ~i_8_136_192_0 & ~i_8_136_1399_0 & i_8_136_1439_0 & ~i_8_136_2177_0))) | (~i_8_136_1599_0 & ((~i_8_136_151_0 & ((~i_8_136_149_0 & i_8_136_1335_0 & i_8_136_1434_0 & ~i_8_136_1481_0) | (~i_8_136_703_0 & ~i_8_136_751_0 & ~i_8_136_752_0 & ~i_8_136_1164_0 & ~i_8_136_1285_0 & ~i_8_136_1357_0 & ~i_8_136_1663_0 & ~i_8_136_1749_0 & ~i_8_136_1773_0 & ~i_8_136_2095_0 & ~i_8_136_2154_0 & ~i_8_136_2258_0))) | (~i_8_136_189_0 & ~i_8_136_530_0 & ~i_8_136_1164_0 & i_8_136_1436_0 & i_8_136_1787_0 & ~i_8_136_2011_0))) | (~i_8_136_189_0 & ~i_8_136_832_0 & ((~i_8_136_149_0 & ~i_8_136_472_0 & ~i_8_136_1164_0 & ~i_8_136_1357_0 & i_8_136_1886_0 & ~i_8_136_2003_0) | (~i_8_136_226_0 & ~i_8_136_453_0 & ~i_8_136_732_0 & ~i_8_136_1285_0 & ~i_8_136_1355_0 & i_8_136_2089_0))) | (~i_8_136_149_0 & ((~i_8_136_147_0 & ~i_8_136_150_0 & i_8_136_454_0 & ~i_8_136_1399_0 & ~i_8_136_1663_0 & ~i_8_136_1773_0) | (~i_8_136_701_0 & ~i_8_136_750_0 & ~i_8_136_1164_0 & i_8_136_1436_0 & ~i_8_136_2012_0))) | (~i_8_136_150_0 & ((i_8_136_483_0 & ~i_8_136_493_0) | (~i_8_136_732_0 & ~i_8_136_1164_0 & i_8_136_1438_0 & ~i_8_136_2012_0 & ~i_8_136_2258_0))) | (~i_8_136_1327_0 & ~i_8_136_1357_0 & ((i_8_136_657_0 & ~i_8_136_1488_0 & i_8_136_2170_0) | (i_8_136_472_0 & i_8_136_602_0 & ~i_8_136_642_0 & ~i_8_136_705_0 & ~i_8_136_1481_0 & ~i_8_136_2257_0))) | (i_8_136_1157_0 & i_8_136_1336_0) | (i_8_136_1439_0 & i_8_136_2119_0 & ~i_8_136_2174_0) | (i_8_136_271_0 & ~i_8_136_703_0 & ~i_8_136_752_0 & ~i_8_136_1355_0 & ~i_8_136_1596_0 & ~i_8_136_1644_0 & ~i_8_136_2177_0 & ~i_8_136_2253_0));
endmodule



// Benchmark "kernel_8_137" written by ABC on Sun Jul 19 10:05:24 2020

module kernel_8_137 ( 
    i_8_137_33_0, i_8_137_85_0, i_8_137_114_0, i_8_137_141_0,
    i_8_137_159_0, i_8_137_165_0, i_8_137_186_0, i_8_137_204_0,
    i_8_137_220_0, i_8_137_222_0, i_8_137_223_0, i_8_137_230_0,
    i_8_137_231_0, i_8_137_240_0, i_8_137_298_0, i_8_137_420_0,
    i_8_137_476_0, i_8_137_501_0, i_8_137_546_0, i_8_137_549_0,
    i_8_137_550_0, i_8_137_609_0, i_8_137_625_0, i_8_137_636_0,
    i_8_137_700_0, i_8_137_762_0, i_8_137_777_0, i_8_137_780_0,
    i_8_137_824_0, i_8_137_825_0, i_8_137_834_0, i_8_137_868_0,
    i_8_137_870_0, i_8_137_877_0, i_8_137_878_0, i_8_137_879_0,
    i_8_137_888_0, i_8_137_895_0, i_8_137_949_0, i_8_137_991_0,
    i_8_137_993_0, i_8_137_994_0, i_8_137_995_0, i_8_137_1015_0,
    i_8_137_1027_0, i_8_137_1030_0, i_8_137_1073_0, i_8_137_1076_0,
    i_8_137_1086_0, i_8_137_1108_0, i_8_137_1112_0, i_8_137_1228_0,
    i_8_137_1266_0, i_8_137_1267_0, i_8_137_1281_0, i_8_137_1282_0,
    i_8_137_1284_0, i_8_137_1308_0, i_8_137_1329_0, i_8_137_1393_0,
    i_8_137_1402_0, i_8_137_1454_0, i_8_137_1470_0, i_8_137_1525_0,
    i_8_137_1527_0, i_8_137_1537_0, i_8_137_1544_0, i_8_137_1552_0,
    i_8_137_1553_0, i_8_137_1559_0, i_8_137_1653_0, i_8_137_1677_0,
    i_8_137_1678_0, i_8_137_1698_0, i_8_137_1705_0, i_8_137_1707_0,
    i_8_137_1721_0, i_8_137_1723_0, i_8_137_1725_0, i_8_137_1726_0,
    i_8_137_1729_0, i_8_137_1747_0, i_8_137_1779_0, i_8_137_1806_0,
    i_8_137_1808_0, i_8_137_1821_0, i_8_137_1834_0, i_8_137_1838_0,
    i_8_137_1867_0, i_8_137_1903_0, i_8_137_1948_0, i_8_137_2011_0,
    i_8_137_2046_0, i_8_137_2121_0, i_8_137_2139_0, i_8_137_2147_0,
    i_8_137_2149_0, i_8_137_2175_0, i_8_137_2214_0, i_8_137_2301_0,
    o_8_137_0_0  );
  input  i_8_137_33_0, i_8_137_85_0, i_8_137_114_0, i_8_137_141_0,
    i_8_137_159_0, i_8_137_165_0, i_8_137_186_0, i_8_137_204_0,
    i_8_137_220_0, i_8_137_222_0, i_8_137_223_0, i_8_137_230_0,
    i_8_137_231_0, i_8_137_240_0, i_8_137_298_0, i_8_137_420_0,
    i_8_137_476_0, i_8_137_501_0, i_8_137_546_0, i_8_137_549_0,
    i_8_137_550_0, i_8_137_609_0, i_8_137_625_0, i_8_137_636_0,
    i_8_137_700_0, i_8_137_762_0, i_8_137_777_0, i_8_137_780_0,
    i_8_137_824_0, i_8_137_825_0, i_8_137_834_0, i_8_137_868_0,
    i_8_137_870_0, i_8_137_877_0, i_8_137_878_0, i_8_137_879_0,
    i_8_137_888_0, i_8_137_895_0, i_8_137_949_0, i_8_137_991_0,
    i_8_137_993_0, i_8_137_994_0, i_8_137_995_0, i_8_137_1015_0,
    i_8_137_1027_0, i_8_137_1030_0, i_8_137_1073_0, i_8_137_1076_0,
    i_8_137_1086_0, i_8_137_1108_0, i_8_137_1112_0, i_8_137_1228_0,
    i_8_137_1266_0, i_8_137_1267_0, i_8_137_1281_0, i_8_137_1282_0,
    i_8_137_1284_0, i_8_137_1308_0, i_8_137_1329_0, i_8_137_1393_0,
    i_8_137_1402_0, i_8_137_1454_0, i_8_137_1470_0, i_8_137_1525_0,
    i_8_137_1527_0, i_8_137_1537_0, i_8_137_1544_0, i_8_137_1552_0,
    i_8_137_1553_0, i_8_137_1559_0, i_8_137_1653_0, i_8_137_1677_0,
    i_8_137_1678_0, i_8_137_1698_0, i_8_137_1705_0, i_8_137_1707_0,
    i_8_137_1721_0, i_8_137_1723_0, i_8_137_1725_0, i_8_137_1726_0,
    i_8_137_1729_0, i_8_137_1747_0, i_8_137_1779_0, i_8_137_1806_0,
    i_8_137_1808_0, i_8_137_1821_0, i_8_137_1834_0, i_8_137_1838_0,
    i_8_137_1867_0, i_8_137_1903_0, i_8_137_1948_0, i_8_137_2011_0,
    i_8_137_2046_0, i_8_137_2121_0, i_8_137_2139_0, i_8_137_2147_0,
    i_8_137_2149_0, i_8_137_2175_0, i_8_137_2214_0, i_8_137_2301_0;
  output o_8_137_0_0;
  assign o_8_137_0_0 = 0;
endmodule



// Benchmark "kernel_8_138" written by ABC on Sun Jul 19 10:05:26 2020

module kernel_8_138 ( 
    i_8_138_34_0, i_8_138_107_0, i_8_138_114_0, i_8_138_115_0,
    i_8_138_143_0, i_8_138_205_0, i_8_138_259_0, i_8_138_296_0,
    i_8_138_380_0, i_8_138_452_0, i_8_138_470_0, i_8_138_492_0,
    i_8_138_528_0, i_8_138_590_0, i_8_138_605_0, i_8_138_660_0,
    i_8_138_662_0, i_8_138_663_0, i_8_138_673_0, i_8_138_681_0,
    i_8_138_682_0, i_8_138_683_0, i_8_138_692_0, i_8_138_736_0,
    i_8_138_870_0, i_8_138_876_0, i_8_138_898_0, i_8_138_899_0,
    i_8_138_994_0, i_8_138_1026_0, i_8_138_1028_0, i_8_138_1075_0,
    i_8_138_1136_0, i_8_138_1157_0, i_8_138_1160_0, i_8_138_1224_0,
    i_8_138_1257_0, i_8_138_1258_0, i_8_138_1264_0, i_8_138_1273_0,
    i_8_138_1274_0, i_8_138_1276_0, i_8_138_1281_0, i_8_138_1340_0,
    i_8_138_1342_0, i_8_138_1343_0, i_8_138_1351_0, i_8_138_1355_0,
    i_8_138_1356_0, i_8_138_1403_0, i_8_138_1437_0, i_8_138_1438_0,
    i_8_138_1439_0, i_8_138_1444_0, i_8_138_1451_0, i_8_138_1489_0,
    i_8_138_1492_0, i_8_138_1503_0, i_8_138_1527_0, i_8_138_1529_0,
    i_8_138_1543_0, i_8_138_1562_0, i_8_138_1592_0, i_8_138_1599_0,
    i_8_138_1601_0, i_8_138_1603_0, i_8_138_1623_0, i_8_138_1625_0,
    i_8_138_1627_0, i_8_138_1628_0, i_8_138_1634_0, i_8_138_1636_0,
    i_8_138_1637_0, i_8_138_1645_0, i_8_138_1651_0, i_8_138_1675_0,
    i_8_138_1714_0, i_8_138_1716_0, i_8_138_1717_0, i_8_138_1748_0,
    i_8_138_1750_0, i_8_138_1751_0, i_8_138_1754_0, i_8_138_1818_0,
    i_8_138_1852_0, i_8_138_1857_0, i_8_138_1946_0, i_8_138_1964_0,
    i_8_138_1966_0, i_8_138_2128_0, i_8_138_2137_0, i_8_138_2138_0,
    i_8_138_2140_0, i_8_138_2141_0, i_8_138_2143_0, i_8_138_2144_0,
    i_8_138_2156_0, i_8_138_2214_0, i_8_138_2242_0, i_8_138_2288_0,
    o_8_138_0_0  );
  input  i_8_138_34_0, i_8_138_107_0, i_8_138_114_0, i_8_138_115_0,
    i_8_138_143_0, i_8_138_205_0, i_8_138_259_0, i_8_138_296_0,
    i_8_138_380_0, i_8_138_452_0, i_8_138_470_0, i_8_138_492_0,
    i_8_138_528_0, i_8_138_590_0, i_8_138_605_0, i_8_138_660_0,
    i_8_138_662_0, i_8_138_663_0, i_8_138_673_0, i_8_138_681_0,
    i_8_138_682_0, i_8_138_683_0, i_8_138_692_0, i_8_138_736_0,
    i_8_138_870_0, i_8_138_876_0, i_8_138_898_0, i_8_138_899_0,
    i_8_138_994_0, i_8_138_1026_0, i_8_138_1028_0, i_8_138_1075_0,
    i_8_138_1136_0, i_8_138_1157_0, i_8_138_1160_0, i_8_138_1224_0,
    i_8_138_1257_0, i_8_138_1258_0, i_8_138_1264_0, i_8_138_1273_0,
    i_8_138_1274_0, i_8_138_1276_0, i_8_138_1281_0, i_8_138_1340_0,
    i_8_138_1342_0, i_8_138_1343_0, i_8_138_1351_0, i_8_138_1355_0,
    i_8_138_1356_0, i_8_138_1403_0, i_8_138_1437_0, i_8_138_1438_0,
    i_8_138_1439_0, i_8_138_1444_0, i_8_138_1451_0, i_8_138_1489_0,
    i_8_138_1492_0, i_8_138_1503_0, i_8_138_1527_0, i_8_138_1529_0,
    i_8_138_1543_0, i_8_138_1562_0, i_8_138_1592_0, i_8_138_1599_0,
    i_8_138_1601_0, i_8_138_1603_0, i_8_138_1623_0, i_8_138_1625_0,
    i_8_138_1627_0, i_8_138_1628_0, i_8_138_1634_0, i_8_138_1636_0,
    i_8_138_1637_0, i_8_138_1645_0, i_8_138_1651_0, i_8_138_1675_0,
    i_8_138_1714_0, i_8_138_1716_0, i_8_138_1717_0, i_8_138_1748_0,
    i_8_138_1750_0, i_8_138_1751_0, i_8_138_1754_0, i_8_138_1818_0,
    i_8_138_1852_0, i_8_138_1857_0, i_8_138_1946_0, i_8_138_1964_0,
    i_8_138_1966_0, i_8_138_2128_0, i_8_138_2137_0, i_8_138_2138_0,
    i_8_138_2140_0, i_8_138_2141_0, i_8_138_2143_0, i_8_138_2144_0,
    i_8_138_2156_0, i_8_138_2214_0, i_8_138_2242_0, i_8_138_2288_0;
  output o_8_138_0_0;
  assign o_8_138_0_0 = ~((i_8_138_114_0 & ((i_8_138_115_0 & ~i_8_138_736_0 & ~i_8_138_870_0 & ~i_8_138_1028_0 & ~i_8_138_1403_0 & ~i_8_138_1637_0 & ~i_8_138_1714_0 & ~i_8_138_1946_0) | (~i_8_138_115_0 & ~i_8_138_663_0 & ~i_8_138_1224_0 & ~i_8_138_1343_0 & ~i_8_138_1603_0 & ~i_8_138_2140_0))) | (~i_8_138_1437_0 & ((~i_8_138_2138_0 & ((~i_8_138_205_0 & ((~i_8_138_692_0 & ~i_8_138_1136_0 & ~i_8_138_1340_0 & ~i_8_138_1342_0 & ~i_8_138_1489_0 & i_8_138_1625_0 & ~i_8_138_2137_0) | (~i_8_138_115_0 & ~i_8_138_1026_0 & ~i_8_138_1343_0 & ~i_8_138_1438_0 & ~i_8_138_1527_0 & ~i_8_138_1562_0 & ~i_8_138_1637_0 & i_8_138_1651_0 & ~i_8_138_1714_0 & ~i_8_138_1852_0 & ~i_8_138_2156_0 & ~i_8_138_2214_0))) | (~i_8_138_1342_0 & i_8_138_1503_0 & i_8_138_1543_0 & i_8_138_1675_0) | (~i_8_138_114_0 & ~i_8_138_380_0 & ~i_8_138_1264_0 & i_8_138_1356_0 & ~i_8_138_1754_0 & ~i_8_138_2156_0))) | (~i_8_138_1603_0 & ((~i_8_138_1342_0 & ((~i_8_138_452_0 & ~i_8_138_1028_0 & ((~i_8_138_470_0 & ~i_8_138_590_0 & ~i_8_138_662_0 & ~i_8_138_663_0 & ~i_8_138_683_0 & ~i_8_138_899_0 & ~i_8_138_994_0 & ~i_8_138_1026_0 & ~i_8_138_1340_0 & ~i_8_138_1562_0 & ~i_8_138_1625_0 & ~i_8_138_1675_0 & ~i_8_138_1748_0) | (~i_8_138_682_0 & ~i_8_138_898_0 & ~i_8_138_1075_0 & i_8_138_1355_0 & ~i_8_138_1503_0 & ~i_8_138_1637_0 & ~i_8_138_2140_0 & ~i_8_138_2156_0))) | (~i_8_138_590_0 & ~i_8_138_663_0 & ~i_8_138_1136_0 & ~i_8_138_1403_0 & ~i_8_138_1492_0 & ~i_8_138_1562_0 & ~i_8_138_1637_0 & ~i_8_138_1675_0 & ~i_8_138_1717_0 & ~i_8_138_1754_0 & ~i_8_138_1946_0 & ~i_8_138_1964_0 & ~i_8_138_1966_0))) | (~i_8_138_1136_0 & ~i_8_138_1281_0 & ~i_8_138_1439_0 & ~i_8_138_1754_0 & i_8_138_1852_0) | (~i_8_138_590_0 & i_8_138_876_0 & ~i_8_138_1224_0 & ~i_8_138_1343_0 & ~i_8_138_1356_0 & ~i_8_138_1444_0 & ~i_8_138_1946_0 & i_8_138_2242_0))) | (~i_8_138_2288_0 & ((~i_8_138_683_0 & ((~i_8_138_605_0 & ~i_8_138_899_0 & ~i_8_138_1026_0 & i_8_138_1492_0 & i_8_138_1645_0) | (~i_8_138_143_0 & ~i_8_138_681_0 & ~i_8_138_994_0 & ~i_8_138_1281_0 & ~i_8_138_1342_0 & ~i_8_138_1451_0 & ~i_8_138_1634_0 & ~i_8_138_1675_0 & ~i_8_138_1754_0 & ~i_8_138_1946_0 & ~i_8_138_1964_0 & ~i_8_138_2140_0 & ~i_8_138_2242_0))) | (~i_8_138_1157_0 & ~i_8_138_1438_0 & ~i_8_138_1439_0 & ~i_8_138_1451_0 & ~i_8_138_1492_0 & ~i_8_138_1543_0 & ~i_8_138_1637_0 & ~i_8_138_1675_0 & ~i_8_138_1717_0 & ~i_8_138_1964_0 & ~i_8_138_2140_0 & i_8_138_2156_0))) | (i_8_138_1264_0 & i_8_138_1503_0 & ~i_8_138_1748_0 & ~i_8_138_2143_0))) | (~i_8_138_114_0 & ((~i_8_138_663_0 & ~i_8_138_682_0 & ~i_8_138_1026_0 & ~i_8_138_1136_0 & i_8_138_1224_0 & ~i_8_138_1489_0 & ~i_8_138_1503_0 & ~i_8_138_1603_0 & ~i_8_138_1966_0) | (i_8_138_115_0 & ~i_8_138_470_0 & ~i_8_138_1281_0 & ~i_8_138_1351_0 & ~i_8_138_1438_0 & ~i_8_138_1562_0 & ~i_8_138_1818_0 & ~i_8_138_2141_0))) | (~i_8_138_660_0 & ((i_8_138_115_0 & ((~i_8_138_662_0 & ~i_8_138_681_0 & ~i_8_138_1028_0 & ~i_8_138_1136_0 & ~i_8_138_1340_0 & ~i_8_138_1529_0 & ~i_8_138_1637_0 & ~i_8_138_1675_0 & ~i_8_138_1716_0) | (~i_8_138_1160_0 & i_8_138_1438_0 & i_8_138_1439_0 & ~i_8_138_1562_0 & ~i_8_138_1636_0 & ~i_8_138_1748_0 & ~i_8_138_1852_0 & ~i_8_138_2214_0))) | (~i_8_138_1750_0 & ((~i_8_138_380_0 & ~i_8_138_1964_0 & ((~i_8_138_876_0 & ~i_8_138_1026_0 & i_8_138_1857_0 & ~i_8_138_2137_0) | (~i_8_138_681_0 & ~i_8_138_870_0 & ~i_8_138_1340_0 & ~i_8_138_1342_0 & ~i_8_138_1438_0 & ~i_8_138_1562_0 & ~i_8_138_1634_0 & ~i_8_138_1675_0 & ~i_8_138_1751_0 & ~i_8_138_1754_0 & ~i_8_138_2140_0))) | (~i_8_138_1637_0 & ((~i_8_138_662_0 & ~i_8_138_681_0 & ~i_8_138_452_0 & ~i_8_138_470_0 & ~i_8_138_1264_0 & ~i_8_138_1342_0 & ~i_8_138_1355_0 & ~i_8_138_1438_0 & ~i_8_138_1444_0 & ~i_8_138_1562_0 & ~i_8_138_1603_0 & ~i_8_138_1636_0 & ~i_8_138_1754_0 & ~i_8_138_2140_0 & ~i_8_138_1651_0 & ~i_8_138_1675_0) | (~i_8_138_736_0 & ~i_8_138_1026_0 & ~i_8_138_1075_0 & ~i_8_138_1343_0 & i_8_138_1966_0 & ~i_8_138_2137_0 & i_8_138_2144_0 & ~i_8_138_2214_0))))) | (~i_8_138_1342_0 & ((i_8_138_876_0 & i_8_138_1750_0 & i_8_138_1857_0 & ~i_8_138_2128_0) | (~i_8_138_107_0 & ~i_8_138_683_0 & ~i_8_138_692_0 & ~i_8_138_1026_0 & ~i_8_138_1224_0 & ~i_8_138_1343_0 & ~i_8_138_1651_0 & i_8_138_2214_0))))) | (~i_8_138_1675_0 & ((~i_8_138_1343_0 & ((~i_8_138_107_0 & ~i_8_138_1342_0 & ((i_8_138_452_0 & ~i_8_138_470_0 & ~i_8_138_1274_0 & ~i_8_138_1492_0 & ~i_8_138_1750_0 & ~i_8_138_2137_0 & i_8_138_2144_0) | (~i_8_138_692_0 & ~i_8_138_898_0 & ~i_8_138_899_0 & ~i_8_138_1026_0 & ~i_8_138_1444_0 & ~i_8_138_1451_0 & ~i_8_138_1529_0 & ~i_8_138_1716_0 & i_8_138_1852_0 & ~i_8_138_1857_0 & ~i_8_138_2288_0))) | (~i_8_138_663_0 & ((~i_8_138_682_0 & ~i_8_138_1451_0 & ~i_8_138_1603_0 & ~i_8_138_1751_0 & ((~i_8_138_605_0 & ~i_8_138_683_0 & ~i_8_138_899_0 & ~i_8_138_1160_0 & ~i_8_138_1340_0 & ~i_8_138_1714_0 & i_8_138_1966_0) | (~i_8_138_870_0 & ~i_8_138_898_0 & ~i_8_138_1351_0 & ~i_8_138_1438_0 & ~i_8_138_1439_0 & ~i_8_138_1750_0 & ~i_8_138_1966_0))) | (~i_8_138_380_0 & i_8_138_1492_0 & ~i_8_138_1562_0 & ~i_8_138_1716_0 & ~i_8_138_1717_0 & ~i_8_138_1754_0 & ~i_8_138_2141_0) | (~i_8_138_899_0 & ~i_8_138_1160_0 & i_8_138_1274_0 & ~i_8_138_1276_0 & ~i_8_138_1637_0 & ~i_8_138_1946_0 & ~i_8_138_2156_0))))) | (~i_8_138_662_0 & ~i_8_138_1562_0 & ((i_8_138_452_0 & ~i_8_138_1451_0 & ~i_8_138_1754_0 & ~i_8_138_1946_0 & ~i_8_138_2137_0 & ~i_8_138_2141_0) | (i_8_138_528_0 & ~i_8_138_870_0 & ~i_8_138_898_0 & ~i_8_138_1157_0 & ~i_8_138_1224_0 & ~i_8_138_1403_0 & ~i_8_138_1503_0 & ~i_8_138_1651_0 & ~i_8_138_1964_0 & ~i_8_138_1966_0 & ~i_8_138_2156_0))) | (~i_8_138_683_0 & ((~i_8_138_452_0 & ~i_8_138_681_0 & ~i_8_138_736_0 & ~i_8_138_870_0 & ~i_8_138_876_0 & ~i_8_138_898_0 & ~i_8_138_1136_0 & ~i_8_138_1157_0 & ~i_8_138_1340_0 & ~i_8_138_1403_0 & ~i_8_138_1492_0 & ~i_8_138_1623_0 & ~i_8_138_1634_0 & ~i_8_138_1716_0 & ~i_8_138_1748_0 & ~i_8_138_1750_0 & ~i_8_138_1751_0 & ~i_8_138_1946_0 & ~i_8_138_1964_0) | (~i_8_138_143_0 & i_8_138_590_0 & ~i_8_138_682_0 & ~i_8_138_692_0 & ~i_8_138_1026_0 & ~i_8_138_1451_0 & ~i_8_138_1714_0 & ~i_8_138_1717_0 & i_8_138_1754_0 & ~i_8_138_2140_0))) | (i_8_138_259_0 & ~i_8_138_380_0 & ~i_8_138_673_0 & ~i_8_138_898_0 & ~i_8_138_1281_0 & ~i_8_138_1342_0 & ~i_8_138_1964_0 & ~i_8_138_2140_0) | (~i_8_138_1439_0 & ~i_8_138_1754_0 & ~i_8_138_1946_0 & i_8_138_2128_0 & i_8_138_2144_0 & ~i_8_138_2288_0))) | (~i_8_138_107_0 & ((~i_8_138_34_0 & ~i_8_138_452_0 & i_8_138_492_0 & ~i_8_138_663_0 & ~i_8_138_683_0 & ~i_8_138_870_0 & i_8_138_1356_0 & ~i_8_138_1451_0 & ~i_8_138_1716_0) | (~i_8_138_1157_0 & i_8_138_1355_0 & ~i_8_138_1492_0 & ~i_8_138_1603_0 & ~i_8_138_1628_0 & ~i_8_138_1634_0 & ~i_8_138_1754_0 & ~i_8_138_1852_0 & ~i_8_138_1946_0 & ~i_8_138_2140_0))) | (~i_8_138_34_0 & ((~i_8_138_115_0 & ~i_8_138_143_0 & ~i_8_138_380_0 & ~i_8_138_662_0 & ~i_8_138_681_0 & ~i_8_138_1276_0 & ~i_8_138_1281_0 & ~i_8_138_1489_0 & i_8_138_1492_0 & ~i_8_138_1751_0 & ~i_8_138_1818_0) | (~i_8_138_663_0 & ~i_8_138_994_0 & ~i_8_138_1028_0 & i_8_138_1750_0 & ~i_8_138_1857_0 & ~i_8_138_1964_0 & i_8_138_1966_0 & i_8_138_2128_0 & ~i_8_138_2288_0))) | (~i_8_138_115_0 & ((~i_8_138_1028_0 & ~i_8_138_1342_0 & i_8_138_1543_0 & ~i_8_138_1750_0 & ~i_8_138_2140_0) | (~i_8_138_1274_0 & ~i_8_138_1281_0 & ~i_8_138_1343_0 & ~i_8_138_1438_0 & ~i_8_138_1717_0 & ~i_8_138_1751_0 & ~i_8_138_1754_0 & ~i_8_138_1857_0 & i_8_138_2128_0 & ~i_8_138_2288_0))) | (~i_8_138_380_0 & i_8_138_2144_0 & ((~i_8_138_590_0 & ~i_8_138_605_0 & ~i_8_138_1028_0 & ~i_8_138_1264_0 & ~i_8_138_1403_0 & ~i_8_138_1503_0 & ~i_8_138_2137_0) | (~i_8_138_899_0 & i_8_138_1273_0 & ~i_8_138_1439_0 & ~i_8_138_1852_0 & ~i_8_138_2141_0))) | (i_8_138_492_0 & ((i_8_138_1257_0 & i_8_138_1258_0 & ~i_8_138_1637_0) | (~i_8_138_1592_0 & i_8_138_1623_0 & ~i_8_138_1636_0 & i_8_138_1857_0 & ~i_8_138_1946_0))) | (~i_8_138_1946_0 & ((~i_8_138_528_0 & ((~i_8_138_470_0 & ~i_8_138_662_0 & ~i_8_138_870_0 & ~i_8_138_899_0 & ~i_8_138_1028_0 & ~i_8_138_1403_0 & ~i_8_138_1439_0 & ~i_8_138_1451_0 & ~i_8_138_1714_0 & ~i_8_138_1716_0 & ~i_8_138_1750_0 & i_8_138_1966_0 & ~i_8_138_2242_0) | (~i_8_138_681_0 & ~i_8_138_682_0 & i_8_138_1543_0 & ~i_8_138_1634_0 & i_8_138_1818_0 & ~i_8_138_2288_0))) | (~i_8_138_143_0 & ~i_8_138_662_0 & ~i_8_138_870_0 & ~i_8_138_1157_0 & ~i_8_138_1281_0 & ~i_8_138_1451_0 & i_8_138_1489_0 & ~i_8_138_1527_0 & ~i_8_138_1562_0 & ~i_8_138_1603_0 & ~i_8_138_2140_0 & ~i_8_138_2288_0))) | (~i_8_138_1343_0 & ((~i_8_138_1451_0 & ((~i_8_138_470_0 & ((~i_8_138_1026_0 & ~i_8_138_1157_0 & ~i_8_138_1264_0 & ~i_8_138_1439_0 & ~i_8_138_1489_0 & ~i_8_138_1750_0 & ~i_8_138_1754_0 & i_8_138_1966_0 & ~i_8_138_2137_0) | (~i_8_138_681_0 & ~i_8_138_899_0 & ~i_8_138_1562_0 & ~i_8_138_1717_0 & i_8_138_2128_0 & i_8_138_2143_0 & ~i_8_138_2288_0))) | (~i_8_138_452_0 & ~i_8_138_663_0 & ~i_8_138_682_0 & ~i_8_138_898_0 & i_8_138_1276_0 & ~i_8_138_1637_0 & ~i_8_138_1716_0) | (~i_8_138_870_0 & ~i_8_138_1028_0 & ~i_8_138_1157_0 & ~i_8_138_1438_0 & ~i_8_138_1489_0 & ~i_8_138_1562_0 & i_8_138_1750_0 & i_8_138_1751_0 & i_8_138_2137_0))) | (~i_8_138_663_0 & ~i_8_138_2138_0 & ((~i_8_138_259_0 & i_8_138_528_0 & ~i_8_138_682_0 & ~i_8_138_876_0 & ~i_8_138_1403_0 & ~i_8_138_1444_0 & ~i_8_138_1527_0 & ~i_8_138_1562_0 & ~i_8_138_1637_0 & ~i_8_138_1748_0 & ~i_8_138_1857_0) | (~i_8_138_1075_0 & ~i_8_138_1603_0 & i_8_138_1675_0 & ~i_8_138_1714_0 & ~i_8_138_1818_0 & i_8_138_2137_0 & ~i_8_138_2242_0 & ~i_8_138_2288_0))))) | (~i_8_138_899_0 & ((~i_8_138_1028_0 & ~i_8_138_1403_0 & ~i_8_138_605_0 & ~i_8_138_683_0 & ~i_8_138_1492_0 & ~i_8_138_1529_0 & i_8_138_1645_0 & ~i_8_138_1966_0) | (~i_8_138_870_0 & i_8_138_1592_0 & ~i_8_138_1748_0 & ~i_8_138_2138_0))) | (~i_8_138_1028_0 & ((~i_8_138_605_0 & ~i_8_138_1754_0 & ((~i_8_138_898_0 & ~i_8_138_994_0 & ~i_8_138_1026_0 & ~i_8_138_1157_0 & i_8_138_1264_0 & ~i_8_138_1340_0 & i_8_138_1489_0 & ~i_8_138_1492_0 & ~i_8_138_1562_0 & ~i_8_138_1637_0) | (i_8_138_1274_0 & ~i_8_138_1603_0 & ~i_8_138_1751_0 & ~i_8_138_2140_0 & ~i_8_138_2288_0))) | (~i_8_138_1751_0 & ((~i_8_138_1274_0 & ~i_8_138_1527_0 & i_8_138_1628_0 & ~i_8_138_1637_0 & ~i_8_138_1714_0 & ~i_8_138_1717_0) | (~i_8_138_470_0 & ~i_8_138_1026_0 & i_8_138_1224_0 & ~i_8_138_1438_0 & ~i_8_138_1716_0 & ~i_8_138_2140_0))))) | (i_8_138_1818_0 & ((~i_8_138_1751_0 & i_8_138_2143_0 & ((~i_8_138_590_0 & ~i_8_138_876_0 & ~i_8_138_1281_0 & ~i_8_138_1451_0 & ~i_8_138_1754_0 & ~i_8_138_2137_0 & ~i_8_138_2140_0) | (~i_8_138_1351_0 & ~i_8_138_1651_0 & ~i_8_138_2242_0))) | (~i_8_138_1342_0 & i_8_138_1437_0 & ~i_8_138_1438_0 & i_8_138_1750_0 & ~i_8_138_2137_0))) | (i_8_138_1257_0 & i_8_138_1651_0 & ~i_8_138_2140_0));
endmodule



// Benchmark "kernel_8_139" written by ABC on Sun Jul 19 10:05:26 2020

module kernel_8_139 ( 
    i_8_139_39_0, i_8_139_42_0, i_8_139_44_0, i_8_139_49_0, i_8_139_66_0,
    i_8_139_69_0, i_8_139_70_0, i_8_139_93_0, i_8_139_105_0, i_8_139_175_0,
    i_8_139_202_0, i_8_139_333_0, i_8_139_355_0, i_8_139_367_0,
    i_8_139_372_0, i_8_139_384_0, i_8_139_426_0, i_8_139_444_0,
    i_8_139_454_0, i_8_139_481_0, i_8_139_484_0, i_8_139_540_0,
    i_8_139_601_0, i_8_139_634_0, i_8_139_652_0, i_8_139_662_0,
    i_8_139_687_0, i_8_139_703_0, i_8_139_769_0, i_8_139_784_0,
    i_8_139_801_0, i_8_139_822_0, i_8_139_866_0, i_8_139_883_0,
    i_8_139_930_0, i_8_139_931_0, i_8_139_939_0, i_8_139_949_0,
    i_8_139_966_0, i_8_139_981_0, i_8_139_1071_0, i_8_139_1081_0,
    i_8_139_1096_0, i_8_139_1110_0, i_8_139_1135_0, i_8_139_1170_0,
    i_8_139_1213_0, i_8_139_1228_0, i_8_139_1233_0, i_8_139_1263_0,
    i_8_139_1267_0, i_8_139_1284_0, i_8_139_1290_0, i_8_139_1294_0,
    i_8_139_1410_0, i_8_139_1425_0, i_8_139_1470_0, i_8_139_1488_0,
    i_8_139_1497_0, i_8_139_1524_0, i_8_139_1596_0, i_8_139_1611_0,
    i_8_139_1648_0, i_8_139_1650_0, i_8_139_1659_0, i_8_139_1678_0,
    i_8_139_1689_0, i_8_139_1696_0, i_8_139_1704_0, i_8_139_1705_0,
    i_8_139_1747_0, i_8_139_1764_0, i_8_139_1777_0, i_8_139_1806_0,
    i_8_139_1807_0, i_8_139_1821_0, i_8_139_1869_0, i_8_139_1875_0,
    i_8_139_1882_0, i_8_139_1918_0, i_8_139_1919_0, i_8_139_1949_0,
    i_8_139_1972_0, i_8_139_1992_0, i_8_139_1995_0, i_8_139_2008_0,
    i_8_139_2010_0, i_8_139_2056_0, i_8_139_2089_0, i_8_139_2146_0,
    i_8_139_2148_0, i_8_139_2172_0, i_8_139_2179_0, i_8_139_2181_0,
    i_8_139_2182_0, i_8_139_2226_0, i_8_139_2241_0, i_8_139_2280_0,
    i_8_139_2281_0, i_8_139_2299_0,
    o_8_139_0_0  );
  input  i_8_139_39_0, i_8_139_42_0, i_8_139_44_0, i_8_139_49_0,
    i_8_139_66_0, i_8_139_69_0, i_8_139_70_0, i_8_139_93_0, i_8_139_105_0,
    i_8_139_175_0, i_8_139_202_0, i_8_139_333_0, i_8_139_355_0,
    i_8_139_367_0, i_8_139_372_0, i_8_139_384_0, i_8_139_426_0,
    i_8_139_444_0, i_8_139_454_0, i_8_139_481_0, i_8_139_484_0,
    i_8_139_540_0, i_8_139_601_0, i_8_139_634_0, i_8_139_652_0,
    i_8_139_662_0, i_8_139_687_0, i_8_139_703_0, i_8_139_769_0,
    i_8_139_784_0, i_8_139_801_0, i_8_139_822_0, i_8_139_866_0,
    i_8_139_883_0, i_8_139_930_0, i_8_139_931_0, i_8_139_939_0,
    i_8_139_949_0, i_8_139_966_0, i_8_139_981_0, i_8_139_1071_0,
    i_8_139_1081_0, i_8_139_1096_0, i_8_139_1110_0, i_8_139_1135_0,
    i_8_139_1170_0, i_8_139_1213_0, i_8_139_1228_0, i_8_139_1233_0,
    i_8_139_1263_0, i_8_139_1267_0, i_8_139_1284_0, i_8_139_1290_0,
    i_8_139_1294_0, i_8_139_1410_0, i_8_139_1425_0, i_8_139_1470_0,
    i_8_139_1488_0, i_8_139_1497_0, i_8_139_1524_0, i_8_139_1596_0,
    i_8_139_1611_0, i_8_139_1648_0, i_8_139_1650_0, i_8_139_1659_0,
    i_8_139_1678_0, i_8_139_1689_0, i_8_139_1696_0, i_8_139_1704_0,
    i_8_139_1705_0, i_8_139_1747_0, i_8_139_1764_0, i_8_139_1777_0,
    i_8_139_1806_0, i_8_139_1807_0, i_8_139_1821_0, i_8_139_1869_0,
    i_8_139_1875_0, i_8_139_1882_0, i_8_139_1918_0, i_8_139_1919_0,
    i_8_139_1949_0, i_8_139_1972_0, i_8_139_1992_0, i_8_139_1995_0,
    i_8_139_2008_0, i_8_139_2010_0, i_8_139_2056_0, i_8_139_2089_0,
    i_8_139_2146_0, i_8_139_2148_0, i_8_139_2172_0, i_8_139_2179_0,
    i_8_139_2181_0, i_8_139_2182_0, i_8_139_2226_0, i_8_139_2241_0,
    i_8_139_2280_0, i_8_139_2281_0, i_8_139_2299_0;
  output o_8_139_0_0;
  assign o_8_139_0_0 = 0;
endmodule



// Benchmark "kernel_8_140" written by ABC on Sun Jul 19 10:05:27 2020

module kernel_8_140 ( 
    i_8_140_31_0, i_8_140_77_0, i_8_140_89_0, i_8_140_161_0, i_8_140_170_0,
    i_8_140_224_0, i_8_140_229_0, i_8_140_233_0, i_8_140_259_0,
    i_8_140_305_0, i_8_140_347_0, i_8_140_359_0, i_8_140_366_0,
    i_8_140_458_0, i_8_140_481_0, i_8_140_493_0, i_8_140_525_0,
    i_8_140_526_0, i_8_140_530_0, i_8_140_557_0, i_8_140_593_0,
    i_8_140_601_0, i_8_140_604_0, i_8_140_663_0, i_8_140_665_0,
    i_8_140_692_0, i_8_140_698_0, i_8_140_699_0, i_8_140_719_0,
    i_8_140_763_0, i_8_140_826_0, i_8_140_827_0, i_8_140_845_0,
    i_8_140_869_0, i_8_140_880_0, i_8_140_896_0, i_8_140_974_0,
    i_8_140_994_0, i_8_140_1016_0, i_8_140_1031_0, i_8_140_1075_0,
    i_8_140_1097_0, i_8_140_1106_0, i_8_140_1115_0, i_8_140_1124_0,
    i_8_140_1133_0, i_8_140_1160_0, i_8_140_1184_0, i_8_140_1196_0,
    i_8_140_1232_0, i_8_140_1270_0, i_8_140_1277_0, i_8_140_1282_0,
    i_8_140_1285_0, i_8_140_1301_0, i_8_140_1349_0, i_8_140_1388_0,
    i_8_140_1441_0, i_8_140_1454_0, i_8_140_1457_0, i_8_140_1471_0,
    i_8_140_1472_0, i_8_140_1475_0, i_8_140_1484_0, i_8_140_1537_0,
    i_8_140_1546_0, i_8_140_1550_0, i_8_140_1553_0, i_8_140_1592_0,
    i_8_140_1633_0, i_8_140_1634_0, i_8_140_1636_0, i_8_140_1642_0,
    i_8_140_1647_0, i_8_140_1655_0, i_8_140_1678_0, i_8_140_1681_0,
    i_8_140_1682_0, i_8_140_1718_0, i_8_140_1733_0, i_8_140_1768_0,
    i_8_140_1807_0, i_8_140_1824_0, i_8_140_1826_0, i_8_140_1834_0,
    i_8_140_1840_0, i_8_140_1844_0, i_8_140_1870_0, i_8_140_1898_0,
    i_8_140_2008_0, i_8_140_2046_0, i_8_140_2111_0, i_8_140_2129_0,
    i_8_140_2132_0, i_8_140_2186_0, i_8_140_2194_0, i_8_140_2204_0,
    i_8_140_2249_0, i_8_140_2291_0, i_8_140_2294_0,
    o_8_140_0_0  );
  input  i_8_140_31_0, i_8_140_77_0, i_8_140_89_0, i_8_140_161_0,
    i_8_140_170_0, i_8_140_224_0, i_8_140_229_0, i_8_140_233_0,
    i_8_140_259_0, i_8_140_305_0, i_8_140_347_0, i_8_140_359_0,
    i_8_140_366_0, i_8_140_458_0, i_8_140_481_0, i_8_140_493_0,
    i_8_140_525_0, i_8_140_526_0, i_8_140_530_0, i_8_140_557_0,
    i_8_140_593_0, i_8_140_601_0, i_8_140_604_0, i_8_140_663_0,
    i_8_140_665_0, i_8_140_692_0, i_8_140_698_0, i_8_140_699_0,
    i_8_140_719_0, i_8_140_763_0, i_8_140_826_0, i_8_140_827_0,
    i_8_140_845_0, i_8_140_869_0, i_8_140_880_0, i_8_140_896_0,
    i_8_140_974_0, i_8_140_994_0, i_8_140_1016_0, i_8_140_1031_0,
    i_8_140_1075_0, i_8_140_1097_0, i_8_140_1106_0, i_8_140_1115_0,
    i_8_140_1124_0, i_8_140_1133_0, i_8_140_1160_0, i_8_140_1184_0,
    i_8_140_1196_0, i_8_140_1232_0, i_8_140_1270_0, i_8_140_1277_0,
    i_8_140_1282_0, i_8_140_1285_0, i_8_140_1301_0, i_8_140_1349_0,
    i_8_140_1388_0, i_8_140_1441_0, i_8_140_1454_0, i_8_140_1457_0,
    i_8_140_1471_0, i_8_140_1472_0, i_8_140_1475_0, i_8_140_1484_0,
    i_8_140_1537_0, i_8_140_1546_0, i_8_140_1550_0, i_8_140_1553_0,
    i_8_140_1592_0, i_8_140_1633_0, i_8_140_1634_0, i_8_140_1636_0,
    i_8_140_1642_0, i_8_140_1647_0, i_8_140_1655_0, i_8_140_1678_0,
    i_8_140_1681_0, i_8_140_1682_0, i_8_140_1718_0, i_8_140_1733_0,
    i_8_140_1768_0, i_8_140_1807_0, i_8_140_1824_0, i_8_140_1826_0,
    i_8_140_1834_0, i_8_140_1840_0, i_8_140_1844_0, i_8_140_1870_0,
    i_8_140_1898_0, i_8_140_2008_0, i_8_140_2046_0, i_8_140_2111_0,
    i_8_140_2129_0, i_8_140_2132_0, i_8_140_2186_0, i_8_140_2194_0,
    i_8_140_2204_0, i_8_140_2249_0, i_8_140_2291_0, i_8_140_2294_0;
  output o_8_140_0_0;
  assign o_8_140_0_0 = 0;
endmodule



// Benchmark "kernel_8_141" written by ABC on Sun Jul 19 10:05:28 2020

module kernel_8_141 ( 
    i_8_141_18_0, i_8_141_34_0, i_8_141_35_0, i_8_141_81_0, i_8_141_84_0,
    i_8_141_93_0, i_8_141_94_0, i_8_141_143_0, i_8_141_221_0,
    i_8_141_244_0, i_8_141_288_0, i_8_141_298_0, i_8_141_301_0,
    i_8_141_344_0, i_8_141_346_0, i_8_141_369_0, i_8_141_374_0,
    i_8_141_383_0, i_8_141_415_0, i_8_141_434_0, i_8_141_459_0,
    i_8_141_460_0, i_8_141_471_0, i_8_141_481_0, i_8_141_482_0,
    i_8_141_485_0, i_8_141_522_0, i_8_141_526_0, i_8_141_550_0,
    i_8_141_613_0, i_8_141_615_0, i_8_141_622_0, i_8_141_715_0,
    i_8_141_756_0, i_8_141_780_0, i_8_141_793_0, i_8_141_812_0,
    i_8_141_844_0, i_8_141_874_0, i_8_141_895_0, i_8_141_946_0,
    i_8_141_977_0, i_8_141_988_0, i_8_141_1028_0, i_8_141_1029_0,
    i_8_141_1113_0, i_8_141_1153_0, i_8_141_1156_0, i_8_141_1216_0,
    i_8_141_1233_0, i_8_141_1235_0, i_8_141_1251_0, i_8_141_1269_0,
    i_8_141_1270_0, i_8_141_1283_0, i_8_141_1300_0, i_8_141_1315_0,
    i_8_141_1337_0, i_8_141_1434_0, i_8_141_1444_0, i_8_141_1468_0,
    i_8_141_1549_0, i_8_141_1584_0, i_8_141_1586_0, i_8_141_1596_0,
    i_8_141_1597_0, i_8_141_1602_0, i_8_141_1612_0, i_8_141_1615_0,
    i_8_141_1630_0, i_8_141_1657_0, i_8_141_1666_0, i_8_141_1678_0,
    i_8_141_1679_0, i_8_141_1707_0, i_8_141_1743_0, i_8_141_1753_0,
    i_8_141_1754_0, i_8_141_1762_0, i_8_141_1780_0, i_8_141_1783_0,
    i_8_141_1794_0, i_8_141_1805_0, i_8_141_1840_0, i_8_141_1858_0,
    i_8_141_1859_0, i_8_141_1918_0, i_8_141_1946_0, i_8_141_1950_0,
    i_8_141_1963_0, i_8_141_2050_0, i_8_141_2073_0, i_8_141_2125_0,
    i_8_141_2126_0, i_8_141_2139_0, i_8_141_2140_0, i_8_141_2179_0,
    i_8_141_2183_0, i_8_141_2227_0, i_8_141_2290_0,
    o_8_141_0_0  );
  input  i_8_141_18_0, i_8_141_34_0, i_8_141_35_0, i_8_141_81_0,
    i_8_141_84_0, i_8_141_93_0, i_8_141_94_0, i_8_141_143_0, i_8_141_221_0,
    i_8_141_244_0, i_8_141_288_0, i_8_141_298_0, i_8_141_301_0,
    i_8_141_344_0, i_8_141_346_0, i_8_141_369_0, i_8_141_374_0,
    i_8_141_383_0, i_8_141_415_0, i_8_141_434_0, i_8_141_459_0,
    i_8_141_460_0, i_8_141_471_0, i_8_141_481_0, i_8_141_482_0,
    i_8_141_485_0, i_8_141_522_0, i_8_141_526_0, i_8_141_550_0,
    i_8_141_613_0, i_8_141_615_0, i_8_141_622_0, i_8_141_715_0,
    i_8_141_756_0, i_8_141_780_0, i_8_141_793_0, i_8_141_812_0,
    i_8_141_844_0, i_8_141_874_0, i_8_141_895_0, i_8_141_946_0,
    i_8_141_977_0, i_8_141_988_0, i_8_141_1028_0, i_8_141_1029_0,
    i_8_141_1113_0, i_8_141_1153_0, i_8_141_1156_0, i_8_141_1216_0,
    i_8_141_1233_0, i_8_141_1235_0, i_8_141_1251_0, i_8_141_1269_0,
    i_8_141_1270_0, i_8_141_1283_0, i_8_141_1300_0, i_8_141_1315_0,
    i_8_141_1337_0, i_8_141_1434_0, i_8_141_1444_0, i_8_141_1468_0,
    i_8_141_1549_0, i_8_141_1584_0, i_8_141_1586_0, i_8_141_1596_0,
    i_8_141_1597_0, i_8_141_1602_0, i_8_141_1612_0, i_8_141_1615_0,
    i_8_141_1630_0, i_8_141_1657_0, i_8_141_1666_0, i_8_141_1678_0,
    i_8_141_1679_0, i_8_141_1707_0, i_8_141_1743_0, i_8_141_1753_0,
    i_8_141_1754_0, i_8_141_1762_0, i_8_141_1780_0, i_8_141_1783_0,
    i_8_141_1794_0, i_8_141_1805_0, i_8_141_1840_0, i_8_141_1858_0,
    i_8_141_1859_0, i_8_141_1918_0, i_8_141_1946_0, i_8_141_1950_0,
    i_8_141_1963_0, i_8_141_2050_0, i_8_141_2073_0, i_8_141_2125_0,
    i_8_141_2126_0, i_8_141_2139_0, i_8_141_2140_0, i_8_141_2179_0,
    i_8_141_2183_0, i_8_141_2227_0, i_8_141_2290_0;
  output o_8_141_0_0;
  assign o_8_141_0_0 = 0;
endmodule



// Benchmark "kernel_8_142" written by ABC on Sun Jul 19 10:05:29 2020

module kernel_8_142 ( 
    i_8_142_12_0, i_8_142_22_0, i_8_142_28_0, i_8_142_52_0, i_8_142_67_0,
    i_8_142_75_0, i_8_142_79_0, i_8_142_136_0, i_8_142_222_0,
    i_8_142_225_0, i_8_142_321_0, i_8_142_333_0, i_8_142_360_0,
    i_8_142_364_0, i_8_142_366_0, i_8_142_367_0, i_8_142_381_0,
    i_8_142_391_0, i_8_142_397_0, i_8_142_398_0, i_8_142_400_0,
    i_8_142_418_0, i_8_142_426_0, i_8_142_427_0, i_8_142_430_0,
    i_8_142_454_0, i_8_142_507_0, i_8_142_516_0, i_8_142_526_0,
    i_8_142_571_0, i_8_142_604_0, i_8_142_634_0, i_8_142_639_0,
    i_8_142_661_0, i_8_142_747_0, i_8_142_750_0, i_8_142_784_0,
    i_8_142_849_0, i_8_142_850_0, i_8_142_860_0, i_8_142_937_0,
    i_8_142_969_0, i_8_142_970_0, i_8_142_971_0, i_8_142_973_0,
    i_8_142_1102_0, i_8_142_1107_0, i_8_142_1109_0, i_8_142_1144_0,
    i_8_142_1153_0, i_8_142_1162_0, i_8_142_1196_0, i_8_142_1201_0,
    i_8_142_1224_0, i_8_142_1297_0, i_8_142_1300_0, i_8_142_1327_0,
    i_8_142_1336_0, i_8_142_1362_0, i_8_142_1365_0, i_8_142_1399_0,
    i_8_142_1422_0, i_8_142_1432_0, i_8_142_1436_0, i_8_142_1441_0,
    i_8_142_1461_0, i_8_142_1471_0, i_8_142_1477_0, i_8_142_1480_0,
    i_8_142_1491_0, i_8_142_1513_0, i_8_142_1558_0, i_8_142_1615_0,
    i_8_142_1633_0, i_8_142_1679_0, i_8_142_1683_0, i_8_142_1692_0,
    i_8_142_1701_0, i_8_142_1705_0, i_8_142_1714_0, i_8_142_1750_0,
    i_8_142_1764_0, i_8_142_1768_0, i_8_142_1774_0, i_8_142_1809_0,
    i_8_142_1839_0, i_8_142_1849_0, i_8_142_1912_0, i_8_142_1917_0,
    i_8_142_1926_0, i_8_142_1935_0, i_8_142_1972_0, i_8_142_2070_0,
    i_8_142_2073_0, i_8_142_2134_0, i_8_142_2145_0, i_8_142_2155_0,
    i_8_142_2169_0, i_8_142_2242_0, i_8_142_2244_0,
    o_8_142_0_0  );
  input  i_8_142_12_0, i_8_142_22_0, i_8_142_28_0, i_8_142_52_0,
    i_8_142_67_0, i_8_142_75_0, i_8_142_79_0, i_8_142_136_0, i_8_142_222_0,
    i_8_142_225_0, i_8_142_321_0, i_8_142_333_0, i_8_142_360_0,
    i_8_142_364_0, i_8_142_366_0, i_8_142_367_0, i_8_142_381_0,
    i_8_142_391_0, i_8_142_397_0, i_8_142_398_0, i_8_142_400_0,
    i_8_142_418_0, i_8_142_426_0, i_8_142_427_0, i_8_142_430_0,
    i_8_142_454_0, i_8_142_507_0, i_8_142_516_0, i_8_142_526_0,
    i_8_142_571_0, i_8_142_604_0, i_8_142_634_0, i_8_142_639_0,
    i_8_142_661_0, i_8_142_747_0, i_8_142_750_0, i_8_142_784_0,
    i_8_142_849_0, i_8_142_850_0, i_8_142_860_0, i_8_142_937_0,
    i_8_142_969_0, i_8_142_970_0, i_8_142_971_0, i_8_142_973_0,
    i_8_142_1102_0, i_8_142_1107_0, i_8_142_1109_0, i_8_142_1144_0,
    i_8_142_1153_0, i_8_142_1162_0, i_8_142_1196_0, i_8_142_1201_0,
    i_8_142_1224_0, i_8_142_1297_0, i_8_142_1300_0, i_8_142_1327_0,
    i_8_142_1336_0, i_8_142_1362_0, i_8_142_1365_0, i_8_142_1399_0,
    i_8_142_1422_0, i_8_142_1432_0, i_8_142_1436_0, i_8_142_1441_0,
    i_8_142_1461_0, i_8_142_1471_0, i_8_142_1477_0, i_8_142_1480_0,
    i_8_142_1491_0, i_8_142_1513_0, i_8_142_1558_0, i_8_142_1615_0,
    i_8_142_1633_0, i_8_142_1679_0, i_8_142_1683_0, i_8_142_1692_0,
    i_8_142_1701_0, i_8_142_1705_0, i_8_142_1714_0, i_8_142_1750_0,
    i_8_142_1764_0, i_8_142_1768_0, i_8_142_1774_0, i_8_142_1809_0,
    i_8_142_1839_0, i_8_142_1849_0, i_8_142_1912_0, i_8_142_1917_0,
    i_8_142_1926_0, i_8_142_1935_0, i_8_142_1972_0, i_8_142_2070_0,
    i_8_142_2073_0, i_8_142_2134_0, i_8_142_2145_0, i_8_142_2155_0,
    i_8_142_2169_0, i_8_142_2242_0, i_8_142_2244_0;
  output o_8_142_0_0;
  assign o_8_142_0_0 = 0;
endmodule



// Benchmark "kernel_8_143" written by ABC on Sun Jul 19 10:05:30 2020

module kernel_8_143 ( 
    i_8_143_41_0, i_8_143_44_0, i_8_143_48_0, i_8_143_54_0, i_8_143_57_0,
    i_8_143_66_0, i_8_143_103_0, i_8_143_108_0, i_8_143_150_0,
    i_8_143_189_0, i_8_143_203_0, i_8_143_225_0, i_8_143_226_0,
    i_8_143_252_0, i_8_143_253_0, i_8_143_297_0, i_8_143_378_0,
    i_8_143_390_0, i_8_143_433_0, i_8_143_534_0, i_8_143_553_0,
    i_8_143_594_0, i_8_143_604_0, i_8_143_610_0, i_8_143_612_0,
    i_8_143_639_0, i_8_143_648_0, i_8_143_652_0, i_8_143_658_0,
    i_8_143_675_0, i_8_143_696_0, i_8_143_699_0, i_8_143_700_0,
    i_8_143_763_0, i_8_143_780_0, i_8_143_846_0, i_8_143_849_0,
    i_8_143_855_0, i_8_143_857_0, i_8_143_858_0, i_8_143_880_0,
    i_8_143_967_0, i_8_143_982_0, i_8_143_988_0, i_8_143_1032_0,
    i_8_143_1059_0, i_8_143_1083_0, i_8_143_1134_0, i_8_143_1137_0,
    i_8_143_1152_0, i_8_143_1157_0, i_8_143_1196_0, i_8_143_1263_0,
    i_8_143_1278_0, i_8_143_1281_0, i_8_143_1300_0, i_8_143_1314_0,
    i_8_143_1326_0, i_8_143_1354_0, i_8_143_1357_0, i_8_143_1383_0,
    i_8_143_1461_0, i_8_143_1473_0, i_8_143_1512_0, i_8_143_1530_0,
    i_8_143_1542_0, i_8_143_1557_0, i_8_143_1558_0, i_8_143_1602_0,
    i_8_143_1605_0, i_8_143_1623_0, i_8_143_1656_0, i_8_143_1674_0,
    i_8_143_1683_0, i_8_143_1695_0, i_8_143_1710_0, i_8_143_1713_0,
    i_8_143_1755_0, i_8_143_1759_0, i_8_143_1773_0, i_8_143_1791_0,
    i_8_143_1803_0, i_8_143_1809_0, i_8_143_1818_0, i_8_143_1885_0,
    i_8_143_1980_0, i_8_143_1990_0, i_8_143_1992_0, i_8_143_1993_0,
    i_8_143_1996_0, i_8_143_2052_0, i_8_143_2076_0, i_8_143_2109_0,
    i_8_143_2156_0, i_8_143_2161_0, i_8_143_2232_0, i_8_143_2233_0,
    i_8_143_2235_0, i_8_143_2244_0, i_8_143_2253_0,
    o_8_143_0_0  );
  input  i_8_143_41_0, i_8_143_44_0, i_8_143_48_0, i_8_143_54_0,
    i_8_143_57_0, i_8_143_66_0, i_8_143_103_0, i_8_143_108_0,
    i_8_143_150_0, i_8_143_189_0, i_8_143_203_0, i_8_143_225_0,
    i_8_143_226_0, i_8_143_252_0, i_8_143_253_0, i_8_143_297_0,
    i_8_143_378_0, i_8_143_390_0, i_8_143_433_0, i_8_143_534_0,
    i_8_143_553_0, i_8_143_594_0, i_8_143_604_0, i_8_143_610_0,
    i_8_143_612_0, i_8_143_639_0, i_8_143_648_0, i_8_143_652_0,
    i_8_143_658_0, i_8_143_675_0, i_8_143_696_0, i_8_143_699_0,
    i_8_143_700_0, i_8_143_763_0, i_8_143_780_0, i_8_143_846_0,
    i_8_143_849_0, i_8_143_855_0, i_8_143_857_0, i_8_143_858_0,
    i_8_143_880_0, i_8_143_967_0, i_8_143_982_0, i_8_143_988_0,
    i_8_143_1032_0, i_8_143_1059_0, i_8_143_1083_0, i_8_143_1134_0,
    i_8_143_1137_0, i_8_143_1152_0, i_8_143_1157_0, i_8_143_1196_0,
    i_8_143_1263_0, i_8_143_1278_0, i_8_143_1281_0, i_8_143_1300_0,
    i_8_143_1314_0, i_8_143_1326_0, i_8_143_1354_0, i_8_143_1357_0,
    i_8_143_1383_0, i_8_143_1461_0, i_8_143_1473_0, i_8_143_1512_0,
    i_8_143_1530_0, i_8_143_1542_0, i_8_143_1557_0, i_8_143_1558_0,
    i_8_143_1602_0, i_8_143_1605_0, i_8_143_1623_0, i_8_143_1656_0,
    i_8_143_1674_0, i_8_143_1683_0, i_8_143_1695_0, i_8_143_1710_0,
    i_8_143_1713_0, i_8_143_1755_0, i_8_143_1759_0, i_8_143_1773_0,
    i_8_143_1791_0, i_8_143_1803_0, i_8_143_1809_0, i_8_143_1818_0,
    i_8_143_1885_0, i_8_143_1980_0, i_8_143_1990_0, i_8_143_1992_0,
    i_8_143_1993_0, i_8_143_1996_0, i_8_143_2052_0, i_8_143_2076_0,
    i_8_143_2109_0, i_8_143_2156_0, i_8_143_2161_0, i_8_143_2232_0,
    i_8_143_2233_0, i_8_143_2235_0, i_8_143_2244_0, i_8_143_2253_0;
  output o_8_143_0_0;
  assign o_8_143_0_0 = ~((~i_8_143_44_0 & ((~i_8_143_57_0 & ~i_8_143_604_0 & ~i_8_143_639_0 & ~i_8_143_1602_0 & ~i_8_143_1605_0 & ~i_8_143_1990_0) | (~i_8_143_297_0 & ~i_8_143_594_0 & ~i_8_143_1134_0 & ~i_8_143_1542_0 & ~i_8_143_1818_0 & ~i_8_143_2156_0 & ~i_8_143_2244_0))) | (~i_8_143_1713_0 & ((~i_8_143_103_0 & ((i_8_143_658_0 & ~i_8_143_1674_0 & ~i_8_143_1980_0) | (~i_8_143_433_0 & i_8_143_612_0 & ~i_8_143_849_0 & ~i_8_143_1512_0 & i_8_143_1818_0 & ~i_8_143_2244_0))) | (~i_8_143_610_0 & ~i_8_143_675_0 & ~i_8_143_1980_0 & ~i_8_143_1992_0))) | (~i_8_143_433_0 & ((~i_8_143_226_0 & ~i_8_143_253_0 & ~i_8_143_1773_0 & ~i_8_143_1992_0) | (~i_8_143_41_0 & ~i_8_143_858_0 & ~i_8_143_1557_0 & ~i_8_143_1759_0 & i_8_143_1992_0 & ~i_8_143_2052_0 & ~i_8_143_2233_0))) | (i_8_143_534_0 & ((~i_8_143_1152_0 & ~i_8_143_1674_0) | (i_8_143_1152_0 & ~i_8_143_1993_0 & ~i_8_143_2156_0))) | (~i_8_143_553_0 & ((~i_8_143_855_0 & ~i_8_143_1152_0 & ~i_8_143_1281_0 & ~i_8_143_1530_0 & i_8_143_1557_0 & i_8_143_1993_0) | (~i_8_143_66_0 & i_8_143_880_0 & ~i_8_143_1300_0 & ~i_8_143_1326_0 & ~i_8_143_1656_0 & ~i_8_143_1683_0 & ~i_8_143_1755_0 & ~i_8_143_2232_0))) | (~i_8_143_849_0 & ((~i_8_143_54_0 & ~i_8_143_982_0 & ~i_8_143_1137_0 & i_8_143_1281_0 & ~i_8_143_1557_0) | (~i_8_143_48_0 & ~i_8_143_1134_0 & ~i_8_143_1558_0 & ~i_8_143_1710_0))) | (~i_8_143_1263_0 & ((~i_8_143_639_0 & ~i_8_143_696_0 & ~i_8_143_1137_0 & ~i_8_143_1152_0 & i_8_143_1326_0 & ~i_8_143_1357_0 & ~i_8_143_1755_0 & ~i_8_143_1996_0) | (~i_8_143_1059_0 & ~i_8_143_1710_0 & ~i_8_143_1990_0 & ~i_8_143_2244_0))) | (~i_8_143_1710_0 & ((~i_8_143_54_0 & ((i_8_143_612_0 & i_8_143_849_0 & ~i_8_143_1032_0 & ~i_8_143_1157_0) | (~i_8_143_612_0 & ~i_8_143_675_0 & ~i_8_143_1557_0))) | (i_8_143_54_0 & ~i_8_143_648_0 & ~i_8_143_855_0 & ~i_8_143_1557_0 & ~i_8_143_1809_0 & ~i_8_143_2233_0))) | (~i_8_143_54_0 & ((~i_8_143_658_0 & ~i_8_143_675_0 & i_8_143_1263_0 & ~i_8_143_1683_0 & ~i_8_143_1980_0) | (i_8_143_189_0 & ~i_8_143_610_0 & ~i_8_143_2233_0))) | (~i_8_143_57_0 & ~i_8_143_594_0 & ~i_8_143_675_0 & ~i_8_143_880_0 & ~i_8_143_1542_0 & ~i_8_143_1759_0 & ~i_8_143_2076_0 & ~i_8_143_2156_0));
endmodule



// Benchmark "kernel_8_144" written by ABC on Sun Jul 19 10:05:31 2020

module kernel_8_144 ( 
    i_8_144_11_0, i_8_144_35_0, i_8_144_49_0, i_8_144_59_0, i_8_144_77_0,
    i_8_144_111_0, i_8_144_226_0, i_8_144_229_0, i_8_144_230_0,
    i_8_144_231_0, i_8_144_282_0, i_8_144_293_0, i_8_144_310_0,
    i_8_144_325_0, i_8_144_337_0, i_8_144_342_0, i_8_144_343_0,
    i_8_144_345_0, i_8_144_364_0, i_8_144_370_0, i_8_144_373_0,
    i_8_144_423_0, i_8_144_443_0, i_8_144_450_0, i_8_144_454_0,
    i_8_144_479_0, i_8_144_481_0, i_8_144_482_0, i_8_144_499_0,
    i_8_144_505_0, i_8_144_522_0, i_8_144_526_0, i_8_144_544_0,
    i_8_144_549_0, i_8_144_554_0, i_8_144_613_0, i_8_144_662_0,
    i_8_144_687_0, i_8_144_688_0, i_8_144_697_0, i_8_144_704_0,
    i_8_144_715_0, i_8_144_769_0, i_8_144_783_0, i_8_144_786_0,
    i_8_144_795_0, i_8_144_815_0, i_8_144_832_0, i_8_144_840_0,
    i_8_144_875_0, i_8_144_931_0, i_8_144_932_0, i_8_144_954_0,
    i_8_144_955_0, i_8_144_973_0, i_8_144_985_0, i_8_144_1047_0,
    i_8_144_1057_0, i_8_144_1090_0, i_8_144_1099_0, i_8_144_1121_0,
    i_8_144_1123_0, i_8_144_1220_0, i_8_144_1243_0, i_8_144_1251_0,
    i_8_144_1266_0, i_8_144_1273_0, i_8_144_1274_0, i_8_144_1282_0,
    i_8_144_1305_0, i_8_144_1306_0, i_8_144_1328_0, i_8_144_1331_0,
    i_8_144_1346_0, i_8_144_1387_0, i_8_144_1401_0, i_8_144_1407_0,
    i_8_144_1537_0, i_8_144_1564_0, i_8_144_1571_0, i_8_144_1588_0,
    i_8_144_1612_0, i_8_144_1621_0, i_8_144_1629_0, i_8_144_1633_0,
    i_8_144_1651_0, i_8_144_1675_0, i_8_144_1721_0, i_8_144_1741_0,
    i_8_144_1804_0, i_8_144_1884_0, i_8_144_2003_0, i_8_144_2109_0,
    i_8_144_2145_0, i_8_144_2148_0, i_8_144_2191_0, i_8_144_2209_0,
    i_8_144_2215_0, i_8_144_2223_0, i_8_144_2289_0,
    o_8_144_0_0  );
  input  i_8_144_11_0, i_8_144_35_0, i_8_144_49_0, i_8_144_59_0,
    i_8_144_77_0, i_8_144_111_0, i_8_144_226_0, i_8_144_229_0,
    i_8_144_230_0, i_8_144_231_0, i_8_144_282_0, i_8_144_293_0,
    i_8_144_310_0, i_8_144_325_0, i_8_144_337_0, i_8_144_342_0,
    i_8_144_343_0, i_8_144_345_0, i_8_144_364_0, i_8_144_370_0,
    i_8_144_373_0, i_8_144_423_0, i_8_144_443_0, i_8_144_450_0,
    i_8_144_454_0, i_8_144_479_0, i_8_144_481_0, i_8_144_482_0,
    i_8_144_499_0, i_8_144_505_0, i_8_144_522_0, i_8_144_526_0,
    i_8_144_544_0, i_8_144_549_0, i_8_144_554_0, i_8_144_613_0,
    i_8_144_662_0, i_8_144_687_0, i_8_144_688_0, i_8_144_697_0,
    i_8_144_704_0, i_8_144_715_0, i_8_144_769_0, i_8_144_783_0,
    i_8_144_786_0, i_8_144_795_0, i_8_144_815_0, i_8_144_832_0,
    i_8_144_840_0, i_8_144_875_0, i_8_144_931_0, i_8_144_932_0,
    i_8_144_954_0, i_8_144_955_0, i_8_144_973_0, i_8_144_985_0,
    i_8_144_1047_0, i_8_144_1057_0, i_8_144_1090_0, i_8_144_1099_0,
    i_8_144_1121_0, i_8_144_1123_0, i_8_144_1220_0, i_8_144_1243_0,
    i_8_144_1251_0, i_8_144_1266_0, i_8_144_1273_0, i_8_144_1274_0,
    i_8_144_1282_0, i_8_144_1305_0, i_8_144_1306_0, i_8_144_1328_0,
    i_8_144_1331_0, i_8_144_1346_0, i_8_144_1387_0, i_8_144_1401_0,
    i_8_144_1407_0, i_8_144_1537_0, i_8_144_1564_0, i_8_144_1571_0,
    i_8_144_1588_0, i_8_144_1612_0, i_8_144_1621_0, i_8_144_1629_0,
    i_8_144_1633_0, i_8_144_1651_0, i_8_144_1675_0, i_8_144_1721_0,
    i_8_144_1741_0, i_8_144_1804_0, i_8_144_1884_0, i_8_144_2003_0,
    i_8_144_2109_0, i_8_144_2145_0, i_8_144_2148_0, i_8_144_2191_0,
    i_8_144_2209_0, i_8_144_2215_0, i_8_144_2223_0, i_8_144_2289_0;
  output o_8_144_0_0;
  assign o_8_144_0_0 = 0;
endmodule



// Benchmark "kernel_8_145" written by ABC on Sun Jul 19 10:05:32 2020

module kernel_8_145 ( 
    i_8_145_24_0, i_8_145_52_0, i_8_145_67_0, i_8_145_165_0, i_8_145_210_0,
    i_8_145_231_0, i_8_145_232_0, i_8_145_301_0, i_8_145_310_0,
    i_8_145_325_0, i_8_145_336_0, i_8_145_342_0, i_8_145_349_0,
    i_8_145_354_0, i_8_145_363_0, i_8_145_366_0, i_8_145_367_0,
    i_8_145_426_0, i_8_145_430_0, i_8_145_475_0, i_8_145_492_0,
    i_8_145_498_0, i_8_145_529_0, i_8_145_552_0, i_8_145_580_0,
    i_8_145_588_0, i_8_145_598_0, i_8_145_604_0, i_8_145_606_0,
    i_8_145_607_0, i_8_145_609_0, i_8_145_610_0, i_8_145_612_0,
    i_8_145_615_0, i_8_145_651_0, i_8_145_660_0, i_8_145_681_0,
    i_8_145_702_0, i_8_145_735_0, i_8_145_768_0, i_8_145_780_0,
    i_8_145_795_0, i_8_145_876_0, i_8_145_921_0, i_8_145_927_0,
    i_8_145_958_0, i_8_145_1020_0, i_8_145_1053_0, i_8_145_1068_0,
    i_8_145_1074_0, i_8_145_1101_0, i_8_145_1156_0, i_8_145_1170_0,
    i_8_145_1173_0, i_8_145_1228_0, i_8_145_1236_0, i_8_145_1251_0,
    i_8_145_1254_0, i_8_145_1291_0, i_8_145_1292_0, i_8_145_1311_0,
    i_8_145_1317_0, i_8_145_1354_0, i_8_145_1454_0, i_8_145_1470_0,
    i_8_145_1489_0, i_8_145_1524_0, i_8_145_1560_0, i_8_145_1623_0,
    i_8_145_1641_0, i_8_145_1649_0, i_8_145_1650_0, i_8_145_1678_0,
    i_8_145_1704_0, i_8_145_1707_0, i_8_145_1800_0, i_8_145_1819_0,
    i_8_145_1821_0, i_8_145_1824_0, i_8_145_1825_0, i_8_145_1861_0,
    i_8_145_1884_0, i_8_145_1941_0, i_8_145_1966_0, i_8_145_2001_0,
    i_8_145_2004_0, i_8_145_2016_0, i_8_145_2019_0, i_8_145_2020_0,
    i_8_145_2037_0, i_8_145_2073_0, i_8_145_2113_0, i_8_145_2146_0,
    i_8_145_2181_0, i_8_145_2199_0, i_8_145_2208_0, i_8_145_2209_0,
    i_8_145_2226_0, i_8_145_2235_0, i_8_145_2244_0,
    o_8_145_0_0  );
  input  i_8_145_24_0, i_8_145_52_0, i_8_145_67_0, i_8_145_165_0,
    i_8_145_210_0, i_8_145_231_0, i_8_145_232_0, i_8_145_301_0,
    i_8_145_310_0, i_8_145_325_0, i_8_145_336_0, i_8_145_342_0,
    i_8_145_349_0, i_8_145_354_0, i_8_145_363_0, i_8_145_366_0,
    i_8_145_367_0, i_8_145_426_0, i_8_145_430_0, i_8_145_475_0,
    i_8_145_492_0, i_8_145_498_0, i_8_145_529_0, i_8_145_552_0,
    i_8_145_580_0, i_8_145_588_0, i_8_145_598_0, i_8_145_604_0,
    i_8_145_606_0, i_8_145_607_0, i_8_145_609_0, i_8_145_610_0,
    i_8_145_612_0, i_8_145_615_0, i_8_145_651_0, i_8_145_660_0,
    i_8_145_681_0, i_8_145_702_0, i_8_145_735_0, i_8_145_768_0,
    i_8_145_780_0, i_8_145_795_0, i_8_145_876_0, i_8_145_921_0,
    i_8_145_927_0, i_8_145_958_0, i_8_145_1020_0, i_8_145_1053_0,
    i_8_145_1068_0, i_8_145_1074_0, i_8_145_1101_0, i_8_145_1156_0,
    i_8_145_1170_0, i_8_145_1173_0, i_8_145_1228_0, i_8_145_1236_0,
    i_8_145_1251_0, i_8_145_1254_0, i_8_145_1291_0, i_8_145_1292_0,
    i_8_145_1311_0, i_8_145_1317_0, i_8_145_1354_0, i_8_145_1454_0,
    i_8_145_1470_0, i_8_145_1489_0, i_8_145_1524_0, i_8_145_1560_0,
    i_8_145_1623_0, i_8_145_1641_0, i_8_145_1649_0, i_8_145_1650_0,
    i_8_145_1678_0, i_8_145_1704_0, i_8_145_1707_0, i_8_145_1800_0,
    i_8_145_1819_0, i_8_145_1821_0, i_8_145_1824_0, i_8_145_1825_0,
    i_8_145_1861_0, i_8_145_1884_0, i_8_145_1941_0, i_8_145_1966_0,
    i_8_145_2001_0, i_8_145_2004_0, i_8_145_2016_0, i_8_145_2019_0,
    i_8_145_2020_0, i_8_145_2037_0, i_8_145_2073_0, i_8_145_2113_0,
    i_8_145_2146_0, i_8_145_2181_0, i_8_145_2199_0, i_8_145_2208_0,
    i_8_145_2209_0, i_8_145_2226_0, i_8_145_2235_0, i_8_145_2244_0;
  output o_8_145_0_0;
  assign o_8_145_0_0 = 0;
endmodule



// Benchmark "kernel_8_146" written by ABC on Sun Jul 19 10:05:33 2020

module kernel_8_146 ( 
    i_8_146_4_0, i_8_146_13_0, i_8_146_22_0, i_8_146_53_0, i_8_146_67_0,
    i_8_146_97_0, i_8_146_184_0, i_8_146_239_0, i_8_146_246_0,
    i_8_146_263_0, i_8_146_298_0, i_8_146_327_0, i_8_146_364_0,
    i_8_146_365_0, i_8_146_368_0, i_8_146_437_0, i_8_146_455_0,
    i_8_146_464_0, i_8_146_473_0, i_8_146_507_0, i_8_146_517_0,
    i_8_146_518_0, i_8_146_534_0, i_8_146_535_0, i_8_146_553_0,
    i_8_146_571_0, i_8_146_589_0, i_8_146_592_0, i_8_146_595_0,
    i_8_146_615_0, i_8_146_624_0, i_8_146_632_0, i_8_146_634_0,
    i_8_146_652_0, i_8_146_660_0, i_8_146_661_0, i_8_146_663_0,
    i_8_146_665_0, i_8_146_682_0, i_8_146_706_0, i_8_146_751_0,
    i_8_146_841_0, i_8_146_869_0, i_8_146_938_0, i_8_146_941_0,
    i_8_146_958_0, i_8_146_965_0, i_8_146_977_0, i_8_146_1039_0,
    i_8_146_1042_0, i_8_146_1079_0, i_8_146_1102_0, i_8_146_1111_0,
    i_8_146_1122_0, i_8_146_1169_0, i_8_146_1210_0, i_8_146_1222_0,
    i_8_146_1223_0, i_8_146_1249_0, i_8_146_1267_0, i_8_146_1303_0,
    i_8_146_1318_0, i_8_146_1354_0, i_8_146_1381_0, i_8_146_1384_0,
    i_8_146_1397_0, i_8_146_1438_0, i_8_146_1456_0, i_8_146_1458_0,
    i_8_146_1469_0, i_8_146_1489_0, i_8_146_1513_0, i_8_146_1528_0,
    i_8_146_1532_0, i_8_146_1564_0, i_8_146_1641_0, i_8_146_1659_0,
    i_8_146_1687_0, i_8_146_1697_0, i_8_146_1729_0, i_8_146_1767_0,
    i_8_146_1774_0, i_8_146_1813_0, i_8_146_1824_0, i_8_146_1825_0,
    i_8_146_1826_0, i_8_146_1884_0, i_8_146_1885_0, i_8_146_1957_0,
    i_8_146_1992_0, i_8_146_1995_0, i_8_146_1996_0, i_8_146_2115_0,
    i_8_146_2119_0, i_8_146_2146_0, i_8_146_2226_0, i_8_146_2236_0,
    i_8_146_2242_0, i_8_146_2248_0, i_8_146_2299_0,
    o_8_146_0_0  );
  input  i_8_146_4_0, i_8_146_13_0, i_8_146_22_0, i_8_146_53_0,
    i_8_146_67_0, i_8_146_97_0, i_8_146_184_0, i_8_146_239_0,
    i_8_146_246_0, i_8_146_263_0, i_8_146_298_0, i_8_146_327_0,
    i_8_146_364_0, i_8_146_365_0, i_8_146_368_0, i_8_146_437_0,
    i_8_146_455_0, i_8_146_464_0, i_8_146_473_0, i_8_146_507_0,
    i_8_146_517_0, i_8_146_518_0, i_8_146_534_0, i_8_146_535_0,
    i_8_146_553_0, i_8_146_571_0, i_8_146_589_0, i_8_146_592_0,
    i_8_146_595_0, i_8_146_615_0, i_8_146_624_0, i_8_146_632_0,
    i_8_146_634_0, i_8_146_652_0, i_8_146_660_0, i_8_146_661_0,
    i_8_146_663_0, i_8_146_665_0, i_8_146_682_0, i_8_146_706_0,
    i_8_146_751_0, i_8_146_841_0, i_8_146_869_0, i_8_146_938_0,
    i_8_146_941_0, i_8_146_958_0, i_8_146_965_0, i_8_146_977_0,
    i_8_146_1039_0, i_8_146_1042_0, i_8_146_1079_0, i_8_146_1102_0,
    i_8_146_1111_0, i_8_146_1122_0, i_8_146_1169_0, i_8_146_1210_0,
    i_8_146_1222_0, i_8_146_1223_0, i_8_146_1249_0, i_8_146_1267_0,
    i_8_146_1303_0, i_8_146_1318_0, i_8_146_1354_0, i_8_146_1381_0,
    i_8_146_1384_0, i_8_146_1397_0, i_8_146_1438_0, i_8_146_1456_0,
    i_8_146_1458_0, i_8_146_1469_0, i_8_146_1489_0, i_8_146_1513_0,
    i_8_146_1528_0, i_8_146_1532_0, i_8_146_1564_0, i_8_146_1641_0,
    i_8_146_1659_0, i_8_146_1687_0, i_8_146_1697_0, i_8_146_1729_0,
    i_8_146_1767_0, i_8_146_1774_0, i_8_146_1813_0, i_8_146_1824_0,
    i_8_146_1825_0, i_8_146_1826_0, i_8_146_1884_0, i_8_146_1885_0,
    i_8_146_1957_0, i_8_146_1992_0, i_8_146_1995_0, i_8_146_1996_0,
    i_8_146_2115_0, i_8_146_2119_0, i_8_146_2146_0, i_8_146_2226_0,
    i_8_146_2236_0, i_8_146_2242_0, i_8_146_2248_0, i_8_146_2299_0;
  output o_8_146_0_0;
  assign o_8_146_0_0 = 0;
endmodule



// Benchmark "kernel_8_147" written by ABC on Sun Jul 19 10:05:34 2020

module kernel_8_147 ( 
    i_8_147_28_0, i_8_147_97_0, i_8_147_98_0, i_8_147_136_0, i_8_147_224_0,
    i_8_147_356_0, i_8_147_370_0, i_8_147_376_0, i_8_147_424_0,
    i_8_147_426_0, i_8_147_427_0, i_8_147_463_0, i_8_147_475_0,
    i_8_147_476_0, i_8_147_488_0, i_8_147_491_0, i_8_147_493_0,
    i_8_147_502_0, i_8_147_563_0, i_8_147_570_0, i_8_147_592_0,
    i_8_147_625_0, i_8_147_632_0, i_8_147_666_0, i_8_147_679_0,
    i_8_147_683_0, i_8_147_696_0, i_8_147_697_0, i_8_147_705_0,
    i_8_147_725_0, i_8_147_757_0, i_8_147_773_0, i_8_147_778_0,
    i_8_147_781_0, i_8_147_783_0, i_8_147_786_0, i_8_147_787_0,
    i_8_147_790_0, i_8_147_812_0, i_8_147_826_0, i_8_147_829_0,
    i_8_147_838_0, i_8_147_841_0, i_8_147_842_0, i_8_147_847_0,
    i_8_147_848_0, i_8_147_869_0, i_8_147_874_0, i_8_147_917_0,
    i_8_147_932_0, i_8_147_1000_0, i_8_147_1057_0, i_8_147_1072_0,
    i_8_147_1135_0, i_8_147_1189_0, i_8_147_1234_0, i_8_147_1271_0,
    i_8_147_1328_0, i_8_147_1363_0, i_8_147_1369_0, i_8_147_1454_0,
    i_8_147_1457_0, i_8_147_1470_0, i_8_147_1524_0, i_8_147_1589_0,
    i_8_147_1607_0, i_8_147_1648_0, i_8_147_1655_0, i_8_147_1684_0,
    i_8_147_1696_0, i_8_147_1700_0, i_8_147_1729_0, i_8_147_1732_0,
    i_8_147_1749_0, i_8_147_1805_0, i_8_147_1846_0, i_8_147_1855_0,
    i_8_147_1856_0, i_8_147_1857_0, i_8_147_1858_0, i_8_147_1859_0,
    i_8_147_1861_0, i_8_147_1867_0, i_8_147_1888_0, i_8_147_1895_0,
    i_8_147_1898_0, i_8_147_1904_0, i_8_147_1981_0, i_8_147_2029_0,
    i_8_147_2072_0, i_8_147_2090_0, i_8_147_2174_0, i_8_147_2182_0,
    i_8_147_2183_0, i_8_147_2185_0, i_8_147_2191_0, i_8_147_2280_0,
    i_8_147_2290_0, i_8_147_2292_0, i_8_147_2294_0,
    o_8_147_0_0  );
  input  i_8_147_28_0, i_8_147_97_0, i_8_147_98_0, i_8_147_136_0,
    i_8_147_224_0, i_8_147_356_0, i_8_147_370_0, i_8_147_376_0,
    i_8_147_424_0, i_8_147_426_0, i_8_147_427_0, i_8_147_463_0,
    i_8_147_475_0, i_8_147_476_0, i_8_147_488_0, i_8_147_491_0,
    i_8_147_493_0, i_8_147_502_0, i_8_147_563_0, i_8_147_570_0,
    i_8_147_592_0, i_8_147_625_0, i_8_147_632_0, i_8_147_666_0,
    i_8_147_679_0, i_8_147_683_0, i_8_147_696_0, i_8_147_697_0,
    i_8_147_705_0, i_8_147_725_0, i_8_147_757_0, i_8_147_773_0,
    i_8_147_778_0, i_8_147_781_0, i_8_147_783_0, i_8_147_786_0,
    i_8_147_787_0, i_8_147_790_0, i_8_147_812_0, i_8_147_826_0,
    i_8_147_829_0, i_8_147_838_0, i_8_147_841_0, i_8_147_842_0,
    i_8_147_847_0, i_8_147_848_0, i_8_147_869_0, i_8_147_874_0,
    i_8_147_917_0, i_8_147_932_0, i_8_147_1000_0, i_8_147_1057_0,
    i_8_147_1072_0, i_8_147_1135_0, i_8_147_1189_0, i_8_147_1234_0,
    i_8_147_1271_0, i_8_147_1328_0, i_8_147_1363_0, i_8_147_1369_0,
    i_8_147_1454_0, i_8_147_1457_0, i_8_147_1470_0, i_8_147_1524_0,
    i_8_147_1589_0, i_8_147_1607_0, i_8_147_1648_0, i_8_147_1655_0,
    i_8_147_1684_0, i_8_147_1696_0, i_8_147_1700_0, i_8_147_1729_0,
    i_8_147_1732_0, i_8_147_1749_0, i_8_147_1805_0, i_8_147_1846_0,
    i_8_147_1855_0, i_8_147_1856_0, i_8_147_1857_0, i_8_147_1858_0,
    i_8_147_1859_0, i_8_147_1861_0, i_8_147_1867_0, i_8_147_1888_0,
    i_8_147_1895_0, i_8_147_1898_0, i_8_147_1904_0, i_8_147_1981_0,
    i_8_147_2029_0, i_8_147_2072_0, i_8_147_2090_0, i_8_147_2174_0,
    i_8_147_2182_0, i_8_147_2183_0, i_8_147_2185_0, i_8_147_2191_0,
    i_8_147_2280_0, i_8_147_2290_0, i_8_147_2292_0, i_8_147_2294_0;
  output o_8_147_0_0;
  assign o_8_147_0_0 = 0;
endmodule



// Benchmark "kernel_8_148" written by ABC on Sun Jul 19 10:05:34 2020

module kernel_8_148 ( 
    i_8_148_9_0, i_8_148_70_0, i_8_148_118_0, i_8_148_123_0, i_8_148_127_0,
    i_8_148_164_0, i_8_148_180_0, i_8_148_218_0, i_8_148_228_0,
    i_8_148_236_0, i_8_148_271_0, i_8_148_313_0, i_8_148_352_0,
    i_8_148_378_0, i_8_148_388_0, i_8_148_425_0, i_8_148_433_0,
    i_8_148_438_0, i_8_148_531_0, i_8_148_551_0, i_8_148_553_0,
    i_8_148_567_0, i_8_148_603_0, i_8_148_621_0, i_8_148_649_0,
    i_8_148_698_0, i_8_148_804_0, i_8_148_831_0, i_8_148_832_0,
    i_8_148_837_0, i_8_148_848_0, i_8_148_878_0, i_8_148_885_0,
    i_8_148_921_0, i_8_148_930_0, i_8_148_981_0, i_8_148_982_0,
    i_8_148_984_0, i_8_148_985_0, i_8_148_990_0, i_8_148_994_0,
    i_8_148_999_0, i_8_148_1011_0, i_8_148_1012_0, i_8_148_1074_0,
    i_8_148_1089_0, i_8_148_1090_0, i_8_148_1128_0, i_8_148_1165_0,
    i_8_148_1183_0, i_8_148_1280_0, i_8_148_1291_0, i_8_148_1308_0,
    i_8_148_1317_0, i_8_148_1320_0, i_8_148_1387_0, i_8_148_1393_0,
    i_8_148_1401_0, i_8_148_1407_0, i_8_148_1424_0, i_8_148_1620_0,
    i_8_148_1621_0, i_8_148_1623_0, i_8_148_1641_0, i_8_148_1651_0,
    i_8_148_1654_0, i_8_148_1683_0, i_8_148_1686_0, i_8_148_1687_0,
    i_8_148_1728_0, i_8_148_1731_0, i_8_148_1734_0, i_8_148_1782_0,
    i_8_148_1794_0, i_8_148_1803_0, i_8_148_1829_0, i_8_148_1858_0,
    i_8_148_1864_0, i_8_148_1882_0, i_8_148_1884_0, i_8_148_1893_0,
    i_8_148_1896_0, i_8_148_1906_0, i_8_148_2055_0, i_8_148_2070_0,
    i_8_148_2073_0, i_8_148_2074_0, i_8_148_2083_0, i_8_148_2086_0,
    i_8_148_2092_0, i_8_148_2097_0, i_8_148_2148_0, i_8_148_2155_0,
    i_8_148_2215_0, i_8_148_2229_0, i_8_148_2232_0, i_8_148_2236_0,
    i_8_148_2247_0, i_8_148_2248_0, i_8_148_2258_0,
    o_8_148_0_0  );
  input  i_8_148_9_0, i_8_148_70_0, i_8_148_118_0, i_8_148_123_0,
    i_8_148_127_0, i_8_148_164_0, i_8_148_180_0, i_8_148_218_0,
    i_8_148_228_0, i_8_148_236_0, i_8_148_271_0, i_8_148_313_0,
    i_8_148_352_0, i_8_148_378_0, i_8_148_388_0, i_8_148_425_0,
    i_8_148_433_0, i_8_148_438_0, i_8_148_531_0, i_8_148_551_0,
    i_8_148_553_0, i_8_148_567_0, i_8_148_603_0, i_8_148_621_0,
    i_8_148_649_0, i_8_148_698_0, i_8_148_804_0, i_8_148_831_0,
    i_8_148_832_0, i_8_148_837_0, i_8_148_848_0, i_8_148_878_0,
    i_8_148_885_0, i_8_148_921_0, i_8_148_930_0, i_8_148_981_0,
    i_8_148_982_0, i_8_148_984_0, i_8_148_985_0, i_8_148_990_0,
    i_8_148_994_0, i_8_148_999_0, i_8_148_1011_0, i_8_148_1012_0,
    i_8_148_1074_0, i_8_148_1089_0, i_8_148_1090_0, i_8_148_1128_0,
    i_8_148_1165_0, i_8_148_1183_0, i_8_148_1280_0, i_8_148_1291_0,
    i_8_148_1308_0, i_8_148_1317_0, i_8_148_1320_0, i_8_148_1387_0,
    i_8_148_1393_0, i_8_148_1401_0, i_8_148_1407_0, i_8_148_1424_0,
    i_8_148_1620_0, i_8_148_1621_0, i_8_148_1623_0, i_8_148_1641_0,
    i_8_148_1651_0, i_8_148_1654_0, i_8_148_1683_0, i_8_148_1686_0,
    i_8_148_1687_0, i_8_148_1728_0, i_8_148_1731_0, i_8_148_1734_0,
    i_8_148_1782_0, i_8_148_1794_0, i_8_148_1803_0, i_8_148_1829_0,
    i_8_148_1858_0, i_8_148_1864_0, i_8_148_1882_0, i_8_148_1884_0,
    i_8_148_1893_0, i_8_148_1896_0, i_8_148_1906_0, i_8_148_2055_0,
    i_8_148_2070_0, i_8_148_2073_0, i_8_148_2074_0, i_8_148_2083_0,
    i_8_148_2086_0, i_8_148_2092_0, i_8_148_2097_0, i_8_148_2148_0,
    i_8_148_2155_0, i_8_148_2215_0, i_8_148_2229_0, i_8_148_2232_0,
    i_8_148_2236_0, i_8_148_2247_0, i_8_148_2248_0, i_8_148_2258_0;
  output o_8_148_0_0;
  assign o_8_148_0_0 = 0;
endmodule



// Benchmark "kernel_8_149" written by ABC on Sun Jul 19 10:05:35 2020

module kernel_8_149 ( 
    i_8_149_34_0, i_8_149_44_0, i_8_149_87_0, i_8_149_106_0, i_8_149_159_0,
    i_8_149_160_0, i_8_149_161_0, i_8_149_168_0, i_8_149_204_0,
    i_8_149_205_0, i_8_149_214_0, i_8_149_222_0, i_8_149_258_0,
    i_8_149_340_0, i_8_149_345_0, i_8_149_417_0, i_8_149_463_0,
    i_8_149_464_0, i_8_149_474_0, i_8_149_478_0, i_8_149_480_0,
    i_8_149_483_0, i_8_149_524_0, i_8_149_526_0, i_8_149_557_0,
    i_8_149_594_0, i_8_149_601_0, i_8_149_619_0, i_8_149_629_0,
    i_8_149_661_0, i_8_149_664_0, i_8_149_718_0, i_8_149_726_0,
    i_8_149_748_0, i_8_149_749_0, i_8_149_764_0, i_8_149_773_0,
    i_8_149_834_0, i_8_149_907_0, i_8_149_925_0, i_8_149_952_0,
    i_8_149_984_0, i_8_149_985_0, i_8_149_988_0, i_8_149_997_0,
    i_8_149_1069_0, i_8_149_1072_0, i_8_149_1086_0, i_8_149_1087_0,
    i_8_149_1114_0, i_8_149_1137_0, i_8_149_1148_0, i_8_149_1174_0,
    i_8_149_1193_0, i_8_149_1199_0, i_8_149_1219_0, i_8_149_1254_0,
    i_8_149_1302_0, i_8_149_1320_0, i_8_149_1338_0, i_8_149_1420_0,
    i_8_149_1423_0, i_8_149_1426_0, i_8_149_1434_0, i_8_149_1484_0,
    i_8_149_1528_0, i_8_149_1537_0, i_8_149_1544_0, i_8_149_1549_0,
    i_8_149_1582_0, i_8_149_1610_0, i_8_149_1614_0, i_8_149_1615_0,
    i_8_149_1617_0, i_8_149_1633_0, i_8_149_1666_0, i_8_149_1680_0,
    i_8_149_1734_0, i_8_149_1735_0, i_8_149_1751_0, i_8_149_1752_0,
    i_8_149_1761_0, i_8_149_1799_0, i_8_149_1836_0, i_8_149_1869_0,
    i_8_149_1932_0, i_8_149_2001_0, i_8_149_2002_0, i_8_149_2004_0,
    i_8_149_2013_0, i_8_149_2014_0, i_8_149_2049_0, i_8_149_2073_0,
    i_8_149_2094_0, i_8_149_2113_0, i_8_149_2156_0, i_8_149_2175_0,
    i_8_149_2182_0, i_8_149_2266_0, i_8_149_2293_0,
    o_8_149_0_0  );
  input  i_8_149_34_0, i_8_149_44_0, i_8_149_87_0, i_8_149_106_0,
    i_8_149_159_0, i_8_149_160_0, i_8_149_161_0, i_8_149_168_0,
    i_8_149_204_0, i_8_149_205_0, i_8_149_214_0, i_8_149_222_0,
    i_8_149_258_0, i_8_149_340_0, i_8_149_345_0, i_8_149_417_0,
    i_8_149_463_0, i_8_149_464_0, i_8_149_474_0, i_8_149_478_0,
    i_8_149_480_0, i_8_149_483_0, i_8_149_524_0, i_8_149_526_0,
    i_8_149_557_0, i_8_149_594_0, i_8_149_601_0, i_8_149_619_0,
    i_8_149_629_0, i_8_149_661_0, i_8_149_664_0, i_8_149_718_0,
    i_8_149_726_0, i_8_149_748_0, i_8_149_749_0, i_8_149_764_0,
    i_8_149_773_0, i_8_149_834_0, i_8_149_907_0, i_8_149_925_0,
    i_8_149_952_0, i_8_149_984_0, i_8_149_985_0, i_8_149_988_0,
    i_8_149_997_0, i_8_149_1069_0, i_8_149_1072_0, i_8_149_1086_0,
    i_8_149_1087_0, i_8_149_1114_0, i_8_149_1137_0, i_8_149_1148_0,
    i_8_149_1174_0, i_8_149_1193_0, i_8_149_1199_0, i_8_149_1219_0,
    i_8_149_1254_0, i_8_149_1302_0, i_8_149_1320_0, i_8_149_1338_0,
    i_8_149_1420_0, i_8_149_1423_0, i_8_149_1426_0, i_8_149_1434_0,
    i_8_149_1484_0, i_8_149_1528_0, i_8_149_1537_0, i_8_149_1544_0,
    i_8_149_1549_0, i_8_149_1582_0, i_8_149_1610_0, i_8_149_1614_0,
    i_8_149_1615_0, i_8_149_1617_0, i_8_149_1633_0, i_8_149_1666_0,
    i_8_149_1680_0, i_8_149_1734_0, i_8_149_1735_0, i_8_149_1751_0,
    i_8_149_1752_0, i_8_149_1761_0, i_8_149_1799_0, i_8_149_1836_0,
    i_8_149_1869_0, i_8_149_1932_0, i_8_149_2001_0, i_8_149_2002_0,
    i_8_149_2004_0, i_8_149_2013_0, i_8_149_2014_0, i_8_149_2049_0,
    i_8_149_2073_0, i_8_149_2094_0, i_8_149_2113_0, i_8_149_2156_0,
    i_8_149_2175_0, i_8_149_2182_0, i_8_149_2266_0, i_8_149_2293_0;
  output o_8_149_0_0;
  assign o_8_149_0_0 = 0;
endmodule



// Benchmark "kernel_8_150" written by ABC on Sun Jul 19 10:05:36 2020

module kernel_8_150 ( 
    i_8_150_147_0, i_8_150_190_0, i_8_150_194_0, i_8_150_228_0,
    i_8_150_229_0, i_8_150_283_0, i_8_150_310_0, i_8_150_318_0,
    i_8_150_346_0, i_8_150_361_0, i_8_150_379_0, i_8_150_418_0,
    i_8_150_450_0, i_8_150_452_0, i_8_150_490_0, i_8_150_571_0,
    i_8_150_598_0, i_8_150_628_0, i_8_150_652_0, i_8_150_658_0,
    i_8_150_693_0, i_8_150_694_0, i_8_150_695_0, i_8_150_700_0,
    i_8_150_705_0, i_8_150_748_0, i_8_150_751_0, i_8_150_778_0,
    i_8_150_838_0, i_8_150_839_0, i_8_150_841_0, i_8_150_874_0,
    i_8_150_876_0, i_8_150_877_0, i_8_150_878_0, i_8_150_966_0,
    i_8_150_967_0, i_8_150_990_0, i_8_150_991_0, i_8_150_1000_0,
    i_8_150_1002_0, i_8_150_1034_0, i_8_150_1036_0, i_8_150_1037_0,
    i_8_150_1039_0, i_8_150_1046_0, i_8_150_1075_0, i_8_150_1147_0,
    i_8_150_1164_0, i_8_150_1226_0, i_8_150_1234_0, i_8_150_1268_0,
    i_8_150_1270_0, i_8_150_1283_0, i_8_150_1354_0, i_8_150_1355_0,
    i_8_150_1399_0, i_8_150_1407_0, i_8_150_1411_0, i_8_150_1452_0,
    i_8_150_1507_0, i_8_150_1524_0, i_8_150_1539_0, i_8_150_1540_0,
    i_8_150_1542_0, i_8_150_1605_0, i_8_150_1621_0, i_8_150_1622_0,
    i_8_150_1625_0, i_8_150_1629_0, i_8_150_1641_0, i_8_150_1642_0,
    i_8_150_1703_0, i_8_150_1729_0, i_8_150_1732_0, i_8_150_1767_0,
    i_8_150_1777_0, i_8_150_1807_0, i_8_150_1821_0, i_8_150_1822_0,
    i_8_150_1894_0, i_8_150_1903_0, i_8_150_1904_0, i_8_150_1936_0,
    i_8_150_1984_0, i_8_150_1992_0, i_8_150_1996_0, i_8_150_2009_0,
    i_8_150_2011_0, i_8_150_2014_0, i_8_150_2055_0, i_8_150_2056_0,
    i_8_150_2082_0, i_8_150_2083_0, i_8_150_2147_0, i_8_150_2151_0,
    i_8_150_2155_0, i_8_150_2170_0, i_8_150_2225_0, i_8_150_2272_0,
    o_8_150_0_0  );
  input  i_8_150_147_0, i_8_150_190_0, i_8_150_194_0, i_8_150_228_0,
    i_8_150_229_0, i_8_150_283_0, i_8_150_310_0, i_8_150_318_0,
    i_8_150_346_0, i_8_150_361_0, i_8_150_379_0, i_8_150_418_0,
    i_8_150_450_0, i_8_150_452_0, i_8_150_490_0, i_8_150_571_0,
    i_8_150_598_0, i_8_150_628_0, i_8_150_652_0, i_8_150_658_0,
    i_8_150_693_0, i_8_150_694_0, i_8_150_695_0, i_8_150_700_0,
    i_8_150_705_0, i_8_150_748_0, i_8_150_751_0, i_8_150_778_0,
    i_8_150_838_0, i_8_150_839_0, i_8_150_841_0, i_8_150_874_0,
    i_8_150_876_0, i_8_150_877_0, i_8_150_878_0, i_8_150_966_0,
    i_8_150_967_0, i_8_150_990_0, i_8_150_991_0, i_8_150_1000_0,
    i_8_150_1002_0, i_8_150_1034_0, i_8_150_1036_0, i_8_150_1037_0,
    i_8_150_1039_0, i_8_150_1046_0, i_8_150_1075_0, i_8_150_1147_0,
    i_8_150_1164_0, i_8_150_1226_0, i_8_150_1234_0, i_8_150_1268_0,
    i_8_150_1270_0, i_8_150_1283_0, i_8_150_1354_0, i_8_150_1355_0,
    i_8_150_1399_0, i_8_150_1407_0, i_8_150_1411_0, i_8_150_1452_0,
    i_8_150_1507_0, i_8_150_1524_0, i_8_150_1539_0, i_8_150_1540_0,
    i_8_150_1542_0, i_8_150_1605_0, i_8_150_1621_0, i_8_150_1622_0,
    i_8_150_1625_0, i_8_150_1629_0, i_8_150_1641_0, i_8_150_1642_0,
    i_8_150_1703_0, i_8_150_1729_0, i_8_150_1732_0, i_8_150_1767_0,
    i_8_150_1777_0, i_8_150_1807_0, i_8_150_1821_0, i_8_150_1822_0,
    i_8_150_1894_0, i_8_150_1903_0, i_8_150_1904_0, i_8_150_1936_0,
    i_8_150_1984_0, i_8_150_1992_0, i_8_150_1996_0, i_8_150_2009_0,
    i_8_150_2011_0, i_8_150_2014_0, i_8_150_2055_0, i_8_150_2056_0,
    i_8_150_2082_0, i_8_150_2083_0, i_8_150_2147_0, i_8_150_2151_0,
    i_8_150_2155_0, i_8_150_2170_0, i_8_150_2225_0, i_8_150_2272_0;
  output o_8_150_0_0;
  assign o_8_150_0_0 = 0;
endmodule



// Benchmark "kernel_8_151" written by ABC on Sun Jul 19 10:05:37 2020

module kernel_8_151 ( 
    i_8_151_11_0, i_8_151_33_0, i_8_151_51_0, i_8_151_67_0, i_8_151_74_0,
    i_8_151_96_0, i_8_151_120_0, i_8_151_137_0, i_8_151_142_0,
    i_8_151_159_0, i_8_151_191_0, i_8_151_254_0, i_8_151_262_0,
    i_8_151_310_0, i_8_151_312_0, i_8_151_346_0, i_8_151_348_0,
    i_8_151_372_0, i_8_151_441_0, i_8_151_448_0, i_8_151_456_0,
    i_8_151_484_0, i_8_151_492_0, i_8_151_524_0, i_8_151_598_0,
    i_8_151_600_0, i_8_151_601_0, i_8_151_690_0, i_8_151_691_0,
    i_8_151_718_0, i_8_151_734_0, i_8_151_735_0, i_8_151_736_0,
    i_8_151_799_0, i_8_151_800_0, i_8_151_826_0, i_8_151_838_0,
    i_8_151_923_0, i_8_151_946_0, i_8_151_1014_0, i_8_151_1015_0,
    i_8_151_1026_0, i_8_151_1060_0, i_8_151_1077_0, i_8_151_1113_0,
    i_8_151_1119_0, i_8_151_1120_0, i_8_151_1188_0, i_8_151_1231_0,
    i_8_151_1258_0, i_8_151_1273_0, i_8_151_1300_0, i_8_151_1305_0,
    i_8_151_1306_0, i_8_151_1324_0, i_8_151_1348_0, i_8_151_1387_0,
    i_8_151_1418_0, i_8_151_1425_0, i_8_151_1506_0, i_8_151_1507_0,
    i_8_151_1525_0, i_8_151_1578_0, i_8_151_1581_0, i_8_151_1582_0,
    i_8_151_1587_0, i_8_151_1588_0, i_8_151_1623_0, i_8_151_1632_0,
    i_8_151_1647_0, i_8_151_1648_0, i_8_151_1677_0, i_8_151_1686_0,
    i_8_151_1699_0, i_8_151_1720_0, i_8_151_1721_0, i_8_151_1740_0,
    i_8_151_1742_0, i_8_151_1749_0, i_8_151_1786_0, i_8_151_1789_0,
    i_8_151_1791_0, i_8_151_1876_0, i_8_151_1905_0, i_8_151_1906_0,
    i_8_151_1907_0, i_8_151_2004_0, i_8_151_2031_0, i_8_151_2049_0,
    i_8_151_2050_0, i_8_151_2092_0, i_8_151_2143_0, i_8_151_2155_0,
    i_8_151_2156_0, i_8_151_2157_0, i_8_151_2158_0, i_8_151_2182_0,
    i_8_151_2214_0, i_8_151_2219_0, i_8_151_2262_0,
    o_8_151_0_0  );
  input  i_8_151_11_0, i_8_151_33_0, i_8_151_51_0, i_8_151_67_0,
    i_8_151_74_0, i_8_151_96_0, i_8_151_120_0, i_8_151_137_0,
    i_8_151_142_0, i_8_151_159_0, i_8_151_191_0, i_8_151_254_0,
    i_8_151_262_0, i_8_151_310_0, i_8_151_312_0, i_8_151_346_0,
    i_8_151_348_0, i_8_151_372_0, i_8_151_441_0, i_8_151_448_0,
    i_8_151_456_0, i_8_151_484_0, i_8_151_492_0, i_8_151_524_0,
    i_8_151_598_0, i_8_151_600_0, i_8_151_601_0, i_8_151_690_0,
    i_8_151_691_0, i_8_151_718_0, i_8_151_734_0, i_8_151_735_0,
    i_8_151_736_0, i_8_151_799_0, i_8_151_800_0, i_8_151_826_0,
    i_8_151_838_0, i_8_151_923_0, i_8_151_946_0, i_8_151_1014_0,
    i_8_151_1015_0, i_8_151_1026_0, i_8_151_1060_0, i_8_151_1077_0,
    i_8_151_1113_0, i_8_151_1119_0, i_8_151_1120_0, i_8_151_1188_0,
    i_8_151_1231_0, i_8_151_1258_0, i_8_151_1273_0, i_8_151_1300_0,
    i_8_151_1305_0, i_8_151_1306_0, i_8_151_1324_0, i_8_151_1348_0,
    i_8_151_1387_0, i_8_151_1418_0, i_8_151_1425_0, i_8_151_1506_0,
    i_8_151_1507_0, i_8_151_1525_0, i_8_151_1578_0, i_8_151_1581_0,
    i_8_151_1582_0, i_8_151_1587_0, i_8_151_1588_0, i_8_151_1623_0,
    i_8_151_1632_0, i_8_151_1647_0, i_8_151_1648_0, i_8_151_1677_0,
    i_8_151_1686_0, i_8_151_1699_0, i_8_151_1720_0, i_8_151_1721_0,
    i_8_151_1740_0, i_8_151_1742_0, i_8_151_1749_0, i_8_151_1786_0,
    i_8_151_1789_0, i_8_151_1791_0, i_8_151_1876_0, i_8_151_1905_0,
    i_8_151_1906_0, i_8_151_1907_0, i_8_151_2004_0, i_8_151_2031_0,
    i_8_151_2049_0, i_8_151_2050_0, i_8_151_2092_0, i_8_151_2143_0,
    i_8_151_2155_0, i_8_151_2156_0, i_8_151_2157_0, i_8_151_2158_0,
    i_8_151_2182_0, i_8_151_2214_0, i_8_151_2219_0, i_8_151_2262_0;
  output o_8_151_0_0;
  assign o_8_151_0_0 = 0;
endmodule



// Benchmark "kernel_8_152" written by ABC on Sun Jul 19 10:05:38 2020

module kernel_8_152 ( 
    i_8_152_4_0, i_8_152_57_0, i_8_152_86_0, i_8_152_95_0, i_8_152_97_0,
    i_8_152_157_0, i_8_152_181_0, i_8_152_184_0, i_8_152_185_0,
    i_8_152_224_0, i_8_152_227_0, i_8_152_233_0, i_8_152_374_0,
    i_8_152_388_0, i_8_152_417_0, i_8_152_436_0, i_8_152_437_0,
    i_8_152_454_0, i_8_152_459_0, i_8_152_462_0, i_8_152_475_0,
    i_8_152_485_0, i_8_152_499_0, i_8_152_505_0, i_8_152_550_0,
    i_8_152_595_0, i_8_152_599_0, i_8_152_610_0, i_8_152_621_0,
    i_8_152_625_0, i_8_152_670_0, i_8_152_671_0, i_8_152_696_0,
    i_8_152_713_0, i_8_152_716_0, i_8_152_758_0, i_8_152_766_0,
    i_8_152_775_0, i_8_152_793_0, i_8_152_820_0, i_8_152_824_0,
    i_8_152_866_0, i_8_152_923_0, i_8_152_1009_0, i_8_152_1031_0,
    i_8_152_1081_0, i_8_152_1118_0, i_8_152_1180_0, i_8_152_1188_0,
    i_8_152_1204_0, i_8_152_1235_0, i_8_152_1255_0, i_8_152_1261_0,
    i_8_152_1269_0, i_8_152_1270_0, i_8_152_1280_0, i_8_152_1282_0,
    i_8_152_1283_0, i_8_152_1298_0, i_8_152_1308_0, i_8_152_1342_0,
    i_8_152_1346_0, i_8_152_1436_0, i_8_152_1450_0, i_8_152_1467_0,
    i_8_152_1469_0, i_8_152_1492_0, i_8_152_1503_0, i_8_152_1504_0,
    i_8_152_1539_0, i_8_152_1571_0, i_8_152_1597_0, i_8_152_1622_0,
    i_8_152_1679_0, i_8_152_1681_0, i_8_152_1746_0, i_8_152_1751_0,
    i_8_152_1752_0, i_8_152_1753_0, i_8_152_1781_0, i_8_152_1787_0,
    i_8_152_1789_0, i_8_152_1800_0, i_8_152_1805_0, i_8_152_1817_0,
    i_8_152_1855_0, i_8_152_1918_0, i_8_152_1948_0, i_8_152_1963_0,
    i_8_152_1966_0, i_8_152_2108_0, i_8_152_2109_0, i_8_152_2110_0,
    i_8_152_2139_0, i_8_152_2147_0, i_8_152_2244_0, i_8_152_2270_0,
    i_8_152_2272_0, i_8_152_2286_0, i_8_152_2290_0,
    o_8_152_0_0  );
  input  i_8_152_4_0, i_8_152_57_0, i_8_152_86_0, i_8_152_95_0,
    i_8_152_97_0, i_8_152_157_0, i_8_152_181_0, i_8_152_184_0,
    i_8_152_185_0, i_8_152_224_0, i_8_152_227_0, i_8_152_233_0,
    i_8_152_374_0, i_8_152_388_0, i_8_152_417_0, i_8_152_436_0,
    i_8_152_437_0, i_8_152_454_0, i_8_152_459_0, i_8_152_462_0,
    i_8_152_475_0, i_8_152_485_0, i_8_152_499_0, i_8_152_505_0,
    i_8_152_550_0, i_8_152_595_0, i_8_152_599_0, i_8_152_610_0,
    i_8_152_621_0, i_8_152_625_0, i_8_152_670_0, i_8_152_671_0,
    i_8_152_696_0, i_8_152_713_0, i_8_152_716_0, i_8_152_758_0,
    i_8_152_766_0, i_8_152_775_0, i_8_152_793_0, i_8_152_820_0,
    i_8_152_824_0, i_8_152_866_0, i_8_152_923_0, i_8_152_1009_0,
    i_8_152_1031_0, i_8_152_1081_0, i_8_152_1118_0, i_8_152_1180_0,
    i_8_152_1188_0, i_8_152_1204_0, i_8_152_1235_0, i_8_152_1255_0,
    i_8_152_1261_0, i_8_152_1269_0, i_8_152_1270_0, i_8_152_1280_0,
    i_8_152_1282_0, i_8_152_1283_0, i_8_152_1298_0, i_8_152_1308_0,
    i_8_152_1342_0, i_8_152_1346_0, i_8_152_1436_0, i_8_152_1450_0,
    i_8_152_1467_0, i_8_152_1469_0, i_8_152_1492_0, i_8_152_1503_0,
    i_8_152_1504_0, i_8_152_1539_0, i_8_152_1571_0, i_8_152_1597_0,
    i_8_152_1622_0, i_8_152_1679_0, i_8_152_1681_0, i_8_152_1746_0,
    i_8_152_1751_0, i_8_152_1752_0, i_8_152_1753_0, i_8_152_1781_0,
    i_8_152_1787_0, i_8_152_1789_0, i_8_152_1800_0, i_8_152_1805_0,
    i_8_152_1817_0, i_8_152_1855_0, i_8_152_1918_0, i_8_152_1948_0,
    i_8_152_1963_0, i_8_152_1966_0, i_8_152_2108_0, i_8_152_2109_0,
    i_8_152_2110_0, i_8_152_2139_0, i_8_152_2147_0, i_8_152_2244_0,
    i_8_152_2270_0, i_8_152_2272_0, i_8_152_2286_0, i_8_152_2290_0;
  output o_8_152_0_0;
  assign o_8_152_0_0 = 0;
endmodule



// Benchmark "kernel_8_153" written by ABC on Sun Jul 19 10:05:40 2020

module kernel_8_153 ( 
    i_8_153_51_0, i_8_153_53_0, i_8_153_124_0, i_8_153_125_0,
    i_8_153_168_0, i_8_153_169_0, i_8_153_170_0, i_8_153_172_0,
    i_8_153_177_0, i_8_153_330_0, i_8_153_341_0, i_8_153_348_0,
    i_8_153_368_0, i_8_153_378_0, i_8_153_379_0, i_8_153_384_0,
    i_8_153_393_0, i_8_153_418_0, i_8_153_420_0, i_8_153_422_0,
    i_8_153_469_0, i_8_153_499_0, i_8_153_598_0, i_8_153_659_0,
    i_8_153_704_0, i_8_153_753_0, i_8_153_778_0, i_8_153_879_0,
    i_8_153_898_0, i_8_153_985_0, i_8_153_987_0, i_8_153_988_0,
    i_8_153_994_0, i_8_153_1015_0, i_8_153_1040_0, i_8_153_1051_0,
    i_8_153_1111_0, i_8_153_1131_0, i_8_153_1132_0, i_8_153_1139_0,
    i_8_153_1140_0, i_8_153_1141_0, i_8_153_1168_0, i_8_153_1228_0,
    i_8_153_1236_0, i_8_153_1237_0, i_8_153_1261_0, i_8_153_1263_0,
    i_8_153_1275_0, i_8_153_1276_0, i_8_153_1277_0, i_8_153_1281_0,
    i_8_153_1284_0, i_8_153_1285_0, i_8_153_1286_0, i_8_153_1331_0,
    i_8_153_1381_0, i_8_153_1434_0, i_8_153_1446_0, i_8_153_1470_0,
    i_8_153_1471_0, i_8_153_1474_0, i_8_153_1475_0, i_8_153_1479_0,
    i_8_153_1482_0, i_8_153_1484_0, i_8_153_1511_0, i_8_153_1520_0,
    i_8_153_1527_0, i_8_153_1529_0, i_8_153_1536_0, i_8_153_1554_0,
    i_8_153_1588_0, i_8_153_1590_0, i_8_153_1635_0, i_8_153_1645_0,
    i_8_153_1654_0, i_8_153_1664_0, i_8_153_1671_0, i_8_153_1672_0,
    i_8_153_1734_0, i_8_153_1735_0, i_8_153_1762_0, i_8_153_1770_0,
    i_8_153_1783_0, i_8_153_1808_0, i_8_153_1862_0, i_8_153_1870_0,
    i_8_153_1969_0, i_8_153_1992_0, i_8_153_1993_0, i_8_153_2013_0,
    i_8_153_2015_0, i_8_153_2038_0, i_8_153_2048_0, i_8_153_2095_0,
    i_8_153_2122_0, i_8_153_2146_0, i_8_153_2147_0, i_8_153_2276_0,
    o_8_153_0_0  );
  input  i_8_153_51_0, i_8_153_53_0, i_8_153_124_0, i_8_153_125_0,
    i_8_153_168_0, i_8_153_169_0, i_8_153_170_0, i_8_153_172_0,
    i_8_153_177_0, i_8_153_330_0, i_8_153_341_0, i_8_153_348_0,
    i_8_153_368_0, i_8_153_378_0, i_8_153_379_0, i_8_153_384_0,
    i_8_153_393_0, i_8_153_418_0, i_8_153_420_0, i_8_153_422_0,
    i_8_153_469_0, i_8_153_499_0, i_8_153_598_0, i_8_153_659_0,
    i_8_153_704_0, i_8_153_753_0, i_8_153_778_0, i_8_153_879_0,
    i_8_153_898_0, i_8_153_985_0, i_8_153_987_0, i_8_153_988_0,
    i_8_153_994_0, i_8_153_1015_0, i_8_153_1040_0, i_8_153_1051_0,
    i_8_153_1111_0, i_8_153_1131_0, i_8_153_1132_0, i_8_153_1139_0,
    i_8_153_1140_0, i_8_153_1141_0, i_8_153_1168_0, i_8_153_1228_0,
    i_8_153_1236_0, i_8_153_1237_0, i_8_153_1261_0, i_8_153_1263_0,
    i_8_153_1275_0, i_8_153_1276_0, i_8_153_1277_0, i_8_153_1281_0,
    i_8_153_1284_0, i_8_153_1285_0, i_8_153_1286_0, i_8_153_1331_0,
    i_8_153_1381_0, i_8_153_1434_0, i_8_153_1446_0, i_8_153_1470_0,
    i_8_153_1471_0, i_8_153_1474_0, i_8_153_1475_0, i_8_153_1479_0,
    i_8_153_1482_0, i_8_153_1484_0, i_8_153_1511_0, i_8_153_1520_0,
    i_8_153_1527_0, i_8_153_1529_0, i_8_153_1536_0, i_8_153_1554_0,
    i_8_153_1588_0, i_8_153_1590_0, i_8_153_1635_0, i_8_153_1645_0,
    i_8_153_1654_0, i_8_153_1664_0, i_8_153_1671_0, i_8_153_1672_0,
    i_8_153_1734_0, i_8_153_1735_0, i_8_153_1762_0, i_8_153_1770_0,
    i_8_153_1783_0, i_8_153_1808_0, i_8_153_1862_0, i_8_153_1870_0,
    i_8_153_1969_0, i_8_153_1992_0, i_8_153_1993_0, i_8_153_2013_0,
    i_8_153_2015_0, i_8_153_2038_0, i_8_153_2048_0, i_8_153_2095_0,
    i_8_153_2122_0, i_8_153_2146_0, i_8_153_2147_0, i_8_153_2276_0;
  output o_8_153_0_0;
  assign o_8_153_0_0 = ~((~i_8_153_1529_0 & ((~i_8_153_1479_0 & ((~i_8_153_2013_0 & ((~i_8_153_1664_0 & ((~i_8_153_341_0 & ((~i_8_153_418_0 & ~i_8_153_1237_0 & ~i_8_153_1277_0 & i_8_153_1281_0 & ~i_8_153_1446_0 & ~i_8_153_1470_0 & ~i_8_153_1734_0) | (~i_8_153_378_0 & ~i_8_153_379_0 & ~i_8_153_420_0 & ~i_8_153_469_0 & ~i_8_153_987_0 & ~i_8_153_1139_0 & ~i_8_153_1520_0 & ~i_8_153_2015_0 & ~i_8_153_2095_0))) | (i_8_153_879_0 & ~i_8_153_994_0 & ~i_8_153_1446_0 & i_8_153_1862_0 & ~i_8_153_1969_0 & ~i_8_153_2122_0))) | (~i_8_153_378_0 & ~i_8_153_420_0 & ~i_8_153_988_0 & ~i_8_153_994_0 & ~i_8_153_1132_0 & ~i_8_153_1277_0 & ~i_8_153_1520_0 & ~i_8_153_1536_0 & ~i_8_153_1654_0 & ~i_8_153_1783_0 & ~i_8_153_1862_0 & ~i_8_153_2015_0 & ~i_8_153_2276_0))) | (~i_8_153_125_0 & ~i_8_153_378_0 & ~i_8_153_422_0 & ~i_8_153_985_0 & ~i_8_153_988_0 & ~i_8_153_1132_0 & ~i_8_153_1139_0 & ~i_8_153_1520_0 & ~i_8_153_1635_0 & ~i_8_153_1770_0))) | (~i_8_153_1139_0 & ((~i_8_153_985_0 & ~i_8_153_1672_0 & ((~i_8_153_125_0 & ~i_8_153_1140_0 & ~i_8_153_1527_0 & ((~i_8_153_379_0 & i_8_153_469_0 & ~i_8_153_988_0 & ~i_8_153_1141_0 & ~i_8_153_1664_0) | (~i_8_153_378_0 & ~i_8_153_422_0 & ~i_8_153_1484_0 & ~i_8_153_1671_0 & ~i_8_153_1770_0 & ~i_8_153_1992_0 & ~i_8_153_1993_0))) | (~i_8_153_378_0 & ~i_8_153_1132_0 & ~i_8_153_1520_0 & ~i_8_153_1554_0 & ~i_8_153_1645_0 & ~i_8_153_1862_0 & ~i_8_153_2013_0 & ~i_8_153_2015_0))) | (~i_8_153_393_0 & ((~i_8_153_125_0 & ~i_8_153_987_0 & ~i_8_153_1131_0 & i_8_153_1993_0 & ~i_8_153_2015_0) | (~i_8_153_379_0 & ~i_8_153_422_0 & ~i_8_153_879_0 & ~i_8_153_1040_0 & ~i_8_153_1168_0 & ~i_8_153_1284_0 & ~i_8_153_1484_0 & ~i_8_153_1635_0 & ~i_8_153_1969_0 & ~i_8_153_2146_0))) | (~i_8_153_418_0 & ~i_8_153_659_0 & i_8_153_1040_0 & ~i_8_153_1671_0 & i_8_153_1969_0 & ~i_8_153_2276_0))) | (~i_8_153_125_0 & ((~i_8_153_994_0 & ~i_8_153_1040_0 & ~i_8_153_1168_0 & i_8_153_1434_0 & ~i_8_153_1482_0) | (~i_8_153_898_0 & ~i_8_153_1051_0 & ~i_8_153_1261_0 & i_8_153_1277_0 & ~i_8_153_1862_0))) | (~i_8_153_1482_0 & ((~i_8_153_1140_0 & i_8_153_1470_0 & ~i_8_153_1664_0) | (i_8_153_778_0 & ~i_8_153_1168_0 & ~i_8_153_1520_0 & ~i_8_153_1536_0 & ~i_8_153_1808_0 & ~i_8_153_2095_0))) | (~i_8_153_987_0 & ~i_8_153_1040_0 & ~i_8_153_1141_0 & i_8_153_1381_0) | (~i_8_153_704_0 & ~i_8_153_1111_0 & ~i_8_153_1277_0 & i_8_153_1331_0 & i_8_153_1808_0))) | (~i_8_153_125_0 & ((~i_8_153_1015_0 & ~i_8_153_1132_0 & ~i_8_153_1141_0 & ~i_8_153_1168_0 & i_8_153_1237_0 & ~i_8_153_1482_0) | (~i_8_153_330_0 & ~i_8_153_987_0 & ~i_8_153_1275_0 & i_8_153_1475_0 & ~i_8_153_1511_0))) | (~i_8_153_378_0 & ((~i_8_153_124_0 & ~i_8_153_379_0 & i_8_153_659_0 & ~i_8_153_879_0 & ~i_8_153_1511_0 & ~i_8_153_1734_0) | (i_8_153_53_0 & ~i_8_153_1168_0 & ~i_8_153_2015_0))) | (i_8_153_598_0 & ((~i_8_153_985_0 & i_8_153_1111_0 & ~i_8_153_1286_0 & ~i_8_153_1527_0 & ~i_8_153_1862_0) | (~i_8_153_469_0 & i_8_153_1131_0 & ~i_8_153_1228_0 & i_8_153_1434_0 & ~i_8_153_1511_0 & ~i_8_153_2095_0))) | (~i_8_153_469_0 & ~i_8_153_2013_0 & ((~i_8_153_598_0 & ~i_8_153_1475_0 & ~i_8_153_1664_0 & ~i_8_153_1671_0 & ~i_8_153_1993_0 & i_8_153_2048_0) | (~i_8_153_330_0 & ~i_8_153_341_0 & ~i_8_153_1111_0 & ~i_8_153_1168_0 & ~i_8_153_1520_0 & i_8_153_2146_0 & ~i_8_153_2276_0))) | (~i_8_153_330_0 & ((i_8_153_469_0 & i_8_153_1261_0 & ~i_8_153_1554_0 & ~i_8_153_1808_0 & ~i_8_153_1969_0) | (~i_8_153_985_0 & ~i_8_153_988_0 & ~i_8_153_1168_0 & ~i_8_153_1285_0 & ~i_8_153_1511_0 & ~i_8_153_1527_0 & ~i_8_153_1664_0 & i_8_153_2147_0))) | (i_8_153_704_0 & ((~i_8_153_985_0 & ~i_8_153_1040_0 & ~i_8_153_1484_0 & ~i_8_153_1520_0 & ~i_8_153_1735_0 & i_8_153_1862_0) | (~i_8_153_422_0 & ~i_8_153_1511_0 & ~i_8_153_1862_0 & ~i_8_153_2095_0))) | (~i_8_153_422_0 & ((~i_8_153_379_0 & i_8_153_1263_0 & ~i_8_153_1554_0) | (~i_8_153_985_0 & i_8_153_1286_0 & i_8_153_1969_0))) | (~i_8_153_994_0 & ((~i_8_153_1111_0 & i_8_153_1434_0 & ~i_8_153_1770_0 & i_8_153_1783_0) | (~i_8_153_598_0 & ~i_8_153_1168_0 & ~i_8_153_1520_0 & ~i_8_153_1527_0 & ~i_8_153_1672_0 & ~i_8_153_1734_0 & i_8_153_1992_0 & ~i_8_153_2276_0))) | (~i_8_153_1168_0 & ((~i_8_153_124_0 & ~i_8_153_341_0 & ~i_8_153_987_0 & i_8_153_1236_0 & i_8_153_1482_0 & ~i_8_153_1770_0) | (i_8_153_379_0 & i_8_153_659_0 & ~i_8_153_1139_0 & ~i_8_153_1783_0 & ~i_8_153_1808_0))) | (~i_8_153_341_0 & ((~i_8_153_124_0 & ~i_8_153_177_0 & ~i_8_153_1139_0 & i_8_153_1474_0 & ~i_8_153_1664_0 & ~i_8_153_1672_0 & ~i_8_153_1783_0) | (i_8_153_499_0 & ~i_8_153_987_0 & ~i_8_153_1479_0 & ~i_8_153_1635_0 & ~i_8_153_2146_0))) | (~i_8_153_124_0 & ((~i_8_153_987_0 & ~i_8_153_1131_0 & i_8_153_1284_0 & ~i_8_153_1511_0 & ~i_8_153_1635_0 & ~i_8_153_1664_0 & ~i_8_153_1783_0) | (i_8_153_1111_0 & ~i_8_153_1139_0 & ~i_8_153_1263_0 & ~i_8_153_1277_0 & ~i_8_153_1434_0 & ~i_8_153_1479_0 & ~i_8_153_1588_0 & ~i_8_153_1770_0 & ~i_8_153_1808_0))) | (~i_8_153_1527_0 & ~i_8_153_1862_0 & ((i_8_153_1263_0 & i_8_153_1434_0 & ~i_8_153_1484_0) | (i_8_153_1236_0 & ~i_8_153_1482_0 & ~i_8_153_1635_0 & ~i_8_153_1672_0))) | (~i_8_153_1484_0 & ((~i_8_153_987_0 & ~i_8_153_1040_0 & i_8_153_1277_0 & ~i_8_153_1554_0) | (~i_8_153_420_0 & ~i_8_153_898_0 & i_8_153_1590_0) | (~i_8_153_1051_0 & ~i_8_153_1139_0 & ~i_8_153_1762_0 & ~i_8_153_1969_0 & i_8_153_2147_0))) | (i_8_153_348_0 & i_8_153_418_0 & i_8_153_1635_0 & ~i_8_153_1671_0) | (i_8_153_1285_0 & i_8_153_1286_0 & ~i_8_153_1446_0 & ~i_8_153_1511_0 & ~i_8_153_2015_0));
endmodule



// Benchmark "kernel_8_154" written by ABC on Sun Jul 19 10:05:40 2020

module kernel_8_154 ( 
    i_8_154_28_0, i_8_154_47_0, i_8_154_64_0, i_8_154_72_0, i_8_154_77_0,
    i_8_154_111_0, i_8_154_181_0, i_8_154_226_0, i_8_154_308_0,
    i_8_154_319_0, i_8_154_320_0, i_8_154_388_0, i_8_154_398_0,
    i_8_154_506_0, i_8_154_536_0, i_8_154_551_0, i_8_154_559_0,
    i_8_154_571_0, i_8_154_572_0, i_8_154_578_0, i_8_154_579_0,
    i_8_154_586_0, i_8_154_587_0, i_8_154_596_0, i_8_154_603_0,
    i_8_154_611_0, i_8_154_630_0, i_8_154_631_0, i_8_154_634_0,
    i_8_154_640_0, i_8_154_649_0, i_8_154_652_0, i_8_154_659_0,
    i_8_154_680_0, i_8_154_707_0, i_8_154_748_0, i_8_154_793_0,
    i_8_154_794_0, i_8_154_837_0, i_8_154_844_0, i_8_154_845_0,
    i_8_154_855_0, i_8_154_859_0, i_8_154_874_0, i_8_154_882_0,
    i_8_154_969_0, i_8_154_973_0, i_8_154_991_0, i_8_154_1073_0,
    i_8_154_1108_0, i_8_154_1128_0, i_8_154_1143_0, i_8_154_1170_0,
    i_8_154_1180_0, i_8_154_1199_0, i_8_154_1226_0, i_8_154_1243_0,
    i_8_154_1261_0, i_8_154_1264_0, i_8_154_1328_0, i_8_154_1405_0,
    i_8_154_1410_0, i_8_154_1459_0, i_8_154_1462_0, i_8_154_1469_0,
    i_8_154_1472_0, i_8_154_1478_0, i_8_154_1523_0, i_8_154_1536_0,
    i_8_154_1544_0, i_8_154_1625_0, i_8_154_1648_0, i_8_154_1650_0,
    i_8_154_1651_0, i_8_154_1682_0, i_8_154_1684_0, i_8_154_1694_0,
    i_8_154_1703_0, i_8_154_1748_0, i_8_154_1765_0, i_8_154_1777_0,
    i_8_154_1781_0, i_8_154_1782_0, i_8_154_1819_0, i_8_154_1820_0,
    i_8_154_1822_0, i_8_154_1823_0, i_8_154_1855_0, i_8_154_1881_0,
    i_8_154_1909_0, i_8_154_1936_0, i_8_154_1954_0, i_8_154_1994_0,
    i_8_154_2146_0, i_8_154_2147_0, i_8_154_2170_0, i_8_154_2191_0,
    i_8_154_2207_0, i_8_154_2225_0, i_8_154_2241_0,
    o_8_154_0_0  );
  input  i_8_154_28_0, i_8_154_47_0, i_8_154_64_0, i_8_154_72_0,
    i_8_154_77_0, i_8_154_111_0, i_8_154_181_0, i_8_154_226_0,
    i_8_154_308_0, i_8_154_319_0, i_8_154_320_0, i_8_154_388_0,
    i_8_154_398_0, i_8_154_506_0, i_8_154_536_0, i_8_154_551_0,
    i_8_154_559_0, i_8_154_571_0, i_8_154_572_0, i_8_154_578_0,
    i_8_154_579_0, i_8_154_586_0, i_8_154_587_0, i_8_154_596_0,
    i_8_154_603_0, i_8_154_611_0, i_8_154_630_0, i_8_154_631_0,
    i_8_154_634_0, i_8_154_640_0, i_8_154_649_0, i_8_154_652_0,
    i_8_154_659_0, i_8_154_680_0, i_8_154_707_0, i_8_154_748_0,
    i_8_154_793_0, i_8_154_794_0, i_8_154_837_0, i_8_154_844_0,
    i_8_154_845_0, i_8_154_855_0, i_8_154_859_0, i_8_154_874_0,
    i_8_154_882_0, i_8_154_969_0, i_8_154_973_0, i_8_154_991_0,
    i_8_154_1073_0, i_8_154_1108_0, i_8_154_1128_0, i_8_154_1143_0,
    i_8_154_1170_0, i_8_154_1180_0, i_8_154_1199_0, i_8_154_1226_0,
    i_8_154_1243_0, i_8_154_1261_0, i_8_154_1264_0, i_8_154_1328_0,
    i_8_154_1405_0, i_8_154_1410_0, i_8_154_1459_0, i_8_154_1462_0,
    i_8_154_1469_0, i_8_154_1472_0, i_8_154_1478_0, i_8_154_1523_0,
    i_8_154_1536_0, i_8_154_1544_0, i_8_154_1625_0, i_8_154_1648_0,
    i_8_154_1650_0, i_8_154_1651_0, i_8_154_1682_0, i_8_154_1684_0,
    i_8_154_1694_0, i_8_154_1703_0, i_8_154_1748_0, i_8_154_1765_0,
    i_8_154_1777_0, i_8_154_1781_0, i_8_154_1782_0, i_8_154_1819_0,
    i_8_154_1820_0, i_8_154_1822_0, i_8_154_1823_0, i_8_154_1855_0,
    i_8_154_1881_0, i_8_154_1909_0, i_8_154_1936_0, i_8_154_1954_0,
    i_8_154_1994_0, i_8_154_2146_0, i_8_154_2147_0, i_8_154_2170_0,
    i_8_154_2191_0, i_8_154_2207_0, i_8_154_2225_0, i_8_154_2241_0;
  output o_8_154_0_0;
  assign o_8_154_0_0 = 0;
endmodule



// Benchmark "kernel_8_155" written by ABC on Sun Jul 19 10:05:41 2020

module kernel_8_155 ( 
    i_8_155_6_0, i_8_155_32_0, i_8_155_43_0, i_8_155_49_0, i_8_155_50_0,
    i_8_155_64_0, i_8_155_67_0, i_8_155_75_0, i_8_155_142_0, i_8_155_151_0,
    i_8_155_169_0, i_8_155_215_0, i_8_155_260_0, i_8_155_337_0,
    i_8_155_338_0, i_8_155_347_0, i_8_155_355_0, i_8_155_363_0,
    i_8_155_385_0, i_8_155_386_0, i_8_155_416_0, i_8_155_427_0,
    i_8_155_453_0, i_8_155_500_0, i_8_155_523_0, i_8_155_527_0,
    i_8_155_538_0, i_8_155_593_0, i_8_155_608_0, i_8_155_613_0,
    i_8_155_614_0, i_8_155_633_0, i_8_155_634_0, i_8_155_664_0,
    i_8_155_703_0, i_8_155_704_0, i_8_155_705_0, i_8_155_706_0,
    i_8_155_763_0, i_8_155_770_0, i_8_155_955_0, i_8_155_958_0,
    i_8_155_964_0, i_8_155_994_0, i_8_155_995_0, i_8_155_1078_0,
    i_8_155_1110_0, i_8_155_1125_0, i_8_155_1139_0, i_8_155_1154_0,
    i_8_155_1174_0, i_8_155_1175_0, i_8_155_1227_0, i_8_155_1228_0,
    i_8_155_1262_0, i_8_155_1299_0, i_8_155_1410_0, i_8_155_1417_0,
    i_8_155_1438_0, i_8_155_1453_0, i_8_155_1456_0, i_8_155_1475_0,
    i_8_155_1525_0, i_8_155_1531_0, i_8_155_1556_0, i_8_155_1600_0,
    i_8_155_1624_0, i_8_155_1648_0, i_8_155_1679_0, i_8_155_1682_0,
    i_8_155_1733_0, i_8_155_1785_0, i_8_155_1818_0, i_8_155_1819_0,
    i_8_155_1821_0, i_8_155_1824_0, i_8_155_1866_0, i_8_155_1877_0,
    i_8_155_1957_0, i_8_155_1967_0, i_8_155_1975_0, i_8_155_1995_0,
    i_8_155_2005_0, i_8_155_2013_0, i_8_155_2048_0, i_8_155_2057_0,
    i_8_155_2065_0, i_8_155_2094_0, i_8_155_2095_0, i_8_155_2143_0,
    i_8_155_2147_0, i_8_155_2148_0, i_8_155_2150_0, i_8_155_2157_0,
    i_8_155_2159_0, i_8_155_2171_0, i_8_155_2183_0, i_8_155_2226_0,
    i_8_155_2231_0, i_8_155_2266_0,
    o_8_155_0_0  );
  input  i_8_155_6_0, i_8_155_32_0, i_8_155_43_0, i_8_155_49_0,
    i_8_155_50_0, i_8_155_64_0, i_8_155_67_0, i_8_155_75_0, i_8_155_142_0,
    i_8_155_151_0, i_8_155_169_0, i_8_155_215_0, i_8_155_260_0,
    i_8_155_337_0, i_8_155_338_0, i_8_155_347_0, i_8_155_355_0,
    i_8_155_363_0, i_8_155_385_0, i_8_155_386_0, i_8_155_416_0,
    i_8_155_427_0, i_8_155_453_0, i_8_155_500_0, i_8_155_523_0,
    i_8_155_527_0, i_8_155_538_0, i_8_155_593_0, i_8_155_608_0,
    i_8_155_613_0, i_8_155_614_0, i_8_155_633_0, i_8_155_634_0,
    i_8_155_664_0, i_8_155_703_0, i_8_155_704_0, i_8_155_705_0,
    i_8_155_706_0, i_8_155_763_0, i_8_155_770_0, i_8_155_955_0,
    i_8_155_958_0, i_8_155_964_0, i_8_155_994_0, i_8_155_995_0,
    i_8_155_1078_0, i_8_155_1110_0, i_8_155_1125_0, i_8_155_1139_0,
    i_8_155_1154_0, i_8_155_1174_0, i_8_155_1175_0, i_8_155_1227_0,
    i_8_155_1228_0, i_8_155_1262_0, i_8_155_1299_0, i_8_155_1410_0,
    i_8_155_1417_0, i_8_155_1438_0, i_8_155_1453_0, i_8_155_1456_0,
    i_8_155_1475_0, i_8_155_1525_0, i_8_155_1531_0, i_8_155_1556_0,
    i_8_155_1600_0, i_8_155_1624_0, i_8_155_1648_0, i_8_155_1679_0,
    i_8_155_1682_0, i_8_155_1733_0, i_8_155_1785_0, i_8_155_1818_0,
    i_8_155_1819_0, i_8_155_1821_0, i_8_155_1824_0, i_8_155_1866_0,
    i_8_155_1877_0, i_8_155_1957_0, i_8_155_1967_0, i_8_155_1975_0,
    i_8_155_1995_0, i_8_155_2005_0, i_8_155_2013_0, i_8_155_2048_0,
    i_8_155_2057_0, i_8_155_2065_0, i_8_155_2094_0, i_8_155_2095_0,
    i_8_155_2143_0, i_8_155_2147_0, i_8_155_2148_0, i_8_155_2150_0,
    i_8_155_2157_0, i_8_155_2159_0, i_8_155_2171_0, i_8_155_2183_0,
    i_8_155_2226_0, i_8_155_2231_0, i_8_155_2266_0;
  output o_8_155_0_0;
  assign o_8_155_0_0 = 0;
endmodule



// Benchmark "kernel_8_156" written by ABC on Sun Jul 19 10:05:43 2020

module kernel_8_156 ( 
    i_8_156_35_0, i_8_156_37_0, i_8_156_77_0, i_8_156_87_0, i_8_156_111_0,
    i_8_156_140_0, i_8_156_229_0, i_8_156_235_0, i_8_156_259_0,
    i_8_156_304_0, i_8_156_355_0, i_8_156_382_0, i_8_156_418_0,
    i_8_156_419_0, i_8_156_442_0, i_8_156_445_0, i_8_156_446_0,
    i_8_156_464_0, i_8_156_490_0, i_8_156_504_0, i_8_156_505_0,
    i_8_156_506_0, i_8_156_507_0, i_8_156_508_0, i_8_156_509_0,
    i_8_156_528_0, i_8_156_610_0, i_8_156_621_0, i_8_156_625_0,
    i_8_156_665_0, i_8_156_698_0, i_8_156_748_0, i_8_156_780_0,
    i_8_156_781_0, i_8_156_845_0, i_8_156_876_0, i_8_156_880_0,
    i_8_156_885_0, i_8_156_967_0, i_8_156_1028_0, i_8_156_1030_0,
    i_8_156_1031_0, i_8_156_1136_0, i_8_156_1158_0, i_8_156_1192_0,
    i_8_156_1200_0, i_8_156_1201_0, i_8_156_1202_0, i_8_156_1225_0,
    i_8_156_1269_0, i_8_156_1281_0, i_8_156_1315_0, i_8_156_1325_0,
    i_8_156_1328_0, i_8_156_1350_0, i_8_156_1355_0, i_8_156_1387_0,
    i_8_156_1398_0, i_8_156_1399_0, i_8_156_1400_0, i_8_156_1437_0,
    i_8_156_1450_0, i_8_156_1453_0, i_8_156_1454_0, i_8_156_1537_0,
    i_8_156_1604_0, i_8_156_1623_0, i_8_156_1630_0, i_8_156_1631_0,
    i_8_156_1634_0, i_8_156_1650_0, i_8_156_1677_0, i_8_156_1678_0,
    i_8_156_1679_0, i_8_156_1701_0, i_8_156_1746_0, i_8_156_1751_0,
    i_8_156_1771_0, i_8_156_1792_0, i_8_156_1793_0, i_8_156_1794_0,
    i_8_156_1795_0, i_8_156_1855_0, i_8_156_1856_0, i_8_156_1858_0,
    i_8_156_1876_0, i_8_156_1877_0, i_8_156_1912_0, i_8_156_1980_0,
    i_8_156_1981_0, i_8_156_1984_0, i_8_156_1985_0, i_8_156_1993_0,
    i_8_156_2056_0, i_8_156_2057_0, i_8_156_2129_0, i_8_156_2143_0,
    i_8_156_2144_0, i_8_156_2156_0, i_8_156_2272_0,
    o_8_156_0_0  );
  input  i_8_156_35_0, i_8_156_37_0, i_8_156_77_0, i_8_156_87_0,
    i_8_156_111_0, i_8_156_140_0, i_8_156_229_0, i_8_156_235_0,
    i_8_156_259_0, i_8_156_304_0, i_8_156_355_0, i_8_156_382_0,
    i_8_156_418_0, i_8_156_419_0, i_8_156_442_0, i_8_156_445_0,
    i_8_156_446_0, i_8_156_464_0, i_8_156_490_0, i_8_156_504_0,
    i_8_156_505_0, i_8_156_506_0, i_8_156_507_0, i_8_156_508_0,
    i_8_156_509_0, i_8_156_528_0, i_8_156_610_0, i_8_156_621_0,
    i_8_156_625_0, i_8_156_665_0, i_8_156_698_0, i_8_156_748_0,
    i_8_156_780_0, i_8_156_781_0, i_8_156_845_0, i_8_156_876_0,
    i_8_156_880_0, i_8_156_885_0, i_8_156_967_0, i_8_156_1028_0,
    i_8_156_1030_0, i_8_156_1031_0, i_8_156_1136_0, i_8_156_1158_0,
    i_8_156_1192_0, i_8_156_1200_0, i_8_156_1201_0, i_8_156_1202_0,
    i_8_156_1225_0, i_8_156_1269_0, i_8_156_1281_0, i_8_156_1315_0,
    i_8_156_1325_0, i_8_156_1328_0, i_8_156_1350_0, i_8_156_1355_0,
    i_8_156_1387_0, i_8_156_1398_0, i_8_156_1399_0, i_8_156_1400_0,
    i_8_156_1437_0, i_8_156_1450_0, i_8_156_1453_0, i_8_156_1454_0,
    i_8_156_1537_0, i_8_156_1604_0, i_8_156_1623_0, i_8_156_1630_0,
    i_8_156_1631_0, i_8_156_1634_0, i_8_156_1650_0, i_8_156_1677_0,
    i_8_156_1678_0, i_8_156_1679_0, i_8_156_1701_0, i_8_156_1746_0,
    i_8_156_1751_0, i_8_156_1771_0, i_8_156_1792_0, i_8_156_1793_0,
    i_8_156_1794_0, i_8_156_1795_0, i_8_156_1855_0, i_8_156_1856_0,
    i_8_156_1858_0, i_8_156_1876_0, i_8_156_1877_0, i_8_156_1912_0,
    i_8_156_1980_0, i_8_156_1981_0, i_8_156_1984_0, i_8_156_1985_0,
    i_8_156_1993_0, i_8_156_2056_0, i_8_156_2057_0, i_8_156_2129_0,
    i_8_156_2143_0, i_8_156_2144_0, i_8_156_2156_0, i_8_156_2272_0;
  output o_8_156_0_0;
  assign o_8_156_0_0 = ~((~i_8_156_1793_0 & ((i_8_156_111_0 & ((~i_8_156_259_0 & ~i_8_156_419_0 & ~i_8_156_445_0 & ~i_8_156_508_0 & ~i_8_156_1158_0 & ~i_8_156_1631_0 & ~i_8_156_1746_0 & ~i_8_156_1794_0) | (~i_8_156_140_0 & ~i_8_156_235_0 & ~i_8_156_355_0 & ~i_8_156_504_0 & ~i_8_156_1201_0 & ~i_8_156_1858_0 & ~i_8_156_1912_0 & i_8_156_1993_0))) | (~i_8_156_507_0 & ((~i_8_156_140_0 & ((~i_8_156_37_0 & ~i_8_156_442_0 & ~i_8_156_464_0 & i_8_156_698_0 & ~i_8_156_1325_0 & ~i_8_156_1328_0 & ~i_8_156_1912_0) | (~i_8_156_77_0 & ~i_8_156_355_0 & ~i_8_156_504_0 & ~i_8_156_508_0 & ~i_8_156_509_0 & ~i_8_156_1136_0 & ~i_8_156_1192_0 & ~i_8_156_1201_0 & ~i_8_156_1679_0 & ~i_8_156_1985_0))) | (~i_8_156_419_0 & ~i_8_156_446_0 & ~i_8_156_880_0 & ~i_8_156_1192_0 & ~i_8_156_1281_0 & ~i_8_156_1325_0 & ~i_8_156_1398_0 & ~i_8_156_1399_0 & ~i_8_156_1701_0 & ~i_8_156_1746_0 & ~i_8_156_1792_0 & ~i_8_156_1877_0 & ~i_8_156_2129_0))) | (~i_8_156_1876_0 & ((~i_8_156_37_0 & ((~i_8_156_446_0 & ~i_8_156_508_0 & i_8_156_780_0) | (i_8_156_304_0 & ~i_8_156_419_0 & ~i_8_156_464_0 & i_8_156_880_0 & ~i_8_156_1200_0 & ~i_8_156_1269_0 & ~i_8_156_1315_0 & ~i_8_156_1325_0 & ~i_8_156_1701_0 & ~i_8_156_1912_0))) | (~i_8_156_464_0 & ~i_8_156_505_0 & ~i_8_156_876_0 & i_8_156_880_0 & ~i_8_156_1028_0 & ~i_8_156_1398_0 & ~i_8_156_1437_0 & ~i_8_156_1771_0 & ~i_8_156_1877_0))) | (~i_8_156_528_0 & ((~i_8_156_77_0 & ((~i_8_156_509_0 & ~i_8_156_967_0 & ~i_8_156_1387_0 & ~i_8_156_1400_0 & ~i_8_156_1701_0 & ~i_8_156_1912_0 & i_8_156_1981_0) | (~i_8_156_419_0 & ~i_8_156_446_0 & ~i_8_156_1201_0 & ~i_8_156_1315_0 & ~i_8_156_1630_0 & ~i_8_156_1746_0 & ~i_8_156_1792_0 & ~i_8_156_1993_0 & ~i_8_156_2144_0))) | (~i_8_156_259_0 & ~i_8_156_504_0 & ~i_8_156_505_0 & ~i_8_156_665_0 & ~i_8_156_781_0 & ~i_8_156_1202_0 & ~i_8_156_1269_0 & ~i_8_156_1328_0 & ~i_8_156_1400_0 & ~i_8_156_1677_0 & ~i_8_156_1751_0 & ~i_8_156_1771_0 & ~i_8_156_1795_0))))) | (~i_8_156_77_0 & ((~i_8_156_445_0 & ~i_8_156_506_0 & ~i_8_156_1325_0 & i_8_156_1678_0 & i_8_156_1858_0) | (~i_8_156_442_0 & ~i_8_156_508_0 & ~i_8_156_509_0 & ~i_8_156_780_0 & ~i_8_156_880_0 & ~i_8_156_1350_0 & ~i_8_156_1387_0 & ~i_8_156_1400_0 & ~i_8_156_1746_0 & ~i_8_156_1792_0 & ~i_8_156_1993_0))) | (~i_8_156_442_0 & ((~i_8_156_418_0 & ~i_8_156_446_0 & ~i_8_156_505_0 & ~i_8_156_507_0 & ~i_8_156_509_0 & ~i_8_156_967_0 & ~i_8_156_1192_0 & ~i_8_156_1631_0 & ~i_8_156_1634_0 & ~i_8_156_1794_0) | (~i_8_156_506_0 & ~i_8_156_1399_0 & ~i_8_156_1630_0 & i_8_156_1856_0))) | (~i_8_156_505_0 & ((~i_8_156_419_0 & ~i_8_156_446_0 & ((~i_8_156_304_0 & ~i_8_156_504_0 & ~i_8_156_1202_0 & ~i_8_156_1877_0 & ((~i_8_156_464_0 & ~i_8_156_490_0 & ~i_8_156_1315_0 & ~i_8_156_1325_0 & ~i_8_156_1350_0 & ~i_8_156_1792_0 & ~i_8_156_1795_0 & ~i_8_156_1980_0 & ~i_8_156_2129_0) | (~i_8_156_37_0 & ~i_8_156_140_0 & ~i_8_156_418_0 & ~i_8_156_507_0 & ~i_8_156_845_0 & ~i_8_156_2143_0))) | (~i_8_156_508_0 & ~i_8_156_509_0 & ~i_8_156_1269_0 & ~i_8_156_1325_0 & ~i_8_156_1355_0 & ~i_8_156_1398_0 & ~i_8_156_1604_0 & ~i_8_156_1701_0 & ~i_8_156_1876_0 & ~i_8_156_2272_0))) | (~i_8_156_1630_0 & ((~i_8_156_508_0 & ~i_8_156_509_0 & ~i_8_156_418_0 & ~i_8_156_507_0 & ~i_8_156_1634_0 & ~i_8_156_1794_0 & ~i_8_156_1328_0 & ~i_8_156_1631_0) | (~i_8_156_445_0 & i_8_156_876_0 & ~i_8_156_1450_0 & ~i_8_156_1751_0 & ~i_8_156_1876_0 & ~i_8_156_1912_0))) | (~i_8_156_355_0 & i_8_156_625_0 & ~i_8_156_1269_0 & ~i_8_156_1701_0 & ~i_8_156_1912_0 & ~i_8_156_1281_0 & i_8_156_1678_0))) | (~i_8_156_504_0 & ((~i_8_156_140_0 & ((~i_8_156_506_0 & i_8_156_1985_0 & i_8_156_2129_0) | (~i_8_156_304_0 & ~i_8_156_464_0 & ~i_8_156_610_0 & ~i_8_156_748_0 & ~i_8_156_1200_0 & ~i_8_156_1269_0 & ~i_8_156_1328_0 & ~i_8_156_1604_0 & ~i_8_156_1792_0 & ~i_8_156_1794_0 & ~i_8_156_1795_0 & ~i_8_156_1876_0 & ~i_8_156_1877_0 & ~i_8_156_1912_0 & ~i_8_156_2144_0))) | (~i_8_156_748_0 & ((~i_8_156_506_0 & ~i_8_156_665_0 & ~i_8_156_1355_0 & ~i_8_156_1398_0 & ~i_8_156_1399_0 & ~i_8_156_1400_0 & ~i_8_156_1604_0 & ~i_8_156_1876_0 & ~i_8_156_1877_0 & ~i_8_156_1993_0) | (~i_8_156_111_0 & ~i_8_156_509_0 & i_8_156_967_0 & ~i_8_156_1136_0 & ~i_8_156_1158_0 & ~i_8_156_1200_0 & ~i_8_156_1315_0 & ~i_8_156_1325_0 & ~i_8_156_1328_0 & ~i_8_156_1792_0 & ~i_8_156_1794_0 & ~i_8_156_2272_0))))) | (~i_8_156_419_0 & ((~i_8_156_355_0 & ~i_8_156_1792_0 & ((~i_8_156_445_0 & ~i_8_156_621_0 & ~i_8_156_748_0 & ~i_8_156_967_0 & ~i_8_156_1225_0 & i_8_156_1281_0 & ~i_8_156_1315_0 & ~i_8_156_1630_0 & ~i_8_156_1634_0 & ~i_8_156_1981_0) | (~i_8_156_509_0 & ~i_8_156_528_0 & i_8_156_610_0 & ~i_8_156_845_0 & ~i_8_156_885_0 & ~i_8_156_1650_0 & ~i_8_156_1701_0 & ~i_8_156_1912_0 & ~i_8_156_2129_0))) | (~i_8_156_610_0 & ~i_8_156_1202_0 & ~i_8_156_1315_0 & ~i_8_156_1701_0 & i_8_156_1858_0 & ~i_8_156_1980_0 & ~i_8_156_2129_0 & ~i_8_156_2156_0))) | (~i_8_156_1634_0 & ((i_8_156_382_0 & ~i_8_156_507_0 & ~i_8_156_1355_0 & ~i_8_156_1630_0 & ~i_8_156_1631_0) | (~i_8_156_1399_0 & i_8_156_1450_0 & i_8_156_1679_0 & i_8_156_2272_0))) | (~i_8_156_507_0 & ((~i_8_156_446_0 & ~i_8_156_1200_0 & ~i_8_156_1328_0 & i_8_156_1678_0 & i_8_156_1984_0) | (i_8_156_1202_0 & ~i_8_156_1387_0 & i_8_156_1454_0 & ~i_8_156_1981_0 & ~i_8_156_1993_0 & ~i_8_156_2057_0))) | (~i_8_156_229_0 & ~i_8_156_845_0 & ~i_8_156_967_0 & ~i_8_156_1269_0 & ~i_8_156_1325_0 & ~i_8_156_1398_0 & ~i_8_156_1400_0 & i_8_156_1678_0 & ~i_8_156_1792_0 & ~i_8_156_1993_0) | (i_8_156_1030_0 & i_8_156_1453_0 & ~i_8_156_1795_0 & ~i_8_156_1912_0));
endmodule



// Benchmark "kernel_8_157" written by ABC on Sun Jul 19 10:05:44 2020

module kernel_8_157 ( 
    i_8_157_25_0, i_8_157_33_0, i_8_157_72_0, i_8_157_96_0, i_8_157_97_0,
    i_8_157_214_0, i_8_157_215_0, i_8_157_220_0, i_8_157_241_0,
    i_8_157_286_0, i_8_157_295_0, i_8_157_301_0, i_8_157_348_0,
    i_8_157_361_0, i_8_157_367_0, i_8_157_376_0, i_8_157_385_0,
    i_8_157_421_0, i_8_157_445_0, i_8_157_457_0, i_8_157_467_0,
    i_8_157_484_0, i_8_157_485_0, i_8_157_525_0, i_8_157_555_0,
    i_8_157_592_0, i_8_157_593_0, i_8_157_610_0, i_8_157_611_0,
    i_8_157_616_0, i_8_157_630_0, i_8_157_715_0, i_8_157_718_0,
    i_8_157_719_0, i_8_157_760_0, i_8_157_763_0, i_8_157_764_0,
    i_8_157_772_0, i_8_157_799_0, i_8_157_838_0, i_8_157_889_0,
    i_8_157_925_0, i_8_157_952_0, i_8_157_991_0, i_8_157_1012_0,
    i_8_157_1015_0, i_8_157_1016_0, i_8_157_1029_0, i_8_157_1030_0,
    i_8_157_1114_0, i_8_157_1124_0, i_8_157_1160_0, i_8_157_1237_0,
    i_8_157_1258_0, i_8_157_1263_0, i_8_157_1264_0, i_8_157_1273_0,
    i_8_157_1300_0, i_8_157_1305_0, i_8_157_1306_0, i_8_157_1331_0,
    i_8_157_1344_0, i_8_157_1363_0, i_8_157_1387_0, i_8_157_1438_0,
    i_8_157_1455_0, i_8_157_1456_0, i_8_157_1544_0, i_8_157_1600_0,
    i_8_157_1601_0, i_8_157_1632_0, i_8_157_1644_0, i_8_157_1680_0,
    i_8_157_1735_0, i_8_157_1748_0, i_8_157_1749_0, i_8_157_1754_0,
    i_8_157_1818_0, i_8_157_1867_0, i_8_157_1869_0, i_8_157_1894_0,
    i_8_157_1897_0, i_8_157_1903_0, i_8_157_1921_0, i_8_157_1922_0,
    i_8_157_1967_0, i_8_157_1969_0, i_8_157_2020_0, i_8_157_2056_0,
    i_8_157_2092_0, i_8_157_2114_0, i_8_157_2131_0, i_8_157_2157_0,
    i_8_157_2218_0, i_8_157_2266_0, i_8_157_2274_0, i_8_157_2275_0,
    i_8_157_2292_0, i_8_157_2293_0, i_8_157_2294_0,
    o_8_157_0_0  );
  input  i_8_157_25_0, i_8_157_33_0, i_8_157_72_0, i_8_157_96_0,
    i_8_157_97_0, i_8_157_214_0, i_8_157_215_0, i_8_157_220_0,
    i_8_157_241_0, i_8_157_286_0, i_8_157_295_0, i_8_157_301_0,
    i_8_157_348_0, i_8_157_361_0, i_8_157_367_0, i_8_157_376_0,
    i_8_157_385_0, i_8_157_421_0, i_8_157_445_0, i_8_157_457_0,
    i_8_157_467_0, i_8_157_484_0, i_8_157_485_0, i_8_157_525_0,
    i_8_157_555_0, i_8_157_592_0, i_8_157_593_0, i_8_157_610_0,
    i_8_157_611_0, i_8_157_616_0, i_8_157_630_0, i_8_157_715_0,
    i_8_157_718_0, i_8_157_719_0, i_8_157_760_0, i_8_157_763_0,
    i_8_157_764_0, i_8_157_772_0, i_8_157_799_0, i_8_157_838_0,
    i_8_157_889_0, i_8_157_925_0, i_8_157_952_0, i_8_157_991_0,
    i_8_157_1012_0, i_8_157_1015_0, i_8_157_1016_0, i_8_157_1029_0,
    i_8_157_1030_0, i_8_157_1114_0, i_8_157_1124_0, i_8_157_1160_0,
    i_8_157_1237_0, i_8_157_1258_0, i_8_157_1263_0, i_8_157_1264_0,
    i_8_157_1273_0, i_8_157_1300_0, i_8_157_1305_0, i_8_157_1306_0,
    i_8_157_1331_0, i_8_157_1344_0, i_8_157_1363_0, i_8_157_1387_0,
    i_8_157_1438_0, i_8_157_1455_0, i_8_157_1456_0, i_8_157_1544_0,
    i_8_157_1600_0, i_8_157_1601_0, i_8_157_1632_0, i_8_157_1644_0,
    i_8_157_1680_0, i_8_157_1735_0, i_8_157_1748_0, i_8_157_1749_0,
    i_8_157_1754_0, i_8_157_1818_0, i_8_157_1867_0, i_8_157_1869_0,
    i_8_157_1894_0, i_8_157_1897_0, i_8_157_1903_0, i_8_157_1921_0,
    i_8_157_1922_0, i_8_157_1967_0, i_8_157_1969_0, i_8_157_2020_0,
    i_8_157_2056_0, i_8_157_2092_0, i_8_157_2114_0, i_8_157_2131_0,
    i_8_157_2157_0, i_8_157_2218_0, i_8_157_2266_0, i_8_157_2274_0,
    i_8_157_2275_0, i_8_157_2292_0, i_8_157_2293_0, i_8_157_2294_0;
  output o_8_157_0_0;
  assign o_8_157_0_0 = 0;
endmodule



// Benchmark "kernel_8_158" written by ABC on Sun Jul 19 10:05:45 2020

module kernel_8_158 ( 
    i_8_158_6_0, i_8_158_76_0, i_8_158_78_0, i_8_158_79_0, i_8_158_114_0,
    i_8_158_157_0, i_8_158_159_0, i_8_158_204_0, i_8_158_205_0,
    i_8_158_240_0, i_8_158_241_0, i_8_158_249_0, i_8_158_256_0,
    i_8_158_259_0, i_8_158_301_0, i_8_158_312_0, i_8_158_313_0,
    i_8_158_327_0, i_8_158_348_0, i_8_158_366_0, i_8_158_429_0,
    i_8_158_453_0, i_8_158_499_0, i_8_158_507_0, i_8_158_553_0,
    i_8_158_570_0, i_8_158_574_0, i_8_158_597_0, i_8_158_600_0,
    i_8_158_606_0, i_8_158_660_0, i_8_158_665_0, i_8_158_687_0,
    i_8_158_690_0, i_8_158_771_0, i_8_158_777_0, i_8_158_778_0,
    i_8_158_783_0, i_8_158_849_0, i_8_158_885_0, i_8_158_943_0,
    i_8_158_993_0, i_8_158_1028_0, i_8_158_1037_0, i_8_158_1048_0,
    i_8_158_1056_0, i_8_158_1059_0, i_8_158_1077_0, i_8_158_1104_0,
    i_8_158_1138_0, i_8_158_1146_0, i_8_158_1182_0, i_8_158_1227_0,
    i_8_158_1228_0, i_8_158_1294_0, i_8_158_1306_0, i_8_158_1371_0,
    i_8_158_1410_0, i_8_158_1436_0, i_8_158_1455_0, i_8_158_1510_0,
    i_8_158_1624_0, i_8_158_1626_0, i_8_158_1629_0, i_8_158_1644_0,
    i_8_158_1653_0, i_8_158_1654_0, i_8_158_1689_0, i_8_158_1705_0,
    i_8_158_1748_0, i_8_158_1750_0, i_8_158_1753_0, i_8_158_1754_0,
    i_8_158_1808_0, i_8_158_1823_0, i_8_158_1837_0, i_8_158_1860_0,
    i_8_158_1861_0, i_8_158_1863_0, i_8_158_1884_0, i_8_158_1887_0,
    i_8_158_1983_0, i_8_158_1984_0, i_8_158_1986_0, i_8_158_2046_0,
    i_8_158_2055_0, i_8_158_2058_0, i_8_158_2073_0, i_8_158_2074_0,
    i_8_158_2076_0, i_8_158_2085_0, i_8_158_2086_0, i_8_158_2141_0,
    i_8_158_2146_0, i_8_158_2150_0, i_8_158_2157_0, i_8_158_2217_0,
    i_8_158_2244_0, i_8_158_2274_0, i_8_158_2275_0,
    o_8_158_0_0  );
  input  i_8_158_6_0, i_8_158_76_0, i_8_158_78_0, i_8_158_79_0,
    i_8_158_114_0, i_8_158_157_0, i_8_158_159_0, i_8_158_204_0,
    i_8_158_205_0, i_8_158_240_0, i_8_158_241_0, i_8_158_249_0,
    i_8_158_256_0, i_8_158_259_0, i_8_158_301_0, i_8_158_312_0,
    i_8_158_313_0, i_8_158_327_0, i_8_158_348_0, i_8_158_366_0,
    i_8_158_429_0, i_8_158_453_0, i_8_158_499_0, i_8_158_507_0,
    i_8_158_553_0, i_8_158_570_0, i_8_158_574_0, i_8_158_597_0,
    i_8_158_600_0, i_8_158_606_0, i_8_158_660_0, i_8_158_665_0,
    i_8_158_687_0, i_8_158_690_0, i_8_158_771_0, i_8_158_777_0,
    i_8_158_778_0, i_8_158_783_0, i_8_158_849_0, i_8_158_885_0,
    i_8_158_943_0, i_8_158_993_0, i_8_158_1028_0, i_8_158_1037_0,
    i_8_158_1048_0, i_8_158_1056_0, i_8_158_1059_0, i_8_158_1077_0,
    i_8_158_1104_0, i_8_158_1138_0, i_8_158_1146_0, i_8_158_1182_0,
    i_8_158_1227_0, i_8_158_1228_0, i_8_158_1294_0, i_8_158_1306_0,
    i_8_158_1371_0, i_8_158_1410_0, i_8_158_1436_0, i_8_158_1455_0,
    i_8_158_1510_0, i_8_158_1624_0, i_8_158_1626_0, i_8_158_1629_0,
    i_8_158_1644_0, i_8_158_1653_0, i_8_158_1654_0, i_8_158_1689_0,
    i_8_158_1705_0, i_8_158_1748_0, i_8_158_1750_0, i_8_158_1753_0,
    i_8_158_1754_0, i_8_158_1808_0, i_8_158_1823_0, i_8_158_1837_0,
    i_8_158_1860_0, i_8_158_1861_0, i_8_158_1863_0, i_8_158_1884_0,
    i_8_158_1887_0, i_8_158_1983_0, i_8_158_1984_0, i_8_158_1986_0,
    i_8_158_2046_0, i_8_158_2055_0, i_8_158_2058_0, i_8_158_2073_0,
    i_8_158_2074_0, i_8_158_2076_0, i_8_158_2085_0, i_8_158_2086_0,
    i_8_158_2141_0, i_8_158_2146_0, i_8_158_2150_0, i_8_158_2157_0,
    i_8_158_2217_0, i_8_158_2244_0, i_8_158_2274_0, i_8_158_2275_0;
  output o_8_158_0_0;
  assign o_8_158_0_0 = ~((~i_8_158_204_0 & ((~i_8_158_943_0 & ~i_8_158_1077_0 & ~i_8_158_1410_0 & ~i_8_158_1689_0 & ~i_8_158_1860_0 & ~i_8_158_2046_0 & ~i_8_158_2085_0) | (~i_8_158_205_0 & ~i_8_158_327_0 & ~i_8_158_366_0 & ~i_8_158_429_0 & ~i_8_158_453_0 & ~i_8_158_1104_0 & ~i_8_158_1624_0 & ~i_8_158_1837_0 & ~i_8_158_2086_0 & ~i_8_158_2141_0))) | (~i_8_158_312_0 & ~i_8_158_348_0 & ((i_8_158_79_0 & ~i_8_158_1059_0) | (~i_8_158_240_0 & i_8_158_1624_0 & ~i_8_158_1689_0 & ~i_8_158_1887_0 & ~i_8_158_2076_0 & ~i_8_158_2085_0))) | (~i_8_158_240_0 & ((~i_8_158_570_0 & ~i_8_158_1059_0 & ~i_8_158_1626_0 & ~i_8_158_1861_0) | (~i_8_158_606_0 & ~i_8_158_885_0 & ~i_8_158_1510_0 & ~i_8_158_1887_0))) | (~i_8_158_327_0 & ((~i_8_158_79_0 & ~i_8_158_690_0 & ~i_8_158_1048_0 & ~i_8_158_1371_0 & i_8_158_2074_0) | (~i_8_158_570_0 & ~i_8_158_574_0 & ~i_8_158_771_0 & i_8_158_1410_0 & ~i_8_158_1689_0 & ~i_8_158_1986_0 & ~i_8_158_2085_0))) | (~i_8_158_690_0 & ((~i_8_158_570_0 & ~i_8_158_606_0 & ~i_8_158_778_0 & ~i_8_158_1048_0 & ~i_8_158_1705_0 & ~i_8_158_1986_0 & i_8_158_2274_0) | (~i_8_158_993_0 & ~i_8_158_1059_0 & ~i_8_158_1146_0 & ~i_8_158_2274_0))) | (~i_8_158_2157_0 & ((i_8_158_366_0 & ~i_8_158_1056_0 & ~i_8_158_1629_0 & ~i_8_158_1653_0) | (i_8_158_553_0 & i_8_158_660_0 & ~i_8_158_778_0 & ~i_8_158_1983_0))) | (~i_8_158_1056_0 & ((~i_8_158_313_0 & ~i_8_158_1048_0 & ~i_8_158_2055_0 & ~i_8_158_2058_0) | (~i_8_158_600_0 & ~i_8_158_1306_0 & ~i_8_158_1689_0 & ~i_8_158_1986_0 & ~i_8_158_2074_0))) | (~i_8_158_1653_0 & ((~i_8_158_114_0 & ~i_8_158_1624_0 & ~i_8_158_1626_0) | (~i_8_158_943_0 & ~i_8_158_1455_0 & ~i_8_158_2073_0 & ~i_8_158_2086_0 & ~i_8_158_2275_0))) | (i_8_158_159_0 & i_8_158_1808_0));
endmodule



// Benchmark "kernel_8_159" written by ABC on Sun Jul 19 10:05:46 2020

module kernel_8_159 ( 
    i_8_159_26_0, i_8_159_50_0, i_8_159_76_0, i_8_159_88_0, i_8_159_93_0,
    i_8_159_106_0, i_8_159_250_0, i_8_159_266_0, i_8_159_282_0,
    i_8_159_286_0, i_8_159_291_0, i_8_159_321_0, i_8_159_383_0,
    i_8_159_384_0, i_8_159_436_0, i_8_159_437_0, i_8_159_453_0,
    i_8_159_454_0, i_8_159_456_0, i_8_159_491_0, i_8_159_555_0,
    i_8_159_624_0, i_8_159_633_0, i_8_159_636_0, i_8_159_642_0,
    i_8_159_643_0, i_8_159_672_0, i_8_159_687_0, i_8_159_696_0,
    i_8_159_703_0, i_8_159_718_0, i_8_159_727_0, i_8_159_728_0,
    i_8_159_730_0, i_8_159_735_0, i_8_159_736_0, i_8_159_782_0,
    i_8_159_814_0, i_8_159_834_0, i_8_159_843_0, i_8_159_848_0,
    i_8_159_852_0, i_8_159_933_0, i_8_159_1074_0, i_8_159_1088_0,
    i_8_159_1138_0, i_8_159_1185_0, i_8_159_1213_0, i_8_159_1221_0,
    i_8_159_1222_0, i_8_159_1227_0, i_8_159_1228_0, i_8_159_1236_0,
    i_8_159_1237_0, i_8_159_1239_0, i_8_159_1266_0, i_8_159_1281_0,
    i_8_159_1290_0, i_8_159_1309_0, i_8_159_1349_0, i_8_159_1384_0,
    i_8_159_1390_0, i_8_159_1446_0, i_8_159_1455_0, i_8_159_1545_0,
    i_8_159_1561_0, i_8_159_1580_0, i_8_159_1617_0, i_8_159_1624_0,
    i_8_159_1653_0, i_8_159_1654_0, i_8_159_1704_0, i_8_159_1706_0,
    i_8_159_1723_0, i_8_159_1770_0, i_8_159_1808_0, i_8_159_1825_0,
    i_8_159_1843_0, i_8_159_1849_0, i_8_159_1860_0, i_8_159_1903_0,
    i_8_159_1989_0, i_8_159_1992_0, i_8_159_1995_0, i_8_159_2010_0,
    i_8_159_2019_0, i_8_159_2031_0, i_8_159_2040_0, i_8_159_2084_0,
    i_8_159_2131_0, i_8_159_2138_0, i_8_159_2147_0, i_8_159_2158_0,
    i_8_159_2173_0, i_8_159_2194_0, i_8_159_2226_0, i_8_159_2247_0,
    i_8_159_2263_0, i_8_159_2284_0, i_8_159_2289_0,
    o_8_159_0_0  );
  input  i_8_159_26_0, i_8_159_50_0, i_8_159_76_0, i_8_159_88_0,
    i_8_159_93_0, i_8_159_106_0, i_8_159_250_0, i_8_159_266_0,
    i_8_159_282_0, i_8_159_286_0, i_8_159_291_0, i_8_159_321_0,
    i_8_159_383_0, i_8_159_384_0, i_8_159_436_0, i_8_159_437_0,
    i_8_159_453_0, i_8_159_454_0, i_8_159_456_0, i_8_159_491_0,
    i_8_159_555_0, i_8_159_624_0, i_8_159_633_0, i_8_159_636_0,
    i_8_159_642_0, i_8_159_643_0, i_8_159_672_0, i_8_159_687_0,
    i_8_159_696_0, i_8_159_703_0, i_8_159_718_0, i_8_159_727_0,
    i_8_159_728_0, i_8_159_730_0, i_8_159_735_0, i_8_159_736_0,
    i_8_159_782_0, i_8_159_814_0, i_8_159_834_0, i_8_159_843_0,
    i_8_159_848_0, i_8_159_852_0, i_8_159_933_0, i_8_159_1074_0,
    i_8_159_1088_0, i_8_159_1138_0, i_8_159_1185_0, i_8_159_1213_0,
    i_8_159_1221_0, i_8_159_1222_0, i_8_159_1227_0, i_8_159_1228_0,
    i_8_159_1236_0, i_8_159_1237_0, i_8_159_1239_0, i_8_159_1266_0,
    i_8_159_1281_0, i_8_159_1290_0, i_8_159_1309_0, i_8_159_1349_0,
    i_8_159_1384_0, i_8_159_1390_0, i_8_159_1446_0, i_8_159_1455_0,
    i_8_159_1545_0, i_8_159_1561_0, i_8_159_1580_0, i_8_159_1617_0,
    i_8_159_1624_0, i_8_159_1653_0, i_8_159_1654_0, i_8_159_1704_0,
    i_8_159_1706_0, i_8_159_1723_0, i_8_159_1770_0, i_8_159_1808_0,
    i_8_159_1825_0, i_8_159_1843_0, i_8_159_1849_0, i_8_159_1860_0,
    i_8_159_1903_0, i_8_159_1989_0, i_8_159_1992_0, i_8_159_1995_0,
    i_8_159_2010_0, i_8_159_2019_0, i_8_159_2031_0, i_8_159_2040_0,
    i_8_159_2084_0, i_8_159_2131_0, i_8_159_2138_0, i_8_159_2147_0,
    i_8_159_2158_0, i_8_159_2173_0, i_8_159_2194_0, i_8_159_2226_0,
    i_8_159_2247_0, i_8_159_2263_0, i_8_159_2284_0, i_8_159_2289_0;
  output o_8_159_0_0;
  assign o_8_159_0_0 = 0;
endmodule



// Benchmark "kernel_8_160" written by ABC on Sun Jul 19 10:05:48 2020

module kernel_8_160 ( 
    i_8_160_31_0, i_8_160_34_0, i_8_160_35_0, i_8_160_46_0, i_8_160_52_0,
    i_8_160_53_0, i_8_160_59_0, i_8_160_80_0, i_8_160_94_0, i_8_160_95_0,
    i_8_160_98_0, i_8_160_115_0, i_8_160_184_0, i_8_160_232_0,
    i_8_160_233_0, i_8_160_304_0, i_8_160_314_0, i_8_160_329_0,
    i_8_160_349_0, i_8_160_381_0, i_8_160_425_0, i_8_160_454_0,
    i_8_160_455_0, i_8_160_503_0, i_8_160_552_0, i_8_160_556_0,
    i_8_160_557_0, i_8_160_614_0, i_8_160_696_0, i_8_160_698_0,
    i_8_160_706_0, i_8_160_956_0, i_8_160_967_0, i_8_160_968_0,
    i_8_160_992_0, i_8_160_994_0, i_8_160_1048_0, i_8_160_1049_0,
    i_8_160_1052_0, i_8_160_1075_0, i_8_160_1094_0, i_8_160_1110_0,
    i_8_160_1115_0, i_8_160_1135_0, i_8_160_1179_0, i_8_160_1183_0,
    i_8_160_1263_0, i_8_160_1271_0, i_8_160_1274_0, i_8_160_1282_0,
    i_8_160_1291_0, i_8_160_1306_0, i_8_160_1307_0, i_8_160_1325_0,
    i_8_160_1339_0, i_8_160_1348_0, i_8_160_1352_0, i_8_160_1355_0,
    i_8_160_1372_0, i_8_160_1388_0, i_8_160_1435_0, i_8_160_1436_0,
    i_8_160_1437_0, i_8_160_1438_0, i_8_160_1439_0, i_8_160_1506_0,
    i_8_160_1507_0, i_8_160_1535_0, i_8_160_1625_0, i_8_160_1627_0,
    i_8_160_1628_0, i_8_160_1636_0, i_8_160_1676_0, i_8_160_1677_0,
    i_8_160_1678_0, i_8_160_1679_0, i_8_160_1682_0, i_8_160_1750_0,
    i_8_160_1764_0, i_8_160_1784_0, i_8_160_1807_0, i_8_160_1822_0,
    i_8_160_1873_0, i_8_160_1876_0, i_8_160_1906_0, i_8_160_1907_0,
    i_8_160_1963_0, i_8_160_1966_0, i_8_160_1981_0, i_8_160_1982_0,
    i_8_160_2006_0, i_8_160_2032_0, i_8_160_2050_0, i_8_160_2093_0,
    i_8_160_2096_0, i_8_160_2109_0, i_8_160_2152_0, i_8_160_2216_0,
    i_8_160_2281_0, i_8_160_2282_0,
    o_8_160_0_0  );
  input  i_8_160_31_0, i_8_160_34_0, i_8_160_35_0, i_8_160_46_0,
    i_8_160_52_0, i_8_160_53_0, i_8_160_59_0, i_8_160_80_0, i_8_160_94_0,
    i_8_160_95_0, i_8_160_98_0, i_8_160_115_0, i_8_160_184_0,
    i_8_160_232_0, i_8_160_233_0, i_8_160_304_0, i_8_160_314_0,
    i_8_160_329_0, i_8_160_349_0, i_8_160_381_0, i_8_160_425_0,
    i_8_160_454_0, i_8_160_455_0, i_8_160_503_0, i_8_160_552_0,
    i_8_160_556_0, i_8_160_557_0, i_8_160_614_0, i_8_160_696_0,
    i_8_160_698_0, i_8_160_706_0, i_8_160_956_0, i_8_160_967_0,
    i_8_160_968_0, i_8_160_992_0, i_8_160_994_0, i_8_160_1048_0,
    i_8_160_1049_0, i_8_160_1052_0, i_8_160_1075_0, i_8_160_1094_0,
    i_8_160_1110_0, i_8_160_1115_0, i_8_160_1135_0, i_8_160_1179_0,
    i_8_160_1183_0, i_8_160_1263_0, i_8_160_1271_0, i_8_160_1274_0,
    i_8_160_1282_0, i_8_160_1291_0, i_8_160_1306_0, i_8_160_1307_0,
    i_8_160_1325_0, i_8_160_1339_0, i_8_160_1348_0, i_8_160_1352_0,
    i_8_160_1355_0, i_8_160_1372_0, i_8_160_1388_0, i_8_160_1435_0,
    i_8_160_1436_0, i_8_160_1437_0, i_8_160_1438_0, i_8_160_1439_0,
    i_8_160_1506_0, i_8_160_1507_0, i_8_160_1535_0, i_8_160_1625_0,
    i_8_160_1627_0, i_8_160_1628_0, i_8_160_1636_0, i_8_160_1676_0,
    i_8_160_1677_0, i_8_160_1678_0, i_8_160_1679_0, i_8_160_1682_0,
    i_8_160_1750_0, i_8_160_1764_0, i_8_160_1784_0, i_8_160_1807_0,
    i_8_160_1822_0, i_8_160_1873_0, i_8_160_1876_0, i_8_160_1906_0,
    i_8_160_1907_0, i_8_160_1963_0, i_8_160_1966_0, i_8_160_1981_0,
    i_8_160_1982_0, i_8_160_2006_0, i_8_160_2032_0, i_8_160_2050_0,
    i_8_160_2093_0, i_8_160_2096_0, i_8_160_2109_0, i_8_160_2152_0,
    i_8_160_2216_0, i_8_160_2281_0, i_8_160_2282_0;
  output o_8_160_0_0;
  assign o_8_160_0_0 = ~((~i_8_160_1907_0 & ((~i_8_160_2281_0 & ((~i_8_160_31_0 & ~i_8_160_454_0 & ((~i_8_160_232_0 & ~i_8_160_968_0 & ~i_8_160_1388_0 & i_8_160_1750_0 & ~i_8_160_2050_0) | (i_8_160_80_0 & ~i_8_160_1271_0 & ~i_8_160_1306_0 & ~i_8_160_1372_0 & ~i_8_160_1625_0 & ~i_8_160_2216_0))) | (i_8_160_46_0 & ~i_8_160_94_0 & ~i_8_160_115_0 & ~i_8_160_329_0 & ~i_8_160_1306_0 & ~i_8_160_1507_0 & ~i_8_160_1676_0 & ~i_8_160_1873_0 & ~i_8_160_2216_0) | (~i_8_160_53_0 & ~i_8_160_95_0 & ~i_8_160_314_0 & ~i_8_160_706_0 & ~i_8_160_1388_0 & i_8_160_1438_0 & ~i_8_160_1822_0 & ~i_8_160_1876_0 & ~i_8_160_2282_0))) | (~i_8_160_1628_0 & ((~i_8_160_59_0 & ~i_8_160_233_0 & ((~i_8_160_232_0 & ~i_8_160_314_0 & ~i_8_160_329_0 & ~i_8_160_1049_0 & ~i_8_160_1052_0 & ~i_8_160_1094_0 & ~i_8_160_1372_0 & i_8_160_2093_0) | (~i_8_160_35_0 & ~i_8_160_115_0 & ~i_8_160_614_0 & i_8_160_1435_0 & ~i_8_160_2006_0 & ~i_8_160_2032_0 & ~i_8_160_2152_0 & ~i_8_160_2282_0))) | (~i_8_160_956_0 & ((~i_8_160_94_0 & ~i_8_160_994_0 & ~i_8_160_1049_0 & ~i_8_160_1052_0 & ~i_8_160_1094_0 & ~i_8_160_1306_0 & ~i_8_160_1372_0 & ~i_8_160_1388_0 & ~i_8_160_1625_0 & ~i_8_160_1627_0 & ~i_8_160_1906_0) | (~i_8_160_381_0 & ~i_8_160_1183_0 & ~i_8_160_1291_0 & i_8_160_1535_0 & i_8_160_1679_0 & ~i_8_160_1807_0 & ~i_8_160_2032_0 & ~i_8_160_2096_0))))) | (~i_8_160_115_0 & ~i_8_160_1049_0 & ((~i_8_160_53_0 & ~i_8_160_98_0 & ~i_8_160_696_0 & ~i_8_160_1075_0 & ~i_8_160_1094_0 & ~i_8_160_1352_0 & ~i_8_160_1507_0 & ~i_8_160_1963_0 & ~i_8_160_1966_0) | (~i_8_160_52_0 & ~i_8_160_454_0 & ~i_8_160_967_0 & ~i_8_160_1306_0 & ~i_8_160_1355_0 & ~i_8_160_1873_0 & ~i_8_160_2109_0 & ~i_8_160_2282_0))) | (~i_8_160_1876_0 & ((~i_8_160_698_0 & ~i_8_160_1274_0 & i_8_160_1676_0 & ~i_8_160_1966_0) | (~i_8_160_34_0 & ~i_8_160_95_0 & i_8_160_425_0 & ~i_8_160_1307_0 & ~i_8_160_1372_0 & ~i_8_160_1388_0 & ~i_8_160_1873_0 & ~i_8_160_2032_0 & ~i_8_160_2093_0) | (~i_8_160_1325_0 & ~i_8_160_1352_0 & i_8_160_1963_0 & ~i_8_160_2006_0 & ~i_8_160_2096_0 & i_8_160_2152_0))) | (~i_8_160_94_0 & ~i_8_160_314_0 & ~i_8_160_329_0 & i_8_160_455_0 & ~i_8_160_696_0 & ~i_8_160_992_0 & ~i_8_160_1306_0 & ~i_8_160_2216_0 & ~i_8_160_2282_0))) | (~i_8_160_115_0 & ((~i_8_160_184_0 & ~i_8_160_425_0 & ~i_8_160_455_0 & i_8_160_967_0 & i_8_160_994_0 & ~i_8_160_1627_0 & ~i_8_160_1682_0 & ~i_8_160_1906_0 & ~i_8_160_2093_0) | (~i_8_160_53_0 & ~i_8_160_956_0 & ~i_8_160_968_0 & ~i_8_160_1052_0 & ~i_8_160_1388_0 & ~i_8_160_1535_0 & ~i_8_160_1628_0 & ~i_8_160_1678_0 & ~i_8_160_1876_0 & ~i_8_160_2096_0 & ~i_8_160_2109_0 & ~i_8_160_2281_0 & ~i_8_160_2282_0))) | (~i_8_160_304_0 & ((~i_8_160_94_0 & ~i_8_160_329_0 & ~i_8_160_956_0 & ~i_8_160_1052_0 & i_8_160_1263_0 & ~i_8_160_1625_0 & ~i_8_160_1628_0 & ~i_8_160_1679_0 & ~i_8_160_1873_0) | (~i_8_160_52_0 & ~i_8_160_233_0 & i_8_160_552_0 & ~i_8_160_698_0 & ~i_8_160_1348_0 & ~i_8_160_1352_0 & ~i_8_160_1636_0 & ~i_8_160_2006_0 & ~i_8_160_2282_0))) | (~i_8_160_52_0 & ((~i_8_160_706_0 & ~i_8_160_968_0 & ~i_8_160_1325_0 & ~i_8_160_1506_0 & ~i_8_160_1507_0 & i_8_160_1678_0 & ~i_8_160_1873_0 & ~i_8_160_1876_0) | (~i_8_160_1274_0 & ~i_8_160_1355_0 & i_8_160_1636_0 & ~i_8_160_1676_0 & ~i_8_160_2281_0))) | (~i_8_160_1388_0 & ((~i_8_160_1873_0 & ((~i_8_160_94_0 & ((~i_8_160_53_0 & ~i_8_160_967_0 & ~i_8_160_968_0 & ~i_8_160_1352_0 & ~i_8_160_1625_0 & i_8_160_1750_0) | (~i_8_160_95_0 & ~i_8_160_98_0 & ~i_8_160_503_0 & ~i_8_160_994_0 & ~i_8_160_1052_0 & ~i_8_160_1094_0 & ~i_8_160_1274_0 & ~i_8_160_1307_0 & ~i_8_160_1372_0 & ~i_8_160_1507_0 & ~i_8_160_1627_0 & ~i_8_160_1906_0))) | (~i_8_160_34_0 & ~i_8_160_95_0 & ~i_8_160_184_0 & ~i_8_160_233_0 & i_8_160_1110_0 & ~i_8_160_1625_0 & ~i_8_160_1627_0 & ~i_8_160_1628_0))) | (~i_8_160_232_0 & ((~i_8_160_314_0 & ~i_8_160_1372_0 & ~i_8_160_2096_0 & ((~i_8_160_59_0 & ~i_8_160_698_0 & i_8_160_967_0 & ~i_8_160_1094_0 & ~i_8_160_1627_0 & ~i_8_160_1906_0 & ~i_8_160_1307_0 & ~i_8_160_1535_0) | (~i_8_160_329_0 & ~i_8_160_967_0 & ~i_8_160_1183_0 & ~i_8_160_1506_0 & ~i_8_160_1507_0 & ~i_8_160_1625_0 & ~i_8_160_1628_0 & ~i_8_160_2032_0 & ~i_8_160_2216_0))) | (~i_8_160_95_0 & ~i_8_160_233_0 & ~i_8_160_614_0 & ~i_8_160_992_0 & i_8_160_1348_0 & ~i_8_160_1507_0 & ~i_8_160_1906_0 & ~i_8_160_2281_0))) | (~i_8_160_706_0 & ~i_8_160_994_0 & ~i_8_160_1052_0 & ~i_8_160_1325_0 & i_8_160_1355_0 & ~i_8_160_1372_0 & ~i_8_160_1506_0 & ~i_8_160_1625_0 & ~i_8_160_1628_0 & ~i_8_160_1807_0 & ~i_8_160_1906_0 & ~i_8_160_2093_0 & ~i_8_160_2096_0))) | (~i_8_160_53_0 & ((i_8_160_52_0 & i_8_160_115_0 & ~i_8_160_454_0 & ~i_8_160_967_0 & ~i_8_160_994_0 & ~i_8_160_1750_0) | (~i_8_160_1094_0 & ~i_8_160_1271_0 & ~i_8_160_1355_0 & ~i_8_160_1372_0 & ~i_8_160_1506_0 & ~i_8_160_1628_0 & ~i_8_160_1876_0 & ~i_8_160_1906_0 & ~i_8_160_2281_0))) | (~i_8_160_95_0 & ((~i_8_160_35_0 & ~i_8_160_967_0 & ~i_8_160_1135_0 & ~i_8_160_1627_0 & i_8_160_1677_0 & ~i_8_160_1873_0 & ~i_8_160_2050_0) | (i_8_160_503_0 & ~i_8_160_1507_0 & i_8_160_1966_0 & ~i_8_160_2282_0))) | (~i_8_160_98_0 & ((i_8_160_614_0 & i_8_160_698_0 & i_8_160_1282_0 & ~i_8_160_1678_0 & ~i_8_160_1876_0 & ~i_8_160_1352_0 & ~i_8_160_1625_0) | (~i_8_160_314_0 & ~i_8_160_552_0 & ~i_8_160_1049_0 & ~i_8_160_1075_0 & ~i_8_160_1306_0 & ~i_8_160_1355_0 & i_8_160_1438_0 & ~i_8_160_2109_0 & ~i_8_160_2281_0))) | (~i_8_160_184_0 & ((~i_8_160_956_0 & ~i_8_160_992_0 & ~i_8_160_994_0 & i_8_160_1049_0 & ~i_8_160_1052_0 & ~i_8_160_1075_0 & ~i_8_160_1094_0 & ~i_8_160_1627_0 & ~i_8_160_1963_0 & ~i_8_160_2281_0) | (~i_8_160_94_0 & ~i_8_160_552_0 & i_8_160_557_0 & ~i_8_160_1873_0 & ~i_8_160_1876_0 & ~i_8_160_1906_0 & ~i_8_160_2096_0 & ~i_8_160_2282_0))) | (~i_8_160_46_0 & i_8_160_556_0 & ~i_8_160_698_0 & ~i_8_160_956_0 & ~i_8_160_1048_0 & ~i_8_160_1325_0 & ~i_8_160_1339_0 & ~i_8_160_1628_0 & ~i_8_160_1981_0) | (i_8_160_696_0 & i_8_160_706_0 & ~i_8_160_1052_0 & ~i_8_160_1271_0 & ~i_8_160_1627_0 & ~i_8_160_1873_0 & ~i_8_160_1963_0 & ~i_8_160_2032_0 & ~i_8_160_2093_0 & ~i_8_160_2109_0) | (~i_8_160_1115_0 & ~i_8_160_1307_0 & ~i_8_160_1355_0 & ~i_8_160_1625_0 & i_8_160_1679_0 & ~i_8_160_1750_0 & ~i_8_160_1764_0 & ~i_8_160_2216_0));
endmodule



// Benchmark "kernel_8_161" written by ABC on Sun Jul 19 10:05:49 2020

module kernel_8_161 ( 
    i_8_161_20_0, i_8_161_23_0, i_8_161_43_0, i_8_161_88_0, i_8_161_121_0,
    i_8_161_131_0, i_8_161_194_0, i_8_161_230_0, i_8_161_232_0,
    i_8_161_247_0, i_8_161_278_0, i_8_161_310_0, i_8_161_311_0,
    i_8_161_314_0, i_8_161_325_0, i_8_161_363_0, i_8_161_367_0,
    i_8_161_393_0, i_8_161_419_0, i_8_161_430_0, i_8_161_473_0,
    i_8_161_492_0, i_8_161_634_0, i_8_161_693_0, i_8_161_706_0,
    i_8_161_709_0, i_8_161_751_0, i_8_161_790_0, i_8_161_799_0,
    i_8_161_825_0, i_8_161_831_0, i_8_161_838_0, i_8_161_842_0,
    i_8_161_844_0, i_8_161_850_0, i_8_161_878_0, i_8_161_879_0,
    i_8_161_880_0, i_8_161_886_0, i_8_161_887_0, i_8_161_953_0,
    i_8_161_964_0, i_8_161_968_0, i_8_161_970_0, i_8_161_986_0,
    i_8_161_994_0, i_8_161_1016_0, i_8_161_1039_0, i_8_161_1040_0,
    i_8_161_1048_0, i_8_161_1063_0, i_8_161_1075_0, i_8_161_1076_0,
    i_8_161_1102_0, i_8_161_1113_0, i_8_161_1127_0, i_8_161_1165_0,
    i_8_161_1239_0, i_8_161_1240_0, i_8_161_1246_0, i_8_161_1318_0,
    i_8_161_1336_0, i_8_161_1372_0, i_8_161_1399_0, i_8_161_1407_0,
    i_8_161_1470_0, i_8_161_1498_0, i_8_161_1528_0, i_8_161_1607_0,
    i_8_161_1609_0, i_8_161_1641_0, i_8_161_1645_0, i_8_161_1653_0,
    i_8_161_1690_0, i_8_161_1691_0, i_8_161_1704_0, i_8_161_1708_0,
    i_8_161_1733_0, i_8_161_1746_0, i_8_161_1751_0, i_8_161_1767_0,
    i_8_161_1769_0, i_8_161_1870_0, i_8_161_1884_0, i_8_161_1896_0,
    i_8_161_1906_0, i_8_161_1984_0, i_8_161_2039_0, i_8_161_2042_0,
    i_8_161_2066_0, i_8_161_2072_0, i_8_161_2075_0, i_8_161_2086_0,
    i_8_161_2089_0, i_8_161_2119_0, i_8_161_2153_0, i_8_161_2174_0,
    i_8_161_2227_0, i_8_161_2232_0, i_8_161_2275_0,
    o_8_161_0_0  );
  input  i_8_161_20_0, i_8_161_23_0, i_8_161_43_0, i_8_161_88_0,
    i_8_161_121_0, i_8_161_131_0, i_8_161_194_0, i_8_161_230_0,
    i_8_161_232_0, i_8_161_247_0, i_8_161_278_0, i_8_161_310_0,
    i_8_161_311_0, i_8_161_314_0, i_8_161_325_0, i_8_161_363_0,
    i_8_161_367_0, i_8_161_393_0, i_8_161_419_0, i_8_161_430_0,
    i_8_161_473_0, i_8_161_492_0, i_8_161_634_0, i_8_161_693_0,
    i_8_161_706_0, i_8_161_709_0, i_8_161_751_0, i_8_161_790_0,
    i_8_161_799_0, i_8_161_825_0, i_8_161_831_0, i_8_161_838_0,
    i_8_161_842_0, i_8_161_844_0, i_8_161_850_0, i_8_161_878_0,
    i_8_161_879_0, i_8_161_880_0, i_8_161_886_0, i_8_161_887_0,
    i_8_161_953_0, i_8_161_964_0, i_8_161_968_0, i_8_161_970_0,
    i_8_161_986_0, i_8_161_994_0, i_8_161_1016_0, i_8_161_1039_0,
    i_8_161_1040_0, i_8_161_1048_0, i_8_161_1063_0, i_8_161_1075_0,
    i_8_161_1076_0, i_8_161_1102_0, i_8_161_1113_0, i_8_161_1127_0,
    i_8_161_1165_0, i_8_161_1239_0, i_8_161_1240_0, i_8_161_1246_0,
    i_8_161_1318_0, i_8_161_1336_0, i_8_161_1372_0, i_8_161_1399_0,
    i_8_161_1407_0, i_8_161_1470_0, i_8_161_1498_0, i_8_161_1528_0,
    i_8_161_1607_0, i_8_161_1609_0, i_8_161_1641_0, i_8_161_1645_0,
    i_8_161_1653_0, i_8_161_1690_0, i_8_161_1691_0, i_8_161_1704_0,
    i_8_161_1708_0, i_8_161_1733_0, i_8_161_1746_0, i_8_161_1751_0,
    i_8_161_1767_0, i_8_161_1769_0, i_8_161_1870_0, i_8_161_1884_0,
    i_8_161_1896_0, i_8_161_1906_0, i_8_161_1984_0, i_8_161_2039_0,
    i_8_161_2042_0, i_8_161_2066_0, i_8_161_2072_0, i_8_161_2075_0,
    i_8_161_2086_0, i_8_161_2089_0, i_8_161_2119_0, i_8_161_2153_0,
    i_8_161_2174_0, i_8_161_2227_0, i_8_161_2232_0, i_8_161_2275_0;
  output o_8_161_0_0;
  assign o_8_161_0_0 = 0;
endmodule



// Benchmark "kernel_8_162" written by ABC on Sun Jul 19 10:05:50 2020

module kernel_8_162 ( 
    i_8_162_23_0, i_8_162_25_0, i_8_162_138_0, i_8_162_139_0,
    i_8_162_140_0, i_8_162_141_0, i_8_162_143_0, i_8_162_194_0,
    i_8_162_228_0, i_8_162_282_0, i_8_162_286_0, i_8_162_287_0,
    i_8_162_318_0, i_8_162_320_0, i_8_162_398_0, i_8_162_404_0,
    i_8_162_440_0, i_8_162_504_0, i_8_162_580_0, i_8_162_583_0,
    i_8_162_641_0, i_8_162_642_0, i_8_162_694_0, i_8_162_727_0,
    i_8_162_823_0, i_8_162_858_0, i_8_162_859_0, i_8_162_873_0,
    i_8_162_877_0, i_8_162_882_0, i_8_162_885_0, i_8_162_972_0,
    i_8_162_973_0, i_8_162_974_0, i_8_162_976_0, i_8_162_977_0,
    i_8_162_979_0, i_8_162_980_0, i_8_162_1030_0, i_8_162_1040_0,
    i_8_162_1187_0, i_8_162_1198_0, i_8_162_1238_0, i_8_162_1362_0,
    i_8_162_1367_0, i_8_162_1410_0, i_8_162_1426_0, i_8_162_1427_0,
    i_8_162_1440_0, i_8_162_1443_0, i_8_162_1444_0, i_8_162_1447_0,
    i_8_162_1462_0, i_8_162_1470_0, i_8_162_1471_0, i_8_162_1525_0,
    i_8_162_1526_0, i_8_162_1529_0, i_8_162_1534_0, i_8_162_1600_0,
    i_8_162_1604_0, i_8_162_1606_0, i_8_162_1641_0, i_8_162_1669_0,
    i_8_162_1679_0, i_8_162_1697_0, i_8_162_1718_0, i_8_162_1726_0,
    i_8_162_1777_0, i_8_162_1808_0, i_8_162_1905_0, i_8_162_1944_0,
    i_8_162_1965_0, i_8_162_1966_0, i_8_162_1967_0, i_8_162_1969_0,
    i_8_162_1970_0, i_8_162_1975_0, i_8_162_1983_0, i_8_162_2011_0,
    i_8_162_2031_0, i_8_162_2052_0, i_8_162_2055_0, i_8_162_2056_0,
    i_8_162_2057_0, i_8_162_2109_0, i_8_162_2110_0, i_8_162_2112_0,
    i_8_162_2137_0, i_8_162_2154_0, i_8_162_2155_0, i_8_162_2159_0,
    i_8_162_2172_0, i_8_162_2173_0, i_8_162_2176_0, i_8_162_2232_0,
    i_8_162_2233_0, i_8_162_2234_0, i_8_162_2246_0, i_8_162_2249_0,
    o_8_162_0_0  );
  input  i_8_162_23_0, i_8_162_25_0, i_8_162_138_0, i_8_162_139_0,
    i_8_162_140_0, i_8_162_141_0, i_8_162_143_0, i_8_162_194_0,
    i_8_162_228_0, i_8_162_282_0, i_8_162_286_0, i_8_162_287_0,
    i_8_162_318_0, i_8_162_320_0, i_8_162_398_0, i_8_162_404_0,
    i_8_162_440_0, i_8_162_504_0, i_8_162_580_0, i_8_162_583_0,
    i_8_162_641_0, i_8_162_642_0, i_8_162_694_0, i_8_162_727_0,
    i_8_162_823_0, i_8_162_858_0, i_8_162_859_0, i_8_162_873_0,
    i_8_162_877_0, i_8_162_882_0, i_8_162_885_0, i_8_162_972_0,
    i_8_162_973_0, i_8_162_974_0, i_8_162_976_0, i_8_162_977_0,
    i_8_162_979_0, i_8_162_980_0, i_8_162_1030_0, i_8_162_1040_0,
    i_8_162_1187_0, i_8_162_1198_0, i_8_162_1238_0, i_8_162_1362_0,
    i_8_162_1367_0, i_8_162_1410_0, i_8_162_1426_0, i_8_162_1427_0,
    i_8_162_1440_0, i_8_162_1443_0, i_8_162_1444_0, i_8_162_1447_0,
    i_8_162_1462_0, i_8_162_1470_0, i_8_162_1471_0, i_8_162_1525_0,
    i_8_162_1526_0, i_8_162_1529_0, i_8_162_1534_0, i_8_162_1600_0,
    i_8_162_1604_0, i_8_162_1606_0, i_8_162_1641_0, i_8_162_1669_0,
    i_8_162_1679_0, i_8_162_1697_0, i_8_162_1718_0, i_8_162_1726_0,
    i_8_162_1777_0, i_8_162_1808_0, i_8_162_1905_0, i_8_162_1944_0,
    i_8_162_1965_0, i_8_162_1966_0, i_8_162_1967_0, i_8_162_1969_0,
    i_8_162_1970_0, i_8_162_1975_0, i_8_162_1983_0, i_8_162_2011_0,
    i_8_162_2031_0, i_8_162_2052_0, i_8_162_2055_0, i_8_162_2056_0,
    i_8_162_2057_0, i_8_162_2109_0, i_8_162_2110_0, i_8_162_2112_0,
    i_8_162_2137_0, i_8_162_2154_0, i_8_162_2155_0, i_8_162_2159_0,
    i_8_162_2172_0, i_8_162_2173_0, i_8_162_2176_0, i_8_162_2232_0,
    i_8_162_2233_0, i_8_162_2234_0, i_8_162_2246_0, i_8_162_2249_0;
  output o_8_162_0_0;
  assign o_8_162_0_0 = ~((~i_8_162_25_0 & ((i_8_162_23_0 & ~i_8_162_141_0 & ~i_8_162_320_0 & ~i_8_162_583_0 & ~i_8_162_974_0 & ~i_8_162_1198_0 & ~i_8_162_1529_0 & ~i_8_162_1726_0) | (~i_8_162_287_0 & ~i_8_162_1187_0 & ~i_8_162_1443_0 & ~i_8_162_1444_0 & ~i_8_162_1447_0 & i_8_162_2056_0 & i_8_162_2155_0))) | (i_8_162_138_0 & ((~i_8_162_318_0 & ~i_8_162_1030_0 & ~i_8_162_1447_0 & i_8_162_1777_0 & ~i_8_162_1969_0 & ~i_8_162_2031_0 & i_8_162_2154_0 & ~i_8_162_2155_0) | (~i_8_162_23_0 & i_8_162_139_0 & ~i_8_162_583_0 & ~i_8_162_641_0 & ~i_8_162_823_0 & ~i_8_162_973_0 & ~i_8_162_1440_0 & i_8_162_1471_0 & ~i_8_162_1526_0 & ~i_8_162_1726_0 & ~i_8_162_2246_0))) | (~i_8_162_2137_0 & ((i_8_162_139_0 & ((~i_8_162_143_0 & ~i_8_162_694_0 & i_8_162_877_0 & ~i_8_162_1443_0 & ~i_8_162_1726_0 & i_8_162_1966_0) | (~i_8_162_320_0 & ~i_8_162_974_0 & i_8_162_1238_0 & ~i_8_162_1367_0 & ~i_8_162_1534_0 & i_8_162_1967_0))) | (~i_8_162_143_0 & ~i_8_162_1526_0 & i_8_162_1679_0 & ~i_8_162_2031_0 & ((~i_8_162_504_0 & ~i_8_162_694_0 & ~i_8_162_823_0 & ~i_8_162_1187_0 & ~i_8_162_1198_0 & ~i_8_162_1808_0 & ~i_8_162_1967_0 & ~i_8_162_2057_0 & ~i_8_162_2159_0) | (~i_8_162_139_0 & ~i_8_162_140_0 & ~i_8_162_320_0 & ~i_8_162_398_0 & ~i_8_162_404_0 & ~i_8_162_641_0 & ~i_8_162_1367_0 & ~i_8_162_1427_0 & ~i_8_162_1440_0 & ~i_8_162_1444_0 & ~i_8_162_1944_0 & ~i_8_162_2233_0))) | (~i_8_162_287_0 & ~i_8_162_398_0 & i_8_162_694_0 & ~i_8_162_823_0 & ~i_8_162_877_0 & ~i_8_162_972_0 & ~i_8_162_974_0 & ~i_8_162_1040_0 & ~i_8_162_1198_0 & ~i_8_162_1238_0 & ~i_8_162_1443_0 & ~i_8_162_1697_0 & ~i_8_162_2057_0) | (~i_8_162_138_0 & i_8_162_873_0 & i_8_162_877_0 & i_8_162_1777_0))) | (~i_8_162_972_0 & ((~i_8_162_141_0 & ((~i_8_162_823_0 & i_8_162_885_0 & ~i_8_162_1944_0) | (~i_8_162_140_0 & i_8_162_194_0 & ~i_8_162_974_0 & ~i_8_162_979_0 & ~i_8_162_980_0 & ~i_8_162_1427_0 & ~i_8_162_1526_0 & ~i_8_162_1905_0 & i_8_162_1969_0))) | (~i_8_162_1443_0 & ((~i_8_162_140_0 & ((~i_8_162_143_0 & ~i_8_162_282_0 & ~i_8_162_398_0 & ~i_8_162_580_0 & ~i_8_162_1470_0 & ~i_8_162_1471_0 & ~i_8_162_1534_0 & ~i_8_162_1669_0 & i_8_162_1777_0 & i_8_162_1965_0 & ~i_8_162_1969_0 & ~i_8_162_2155_0 & ~i_8_162_2159_0) | (~i_8_162_823_0 & i_8_162_882_0 & ~i_8_162_1238_0 & ~i_8_162_2011_0 & ~i_8_162_2176_0))) | (~i_8_162_320_0 & ~i_8_162_823_0 & ~i_8_162_973_0 & ~i_8_162_1187_0 & ~i_8_162_1427_0 & ~i_8_162_1718_0 & ~i_8_162_1905_0 & ~i_8_162_2011_0 & ~i_8_162_2031_0 & i_8_162_2233_0 & ~i_8_162_2246_0))) | (~i_8_162_642_0 & ((i_8_162_228_0 & ~i_8_162_318_0 & ~i_8_162_580_0 & i_8_162_877_0 & ~i_8_162_1447_0 & ~i_8_162_1525_0 & ~i_8_162_2031_0) | (~i_8_162_641_0 & ~i_8_162_823_0 & ~i_8_162_973_0 & ~i_8_162_974_0 & ~i_8_162_1444_0 & i_8_162_1534_0 & ~i_8_162_1679_0 & ~i_8_162_1726_0 & ~i_8_162_1969_0 & ~i_8_162_2234_0))) | (~i_8_162_973_0 & ((~i_8_162_404_0 & ~i_8_162_583_0 & ~i_8_162_727_0 & i_8_162_1969_0 & ~i_8_162_2011_0 & i_8_162_2112_0) | (i_8_162_194_0 & i_8_162_504_0 & ~i_8_162_885_0 & ~i_8_162_977_0 & ~i_8_162_1238_0 & ~i_8_162_1905_0 & ~i_8_162_1970_0 & ~i_8_162_2159_0))) | (~i_8_162_979_0 & ~i_8_162_1040_0 & ~i_8_162_1198_0 & ~i_8_162_1444_0 & ~i_8_162_1905_0 & ~i_8_162_2031_0 & i_8_162_2112_0))) | (i_8_162_228_0 & ((~i_8_162_1426_0 & ~i_8_162_1443_0 & ~i_8_162_1447_0 & i_8_162_1470_0 & ~i_8_162_1529_0 & ~i_8_162_2031_0) | (i_8_162_2109_0 & i_8_162_2172_0))) | (~i_8_162_580_0 & ((~i_8_162_139_0 & ~i_8_162_1426_0 & ~i_8_162_1427_0 & i_8_162_1966_0 & i_8_162_2233_0) | (~i_8_162_398_0 & ~i_8_162_504_0 & ~i_8_162_976_0 & ~i_8_162_1529_0 & ~i_8_162_1726_0 & i_8_162_1967_0 & ~i_8_162_2031_0 & i_8_162_2234_0))) | (~i_8_162_1526_0 & ((~i_8_162_398_0 & ((~i_8_162_141_0 & ~i_8_162_320_0 & ~i_8_162_727_0 & ~i_8_162_977_0 & ~i_8_162_980_0 & ~i_8_162_1030_0 & ~i_8_162_1187_0 & ~i_8_162_1726_0 & ~i_8_162_1777_0 & i_8_162_2056_0) | (~i_8_162_641_0 & ~i_8_162_979_0 & ~i_8_162_1427_0 & ~i_8_162_1965_0 & i_8_162_1967_0 & ~i_8_162_2031_0 & i_8_162_2057_0))) | (~i_8_162_139_0 & ~i_8_162_143_0 & ~i_8_162_1808_0 & ~i_8_162_1967_0 & ~i_8_162_1970_0 & ~i_8_162_2155_0 & ~i_8_162_2246_0 & i_8_162_2249_0) | (~i_8_162_138_0 & ~i_8_162_504_0 & ~i_8_162_727_0 & i_8_162_1669_0 & i_8_162_2155_0 & ~i_8_162_2249_0))) | (~i_8_162_1198_0 & ((~i_8_162_140_0 & ((~i_8_162_398_0 & ((~i_8_162_440_0 & ~i_8_162_823_0 & ~i_8_162_980_0 & ~i_8_162_1040_0 & ~i_8_162_1187_0 & ~i_8_162_1367_0 & ~i_8_162_1726_0 & ~i_8_162_1944_0 & i_8_162_1970_0) | (~i_8_162_143_0 & ~i_8_162_641_0 & ~i_8_162_1238_0 & i_8_162_2234_0))) | (~i_8_162_641_0 & ~i_8_162_823_0 & ~i_8_162_974_0 & i_8_162_1604_0 & ~i_8_162_1669_0) | (~i_8_162_139_0 & ~i_8_162_141_0 & ~i_8_162_504_0 & ~i_8_162_1030_0 & ~i_8_162_1426_0 & i_8_162_1444_0 & ~i_8_162_2246_0 & ~i_8_162_2249_0))) | (~i_8_162_141_0 & ((~i_8_162_504_0 & ~i_8_162_873_0 & ~i_8_162_1726_0 & ~i_8_162_1969_0 & ~i_8_162_2031_0 & i_8_162_2052_0) | (~i_8_162_143_0 & ~i_8_162_642_0 & ~i_8_162_1529_0 & ~i_8_162_1679_0 & i_8_162_1965_0 & i_8_162_2176_0))) | (~i_8_162_823_0 & ((~i_8_162_1362_0 & i_8_162_1444_0 & i_8_162_1983_0 & ~i_8_162_2172_0) | (~i_8_162_885_0 & ~i_8_162_1238_0 & ~i_8_162_1447_0 & ~i_8_162_1525_0 & ~i_8_162_1726_0 & ~i_8_162_1966_0 & i_8_162_2011_0 & ~i_8_162_2249_0))) | (~i_8_162_1529_0 & ((~i_8_162_976_0 & ((~i_8_162_286_0 & ~i_8_162_504_0 & ~i_8_162_977_0 & ~i_8_162_1726_0 & ~i_8_162_2031_0 & i_8_162_2055_0) | (~i_8_162_404_0 & ~i_8_162_882_0 & ~i_8_162_974_0 & ~i_8_162_980_0 & ~i_8_162_1426_0 & ~i_8_162_1447_0 & i_8_162_1679_0 & i_8_162_1970_0 & ~i_8_162_2172_0))) | (~i_8_162_977_0 & ((~i_8_162_320_0 & i_8_162_1534_0 & i_8_162_1679_0) | (~i_8_162_1040_0 & ~i_8_162_1967_0 & i_8_162_1969_0 & ~i_8_162_2011_0 & i_8_162_2057_0))))) | (~i_8_162_1669_0 & ((~i_8_162_1040_0 & i_8_162_1604_0 & ~i_8_162_1679_0 & ~i_8_162_1966_0 & ~i_8_162_1967_0) | (~i_8_162_138_0 & ~i_8_162_143_0 & ~i_8_162_583_0 & ~i_8_162_1426_0 & ~i_8_162_1440_0 & ~i_8_162_1944_0 & i_8_162_1983_0) | (i_8_162_882_0 & ~i_8_162_1606_0 & i_8_162_2052_0))))) | (~i_8_162_140_0 & ((~i_8_162_139_0 & ~i_8_162_282_0 & ~i_8_162_404_0 & ~i_8_162_973_0 & ~i_8_162_1367_0 & ~i_8_162_1462_0 & ~i_8_162_1718_0 & ~i_8_162_1726_0 & ~i_8_162_1905_0 & i_8_162_1965_0 & i_8_162_1969_0) | (i_8_162_877_0 & ~i_8_162_1040_0 & ~i_8_162_1777_0 & ~i_8_162_1966_0 & ~i_8_162_2031_0 & i_8_162_2155_0))) | (~i_8_162_1440_0 & ((~i_8_162_139_0 & ((~i_8_162_286_0 & ~i_8_162_398_0 & ~i_8_162_1410_0 & i_8_162_1777_0 & i_8_162_2057_0) | (~i_8_162_143_0 & ~i_8_162_823_0 & ~i_8_162_973_0 & ~i_8_162_1040_0 & ~i_8_162_1187_0 & ~i_8_162_1238_0 & ~i_8_162_1447_0 & ~i_8_162_1529_0 & ~i_8_162_1726_0 & i_8_162_1966_0 & ~i_8_162_1967_0 & ~i_8_162_1969_0 & ~i_8_162_2057_0 & ~i_8_162_2246_0))) | (~i_8_162_980_0 & ~i_8_162_1726_0 & ((i_8_162_25_0 & ~i_8_162_286_0 & ~i_8_162_320_0 & ~i_8_162_974_0 & ~i_8_162_1187_0 & ~i_8_162_1427_0 & i_8_162_1970_0) | (i_8_162_873_0 & ~i_8_162_1367_0 & ~i_8_162_1462_0 & ~i_8_162_1905_0 & i_8_162_2052_0))) | (~i_8_162_398_0 & ~i_8_162_977_0 & ~i_8_162_1187_0 & i_8_162_1965_0 & i_8_162_1967_0 & ~i_8_162_1969_0 & ~i_8_162_2176_0))) | (~i_8_162_138_0 & ((~i_8_162_143_0 & ((~i_8_162_139_0 & ~i_8_162_320_0 & ~i_8_162_1427_0 & ((~i_8_162_287_0 & ~i_8_162_318_0 & ~i_8_162_440_0 & ~i_8_162_973_0 & ~i_8_162_1238_0 & ~i_8_162_1367_0 & i_8_162_1471_0 & ~i_8_162_1529_0 & ~i_8_162_2246_0) | (~i_8_162_641_0 & ~i_8_162_977_0 & ~i_8_162_1187_0 & ~i_8_162_1525_0 & ~i_8_162_1534_0 & ~i_8_162_1965_0 & i_8_162_1967_0 & ~i_8_162_2172_0 & ~i_8_162_2249_0))) | (~i_8_162_141_0 & ~i_8_162_1187_0 & ~i_8_162_1447_0 & ~i_8_162_2031_0 & i_8_162_2154_0 & i_8_162_2155_0))) | (~i_8_162_1443_0 & i_8_162_1777_0 & i_8_162_2112_0) | (i_8_162_885_0 & ~i_8_162_973_0 & i_8_162_2172_0))) | (~i_8_162_139_0 & ((~i_8_162_141_0 & ~i_8_162_404_0 & ~i_8_162_642_0 & ~i_8_162_1187_0 & ~i_8_162_1444_0 & ~i_8_162_1718_0 & i_8_162_1969_0 & i_8_162_2173_0) | (~i_8_162_143_0 & ~i_8_162_858_0 & ~i_8_162_1362_0 & i_8_162_1410_0 & ~i_8_162_1426_0 & ~i_8_162_1529_0 & ~i_8_162_1534_0 & ~i_8_162_1969_0 & ~i_8_162_2031_0 & ~i_8_162_2056_0 & ~i_8_162_2233_0))) | (~i_8_162_1362_0 & ((~i_8_162_1444_0 & ~i_8_162_1447_0 & ~i_8_162_1040_0 & ~i_8_162_1443_0 & ~i_8_162_2031_0 & i_8_162_2112_0 & ~i_8_162_1471_0 & ~i_8_162_1726_0) | (~i_8_162_286_0 & i_8_162_1470_0 & i_8_162_2109_0 & ~i_8_162_2246_0))) | (~i_8_162_1970_0 & ((~i_8_162_1447_0 & ((~i_8_162_1470_0 & i_8_162_2154_0 & i_8_162_2232_0) | (~i_8_162_141_0 & ~i_8_162_143_0 & ~i_8_162_404_0 & ~i_8_162_1187_0 & ~i_8_162_1529_0 & ~i_8_162_1679_0 & i_8_162_1808_0 & ~i_8_162_1905_0 & ~i_8_162_2056_0 & ~i_8_162_2246_0))) | (~i_8_162_440_0 & i_8_162_1808_0 & i_8_162_1966_0 & i_8_162_1969_0 & i_8_162_2246_0))) | (i_8_162_1965_0 & ((~i_8_162_504_0 & ~i_8_162_1238_0 & ~i_8_162_1427_0 & ~i_8_162_1447_0 & ~i_8_162_1726_0 & i_8_162_2055_0) | (~i_8_162_877_0 & ~i_8_162_980_0 & ~i_8_162_1777_0 & ~i_8_162_1905_0 & i_8_162_2154_0 & ~i_8_162_2173_0))) | (~i_8_162_642_0 & ~i_8_162_1471_0 & i_8_162_1641_0 & i_8_162_2232_0));
endmodule



// Benchmark "kernel_8_163" written by ABC on Sun Jul 19 10:05:51 2020

module kernel_8_163 ( 
    i_8_163_103_0, i_8_163_140_0, i_8_163_220_0, i_8_163_226_0,
    i_8_163_230_0, i_8_163_247_0, i_8_163_256_0, i_8_163_262_0,
    i_8_163_299_0, i_8_163_304_0, i_8_163_314_0, i_8_163_316_0,
    i_8_163_326_0, i_8_163_363_0, i_8_163_367_0, i_8_163_381_0,
    i_8_163_418_0, i_8_163_428_0, i_8_163_454_0, i_8_163_455_0,
    i_8_163_553_0, i_8_163_581_0, i_8_163_582_0, i_8_163_584_0,
    i_8_163_599_0, i_8_163_635_0, i_8_163_793_0, i_8_163_823_0,
    i_8_163_839_0, i_8_163_840_0, i_8_163_844_0, i_8_163_845_0,
    i_8_163_859_0, i_8_163_874_0, i_8_163_881_0, i_8_163_882_0,
    i_8_163_891_0, i_8_163_994_0, i_8_163_1145_0, i_8_163_1147_0,
    i_8_163_1226_0, i_8_163_1229_0, i_8_163_1268_0, i_8_163_1282_0,
    i_8_163_1286_0, i_8_163_1319_0, i_8_163_1399_0, i_8_163_1403_0,
    i_8_163_1432_0, i_8_163_1435_0, i_8_163_1436_0, i_8_163_1438_0,
    i_8_163_1463_0, i_8_163_1470_0, i_8_163_1510_0, i_8_163_1562_0,
    i_8_163_1574_0, i_8_163_1668_0, i_8_163_1688_0, i_8_163_1690_0,
    i_8_163_1704_0, i_8_163_1774_0, i_8_163_1779_0, i_8_163_1786_0,
    i_8_163_1787_0, i_8_163_1805_0, i_8_163_1810_0, i_8_163_1819_0,
    i_8_163_1894_0, i_8_163_1963_0, i_8_163_1971_0, i_8_163_1975_0,
    i_8_163_1981_0, i_8_163_1983_0, i_8_163_1984_0, i_8_163_1994_0,
    i_8_163_2053_0, i_8_163_2056_0, i_8_163_2107_0, i_8_163_2108_0,
    i_8_163_2110_0, i_8_163_2134_0, i_8_163_2145_0, i_8_163_2146_0,
    i_8_163_2147_0, i_8_163_2148_0, i_8_163_2149_0, i_8_163_2155_0,
    i_8_163_2156_0, i_8_163_2158_0, i_8_163_2159_0, i_8_163_2169_0,
    i_8_163_2170_0, i_8_163_2223_0, i_8_163_2228_0, i_8_163_2229_0,
    i_8_163_2230_0, i_8_163_2234_0, i_8_163_2248_0, i_8_163_2263_0,
    o_8_163_0_0  );
  input  i_8_163_103_0, i_8_163_140_0, i_8_163_220_0, i_8_163_226_0,
    i_8_163_230_0, i_8_163_247_0, i_8_163_256_0, i_8_163_262_0,
    i_8_163_299_0, i_8_163_304_0, i_8_163_314_0, i_8_163_316_0,
    i_8_163_326_0, i_8_163_363_0, i_8_163_367_0, i_8_163_381_0,
    i_8_163_418_0, i_8_163_428_0, i_8_163_454_0, i_8_163_455_0,
    i_8_163_553_0, i_8_163_581_0, i_8_163_582_0, i_8_163_584_0,
    i_8_163_599_0, i_8_163_635_0, i_8_163_793_0, i_8_163_823_0,
    i_8_163_839_0, i_8_163_840_0, i_8_163_844_0, i_8_163_845_0,
    i_8_163_859_0, i_8_163_874_0, i_8_163_881_0, i_8_163_882_0,
    i_8_163_891_0, i_8_163_994_0, i_8_163_1145_0, i_8_163_1147_0,
    i_8_163_1226_0, i_8_163_1229_0, i_8_163_1268_0, i_8_163_1282_0,
    i_8_163_1286_0, i_8_163_1319_0, i_8_163_1399_0, i_8_163_1403_0,
    i_8_163_1432_0, i_8_163_1435_0, i_8_163_1436_0, i_8_163_1438_0,
    i_8_163_1463_0, i_8_163_1470_0, i_8_163_1510_0, i_8_163_1562_0,
    i_8_163_1574_0, i_8_163_1668_0, i_8_163_1688_0, i_8_163_1690_0,
    i_8_163_1704_0, i_8_163_1774_0, i_8_163_1779_0, i_8_163_1786_0,
    i_8_163_1787_0, i_8_163_1805_0, i_8_163_1810_0, i_8_163_1819_0,
    i_8_163_1894_0, i_8_163_1963_0, i_8_163_1971_0, i_8_163_1975_0,
    i_8_163_1981_0, i_8_163_1983_0, i_8_163_1984_0, i_8_163_1994_0,
    i_8_163_2053_0, i_8_163_2056_0, i_8_163_2107_0, i_8_163_2108_0,
    i_8_163_2110_0, i_8_163_2134_0, i_8_163_2145_0, i_8_163_2146_0,
    i_8_163_2147_0, i_8_163_2148_0, i_8_163_2149_0, i_8_163_2155_0,
    i_8_163_2156_0, i_8_163_2158_0, i_8_163_2159_0, i_8_163_2169_0,
    i_8_163_2170_0, i_8_163_2223_0, i_8_163_2228_0, i_8_163_2229_0,
    i_8_163_2230_0, i_8_163_2234_0, i_8_163_2248_0, i_8_163_2263_0;
  output o_8_163_0_0;
  assign o_8_163_0_0 = 0;
endmodule



// Benchmark "kernel_8_164" written by ABC on Sun Jul 19 10:05:52 2020

module kernel_8_164 ( 
    i_8_164_21_0, i_8_164_33_0, i_8_164_34_0, i_8_164_35_0, i_8_164_85_0,
    i_8_164_93_0, i_8_164_96_0, i_8_164_156_0, i_8_164_165_0,
    i_8_164_202_0, i_8_164_220_0, i_8_164_222_0, i_8_164_223_0,
    i_8_164_255_0, i_8_164_262_0, i_8_164_277_0, i_8_164_291_0,
    i_8_164_300_0, i_8_164_301_0, i_8_164_345_0, i_8_164_393_0,
    i_8_164_420_0, i_8_164_474_0, i_8_164_475_0, i_8_164_493_0,
    i_8_164_500_0, i_8_164_501_0, i_8_164_503_0, i_8_164_547_0,
    i_8_164_552_0, i_8_164_555_0, i_8_164_588_0, i_8_164_589_0,
    i_8_164_624_0, i_8_164_657_0, i_8_164_670_0, i_8_164_715_0,
    i_8_164_716_0, i_8_164_723_0, i_8_164_759_0, i_8_164_768_0,
    i_8_164_781_0, i_8_164_823_0, i_8_164_877_0, i_8_164_1011_0,
    i_8_164_1029_0, i_8_164_1114_0, i_8_164_1115_0, i_8_164_1119_0,
    i_8_164_1128_0, i_8_164_1156_0, i_8_164_1159_0, i_8_164_1191_0,
    i_8_164_1254_0, i_8_164_1257_0, i_8_164_1258_0, i_8_164_1282_0,
    i_8_164_1344_0, i_8_164_1345_0, i_8_164_1347_0, i_8_164_1452_0,
    i_8_164_1453_0, i_8_164_1542_0, i_8_164_1551_0, i_8_164_1555_0,
    i_8_164_1587_0, i_8_164_1596_0, i_8_164_1597_0, i_8_164_1600_0,
    i_8_164_1611_0, i_8_164_1626_0, i_8_164_1651_0, i_8_164_1668_0,
    i_8_164_1680_0, i_8_164_1682_0, i_8_164_1708_0, i_8_164_1743_0,
    i_8_164_1760_0, i_8_164_1761_0, i_8_164_1762_0, i_8_164_1782_0,
    i_8_164_1804_0, i_8_164_1806_0, i_8_164_1839_0, i_8_164_1849_0,
    i_8_164_1867_0, i_8_164_1893_0, i_8_164_1894_0, i_8_164_1952_0,
    i_8_164_1992_0, i_8_164_1995_0, i_8_164_2031_0, i_8_164_2049_0,
    i_8_164_2110_0, i_8_164_2128_0, i_8_164_2190_0, i_8_164_2214_0,
    i_8_164_2215_0, i_8_164_2287_0, i_8_164_2289_0,
    o_8_164_0_0  );
  input  i_8_164_21_0, i_8_164_33_0, i_8_164_34_0, i_8_164_35_0,
    i_8_164_85_0, i_8_164_93_0, i_8_164_96_0, i_8_164_156_0, i_8_164_165_0,
    i_8_164_202_0, i_8_164_220_0, i_8_164_222_0, i_8_164_223_0,
    i_8_164_255_0, i_8_164_262_0, i_8_164_277_0, i_8_164_291_0,
    i_8_164_300_0, i_8_164_301_0, i_8_164_345_0, i_8_164_393_0,
    i_8_164_420_0, i_8_164_474_0, i_8_164_475_0, i_8_164_493_0,
    i_8_164_500_0, i_8_164_501_0, i_8_164_503_0, i_8_164_547_0,
    i_8_164_552_0, i_8_164_555_0, i_8_164_588_0, i_8_164_589_0,
    i_8_164_624_0, i_8_164_657_0, i_8_164_670_0, i_8_164_715_0,
    i_8_164_716_0, i_8_164_723_0, i_8_164_759_0, i_8_164_768_0,
    i_8_164_781_0, i_8_164_823_0, i_8_164_877_0, i_8_164_1011_0,
    i_8_164_1029_0, i_8_164_1114_0, i_8_164_1115_0, i_8_164_1119_0,
    i_8_164_1128_0, i_8_164_1156_0, i_8_164_1159_0, i_8_164_1191_0,
    i_8_164_1254_0, i_8_164_1257_0, i_8_164_1258_0, i_8_164_1282_0,
    i_8_164_1344_0, i_8_164_1345_0, i_8_164_1347_0, i_8_164_1452_0,
    i_8_164_1453_0, i_8_164_1542_0, i_8_164_1551_0, i_8_164_1555_0,
    i_8_164_1587_0, i_8_164_1596_0, i_8_164_1597_0, i_8_164_1600_0,
    i_8_164_1611_0, i_8_164_1626_0, i_8_164_1651_0, i_8_164_1668_0,
    i_8_164_1680_0, i_8_164_1682_0, i_8_164_1708_0, i_8_164_1743_0,
    i_8_164_1760_0, i_8_164_1761_0, i_8_164_1762_0, i_8_164_1782_0,
    i_8_164_1804_0, i_8_164_1806_0, i_8_164_1839_0, i_8_164_1849_0,
    i_8_164_1867_0, i_8_164_1893_0, i_8_164_1894_0, i_8_164_1952_0,
    i_8_164_1992_0, i_8_164_1995_0, i_8_164_2031_0, i_8_164_2049_0,
    i_8_164_2110_0, i_8_164_2128_0, i_8_164_2190_0, i_8_164_2214_0,
    i_8_164_2215_0, i_8_164_2287_0, i_8_164_2289_0;
  output o_8_164_0_0;
  assign o_8_164_0_0 = 0;
endmodule



// Benchmark "kernel_8_165" written by ABC on Sun Jul 19 10:05:53 2020

module kernel_8_165 ( 
    i_8_165_20_0, i_8_165_38_0, i_8_165_44_0, i_8_165_106_0, i_8_165_184_0,
    i_8_165_214_0, i_8_165_226_0, i_8_165_257_0, i_8_165_263_0,
    i_8_165_270_0, i_8_165_288_0, i_8_165_289_0, i_8_165_297_0,
    i_8_165_344_0, i_8_165_353_0, i_8_165_370_0, i_8_165_380_0,
    i_8_165_388_0, i_8_165_416_0, i_8_165_443_0, i_8_165_452_0,
    i_8_165_462_0, i_8_165_475_0, i_8_165_535_0, i_8_165_625_0,
    i_8_165_627_0, i_8_165_638_0, i_8_165_661_0, i_8_165_663_0,
    i_8_165_665_0, i_8_165_695_0, i_8_165_696_0, i_8_165_713_0,
    i_8_165_724_0, i_8_165_756_0, i_8_165_759_0, i_8_165_792_0,
    i_8_165_793_0, i_8_165_817_0, i_8_165_869_0, i_8_165_875_0,
    i_8_165_876_0, i_8_165_927_0, i_8_165_971_0, i_8_165_982_0,
    i_8_165_988_0, i_8_165_992_0, i_8_165_999_0, i_8_165_1051_0,
    i_8_165_1110_0, i_8_165_1127_0, i_8_165_1156_0, i_8_165_1161_0,
    i_8_165_1217_0, i_8_165_1224_0, i_8_165_1236_0, i_8_165_1246_0,
    i_8_165_1252_0, i_8_165_1271_0, i_8_165_1281_0, i_8_165_1300_0,
    i_8_165_1341_0, i_8_165_1363_0, i_8_165_1367_0, i_8_165_1424_0,
    i_8_165_1427_0, i_8_165_1453_0, i_8_165_1469_0, i_8_165_1504_0,
    i_8_165_1560_0, i_8_165_1603_0, i_8_165_1604_0, i_8_165_1613_0,
    i_8_165_1631_0, i_8_165_1674_0, i_8_165_1687_0, i_8_165_1699_0,
    i_8_165_1714_0, i_8_165_1733_0, i_8_165_1750_0, i_8_165_1758_0,
    i_8_165_1762_0, i_8_165_1780_0, i_8_165_1791_0, i_8_165_1807_0,
    i_8_165_1838_0, i_8_165_1854_0, i_8_165_1920_0, i_8_165_1996_0,
    i_8_165_2018_0, i_8_165_2054_0, i_8_165_2056_0, i_8_165_2124_0,
    i_8_165_2129_0, i_8_165_2170_0, i_8_165_2171_0, i_8_165_2188_0,
    i_8_165_2223_0, i_8_165_2261_0, i_8_165_2270_0,
    o_8_165_0_0  );
  input  i_8_165_20_0, i_8_165_38_0, i_8_165_44_0, i_8_165_106_0,
    i_8_165_184_0, i_8_165_214_0, i_8_165_226_0, i_8_165_257_0,
    i_8_165_263_0, i_8_165_270_0, i_8_165_288_0, i_8_165_289_0,
    i_8_165_297_0, i_8_165_344_0, i_8_165_353_0, i_8_165_370_0,
    i_8_165_380_0, i_8_165_388_0, i_8_165_416_0, i_8_165_443_0,
    i_8_165_452_0, i_8_165_462_0, i_8_165_475_0, i_8_165_535_0,
    i_8_165_625_0, i_8_165_627_0, i_8_165_638_0, i_8_165_661_0,
    i_8_165_663_0, i_8_165_665_0, i_8_165_695_0, i_8_165_696_0,
    i_8_165_713_0, i_8_165_724_0, i_8_165_756_0, i_8_165_759_0,
    i_8_165_792_0, i_8_165_793_0, i_8_165_817_0, i_8_165_869_0,
    i_8_165_875_0, i_8_165_876_0, i_8_165_927_0, i_8_165_971_0,
    i_8_165_982_0, i_8_165_988_0, i_8_165_992_0, i_8_165_999_0,
    i_8_165_1051_0, i_8_165_1110_0, i_8_165_1127_0, i_8_165_1156_0,
    i_8_165_1161_0, i_8_165_1217_0, i_8_165_1224_0, i_8_165_1236_0,
    i_8_165_1246_0, i_8_165_1252_0, i_8_165_1271_0, i_8_165_1281_0,
    i_8_165_1300_0, i_8_165_1341_0, i_8_165_1363_0, i_8_165_1367_0,
    i_8_165_1424_0, i_8_165_1427_0, i_8_165_1453_0, i_8_165_1469_0,
    i_8_165_1504_0, i_8_165_1560_0, i_8_165_1603_0, i_8_165_1604_0,
    i_8_165_1613_0, i_8_165_1631_0, i_8_165_1674_0, i_8_165_1687_0,
    i_8_165_1699_0, i_8_165_1714_0, i_8_165_1733_0, i_8_165_1750_0,
    i_8_165_1758_0, i_8_165_1762_0, i_8_165_1780_0, i_8_165_1791_0,
    i_8_165_1807_0, i_8_165_1838_0, i_8_165_1854_0, i_8_165_1920_0,
    i_8_165_1996_0, i_8_165_2018_0, i_8_165_2054_0, i_8_165_2056_0,
    i_8_165_2124_0, i_8_165_2129_0, i_8_165_2170_0, i_8_165_2171_0,
    i_8_165_2188_0, i_8_165_2223_0, i_8_165_2261_0, i_8_165_2270_0;
  output o_8_165_0_0;
  assign o_8_165_0_0 = 0;
endmodule



// Benchmark "kernel_8_166" written by ABC on Sun Jul 19 10:05:54 2020

module kernel_8_166 ( 
    i_8_166_13_0, i_8_166_28_0, i_8_166_44_0, i_8_166_79_0, i_8_166_80_0,
    i_8_166_106_0, i_8_166_115_0, i_8_166_140_0, i_8_166_185_0,
    i_8_166_227_0, i_8_166_320_0, i_8_166_322_0, i_8_166_323_0,
    i_8_166_349_0, i_8_166_391_0, i_8_166_401_0, i_8_166_421_0,
    i_8_166_431_0, i_8_166_455_0, i_8_166_486_0, i_8_166_500_0,
    i_8_166_536_0, i_8_166_556_0, i_8_166_557_0, i_8_166_572_0,
    i_8_166_607_0, i_8_166_623_0, i_8_166_635_0, i_8_166_653_0,
    i_8_166_655_0, i_8_166_656_0, i_8_166_670_0, i_8_166_674_0,
    i_8_166_702_0, i_8_166_703_0, i_8_166_826_0, i_8_166_827_0,
    i_8_166_838_0, i_8_166_839_0, i_8_166_877_0, i_8_166_881_0,
    i_8_166_896_0, i_8_166_956_0, i_8_166_970_0, i_8_166_971_0,
    i_8_166_991_0, i_8_166_1055_0, i_8_166_1111_0, i_8_166_1154_0,
    i_8_166_1202_0, i_8_166_1300_0, i_8_166_1301_0, i_8_166_1331_0,
    i_8_166_1336_0, i_8_166_1337_0, i_8_166_1366_0, i_8_166_1367_0,
    i_8_166_1400_0, i_8_166_1402_0, i_8_166_1435_0, i_8_166_1465_0,
    i_8_166_1474_0, i_8_166_1489_0, i_8_166_1493_0, i_8_166_1510_0,
    i_8_166_1517_0, i_8_166_1525_0, i_8_166_1526_0, i_8_166_1529_0,
    i_8_166_1548_0, i_8_166_1550_0, i_8_166_1553_0, i_8_166_1574_0,
    i_8_166_1622_0, i_8_166_1625_0, i_8_166_1630_0, i_8_166_1634_0,
    i_8_166_1651_0, i_8_166_1672_0, i_8_166_1753_0, i_8_166_1771_0,
    i_8_166_1774_0, i_8_166_1784_0, i_8_166_1795_0, i_8_166_1824_0,
    i_8_166_1825_0, i_8_166_1849_0, i_8_166_1886_0, i_8_166_1888_0,
    i_8_166_1937_0, i_8_166_1960_0, i_8_166_1968_0, i_8_166_1975_0,
    i_8_166_1995_0, i_8_166_2057_0, i_8_166_2072_0, i_8_166_2125_0,
    i_8_166_2146_0, i_8_166_2242_0, i_8_166_2285_0,
    o_8_166_0_0  );
  input  i_8_166_13_0, i_8_166_28_0, i_8_166_44_0, i_8_166_79_0,
    i_8_166_80_0, i_8_166_106_0, i_8_166_115_0, i_8_166_140_0,
    i_8_166_185_0, i_8_166_227_0, i_8_166_320_0, i_8_166_322_0,
    i_8_166_323_0, i_8_166_349_0, i_8_166_391_0, i_8_166_401_0,
    i_8_166_421_0, i_8_166_431_0, i_8_166_455_0, i_8_166_486_0,
    i_8_166_500_0, i_8_166_536_0, i_8_166_556_0, i_8_166_557_0,
    i_8_166_572_0, i_8_166_607_0, i_8_166_623_0, i_8_166_635_0,
    i_8_166_653_0, i_8_166_655_0, i_8_166_656_0, i_8_166_670_0,
    i_8_166_674_0, i_8_166_702_0, i_8_166_703_0, i_8_166_826_0,
    i_8_166_827_0, i_8_166_838_0, i_8_166_839_0, i_8_166_877_0,
    i_8_166_881_0, i_8_166_896_0, i_8_166_956_0, i_8_166_970_0,
    i_8_166_971_0, i_8_166_991_0, i_8_166_1055_0, i_8_166_1111_0,
    i_8_166_1154_0, i_8_166_1202_0, i_8_166_1300_0, i_8_166_1301_0,
    i_8_166_1331_0, i_8_166_1336_0, i_8_166_1337_0, i_8_166_1366_0,
    i_8_166_1367_0, i_8_166_1400_0, i_8_166_1402_0, i_8_166_1435_0,
    i_8_166_1465_0, i_8_166_1474_0, i_8_166_1489_0, i_8_166_1493_0,
    i_8_166_1510_0, i_8_166_1517_0, i_8_166_1525_0, i_8_166_1526_0,
    i_8_166_1529_0, i_8_166_1548_0, i_8_166_1550_0, i_8_166_1553_0,
    i_8_166_1574_0, i_8_166_1622_0, i_8_166_1625_0, i_8_166_1630_0,
    i_8_166_1634_0, i_8_166_1651_0, i_8_166_1672_0, i_8_166_1753_0,
    i_8_166_1771_0, i_8_166_1774_0, i_8_166_1784_0, i_8_166_1795_0,
    i_8_166_1824_0, i_8_166_1825_0, i_8_166_1849_0, i_8_166_1886_0,
    i_8_166_1888_0, i_8_166_1937_0, i_8_166_1960_0, i_8_166_1968_0,
    i_8_166_1975_0, i_8_166_1995_0, i_8_166_2057_0, i_8_166_2072_0,
    i_8_166_2125_0, i_8_166_2146_0, i_8_166_2242_0, i_8_166_2285_0;
  output o_8_166_0_0;
  assign o_8_166_0_0 = 0;
endmodule



// Benchmark "kernel_8_167" written by ABC on Sun Jul 19 10:05:55 2020

module kernel_8_167 ( 
    i_8_167_76_0, i_8_167_115_0, i_8_167_137_0, i_8_167_184_0,
    i_8_167_279_0, i_8_167_299_0, i_8_167_320_0, i_8_167_322_0,
    i_8_167_392_0, i_8_167_423_0, i_8_167_427_0, i_8_167_429_0,
    i_8_167_483_0, i_8_167_487_0, i_8_167_489_0, i_8_167_496_0,
    i_8_167_553_0, i_8_167_574_0, i_8_167_580_0, i_8_167_581_0,
    i_8_167_588_0, i_8_167_606_0, i_8_167_607_0, i_8_167_630_0,
    i_8_167_633_0, i_8_167_640_0, i_8_167_641_0, i_8_167_651_0,
    i_8_167_655_0, i_8_167_661_0, i_8_167_676_0, i_8_167_703_0,
    i_8_167_706_0, i_8_167_742_0, i_8_167_744_0, i_8_167_755_0,
    i_8_167_841_0, i_8_167_842_0, i_8_167_895_0, i_8_167_971_0,
    i_8_167_973_0, i_8_167_974_0, i_8_167_1010_0, i_8_167_1020_0,
    i_8_167_1036_0, i_8_167_1039_0, i_8_167_1107_0, i_8_167_1109_0,
    i_8_167_1200_0, i_8_167_1201_0, i_8_167_1246_0, i_8_167_1247_0,
    i_8_167_1264_0, i_8_167_1267_0, i_8_167_1297_0, i_8_167_1315_0,
    i_8_167_1351_0, i_8_167_1363_0, i_8_167_1365_0, i_8_167_1382_0,
    i_8_167_1383_0, i_8_167_1416_0, i_8_167_1434_0, i_8_167_1435_0,
    i_8_167_1436_0, i_8_167_1438_0, i_8_167_1461_0, i_8_167_1462_0,
    i_8_167_1465_0, i_8_167_1469_0, i_8_167_1477_0, i_8_167_1487_0,
    i_8_167_1512_0, i_8_167_1547_0, i_8_167_1607_0, i_8_167_1630_0,
    i_8_167_1638_0, i_8_167_1707_0, i_8_167_1720_0, i_8_167_1802_0,
    i_8_167_1809_0, i_8_167_1825_0, i_8_167_1837_0, i_8_167_1838_0,
    i_8_167_1840_0, i_8_167_1912_0, i_8_167_1957_0, i_8_167_1981_0,
    i_8_167_1992_0, i_8_167_1994_0, i_8_167_1997_0, i_8_167_2119_0,
    i_8_167_2146_0, i_8_167_2147_0, i_8_167_2169_0, i_8_167_2170_0,
    i_8_167_2227_0, i_8_167_2247_0, i_8_167_2248_0, i_8_167_2289_0,
    o_8_167_0_0  );
  input  i_8_167_76_0, i_8_167_115_0, i_8_167_137_0, i_8_167_184_0,
    i_8_167_279_0, i_8_167_299_0, i_8_167_320_0, i_8_167_322_0,
    i_8_167_392_0, i_8_167_423_0, i_8_167_427_0, i_8_167_429_0,
    i_8_167_483_0, i_8_167_487_0, i_8_167_489_0, i_8_167_496_0,
    i_8_167_553_0, i_8_167_574_0, i_8_167_580_0, i_8_167_581_0,
    i_8_167_588_0, i_8_167_606_0, i_8_167_607_0, i_8_167_630_0,
    i_8_167_633_0, i_8_167_640_0, i_8_167_641_0, i_8_167_651_0,
    i_8_167_655_0, i_8_167_661_0, i_8_167_676_0, i_8_167_703_0,
    i_8_167_706_0, i_8_167_742_0, i_8_167_744_0, i_8_167_755_0,
    i_8_167_841_0, i_8_167_842_0, i_8_167_895_0, i_8_167_971_0,
    i_8_167_973_0, i_8_167_974_0, i_8_167_1010_0, i_8_167_1020_0,
    i_8_167_1036_0, i_8_167_1039_0, i_8_167_1107_0, i_8_167_1109_0,
    i_8_167_1200_0, i_8_167_1201_0, i_8_167_1246_0, i_8_167_1247_0,
    i_8_167_1264_0, i_8_167_1267_0, i_8_167_1297_0, i_8_167_1315_0,
    i_8_167_1351_0, i_8_167_1363_0, i_8_167_1365_0, i_8_167_1382_0,
    i_8_167_1383_0, i_8_167_1416_0, i_8_167_1434_0, i_8_167_1435_0,
    i_8_167_1436_0, i_8_167_1438_0, i_8_167_1461_0, i_8_167_1462_0,
    i_8_167_1465_0, i_8_167_1469_0, i_8_167_1477_0, i_8_167_1487_0,
    i_8_167_1512_0, i_8_167_1547_0, i_8_167_1607_0, i_8_167_1630_0,
    i_8_167_1638_0, i_8_167_1707_0, i_8_167_1720_0, i_8_167_1802_0,
    i_8_167_1809_0, i_8_167_1825_0, i_8_167_1837_0, i_8_167_1838_0,
    i_8_167_1840_0, i_8_167_1912_0, i_8_167_1957_0, i_8_167_1981_0,
    i_8_167_1992_0, i_8_167_1994_0, i_8_167_1997_0, i_8_167_2119_0,
    i_8_167_2146_0, i_8_167_2147_0, i_8_167_2169_0, i_8_167_2170_0,
    i_8_167_2227_0, i_8_167_2247_0, i_8_167_2248_0, i_8_167_2289_0;
  output o_8_167_0_0;
  assign o_8_167_0_0 = 0;
endmodule



// Benchmark "kernel_8_168" written by ABC on Sun Jul 19 10:05:56 2020

module kernel_8_168 ( 
    i_8_168_19_0, i_8_168_20_0, i_8_168_58_0, i_8_168_78_0, i_8_168_79_0,
    i_8_168_94_0, i_8_168_114_0, i_8_168_289_0, i_8_168_298_0,
    i_8_168_325_0, i_8_168_353_0, i_8_168_360_0, i_8_168_370_0,
    i_8_168_383_0, i_8_168_417_0, i_8_168_459_0, i_8_168_460_0,
    i_8_168_461_0, i_8_168_482_0, i_8_168_490_0, i_8_168_526_0,
    i_8_168_549_0, i_8_168_553_0, i_8_168_615_0, i_8_168_621_0,
    i_8_168_622_0, i_8_168_623_0, i_8_168_627_0, i_8_168_628_0,
    i_8_168_629_0, i_8_168_661_0, i_8_168_667_0, i_8_168_696_0,
    i_8_168_703_0, i_8_168_712_0, i_8_168_779_0, i_8_168_792_0,
    i_8_168_830_0, i_8_168_832_0, i_8_168_841_0, i_8_168_885_0,
    i_8_168_938_0, i_8_168_971_0, i_8_168_977_0, i_8_168_990_0,
    i_8_168_992_0, i_8_168_997_0, i_8_168_1010_0, i_8_168_1110_0,
    i_8_168_1118_0, i_8_168_1127_0, i_8_168_1128_0, i_8_168_1225_0,
    i_8_168_1234_0, i_8_168_1278_0, i_8_168_1280_0, i_8_168_1316_0,
    i_8_168_1324_0, i_8_168_1341_0, i_8_168_1408_0, i_8_168_1411_0,
    i_8_168_1449_0, i_8_168_1450_0, i_8_168_1451_0, i_8_168_1504_0,
    i_8_168_1532_0, i_8_168_1533_0, i_8_168_1548_0, i_8_168_1549_0,
    i_8_168_1553_0, i_8_168_1594_0, i_8_168_1650_0, i_8_168_1749_0,
    i_8_168_1750_0, i_8_168_1758_0, i_8_168_1759_0, i_8_168_1775_0,
    i_8_168_1801_0, i_8_168_1838_0, i_8_168_1864_0, i_8_168_1865_0,
    i_8_168_1891_0, i_8_168_1909_0, i_8_168_1919_0, i_8_168_1963_0,
    i_8_168_1967_0, i_8_168_1985_0, i_8_168_1990_0, i_8_168_2106_0,
    i_8_168_2107_0, i_8_168_2126_0, i_8_168_2141_0, i_8_168_2142_0,
    i_8_168_2188_0, i_8_168_2224_0, i_8_168_2269_0, i_8_168_2270_0,
    i_8_168_2273_0, i_8_168_2286_0, i_8_168_2288_0,
    o_8_168_0_0  );
  input  i_8_168_19_0, i_8_168_20_0, i_8_168_58_0, i_8_168_78_0,
    i_8_168_79_0, i_8_168_94_0, i_8_168_114_0, i_8_168_289_0,
    i_8_168_298_0, i_8_168_325_0, i_8_168_353_0, i_8_168_360_0,
    i_8_168_370_0, i_8_168_383_0, i_8_168_417_0, i_8_168_459_0,
    i_8_168_460_0, i_8_168_461_0, i_8_168_482_0, i_8_168_490_0,
    i_8_168_526_0, i_8_168_549_0, i_8_168_553_0, i_8_168_615_0,
    i_8_168_621_0, i_8_168_622_0, i_8_168_623_0, i_8_168_627_0,
    i_8_168_628_0, i_8_168_629_0, i_8_168_661_0, i_8_168_667_0,
    i_8_168_696_0, i_8_168_703_0, i_8_168_712_0, i_8_168_779_0,
    i_8_168_792_0, i_8_168_830_0, i_8_168_832_0, i_8_168_841_0,
    i_8_168_885_0, i_8_168_938_0, i_8_168_971_0, i_8_168_977_0,
    i_8_168_990_0, i_8_168_992_0, i_8_168_997_0, i_8_168_1010_0,
    i_8_168_1110_0, i_8_168_1118_0, i_8_168_1127_0, i_8_168_1128_0,
    i_8_168_1225_0, i_8_168_1234_0, i_8_168_1278_0, i_8_168_1280_0,
    i_8_168_1316_0, i_8_168_1324_0, i_8_168_1341_0, i_8_168_1408_0,
    i_8_168_1411_0, i_8_168_1449_0, i_8_168_1450_0, i_8_168_1451_0,
    i_8_168_1504_0, i_8_168_1532_0, i_8_168_1533_0, i_8_168_1548_0,
    i_8_168_1549_0, i_8_168_1553_0, i_8_168_1594_0, i_8_168_1650_0,
    i_8_168_1749_0, i_8_168_1750_0, i_8_168_1758_0, i_8_168_1759_0,
    i_8_168_1775_0, i_8_168_1801_0, i_8_168_1838_0, i_8_168_1864_0,
    i_8_168_1865_0, i_8_168_1891_0, i_8_168_1909_0, i_8_168_1919_0,
    i_8_168_1963_0, i_8_168_1967_0, i_8_168_1985_0, i_8_168_1990_0,
    i_8_168_2106_0, i_8_168_2107_0, i_8_168_2126_0, i_8_168_2141_0,
    i_8_168_2142_0, i_8_168_2188_0, i_8_168_2224_0, i_8_168_2269_0,
    i_8_168_2270_0, i_8_168_2273_0, i_8_168_2286_0, i_8_168_2288_0;
  output o_8_168_0_0;
  assign o_8_168_0_0 = 0;
endmodule



// Benchmark "kernel_8_169" written by ABC on Sun Jul 19 10:05:57 2020

module kernel_8_169 ( 
    i_8_169_10_0, i_8_169_80_0, i_8_169_226_0, i_8_169_230_0,
    i_8_169_233_0, i_8_169_260_0, i_8_169_298_0, i_8_169_301_0,
    i_8_169_314_0, i_8_169_316_0, i_8_169_367_0, i_8_169_419_0,
    i_8_169_469_0, i_8_169_526_0, i_8_169_530_0, i_8_169_604_0,
    i_8_169_605_0, i_8_169_607_0, i_8_169_616_0, i_8_169_629_0,
    i_8_169_649_0, i_8_169_657_0, i_8_169_665_0, i_8_169_691_0,
    i_8_169_692_0, i_8_169_696_0, i_8_169_697_0, i_8_169_700_0,
    i_8_169_701_0, i_8_169_705_0, i_8_169_709_0, i_8_169_836_0,
    i_8_169_843_0, i_8_169_844_0, i_8_169_855_0, i_8_169_863_0,
    i_8_169_881_0, i_8_169_890_0, i_8_169_976_0, i_8_169_988_0,
    i_8_169_989_0, i_8_169_994_0, i_8_169_1006_0, i_8_169_1043_0,
    i_8_169_1052_0, i_8_169_1060_0, i_8_169_1097_0, i_8_169_1105_0,
    i_8_169_1150_0, i_8_169_1168_0, i_8_169_1219_0, i_8_169_1297_0,
    i_8_169_1325_0, i_8_169_1351_0, i_8_169_1411_0, i_8_169_1434_0,
    i_8_169_1462_0, i_8_169_1492_0, i_8_169_1504_0, i_8_169_1544_0,
    i_8_169_1551_0, i_8_169_1555_0, i_8_169_1565_0, i_8_169_1567_0,
    i_8_169_1609_0, i_8_169_1627_0, i_8_169_1628_0, i_8_169_1652_0,
    i_8_169_1663_0, i_8_169_1669_0, i_8_169_1674_0, i_8_169_1693_0,
    i_8_169_1709_0, i_8_169_1766_0, i_8_169_1780_0, i_8_169_1792_0,
    i_8_169_1798_0, i_8_169_1826_0, i_8_169_1837_0, i_8_169_1855_0,
    i_8_169_1858_0, i_8_169_1867_0, i_8_169_1880_0, i_8_169_1885_0,
    i_8_169_1888_0, i_8_169_1894_0, i_8_169_1897_0, i_8_169_1954_0,
    i_8_169_1990_0, i_8_169_2015_0, i_8_169_2071_0, i_8_169_2077_0,
    i_8_169_2078_0, i_8_169_2093_0, i_8_169_2095_0, i_8_169_2105_0,
    i_8_169_2136_0, i_8_169_2170_0, i_8_169_2259_0, i_8_169_2275_0,
    o_8_169_0_0  );
  input  i_8_169_10_0, i_8_169_80_0, i_8_169_226_0, i_8_169_230_0,
    i_8_169_233_0, i_8_169_260_0, i_8_169_298_0, i_8_169_301_0,
    i_8_169_314_0, i_8_169_316_0, i_8_169_367_0, i_8_169_419_0,
    i_8_169_469_0, i_8_169_526_0, i_8_169_530_0, i_8_169_604_0,
    i_8_169_605_0, i_8_169_607_0, i_8_169_616_0, i_8_169_629_0,
    i_8_169_649_0, i_8_169_657_0, i_8_169_665_0, i_8_169_691_0,
    i_8_169_692_0, i_8_169_696_0, i_8_169_697_0, i_8_169_700_0,
    i_8_169_701_0, i_8_169_705_0, i_8_169_709_0, i_8_169_836_0,
    i_8_169_843_0, i_8_169_844_0, i_8_169_855_0, i_8_169_863_0,
    i_8_169_881_0, i_8_169_890_0, i_8_169_976_0, i_8_169_988_0,
    i_8_169_989_0, i_8_169_994_0, i_8_169_1006_0, i_8_169_1043_0,
    i_8_169_1052_0, i_8_169_1060_0, i_8_169_1097_0, i_8_169_1105_0,
    i_8_169_1150_0, i_8_169_1168_0, i_8_169_1219_0, i_8_169_1297_0,
    i_8_169_1325_0, i_8_169_1351_0, i_8_169_1411_0, i_8_169_1434_0,
    i_8_169_1462_0, i_8_169_1492_0, i_8_169_1504_0, i_8_169_1544_0,
    i_8_169_1551_0, i_8_169_1555_0, i_8_169_1565_0, i_8_169_1567_0,
    i_8_169_1609_0, i_8_169_1627_0, i_8_169_1628_0, i_8_169_1652_0,
    i_8_169_1663_0, i_8_169_1669_0, i_8_169_1674_0, i_8_169_1693_0,
    i_8_169_1709_0, i_8_169_1766_0, i_8_169_1780_0, i_8_169_1792_0,
    i_8_169_1798_0, i_8_169_1826_0, i_8_169_1837_0, i_8_169_1855_0,
    i_8_169_1858_0, i_8_169_1867_0, i_8_169_1880_0, i_8_169_1885_0,
    i_8_169_1888_0, i_8_169_1894_0, i_8_169_1897_0, i_8_169_1954_0,
    i_8_169_1990_0, i_8_169_2015_0, i_8_169_2071_0, i_8_169_2077_0,
    i_8_169_2078_0, i_8_169_2093_0, i_8_169_2095_0, i_8_169_2105_0,
    i_8_169_2136_0, i_8_169_2170_0, i_8_169_2259_0, i_8_169_2275_0;
  output o_8_169_0_0;
  assign o_8_169_0_0 = 0;
endmodule



// Benchmark "kernel_8_170" written by ABC on Sun Jul 19 10:05:58 2020

module kernel_8_170 ( 
    i_8_170_3_0, i_8_170_6_0, i_8_170_9_0, i_8_170_54_0, i_8_170_115_0,
    i_8_170_210_0, i_8_170_219_0, i_8_170_249_0, i_8_170_258_0,
    i_8_170_295_0, i_8_170_298_0, i_8_170_350_0, i_8_170_358_0,
    i_8_170_363_0, i_8_170_365_0, i_8_170_421_0, i_8_170_448_0,
    i_8_170_454_0, i_8_170_466_0, i_8_170_490_0, i_8_170_516_0,
    i_8_170_523_0, i_8_170_574_0, i_8_170_598_0, i_8_170_601_0,
    i_8_170_606_0, i_8_170_607_0, i_8_170_610_0, i_8_170_661_0,
    i_8_170_672_0, i_8_170_699_0, i_8_170_717_0, i_8_170_718_0,
    i_8_170_726_0, i_8_170_736_0, i_8_170_789_0, i_8_170_813_0,
    i_8_170_816_0, i_8_170_817_0, i_8_170_835_0, i_8_170_836_0,
    i_8_170_842_0, i_8_170_852_0, i_8_170_853_0, i_8_170_889_0,
    i_8_170_1015_0, i_8_170_1029_0, i_8_170_1031_0, i_8_170_1044_0,
    i_8_170_1074_0, i_8_170_1078_0, i_8_170_1087_0, i_8_170_1156_0,
    i_8_170_1204_0, i_8_170_1285_0, i_8_170_1308_0, i_8_170_1317_0,
    i_8_170_1392_0, i_8_170_1393_0, i_8_170_1394_0, i_8_170_1437_0,
    i_8_170_1446_0, i_8_170_1500_0, i_8_170_1636_0, i_8_170_1662_0,
    i_8_170_1695_0, i_8_170_1699_0, i_8_170_1763_0, i_8_170_1798_0,
    i_8_170_1808_0, i_8_170_1824_0, i_8_170_1848_0, i_8_170_1851_0,
    i_8_170_1858_0, i_8_170_1866_0, i_8_170_1870_0, i_8_170_1879_0,
    i_8_170_1881_0, i_8_170_1897_0, i_8_170_1920_0, i_8_170_2031_0,
    i_8_170_2059_0, i_8_170_2067_0, i_8_170_2068_0, i_8_170_2073_0,
    i_8_170_2074_0, i_8_170_2076_0, i_8_170_2077_0, i_8_170_2092_0,
    i_8_170_2112_0, i_8_170_2118_0, i_8_170_2121_0, i_8_170_2122_0,
    i_8_170_2154_0, i_8_170_2215_0, i_8_170_2235_0, i_8_170_2246_0,
    i_8_170_2283_0, i_8_170_2284_0, i_8_170_2293_0,
    o_8_170_0_0  );
  input  i_8_170_3_0, i_8_170_6_0, i_8_170_9_0, i_8_170_54_0,
    i_8_170_115_0, i_8_170_210_0, i_8_170_219_0, i_8_170_249_0,
    i_8_170_258_0, i_8_170_295_0, i_8_170_298_0, i_8_170_350_0,
    i_8_170_358_0, i_8_170_363_0, i_8_170_365_0, i_8_170_421_0,
    i_8_170_448_0, i_8_170_454_0, i_8_170_466_0, i_8_170_490_0,
    i_8_170_516_0, i_8_170_523_0, i_8_170_574_0, i_8_170_598_0,
    i_8_170_601_0, i_8_170_606_0, i_8_170_607_0, i_8_170_610_0,
    i_8_170_661_0, i_8_170_672_0, i_8_170_699_0, i_8_170_717_0,
    i_8_170_718_0, i_8_170_726_0, i_8_170_736_0, i_8_170_789_0,
    i_8_170_813_0, i_8_170_816_0, i_8_170_817_0, i_8_170_835_0,
    i_8_170_836_0, i_8_170_842_0, i_8_170_852_0, i_8_170_853_0,
    i_8_170_889_0, i_8_170_1015_0, i_8_170_1029_0, i_8_170_1031_0,
    i_8_170_1044_0, i_8_170_1074_0, i_8_170_1078_0, i_8_170_1087_0,
    i_8_170_1156_0, i_8_170_1204_0, i_8_170_1285_0, i_8_170_1308_0,
    i_8_170_1317_0, i_8_170_1392_0, i_8_170_1393_0, i_8_170_1394_0,
    i_8_170_1437_0, i_8_170_1446_0, i_8_170_1500_0, i_8_170_1636_0,
    i_8_170_1662_0, i_8_170_1695_0, i_8_170_1699_0, i_8_170_1763_0,
    i_8_170_1798_0, i_8_170_1808_0, i_8_170_1824_0, i_8_170_1848_0,
    i_8_170_1851_0, i_8_170_1858_0, i_8_170_1866_0, i_8_170_1870_0,
    i_8_170_1879_0, i_8_170_1881_0, i_8_170_1897_0, i_8_170_1920_0,
    i_8_170_2031_0, i_8_170_2059_0, i_8_170_2067_0, i_8_170_2068_0,
    i_8_170_2073_0, i_8_170_2074_0, i_8_170_2076_0, i_8_170_2077_0,
    i_8_170_2092_0, i_8_170_2112_0, i_8_170_2118_0, i_8_170_2121_0,
    i_8_170_2122_0, i_8_170_2154_0, i_8_170_2215_0, i_8_170_2235_0,
    i_8_170_2246_0, i_8_170_2283_0, i_8_170_2284_0, i_8_170_2293_0;
  output o_8_170_0_0;
  assign o_8_170_0_0 = ~((~i_8_170_298_0 & ((~i_8_170_448_0 & ~i_8_170_889_0 & i_8_170_1015_0 & ~i_8_170_1392_0 & ~i_8_170_1699_0 & ~i_8_170_1824_0 & ~i_8_170_1851_0) | (~i_8_170_295_0 & ~i_8_170_516_0 & ~i_8_170_835_0 & ~i_8_170_836_0 & ~i_8_170_1031_0 & i_8_170_1078_0 & ~i_8_170_1808_0 & ~i_8_170_2068_0 & ~i_8_170_2112_0 & ~i_8_170_2121_0 & ~i_8_170_2283_0))) | (~i_8_170_1392_0 & ((~i_8_170_598_0 & ~i_8_170_1204_0 & ((~i_8_170_6_0 & ~i_8_170_813_0 & ~i_8_170_1074_0 & ~i_8_170_1393_0 & ~i_8_170_1500_0 & ~i_8_170_1870_0) | (~i_8_170_672_0 & ~i_8_170_817_0 & ~i_8_170_853_0 & ~i_8_170_2067_0))) | (~i_8_170_6_0 & ~i_8_170_1393_0 & ((~i_8_170_115_0 & ~i_8_170_601_0 & ~i_8_170_672_0 & ~i_8_170_817_0 & ~i_8_170_1087_0 & ~i_8_170_1798_0) | (~i_8_170_448_0 & ~i_8_170_516_0 & ~i_8_170_836_0 & ~i_8_170_1317_0 & ~i_8_170_1866_0 & ~i_8_170_1879_0 & ~i_8_170_2031_0 & ~i_8_170_2284_0))) | (~i_8_170_1500_0 & ((~i_8_170_295_0 & ~i_8_170_699_0 & ~i_8_170_718_0 & ~i_8_170_1870_0 & ~i_8_170_1879_0 & ~i_8_170_2092_0 & ~i_8_170_2118_0) | (~i_8_170_249_0 & ~i_8_170_1078_0 & ~i_8_170_1308_0 & ~i_8_170_1394_0 & ~i_8_170_1446_0 & ~i_8_170_2067_0 & ~i_8_170_2122_0 & ~i_8_170_2283_0))))) | (~i_8_170_249_0 & ((i_8_170_490_0 & ~i_8_170_816_0 & ~i_8_170_1074_0 & ~i_8_170_1078_0 & ~i_8_170_1394_0 & ~i_8_170_1636_0 & ~i_8_170_2121_0) | (~i_8_170_672_0 & ~i_8_170_836_0 & ~i_8_170_853_0 & ~i_8_170_889_0 & ~i_8_170_1308_0 & ~i_8_170_1662_0 & ~i_8_170_2031_0 & ~i_8_170_2283_0))) | (~i_8_170_1851_0 & ((~i_8_170_295_0 & ((~i_8_170_6_0 & ~i_8_170_601_0 & ~i_8_170_816_0 & ~i_8_170_1636_0 & ~i_8_170_1848_0 & ~i_8_170_2068_0) | (~i_8_170_490_0 & ~i_8_170_672_0 & ~i_8_170_717_0 & ~i_8_170_1204_0 & ~i_8_170_1394_0 & ~i_8_170_1879_0 & ~i_8_170_1881_0 & ~i_8_170_2092_0))) | (~i_8_170_516_0 & i_8_170_699_0 & ~i_8_170_852_0 & i_8_170_1285_0 & ~i_8_170_1500_0 & ~i_8_170_1866_0) | (i_8_170_598_0 & i_8_170_601_0 & ~i_8_170_1087_0 & ~i_8_170_1156_0 & ~i_8_170_1308_0 & ~i_8_170_1394_0 & ~i_8_170_1848_0 & ~i_8_170_1879_0 & ~i_8_170_2067_0 & ~i_8_170_2283_0))) | (~i_8_170_516_0 & ~i_8_170_1394_0 & ((~i_8_170_6_0 & i_8_170_661_0 & ~i_8_170_726_0 & ~i_8_170_1204_0 & i_8_170_1824_0 & ~i_8_170_2118_0) | (~i_8_170_789_0 & ~i_8_170_816_0 & ~i_8_170_853_0 & ~i_8_170_1087_0 & ~i_8_170_1393_0 & ~i_8_170_1662_0 & ~i_8_170_1798_0 & ~i_8_170_2031_0 & ~i_8_170_2121_0 & ~i_8_170_2284_0))) | (~i_8_170_6_0 & ((~i_8_170_699_0 & ~i_8_170_835_0 & ~i_8_170_1087_0 & i_8_170_1204_0 & ~i_8_170_1308_0 & ~i_8_170_1393_0 & ~i_8_170_1662_0) | (~i_8_170_258_0 & i_8_170_295_0 & ~i_8_170_836_0 & i_8_170_1285_0 & ~i_8_170_2215_0 & ~i_8_170_2283_0))) | (i_8_170_699_0 & i_8_170_1015_0 & i_8_170_1437_0 & ~i_8_170_2031_0) | (i_8_170_606_0 & ~i_8_170_817_0 & i_8_170_2073_0));
endmodule



// Benchmark "kernel_8_171" written by ABC on Sun Jul 19 10:06:00 2020

module kernel_8_171 ( 
    i_8_171_53_0, i_8_171_58_0, i_8_171_62_0, i_8_171_83_0, i_8_171_115_0,
    i_8_171_136_0, i_8_171_142_0, i_8_171_143_0, i_8_171_147_0,
    i_8_171_195_0, i_8_171_225_0, i_8_171_227_0, i_8_171_238_0,
    i_8_171_262_0, i_8_171_364_0, i_8_171_418_0, i_8_171_491_0,
    i_8_171_493_0, i_8_171_555_0, i_8_171_556_0, i_8_171_557_0,
    i_8_171_575_0, i_8_171_781_0, i_8_171_782_0, i_8_171_786_0,
    i_8_171_964_0, i_8_171_976_0, i_8_171_993_0, i_8_171_994_0,
    i_8_171_996_0, i_8_171_1008_0, i_8_171_1051_0, i_8_171_1110_0,
    i_8_171_1111_0, i_8_171_1120_0, i_8_171_1121_0, i_8_171_1124_0,
    i_8_171_1191_0, i_8_171_1263_0, i_8_171_1281_0, i_8_171_1282_0,
    i_8_171_1284_0, i_8_171_1285_0, i_8_171_1305_0, i_8_171_1306_0,
    i_8_171_1307_0, i_8_171_1315_0, i_8_171_1330_0, i_8_171_1331_0,
    i_8_171_1344_0, i_8_171_1408_0, i_8_171_1409_0, i_8_171_1411_0,
    i_8_171_1435_0, i_8_171_1436_0, i_8_171_1437_0, i_8_171_1470_0,
    i_8_171_1474_0, i_8_171_1506_0, i_8_171_1507_0, i_8_171_1509_0,
    i_8_171_1545_0, i_8_171_1565_0, i_8_171_1573_0, i_8_171_1574_0,
    i_8_171_1590_0, i_8_171_1629_0, i_8_171_1653_0, i_8_171_1655_0,
    i_8_171_1682_0, i_8_171_1687_0, i_8_171_1700_0, i_8_171_1723_0,
    i_8_171_1740_0, i_8_171_1747_0, i_8_171_1804_0, i_8_171_1807_0,
    i_8_171_1875_0, i_8_171_1876_0, i_8_171_1888_0, i_8_171_1903_0,
    i_8_171_1925_0, i_8_171_1990_0, i_8_171_1991_0, i_8_171_1992_0,
    i_8_171_2005_0, i_8_171_2093_0, i_8_171_2102_0, i_8_171_2133_0,
    i_8_171_2147_0, i_8_171_2152_0, i_8_171_2155_0, i_8_171_2214_0,
    i_8_171_2215_0, i_8_171_2216_0, i_8_171_2242_0, i_8_171_2245_0,
    i_8_171_2246_0, i_8_171_2249_0, i_8_171_2260_0,
    o_8_171_0_0  );
  input  i_8_171_53_0, i_8_171_58_0, i_8_171_62_0, i_8_171_83_0,
    i_8_171_115_0, i_8_171_136_0, i_8_171_142_0, i_8_171_143_0,
    i_8_171_147_0, i_8_171_195_0, i_8_171_225_0, i_8_171_227_0,
    i_8_171_238_0, i_8_171_262_0, i_8_171_364_0, i_8_171_418_0,
    i_8_171_491_0, i_8_171_493_0, i_8_171_555_0, i_8_171_556_0,
    i_8_171_557_0, i_8_171_575_0, i_8_171_781_0, i_8_171_782_0,
    i_8_171_786_0, i_8_171_964_0, i_8_171_976_0, i_8_171_993_0,
    i_8_171_994_0, i_8_171_996_0, i_8_171_1008_0, i_8_171_1051_0,
    i_8_171_1110_0, i_8_171_1111_0, i_8_171_1120_0, i_8_171_1121_0,
    i_8_171_1124_0, i_8_171_1191_0, i_8_171_1263_0, i_8_171_1281_0,
    i_8_171_1282_0, i_8_171_1284_0, i_8_171_1285_0, i_8_171_1305_0,
    i_8_171_1306_0, i_8_171_1307_0, i_8_171_1315_0, i_8_171_1330_0,
    i_8_171_1331_0, i_8_171_1344_0, i_8_171_1408_0, i_8_171_1409_0,
    i_8_171_1411_0, i_8_171_1435_0, i_8_171_1436_0, i_8_171_1437_0,
    i_8_171_1470_0, i_8_171_1474_0, i_8_171_1506_0, i_8_171_1507_0,
    i_8_171_1509_0, i_8_171_1545_0, i_8_171_1565_0, i_8_171_1573_0,
    i_8_171_1574_0, i_8_171_1590_0, i_8_171_1629_0, i_8_171_1653_0,
    i_8_171_1655_0, i_8_171_1682_0, i_8_171_1687_0, i_8_171_1700_0,
    i_8_171_1723_0, i_8_171_1740_0, i_8_171_1747_0, i_8_171_1804_0,
    i_8_171_1807_0, i_8_171_1875_0, i_8_171_1876_0, i_8_171_1888_0,
    i_8_171_1903_0, i_8_171_1925_0, i_8_171_1990_0, i_8_171_1991_0,
    i_8_171_1992_0, i_8_171_2005_0, i_8_171_2093_0, i_8_171_2102_0,
    i_8_171_2133_0, i_8_171_2147_0, i_8_171_2152_0, i_8_171_2155_0,
    i_8_171_2214_0, i_8_171_2215_0, i_8_171_2216_0, i_8_171_2242_0,
    i_8_171_2245_0, i_8_171_2246_0, i_8_171_2249_0, i_8_171_2260_0;
  output o_8_171_0_0;
  assign o_8_171_0_0 = ~((~i_8_171_1470_0 & ((i_8_171_83_0 & ((~i_8_171_1121_0 & ~i_8_171_1474_0 & i_8_171_1747_0) | (~i_8_171_143_0 & ~i_8_171_1306_0 & ~i_8_171_2093_0 & ~i_8_171_2215_0))) | (~i_8_171_58_0 & ~i_8_171_227_0 & ~i_8_171_238_0 & ~i_8_171_418_0 & i_8_171_1282_0 & ~i_8_171_1307_0 & ~i_8_171_1330_0 & ~i_8_171_1565_0 & ~i_8_171_1574_0 & ~i_8_171_2152_0 & ~i_8_171_2215_0))) | (~i_8_171_147_0 & ((~i_8_171_143_0 & ~i_8_171_786_0 & ~i_8_171_993_0 & i_8_171_1111_0 & i_8_171_1408_0) | (~i_8_171_491_0 & ~i_8_171_1545_0 & ~i_8_171_1574_0 & ~i_8_171_1876_0 & i_8_171_2245_0))) | (~i_8_171_996_0 & ((~i_8_171_225_0 & ~i_8_171_993_0 & i_8_171_1110_0 & ~i_8_171_1307_0 & ~i_8_171_1409_0) | (~i_8_171_227_0 & ~i_8_171_1191_0 & i_8_171_1411_0 & ~i_8_171_2005_0 & ~i_8_171_2214_0))) | (~i_8_171_1124_0 & ((~i_8_171_993_0 & i_8_171_1436_0 & ~i_8_171_1573_0 & ~i_8_171_1574_0 & ~i_8_171_1687_0) | (~i_8_171_364_0 & i_8_171_491_0 & ~i_8_171_994_0 & ~i_8_171_1315_0 & i_8_171_1409_0 & ~i_8_171_1509_0 & ~i_8_171_1565_0 & ~i_8_171_1991_0 & ~i_8_171_2215_0 & ~i_8_171_2216_0))) | (i_8_171_1263_0 & ((~i_8_171_786_0 & ~i_8_171_994_0 & ~i_8_171_1315_0 & ~i_8_171_1408_0) | (i_8_171_1408_0 & ~i_8_171_2215_0))) | (~i_8_171_2214_0 & ((~i_8_171_964_0 & ((~i_8_171_136_0 & ~i_8_171_2152_0 & ((i_8_171_364_0 & ~i_8_171_786_0 & ~i_8_171_1111_0 & ~i_8_171_1191_0 & ~i_8_171_1305_0) | (~i_8_171_62_0 & ~i_8_171_225_0 & ~i_8_171_491_0 & ~i_8_171_1315_0 & ~i_8_171_1506_0 & ~i_8_171_1507_0 & ~i_8_171_1509_0 & ~i_8_171_1574_0 & ~i_8_171_1925_0 & ~i_8_171_1990_0 & ~i_8_171_1991_0 & ~i_8_171_2155_0 & ~i_8_171_2215_0))) | (i_8_171_1281_0 & ~i_8_171_1315_0 & ~i_8_171_1331_0 & ~i_8_171_1506_0 & ~i_8_171_1507_0))) | (i_8_171_493_0 & ~i_8_171_786_0 & ~i_8_171_1331_0 & ~i_8_171_1509_0 & ~i_8_171_1565_0 & ~i_8_171_1875_0 & ~i_8_171_2215_0) | (~i_8_171_993_0 & ~i_8_171_1191_0 & i_8_171_1747_0 & i_8_171_2155_0))) | (~i_8_171_2152_0 & ((~i_8_171_62_0 & ((~i_8_171_994_0 & ~i_8_171_1121_0 & ~i_8_171_1574_0 & ~i_8_171_1629_0 & i_8_171_1682_0) | (~i_8_171_53_0 & ~i_8_171_83_0 & ~i_8_171_418_0 & ~i_8_171_1306_0 & i_8_171_1507_0 & ~i_8_171_1545_0 & ~i_8_171_1573_0 & ~i_8_171_1875_0 & ~i_8_171_2215_0 & ~i_8_171_2216_0))) | (~i_8_171_491_0 & ((~i_8_171_143_0 & ~i_8_171_1051_0 & i_8_171_1111_0 & ~i_8_171_1990_0) | (i_8_171_1282_0 & ~i_8_171_1474_0 & ~i_8_171_1509_0 & ~i_8_171_1991_0 & ~i_8_171_2102_0))))) | (~i_8_171_227_0 & ((~i_8_171_53_0 & ((i_8_171_1437_0 & ~i_8_171_1687_0 & ~i_8_171_1875_0) | (~i_8_171_964_0 & ~i_8_171_1306_0 & ~i_8_171_1990_0 & ~i_8_171_2093_0 & i_8_171_2147_0))) | (~i_8_171_493_0 & ~i_8_171_1545_0 & ~i_8_171_1740_0 & i_8_171_2133_0) | (~i_8_171_1051_0 & ~i_8_171_1315_0 & ~i_8_171_1409_0 & ~i_8_171_1435_0 & ~i_8_171_1574_0 & i_8_171_2147_0 & ~i_8_171_2155_0))) | (~i_8_171_225_0 & ((i_8_171_115_0 & ~i_8_171_195_0 & ~i_8_171_1474_0 & ~i_8_171_1573_0 & i_8_171_1888_0) | (~i_8_171_58_0 & i_8_171_556_0 & ~i_8_171_1436_0 & ~i_8_171_2155_0))) | (~i_8_171_195_0 & ((~i_8_171_143_0 & ~i_8_171_491_0 & ~i_8_171_1281_0 & ~i_8_171_1284_0 & ~i_8_171_1305_0 & i_8_171_1411_0 & ~i_8_171_1740_0 & ~i_8_171_1888_0) | (~i_8_171_964_0 & ~i_8_171_1191_0 & i_8_171_1807_0 & ~i_8_171_1990_0))) | (~i_8_171_1307_0 & ((~i_8_171_994_0 & ~i_8_171_1565_0 & i_8_171_1991_0 & (i_8_171_227_0 | (~i_8_171_993_0 & ~i_8_171_1315_0 & i_8_171_1990_0))) | (i_8_171_1285_0 & ~i_8_171_1409_0 & ~i_8_171_1655_0 & ~i_8_171_1875_0))) | (~i_8_171_2215_0 & ((~i_8_171_143_0 & ((~i_8_171_993_0 & i_8_171_1435_0) | (i_8_171_781_0 & ~i_8_171_1331_0 & ~i_8_171_1507_0 & ~i_8_171_1925_0))) | (i_8_171_1282_0 & ((~i_8_171_142_0 & i_8_171_1747_0) | (~i_8_171_58_0 & ~i_8_171_1315_0 & i_8_171_1991_0))) | (~i_8_171_2216_0 & ((~i_8_171_993_0 & i_8_171_1110_0 & ~i_8_171_1191_0 & ~i_8_171_1509_0 & i_8_171_1992_0) | (i_8_171_1344_0 & ~i_8_171_1653_0 & ~i_8_171_1875_0 & ~i_8_171_2093_0))) | (~i_8_171_781_0 & ~i_8_171_1284_0 & ~i_8_171_1687_0 & i_8_171_1807_0 & ~i_8_171_2246_0))) | (~i_8_171_58_0 & ((~i_8_171_1474_0 & ~i_8_171_1545_0 & i_8_171_2246_0) | (~i_8_171_143_0 & ~i_8_171_1051_0 & ~i_8_171_1120_0 & ~i_8_171_1991_0 & i_8_171_2093_0 & i_8_171_2216_0 & ~i_8_171_2249_0))) | (~i_8_171_142_0 & ((i_8_171_1307_0 & i_8_171_1408_0 & ~i_8_171_1506_0 & ~i_8_171_1903_0) | (~i_8_171_136_0 & i_8_171_993_0 & i_8_171_994_0 & ~i_8_171_1191_0 & ~i_8_171_1408_0 & ~i_8_171_1875_0 & ~i_8_171_2102_0 & ~i_8_171_2147_0))) | (~i_8_171_1306_0 & ((~i_8_171_1120_0 & i_8_171_1653_0 & i_8_171_1903_0) | (i_8_171_58_0 & i_8_171_136_0 & ~i_8_171_1051_0 & ~i_8_171_1747_0 & ~i_8_171_2093_0))) | (~i_8_171_1120_0 & ((i_8_171_1281_0 & ~i_8_171_1411_0 & i_8_171_1990_0) | (~i_8_171_1331_0 & ~i_8_171_1408_0 & ~i_8_171_1747_0 & i_8_171_1888_0 & ~i_8_171_1992_0))) | (~i_8_171_1315_0 & ((i_8_171_1435_0 & ~i_8_171_1509_0 & ~i_8_171_1565_0 & ~i_8_171_1573_0) | (~i_8_171_1506_0 & ~i_8_171_1876_0 & i_8_171_1990_0 & ~i_8_171_1991_0 & ~i_8_171_1992_0 & ~i_8_171_2093_0 & ~i_8_171_2242_0))) | (~i_8_171_1875_0 & ((~i_8_171_557_0 & i_8_171_1285_0 & ~i_8_171_1655_0 & i_8_171_1682_0) | (i_8_171_1284_0 & i_8_171_2155_0) | (~i_8_171_1330_0 & ~i_8_171_1687_0 & i_8_171_2245_0))) | (~i_8_171_1506_0 & ~i_8_171_1507_0 & i_8_171_1629_0 & i_8_171_1747_0 & ~i_8_171_2102_0) | (i_8_171_557_0 & ~i_8_171_2216_0));
endmodule



// Benchmark "kernel_8_172" written by ABC on Sun Jul 19 10:06:01 2020

module kernel_8_172 ( 
    i_8_172_53_0, i_8_172_59_0, i_8_172_62_0, i_8_172_63_0, i_8_172_98_0,
    i_8_172_139_0, i_8_172_143_0, i_8_172_188_0, i_8_172_259_0,
    i_8_172_260_0, i_8_172_287_0, i_8_172_304_0, i_8_172_346_0,
    i_8_172_360_0, i_8_172_366_0, i_8_172_376_0, i_8_172_385_0,
    i_8_172_422_0, i_8_172_438_0, i_8_172_448_0, i_8_172_457_0,
    i_8_172_460_0, i_8_172_461_0, i_8_172_485_0, i_8_172_502_0,
    i_8_172_508_0, i_8_172_511_0, i_8_172_512_0, i_8_172_529_0,
    i_8_172_587_0, i_8_172_599_0, i_8_172_749_0, i_8_172_763_0,
    i_8_172_764_0, i_8_172_790_0, i_8_172_824_0, i_8_172_851_0,
    i_8_172_854_0, i_8_172_880_0, i_8_172_958_0, i_8_172_994_0,
    i_8_172_995_0, i_8_172_997_0, i_8_172_1016_0, i_8_172_1051_0,
    i_8_172_1052_0, i_8_172_1075_0, i_8_172_1078_0, i_8_172_1079_0,
    i_8_172_1094_0, i_8_172_1103_0, i_8_172_1105_0, i_8_172_1114_0,
    i_8_172_1124_0, i_8_172_1130_0, i_8_172_1192_0, i_8_172_1193_0,
    i_8_172_1267_0, i_8_172_1306_0, i_8_172_1307_0, i_8_172_1310_0,
    i_8_172_1315_0, i_8_172_1350_0, i_8_172_1391_0, i_8_172_1394_0,
    i_8_172_1407_0, i_8_172_1508_0, i_8_172_1546_0, i_8_172_1553_0,
    i_8_172_1573_0, i_8_172_1574_0, i_8_172_1633_0, i_8_172_1653_0,
    i_8_172_1681_0, i_8_172_1690_0, i_8_172_1724_0, i_8_172_1726_0,
    i_8_172_1727_0, i_8_172_1753_0, i_8_172_1763_0, i_8_172_1837_0,
    i_8_172_1859_0, i_8_172_1862_0, i_8_172_1870_0, i_8_172_1879_0,
    i_8_172_1880_0, i_8_172_1888_0, i_8_172_1907_0, i_8_172_2002_0,
    i_8_172_2006_0, i_8_172_2033_0, i_8_172_2139_0, i_8_172_2154_0,
    i_8_172_2155_0, i_8_172_2170_0, i_8_172_2187_0, i_8_172_2197_0,
    i_8_172_2215_0, i_8_172_2237_0, i_8_172_2247_0,
    o_8_172_0_0  );
  input  i_8_172_53_0, i_8_172_59_0, i_8_172_62_0, i_8_172_63_0,
    i_8_172_98_0, i_8_172_139_0, i_8_172_143_0, i_8_172_188_0,
    i_8_172_259_0, i_8_172_260_0, i_8_172_287_0, i_8_172_304_0,
    i_8_172_346_0, i_8_172_360_0, i_8_172_366_0, i_8_172_376_0,
    i_8_172_385_0, i_8_172_422_0, i_8_172_438_0, i_8_172_448_0,
    i_8_172_457_0, i_8_172_460_0, i_8_172_461_0, i_8_172_485_0,
    i_8_172_502_0, i_8_172_508_0, i_8_172_511_0, i_8_172_512_0,
    i_8_172_529_0, i_8_172_587_0, i_8_172_599_0, i_8_172_749_0,
    i_8_172_763_0, i_8_172_764_0, i_8_172_790_0, i_8_172_824_0,
    i_8_172_851_0, i_8_172_854_0, i_8_172_880_0, i_8_172_958_0,
    i_8_172_994_0, i_8_172_995_0, i_8_172_997_0, i_8_172_1016_0,
    i_8_172_1051_0, i_8_172_1052_0, i_8_172_1075_0, i_8_172_1078_0,
    i_8_172_1079_0, i_8_172_1094_0, i_8_172_1103_0, i_8_172_1105_0,
    i_8_172_1114_0, i_8_172_1124_0, i_8_172_1130_0, i_8_172_1192_0,
    i_8_172_1193_0, i_8_172_1267_0, i_8_172_1306_0, i_8_172_1307_0,
    i_8_172_1310_0, i_8_172_1315_0, i_8_172_1350_0, i_8_172_1391_0,
    i_8_172_1394_0, i_8_172_1407_0, i_8_172_1508_0, i_8_172_1546_0,
    i_8_172_1553_0, i_8_172_1573_0, i_8_172_1574_0, i_8_172_1633_0,
    i_8_172_1653_0, i_8_172_1681_0, i_8_172_1690_0, i_8_172_1724_0,
    i_8_172_1726_0, i_8_172_1727_0, i_8_172_1753_0, i_8_172_1763_0,
    i_8_172_1837_0, i_8_172_1859_0, i_8_172_1862_0, i_8_172_1870_0,
    i_8_172_1879_0, i_8_172_1880_0, i_8_172_1888_0, i_8_172_1907_0,
    i_8_172_2002_0, i_8_172_2006_0, i_8_172_2033_0, i_8_172_2139_0,
    i_8_172_2154_0, i_8_172_2155_0, i_8_172_2170_0, i_8_172_2187_0,
    i_8_172_2197_0, i_8_172_2215_0, i_8_172_2237_0, i_8_172_2247_0;
  output o_8_172_0_0;
  assign o_8_172_0_0 = 0;
endmodule



// Benchmark "kernel_8_173" written by ABC on Sun Jul 19 10:06:02 2020

module kernel_8_173 ( 
    i_8_173_25_0, i_8_173_40_0, i_8_173_42_0, i_8_173_250_0, i_8_173_257_0,
    i_8_173_277_0, i_8_173_303_0, i_8_173_367_0, i_8_173_374_0,
    i_8_173_426_0, i_8_173_445_0, i_8_173_471_0, i_8_173_493_0,
    i_8_173_499_0, i_8_173_552_0, i_8_173_553_0, i_8_173_555_0,
    i_8_173_592_0, i_8_173_593_0, i_8_173_597_0, i_8_173_604_0,
    i_8_173_610_0, i_8_173_635_0, i_8_173_653_0, i_8_173_673_0,
    i_8_173_674_0, i_8_173_677_0, i_8_173_718_0, i_8_173_719_0,
    i_8_173_729_0, i_8_173_841_0, i_8_173_852_0, i_8_173_853_0,
    i_8_173_868_0, i_8_173_877_0, i_8_173_880_0, i_8_173_881_0,
    i_8_173_958_0, i_8_173_959_0, i_8_173_994_0, i_8_173_1035_0,
    i_8_173_1075_0, i_8_173_1078_0, i_8_173_1105_0, i_8_173_1113_0,
    i_8_173_1114_0, i_8_173_1186_0, i_8_173_1201_0, i_8_173_1203_0,
    i_8_173_1227_0, i_8_173_1230_0, i_8_173_1246_0, i_8_173_1263_0,
    i_8_173_1320_0, i_8_173_1345_0, i_8_173_1410_0, i_8_173_1411_0,
    i_8_173_1423_0, i_8_173_1440_0, i_8_173_1482_0, i_8_173_1483_0,
    i_8_173_1485_0, i_8_173_1488_0, i_8_173_1498_0, i_8_173_1529_0,
    i_8_173_1534_0, i_8_173_1536_0, i_8_173_1600_0, i_8_173_1601_0,
    i_8_173_1605_0, i_8_173_1644_0, i_8_173_1705_0, i_8_173_1715_0,
    i_8_173_1749_0, i_8_173_1813_0, i_8_173_1826_0, i_8_173_1853_0,
    i_8_173_1869_0, i_8_173_1870_0, i_8_173_1875_0, i_8_173_1878_0,
    i_8_173_1888_0, i_8_173_1918_0, i_8_173_1921_0, i_8_173_1951_0,
    i_8_173_1965_0, i_8_173_1974_0, i_8_173_1975_0, i_8_173_1983_0,
    i_8_173_1987_0, i_8_173_1997_0, i_8_173_2007_0, i_8_173_2049_0,
    i_8_173_2065_0, i_8_173_2068_0, i_8_173_2229_0, i_8_173_2231_0,
    i_8_173_2239_0, i_8_173_2242_0, i_8_173_2257_0,
    o_8_173_0_0  );
  input  i_8_173_25_0, i_8_173_40_0, i_8_173_42_0, i_8_173_250_0,
    i_8_173_257_0, i_8_173_277_0, i_8_173_303_0, i_8_173_367_0,
    i_8_173_374_0, i_8_173_426_0, i_8_173_445_0, i_8_173_471_0,
    i_8_173_493_0, i_8_173_499_0, i_8_173_552_0, i_8_173_553_0,
    i_8_173_555_0, i_8_173_592_0, i_8_173_593_0, i_8_173_597_0,
    i_8_173_604_0, i_8_173_610_0, i_8_173_635_0, i_8_173_653_0,
    i_8_173_673_0, i_8_173_674_0, i_8_173_677_0, i_8_173_718_0,
    i_8_173_719_0, i_8_173_729_0, i_8_173_841_0, i_8_173_852_0,
    i_8_173_853_0, i_8_173_868_0, i_8_173_877_0, i_8_173_880_0,
    i_8_173_881_0, i_8_173_958_0, i_8_173_959_0, i_8_173_994_0,
    i_8_173_1035_0, i_8_173_1075_0, i_8_173_1078_0, i_8_173_1105_0,
    i_8_173_1113_0, i_8_173_1114_0, i_8_173_1186_0, i_8_173_1201_0,
    i_8_173_1203_0, i_8_173_1227_0, i_8_173_1230_0, i_8_173_1246_0,
    i_8_173_1263_0, i_8_173_1320_0, i_8_173_1345_0, i_8_173_1410_0,
    i_8_173_1411_0, i_8_173_1423_0, i_8_173_1440_0, i_8_173_1482_0,
    i_8_173_1483_0, i_8_173_1485_0, i_8_173_1488_0, i_8_173_1498_0,
    i_8_173_1529_0, i_8_173_1534_0, i_8_173_1536_0, i_8_173_1600_0,
    i_8_173_1601_0, i_8_173_1605_0, i_8_173_1644_0, i_8_173_1705_0,
    i_8_173_1715_0, i_8_173_1749_0, i_8_173_1813_0, i_8_173_1826_0,
    i_8_173_1853_0, i_8_173_1869_0, i_8_173_1870_0, i_8_173_1875_0,
    i_8_173_1878_0, i_8_173_1888_0, i_8_173_1918_0, i_8_173_1921_0,
    i_8_173_1951_0, i_8_173_1965_0, i_8_173_1974_0, i_8_173_1975_0,
    i_8_173_1983_0, i_8_173_1987_0, i_8_173_1997_0, i_8_173_2007_0,
    i_8_173_2049_0, i_8_173_2065_0, i_8_173_2068_0, i_8_173_2229_0,
    i_8_173_2231_0, i_8_173_2239_0, i_8_173_2242_0, i_8_173_2257_0;
  output o_8_173_0_0;
  assign o_8_173_0_0 = 0;
endmodule



// Benchmark "kernel_8_174" written by ABC on Sun Jul 19 10:06:03 2020

module kernel_8_174 ( 
    i_8_174_9_0, i_8_174_10_0, i_8_174_73_0, i_8_174_91_0, i_8_174_102_0,
    i_8_174_112_0, i_8_174_143_0, i_8_174_165_0, i_8_174_181_0,
    i_8_174_205_0, i_8_174_208_0, i_8_174_230_0, i_8_174_238_0,
    i_8_174_248_0, i_8_174_265_0, i_8_174_274_0, i_8_174_284_0,
    i_8_174_292_0, i_8_174_324_0, i_8_174_343_0, i_8_174_366_0,
    i_8_174_371_0, i_8_174_491_0, i_8_174_537_0, i_8_174_568_0,
    i_8_174_609_0, i_8_174_625_0, i_8_174_626_0, i_8_174_631_0,
    i_8_174_640_0, i_8_174_662_0, i_8_174_688_0, i_8_174_705_0,
    i_8_174_724_0, i_8_174_780_0, i_8_174_811_0, i_8_174_838_0,
    i_8_174_878_0, i_8_174_929_0, i_8_174_940_0, i_8_174_970_0,
    i_8_174_982_0, i_8_174_1009_0, i_8_174_1019_0, i_8_174_1053_0,
    i_8_174_1073_0, i_8_174_1100_0, i_8_174_1102_0, i_8_174_1104_0,
    i_8_174_1113_0, i_8_174_1152_0, i_8_174_1171_0, i_8_174_1172_0,
    i_8_174_1173_0, i_8_174_1192_0, i_8_174_1245_0, i_8_174_1258_0,
    i_8_174_1281_0, i_8_174_1297_0, i_8_174_1306_0, i_8_174_1312_0,
    i_8_174_1336_0, i_8_174_1368_0, i_8_174_1404_0, i_8_174_1475_0,
    i_8_174_1539_0, i_8_174_1554_0, i_8_174_1589_0, i_8_174_1668_0,
    i_8_174_1672_0, i_8_174_1675_0, i_8_174_1687_0, i_8_174_1690_0,
    i_8_174_1733_0, i_8_174_1758_0, i_8_174_1759_0, i_8_174_1789_0,
    i_8_174_1804_0, i_8_174_1831_0, i_8_174_1842_0, i_8_174_1846_0,
    i_8_174_1868_0, i_8_174_1873_0, i_8_174_1881_0, i_8_174_1889_0,
    i_8_174_1907_0, i_8_174_1937_0, i_8_174_1992_0, i_8_174_2070_0,
    i_8_174_2100_0, i_8_174_2129_0, i_8_174_2150_0, i_8_174_2151_0,
    i_8_174_2161_0, i_8_174_2205_0, i_8_174_2223_0, i_8_174_2241_0,
    i_8_174_2261_0, i_8_174_2287_0, i_8_174_2296_0,
    o_8_174_0_0  );
  input  i_8_174_9_0, i_8_174_10_0, i_8_174_73_0, i_8_174_91_0,
    i_8_174_102_0, i_8_174_112_0, i_8_174_143_0, i_8_174_165_0,
    i_8_174_181_0, i_8_174_205_0, i_8_174_208_0, i_8_174_230_0,
    i_8_174_238_0, i_8_174_248_0, i_8_174_265_0, i_8_174_274_0,
    i_8_174_284_0, i_8_174_292_0, i_8_174_324_0, i_8_174_343_0,
    i_8_174_366_0, i_8_174_371_0, i_8_174_491_0, i_8_174_537_0,
    i_8_174_568_0, i_8_174_609_0, i_8_174_625_0, i_8_174_626_0,
    i_8_174_631_0, i_8_174_640_0, i_8_174_662_0, i_8_174_688_0,
    i_8_174_705_0, i_8_174_724_0, i_8_174_780_0, i_8_174_811_0,
    i_8_174_838_0, i_8_174_878_0, i_8_174_929_0, i_8_174_940_0,
    i_8_174_970_0, i_8_174_982_0, i_8_174_1009_0, i_8_174_1019_0,
    i_8_174_1053_0, i_8_174_1073_0, i_8_174_1100_0, i_8_174_1102_0,
    i_8_174_1104_0, i_8_174_1113_0, i_8_174_1152_0, i_8_174_1171_0,
    i_8_174_1172_0, i_8_174_1173_0, i_8_174_1192_0, i_8_174_1245_0,
    i_8_174_1258_0, i_8_174_1281_0, i_8_174_1297_0, i_8_174_1306_0,
    i_8_174_1312_0, i_8_174_1336_0, i_8_174_1368_0, i_8_174_1404_0,
    i_8_174_1475_0, i_8_174_1539_0, i_8_174_1554_0, i_8_174_1589_0,
    i_8_174_1668_0, i_8_174_1672_0, i_8_174_1675_0, i_8_174_1687_0,
    i_8_174_1690_0, i_8_174_1733_0, i_8_174_1758_0, i_8_174_1759_0,
    i_8_174_1789_0, i_8_174_1804_0, i_8_174_1831_0, i_8_174_1842_0,
    i_8_174_1846_0, i_8_174_1868_0, i_8_174_1873_0, i_8_174_1881_0,
    i_8_174_1889_0, i_8_174_1907_0, i_8_174_1937_0, i_8_174_1992_0,
    i_8_174_2070_0, i_8_174_2100_0, i_8_174_2129_0, i_8_174_2150_0,
    i_8_174_2151_0, i_8_174_2161_0, i_8_174_2205_0, i_8_174_2223_0,
    i_8_174_2241_0, i_8_174_2261_0, i_8_174_2287_0, i_8_174_2296_0;
  output o_8_174_0_0;
  assign o_8_174_0_0 = 0;
endmodule



// Benchmark "kernel_8_175" written by ABC on Sun Jul 19 10:06:04 2020

module kernel_8_175 ( 
    i_8_175_42_0, i_8_175_176_0, i_8_175_189_0, i_8_175_190_0,
    i_8_175_242_0, i_8_175_246_0, i_8_175_311_0, i_8_175_366_0,
    i_8_175_369_0, i_8_175_394_0, i_8_175_462_0, i_8_175_466_0,
    i_8_175_525_0, i_8_175_535_0, i_8_175_555_0, i_8_175_595_0,
    i_8_175_596_0, i_8_175_613_0, i_8_175_660_0, i_8_175_661_0,
    i_8_175_696_0, i_8_175_702_0, i_8_175_706_0, i_8_175_729_0,
    i_8_175_730_0, i_8_175_747_0, i_8_175_748_0, i_8_175_814_0,
    i_8_175_825_0, i_8_175_837_0, i_8_175_838_0, i_8_175_859_0,
    i_8_175_915_0, i_8_175_940_0, i_8_175_1126_0, i_8_175_1174_0,
    i_8_175_1182_0, i_8_175_1183_0, i_8_175_1198_0, i_8_175_1239_0,
    i_8_175_1241_0, i_8_175_1273_0, i_8_175_1282_0, i_8_175_1284_0,
    i_8_175_1299_0, i_8_175_1306_0, i_8_175_1318_0, i_8_175_1338_0,
    i_8_175_1434_0, i_8_175_1435_0, i_8_175_1442_0, i_8_175_1471_0,
    i_8_175_1479_0, i_8_175_1498_0, i_8_175_1509_0, i_8_175_1524_0,
    i_8_175_1525_0, i_8_175_1533_0, i_8_175_1540_0, i_8_175_1546_0,
    i_8_175_1606_0, i_8_175_1633_0, i_8_175_1641_0, i_8_175_1642_0,
    i_8_175_1647_0, i_8_175_1648_0, i_8_175_1687_0, i_8_175_1818_0,
    i_8_175_1821_0, i_8_175_1854_0, i_8_175_1858_0, i_8_175_1909_0,
    i_8_175_1915_0, i_8_175_1917_0, i_8_175_1930_0, i_8_175_1948_0,
    i_8_175_1962_0, i_8_175_1969_0, i_8_175_1992_0, i_8_175_2038_0,
    i_8_175_2047_0, i_8_175_2058_0, i_8_175_2065_0, i_8_175_2066_0,
    i_8_175_2089_0, i_8_175_2091_0, i_8_175_2119_0, i_8_175_2122_0,
    i_8_175_2136_0, i_8_175_2170_0, i_8_175_2172_0, i_8_175_2173_0,
    i_8_175_2200_0, i_8_175_2218_0, i_8_175_2221_0, i_8_175_2233_0,
    i_8_175_2248_0, i_8_175_2253_0, i_8_175_2274_0, i_8_175_2286_0,
    o_8_175_0_0  );
  input  i_8_175_42_0, i_8_175_176_0, i_8_175_189_0, i_8_175_190_0,
    i_8_175_242_0, i_8_175_246_0, i_8_175_311_0, i_8_175_366_0,
    i_8_175_369_0, i_8_175_394_0, i_8_175_462_0, i_8_175_466_0,
    i_8_175_525_0, i_8_175_535_0, i_8_175_555_0, i_8_175_595_0,
    i_8_175_596_0, i_8_175_613_0, i_8_175_660_0, i_8_175_661_0,
    i_8_175_696_0, i_8_175_702_0, i_8_175_706_0, i_8_175_729_0,
    i_8_175_730_0, i_8_175_747_0, i_8_175_748_0, i_8_175_814_0,
    i_8_175_825_0, i_8_175_837_0, i_8_175_838_0, i_8_175_859_0,
    i_8_175_915_0, i_8_175_940_0, i_8_175_1126_0, i_8_175_1174_0,
    i_8_175_1182_0, i_8_175_1183_0, i_8_175_1198_0, i_8_175_1239_0,
    i_8_175_1241_0, i_8_175_1273_0, i_8_175_1282_0, i_8_175_1284_0,
    i_8_175_1299_0, i_8_175_1306_0, i_8_175_1318_0, i_8_175_1338_0,
    i_8_175_1434_0, i_8_175_1435_0, i_8_175_1442_0, i_8_175_1471_0,
    i_8_175_1479_0, i_8_175_1498_0, i_8_175_1509_0, i_8_175_1524_0,
    i_8_175_1525_0, i_8_175_1533_0, i_8_175_1540_0, i_8_175_1546_0,
    i_8_175_1606_0, i_8_175_1633_0, i_8_175_1641_0, i_8_175_1642_0,
    i_8_175_1647_0, i_8_175_1648_0, i_8_175_1687_0, i_8_175_1818_0,
    i_8_175_1821_0, i_8_175_1854_0, i_8_175_1858_0, i_8_175_1909_0,
    i_8_175_1915_0, i_8_175_1917_0, i_8_175_1930_0, i_8_175_1948_0,
    i_8_175_1962_0, i_8_175_1969_0, i_8_175_1992_0, i_8_175_2038_0,
    i_8_175_2047_0, i_8_175_2058_0, i_8_175_2065_0, i_8_175_2066_0,
    i_8_175_2089_0, i_8_175_2091_0, i_8_175_2119_0, i_8_175_2122_0,
    i_8_175_2136_0, i_8_175_2170_0, i_8_175_2172_0, i_8_175_2173_0,
    i_8_175_2200_0, i_8_175_2218_0, i_8_175_2221_0, i_8_175_2233_0,
    i_8_175_2248_0, i_8_175_2253_0, i_8_175_2274_0, i_8_175_2286_0;
  output o_8_175_0_0;
  assign o_8_175_0_0 = 0;
endmodule



// Benchmark "kernel_8_176" written by ABC on Sun Jul 19 10:06:06 2020

module kernel_8_176 ( 
    i_8_176_7_0, i_8_176_35_0, i_8_176_78_0, i_8_176_84_0, i_8_176_87_0,
    i_8_176_88_0, i_8_176_135_0, i_8_176_191_0, i_8_176_230_0,
    i_8_176_231_0, i_8_176_233_0, i_8_176_242_0, i_8_176_249_0,
    i_8_176_259_0, i_8_176_260_0, i_8_176_264_0, i_8_176_267_0,
    i_8_176_285_0, i_8_176_340_0, i_8_176_381_0, i_8_176_395_0,
    i_8_176_462_0, i_8_176_464_0, i_8_176_466_0, i_8_176_489_0,
    i_8_176_490_0, i_8_176_553_0, i_8_176_556_0, i_8_176_592_0,
    i_8_176_599_0, i_8_176_673_0, i_8_176_674_0, i_8_176_690_0,
    i_8_176_691_0, i_8_176_698_0, i_8_176_717_0, i_8_176_719_0,
    i_8_176_736_0, i_8_176_737_0, i_8_176_825_0, i_8_176_838_0,
    i_8_176_895_0, i_8_176_927_0, i_8_176_971_0, i_8_176_991_0,
    i_8_176_993_0, i_8_176_994_0, i_8_176_995_0, i_8_176_997_0,
    i_8_176_998_0, i_8_176_1047_0, i_8_176_1056_0, i_8_176_1060_0,
    i_8_176_1131_0, i_8_176_1132_0, i_8_176_1133_0, i_8_176_1137_0,
    i_8_176_1139_0, i_8_176_1186_0, i_8_176_1203_0, i_8_176_1204_0,
    i_8_176_1205_0, i_8_176_1236_0, i_8_176_1266_0, i_8_176_1293_0,
    i_8_176_1306_0, i_8_176_1315_0, i_8_176_1365_0, i_8_176_1385_0,
    i_8_176_1446_0, i_8_176_1457_0, i_8_176_1475_0, i_8_176_1547_0,
    i_8_176_1606_0, i_8_176_1623_0, i_8_176_1797_0, i_8_176_1798_0,
    i_8_176_1844_0, i_8_176_1911_0, i_8_176_1916_0, i_8_176_1918_0,
    i_8_176_1922_0, i_8_176_1981_0, i_8_176_1983_0, i_8_176_1985_0,
    i_8_176_2005_0, i_8_176_2053_0, i_8_176_2055_0, i_8_176_2059_0,
    i_8_176_2060_0, i_8_176_2069_0, i_8_176_2100_0, i_8_176_2145_0,
    i_8_176_2156_0, i_8_176_2175_0, i_8_176_2193_0, i_8_176_2195_0,
    i_8_176_2226_0, i_8_176_2263_0, i_8_176_2291_0,
    o_8_176_0_0  );
  input  i_8_176_7_0, i_8_176_35_0, i_8_176_78_0, i_8_176_84_0,
    i_8_176_87_0, i_8_176_88_0, i_8_176_135_0, i_8_176_191_0,
    i_8_176_230_0, i_8_176_231_0, i_8_176_233_0, i_8_176_242_0,
    i_8_176_249_0, i_8_176_259_0, i_8_176_260_0, i_8_176_264_0,
    i_8_176_267_0, i_8_176_285_0, i_8_176_340_0, i_8_176_381_0,
    i_8_176_395_0, i_8_176_462_0, i_8_176_464_0, i_8_176_466_0,
    i_8_176_489_0, i_8_176_490_0, i_8_176_553_0, i_8_176_556_0,
    i_8_176_592_0, i_8_176_599_0, i_8_176_673_0, i_8_176_674_0,
    i_8_176_690_0, i_8_176_691_0, i_8_176_698_0, i_8_176_717_0,
    i_8_176_719_0, i_8_176_736_0, i_8_176_737_0, i_8_176_825_0,
    i_8_176_838_0, i_8_176_895_0, i_8_176_927_0, i_8_176_971_0,
    i_8_176_991_0, i_8_176_993_0, i_8_176_994_0, i_8_176_995_0,
    i_8_176_997_0, i_8_176_998_0, i_8_176_1047_0, i_8_176_1056_0,
    i_8_176_1060_0, i_8_176_1131_0, i_8_176_1132_0, i_8_176_1133_0,
    i_8_176_1137_0, i_8_176_1139_0, i_8_176_1186_0, i_8_176_1203_0,
    i_8_176_1204_0, i_8_176_1205_0, i_8_176_1236_0, i_8_176_1266_0,
    i_8_176_1293_0, i_8_176_1306_0, i_8_176_1315_0, i_8_176_1365_0,
    i_8_176_1385_0, i_8_176_1446_0, i_8_176_1457_0, i_8_176_1475_0,
    i_8_176_1547_0, i_8_176_1606_0, i_8_176_1623_0, i_8_176_1797_0,
    i_8_176_1798_0, i_8_176_1844_0, i_8_176_1911_0, i_8_176_1916_0,
    i_8_176_1918_0, i_8_176_1922_0, i_8_176_1981_0, i_8_176_1983_0,
    i_8_176_1985_0, i_8_176_2005_0, i_8_176_2053_0, i_8_176_2055_0,
    i_8_176_2059_0, i_8_176_2060_0, i_8_176_2069_0, i_8_176_2100_0,
    i_8_176_2145_0, i_8_176_2156_0, i_8_176_2175_0, i_8_176_2193_0,
    i_8_176_2195_0, i_8_176_2226_0, i_8_176_2263_0, i_8_176_2291_0;
  output o_8_176_0_0;
  assign o_8_176_0_0 = ~((~i_8_176_135_0 & ((i_8_176_462_0 & ~i_8_176_490_0 & ~i_8_176_556_0 & i_8_176_1315_0 & i_8_176_1918_0) | (~i_8_176_191_0 & ~i_8_176_462_0 & i_8_176_592_0 & ~i_8_176_698_0 & ~i_8_176_825_0 & ~i_8_176_971_0 & ~i_8_176_1186_0 & ~i_8_176_1306_0 & ~i_8_176_1365_0 & ~i_8_176_1457_0 & ~i_8_176_1606_0 & ~i_8_176_1916_0 & ~i_8_176_2055_0 & ~i_8_176_2145_0 & ~i_8_176_2156_0 & ~i_8_176_2226_0))) | (~i_8_176_466_0 & ((~i_8_176_249_0 & ((~i_8_176_230_0 & i_8_176_340_0 & ~i_8_176_381_0 & ~i_8_176_464_0 & ~i_8_176_1132_0 & ~i_8_176_1137_0 & ~i_8_176_1306_0 & ~i_8_176_1315_0 & ~i_8_176_1606_0 & ~i_8_176_1797_0 & ~i_8_176_2069_0 & ~i_8_176_2193_0 & ~i_8_176_2195_0) | (~i_8_176_553_0 & ~i_8_176_599_0 & ~i_8_176_674_0 & ~i_8_176_698_0 & ~i_8_176_1236_0 & ~i_8_176_1911_0 & ~i_8_176_2100_0 & i_8_176_2291_0))) | (~i_8_176_462_0 & ((~i_8_176_267_0 & ~i_8_176_1797_0 & ((~i_8_176_191_0 & ~i_8_176_673_0 & ~i_8_176_737_0 & ~i_8_176_1922_0 & ((~i_8_176_285_0 & ~i_8_176_592_0 & ~i_8_176_717_0 & ~i_8_176_719_0 & ~i_8_176_1133_0 & ~i_8_176_1205_0 & ~i_8_176_1547_0 & ~i_8_176_2145_0) | (~i_8_176_464_0 & i_8_176_592_0 & ~i_8_176_927_0 & ~i_8_176_994_0 & ~i_8_176_2193_0 & ~i_8_176_2195_0))) | (~i_8_176_84_0 & ~i_8_176_264_0 & ~i_8_176_464_0 & ~i_8_176_719_0 & ~i_8_176_825_0 & ~i_8_176_971_0 & ~i_8_176_1133_0 & ~i_8_176_1186_0 & ~i_8_176_1203_0 & ~i_8_176_1204_0))) | (~i_8_176_264_0 & ~i_8_176_381_0 & ~i_8_176_553_0 & ~i_8_176_592_0 & ~i_8_176_674_0 & ~i_8_176_736_0 & ~i_8_176_737_0 & ~i_8_176_1132_0 & ~i_8_176_1205_0 & ~i_8_176_1446_0 & ~i_8_176_1911_0 & ~i_8_176_1922_0 & ~i_8_176_2195_0 & ~i_8_176_2291_0))) | (~i_8_176_78_0 & ~i_8_176_191_0 & i_8_176_691_0 & ~i_8_176_698_0 & ~i_8_176_1446_0 & ~i_8_176_1916_0 & ~i_8_176_1985_0 & ~i_8_176_2060_0) | (~i_8_176_717_0 & i_8_176_995_0 & ~i_8_176_1205_0 & ~i_8_176_1306_0 & ~i_8_176_1798_0 & ~i_8_176_2195_0 & ~i_8_176_2226_0))) | (~i_8_176_674_0 & ((~i_8_176_84_0 & ((~i_8_176_462_0 & i_8_176_991_0 & ~i_8_176_1797_0 & ~i_8_176_2195_0) | (~i_8_176_87_0 & ~i_8_176_395_0 & i_8_176_1047_0 & ~i_8_176_1385_0 & ~i_8_176_1446_0 & ~i_8_176_1911_0 & ~i_8_176_2053_0 & ~i_8_176_2060_0 & ~i_8_176_2100_0 & ~i_8_176_2291_0))) | (~i_8_176_191_0 & ((~i_8_176_267_0 & i_8_176_2100_0 & ((~i_8_176_87_0 & ~i_8_176_285_0 & ~i_8_176_599_0 & ~i_8_176_673_0 & ~i_8_176_927_0 & ~i_8_176_1205_0 & ~i_8_176_1306_0 & ~i_8_176_1385_0 & ~i_8_176_1446_0 & ~i_8_176_1911_0 & ~i_8_176_1985_0) | (~i_8_176_736_0 & i_8_176_991_0 & ~i_8_176_1365_0 & ~i_8_176_1547_0 & ~i_8_176_2193_0))) | (~i_8_176_78_0 & ~i_8_176_230_0 & ~i_8_176_489_0 & ~i_8_176_825_0 & i_8_176_838_0 & ~i_8_176_1306_0 & ~i_8_176_1797_0 & ~i_8_176_1844_0 & ~i_8_176_2053_0 & ~i_8_176_2195_0 & ~i_8_176_2226_0))) | (~i_8_176_462_0 & ~i_8_176_2193_0 & ((~i_8_176_264_0 & i_8_176_1056_0 & ~i_8_176_1385_0 & ~i_8_176_1457_0 & ~i_8_176_1797_0 & ~i_8_176_1798_0 & ~i_8_176_1911_0) | (~i_8_176_698_0 & ~i_8_176_1056_0 & ~i_8_176_1315_0 & i_8_176_2060_0 & ~i_8_176_2069_0))))) | (~i_8_176_489_0 & ~i_8_176_2055_0 & ((~i_8_176_230_0 & ~i_8_176_462_0 & ~i_8_176_737_0 & ~i_8_176_1446_0 & ~i_8_176_1547_0 & ~i_8_176_1844_0 & ~i_8_176_2069_0 & ~i_8_176_2100_0 & i_8_176_2156_0 & ~i_8_176_2195_0) | (~i_8_176_7_0 & i_8_176_135_0 & ~i_8_176_464_0 & ~i_8_176_673_0 & ~i_8_176_719_0 & ~i_8_176_1315_0 & ~i_8_176_1365_0 & ~i_8_176_2145_0 & ~i_8_176_2226_0 & ~i_8_176_2291_0))) | (~i_8_176_1131_0 & ((~i_8_176_7_0 & ((~i_8_176_264_0 & ~i_8_176_464_0 & ~i_8_176_553_0 & ~i_8_176_927_0 & ~i_8_176_1203_0 & ~i_8_176_1446_0 & i_8_176_1983_0) | (~i_8_176_592_0 & ~i_8_176_673_0 & ~i_8_176_825_0 & ~i_8_176_1797_0 & ~i_8_176_1798_0 & ~i_8_176_1911_0 & ~i_8_176_1916_0 & ~i_8_176_1918_0 & i_8_176_2156_0 & ~i_8_176_2195_0))) | (~i_8_176_462_0 & ~i_8_176_1204_0 & ~i_8_176_2193_0 & ((i_8_176_489_0 & ~i_8_176_553_0 & ~i_8_176_556_0 & ~i_8_176_719_0 & ~i_8_176_1056_0 & ~i_8_176_1203_0 & ~i_8_176_1306_0 & ~i_8_176_1446_0 & ~i_8_176_1985_0) | (~i_8_176_1133_0 & i_8_176_1985_0 & ~i_8_176_2195_0 & ~i_8_176_2263_0))))) | (~i_8_176_264_0 & ((~i_8_176_340_0 & ~i_8_176_599_0 & ~i_8_176_1132_0 & ~i_8_176_1985_0 & i_8_176_2005_0) | (~i_8_176_285_0 & i_8_176_838_0 & i_8_176_1047_0 & ~i_8_176_1203_0 & ~i_8_176_1385_0 & ~i_8_176_2069_0 & ~i_8_176_2193_0))) | (~i_8_176_599_0 & ((~i_8_176_673_0 & ((~i_8_176_285_0 & ~i_8_176_1132_0 & ((~i_8_176_340_0 & ~i_8_176_462_0 & ~i_8_176_592_0 & ~i_8_176_1446_0 & i_8_176_2175_0) | (~i_8_176_381_0 & ~i_8_176_1133_0 & i_8_176_1315_0 & ~i_8_176_1911_0 & ~i_8_176_2053_0 & ~i_8_176_2069_0 & ~i_8_176_2193_0))) | (~i_8_176_35_0 & ~i_8_176_87_0 & i_8_176_242_0 & ~i_8_176_2195_0 & ~i_8_176_2263_0 & ~i_8_176_825_0 & ~i_8_176_2193_0))) | (~i_8_176_78_0 & ~i_8_176_191_0 & ~i_8_176_395_0 & ~i_8_176_462_0 & ~i_8_176_556_0 & ~i_8_176_719_0 & ~i_8_176_825_0 & ~i_8_176_1205_0 & ~i_8_176_1266_0 & ~i_8_176_2195_0 & ~i_8_176_2291_0 & ~i_8_176_1918_0 & ~i_8_176_2156_0))) | (~i_8_176_78_0 & ~i_8_176_395_0 & ((~i_8_176_87_0 & i_8_176_88_0 & ~i_8_176_737_0 & ~i_8_176_995_0 & i_8_176_1922_0 & ~i_8_176_2145_0 & ~i_8_176_2156_0) | (~i_8_176_260_0 & ~i_8_176_825_0 & ~i_8_176_971_0 & ~i_8_176_1203_0 & ~i_8_176_1205_0 & ~i_8_176_1236_0 & ~i_8_176_1911_0 & ~i_8_176_1918_0 & ~i_8_176_2193_0 & ~i_8_176_2195_0))) | (~i_8_176_719_0 & ((~i_8_176_993_0 & i_8_176_2263_0 & i_8_176_2291_0) | (~i_8_176_895_0 & ~i_8_176_927_0 & ~i_8_176_1139_0 & ~i_8_176_1203_0 & ~i_8_176_1205_0 & ~i_8_176_1315_0 & i_8_176_1981_0 & ~i_8_176_2175_0 & ~i_8_176_2291_0))) | (i_8_176_998_0 & ((~i_8_176_340_0 & ~i_8_176_464_0 & ~i_8_176_592_0 & ~i_8_176_1204_0 & ~i_8_176_1606_0 & ~i_8_176_1916_0 & ~i_8_176_1205_0 & ~i_8_176_1315_0) | (~i_8_176_673_0 & i_8_176_1457_0 & ~i_8_176_1798_0 & ~i_8_176_1981_0 & ~i_8_176_2060_0 & ~i_8_176_2226_0))) | (~i_8_176_464_0 & ((i_8_176_230_0 & i_8_176_737_0 & ~i_8_176_1205_0 & ~i_8_176_1798_0 & ~i_8_176_1916_0 & ~i_8_176_1922_0) | (~i_8_176_825_0 & i_8_176_993_0 & i_8_176_1983_0))) | (~i_8_176_2069_0 & ((~i_8_176_462_0 & i_8_176_997_0 & ~i_8_176_1203_0 & ~i_8_176_1205_0 & ~i_8_176_1446_0 & ~i_8_176_1457_0 & ~i_8_176_1606_0) | (~i_8_176_2145_0 & ~i_8_176_2156_0 & i_8_176_1047_0 & i_8_176_1266_0))) | (~i_8_176_87_0 & i_8_176_994_0 & ~i_8_176_1133_0 & ~i_8_176_1911_0 & ~i_8_176_1916_0 & ~i_8_176_1236_0 & ~i_8_176_1797_0));
endmodule



// Benchmark "kernel_8_177" written by ABC on Sun Jul 19 10:06:07 2020

module kernel_8_177 ( 
    i_8_177_54_0, i_8_177_77_0, i_8_177_242_0, i_8_177_256_0,
    i_8_177_329_0, i_8_177_337_0, i_8_177_344_0, i_8_177_347_0,
    i_8_177_377_0, i_8_177_480_0, i_8_177_483_0, i_8_177_523_0,
    i_8_177_525_0, i_8_177_527_0, i_8_177_553_0, i_8_177_608_0,
    i_8_177_634_0, i_8_177_672_0, i_8_177_679_0, i_8_177_688_0,
    i_8_177_689_0, i_8_177_760_0, i_8_177_762_0, i_8_177_763_0,
    i_8_177_764_0, i_8_177_787_0, i_8_177_796_0, i_8_177_930_0,
    i_8_177_944_0, i_8_177_986_0, i_8_177_1030_0, i_8_177_1048_0,
    i_8_177_1049_0, i_8_177_1050_0, i_8_177_1051_0, i_8_177_1093_0,
    i_8_177_1112_0, i_8_177_1124_0, i_8_177_1227_0, i_8_177_1229_0,
    i_8_177_1236_0, i_8_177_1237_0, i_8_177_1268_0, i_8_177_1274_0,
    i_8_177_1281_0, i_8_177_1286_0, i_8_177_1295_0, i_8_177_1305_0,
    i_8_177_1307_0, i_8_177_1309_0, i_8_177_1317_0, i_8_177_1323_0,
    i_8_177_1328_0, i_8_177_1412_0, i_8_177_1435_0, i_8_177_1439_0,
    i_8_177_1537_0, i_8_177_1546_0, i_8_177_1547_0, i_8_177_1624_0,
    i_8_177_1643_0, i_8_177_1651_0, i_8_177_1679_0, i_8_177_1682_0,
    i_8_177_1696_0, i_8_177_1700_0, i_8_177_1720_0, i_8_177_1723_0,
    i_8_177_1724_0, i_8_177_1733_0, i_8_177_1742_0, i_8_177_1744_0,
    i_8_177_1745_0, i_8_177_1749_0, i_8_177_1750_0, i_8_177_1762_0,
    i_8_177_1763_0, i_8_177_1822_0, i_8_177_1832_0, i_8_177_1876_0,
    i_8_177_1877_0, i_8_177_1889_0, i_8_177_1903_0, i_8_177_1981_0,
    i_8_177_1984_0, i_8_177_1985_0, i_8_177_2041_0, i_8_177_2048_0,
    i_8_177_2057_0, i_8_177_2075_0, i_8_177_2084_0, i_8_177_2093_0,
    i_8_177_2148_0, i_8_177_2158_0, i_8_177_2164_0, i_8_177_2174_0,
    i_8_177_2216_0, i_8_177_2219_0, i_8_177_2230_0, i_8_177_2263_0,
    o_8_177_0_0  );
  input  i_8_177_54_0, i_8_177_77_0, i_8_177_242_0, i_8_177_256_0,
    i_8_177_329_0, i_8_177_337_0, i_8_177_344_0, i_8_177_347_0,
    i_8_177_377_0, i_8_177_480_0, i_8_177_483_0, i_8_177_523_0,
    i_8_177_525_0, i_8_177_527_0, i_8_177_553_0, i_8_177_608_0,
    i_8_177_634_0, i_8_177_672_0, i_8_177_679_0, i_8_177_688_0,
    i_8_177_689_0, i_8_177_760_0, i_8_177_762_0, i_8_177_763_0,
    i_8_177_764_0, i_8_177_787_0, i_8_177_796_0, i_8_177_930_0,
    i_8_177_944_0, i_8_177_986_0, i_8_177_1030_0, i_8_177_1048_0,
    i_8_177_1049_0, i_8_177_1050_0, i_8_177_1051_0, i_8_177_1093_0,
    i_8_177_1112_0, i_8_177_1124_0, i_8_177_1227_0, i_8_177_1229_0,
    i_8_177_1236_0, i_8_177_1237_0, i_8_177_1268_0, i_8_177_1274_0,
    i_8_177_1281_0, i_8_177_1286_0, i_8_177_1295_0, i_8_177_1305_0,
    i_8_177_1307_0, i_8_177_1309_0, i_8_177_1317_0, i_8_177_1323_0,
    i_8_177_1328_0, i_8_177_1412_0, i_8_177_1435_0, i_8_177_1439_0,
    i_8_177_1537_0, i_8_177_1546_0, i_8_177_1547_0, i_8_177_1624_0,
    i_8_177_1643_0, i_8_177_1651_0, i_8_177_1679_0, i_8_177_1682_0,
    i_8_177_1696_0, i_8_177_1700_0, i_8_177_1720_0, i_8_177_1723_0,
    i_8_177_1724_0, i_8_177_1733_0, i_8_177_1742_0, i_8_177_1744_0,
    i_8_177_1745_0, i_8_177_1749_0, i_8_177_1750_0, i_8_177_1762_0,
    i_8_177_1763_0, i_8_177_1822_0, i_8_177_1832_0, i_8_177_1876_0,
    i_8_177_1877_0, i_8_177_1889_0, i_8_177_1903_0, i_8_177_1981_0,
    i_8_177_1984_0, i_8_177_1985_0, i_8_177_2041_0, i_8_177_2048_0,
    i_8_177_2057_0, i_8_177_2075_0, i_8_177_2084_0, i_8_177_2093_0,
    i_8_177_2148_0, i_8_177_2158_0, i_8_177_2164_0, i_8_177_2174_0,
    i_8_177_2216_0, i_8_177_2219_0, i_8_177_2230_0, i_8_177_2263_0;
  output o_8_177_0_0;
  assign o_8_177_0_0 = 0;
endmodule



// Benchmark "kernel_8_178" written by ABC on Sun Jul 19 10:06:08 2020

module kernel_8_178 ( 
    i_8_178_14_0, i_8_178_31_0, i_8_178_32_0, i_8_178_51_0, i_8_178_52_0,
    i_8_178_55_0, i_8_178_59_0, i_8_178_77_0, i_8_178_201_0, i_8_178_229_0,
    i_8_178_255_0, i_8_178_256_0, i_8_178_378_0, i_8_178_385_0,
    i_8_178_387_0, i_8_178_388_0, i_8_178_390_0, i_8_178_391_0,
    i_8_178_392_0, i_8_178_415_0, i_8_178_417_0, i_8_178_426_0,
    i_8_178_450_0, i_8_178_493_0, i_8_178_508_0, i_8_178_509_0,
    i_8_178_534_0, i_8_178_536_0, i_8_178_608_0, i_8_178_630_0,
    i_8_178_634_0, i_8_178_658_0, i_8_178_676_0, i_8_178_748_0,
    i_8_178_750_0, i_8_178_752_0, i_8_178_880_0, i_8_178_1010_0,
    i_8_178_1030_0, i_8_178_1127_0, i_8_178_1128_0, i_8_178_1129_0,
    i_8_178_1130_0, i_8_178_1200_0, i_8_178_1228_0, i_8_178_1234_0,
    i_8_178_1261_0, i_8_178_1282_0, i_8_178_1289_0, i_8_178_1328_0,
    i_8_178_1355_0, i_8_178_1358_0, i_8_178_1385_0, i_8_178_1405_0,
    i_8_178_1476_0, i_8_178_1477_0, i_8_178_1478_0, i_8_178_1479_0,
    i_8_178_1480_0, i_8_178_1486_0, i_8_178_1490_0, i_8_178_1506_0,
    i_8_178_1510_0, i_8_178_1540_0, i_8_178_1548_0, i_8_178_1550_0,
    i_8_178_1559_0, i_8_178_1603_0, i_8_178_1605_0, i_8_178_1607_0,
    i_8_178_1627_0, i_8_178_1677_0, i_8_178_1713_0, i_8_178_1810_0,
    i_8_178_1813_0, i_8_178_1822_0, i_8_178_1836_0, i_8_178_1841_0,
    i_8_178_1873_0, i_8_178_1882_0, i_8_178_1890_0, i_8_178_1891_0,
    i_8_178_1892_0, i_8_178_1893_0, i_8_178_1894_0, i_8_178_1895_0,
    i_8_178_1939_0, i_8_178_1984_0, i_8_178_1996_0, i_8_178_2053_0,
    i_8_178_2057_0, i_8_178_2089_0, i_8_178_2146_0, i_8_178_2147_0,
    i_8_178_2150_0, i_8_178_2151_0, i_8_178_2155_0, i_8_178_2261_0,
    i_8_178_2263_0, i_8_178_2276_0,
    o_8_178_0_0  );
  input  i_8_178_14_0, i_8_178_31_0, i_8_178_32_0, i_8_178_51_0,
    i_8_178_52_0, i_8_178_55_0, i_8_178_59_0, i_8_178_77_0, i_8_178_201_0,
    i_8_178_229_0, i_8_178_255_0, i_8_178_256_0, i_8_178_378_0,
    i_8_178_385_0, i_8_178_387_0, i_8_178_388_0, i_8_178_390_0,
    i_8_178_391_0, i_8_178_392_0, i_8_178_415_0, i_8_178_417_0,
    i_8_178_426_0, i_8_178_450_0, i_8_178_493_0, i_8_178_508_0,
    i_8_178_509_0, i_8_178_534_0, i_8_178_536_0, i_8_178_608_0,
    i_8_178_630_0, i_8_178_634_0, i_8_178_658_0, i_8_178_676_0,
    i_8_178_748_0, i_8_178_750_0, i_8_178_752_0, i_8_178_880_0,
    i_8_178_1010_0, i_8_178_1030_0, i_8_178_1127_0, i_8_178_1128_0,
    i_8_178_1129_0, i_8_178_1130_0, i_8_178_1200_0, i_8_178_1228_0,
    i_8_178_1234_0, i_8_178_1261_0, i_8_178_1282_0, i_8_178_1289_0,
    i_8_178_1328_0, i_8_178_1355_0, i_8_178_1358_0, i_8_178_1385_0,
    i_8_178_1405_0, i_8_178_1476_0, i_8_178_1477_0, i_8_178_1478_0,
    i_8_178_1479_0, i_8_178_1480_0, i_8_178_1486_0, i_8_178_1490_0,
    i_8_178_1506_0, i_8_178_1510_0, i_8_178_1540_0, i_8_178_1548_0,
    i_8_178_1550_0, i_8_178_1559_0, i_8_178_1603_0, i_8_178_1605_0,
    i_8_178_1607_0, i_8_178_1627_0, i_8_178_1677_0, i_8_178_1713_0,
    i_8_178_1810_0, i_8_178_1813_0, i_8_178_1822_0, i_8_178_1836_0,
    i_8_178_1841_0, i_8_178_1873_0, i_8_178_1882_0, i_8_178_1890_0,
    i_8_178_1891_0, i_8_178_1892_0, i_8_178_1893_0, i_8_178_1894_0,
    i_8_178_1895_0, i_8_178_1939_0, i_8_178_1984_0, i_8_178_1996_0,
    i_8_178_2053_0, i_8_178_2057_0, i_8_178_2089_0, i_8_178_2146_0,
    i_8_178_2147_0, i_8_178_2150_0, i_8_178_2151_0, i_8_178_2155_0,
    i_8_178_2261_0, i_8_178_2263_0, i_8_178_2276_0;
  output o_8_178_0_0;
  assign o_8_178_0_0 = ~((~i_8_178_1893_0 & ((~i_8_178_1892_0 & ((~i_8_178_77_0 & ((~i_8_178_14_0 & ~i_8_178_388_0 & ~i_8_178_534_0 & i_8_178_1030_0 & ~i_8_178_1234_0 & ~i_8_178_1328_0 & ~i_8_178_1479_0 & ~i_8_178_1548_0 & ~i_8_178_1822_0 & ~i_8_178_1894_0) | (~i_8_178_387_0 & ~i_8_178_417_0 & ~i_8_178_509_0 & ~i_8_178_752_0 & ~i_8_178_1261_0 & ~i_8_178_1385_0 & ~i_8_178_1506_0 & ~i_8_178_1550_0 & ~i_8_178_1627_0 & ~i_8_178_1813_0 & ~i_8_178_1836_0 & ~i_8_178_1841_0 & ~i_8_178_1890_0 & ~i_8_178_2146_0 & ~i_8_178_2147_0 & ~i_8_178_2151_0))) | (~i_8_178_387_0 & ~i_8_178_752_0 & ((~i_8_178_229_0 & ~i_8_178_256_0 & ~i_8_178_390_0 & ~i_8_178_536_0 & i_8_178_634_0 & ~i_8_178_1128_0 & ~i_8_178_1477_0 & ~i_8_178_1478_0 & ~i_8_178_1480_0 & ~i_8_178_1486_0 & ~i_8_178_1836_0) | (i_8_178_229_0 & ~i_8_178_392_0 & ~i_8_178_426_0 & ~i_8_178_534_0 & ~i_8_178_1890_0 & ~i_8_178_1894_0 & ~i_8_178_1939_0 & ~i_8_178_2147_0))))) | (~i_8_178_14_0 & ((~i_8_178_750_0 & ((~i_8_178_388_0 & ~i_8_178_1130_0 & ~i_8_178_1486_0 & ((~i_8_178_201_0 & ~i_8_178_387_0 & ~i_8_178_390_0 & ~i_8_178_391_0 & ~i_8_178_1127_0 & ~i_8_178_1358_0 & ~i_8_178_1506_0 & ~i_8_178_1607_0 & ~i_8_178_1890_0 & ~i_8_178_1996_0) | (~i_8_178_392_0 & ~i_8_178_534_0 & ~i_8_178_658_0 & ~i_8_178_748_0 & ~i_8_178_1010_0 & ~i_8_178_1030_0 & ~i_8_178_1355_0 & ~i_8_178_1540_0 & ~i_8_178_1548_0 & ~i_8_178_1810_0 & ~i_8_178_2146_0))) | (~i_8_178_51_0 & ~i_8_178_391_0 & ~i_8_178_536_0 & ~i_8_178_1010_0 & ~i_8_178_1385_0 & ~i_8_178_1405_0 & ~i_8_178_1510_0 & ~i_8_178_1548_0 & ~i_8_178_1822_0 & ~i_8_178_1836_0 & ~i_8_178_1895_0 & ~i_8_178_1996_0 & ~i_8_178_2089_0 & ~i_8_178_2147_0))) | (~i_8_178_390_0 & ~i_8_178_534_0 & ~i_8_178_630_0 & ~i_8_178_676_0 & i_8_178_1282_0 & ~i_8_178_1328_0 & i_8_178_1486_0 & ~i_8_178_2089_0 & ~i_8_178_2147_0))) | (~i_8_178_2146_0 & ((~i_8_178_388_0 & ~i_8_178_493_0 & ~i_8_178_1130_0 & ((~i_8_178_508_0 & ~i_8_178_534_0 & ~i_8_178_1200_0 & ~i_8_178_1282_0 & ~i_8_178_1355_0 & ~i_8_178_1476_0 & ~i_8_178_1478_0 & ~i_8_178_1486_0 & ~i_8_178_1490_0 & ~i_8_178_1510_0 & ~i_8_178_1540_0 & ~i_8_178_1836_0) | (~i_8_178_59_0 & ~i_8_178_378_0 & ~i_8_178_426_0 & ~i_8_178_630_0 & ~i_8_178_634_0 & ~i_8_178_750_0 & ~i_8_178_1127_0 & ~i_8_178_1129_0 & ~i_8_178_1228_0 & ~i_8_178_1550_0 & ~i_8_178_1605_0 & ~i_8_178_1813_0 & ~i_8_178_1890_0 & ~i_8_178_1891_0 & ~i_8_178_1894_0))) | (~i_8_178_1891_0 & ((~i_8_178_417_0 & ~i_8_178_534_0 & ~i_8_178_536_0 & ~i_8_178_608_0 & ~i_8_178_1127_0 & ~i_8_178_1228_0 & ~i_8_178_1328_0 & ~i_8_178_1358_0 & ~i_8_178_1405_0 & ~i_8_178_1479_0 & ~i_8_178_1486_0 & ~i_8_178_1890_0 & ~i_8_178_1996_0 & ~i_8_178_2151_0) | (~i_8_178_390_0 & ~i_8_178_509_0 & ~i_8_178_1550_0 & i_8_178_1677_0 & i_8_178_1984_0 & ~i_8_178_2147_0 & ~i_8_178_2263_0))))) | (~i_8_178_493_0 & ~i_8_178_536_0 & ~i_8_178_1128_0 & ~i_8_178_1129_0 & ~i_8_178_1477_0 & ~i_8_178_1479_0 & i_8_178_1510_0 & ~i_8_178_1540_0 & ~i_8_178_1550_0 & ~i_8_178_1713_0 & ~i_8_178_1836_0 & ~i_8_178_1895_0))) | (~i_8_178_1550_0 & ((~i_8_178_1478_0 & ((~i_8_178_14_0 & ~i_8_178_1490_0 & ((~i_8_178_229_0 & ~i_8_178_390_0 & ~i_8_178_608_0 & ~i_8_178_634_0 & ~i_8_178_880_0 & ~i_8_178_1128_0 & ~i_8_178_1476_0 & ~i_8_178_1479_0 & ~i_8_178_1822_0 & ~i_8_178_1841_0 & ~i_8_178_1882_0 & ~i_8_178_1891_0 & ~i_8_178_1894_0 & ~i_8_178_2089_0 & ~i_8_178_2155_0) | (~i_8_178_1010_0 & ~i_8_178_1200_0 & i_8_178_1328_0 & ~i_8_178_1548_0 & ~i_8_178_2276_0))) | (~i_8_178_390_0 & ~i_8_178_426_0 & ~i_8_178_750_0 & ~i_8_178_1128_0 & ~i_8_178_1129_0 & ~i_8_178_1130_0 & ~i_8_178_1328_0 & ~i_8_178_1355_0 & ~i_8_178_1358_0 & ~i_8_178_1476_0 & ~i_8_178_1477_0 & ~i_8_178_1479_0 & ~i_8_178_1510_0 & ~i_8_178_1548_0 & ~i_8_178_1892_0))) | (~i_8_178_387_0 & ((~i_8_178_536_0 & ((~i_8_178_390_0 & ~i_8_178_1510_0 & ((~i_8_178_255_0 & ~i_8_178_391_0 & ~i_8_178_392_0 & ~i_8_178_509_0 & ~i_8_178_750_0 & ~i_8_178_752_0 & ~i_8_178_1129_0 & ~i_8_178_1677_0 & ~i_8_178_1810_0 & ~i_8_178_1836_0 & ~i_8_178_1890_0 & ~i_8_178_1892_0 & ~i_8_178_2089_0) | (~i_8_178_388_0 & ~i_8_178_415_0 & ~i_8_178_534_0 & ~i_8_178_1127_0 & ~i_8_178_1128_0 & ~i_8_178_1385_0 & ~i_8_178_1405_0 & ~i_8_178_1479_0 & ~i_8_178_1841_0 & ~i_8_178_1894_0 & ~i_8_178_2147_0))) | (~i_8_178_391_0 & ~i_8_178_426_0 & ~i_8_178_493_0 & ~i_8_178_534_0 & ~i_8_178_1010_0 & ~i_8_178_1128_0 & ~i_8_178_1130_0 & ~i_8_178_1228_0 & ~i_8_178_1506_0 & ~i_8_178_1836_0 & ~i_8_178_1892_0 & ~i_8_178_2089_0))) | (i_8_178_426_0 & ~i_8_178_1010_0 & ~i_8_178_1127_0 & ~i_8_178_1130_0 & ~i_8_178_1200_0 & ~i_8_178_1477_0 & ~i_8_178_1479_0 & ~i_8_178_1490_0 & ~i_8_178_1506_0 & ~i_8_178_1836_0 & ~i_8_178_1894_0))) | (~i_8_178_229_0 & i_8_178_880_0 & ~i_8_178_1129_0 & ~i_8_178_1228_0 & ~i_8_178_1476_0 & i_8_178_2276_0))) | (~i_8_178_388_0 & ((~i_8_178_52_0 & i_8_178_229_0 & ~i_8_178_387_0 & i_8_178_634_0 & ~i_8_178_750_0 & ~i_8_178_1129_0 & ~i_8_178_1477_0) | (~i_8_178_1127_0 & ~i_8_178_1130_0 & ~i_8_178_1486_0 & ~i_8_178_1548_0 & i_8_178_1559_0 & ~i_8_178_1939_0))) | (~i_8_178_391_0 & i_8_178_493_0 & ((~i_8_178_748_0 & ~i_8_178_1010_0 & ~i_8_178_1490_0 & ~i_8_178_1892_0 & ~i_8_178_1894_0 & i_8_178_2057_0) | (~i_8_178_415_0 & ~i_8_178_534_0 & ~i_8_178_750_0 & ~i_8_178_1130_0 & ~i_8_178_1328_0 & ~i_8_178_1355_0 & ~i_8_178_1603_0 & ~i_8_178_1713_0 & ~i_8_178_2089_0))) | (~i_8_178_1130_0 & ((~i_8_178_1128_0 & ((~i_8_178_390_0 & ~i_8_178_1328_0 & ~i_8_178_1890_0 & ((~i_8_178_415_0 & ~i_8_178_426_0 & ~i_8_178_508_0 & ~i_8_178_534_0 & ~i_8_178_752_0 & ~i_8_178_1405_0 & ~i_8_178_1478_0 & ~i_8_178_1540_0 & ~i_8_178_1603_0 & ~i_8_178_1607_0) | (~i_8_178_385_0 & ~i_8_178_417_0 & i_8_178_880_0 & ~i_8_178_1228_0 & ~i_8_178_1355_0 & ~i_8_178_1477_0 & ~i_8_178_1479_0 & ~i_8_178_1892_0 & ~i_8_178_2276_0))) | (~i_8_178_55_0 & ~i_8_178_201_0 & ~i_8_178_387_0 & ~i_8_178_534_0 & ~i_8_178_536_0 & ~i_8_178_748_0 & ~i_8_178_752_0 & ~i_8_178_1030_0 & ~i_8_178_1355_0 & ~i_8_178_1479_0 & ~i_8_178_1540_0 & ~i_8_178_1605_0 & ~i_8_178_1822_0 & ~i_8_178_1892_0 & ~i_8_178_1996_0 & ~i_8_178_2155_0 & ~i_8_178_2263_0))) | (~i_8_178_748_0 & ~i_8_178_1010_0 & ~i_8_178_1200_0 & ((~i_8_178_392_0 & ~i_8_178_509_0 & ~i_8_178_750_0 & ~i_8_178_1328_0 & i_8_178_1355_0 & ~i_8_178_1479_0 & ~i_8_178_1480_0 & ~i_8_178_1540_0 & ~i_8_178_1713_0 & ~i_8_178_1892_0) | (~i_8_178_534_0 & ~i_8_178_1129_0 & ~i_8_178_1282_0 & ~i_8_178_1478_0 & ~i_8_178_1506_0 & ~i_8_178_1548_0 & ~i_8_178_1836_0 & ~i_8_178_1891_0 & ~i_8_178_1894_0 & i_8_178_2146_0))) | (~i_8_178_415_0 & ~i_8_178_1129_0 & i_8_178_1282_0 & ~i_8_178_1476_0 & ~i_8_178_1477_0 & ~i_8_178_1627_0 & i_8_178_1810_0 & ~i_8_178_1891_0 & ~i_8_178_1894_0 & ~i_8_178_2089_0))) | (~i_8_178_1895_0 & ((~i_8_178_387_0 & ((~i_8_178_534_0 & ~i_8_178_536_0 & ~i_8_178_750_0 & ~i_8_178_1010_0 & ~i_8_178_1127_0 & ~i_8_178_1129_0 & i_8_178_1261_0 & ~i_8_178_1478_0 & ~i_8_178_1540_0 & ~i_8_178_1605_0 & ~i_8_178_1873_0) | (~i_8_178_392_0 & i_8_178_880_0 & ~i_8_178_1128_0 & ~i_8_178_1476_0 & ~i_8_178_1486_0 & ~i_8_178_1894_0 & i_8_178_2151_0))) | (~i_8_178_390_0 & ~i_8_178_392_0 & ~i_8_178_534_0 & ~i_8_178_750_0 & ~i_8_178_1010_0 & ~i_8_178_1127_0 & ~i_8_178_1228_0 & ~i_8_178_1282_0 & ~i_8_178_1540_0 & ~i_8_178_1836_0 & ~i_8_178_1328_0 & ~i_8_178_1405_0 & ~i_8_178_1890_0 & ~i_8_178_1892_0 & ~i_8_178_1894_0 & ~i_8_178_2146_0 & ~i_8_178_2150_0))) | (~i_8_178_1128_0 & ((~i_8_178_390_0 & ~i_8_178_752_0 & ~i_8_178_1129_0 & ~i_8_178_1478_0 & ~i_8_178_1480_0 & ~i_8_178_1506_0 & i_8_178_1813_0 & ~i_8_178_1890_0) | (~i_8_178_1605_0 & i_8_178_1627_0 & ~i_8_178_1822_0 & i_8_178_1893_0))));
endmodule



// Benchmark "kernel_8_179" written by ABC on Sun Jul 19 10:06:09 2020

module kernel_8_179 ( 
    i_8_179_30_0, i_8_179_31_0, i_8_179_40_0, i_8_179_51_0, i_8_179_75_0,
    i_8_179_78_0, i_8_179_81_0, i_8_179_102_0, i_8_179_120_0,
    i_8_179_165_0, i_8_179_166_0, i_8_179_363_0, i_8_179_364_0,
    i_8_179_373_0, i_8_179_426_0, i_8_179_450_0, i_8_179_492_0,
    i_8_179_582_0, i_8_179_588_0, i_8_179_607_0, i_8_179_612_0,
    i_8_179_633_0, i_8_179_654_0, i_8_179_660_0, i_8_179_665_0,
    i_8_179_676_0, i_8_179_696_0, i_8_179_699_0, i_8_179_700_0,
    i_8_179_714_0, i_8_179_723_0, i_8_179_754_0, i_8_179_804_0,
    i_8_179_807_0, i_8_179_822_0, i_8_179_825_0, i_8_179_832_0,
    i_8_179_841_0, i_8_179_865_0, i_8_179_877_0, i_8_179_930_0,
    i_8_179_941_0, i_8_179_964_0, i_8_179_966_0, i_8_179_993_0,
    i_8_179_994_0, i_8_179_1050_0, i_8_179_1056_0, i_8_179_1065_0,
    i_8_179_1071_0, i_8_179_1093_0, i_8_179_1108_0, i_8_179_1111_0,
    i_8_179_1138_0, i_8_179_1182_0, i_8_179_1201_0, i_8_179_1217_0,
    i_8_179_1273_0, i_8_179_1281_0, i_8_179_1326_0, i_8_179_1337_0,
    i_8_179_1351_0, i_8_179_1359_0, i_8_179_1372_0, i_8_179_1386_0,
    i_8_179_1432_0, i_8_179_1515_0, i_8_179_1542_0, i_8_179_1545_0,
    i_8_179_1563_0, i_8_179_1565_0, i_8_179_1587_0, i_8_179_1621_0,
    i_8_179_1632_0, i_8_179_1668_0, i_8_179_1677_0, i_8_179_1698_0,
    i_8_179_1699_0, i_8_179_1704_0, i_8_179_1716_0, i_8_179_1747_0,
    i_8_179_1752_0, i_8_179_1804_0, i_8_179_1819_0, i_8_179_1821_0,
    i_8_179_1845_0, i_8_179_1946_0, i_8_179_1981_0, i_8_179_1992_0,
    i_8_179_1995_0, i_8_179_1997_0, i_8_179_2045_0, i_8_179_2115_0,
    i_8_179_2118_0, i_8_179_2146_0, i_8_179_2149_0, i_8_179_2190_0,
    i_8_179_2226_0, i_8_179_2235_0, i_8_179_2259_0,
    o_8_179_0_0  );
  input  i_8_179_30_0, i_8_179_31_0, i_8_179_40_0, i_8_179_51_0,
    i_8_179_75_0, i_8_179_78_0, i_8_179_81_0, i_8_179_102_0, i_8_179_120_0,
    i_8_179_165_0, i_8_179_166_0, i_8_179_363_0, i_8_179_364_0,
    i_8_179_373_0, i_8_179_426_0, i_8_179_450_0, i_8_179_492_0,
    i_8_179_582_0, i_8_179_588_0, i_8_179_607_0, i_8_179_612_0,
    i_8_179_633_0, i_8_179_654_0, i_8_179_660_0, i_8_179_665_0,
    i_8_179_676_0, i_8_179_696_0, i_8_179_699_0, i_8_179_700_0,
    i_8_179_714_0, i_8_179_723_0, i_8_179_754_0, i_8_179_804_0,
    i_8_179_807_0, i_8_179_822_0, i_8_179_825_0, i_8_179_832_0,
    i_8_179_841_0, i_8_179_865_0, i_8_179_877_0, i_8_179_930_0,
    i_8_179_941_0, i_8_179_964_0, i_8_179_966_0, i_8_179_993_0,
    i_8_179_994_0, i_8_179_1050_0, i_8_179_1056_0, i_8_179_1065_0,
    i_8_179_1071_0, i_8_179_1093_0, i_8_179_1108_0, i_8_179_1111_0,
    i_8_179_1138_0, i_8_179_1182_0, i_8_179_1201_0, i_8_179_1217_0,
    i_8_179_1273_0, i_8_179_1281_0, i_8_179_1326_0, i_8_179_1337_0,
    i_8_179_1351_0, i_8_179_1359_0, i_8_179_1372_0, i_8_179_1386_0,
    i_8_179_1432_0, i_8_179_1515_0, i_8_179_1542_0, i_8_179_1545_0,
    i_8_179_1563_0, i_8_179_1565_0, i_8_179_1587_0, i_8_179_1621_0,
    i_8_179_1632_0, i_8_179_1668_0, i_8_179_1677_0, i_8_179_1698_0,
    i_8_179_1699_0, i_8_179_1704_0, i_8_179_1716_0, i_8_179_1747_0,
    i_8_179_1752_0, i_8_179_1804_0, i_8_179_1819_0, i_8_179_1821_0,
    i_8_179_1845_0, i_8_179_1946_0, i_8_179_1981_0, i_8_179_1992_0,
    i_8_179_1995_0, i_8_179_1997_0, i_8_179_2045_0, i_8_179_2115_0,
    i_8_179_2118_0, i_8_179_2146_0, i_8_179_2149_0, i_8_179_2190_0,
    i_8_179_2226_0, i_8_179_2235_0, i_8_179_2259_0;
  output o_8_179_0_0;
  assign o_8_179_0_0 = 0;
endmodule



// Benchmark "kernel_8_180" written by ABC on Sun Jul 19 10:06:10 2020

module kernel_8_180 ( 
    i_8_180_39_0, i_8_180_76_0, i_8_180_85_0, i_8_180_138_0, i_8_180_139_0,
    i_8_180_169_0, i_8_180_183_0, i_8_180_190_0, i_8_180_222_0,
    i_8_180_226_0, i_8_180_300_0, i_8_180_318_0, i_8_180_333_0,
    i_8_180_360_0, i_8_180_363_0, i_8_180_382_0, i_8_180_384_0,
    i_8_180_389_0, i_8_180_400_0, i_8_180_507_0, i_8_180_508_0,
    i_8_180_510_0, i_8_180_525_0, i_8_180_571_0, i_8_180_591_0,
    i_8_180_606_0, i_8_180_631_0, i_8_180_659_0, i_8_180_672_0,
    i_8_180_678_0, i_8_180_679_0, i_8_180_695_0, i_8_180_697_0,
    i_8_180_841_0, i_8_180_844_0, i_8_180_876_0, i_8_180_895_0,
    i_8_180_955_0, i_8_180_1039_0, i_8_180_1056_0, i_8_180_1102_0,
    i_8_180_1105_0, i_8_180_1156_0, i_8_180_1166_0, i_8_180_1246_0,
    i_8_180_1276_0, i_8_180_1282_0, i_8_180_1304_0, i_8_180_1306_0,
    i_8_180_1317_0, i_8_180_1318_0, i_8_180_1321_0, i_8_180_1327_0,
    i_8_180_1330_0, i_8_180_1339_0, i_8_180_1383_0, i_8_180_1423_0,
    i_8_180_1426_0, i_8_180_1438_0, i_8_180_1461_0, i_8_180_1464_0,
    i_8_180_1506_0, i_8_180_1509_0, i_8_180_1511_0, i_8_180_1516_0,
    i_8_180_1519_0, i_8_180_1606_0, i_8_180_1630_0, i_8_180_1632_0,
    i_8_180_1633_0, i_8_180_1636_0, i_8_180_1642_0, i_8_180_1651_0,
    i_8_180_1681_0, i_8_180_1686_0, i_8_180_1687_0, i_8_180_1722_0,
    i_8_180_1723_0, i_8_180_1749_0, i_8_180_1770_0, i_8_180_1781_0,
    i_8_180_1794_0, i_8_180_1837_0, i_8_180_1849_0, i_8_180_1858_0,
    i_8_180_1890_0, i_8_180_1938_0, i_8_180_1939_0, i_8_180_1956_0,
    i_8_180_1957_0, i_8_180_1965_0, i_8_180_1996_0, i_8_180_2054_0,
    i_8_180_2059_0, i_8_180_2155_0, i_8_180_2174_0, i_8_180_2233_0,
    i_8_180_2244_0, i_8_180_2262_0, i_8_180_2272_0,
    o_8_180_0_0  );
  input  i_8_180_39_0, i_8_180_76_0, i_8_180_85_0, i_8_180_138_0,
    i_8_180_139_0, i_8_180_169_0, i_8_180_183_0, i_8_180_190_0,
    i_8_180_222_0, i_8_180_226_0, i_8_180_300_0, i_8_180_318_0,
    i_8_180_333_0, i_8_180_360_0, i_8_180_363_0, i_8_180_382_0,
    i_8_180_384_0, i_8_180_389_0, i_8_180_400_0, i_8_180_507_0,
    i_8_180_508_0, i_8_180_510_0, i_8_180_525_0, i_8_180_571_0,
    i_8_180_591_0, i_8_180_606_0, i_8_180_631_0, i_8_180_659_0,
    i_8_180_672_0, i_8_180_678_0, i_8_180_679_0, i_8_180_695_0,
    i_8_180_697_0, i_8_180_841_0, i_8_180_844_0, i_8_180_876_0,
    i_8_180_895_0, i_8_180_955_0, i_8_180_1039_0, i_8_180_1056_0,
    i_8_180_1102_0, i_8_180_1105_0, i_8_180_1156_0, i_8_180_1166_0,
    i_8_180_1246_0, i_8_180_1276_0, i_8_180_1282_0, i_8_180_1304_0,
    i_8_180_1306_0, i_8_180_1317_0, i_8_180_1318_0, i_8_180_1321_0,
    i_8_180_1327_0, i_8_180_1330_0, i_8_180_1339_0, i_8_180_1383_0,
    i_8_180_1423_0, i_8_180_1426_0, i_8_180_1438_0, i_8_180_1461_0,
    i_8_180_1464_0, i_8_180_1506_0, i_8_180_1509_0, i_8_180_1511_0,
    i_8_180_1516_0, i_8_180_1519_0, i_8_180_1606_0, i_8_180_1630_0,
    i_8_180_1632_0, i_8_180_1633_0, i_8_180_1636_0, i_8_180_1642_0,
    i_8_180_1651_0, i_8_180_1681_0, i_8_180_1686_0, i_8_180_1687_0,
    i_8_180_1722_0, i_8_180_1723_0, i_8_180_1749_0, i_8_180_1770_0,
    i_8_180_1781_0, i_8_180_1794_0, i_8_180_1837_0, i_8_180_1849_0,
    i_8_180_1858_0, i_8_180_1890_0, i_8_180_1938_0, i_8_180_1939_0,
    i_8_180_1956_0, i_8_180_1957_0, i_8_180_1965_0, i_8_180_1996_0,
    i_8_180_2054_0, i_8_180_2059_0, i_8_180_2155_0, i_8_180_2174_0,
    i_8_180_2233_0, i_8_180_2244_0, i_8_180_2262_0, i_8_180_2272_0;
  output o_8_180_0_0;
  assign o_8_180_0_0 = ~((~i_8_180_139_0 & ((~i_8_180_1426_0 & ~i_8_180_1686_0 & ~i_8_180_1770_0) | (i_8_180_841_0 & ~i_8_180_1630_0 & ~i_8_180_1749_0 & ~i_8_180_1938_0))) | (~i_8_180_400_0 & ((~i_8_180_76_0 & ~i_8_180_571_0 & ~i_8_180_955_0 & ~i_8_180_1102_0 & ~i_8_180_1105_0 & ~i_8_180_1304_0 & ~i_8_180_1642_0) | (~i_8_180_508_0 & ~i_8_180_1506_0 & ~i_8_180_1509_0 & ~i_8_180_1722_0))) | (~i_8_180_510_0 & ((~i_8_180_507_0 & ~i_8_180_508_0 & ~i_8_180_2174_0) | (~i_8_180_138_0 & ~i_8_180_679_0 & i_8_180_2272_0))) | (~i_8_180_1318_0 & ((~i_8_180_1039_0 & ~i_8_180_1321_0 & ~i_8_180_1327_0 & ~i_8_180_1519_0 & ~i_8_180_1939_0) | (~i_8_180_39_0 & ~i_8_180_318_0 & ~i_8_180_1156_0 & ~i_8_180_1957_0))) | (~i_8_180_1330_0 & ((~i_8_180_1105_0 & ~i_8_180_1321_0 & ~i_8_180_1423_0 & ~i_8_180_1461_0 & ~i_8_180_1636_0) | (~i_8_180_571_0 & ~i_8_180_1438_0 & ~i_8_180_1511_0 & i_8_180_1633_0 & ~i_8_180_1722_0 & i_8_180_1996_0))) | (~i_8_180_895_0 & i_8_180_1321_0 & ~i_8_180_1339_0 & ~i_8_180_1423_0 & ~i_8_180_1461_0) | (~i_8_180_1317_0 & ~i_8_180_1516_0 & ~i_8_180_1686_0 & ~i_8_180_1837_0 & ~i_8_180_1956_0) | (~i_8_180_333_0 & ~i_8_180_1276_0 & ~i_8_180_1304_0 & ~i_8_180_1509_0 & ~i_8_180_1511_0 & ~i_8_180_1519_0 & ~i_8_180_1632_0 & ~i_8_180_2174_0) | (i_8_180_1858_0 & i_8_180_2262_0));
endmodule



// Benchmark "kernel_8_181" written by ABC on Sun Jul 19 10:06:11 2020

module kernel_8_181 ( 
    i_8_181_38_0, i_8_181_65_0, i_8_181_86_0, i_8_181_143_0, i_8_181_163_0,
    i_8_181_184_0, i_8_181_190_0, i_8_181_230_0, i_8_181_300_0,
    i_8_181_305_0, i_8_181_334_0, i_8_181_347_0, i_8_181_362_0,
    i_8_181_364_0, i_8_181_382_0, i_8_181_416_0, i_8_181_429_0,
    i_8_181_442_0, i_8_181_451_0, i_8_181_454_0, i_8_181_493_0,
    i_8_181_524_0, i_8_181_536_0, i_8_181_572_0, i_8_181_611_0,
    i_8_181_653_0, i_8_181_658_0, i_8_181_662_0, i_8_181_665_0,
    i_8_181_680_0, i_8_181_693_0, i_8_181_696_0, i_8_181_698_0,
    i_8_181_699_0, i_8_181_704_0, i_8_181_706_0, i_8_181_710_0,
    i_8_181_716_0, i_8_181_751_0, i_8_181_773_0, i_8_181_799_0,
    i_8_181_823_0, i_8_181_850_0, i_8_181_866_0, i_8_181_881_0,
    i_8_181_964_0, i_8_181_965_0, i_8_181_967_0, i_8_181_977_0,
    i_8_181_1103_0, i_8_181_1180_0, i_8_181_1181_0, i_8_181_1192_0,
    i_8_181_1198_0, i_8_181_1226_0, i_8_181_1247_0, i_8_181_1266_0,
    i_8_181_1267_0, i_8_181_1283_0, i_8_181_1289_0, i_8_181_1295_0,
    i_8_181_1318_0, i_8_181_1328_0, i_8_181_1344_0, i_8_181_1364_0,
    i_8_181_1372_0, i_8_181_1400_0, i_8_181_1403_0, i_8_181_1404_0,
    i_8_181_1408_0, i_8_181_1410_0, i_8_181_1438_0, i_8_181_1450_0,
    i_8_181_1453_0, i_8_181_1562_0, i_8_181_1564_0, i_8_181_1655_0,
    i_8_181_1681_0, i_8_181_1690_0, i_8_181_1706_0, i_8_181_1777_0,
    i_8_181_1780_0, i_8_181_1784_0, i_8_181_1792_0, i_8_181_1825_0,
    i_8_181_1886_0, i_8_181_1903_0, i_8_181_1907_0, i_8_181_1975_0,
    i_8_181_1981_0, i_8_181_1993_0, i_8_181_1996_0, i_8_181_2056_0,
    i_8_181_2075_0, i_8_181_2146_0, i_8_181_2156_0, i_8_181_2165_0,
    i_8_181_2197_0, i_8_181_2229_0, i_8_181_2257_0,
    o_8_181_0_0  );
  input  i_8_181_38_0, i_8_181_65_0, i_8_181_86_0, i_8_181_143_0,
    i_8_181_163_0, i_8_181_184_0, i_8_181_190_0, i_8_181_230_0,
    i_8_181_300_0, i_8_181_305_0, i_8_181_334_0, i_8_181_347_0,
    i_8_181_362_0, i_8_181_364_0, i_8_181_382_0, i_8_181_416_0,
    i_8_181_429_0, i_8_181_442_0, i_8_181_451_0, i_8_181_454_0,
    i_8_181_493_0, i_8_181_524_0, i_8_181_536_0, i_8_181_572_0,
    i_8_181_611_0, i_8_181_653_0, i_8_181_658_0, i_8_181_662_0,
    i_8_181_665_0, i_8_181_680_0, i_8_181_693_0, i_8_181_696_0,
    i_8_181_698_0, i_8_181_699_0, i_8_181_704_0, i_8_181_706_0,
    i_8_181_710_0, i_8_181_716_0, i_8_181_751_0, i_8_181_773_0,
    i_8_181_799_0, i_8_181_823_0, i_8_181_850_0, i_8_181_866_0,
    i_8_181_881_0, i_8_181_964_0, i_8_181_965_0, i_8_181_967_0,
    i_8_181_977_0, i_8_181_1103_0, i_8_181_1180_0, i_8_181_1181_0,
    i_8_181_1192_0, i_8_181_1198_0, i_8_181_1226_0, i_8_181_1247_0,
    i_8_181_1266_0, i_8_181_1267_0, i_8_181_1283_0, i_8_181_1289_0,
    i_8_181_1295_0, i_8_181_1318_0, i_8_181_1328_0, i_8_181_1344_0,
    i_8_181_1364_0, i_8_181_1372_0, i_8_181_1400_0, i_8_181_1403_0,
    i_8_181_1404_0, i_8_181_1408_0, i_8_181_1410_0, i_8_181_1438_0,
    i_8_181_1450_0, i_8_181_1453_0, i_8_181_1562_0, i_8_181_1564_0,
    i_8_181_1655_0, i_8_181_1681_0, i_8_181_1690_0, i_8_181_1706_0,
    i_8_181_1777_0, i_8_181_1780_0, i_8_181_1784_0, i_8_181_1792_0,
    i_8_181_1825_0, i_8_181_1886_0, i_8_181_1903_0, i_8_181_1907_0,
    i_8_181_1975_0, i_8_181_1981_0, i_8_181_1993_0, i_8_181_1996_0,
    i_8_181_2056_0, i_8_181_2075_0, i_8_181_2146_0, i_8_181_2156_0,
    i_8_181_2165_0, i_8_181_2197_0, i_8_181_2229_0, i_8_181_2257_0;
  output o_8_181_0_0;
  assign o_8_181_0_0 = 0;
endmodule



// Benchmark "kernel_8_182" written by ABC on Sun Jul 19 10:06:13 2020

module kernel_8_182 ( 
    i_8_182_0_0, i_8_182_1_0, i_8_182_3_0, i_8_182_73_0, i_8_182_81_0,
    i_8_182_82_0, i_8_182_111_0, i_8_182_112_0, i_8_182_153_0,
    i_8_182_198_0, i_8_182_227_0, i_8_182_243_0, i_8_182_279_0,
    i_8_182_283_0, i_8_182_318_0, i_8_182_342_0, i_8_182_345_0,
    i_8_182_363_0, i_8_182_364_0, i_8_182_434_0, i_8_182_436_0,
    i_8_182_450_0, i_8_182_486_0, i_8_182_568_0, i_8_182_604_0,
    i_8_182_626_0, i_8_182_630_0, i_8_182_666_0, i_8_182_673_0,
    i_8_182_705_0, i_8_182_710_0, i_8_182_729_0, i_8_182_811_0,
    i_8_182_829_0, i_8_182_832_0, i_8_182_833_0, i_8_182_865_0,
    i_8_182_892_0, i_8_182_992_0, i_8_182_1028_0, i_8_182_1030_0,
    i_8_182_1033_0, i_8_182_1035_0, i_8_182_1081_0, i_8_182_1091_0,
    i_8_182_1172_0, i_8_182_1182_0, i_8_182_1198_0, i_8_182_1228_0,
    i_8_182_1233_0, i_8_182_1270_0, i_8_182_1293_0, i_8_182_1296_0,
    i_8_182_1299_0, i_8_182_1314_0, i_8_182_1351_0, i_8_182_1386_0,
    i_8_182_1404_0, i_8_182_1434_0, i_8_182_1506_0, i_8_182_1561_0,
    i_8_182_1587_0, i_8_182_1633_0, i_8_182_1641_0, i_8_182_1677_0,
    i_8_182_1720_0, i_8_182_1746_0, i_8_182_1749_0, i_8_182_1777_0,
    i_8_182_1780_0, i_8_182_1791_0, i_8_182_1801_0, i_8_182_1804_0,
    i_8_182_1813_0, i_8_182_1845_0, i_8_182_1846_0, i_8_182_1881_0,
    i_8_182_1890_0, i_8_182_1893_0, i_8_182_1912_0, i_8_182_1923_0,
    i_8_182_1935_0, i_8_182_1966_0, i_8_182_1971_0, i_8_182_1980_0,
    i_8_182_1992_0, i_8_182_2025_0, i_8_182_2034_0, i_8_182_2035_0,
    i_8_182_2055_0, i_8_182_2074_0, i_8_182_2115_0, i_8_182_2116_0,
    i_8_182_2128_0, i_8_182_2133_0, i_8_182_2134_0, i_8_182_2142_0,
    i_8_182_2145_0, i_8_182_2157_0, i_8_182_2274_0,
    o_8_182_0_0  );
  input  i_8_182_0_0, i_8_182_1_0, i_8_182_3_0, i_8_182_73_0,
    i_8_182_81_0, i_8_182_82_0, i_8_182_111_0, i_8_182_112_0,
    i_8_182_153_0, i_8_182_198_0, i_8_182_227_0, i_8_182_243_0,
    i_8_182_279_0, i_8_182_283_0, i_8_182_318_0, i_8_182_342_0,
    i_8_182_345_0, i_8_182_363_0, i_8_182_364_0, i_8_182_434_0,
    i_8_182_436_0, i_8_182_450_0, i_8_182_486_0, i_8_182_568_0,
    i_8_182_604_0, i_8_182_626_0, i_8_182_630_0, i_8_182_666_0,
    i_8_182_673_0, i_8_182_705_0, i_8_182_710_0, i_8_182_729_0,
    i_8_182_811_0, i_8_182_829_0, i_8_182_832_0, i_8_182_833_0,
    i_8_182_865_0, i_8_182_892_0, i_8_182_992_0, i_8_182_1028_0,
    i_8_182_1030_0, i_8_182_1033_0, i_8_182_1035_0, i_8_182_1081_0,
    i_8_182_1091_0, i_8_182_1172_0, i_8_182_1182_0, i_8_182_1198_0,
    i_8_182_1228_0, i_8_182_1233_0, i_8_182_1270_0, i_8_182_1293_0,
    i_8_182_1296_0, i_8_182_1299_0, i_8_182_1314_0, i_8_182_1351_0,
    i_8_182_1386_0, i_8_182_1404_0, i_8_182_1434_0, i_8_182_1506_0,
    i_8_182_1561_0, i_8_182_1587_0, i_8_182_1633_0, i_8_182_1641_0,
    i_8_182_1677_0, i_8_182_1720_0, i_8_182_1746_0, i_8_182_1749_0,
    i_8_182_1777_0, i_8_182_1780_0, i_8_182_1791_0, i_8_182_1801_0,
    i_8_182_1804_0, i_8_182_1813_0, i_8_182_1845_0, i_8_182_1846_0,
    i_8_182_1881_0, i_8_182_1890_0, i_8_182_1893_0, i_8_182_1912_0,
    i_8_182_1923_0, i_8_182_1935_0, i_8_182_1966_0, i_8_182_1971_0,
    i_8_182_1980_0, i_8_182_1992_0, i_8_182_2025_0, i_8_182_2034_0,
    i_8_182_2035_0, i_8_182_2055_0, i_8_182_2074_0, i_8_182_2115_0,
    i_8_182_2116_0, i_8_182_2128_0, i_8_182_2133_0, i_8_182_2134_0,
    i_8_182_2142_0, i_8_182_2145_0, i_8_182_2157_0, i_8_182_2274_0;
  output o_8_182_0_0;
  assign o_8_182_0_0 = ~((~i_8_182_0_0 & ((~i_8_182_1_0 & ~i_8_182_3_0 & ~i_8_182_81_0 & ~i_8_182_82_0 & ~i_8_182_1386_0 & ~i_8_182_2134_0) | (~i_8_182_112_0 & ~i_8_182_673_0 & ~i_8_182_829_0 & ~i_8_182_1270_0 & ~i_8_182_2116_0 & ~i_8_182_2142_0))) | (~i_8_182_73_0 & ((~i_8_182_82_0 & ~i_8_182_434_0 & i_8_182_705_0 & ~i_8_182_2116_0) | (~i_8_182_198_0 & ~i_8_182_1198_0 & ~i_8_182_1992_0 & ~i_8_182_2025_0 & ~i_8_182_2142_0))) | (~i_8_182_111_0 & ((~i_8_182_279_0 & ~i_8_182_318_0 & ~i_8_182_832_0 & ~i_8_182_1033_0 & ~i_8_182_1182_0 & ~i_8_182_1299_0 & ~i_8_182_1587_0 & ~i_8_182_1923_0 & ~i_8_182_2035_0) | (~i_8_182_243_0 & ~i_8_182_892_0 & ~i_8_182_1081_0 & i_8_182_1813_0 & ~i_8_182_2274_0))) | (~i_8_182_198_0 & ((~i_8_182_1_0 & ~i_8_182_673_0 & i_8_182_1749_0 & ~i_8_182_1845_0) | (~i_8_182_666_0 & i_8_182_705_0 & ~i_8_182_1172_0 & ~i_8_182_1386_0 & i_8_182_1801_0 & ~i_8_182_1923_0 & ~i_8_182_2157_0))) | (~i_8_182_1846_0 & ((~i_8_182_1_0 & ~i_8_182_729_0 & ((~i_8_182_153_0 & ~i_8_182_279_0 & ~i_8_182_604_0 & ~i_8_182_1028_0 & ~i_8_182_1587_0 & ~i_8_182_1791_0) | (~i_8_182_283_0 & ~i_8_182_630_0 & ~i_8_182_1633_0 & ~i_8_182_1845_0 & ~i_8_182_2157_0 & ~i_8_182_2274_0))) | (~i_8_182_829_0 & ~i_8_182_892_0 & ~i_8_182_1028_0 & ~i_8_182_1386_0 & ~i_8_182_1813_0 & ~i_8_182_1845_0 & ~i_8_182_2116_0))) | (~i_8_182_243_0 & ((~i_8_182_434_0 & ~i_8_182_486_0 & ~i_8_182_666_0 & ~i_8_182_1182_0 & ~i_8_182_1351_0 & ~i_8_182_2142_0) | (i_8_182_82_0 & ~i_8_182_279_0 & ~i_8_182_829_0 & ~i_8_182_2025_0 & ~i_8_182_2133_0 & ~i_8_182_2274_0))) | (~i_8_182_1386_0 & ((~i_8_182_434_0 & i_8_182_832_0 & ~i_8_182_865_0 & ~i_8_182_1677_0 & ~i_8_182_1845_0 & ~i_8_182_2025_0 & ~i_8_182_2128_0) | (~i_8_182_227_0 & ~i_8_182_1081_0 & ~i_8_182_1587_0 & ~i_8_182_1801_0 & ~i_8_182_2115_0 & ~i_8_182_2116_0 & ~i_8_182_2157_0))) | (~i_8_182_1845_0 & ((~i_8_182_436_0 & i_8_182_1677_0 & ~i_8_182_1881_0) | (~i_8_182_81_0 & i_8_182_604_0 & ~i_8_182_2116_0))) | (~i_8_182_283_0 & i_8_182_450_0 & ~i_8_182_673_0 & ~i_8_182_1270_0 & ~i_8_182_1351_0 & i_8_182_1434_0 & ~i_8_182_1912_0 & ~i_8_182_1992_0));
endmodule



// Benchmark "kernel_8_183" written by ABC on Sun Jul 19 10:06:14 2020

module kernel_8_183 ( 
    i_8_183_1_0, i_8_183_95_0, i_8_183_103_0, i_8_183_104_0, i_8_183_106_0,
    i_8_183_143_0, i_8_183_214_0, i_8_183_219_0, i_8_183_220_0,
    i_8_183_243_0, i_8_183_244_0, i_8_183_265_0, i_8_183_310_0,
    i_8_183_346_0, i_8_183_377_0, i_8_183_395_0, i_8_183_419_0,
    i_8_183_422_0, i_8_183_427_0, i_8_183_438_0, i_8_183_440_0,
    i_8_183_446_0, i_8_183_460_0, i_8_183_474_0, i_8_183_484_0,
    i_8_183_505_0, i_8_183_522_0, i_8_183_584_0, i_8_183_599_0,
    i_8_183_627_0, i_8_183_689_0, i_8_183_691_0, i_8_183_706_0,
    i_8_183_707_0, i_8_183_718_0, i_8_183_780_0, i_8_183_872_0,
    i_8_183_926_0, i_8_183_931_0, i_8_183_932_0, i_8_183_978_0,
    i_8_183_1021_0, i_8_183_1030_0, i_8_183_1070_0, i_8_183_1074_0,
    i_8_183_1107_0, i_8_183_1108_0, i_8_183_1137_0, i_8_183_1159_0,
    i_8_183_1233_0, i_8_183_1265_0, i_8_183_1267_0, i_8_183_1364_0,
    i_8_183_1376_0, i_8_183_1382_0, i_8_183_1414_0, i_8_183_1434_0,
    i_8_183_1453_0, i_8_183_1531_0, i_8_183_1532_0, i_8_183_1533_0,
    i_8_183_1539_0, i_8_183_1548_0, i_8_183_1555_0, i_8_183_1592_0,
    i_8_183_1633_0, i_8_183_1642_0, i_8_183_1648_0, i_8_183_1677_0,
    i_8_183_1703_0, i_8_183_1706_0, i_8_183_1723_0, i_8_183_1758_0,
    i_8_183_1761_0, i_8_183_1819_0, i_8_183_1857_0, i_8_183_1889_0,
    i_8_183_1918_0, i_8_183_1963_0, i_8_183_2003_0, i_8_183_2010_0,
    i_8_183_2011_0, i_8_183_2028_0, i_8_183_2049_0, i_8_183_2057_0,
    i_8_183_2093_0, i_8_183_2114_0, i_8_183_2153_0, i_8_183_2154_0,
    i_8_183_2156_0, i_8_183_2165_0, i_8_183_2182_0, i_8_183_2183_0,
    i_8_183_2190_0, i_8_183_2214_0, i_8_183_2240_0, i_8_183_2270_0,
    i_8_183_2273_0, i_8_183_2294_0, i_8_183_2300_0,
    o_8_183_0_0  );
  input  i_8_183_1_0, i_8_183_95_0, i_8_183_103_0, i_8_183_104_0,
    i_8_183_106_0, i_8_183_143_0, i_8_183_214_0, i_8_183_219_0,
    i_8_183_220_0, i_8_183_243_0, i_8_183_244_0, i_8_183_265_0,
    i_8_183_310_0, i_8_183_346_0, i_8_183_377_0, i_8_183_395_0,
    i_8_183_419_0, i_8_183_422_0, i_8_183_427_0, i_8_183_438_0,
    i_8_183_440_0, i_8_183_446_0, i_8_183_460_0, i_8_183_474_0,
    i_8_183_484_0, i_8_183_505_0, i_8_183_522_0, i_8_183_584_0,
    i_8_183_599_0, i_8_183_627_0, i_8_183_689_0, i_8_183_691_0,
    i_8_183_706_0, i_8_183_707_0, i_8_183_718_0, i_8_183_780_0,
    i_8_183_872_0, i_8_183_926_0, i_8_183_931_0, i_8_183_932_0,
    i_8_183_978_0, i_8_183_1021_0, i_8_183_1030_0, i_8_183_1070_0,
    i_8_183_1074_0, i_8_183_1107_0, i_8_183_1108_0, i_8_183_1137_0,
    i_8_183_1159_0, i_8_183_1233_0, i_8_183_1265_0, i_8_183_1267_0,
    i_8_183_1364_0, i_8_183_1376_0, i_8_183_1382_0, i_8_183_1414_0,
    i_8_183_1434_0, i_8_183_1453_0, i_8_183_1531_0, i_8_183_1532_0,
    i_8_183_1533_0, i_8_183_1539_0, i_8_183_1548_0, i_8_183_1555_0,
    i_8_183_1592_0, i_8_183_1633_0, i_8_183_1642_0, i_8_183_1648_0,
    i_8_183_1677_0, i_8_183_1703_0, i_8_183_1706_0, i_8_183_1723_0,
    i_8_183_1758_0, i_8_183_1761_0, i_8_183_1819_0, i_8_183_1857_0,
    i_8_183_1889_0, i_8_183_1918_0, i_8_183_1963_0, i_8_183_2003_0,
    i_8_183_2010_0, i_8_183_2011_0, i_8_183_2028_0, i_8_183_2049_0,
    i_8_183_2057_0, i_8_183_2093_0, i_8_183_2114_0, i_8_183_2153_0,
    i_8_183_2154_0, i_8_183_2156_0, i_8_183_2165_0, i_8_183_2182_0,
    i_8_183_2183_0, i_8_183_2190_0, i_8_183_2214_0, i_8_183_2240_0,
    i_8_183_2270_0, i_8_183_2273_0, i_8_183_2294_0, i_8_183_2300_0;
  output o_8_183_0_0;
  assign o_8_183_0_0 = 0;
endmodule



// Benchmark "kernel_8_184" written by ABC on Sun Jul 19 10:06:15 2020

module kernel_8_184 ( 
    i_8_184_33_0, i_8_184_102_0, i_8_184_105_0, i_8_184_107_0,
    i_8_184_154_0, i_8_184_158_0, i_8_184_247_0, i_8_184_302_0,
    i_8_184_348_0, i_8_184_349_0, i_8_184_363_0, i_8_184_364_0,
    i_8_184_428_0, i_8_184_621_0, i_8_184_622_0, i_8_184_623_0,
    i_8_184_624_0, i_8_184_632_0, i_8_184_660_0, i_8_184_662_0,
    i_8_184_687_0, i_8_184_688_0, i_8_184_692_0, i_8_184_699_0,
    i_8_184_723_0, i_8_184_780_0, i_8_184_781_0, i_8_184_782_0,
    i_8_184_822_0, i_8_184_824_0, i_8_184_825_0, i_8_184_840_0,
    i_8_184_867_0, i_8_184_869_0, i_8_184_870_0, i_8_184_871_0,
    i_8_184_872_0, i_8_184_886_0, i_8_184_967_0, i_8_184_1008_0,
    i_8_184_1011_0, i_8_184_1026_0, i_8_184_1054_0, i_8_184_1056_0,
    i_8_184_1058_0, i_8_184_1060_0, i_8_184_1108_0, i_8_184_1192_0,
    i_8_184_1272_0, i_8_184_1274_0, i_8_184_1305_0, i_8_184_1306_0,
    i_8_184_1307_0, i_8_184_1341_0, i_8_184_1342_0, i_8_184_1407_0,
    i_8_184_1408_0, i_8_184_1409_0, i_8_184_1411_0, i_8_184_1431_0,
    i_8_184_1434_0, i_8_184_1437_0, i_8_184_1439_0, i_8_184_1449_0,
    i_8_184_1474_0, i_8_184_1625_0, i_8_184_1641_0, i_8_184_1642_0,
    i_8_184_1644_0, i_8_184_1648_0, i_8_184_1650_0, i_8_184_1652_0,
    i_8_184_1654_0, i_8_184_1676_0, i_8_184_1679_0, i_8_184_1681_0,
    i_8_184_1713_0, i_8_184_1716_0, i_8_184_1717_0, i_8_184_1720_0,
    i_8_184_1722_0, i_8_184_1723_0, i_8_184_1741_0, i_8_184_1750_0,
    i_8_184_1751_0, i_8_184_1758_0, i_8_184_1812_0, i_8_184_1828_0,
    i_8_184_1881_0, i_8_184_1882_0, i_8_184_1884_0, i_8_184_2088_0,
    i_8_184_2133_0, i_8_184_2136_0, i_8_184_2138_0, i_8_184_2143_0,
    i_8_184_2242_0, i_8_184_2249_0, i_8_184_2272_0, i_8_184_2288_0,
    o_8_184_0_0  );
  input  i_8_184_33_0, i_8_184_102_0, i_8_184_105_0, i_8_184_107_0,
    i_8_184_154_0, i_8_184_158_0, i_8_184_247_0, i_8_184_302_0,
    i_8_184_348_0, i_8_184_349_0, i_8_184_363_0, i_8_184_364_0,
    i_8_184_428_0, i_8_184_621_0, i_8_184_622_0, i_8_184_623_0,
    i_8_184_624_0, i_8_184_632_0, i_8_184_660_0, i_8_184_662_0,
    i_8_184_687_0, i_8_184_688_0, i_8_184_692_0, i_8_184_699_0,
    i_8_184_723_0, i_8_184_780_0, i_8_184_781_0, i_8_184_782_0,
    i_8_184_822_0, i_8_184_824_0, i_8_184_825_0, i_8_184_840_0,
    i_8_184_867_0, i_8_184_869_0, i_8_184_870_0, i_8_184_871_0,
    i_8_184_872_0, i_8_184_886_0, i_8_184_967_0, i_8_184_1008_0,
    i_8_184_1011_0, i_8_184_1026_0, i_8_184_1054_0, i_8_184_1056_0,
    i_8_184_1058_0, i_8_184_1060_0, i_8_184_1108_0, i_8_184_1192_0,
    i_8_184_1272_0, i_8_184_1274_0, i_8_184_1305_0, i_8_184_1306_0,
    i_8_184_1307_0, i_8_184_1341_0, i_8_184_1342_0, i_8_184_1407_0,
    i_8_184_1408_0, i_8_184_1409_0, i_8_184_1411_0, i_8_184_1431_0,
    i_8_184_1434_0, i_8_184_1437_0, i_8_184_1439_0, i_8_184_1449_0,
    i_8_184_1474_0, i_8_184_1625_0, i_8_184_1641_0, i_8_184_1642_0,
    i_8_184_1644_0, i_8_184_1648_0, i_8_184_1650_0, i_8_184_1652_0,
    i_8_184_1654_0, i_8_184_1676_0, i_8_184_1679_0, i_8_184_1681_0,
    i_8_184_1713_0, i_8_184_1716_0, i_8_184_1717_0, i_8_184_1720_0,
    i_8_184_1722_0, i_8_184_1723_0, i_8_184_1741_0, i_8_184_1750_0,
    i_8_184_1751_0, i_8_184_1758_0, i_8_184_1812_0, i_8_184_1828_0,
    i_8_184_1881_0, i_8_184_1882_0, i_8_184_1884_0, i_8_184_2088_0,
    i_8_184_2133_0, i_8_184_2136_0, i_8_184_2138_0, i_8_184_2143_0,
    i_8_184_2242_0, i_8_184_2249_0, i_8_184_2272_0, i_8_184_2288_0;
  output o_8_184_0_0;
  assign o_8_184_0_0 = ~((~i_8_184_624_0 & ((~i_8_184_107_0 & ((~i_8_184_870_0 & ((~i_8_184_824_0 & ~i_8_184_872_0 & ((~i_8_184_102_0 & ~i_8_184_1008_0 & ~i_8_184_1342_0 & ~i_8_184_1812_0 & ((~i_8_184_33_0 & ~i_8_184_247_0 & ~i_8_184_349_0 & ~i_8_184_428_0 & ~i_8_184_692_0 & ~i_8_184_781_0 & ~i_8_184_782_0 & ~i_8_184_822_0 & ~i_8_184_867_0 & ~i_8_184_1011_0 & ~i_8_184_1108_0 & ~i_8_184_1676_0 & ~i_8_184_1679_0 & ~i_8_184_1716_0 & ~i_8_184_2136_0) | (~i_8_184_105_0 & ~i_8_184_621_0 & ~i_8_184_622_0 & ~i_8_184_780_0 & ~i_8_184_1274_0 & ~i_8_184_1341_0 & i_8_184_1434_0 & ~i_8_184_2143_0 & ~i_8_184_2242_0 & ~i_8_184_2288_0))) | (~i_8_184_621_0 & ~i_8_184_623_0 & ~i_8_184_632_0 & ~i_8_184_699_0 & ~i_8_184_780_0 & ~i_8_184_782_0 & ~i_8_184_871_0 & ~i_8_184_1341_0 & ~i_8_184_1434_0 & ~i_8_184_1449_0 & ~i_8_184_1679_0 & ~i_8_184_1716_0 & ~i_8_184_2138_0 & ~i_8_184_2249_0 & ~i_8_184_2288_0))) | (~i_8_184_302_0 & ~i_8_184_621_0 & ~i_8_184_662_0 & i_8_184_687_0 & ~i_8_184_825_0 & ~i_8_184_871_0 & ~i_8_184_1341_0 & ~i_8_184_2136_0))) | (~i_8_184_302_0 & ~i_8_184_621_0 & ~i_8_184_781_0 & ~i_8_184_840_0 & ~i_8_184_869_0 & ~i_8_184_872_0 & ~i_8_184_1026_0 & ~i_8_184_1056_0 & ~i_8_184_1342_0 & ~i_8_184_1437_0 & ~i_8_184_1449_0 & ~i_8_184_1474_0 & ~i_8_184_1652_0 & ~i_8_184_1713_0 & ~i_8_184_1716_0 & ~i_8_184_1751_0 & ~i_8_184_2138_0 & ~i_8_184_2143_0 & ~i_8_184_2249_0))) | (~i_8_184_348_0 & ~i_8_184_780_0 & ((~i_8_184_621_0 & ~i_8_184_660_0 & ~i_8_184_822_0 & ~i_8_184_867_0 & ~i_8_184_1008_0 & ~i_8_184_1026_0 & ~i_8_184_1409_0 & ~i_8_184_1449_0 & ~i_8_184_1644_0 & i_8_184_2133_0 & ~i_8_184_2138_0) | (~i_8_184_428_0 & ~i_8_184_622_0 & i_8_184_688_0 & ~i_8_184_781_0 & ~i_8_184_870_0 & ~i_8_184_872_0 & ~i_8_184_1108_0 & ~i_8_184_2288_0))) | (~i_8_184_660_0 & ~i_8_184_825_0 & ~i_8_184_871_0 & i_8_184_1054_0 & ~i_8_184_1108_0 & ~i_8_184_1439_0 & ~i_8_184_2133_0 & ~i_8_184_2242_0 & ~i_8_184_2249_0))) | (~i_8_184_2288_0 & ((~i_8_184_871_0 & ((~i_8_184_33_0 & ((~i_8_184_107_0 & ~i_8_184_867_0 & ~i_8_184_870_0 & i_8_184_1056_0 & ~i_8_184_1676_0 & ~i_8_184_1713_0 & ~i_8_184_1812_0 & ~i_8_184_2133_0) | (~i_8_184_105_0 & ~i_8_184_154_0 & ~i_8_184_302_0 & ~i_8_184_781_0 & ~i_8_184_824_0 & ~i_8_184_872_0 & ~i_8_184_1342_0 & i_8_184_1648_0 & ~i_8_184_1828_0 & ~i_8_184_2136_0))) | (~i_8_184_872_0 & ((~i_8_184_302_0 & ~i_8_184_621_0 & ~i_8_184_780_0 & ~i_8_184_782_0 & i_8_184_1407_0 & ~i_8_184_1434_0) | (~i_8_184_363_0 & ~i_8_184_824_0 & ~i_8_184_825_0 & ~i_8_184_869_0 & ~i_8_184_1026_0 & i_8_184_1306_0 & ~i_8_184_1342_0 & ~i_8_184_2272_0))))) | (~i_8_184_781_0 & ((~i_8_184_102_0 & ~i_8_184_1341_0 & ~i_8_184_1758_0 & ((~i_8_184_158_0 & ~i_8_184_622_0 & ~i_8_184_623_0 & ~i_8_184_688_0 & ~i_8_184_825_0 & ~i_8_184_872_0 & ~i_8_184_1054_0 & ~i_8_184_1307_0 & ~i_8_184_1716_0 & ~i_8_184_1717_0 & i_8_184_1750_0 & ~i_8_184_2133_0 & ~i_8_184_2143_0) | (~i_8_184_247_0 & ~i_8_184_302_0 & ~i_8_184_662_0 & ~i_8_184_782_0 & ~i_8_184_824_0 & i_8_184_1439_0 & ~i_8_184_2249_0))) | (~i_8_184_158_0 & ~i_8_184_662_0 & i_8_184_1274_0 & ~i_8_184_1751_0 & ~i_8_184_2136_0))) | (~i_8_184_107_0 & ((~i_8_184_302_0 & ~i_8_184_660_0 & ~i_8_184_886_0 & ~i_8_184_1449_0 & i_8_184_1652_0 & ~i_8_184_1681_0 & ~i_8_184_1741_0) | (~i_8_184_154_0 & ~i_8_184_247_0 & ~i_8_184_349_0 & ~i_8_184_428_0 & ~i_8_184_782_0 & ~i_8_184_870_0 & i_8_184_967_0 & ~i_8_184_1026_0 & ~i_8_184_1272_0 & ~i_8_184_1342_0 & ~i_8_184_1439_0 & ~i_8_184_1716_0 & ~i_8_184_1717_0 & ~i_8_184_1750_0 & ~i_8_184_1751_0 & ~i_8_184_1828_0 & ~i_8_184_1881_0 & ~i_8_184_1882_0 & ~i_8_184_2138_0))) | (~i_8_184_825_0 & ~i_8_184_1437_0 & ((~i_8_184_105_0 & ~i_8_184_302_0 & i_8_184_692_0 & ~i_8_184_869_0 & ~i_8_184_1342_0 & ~i_8_184_1648_0 & ~i_8_184_1758_0) | (~i_8_184_349_0 & ~i_8_184_870_0 & ~i_8_184_1026_0 & i_8_184_1641_0 & ~i_8_184_1716_0 & ~i_8_184_1717_0 & ~i_8_184_1828_0))))) | (~i_8_184_1108_0 & ((~i_8_184_33_0 & ((~i_8_184_107_0 & i_8_184_348_0 & ~i_8_184_632_0 & ~i_8_184_780_0 & ~i_8_184_825_0 & ~i_8_184_1342_0) | (~i_8_184_782_0 & ~i_8_184_870_0 & ~i_8_184_872_0 & i_8_184_1058_0 & ~i_8_184_1758_0 & ~i_8_184_1812_0 & ~i_8_184_2136_0))) | (~i_8_184_107_0 & ~i_8_184_692_0 & ((~i_8_184_662_0 & ~i_8_184_869_0 & i_8_184_1411_0 & ~i_8_184_1437_0 & i_8_184_1654_0 & ~i_8_184_1713_0) | (i_8_184_428_0 & ~i_8_184_622_0 & ~i_8_184_781_0 & ~i_8_184_1679_0 & ~i_8_184_1750_0 & ~i_8_184_1751_0 & ~i_8_184_1758_0 & ~i_8_184_2249_0))) | (~i_8_184_1431_0 & ((~i_8_184_302_0 & ~i_8_184_363_0 & ~i_8_184_622_0 & ~i_8_184_782_0 & ~i_8_184_824_0 & ~i_8_184_1751_0 & i_8_184_2143_0) | (~i_8_184_158_0 & ~i_8_184_247_0 & ~i_8_184_662_0 & ~i_8_184_699_0 & ~i_8_184_780_0 & ~i_8_184_822_0 & ~i_8_184_872_0 & ~i_8_184_2136_0 & i_8_184_2242_0))))) | (~i_8_184_1008_0 & ((~i_8_184_1717_0 & ((~i_8_184_102_0 & ~i_8_184_1713_0 & ~i_8_184_2242_0 & ((~i_8_184_105_0 & ~i_8_184_662_0 & ~i_8_184_692_0 & ~i_8_184_824_0 & ~i_8_184_870_0 & i_8_184_1411_0 & ~i_8_184_1449_0 & ~i_8_184_1644_0 & ~i_8_184_1716_0 & ~i_8_184_1751_0 & ~i_8_184_1812_0) | (~i_8_184_621_0 & ~i_8_184_687_0 & ~i_8_184_871_0 & ~i_8_184_1274_0 & i_8_184_1644_0 & ~i_8_184_2138_0))) | (~i_8_184_621_0 & ~i_8_184_781_0 & ~i_8_184_825_0 & ~i_8_184_869_0 & ~i_8_184_872_0 & i_8_184_967_0 & ~i_8_184_1341_0 & ~i_8_184_1439_0 & ~i_8_184_1449_0 & ~i_8_184_1625_0 & ~i_8_184_1679_0))) | (~i_8_184_105_0 & ~i_8_184_158_0 & ~i_8_184_363_0 & ~i_8_184_623_0 & ~i_8_184_688_0 & ~i_8_184_840_0 & ~i_8_184_886_0 & ~i_8_184_967_0 & i_8_184_1108_0 & ~i_8_184_1274_0 & ~i_8_184_1341_0 & ~i_8_184_1652_0 & ~i_8_184_1751_0))) | (~i_8_184_428_0 & ((i_8_184_302_0 & ~i_8_184_662_0 & ~i_8_184_781_0 & i_8_184_1409_0 & ~i_8_184_1434_0 & ~i_8_184_1751_0) | (~i_8_184_967_0 & i_8_184_1054_0 & i_8_184_1272_0 & ~i_8_184_1681_0 & ~i_8_184_1828_0))) | (~i_8_184_621_0 & ((~i_8_184_302_0 & ~i_8_184_660_0 & ~i_8_184_871_0 & ~i_8_184_1011_0 & ~i_8_184_1306_0 & i_8_184_1431_0 & ~i_8_184_1449_0 & i_8_184_1648_0 & ~i_8_184_1812_0 & ~i_8_184_2088_0) | (~i_8_184_158_0 & ~i_8_184_623_0 & ~i_8_184_782_0 & ~i_8_184_869_0 & ~i_8_184_870_0 & ~i_8_184_1431_0 & ~i_8_184_1750_0 & ~i_8_184_2138_0 & i_8_184_2143_0))) | (~i_8_184_302_0 & ((~i_8_184_107_0 & ~i_8_184_154_0 & ~i_8_184_623_0 & ~i_8_184_782_0 & ~i_8_184_824_0 & ~i_8_184_840_0 & ~i_8_184_872_0 & ~i_8_184_1192_0 & ~i_8_184_1676_0 & ~i_8_184_1679_0 & ~i_8_184_1341_0 & ~i_8_184_1437_0 & ~i_8_184_1716_0 & ~i_8_184_1812_0 & ~i_8_184_2136_0 & ~i_8_184_2138_0) | (i_8_184_632_0 & i_8_184_1679_0 & i_8_184_2138_0 & i_8_184_2143_0))) | (~i_8_184_871_0 & ((~i_8_184_107_0 & ~i_8_184_872_0 & ((~i_8_184_824_0 & ~i_8_184_870_0 & ~i_8_184_154_0 & ~i_8_184_687_0 & i_8_184_1058_0 & ~i_8_184_1411_0 & ~i_8_184_1474_0 & ~i_8_184_1641_0 & ~i_8_184_2138_0) | (~i_8_184_781_0 & ~i_8_184_822_0 & ~i_8_184_825_0 & ~i_8_184_867_0 & ~i_8_184_1341_0 & i_8_184_1408_0 & ~i_8_184_2136_0 & ~i_8_184_2249_0))) | (~i_8_184_782_0 & ((~i_8_184_158_0 & i_8_184_349_0 & ~i_8_184_780_0 & ~i_8_184_1272_0 & ~i_8_184_1341_0 & ~i_8_184_1449_0 & ~i_8_184_1648_0 & ~i_8_184_1713_0 & ~i_8_184_1812_0) | (~i_8_184_824_0 & ~i_8_184_840_0 & ~i_8_184_632_0 & ~i_8_184_781_0 & i_8_184_1652_0 & ~i_8_184_1676_0 & ~i_8_184_1758_0 & ~i_8_184_2242_0))))) | (~i_8_184_158_0 & ~i_8_184_1341_0 & ((~i_8_184_154_0 & ~i_8_184_247_0 & i_8_184_624_0 & ~i_8_184_660_0 & ~i_8_184_822_0 & ~i_8_184_1272_0 & ~i_8_184_1713_0 & ~i_8_184_1751_0 & ~i_8_184_1812_0 & ~i_8_184_2133_0 & i_8_184_2136_0) | (i_8_184_1056_0 & i_8_184_1407_0 & i_8_184_1884_0 & ~i_8_184_2138_0))) | (i_8_184_1408_0 & ((~i_8_184_363_0 & ~i_8_184_688_0 & ~i_8_184_782_0 & ~i_8_184_825_0 & i_8_184_1108_0 & ~i_8_184_1449_0 & ~i_8_184_1722_0) | (~i_8_184_1011_0 & ~i_8_184_1026_0 & ~i_8_184_1411_0 & ~i_8_184_1434_0 & i_8_184_1882_0 & i_8_184_2136_0))) | (~i_8_184_2136_0 & ((i_8_184_428_0 & ~i_8_184_1307_0 & ~i_8_184_1431_0 & ~i_8_184_1439_0 & i_8_184_1648_0 & ~i_8_184_1828_0 & ~i_8_184_2249_0) | (~i_8_184_781_0 & ~i_8_184_869_0 & i_8_184_967_0 & ~i_8_184_1408_0 & ~i_8_184_1625_0 & ~i_8_184_1676_0 & ~i_8_184_1750_0 & i_8_184_2138_0 & ~i_8_184_2272_0))) | (~i_8_184_1751_0 & i_8_184_1884_0 & ~i_8_184_2143_0 & i_8_184_2249_0 & ~i_8_184_2272_0));
endmodule



// Benchmark "kernel_8_185" written by ABC on Sun Jul 19 10:06:16 2020

module kernel_8_185 ( 
    i_8_185_19_0, i_8_185_43_0, i_8_185_44_0, i_8_185_99_0, i_8_185_136_0,
    i_8_185_138_0, i_8_185_187_0, i_8_185_225_0, i_8_185_262_0,
    i_8_185_334_0, i_8_185_336_0, i_8_185_365_0, i_8_185_369_0,
    i_8_185_370_0, i_8_185_379_0, i_8_185_423_0, i_8_185_427_0,
    i_8_185_439_0, i_8_185_492_0, i_8_185_497_0, i_8_185_505_0,
    i_8_185_554_0, i_8_185_568_0, i_8_185_588_0, i_8_185_594_0,
    i_8_185_597_0, i_8_185_604_0, i_8_185_630_0, i_8_185_639_0,
    i_8_185_652_0, i_8_185_661_0, i_8_185_675_0, i_8_185_678_0,
    i_8_185_695_0, i_8_185_705_0, i_8_185_833_0, i_8_185_837_0,
    i_8_185_846_0, i_8_185_850_0, i_8_185_855_0, i_8_185_882_0,
    i_8_185_883_0, i_8_185_937_0, i_8_185_966_0, i_8_185_1062_0,
    i_8_185_1071_0, i_8_185_1107_0, i_8_185_1110_0, i_8_185_1117_0,
    i_8_185_1135_0, i_8_185_1153_0, i_8_185_1191_0, i_8_185_1215_0,
    i_8_185_1226_0, i_8_185_1243_0, i_8_185_1269_0, i_8_185_1297_0,
    i_8_185_1351_0, i_8_185_1354_0, i_8_185_1355_0, i_8_185_1431_0,
    i_8_185_1434_0, i_8_185_1474_0, i_8_185_1486_0, i_8_185_1503_0,
    i_8_185_1602_0, i_8_185_1611_0, i_8_185_1629_0, i_8_185_1671_0,
    i_8_185_1681_0, i_8_185_1682_0, i_8_185_1696_0, i_8_185_1710_0,
    i_8_185_1711_0, i_8_185_1746_0, i_8_185_1755_0, i_8_185_1756_0,
    i_8_185_1767_0, i_8_185_1809_0, i_8_185_1812_0, i_8_185_1824_0,
    i_8_185_1836_0, i_8_185_1840_0, i_8_185_1867_0, i_8_185_1881_0,
    i_8_185_1882_0, i_8_185_1891_0, i_8_185_1945_0, i_8_185_1962_0,
    i_8_185_1963_0, i_8_185_1980_0, i_8_185_2038_0, i_8_185_2106_0,
    i_8_185_2107_0, i_8_185_2125_0, i_8_185_2149_0, i_8_185_2152_0,
    i_8_185_2156_0, i_8_185_2169_0, i_8_185_2242_0,
    o_8_185_0_0  );
  input  i_8_185_19_0, i_8_185_43_0, i_8_185_44_0, i_8_185_99_0,
    i_8_185_136_0, i_8_185_138_0, i_8_185_187_0, i_8_185_225_0,
    i_8_185_262_0, i_8_185_334_0, i_8_185_336_0, i_8_185_365_0,
    i_8_185_369_0, i_8_185_370_0, i_8_185_379_0, i_8_185_423_0,
    i_8_185_427_0, i_8_185_439_0, i_8_185_492_0, i_8_185_497_0,
    i_8_185_505_0, i_8_185_554_0, i_8_185_568_0, i_8_185_588_0,
    i_8_185_594_0, i_8_185_597_0, i_8_185_604_0, i_8_185_630_0,
    i_8_185_639_0, i_8_185_652_0, i_8_185_661_0, i_8_185_675_0,
    i_8_185_678_0, i_8_185_695_0, i_8_185_705_0, i_8_185_833_0,
    i_8_185_837_0, i_8_185_846_0, i_8_185_850_0, i_8_185_855_0,
    i_8_185_882_0, i_8_185_883_0, i_8_185_937_0, i_8_185_966_0,
    i_8_185_1062_0, i_8_185_1071_0, i_8_185_1107_0, i_8_185_1110_0,
    i_8_185_1117_0, i_8_185_1135_0, i_8_185_1153_0, i_8_185_1191_0,
    i_8_185_1215_0, i_8_185_1226_0, i_8_185_1243_0, i_8_185_1269_0,
    i_8_185_1297_0, i_8_185_1351_0, i_8_185_1354_0, i_8_185_1355_0,
    i_8_185_1431_0, i_8_185_1434_0, i_8_185_1474_0, i_8_185_1486_0,
    i_8_185_1503_0, i_8_185_1602_0, i_8_185_1611_0, i_8_185_1629_0,
    i_8_185_1671_0, i_8_185_1681_0, i_8_185_1682_0, i_8_185_1696_0,
    i_8_185_1710_0, i_8_185_1711_0, i_8_185_1746_0, i_8_185_1755_0,
    i_8_185_1756_0, i_8_185_1767_0, i_8_185_1809_0, i_8_185_1812_0,
    i_8_185_1824_0, i_8_185_1836_0, i_8_185_1840_0, i_8_185_1867_0,
    i_8_185_1881_0, i_8_185_1882_0, i_8_185_1891_0, i_8_185_1945_0,
    i_8_185_1962_0, i_8_185_1963_0, i_8_185_1980_0, i_8_185_2038_0,
    i_8_185_2106_0, i_8_185_2107_0, i_8_185_2125_0, i_8_185_2149_0,
    i_8_185_2152_0, i_8_185_2156_0, i_8_185_2169_0, i_8_185_2242_0;
  output o_8_185_0_0;
  assign o_8_185_0_0 = 0;
endmodule



// Benchmark "kernel_8_186" written by ABC on Sun Jul 19 10:06:17 2020

module kernel_8_186 ( 
    i_8_186_22_0, i_8_186_34_0, i_8_186_98_0, i_8_186_107_0, i_8_186_114_0,
    i_8_186_130_0, i_8_186_131_0, i_8_186_165_0, i_8_186_166_0,
    i_8_186_256_0, i_8_186_320_0, i_8_186_322_0, i_8_186_345_0,
    i_8_186_375_0, i_8_186_390_0, i_8_186_397_0, i_8_186_398_0,
    i_8_186_439_0, i_8_186_450_0, i_8_186_451_0, i_8_186_457_0,
    i_8_186_492_0, i_8_186_508_0, i_8_186_530_0, i_8_186_580_0,
    i_8_186_606_0, i_8_186_608_0, i_8_186_626_0, i_8_186_639_0,
    i_8_186_643_0, i_8_186_660_0, i_8_186_665_0, i_8_186_675_0,
    i_8_186_707_0, i_8_186_748_0, i_8_186_750_0, i_8_186_778_0,
    i_8_186_811_0, i_8_186_838_0, i_8_186_853_0, i_8_186_883_0,
    i_8_186_888_0, i_8_186_921_0, i_8_186_955_0, i_8_186_1099_0,
    i_8_186_1102_0, i_8_186_1108_0, i_8_186_1134_0, i_8_186_1135_0,
    i_8_186_1231_0, i_8_186_1233_0, i_8_186_1236_0, i_8_186_1263_0,
    i_8_186_1273_0, i_8_186_1286_0, i_8_186_1300_0, i_8_186_1352_0,
    i_8_186_1360_0, i_8_186_1362_0, i_8_186_1384_0, i_8_186_1423_0,
    i_8_186_1441_0, i_8_186_1442_0, i_8_186_1461_0, i_8_186_1462_0,
    i_8_186_1471_0, i_8_186_1512_0, i_8_186_1559_0, i_8_186_1569_0,
    i_8_186_1570_0, i_8_186_1603_0, i_8_186_1615_0, i_8_186_1616_0,
    i_8_186_1618_0, i_8_186_1642_0, i_8_186_1643_0, i_8_186_1644_0,
    i_8_186_1719_0, i_8_186_1781_0, i_8_186_1783_0, i_8_186_1787_0,
    i_8_186_1822_0, i_8_186_1836_0, i_8_186_1849_0, i_8_186_1852_0,
    i_8_186_1935_0, i_8_186_1954_0, i_8_186_1958_0, i_8_186_1981_0,
    i_8_186_1993_0, i_8_186_2055_0, i_8_186_2077_0, i_8_186_2088_0,
    i_8_186_2120_0, i_8_186_2151_0, i_8_186_2163_0, i_8_186_2169_0,
    i_8_186_2170_0, i_8_186_2212_0, i_8_186_2296_0,
    o_8_186_0_0  );
  input  i_8_186_22_0, i_8_186_34_0, i_8_186_98_0, i_8_186_107_0,
    i_8_186_114_0, i_8_186_130_0, i_8_186_131_0, i_8_186_165_0,
    i_8_186_166_0, i_8_186_256_0, i_8_186_320_0, i_8_186_322_0,
    i_8_186_345_0, i_8_186_375_0, i_8_186_390_0, i_8_186_397_0,
    i_8_186_398_0, i_8_186_439_0, i_8_186_450_0, i_8_186_451_0,
    i_8_186_457_0, i_8_186_492_0, i_8_186_508_0, i_8_186_530_0,
    i_8_186_580_0, i_8_186_606_0, i_8_186_608_0, i_8_186_626_0,
    i_8_186_639_0, i_8_186_643_0, i_8_186_660_0, i_8_186_665_0,
    i_8_186_675_0, i_8_186_707_0, i_8_186_748_0, i_8_186_750_0,
    i_8_186_778_0, i_8_186_811_0, i_8_186_838_0, i_8_186_853_0,
    i_8_186_883_0, i_8_186_888_0, i_8_186_921_0, i_8_186_955_0,
    i_8_186_1099_0, i_8_186_1102_0, i_8_186_1108_0, i_8_186_1134_0,
    i_8_186_1135_0, i_8_186_1231_0, i_8_186_1233_0, i_8_186_1236_0,
    i_8_186_1263_0, i_8_186_1273_0, i_8_186_1286_0, i_8_186_1300_0,
    i_8_186_1352_0, i_8_186_1360_0, i_8_186_1362_0, i_8_186_1384_0,
    i_8_186_1423_0, i_8_186_1441_0, i_8_186_1442_0, i_8_186_1461_0,
    i_8_186_1462_0, i_8_186_1471_0, i_8_186_1512_0, i_8_186_1559_0,
    i_8_186_1569_0, i_8_186_1570_0, i_8_186_1603_0, i_8_186_1615_0,
    i_8_186_1616_0, i_8_186_1618_0, i_8_186_1642_0, i_8_186_1643_0,
    i_8_186_1644_0, i_8_186_1719_0, i_8_186_1781_0, i_8_186_1783_0,
    i_8_186_1787_0, i_8_186_1822_0, i_8_186_1836_0, i_8_186_1849_0,
    i_8_186_1852_0, i_8_186_1935_0, i_8_186_1954_0, i_8_186_1958_0,
    i_8_186_1981_0, i_8_186_1993_0, i_8_186_2055_0, i_8_186_2077_0,
    i_8_186_2088_0, i_8_186_2120_0, i_8_186_2151_0, i_8_186_2163_0,
    i_8_186_2169_0, i_8_186_2170_0, i_8_186_2212_0, i_8_186_2296_0;
  output o_8_186_0_0;
  assign o_8_186_0_0 = 0;
endmodule



// Benchmark "kernel_8_187" written by ABC on Sun Jul 19 10:06:18 2020

module kernel_8_187 ( 
    i_8_187_23_0, i_8_187_52_0, i_8_187_81_0, i_8_187_93_0, i_8_187_111_0,
    i_8_187_114_0, i_8_187_115_0, i_8_187_117_0, i_8_187_118_0,
    i_8_187_162_0, i_8_187_165_0, i_8_187_166_0, i_8_187_173_0,
    i_8_187_279_0, i_8_187_318_0, i_8_187_346_0, i_8_187_349_0,
    i_8_187_382_0, i_8_187_392_0, i_8_187_433_0, i_8_187_486_0,
    i_8_187_493_0, i_8_187_556_0, i_8_187_562_0, i_8_187_621_0,
    i_8_187_628_0, i_8_187_630_0, i_8_187_666_0, i_8_187_696_0,
    i_8_187_697_0, i_8_187_712_0, i_8_187_715_0, i_8_187_716_0,
    i_8_187_718_0, i_8_187_720_0, i_8_187_762_0, i_8_187_819_0,
    i_8_187_826_0, i_8_187_845_0, i_8_187_846_0, i_8_187_928_0,
    i_8_187_956_0, i_8_187_985_0, i_8_187_996_0, i_8_187_1026_0,
    i_8_187_1057_0, i_8_187_1059_0, i_8_187_1060_0, i_8_187_1061_0,
    i_8_187_1065_0, i_8_187_1080_0, i_8_187_1114_0, i_8_187_1158_0,
    i_8_187_1164_0, i_8_187_1183_0, i_8_187_1226_0, i_8_187_1229_0,
    i_8_187_1258_0, i_8_187_1315_0, i_8_187_1353_0, i_8_187_1359_0,
    i_8_187_1467_0, i_8_187_1471_0, i_8_187_1565_0, i_8_187_1587_0,
    i_8_187_1608_0, i_8_187_1621_0, i_8_187_1642_0, i_8_187_1696_0,
    i_8_187_1699_0, i_8_187_1703_0, i_8_187_1704_0, i_8_187_1705_0,
    i_8_187_1728_0, i_8_187_1734_0, i_8_187_1752_0, i_8_187_1773_0,
    i_8_187_1800_0, i_8_187_1857_0, i_8_187_1860_0, i_8_187_1867_0,
    i_8_187_1885_0, i_8_187_1962_0, i_8_187_1967_0, i_8_187_1983_0,
    i_8_187_1984_0, i_8_187_1986_0, i_8_187_2017_0, i_8_187_2061_0,
    i_8_187_2115_0, i_8_187_2125_0, i_8_187_2142_0, i_8_187_2143_0,
    i_8_187_2145_0, i_8_187_2187_0, i_8_187_2192_0, i_8_187_2224_0,
    i_8_187_2225_0, i_8_187_2282_0, i_8_187_2292_0,
    o_8_187_0_0  );
  input  i_8_187_23_0, i_8_187_52_0, i_8_187_81_0, i_8_187_93_0,
    i_8_187_111_0, i_8_187_114_0, i_8_187_115_0, i_8_187_117_0,
    i_8_187_118_0, i_8_187_162_0, i_8_187_165_0, i_8_187_166_0,
    i_8_187_173_0, i_8_187_279_0, i_8_187_318_0, i_8_187_346_0,
    i_8_187_349_0, i_8_187_382_0, i_8_187_392_0, i_8_187_433_0,
    i_8_187_486_0, i_8_187_493_0, i_8_187_556_0, i_8_187_562_0,
    i_8_187_621_0, i_8_187_628_0, i_8_187_630_0, i_8_187_666_0,
    i_8_187_696_0, i_8_187_697_0, i_8_187_712_0, i_8_187_715_0,
    i_8_187_716_0, i_8_187_718_0, i_8_187_720_0, i_8_187_762_0,
    i_8_187_819_0, i_8_187_826_0, i_8_187_845_0, i_8_187_846_0,
    i_8_187_928_0, i_8_187_956_0, i_8_187_985_0, i_8_187_996_0,
    i_8_187_1026_0, i_8_187_1057_0, i_8_187_1059_0, i_8_187_1060_0,
    i_8_187_1061_0, i_8_187_1065_0, i_8_187_1080_0, i_8_187_1114_0,
    i_8_187_1158_0, i_8_187_1164_0, i_8_187_1183_0, i_8_187_1226_0,
    i_8_187_1229_0, i_8_187_1258_0, i_8_187_1315_0, i_8_187_1353_0,
    i_8_187_1359_0, i_8_187_1467_0, i_8_187_1471_0, i_8_187_1565_0,
    i_8_187_1587_0, i_8_187_1608_0, i_8_187_1621_0, i_8_187_1642_0,
    i_8_187_1696_0, i_8_187_1699_0, i_8_187_1703_0, i_8_187_1704_0,
    i_8_187_1705_0, i_8_187_1728_0, i_8_187_1734_0, i_8_187_1752_0,
    i_8_187_1773_0, i_8_187_1800_0, i_8_187_1857_0, i_8_187_1860_0,
    i_8_187_1867_0, i_8_187_1885_0, i_8_187_1962_0, i_8_187_1967_0,
    i_8_187_1983_0, i_8_187_1984_0, i_8_187_1986_0, i_8_187_2017_0,
    i_8_187_2061_0, i_8_187_2115_0, i_8_187_2125_0, i_8_187_2142_0,
    i_8_187_2143_0, i_8_187_2145_0, i_8_187_2187_0, i_8_187_2192_0,
    i_8_187_2224_0, i_8_187_2225_0, i_8_187_2282_0, i_8_187_2292_0;
  output o_8_187_0_0;
  assign o_8_187_0_0 = 0;
endmodule



// Benchmark "kernel_8_188" written by ABC on Sun Jul 19 10:06:19 2020

module kernel_8_188 ( 
    i_8_188_33_0, i_8_188_53_0, i_8_188_55_0, i_8_188_57_0, i_8_188_63_0,
    i_8_188_86_0, i_8_188_97_0, i_8_188_98_0, i_8_188_141_0, i_8_188_223_0,
    i_8_188_256_0, i_8_188_260_0, i_8_188_313_0, i_8_188_314_0,
    i_8_188_328_0, i_8_188_346_0, i_8_188_362_0, i_8_188_363_0,
    i_8_188_373_0, i_8_188_379_0, i_8_188_439_0, i_8_188_481_0,
    i_8_188_507_0, i_8_188_525_0, i_8_188_528_0, i_8_188_529_0,
    i_8_188_530_0, i_8_188_553_0, i_8_188_556_0, i_8_188_557_0,
    i_8_188_598_0, i_8_188_602_0, i_8_188_633_0, i_8_188_657_0,
    i_8_188_658_0, i_8_188_691_0, i_8_188_692_0, i_8_188_703_0,
    i_8_188_705_0, i_8_188_789_0, i_8_188_800_0, i_8_188_853_0,
    i_8_188_854_0, i_8_188_855_0, i_8_188_880_0, i_8_188_946_0,
    i_8_188_1050_0, i_8_188_1072_0, i_8_188_1113_0, i_8_188_1120_0,
    i_8_188_1123_0, i_8_188_1124_0, i_8_188_1191_0, i_8_188_1223_0,
    i_8_188_1232_0, i_8_188_1263_0, i_8_188_1264_0, i_8_188_1274_0,
    i_8_188_1299_0, i_8_188_1305_0, i_8_188_1307_0, i_8_188_1309_0,
    i_8_188_1317_0, i_8_188_1318_0, i_8_188_1327_0, i_8_188_1331_0,
    i_8_188_1407_0, i_8_188_1450_0, i_8_188_1467_0, i_8_188_1470_0,
    i_8_188_1540_0, i_8_188_1545_0, i_8_188_1564_0, i_8_188_1573_0,
    i_8_188_1574_0, i_8_188_1576_0, i_8_188_1637_0, i_8_188_1675_0,
    i_8_188_1677_0, i_8_188_1678_0, i_8_188_1680_0, i_8_188_1741_0,
    i_8_188_1749_0, i_8_188_1790_0, i_8_188_1795_0, i_8_188_1808_0,
    i_8_188_1879_0, i_8_188_1884_0, i_8_188_1907_0, i_8_188_1995_0,
    i_8_188_1997_0, i_8_188_2031_0, i_8_188_2032_0, i_8_188_2095_0,
    i_8_188_2096_0, i_8_188_2104_0, i_8_188_2105_0, i_8_188_2222_0,
    i_8_188_2260_0, i_8_188_2275_0,
    o_8_188_0_0  );
  input  i_8_188_33_0, i_8_188_53_0, i_8_188_55_0, i_8_188_57_0,
    i_8_188_63_0, i_8_188_86_0, i_8_188_97_0, i_8_188_98_0, i_8_188_141_0,
    i_8_188_223_0, i_8_188_256_0, i_8_188_260_0, i_8_188_313_0,
    i_8_188_314_0, i_8_188_328_0, i_8_188_346_0, i_8_188_362_0,
    i_8_188_363_0, i_8_188_373_0, i_8_188_379_0, i_8_188_439_0,
    i_8_188_481_0, i_8_188_507_0, i_8_188_525_0, i_8_188_528_0,
    i_8_188_529_0, i_8_188_530_0, i_8_188_553_0, i_8_188_556_0,
    i_8_188_557_0, i_8_188_598_0, i_8_188_602_0, i_8_188_633_0,
    i_8_188_657_0, i_8_188_658_0, i_8_188_691_0, i_8_188_692_0,
    i_8_188_703_0, i_8_188_705_0, i_8_188_789_0, i_8_188_800_0,
    i_8_188_853_0, i_8_188_854_0, i_8_188_855_0, i_8_188_880_0,
    i_8_188_946_0, i_8_188_1050_0, i_8_188_1072_0, i_8_188_1113_0,
    i_8_188_1120_0, i_8_188_1123_0, i_8_188_1124_0, i_8_188_1191_0,
    i_8_188_1223_0, i_8_188_1232_0, i_8_188_1263_0, i_8_188_1264_0,
    i_8_188_1274_0, i_8_188_1299_0, i_8_188_1305_0, i_8_188_1307_0,
    i_8_188_1309_0, i_8_188_1317_0, i_8_188_1318_0, i_8_188_1327_0,
    i_8_188_1331_0, i_8_188_1407_0, i_8_188_1450_0, i_8_188_1467_0,
    i_8_188_1470_0, i_8_188_1540_0, i_8_188_1545_0, i_8_188_1564_0,
    i_8_188_1573_0, i_8_188_1574_0, i_8_188_1576_0, i_8_188_1637_0,
    i_8_188_1675_0, i_8_188_1677_0, i_8_188_1678_0, i_8_188_1680_0,
    i_8_188_1741_0, i_8_188_1749_0, i_8_188_1790_0, i_8_188_1795_0,
    i_8_188_1808_0, i_8_188_1879_0, i_8_188_1884_0, i_8_188_1907_0,
    i_8_188_1995_0, i_8_188_1997_0, i_8_188_2031_0, i_8_188_2032_0,
    i_8_188_2095_0, i_8_188_2096_0, i_8_188_2104_0, i_8_188_2105_0,
    i_8_188_2222_0, i_8_188_2260_0, i_8_188_2275_0;
  output o_8_188_0_0;
  assign o_8_188_0_0 = 0;
endmodule



// Benchmark "kernel_8_189" written by ABC on Sun Jul 19 10:06:20 2020

module kernel_8_189 ( 
    i_8_189_61_0, i_8_189_80_0, i_8_189_87_0, i_8_189_88_0, i_8_189_160_0,
    i_8_189_165_0, i_8_189_174_0, i_8_189_177_0, i_8_189_196_0,
    i_8_189_256_0, i_8_189_268_0, i_8_189_309_0, i_8_189_312_0,
    i_8_189_313_0, i_8_189_331_0, i_8_189_356_0, i_8_189_376_0,
    i_8_189_395_0, i_8_189_418_0, i_8_189_517_0, i_8_189_520_0,
    i_8_189_522_0, i_8_189_529_0, i_8_189_530_0, i_8_189_535_0,
    i_8_189_550_0, i_8_189_652_0, i_8_189_696_0, i_8_189_701_0,
    i_8_189_704_0, i_8_189_709_0, i_8_189_718_0, i_8_189_751_0,
    i_8_189_832_0, i_8_189_835_0, i_8_189_841_0, i_8_189_853_0,
    i_8_189_862_0, i_8_189_873_0, i_8_189_916_0, i_8_189_933_0,
    i_8_189_940_0, i_8_189_1014_0, i_8_189_1043_0, i_8_189_1067_0,
    i_8_189_1111_0, i_8_189_1131_0, i_8_189_1158_0, i_8_189_1177_0,
    i_8_189_1204_0, i_8_189_1264_0, i_8_189_1273_0, i_8_189_1299_0,
    i_8_189_1300_0, i_8_189_1309_0, i_8_189_1317_0, i_8_189_1321_0,
    i_8_189_1348_0, i_8_189_1353_0, i_8_189_1366_0, i_8_189_1375_0,
    i_8_189_1381_0, i_8_189_1434_0, i_8_189_1446_0, i_8_189_1454_0,
    i_8_189_1498_0, i_8_189_1537_0, i_8_189_1553_0, i_8_189_1560_0,
    i_8_189_1618_0, i_8_189_1619_0, i_8_189_1668_0, i_8_189_1690_0,
    i_8_189_1707_0, i_8_189_1709_0, i_8_189_1768_0, i_8_189_1771_0,
    i_8_189_1818_0, i_8_189_1822_0, i_8_189_1824_0, i_8_189_1826_0,
    i_8_189_1840_0, i_8_189_1864_0, i_8_189_1870_0, i_8_189_1871_0,
    i_8_189_1995_0, i_8_189_2058_0, i_8_189_2112_0, i_8_189_2137_0,
    i_8_189_2139_0, i_8_189_2141_0, i_8_189_2147_0, i_8_189_2148_0,
    i_8_189_2151_0, i_8_189_2174_0, i_8_189_2185_0, i_8_189_2229_0,
    i_8_189_2240_0, i_8_189_2258_0, i_8_189_2274_0,
    o_8_189_0_0  );
  input  i_8_189_61_0, i_8_189_80_0, i_8_189_87_0, i_8_189_88_0,
    i_8_189_160_0, i_8_189_165_0, i_8_189_174_0, i_8_189_177_0,
    i_8_189_196_0, i_8_189_256_0, i_8_189_268_0, i_8_189_309_0,
    i_8_189_312_0, i_8_189_313_0, i_8_189_331_0, i_8_189_356_0,
    i_8_189_376_0, i_8_189_395_0, i_8_189_418_0, i_8_189_517_0,
    i_8_189_520_0, i_8_189_522_0, i_8_189_529_0, i_8_189_530_0,
    i_8_189_535_0, i_8_189_550_0, i_8_189_652_0, i_8_189_696_0,
    i_8_189_701_0, i_8_189_704_0, i_8_189_709_0, i_8_189_718_0,
    i_8_189_751_0, i_8_189_832_0, i_8_189_835_0, i_8_189_841_0,
    i_8_189_853_0, i_8_189_862_0, i_8_189_873_0, i_8_189_916_0,
    i_8_189_933_0, i_8_189_940_0, i_8_189_1014_0, i_8_189_1043_0,
    i_8_189_1067_0, i_8_189_1111_0, i_8_189_1131_0, i_8_189_1158_0,
    i_8_189_1177_0, i_8_189_1204_0, i_8_189_1264_0, i_8_189_1273_0,
    i_8_189_1299_0, i_8_189_1300_0, i_8_189_1309_0, i_8_189_1317_0,
    i_8_189_1321_0, i_8_189_1348_0, i_8_189_1353_0, i_8_189_1366_0,
    i_8_189_1375_0, i_8_189_1381_0, i_8_189_1434_0, i_8_189_1446_0,
    i_8_189_1454_0, i_8_189_1498_0, i_8_189_1537_0, i_8_189_1553_0,
    i_8_189_1560_0, i_8_189_1618_0, i_8_189_1619_0, i_8_189_1668_0,
    i_8_189_1690_0, i_8_189_1707_0, i_8_189_1709_0, i_8_189_1768_0,
    i_8_189_1771_0, i_8_189_1818_0, i_8_189_1822_0, i_8_189_1824_0,
    i_8_189_1826_0, i_8_189_1840_0, i_8_189_1864_0, i_8_189_1870_0,
    i_8_189_1871_0, i_8_189_1995_0, i_8_189_2058_0, i_8_189_2112_0,
    i_8_189_2137_0, i_8_189_2139_0, i_8_189_2141_0, i_8_189_2147_0,
    i_8_189_2148_0, i_8_189_2151_0, i_8_189_2174_0, i_8_189_2185_0,
    i_8_189_2229_0, i_8_189_2240_0, i_8_189_2258_0, i_8_189_2274_0;
  output o_8_189_0_0;
  assign o_8_189_0_0 = 0;
endmodule



// Benchmark "kernel_8_190" written by ABC on Sun Jul 19 10:06:21 2020

module kernel_8_190 ( 
    i_8_190_71_0, i_8_190_142_0, i_8_190_143_0, i_8_190_154_0,
    i_8_190_173_0, i_8_190_202_0, i_8_190_203_0, i_8_190_205_0,
    i_8_190_208_0, i_8_190_268_0, i_8_190_275_0, i_8_190_278_0,
    i_8_190_341_0, i_8_190_345_0, i_8_190_346_0, i_8_190_348_0,
    i_8_190_377_0, i_8_190_380_0, i_8_190_495_0, i_8_190_496_0,
    i_8_190_497_0, i_8_190_522_0, i_8_190_523_0, i_8_190_524_0,
    i_8_190_553_0, i_8_190_555_0, i_8_190_607_0, i_8_190_609_0,
    i_8_190_620_0, i_8_190_652_0, i_8_190_696_0, i_8_190_700_0,
    i_8_190_837_0, i_8_190_838_0, i_8_190_839_0, i_8_190_841_0,
    i_8_190_868_0, i_8_190_879_0, i_8_190_881_0, i_8_190_980_0,
    i_8_190_1033_0, i_8_190_1049_0, i_8_190_1057_0, i_8_190_1088_0,
    i_8_190_1110_0, i_8_190_1128_0, i_8_190_1204_0, i_8_190_1281_0,
    i_8_190_1284_0, i_8_190_1285_0, i_8_190_1286_0, i_8_190_1302_0,
    i_8_190_1303_0, i_8_190_1322_0, i_8_190_1343_0, i_8_190_1396_0,
    i_8_190_1402_0, i_8_190_1430_0, i_8_190_1436_0, i_8_190_1528_0,
    i_8_190_1620_0, i_8_190_1708_0, i_8_190_1714_0, i_8_190_1727_0,
    i_8_190_1747_0, i_8_190_1762_0, i_8_190_1766_0, i_8_190_1778_0,
    i_8_190_1795_0, i_8_190_1798_0, i_8_190_1799_0, i_8_190_1800_0,
    i_8_190_1802_0, i_8_190_1803_0, i_8_190_1804_0, i_8_190_1805_0,
    i_8_190_1808_0, i_8_190_1826_0, i_8_190_1858_0, i_8_190_1861_0,
    i_8_190_1864_0, i_8_190_1865_0, i_8_190_1914_0, i_8_190_1915_0,
    i_8_190_1964_0, i_8_190_1970_0, i_8_190_1980_0, i_8_190_1983_0,
    i_8_190_2046_0, i_8_190_2047_0, i_8_190_2049_0, i_8_190_2065_0,
    i_8_190_2073_0, i_8_190_2125_0, i_8_190_2128_0, i_8_190_2237_0,
    i_8_190_2244_0, i_8_190_2286_0, i_8_190_2287_0, i_8_190_2289_0,
    o_8_190_0_0  );
  input  i_8_190_71_0, i_8_190_142_0, i_8_190_143_0, i_8_190_154_0,
    i_8_190_173_0, i_8_190_202_0, i_8_190_203_0, i_8_190_205_0,
    i_8_190_208_0, i_8_190_268_0, i_8_190_275_0, i_8_190_278_0,
    i_8_190_341_0, i_8_190_345_0, i_8_190_346_0, i_8_190_348_0,
    i_8_190_377_0, i_8_190_380_0, i_8_190_495_0, i_8_190_496_0,
    i_8_190_497_0, i_8_190_522_0, i_8_190_523_0, i_8_190_524_0,
    i_8_190_553_0, i_8_190_555_0, i_8_190_607_0, i_8_190_609_0,
    i_8_190_620_0, i_8_190_652_0, i_8_190_696_0, i_8_190_700_0,
    i_8_190_837_0, i_8_190_838_0, i_8_190_839_0, i_8_190_841_0,
    i_8_190_868_0, i_8_190_879_0, i_8_190_881_0, i_8_190_980_0,
    i_8_190_1033_0, i_8_190_1049_0, i_8_190_1057_0, i_8_190_1088_0,
    i_8_190_1110_0, i_8_190_1128_0, i_8_190_1204_0, i_8_190_1281_0,
    i_8_190_1284_0, i_8_190_1285_0, i_8_190_1286_0, i_8_190_1302_0,
    i_8_190_1303_0, i_8_190_1322_0, i_8_190_1343_0, i_8_190_1396_0,
    i_8_190_1402_0, i_8_190_1430_0, i_8_190_1436_0, i_8_190_1528_0,
    i_8_190_1620_0, i_8_190_1708_0, i_8_190_1714_0, i_8_190_1727_0,
    i_8_190_1747_0, i_8_190_1762_0, i_8_190_1766_0, i_8_190_1778_0,
    i_8_190_1795_0, i_8_190_1798_0, i_8_190_1799_0, i_8_190_1800_0,
    i_8_190_1802_0, i_8_190_1803_0, i_8_190_1804_0, i_8_190_1805_0,
    i_8_190_1808_0, i_8_190_1826_0, i_8_190_1858_0, i_8_190_1861_0,
    i_8_190_1864_0, i_8_190_1865_0, i_8_190_1914_0, i_8_190_1915_0,
    i_8_190_1964_0, i_8_190_1970_0, i_8_190_1980_0, i_8_190_1983_0,
    i_8_190_2046_0, i_8_190_2047_0, i_8_190_2049_0, i_8_190_2065_0,
    i_8_190_2073_0, i_8_190_2125_0, i_8_190_2128_0, i_8_190_2237_0,
    i_8_190_2244_0, i_8_190_2286_0, i_8_190_2287_0, i_8_190_2289_0;
  output o_8_190_0_0;
  assign o_8_190_0_0 = ~((~i_8_190_1865_0 & ((~i_8_190_1088_0 & ((~i_8_190_143_0 & ~i_8_190_154_0 & ~i_8_190_1803_0 & ((~i_8_190_173_0 & ~i_8_190_202_0 & ~i_8_190_275_0 & ~i_8_190_278_0 & ~i_8_190_380_0 & ~i_8_190_496_0 & ~i_8_190_555_0 & ~i_8_190_980_0 & ~i_8_190_1322_0 & ~i_8_190_1708_0 & ~i_8_190_1727_0 & ~i_8_190_1915_0) | (~i_8_190_497_0 & i_8_190_838_0 & ~i_8_190_1302_0 & ~i_8_190_1528_0 & ~i_8_190_1795_0 & ~i_8_190_1799_0 & ~i_8_190_2046_0 & ~i_8_190_2047_0))) | (i_8_190_1284_0 & ~i_8_190_1915_0 & ((~i_8_190_208_0 & ~i_8_190_268_0 & ~i_8_190_1528_0 & i_8_190_1762_0 & ~i_8_190_1799_0 & ~i_8_190_1864_0 & ~i_8_190_1914_0 & ~i_8_190_2047_0) | (~i_8_190_523_0 & ~i_8_190_1430_0 & ~i_8_190_1727_0 & ~i_8_190_1798_0 & ~i_8_190_1805_0 & ~i_8_190_2065_0))) | (~i_8_190_142_0 & ~i_8_190_496_0 & ~i_8_190_700_0 & ~i_8_190_1110_0 & ~i_8_190_1303_0 & i_8_190_1436_0 & ~i_8_190_1727_0 & ~i_8_190_1762_0 & ~i_8_190_1980_0))) | (~i_8_190_202_0 & ((~i_8_190_523_0 & ~i_8_190_524_0 & i_8_190_607_0 & ~i_8_190_620_0 & i_8_190_1747_0) | (~i_8_190_205_0 & ~i_8_190_268_0 & ~i_8_190_275_0 & ~i_8_190_495_0 & ~i_8_190_555_0 & ~i_8_190_839_0 & ~i_8_190_1286_0 & ~i_8_190_1430_0 & ~i_8_190_1727_0 & ~i_8_190_1799_0 & i_8_190_1804_0 & ~i_8_190_1914_0 & ~i_8_190_1915_0 & ~i_8_190_1964_0 & ~i_8_190_2065_0 & ~i_8_190_2287_0))) | (~i_8_190_203_0 & ((i_8_190_837_0 & ~i_8_190_1430_0 & ~i_8_190_1795_0 & ~i_8_190_1799_0 & ~i_8_190_1864_0 & ~i_8_190_2049_0) | (~i_8_190_208_0 & i_8_190_553_0 & i_8_190_1285_0 & i_8_190_1436_0 & ~i_8_190_1528_0 & i_8_190_1778_0 & ~i_8_190_1800_0 & ~i_8_190_2065_0 & ~i_8_190_2289_0))) | (~i_8_190_1343_0 & ~i_8_190_1798_0 & ~i_8_190_1799_0 & ~i_8_190_1914_0 & ~i_8_190_2049_0 & ((~i_8_190_205_0 & ~i_8_190_208_0 & ~i_8_190_275_0 & ~i_8_190_278_0 & ~i_8_190_620_0 & ~i_8_190_980_0 & ~i_8_190_1284_0 & ~i_8_190_1402_0 & ~i_8_190_1620_0 & ~i_8_190_1714_0 & ~i_8_190_1747_0 & ~i_8_190_1795_0 & ~i_8_190_1864_0 & ~i_8_190_1980_0 & ~i_8_190_2046_0 & ~i_8_190_2073_0 & ~i_8_190_2237_0 & ~i_8_190_2286_0) | (~i_8_190_71_0 & ~i_8_190_341_0 & ~i_8_190_495_0 & ~i_8_190_497_0 & ~i_8_190_1110_0 & ~i_8_190_1204_0 & ~i_8_190_1805_0 & ~i_8_190_2287_0))))) | (~i_8_190_203_0 & ((~i_8_190_142_0 & ((~i_8_190_71_0 & ~i_8_190_173_0 & ~i_8_190_341_0 & ~i_8_190_523_0 & ~i_8_190_555_0 & ~i_8_190_607_0 & ~i_8_190_1088_0 & ~i_8_190_1204_0 & ~i_8_190_1343_0 & ~i_8_190_1714_0 & ~i_8_190_1800_0 & ~i_8_190_1803_0 & ~i_8_190_2065_0) | (~i_8_190_495_0 & i_8_190_839_0 & i_8_190_2125_0 & ~i_8_190_2286_0))) | (~i_8_190_278_0 & ~i_8_190_497_0 & ~i_8_190_1799_0 & ((~i_8_190_495_0 & ~i_8_190_553_0 & ~i_8_190_696_0 & ~i_8_190_838_0 & i_8_190_1057_0 & ~i_8_190_1285_0 & ~i_8_190_1798_0 & ~i_8_190_1914_0) | (~i_8_190_275_0 & ~i_8_190_380_0 & ~i_8_190_522_0 & ~i_8_190_555_0 & ~i_8_190_980_0 & ~i_8_190_1302_0 & ~i_8_190_1343_0 & ~i_8_190_1620_0 & ~i_8_190_1804_0 & ~i_8_190_1808_0 & ~i_8_190_1915_0 & ~i_8_190_2046_0 & ~i_8_190_2289_0))))) | (~i_8_190_275_0 & ((~i_8_190_71_0 & ((~i_8_190_202_0 & ~i_8_190_522_0 & i_8_190_881_0 & i_8_190_1286_0 & ~i_8_190_1396_0 & ~i_8_190_1800_0 & ~i_8_190_2047_0) | (~i_8_190_205_0 & ~i_8_190_268_0 & ~i_8_190_523_0 & ~i_8_190_553_0 & ~i_8_190_838_0 & ~i_8_190_1057_0 & ~i_8_190_1303_0 & ~i_8_190_1708_0 & ~i_8_190_1747_0 & ~i_8_190_1766_0 & ~i_8_190_1802_0 & ~i_8_190_1805_0 & ~i_8_190_1808_0 & ~i_8_190_1914_0 & ~i_8_190_1980_0 & ~i_8_190_2073_0))) | (~i_8_190_268_0 & ~i_8_190_2065_0 & ((~i_8_190_341_0 & ~i_8_190_497_0 & ~i_8_190_1088_0 & ~i_8_190_1322_0 & i_8_190_1396_0 & ~i_8_190_1436_0 & ~i_8_190_1803_0) | (~i_8_190_173_0 & ~i_8_190_524_0 & ~i_8_190_620_0 & ~i_8_190_700_0 & ~i_8_190_980_0 & ~i_8_190_1057_0 & ~i_8_190_1110_0 & ~i_8_190_1128_0 & ~i_8_190_1281_0 & ~i_8_190_1430_0 & ~i_8_190_1528_0 & ~i_8_190_1808_0 & ~i_8_190_2237_0 & ~i_8_190_2244_0))) | (~i_8_190_497_0 & ~i_8_190_1322_0 & ~i_8_190_1861_0 & ((~i_8_190_202_0 & ~i_8_190_496_0 & i_8_190_523_0 & ~i_8_190_609_0 & ~i_8_190_838_0 & ~i_8_190_868_0 & ~i_8_190_1281_0 & ~i_8_190_1343_0 & ~i_8_190_1396_0 & ~i_8_190_1799_0 & ~i_8_190_2049_0) | (i_8_190_609_0 & ~i_8_190_1033_0 & i_8_190_1128_0 & ~i_8_190_1620_0 & ~i_8_190_1766_0 & ~i_8_190_1915_0 & ~i_8_190_2287_0))))) | (i_8_190_522_0 & ((~i_8_190_380_0 & ~i_8_190_497_0 & ~i_8_190_553_0 & ~i_8_190_1747_0 & i_8_190_1858_0) | (~i_8_190_524_0 & i_8_190_609_0 & i_8_190_879_0 & ~i_8_190_1858_0 & ~i_8_190_2065_0 & ~i_8_190_2286_0))) | (~i_8_190_380_0 & ~i_8_190_838_0 & ~i_8_190_1778_0 & ((~i_8_190_205_0 & i_8_190_700_0 & ~i_8_190_881_0 & ~i_8_190_1281_0 & i_8_190_1286_0 & i_8_190_1970_0) | (~i_8_190_278_0 & ~i_8_190_1204_0 & i_8_190_1281_0 & ~i_8_190_1302_0 & ~i_8_190_1708_0 & ~i_8_190_1799_0 & ~i_8_190_2065_0 & ~i_8_190_2073_0 & ~i_8_190_2286_0 & ~i_8_190_2289_0))) | (~i_8_190_1799_0 & ((~i_8_190_495_0 & ((~i_8_190_173_0 & ~i_8_190_620_0 & i_8_190_841_0 & i_8_190_1049_0 & ~i_8_190_1798_0 & ~i_8_190_1980_0 & ~i_8_190_2125_0) | (~i_8_190_205_0 & ~i_8_190_278_0 & ~i_8_190_1128_0 & ~i_8_190_1303_0 & ~i_8_190_1402_0 & ~i_8_190_1714_0 & ~i_8_190_1864_0 & i_8_190_2244_0))) | (~i_8_190_173_0 & ~i_8_190_1802_0 & ~i_8_190_2046_0 & ((~i_8_190_71_0 & ~i_8_190_143_0 & ~i_8_190_496_0 & ~i_8_190_607_0 & ~i_8_190_696_0 & ~i_8_190_881_0 & ~i_8_190_1057_0 & ~i_8_190_1204_0 & ~i_8_190_1281_0 & ~i_8_190_1727_0 & ~i_8_190_1804_0 & ~i_8_190_1861_0 & ~i_8_190_2049_0 & ~i_8_190_2065_0) | (~i_8_190_522_0 & ~i_8_190_620_0 & ~i_8_190_1303_0 & ~i_8_190_1343_0 & ~i_8_190_1714_0 & ~i_8_190_1803_0 & i_8_190_1861_0 & ~i_8_190_1915_0 & ~i_8_190_2289_0))) | (~i_8_190_278_0 & ~i_8_190_497_0 & ~i_8_190_1088_0 & ((~i_8_190_208_0 & i_8_190_1286_0 & ~i_8_190_1322_0 & ~i_8_190_1803_0 & i_8_190_1861_0 & ~i_8_190_2049_0) | (~i_8_190_524_0 & i_8_190_881_0 & ~i_8_190_1343_0 & ~i_8_190_1430_0 & ~i_8_190_1708_0 & ~i_8_190_1795_0 & ~i_8_190_1798_0 & ~i_8_190_2065_0 & ~i_8_190_2128_0))))) | (~i_8_190_205_0 & ((i_8_190_345_0 & i_8_190_696_0 & ~i_8_190_1343_0 & ~i_8_190_1396_0 & ~i_8_190_1915_0 & ~i_8_190_2047_0) | (~i_8_190_497_0 & i_8_190_607_0 & ~i_8_190_841_0 & ~i_8_190_868_0 & ~i_8_190_1204_0 & ~i_8_190_1805_0 & ~i_8_190_1826_0 & ~i_8_190_1864_0 & ~i_8_190_1914_0 & ~i_8_190_2065_0))) | (~i_8_190_523_0 & ((~i_8_190_278_0 & ~i_8_190_1057_0 & ((~i_8_190_377_0 & ~i_8_190_497_0 & ~i_8_190_841_0 & ~i_8_190_1430_0 & ~i_8_190_1804_0 & i_8_190_1805_0) | (i_8_190_143_0 & ~i_8_190_881_0 & i_8_190_980_0 & ~i_8_190_1302_0 & ~i_8_190_1528_0 & ~i_8_190_1805_0))) | (~i_8_190_497_0 & ~i_8_190_1795_0 & i_8_190_1983_0 & ~i_8_190_2049_0))) | (~i_8_190_2046_0 & ((i_8_190_346_0 & ~i_8_190_495_0 & ~i_8_190_700_0 & ~i_8_190_1204_0 & ~i_8_190_1322_0 & ~i_8_190_1804_0 & ~i_8_190_1808_0 & ~i_8_190_1858_0 & ~i_8_190_1964_0 & ~i_8_190_2047_0 & ~i_8_190_2049_0) | (~i_8_190_1864_0 & i_8_190_2065_0 & i_8_190_2073_0 & i_8_190_2286_0))));
endmodule



// Benchmark "kernel_8_191" written by ABC on Sun Jul 19 10:06:22 2020

module kernel_8_191 ( 
    i_8_191_22_0, i_8_191_25_0, i_8_191_52_0, i_8_191_54_0, i_8_191_60_0,
    i_8_191_138_0, i_8_191_160_0, i_8_191_193_0, i_8_191_262_0,
    i_8_191_336_0, i_8_191_341_0, i_8_191_354_0, i_8_191_376_0,
    i_8_191_385_0, i_8_191_403_0, i_8_191_457_0, i_8_191_499_0,
    i_8_191_529_0, i_8_191_555_0, i_8_191_573_0, i_8_191_604_0,
    i_8_191_607_0, i_8_191_609_0, i_8_191_653_0, i_8_191_675_0,
    i_8_191_678_0, i_8_191_688_0, i_8_191_798_0, i_8_191_799_0,
    i_8_191_837_0, i_8_191_838_0, i_8_191_843_0, i_8_191_849_0,
    i_8_191_881_0, i_8_191_922_0, i_8_191_924_0, i_8_191_933_0,
    i_8_191_968_0, i_8_191_970_0, i_8_191_991_0, i_8_191_993_0,
    i_8_191_995_0, i_8_191_1024_0, i_8_191_1043_0, i_8_191_1072_0,
    i_8_191_1075_0, i_8_191_1101_0, i_8_191_1112_0, i_8_191_1140_0,
    i_8_191_1155_0, i_8_191_1173_0, i_8_191_1194_0, i_8_191_1229_0,
    i_8_191_1263_0, i_8_191_1267_0, i_8_191_1284_0, i_8_191_1300_0,
    i_8_191_1301_0, i_8_191_1328_0, i_8_191_1331_0, i_8_191_1372_0,
    i_8_191_1384_0, i_8_191_1430_0, i_8_191_1442_0, i_8_191_1470_0,
    i_8_191_1473_0, i_8_191_1488_0, i_8_191_1527_0, i_8_191_1569_0,
    i_8_191_1570_0, i_8_191_1579_0, i_8_191_1609_0, i_8_191_1610_0,
    i_8_191_1624_0, i_8_191_1625_0, i_8_191_1629_0, i_8_191_1632_0,
    i_8_191_1644_0, i_8_191_1649_0, i_8_191_1700_0, i_8_191_1766_0,
    i_8_191_1788_0, i_8_191_1797_0, i_8_191_1818_0, i_8_191_1824_0,
    i_8_191_1828_0, i_8_191_1839_0, i_8_191_1893_0, i_8_191_1894_0,
    i_8_191_1942_0, i_8_191_1996_0, i_8_191_2019_0, i_8_191_2028_0,
    i_8_191_2112_0, i_8_191_2113_0, i_8_191_2152_0, i_8_191_2167_0,
    i_8_191_2231_0, i_8_191_2235_0, i_8_191_2241_0,
    o_8_191_0_0  );
  input  i_8_191_22_0, i_8_191_25_0, i_8_191_52_0, i_8_191_54_0,
    i_8_191_60_0, i_8_191_138_0, i_8_191_160_0, i_8_191_193_0,
    i_8_191_262_0, i_8_191_336_0, i_8_191_341_0, i_8_191_354_0,
    i_8_191_376_0, i_8_191_385_0, i_8_191_403_0, i_8_191_457_0,
    i_8_191_499_0, i_8_191_529_0, i_8_191_555_0, i_8_191_573_0,
    i_8_191_604_0, i_8_191_607_0, i_8_191_609_0, i_8_191_653_0,
    i_8_191_675_0, i_8_191_678_0, i_8_191_688_0, i_8_191_798_0,
    i_8_191_799_0, i_8_191_837_0, i_8_191_838_0, i_8_191_843_0,
    i_8_191_849_0, i_8_191_881_0, i_8_191_922_0, i_8_191_924_0,
    i_8_191_933_0, i_8_191_968_0, i_8_191_970_0, i_8_191_991_0,
    i_8_191_993_0, i_8_191_995_0, i_8_191_1024_0, i_8_191_1043_0,
    i_8_191_1072_0, i_8_191_1075_0, i_8_191_1101_0, i_8_191_1112_0,
    i_8_191_1140_0, i_8_191_1155_0, i_8_191_1173_0, i_8_191_1194_0,
    i_8_191_1229_0, i_8_191_1263_0, i_8_191_1267_0, i_8_191_1284_0,
    i_8_191_1300_0, i_8_191_1301_0, i_8_191_1328_0, i_8_191_1331_0,
    i_8_191_1372_0, i_8_191_1384_0, i_8_191_1430_0, i_8_191_1442_0,
    i_8_191_1470_0, i_8_191_1473_0, i_8_191_1488_0, i_8_191_1527_0,
    i_8_191_1569_0, i_8_191_1570_0, i_8_191_1579_0, i_8_191_1609_0,
    i_8_191_1610_0, i_8_191_1624_0, i_8_191_1625_0, i_8_191_1629_0,
    i_8_191_1632_0, i_8_191_1644_0, i_8_191_1649_0, i_8_191_1700_0,
    i_8_191_1766_0, i_8_191_1788_0, i_8_191_1797_0, i_8_191_1818_0,
    i_8_191_1824_0, i_8_191_1828_0, i_8_191_1839_0, i_8_191_1893_0,
    i_8_191_1894_0, i_8_191_1942_0, i_8_191_1996_0, i_8_191_2019_0,
    i_8_191_2028_0, i_8_191_2112_0, i_8_191_2113_0, i_8_191_2152_0,
    i_8_191_2167_0, i_8_191_2231_0, i_8_191_2235_0, i_8_191_2241_0;
  output o_8_191_0_0;
  assign o_8_191_0_0 = 0;
endmodule



// Benchmark "kernel_8_192" written by ABC on Sun Jul 19 10:06:23 2020

module kernel_8_192 ( 
    i_8_192_33_0, i_8_192_88_0, i_8_192_114_0, i_8_192_266_0,
    i_8_192_293_0, i_8_192_374_0, i_8_192_377_0, i_8_192_383_0,
    i_8_192_386_0, i_8_192_440_0, i_8_192_463_0, i_8_192_476_0,
    i_8_192_482_0, i_8_192_485_0, i_8_192_500_0, i_8_192_524_0,
    i_8_192_530_0, i_8_192_571_0, i_8_192_574_0, i_8_192_616_0,
    i_8_192_617_0, i_8_192_624_0, i_8_192_634_0, i_8_192_674_0,
    i_8_192_760_0, i_8_192_762_0, i_8_192_781_0, i_8_192_787_0,
    i_8_192_826_0, i_8_192_841_0, i_8_192_878_0, i_8_192_886_0,
    i_8_192_895_0, i_8_192_936_0, i_8_192_939_0, i_8_192_945_0,
    i_8_192_946_0, i_8_192_995_0, i_8_192_1011_0, i_8_192_1013_0,
    i_8_192_1030_0, i_8_192_1114_0, i_8_192_1124_0, i_8_192_1140_0,
    i_8_192_1159_0, i_8_192_1192_0, i_8_192_1222_0, i_8_192_1237_0,
    i_8_192_1259_0, i_8_192_1264_0, i_8_192_1282_0, i_8_192_1283_0,
    i_8_192_1284_0, i_8_192_1285_0, i_8_192_1305_0, i_8_192_1306_0,
    i_8_192_1328_0, i_8_192_1331_0, i_8_192_1346_0, i_8_192_1438_0,
    i_8_192_1439_0, i_8_192_1441_0, i_8_192_1453_0, i_8_192_1470_0,
    i_8_192_1509_0, i_8_192_1534_0, i_8_192_1535_0, i_8_192_1544_0,
    i_8_192_1565_0, i_8_192_1632_0, i_8_192_1655_0, i_8_192_1681_0,
    i_8_192_1706_0, i_8_192_1732_0, i_8_192_1733_0, i_8_192_1742_0,
    i_8_192_1787_0, i_8_192_1841_0, i_8_192_1857_0, i_8_192_1859_0,
    i_8_192_1866_0, i_8_192_1867_0, i_8_192_1884_0, i_8_192_1885_0,
    i_8_192_1918_0, i_8_192_1919_0, i_8_192_1949_0, i_8_192_1952_0,
    i_8_192_1966_0, i_8_192_1967_0, i_8_192_2056_0, i_8_192_2111_0,
    i_8_192_2127_0, i_8_192_2128_0, i_8_192_2143_0, i_8_192_2156_0,
    i_8_192_2191_0, i_8_192_2192_0, i_8_192_2214_0, i_8_192_2276_0,
    o_8_192_0_0  );
  input  i_8_192_33_0, i_8_192_88_0, i_8_192_114_0, i_8_192_266_0,
    i_8_192_293_0, i_8_192_374_0, i_8_192_377_0, i_8_192_383_0,
    i_8_192_386_0, i_8_192_440_0, i_8_192_463_0, i_8_192_476_0,
    i_8_192_482_0, i_8_192_485_0, i_8_192_500_0, i_8_192_524_0,
    i_8_192_530_0, i_8_192_571_0, i_8_192_574_0, i_8_192_616_0,
    i_8_192_617_0, i_8_192_624_0, i_8_192_634_0, i_8_192_674_0,
    i_8_192_760_0, i_8_192_762_0, i_8_192_781_0, i_8_192_787_0,
    i_8_192_826_0, i_8_192_841_0, i_8_192_878_0, i_8_192_886_0,
    i_8_192_895_0, i_8_192_936_0, i_8_192_939_0, i_8_192_945_0,
    i_8_192_946_0, i_8_192_995_0, i_8_192_1011_0, i_8_192_1013_0,
    i_8_192_1030_0, i_8_192_1114_0, i_8_192_1124_0, i_8_192_1140_0,
    i_8_192_1159_0, i_8_192_1192_0, i_8_192_1222_0, i_8_192_1237_0,
    i_8_192_1259_0, i_8_192_1264_0, i_8_192_1282_0, i_8_192_1283_0,
    i_8_192_1284_0, i_8_192_1285_0, i_8_192_1305_0, i_8_192_1306_0,
    i_8_192_1328_0, i_8_192_1331_0, i_8_192_1346_0, i_8_192_1438_0,
    i_8_192_1439_0, i_8_192_1441_0, i_8_192_1453_0, i_8_192_1470_0,
    i_8_192_1509_0, i_8_192_1534_0, i_8_192_1535_0, i_8_192_1544_0,
    i_8_192_1565_0, i_8_192_1632_0, i_8_192_1655_0, i_8_192_1681_0,
    i_8_192_1706_0, i_8_192_1732_0, i_8_192_1733_0, i_8_192_1742_0,
    i_8_192_1787_0, i_8_192_1841_0, i_8_192_1857_0, i_8_192_1859_0,
    i_8_192_1866_0, i_8_192_1867_0, i_8_192_1884_0, i_8_192_1885_0,
    i_8_192_1918_0, i_8_192_1919_0, i_8_192_1949_0, i_8_192_1952_0,
    i_8_192_1966_0, i_8_192_1967_0, i_8_192_2056_0, i_8_192_2111_0,
    i_8_192_2127_0, i_8_192_2128_0, i_8_192_2143_0, i_8_192_2156_0,
    i_8_192_2191_0, i_8_192_2192_0, i_8_192_2214_0, i_8_192_2276_0;
  output o_8_192_0_0;
  assign o_8_192_0_0 = 0;
endmodule



// Benchmark "kernel_8_193" written by ABC on Sun Jul 19 10:06:24 2020

module kernel_8_193 ( 
    i_8_193_33_0, i_8_193_39_0, i_8_193_45_0, i_8_193_55_0, i_8_193_104_0,
    i_8_193_114_0, i_8_193_119_0, i_8_193_190_0, i_8_193_226_0,
    i_8_193_327_0, i_8_193_364_0, i_8_193_367_0, i_8_193_423_0,
    i_8_193_426_0, i_8_193_450_0, i_8_193_481_0, i_8_193_525_0,
    i_8_193_526_0, i_8_193_530_0, i_8_193_549_0, i_8_193_570_0,
    i_8_193_588_0, i_8_193_612_0, i_8_193_659_0, i_8_193_661_0,
    i_8_193_665_0, i_8_193_684_0, i_8_193_695_0, i_8_193_697_0,
    i_8_193_700_0, i_8_193_706_0, i_8_193_747_0, i_8_193_769_0,
    i_8_193_777_0, i_8_193_792_0, i_8_193_832_0, i_8_193_877_0,
    i_8_193_882_0, i_8_193_981_0, i_8_193_990_0, i_8_193_996_0,
    i_8_193_1032_0, i_8_193_1044_0, i_8_193_1128_0, i_8_193_1135_0,
    i_8_193_1138_0, i_8_193_1143_0, i_8_193_1144_0, i_8_193_1148_0,
    i_8_193_1152_0, i_8_193_1188_0, i_8_193_1270_0, i_8_193_1278_0,
    i_8_193_1330_0, i_8_193_1360_0, i_8_193_1362_0, i_8_193_1368_0,
    i_8_193_1393_0, i_8_193_1404_0, i_8_193_1408_0, i_8_193_1413_0,
    i_8_193_1442_0, i_8_193_1480_0, i_8_193_1506_0, i_8_193_1530_0,
    i_8_193_1543_0, i_8_193_1620_0, i_8_193_1630_0, i_8_193_1632_0,
    i_8_193_1639_0, i_8_193_1648_0, i_8_193_1650_0, i_8_193_1668_0,
    i_8_193_1674_0, i_8_193_1701_0, i_8_193_1714_0, i_8_193_1719_0,
    i_8_193_1728_0, i_8_193_1764_0, i_8_193_1777_0, i_8_193_1821_0,
    i_8_193_1881_0, i_8_193_1900_0, i_8_193_1903_0, i_8_193_1935_0,
    i_8_193_1967_0, i_8_193_1971_0, i_8_193_1983_0, i_8_193_1984_0,
    i_8_193_2070_0, i_8_193_2108_0, i_8_193_2133_0, i_8_193_2146_0,
    i_8_193_2149_0, i_8_193_2150_0, i_8_193_2152_0, i_8_193_2227_0,
    i_8_193_2242_0, i_8_193_2244_0, i_8_193_2269_0,
    o_8_193_0_0  );
  input  i_8_193_33_0, i_8_193_39_0, i_8_193_45_0, i_8_193_55_0,
    i_8_193_104_0, i_8_193_114_0, i_8_193_119_0, i_8_193_190_0,
    i_8_193_226_0, i_8_193_327_0, i_8_193_364_0, i_8_193_367_0,
    i_8_193_423_0, i_8_193_426_0, i_8_193_450_0, i_8_193_481_0,
    i_8_193_525_0, i_8_193_526_0, i_8_193_530_0, i_8_193_549_0,
    i_8_193_570_0, i_8_193_588_0, i_8_193_612_0, i_8_193_659_0,
    i_8_193_661_0, i_8_193_665_0, i_8_193_684_0, i_8_193_695_0,
    i_8_193_697_0, i_8_193_700_0, i_8_193_706_0, i_8_193_747_0,
    i_8_193_769_0, i_8_193_777_0, i_8_193_792_0, i_8_193_832_0,
    i_8_193_877_0, i_8_193_882_0, i_8_193_981_0, i_8_193_990_0,
    i_8_193_996_0, i_8_193_1032_0, i_8_193_1044_0, i_8_193_1128_0,
    i_8_193_1135_0, i_8_193_1138_0, i_8_193_1143_0, i_8_193_1144_0,
    i_8_193_1148_0, i_8_193_1152_0, i_8_193_1188_0, i_8_193_1270_0,
    i_8_193_1278_0, i_8_193_1330_0, i_8_193_1360_0, i_8_193_1362_0,
    i_8_193_1368_0, i_8_193_1393_0, i_8_193_1404_0, i_8_193_1408_0,
    i_8_193_1413_0, i_8_193_1442_0, i_8_193_1480_0, i_8_193_1506_0,
    i_8_193_1530_0, i_8_193_1543_0, i_8_193_1620_0, i_8_193_1630_0,
    i_8_193_1632_0, i_8_193_1639_0, i_8_193_1648_0, i_8_193_1650_0,
    i_8_193_1668_0, i_8_193_1674_0, i_8_193_1701_0, i_8_193_1714_0,
    i_8_193_1719_0, i_8_193_1728_0, i_8_193_1764_0, i_8_193_1777_0,
    i_8_193_1821_0, i_8_193_1881_0, i_8_193_1900_0, i_8_193_1903_0,
    i_8_193_1935_0, i_8_193_1967_0, i_8_193_1971_0, i_8_193_1983_0,
    i_8_193_1984_0, i_8_193_2070_0, i_8_193_2108_0, i_8_193_2133_0,
    i_8_193_2146_0, i_8_193_2149_0, i_8_193_2150_0, i_8_193_2152_0,
    i_8_193_2227_0, i_8_193_2242_0, i_8_193_2244_0, i_8_193_2269_0;
  output o_8_193_0_0;
  assign o_8_193_0_0 = 0;
endmodule



// Benchmark "kernel_8_194" written by ABC on Sun Jul 19 10:06:25 2020

module kernel_8_194 ( 
    i_8_194_21_0, i_8_194_42_0, i_8_194_52_0, i_8_194_55_0, i_8_194_58_0,
    i_8_194_89_0, i_8_194_120_0, i_8_194_129_0, i_8_194_183_0,
    i_8_194_184_0, i_8_194_211_0, i_8_194_218_0, i_8_194_241_0,
    i_8_194_262_0, i_8_194_319_0, i_8_194_365_0, i_8_194_369_0,
    i_8_194_427_0, i_8_194_456_0, i_8_194_478_0, i_8_194_535_0,
    i_8_194_543_0, i_8_194_549_0, i_8_194_551_0, i_8_194_593_0,
    i_8_194_611_0, i_8_194_612_0, i_8_194_613_0, i_8_194_634_0,
    i_8_194_643_0, i_8_194_656_0, i_8_194_662_0, i_8_194_665_0,
    i_8_194_730_0, i_8_194_787_0, i_8_194_802_0, i_8_194_804_0,
    i_8_194_832_0, i_8_194_851_0, i_8_194_865_0, i_8_194_876_0,
    i_8_194_891_0, i_8_194_895_0, i_8_194_931_0, i_8_194_945_0,
    i_8_194_994_0, i_8_194_1101_0, i_8_194_1104_0, i_8_194_1115_0,
    i_8_194_1129_0, i_8_194_1240_0, i_8_194_1251_0, i_8_194_1256_0,
    i_8_194_1267_0, i_8_194_1268_0, i_8_194_1271_0, i_8_194_1291_0,
    i_8_194_1296_0, i_8_194_1329_0, i_8_194_1366_0, i_8_194_1378_0,
    i_8_194_1407_0, i_8_194_1435_0, i_8_194_1461_0, i_8_194_1465_0,
    i_8_194_1482_0, i_8_194_1544_0, i_8_194_1608_0, i_8_194_1620_0,
    i_8_194_1627_0, i_8_194_1651_0, i_8_194_1740_0, i_8_194_1747_0,
    i_8_194_1750_0, i_8_194_1760_0, i_8_194_1784_0, i_8_194_1787_0,
    i_8_194_1788_0, i_8_194_1789_0, i_8_194_1810_0, i_8_194_1840_0,
    i_8_194_1867_0, i_8_194_1899_0, i_8_194_1963_0, i_8_194_1966_0,
    i_8_194_1983_0, i_8_194_1984_0, i_8_194_1992_0, i_8_194_2068_0,
    i_8_194_2091_0, i_8_194_2104_0, i_8_194_2127_0, i_8_194_2158_0,
    i_8_194_2191_0, i_8_194_2216_0, i_8_194_2236_0, i_8_194_2240_0,
    i_8_194_2241_0, i_8_194_2246_0, i_8_194_2248_0,
    o_8_194_0_0  );
  input  i_8_194_21_0, i_8_194_42_0, i_8_194_52_0, i_8_194_55_0,
    i_8_194_58_0, i_8_194_89_0, i_8_194_120_0, i_8_194_129_0,
    i_8_194_183_0, i_8_194_184_0, i_8_194_211_0, i_8_194_218_0,
    i_8_194_241_0, i_8_194_262_0, i_8_194_319_0, i_8_194_365_0,
    i_8_194_369_0, i_8_194_427_0, i_8_194_456_0, i_8_194_478_0,
    i_8_194_535_0, i_8_194_543_0, i_8_194_549_0, i_8_194_551_0,
    i_8_194_593_0, i_8_194_611_0, i_8_194_612_0, i_8_194_613_0,
    i_8_194_634_0, i_8_194_643_0, i_8_194_656_0, i_8_194_662_0,
    i_8_194_665_0, i_8_194_730_0, i_8_194_787_0, i_8_194_802_0,
    i_8_194_804_0, i_8_194_832_0, i_8_194_851_0, i_8_194_865_0,
    i_8_194_876_0, i_8_194_891_0, i_8_194_895_0, i_8_194_931_0,
    i_8_194_945_0, i_8_194_994_0, i_8_194_1101_0, i_8_194_1104_0,
    i_8_194_1115_0, i_8_194_1129_0, i_8_194_1240_0, i_8_194_1251_0,
    i_8_194_1256_0, i_8_194_1267_0, i_8_194_1268_0, i_8_194_1271_0,
    i_8_194_1291_0, i_8_194_1296_0, i_8_194_1329_0, i_8_194_1366_0,
    i_8_194_1378_0, i_8_194_1407_0, i_8_194_1435_0, i_8_194_1461_0,
    i_8_194_1465_0, i_8_194_1482_0, i_8_194_1544_0, i_8_194_1608_0,
    i_8_194_1620_0, i_8_194_1627_0, i_8_194_1651_0, i_8_194_1740_0,
    i_8_194_1747_0, i_8_194_1750_0, i_8_194_1760_0, i_8_194_1784_0,
    i_8_194_1787_0, i_8_194_1788_0, i_8_194_1789_0, i_8_194_1810_0,
    i_8_194_1840_0, i_8_194_1867_0, i_8_194_1899_0, i_8_194_1963_0,
    i_8_194_1966_0, i_8_194_1983_0, i_8_194_1984_0, i_8_194_1992_0,
    i_8_194_2068_0, i_8_194_2091_0, i_8_194_2104_0, i_8_194_2127_0,
    i_8_194_2158_0, i_8_194_2191_0, i_8_194_2216_0, i_8_194_2236_0,
    i_8_194_2240_0, i_8_194_2241_0, i_8_194_2246_0, i_8_194_2248_0;
  output o_8_194_0_0;
  assign o_8_194_0_0 = 0;
endmodule



// Benchmark "kernel_8_195" written by ABC on Sun Jul 19 10:06:26 2020

module kernel_8_195 ( 
    i_8_195_21_0, i_8_195_79_0, i_8_195_129_0, i_8_195_138_0,
    i_8_195_192_0, i_8_195_195_0, i_8_195_228_0, i_8_195_256_0,
    i_8_195_345_0, i_8_195_347_0, i_8_195_349_0, i_8_195_354_0,
    i_8_195_362_0, i_8_195_368_0, i_8_195_382_0, i_8_195_428_0,
    i_8_195_477_0, i_8_195_525_0, i_8_195_529_0, i_8_195_552_0,
    i_8_195_555_0, i_8_195_567_0, i_8_195_570_0, i_8_195_651_0,
    i_8_195_654_0, i_8_195_662_0, i_8_195_675_0, i_8_195_688_0,
    i_8_195_696_0, i_8_195_703_0, i_8_195_705_0, i_8_195_729_0,
    i_8_195_732_0, i_8_195_750_0, i_8_195_751_0, i_8_195_774_0,
    i_8_195_775_0, i_8_195_789_0, i_8_195_801_0, i_8_195_832_0,
    i_8_195_859_0, i_8_195_885_0, i_8_195_886_0, i_8_195_969_0,
    i_8_195_984_0, i_8_195_1002_0, i_8_195_1038_0, i_8_195_1051_0,
    i_8_195_1101_0, i_8_195_1119_0, i_8_195_1130_0, i_8_195_1137_0,
    i_8_195_1146_0, i_8_195_1164_0, i_8_195_1191_0, i_8_195_1356_0,
    i_8_195_1371_0, i_8_195_1395_0, i_8_195_1405_0, i_8_195_1435_0,
    i_8_195_1507_0, i_8_195_1524_0, i_8_195_1546_0, i_8_195_1547_0,
    i_8_195_1597_0, i_8_195_1606_0, i_8_195_1610_0, i_8_195_1626_0,
    i_8_195_1632_0, i_8_195_1650_0, i_8_195_1659_0, i_8_195_1677_0,
    i_8_195_1683_0, i_8_195_1722_0, i_8_195_1728_0, i_8_195_1731_0,
    i_8_195_1767_0, i_8_195_1768_0, i_8_195_1779_0, i_8_195_1780_0,
    i_8_195_1825_0, i_8_195_1858_0, i_8_195_1888_0, i_8_195_1938_0,
    i_8_195_1947_0, i_8_195_1978_0, i_8_195_1992_0, i_8_195_2056_0,
    i_8_195_2073_0, i_8_195_2091_0, i_8_195_2092_0, i_8_195_2097_0,
    i_8_195_2100_0, i_8_195_2142_0, i_8_195_2146_0, i_8_195_2172_0,
    i_8_195_2215_0, i_8_195_2258_0, i_8_195_2284_0, i_8_195_2298_0,
    o_8_195_0_0  );
  input  i_8_195_21_0, i_8_195_79_0, i_8_195_129_0, i_8_195_138_0,
    i_8_195_192_0, i_8_195_195_0, i_8_195_228_0, i_8_195_256_0,
    i_8_195_345_0, i_8_195_347_0, i_8_195_349_0, i_8_195_354_0,
    i_8_195_362_0, i_8_195_368_0, i_8_195_382_0, i_8_195_428_0,
    i_8_195_477_0, i_8_195_525_0, i_8_195_529_0, i_8_195_552_0,
    i_8_195_555_0, i_8_195_567_0, i_8_195_570_0, i_8_195_651_0,
    i_8_195_654_0, i_8_195_662_0, i_8_195_675_0, i_8_195_688_0,
    i_8_195_696_0, i_8_195_703_0, i_8_195_705_0, i_8_195_729_0,
    i_8_195_732_0, i_8_195_750_0, i_8_195_751_0, i_8_195_774_0,
    i_8_195_775_0, i_8_195_789_0, i_8_195_801_0, i_8_195_832_0,
    i_8_195_859_0, i_8_195_885_0, i_8_195_886_0, i_8_195_969_0,
    i_8_195_984_0, i_8_195_1002_0, i_8_195_1038_0, i_8_195_1051_0,
    i_8_195_1101_0, i_8_195_1119_0, i_8_195_1130_0, i_8_195_1137_0,
    i_8_195_1146_0, i_8_195_1164_0, i_8_195_1191_0, i_8_195_1356_0,
    i_8_195_1371_0, i_8_195_1395_0, i_8_195_1405_0, i_8_195_1435_0,
    i_8_195_1507_0, i_8_195_1524_0, i_8_195_1546_0, i_8_195_1547_0,
    i_8_195_1597_0, i_8_195_1606_0, i_8_195_1610_0, i_8_195_1626_0,
    i_8_195_1632_0, i_8_195_1650_0, i_8_195_1659_0, i_8_195_1677_0,
    i_8_195_1683_0, i_8_195_1722_0, i_8_195_1728_0, i_8_195_1731_0,
    i_8_195_1767_0, i_8_195_1768_0, i_8_195_1779_0, i_8_195_1780_0,
    i_8_195_1825_0, i_8_195_1858_0, i_8_195_1888_0, i_8_195_1938_0,
    i_8_195_1947_0, i_8_195_1978_0, i_8_195_1992_0, i_8_195_2056_0,
    i_8_195_2073_0, i_8_195_2091_0, i_8_195_2092_0, i_8_195_2097_0,
    i_8_195_2100_0, i_8_195_2142_0, i_8_195_2146_0, i_8_195_2172_0,
    i_8_195_2215_0, i_8_195_2258_0, i_8_195_2284_0, i_8_195_2298_0;
  output o_8_195_0_0;
  assign o_8_195_0_0 = 0;
endmodule



// Benchmark "kernel_8_196" written by ABC on Sun Jul 19 10:06:27 2020

module kernel_8_196 ( 
    i_8_196_0_0, i_8_196_3_0, i_8_196_67_0, i_8_196_73_0, i_8_196_75_0,
    i_8_196_84_0, i_8_196_111_0, i_8_196_114_0, i_8_196_126_0,
    i_8_196_184_0, i_8_196_192_0, i_8_196_194_0, i_8_196_246_0,
    i_8_196_274_0, i_8_196_301_0, i_8_196_305_0, i_8_196_345_0,
    i_8_196_354_0, i_8_196_364_0, i_8_196_388_0, i_8_196_397_0,
    i_8_196_418_0, i_8_196_453_0, i_8_196_462_0, i_8_196_463_0,
    i_8_196_495_0, i_8_196_572_0, i_8_196_578_0, i_8_196_588_0,
    i_8_196_592_0, i_8_196_604_0, i_8_196_615_0, i_8_196_641_0,
    i_8_196_642_0, i_8_196_648_0, i_8_196_652_0, i_8_196_659_0,
    i_8_196_669_0, i_8_196_676_0, i_8_196_699_0, i_8_196_733_0,
    i_8_196_748_0, i_8_196_756_0, i_8_196_833_0, i_8_196_841_0,
    i_8_196_866_0, i_8_196_886_0, i_8_196_913_0, i_8_196_1107_0,
    i_8_196_1201_0, i_8_196_1219_0, i_8_196_1225_0, i_8_196_1226_0,
    i_8_196_1234_0, i_8_196_1240_0, i_8_196_1279_0, i_8_196_1315_0,
    i_8_196_1335_0, i_8_196_1336_0, i_8_196_1353_0, i_8_196_1355_0,
    i_8_196_1363_0, i_8_196_1366_0, i_8_196_1375_0, i_8_196_1389_0,
    i_8_196_1390_0, i_8_196_1436_0, i_8_196_1492_0, i_8_196_1494_0,
    i_8_196_1508_0, i_8_196_1509_0, i_8_196_1533_0, i_8_196_1606_0,
    i_8_196_1633_0, i_8_196_1638_0, i_8_196_1641_0, i_8_196_1682_0,
    i_8_196_1697_0, i_8_196_1703_0, i_8_196_1747_0, i_8_196_1765_0,
    i_8_196_1787_0, i_8_196_1819_0, i_8_196_1820_0, i_8_196_1843_0,
    i_8_196_1848_0, i_8_196_1863_0, i_8_196_1866_0, i_8_196_1881_0,
    i_8_196_1884_0, i_8_196_1918_0, i_8_196_1927_0, i_8_196_2064_0,
    i_8_196_2133_0, i_8_196_2224_0, i_8_196_2232_0, i_8_196_2242_0,
    i_8_196_2245_0, i_8_196_2246_0, i_8_196_2281_0,
    o_8_196_0_0  );
  input  i_8_196_0_0, i_8_196_3_0, i_8_196_67_0, i_8_196_73_0,
    i_8_196_75_0, i_8_196_84_0, i_8_196_111_0, i_8_196_114_0,
    i_8_196_126_0, i_8_196_184_0, i_8_196_192_0, i_8_196_194_0,
    i_8_196_246_0, i_8_196_274_0, i_8_196_301_0, i_8_196_305_0,
    i_8_196_345_0, i_8_196_354_0, i_8_196_364_0, i_8_196_388_0,
    i_8_196_397_0, i_8_196_418_0, i_8_196_453_0, i_8_196_462_0,
    i_8_196_463_0, i_8_196_495_0, i_8_196_572_0, i_8_196_578_0,
    i_8_196_588_0, i_8_196_592_0, i_8_196_604_0, i_8_196_615_0,
    i_8_196_641_0, i_8_196_642_0, i_8_196_648_0, i_8_196_652_0,
    i_8_196_659_0, i_8_196_669_0, i_8_196_676_0, i_8_196_699_0,
    i_8_196_733_0, i_8_196_748_0, i_8_196_756_0, i_8_196_833_0,
    i_8_196_841_0, i_8_196_866_0, i_8_196_886_0, i_8_196_913_0,
    i_8_196_1107_0, i_8_196_1201_0, i_8_196_1219_0, i_8_196_1225_0,
    i_8_196_1226_0, i_8_196_1234_0, i_8_196_1240_0, i_8_196_1279_0,
    i_8_196_1315_0, i_8_196_1335_0, i_8_196_1336_0, i_8_196_1353_0,
    i_8_196_1355_0, i_8_196_1363_0, i_8_196_1366_0, i_8_196_1375_0,
    i_8_196_1389_0, i_8_196_1390_0, i_8_196_1436_0, i_8_196_1492_0,
    i_8_196_1494_0, i_8_196_1508_0, i_8_196_1509_0, i_8_196_1533_0,
    i_8_196_1606_0, i_8_196_1633_0, i_8_196_1638_0, i_8_196_1641_0,
    i_8_196_1682_0, i_8_196_1697_0, i_8_196_1703_0, i_8_196_1747_0,
    i_8_196_1765_0, i_8_196_1787_0, i_8_196_1819_0, i_8_196_1820_0,
    i_8_196_1843_0, i_8_196_1848_0, i_8_196_1863_0, i_8_196_1866_0,
    i_8_196_1881_0, i_8_196_1884_0, i_8_196_1918_0, i_8_196_1927_0,
    i_8_196_2064_0, i_8_196_2133_0, i_8_196_2224_0, i_8_196_2232_0,
    i_8_196_2242_0, i_8_196_2245_0, i_8_196_2246_0, i_8_196_2281_0;
  output o_8_196_0_0;
  assign o_8_196_0_0 = 0;
endmodule



// Benchmark "kernel_8_197" written by ABC on Sun Jul 19 10:06:28 2020

module kernel_8_197 ( 
    i_8_197_66_0, i_8_197_75_0, i_8_197_88_0, i_8_197_114_0, i_8_197_148_0,
    i_8_197_165_0, i_8_197_174_0, i_8_197_193_0, i_8_197_202_0,
    i_8_197_228_0, i_8_197_300_0, i_8_197_312_0, i_8_197_336_0,
    i_8_197_349_0, i_8_197_354_0, i_8_197_366_0, i_8_197_418_0,
    i_8_197_426_0, i_8_197_429_0, i_8_197_453_0, i_8_197_489_0,
    i_8_197_508_0, i_8_197_522_0, i_8_197_535_0, i_8_197_574_0,
    i_8_197_582_0, i_8_197_606_0, i_8_197_608_0, i_8_197_615_0,
    i_8_197_657_0, i_8_197_665_0, i_8_197_700_0, i_8_197_701_0,
    i_8_197_705_0, i_8_197_730_0, i_8_197_759_0, i_8_197_772_0,
    i_8_197_835_0, i_8_197_840_0, i_8_197_841_0, i_8_197_858_0,
    i_8_197_865_0, i_8_197_870_0, i_8_197_912_0, i_8_197_921_0,
    i_8_197_969_0, i_8_197_1029_0, i_8_197_1034_0, i_8_197_1038_0,
    i_8_197_1068_0, i_8_197_1114_0, i_8_197_1123_0, i_8_197_1132_0,
    i_8_197_1134_0, i_8_197_1227_0, i_8_197_1232_0, i_8_197_1281_0,
    i_8_197_1305_0, i_8_197_1323_0, i_8_197_1372_0, i_8_197_1398_0,
    i_8_197_1470_0, i_8_197_1548_0, i_8_197_1571_0, i_8_197_1587_0,
    i_8_197_1623_0, i_8_197_1633_0, i_8_197_1686_0, i_8_197_1696_0,
    i_8_197_1699_0, i_8_197_1767_0, i_8_197_1773_0, i_8_197_1790_0,
    i_8_197_1794_0, i_8_197_1806_0, i_8_197_1822_0, i_8_197_1824_0,
    i_8_197_1840_0, i_8_197_1869_0, i_8_197_1929_0, i_8_197_1938_0,
    i_8_197_2004_0, i_8_197_2008_0, i_8_197_2010_0, i_8_197_2019_0,
    i_8_197_2073_0, i_8_197_2103_0, i_8_197_2109_0, i_8_197_2134_0,
    i_8_197_2144_0, i_8_197_2145_0, i_8_197_2147_0, i_8_197_2154_0,
    i_8_197_2158_0, i_8_197_2225_0, i_8_197_2226_0, i_8_197_2227_0,
    i_8_197_2229_0, i_8_197_2271_0, i_8_197_2281_0,
    o_8_197_0_0  );
  input  i_8_197_66_0, i_8_197_75_0, i_8_197_88_0, i_8_197_114_0,
    i_8_197_148_0, i_8_197_165_0, i_8_197_174_0, i_8_197_193_0,
    i_8_197_202_0, i_8_197_228_0, i_8_197_300_0, i_8_197_312_0,
    i_8_197_336_0, i_8_197_349_0, i_8_197_354_0, i_8_197_366_0,
    i_8_197_418_0, i_8_197_426_0, i_8_197_429_0, i_8_197_453_0,
    i_8_197_489_0, i_8_197_508_0, i_8_197_522_0, i_8_197_535_0,
    i_8_197_574_0, i_8_197_582_0, i_8_197_606_0, i_8_197_608_0,
    i_8_197_615_0, i_8_197_657_0, i_8_197_665_0, i_8_197_700_0,
    i_8_197_701_0, i_8_197_705_0, i_8_197_730_0, i_8_197_759_0,
    i_8_197_772_0, i_8_197_835_0, i_8_197_840_0, i_8_197_841_0,
    i_8_197_858_0, i_8_197_865_0, i_8_197_870_0, i_8_197_912_0,
    i_8_197_921_0, i_8_197_969_0, i_8_197_1029_0, i_8_197_1034_0,
    i_8_197_1038_0, i_8_197_1068_0, i_8_197_1114_0, i_8_197_1123_0,
    i_8_197_1132_0, i_8_197_1134_0, i_8_197_1227_0, i_8_197_1232_0,
    i_8_197_1281_0, i_8_197_1305_0, i_8_197_1323_0, i_8_197_1372_0,
    i_8_197_1398_0, i_8_197_1470_0, i_8_197_1548_0, i_8_197_1571_0,
    i_8_197_1587_0, i_8_197_1623_0, i_8_197_1633_0, i_8_197_1686_0,
    i_8_197_1696_0, i_8_197_1699_0, i_8_197_1767_0, i_8_197_1773_0,
    i_8_197_1790_0, i_8_197_1794_0, i_8_197_1806_0, i_8_197_1822_0,
    i_8_197_1824_0, i_8_197_1840_0, i_8_197_1869_0, i_8_197_1929_0,
    i_8_197_1938_0, i_8_197_2004_0, i_8_197_2008_0, i_8_197_2010_0,
    i_8_197_2019_0, i_8_197_2073_0, i_8_197_2103_0, i_8_197_2109_0,
    i_8_197_2134_0, i_8_197_2144_0, i_8_197_2145_0, i_8_197_2147_0,
    i_8_197_2154_0, i_8_197_2158_0, i_8_197_2225_0, i_8_197_2226_0,
    i_8_197_2227_0, i_8_197_2229_0, i_8_197_2271_0, i_8_197_2281_0;
  output o_8_197_0_0;
  assign o_8_197_0_0 = 0;
endmodule



// Benchmark "kernel_8_198" written by ABC on Sun Jul 19 10:06:28 2020

module kernel_8_198 ( 
    i_8_198_58_0, i_8_198_73_0, i_8_198_76_0, i_8_198_77_0, i_8_198_115_0,
    i_8_198_116_0, i_8_198_137_0, i_8_198_140_0, i_8_198_181_0,
    i_8_198_184_0, i_8_198_221_0, i_8_198_231_0, i_8_198_256_0,
    i_8_198_301_0, i_8_198_320_0, i_8_198_389_0, i_8_198_419_0,
    i_8_198_431_0, i_8_198_482_0, i_8_198_496_0, i_8_198_509_0,
    i_8_198_524_0, i_8_198_526_0, i_8_198_527_0, i_8_198_572_0,
    i_8_198_590_0, i_8_198_608_0, i_8_198_611_0, i_8_198_655_0,
    i_8_198_658_0, i_8_198_694_0, i_8_198_696_0, i_8_198_737_0,
    i_8_198_760_0, i_8_198_761_0, i_8_198_776_0, i_8_198_824_0,
    i_8_198_837_0, i_8_198_838_0, i_8_198_850_0, i_8_198_928_0,
    i_8_198_1010_0, i_8_198_1100_0, i_8_198_1103_0, i_8_198_1129_0,
    i_8_198_1130_0, i_8_198_1229_0, i_8_198_1247_0, i_8_198_1268_0,
    i_8_198_1279_0, i_8_198_1295_0, i_8_198_1316_0, i_8_198_1319_0,
    i_8_198_1327_0, i_8_198_1334_0, i_8_198_1397_0, i_8_198_1423_0,
    i_8_198_1424_0, i_8_198_1442_0, i_8_198_1462_0, i_8_198_1463_0,
    i_8_198_1472_0, i_8_198_1478_0, i_8_198_1481_0, i_8_198_1493_0,
    i_8_198_1511_0, i_8_198_1514_0, i_8_198_1525_0, i_8_198_1526_0,
    i_8_198_1549_0, i_8_198_1550_0, i_8_198_1551_0, i_8_198_1559_0,
    i_8_198_1640_0, i_8_198_1643_0, i_8_198_1675_0, i_8_198_1676_0,
    i_8_198_1679_0, i_8_198_1684_0, i_8_198_1697_0, i_8_198_1700_0,
    i_8_198_1706_0, i_8_198_1721_0, i_8_198_1747_0, i_8_198_1780_0,
    i_8_198_1781_0, i_8_198_1787_0, i_8_198_1793_0, i_8_198_1810_0,
    i_8_198_1838_0, i_8_198_1840_0, i_8_198_1841_0, i_8_198_1885_0,
    i_8_198_1937_0, i_8_198_1949_0, i_8_198_1954_0, i_8_198_1968_0,
    i_8_198_2075_0, i_8_198_2135_0, i_8_198_2297_0,
    o_8_198_0_0  );
  input  i_8_198_58_0, i_8_198_73_0, i_8_198_76_0, i_8_198_77_0,
    i_8_198_115_0, i_8_198_116_0, i_8_198_137_0, i_8_198_140_0,
    i_8_198_181_0, i_8_198_184_0, i_8_198_221_0, i_8_198_231_0,
    i_8_198_256_0, i_8_198_301_0, i_8_198_320_0, i_8_198_389_0,
    i_8_198_419_0, i_8_198_431_0, i_8_198_482_0, i_8_198_496_0,
    i_8_198_509_0, i_8_198_524_0, i_8_198_526_0, i_8_198_527_0,
    i_8_198_572_0, i_8_198_590_0, i_8_198_608_0, i_8_198_611_0,
    i_8_198_655_0, i_8_198_658_0, i_8_198_694_0, i_8_198_696_0,
    i_8_198_737_0, i_8_198_760_0, i_8_198_761_0, i_8_198_776_0,
    i_8_198_824_0, i_8_198_837_0, i_8_198_838_0, i_8_198_850_0,
    i_8_198_928_0, i_8_198_1010_0, i_8_198_1100_0, i_8_198_1103_0,
    i_8_198_1129_0, i_8_198_1130_0, i_8_198_1229_0, i_8_198_1247_0,
    i_8_198_1268_0, i_8_198_1279_0, i_8_198_1295_0, i_8_198_1316_0,
    i_8_198_1319_0, i_8_198_1327_0, i_8_198_1334_0, i_8_198_1397_0,
    i_8_198_1423_0, i_8_198_1424_0, i_8_198_1442_0, i_8_198_1462_0,
    i_8_198_1463_0, i_8_198_1472_0, i_8_198_1478_0, i_8_198_1481_0,
    i_8_198_1493_0, i_8_198_1511_0, i_8_198_1514_0, i_8_198_1525_0,
    i_8_198_1526_0, i_8_198_1549_0, i_8_198_1550_0, i_8_198_1551_0,
    i_8_198_1559_0, i_8_198_1640_0, i_8_198_1643_0, i_8_198_1675_0,
    i_8_198_1676_0, i_8_198_1679_0, i_8_198_1684_0, i_8_198_1697_0,
    i_8_198_1700_0, i_8_198_1706_0, i_8_198_1721_0, i_8_198_1747_0,
    i_8_198_1780_0, i_8_198_1781_0, i_8_198_1787_0, i_8_198_1793_0,
    i_8_198_1810_0, i_8_198_1838_0, i_8_198_1840_0, i_8_198_1841_0,
    i_8_198_1885_0, i_8_198_1937_0, i_8_198_1949_0, i_8_198_1954_0,
    i_8_198_1968_0, i_8_198_2075_0, i_8_198_2135_0, i_8_198_2297_0;
  output o_8_198_0_0;
  assign o_8_198_0_0 = 0;
endmodule



// Benchmark "kernel_8_199" written by ABC on Sun Jul 19 10:06:30 2020

module kernel_8_199 ( 
    i_8_199_1_0, i_8_199_49_0, i_8_199_76_0, i_8_199_86_0, i_8_199_118_0,
    i_8_199_119_0, i_8_199_164_0, i_8_199_167_0, i_8_199_226_0,
    i_8_199_244_0, i_8_199_300_0, i_8_199_326_0, i_8_199_350_0,
    i_8_199_425_0, i_8_199_452_0, i_8_199_464_0, i_8_199_487_0,
    i_8_199_490_0, i_8_199_496_0, i_8_199_497_0, i_8_199_500_0,
    i_8_199_530_0, i_8_199_556_0, i_8_199_589_0, i_8_199_605_0,
    i_8_199_653_0, i_8_199_695_0, i_8_199_698_0, i_8_199_707_0,
    i_8_199_823_0, i_8_199_824_0, i_8_199_838_0, i_8_199_839_0,
    i_8_199_841_0, i_8_199_875_0, i_8_199_884_0, i_8_199_929_0,
    i_8_199_968_0, i_8_199_992_0, i_8_199_1001_0, i_8_199_1036_0,
    i_8_199_1037_0, i_8_199_1046_0, i_8_199_1052_0, i_8_199_1072_0,
    i_8_199_1075_0, i_8_199_1076_0, i_8_199_1163_0, i_8_199_1166_0,
    i_8_199_1226_0, i_8_199_1233_0, i_8_199_1270_0, i_8_199_1274_0,
    i_8_199_1280_0, i_8_199_1281_0, i_8_199_1282_0, i_8_199_1298_0,
    i_8_199_1318_0, i_8_199_1321_0, i_8_199_1327_0, i_8_199_1408_0,
    i_8_199_1432_0, i_8_199_1435_0, i_8_199_1436_0, i_8_199_1467_0,
    i_8_199_1468_0, i_8_199_1478_0, i_8_199_1496_0, i_8_199_1534_0,
    i_8_199_1543_0, i_8_199_1544_0, i_8_199_1657_0, i_8_199_1703_0,
    i_8_199_1733_0, i_8_199_1749_0, i_8_199_1751_0, i_8_199_1754_0,
    i_8_199_1760_0, i_8_199_1766_0, i_8_199_1769_0, i_8_199_1777_0,
    i_8_199_1811_0, i_8_199_1822_0, i_8_199_1850_0, i_8_199_1868_0,
    i_8_199_1974_0, i_8_199_1976_0, i_8_199_1982_0, i_8_199_1993_0,
    i_8_199_1994_0, i_8_199_2057_0, i_8_199_2102_0, i_8_199_2125_0,
    i_8_199_2135_0, i_8_199_2143_0, i_8_199_2153_0, i_8_199_2223_0,
    i_8_199_2225_0, i_8_199_2269_0, i_8_199_2273_0,
    o_8_199_0_0  );
  input  i_8_199_1_0, i_8_199_49_0, i_8_199_76_0, i_8_199_86_0,
    i_8_199_118_0, i_8_199_119_0, i_8_199_164_0, i_8_199_167_0,
    i_8_199_226_0, i_8_199_244_0, i_8_199_300_0, i_8_199_326_0,
    i_8_199_350_0, i_8_199_425_0, i_8_199_452_0, i_8_199_464_0,
    i_8_199_487_0, i_8_199_490_0, i_8_199_496_0, i_8_199_497_0,
    i_8_199_500_0, i_8_199_530_0, i_8_199_556_0, i_8_199_589_0,
    i_8_199_605_0, i_8_199_653_0, i_8_199_695_0, i_8_199_698_0,
    i_8_199_707_0, i_8_199_823_0, i_8_199_824_0, i_8_199_838_0,
    i_8_199_839_0, i_8_199_841_0, i_8_199_875_0, i_8_199_884_0,
    i_8_199_929_0, i_8_199_968_0, i_8_199_992_0, i_8_199_1001_0,
    i_8_199_1036_0, i_8_199_1037_0, i_8_199_1046_0, i_8_199_1052_0,
    i_8_199_1072_0, i_8_199_1075_0, i_8_199_1076_0, i_8_199_1163_0,
    i_8_199_1166_0, i_8_199_1226_0, i_8_199_1233_0, i_8_199_1270_0,
    i_8_199_1274_0, i_8_199_1280_0, i_8_199_1281_0, i_8_199_1282_0,
    i_8_199_1298_0, i_8_199_1318_0, i_8_199_1321_0, i_8_199_1327_0,
    i_8_199_1408_0, i_8_199_1432_0, i_8_199_1435_0, i_8_199_1436_0,
    i_8_199_1467_0, i_8_199_1468_0, i_8_199_1478_0, i_8_199_1496_0,
    i_8_199_1534_0, i_8_199_1543_0, i_8_199_1544_0, i_8_199_1657_0,
    i_8_199_1703_0, i_8_199_1733_0, i_8_199_1749_0, i_8_199_1751_0,
    i_8_199_1754_0, i_8_199_1760_0, i_8_199_1766_0, i_8_199_1769_0,
    i_8_199_1777_0, i_8_199_1811_0, i_8_199_1822_0, i_8_199_1850_0,
    i_8_199_1868_0, i_8_199_1974_0, i_8_199_1976_0, i_8_199_1982_0,
    i_8_199_1993_0, i_8_199_1994_0, i_8_199_2057_0, i_8_199_2102_0,
    i_8_199_2125_0, i_8_199_2135_0, i_8_199_2143_0, i_8_199_2153_0,
    i_8_199_2223_0, i_8_199_2225_0, i_8_199_2269_0, i_8_199_2273_0;
  output o_8_199_0_0;
  assign o_8_199_0_0 = ~((~i_8_199_1_0 & ((~i_8_199_49_0 & ~i_8_199_118_0 & ~i_8_199_556_0 & ~i_8_199_1166_0 & i_8_199_1226_0 & ~i_8_199_1544_0 & ~i_8_199_1733_0 & ~i_8_199_1769_0) | (~i_8_199_326_0 & ~i_8_199_530_0 & ~i_8_199_838_0 & ~i_8_199_1052_0 & ~i_8_199_1754_0 & i_8_199_1777_0 & ~i_8_199_2125_0))) | (i_8_199_452_0 & ((i_8_199_164_0 & ~i_8_199_707_0 & i_8_199_968_0 & ~i_8_199_1318_0) | (~i_8_199_490_0 & ~i_8_199_556_0 & ~i_8_199_823_0 & ~i_8_199_929_0 & ~i_8_199_1037_0 & ~i_8_199_1163_0 & ~i_8_199_1657_0 & ~i_8_199_2143_0))) | (~i_8_199_1046_0 & ((~i_8_199_496_0 & ((~i_8_199_487_0 & ~i_8_199_875_0 & ~i_8_199_1282_0 & ~i_8_199_1534_0 & ~i_8_199_1733_0 & i_8_199_1822_0) | (~i_8_199_76_0 & i_8_199_300_0 & ~i_8_199_589_0 & ~i_8_199_1036_0 & ~i_8_199_1318_0 & ~i_8_199_1822_0))) | (i_8_199_589_0 & ~i_8_199_605_0 & i_8_199_823_0 & ~i_8_199_1036_0 & ~i_8_199_1657_0) | (~i_8_199_1001_0 & i_8_199_1327_0 & ~i_8_199_1760_0))) | (~i_8_199_530_0 & ((~i_8_199_1001_0 & i_8_199_1534_0 & ~i_8_199_1543_0 & ~i_8_199_2102_0 & ~i_8_199_2125_0) | (~i_8_199_487_0 & i_8_199_605_0 & ~i_8_199_1072_0 & i_8_199_1281_0 & i_8_199_1432_0 & ~i_8_199_2269_0))) | (~i_8_199_487_0 & ((~i_8_199_653_0 & i_8_199_841_0 & i_8_199_1408_0 & ~i_8_199_1543_0) | (~i_8_199_425_0 & ~i_8_199_1769_0 & i_8_199_1777_0 & ~i_8_199_1993_0))) | (~i_8_199_425_0 & ((i_8_199_698_0 & ~i_8_199_875_0 & ~i_8_199_1036_0 & ~i_8_199_1037_0 & ~i_8_199_1166_0 & ~i_8_199_1233_0 & ~i_8_199_1281_0 & ~i_8_199_1543_0) | (~i_8_199_838_0 & ~i_8_199_968_0 & ~i_8_199_1993_0 & ~i_8_199_2057_0))) | (i_8_199_556_0 & ((~i_8_199_707_0 & ~i_8_199_1543_0) | (i_8_199_1657_0 & ~i_8_199_1822_0))) | (i_8_199_589_0 & ((~i_8_199_226_0 & ~i_8_199_300_0 & ~i_8_199_1233_0 & i_8_199_1282_0 & ~i_8_199_1408_0 & i_8_199_1544_0 & ~i_8_199_1703_0) | (~i_8_199_490_0 & ~i_8_199_497_0 & ~i_8_199_605_0 & i_8_199_1435_0 & ~i_8_199_1657_0 & ~i_8_199_2102_0))) | (~i_8_199_695_0 & ((~i_8_199_167_0 & ~i_8_199_452_0 & ~i_8_199_838_0 & ~i_8_199_992_0 & ~i_8_199_1037_0 & ~i_8_199_1166_0 & ~i_8_199_1226_0 & ~i_8_199_1543_0 & ~i_8_199_2135_0) | (~i_8_199_226_0 & ~i_8_199_1036_0 & i_8_199_1281_0 & ~i_8_199_1749_0 & ~i_8_199_1769_0 & ~i_8_199_1822_0 & ~i_8_199_2223_0 & ~i_8_199_2225_0))) | (~i_8_199_2143_0 & ((~i_8_199_838_0 & ((~i_8_199_118_0 & ~i_8_199_824_0 & ~i_8_199_1037_0 & ~i_8_199_1318_0 & ~i_8_199_1544_0 & i_8_199_2102_0) | (~i_8_199_326_0 & ~i_8_199_589_0 & ~i_8_199_839_0 & ~i_8_199_1993_0 & ~i_8_199_2273_0))) | (i_8_199_76_0 & ~i_8_199_653_0 & ~i_8_199_1408_0))) | (i_8_199_76_0 & ((~i_8_199_556_0 & ~i_8_199_653_0 & ~i_8_199_1281_0 & ~i_8_199_1749_0 & ~i_8_199_1822_0) | (~i_8_199_350_0 & ~i_8_199_490_0 & ~i_8_199_1037_0 & i_8_199_1436_0 & ~i_8_199_2125_0))) | (~i_8_199_326_0 & ((~i_8_199_992_0 & i_8_199_1233_0 & ~i_8_199_1496_0 & ~i_8_199_1543_0) | (i_8_199_500_0 & ~i_8_199_1544_0))) | (~i_8_199_490_0 & ((~i_8_199_119_0 & ~i_8_199_841_0 & ~i_8_199_1163_0 & ~i_8_199_1769_0 & ~i_8_199_2135_0) | (~i_8_199_653_0 & ~i_8_199_839_0 & ~i_8_199_968_0 & ~i_8_199_1543_0 & ~i_8_199_1777_0 & ~i_8_199_2269_0))) | (~i_8_199_119_0 & ((i_8_199_707_0 & ~i_8_199_992_0 & ~i_8_199_1163_0 & i_8_199_1282_0 & ~i_8_199_1327_0 & ~i_8_199_1543_0 & ~i_8_199_1766_0) | (i_8_199_49_0 & i_8_199_490_0 & ~i_8_199_653_0 & i_8_199_1822_0))) | (~i_8_199_653_0 & ((~i_8_199_884_0 & i_8_199_1075_0 & ~i_8_199_1822_0) | (~i_8_199_226_0 & ~i_8_199_875_0 & ~i_8_199_1327_0 & ~i_8_199_1408_0 & ~i_8_199_1478_0 & ~i_8_199_1543_0 & ~i_8_199_1703_0 & ~i_8_199_2135_0 & ~i_8_199_2273_0))) | (~i_8_199_226_0 & ((~i_8_199_589_0 & ~i_8_199_1163_0 & i_8_199_1280_0 & ~i_8_199_1432_0 & ~i_8_199_1534_0 & ~i_8_199_1544_0 & ~i_8_199_1769_0) | (~i_8_199_1166_0 & i_8_199_1436_0 & i_8_199_1751_0 & ~i_8_199_1850_0 & ~i_8_199_2057_0))) | (~i_8_199_875_0 & ~i_8_199_1435_0 & ((~i_8_199_698_0 & i_8_199_1036_0 & ~i_8_199_1281_0 & i_8_199_1432_0) | (~i_8_199_929_0 & ~i_8_199_992_0 & ~i_8_199_1052_0 & ~i_8_199_1468_0 & ~i_8_199_1496_0 & ~i_8_199_1543_0 & ~i_8_199_1544_0 & i_8_199_1822_0 & ~i_8_199_2269_0))) | (~i_8_199_698_0 & ((i_8_199_1754_0 & ~i_8_199_1982_0 & ~i_8_199_2057_0) | (~i_8_199_1777_0 & ~i_8_199_1994_0 & ~i_8_199_2125_0 & i_8_199_2269_0))) | (i_8_199_1233_0 & ((~i_8_199_884_0 & ~i_8_199_1163_0 & ~i_8_199_1657_0 & ~i_8_199_1777_0) | (i_8_199_1281_0 & ~i_8_199_2135_0))) | (i_8_199_1467_0 & ((~i_8_199_968_0 & ~i_8_199_1543_0) | (~i_8_199_1432_0 & ~i_8_199_1657_0))) | (~i_8_199_1543_0 & ((~i_8_199_1327_0 & i_8_199_1435_0 & ~i_8_199_1544_0 & ~i_8_199_1994_0) | (~i_8_199_839_0 & i_8_199_1318_0 & ~i_8_199_2273_0))) | (i_8_199_1777_0 & ((~i_8_199_707_0 & i_8_199_1321_0 & ~i_8_199_1822_0) | (~i_8_199_589_0 & ~i_8_199_1166_0 & ~i_8_199_1281_0 & ~i_8_199_1408_0 & ~i_8_199_1993_0))) | (~i_8_199_589_0 & ((i_8_199_1468_0 & ~i_8_199_1534_0 & ~i_8_199_1766_0) | (i_8_199_1408_0 & ~i_8_199_1467_0 & i_8_199_1749_0 & ~i_8_199_1993_0 & ~i_8_199_2225_0))) | (i_8_199_226_0 & ~i_8_199_1544_0 & i_8_199_1657_0 & ~i_8_199_2125_0));
endmodule



// Benchmark "kernel_8_200" written by ABC on Sun Jul 19 10:06:32 2020

module kernel_8_200 ( 
    i_8_200_25_0, i_8_200_50_0, i_8_200_53_0, i_8_200_111_0, i_8_200_114_0,
    i_8_200_115_0, i_8_200_116_0, i_8_200_123_0, i_8_200_124_0,
    i_8_200_175_0, i_8_200_179_0, i_8_200_219_0, i_8_200_220_0,
    i_8_200_221_0, i_8_200_224_0, i_8_200_257_0, i_8_200_383_0,
    i_8_200_453_0, i_8_200_455_0, i_8_200_457_0, i_8_200_458_0,
    i_8_200_523_0, i_8_200_571_0, i_8_200_572_0, i_8_200_575_0,
    i_8_200_601_0, i_8_200_602_0, i_8_200_607_0, i_8_200_657_0,
    i_8_200_658_0, i_8_200_689_0, i_8_200_702_0, i_8_200_703_0,
    i_8_200_704_0, i_8_200_768_0, i_8_200_775_0, i_8_200_776_0,
    i_8_200_798_0, i_8_200_883_0, i_8_200_887_0, i_8_200_888_0,
    i_8_200_932_0, i_8_200_959_0, i_8_200_961_0, i_8_200_966_0,
    i_8_200_1072_0, i_8_200_1167_0, i_8_200_1178_0, i_8_200_1179_0,
    i_8_200_1180_0, i_8_200_1227_0, i_8_200_1228_0, i_8_200_1229_0,
    i_8_200_1262_0, i_8_200_1263_0, i_8_200_1278_0, i_8_200_1296_0,
    i_8_200_1470_0, i_8_200_1474_0, i_8_200_1487_0, i_8_200_1490_0,
    i_8_200_1560_0, i_8_200_1563_0, i_8_200_1564_0, i_8_200_1584_0,
    i_8_200_1585_0, i_8_200_1587_0, i_8_200_1588_0, i_8_200_1623_0,
    i_8_200_1632_0, i_8_200_1683_0, i_8_200_1695_0, i_8_200_1696_0,
    i_8_200_1699_0, i_8_200_1700_0, i_8_200_1738_0, i_8_200_1746_0,
    i_8_200_1758_0, i_8_200_1770_0, i_8_200_1772_0, i_8_200_1787_0,
    i_8_200_1789_0, i_8_200_1818_0, i_8_200_1820_0, i_8_200_1821_0,
    i_8_200_1854_0, i_8_200_1857_0, i_8_200_1969_0, i_8_200_2009_0,
    i_8_200_2073_0, i_8_200_2129_0, i_8_200_2222_0, i_8_200_2224_0,
    i_8_200_2226_0, i_8_200_2237_0, i_8_200_2247_0, i_8_200_2248_0,
    i_8_200_2249_0, i_8_200_2261_0, i_8_200_2293_0,
    o_8_200_0_0  );
  input  i_8_200_25_0, i_8_200_50_0, i_8_200_53_0, i_8_200_111_0,
    i_8_200_114_0, i_8_200_115_0, i_8_200_116_0, i_8_200_123_0,
    i_8_200_124_0, i_8_200_175_0, i_8_200_179_0, i_8_200_219_0,
    i_8_200_220_0, i_8_200_221_0, i_8_200_224_0, i_8_200_257_0,
    i_8_200_383_0, i_8_200_453_0, i_8_200_455_0, i_8_200_457_0,
    i_8_200_458_0, i_8_200_523_0, i_8_200_571_0, i_8_200_572_0,
    i_8_200_575_0, i_8_200_601_0, i_8_200_602_0, i_8_200_607_0,
    i_8_200_657_0, i_8_200_658_0, i_8_200_689_0, i_8_200_702_0,
    i_8_200_703_0, i_8_200_704_0, i_8_200_768_0, i_8_200_775_0,
    i_8_200_776_0, i_8_200_798_0, i_8_200_883_0, i_8_200_887_0,
    i_8_200_888_0, i_8_200_932_0, i_8_200_959_0, i_8_200_961_0,
    i_8_200_966_0, i_8_200_1072_0, i_8_200_1167_0, i_8_200_1178_0,
    i_8_200_1179_0, i_8_200_1180_0, i_8_200_1227_0, i_8_200_1228_0,
    i_8_200_1229_0, i_8_200_1262_0, i_8_200_1263_0, i_8_200_1278_0,
    i_8_200_1296_0, i_8_200_1470_0, i_8_200_1474_0, i_8_200_1487_0,
    i_8_200_1490_0, i_8_200_1560_0, i_8_200_1563_0, i_8_200_1564_0,
    i_8_200_1584_0, i_8_200_1585_0, i_8_200_1587_0, i_8_200_1588_0,
    i_8_200_1623_0, i_8_200_1632_0, i_8_200_1683_0, i_8_200_1695_0,
    i_8_200_1696_0, i_8_200_1699_0, i_8_200_1700_0, i_8_200_1738_0,
    i_8_200_1746_0, i_8_200_1758_0, i_8_200_1770_0, i_8_200_1772_0,
    i_8_200_1787_0, i_8_200_1789_0, i_8_200_1818_0, i_8_200_1820_0,
    i_8_200_1821_0, i_8_200_1854_0, i_8_200_1857_0, i_8_200_1969_0,
    i_8_200_2009_0, i_8_200_2073_0, i_8_200_2129_0, i_8_200_2222_0,
    i_8_200_2224_0, i_8_200_2226_0, i_8_200_2237_0, i_8_200_2247_0,
    i_8_200_2248_0, i_8_200_2249_0, i_8_200_2261_0, i_8_200_2293_0;
  output o_8_200_0_0;
  assign o_8_200_0_0 = ~((i_8_200_50_0 & ((i_8_200_115_0 & ~i_8_200_575_0 & ~i_8_200_888_0 & ~i_8_200_1585_0 & ~i_8_200_1696_0 & ~i_8_200_1789_0) | (~i_8_200_887_0 & ~i_8_200_1179_0 & ~i_8_200_1487_0 & ~i_8_200_1587_0 & ~i_8_200_1588_0 & ~i_8_200_1632_0 & ~i_8_200_1695_0 & i_8_200_1787_0 & ~i_8_200_2073_0))) | (~i_8_200_219_0 & ((~i_8_200_575_0 & ~i_8_200_887_0 & ~i_8_200_1263_0 & ~i_8_200_1560_0 & i_8_200_1564_0 & ~i_8_200_1632_0 & ~i_8_200_1683_0 & ~i_8_200_1818_0 & ~i_8_200_1854_0) | (~i_8_200_224_0 & i_8_200_961_0 & ~i_8_200_966_0 & ~i_8_200_1585_0 & ~i_8_200_1699_0 & ~i_8_200_1857_0 & ~i_8_200_2129_0))) | (~i_8_200_123_0 & ((~i_8_200_1585_0 & ((~i_8_200_776_0 & ~i_8_200_1695_0 & ((~i_8_200_114_0 & ((i_8_200_219_0 & ~i_8_200_575_0 & ~i_8_200_1587_0 & ~i_8_200_1699_0 & ~i_8_200_1854_0 & ~i_8_200_1857_0) | (~i_8_200_116_0 & ~i_8_200_224_0 & ~i_8_200_1584_0 & ~i_8_200_1588_0 & ~i_8_200_1818_0 & ~i_8_200_2129_0 & ~i_8_200_2222_0 & ~i_8_200_2247_0))) | (~i_8_200_224_0 & ~i_8_200_1262_0 & i_8_200_1263_0 & ~i_8_200_1490_0 & ~i_8_200_1584_0 & ~i_8_200_1587_0 & ~i_8_200_1738_0 & ~i_8_200_2248_0))) | (~i_8_200_1587_0 & ((~i_8_200_220_0 & ~i_8_200_571_0 & ~i_8_200_888_0 & ~i_8_200_1167_0 & i_8_200_1623_0 & ~i_8_200_1758_0 & ~i_8_200_1770_0) | (~i_8_200_1179_0 & ~i_8_200_1227_0 & ~i_8_200_1262_0 & i_8_200_1263_0 & ~i_8_200_1490_0 & ~i_8_200_1623_0 & ~i_8_200_1746_0 & ~i_8_200_1772_0 & ~i_8_200_1787_0 & ~i_8_200_1789_0))))) | (~i_8_200_1738_0 & ((~i_8_200_116_0 & ((i_8_200_798_0 & i_8_200_1470_0 & ~i_8_200_2248_0) | (i_8_200_224_0 & ~i_8_200_798_0 & ~i_8_200_1180_0 & ~i_8_200_1584_0 & ~i_8_200_1695_0 & ~i_8_200_1772_0 & ~i_8_200_2009_0 & ~i_8_200_2293_0))) | (~i_8_200_111_0 & ~i_8_200_220_0 & ~i_8_200_257_0 & ~i_8_200_383_0 & ~i_8_200_455_0 & ~i_8_200_575_0 & i_8_200_1262_0 & ~i_8_200_1700_0 & ~i_8_200_2129_0 & ~i_8_200_2224_0))) | (~i_8_200_1584_0 & ((~i_8_200_1588_0 & ((~i_8_200_115_0 & ~i_8_200_966_0 & ~i_8_200_1758_0 & i_8_200_1770_0 & ~i_8_200_2073_0 & ~i_8_200_2129_0) | (~i_8_200_575_0 & ~i_8_200_1167_0 & ~i_8_200_1490_0 & ~i_8_200_1623_0 & i_8_200_1758_0 & ~i_8_200_1857_0 & ~i_8_200_2247_0))) | (~i_8_200_571_0 & ~i_8_200_888_0 & ~i_8_200_1179_0 & ~i_8_200_1587_0 & ~i_8_200_1699_0 & i_8_200_1821_0))) | (i_8_200_221_0 & i_8_200_888_0 & i_8_200_2222_0))) | (~i_8_200_1585_0 & ((~i_8_200_1490_0 & ((~i_8_200_1584_0 & ((~i_8_200_111_0 & ((~i_8_200_114_0 & ~i_8_200_115_0 & ~i_8_200_575_0 & ~i_8_200_776_0 & ~i_8_200_888_0 & ~i_8_200_1179_0 & ~i_8_200_1262_0 & ~i_8_200_1623_0 & ~i_8_200_1770_0 & ~i_8_200_2129_0) | (i_8_200_219_0 & ~i_8_200_1167_0 & ~i_8_200_1487_0 & ~i_8_200_1695_0 & ~i_8_200_1700_0 & ~i_8_200_2222_0))) | (~i_8_200_114_0 & ~i_8_200_224_0 & ~i_8_200_571_0 & ~i_8_200_575_0 & ~i_8_200_776_0 & ~i_8_200_888_0 & ~i_8_200_1167_0 & ~i_8_200_1179_0 & ~i_8_200_1180_0 & ~i_8_200_1263_0 & ~i_8_200_1587_0 & ~i_8_200_1588_0 & ~i_8_200_1696_0 & ~i_8_200_1758_0 & ~i_8_200_2222_0))) | (~i_8_200_114_0 & i_8_200_703_0 & ~i_8_200_888_0 & ~i_8_200_1278_0 & ~i_8_200_1758_0 & ~i_8_200_2073_0))) | (~i_8_200_1695_0 & ((i_8_200_220_0 & ~i_8_200_572_0 & ((~i_8_200_50_0 & ~i_8_200_775_0 & ~i_8_200_888_0 & ~i_8_200_959_0 & ~i_8_200_1699_0 & ~i_8_200_1772_0) | (~i_8_200_116_0 & ~i_8_200_607_0 & ~i_8_200_1167_0 & ~i_8_200_1179_0 & ~i_8_200_1683_0 & ~i_8_200_1758_0 & ~i_8_200_2249_0))) | (i_8_200_775_0 & ~i_8_200_776_0 & ~i_8_200_959_0 & ~i_8_200_966_0 & ~i_8_200_1263_0 & ~i_8_200_1696_0 & ~i_8_200_1746_0 & ~i_8_200_1770_0))) | (~i_8_200_1587_0 & ((i_8_200_111_0 & ~i_8_200_601_0 & i_8_200_703_0 & ~i_8_200_1278_0 & i_8_200_1818_0 & i_8_200_1821_0) | (i_8_200_221_0 & ~i_8_200_689_0 & i_8_200_2261_0))) | (i_8_200_219_0 & i_8_200_657_0 & ~i_8_200_1857_0 & i_8_200_2247_0) | (~i_8_200_455_0 & ~i_8_200_775_0 & ~i_8_200_887_0 & ~i_8_200_1487_0 & ~i_8_200_1588_0 & ~i_8_200_1683_0 & ~i_8_200_1696_0 & i_8_200_1820_0 & ~i_8_200_2249_0))) | (~i_8_200_124_0 & ((~i_8_200_111_0 & ((~i_8_200_115_0 & i_8_200_383_0 & ~i_8_200_572_0 & ~i_8_200_887_0 & ~i_8_200_1072_0 & ~i_8_200_1178_0 & ~i_8_200_1262_0 & ~i_8_200_1632_0 & ~i_8_200_2129_0 & ~i_8_200_2226_0) | (i_8_200_523_0 & ~i_8_200_1167_0 & ~i_8_200_1487_0 & ~i_8_200_1588_0 & i_8_200_1632_0 & ~i_8_200_2293_0))) | (~i_8_200_114_0 & ~i_8_200_1584_0 & ~i_8_200_1623_0 & ((~i_8_200_523_0 & ~i_8_200_575_0 & i_8_200_2226_0) | (~i_8_200_116_0 & ~i_8_200_572_0 & ~i_8_200_607_0 & ~i_8_200_775_0 & ~i_8_200_1179_0 & ~i_8_200_1490_0 & ~i_8_200_1738_0 & ~i_8_200_1758_0 & ~i_8_200_2129_0 & ~i_8_200_2222_0 & ~i_8_200_2247_0))) | (~i_8_200_1738_0 & ~i_8_200_2247_0 & ((~i_8_200_116_0 & ~i_8_200_575_0 & ~i_8_200_776_0 & ~i_8_200_1072_0 & ~i_8_200_1179_0 & ~i_8_200_1262_0 & ~i_8_200_1263_0 & ~i_8_200_1490_0 & ~i_8_200_1683_0 & ~i_8_200_1695_0 & ~i_8_200_1699_0 & ~i_8_200_1746_0 & ~i_8_200_1854_0 & ~i_8_200_1857_0 & ~i_8_200_1758_0 & ~i_8_200_1821_0) | (~i_8_200_25_0 & i_8_200_657_0 & i_8_200_1072_0 & ~i_8_200_1588_0 & ~i_8_200_2129_0))))) | (~i_8_200_115_0 & ((~i_8_200_116_0 & ~i_8_200_455_0 & ~i_8_200_571_0 & ~i_8_200_575_0 & ~i_8_200_607_0 & ~i_8_200_776_0 & ~i_8_200_883_0 & ~i_8_200_888_0 & ~i_8_200_1180_0 & ~i_8_200_1584_0 & ~i_8_200_1696_0 & ~i_8_200_1699_0 & ~i_8_200_1700_0 & ~i_8_200_1758_0 & ~i_8_200_1854_0 & ~i_8_200_2073_0 & ~i_8_200_2247_0 & ~i_8_200_2248_0) | (~i_8_200_114_0 & ~i_8_200_602_0 & ~i_8_200_1787_0 & i_8_200_1969_0 & i_8_200_2249_0))) | (~i_8_200_887_0 & ((~i_8_200_114_0 & ~i_8_200_1262_0 & ((~i_8_200_572_0 & ~i_8_200_575_0 & ~i_8_200_601_0 & ~i_8_200_966_0 & ~i_8_200_1167_0 & ~i_8_200_1180_0 & ~i_8_200_1263_0 & ~i_8_200_1296_0 & ~i_8_200_1588_0 & ~i_8_200_1695_0 & ~i_8_200_1696_0 & ~i_8_200_1746_0 & ~i_8_200_1818_0 & ~i_8_200_1857_0 & ~i_8_200_2129_0 & ~i_8_200_2247_0) | (i_8_200_602_0 & ~i_8_200_888_0 & ~i_8_200_1278_0 & ~i_8_200_2293_0))) | (~i_8_200_1772_0 & ((~i_8_200_703_0 & ~i_8_200_966_0 & ~i_8_200_1180_0 & ~i_8_200_1263_0 & ~i_8_200_1588_0 & i_8_200_2009_0) | (i_8_200_25_0 & ~i_8_200_571_0 & ~i_8_200_888_0 & ~i_8_200_1487_0 & ~i_8_200_1584_0 & ~i_8_200_2248_0))))) | (~i_8_200_1263_0 & ((~i_8_200_116_0 & ((~i_8_200_658_0 & i_8_200_689_0 & ~i_8_200_798_0 & ~i_8_200_959_0 & ~i_8_200_961_0 & ~i_8_200_1587_0 & ~i_8_200_1588_0 & ~i_8_200_1696_0 & ~i_8_200_2073_0) | (~i_8_200_1584_0 & ~i_8_200_1623_0 & i_8_200_1632_0 & ~i_8_200_2222_0))) | (~i_8_200_575_0 & i_8_200_704_0 & i_8_200_887_0 & ~i_8_200_959_0 & ~i_8_200_1178_0 & ~i_8_200_1180_0 & ~i_8_200_2009_0 & ~i_8_200_2222_0) | (i_8_200_1470_0 & ~i_8_200_1696_0 & i_8_200_1746_0 & ~i_8_200_1772_0 & ~i_8_200_1818_0 & ~i_8_200_2129_0))) | (i_8_200_220_0 & i_8_200_221_0 & ((~i_8_200_572_0 & i_8_200_1227_0 & ~i_8_200_1623_0) | (i_8_200_224_0 & i_8_200_1229_0 & ~i_8_200_1584_0 & ~i_8_200_1587_0 & ~i_8_200_1738_0 & ~i_8_200_1758_0))) | (i_8_200_455_0 & ~i_8_200_1180_0 & ((~i_8_200_775_0 & i_8_200_959_0) | (~i_8_200_523_0 & ~i_8_200_959_0 & ~i_8_200_1487_0 & ~i_8_200_1564_0 & ~i_8_200_1623_0 & ~i_8_200_1700_0))) | (~i_8_200_575_0 & ((~i_8_200_658_0 & i_8_200_1228_0 & i_8_200_1229_0 & ~i_8_200_2222_0) | (i_8_200_224_0 & ~i_8_200_704_0 & ~i_8_200_776_0 & ~i_8_200_1167_0 & ~i_8_200_1278_0 & ~i_8_200_1487_0 & ~i_8_200_1696_0 & ~i_8_200_1969_0 & ~i_8_200_2226_0 & ~i_8_200_2248_0))) | (~i_8_200_1695_0 & ((i_8_200_1227_0 & ((~i_8_200_1179_0 & i_8_200_1560_0) | (~i_8_200_1588_0 & i_8_200_1623_0 & i_8_200_1699_0 & ~i_8_200_2226_0))) | (i_8_200_2129_0 & ((~i_8_200_1789_0 & i_8_200_1818_0 & ~i_8_200_1820_0) | (~i_8_200_1262_0 & ~i_8_200_1490_0 & i_8_200_2224_0))) | (i_8_200_523_0 & ~i_8_200_572_0 & ~i_8_200_776_0 & ~i_8_200_1588_0 & i_8_200_1820_0 & ~i_8_200_2247_0 & ~i_8_200_2248_0 & ~i_8_200_2261_0))) | (~i_8_200_453_0 & ~i_8_200_523_0 & i_8_200_966_0 & ~i_8_200_1584_0 & ~i_8_200_1623_0 & i_8_200_1696_0 & ~i_8_200_1700_0 & ~i_8_200_1738_0 & ~i_8_200_2073_0) | (~i_8_200_775_0 & ~i_8_200_966_0 & i_8_200_1229_0 & ~i_8_200_1490_0 & ~i_8_200_1564_0 & ~i_8_200_2247_0) | (~i_8_200_224_0 & i_8_200_383_0 & ~i_8_200_458_0 & ~i_8_200_689_0 & i_8_200_1262_0 & i_8_200_1487_0 & ~i_8_200_2248_0));
endmodule



// Benchmark "kernel_8_201" written by ABC on Sun Jul 19 10:06:33 2020

module kernel_8_201 ( 
    i_8_201_21_0, i_8_201_25_0, i_8_201_33_0, i_8_201_34_0, i_8_201_85_0,
    i_8_201_183_0, i_8_201_190_0, i_8_201_294_0, i_8_201_300_0,
    i_8_201_373_0, i_8_201_386_0, i_8_201_420_0, i_8_201_481_0,
    i_8_201_483_0, i_8_201_508_0, i_8_201_510_0, i_8_201_529_0,
    i_8_201_530_0, i_8_201_589_0, i_8_201_592_0, i_8_201_594_0,
    i_8_201_595_0, i_8_201_598_0, i_8_201_601_0, i_8_201_607_0,
    i_8_201_634_0, i_8_201_636_0, i_8_201_691_0, i_8_201_714_0,
    i_8_201_715_0, i_8_201_717_0, i_8_201_759_0, i_8_201_777_0,
    i_8_201_778_0, i_8_201_789_0, i_8_201_790_0, i_8_201_800_0,
    i_8_201_810_0, i_8_201_838_0, i_8_201_852_0, i_8_201_853_0,
    i_8_201_912_0, i_8_201_933_0, i_8_201_997_0, i_8_201_1005_0,
    i_8_201_1059_0, i_8_201_1093_0, i_8_201_1114_0, i_8_201_1123_0,
    i_8_201_1129_0, i_8_201_1159_0, i_8_201_1222_0, i_8_201_1277_0,
    i_8_201_1282_0, i_8_201_1285_0, i_8_201_1286_0, i_8_201_1307_0,
    i_8_201_1320_0, i_8_201_1321_0, i_8_201_1330_0, i_8_201_1366_0,
    i_8_201_1431_0, i_8_201_1451_0, i_8_201_1470_0, i_8_201_1471_0,
    i_8_201_1473_0, i_8_201_1474_0, i_8_201_1537_0, i_8_201_1543_0,
    i_8_201_1545_0, i_8_201_1548_0, i_8_201_1563_0, i_8_201_1570_0,
    i_8_201_1590_0, i_8_201_1668_0, i_8_201_1671_0, i_8_201_1681_0,
    i_8_201_1682_0, i_8_201_1723_0, i_8_201_1743_0, i_8_201_1749_0,
    i_8_201_1750_0, i_8_201_1753_0, i_8_201_1875_0, i_8_201_1876_0,
    i_8_201_1878_0, i_8_201_1920_0, i_8_201_1959_0, i_8_201_1960_0,
    i_8_201_1965_0, i_8_201_1969_0, i_8_201_1971_0, i_8_201_1995_0,
    i_8_201_2011_0, i_8_201_2137_0, i_8_201_2235_0, i_8_201_2253_0,
    i_8_201_2277_0, i_8_201_2284_0, i_8_201_2292_0,
    o_8_201_0_0  );
  input  i_8_201_21_0, i_8_201_25_0, i_8_201_33_0, i_8_201_34_0,
    i_8_201_85_0, i_8_201_183_0, i_8_201_190_0, i_8_201_294_0,
    i_8_201_300_0, i_8_201_373_0, i_8_201_386_0, i_8_201_420_0,
    i_8_201_481_0, i_8_201_483_0, i_8_201_508_0, i_8_201_510_0,
    i_8_201_529_0, i_8_201_530_0, i_8_201_589_0, i_8_201_592_0,
    i_8_201_594_0, i_8_201_595_0, i_8_201_598_0, i_8_201_601_0,
    i_8_201_607_0, i_8_201_634_0, i_8_201_636_0, i_8_201_691_0,
    i_8_201_714_0, i_8_201_715_0, i_8_201_717_0, i_8_201_759_0,
    i_8_201_777_0, i_8_201_778_0, i_8_201_789_0, i_8_201_790_0,
    i_8_201_800_0, i_8_201_810_0, i_8_201_838_0, i_8_201_852_0,
    i_8_201_853_0, i_8_201_912_0, i_8_201_933_0, i_8_201_997_0,
    i_8_201_1005_0, i_8_201_1059_0, i_8_201_1093_0, i_8_201_1114_0,
    i_8_201_1123_0, i_8_201_1129_0, i_8_201_1159_0, i_8_201_1222_0,
    i_8_201_1277_0, i_8_201_1282_0, i_8_201_1285_0, i_8_201_1286_0,
    i_8_201_1307_0, i_8_201_1320_0, i_8_201_1321_0, i_8_201_1330_0,
    i_8_201_1366_0, i_8_201_1431_0, i_8_201_1451_0, i_8_201_1470_0,
    i_8_201_1471_0, i_8_201_1473_0, i_8_201_1474_0, i_8_201_1537_0,
    i_8_201_1543_0, i_8_201_1545_0, i_8_201_1548_0, i_8_201_1563_0,
    i_8_201_1570_0, i_8_201_1590_0, i_8_201_1668_0, i_8_201_1671_0,
    i_8_201_1681_0, i_8_201_1682_0, i_8_201_1723_0, i_8_201_1743_0,
    i_8_201_1749_0, i_8_201_1750_0, i_8_201_1753_0, i_8_201_1875_0,
    i_8_201_1876_0, i_8_201_1878_0, i_8_201_1920_0, i_8_201_1959_0,
    i_8_201_1960_0, i_8_201_1965_0, i_8_201_1969_0, i_8_201_1971_0,
    i_8_201_1995_0, i_8_201_2011_0, i_8_201_2137_0, i_8_201_2235_0,
    i_8_201_2253_0, i_8_201_2277_0, i_8_201_2284_0, i_8_201_2292_0;
  output o_8_201_0_0;
  assign o_8_201_0_0 = 0;
endmodule



// Benchmark "kernel_8_202" written by ABC on Sun Jul 19 10:06:34 2020

module kernel_8_202 ( 
    i_8_202_1_0, i_8_202_19_0, i_8_202_73_0, i_8_202_76_0, i_8_202_82_0,
    i_8_202_188_0, i_8_202_202_0, i_8_202_244_0, i_8_202_268_0,
    i_8_202_274_0, i_8_202_275_0, i_8_202_325_0, i_8_202_335_0,
    i_8_202_343_0, i_8_202_352_0, i_8_202_353_0, i_8_202_373_0,
    i_8_202_426_0, i_8_202_459_0, i_8_202_478_0, i_8_202_500_0,
    i_8_202_513_0, i_8_202_514_0, i_8_202_515_0, i_8_202_523_0,
    i_8_202_613_0, i_8_202_631_0, i_8_202_662_0, i_8_202_663_0,
    i_8_202_729_0, i_8_202_731_0, i_8_202_751_0, i_8_202_756_0,
    i_8_202_811_0, i_8_202_812_0, i_8_202_819_0, i_8_202_864_0,
    i_8_202_910_0, i_8_202_950_0, i_8_202_973_0, i_8_202_1029_0,
    i_8_202_1057_0, i_8_202_1072_0, i_8_202_1108_0, i_8_202_1170_0,
    i_8_202_1187_0, i_8_202_1188_0, i_8_202_1225_0, i_8_202_1226_0,
    i_8_202_1238_0, i_8_202_1261_0, i_8_202_1330_0, i_8_202_1355_0,
    i_8_202_1408_0, i_8_202_1429_0, i_8_202_1454_0, i_8_202_1468_0,
    i_8_202_1471_0, i_8_202_1494_0, i_8_202_1495_0, i_8_202_1496_0,
    i_8_202_1507_0, i_8_202_1509_0, i_8_202_1542_0, i_8_202_1561_0,
    i_8_202_1624_0, i_8_202_1641_0, i_8_202_1649_0, i_8_202_1656_0,
    i_8_202_1694_0, i_8_202_1702_0, i_8_202_1751_0, i_8_202_1800_0,
    i_8_202_1804_0, i_8_202_1810_0, i_8_202_1855_0, i_8_202_1864_0,
    i_8_202_1865_0, i_8_202_1873_0, i_8_202_1874_0, i_8_202_1963_0,
    i_8_202_1968_0, i_8_202_1973_0, i_8_202_1992_0, i_8_202_1994_0,
    i_8_202_2008_0, i_8_202_2045_0, i_8_202_2056_0, i_8_202_2062_0,
    i_8_202_2063_0, i_8_202_2071_0, i_8_202_2116_0, i_8_202_2117_0,
    i_8_202_2118_0, i_8_202_2130_0, i_8_202_2143_0, i_8_202_2170_0,
    i_8_202_2228_0, i_8_202_2234_0, i_8_202_2253_0,
    o_8_202_0_0  );
  input  i_8_202_1_0, i_8_202_19_0, i_8_202_73_0, i_8_202_76_0,
    i_8_202_82_0, i_8_202_188_0, i_8_202_202_0, i_8_202_244_0,
    i_8_202_268_0, i_8_202_274_0, i_8_202_275_0, i_8_202_325_0,
    i_8_202_335_0, i_8_202_343_0, i_8_202_352_0, i_8_202_353_0,
    i_8_202_373_0, i_8_202_426_0, i_8_202_459_0, i_8_202_478_0,
    i_8_202_500_0, i_8_202_513_0, i_8_202_514_0, i_8_202_515_0,
    i_8_202_523_0, i_8_202_613_0, i_8_202_631_0, i_8_202_662_0,
    i_8_202_663_0, i_8_202_729_0, i_8_202_731_0, i_8_202_751_0,
    i_8_202_756_0, i_8_202_811_0, i_8_202_812_0, i_8_202_819_0,
    i_8_202_864_0, i_8_202_910_0, i_8_202_950_0, i_8_202_973_0,
    i_8_202_1029_0, i_8_202_1057_0, i_8_202_1072_0, i_8_202_1108_0,
    i_8_202_1170_0, i_8_202_1187_0, i_8_202_1188_0, i_8_202_1225_0,
    i_8_202_1226_0, i_8_202_1238_0, i_8_202_1261_0, i_8_202_1330_0,
    i_8_202_1355_0, i_8_202_1408_0, i_8_202_1429_0, i_8_202_1454_0,
    i_8_202_1468_0, i_8_202_1471_0, i_8_202_1494_0, i_8_202_1495_0,
    i_8_202_1496_0, i_8_202_1507_0, i_8_202_1509_0, i_8_202_1542_0,
    i_8_202_1561_0, i_8_202_1624_0, i_8_202_1641_0, i_8_202_1649_0,
    i_8_202_1656_0, i_8_202_1694_0, i_8_202_1702_0, i_8_202_1751_0,
    i_8_202_1800_0, i_8_202_1804_0, i_8_202_1810_0, i_8_202_1855_0,
    i_8_202_1864_0, i_8_202_1865_0, i_8_202_1873_0, i_8_202_1874_0,
    i_8_202_1963_0, i_8_202_1968_0, i_8_202_1973_0, i_8_202_1992_0,
    i_8_202_1994_0, i_8_202_2008_0, i_8_202_2045_0, i_8_202_2056_0,
    i_8_202_2062_0, i_8_202_2063_0, i_8_202_2071_0, i_8_202_2116_0,
    i_8_202_2117_0, i_8_202_2118_0, i_8_202_2130_0, i_8_202_2143_0,
    i_8_202_2170_0, i_8_202_2228_0, i_8_202_2234_0, i_8_202_2253_0;
  output o_8_202_0_0;
  assign o_8_202_0_0 = ~((~i_8_202_1_0 & ((~i_8_202_244_0 & ~i_8_202_353_0 & ~i_8_202_751_0 & ~i_8_202_1261_0 & ~i_8_202_1355_0 & ~i_8_202_1494_0 & ~i_8_202_1641_0 & ~i_8_202_1994_0 & ~i_8_202_2116_0) | (~i_8_202_729_0 & ~i_8_202_1226_0 & ~i_8_202_1542_0 & ~i_8_202_1992_0 & ~i_8_202_2045_0 & ~i_8_202_2063_0 & ~i_8_202_2228_0))) | (~i_8_202_352_0 & ((~i_8_202_82_0 & ~i_8_202_514_0 & ~i_8_202_756_0 & ~i_8_202_811_0 & ~i_8_202_812_0 & ~i_8_202_1238_0 & ~i_8_202_1865_0) | (i_8_202_500_0 & ~i_8_202_1408_0 & ~i_8_202_2062_0 & i_8_202_2234_0))) | (~i_8_202_515_0 & ((~i_8_202_19_0 & ~i_8_202_514_0 & ~i_8_202_1496_0 & ~i_8_202_1641_0 & ~i_8_202_1804_0 & ~i_8_202_1864_0) | (~i_8_202_1330_0 & ~i_8_202_1509_0 & ~i_8_202_1874_0 & ~i_8_202_2063_0 & i_8_202_2071_0 & ~i_8_202_2116_0 & ~i_8_202_2228_0))) | (~i_8_202_812_0 & ~i_8_202_2045_0 & ((~i_8_202_1468_0 & ~i_8_202_1495_0 & ~i_8_202_1656_0 & ~i_8_202_1865_0 & ~i_8_202_1873_0 & ~i_8_202_1874_0 & ~i_8_202_2008_0) | (~i_8_202_729_0 & ~i_8_202_1429_0 & ~i_8_202_1542_0 & ~i_8_202_1694_0 & ~i_8_202_2116_0 & i_8_202_2228_0))) | (~i_8_202_2062_0 & ((~i_8_202_1170_0 & ~i_8_202_1225_0 & ((~i_8_202_631_0 & ~i_8_202_1072_0 & ~i_8_202_1496_0 & ~i_8_202_2008_0 & ~i_8_202_2118_0) | (~i_8_202_1494_0 & ~i_8_202_1865_0 & ~i_8_202_2234_0))) | (i_8_202_613_0 & ~i_8_202_731_0 & ~i_8_202_1509_0 & i_8_202_1694_0))) | (~i_8_202_514_0 & ((~i_8_202_731_0 & ((~i_8_202_343_0 & ~i_8_202_663_0 & ~i_8_202_1494_0 & ~i_8_202_1495_0 & ~i_8_202_1624_0 & ~i_8_202_1656_0 & ~i_8_202_1874_0 & ~i_8_202_2063_0) | (~i_8_202_353_0 & ~i_8_202_1226_0 & ~i_8_202_1542_0 & ~i_8_202_1865_0 & ~i_8_202_2118_0 & ~i_8_202_2170_0))) | (~i_8_202_662_0 & i_8_202_1225_0 & ~i_8_202_1454_0 & ~i_8_202_1494_0 & ~i_8_202_1507_0 & ~i_8_202_1800_0 & ~i_8_202_1804_0 & ~i_8_202_2117_0))) | (i_8_202_515_0 & i_8_202_1542_0 & i_8_202_2056_0) | (~i_8_202_500_0 & ~i_8_202_613_0 & ~i_8_202_1496_0 & ~i_8_202_1656_0 & ~i_8_202_1800_0 & ~i_8_202_1810_0 & ~i_8_202_2056_0));
endmodule



// Benchmark "kernel_8_203" written by ABC on Sun Jul 19 10:06:35 2020

module kernel_8_203 ( 
    i_8_203_25_0, i_8_203_27_0, i_8_203_46_0, i_8_203_54_0, i_8_203_57_0,
    i_8_203_70_0, i_8_203_104_0, i_8_203_171_0, i_8_203_172_0,
    i_8_203_197_0, i_8_203_337_0, i_8_203_372_0, i_8_203_415_0,
    i_8_203_423_0, i_8_203_427_0, i_8_203_450_0, i_8_203_453_0,
    i_8_203_549_0, i_8_203_571_0, i_8_203_586_0, i_8_203_594_0,
    i_8_203_598_0, i_8_203_599_0, i_8_203_604_0, i_8_203_632_0,
    i_8_203_633_0, i_8_203_640_0, i_8_203_658_0, i_8_203_662_0,
    i_8_203_679_0, i_8_203_695_0, i_8_203_704_0, i_8_203_778_0,
    i_8_203_781_0, i_8_203_835_0, i_8_203_837_0, i_8_203_865_0,
    i_8_203_880_0, i_8_203_993_0, i_8_203_1035_0, i_8_203_1063_0,
    i_8_203_1137_0, i_8_203_1154_0, i_8_203_1178_0, i_8_203_1264_0,
    i_8_203_1281_0, i_8_203_1297_0, i_8_203_1298_0, i_8_203_1299_0,
    i_8_203_1367_0, i_8_203_1406_0, i_8_203_1470_0, i_8_203_1471_0,
    i_8_203_1557_0, i_8_203_1558_0, i_8_203_1559_0, i_8_203_1571_0,
    i_8_203_1602_0, i_8_203_1603_0, i_8_203_1611_0, i_8_203_1612_0,
    i_8_203_1629_0, i_8_203_1635_0, i_8_203_1646_0, i_8_203_1655_0,
    i_8_203_1686_0, i_8_203_1690_0, i_8_203_1710_0, i_8_203_1711_0,
    i_8_203_1713_0, i_8_203_1750_0, i_8_203_1753_0, i_8_203_1754_0,
    i_8_203_1755_0, i_8_203_1758_0, i_8_203_1759_0, i_8_203_1774_0,
    i_8_203_1780_0, i_8_203_1809_0, i_8_203_1819_0, i_8_203_1824_0,
    i_8_203_1889_0, i_8_203_1971_0, i_8_203_1980_0, i_8_203_1989_0,
    i_8_203_1993_0, i_8_203_1994_0, i_8_203_1996_0, i_8_203_2052_0,
    i_8_203_2053_0, i_8_203_2069_0, i_8_203_2106_0, i_8_203_2116_0,
    i_8_203_2147_0, i_8_203_2149_0, i_8_203_2223_0, i_8_203_2233_0,
    i_8_203_2235_0, i_8_203_2244_0, i_8_203_2259_0,
    o_8_203_0_0  );
  input  i_8_203_25_0, i_8_203_27_0, i_8_203_46_0, i_8_203_54_0,
    i_8_203_57_0, i_8_203_70_0, i_8_203_104_0, i_8_203_171_0,
    i_8_203_172_0, i_8_203_197_0, i_8_203_337_0, i_8_203_372_0,
    i_8_203_415_0, i_8_203_423_0, i_8_203_427_0, i_8_203_450_0,
    i_8_203_453_0, i_8_203_549_0, i_8_203_571_0, i_8_203_586_0,
    i_8_203_594_0, i_8_203_598_0, i_8_203_599_0, i_8_203_604_0,
    i_8_203_632_0, i_8_203_633_0, i_8_203_640_0, i_8_203_658_0,
    i_8_203_662_0, i_8_203_679_0, i_8_203_695_0, i_8_203_704_0,
    i_8_203_778_0, i_8_203_781_0, i_8_203_835_0, i_8_203_837_0,
    i_8_203_865_0, i_8_203_880_0, i_8_203_993_0, i_8_203_1035_0,
    i_8_203_1063_0, i_8_203_1137_0, i_8_203_1154_0, i_8_203_1178_0,
    i_8_203_1264_0, i_8_203_1281_0, i_8_203_1297_0, i_8_203_1298_0,
    i_8_203_1299_0, i_8_203_1367_0, i_8_203_1406_0, i_8_203_1470_0,
    i_8_203_1471_0, i_8_203_1557_0, i_8_203_1558_0, i_8_203_1559_0,
    i_8_203_1571_0, i_8_203_1602_0, i_8_203_1603_0, i_8_203_1611_0,
    i_8_203_1612_0, i_8_203_1629_0, i_8_203_1635_0, i_8_203_1646_0,
    i_8_203_1655_0, i_8_203_1686_0, i_8_203_1690_0, i_8_203_1710_0,
    i_8_203_1711_0, i_8_203_1713_0, i_8_203_1750_0, i_8_203_1753_0,
    i_8_203_1754_0, i_8_203_1755_0, i_8_203_1758_0, i_8_203_1759_0,
    i_8_203_1774_0, i_8_203_1780_0, i_8_203_1809_0, i_8_203_1819_0,
    i_8_203_1824_0, i_8_203_1889_0, i_8_203_1971_0, i_8_203_1980_0,
    i_8_203_1989_0, i_8_203_1993_0, i_8_203_1994_0, i_8_203_1996_0,
    i_8_203_2052_0, i_8_203_2053_0, i_8_203_2069_0, i_8_203_2106_0,
    i_8_203_2116_0, i_8_203_2147_0, i_8_203_2149_0, i_8_203_2223_0,
    i_8_203_2233_0, i_8_203_2235_0, i_8_203_2244_0, i_8_203_2259_0;
  output o_8_203_0_0;
  assign o_8_203_0_0 = 0;
endmodule



// Benchmark "kernel_8_204" written by ABC on Sun Jul 19 10:06:36 2020

module kernel_8_204 ( 
    i_8_204_32_0, i_8_204_73_0, i_8_204_82_0, i_8_204_88_0, i_8_204_90_0,
    i_8_204_104_0, i_8_204_182_0, i_8_204_216_0, i_8_204_217_0,
    i_8_204_220_0, i_8_204_244_0, i_8_204_300_0, i_8_204_319_0,
    i_8_204_349_0, i_8_204_364_0, i_8_204_369_0, i_8_204_380_0,
    i_8_204_385_0, i_8_204_388_0, i_8_204_460_0, i_8_204_471_0,
    i_8_204_496_0, i_8_204_515_0, i_8_204_528_0, i_8_204_552_0,
    i_8_204_555_0, i_8_204_623_0, i_8_204_657_0, i_8_204_659_0,
    i_8_204_664_0, i_8_204_665_0, i_8_204_693_0, i_8_204_711_0,
    i_8_204_737_0, i_8_204_778_0, i_8_204_779_0, i_8_204_783_0,
    i_8_204_793_0, i_8_204_830_0, i_8_204_844_0, i_8_204_874_0,
    i_8_204_967_0, i_8_204_970_0, i_8_204_998_0, i_8_204_1042_0,
    i_8_204_1071_0, i_8_204_1079_0, i_8_204_1104_0, i_8_204_1105_0,
    i_8_204_1110_0, i_8_204_1111_0, i_8_204_1151_0, i_8_204_1224_0,
    i_8_204_1225_0, i_8_204_1246_0, i_8_204_1260_0, i_8_204_1279_0,
    i_8_204_1281_0, i_8_204_1283_0, i_8_204_1306_0, i_8_204_1359_0,
    i_8_204_1397_0, i_8_204_1477_0, i_8_204_1486_0, i_8_204_1487_0,
    i_8_204_1522_0, i_8_204_1537_0, i_8_204_1538_0, i_8_204_1541_0,
    i_8_204_1549_0, i_8_204_1567_0, i_8_204_1594_0, i_8_204_1602_0,
    i_8_204_1649_0, i_8_204_1670_0, i_8_204_1680_0, i_8_204_1719_0,
    i_8_204_1720_0, i_8_204_1746_0, i_8_204_1752_0, i_8_204_1800_0,
    i_8_204_1803_0, i_8_204_1815_0, i_8_204_1816_0, i_8_204_1891_0,
    i_8_204_1910_0, i_8_204_1948_0, i_8_204_1962_0, i_8_204_1963_0,
    i_8_204_1969_0, i_8_204_1972_0, i_8_204_1989_0, i_8_204_2047_0,
    i_8_204_2071_0, i_8_204_2106_0, i_8_204_2107_0, i_8_204_2113_0,
    i_8_204_2133_0, i_8_204_2140_0, i_8_204_2141_0,
    o_8_204_0_0  );
  input  i_8_204_32_0, i_8_204_73_0, i_8_204_82_0, i_8_204_88_0,
    i_8_204_90_0, i_8_204_104_0, i_8_204_182_0, i_8_204_216_0,
    i_8_204_217_0, i_8_204_220_0, i_8_204_244_0, i_8_204_300_0,
    i_8_204_319_0, i_8_204_349_0, i_8_204_364_0, i_8_204_369_0,
    i_8_204_380_0, i_8_204_385_0, i_8_204_388_0, i_8_204_460_0,
    i_8_204_471_0, i_8_204_496_0, i_8_204_515_0, i_8_204_528_0,
    i_8_204_552_0, i_8_204_555_0, i_8_204_623_0, i_8_204_657_0,
    i_8_204_659_0, i_8_204_664_0, i_8_204_665_0, i_8_204_693_0,
    i_8_204_711_0, i_8_204_737_0, i_8_204_778_0, i_8_204_779_0,
    i_8_204_783_0, i_8_204_793_0, i_8_204_830_0, i_8_204_844_0,
    i_8_204_874_0, i_8_204_967_0, i_8_204_970_0, i_8_204_998_0,
    i_8_204_1042_0, i_8_204_1071_0, i_8_204_1079_0, i_8_204_1104_0,
    i_8_204_1105_0, i_8_204_1110_0, i_8_204_1111_0, i_8_204_1151_0,
    i_8_204_1224_0, i_8_204_1225_0, i_8_204_1246_0, i_8_204_1260_0,
    i_8_204_1279_0, i_8_204_1281_0, i_8_204_1283_0, i_8_204_1306_0,
    i_8_204_1359_0, i_8_204_1397_0, i_8_204_1477_0, i_8_204_1486_0,
    i_8_204_1487_0, i_8_204_1522_0, i_8_204_1537_0, i_8_204_1538_0,
    i_8_204_1541_0, i_8_204_1549_0, i_8_204_1567_0, i_8_204_1594_0,
    i_8_204_1602_0, i_8_204_1649_0, i_8_204_1670_0, i_8_204_1680_0,
    i_8_204_1719_0, i_8_204_1720_0, i_8_204_1746_0, i_8_204_1752_0,
    i_8_204_1800_0, i_8_204_1803_0, i_8_204_1815_0, i_8_204_1816_0,
    i_8_204_1891_0, i_8_204_1910_0, i_8_204_1948_0, i_8_204_1962_0,
    i_8_204_1963_0, i_8_204_1969_0, i_8_204_1972_0, i_8_204_1989_0,
    i_8_204_2047_0, i_8_204_2071_0, i_8_204_2106_0, i_8_204_2107_0,
    i_8_204_2113_0, i_8_204_2133_0, i_8_204_2140_0, i_8_204_2141_0;
  output o_8_204_0_0;
  assign o_8_204_0_0 = 0;
endmodule



// Benchmark "kernel_8_205" written by ABC on Sun Jul 19 10:06:37 2020

module kernel_8_205 ( 
    i_8_205_34_0, i_8_205_85_0, i_8_205_158_0, i_8_205_181_0,
    i_8_205_184_0, i_8_205_203_0, i_8_205_217_0, i_8_205_220_0,
    i_8_205_233_0, i_8_205_237_0, i_8_205_238_0, i_8_205_255_0,
    i_8_205_304_0, i_8_205_371_0, i_8_205_374_0, i_8_205_380_0,
    i_8_205_382_0, i_8_205_385_0, i_8_205_423_0, i_8_205_437_0,
    i_8_205_453_0, i_8_205_477_0, i_8_205_478_0, i_8_205_481_0,
    i_8_205_482_0, i_8_205_484_0, i_8_205_485_0, i_8_205_498_0,
    i_8_205_499_0, i_8_205_505_0, i_8_205_523_0, i_8_205_526_0,
    i_8_205_532_0, i_8_205_564_0, i_8_205_634_0, i_8_205_661_0,
    i_8_205_684_0, i_8_205_703_0, i_8_205_757_0, i_8_205_759_0,
    i_8_205_760_0, i_8_205_761_0, i_8_205_767_0, i_8_205_780_0,
    i_8_205_811_0, i_8_205_823_0, i_8_205_830_0, i_8_205_869_0,
    i_8_205_892_0, i_8_205_904_0, i_8_205_1013_0, i_8_205_1030_0,
    i_8_205_1111_0, i_8_205_1112_0, i_8_205_1135_0, i_8_205_1174_0,
    i_8_205_1282_0, i_8_205_1294_0, i_8_205_1309_0, i_8_205_1328_0,
    i_8_205_1363_0, i_8_205_1366_0, i_8_205_1398_0, i_8_205_1506_0,
    i_8_205_1522_0, i_8_205_1537_0, i_8_205_1552_0, i_8_205_1565_0,
    i_8_205_1577_0, i_8_205_1605_0, i_8_205_1676_0, i_8_205_1678_0,
    i_8_205_1711_0, i_8_205_1723_0, i_8_205_1729_0, i_8_205_1730_0,
    i_8_205_1749_0, i_8_205_1752_0, i_8_205_1760_0, i_8_205_1805_0,
    i_8_205_1807_0, i_8_205_1818_0, i_8_205_1855_0, i_8_205_1903_0,
    i_8_205_1920_0, i_8_205_1947_0, i_8_205_1980_0, i_8_205_2020_0,
    i_8_205_2037_0, i_8_205_2038_0, i_8_205_2070_0, i_8_205_2093_0,
    i_8_205_2109_0, i_8_205_2150_0, i_8_205_2170_0, i_8_205_2218_0,
    i_8_205_2224_0, i_8_205_2237_0, i_8_205_2271_0, i_8_205_2286_0,
    o_8_205_0_0  );
  input  i_8_205_34_0, i_8_205_85_0, i_8_205_158_0, i_8_205_181_0,
    i_8_205_184_0, i_8_205_203_0, i_8_205_217_0, i_8_205_220_0,
    i_8_205_233_0, i_8_205_237_0, i_8_205_238_0, i_8_205_255_0,
    i_8_205_304_0, i_8_205_371_0, i_8_205_374_0, i_8_205_380_0,
    i_8_205_382_0, i_8_205_385_0, i_8_205_423_0, i_8_205_437_0,
    i_8_205_453_0, i_8_205_477_0, i_8_205_478_0, i_8_205_481_0,
    i_8_205_482_0, i_8_205_484_0, i_8_205_485_0, i_8_205_498_0,
    i_8_205_499_0, i_8_205_505_0, i_8_205_523_0, i_8_205_526_0,
    i_8_205_532_0, i_8_205_564_0, i_8_205_634_0, i_8_205_661_0,
    i_8_205_684_0, i_8_205_703_0, i_8_205_757_0, i_8_205_759_0,
    i_8_205_760_0, i_8_205_761_0, i_8_205_767_0, i_8_205_780_0,
    i_8_205_811_0, i_8_205_823_0, i_8_205_830_0, i_8_205_869_0,
    i_8_205_892_0, i_8_205_904_0, i_8_205_1013_0, i_8_205_1030_0,
    i_8_205_1111_0, i_8_205_1112_0, i_8_205_1135_0, i_8_205_1174_0,
    i_8_205_1282_0, i_8_205_1294_0, i_8_205_1309_0, i_8_205_1328_0,
    i_8_205_1363_0, i_8_205_1366_0, i_8_205_1398_0, i_8_205_1506_0,
    i_8_205_1522_0, i_8_205_1537_0, i_8_205_1552_0, i_8_205_1565_0,
    i_8_205_1577_0, i_8_205_1605_0, i_8_205_1676_0, i_8_205_1678_0,
    i_8_205_1711_0, i_8_205_1723_0, i_8_205_1729_0, i_8_205_1730_0,
    i_8_205_1749_0, i_8_205_1752_0, i_8_205_1760_0, i_8_205_1805_0,
    i_8_205_1807_0, i_8_205_1818_0, i_8_205_1855_0, i_8_205_1903_0,
    i_8_205_1920_0, i_8_205_1947_0, i_8_205_1980_0, i_8_205_2020_0,
    i_8_205_2037_0, i_8_205_2038_0, i_8_205_2070_0, i_8_205_2093_0,
    i_8_205_2109_0, i_8_205_2150_0, i_8_205_2170_0, i_8_205_2218_0,
    i_8_205_2224_0, i_8_205_2237_0, i_8_205_2271_0, i_8_205_2286_0;
  output o_8_205_0_0;
  assign o_8_205_0_0 = 0;
endmodule



// Benchmark "kernel_8_206" written by ABC on Sun Jul 19 10:06:38 2020

module kernel_8_206 ( 
    i_8_206_22_0, i_8_206_41_0, i_8_206_52_0, i_8_206_53_0, i_8_206_76_0,
    i_8_206_103_0, i_8_206_130_0, i_8_206_138_0, i_8_206_168_0,
    i_8_206_169_0, i_8_206_319_0, i_8_206_354_0, i_8_206_365_0,
    i_8_206_373_0, i_8_206_382_0, i_8_206_386_0, i_8_206_394_0,
    i_8_206_429_0, i_8_206_430_0, i_8_206_454_0, i_8_206_492_0,
    i_8_206_493_0, i_8_206_495_0, i_8_206_507_0, i_8_206_538_0,
    i_8_206_544_0, i_8_206_556_0, i_8_206_565_0, i_8_206_610_0,
    i_8_206_637_0, i_8_206_679_0, i_8_206_694_0, i_8_206_724_0,
    i_8_206_747_0, i_8_206_766_0, i_8_206_823_0, i_8_206_835_0,
    i_8_206_847_0, i_8_206_962_0, i_8_206_970_0, i_8_206_1052_0,
    i_8_206_1065_0, i_8_206_1114_0, i_8_206_1115_0, i_8_206_1254_0,
    i_8_206_1257_0, i_8_206_1264_0, i_8_206_1265_0, i_8_206_1283_0,
    i_8_206_1315_0, i_8_206_1318_0, i_8_206_1354_0, i_8_206_1362_0,
    i_8_206_1363_0, i_8_206_1381_0, i_8_206_1384_0, i_8_206_1410_0,
    i_8_206_1413_0, i_8_206_1440_0, i_8_206_1455_0, i_8_206_1465_0,
    i_8_206_1467_0, i_8_206_1539_0, i_8_206_1542_0, i_8_206_1545_0,
    i_8_206_1553_0, i_8_206_1583_0, i_8_206_1669_0, i_8_206_1672_0,
    i_8_206_1687_0, i_8_206_1699_0, i_8_206_1731_0, i_8_206_1750_0,
    i_8_206_1801_0, i_8_206_1819_0, i_8_206_1823_0, i_8_206_1826_0,
    i_8_206_1850_0, i_8_206_1855_0, i_8_206_1859_0, i_8_206_1883_0,
    i_8_206_1972_0, i_8_206_1980_0, i_8_206_1986_0, i_8_206_2023_0,
    i_8_206_2073_0, i_8_206_2083_0, i_8_206_2126_0, i_8_206_2138_0,
    i_8_206_2146_0, i_8_206_2147_0, i_8_206_2191_0, i_8_206_2193_0,
    i_8_206_2224_0, i_8_206_2227_0, i_8_206_2243_0, i_8_206_2262_0,
    i_8_206_2278_0, i_8_206_2289_0, i_8_206_2292_0,
    o_8_206_0_0  );
  input  i_8_206_22_0, i_8_206_41_0, i_8_206_52_0, i_8_206_53_0,
    i_8_206_76_0, i_8_206_103_0, i_8_206_130_0, i_8_206_138_0,
    i_8_206_168_0, i_8_206_169_0, i_8_206_319_0, i_8_206_354_0,
    i_8_206_365_0, i_8_206_373_0, i_8_206_382_0, i_8_206_386_0,
    i_8_206_394_0, i_8_206_429_0, i_8_206_430_0, i_8_206_454_0,
    i_8_206_492_0, i_8_206_493_0, i_8_206_495_0, i_8_206_507_0,
    i_8_206_538_0, i_8_206_544_0, i_8_206_556_0, i_8_206_565_0,
    i_8_206_610_0, i_8_206_637_0, i_8_206_679_0, i_8_206_694_0,
    i_8_206_724_0, i_8_206_747_0, i_8_206_766_0, i_8_206_823_0,
    i_8_206_835_0, i_8_206_847_0, i_8_206_962_0, i_8_206_970_0,
    i_8_206_1052_0, i_8_206_1065_0, i_8_206_1114_0, i_8_206_1115_0,
    i_8_206_1254_0, i_8_206_1257_0, i_8_206_1264_0, i_8_206_1265_0,
    i_8_206_1283_0, i_8_206_1315_0, i_8_206_1318_0, i_8_206_1354_0,
    i_8_206_1362_0, i_8_206_1363_0, i_8_206_1381_0, i_8_206_1384_0,
    i_8_206_1410_0, i_8_206_1413_0, i_8_206_1440_0, i_8_206_1455_0,
    i_8_206_1465_0, i_8_206_1467_0, i_8_206_1539_0, i_8_206_1542_0,
    i_8_206_1545_0, i_8_206_1553_0, i_8_206_1583_0, i_8_206_1669_0,
    i_8_206_1672_0, i_8_206_1687_0, i_8_206_1699_0, i_8_206_1731_0,
    i_8_206_1750_0, i_8_206_1801_0, i_8_206_1819_0, i_8_206_1823_0,
    i_8_206_1826_0, i_8_206_1850_0, i_8_206_1855_0, i_8_206_1859_0,
    i_8_206_1883_0, i_8_206_1972_0, i_8_206_1980_0, i_8_206_1986_0,
    i_8_206_2023_0, i_8_206_2073_0, i_8_206_2083_0, i_8_206_2126_0,
    i_8_206_2138_0, i_8_206_2146_0, i_8_206_2147_0, i_8_206_2191_0,
    i_8_206_2193_0, i_8_206_2224_0, i_8_206_2227_0, i_8_206_2243_0,
    i_8_206_2262_0, i_8_206_2278_0, i_8_206_2289_0, i_8_206_2292_0;
  output o_8_206_0_0;
  assign o_8_206_0_0 = 0;
endmodule



// Benchmark "kernel_8_207" written by ABC on Sun Jul 19 10:06:39 2020

module kernel_8_207 ( 
    i_8_207_18_0, i_8_207_37_0, i_8_207_39_0, i_8_207_49_0, i_8_207_63_0,
    i_8_207_81_0, i_8_207_102_0, i_8_207_147_0, i_8_207_175_0,
    i_8_207_189_0, i_8_207_198_0, i_8_207_220_0, i_8_207_252_0,
    i_8_207_261_0, i_8_207_270_0, i_8_207_297_0, i_8_207_302_0,
    i_8_207_306_0, i_8_207_363_0, i_8_207_426_0, i_8_207_489_0,
    i_8_207_531_0, i_8_207_534_0, i_8_207_539_0, i_8_207_552_0,
    i_8_207_568_0, i_8_207_634_0, i_8_207_639_0, i_8_207_648_0,
    i_8_207_651_0, i_8_207_666_0, i_8_207_674_0, i_8_207_679_0,
    i_8_207_697_0, i_8_207_712_0, i_8_207_748_0, i_8_207_823_0,
    i_8_207_841_0, i_8_207_844_0, i_8_207_862_0, i_8_207_865_0,
    i_8_207_891_0, i_8_207_963_0, i_8_207_966_0, i_8_207_1080_0,
    i_8_207_1098_0, i_8_207_1128_0, i_8_207_1133_0, i_8_207_1170_0,
    i_8_207_1171_0, i_8_207_1179_0, i_8_207_1224_0, i_8_207_1227_0,
    i_8_207_1233_0, i_8_207_1236_0, i_8_207_1237_0, i_8_207_1263_0,
    i_8_207_1281_0, i_8_207_1297_0, i_8_207_1326_0, i_8_207_1377_0,
    i_8_207_1381_0, i_8_207_1386_0, i_8_207_1395_0, i_8_207_1431_0,
    i_8_207_1458_0, i_8_207_1506_0, i_8_207_1534_0, i_8_207_1560_0,
    i_8_207_1630_0, i_8_207_1639_0, i_8_207_1647_0, i_8_207_1650_0,
    i_8_207_1651_0, i_8_207_1674_0, i_8_207_1696_0, i_8_207_1754_0,
    i_8_207_1764_0, i_8_207_1767_0, i_8_207_1803_0, i_8_207_1804_0,
    i_8_207_1818_0, i_8_207_1864_0, i_8_207_1866_0, i_8_207_1910_0,
    i_8_207_1918_0, i_8_207_1927_0, i_8_207_1947_0, i_8_207_1966_0,
    i_8_207_1988_0, i_8_207_2034_0, i_8_207_2043_0, i_8_207_2062_0,
    i_8_207_2142_0, i_8_207_2146_0, i_8_207_2169_0, i_8_207_2177_0,
    i_8_207_2232_0, i_8_207_2268_0, i_8_207_2289_0,
    o_8_207_0_0  );
  input  i_8_207_18_0, i_8_207_37_0, i_8_207_39_0, i_8_207_49_0,
    i_8_207_63_0, i_8_207_81_0, i_8_207_102_0, i_8_207_147_0,
    i_8_207_175_0, i_8_207_189_0, i_8_207_198_0, i_8_207_220_0,
    i_8_207_252_0, i_8_207_261_0, i_8_207_270_0, i_8_207_297_0,
    i_8_207_302_0, i_8_207_306_0, i_8_207_363_0, i_8_207_426_0,
    i_8_207_489_0, i_8_207_531_0, i_8_207_534_0, i_8_207_539_0,
    i_8_207_552_0, i_8_207_568_0, i_8_207_634_0, i_8_207_639_0,
    i_8_207_648_0, i_8_207_651_0, i_8_207_666_0, i_8_207_674_0,
    i_8_207_679_0, i_8_207_697_0, i_8_207_712_0, i_8_207_748_0,
    i_8_207_823_0, i_8_207_841_0, i_8_207_844_0, i_8_207_862_0,
    i_8_207_865_0, i_8_207_891_0, i_8_207_963_0, i_8_207_966_0,
    i_8_207_1080_0, i_8_207_1098_0, i_8_207_1128_0, i_8_207_1133_0,
    i_8_207_1170_0, i_8_207_1171_0, i_8_207_1179_0, i_8_207_1224_0,
    i_8_207_1227_0, i_8_207_1233_0, i_8_207_1236_0, i_8_207_1237_0,
    i_8_207_1263_0, i_8_207_1281_0, i_8_207_1297_0, i_8_207_1326_0,
    i_8_207_1377_0, i_8_207_1381_0, i_8_207_1386_0, i_8_207_1395_0,
    i_8_207_1431_0, i_8_207_1458_0, i_8_207_1506_0, i_8_207_1534_0,
    i_8_207_1560_0, i_8_207_1630_0, i_8_207_1639_0, i_8_207_1647_0,
    i_8_207_1650_0, i_8_207_1651_0, i_8_207_1674_0, i_8_207_1696_0,
    i_8_207_1754_0, i_8_207_1764_0, i_8_207_1767_0, i_8_207_1803_0,
    i_8_207_1804_0, i_8_207_1818_0, i_8_207_1864_0, i_8_207_1866_0,
    i_8_207_1910_0, i_8_207_1918_0, i_8_207_1927_0, i_8_207_1947_0,
    i_8_207_1966_0, i_8_207_1988_0, i_8_207_2034_0, i_8_207_2043_0,
    i_8_207_2062_0, i_8_207_2142_0, i_8_207_2146_0, i_8_207_2169_0,
    i_8_207_2177_0, i_8_207_2232_0, i_8_207_2268_0, i_8_207_2289_0;
  output o_8_207_0_0;
  assign o_8_207_0_0 = 0;
endmodule



// Benchmark "kernel_8_208" written by ABC on Sun Jul 19 10:06:40 2020

module kernel_8_208 ( 
    i_8_208_7_0, i_8_208_26_0, i_8_208_88_0, i_8_208_179_0, i_8_208_219_0,
    i_8_208_232_0, i_8_208_240_0, i_8_208_250_0, i_8_208_266_0,
    i_8_208_287_0, i_8_208_292_0, i_8_208_332_0, i_8_208_348_0,
    i_8_208_349_0, i_8_208_386_0, i_8_208_463_0, i_8_208_466_0,
    i_8_208_467_0, i_8_208_502_0, i_8_208_520_0, i_8_208_526_0,
    i_8_208_527_0, i_8_208_556_0, i_8_208_594_0, i_8_208_610_0,
    i_8_208_627_0, i_8_208_656_0, i_8_208_662_0, i_8_208_672_0,
    i_8_208_673_0, i_8_208_698_0, i_8_208_717_0, i_8_208_718_0,
    i_8_208_754_0, i_8_208_782_0, i_8_208_798_0, i_8_208_799_0,
    i_8_208_808_0, i_8_208_843_0, i_8_208_879_0, i_8_208_926_0,
    i_8_208_992_0, i_8_208_994_0, i_8_208_995_0, i_8_208_997_0,
    i_8_208_998_0, i_8_208_1060_0, i_8_208_1077_0, i_8_208_1093_0,
    i_8_208_1139_0, i_8_208_1194_0, i_8_208_1205_0, i_8_208_1222_0,
    i_8_208_1258_0, i_8_208_1285_0, i_8_208_1286_0, i_8_208_1308_0,
    i_8_208_1316_0, i_8_208_1342_0, i_8_208_1357_0, i_8_208_1457_0,
    i_8_208_1474_0, i_8_208_1509_0, i_8_208_1538_0, i_8_208_1545_0,
    i_8_208_1546_0, i_8_208_1553_0, i_8_208_1555_0, i_8_208_1599_0,
    i_8_208_1601_0, i_8_208_1610_0, i_8_208_1647_0, i_8_208_1727_0,
    i_8_208_1751_0, i_8_208_1770_0, i_8_208_1832_0, i_8_208_1852_0,
    i_8_208_1853_0, i_8_208_1870_0, i_8_208_1897_0, i_8_208_1898_0,
    i_8_208_1921_0, i_8_208_1922_0, i_8_208_1925_0, i_8_208_1969_0,
    i_8_208_2014_0, i_8_208_2032_0, i_8_208_2074_0, i_8_208_2078_0,
    i_8_208_2113_0, i_8_208_2122_0, i_8_208_2131_0, i_8_208_2132_0,
    i_8_208_2150_0, i_8_208_2183_0, i_8_208_2219_0, i_8_208_2238_0,
    i_8_208_2249_0, i_8_208_2275_0, i_8_208_2293_0,
    o_8_208_0_0  );
  input  i_8_208_7_0, i_8_208_26_0, i_8_208_88_0, i_8_208_179_0,
    i_8_208_219_0, i_8_208_232_0, i_8_208_240_0, i_8_208_250_0,
    i_8_208_266_0, i_8_208_287_0, i_8_208_292_0, i_8_208_332_0,
    i_8_208_348_0, i_8_208_349_0, i_8_208_386_0, i_8_208_463_0,
    i_8_208_466_0, i_8_208_467_0, i_8_208_502_0, i_8_208_520_0,
    i_8_208_526_0, i_8_208_527_0, i_8_208_556_0, i_8_208_594_0,
    i_8_208_610_0, i_8_208_627_0, i_8_208_656_0, i_8_208_662_0,
    i_8_208_672_0, i_8_208_673_0, i_8_208_698_0, i_8_208_717_0,
    i_8_208_718_0, i_8_208_754_0, i_8_208_782_0, i_8_208_798_0,
    i_8_208_799_0, i_8_208_808_0, i_8_208_843_0, i_8_208_879_0,
    i_8_208_926_0, i_8_208_992_0, i_8_208_994_0, i_8_208_995_0,
    i_8_208_997_0, i_8_208_998_0, i_8_208_1060_0, i_8_208_1077_0,
    i_8_208_1093_0, i_8_208_1139_0, i_8_208_1194_0, i_8_208_1205_0,
    i_8_208_1222_0, i_8_208_1258_0, i_8_208_1285_0, i_8_208_1286_0,
    i_8_208_1308_0, i_8_208_1316_0, i_8_208_1342_0, i_8_208_1357_0,
    i_8_208_1457_0, i_8_208_1474_0, i_8_208_1509_0, i_8_208_1538_0,
    i_8_208_1545_0, i_8_208_1546_0, i_8_208_1553_0, i_8_208_1555_0,
    i_8_208_1599_0, i_8_208_1601_0, i_8_208_1610_0, i_8_208_1647_0,
    i_8_208_1727_0, i_8_208_1751_0, i_8_208_1770_0, i_8_208_1832_0,
    i_8_208_1852_0, i_8_208_1853_0, i_8_208_1870_0, i_8_208_1897_0,
    i_8_208_1898_0, i_8_208_1921_0, i_8_208_1922_0, i_8_208_1925_0,
    i_8_208_1969_0, i_8_208_2014_0, i_8_208_2032_0, i_8_208_2074_0,
    i_8_208_2078_0, i_8_208_2113_0, i_8_208_2122_0, i_8_208_2131_0,
    i_8_208_2132_0, i_8_208_2150_0, i_8_208_2183_0, i_8_208_2219_0,
    i_8_208_2238_0, i_8_208_2249_0, i_8_208_2275_0, i_8_208_2293_0;
  output o_8_208_0_0;
  assign o_8_208_0_0 = 0;
endmodule



// Benchmark "kernel_8_209" written by ABC on Sun Jul 19 10:06:41 2020

module kernel_8_209 ( 
    i_8_209_33_0, i_8_209_52_0, i_8_209_155_0, i_8_209_221_0,
    i_8_209_256_0, i_8_209_289_0, i_8_209_297_0, i_8_209_298_0,
    i_8_209_342_0, i_8_209_343_0, i_8_209_369_0, i_8_209_370_0,
    i_8_209_371_0, i_8_209_378_0, i_8_209_379_0, i_8_209_388_0,
    i_8_209_389_0, i_8_209_415_0, i_8_209_441_0, i_8_209_453_0,
    i_8_209_459_0, i_8_209_460_0, i_8_209_461_0, i_8_209_472_0,
    i_8_209_544_0, i_8_209_549_0, i_8_209_604_0, i_8_209_609_0,
    i_8_209_610_0, i_8_209_613_0, i_8_209_625_0, i_8_209_711_0,
    i_8_209_712_0, i_8_209_715_0, i_8_209_756_0, i_8_209_782_0,
    i_8_209_783_0, i_8_209_792_0, i_8_209_793_0, i_8_209_846_0,
    i_8_209_867_0, i_8_209_998_0, i_8_209_1008_0, i_8_209_1013_0,
    i_8_209_1027_0, i_8_209_1117_0, i_8_209_1118_0, i_8_209_1125_0,
    i_8_209_1128_0, i_8_209_1130_0, i_8_209_1156_0, i_8_209_1233_0,
    i_8_209_1246_0, i_8_209_1249_0, i_8_209_1324_0, i_8_209_1333_0,
    i_8_209_1343_0, i_8_209_1419_0, i_8_209_1420_0, i_8_209_1421_0,
    i_8_209_1467_0, i_8_209_1488_0, i_8_209_1531_0, i_8_209_1532_0,
    i_8_209_1537_0, i_8_209_1539_0, i_8_209_1540_0, i_8_209_1565_0,
    i_8_209_1579_0, i_8_209_1594_0, i_8_209_1595_0, i_8_209_1609_0,
    i_8_209_1611_0, i_8_209_1649_0, i_8_209_1676_0, i_8_209_1731_0,
    i_8_209_1738_0, i_8_209_1750_0, i_8_209_1783_0, i_8_209_1793_0,
    i_8_209_1801_0, i_8_209_1802_0, i_8_209_1864_0, i_8_209_1866_0,
    i_8_209_1869_0, i_8_209_1885_0, i_8_209_1926_0, i_8_209_1947_0,
    i_8_209_1992_0, i_8_209_2124_0, i_8_209_2125_0, i_8_209_2136_0,
    i_8_209_2141_0, i_8_209_2179_0, i_8_209_2180_0, i_8_209_2187_0,
    i_8_209_2188_0, i_8_209_2273_0, i_8_209_2287_0, i_8_209_2298_0,
    o_8_209_0_0  );
  input  i_8_209_33_0, i_8_209_52_0, i_8_209_155_0, i_8_209_221_0,
    i_8_209_256_0, i_8_209_289_0, i_8_209_297_0, i_8_209_298_0,
    i_8_209_342_0, i_8_209_343_0, i_8_209_369_0, i_8_209_370_0,
    i_8_209_371_0, i_8_209_378_0, i_8_209_379_0, i_8_209_388_0,
    i_8_209_389_0, i_8_209_415_0, i_8_209_441_0, i_8_209_453_0,
    i_8_209_459_0, i_8_209_460_0, i_8_209_461_0, i_8_209_472_0,
    i_8_209_544_0, i_8_209_549_0, i_8_209_604_0, i_8_209_609_0,
    i_8_209_610_0, i_8_209_613_0, i_8_209_625_0, i_8_209_711_0,
    i_8_209_712_0, i_8_209_715_0, i_8_209_756_0, i_8_209_782_0,
    i_8_209_783_0, i_8_209_792_0, i_8_209_793_0, i_8_209_846_0,
    i_8_209_867_0, i_8_209_998_0, i_8_209_1008_0, i_8_209_1013_0,
    i_8_209_1027_0, i_8_209_1117_0, i_8_209_1118_0, i_8_209_1125_0,
    i_8_209_1128_0, i_8_209_1130_0, i_8_209_1156_0, i_8_209_1233_0,
    i_8_209_1246_0, i_8_209_1249_0, i_8_209_1324_0, i_8_209_1333_0,
    i_8_209_1343_0, i_8_209_1419_0, i_8_209_1420_0, i_8_209_1421_0,
    i_8_209_1467_0, i_8_209_1488_0, i_8_209_1531_0, i_8_209_1532_0,
    i_8_209_1537_0, i_8_209_1539_0, i_8_209_1540_0, i_8_209_1565_0,
    i_8_209_1579_0, i_8_209_1594_0, i_8_209_1595_0, i_8_209_1609_0,
    i_8_209_1611_0, i_8_209_1649_0, i_8_209_1676_0, i_8_209_1731_0,
    i_8_209_1738_0, i_8_209_1750_0, i_8_209_1783_0, i_8_209_1793_0,
    i_8_209_1801_0, i_8_209_1802_0, i_8_209_1864_0, i_8_209_1866_0,
    i_8_209_1869_0, i_8_209_1885_0, i_8_209_1926_0, i_8_209_1947_0,
    i_8_209_1992_0, i_8_209_2124_0, i_8_209_2125_0, i_8_209_2136_0,
    i_8_209_2141_0, i_8_209_2179_0, i_8_209_2180_0, i_8_209_2187_0,
    i_8_209_2188_0, i_8_209_2273_0, i_8_209_2287_0, i_8_209_2298_0;
  output o_8_209_0_0;
  assign o_8_209_0_0 = 0;
endmodule



// Benchmark "kernel_8_210" written by ABC on Sun Jul 19 10:06:41 2020

module kernel_8_210 ( 
    i_8_210_32_0, i_8_210_47_0, i_8_210_49_0, i_8_210_65_0, i_8_210_91_0,
    i_8_210_92_0, i_8_210_103_0, i_8_210_236_0, i_8_210_320_0,
    i_8_210_326_0, i_8_210_362_0, i_8_210_380_0, i_8_210_383_0,
    i_8_210_388_0, i_8_210_417_0, i_8_210_424_0, i_8_210_452_0,
    i_8_210_490_0, i_8_210_493_0, i_8_210_512_0, i_8_210_578_0,
    i_8_210_604_0, i_8_210_635_0, i_8_210_640_0, i_8_210_658_0,
    i_8_210_668_0, i_8_210_676_0, i_8_210_677_0, i_8_210_686_0,
    i_8_210_701_0, i_8_210_703_0, i_8_210_705_0, i_8_210_731_0,
    i_8_210_767_0, i_8_210_778_0, i_8_210_841_0, i_8_210_844_0,
    i_8_210_929_0, i_8_210_955_0, i_8_210_967_0, i_8_210_968_0,
    i_8_210_1057_0, i_8_210_1112_0, i_8_210_1226_0, i_8_210_1261_0,
    i_8_210_1280_0, i_8_210_1316_0, i_8_210_1334_0, i_8_210_1352_0,
    i_8_210_1404_0, i_8_210_1442_0, i_8_210_1456_0, i_8_210_1468_0,
    i_8_210_1469_0, i_8_210_1473_0, i_8_210_1514_0, i_8_210_1530_0,
    i_8_210_1559_0, i_8_210_1604_0, i_8_210_1607_0, i_8_210_1612_0,
    i_8_210_1621_0, i_8_210_1622_0, i_8_210_1631_0, i_8_210_1648_0,
    i_8_210_1669_0, i_8_210_1678_0, i_8_210_1680_0, i_8_210_1684_0,
    i_8_210_1685_0, i_8_210_1693_0, i_8_210_1724_0, i_8_210_1730_0,
    i_8_210_1757_0, i_8_210_1768_0, i_8_210_1778_0, i_8_210_1783_0,
    i_8_210_1784_0, i_8_210_1818_0, i_8_210_1825_0, i_8_210_1864_0,
    i_8_210_1882_0, i_8_210_1946_0, i_8_210_1981_0, i_8_210_2000_0,
    i_8_210_2071_0, i_8_210_2075_0, i_8_210_2107_0, i_8_210_2133_0,
    i_8_210_2134_0, i_8_210_2147_0, i_8_210_2154_0, i_8_210_2156_0,
    i_8_210_2197_0, i_8_210_2198_0, i_8_210_2206_0, i_8_210_2224_0,
    i_8_210_2233_0, i_8_210_2260_0, i_8_210_2273_0,
    o_8_210_0_0  );
  input  i_8_210_32_0, i_8_210_47_0, i_8_210_49_0, i_8_210_65_0,
    i_8_210_91_0, i_8_210_92_0, i_8_210_103_0, i_8_210_236_0,
    i_8_210_320_0, i_8_210_326_0, i_8_210_362_0, i_8_210_380_0,
    i_8_210_383_0, i_8_210_388_0, i_8_210_417_0, i_8_210_424_0,
    i_8_210_452_0, i_8_210_490_0, i_8_210_493_0, i_8_210_512_0,
    i_8_210_578_0, i_8_210_604_0, i_8_210_635_0, i_8_210_640_0,
    i_8_210_658_0, i_8_210_668_0, i_8_210_676_0, i_8_210_677_0,
    i_8_210_686_0, i_8_210_701_0, i_8_210_703_0, i_8_210_705_0,
    i_8_210_731_0, i_8_210_767_0, i_8_210_778_0, i_8_210_841_0,
    i_8_210_844_0, i_8_210_929_0, i_8_210_955_0, i_8_210_967_0,
    i_8_210_968_0, i_8_210_1057_0, i_8_210_1112_0, i_8_210_1226_0,
    i_8_210_1261_0, i_8_210_1280_0, i_8_210_1316_0, i_8_210_1334_0,
    i_8_210_1352_0, i_8_210_1404_0, i_8_210_1442_0, i_8_210_1456_0,
    i_8_210_1468_0, i_8_210_1469_0, i_8_210_1473_0, i_8_210_1514_0,
    i_8_210_1530_0, i_8_210_1559_0, i_8_210_1604_0, i_8_210_1607_0,
    i_8_210_1612_0, i_8_210_1621_0, i_8_210_1622_0, i_8_210_1631_0,
    i_8_210_1648_0, i_8_210_1669_0, i_8_210_1678_0, i_8_210_1680_0,
    i_8_210_1684_0, i_8_210_1685_0, i_8_210_1693_0, i_8_210_1724_0,
    i_8_210_1730_0, i_8_210_1757_0, i_8_210_1768_0, i_8_210_1778_0,
    i_8_210_1783_0, i_8_210_1784_0, i_8_210_1818_0, i_8_210_1825_0,
    i_8_210_1864_0, i_8_210_1882_0, i_8_210_1946_0, i_8_210_1981_0,
    i_8_210_2000_0, i_8_210_2071_0, i_8_210_2075_0, i_8_210_2107_0,
    i_8_210_2133_0, i_8_210_2134_0, i_8_210_2147_0, i_8_210_2154_0,
    i_8_210_2156_0, i_8_210_2197_0, i_8_210_2198_0, i_8_210_2206_0,
    i_8_210_2224_0, i_8_210_2233_0, i_8_210_2260_0, i_8_210_2273_0;
  output o_8_210_0_0;
  assign o_8_210_0_0 = 0;
endmodule



// Benchmark "kernel_8_211" written by ABC on Sun Jul 19 10:06:42 2020

module kernel_8_211 ( 
    i_8_211_13_0, i_8_211_21_0, i_8_211_28_0, i_8_211_41_0, i_8_211_55_0,
    i_8_211_58_0, i_8_211_72_0, i_8_211_169_0, i_8_211_172_0,
    i_8_211_199_0, i_8_211_221_0, i_8_211_226_0, i_8_211_253_0,
    i_8_211_304_0, i_8_211_415_0, i_8_211_416_0, i_8_211_419_0,
    i_8_211_451_0, i_8_211_489_0, i_8_211_505_0, i_8_211_506_0,
    i_8_211_533_0, i_8_211_549_0, i_8_211_572_0, i_8_211_595_0,
    i_8_211_598_0, i_8_211_602_0, i_8_211_610_0, i_8_211_624_0,
    i_8_211_626_0, i_8_211_630_0, i_8_211_662_0, i_8_211_675_0,
    i_8_211_689_0, i_8_211_693_0, i_8_211_712_0, i_8_211_730_0,
    i_8_211_775_0, i_8_211_841_0, i_8_211_850_0, i_8_211_866_0,
    i_8_211_877_0, i_8_211_980_0, i_8_211_1073_0, i_8_211_1107_0,
    i_8_211_1135_0, i_8_211_1143_0, i_8_211_1199_0, i_8_211_1234_0,
    i_8_211_1260_0, i_8_211_1270_0, i_8_211_1278_0, i_8_211_1279_0,
    i_8_211_1282_0, i_8_211_1286_0, i_8_211_1298_0, i_8_211_1316_0,
    i_8_211_1387_0, i_8_211_1407_0, i_8_211_1408_0, i_8_211_1424_0,
    i_8_211_1438_0, i_8_211_1452_0, i_8_211_1470_0, i_8_211_1478_0,
    i_8_211_1481_0, i_8_211_1558_0, i_8_211_1607_0, i_8_211_1631_0,
    i_8_211_1632_0, i_8_211_1659_0, i_8_211_1684_0, i_8_211_1710_0,
    i_8_211_1747_0, i_8_211_1748_0, i_8_211_1766_0, i_8_211_1820_0,
    i_8_211_1821_0, i_8_211_1823_0, i_8_211_1854_0, i_8_211_1873_0,
    i_8_211_1882_0, i_8_211_1883_0, i_8_211_1885_0, i_8_211_1962_0,
    i_8_211_1966_0, i_8_211_1980_0, i_8_211_2017_0, i_8_211_2044_0,
    i_8_211_2088_0, i_8_211_2125_0, i_8_211_2135_0, i_8_211_2140_0,
    i_8_211_2151_0, i_8_211_2169_0, i_8_211_2232_0, i_8_211_2234_0,
    i_8_211_2261_0, i_8_211_2273_0, i_8_211_2296_0,
    o_8_211_0_0  );
  input  i_8_211_13_0, i_8_211_21_0, i_8_211_28_0, i_8_211_41_0,
    i_8_211_55_0, i_8_211_58_0, i_8_211_72_0, i_8_211_169_0, i_8_211_172_0,
    i_8_211_199_0, i_8_211_221_0, i_8_211_226_0, i_8_211_253_0,
    i_8_211_304_0, i_8_211_415_0, i_8_211_416_0, i_8_211_419_0,
    i_8_211_451_0, i_8_211_489_0, i_8_211_505_0, i_8_211_506_0,
    i_8_211_533_0, i_8_211_549_0, i_8_211_572_0, i_8_211_595_0,
    i_8_211_598_0, i_8_211_602_0, i_8_211_610_0, i_8_211_624_0,
    i_8_211_626_0, i_8_211_630_0, i_8_211_662_0, i_8_211_675_0,
    i_8_211_689_0, i_8_211_693_0, i_8_211_712_0, i_8_211_730_0,
    i_8_211_775_0, i_8_211_841_0, i_8_211_850_0, i_8_211_866_0,
    i_8_211_877_0, i_8_211_980_0, i_8_211_1073_0, i_8_211_1107_0,
    i_8_211_1135_0, i_8_211_1143_0, i_8_211_1199_0, i_8_211_1234_0,
    i_8_211_1260_0, i_8_211_1270_0, i_8_211_1278_0, i_8_211_1279_0,
    i_8_211_1282_0, i_8_211_1286_0, i_8_211_1298_0, i_8_211_1316_0,
    i_8_211_1387_0, i_8_211_1407_0, i_8_211_1408_0, i_8_211_1424_0,
    i_8_211_1438_0, i_8_211_1452_0, i_8_211_1470_0, i_8_211_1478_0,
    i_8_211_1481_0, i_8_211_1558_0, i_8_211_1607_0, i_8_211_1631_0,
    i_8_211_1632_0, i_8_211_1659_0, i_8_211_1684_0, i_8_211_1710_0,
    i_8_211_1747_0, i_8_211_1748_0, i_8_211_1766_0, i_8_211_1820_0,
    i_8_211_1821_0, i_8_211_1823_0, i_8_211_1854_0, i_8_211_1873_0,
    i_8_211_1882_0, i_8_211_1883_0, i_8_211_1885_0, i_8_211_1962_0,
    i_8_211_1966_0, i_8_211_1980_0, i_8_211_2017_0, i_8_211_2044_0,
    i_8_211_2088_0, i_8_211_2125_0, i_8_211_2135_0, i_8_211_2140_0,
    i_8_211_2151_0, i_8_211_2169_0, i_8_211_2232_0, i_8_211_2234_0,
    i_8_211_2261_0, i_8_211_2273_0, i_8_211_2296_0;
  output o_8_211_0_0;
  assign o_8_211_0_0 = 0;
endmodule



// Benchmark "kernel_8_212" written by ABC on Sun Jul 19 10:06:44 2020

module kernel_8_212 ( 
    i_8_212_13_0, i_8_212_16_0, i_8_212_31_0, i_8_212_57_0, i_8_212_66_0,
    i_8_212_75_0, i_8_212_94_0, i_8_212_98_0, i_8_212_124_0, i_8_212_188_0,
    i_8_212_229_0, i_8_212_232_0, i_8_212_304_0, i_8_212_339_0,
    i_8_212_360_0, i_8_212_367_0, i_8_212_384_0, i_8_212_385_0,
    i_8_212_399_0, i_8_212_400_0, i_8_212_420_0, i_8_212_466_0,
    i_8_212_525_0, i_8_212_574_0, i_8_212_591_0, i_8_212_592_0,
    i_8_212_608_0, i_8_212_655_0, i_8_212_678_0, i_8_212_681_0,
    i_8_212_750_0, i_8_212_817_0, i_8_212_843_0, i_8_212_844_0,
    i_8_212_852_0, i_8_212_853_0, i_8_212_861_0, i_8_212_879_0,
    i_8_212_883_0, i_8_212_961_0, i_8_212_967_0, i_8_212_1012_0,
    i_8_212_1128_0, i_8_212_1140_0, i_8_212_1141_0, i_8_212_1149_0,
    i_8_212_1150_0, i_8_212_1158_0, i_8_212_1186_0, i_8_212_1228_0,
    i_8_212_1231_0, i_8_212_1236_0, i_8_212_1263_0, i_8_212_1302_0,
    i_8_212_1317_0, i_8_212_1320_0, i_8_212_1321_0, i_8_212_1330_0,
    i_8_212_1331_0, i_8_212_1482_0, i_8_212_1553_0, i_8_212_1561_0,
    i_8_212_1606_0, i_8_212_1608_0, i_8_212_1636_0, i_8_212_1677_0,
    i_8_212_1680_0, i_8_212_1716_0, i_8_212_1722_0, i_8_212_1752_0,
    i_8_212_1763_0, i_8_212_1789_0, i_8_212_1795_0, i_8_212_1813_0,
    i_8_212_1816_0, i_8_212_1818_0, i_8_212_1860_0, i_8_212_1922_0,
    i_8_212_1951_0, i_8_212_1960_0, i_8_212_1995_0, i_8_212_2004_0,
    i_8_212_2058_0, i_8_212_2076_0, i_8_212_2094_0, i_8_212_2109_0,
    i_8_212_2136_0, i_8_212_2137_0, i_8_212_2142_0, i_8_212_2145_0,
    i_8_212_2147_0, i_8_212_2158_0, i_8_212_2176_0, i_8_212_2190_0,
    i_8_212_2238_0, i_8_212_2239_0, i_8_212_2244_0, i_8_212_2246_0,
    i_8_212_2248_0, i_8_212_2266_0,
    o_8_212_0_0  );
  input  i_8_212_13_0, i_8_212_16_0, i_8_212_31_0, i_8_212_57_0,
    i_8_212_66_0, i_8_212_75_0, i_8_212_94_0, i_8_212_98_0, i_8_212_124_0,
    i_8_212_188_0, i_8_212_229_0, i_8_212_232_0, i_8_212_304_0,
    i_8_212_339_0, i_8_212_360_0, i_8_212_367_0, i_8_212_384_0,
    i_8_212_385_0, i_8_212_399_0, i_8_212_400_0, i_8_212_420_0,
    i_8_212_466_0, i_8_212_525_0, i_8_212_574_0, i_8_212_591_0,
    i_8_212_592_0, i_8_212_608_0, i_8_212_655_0, i_8_212_678_0,
    i_8_212_681_0, i_8_212_750_0, i_8_212_817_0, i_8_212_843_0,
    i_8_212_844_0, i_8_212_852_0, i_8_212_853_0, i_8_212_861_0,
    i_8_212_879_0, i_8_212_883_0, i_8_212_961_0, i_8_212_967_0,
    i_8_212_1012_0, i_8_212_1128_0, i_8_212_1140_0, i_8_212_1141_0,
    i_8_212_1149_0, i_8_212_1150_0, i_8_212_1158_0, i_8_212_1186_0,
    i_8_212_1228_0, i_8_212_1231_0, i_8_212_1236_0, i_8_212_1263_0,
    i_8_212_1302_0, i_8_212_1317_0, i_8_212_1320_0, i_8_212_1321_0,
    i_8_212_1330_0, i_8_212_1331_0, i_8_212_1482_0, i_8_212_1553_0,
    i_8_212_1561_0, i_8_212_1606_0, i_8_212_1608_0, i_8_212_1636_0,
    i_8_212_1677_0, i_8_212_1680_0, i_8_212_1716_0, i_8_212_1722_0,
    i_8_212_1752_0, i_8_212_1763_0, i_8_212_1789_0, i_8_212_1795_0,
    i_8_212_1813_0, i_8_212_1816_0, i_8_212_1818_0, i_8_212_1860_0,
    i_8_212_1922_0, i_8_212_1951_0, i_8_212_1960_0, i_8_212_1995_0,
    i_8_212_2004_0, i_8_212_2058_0, i_8_212_2076_0, i_8_212_2094_0,
    i_8_212_2109_0, i_8_212_2136_0, i_8_212_2137_0, i_8_212_2142_0,
    i_8_212_2145_0, i_8_212_2147_0, i_8_212_2158_0, i_8_212_2176_0,
    i_8_212_2190_0, i_8_212_2238_0, i_8_212_2239_0, i_8_212_2244_0,
    i_8_212_2246_0, i_8_212_2248_0, i_8_212_2266_0;
  output o_8_212_0_0;
  assign o_8_212_0_0 = ~((~i_8_212_1561_0 & ((i_8_212_75_0 & ((i_8_212_591_0 & ~i_8_212_1331_0 & ~i_8_212_1606_0 & ~i_8_212_1816_0 & ~i_8_212_2058_0) | (~i_8_212_1150_0 & ~i_8_212_1186_0 & ~i_8_212_1677_0 & ~i_8_212_1716_0 & ~i_8_212_1752_0 & ~i_8_212_1763_0 & i_8_212_2137_0))) | (~i_8_212_232_0 & ~i_8_212_2266_0 & ((~i_8_212_57_0 & ~i_8_212_852_0 & ~i_8_212_1140_0 & ~i_8_212_1231_0 & ~i_8_212_1302_0 & ~i_8_212_2004_0 & ~i_8_212_2176_0 & ~i_8_212_2238_0) | (~i_8_212_399_0 & i_8_212_420_0 & ~i_8_212_2158_0 & i_8_212_2244_0))))) | (~i_8_212_98_0 & ((~i_8_212_304_0 & ~i_8_212_861_0 & i_8_212_967_0 & ~i_8_212_1636_0 & ~i_8_212_1763_0 & ~i_8_212_1951_0 & ~i_8_212_2058_0) | (~i_8_212_31_0 & ~i_8_212_57_0 & ~i_8_212_655_0 & ~i_8_212_843_0 & ~i_8_212_853_0 & ~i_8_212_1813_0 & ~i_8_212_1816_0 & ~i_8_212_2109_0))) | (~i_8_212_31_0 & ((~i_8_212_384_0 & ~i_8_212_655_0 & ~i_8_212_853_0 & ~i_8_212_1149_0 & ~i_8_212_1302_0 & ~i_8_212_1995_0) | (~i_8_212_385_0 & ~i_8_212_592_0 & i_8_212_655_0 & ~i_8_212_843_0 & ~i_8_212_1228_0 & ~i_8_212_1263_0 & ~i_8_212_2058_0 & ~i_8_212_2136_0))) | (~i_8_212_592_0 & ((i_8_212_367_0 & ((~i_8_212_678_0 & ~i_8_212_861_0 & i_8_212_1860_0 & ~i_8_212_2094_0 & ~i_8_212_2158_0) | (~i_8_212_57_0 & ~i_8_212_879_0 & ~i_8_212_1140_0 & i_8_212_1553_0 & ~i_8_212_1752_0 & ~i_8_212_2266_0))) | (~i_8_212_385_0 & ~i_8_212_574_0 & ~i_8_212_608_0 & ~i_8_212_843_0 & ~i_8_212_853_0 & ~i_8_212_1150_0 & ~i_8_212_1320_0))) | (~i_8_212_1951_0 & ((~i_8_212_57_0 & ((~i_8_212_420_0 & ~i_8_212_574_0 & ~i_8_212_681_0 & i_8_212_1228_0 & ~i_8_212_1636_0 & i_8_212_1813_0 & i_8_212_1922_0 & ~i_8_212_2058_0 & i_8_212_2137_0 & ~i_8_212_2158_0) | (~i_8_212_124_0 & ~i_8_212_853_0 & ~i_8_212_883_0 & ~i_8_212_1150_0 & ~i_8_212_1608_0 & ~i_8_212_1677_0 & ~i_8_212_2239_0))) | (~i_8_212_188_0 & ~i_8_212_304_0 & i_8_212_843_0 & ~i_8_212_1140_0 & ~i_8_212_1716_0 & ~i_8_212_1763_0 & ~i_8_212_1816_0 & ~i_8_212_2004_0 & ~i_8_212_2137_0))) | (~i_8_212_399_0 & ((~i_8_212_655_0 & ~i_8_212_853_0 & ~i_8_212_1012_0 & ~i_8_212_1482_0 & ~i_8_212_1606_0 & ~i_8_212_1752_0 & i_8_212_2145_0) | (~i_8_212_844_0 & ~i_8_212_1231_0 & i_8_212_1677_0 & ~i_8_212_1813_0 & ~i_8_212_2238_0 & ~i_8_212_2239_0))) | (~i_8_212_1140_0 & ((~i_8_212_400_0 & ((i_8_212_525_0 & ~i_8_212_853_0 & ~i_8_212_2145_0) | (~i_8_212_655_0 & ~i_8_212_961_0 & ~i_8_212_1606_0 & ~i_8_212_1608_0 & ~i_8_212_1922_0 & ~i_8_212_2158_0 & ~i_8_212_2248_0))) | (~i_8_212_124_0 & ~i_8_212_367_0 & ~i_8_212_420_0 & ~i_8_212_1141_0 & ~i_8_212_1608_0 & ~i_8_212_1716_0 & ~i_8_212_1763_0 & ~i_8_212_2137_0 & ~i_8_212_2147_0))) | (~i_8_212_1816_0 & ((~i_8_212_678_0 & ~i_8_212_1763_0 & ((~i_8_212_66_0 & ~i_8_212_124_0 & ~i_8_212_681_0 & ~i_8_212_883_0 & ~i_8_212_1150_0 & ~i_8_212_1553_0 & ~i_8_212_1608_0 & ~i_8_212_2004_0 & ~i_8_212_2058_0) | (~i_8_212_75_0 & ~i_8_212_339_0 & ~i_8_212_591_0 & ~i_8_212_655_0 & ~i_8_212_861_0 & ~i_8_212_1141_0 & ~i_8_212_1320_0 & ~i_8_212_2246_0))) | (~i_8_212_1302_0 & ~i_8_212_2136_0 & ((~i_8_212_384_0 & ~i_8_212_883_0 & ~i_8_212_961_0 & ~i_8_212_1149_0 & ~i_8_212_1158_0 & ~i_8_212_1818_0 & ~i_8_212_2158_0) | (~i_8_212_1231_0 & i_8_212_2109_0 & ~i_8_212_2266_0))))) | (~i_8_212_124_0 & ((~i_8_212_16_0 & ~i_8_212_1149_0 & i_8_212_1228_0 & ~i_8_212_1331_0 & ~i_8_212_1763_0 & ~i_8_212_1860_0 & i_8_212_2145_0 & ~i_8_212_2158_0) | (i_8_212_1331_0 & ~i_8_212_1813_0 & ~i_8_212_2266_0))) | (~i_8_212_681_0 & ((~i_8_212_655_0 & ~i_8_212_861_0 & ~i_8_212_1482_0 & ~i_8_212_1763_0 & ~i_8_212_2137_0 & i_8_212_2147_0) | (~i_8_212_360_0 & ~i_8_212_1141_0 & ~i_8_212_1228_0 & ~i_8_212_1606_0 & i_8_212_1636_0 & i_8_212_1752_0 & ~i_8_212_2058_0 & ~i_8_212_2244_0))) | (~i_8_212_1150_0 & ((~i_8_212_655_0 & ((~i_8_212_385_0 & i_8_212_1012_0) | (~i_8_212_750_0 & ~i_8_212_861_0 & ~i_8_212_1228_0 & i_8_212_1922_0 & ~i_8_212_2004_0))) | (~i_8_212_844_0 & ~i_8_212_1149_0 & ~i_8_212_1263_0 & ~i_8_212_1995_0 & ~i_8_212_2137_0 & ~i_8_212_2246_0))) | (i_8_212_1231_0 & i_8_212_1331_0 & i_8_212_1553_0 & ~i_8_212_1608_0 & ~i_8_212_2094_0) | (i_8_212_420_0 & i_8_212_655_0 & ~i_8_212_678_0 & i_8_212_1012_0 & ~i_8_212_1813_0 & i_8_212_1995_0 & ~i_8_212_2246_0));
endmodule



// Benchmark "kernel_8_213" written by ABC on Sun Jul 19 10:06:45 2020

module kernel_8_213 ( 
    i_8_213_9_0, i_8_213_18_0, i_8_213_37_0, i_8_213_73_0, i_8_213_102_0,
    i_8_213_135_0, i_8_213_183_0, i_8_213_225_0, i_8_213_226_0,
    i_8_213_252_0, i_8_213_255_0, i_8_213_259_0, i_8_213_279_0,
    i_8_213_321_0, i_8_213_364_0, i_8_213_365_0, i_8_213_370_0,
    i_8_213_399_0, i_8_213_495_0, i_8_213_499_0, i_8_213_534_0,
    i_8_213_540_0, i_8_213_567_0, i_8_213_570_0, i_8_213_594_0,
    i_8_213_604_0, i_8_213_639_0, i_8_213_659_0, i_8_213_660_0,
    i_8_213_675_0, i_8_213_678_0, i_8_213_777_0, i_8_213_783_0,
    i_8_213_810_0, i_8_213_841_0, i_8_213_864_0, i_8_213_868_0,
    i_8_213_891_0, i_8_213_937_0, i_8_213_954_0, i_8_213_966_0,
    i_8_213_969_0, i_8_213_975_0, i_8_213_1036_0, i_8_213_1107_0,
    i_8_213_1110_0, i_8_213_1111_0, i_8_213_1125_0, i_8_213_1138_0,
    i_8_213_1179_0, i_8_213_1197_0, i_8_213_1225_0, i_8_213_1236_0,
    i_8_213_1242_0, i_8_213_1246_0, i_8_213_1261_0, i_8_213_1263_0,
    i_8_213_1264_0, i_8_213_1314_0, i_8_213_1335_0, i_8_213_1338_0,
    i_8_213_1342_0, i_8_213_1344_0, i_8_213_1377_0, i_8_213_1422_0,
    i_8_213_1424_0, i_8_213_1434_0, i_8_213_1435_0, i_8_213_1467_0,
    i_8_213_1468_0, i_8_213_1476_0, i_8_213_1480_0, i_8_213_1512_0,
    i_8_213_1516_0, i_8_213_1524_0, i_8_213_1539_0, i_8_213_1542_0,
    i_8_213_1555_0, i_8_213_1557_0, i_8_213_1629_0, i_8_213_1651_0,
    i_8_213_1705_0, i_8_213_1753_0, i_8_213_1755_0, i_8_213_1758_0,
    i_8_213_1759_0, i_8_213_1767_0, i_8_213_1773_0, i_8_213_1776_0,
    i_8_213_1789_0, i_8_213_1790_0, i_8_213_1950_0, i_8_213_1989_0,
    i_8_213_1996_0, i_8_213_2133_0, i_8_213_2145_0, i_8_213_2196_0,
    i_8_213_2232_0, i_8_213_2233_0, i_8_213_2271_0,
    o_8_213_0_0  );
  input  i_8_213_9_0, i_8_213_18_0, i_8_213_37_0, i_8_213_73_0,
    i_8_213_102_0, i_8_213_135_0, i_8_213_183_0, i_8_213_225_0,
    i_8_213_226_0, i_8_213_252_0, i_8_213_255_0, i_8_213_259_0,
    i_8_213_279_0, i_8_213_321_0, i_8_213_364_0, i_8_213_365_0,
    i_8_213_370_0, i_8_213_399_0, i_8_213_495_0, i_8_213_499_0,
    i_8_213_534_0, i_8_213_540_0, i_8_213_567_0, i_8_213_570_0,
    i_8_213_594_0, i_8_213_604_0, i_8_213_639_0, i_8_213_659_0,
    i_8_213_660_0, i_8_213_675_0, i_8_213_678_0, i_8_213_777_0,
    i_8_213_783_0, i_8_213_810_0, i_8_213_841_0, i_8_213_864_0,
    i_8_213_868_0, i_8_213_891_0, i_8_213_937_0, i_8_213_954_0,
    i_8_213_966_0, i_8_213_969_0, i_8_213_975_0, i_8_213_1036_0,
    i_8_213_1107_0, i_8_213_1110_0, i_8_213_1111_0, i_8_213_1125_0,
    i_8_213_1138_0, i_8_213_1179_0, i_8_213_1197_0, i_8_213_1225_0,
    i_8_213_1236_0, i_8_213_1242_0, i_8_213_1246_0, i_8_213_1261_0,
    i_8_213_1263_0, i_8_213_1264_0, i_8_213_1314_0, i_8_213_1335_0,
    i_8_213_1338_0, i_8_213_1342_0, i_8_213_1344_0, i_8_213_1377_0,
    i_8_213_1422_0, i_8_213_1424_0, i_8_213_1434_0, i_8_213_1435_0,
    i_8_213_1467_0, i_8_213_1468_0, i_8_213_1476_0, i_8_213_1480_0,
    i_8_213_1512_0, i_8_213_1516_0, i_8_213_1524_0, i_8_213_1539_0,
    i_8_213_1542_0, i_8_213_1555_0, i_8_213_1557_0, i_8_213_1629_0,
    i_8_213_1651_0, i_8_213_1705_0, i_8_213_1753_0, i_8_213_1755_0,
    i_8_213_1758_0, i_8_213_1759_0, i_8_213_1767_0, i_8_213_1773_0,
    i_8_213_1776_0, i_8_213_1789_0, i_8_213_1790_0, i_8_213_1950_0,
    i_8_213_1989_0, i_8_213_1996_0, i_8_213_2133_0, i_8_213_2145_0,
    i_8_213_2196_0, i_8_213_2232_0, i_8_213_2233_0, i_8_213_2271_0;
  output o_8_213_0_0;
  assign o_8_213_0_0 = 0;
endmodule



// Benchmark "kernel_8_214" written by ABC on Sun Jul 19 10:06:47 2020

module kernel_8_214 ( 
    i_8_214_18_0, i_8_214_21_0, i_8_214_57_0, i_8_214_120_0, i_8_214_141_0,
    i_8_214_142_0, i_8_214_169_0, i_8_214_192_0, i_8_214_237_0,
    i_8_214_266_0, i_8_214_269_0, i_8_214_285_0, i_8_214_348_0,
    i_8_214_385_0, i_8_214_426_0, i_8_214_430_0, i_8_214_492_0,
    i_8_214_527_0, i_8_214_530_0, i_8_214_555_0, i_8_214_580_0,
    i_8_214_611_0, i_8_214_637_0, i_8_214_642_0, i_8_214_665_0,
    i_8_214_696_0, i_8_214_706_0, i_8_214_709_0, i_8_214_734_0,
    i_8_214_772_0, i_8_214_832_0, i_8_214_839_0, i_8_214_843_0,
    i_8_214_867_0, i_8_214_957_0, i_8_214_958_0, i_8_214_966_0,
    i_8_214_1041_0, i_8_214_1042_0, i_8_214_1072_0, i_8_214_1130_0,
    i_8_214_1146_0, i_8_214_1149_0, i_8_214_1160_0, i_8_214_1167_0,
    i_8_214_1182_0, i_8_214_1227_0, i_8_214_1237_0, i_8_214_1284_0,
    i_8_214_1285_0, i_8_214_1299_0, i_8_214_1318_0, i_8_214_1358_0,
    i_8_214_1362_0, i_8_214_1443_0, i_8_214_1447_0, i_8_214_1479_0,
    i_8_214_1480_0, i_8_214_1483_0, i_8_214_1488_0, i_8_214_1489_0,
    i_8_214_1490_0, i_8_214_1560_0, i_8_214_1565_0, i_8_214_1605_0,
    i_8_214_1608_0, i_8_214_1679_0, i_8_214_1686_0, i_8_214_1719_0,
    i_8_214_1725_0, i_8_214_1770_0, i_8_214_1785_0, i_8_214_1812_0,
    i_8_214_1824_0, i_8_214_1825_0, i_8_214_1947_0, i_8_214_1956_0,
    i_8_214_1959_0, i_8_214_1983_0, i_8_214_2056_0, i_8_214_2070_0,
    i_8_214_2074_0, i_8_214_2112_0, i_8_214_2113_0, i_8_214_2139_0,
    i_8_214_2140_0, i_8_214_2147_0, i_8_214_2154_0, i_8_214_2158_0,
    i_8_214_2193_0, i_8_214_2203_0, i_8_214_2227_0, i_8_214_2229_0,
    i_8_214_2232_0, i_8_214_2235_0, i_8_214_2239_0, i_8_214_2262_0,
    i_8_214_2263_0, i_8_214_2289_0, i_8_214_2292_0,
    o_8_214_0_0  );
  input  i_8_214_18_0, i_8_214_21_0, i_8_214_57_0, i_8_214_120_0,
    i_8_214_141_0, i_8_214_142_0, i_8_214_169_0, i_8_214_192_0,
    i_8_214_237_0, i_8_214_266_0, i_8_214_269_0, i_8_214_285_0,
    i_8_214_348_0, i_8_214_385_0, i_8_214_426_0, i_8_214_430_0,
    i_8_214_492_0, i_8_214_527_0, i_8_214_530_0, i_8_214_555_0,
    i_8_214_580_0, i_8_214_611_0, i_8_214_637_0, i_8_214_642_0,
    i_8_214_665_0, i_8_214_696_0, i_8_214_706_0, i_8_214_709_0,
    i_8_214_734_0, i_8_214_772_0, i_8_214_832_0, i_8_214_839_0,
    i_8_214_843_0, i_8_214_867_0, i_8_214_957_0, i_8_214_958_0,
    i_8_214_966_0, i_8_214_1041_0, i_8_214_1042_0, i_8_214_1072_0,
    i_8_214_1130_0, i_8_214_1146_0, i_8_214_1149_0, i_8_214_1160_0,
    i_8_214_1167_0, i_8_214_1182_0, i_8_214_1227_0, i_8_214_1237_0,
    i_8_214_1284_0, i_8_214_1285_0, i_8_214_1299_0, i_8_214_1318_0,
    i_8_214_1358_0, i_8_214_1362_0, i_8_214_1443_0, i_8_214_1447_0,
    i_8_214_1479_0, i_8_214_1480_0, i_8_214_1483_0, i_8_214_1488_0,
    i_8_214_1489_0, i_8_214_1490_0, i_8_214_1560_0, i_8_214_1565_0,
    i_8_214_1605_0, i_8_214_1608_0, i_8_214_1679_0, i_8_214_1686_0,
    i_8_214_1719_0, i_8_214_1725_0, i_8_214_1770_0, i_8_214_1785_0,
    i_8_214_1812_0, i_8_214_1824_0, i_8_214_1825_0, i_8_214_1947_0,
    i_8_214_1956_0, i_8_214_1959_0, i_8_214_1983_0, i_8_214_2056_0,
    i_8_214_2070_0, i_8_214_2074_0, i_8_214_2112_0, i_8_214_2113_0,
    i_8_214_2139_0, i_8_214_2140_0, i_8_214_2147_0, i_8_214_2154_0,
    i_8_214_2158_0, i_8_214_2193_0, i_8_214_2203_0, i_8_214_2227_0,
    i_8_214_2229_0, i_8_214_2232_0, i_8_214_2235_0, i_8_214_2239_0,
    i_8_214_2262_0, i_8_214_2263_0, i_8_214_2289_0, i_8_214_2292_0;
  output o_8_214_0_0;
  assign o_8_214_0_0 = ~((~i_8_214_2263_0 & ((i_8_214_57_0 & ((~i_8_214_18_0 & ~i_8_214_839_0 & ~i_8_214_957_0 & ~i_8_214_1284_0 & ~i_8_214_1824_0 & ~i_8_214_1825_0 & ~i_8_214_1947_0 & ~i_8_214_2158_0) | (~i_8_214_348_0 & ~i_8_214_1227_0 & ~i_8_214_1560_0 & ~i_8_214_1608_0 & ~i_8_214_2203_0 & ~i_8_214_2232_0 & ~i_8_214_2289_0))) | (~i_8_214_57_0 & ((~i_8_214_18_0 & ((i_8_214_142_0 & ~i_8_214_1146_0 & ~i_8_214_1362_0 & ~i_8_214_1812_0 & ~i_8_214_2113_0 & ~i_8_214_2158_0) | (~i_8_214_237_0 & i_8_214_426_0 & ~i_8_214_709_0 & ~i_8_214_1167_0 & ~i_8_214_1284_0 & ~i_8_214_1560_0 & ~i_8_214_1679_0 & ~i_8_214_2056_0 & ~i_8_214_2112_0 & ~i_8_214_2154_0 & ~i_8_214_2289_0))) | (i_8_214_21_0 & ~i_8_214_385_0 & ~i_8_214_580_0 & ~i_8_214_843_0 & ~i_8_214_958_0 & ~i_8_214_1149_0 & ~i_8_214_1318_0 & ~i_8_214_1447_0 & ~i_8_214_1785_0 & ~i_8_214_2227_0))) | (~i_8_214_1146_0 & ((i_8_214_192_0 & i_8_214_696_0 & ~i_8_214_1443_0 & ~i_8_214_1725_0 & ~i_8_214_1812_0 & ~i_8_214_2239_0) | (~i_8_214_1160_0 & i_8_214_1358_0 & ~i_8_214_1770_0 & ~i_8_214_2203_0 & ~i_8_214_2229_0 & ~i_8_214_2262_0 & ~i_8_214_2292_0))) | (~i_8_214_2112_0 & ((~i_8_214_839_0 & i_8_214_1237_0 & i_8_214_1358_0 & ~i_8_214_2262_0) | (~i_8_214_1237_0 & i_8_214_1488_0 & ~i_8_214_1560_0 & ~i_8_214_1679_0 & i_8_214_1785_0 & ~i_8_214_2292_0))))) | (~i_8_214_492_0 & ((~i_8_214_18_0 & ~i_8_214_2113_0 & ((~i_8_214_57_0 & ~i_8_214_430_0 & ~i_8_214_1146_0 & ~i_8_214_1149_0 & ~i_8_214_1227_0 & ~i_8_214_1605_0 & ~i_8_214_1947_0 & ~i_8_214_2056_0 & ~i_8_214_2112_0) | (~i_8_214_734_0 & ~i_8_214_1167_0 & ~i_8_214_1284_0 & i_8_214_1679_0 & ~i_8_214_2203_0 & ~i_8_214_2239_0 & ~i_8_214_2289_0))) | (~i_8_214_57_0 & i_8_214_611_0 & ~i_8_214_709_0 & ~i_8_214_1447_0 & ~i_8_214_1785_0 & ~i_8_214_2229_0))) | (~i_8_214_2113_0 & ((~i_8_214_18_0 & ~i_8_214_839_0 & ((~i_8_214_966_0 & ~i_8_214_1160_0 & ~i_8_214_1284_0 & ~i_8_214_1608_0 & ~i_8_214_1825_0 & ~i_8_214_1947_0 & ~i_8_214_1983_0 & ~i_8_214_2235_0 & ~i_8_214_2239_0) | (i_8_214_192_0 & ~i_8_214_665_0 & ~i_8_214_1072_0 & ~i_8_214_1812_0 & ~i_8_214_2158_0 & ~i_8_214_2229_0 & ~i_8_214_2232_0 & ~i_8_214_2262_0))) | (~i_8_214_192_0 & ~i_8_214_1565_0 & ((~i_8_214_348_0 & i_8_214_843_0 & ~i_8_214_1227_0 & ~i_8_214_1983_0 & ~i_8_214_2074_0 & ~i_8_214_2139_0) | (~i_8_214_237_0 & ~i_8_214_426_0 & i_8_214_696_0 & ~i_8_214_1947_0 & ~i_8_214_2070_0 & ~i_8_214_2112_0 & ~i_8_214_2227_0 & ~i_8_214_2232_0 & ~i_8_214_2235_0 & ~i_8_214_2262_0))) | (~i_8_214_237_0 & ~i_8_214_1605_0 & ((~i_8_214_527_0 & ~i_8_214_772_0 & i_8_214_1041_0 & ~i_8_214_2112_0 & i_8_214_2139_0 & ~i_8_214_2227_0) | (~i_8_214_1160_0 & i_8_214_1785_0 & i_8_214_2056_0 & ~i_8_214_2229_0 & ~i_8_214_2232_0 & ~i_8_214_2235_0))) | (~i_8_214_21_0 & ~i_8_214_426_0 & i_8_214_527_0 & ~i_8_214_2203_0))) | (i_8_214_385_0 & ((~i_8_214_527_0 & i_8_214_665_0 & ~i_8_214_772_0 & ~i_8_214_1160_0 & i_8_214_1565_0 & ~i_8_214_2074_0 & i_8_214_2158_0 & ~i_8_214_2229_0) | (~i_8_214_120_0 & ~i_8_214_237_0 & ~i_8_214_958_0 & ~i_8_214_1149_0 & ~i_8_214_1299_0 & i_8_214_2289_0))) | (~i_8_214_1983_0 & ((~i_8_214_237_0 & ((~i_8_214_285_0 & i_8_214_430_0 & i_8_214_1042_0 & ~i_8_214_1227_0 & ~i_8_214_1488_0 & ~i_8_214_1679_0 & i_8_214_1825_0 & ~i_8_214_1956_0 & ~i_8_214_2154_0) | (i_8_214_348_0 & ~i_8_214_706_0 & ~i_8_214_772_0 & ~i_8_214_843_0 & ~i_8_214_2056_0 & ~i_8_214_2112_0 & ~i_8_214_2232_0 & ~i_8_214_2262_0))) | (~i_8_214_348_0 & ((i_8_214_141_0 & ~i_8_214_1299_0 & ~i_8_214_1608_0 & ~i_8_214_1947_0 & ~i_8_214_1959_0 & ~i_8_214_2056_0 & ~i_8_214_2112_0 & ~i_8_214_2239_0) | (~i_8_214_285_0 & i_8_214_696_0 & i_8_214_832_0 & ~i_8_214_867_0 & i_8_214_966_0 & ~i_8_214_1560_0 & ~i_8_214_2289_0))) | (~i_8_214_18_0 & ~i_8_214_696_0 & ~i_8_214_1285_0 & ~i_8_214_1318_0 & ~i_8_214_1560_0 & ~i_8_214_1608_0 & ~i_8_214_1824_0 & ~i_8_214_1959_0 & ~i_8_214_2056_0 & ~i_8_214_2147_0 & ~i_8_214_2232_0 & ~i_8_214_2239_0))) | (~i_8_214_2112_0 & ((~i_8_214_18_0 & ((~i_8_214_385_0 & ((~i_8_214_21_0 & ((~i_8_214_843_0 & ~i_8_214_1149_0 & ~i_8_214_1227_0 & ~i_8_214_1605_0 & i_8_214_2154_0 & ~i_8_214_2227_0) | (~i_8_214_430_0 & ~i_8_214_1560_0 & ~i_8_214_1608_0 & ~i_8_214_1785_0 & ~i_8_214_1812_0 & ~i_8_214_1947_0 & ~i_8_214_2203_0 & ~i_8_214_2232_0 & ~i_8_214_2239_0))) | (~i_8_214_426_0 & ~i_8_214_1146_0 & ~i_8_214_1565_0 & ~i_8_214_2154_0 & ~i_8_214_2158_0 & ~i_8_214_2203_0 & ~i_8_214_2227_0 & ~i_8_214_2235_0))) | (~i_8_214_1299_0 & i_8_214_1719_0 & ~i_8_214_2227_0) | (~i_8_214_285_0 & i_8_214_426_0 & ~i_8_214_772_0 & i_8_214_1042_0 & ~i_8_214_1605_0 & ~i_8_214_1812_0 & ~i_8_214_2154_0 & ~i_8_214_2262_0))) | (~i_8_214_2289_0 & ((~i_8_214_966_0 & ((i_8_214_426_0 & ~i_8_214_709_0 & ~i_8_214_839_0 & ~i_8_214_1299_0 & ~i_8_214_1608_0 & i_8_214_1947_0 & ~i_8_214_2232_0) | (~i_8_214_957_0 & ~i_8_214_1149_0 & i_8_214_1489_0 & ~i_8_214_2262_0))) | (~i_8_214_772_0 & i_8_214_1149_0 & ~i_8_214_1160_0 & ~i_8_214_1488_0 & ~i_8_214_1608_0 & ~i_8_214_1686_0 & ~i_8_214_1770_0 & i_8_214_2227_0))))) | (~i_8_214_18_0 & ~i_8_214_1318_0 & ((~i_8_214_839_0 & ~i_8_214_1284_0 & ~i_8_214_1362_0 & i_8_214_1479_0 & ~i_8_214_1605_0) | (~i_8_214_21_0 & ~i_8_214_958_0 & i_8_214_1488_0 & ~i_8_214_1560_0 & ~i_8_214_1770_0 & ~i_8_214_2158_0 & ~i_8_214_2292_0))) | (~i_8_214_2203_0 & ((~i_8_214_21_0 & ~i_8_214_1812_0 & ((~i_8_214_348_0 & ~i_8_214_665_0 & ~i_8_214_966_0 & ~i_8_214_1042_0 & ~i_8_214_1072_0 & ~i_8_214_1227_0 & ~i_8_214_1299_0 & ~i_8_214_1560_0 & ~i_8_214_1686_0 & ~i_8_214_1719_0 & ~i_8_214_2154_0 & ~i_8_214_2158_0 & ~i_8_214_2227_0 & ~i_8_214_2232_0) | (~i_8_214_957_0 & ~i_8_214_958_0 & ~i_8_214_1284_0 & i_8_214_2147_0 & ~i_8_214_2235_0 & ~i_8_214_2239_0))) | (~i_8_214_2232_0 & ((i_8_214_1488_0 & i_8_214_1489_0 & ~i_8_214_1608_0) | (~i_8_214_385_0 & ~i_8_214_426_0 & ~i_8_214_696_0 & ~i_8_214_958_0 & ~i_8_214_1149_0 & ~i_8_214_1160_0 & ~i_8_214_1299_0 & ~i_8_214_1443_0 & ~i_8_214_1565_0 & ~i_8_214_1947_0 & ~i_8_214_2229_0 & ~i_8_214_2292_0))))) | (~i_8_214_348_0 & ((i_8_214_120_0 & i_8_214_696_0 & ~i_8_214_839_0 & ~i_8_214_1284_0 & i_8_214_1299_0 & ~i_8_214_2289_0) | (~i_8_214_426_0 & ~i_8_214_430_0 & ~i_8_214_1146_0 & ~i_8_214_1947_0 & i_8_214_2292_0))) | (~i_8_214_1560_0 & ((~i_8_214_665_0 & ~i_8_214_1146_0 & i_8_214_1490_0 & ~i_8_214_1605_0) | (~i_8_214_385_0 & ~i_8_214_867_0 & ~i_8_214_957_0 & ~i_8_214_966_0 & ~i_8_214_1072_0 & ~i_8_214_1284_0 & ~i_8_214_1947_0 & ~i_8_214_1956_0 & i_8_214_1983_0 & ~i_8_214_2147_0 & ~i_8_214_2292_0))) | (~i_8_214_385_0 & ~i_8_214_2070_0 & ((~i_8_214_1237_0 & ~i_8_214_1284_0 & ~i_8_214_1285_0 & ~i_8_214_1362_0 & i_8_214_1959_0 & i_8_214_2235_0) | (~i_8_214_1227_0 & ~i_8_214_2154_0 & ~i_8_214_2235_0 & ~i_8_214_2239_0 & i_8_214_2292_0))) | (~i_8_214_2154_0 & ((i_8_214_237_0 & ~i_8_214_706_0 & ~i_8_214_1284_0 & i_8_214_1560_0 & ~i_8_214_1605_0) | (i_8_214_706_0 & i_8_214_1480_0 & i_8_214_1770_0))) | (~i_8_214_2056_0 & i_8_214_2147_0 & i_8_214_2154_0 & i_8_214_2263_0 & ~i_8_214_2289_0));
endmodule



// Benchmark "kernel_8_215" written by ABC on Sun Jul 19 10:06:47 2020

module kernel_8_215 ( 
    i_8_215_53_0, i_8_215_58_0, i_8_215_101_0, i_8_215_107_0,
    i_8_215_210_0, i_8_215_227_0, i_8_215_232_0, i_8_215_256_0,
    i_8_215_323_0, i_8_215_361_0, i_8_215_362_0, i_8_215_364_0,
    i_8_215_365_0, i_8_215_373_0, i_8_215_400_0, i_8_215_426_0,
    i_8_215_442_0, i_8_215_454_0, i_8_215_553_0, i_8_215_571_0,
    i_8_215_660_0, i_8_215_676_0, i_8_215_679_0, i_8_215_699_0,
    i_8_215_700_0, i_8_215_703_0, i_8_215_710_0, i_8_215_759_0,
    i_8_215_838_0, i_8_215_841_0, i_8_215_859_0, i_8_215_877_0,
    i_8_215_887_0, i_8_215_968_0, i_8_215_970_0, i_8_215_1017_0,
    i_8_215_1067_0, i_8_215_1147_0, i_8_215_1189_0, i_8_215_1228_0,
    i_8_215_1229_0, i_8_215_1231_0, i_8_215_1281_0, i_8_215_1297_0,
    i_8_215_1300_0, i_8_215_1301_0, i_8_215_1308_0, i_8_215_1318_0,
    i_8_215_1339_0, i_8_215_1343_0, i_8_215_1344_0, i_8_215_1345_0,
    i_8_215_1363_0, i_8_215_1397_0, i_8_215_1400_0, i_8_215_1441_0,
    i_8_215_1467_0, i_8_215_1486_0, i_8_215_1489_0, i_8_215_1526_0,
    i_8_215_1559_0, i_8_215_1562_0, i_8_215_1574_0, i_8_215_1606_0,
    i_8_215_1607_0, i_8_215_1633_0, i_8_215_1672_0, i_8_215_1677_0,
    i_8_215_1678_0, i_8_215_1718_0, i_8_215_1720_0, i_8_215_1731_0,
    i_8_215_1738_0, i_8_215_1747_0, i_8_215_1748_0, i_8_215_1760_0,
    i_8_215_1763_0, i_8_215_1820_0, i_8_215_1834_0, i_8_215_1972_0,
    i_8_215_1982_0, i_8_215_1989_0, i_8_215_1996_0, i_8_215_2055_0,
    i_8_215_2056_0, i_8_215_2057_0, i_8_215_2107_0, i_8_215_2110_0,
    i_8_215_2111_0, i_8_215_2126_0, i_8_215_2147_0, i_8_215_2156_0,
    i_8_215_2172_0, i_8_215_2225_0, i_8_215_2226_0, i_8_215_2227_0,
    i_8_215_2230_0, i_8_215_2242_0, i_8_215_2248_0, i_8_215_2286_0,
    o_8_215_0_0  );
  input  i_8_215_53_0, i_8_215_58_0, i_8_215_101_0, i_8_215_107_0,
    i_8_215_210_0, i_8_215_227_0, i_8_215_232_0, i_8_215_256_0,
    i_8_215_323_0, i_8_215_361_0, i_8_215_362_0, i_8_215_364_0,
    i_8_215_365_0, i_8_215_373_0, i_8_215_400_0, i_8_215_426_0,
    i_8_215_442_0, i_8_215_454_0, i_8_215_553_0, i_8_215_571_0,
    i_8_215_660_0, i_8_215_676_0, i_8_215_679_0, i_8_215_699_0,
    i_8_215_700_0, i_8_215_703_0, i_8_215_710_0, i_8_215_759_0,
    i_8_215_838_0, i_8_215_841_0, i_8_215_859_0, i_8_215_877_0,
    i_8_215_887_0, i_8_215_968_0, i_8_215_970_0, i_8_215_1017_0,
    i_8_215_1067_0, i_8_215_1147_0, i_8_215_1189_0, i_8_215_1228_0,
    i_8_215_1229_0, i_8_215_1231_0, i_8_215_1281_0, i_8_215_1297_0,
    i_8_215_1300_0, i_8_215_1301_0, i_8_215_1308_0, i_8_215_1318_0,
    i_8_215_1339_0, i_8_215_1343_0, i_8_215_1344_0, i_8_215_1345_0,
    i_8_215_1363_0, i_8_215_1397_0, i_8_215_1400_0, i_8_215_1441_0,
    i_8_215_1467_0, i_8_215_1486_0, i_8_215_1489_0, i_8_215_1526_0,
    i_8_215_1559_0, i_8_215_1562_0, i_8_215_1574_0, i_8_215_1606_0,
    i_8_215_1607_0, i_8_215_1633_0, i_8_215_1672_0, i_8_215_1677_0,
    i_8_215_1678_0, i_8_215_1718_0, i_8_215_1720_0, i_8_215_1731_0,
    i_8_215_1738_0, i_8_215_1747_0, i_8_215_1748_0, i_8_215_1760_0,
    i_8_215_1763_0, i_8_215_1820_0, i_8_215_1834_0, i_8_215_1972_0,
    i_8_215_1982_0, i_8_215_1989_0, i_8_215_1996_0, i_8_215_2055_0,
    i_8_215_2056_0, i_8_215_2057_0, i_8_215_2107_0, i_8_215_2110_0,
    i_8_215_2111_0, i_8_215_2126_0, i_8_215_2147_0, i_8_215_2156_0,
    i_8_215_2172_0, i_8_215_2225_0, i_8_215_2226_0, i_8_215_2227_0,
    i_8_215_2230_0, i_8_215_2242_0, i_8_215_2248_0, i_8_215_2286_0;
  output o_8_215_0_0;
  assign o_8_215_0_0 = 0;
endmodule



// Benchmark "kernel_8_216" written by ABC on Sun Jul 19 10:06:49 2020

module kernel_8_216 ( 
    i_8_216_2_0, i_8_216_6_0, i_8_216_7_0, i_8_216_34_0, i_8_216_106_0,
    i_8_216_108_0, i_8_216_169_0, i_8_216_260_0, i_8_216_285_0,
    i_8_216_286_0, i_8_216_294_0, i_8_216_295_0, i_8_216_323_0,
    i_8_216_328_0, i_8_216_337_0, i_8_216_347_0, i_8_216_431_0,
    i_8_216_439_0, i_8_216_440_0, i_8_216_547_0, i_8_216_583_0,
    i_8_216_602_0, i_8_216_609_0, i_8_216_628_0, i_8_216_654_0,
    i_8_216_705_0, i_8_216_715_0, i_8_216_719_0, i_8_216_726_0,
    i_8_216_781_0, i_8_216_789_0, i_8_216_808_0, i_8_216_814_0,
    i_8_216_817_0, i_8_216_819_0, i_8_216_826_0, i_8_216_850_0,
    i_8_216_851_0, i_8_216_853_0, i_8_216_879_0, i_8_216_899_0,
    i_8_216_925_0, i_8_216_933_0, i_8_216_969_0, i_8_216_970_0,
    i_8_216_975_0, i_8_216_1074_0, i_8_216_1115_0, i_8_216_1133_0,
    i_8_216_1149_0, i_8_216_1185_0, i_8_216_1186_0, i_8_216_1192_0,
    i_8_216_1201_0, i_8_216_1267_0, i_8_216_1273_0, i_8_216_1281_0,
    i_8_216_1282_0, i_8_216_1284_0, i_8_216_1295_0, i_8_216_1300_0,
    i_8_216_1302_0, i_8_216_1339_0, i_8_216_1354_0, i_8_216_1385_0,
    i_8_216_1390_0, i_8_216_1411_0, i_8_216_1440_0, i_8_216_1444_0,
    i_8_216_1473_0, i_8_216_1489_0, i_8_216_1591_0, i_8_216_1614_0,
    i_8_216_1617_0, i_8_216_1628_0, i_8_216_1648_0, i_8_216_1653_0,
    i_8_216_1655_0, i_8_216_1663_0, i_8_216_1678_0, i_8_216_1754_0,
    i_8_216_1792_0, i_8_216_1849_0, i_8_216_1891_0, i_8_216_1898_0,
    i_8_216_2028_0, i_8_216_2031_0, i_8_216_2070_0, i_8_216_2137_0,
    i_8_216_2139_0, i_8_216_2140_0, i_8_216_2141_0, i_8_216_2147_0,
    i_8_216_2148_0, i_8_216_2150_0, i_8_216_2151_0, i_8_216_2154_0,
    i_8_216_2205_0, i_8_216_2220_0, i_8_216_2247_0,
    o_8_216_0_0  );
  input  i_8_216_2_0, i_8_216_6_0, i_8_216_7_0, i_8_216_34_0,
    i_8_216_106_0, i_8_216_108_0, i_8_216_169_0, i_8_216_260_0,
    i_8_216_285_0, i_8_216_286_0, i_8_216_294_0, i_8_216_295_0,
    i_8_216_323_0, i_8_216_328_0, i_8_216_337_0, i_8_216_347_0,
    i_8_216_431_0, i_8_216_439_0, i_8_216_440_0, i_8_216_547_0,
    i_8_216_583_0, i_8_216_602_0, i_8_216_609_0, i_8_216_628_0,
    i_8_216_654_0, i_8_216_705_0, i_8_216_715_0, i_8_216_719_0,
    i_8_216_726_0, i_8_216_781_0, i_8_216_789_0, i_8_216_808_0,
    i_8_216_814_0, i_8_216_817_0, i_8_216_819_0, i_8_216_826_0,
    i_8_216_850_0, i_8_216_851_0, i_8_216_853_0, i_8_216_879_0,
    i_8_216_899_0, i_8_216_925_0, i_8_216_933_0, i_8_216_969_0,
    i_8_216_970_0, i_8_216_975_0, i_8_216_1074_0, i_8_216_1115_0,
    i_8_216_1133_0, i_8_216_1149_0, i_8_216_1185_0, i_8_216_1186_0,
    i_8_216_1192_0, i_8_216_1201_0, i_8_216_1267_0, i_8_216_1273_0,
    i_8_216_1281_0, i_8_216_1282_0, i_8_216_1284_0, i_8_216_1295_0,
    i_8_216_1300_0, i_8_216_1302_0, i_8_216_1339_0, i_8_216_1354_0,
    i_8_216_1385_0, i_8_216_1390_0, i_8_216_1411_0, i_8_216_1440_0,
    i_8_216_1444_0, i_8_216_1473_0, i_8_216_1489_0, i_8_216_1591_0,
    i_8_216_1614_0, i_8_216_1617_0, i_8_216_1628_0, i_8_216_1648_0,
    i_8_216_1653_0, i_8_216_1655_0, i_8_216_1663_0, i_8_216_1678_0,
    i_8_216_1754_0, i_8_216_1792_0, i_8_216_1849_0, i_8_216_1891_0,
    i_8_216_1898_0, i_8_216_2028_0, i_8_216_2031_0, i_8_216_2070_0,
    i_8_216_2137_0, i_8_216_2139_0, i_8_216_2140_0, i_8_216_2141_0,
    i_8_216_2147_0, i_8_216_2148_0, i_8_216_2150_0, i_8_216_2151_0,
    i_8_216_2154_0, i_8_216_2205_0, i_8_216_2220_0, i_8_216_2247_0;
  output o_8_216_0_0;
  assign o_8_216_0_0 = ~((~i_8_216_726_0 & ((~i_8_216_933_0 & ~i_8_216_1185_0 & ~i_8_216_1390_0 & ~i_8_216_1614_0) | (~i_8_216_285_0 & ~i_8_216_440_0 & ~i_8_216_899_0 & ~i_8_216_2031_0))) | (~i_8_216_1201_0 & ((~i_8_216_439_0 & ~i_8_216_850_0 & ~i_8_216_1192_0 & ~i_8_216_1628_0 & ~i_8_216_1648_0) | (~i_8_216_6_0 & ~i_8_216_169_0 & ~i_8_216_817_0 & ~i_8_216_925_0 & ~i_8_216_2205_0))) | (~i_8_216_169_0 & ((~i_8_216_814_0 & ~i_8_216_933_0 & i_8_216_1267_0) | (~i_8_216_34_0 & ~i_8_216_1591_0 & i_8_216_2150_0))) | (~i_8_216_1339_0 & ((~i_8_216_851_0 & ~i_8_216_975_0 & ~i_8_216_1489_0 & ~i_8_216_1628_0 & ~i_8_216_2031_0) | (~i_8_216_295_0 & ~i_8_216_337_0 & ~i_8_216_899_0 & ~i_8_216_1385_0 & ~i_8_216_1440_0 & ~i_8_216_1898_0 & ~i_8_216_2154_0))) | (~i_8_216_826_0 & ~i_8_216_1614_0) | (~i_8_216_106_0 & ~i_8_216_1186_0 & ~i_8_216_1267_0 & ~i_8_216_1754_0));
endmodule



// Benchmark "kernel_8_217" written by ABC on Sun Jul 19 10:06:49 2020

module kernel_8_217 ( 
    i_8_217_15_0, i_8_217_20_0, i_8_217_21_0, i_8_217_41_0, i_8_217_65_0,
    i_8_217_115_0, i_8_217_226_0, i_8_217_299_0, i_8_217_316_0,
    i_8_217_319_0, i_8_217_363_0, i_8_217_415_0, i_8_217_418_0,
    i_8_217_447_0, i_8_217_460_0, i_8_217_483_0, i_8_217_495_0,
    i_8_217_497_0, i_8_217_532_0, i_8_217_550_0, i_8_217_553_0,
    i_8_217_568_0, i_8_217_577_0, i_8_217_596_0, i_8_217_608_0,
    i_8_217_635_0, i_8_217_650_0, i_8_217_705_0, i_8_217_729_0,
    i_8_217_760_0, i_8_217_818_0, i_8_217_859_0, i_8_217_879_0,
    i_8_217_880_0, i_8_217_918_0, i_8_217_968_0, i_8_217_976_0,
    i_8_217_1126_0, i_8_217_1132_0, i_8_217_1153_0, i_8_217_1171_0,
    i_8_217_1188_0, i_8_217_1198_0, i_8_217_1202_0, i_8_217_1226_0,
    i_8_217_1231_0, i_8_217_1234_0, i_8_217_1235_0, i_8_217_1261_0,
    i_8_217_1276_0, i_8_217_1324_0, i_8_217_1325_0, i_8_217_1328_0,
    i_8_217_1342_0, i_8_217_1353_0, i_8_217_1360_0, i_8_217_1378_0,
    i_8_217_1388_0, i_8_217_1396_0, i_8_217_1397_0, i_8_217_1432_0,
    i_8_217_1436_0, i_8_217_1459_0, i_8_217_1463_0, i_8_217_1468_0,
    i_8_217_1491_0, i_8_217_1511_0, i_8_217_1541_0, i_8_217_1556_0,
    i_8_217_1630_0, i_8_217_1643_0, i_8_217_1648_0, i_8_217_1679_0,
    i_8_217_1694_0, i_8_217_1714_0, i_8_217_1759_0, i_8_217_1778_0,
    i_8_217_1792_0, i_8_217_1819_0, i_8_217_1826_0, i_8_217_1838_0,
    i_8_217_1861_0, i_8_217_1873_0, i_8_217_1883_0, i_8_217_1946_0,
    i_8_217_1947_0, i_8_217_1972_0, i_8_217_1990_0, i_8_217_2061_0,
    i_8_217_2062_0, i_8_217_2065_0, i_8_217_2144_0, i_8_217_2145_0,
    i_8_217_2169_0, i_8_217_2170_0, i_8_217_2224_0, i_8_217_2242_0,
    i_8_217_2268_0, i_8_217_2269_0, i_8_217_2273_0,
    o_8_217_0_0  );
  input  i_8_217_15_0, i_8_217_20_0, i_8_217_21_0, i_8_217_41_0,
    i_8_217_65_0, i_8_217_115_0, i_8_217_226_0, i_8_217_299_0,
    i_8_217_316_0, i_8_217_319_0, i_8_217_363_0, i_8_217_415_0,
    i_8_217_418_0, i_8_217_447_0, i_8_217_460_0, i_8_217_483_0,
    i_8_217_495_0, i_8_217_497_0, i_8_217_532_0, i_8_217_550_0,
    i_8_217_553_0, i_8_217_568_0, i_8_217_577_0, i_8_217_596_0,
    i_8_217_608_0, i_8_217_635_0, i_8_217_650_0, i_8_217_705_0,
    i_8_217_729_0, i_8_217_760_0, i_8_217_818_0, i_8_217_859_0,
    i_8_217_879_0, i_8_217_880_0, i_8_217_918_0, i_8_217_968_0,
    i_8_217_976_0, i_8_217_1126_0, i_8_217_1132_0, i_8_217_1153_0,
    i_8_217_1171_0, i_8_217_1188_0, i_8_217_1198_0, i_8_217_1202_0,
    i_8_217_1226_0, i_8_217_1231_0, i_8_217_1234_0, i_8_217_1235_0,
    i_8_217_1261_0, i_8_217_1276_0, i_8_217_1324_0, i_8_217_1325_0,
    i_8_217_1328_0, i_8_217_1342_0, i_8_217_1353_0, i_8_217_1360_0,
    i_8_217_1378_0, i_8_217_1388_0, i_8_217_1396_0, i_8_217_1397_0,
    i_8_217_1432_0, i_8_217_1436_0, i_8_217_1459_0, i_8_217_1463_0,
    i_8_217_1468_0, i_8_217_1491_0, i_8_217_1511_0, i_8_217_1541_0,
    i_8_217_1556_0, i_8_217_1630_0, i_8_217_1643_0, i_8_217_1648_0,
    i_8_217_1679_0, i_8_217_1694_0, i_8_217_1714_0, i_8_217_1759_0,
    i_8_217_1778_0, i_8_217_1792_0, i_8_217_1819_0, i_8_217_1826_0,
    i_8_217_1838_0, i_8_217_1861_0, i_8_217_1873_0, i_8_217_1883_0,
    i_8_217_1946_0, i_8_217_1947_0, i_8_217_1972_0, i_8_217_1990_0,
    i_8_217_2061_0, i_8_217_2062_0, i_8_217_2065_0, i_8_217_2144_0,
    i_8_217_2145_0, i_8_217_2169_0, i_8_217_2170_0, i_8_217_2224_0,
    i_8_217_2242_0, i_8_217_2268_0, i_8_217_2269_0, i_8_217_2273_0;
  output o_8_217_0_0;
  assign o_8_217_0_0 = 0;
endmodule



// Benchmark "kernel_8_218" written by ABC on Sun Jul 19 10:06:50 2020

module kernel_8_218 ( 
    i_8_218_11_0, i_8_218_13_0, i_8_218_19_0, i_8_218_23_0, i_8_218_28_0,
    i_8_218_68_0, i_8_218_86_0, i_8_218_100_0, i_8_218_114_0,
    i_8_218_115_0, i_8_218_116_0, i_8_218_117_0, i_8_218_142_0,
    i_8_218_194_0, i_8_218_210_0, i_8_218_274_0, i_8_218_279_0,
    i_8_218_348_0, i_8_218_378_0, i_8_218_379_0, i_8_218_391_0,
    i_8_218_428_0, i_8_218_507_0, i_8_218_508_0, i_8_218_544_0,
    i_8_218_589_0, i_8_218_622_0, i_8_218_642_0, i_8_218_650_0,
    i_8_218_693_0, i_8_218_694_0, i_8_218_708_0, i_8_218_732_0,
    i_8_218_733_0, i_8_218_764_0, i_8_218_781_0, i_8_218_851_0,
    i_8_218_872_0, i_8_218_874_0, i_8_218_880_0, i_8_218_896_0,
    i_8_218_921_0, i_8_218_937_0, i_8_218_955_0, i_8_218_990_0,
    i_8_218_1027_0, i_8_218_1107_0, i_8_218_1114_0, i_8_218_1130_0,
    i_8_218_1134_0, i_8_218_1137_0, i_8_218_1139_0, i_8_218_1146_0,
    i_8_218_1224_0, i_8_218_1225_0, i_8_218_1260_0, i_8_218_1261_0,
    i_8_218_1264_0, i_8_218_1300_0, i_8_218_1315_0, i_8_218_1396_0,
    i_8_218_1400_0, i_8_218_1410_0, i_8_218_1422_0, i_8_218_1432_0,
    i_8_218_1492_0, i_8_218_1549_0, i_8_218_1611_0, i_8_218_1612_0,
    i_8_218_1633_0, i_8_218_1648_0, i_8_218_1668_0, i_8_218_1671_0,
    i_8_218_1681_0, i_8_218_1710_0, i_8_218_1718_0, i_8_218_1723_0,
    i_8_218_1751_0, i_8_218_1756_0, i_8_218_1775_0, i_8_218_1778_0,
    i_8_218_1803_0, i_8_218_1824_0, i_8_218_1840_0, i_8_218_1859_0,
    i_8_218_1868_0, i_8_218_1869_0, i_8_218_1884_0, i_8_218_1945_0,
    i_8_218_1946_0, i_8_218_1957_0, i_8_218_1989_0, i_8_218_2001_0,
    i_8_218_2053_0, i_8_218_2099_0, i_8_218_2138_0, i_8_218_2152_0,
    i_8_218_2197_0, i_8_218_2215_0, i_8_218_2263_0,
    o_8_218_0_0  );
  input  i_8_218_11_0, i_8_218_13_0, i_8_218_19_0, i_8_218_23_0,
    i_8_218_28_0, i_8_218_68_0, i_8_218_86_0, i_8_218_100_0, i_8_218_114_0,
    i_8_218_115_0, i_8_218_116_0, i_8_218_117_0, i_8_218_142_0,
    i_8_218_194_0, i_8_218_210_0, i_8_218_274_0, i_8_218_279_0,
    i_8_218_348_0, i_8_218_378_0, i_8_218_379_0, i_8_218_391_0,
    i_8_218_428_0, i_8_218_507_0, i_8_218_508_0, i_8_218_544_0,
    i_8_218_589_0, i_8_218_622_0, i_8_218_642_0, i_8_218_650_0,
    i_8_218_693_0, i_8_218_694_0, i_8_218_708_0, i_8_218_732_0,
    i_8_218_733_0, i_8_218_764_0, i_8_218_781_0, i_8_218_851_0,
    i_8_218_872_0, i_8_218_874_0, i_8_218_880_0, i_8_218_896_0,
    i_8_218_921_0, i_8_218_937_0, i_8_218_955_0, i_8_218_990_0,
    i_8_218_1027_0, i_8_218_1107_0, i_8_218_1114_0, i_8_218_1130_0,
    i_8_218_1134_0, i_8_218_1137_0, i_8_218_1139_0, i_8_218_1146_0,
    i_8_218_1224_0, i_8_218_1225_0, i_8_218_1260_0, i_8_218_1261_0,
    i_8_218_1264_0, i_8_218_1300_0, i_8_218_1315_0, i_8_218_1396_0,
    i_8_218_1400_0, i_8_218_1410_0, i_8_218_1422_0, i_8_218_1432_0,
    i_8_218_1492_0, i_8_218_1549_0, i_8_218_1611_0, i_8_218_1612_0,
    i_8_218_1633_0, i_8_218_1648_0, i_8_218_1668_0, i_8_218_1671_0,
    i_8_218_1681_0, i_8_218_1710_0, i_8_218_1718_0, i_8_218_1723_0,
    i_8_218_1751_0, i_8_218_1756_0, i_8_218_1775_0, i_8_218_1778_0,
    i_8_218_1803_0, i_8_218_1824_0, i_8_218_1840_0, i_8_218_1859_0,
    i_8_218_1868_0, i_8_218_1869_0, i_8_218_1884_0, i_8_218_1945_0,
    i_8_218_1946_0, i_8_218_1957_0, i_8_218_1989_0, i_8_218_2001_0,
    i_8_218_2053_0, i_8_218_2099_0, i_8_218_2138_0, i_8_218_2152_0,
    i_8_218_2197_0, i_8_218_2215_0, i_8_218_2263_0;
  output o_8_218_0_0;
  assign o_8_218_0_0 = 0;
endmodule



// Benchmark "kernel_8_219" written by ABC on Sun Jul 19 10:06:51 2020

module kernel_8_219 ( 
    i_8_219_22_0, i_8_219_24_0, i_8_219_34_0, i_8_219_39_0, i_8_219_67_0,
    i_8_219_158_0, i_8_219_180_0, i_8_219_223_0, i_8_219_229_0,
    i_8_219_262_0, i_8_219_300_0, i_8_219_370_0, i_8_219_379_0,
    i_8_219_381_0, i_8_219_426_0, i_8_219_440_0, i_8_219_534_0,
    i_8_219_535_0, i_8_219_592_0, i_8_219_602_0, i_8_219_610_0,
    i_8_219_613_0, i_8_219_628_0, i_8_219_655_0, i_8_219_660_0,
    i_8_219_695_0, i_8_219_703_0, i_8_219_704_0, i_8_219_706_0,
    i_8_219_727_0, i_8_219_753_0, i_8_219_771_0, i_8_219_816_0,
    i_8_219_838_0, i_8_219_840_0, i_8_219_843_0, i_8_219_849_0,
    i_8_219_850_0, i_8_219_853_0, i_8_219_869_0, i_8_219_876_0,
    i_8_219_877_0, i_8_219_940_0, i_8_219_979_0, i_8_219_980_0,
    i_8_219_984_0, i_8_219_993_0, i_8_219_1074_0, i_8_219_1126_0,
    i_8_219_1137_0, i_8_219_1157_0, i_8_219_1224_0, i_8_219_1225_0,
    i_8_219_1226_0, i_8_219_1227_0, i_8_219_1234_0, i_8_219_1263_0,
    i_8_219_1338_0, i_8_219_1346_0, i_8_219_1362_0, i_8_219_1379_0,
    i_8_219_1427_0, i_8_219_1467_0, i_8_219_1470_0, i_8_219_1506_0,
    i_8_219_1547_0, i_8_219_1549_0, i_8_219_1560_0, i_8_219_1574_0,
    i_8_219_1606_0, i_8_219_1615_0, i_8_219_1617_0, i_8_219_1650_0,
    i_8_219_1677_0, i_8_219_1686_0, i_8_219_1706_0, i_8_219_1729_0,
    i_8_219_1755_0, i_8_219_1759_0, i_8_219_1760_0, i_8_219_1787_0,
    i_8_219_1813_0, i_8_219_1824_0, i_8_219_1885_0, i_8_219_1974_0,
    i_8_219_1976_0, i_8_219_1983_0, i_8_219_1989_0, i_8_219_2002_0,
    i_8_219_2136_0, i_8_219_2143_0, i_8_219_2144_0, i_8_219_2146_0,
    i_8_219_2149_0, i_8_219_2158_0, i_8_219_2190_0, i_8_219_2191_0,
    i_8_219_2215_0, i_8_219_2226_0, i_8_219_2236_0,
    o_8_219_0_0  );
  input  i_8_219_22_0, i_8_219_24_0, i_8_219_34_0, i_8_219_39_0,
    i_8_219_67_0, i_8_219_158_0, i_8_219_180_0, i_8_219_223_0,
    i_8_219_229_0, i_8_219_262_0, i_8_219_300_0, i_8_219_370_0,
    i_8_219_379_0, i_8_219_381_0, i_8_219_426_0, i_8_219_440_0,
    i_8_219_534_0, i_8_219_535_0, i_8_219_592_0, i_8_219_602_0,
    i_8_219_610_0, i_8_219_613_0, i_8_219_628_0, i_8_219_655_0,
    i_8_219_660_0, i_8_219_695_0, i_8_219_703_0, i_8_219_704_0,
    i_8_219_706_0, i_8_219_727_0, i_8_219_753_0, i_8_219_771_0,
    i_8_219_816_0, i_8_219_838_0, i_8_219_840_0, i_8_219_843_0,
    i_8_219_849_0, i_8_219_850_0, i_8_219_853_0, i_8_219_869_0,
    i_8_219_876_0, i_8_219_877_0, i_8_219_940_0, i_8_219_979_0,
    i_8_219_980_0, i_8_219_984_0, i_8_219_993_0, i_8_219_1074_0,
    i_8_219_1126_0, i_8_219_1137_0, i_8_219_1157_0, i_8_219_1224_0,
    i_8_219_1225_0, i_8_219_1226_0, i_8_219_1227_0, i_8_219_1234_0,
    i_8_219_1263_0, i_8_219_1338_0, i_8_219_1346_0, i_8_219_1362_0,
    i_8_219_1379_0, i_8_219_1427_0, i_8_219_1467_0, i_8_219_1470_0,
    i_8_219_1506_0, i_8_219_1547_0, i_8_219_1549_0, i_8_219_1560_0,
    i_8_219_1574_0, i_8_219_1606_0, i_8_219_1615_0, i_8_219_1617_0,
    i_8_219_1650_0, i_8_219_1677_0, i_8_219_1686_0, i_8_219_1706_0,
    i_8_219_1729_0, i_8_219_1755_0, i_8_219_1759_0, i_8_219_1760_0,
    i_8_219_1787_0, i_8_219_1813_0, i_8_219_1824_0, i_8_219_1885_0,
    i_8_219_1974_0, i_8_219_1976_0, i_8_219_1983_0, i_8_219_1989_0,
    i_8_219_2002_0, i_8_219_2136_0, i_8_219_2143_0, i_8_219_2144_0,
    i_8_219_2146_0, i_8_219_2149_0, i_8_219_2158_0, i_8_219_2190_0,
    i_8_219_2191_0, i_8_219_2215_0, i_8_219_2226_0, i_8_219_2236_0;
  output o_8_219_0_0;
  assign o_8_219_0_0 = 0;
endmodule



// Benchmark "kernel_8_220" written by ABC on Sun Jul 19 10:06:52 2020

module kernel_8_220 ( 
    i_8_220_5_0, i_8_220_20_0, i_8_220_89_0, i_8_220_194_0, i_8_220_197_0,
    i_8_220_220_0, i_8_220_224_0, i_8_220_227_0, i_8_220_302_0,
    i_8_220_328_0, i_8_220_346_0, i_8_220_356_0, i_8_220_376_0,
    i_8_220_383_0, i_8_220_385_0, i_8_220_386_0, i_8_220_445_0,
    i_8_220_455_0, i_8_220_464_0, i_8_220_476_0, i_8_220_499_0,
    i_8_220_500_0, i_8_220_508_0, i_8_220_525_0, i_8_220_526_0,
    i_8_220_529_0, i_8_220_553_0, i_8_220_589_0, i_8_220_593_0,
    i_8_220_607_0, i_8_220_625_0, i_8_220_662_0, i_8_220_665_0,
    i_8_220_671_0, i_8_220_715_0, i_8_220_716_0, i_8_220_725_0,
    i_8_220_780_0, i_8_220_781_0, i_8_220_782_0, i_8_220_787_0,
    i_8_220_789_0, i_8_220_795_0, i_8_220_796_0, i_8_220_814_0,
    i_8_220_825_0, i_8_220_877_0, i_8_220_904_0, i_8_220_1012_0,
    i_8_220_1015_0, i_8_220_1030_0, i_8_220_1031_0, i_8_220_1086_0,
    i_8_220_1087_0, i_8_220_1132_0, i_8_220_1190_0, i_8_220_1193_0,
    i_8_220_1237_0, i_8_220_1256_0, i_8_220_1345_0, i_8_220_1436_0,
    i_8_220_1456_0, i_8_220_1457_0, i_8_220_1471_0, i_8_220_1540_0,
    i_8_220_1542_0, i_8_220_1544_0, i_8_220_1552_0, i_8_220_1579_0,
    i_8_220_1588_0, i_8_220_1598_0, i_8_220_1601_0, i_8_220_1607_0,
    i_8_220_1633_0, i_8_220_1636_0, i_8_220_1679_0, i_8_220_1714_0,
    i_8_220_1717_0, i_8_220_1732_0, i_8_220_1742_0, i_8_220_1754_0,
    i_8_220_1763_0, i_8_220_1894_0, i_8_220_1895_0, i_8_220_1918_0,
    i_8_220_1919_0, i_8_220_1933_0, i_8_220_1951_0, i_8_220_1967_0,
    i_8_220_1981_0, i_8_220_2005_0, i_8_220_2029_0, i_8_220_2047_0,
    i_8_220_2109_0, i_8_220_2112_0, i_8_220_2129_0, i_8_220_2171_0,
    i_8_220_2196_0, i_8_220_2289_0, i_8_220_2290_0,
    o_8_220_0_0  );
  input  i_8_220_5_0, i_8_220_20_0, i_8_220_89_0, i_8_220_194_0,
    i_8_220_197_0, i_8_220_220_0, i_8_220_224_0, i_8_220_227_0,
    i_8_220_302_0, i_8_220_328_0, i_8_220_346_0, i_8_220_356_0,
    i_8_220_376_0, i_8_220_383_0, i_8_220_385_0, i_8_220_386_0,
    i_8_220_445_0, i_8_220_455_0, i_8_220_464_0, i_8_220_476_0,
    i_8_220_499_0, i_8_220_500_0, i_8_220_508_0, i_8_220_525_0,
    i_8_220_526_0, i_8_220_529_0, i_8_220_553_0, i_8_220_589_0,
    i_8_220_593_0, i_8_220_607_0, i_8_220_625_0, i_8_220_662_0,
    i_8_220_665_0, i_8_220_671_0, i_8_220_715_0, i_8_220_716_0,
    i_8_220_725_0, i_8_220_780_0, i_8_220_781_0, i_8_220_782_0,
    i_8_220_787_0, i_8_220_789_0, i_8_220_795_0, i_8_220_796_0,
    i_8_220_814_0, i_8_220_825_0, i_8_220_877_0, i_8_220_904_0,
    i_8_220_1012_0, i_8_220_1015_0, i_8_220_1030_0, i_8_220_1031_0,
    i_8_220_1086_0, i_8_220_1087_0, i_8_220_1132_0, i_8_220_1190_0,
    i_8_220_1193_0, i_8_220_1237_0, i_8_220_1256_0, i_8_220_1345_0,
    i_8_220_1436_0, i_8_220_1456_0, i_8_220_1457_0, i_8_220_1471_0,
    i_8_220_1540_0, i_8_220_1542_0, i_8_220_1544_0, i_8_220_1552_0,
    i_8_220_1579_0, i_8_220_1588_0, i_8_220_1598_0, i_8_220_1601_0,
    i_8_220_1607_0, i_8_220_1633_0, i_8_220_1636_0, i_8_220_1679_0,
    i_8_220_1714_0, i_8_220_1717_0, i_8_220_1732_0, i_8_220_1742_0,
    i_8_220_1754_0, i_8_220_1763_0, i_8_220_1894_0, i_8_220_1895_0,
    i_8_220_1918_0, i_8_220_1919_0, i_8_220_1933_0, i_8_220_1951_0,
    i_8_220_1967_0, i_8_220_1981_0, i_8_220_2005_0, i_8_220_2029_0,
    i_8_220_2047_0, i_8_220_2109_0, i_8_220_2112_0, i_8_220_2129_0,
    i_8_220_2171_0, i_8_220_2196_0, i_8_220_2289_0, i_8_220_2290_0;
  output o_8_220_0_0;
  assign o_8_220_0_0 = 0;
endmodule



// Benchmark "kernel_8_221" written by ABC on Sun Jul 19 10:06:53 2020

module kernel_8_221 ( 
    i_8_221_26_0, i_8_221_31_0, i_8_221_41_0, i_8_221_57_0, i_8_221_68_0,
    i_8_221_95_0, i_8_221_98_0, i_8_221_107_0, i_8_221_166_0,
    i_8_221_167_0, i_8_221_176_0, i_8_221_179_0, i_8_221_215_0,
    i_8_221_227_0, i_8_221_229_0, i_8_221_260_0, i_8_221_266_0,
    i_8_221_314_0, i_8_221_338_0, i_8_221_359_0, i_8_221_363_0,
    i_8_221_374_0, i_8_221_386_0, i_8_221_427_0, i_8_221_428_0,
    i_8_221_431_0, i_8_221_449_0, i_8_221_455_0, i_8_221_487_0,
    i_8_221_494_0, i_8_221_522_0, i_8_221_539_0, i_8_221_589_0,
    i_8_221_593_0, i_8_221_653_0, i_8_221_656_0, i_8_221_661_0,
    i_8_221_665_0, i_8_221_693_0, i_8_221_694_0, i_8_221_699_0,
    i_8_221_702_0, i_8_221_706_0, i_8_221_710_0, i_8_221_771_0,
    i_8_221_809_0, i_8_221_838_0, i_8_221_842_0, i_8_221_869_0,
    i_8_221_881_0, i_8_221_948_0, i_8_221_959_0, i_8_221_965_0,
    i_8_221_966_0, i_8_221_1022_0, i_8_221_1024_0, i_8_221_1129_0,
    i_8_221_1166_0, i_8_221_1175_0, i_8_221_1231_0, i_8_221_1241_0,
    i_8_221_1268_0, i_8_221_1321_0, i_8_221_1337_0, i_8_221_1373_0,
    i_8_221_1376_0, i_8_221_1402_0, i_8_221_1419_0, i_8_221_1435_0,
    i_8_221_1453_0, i_8_221_1456_0, i_8_221_1472_0, i_8_221_1526_0,
    i_8_221_1546_0, i_8_221_1562_0, i_8_221_1646_0, i_8_221_1655_0,
    i_8_221_1672_0, i_8_221_1673_0, i_8_221_1691_0, i_8_221_1706_0,
    i_8_221_1790_0, i_8_221_1821_0, i_8_221_1822_0, i_8_221_1823_0,
    i_8_221_1825_0, i_8_221_1832_0, i_8_221_1868_0, i_8_221_1870_0,
    i_8_221_1930_0, i_8_221_1965_0, i_8_221_2077_0, i_8_221_2078_0,
    i_8_221_2113_0, i_8_221_2145_0, i_8_221_2227_0, i_8_221_2249_0,
    i_8_221_2267_0, i_8_221_2276_0, i_8_221_2285_0,
    o_8_221_0_0  );
  input  i_8_221_26_0, i_8_221_31_0, i_8_221_41_0, i_8_221_57_0,
    i_8_221_68_0, i_8_221_95_0, i_8_221_98_0, i_8_221_107_0, i_8_221_166_0,
    i_8_221_167_0, i_8_221_176_0, i_8_221_179_0, i_8_221_215_0,
    i_8_221_227_0, i_8_221_229_0, i_8_221_260_0, i_8_221_266_0,
    i_8_221_314_0, i_8_221_338_0, i_8_221_359_0, i_8_221_363_0,
    i_8_221_374_0, i_8_221_386_0, i_8_221_427_0, i_8_221_428_0,
    i_8_221_431_0, i_8_221_449_0, i_8_221_455_0, i_8_221_487_0,
    i_8_221_494_0, i_8_221_522_0, i_8_221_539_0, i_8_221_589_0,
    i_8_221_593_0, i_8_221_653_0, i_8_221_656_0, i_8_221_661_0,
    i_8_221_665_0, i_8_221_693_0, i_8_221_694_0, i_8_221_699_0,
    i_8_221_702_0, i_8_221_706_0, i_8_221_710_0, i_8_221_771_0,
    i_8_221_809_0, i_8_221_838_0, i_8_221_842_0, i_8_221_869_0,
    i_8_221_881_0, i_8_221_948_0, i_8_221_959_0, i_8_221_965_0,
    i_8_221_966_0, i_8_221_1022_0, i_8_221_1024_0, i_8_221_1129_0,
    i_8_221_1166_0, i_8_221_1175_0, i_8_221_1231_0, i_8_221_1241_0,
    i_8_221_1268_0, i_8_221_1321_0, i_8_221_1337_0, i_8_221_1373_0,
    i_8_221_1376_0, i_8_221_1402_0, i_8_221_1419_0, i_8_221_1435_0,
    i_8_221_1453_0, i_8_221_1456_0, i_8_221_1472_0, i_8_221_1526_0,
    i_8_221_1546_0, i_8_221_1562_0, i_8_221_1646_0, i_8_221_1655_0,
    i_8_221_1672_0, i_8_221_1673_0, i_8_221_1691_0, i_8_221_1706_0,
    i_8_221_1790_0, i_8_221_1821_0, i_8_221_1822_0, i_8_221_1823_0,
    i_8_221_1825_0, i_8_221_1832_0, i_8_221_1868_0, i_8_221_1870_0,
    i_8_221_1930_0, i_8_221_1965_0, i_8_221_2077_0, i_8_221_2078_0,
    i_8_221_2113_0, i_8_221_2145_0, i_8_221_2227_0, i_8_221_2249_0,
    i_8_221_2267_0, i_8_221_2276_0, i_8_221_2285_0;
  output o_8_221_0_0;
  assign o_8_221_0_0 = 0;
endmodule



// Benchmark "kernel_8_222" written by ABC on Sun Jul 19 10:06:54 2020

module kernel_8_222 ( 
    i_8_222_33_0, i_8_222_35_0, i_8_222_98_0, i_8_222_157_0, i_8_222_160_0,
    i_8_222_161_0, i_8_222_221_0, i_8_222_224_0, i_8_222_301_0,
    i_8_222_354_0, i_8_222_369_0, i_8_222_373_0, i_8_222_374_0,
    i_8_222_433_0, i_8_222_434_0, i_8_222_440_0, i_8_222_462_0,
    i_8_222_463_0, i_8_222_475_0, i_8_222_476_0, i_8_222_478_0,
    i_8_222_498_0, i_8_222_508_0, i_8_222_526_0, i_8_222_530_0,
    i_8_222_548_0, i_8_222_595_0, i_8_222_660_0, i_8_222_707_0,
    i_8_222_715_0, i_8_222_716_0, i_8_222_735_0, i_8_222_777_0,
    i_8_222_781_0, i_8_222_793_0, i_8_222_796_0, i_8_222_823_0,
    i_8_222_880_0, i_8_222_985_0, i_8_222_996_0, i_8_222_1009_0,
    i_8_222_1011_0, i_8_222_1012_0, i_8_222_1027_0, i_8_222_1085_0,
    i_8_222_1120_0, i_8_222_1121_0, i_8_222_1249_0, i_8_222_1256_0,
    i_8_222_1273_0, i_8_222_1285_0, i_8_222_1300_0, i_8_222_1344_0,
    i_8_222_1453_0, i_8_222_1456_0, i_8_222_1469_0, i_8_222_1471_0,
    i_8_222_1536_0, i_8_222_1540_0, i_8_222_1543_0, i_8_222_1544_0,
    i_8_222_1552_0, i_8_222_1553_0, i_8_222_1558_0, i_8_222_1574_0,
    i_8_222_1579_0, i_8_222_1587_0, i_8_222_1589_0, i_8_222_1597_0,
    i_8_222_1598_0, i_8_222_1629_0, i_8_222_1669_0, i_8_222_1714_0,
    i_8_222_1752_0, i_8_222_1780_0, i_8_222_1781_0, i_8_222_1783_0,
    i_8_222_1785_0, i_8_222_1807_0, i_8_222_1821_0, i_8_222_1840_0,
    i_8_222_1857_0, i_8_222_1858_0, i_8_222_1894_0, i_8_222_1895_0,
    i_8_222_1930_0, i_8_222_1950_0, i_8_222_1951_0, i_8_222_1974_0,
    i_8_222_1975_0, i_8_222_2102_0, i_8_222_2111_0, i_8_222_2128_0,
    i_8_222_2183_0, i_8_222_2191_0, i_8_222_2216_0, i_8_222_2224_0,
    i_8_222_2275_0, i_8_222_2289_0, i_8_222_2295_0,
    o_8_222_0_0  );
  input  i_8_222_33_0, i_8_222_35_0, i_8_222_98_0, i_8_222_157_0,
    i_8_222_160_0, i_8_222_161_0, i_8_222_221_0, i_8_222_224_0,
    i_8_222_301_0, i_8_222_354_0, i_8_222_369_0, i_8_222_373_0,
    i_8_222_374_0, i_8_222_433_0, i_8_222_434_0, i_8_222_440_0,
    i_8_222_462_0, i_8_222_463_0, i_8_222_475_0, i_8_222_476_0,
    i_8_222_478_0, i_8_222_498_0, i_8_222_508_0, i_8_222_526_0,
    i_8_222_530_0, i_8_222_548_0, i_8_222_595_0, i_8_222_660_0,
    i_8_222_707_0, i_8_222_715_0, i_8_222_716_0, i_8_222_735_0,
    i_8_222_777_0, i_8_222_781_0, i_8_222_793_0, i_8_222_796_0,
    i_8_222_823_0, i_8_222_880_0, i_8_222_985_0, i_8_222_996_0,
    i_8_222_1009_0, i_8_222_1011_0, i_8_222_1012_0, i_8_222_1027_0,
    i_8_222_1085_0, i_8_222_1120_0, i_8_222_1121_0, i_8_222_1249_0,
    i_8_222_1256_0, i_8_222_1273_0, i_8_222_1285_0, i_8_222_1300_0,
    i_8_222_1344_0, i_8_222_1453_0, i_8_222_1456_0, i_8_222_1469_0,
    i_8_222_1471_0, i_8_222_1536_0, i_8_222_1540_0, i_8_222_1543_0,
    i_8_222_1544_0, i_8_222_1552_0, i_8_222_1553_0, i_8_222_1558_0,
    i_8_222_1574_0, i_8_222_1579_0, i_8_222_1587_0, i_8_222_1589_0,
    i_8_222_1597_0, i_8_222_1598_0, i_8_222_1629_0, i_8_222_1669_0,
    i_8_222_1714_0, i_8_222_1752_0, i_8_222_1780_0, i_8_222_1781_0,
    i_8_222_1783_0, i_8_222_1785_0, i_8_222_1807_0, i_8_222_1821_0,
    i_8_222_1840_0, i_8_222_1857_0, i_8_222_1858_0, i_8_222_1894_0,
    i_8_222_1895_0, i_8_222_1930_0, i_8_222_1950_0, i_8_222_1951_0,
    i_8_222_1974_0, i_8_222_1975_0, i_8_222_2102_0, i_8_222_2111_0,
    i_8_222_2128_0, i_8_222_2183_0, i_8_222_2191_0, i_8_222_2216_0,
    i_8_222_2224_0, i_8_222_2275_0, i_8_222_2289_0, i_8_222_2295_0;
  output o_8_222_0_0;
  assign o_8_222_0_0 = 0;
endmodule



// Benchmark "kernel_8_223" written by ABC on Sun Jul 19 10:06:56 2020

module kernel_8_223 ( 
    i_8_223_11_0, i_8_223_52_0, i_8_223_53_0, i_8_223_70_0, i_8_223_79_0,
    i_8_223_95_0, i_8_223_111_0, i_8_223_112_0, i_8_223_188_0,
    i_8_223_221_0, i_8_223_250_0, i_8_223_256_0, i_8_223_297_0,
    i_8_223_301_0, i_8_223_305_0, i_8_223_346_0, i_8_223_348_0,
    i_8_223_349_0, i_8_223_360_0, i_8_223_362_0, i_8_223_363_0,
    i_8_223_364_0, i_8_223_365_0, i_8_223_366_0, i_8_223_368_0,
    i_8_223_479_0, i_8_223_555_0, i_8_223_557_0, i_8_223_615_0,
    i_8_223_625_0, i_8_223_635_0, i_8_223_658_0, i_8_223_688_0,
    i_8_223_762_0, i_8_223_770_0, i_8_223_816_0, i_8_223_817_0,
    i_8_223_837_0, i_8_223_838_0, i_8_223_843_0, i_8_223_844_0,
    i_8_223_859_0, i_8_223_860_0, i_8_223_862_0, i_8_223_863_0,
    i_8_223_877_0, i_8_223_879_0, i_8_223_880_0, i_8_223_881_0,
    i_8_223_938_0, i_8_223_942_0, i_8_223_943_0, i_8_223_944_0,
    i_8_223_978_0, i_8_223_1030_0, i_8_223_1045_0, i_8_223_1086_0,
    i_8_223_1087_0, i_8_223_1113_0, i_8_223_1138_0, i_8_223_1148_0,
    i_8_223_1203_0, i_8_223_1301_0, i_8_223_1302_0, i_8_223_1306_0,
    i_8_223_1307_0, i_8_223_1410_0, i_8_223_1455_0, i_8_223_1456_0,
    i_8_223_1511_0, i_8_223_1533_0, i_8_223_1535_0, i_8_223_1543_0,
    i_8_223_1546_0, i_8_223_1649_0, i_8_223_1651_0, i_8_223_1764_0,
    i_8_223_1807_0, i_8_223_1888_0, i_8_223_1915_0, i_8_223_1918_0,
    i_8_223_1997_0, i_8_223_2013_0, i_8_223_2046_0, i_8_223_2048_0,
    i_8_223_2051_0, i_8_223_2111_0, i_8_223_2112_0, i_8_223_2113_0,
    i_8_223_2119_0, i_8_223_2121_0, i_8_223_2123_0, i_8_223_2132_0,
    i_8_223_2140_0, i_8_223_2213_0, i_8_223_2215_0, i_8_223_2216_0,
    i_8_223_2298_0, i_8_223_2299_0, i_8_223_2300_0,
    o_8_223_0_0  );
  input  i_8_223_11_0, i_8_223_52_0, i_8_223_53_0, i_8_223_70_0,
    i_8_223_79_0, i_8_223_95_0, i_8_223_111_0, i_8_223_112_0,
    i_8_223_188_0, i_8_223_221_0, i_8_223_250_0, i_8_223_256_0,
    i_8_223_297_0, i_8_223_301_0, i_8_223_305_0, i_8_223_346_0,
    i_8_223_348_0, i_8_223_349_0, i_8_223_360_0, i_8_223_362_0,
    i_8_223_363_0, i_8_223_364_0, i_8_223_365_0, i_8_223_366_0,
    i_8_223_368_0, i_8_223_479_0, i_8_223_555_0, i_8_223_557_0,
    i_8_223_615_0, i_8_223_625_0, i_8_223_635_0, i_8_223_658_0,
    i_8_223_688_0, i_8_223_762_0, i_8_223_770_0, i_8_223_816_0,
    i_8_223_817_0, i_8_223_837_0, i_8_223_838_0, i_8_223_843_0,
    i_8_223_844_0, i_8_223_859_0, i_8_223_860_0, i_8_223_862_0,
    i_8_223_863_0, i_8_223_877_0, i_8_223_879_0, i_8_223_880_0,
    i_8_223_881_0, i_8_223_938_0, i_8_223_942_0, i_8_223_943_0,
    i_8_223_944_0, i_8_223_978_0, i_8_223_1030_0, i_8_223_1045_0,
    i_8_223_1086_0, i_8_223_1087_0, i_8_223_1113_0, i_8_223_1138_0,
    i_8_223_1148_0, i_8_223_1203_0, i_8_223_1301_0, i_8_223_1302_0,
    i_8_223_1306_0, i_8_223_1307_0, i_8_223_1410_0, i_8_223_1455_0,
    i_8_223_1456_0, i_8_223_1511_0, i_8_223_1533_0, i_8_223_1535_0,
    i_8_223_1543_0, i_8_223_1546_0, i_8_223_1649_0, i_8_223_1651_0,
    i_8_223_1764_0, i_8_223_1807_0, i_8_223_1888_0, i_8_223_1915_0,
    i_8_223_1918_0, i_8_223_1997_0, i_8_223_2013_0, i_8_223_2046_0,
    i_8_223_2048_0, i_8_223_2051_0, i_8_223_2111_0, i_8_223_2112_0,
    i_8_223_2113_0, i_8_223_2119_0, i_8_223_2121_0, i_8_223_2123_0,
    i_8_223_2132_0, i_8_223_2140_0, i_8_223_2213_0, i_8_223_2215_0,
    i_8_223_2216_0, i_8_223_2298_0, i_8_223_2299_0, i_8_223_2300_0;
  output o_8_223_0_0;
  assign o_8_223_0_0 = ~((~i_8_223_2048_0 & ((~i_8_223_53_0 & ((~i_8_223_11_0 & ~i_8_223_555_0 & ~i_8_223_615_0 & ~i_8_223_859_0 & ~i_8_223_938_0 & ~i_8_223_1045_0 & ~i_8_223_1301_0 & i_8_223_1535_0 & ~i_8_223_1915_0 & ~i_8_223_2051_0 & ~i_8_223_2140_0) | (~i_8_223_368_0 & ~i_8_223_770_0 & ~i_8_223_877_0 & ~i_8_223_943_0 & ~i_8_223_1535_0 & ~i_8_223_1807_0 & ~i_8_223_2299_0 & i_8_223_2300_0))) | (~i_8_223_70_0 & ((~i_8_223_11_0 & ~i_8_223_635_0 & ~i_8_223_860_0 & ~i_8_223_862_0 & ~i_8_223_863_0 & ~i_8_223_938_0 & ~i_8_223_942_0 & ~i_8_223_1045_0 & ~i_8_223_1086_0 & ~i_8_223_1307_0 & ~i_8_223_1511_0 & ~i_8_223_1807_0 & ~i_8_223_2046_0 & ~i_8_223_2121_0 & ~i_8_223_2123_0 & ~i_8_223_2215_0) | (i_8_223_349_0 & ~i_8_223_944_0 & ~i_8_223_1301_0 & ~i_8_223_1302_0 & ~i_8_223_1915_0 & ~i_8_223_2298_0))) | (~i_8_223_2051_0 & ((~i_8_223_557_0 & ~i_8_223_2300_0 & ((~i_8_223_11_0 & ~i_8_223_479_0 & ((~i_8_223_112_0 & ~i_8_223_635_0 & ~i_8_223_860_0 & ~i_8_223_944_0 & ~i_8_223_1045_0 & ~i_8_223_1086_0 & ~i_8_223_1087_0 & ~i_8_223_1410_0 & ~i_8_223_2123_0 & ~i_8_223_2298_0) | (~i_8_223_816_0 & ~i_8_223_817_0 & ~i_8_223_863_0 & ~i_8_223_938_0 & ~i_8_223_942_0 & ~i_8_223_943_0 & ~i_8_223_1302_0 & ~i_8_223_1306_0 & ~i_8_223_1307_0 & ~i_8_223_2046_0 & ~i_8_223_2216_0 & ~i_8_223_2299_0))) | (~i_8_223_221_0 & ~i_8_223_250_0 & ~i_8_223_256_0 & ~i_8_223_297_0 & ~i_8_223_346_0 & ~i_8_223_635_0 & ~i_8_223_860_0 & ~i_8_223_943_0 & ~i_8_223_1045_0 & ~i_8_223_1306_0 & ~i_8_223_1307_0 & ~i_8_223_1533_0 & ~i_8_223_1535_0 & ~i_8_223_1651_0 & ~i_8_223_2121_0 & ~i_8_223_2216_0))) | (~i_8_223_938_0 & ((~i_8_223_297_0 & ~i_8_223_362_0 & ~i_8_223_615_0 & ~i_8_223_1148_0 & ~i_8_223_1307_0 & ~i_8_223_1535_0 & i_8_223_1918_0 & ~i_8_223_1997_0 & ~i_8_223_2215_0 & ~i_8_223_2216_0) | (i_8_223_301_0 & ~i_8_223_349_0 & ~i_8_223_635_0 & ~i_8_223_862_0 & ~i_8_223_881_0 & ~i_8_223_942_0 & ~i_8_223_1301_0 & ~i_8_223_1456_0 & ~i_8_223_1915_0 & ~i_8_223_2299_0))))) | (~i_8_223_635_0 & ((~i_8_223_305_0 & i_8_223_877_0 & ~i_8_223_938_0 & ~i_8_223_1203_0 & ~i_8_223_1302_0 & ~i_8_223_1651_0 & ~i_8_223_1997_0 & ~i_8_223_2121_0 & ~i_8_223_2123_0 & ~i_8_223_2215_0 & ~i_8_223_2298_0) | (~i_8_223_615_0 & i_8_223_880_0 & ~i_8_223_1086_0 & ~i_8_223_1138_0 & ~i_8_223_1511_0 & ~i_8_223_1807_0 & ~i_8_223_1888_0 & ~i_8_223_2046_0 & ~i_8_223_2300_0))) | (~i_8_223_860_0 & ((~i_8_223_250_0 & i_8_223_346_0 & ~i_8_223_688_0 & ~i_8_223_816_0 & ~i_8_223_817_0 & ~i_8_223_862_0 & ~i_8_223_1087_0 & ~i_8_223_1649_0 & ~i_8_223_2111_0) | (~i_8_223_363_0 & i_8_223_368_0 & ~i_8_223_555_0 & ~i_8_223_557_0 & ~i_8_223_762_0 & ~i_8_223_938_0 & ~i_8_223_944_0 & ~i_8_223_1030_0 & ~i_8_223_1045_0 & ~i_8_223_1511_0 & ~i_8_223_2121_0 & ~i_8_223_2123_0))) | (i_8_223_53_0 & ~i_8_223_221_0 & ~i_8_223_863_0 & ~i_8_223_1302_0 & ~i_8_223_1511_0 & ~i_8_223_1535_0 & ~i_8_223_1651_0 & ~i_8_223_2013_0 & ~i_8_223_2123_0))) | (~i_8_223_1807_0 & ((~i_8_223_2051_0 & ((~i_8_223_221_0 & ~i_8_223_1113_0 & ~i_8_223_2046_0 & ~i_8_223_2300_0 & ((~i_8_223_479_0 & ~i_8_223_635_0 & ~i_8_223_688_0 & ~i_8_223_862_0 & i_8_223_877_0) | (~i_8_223_79_0 & ~i_8_223_297_0 & ~i_8_223_368_0 & ~i_8_223_816_0 & ~i_8_223_817_0 & ~i_8_223_938_0 & ~i_8_223_942_0 & ~i_8_223_1301_0 & ~i_8_223_1535_0 & ~i_8_223_2123_0 & ~i_8_223_2132_0 & ~i_8_223_2215_0))) | (~i_8_223_368_0 & ~i_8_223_615_0 & i_8_223_1511_0 & i_8_223_1997_0) | (~i_8_223_688_0 & ~i_8_223_844_0 & ~i_8_223_860_0 & ~i_8_223_938_0 & ~i_8_223_1030_0 & ~i_8_223_1301_0 & ~i_8_223_1456_0 & ~i_8_223_1511_0 & ~i_8_223_1535_0 & ~i_8_223_1651_0 & ~i_8_223_1918_0 & ~i_8_223_2121_0 & ~i_8_223_2123_0 & ~i_8_223_2299_0))) | (i_8_223_301_0 & i_8_223_479_0 & i_8_223_635_0 & ~i_8_223_1045_0) | (~i_8_223_112_0 & ~i_8_223_305_0 & ~i_8_223_557_0 & ~i_8_223_635_0 & ~i_8_223_1306_0 & ~i_8_223_1649_0 & ~i_8_223_1651_0 & ~i_8_223_1918_0 & ~i_8_223_1997_0 & ~i_8_223_2013_0 & ~i_8_223_2112_0 & ~i_8_223_2113_0 & ~i_8_223_2123_0 & ~i_8_223_2213_0))) | (~i_8_223_256_0 & ((~i_8_223_79_0 & ((~i_8_223_555_0 & ~i_8_223_1086_0 & i_8_223_2112_0) | (i_8_223_221_0 & ~i_8_223_250_0 & i_8_223_301_0 & ~i_8_223_2051_0 & ~i_8_223_2140_0 & ~i_8_223_860_0 & ~i_8_223_2013_0))) | (~i_8_223_112_0 & ~i_8_223_635_0 & ~i_8_223_816_0 & ~i_8_223_860_0 & ~i_8_223_1203_0 & ~i_8_223_1301_0 & ~i_8_223_1410_0 & ~i_8_223_1511_0 & ~i_8_223_1888_0 & ~i_8_223_2132_0 & i_8_223_2215_0 & ~i_8_223_2300_0))) | (~i_8_223_112_0 & ((i_8_223_221_0 & ~i_8_223_297_0 & i_8_223_479_0 & ~i_8_223_635_0 & ~i_8_223_860_0 & ~i_8_223_943_0 & ~i_8_223_1764_0 & ~i_8_223_1915_0) | (i_8_223_635_0 & ~i_8_223_1307_0 & ~i_8_223_1533_0 & i_8_223_2216_0 & ~i_8_223_2299_0 & i_8_223_2300_0))) | (~i_8_223_250_0 & ~i_8_223_555_0 & ((~i_8_223_11_0 & i_8_223_111_0 & ~i_8_223_762_0 & ~i_8_223_860_0 & ~i_8_223_938_0 & ~i_8_223_942_0 & ~i_8_223_1203_0 & ~i_8_223_1410_0 & ~i_8_223_2215_0) | (i_8_223_221_0 & ~i_8_223_305_0 & i_8_223_635_0 & ~i_8_223_943_0 & ~i_8_223_944_0 & ~i_8_223_1543_0 & i_8_223_2299_0))) | (i_8_223_365_0 & ~i_8_223_938_0 & ((~i_8_223_1086_0 & ~i_8_223_1087_0 & ~i_8_223_863_0 & ~i_8_223_944_0 & ~i_8_223_1302_0 & ~i_8_223_1535_0 & ~i_8_223_2216_0 & ~i_8_223_2298_0) | (~i_8_223_978_0 & ~i_8_223_1888_0 & ~i_8_223_2123_0 & ~i_8_223_2132_0 & ~i_8_223_2299_0 & ~i_8_223_2300_0))) | (~i_8_223_557_0 & ((i_8_223_363_0 & ~i_8_223_816_0 & ~i_8_223_862_0 & ~i_8_223_1086_0 & ~i_8_223_1087_0 & ~i_8_223_2119_0) | (i_8_223_364_0 & ~i_8_223_368_0 & ~i_8_223_942_0 & ~i_8_223_1203_0 & ~i_8_223_2299_0))) | (~i_8_223_862_0 & ((i_8_223_625_0 & ((~i_8_223_688_0 & ~i_8_223_1087_0 & ~i_8_223_1410_0 & i_8_223_1807_0 & ~i_8_223_2051_0) | (~i_8_223_817_0 & ~i_8_223_1302_0 & ~i_8_223_2121_0 & ~i_8_223_2216_0 & ~i_8_223_2298_0))) | (~i_8_223_2299_0 & ((i_8_223_881_0 & ~i_8_223_944_0 & ~i_8_223_1086_0 & ~i_8_223_1651_0 & ~i_8_223_2013_0 & i_8_223_2140_0) | (~i_8_223_859_0 & i_8_223_877_0 & i_8_223_1543_0 & ~i_8_223_2140_0))))) | (~i_8_223_817_0 & ((~i_8_223_880_0 & ~i_8_223_944_0 & ~i_8_223_978_0 & ~i_8_223_1301_0 & ~i_8_223_1307_0 & ~i_8_223_1410_0 & ~i_8_223_1535_0 & i_8_223_2132_0) | (i_8_223_112_0 & ~i_8_223_349_0 & i_8_223_844_0 & ~i_8_223_1086_0 & ~i_8_223_1113_0 & ~i_8_223_1306_0 & ~i_8_223_2123_0 & ~i_8_223_2300_0))) | (~i_8_223_2119_0 & ((~i_8_223_942_0 & ((~i_8_223_635_0 & ~i_8_223_762_0 & i_8_223_879_0 & ~i_8_223_978_0 & ~i_8_223_1086_0 & ~i_8_223_1301_0) | (i_8_223_362_0 & ~i_8_223_944_0 & ~i_8_223_2300_0))) | (~i_8_223_1997_0 & ~i_8_223_2121_0 & i_8_223_188_0 & ~i_8_223_1535_0))) | (~i_8_223_1307_0 & ((~i_8_223_1087_0 & ((i_8_223_1148_0 & ~i_8_223_1410_0 & ~i_8_223_2123_0) | (~i_8_223_111_0 & i_8_223_256_0 & ~i_8_223_978_0 & ~i_8_223_1511_0 & ~i_8_223_2213_0))) | (~i_8_223_658_0 & ~i_8_223_863_0 & i_8_223_1030_0 & ~i_8_223_1113_0))) | (~i_8_223_863_0 & ~i_8_223_1535_0 & ((i_8_223_349_0 & ~i_8_223_1511_0 & i_8_223_2051_0) | (i_8_223_838_0 & ~i_8_223_1915_0 & ~i_8_223_2013_0 & ~i_8_223_2123_0 & ~i_8_223_2298_0))) | (i_8_223_843_0 & i_8_223_1543_0));
endmodule



// Benchmark "kernel_8_224" written by ABC on Sun Jul 19 10:06:57 2020

module kernel_8_224 ( 
    i_8_224_38_0, i_8_224_58_0, i_8_224_71_0, i_8_224_76_0, i_8_224_83_0,
    i_8_224_181_0, i_8_224_185_0, i_8_224_244_0, i_8_224_305_0,
    i_8_224_317_0, i_8_224_320_0, i_8_224_322_0, i_8_224_323_0,
    i_8_224_365_0, i_8_224_424_0, i_8_224_425_0, i_8_224_426_0,
    i_8_224_525_0, i_8_224_532_0, i_8_224_534_0, i_8_224_542_0,
    i_8_224_556_0, i_8_224_603_0, i_8_224_610_0, i_8_224_614_0,
    i_8_224_634_0, i_8_224_635_0, i_8_224_638_0, i_8_224_657_0,
    i_8_224_676_0, i_8_224_679_0, i_8_224_697_0, i_8_224_703_0,
    i_8_224_706_0, i_8_224_707_0, i_8_224_752_0, i_8_224_753_0,
    i_8_224_790_0, i_8_224_806_0, i_8_224_844_0, i_8_224_866_0,
    i_8_224_889_0, i_8_224_890_0, i_8_224_951_0, i_8_224_956_0,
    i_8_224_974_0, i_8_224_984_0, i_8_224_987_0, i_8_224_1003_0,
    i_8_224_1056_0, i_8_224_1060_0, i_8_224_1115_0, i_8_224_1138_0,
    i_8_224_1152_0, i_8_224_1166_0, i_8_224_1167_0, i_8_224_1190_0,
    i_8_224_1201_0, i_8_224_1225_0, i_8_224_1238_0, i_8_224_1247_0,
    i_8_224_1273_0, i_8_224_1282_0, i_8_224_1399_0, i_8_224_1415_0,
    i_8_224_1433_0, i_8_224_1439_0, i_8_224_1456_0, i_8_224_1463_0,
    i_8_224_1491_0, i_8_224_1507_0, i_8_224_1527_0, i_8_224_1546_0,
    i_8_224_1561_0, i_8_224_1606_0, i_8_224_1617_0, i_8_224_1678_0,
    i_8_224_1714_0, i_8_224_1722_0, i_8_224_1744_0, i_8_224_1784_0,
    i_8_224_1787_0, i_8_224_1791_0, i_8_224_1822_0, i_8_224_1826_0,
    i_8_224_1949_0, i_8_224_1957_0, i_8_224_1966_0, i_8_224_1967_0,
    i_8_224_1982_0, i_8_224_1985_0, i_8_224_1996_0, i_8_224_2047_0,
    i_8_224_2144_0, i_8_224_2153_0, i_8_224_2156_0, i_8_224_2188_0,
    i_8_224_2200_0, i_8_224_2226_0, i_8_224_2302_0,
    o_8_224_0_0  );
  input  i_8_224_38_0, i_8_224_58_0, i_8_224_71_0, i_8_224_76_0,
    i_8_224_83_0, i_8_224_181_0, i_8_224_185_0, i_8_224_244_0,
    i_8_224_305_0, i_8_224_317_0, i_8_224_320_0, i_8_224_322_0,
    i_8_224_323_0, i_8_224_365_0, i_8_224_424_0, i_8_224_425_0,
    i_8_224_426_0, i_8_224_525_0, i_8_224_532_0, i_8_224_534_0,
    i_8_224_542_0, i_8_224_556_0, i_8_224_603_0, i_8_224_610_0,
    i_8_224_614_0, i_8_224_634_0, i_8_224_635_0, i_8_224_638_0,
    i_8_224_657_0, i_8_224_676_0, i_8_224_679_0, i_8_224_697_0,
    i_8_224_703_0, i_8_224_706_0, i_8_224_707_0, i_8_224_752_0,
    i_8_224_753_0, i_8_224_790_0, i_8_224_806_0, i_8_224_844_0,
    i_8_224_866_0, i_8_224_889_0, i_8_224_890_0, i_8_224_951_0,
    i_8_224_956_0, i_8_224_974_0, i_8_224_984_0, i_8_224_987_0,
    i_8_224_1003_0, i_8_224_1056_0, i_8_224_1060_0, i_8_224_1115_0,
    i_8_224_1138_0, i_8_224_1152_0, i_8_224_1166_0, i_8_224_1167_0,
    i_8_224_1190_0, i_8_224_1201_0, i_8_224_1225_0, i_8_224_1238_0,
    i_8_224_1247_0, i_8_224_1273_0, i_8_224_1282_0, i_8_224_1399_0,
    i_8_224_1415_0, i_8_224_1433_0, i_8_224_1439_0, i_8_224_1456_0,
    i_8_224_1463_0, i_8_224_1491_0, i_8_224_1507_0, i_8_224_1527_0,
    i_8_224_1546_0, i_8_224_1561_0, i_8_224_1606_0, i_8_224_1617_0,
    i_8_224_1678_0, i_8_224_1714_0, i_8_224_1722_0, i_8_224_1744_0,
    i_8_224_1784_0, i_8_224_1787_0, i_8_224_1791_0, i_8_224_1822_0,
    i_8_224_1826_0, i_8_224_1949_0, i_8_224_1957_0, i_8_224_1966_0,
    i_8_224_1967_0, i_8_224_1982_0, i_8_224_1985_0, i_8_224_1996_0,
    i_8_224_2047_0, i_8_224_2144_0, i_8_224_2153_0, i_8_224_2156_0,
    i_8_224_2188_0, i_8_224_2200_0, i_8_224_2226_0, i_8_224_2302_0;
  output o_8_224_0_0;
  assign o_8_224_0_0 = 0;
endmodule



// Benchmark "kernel_8_225" written by ABC on Sun Jul 19 10:06:58 2020

module kernel_8_225 ( 
    i_8_225_12_0, i_8_225_58_0, i_8_225_111_0, i_8_225_137_0,
    i_8_225_142_0, i_8_225_190_0, i_8_225_193_0, i_8_225_198_0,
    i_8_225_238_0, i_8_225_254_0, i_8_225_289_0, i_8_225_311_0,
    i_8_225_346_0, i_8_225_373_0, i_8_225_379_0, i_8_225_390_0,
    i_8_225_414_0, i_8_225_417_0, i_8_225_439_0, i_8_225_450_0,
    i_8_225_487_0, i_8_225_493_0, i_8_225_555_0, i_8_225_596_0,
    i_8_225_610_0, i_8_225_642_0, i_8_225_645_0, i_8_225_649_0,
    i_8_225_660_0, i_8_225_679_0, i_8_225_695_0, i_8_225_699_0,
    i_8_225_705_0, i_8_225_766_0, i_8_225_783_0, i_8_225_786_0,
    i_8_225_840_0, i_8_225_844_0, i_8_225_845_0, i_8_225_876_0,
    i_8_225_929_0, i_8_225_967_0, i_8_225_970_0, i_8_225_995_0,
    i_8_225_1064_0, i_8_225_1182_0, i_8_225_1185_0, i_8_225_1224_0,
    i_8_225_1226_0, i_8_225_1240_0, i_8_225_1255_0, i_8_225_1285_0,
    i_8_225_1288_0, i_8_225_1289_0, i_8_225_1300_0, i_8_225_1310_0,
    i_8_225_1314_0, i_8_225_1351_0, i_8_225_1354_0, i_8_225_1362_0,
    i_8_225_1381_0, i_8_225_1387_0, i_8_225_1461_0, i_8_225_1472_0,
    i_8_225_1481_0, i_8_225_1515_0, i_8_225_1540_0, i_8_225_1542_0,
    i_8_225_1545_0, i_8_225_1546_0, i_8_225_1632_0, i_8_225_1666_0,
    i_8_225_1671_0, i_8_225_1684_0, i_8_225_1693_0, i_8_225_1694_0,
    i_8_225_1699_0, i_8_225_1706_0, i_8_225_1747_0, i_8_225_1749_0,
    i_8_225_1758_0, i_8_225_1807_0, i_8_225_1826_0, i_8_225_1831_0,
    i_8_225_1855_0, i_8_225_1867_0, i_8_225_1887_0, i_8_225_1992_0,
    i_8_225_1993_0, i_8_225_2014_0, i_8_225_2071_0, i_8_225_2133_0,
    i_8_225_2142_0, i_8_225_2146_0, i_8_225_2151_0, i_8_225_2158_0,
    i_8_225_2226_0, i_8_225_2244_0, i_8_225_2278_0, i_8_225_2290_0,
    o_8_225_0_0  );
  input  i_8_225_12_0, i_8_225_58_0, i_8_225_111_0, i_8_225_137_0,
    i_8_225_142_0, i_8_225_190_0, i_8_225_193_0, i_8_225_198_0,
    i_8_225_238_0, i_8_225_254_0, i_8_225_289_0, i_8_225_311_0,
    i_8_225_346_0, i_8_225_373_0, i_8_225_379_0, i_8_225_390_0,
    i_8_225_414_0, i_8_225_417_0, i_8_225_439_0, i_8_225_450_0,
    i_8_225_487_0, i_8_225_493_0, i_8_225_555_0, i_8_225_596_0,
    i_8_225_610_0, i_8_225_642_0, i_8_225_645_0, i_8_225_649_0,
    i_8_225_660_0, i_8_225_679_0, i_8_225_695_0, i_8_225_699_0,
    i_8_225_705_0, i_8_225_766_0, i_8_225_783_0, i_8_225_786_0,
    i_8_225_840_0, i_8_225_844_0, i_8_225_845_0, i_8_225_876_0,
    i_8_225_929_0, i_8_225_967_0, i_8_225_970_0, i_8_225_995_0,
    i_8_225_1064_0, i_8_225_1182_0, i_8_225_1185_0, i_8_225_1224_0,
    i_8_225_1226_0, i_8_225_1240_0, i_8_225_1255_0, i_8_225_1285_0,
    i_8_225_1288_0, i_8_225_1289_0, i_8_225_1300_0, i_8_225_1310_0,
    i_8_225_1314_0, i_8_225_1351_0, i_8_225_1354_0, i_8_225_1362_0,
    i_8_225_1381_0, i_8_225_1387_0, i_8_225_1461_0, i_8_225_1472_0,
    i_8_225_1481_0, i_8_225_1515_0, i_8_225_1540_0, i_8_225_1542_0,
    i_8_225_1545_0, i_8_225_1546_0, i_8_225_1632_0, i_8_225_1666_0,
    i_8_225_1671_0, i_8_225_1684_0, i_8_225_1693_0, i_8_225_1694_0,
    i_8_225_1699_0, i_8_225_1706_0, i_8_225_1747_0, i_8_225_1749_0,
    i_8_225_1758_0, i_8_225_1807_0, i_8_225_1826_0, i_8_225_1831_0,
    i_8_225_1855_0, i_8_225_1867_0, i_8_225_1887_0, i_8_225_1992_0,
    i_8_225_1993_0, i_8_225_2014_0, i_8_225_2071_0, i_8_225_2133_0,
    i_8_225_2142_0, i_8_225_2146_0, i_8_225_2151_0, i_8_225_2158_0,
    i_8_225_2226_0, i_8_225_2244_0, i_8_225_2278_0, i_8_225_2290_0;
  output o_8_225_0_0;
  assign o_8_225_0_0 = 0;
endmodule



// Benchmark "kernel_8_226" written by ABC on Sun Jul 19 10:07:00 2020

module kernel_8_226 ( 
    i_8_226_53_0, i_8_226_80_0, i_8_226_114_0, i_8_226_115_0,
    i_8_226_120_0, i_8_226_123_0, i_8_226_228_0, i_8_226_371_0,
    i_8_226_381_0, i_8_226_382_0, i_8_226_428_0, i_8_226_451_0,
    i_8_226_454_0, i_8_226_481_0, i_8_226_511_0, i_8_226_570_0,
    i_8_226_571_0, i_8_226_575_0, i_8_226_590_0, i_8_226_599_0,
    i_8_226_605_0, i_8_226_636_0, i_8_226_658_0, i_8_226_660_0,
    i_8_226_663_0, i_8_226_747_0, i_8_226_835_0, i_8_226_873_0,
    i_8_226_886_0, i_8_226_887_0, i_8_226_990_0, i_8_226_1028_0,
    i_8_226_1031_0, i_8_226_1044_0, i_8_226_1048_0, i_8_226_1061_0,
    i_8_226_1072_0, i_8_226_1073_0, i_8_226_1074_0, i_8_226_1111_0,
    i_8_226_1164_0, i_8_226_1187_0, i_8_226_1227_0, i_8_226_1228_0,
    i_8_226_1229_0, i_8_226_1230_0, i_8_226_1231_0, i_8_226_1309_0,
    i_8_226_1331_0, i_8_226_1338_0, i_8_226_1356_0, i_8_226_1370_0,
    i_8_226_1403_0, i_8_226_1411_0, i_8_226_1434_0, i_8_226_1467_0,
    i_8_226_1470_0, i_8_226_1472_0, i_8_226_1474_0, i_8_226_1489_0,
    i_8_226_1556_0, i_8_226_1621_0, i_8_226_1632_0, i_8_226_1633_0,
    i_8_226_1635_0, i_8_226_1637_0, i_8_226_1654_0, i_8_226_1655_0,
    i_8_226_1659_0, i_8_226_1702_0, i_8_226_1704_0, i_8_226_1705_0,
    i_8_226_1736_0, i_8_226_1746_0, i_8_226_1747_0, i_8_226_1749_0,
    i_8_226_1751_0, i_8_226_1752_0, i_8_226_1764_0, i_8_226_1803_0,
    i_8_226_1820_0, i_8_226_1823_0, i_8_226_1857_0, i_8_226_1862_0,
    i_8_226_1945_0, i_8_226_1950_0, i_8_226_1983_0, i_8_226_1984_0,
    i_8_226_1985_0, i_8_226_2058_0, i_8_226_2073_0, i_8_226_2078_0,
    i_8_226_2125_0, i_8_226_2144_0, i_8_226_2172_0, i_8_226_2173_0,
    i_8_226_2218_0, i_8_226_2227_0, i_8_226_2248_0, i_8_226_2276_0,
    o_8_226_0_0  );
  input  i_8_226_53_0, i_8_226_80_0, i_8_226_114_0, i_8_226_115_0,
    i_8_226_120_0, i_8_226_123_0, i_8_226_228_0, i_8_226_371_0,
    i_8_226_381_0, i_8_226_382_0, i_8_226_428_0, i_8_226_451_0,
    i_8_226_454_0, i_8_226_481_0, i_8_226_511_0, i_8_226_570_0,
    i_8_226_571_0, i_8_226_575_0, i_8_226_590_0, i_8_226_599_0,
    i_8_226_605_0, i_8_226_636_0, i_8_226_658_0, i_8_226_660_0,
    i_8_226_663_0, i_8_226_747_0, i_8_226_835_0, i_8_226_873_0,
    i_8_226_886_0, i_8_226_887_0, i_8_226_990_0, i_8_226_1028_0,
    i_8_226_1031_0, i_8_226_1044_0, i_8_226_1048_0, i_8_226_1061_0,
    i_8_226_1072_0, i_8_226_1073_0, i_8_226_1074_0, i_8_226_1111_0,
    i_8_226_1164_0, i_8_226_1187_0, i_8_226_1227_0, i_8_226_1228_0,
    i_8_226_1229_0, i_8_226_1230_0, i_8_226_1231_0, i_8_226_1309_0,
    i_8_226_1331_0, i_8_226_1338_0, i_8_226_1356_0, i_8_226_1370_0,
    i_8_226_1403_0, i_8_226_1411_0, i_8_226_1434_0, i_8_226_1467_0,
    i_8_226_1470_0, i_8_226_1472_0, i_8_226_1474_0, i_8_226_1489_0,
    i_8_226_1556_0, i_8_226_1621_0, i_8_226_1632_0, i_8_226_1633_0,
    i_8_226_1635_0, i_8_226_1637_0, i_8_226_1654_0, i_8_226_1655_0,
    i_8_226_1659_0, i_8_226_1702_0, i_8_226_1704_0, i_8_226_1705_0,
    i_8_226_1736_0, i_8_226_1746_0, i_8_226_1747_0, i_8_226_1749_0,
    i_8_226_1751_0, i_8_226_1752_0, i_8_226_1764_0, i_8_226_1803_0,
    i_8_226_1820_0, i_8_226_1823_0, i_8_226_1857_0, i_8_226_1862_0,
    i_8_226_1945_0, i_8_226_1950_0, i_8_226_1983_0, i_8_226_1984_0,
    i_8_226_1985_0, i_8_226_2058_0, i_8_226_2073_0, i_8_226_2078_0,
    i_8_226_2125_0, i_8_226_2144_0, i_8_226_2172_0, i_8_226_2173_0,
    i_8_226_2218_0, i_8_226_2227_0, i_8_226_2248_0, i_8_226_2276_0;
  output o_8_226_0_0;
  assign o_8_226_0_0 = ~((~i_8_226_1061_0 & ((~i_8_226_228_0 & ((~i_8_226_451_0 & i_8_226_590_0 & ~i_8_226_873_0 & ~i_8_226_990_0 & ~i_8_226_1031_0 & ~i_8_226_1331_0 & ~i_8_226_1702_0 & ~i_8_226_1736_0 & ~i_8_226_1862_0) | (~i_8_226_570_0 & ~i_8_226_575_0 & ~i_8_226_1164_0 & ~i_8_226_1411_0 & i_8_226_1434_0 & ~i_8_226_1746_0 & ~i_8_226_1751_0 & ~i_8_226_1764_0 & ~i_8_226_1984_0 & ~i_8_226_2078_0 & ~i_8_226_2227_0))) | (~i_8_226_123_0 & ~i_8_226_605_0 & ~i_8_226_835_0 & ~i_8_226_1164_0 & ~i_8_226_1633_0 & ~i_8_226_1764_0 & i_8_226_1820_0) | (~i_8_226_120_0 & ~i_8_226_371_0 & ~i_8_226_575_0 & ~i_8_226_887_0 & ~i_8_226_1048_0 & ~i_8_226_1621_0 & ~i_8_226_1702_0 & ~i_8_226_1736_0 & ~i_8_226_1803_0 & ~i_8_226_1857_0 & ~i_8_226_1983_0 & ~i_8_226_1984_0 & ~i_8_226_2172_0 & ~i_8_226_2218_0))) | (i_8_226_381_0 & ((~i_8_226_114_0 & i_8_226_382_0 & ~i_8_226_1044_0 & ~i_8_226_1227_0 & ~i_8_226_1356_0 & ~i_8_226_1820_0) | (~i_8_226_570_0 & ~i_8_226_571_0 & ~i_8_226_835_0 & ~i_8_226_1803_0 & ~i_8_226_1950_0 & ~i_8_226_2125_0 & ~i_8_226_2276_0))) | (~i_8_226_1621_0 & ((~i_8_226_1356_0 & ((~i_8_226_382_0 & ((~i_8_226_747_0 & ~i_8_226_1309_0 & ~i_8_226_1338_0 & ~i_8_226_1411_0 & ~i_8_226_1655_0 & i_8_226_1823_0) | (~i_8_226_570_0 & ~i_8_226_636_0 & ~i_8_226_835_0 & ~i_8_226_990_0 & ~i_8_226_1048_0 & ~i_8_226_1164_0 & ~i_8_226_1187_0 & ~i_8_226_1230_0 & ~i_8_226_1403_0 & ~i_8_226_1489_0 & ~i_8_226_1556_0 & ~i_8_226_1635_0 & ~i_8_226_1704_0 & ~i_8_226_1705_0 & ~i_8_226_1736_0 & ~i_8_226_1747_0 & ~i_8_226_1764_0 & ~i_8_226_1950_0 & ~i_8_226_2248_0))) | (i_8_226_511_0 & ~i_8_226_1857_0 & ~i_8_226_2058_0 & ~i_8_226_2078_0))) | (~i_8_226_575_0 & ((~i_8_226_887_0 & ~i_8_226_1164_0 & i_8_226_1751_0 & ~i_8_226_1764_0) | (i_8_226_454_0 & ~i_8_226_663_0 & ~i_8_226_1044_0 & ~i_8_226_1187_0 & ~i_8_226_1309_0 & ~i_8_226_2073_0 & ~i_8_226_2218_0))) | (~i_8_226_2276_0 & ((i_8_226_371_0 & ~i_8_226_451_0 & ~i_8_226_886_0 & ~i_8_226_1556_0) | (i_8_226_599_0 & ~i_8_226_1803_0 & ~i_8_226_1984_0 & ~i_8_226_2058_0 & ~i_8_226_2078_0))) | (i_8_226_663_0 & ~i_8_226_747_0 & ~i_8_226_1187_0 & ~i_8_226_1659_0 & i_8_226_1752_0) | (~i_8_226_114_0 & ~i_8_226_115_0 & ~i_8_226_873_0 & i_8_226_1434_0 & ~i_8_226_1747_0 & ~i_8_226_1764_0 & ~i_8_226_1985_0 & ~i_8_226_2073_0 & ~i_8_226_2218_0))) | (~i_8_226_575_0 & ((~i_8_226_123_0 & ((~i_8_226_114_0 & ~i_8_226_571_0 & ~i_8_226_873_0 & ~i_8_226_990_0 & ~i_8_226_1187_0 & ~i_8_226_1736_0 & i_8_226_1823_0 & ~i_8_226_1857_0 & ~i_8_226_1984_0 & ~i_8_226_2058_0) | (i_8_226_53_0 & ~i_8_226_663_0 & ~i_8_226_1044_0 & ~i_8_226_1048_0 & ~i_8_226_1655_0 & ~i_8_226_2078_0))) | (~i_8_226_481_0 & ((~i_8_226_1044_0 & ~i_8_226_1338_0 & i_8_226_1474_0 & ~i_8_226_1659_0) | (~i_8_226_571_0 & ~i_8_226_835_0 & ~i_8_226_990_0 & ~i_8_226_1736_0 & ~i_8_226_1857_0 & ~i_8_226_1862_0 & i_8_226_1985_0))) | (~i_8_226_571_0 & ((~i_8_226_120_0 & ~i_8_226_990_0 & ~i_8_226_1655_0 & ~i_8_226_1764_0 & i_8_226_1820_0 & ~i_8_226_1857_0) | (~i_8_226_511_0 & ~i_8_226_599_0 & ~i_8_226_605_0 & ~i_8_226_747_0 & ~i_8_226_887_0 & ~i_8_226_1164_0 & ~i_8_226_1489_0 & i_8_226_1621_0 & ~i_8_226_1747_0 & ~i_8_226_2125_0))) | (~i_8_226_120_0 & ((~i_8_226_1048_0 & ~i_8_226_1309_0 & ~i_8_226_1411_0 & i_8_226_1823_0) | (~i_8_226_115_0 & ~i_8_226_873_0 & i_8_226_1111_0 & ~i_8_226_1489_0 & ~i_8_226_1659_0 & ~i_8_226_1857_0 & ~i_8_226_1983_0 & ~i_8_226_2218_0))) | (~i_8_226_570_0 & ~i_8_226_605_0 & ~i_8_226_636_0 & ~i_8_226_873_0 & ~i_8_226_1044_0 & ~i_8_226_1164_0 & ~i_8_226_1411_0 & ~i_8_226_1489_0 & ~i_8_226_1654_0 & ~i_8_226_1736_0 & ~i_8_226_1752_0 & ~i_8_226_1862_0 & ~i_8_226_2125_0 & ~i_8_226_2144_0 & ~i_8_226_2218_0))) | (~i_8_226_571_0 & ((i_8_226_887_0 & ~i_8_226_1187_0 & i_8_226_1637_0 & ~i_8_226_1823_0) | (~i_8_226_599_0 & ~i_8_226_835_0 & i_8_226_1031_0 & ~i_8_226_1655_0 & ~i_8_226_1820_0 & ~i_8_226_1857_0))) | (~i_8_226_660_0 & ((~i_8_226_663_0 & ~i_8_226_1031_0 & ~i_8_226_1164_0 & i_8_226_1227_0 & ~i_8_226_1764_0 & ~i_8_226_1985_0) | (~i_8_226_120_0 & ~i_8_226_990_0 & ~i_8_226_1370_0 & ~i_8_226_1736_0 & ~i_8_226_2125_0 & i_8_226_2144_0))) | (~i_8_226_747_0 & ((~i_8_226_663_0 & ~i_8_226_1411_0 & i_8_226_1746_0 & ~i_8_226_1983_0 & ~i_8_226_2058_0) | (~i_8_226_570_0 & ~i_8_226_886_0 & i_8_226_1749_0 & ~i_8_226_1764_0 & ~i_8_226_2125_0))) | (~i_8_226_886_0 & ((~i_8_226_114_0 & i_8_226_1111_0 & ~i_8_226_1702_0 & i_8_226_1945_0 & ~i_8_226_2125_0) | (~i_8_226_570_0 & i_8_226_660_0 & i_8_226_1074_0 & ~i_8_226_2218_0))) | (~i_8_226_1111_0 & ((~i_8_226_990_0 & i_8_226_1048_0 & i_8_226_1621_0 & ~i_8_226_1702_0 & ~i_8_226_1764_0 & ~i_8_226_1820_0 & ~i_8_226_2058_0 & ~i_8_226_2173_0) | (~i_8_226_114_0 & ~i_8_226_115_0 & ~i_8_226_123_0 & ~i_8_226_835_0 & ~i_8_226_887_0 & ~i_8_226_1044_0 & i_8_226_1309_0 & ~i_8_226_1857_0 & ~i_8_226_1862_0 & ~i_8_226_1983_0 & ~i_8_226_1985_0 & i_8_226_2218_0 & ~i_8_226_2248_0))) | (~i_8_226_114_0 & ((~i_8_226_990_0 & ~i_8_226_1074_0 & ~i_8_226_1164_0 & ~i_8_226_1411_0 & i_8_226_1749_0) | (~i_8_226_120_0 & i_8_226_1230_0 & i_8_226_1803_0 & ~i_8_226_1820_0))) | (~i_8_226_1164_0 & ((~i_8_226_835_0 & ((~i_8_226_115_0 & ~i_8_226_1187_0 & ~i_8_226_2058_0 & ((~i_8_226_570_0 & ~i_8_226_990_0 & ~i_8_226_1370_0 & ~i_8_226_1556_0 & ~i_8_226_1659_0 & i_8_226_1803_0 & ~i_8_226_1984_0) | (~i_8_226_123_0 & i_8_226_382_0 & ~i_8_226_1764_0 & ~i_8_226_2173_0))) | (~i_8_226_120_0 & i_8_226_382_0 & ~i_8_226_1338_0 & ~i_8_226_1411_0 & ~i_8_226_1736_0 & ~i_8_226_1803_0))) | (~i_8_226_887_0 & ~i_8_226_1031_0 & ~i_8_226_1044_0 & i_8_226_1403_0 & ~i_8_226_2218_0) | (i_8_226_382_0 & ~i_8_226_990_0 & ~i_8_226_1074_0 & ~i_8_226_1632_0 & ~i_8_226_1635_0 & ~i_8_226_1736_0 & ~i_8_226_1803_0 & ~i_8_226_1823_0 & ~i_8_226_1857_0 & ~i_8_226_2073_0 & ~i_8_226_2248_0))) | (~i_8_226_2218_0 & ((~i_8_226_570_0 & ((~i_8_226_1074_0 & i_8_226_1230_0 & i_8_226_1231_0 & ~i_8_226_1489_0) | (~i_8_226_123_0 & i_8_226_636_0 & ~i_8_226_873_0 & ~i_8_226_1073_0 & ~i_8_226_1654_0 & ~i_8_226_1945_0 & ~i_8_226_1985_0 & ~i_8_226_2173_0))) | (~i_8_226_120_0 & ~i_8_226_835_0 & ~i_8_226_1044_0 & i_8_226_1632_0 & ~i_8_226_1655_0 & ~i_8_226_1736_0) | (~i_8_226_658_0 & i_8_226_1746_0 & ~i_8_226_1945_0 & ~i_8_226_1985_0 & ~i_8_226_2058_0 & ~i_8_226_2125_0 & ~i_8_226_2173_0))) | (~i_8_226_120_0 & ((~i_8_226_1736_0 & ~i_8_226_1862_0 & i_8_226_80_0 & i_8_226_1556_0) | (~i_8_226_1044_0 & ~i_8_226_1338_0 & ~i_8_226_1356_0 & i_8_226_1747_0 & ~i_8_226_1764_0 & ~i_8_226_2248_0))) | (~i_8_226_123_0 & i_8_226_1752_0 & (i_8_226_1632_0 | (~i_8_226_1764_0 & ~i_8_226_1857_0 & i_8_226_2058_0))) | (~i_8_226_1556_0 & ((i_8_226_1187_0 & i_8_226_1331_0) | (~i_8_226_1187_0 & i_8_226_1472_0 & ~i_8_226_1633_0 & ~i_8_226_1637_0 & ~i_8_226_1659_0 & ~i_8_226_1945_0))) | (i_8_226_990_0 & i_8_226_1111_0 & i_8_226_1434_0 & ~i_8_226_1752_0 & ~i_8_226_1857_0 & i_8_226_1984_0 & ~i_8_226_2058_0) | (i_8_226_1073_0 & ~i_8_226_1985_0 & ~i_8_226_2125_0 & ~i_8_226_2172_0) | (i_8_226_1655_0 & ~i_8_226_1736_0 & i_8_226_2058_0 & i_8_226_2218_0 & ~i_8_226_2248_0) | (~i_8_226_887_0 & ~i_8_226_1044_0 & i_8_226_1227_0 & i_8_226_1556_0 & ~i_8_226_2276_0));
endmodule



// Benchmark "kernel_8_227" written by ABC on Sun Jul 19 10:07:01 2020

module kernel_8_227 ( 
    i_8_227_65_0, i_8_227_107_0, i_8_227_115_0, i_8_227_140_0,
    i_8_227_172_0, i_8_227_173_0, i_8_227_269_0, i_8_227_284_0,
    i_8_227_293_0, i_8_227_323_0, i_8_227_353_0, i_8_227_360_0,
    i_8_227_368_0, i_8_227_382_0, i_8_227_398_0, i_8_227_452_0,
    i_8_227_489_0, i_8_227_490_0, i_8_227_492_0, i_8_227_530_0,
    i_8_227_590_0, i_8_227_614_0, i_8_227_634_0, i_8_227_706_0,
    i_8_227_707_0, i_8_227_764_0, i_8_227_797_0, i_8_227_833_0,
    i_8_227_845_0, i_8_227_858_0, i_8_227_859_0, i_8_227_868_0,
    i_8_227_922_0, i_8_227_969_0, i_8_227_1057_0, i_8_227_1058_0,
    i_8_227_1073_0, i_8_227_1100_0, i_8_227_1127_0, i_8_227_1129_0,
    i_8_227_1225_0, i_8_227_1226_0, i_8_227_1229_0, i_8_227_1262_0,
    i_8_227_1264_0, i_8_227_1298_0, i_8_227_1317_0, i_8_227_1325_0,
    i_8_227_1328_0, i_8_227_1366_0, i_8_227_1405_0, i_8_227_1406_0,
    i_8_227_1411_0, i_8_227_1435_0, i_8_227_1436_0, i_8_227_1456_0,
    i_8_227_1462_0, i_8_227_1463_0, i_8_227_1473_0, i_8_227_1522_0,
    i_8_227_1547_0, i_8_227_1549_0, i_8_227_1556_0, i_8_227_1622_0,
    i_8_227_1623_0, i_8_227_1633_0, i_8_227_1640_0, i_8_227_1730_0,
    i_8_227_1748_0, i_8_227_1757_0, i_8_227_1777_0, i_8_227_1784_0,
    i_8_227_1796_0, i_8_227_1823_0, i_8_227_1825_0, i_8_227_1832_0,
    i_8_227_1849_0, i_8_227_1867_0, i_8_227_1904_0, i_8_227_1957_0,
    i_8_227_1958_0, i_8_227_1975_0, i_8_227_1994_0, i_8_227_1996_0,
    i_8_227_1997_0, i_8_227_2003_0, i_8_227_2017_0, i_8_227_2020_0,
    i_8_227_2099_0, i_8_227_2117_0, i_8_227_2144_0, i_8_227_2150_0,
    i_8_227_2201_0, i_8_227_2225_0, i_8_227_2226_0, i_8_227_2244_0,
    i_8_227_2246_0, i_8_227_2249_0, i_8_227_2260_0, i_8_227_2287_0,
    o_8_227_0_0  );
  input  i_8_227_65_0, i_8_227_107_0, i_8_227_115_0, i_8_227_140_0,
    i_8_227_172_0, i_8_227_173_0, i_8_227_269_0, i_8_227_284_0,
    i_8_227_293_0, i_8_227_323_0, i_8_227_353_0, i_8_227_360_0,
    i_8_227_368_0, i_8_227_382_0, i_8_227_398_0, i_8_227_452_0,
    i_8_227_489_0, i_8_227_490_0, i_8_227_492_0, i_8_227_530_0,
    i_8_227_590_0, i_8_227_614_0, i_8_227_634_0, i_8_227_706_0,
    i_8_227_707_0, i_8_227_764_0, i_8_227_797_0, i_8_227_833_0,
    i_8_227_845_0, i_8_227_858_0, i_8_227_859_0, i_8_227_868_0,
    i_8_227_922_0, i_8_227_969_0, i_8_227_1057_0, i_8_227_1058_0,
    i_8_227_1073_0, i_8_227_1100_0, i_8_227_1127_0, i_8_227_1129_0,
    i_8_227_1225_0, i_8_227_1226_0, i_8_227_1229_0, i_8_227_1262_0,
    i_8_227_1264_0, i_8_227_1298_0, i_8_227_1317_0, i_8_227_1325_0,
    i_8_227_1328_0, i_8_227_1366_0, i_8_227_1405_0, i_8_227_1406_0,
    i_8_227_1411_0, i_8_227_1435_0, i_8_227_1436_0, i_8_227_1456_0,
    i_8_227_1462_0, i_8_227_1463_0, i_8_227_1473_0, i_8_227_1522_0,
    i_8_227_1547_0, i_8_227_1549_0, i_8_227_1556_0, i_8_227_1622_0,
    i_8_227_1623_0, i_8_227_1633_0, i_8_227_1640_0, i_8_227_1730_0,
    i_8_227_1748_0, i_8_227_1757_0, i_8_227_1777_0, i_8_227_1784_0,
    i_8_227_1796_0, i_8_227_1823_0, i_8_227_1825_0, i_8_227_1832_0,
    i_8_227_1849_0, i_8_227_1867_0, i_8_227_1904_0, i_8_227_1957_0,
    i_8_227_1958_0, i_8_227_1975_0, i_8_227_1994_0, i_8_227_1996_0,
    i_8_227_1997_0, i_8_227_2003_0, i_8_227_2017_0, i_8_227_2020_0,
    i_8_227_2099_0, i_8_227_2117_0, i_8_227_2144_0, i_8_227_2150_0,
    i_8_227_2201_0, i_8_227_2225_0, i_8_227_2226_0, i_8_227_2244_0,
    i_8_227_2246_0, i_8_227_2249_0, i_8_227_2260_0, i_8_227_2287_0;
  output o_8_227_0_0;
  assign o_8_227_0_0 = 0;
endmodule



// Benchmark "kernel_8_228" written by ABC on Sun Jul 19 10:07:01 2020

module kernel_8_228 ( 
    i_8_228_21_0, i_8_228_25_0, i_8_228_44_0, i_8_228_79_0, i_8_228_84_0,
    i_8_228_247_0, i_8_228_248_0, i_8_228_265_0, i_8_228_320_0,
    i_8_228_323_0, i_8_228_338_0, i_8_228_367_0, i_8_228_368_0,
    i_8_228_395_0, i_8_228_422_0, i_8_228_430_0, i_8_228_469_0,
    i_8_228_511_0, i_8_228_516_0, i_8_228_517_0, i_8_228_527_0,
    i_8_228_552_0, i_8_228_571_0, i_8_228_574_0, i_8_228_575_0,
    i_8_228_584_0, i_8_228_591_0, i_8_228_593_0, i_8_228_597_0,
    i_8_228_599_0, i_8_228_611_0, i_8_228_634_0, i_8_228_647_0,
    i_8_228_683_0, i_8_228_704_0, i_8_228_710_0, i_8_228_733_0,
    i_8_228_763_0, i_8_228_788_0, i_8_228_824_0, i_8_228_832_0,
    i_8_228_842_0, i_8_228_858_0, i_8_228_861_0, i_8_228_941_0,
    i_8_228_971_0, i_8_228_1016_0, i_8_228_1106_0, i_8_228_1114_0,
    i_8_228_1129_0, i_8_228_1189_0, i_8_228_1205_0, i_8_228_1240_0,
    i_8_228_1267_0, i_8_228_1300_0, i_8_228_1304_0, i_8_228_1305_0,
    i_8_228_1366_0, i_8_228_1367_0, i_8_228_1403_0, i_8_228_1408_0,
    i_8_228_1410_0, i_8_228_1465_0, i_8_228_1466_0, i_8_228_1516_0,
    i_8_228_1517_0, i_8_228_1528_0, i_8_228_1533_0, i_8_228_1540_0,
    i_8_228_1588_0, i_8_228_1591_0, i_8_228_1653_0, i_8_228_1654_0,
    i_8_228_1691_0, i_8_228_1700_0, i_8_228_1750_0, i_8_228_1843_0,
    i_8_228_1844_0, i_8_228_1857_0, i_8_228_1868_0, i_8_228_1873_0,
    i_8_228_1876_0, i_8_228_1878_0, i_8_228_1886_0, i_8_228_1898_0,
    i_8_228_1916_0, i_8_228_1917_0, i_8_228_2011_0, i_8_228_2040_0,
    i_8_228_2048_0, i_8_228_2065_0, i_8_228_2128_0, i_8_228_2163_0,
    i_8_228_2173_0, i_8_228_2214_0, i_8_228_2231_0, i_8_228_2244_0,
    i_8_228_2245_0, i_8_228_2290_0, i_8_228_2298_0,
    o_8_228_0_0  );
  input  i_8_228_21_0, i_8_228_25_0, i_8_228_44_0, i_8_228_79_0,
    i_8_228_84_0, i_8_228_247_0, i_8_228_248_0, i_8_228_265_0,
    i_8_228_320_0, i_8_228_323_0, i_8_228_338_0, i_8_228_367_0,
    i_8_228_368_0, i_8_228_395_0, i_8_228_422_0, i_8_228_430_0,
    i_8_228_469_0, i_8_228_511_0, i_8_228_516_0, i_8_228_517_0,
    i_8_228_527_0, i_8_228_552_0, i_8_228_571_0, i_8_228_574_0,
    i_8_228_575_0, i_8_228_584_0, i_8_228_591_0, i_8_228_593_0,
    i_8_228_597_0, i_8_228_599_0, i_8_228_611_0, i_8_228_634_0,
    i_8_228_647_0, i_8_228_683_0, i_8_228_704_0, i_8_228_710_0,
    i_8_228_733_0, i_8_228_763_0, i_8_228_788_0, i_8_228_824_0,
    i_8_228_832_0, i_8_228_842_0, i_8_228_858_0, i_8_228_861_0,
    i_8_228_941_0, i_8_228_971_0, i_8_228_1016_0, i_8_228_1106_0,
    i_8_228_1114_0, i_8_228_1129_0, i_8_228_1189_0, i_8_228_1205_0,
    i_8_228_1240_0, i_8_228_1267_0, i_8_228_1300_0, i_8_228_1304_0,
    i_8_228_1305_0, i_8_228_1366_0, i_8_228_1367_0, i_8_228_1403_0,
    i_8_228_1408_0, i_8_228_1410_0, i_8_228_1465_0, i_8_228_1466_0,
    i_8_228_1516_0, i_8_228_1517_0, i_8_228_1528_0, i_8_228_1533_0,
    i_8_228_1540_0, i_8_228_1588_0, i_8_228_1591_0, i_8_228_1653_0,
    i_8_228_1654_0, i_8_228_1691_0, i_8_228_1700_0, i_8_228_1750_0,
    i_8_228_1843_0, i_8_228_1844_0, i_8_228_1857_0, i_8_228_1868_0,
    i_8_228_1873_0, i_8_228_1876_0, i_8_228_1878_0, i_8_228_1886_0,
    i_8_228_1898_0, i_8_228_1916_0, i_8_228_1917_0, i_8_228_2011_0,
    i_8_228_2040_0, i_8_228_2048_0, i_8_228_2065_0, i_8_228_2128_0,
    i_8_228_2163_0, i_8_228_2173_0, i_8_228_2214_0, i_8_228_2231_0,
    i_8_228_2244_0, i_8_228_2245_0, i_8_228_2290_0, i_8_228_2298_0;
  output o_8_228_0_0;
  assign o_8_228_0_0 = 0;
endmodule



// Benchmark "kernel_8_229" written by ABC on Sun Jul 19 10:07:02 2020

module kernel_8_229 ( 
    i_8_229_40_0, i_8_229_59_0, i_8_229_64_0, i_8_229_83_0, i_8_229_104_0,
    i_8_229_140_0, i_8_229_163_0, i_8_229_220_0, i_8_229_221_0,
    i_8_229_229_0, i_8_229_247_0, i_8_229_281_0, i_8_229_283_0,
    i_8_229_326_0, i_8_229_363_0, i_8_229_364_0, i_8_229_381_0,
    i_8_229_434_0, i_8_229_451_0, i_8_229_481_0, i_8_229_487_0,
    i_8_229_504_0, i_8_229_505_0, i_8_229_522_0, i_8_229_524_0,
    i_8_229_526_0, i_8_229_527_0, i_8_229_528_0, i_8_229_589_0,
    i_8_229_594_0, i_8_229_598_0, i_8_229_609_0, i_8_229_610_0,
    i_8_229_623_0, i_8_229_659_0, i_8_229_662_0, i_8_229_685_0,
    i_8_229_689_0, i_8_229_694_0, i_8_229_696_0, i_8_229_706_0,
    i_8_229_716_0, i_8_229_725_0, i_8_229_760_0, i_8_229_823_0,
    i_8_229_838_0, i_8_229_845_0, i_8_229_996_0, i_8_229_1072_0,
    i_8_229_1100_0, i_8_229_1103_0, i_8_229_1180_0, i_8_229_1225_0,
    i_8_229_1234_0, i_8_229_1300_0, i_8_229_1309_0, i_8_229_1310_0,
    i_8_229_1352_0, i_8_229_1434_0, i_8_229_1438_0, i_8_229_1439_0,
    i_8_229_1589_0, i_8_229_1616_0, i_8_229_1625_0, i_8_229_1643_0,
    i_8_229_1674_0, i_8_229_1682_0, i_8_229_1720_0, i_8_229_1751_0,
    i_8_229_1752_0, i_8_229_1753_0, i_8_229_1771_0, i_8_229_1778_0,
    i_8_229_1810_0, i_8_229_1840_0, i_8_229_1856_0, i_8_229_1885_0,
    i_8_229_1901_0, i_8_229_1936_0, i_8_229_1949_0, i_8_229_1950_0,
    i_8_229_1968_0, i_8_229_1969_0, i_8_229_1990_0, i_8_229_2029_0,
    i_8_229_2041_0, i_8_229_2068_0, i_8_229_2089_0, i_8_229_2092_0,
    i_8_229_2129_0, i_8_229_2152_0, i_8_229_2153_0, i_8_229_2171_0,
    i_8_229_2173_0, i_8_229_2236_0, i_8_229_2237_0, i_8_229_2241_0,
    i_8_229_2246_0, i_8_229_2260_0, i_8_229_2261_0,
    o_8_229_0_0  );
  input  i_8_229_40_0, i_8_229_59_0, i_8_229_64_0, i_8_229_83_0,
    i_8_229_104_0, i_8_229_140_0, i_8_229_163_0, i_8_229_220_0,
    i_8_229_221_0, i_8_229_229_0, i_8_229_247_0, i_8_229_281_0,
    i_8_229_283_0, i_8_229_326_0, i_8_229_363_0, i_8_229_364_0,
    i_8_229_381_0, i_8_229_434_0, i_8_229_451_0, i_8_229_481_0,
    i_8_229_487_0, i_8_229_504_0, i_8_229_505_0, i_8_229_522_0,
    i_8_229_524_0, i_8_229_526_0, i_8_229_527_0, i_8_229_528_0,
    i_8_229_589_0, i_8_229_594_0, i_8_229_598_0, i_8_229_609_0,
    i_8_229_610_0, i_8_229_623_0, i_8_229_659_0, i_8_229_662_0,
    i_8_229_685_0, i_8_229_689_0, i_8_229_694_0, i_8_229_696_0,
    i_8_229_706_0, i_8_229_716_0, i_8_229_725_0, i_8_229_760_0,
    i_8_229_823_0, i_8_229_838_0, i_8_229_845_0, i_8_229_996_0,
    i_8_229_1072_0, i_8_229_1100_0, i_8_229_1103_0, i_8_229_1180_0,
    i_8_229_1225_0, i_8_229_1234_0, i_8_229_1300_0, i_8_229_1309_0,
    i_8_229_1310_0, i_8_229_1352_0, i_8_229_1434_0, i_8_229_1438_0,
    i_8_229_1439_0, i_8_229_1589_0, i_8_229_1616_0, i_8_229_1625_0,
    i_8_229_1643_0, i_8_229_1674_0, i_8_229_1682_0, i_8_229_1720_0,
    i_8_229_1751_0, i_8_229_1752_0, i_8_229_1753_0, i_8_229_1771_0,
    i_8_229_1778_0, i_8_229_1810_0, i_8_229_1840_0, i_8_229_1856_0,
    i_8_229_1885_0, i_8_229_1901_0, i_8_229_1936_0, i_8_229_1949_0,
    i_8_229_1950_0, i_8_229_1968_0, i_8_229_1969_0, i_8_229_1990_0,
    i_8_229_2029_0, i_8_229_2041_0, i_8_229_2068_0, i_8_229_2089_0,
    i_8_229_2092_0, i_8_229_2129_0, i_8_229_2152_0, i_8_229_2153_0,
    i_8_229_2171_0, i_8_229_2173_0, i_8_229_2236_0, i_8_229_2237_0,
    i_8_229_2241_0, i_8_229_2246_0, i_8_229_2260_0, i_8_229_2261_0;
  output o_8_229_0_0;
  assign o_8_229_0_0 = 0;
endmodule



// Benchmark "kernel_8_230" written by ABC on Sun Jul 19 10:07:04 2020

module kernel_8_230 ( 
    i_8_230_43_0, i_8_230_96_0, i_8_230_114_0, i_8_230_140_0,
    i_8_230_143_0, i_8_230_156_0, i_8_230_158_0, i_8_230_185_0,
    i_8_230_188_0, i_8_230_217_0, i_8_230_218_0, i_8_230_224_0,
    i_8_230_227_0, i_8_230_253_0, i_8_230_301_0, i_8_230_329_0,
    i_8_230_414_0, i_8_230_461_0, i_8_230_482_0, i_8_230_485_0,
    i_8_230_489_0, i_8_230_496_0, i_8_230_505_0, i_8_230_522_0,
    i_8_230_523_0, i_8_230_524_0, i_8_230_525_0, i_8_230_528_0,
    i_8_230_530_0, i_8_230_592_0, i_8_230_609_0, i_8_230_614_0,
    i_8_230_624_0, i_8_230_630_0, i_8_230_632_0, i_8_230_661_0,
    i_8_230_696_0, i_8_230_697_0, i_8_230_700_0, i_8_230_701_0,
    i_8_230_711_0, i_8_230_713_0, i_8_230_714_0, i_8_230_715_0,
    i_8_230_716_0, i_8_230_719_0, i_8_230_768_0, i_8_230_812_0,
    i_8_230_837_0, i_8_230_839_0, i_8_230_840_0, i_8_230_1012_0,
    i_8_230_1121_0, i_8_230_1180_0, i_8_230_1181_0, i_8_230_1263_0,
    i_8_230_1284_0, i_8_230_1286_0, i_8_230_1297_0, i_8_230_1346_0,
    i_8_230_1382_0, i_8_230_1407_0, i_8_230_1411_0, i_8_230_1412_0,
    i_8_230_1504_0, i_8_230_1506_0, i_8_230_1624_0, i_8_230_1649_0,
    i_8_230_1651_0, i_8_230_1652_0, i_8_230_1655_0, i_8_230_1678_0,
    i_8_230_1747_0, i_8_230_1748_0, i_8_230_1749_0, i_8_230_1754_0,
    i_8_230_1825_0, i_8_230_1855_0, i_8_230_1881_0, i_8_230_1882_0,
    i_8_230_1901_0, i_8_230_1903_0, i_8_230_1981_0, i_8_230_1985_0,
    i_8_230_1992_0, i_8_230_1997_0, i_8_230_1999_0, i_8_230_2031_0,
    i_8_230_2037_0, i_8_230_2053_0, i_8_230_2056_0, i_8_230_2057_0,
    i_8_230_2089_0, i_8_230_2090_0, i_8_230_2143_0, i_8_230_2144_0,
    i_8_230_2150_0, i_8_230_2174_0, i_8_230_2218_0, i_8_230_2246_0,
    o_8_230_0_0  );
  input  i_8_230_43_0, i_8_230_96_0, i_8_230_114_0, i_8_230_140_0,
    i_8_230_143_0, i_8_230_156_0, i_8_230_158_0, i_8_230_185_0,
    i_8_230_188_0, i_8_230_217_0, i_8_230_218_0, i_8_230_224_0,
    i_8_230_227_0, i_8_230_253_0, i_8_230_301_0, i_8_230_329_0,
    i_8_230_414_0, i_8_230_461_0, i_8_230_482_0, i_8_230_485_0,
    i_8_230_489_0, i_8_230_496_0, i_8_230_505_0, i_8_230_522_0,
    i_8_230_523_0, i_8_230_524_0, i_8_230_525_0, i_8_230_528_0,
    i_8_230_530_0, i_8_230_592_0, i_8_230_609_0, i_8_230_614_0,
    i_8_230_624_0, i_8_230_630_0, i_8_230_632_0, i_8_230_661_0,
    i_8_230_696_0, i_8_230_697_0, i_8_230_700_0, i_8_230_701_0,
    i_8_230_711_0, i_8_230_713_0, i_8_230_714_0, i_8_230_715_0,
    i_8_230_716_0, i_8_230_719_0, i_8_230_768_0, i_8_230_812_0,
    i_8_230_837_0, i_8_230_839_0, i_8_230_840_0, i_8_230_1012_0,
    i_8_230_1121_0, i_8_230_1180_0, i_8_230_1181_0, i_8_230_1263_0,
    i_8_230_1284_0, i_8_230_1286_0, i_8_230_1297_0, i_8_230_1346_0,
    i_8_230_1382_0, i_8_230_1407_0, i_8_230_1411_0, i_8_230_1412_0,
    i_8_230_1504_0, i_8_230_1506_0, i_8_230_1624_0, i_8_230_1649_0,
    i_8_230_1651_0, i_8_230_1652_0, i_8_230_1655_0, i_8_230_1678_0,
    i_8_230_1747_0, i_8_230_1748_0, i_8_230_1749_0, i_8_230_1754_0,
    i_8_230_1825_0, i_8_230_1855_0, i_8_230_1881_0, i_8_230_1882_0,
    i_8_230_1901_0, i_8_230_1903_0, i_8_230_1981_0, i_8_230_1985_0,
    i_8_230_1992_0, i_8_230_1997_0, i_8_230_1999_0, i_8_230_2031_0,
    i_8_230_2037_0, i_8_230_2053_0, i_8_230_2056_0, i_8_230_2057_0,
    i_8_230_2089_0, i_8_230_2090_0, i_8_230_2143_0, i_8_230_2144_0,
    i_8_230_2150_0, i_8_230_2174_0, i_8_230_2218_0, i_8_230_2246_0;
  output o_8_230_0_0;
  assign o_8_230_0_0 = ~((~i_8_230_96_0 & ((i_8_230_114_0 & ((~i_8_230_414_0 & ~i_8_230_496_0 & ~i_8_230_714_0 & ~i_8_230_716_0 & ~i_8_230_768_0 & ~i_8_230_839_0 & ~i_8_230_1649_0) | (~i_8_230_217_0 & ~i_8_230_1749_0 & ~i_8_230_1754_0 & ~i_8_230_2089_0))) | (~i_8_230_2218_0 & ((~i_8_230_143_0 & ~i_8_230_1747_0 & ~i_8_230_2090_0 & ((~i_8_230_156_0 & ~i_8_230_218_0 & ~i_8_230_301_0 & ~i_8_230_414_0 & ~i_8_230_530_0 & ~i_8_230_661_0 & ~i_8_230_713_0 & ~i_8_230_716_0 & ~i_8_230_719_0 & ~i_8_230_1504_0 & ~i_8_230_2037_0 & ~i_8_230_2057_0) | (~i_8_230_224_0 & ~i_8_230_496_0 & ~i_8_230_523_0 & ~i_8_230_711_0 & ~i_8_230_768_0 & i_8_230_1263_0 & ~i_8_230_1749_0 & ~i_8_230_1903_0 & ~i_8_230_2031_0 & ~i_8_230_2089_0))) | (~i_8_230_156_0 & ~i_8_230_485_0 & ~i_8_230_496_0 & ~i_8_230_522_0 & ~i_8_230_523_0 & ~i_8_230_711_0 & ~i_8_230_713_0 & ~i_8_230_714_0 & ~i_8_230_716_0 & ~i_8_230_1754_0))) | (~i_8_230_414_0 & ~i_8_230_2031_0 & ((~i_8_230_624_0 & ((~i_8_230_329_0 & ~i_8_230_505_0 & ~i_8_230_614_0 & ~i_8_230_1286_0 & i_8_230_1407_0) | (~i_8_230_43_0 & ~i_8_230_140_0 & ~i_8_230_485_0 & ~i_8_230_524_0 & ~i_8_230_632_0 & ~i_8_230_711_0 & ~i_8_230_768_0 & ~i_8_230_812_0 & ~i_8_230_1012_0 & ~i_8_230_1506_0 & ~i_8_230_1748_0 & ~i_8_230_1754_0 & ~i_8_230_2057_0))) | (~i_8_230_224_0 & ~i_8_230_714_0 & ~i_8_230_719_0 & ~i_8_230_1263_0 & ~i_8_230_1346_0 & i_8_230_2053_0 & ~i_8_230_2057_0))) | (~i_8_230_158_0 & ~i_8_230_218_0 & ~i_8_230_714_0 & ~i_8_230_1506_0 & ~i_8_230_1999_0 & i_8_230_2056_0 & i_8_230_2057_0))) | (~i_8_230_218_0 & ((~i_8_230_140_0 & ~i_8_230_156_0 & ~i_8_230_301_0 & ~i_8_230_414_0 & ~i_8_230_482_0 & ~i_8_230_522_0 & ~i_8_230_528_0 & ~i_8_230_715_0 & ~i_8_230_719_0 & ~i_8_230_1346_0 & ~i_8_230_1506_0 & ~i_8_230_1747_0) | (~i_8_230_188_0 & ~i_8_230_524_0 & ~i_8_230_592_0 & ~i_8_230_1903_0 & i_8_230_2246_0))) | (~i_8_230_253_0 & ((~i_8_230_414_0 & i_8_230_696_0 & i_8_230_711_0 & ~i_8_230_840_0 & i_8_230_1882_0) | (~i_8_230_188_0 & i_8_230_632_0 & ~i_8_230_711_0 & ~i_8_230_715_0 & ~i_8_230_1901_0))) | (~i_8_230_301_0 & ((~i_8_230_227_0 & ~i_8_230_711_0 & ~i_8_230_714_0 & ~i_8_230_768_0 & ~i_8_230_1748_0 & i_8_230_1749_0 & ~i_8_230_1754_0 & ~i_8_230_1903_0) | (~i_8_230_485_0 & i_8_230_489_0 & i_8_230_1407_0 & i_8_230_2089_0))) | (~i_8_230_329_0 & ((~i_8_230_143_0 & ~i_8_230_156_0 & ~i_8_230_158_0 & i_8_230_1655_0 & ~i_8_230_1981_0) | (~i_8_230_482_0 & ~i_8_230_528_0 & ~i_8_230_715_0 & ~i_8_230_716_0 & ~i_8_230_1346_0 & ~i_8_230_1412_0 & ~i_8_230_1747_0 & i_8_230_1754_0 & ~i_8_230_2056_0 & ~i_8_230_2218_0))) | (~i_8_230_482_0 & ((~i_8_230_143_0 & ((~i_8_230_158_0 & ~i_8_230_524_0 & i_8_230_592_0 & ~i_8_230_715_0 & i_8_230_719_0 & ~i_8_230_1749_0 & ~i_8_230_2056_0) | (~i_8_230_217_0 & ~i_8_230_711_0 & ~i_8_230_719_0 & i_8_230_1997_0 & ~i_8_230_2057_0))) | (~i_8_230_711_0 & ((~i_8_230_156_0 & i_8_230_614_0 & ~i_8_230_624_0 & ~i_8_230_2057_0) | (~i_8_230_505_0 & i_8_230_700_0 & ~i_8_230_1412_0 & ~i_8_230_1749_0 & ~i_8_230_2090_0))) | (~i_8_230_485_0 & ~i_8_230_696_0 & ~i_8_230_714_0 & ~i_8_230_1346_0 & ~i_8_230_1747_0 & ~i_8_230_2090_0 & i_8_230_2143_0 & ~i_8_230_2174_0))) | (~i_8_230_768_0 & ((~i_8_230_140_0 & ((~i_8_230_217_0 & ~i_8_230_224_0 & ~i_8_230_525_0 & ~i_8_230_530_0 & ~i_8_230_624_0 & ~i_8_230_713_0 & ~i_8_230_714_0 & ~i_8_230_1747_0 & ~i_8_230_2031_0 & ~i_8_230_2089_0) | (~i_8_230_485_0 & i_8_230_839_0 & ~i_8_230_1749_0 & i_8_230_2090_0))) | (~i_8_230_158_0 & ((~i_8_230_496_0 & ~i_8_230_524_0 & ~i_8_230_711_0 & ~i_8_230_719_0 & i_8_230_839_0) | (~i_8_230_485_0 & i_8_230_1411_0 & ~i_8_230_1747_0 & ~i_8_230_1749_0 & ~i_8_230_2031_0 & ~i_8_230_2090_0))) | (~i_8_230_217_0 & ((i_8_230_697_0 & i_8_230_700_0) | (~i_8_230_461_0 & ~i_8_230_661_0 & ~i_8_230_714_0 & ~i_8_230_719_0 & i_8_230_1263_0 & ~i_8_230_1649_0))) | (~i_8_230_530_0 & i_8_230_840_0 & i_8_230_1825_0) | (~i_8_230_114_0 & i_8_230_489_0 & ~i_8_230_523_0 & ~i_8_230_614_0 & ~i_8_230_2031_0 & ~i_8_230_2090_0 & ~i_8_230_711_0 & ~i_8_230_716_0))) | (~i_8_230_224_0 & ((~i_8_230_592_0 & ~i_8_230_715_0 & i_8_230_1412_0 & ~i_8_230_1754_0) | (~i_8_230_485_0 & ~i_8_230_496_0 & ~i_8_230_713_0 & ~i_8_230_714_0 & ~i_8_230_716_0 & ~i_8_230_1506_0 & ~i_8_230_1747_0 & ~i_8_230_1748_0 & ~i_8_230_2031_0 & ~i_8_230_2089_0 & ~i_8_230_2218_0))) | (~i_8_230_485_0 & ((~i_8_230_489_0 & ~i_8_230_523_0 & i_8_230_592_0 & ~i_8_230_840_0 & i_8_230_1825_0) | (~i_8_230_43_0 & ~i_8_230_140_0 & ~i_8_230_505_0 & ~i_8_230_525_0 & ~i_8_230_614_0 & ~i_8_230_661_0 & ~i_8_230_700_0 & ~i_8_230_713_0 & ~i_8_230_839_0 & ~i_8_230_1411_0 & ~i_8_230_1678_0 & ~i_8_230_1749_0 & ~i_8_230_1985_0 & ~i_8_230_1997_0 & ~i_8_230_2031_0))) | (~i_8_230_2090_0 & ((~i_8_230_43_0 & ((~i_8_230_217_0 & ~i_8_230_522_0 & ~i_8_230_525_0 & ~i_8_230_716_0 & i_8_230_1284_0 & ~i_8_230_1506_0) | (~i_8_230_188_0 & i_8_230_530_0 & ~i_8_230_713_0 & i_8_230_1286_0 & ~i_8_230_1346_0 & ~i_8_230_1903_0))) | (~i_8_230_525_0 & ~i_8_230_661_0 & ~i_8_230_1121_0 & ~i_8_230_1382_0 & ~i_8_230_1855_0 & i_8_230_1981_0 & ~i_8_230_2246_0))) | (~i_8_230_188_0 & ((~i_8_230_489_0 & ~i_8_230_523_0 & ~i_8_230_715_0 & i_8_230_839_0 & ~i_8_230_1263_0 & ~i_8_230_1985_0) | (~i_8_230_530_0 & i_8_230_696_0 & ~i_8_230_1992_0 & i_8_230_2037_0))) | (~i_8_230_713_0 & ((~i_8_230_530_0 & ~i_8_230_2089_0 & ((i_8_230_701_0 & ~i_8_230_715_0) | (~i_8_230_624_0 & ~i_8_230_1506_0 & ~i_8_230_1855_0 & i_8_230_1992_0 & ~i_8_230_2218_0))) | (~i_8_230_43_0 & ~i_8_230_1121_0 & i_8_230_1297_0 & i_8_230_2143_0 & ~i_8_230_2174_0))) | (~i_8_230_716_0 & ((i_8_230_485_0 & ~i_8_230_1346_0 & ~i_8_230_1504_0 & i_8_230_1655_0) | (~i_8_230_715_0 & i_8_230_1181_0 & ~i_8_230_1649_0 & ~i_8_230_1855_0))) | (~i_8_230_156_0 & i_8_230_696_0 & ~i_8_230_839_0 & i_8_230_840_0 & ~i_8_230_1504_0 & ~i_8_230_2031_0 & ~i_8_230_2053_0));
endmodule



// Benchmark "kernel_8_231" written by ABC on Sun Jul 19 10:07:05 2020

module kernel_8_231 ( 
    i_8_231_27_0, i_8_231_28_0, i_8_231_49_0, i_8_231_70_0, i_8_231_94_0,
    i_8_231_147_0, i_8_231_166_0, i_8_231_184_0, i_8_231_196_0,
    i_8_231_233_0, i_8_231_241_0, i_8_231_311_0, i_8_231_322_0,
    i_8_231_337_0, i_8_231_346_0, i_8_231_381_0, i_8_231_431_0,
    i_8_231_447_0, i_8_231_454_0, i_8_231_492_0, i_8_231_493_0,
    i_8_231_570_0, i_8_231_583_0, i_8_231_609_0, i_8_231_610_0,
    i_8_231_634_0, i_8_231_659_0, i_8_231_699_0, i_8_231_701_0,
    i_8_231_732_0, i_8_231_735_0, i_8_231_753_0, i_8_231_777_0,
    i_8_231_798_0, i_8_231_799_0, i_8_231_834_0, i_8_231_835_0,
    i_8_231_843_0, i_8_231_925_0, i_8_231_931_0, i_8_231_959_0,
    i_8_231_967_0, i_8_231_973_0, i_8_231_990_0, i_8_231_991_0,
    i_8_231_1020_0, i_8_231_1033_0, i_8_231_1059_0, i_8_231_1060_0,
    i_8_231_1102_0, i_8_231_1156_0, i_8_231_1236_0, i_8_231_1237_0,
    i_8_231_1263_0, i_8_231_1273_0, i_8_231_1296_0, i_8_231_1300_0,
    i_8_231_1373_0, i_8_231_1381_0, i_8_231_1407_0, i_8_231_1474_0,
    i_8_231_1488_0, i_8_231_1489_0, i_8_231_1491_0, i_8_231_1501_0,
    i_8_231_1564_0, i_8_231_1605_0, i_8_231_1606_0, i_8_231_1627_0,
    i_8_231_1628_0, i_8_231_1650_0, i_8_231_1661_0, i_8_231_1681_0,
    i_8_231_1705_0, i_8_231_1722_0, i_8_231_1758_0, i_8_231_1770_0,
    i_8_231_1826_0, i_8_231_1857_0, i_8_231_1884_0, i_8_231_1906_0,
    i_8_231_1969_0, i_8_231_2002_0, i_8_231_2004_0, i_8_231_2016_0,
    i_8_231_2046_0, i_8_231_2047_0, i_8_231_2102_0, i_8_231_2112_0,
    i_8_231_2145_0, i_8_231_2149_0, i_8_231_2163_0, i_8_231_2167_0,
    i_8_231_2173_0, i_8_231_2174_0, i_8_231_2208_0, i_8_231_2275_0,
    i_8_231_2281_0, i_8_231_2289_0, i_8_231_2298_0,
    o_8_231_0_0  );
  input  i_8_231_27_0, i_8_231_28_0, i_8_231_49_0, i_8_231_70_0,
    i_8_231_94_0, i_8_231_147_0, i_8_231_166_0, i_8_231_184_0,
    i_8_231_196_0, i_8_231_233_0, i_8_231_241_0, i_8_231_311_0,
    i_8_231_322_0, i_8_231_337_0, i_8_231_346_0, i_8_231_381_0,
    i_8_231_431_0, i_8_231_447_0, i_8_231_454_0, i_8_231_492_0,
    i_8_231_493_0, i_8_231_570_0, i_8_231_583_0, i_8_231_609_0,
    i_8_231_610_0, i_8_231_634_0, i_8_231_659_0, i_8_231_699_0,
    i_8_231_701_0, i_8_231_732_0, i_8_231_735_0, i_8_231_753_0,
    i_8_231_777_0, i_8_231_798_0, i_8_231_799_0, i_8_231_834_0,
    i_8_231_835_0, i_8_231_843_0, i_8_231_925_0, i_8_231_931_0,
    i_8_231_959_0, i_8_231_967_0, i_8_231_973_0, i_8_231_990_0,
    i_8_231_991_0, i_8_231_1020_0, i_8_231_1033_0, i_8_231_1059_0,
    i_8_231_1060_0, i_8_231_1102_0, i_8_231_1156_0, i_8_231_1236_0,
    i_8_231_1237_0, i_8_231_1263_0, i_8_231_1273_0, i_8_231_1296_0,
    i_8_231_1300_0, i_8_231_1373_0, i_8_231_1381_0, i_8_231_1407_0,
    i_8_231_1474_0, i_8_231_1488_0, i_8_231_1489_0, i_8_231_1491_0,
    i_8_231_1501_0, i_8_231_1564_0, i_8_231_1605_0, i_8_231_1606_0,
    i_8_231_1627_0, i_8_231_1628_0, i_8_231_1650_0, i_8_231_1661_0,
    i_8_231_1681_0, i_8_231_1705_0, i_8_231_1722_0, i_8_231_1758_0,
    i_8_231_1770_0, i_8_231_1826_0, i_8_231_1857_0, i_8_231_1884_0,
    i_8_231_1906_0, i_8_231_1969_0, i_8_231_2002_0, i_8_231_2004_0,
    i_8_231_2016_0, i_8_231_2046_0, i_8_231_2047_0, i_8_231_2102_0,
    i_8_231_2112_0, i_8_231_2145_0, i_8_231_2149_0, i_8_231_2163_0,
    i_8_231_2167_0, i_8_231_2173_0, i_8_231_2174_0, i_8_231_2208_0,
    i_8_231_2275_0, i_8_231_2281_0, i_8_231_2289_0, i_8_231_2298_0;
  output o_8_231_0_0;
  assign o_8_231_0_0 = 0;
endmodule



// Benchmark "kernel_8_232" written by ABC on Sun Jul 19 10:07:06 2020

module kernel_8_232 ( 
    i_8_232_22_0, i_8_232_23_0, i_8_232_31_0, i_8_232_34_0, i_8_232_35_0,
    i_8_232_85_0, i_8_232_106_0, i_8_232_107_0, i_8_232_232_0,
    i_8_232_247_0, i_8_232_295_0, i_8_232_345_0, i_8_232_346_0,
    i_8_232_348_0, i_8_232_386_0, i_8_232_394_0, i_8_232_426_0,
    i_8_232_443_0, i_8_232_458_0, i_8_232_480_0, i_8_232_482_0,
    i_8_232_524_0, i_8_232_526_0, i_8_232_527_0, i_8_232_529_0,
    i_8_232_554_0, i_8_232_555_0, i_8_232_602_0, i_8_232_609_0,
    i_8_232_611_0, i_8_232_628_0, i_8_232_631_0, i_8_232_633_0,
    i_8_232_634_0, i_8_232_707_0, i_8_232_732_0, i_8_232_761_0,
    i_8_232_763_0, i_8_232_771_0, i_8_232_783_0, i_8_232_799_0,
    i_8_232_800_0, i_8_232_811_0, i_8_232_814_0, i_8_232_815_0,
    i_8_232_838_0, i_8_232_931_0, i_8_232_934_0, i_8_232_965_0,
    i_8_232_986_0, i_8_232_991_0, i_8_232_1120_0, i_8_232_1189_0,
    i_8_232_1194_0, i_8_232_1219_0, i_8_232_1220_0, i_8_232_1223_0,
    i_8_232_1266_0, i_8_232_1267_0, i_8_232_1284_0, i_8_232_1311_0,
    i_8_232_1388_0, i_8_232_1391_0, i_8_232_1441_0, i_8_232_1525_0,
    i_8_232_1526_0, i_8_232_1535_0, i_8_232_1544_0, i_8_232_1545_0,
    i_8_232_1550_0, i_8_232_1554_0, i_8_232_1561_0, i_8_232_1633_0,
    i_8_232_1651_0, i_8_232_1676_0, i_8_232_1699_0, i_8_232_1722_0,
    i_8_232_1726_0, i_8_232_1733_0, i_8_232_1738_0, i_8_232_1740_0,
    i_8_232_1741_0, i_8_232_1748_0, i_8_232_1749_0, i_8_232_1753_0,
    i_8_232_1807_0, i_8_232_1819_0, i_8_232_1858_0, i_8_232_1867_0,
    i_8_232_1876_0, i_8_232_1897_0, i_8_232_1906_0, i_8_232_1956_0,
    i_8_232_1957_0, i_8_232_2150_0, i_8_232_2154_0, i_8_232_2215_0,
    i_8_232_2216_0, i_8_232_2218_0, i_8_232_2292_0,
    o_8_232_0_0  );
  input  i_8_232_22_0, i_8_232_23_0, i_8_232_31_0, i_8_232_34_0,
    i_8_232_35_0, i_8_232_85_0, i_8_232_106_0, i_8_232_107_0,
    i_8_232_232_0, i_8_232_247_0, i_8_232_295_0, i_8_232_345_0,
    i_8_232_346_0, i_8_232_348_0, i_8_232_386_0, i_8_232_394_0,
    i_8_232_426_0, i_8_232_443_0, i_8_232_458_0, i_8_232_480_0,
    i_8_232_482_0, i_8_232_524_0, i_8_232_526_0, i_8_232_527_0,
    i_8_232_529_0, i_8_232_554_0, i_8_232_555_0, i_8_232_602_0,
    i_8_232_609_0, i_8_232_611_0, i_8_232_628_0, i_8_232_631_0,
    i_8_232_633_0, i_8_232_634_0, i_8_232_707_0, i_8_232_732_0,
    i_8_232_761_0, i_8_232_763_0, i_8_232_771_0, i_8_232_783_0,
    i_8_232_799_0, i_8_232_800_0, i_8_232_811_0, i_8_232_814_0,
    i_8_232_815_0, i_8_232_838_0, i_8_232_931_0, i_8_232_934_0,
    i_8_232_965_0, i_8_232_986_0, i_8_232_991_0, i_8_232_1120_0,
    i_8_232_1189_0, i_8_232_1194_0, i_8_232_1219_0, i_8_232_1220_0,
    i_8_232_1223_0, i_8_232_1266_0, i_8_232_1267_0, i_8_232_1284_0,
    i_8_232_1311_0, i_8_232_1388_0, i_8_232_1391_0, i_8_232_1441_0,
    i_8_232_1525_0, i_8_232_1526_0, i_8_232_1535_0, i_8_232_1544_0,
    i_8_232_1545_0, i_8_232_1550_0, i_8_232_1554_0, i_8_232_1561_0,
    i_8_232_1633_0, i_8_232_1651_0, i_8_232_1676_0, i_8_232_1699_0,
    i_8_232_1722_0, i_8_232_1726_0, i_8_232_1733_0, i_8_232_1738_0,
    i_8_232_1740_0, i_8_232_1741_0, i_8_232_1748_0, i_8_232_1749_0,
    i_8_232_1753_0, i_8_232_1807_0, i_8_232_1819_0, i_8_232_1858_0,
    i_8_232_1867_0, i_8_232_1876_0, i_8_232_1897_0, i_8_232_1906_0,
    i_8_232_1956_0, i_8_232_1957_0, i_8_232_2150_0, i_8_232_2154_0,
    i_8_232_2215_0, i_8_232_2216_0, i_8_232_2218_0, i_8_232_2292_0;
  output o_8_232_0_0;
  assign o_8_232_0_0 = 0;
endmodule



// Benchmark "kernel_8_233" written by ABC on Sun Jul 19 10:07:07 2020

module kernel_8_233 ( 
    i_8_233_31_0, i_8_233_41_0, i_8_233_88_0, i_8_233_89_0, i_8_233_187_0,
    i_8_233_212_0, i_8_233_223_0, i_8_233_256_0, i_8_233_266_0,
    i_8_233_269_0, i_8_233_283_0, i_8_233_293_0, i_8_233_302_0,
    i_8_233_337_0, i_8_233_349_0, i_8_233_353_0, i_8_233_374_0,
    i_8_233_453_0, i_8_233_494_0, i_8_233_538_0, i_8_233_539_0,
    i_8_233_547_0, i_8_233_556_0, i_8_233_565_0, i_8_233_593_0,
    i_8_233_602_0, i_8_233_607_0, i_8_233_658_0, i_8_233_661_0,
    i_8_233_716_0, i_8_233_744_0, i_8_233_763_0, i_8_233_766_0,
    i_8_233_767_0, i_8_233_773_0, i_8_233_797_0, i_8_233_826_0,
    i_8_233_827_0, i_8_233_849_0, i_8_233_853_0, i_8_233_877_0,
    i_8_233_878_0, i_8_233_935_0, i_8_233_980_0, i_8_233_985_0,
    i_8_233_988_0, i_8_233_1012_0, i_8_233_1018_0, i_8_233_1030_0,
    i_8_233_1033_0, i_8_233_1041_0, i_8_233_1051_0, i_8_233_1069_0,
    i_8_233_1075_0, i_8_233_1091_0, i_8_233_1128_0, i_8_233_1129_0,
    i_8_233_1133_0, i_8_233_1139_0, i_8_233_1157_0, i_8_233_1226_0,
    i_8_233_1231_0, i_8_233_1237_0, i_8_233_1238_0, i_8_233_1249_0,
    i_8_233_1256_0, i_8_233_1262_0, i_8_233_1281_0, i_8_233_1318_0,
    i_8_233_1358_0, i_8_233_1363_0, i_8_233_1385_0, i_8_233_1453_0,
    i_8_233_1457_0, i_8_233_1543_0, i_8_233_1581_0, i_8_233_1627_0,
    i_8_233_1640_0, i_8_233_1652_0, i_8_233_1666_0, i_8_233_1700_0,
    i_8_233_1705_0, i_8_233_1708_0, i_8_233_1806_0, i_8_233_1855_0,
    i_8_233_1858_0, i_8_233_1868_0, i_8_233_1966_0, i_8_233_1995_0,
    i_8_233_1996_0, i_8_233_1997_0, i_8_233_2142_0, i_8_233_2158_0,
    i_8_233_2233_0, i_8_233_2268_0, i_8_233_2272_0, i_8_233_2273_0,
    i_8_233_2278_0, i_8_233_2282_0, i_8_233_2290_0,
    o_8_233_0_0  );
  input  i_8_233_31_0, i_8_233_41_0, i_8_233_88_0, i_8_233_89_0,
    i_8_233_187_0, i_8_233_212_0, i_8_233_223_0, i_8_233_256_0,
    i_8_233_266_0, i_8_233_269_0, i_8_233_283_0, i_8_233_293_0,
    i_8_233_302_0, i_8_233_337_0, i_8_233_349_0, i_8_233_353_0,
    i_8_233_374_0, i_8_233_453_0, i_8_233_494_0, i_8_233_538_0,
    i_8_233_539_0, i_8_233_547_0, i_8_233_556_0, i_8_233_565_0,
    i_8_233_593_0, i_8_233_602_0, i_8_233_607_0, i_8_233_658_0,
    i_8_233_661_0, i_8_233_716_0, i_8_233_744_0, i_8_233_763_0,
    i_8_233_766_0, i_8_233_767_0, i_8_233_773_0, i_8_233_797_0,
    i_8_233_826_0, i_8_233_827_0, i_8_233_849_0, i_8_233_853_0,
    i_8_233_877_0, i_8_233_878_0, i_8_233_935_0, i_8_233_980_0,
    i_8_233_985_0, i_8_233_988_0, i_8_233_1012_0, i_8_233_1018_0,
    i_8_233_1030_0, i_8_233_1033_0, i_8_233_1041_0, i_8_233_1051_0,
    i_8_233_1069_0, i_8_233_1075_0, i_8_233_1091_0, i_8_233_1128_0,
    i_8_233_1129_0, i_8_233_1133_0, i_8_233_1139_0, i_8_233_1157_0,
    i_8_233_1226_0, i_8_233_1231_0, i_8_233_1237_0, i_8_233_1238_0,
    i_8_233_1249_0, i_8_233_1256_0, i_8_233_1262_0, i_8_233_1281_0,
    i_8_233_1318_0, i_8_233_1358_0, i_8_233_1363_0, i_8_233_1385_0,
    i_8_233_1453_0, i_8_233_1457_0, i_8_233_1543_0, i_8_233_1581_0,
    i_8_233_1627_0, i_8_233_1640_0, i_8_233_1652_0, i_8_233_1666_0,
    i_8_233_1700_0, i_8_233_1705_0, i_8_233_1708_0, i_8_233_1806_0,
    i_8_233_1855_0, i_8_233_1858_0, i_8_233_1868_0, i_8_233_1966_0,
    i_8_233_1995_0, i_8_233_1996_0, i_8_233_1997_0, i_8_233_2142_0,
    i_8_233_2158_0, i_8_233_2233_0, i_8_233_2268_0, i_8_233_2272_0,
    i_8_233_2273_0, i_8_233_2278_0, i_8_233_2282_0, i_8_233_2290_0;
  output o_8_233_0_0;
  assign o_8_233_0_0 = 0;
endmodule



// Benchmark "kernel_8_234" written by ABC on Sun Jul 19 10:07:08 2020

module kernel_8_234 ( 
    i_8_234_3_0, i_8_234_4_0, i_8_234_23_0, i_8_234_31_0, i_8_234_76_0,
    i_8_234_85_0, i_8_234_86_0, i_8_234_89_0, i_8_234_116_0, i_8_234_244_0,
    i_8_234_247_0, i_8_234_265_0, i_8_234_292_0, i_8_234_301_0,
    i_8_234_322_0, i_8_234_361_0, i_8_234_366_0, i_8_234_387_0,
    i_8_234_440_0, i_8_234_463_0, i_8_234_481_0, i_8_234_516_0,
    i_8_234_517_0, i_8_234_527_0, i_8_234_538_0, i_8_234_571_0,
    i_8_234_588_0, i_8_234_594_0, i_8_234_598_0, i_8_234_599_0,
    i_8_234_611_0, i_8_234_634_0, i_8_234_642_0, i_8_234_651_0,
    i_8_234_658_0, i_8_234_669_0, i_8_234_678_0, i_8_234_727_0,
    i_8_234_778_0, i_8_234_804_0, i_8_234_823_0, i_8_234_859_0,
    i_8_234_877_0, i_8_234_913_0, i_8_234_958_0, i_8_234_1012_0,
    i_8_234_1070_0, i_8_234_1210_0, i_8_234_1228_0, i_8_234_1239_0,
    i_8_234_1270_0, i_8_234_1390_0, i_8_234_1438_0, i_8_234_1439_0,
    i_8_234_1471_0, i_8_234_1489_0, i_8_234_1517_0, i_8_234_1533_0,
    i_8_234_1534_0, i_8_234_1571_0, i_8_234_1587_0, i_8_234_1588_0,
    i_8_234_1651_0, i_8_234_1659_0, i_8_234_1679_0, i_8_234_1702_0,
    i_8_234_1703_0, i_8_234_1706_0, i_8_234_1759_0, i_8_234_1763_0,
    i_8_234_1794_0, i_8_234_1795_0, i_8_234_1798_0, i_8_234_1820_0,
    i_8_234_1821_0, i_8_234_1822_0, i_8_234_1823_0, i_8_234_1840_0,
    i_8_234_1849_0, i_8_234_1876_0, i_8_234_1885_0, i_8_234_1903_0,
    i_8_234_1918_0, i_8_234_1948_0, i_8_234_1966_0, i_8_234_1967_0,
    i_8_234_1995_0, i_8_234_2028_0, i_8_234_2037_0, i_8_234_2053_0,
    i_8_234_2065_0, i_8_234_2119_0, i_8_234_2120_0, i_8_234_2154_0,
    i_8_234_2225_0, i_8_234_2226_0, i_8_234_2229_0, i_8_234_2256_0,
    i_8_234_2257_0, i_8_234_2281_0,
    o_8_234_0_0  );
  input  i_8_234_3_0, i_8_234_4_0, i_8_234_23_0, i_8_234_31_0,
    i_8_234_76_0, i_8_234_85_0, i_8_234_86_0, i_8_234_89_0, i_8_234_116_0,
    i_8_234_244_0, i_8_234_247_0, i_8_234_265_0, i_8_234_292_0,
    i_8_234_301_0, i_8_234_322_0, i_8_234_361_0, i_8_234_366_0,
    i_8_234_387_0, i_8_234_440_0, i_8_234_463_0, i_8_234_481_0,
    i_8_234_516_0, i_8_234_517_0, i_8_234_527_0, i_8_234_538_0,
    i_8_234_571_0, i_8_234_588_0, i_8_234_594_0, i_8_234_598_0,
    i_8_234_599_0, i_8_234_611_0, i_8_234_634_0, i_8_234_642_0,
    i_8_234_651_0, i_8_234_658_0, i_8_234_669_0, i_8_234_678_0,
    i_8_234_727_0, i_8_234_778_0, i_8_234_804_0, i_8_234_823_0,
    i_8_234_859_0, i_8_234_877_0, i_8_234_913_0, i_8_234_958_0,
    i_8_234_1012_0, i_8_234_1070_0, i_8_234_1210_0, i_8_234_1228_0,
    i_8_234_1239_0, i_8_234_1270_0, i_8_234_1390_0, i_8_234_1438_0,
    i_8_234_1439_0, i_8_234_1471_0, i_8_234_1489_0, i_8_234_1517_0,
    i_8_234_1533_0, i_8_234_1534_0, i_8_234_1571_0, i_8_234_1587_0,
    i_8_234_1588_0, i_8_234_1651_0, i_8_234_1659_0, i_8_234_1679_0,
    i_8_234_1702_0, i_8_234_1703_0, i_8_234_1706_0, i_8_234_1759_0,
    i_8_234_1763_0, i_8_234_1794_0, i_8_234_1795_0, i_8_234_1798_0,
    i_8_234_1820_0, i_8_234_1821_0, i_8_234_1822_0, i_8_234_1823_0,
    i_8_234_1840_0, i_8_234_1849_0, i_8_234_1876_0, i_8_234_1885_0,
    i_8_234_1903_0, i_8_234_1918_0, i_8_234_1948_0, i_8_234_1966_0,
    i_8_234_1967_0, i_8_234_1995_0, i_8_234_2028_0, i_8_234_2037_0,
    i_8_234_2053_0, i_8_234_2065_0, i_8_234_2119_0, i_8_234_2120_0,
    i_8_234_2154_0, i_8_234_2225_0, i_8_234_2226_0, i_8_234_2229_0,
    i_8_234_2256_0, i_8_234_2257_0, i_8_234_2281_0;
  output o_8_234_0_0;
  assign o_8_234_0_0 = 0;
endmodule



// Benchmark "kernel_8_235" written by ABC on Sun Jul 19 10:07:09 2020

module kernel_8_235 ( 
    i_8_235_16_0, i_8_235_53_0, i_8_235_111_0, i_8_235_148_0,
    i_8_235_194_0, i_8_235_227_0, i_8_235_230_0, i_8_235_259_0,
    i_8_235_260_0, i_8_235_283_0, i_8_235_383_0, i_8_235_401_0,
    i_8_235_417_0, i_8_235_427_0, i_8_235_493_0, i_8_235_508_0,
    i_8_235_556_0, i_8_235_574_0, i_8_235_575_0, i_8_235_579_0,
    i_8_235_591_0, i_8_235_592_0, i_8_235_598_0, i_8_235_599_0,
    i_8_235_665_0, i_8_235_706_0, i_8_235_751_0, i_8_235_786_0,
    i_8_235_798_0, i_8_235_826_0, i_8_235_838_0, i_8_235_841_0,
    i_8_235_977_0, i_8_235_984_0, i_8_235_1101_0, i_8_235_1102_0,
    i_8_235_1105_0, i_8_235_1108_0, i_8_235_1240_0, i_8_235_1270_0,
    i_8_235_1273_0, i_8_235_1274_0, i_8_235_1302_0, i_8_235_1330_0,
    i_8_235_1384_0, i_8_235_1385_0, i_8_235_1392_0, i_8_235_1396_0,
    i_8_235_1409_0, i_8_235_1433_0, i_8_235_1437_0, i_8_235_1439_0,
    i_8_235_1464_0, i_8_235_1483_0, i_8_235_1513_0, i_8_235_1519_0,
    i_8_235_1528_0, i_8_235_1552_0, i_8_235_1573_0, i_8_235_1574_0,
    i_8_235_1605_0, i_8_235_1606_0, i_8_235_1631_0, i_8_235_1632_0,
    i_8_235_1642_0, i_8_235_1671_0, i_8_235_1696_0, i_8_235_1699_0,
    i_8_235_1704_0, i_8_235_1707_0, i_8_235_1716_0, i_8_235_1732_0,
    i_8_235_1750_0, i_8_235_1768_0, i_8_235_1770_0, i_8_235_1791_0,
    i_8_235_1807_0, i_8_235_1813_0, i_8_235_1820_0, i_8_235_1888_0,
    i_8_235_1944_0, i_8_235_1945_0, i_8_235_1950_0, i_8_235_1954_0,
    i_8_235_1957_0, i_8_235_1960_0, i_8_235_1966_0, i_8_235_1975_0,
    i_8_235_1996_0, i_8_235_2056_0, i_8_235_2059_0, i_8_235_2093_0,
    i_8_235_2096_0, i_8_235_2134_0, i_8_235_2135_0, i_8_235_2157_0,
    i_8_235_2164_0, i_8_235_2214_0, i_8_235_2219_0, i_8_235_2257_0,
    o_8_235_0_0  );
  input  i_8_235_16_0, i_8_235_53_0, i_8_235_111_0, i_8_235_148_0,
    i_8_235_194_0, i_8_235_227_0, i_8_235_230_0, i_8_235_259_0,
    i_8_235_260_0, i_8_235_283_0, i_8_235_383_0, i_8_235_401_0,
    i_8_235_417_0, i_8_235_427_0, i_8_235_493_0, i_8_235_508_0,
    i_8_235_556_0, i_8_235_574_0, i_8_235_575_0, i_8_235_579_0,
    i_8_235_591_0, i_8_235_592_0, i_8_235_598_0, i_8_235_599_0,
    i_8_235_665_0, i_8_235_706_0, i_8_235_751_0, i_8_235_786_0,
    i_8_235_798_0, i_8_235_826_0, i_8_235_838_0, i_8_235_841_0,
    i_8_235_977_0, i_8_235_984_0, i_8_235_1101_0, i_8_235_1102_0,
    i_8_235_1105_0, i_8_235_1108_0, i_8_235_1240_0, i_8_235_1270_0,
    i_8_235_1273_0, i_8_235_1274_0, i_8_235_1302_0, i_8_235_1330_0,
    i_8_235_1384_0, i_8_235_1385_0, i_8_235_1392_0, i_8_235_1396_0,
    i_8_235_1409_0, i_8_235_1433_0, i_8_235_1437_0, i_8_235_1439_0,
    i_8_235_1464_0, i_8_235_1483_0, i_8_235_1513_0, i_8_235_1519_0,
    i_8_235_1528_0, i_8_235_1552_0, i_8_235_1573_0, i_8_235_1574_0,
    i_8_235_1605_0, i_8_235_1606_0, i_8_235_1631_0, i_8_235_1632_0,
    i_8_235_1642_0, i_8_235_1671_0, i_8_235_1696_0, i_8_235_1699_0,
    i_8_235_1704_0, i_8_235_1707_0, i_8_235_1716_0, i_8_235_1732_0,
    i_8_235_1750_0, i_8_235_1768_0, i_8_235_1770_0, i_8_235_1791_0,
    i_8_235_1807_0, i_8_235_1813_0, i_8_235_1820_0, i_8_235_1888_0,
    i_8_235_1944_0, i_8_235_1945_0, i_8_235_1950_0, i_8_235_1954_0,
    i_8_235_1957_0, i_8_235_1960_0, i_8_235_1966_0, i_8_235_1975_0,
    i_8_235_1996_0, i_8_235_2056_0, i_8_235_2059_0, i_8_235_2093_0,
    i_8_235_2096_0, i_8_235_2134_0, i_8_235_2135_0, i_8_235_2157_0,
    i_8_235_2164_0, i_8_235_2214_0, i_8_235_2219_0, i_8_235_2257_0;
  output o_8_235_0_0;
  assign o_8_235_0_0 = 0;
endmodule



// Benchmark "kernel_8_236" written by ABC on Sun Jul 19 10:07:11 2020

module kernel_8_236 ( 
    i_8_236_36_0, i_8_236_37_0, i_8_236_64_0, i_8_236_112_0, i_8_236_166_0,
    i_8_236_167_0, i_8_236_193_0, i_8_236_194_0, i_8_236_221_0,
    i_8_236_226_0, i_8_236_300_0, i_8_236_362_0, i_8_236_373_0,
    i_8_236_385_0, i_8_236_397_0, i_8_236_420_0, i_8_236_421_0,
    i_8_236_484_0, i_8_236_489_0, i_8_236_493_0, i_8_236_522_0,
    i_8_236_525_0, i_8_236_526_0, i_8_236_529_0, i_8_236_606_0,
    i_8_236_607_0, i_8_236_608_0, i_8_236_613_0, i_8_236_662_0,
    i_8_236_698_0, i_8_236_700_0, i_8_236_701_0, i_8_236_707_0,
    i_8_236_710_0, i_8_236_801_0, i_8_236_802_0, i_8_236_803_0,
    i_8_236_806_0, i_8_236_809_0, i_8_236_843_0, i_8_236_844_0,
    i_8_236_854_0, i_8_236_932_0, i_8_236_935_0, i_8_236_972_0,
    i_8_236_993_0, i_8_236_995_0, i_8_236_1040_0, i_8_236_1047_0,
    i_8_236_1078_0, i_8_236_1113_0, i_8_236_1114_0, i_8_236_1115_0,
    i_8_236_1134_0, i_8_236_1233_0, i_8_236_1234_0, i_8_236_1259_0,
    i_8_236_1269_0, i_8_236_1271_0, i_8_236_1283_0, i_8_236_1286_0,
    i_8_236_1404_0, i_8_236_1489_0, i_8_236_1490_0, i_8_236_1507_0,
    i_8_236_1529_0, i_8_236_1585_0, i_8_236_1621_0, i_8_236_1624_0,
    i_8_236_1634_0, i_8_236_1650_0, i_8_236_1668_0, i_8_236_1678_0,
    i_8_236_1682_0, i_8_236_1710_0, i_8_236_1711_0, i_8_236_1748_0,
    i_8_236_1766_0, i_8_236_1775_0, i_8_236_1776_0, i_8_236_1777_0,
    i_8_236_1824_0, i_8_236_1854_0, i_8_236_1855_0, i_8_236_1862_0,
    i_8_236_1868_0, i_8_236_1881_0, i_8_236_1984_0, i_8_236_2021_0,
    i_8_236_2034_0, i_8_236_2035_0, i_8_236_2037_0, i_8_236_2039_0,
    i_8_236_2041_0, i_8_236_2092_0, i_8_236_2099_0, i_8_236_2147_0,
    i_8_236_2174_0, i_8_236_2237_0, i_8_236_2268_0,
    o_8_236_0_0  );
  input  i_8_236_36_0, i_8_236_37_0, i_8_236_64_0, i_8_236_112_0,
    i_8_236_166_0, i_8_236_167_0, i_8_236_193_0, i_8_236_194_0,
    i_8_236_221_0, i_8_236_226_0, i_8_236_300_0, i_8_236_362_0,
    i_8_236_373_0, i_8_236_385_0, i_8_236_397_0, i_8_236_420_0,
    i_8_236_421_0, i_8_236_484_0, i_8_236_489_0, i_8_236_493_0,
    i_8_236_522_0, i_8_236_525_0, i_8_236_526_0, i_8_236_529_0,
    i_8_236_606_0, i_8_236_607_0, i_8_236_608_0, i_8_236_613_0,
    i_8_236_662_0, i_8_236_698_0, i_8_236_700_0, i_8_236_701_0,
    i_8_236_707_0, i_8_236_710_0, i_8_236_801_0, i_8_236_802_0,
    i_8_236_803_0, i_8_236_806_0, i_8_236_809_0, i_8_236_843_0,
    i_8_236_844_0, i_8_236_854_0, i_8_236_932_0, i_8_236_935_0,
    i_8_236_972_0, i_8_236_993_0, i_8_236_995_0, i_8_236_1040_0,
    i_8_236_1047_0, i_8_236_1078_0, i_8_236_1113_0, i_8_236_1114_0,
    i_8_236_1115_0, i_8_236_1134_0, i_8_236_1233_0, i_8_236_1234_0,
    i_8_236_1259_0, i_8_236_1269_0, i_8_236_1271_0, i_8_236_1283_0,
    i_8_236_1286_0, i_8_236_1404_0, i_8_236_1489_0, i_8_236_1490_0,
    i_8_236_1507_0, i_8_236_1529_0, i_8_236_1585_0, i_8_236_1621_0,
    i_8_236_1624_0, i_8_236_1634_0, i_8_236_1650_0, i_8_236_1668_0,
    i_8_236_1678_0, i_8_236_1682_0, i_8_236_1710_0, i_8_236_1711_0,
    i_8_236_1748_0, i_8_236_1766_0, i_8_236_1775_0, i_8_236_1776_0,
    i_8_236_1777_0, i_8_236_1824_0, i_8_236_1854_0, i_8_236_1855_0,
    i_8_236_1862_0, i_8_236_1868_0, i_8_236_1881_0, i_8_236_1984_0,
    i_8_236_2021_0, i_8_236_2034_0, i_8_236_2035_0, i_8_236_2037_0,
    i_8_236_2039_0, i_8_236_2041_0, i_8_236_2092_0, i_8_236_2099_0,
    i_8_236_2147_0, i_8_236_2174_0, i_8_236_2237_0, i_8_236_2268_0;
  output o_8_236_0_0;
  assign o_8_236_0_0 = ~((~i_8_236_1233_0 & ((~i_8_236_801_0 & ((~i_8_236_37_0 & ~i_8_236_64_0 & ~i_8_236_698_0 & ~i_8_236_701_0 & ((~i_8_236_489_0 & ~i_8_236_803_0 & ~i_8_236_806_0 & ~i_8_236_809_0 & ~i_8_236_843_0 & ~i_8_236_993_0 & ~i_8_236_1650_0 & ~i_8_236_1777_0 & ~i_8_236_2037_0) | (~i_8_236_385_0 & ~i_8_236_493_0 & ~i_8_236_700_0 & ~i_8_236_802_0 & ~i_8_236_935_0 & ~i_8_236_972_0 & ~i_8_236_1668_0 & ~i_8_236_1776_0 & ~i_8_236_2035_0 & ~i_8_236_2041_0))) | (~i_8_236_935_0 & ((~i_8_236_167_0 & i_8_236_526_0 & ~i_8_236_710_0 & ~i_8_236_806_0 & ~i_8_236_932_0 & ~i_8_236_1078_0 & ~i_8_236_1748_0 & ~i_8_236_1868_0) | (i_8_236_193_0 & ~i_8_236_489_0 & ~i_8_236_809_0 & ~i_8_236_972_0 & ~i_8_236_1624_0 & ~i_8_236_1855_0 & ~i_8_236_2037_0))) | (~i_8_236_36_0 & i_8_236_112_0 & ~i_8_236_700_0 & i_8_236_1047_0 & i_8_236_1678_0) | (~i_8_236_397_0 & ~i_8_236_802_0 & ~i_8_236_803_0 & ~i_8_236_843_0 & ~i_8_236_854_0 & ~i_8_236_1078_0 & ~i_8_236_1259_0 & ~i_8_236_1668_0 & ~i_8_236_1862_0 & i_8_236_1984_0 & ~i_8_236_2021_0 & ~i_8_236_2039_0 & ~i_8_236_2099_0 & ~i_8_236_2237_0))) | (~i_8_236_2041_0 & ((i_8_236_112_0 & i_8_236_484_0 & ~i_8_236_1624_0) | (~i_8_236_37_0 & ~i_8_236_385_0 & i_8_236_993_0 & ~i_8_236_1234_0 & ~i_8_236_1775_0 & ~i_8_236_1854_0 & ~i_8_236_2035_0 & ~i_8_236_2237_0))) | (~i_8_236_806_0 & ~i_8_236_843_0 & ~i_8_236_1283_0 & ~i_8_236_1621_0 & ~i_8_236_1984_0 & i_8_236_2099_0) | (~i_8_236_493_0 & i_8_236_608_0 & ~i_8_236_802_0 & ~i_8_236_932_0 & ~i_8_236_1862_0 & ~i_8_236_1881_0 & ~i_8_236_2021_0 & ~i_8_236_2147_0))) | (~i_8_236_801_0 & ((~i_8_236_112_0 & ~i_8_236_2034_0 & ((~i_8_236_37_0 & ~i_8_236_167_0 & ~i_8_236_843_0 & ~i_8_236_1881_0 & ~i_8_236_2039_0 & ((~i_8_236_166_0 & ~i_8_236_700_0 & ~i_8_236_806_0 & ~i_8_236_935_0 & ~i_8_236_1078_0 & ~i_8_236_1234_0 & ~i_8_236_1259_0 & ~i_8_236_1585_0 & ~i_8_236_1650_0 & ~i_8_236_1984_0 & ~i_8_236_2035_0) | (~i_8_236_64_0 & ~i_8_236_373_0 & ~i_8_236_385_0 & ~i_8_236_484_0 & ~i_8_236_489_0 & ~i_8_236_613_0 & ~i_8_236_662_0 & ~i_8_236_854_0 & ~i_8_236_932_0 & ~i_8_236_1854_0 & ~i_8_236_2099_0 & ~i_8_236_2147_0))) | (~i_8_236_36_0 & ~i_8_236_166_0 & ~i_8_236_385_0 & ~i_8_236_1234_0 & i_8_236_1776_0 & ~i_8_236_2037_0))) | (~i_8_236_385_0 & ((i_8_236_193_0 & ~i_8_236_2037_0 & ~i_8_236_2039_0 & ((~i_8_236_36_0 & ~i_8_236_489_0 & ~i_8_236_972_0 & ~i_8_236_1259_0 & ~i_8_236_1269_0 & ~i_8_236_1711_0) | (~i_8_236_522_0 & ~i_8_236_525_0 & ~i_8_236_606_0 & ~i_8_236_993_0 & ~i_8_236_1114_0 & ~i_8_236_1286_0 & ~i_8_236_1585_0 & ~i_8_236_1621_0 & ~i_8_236_1776_0 & ~i_8_236_2041_0))) | (i_8_236_300_0 & ~i_8_236_373_0 & ~i_8_236_993_0 & ~i_8_236_1286_0 & ~i_8_236_1585_0 & ~i_8_236_1621_0 & ~i_8_236_1650_0 & ~i_8_236_1682_0 & ~i_8_236_1748_0))) | (~i_8_236_36_0 & i_8_236_1678_0 & ((~i_8_236_489_0 & ~i_8_236_493_0 & i_8_236_1777_0 & ~i_8_236_1881_0) | (~i_8_236_37_0 & ~i_8_236_300_0 & i_8_236_489_0 & ~i_8_236_843_0 & ~i_8_236_972_0 & ~i_8_236_1585_0 & ~i_8_236_1824_0 & ~i_8_236_2021_0 & ~i_8_236_2041_0))))) | (~i_8_236_36_0 & ((~i_8_236_37_0 & ~i_8_236_809_0 & ((~i_8_236_167_0 & ~i_8_236_385_0 & i_8_236_698_0 & i_8_236_707_0 & ~i_8_236_802_0 & ~i_8_236_803_0 & ~i_8_236_932_0 & ~i_8_236_1078_0 & ~i_8_236_1711_0 & ~i_8_236_1854_0) | (~i_8_236_64_0 & ~i_8_236_362_0 & ~i_8_236_484_0 & ~i_8_236_489_0 & ~i_8_236_662_0 & ~i_8_236_843_0 & ~i_8_236_1047_0 & ~i_8_236_1259_0 & ~i_8_236_1269_0 & ~i_8_236_1271_0 & ~i_8_236_1775_0 & ~i_8_236_1868_0 & ~i_8_236_1984_0 & ~i_8_236_2034_0 & ~i_8_236_2037_0 & ~i_8_236_2041_0))) | (~i_8_236_844_0 & ((~i_8_236_803_0 & ~i_8_236_1269_0 & ~i_8_236_1283_0 & i_8_236_1404_0 & ~i_8_236_2035_0 & ~i_8_236_2041_0 & i_8_236_2092_0) | (i_8_236_529_0 & ~i_8_236_701_0 & ~i_8_236_1621_0 & ~i_8_236_2099_0))) | (~i_8_236_1078_0 & ~i_8_236_1234_0 & ~i_8_236_1259_0 & ~i_8_236_1271_0 & i_8_236_1748_0 & ~i_8_236_1854_0 & ~i_8_236_1855_0 & ~i_8_236_2035_0) | (~i_8_236_385_0 & i_8_236_526_0 & ~i_8_236_802_0 & i_8_236_1824_0 & ~i_8_236_1868_0) | (~i_8_236_972_0 & i_8_236_1134_0 & i_8_236_1776_0 & ~i_8_236_1824_0 & ~i_8_236_2037_0 & i_8_236_2268_0))) | (~i_8_236_300_0 & ~i_8_236_1078_0 & ((~i_8_236_64_0 & ~i_8_236_698_0 & ~i_8_236_700_0 & ~i_8_236_843_0 & ~i_8_236_993_0 & ~i_8_236_1234_0 & ~i_8_236_1259_0 & ~i_8_236_1269_0 & ~i_8_236_1283_0 & ~i_8_236_1650_0 & ~i_8_236_1776_0 & ~i_8_236_1824_0 & ~i_8_236_1881_0 & ~i_8_236_2035_0 & ~i_8_236_2037_0) | (~i_8_236_613_0 & i_8_236_698_0 & ~i_8_236_803_0 & ~i_8_236_809_0 & i_8_236_1682_0 & ~i_8_236_1855_0 & i_8_236_2147_0))) | (i_8_236_525_0 & ((~i_8_236_489_0 & ~i_8_236_606_0 & i_8_236_1489_0) | (i_8_236_493_0 & i_8_236_844_0 & ~i_8_236_1047_0 & ~i_8_236_1259_0 & ~i_8_236_1777_0 & ~i_8_236_1984_0 & ~i_8_236_2268_0))) | (~i_8_236_803_0 & ((~i_8_236_397_0 & ((i_8_236_221_0 & ~i_8_236_698_0 & ~i_8_236_802_0 & ~i_8_236_806_0 & ~i_8_236_935_0 & ~i_8_236_2034_0 & ~i_8_236_2035_0) | (~i_8_236_1047_0 & i_8_236_1490_0 & ~i_8_236_1855_0 & i_8_236_2092_0))) | (~i_8_236_1404_0 & ((~i_8_236_489_0 & ((~i_8_236_1134_0 & i_8_236_1634_0 & ~i_8_236_1650_0 & ~i_8_236_1855_0 & ~i_8_236_2021_0) | (i_8_236_300_0 & ~i_8_236_809_0 & ~i_8_236_935_0 & ~i_8_236_972_0 & ~i_8_236_1507_0 & ~i_8_236_1624_0 & ~i_8_236_1634_0 & ~i_8_236_2034_0 & ~i_8_236_2037_0))) | (~i_8_236_193_0 & ~i_8_236_522_0 & ~i_8_236_710_0 & ~i_8_236_806_0 & ~i_8_236_993_0 & ~i_8_236_1269_0 & ~i_8_236_1624_0 & ~i_8_236_1682_0 & i_8_236_1775_0 & ~i_8_236_1854_0 & ~i_8_236_2268_0))) | (~i_8_236_64_0 & ~i_8_236_194_0 & ~i_8_236_608_0 & ~i_8_236_806_0 & ~i_8_236_844_0 & ~i_8_236_932_0 & ~i_8_236_1259_0 & ~i_8_236_1777_0 & ~i_8_236_1881_0 & i_8_236_2099_0))) | (~i_8_236_64_0 & ((~i_8_236_221_0 & i_8_236_526_0 & ~i_8_236_843_0 & ~i_8_236_844_0 & ~i_8_236_1668_0 & ~i_8_236_1766_0 & i_8_236_1881_0) | (i_8_236_606_0 & ~i_8_236_700_0 & ~i_8_236_972_0 & ~i_8_236_1624_0 & i_8_236_1776_0 & i_8_236_1777_0 & ~i_8_236_2035_0))) | (~i_8_236_1984_0 & ((~i_8_236_613_0 & ((i_8_236_844_0 & ~i_8_236_1234_0 & ~i_8_236_1621_0 & ~i_8_236_1678_0 & ~i_8_236_1776_0 & i_8_236_1777_0 & ~i_8_236_2092_0 & ~i_8_236_2147_0) | (~i_8_236_806_0 & ~i_8_236_843_0 & ~i_8_236_993_0 & i_8_236_1114_0 & ~i_8_236_1259_0 & ~i_8_236_1269_0 & ~i_8_236_1766_0 & ~i_8_236_1868_0 & ~i_8_236_2037_0 & ~i_8_236_2268_0))) | (~i_8_236_1269_0 & i_8_236_1777_0 & ~i_8_236_1824_0 & i_8_236_2037_0 & ~i_8_236_2268_0))) | (~i_8_236_1271_0 & ((~i_8_236_1040_0 & ~i_8_236_2041_0 & ((i_8_236_362_0 & ~i_8_236_932_0 & ~i_8_236_1114_0 & ~i_8_236_2034_0 & ~i_8_236_2035_0 & ~i_8_236_1710_0 & i_8_236_1775_0) | (i_8_236_373_0 & ~i_8_236_397_0 & ~i_8_236_698_0 & ~i_8_236_701_0 & ~i_8_236_993_0 & ~i_8_236_1621_0 & ~i_8_236_2037_0 & ~i_8_236_2237_0))) | (i_8_236_608_0 & i_8_236_1490_0))) | (~i_8_236_1234_0 & ((~i_8_236_972_0 & i_8_236_1113_0 & ~i_8_236_1766_0 & i_8_236_1776_0 & ~i_8_236_2034_0) | (~i_8_236_167_0 & ~i_8_236_662_0 & i_8_236_701_0 & ~i_8_236_854_0 & ~i_8_236_935_0 & ~i_8_236_1259_0 & ~i_8_236_1404_0 & ~i_8_236_1678_0 & ~i_8_236_2147_0))) | (i_8_236_193_0 & i_8_236_484_0 & i_8_236_1824_0 & ~i_8_236_1862_0) | (~i_8_236_806_0 & ~i_8_236_1286_0 & ~i_8_236_1855_0 & ~i_8_236_1881_0 & i_8_236_2174_0));
endmodule



// Benchmark "kernel_8_237" written by ABC on Sun Jul 19 10:07:12 2020

module kernel_8_237 ( 
    i_8_237_23_0, i_8_237_31_0, i_8_237_136_0, i_8_237_189_0,
    i_8_237_262_0, i_8_237_265_0, i_8_237_266_0, i_8_237_340_0,
    i_8_237_373_0, i_8_237_381_0, i_8_237_394_0, i_8_237_421_0,
    i_8_237_426_0, i_8_237_430_0, i_8_237_453_0, i_8_237_454_0,
    i_8_237_455_0, i_8_237_492_0, i_8_237_528_0, i_8_237_547_0,
    i_8_237_554_0, i_8_237_604_0, i_8_237_616_0, i_8_237_633_0,
    i_8_237_634_0, i_8_237_654_0, i_8_237_658_0, i_8_237_660_0,
    i_8_237_661_0, i_8_237_663_0, i_8_237_706_0, i_8_237_717_0,
    i_8_237_719_0, i_8_237_778_0, i_8_237_840_0, i_8_237_841_0,
    i_8_237_880_0, i_8_237_881_0, i_8_237_903_0, i_8_237_967_0,
    i_8_237_970_0, i_8_237_994_0, i_8_237_1024_0, i_8_237_1074_0,
    i_8_237_1081_0, i_8_237_1111_0, i_8_237_1121_0, i_8_237_1122_0,
    i_8_237_1129_0, i_8_237_1131_0, i_8_237_1198_0, i_8_237_1237_0,
    i_8_237_1249_0, i_8_237_1289_0, i_8_237_1292_0, i_8_237_1294_0,
    i_8_237_1321_0, i_8_237_1326_0, i_8_237_1357_0, i_8_237_1431_0,
    i_8_237_1434_0, i_8_237_1450_0, i_8_237_1471_0, i_8_237_1484_0,
    i_8_237_1489_0, i_8_237_1504_0, i_8_237_1519_0, i_8_237_1538_0,
    i_8_237_1542_0, i_8_237_1605_0, i_8_237_1625_0, i_8_237_1630_0,
    i_8_237_1632_0, i_8_237_1705_0, i_8_237_1743_0, i_8_237_1745_0,
    i_8_237_1749_0, i_8_237_1752_0, i_8_237_1753_0, i_8_237_1790_0,
    i_8_237_1804_0, i_8_237_1805_0, i_8_237_1813_0, i_8_237_1822_0,
    i_8_237_1823_0, i_8_237_1843_0, i_8_237_1849_0, i_8_237_1894_0,
    i_8_237_1922_0, i_8_237_1927_0, i_8_237_1947_0, i_8_237_1965_0,
    i_8_237_1992_0, i_8_237_2044_0, i_8_237_2093_0, i_8_237_2101_0,
    i_8_237_2146_0, i_8_237_2271_0, i_8_237_2289_0, i_8_237_2302_0,
    o_8_237_0_0  );
  input  i_8_237_23_0, i_8_237_31_0, i_8_237_136_0, i_8_237_189_0,
    i_8_237_262_0, i_8_237_265_0, i_8_237_266_0, i_8_237_340_0,
    i_8_237_373_0, i_8_237_381_0, i_8_237_394_0, i_8_237_421_0,
    i_8_237_426_0, i_8_237_430_0, i_8_237_453_0, i_8_237_454_0,
    i_8_237_455_0, i_8_237_492_0, i_8_237_528_0, i_8_237_547_0,
    i_8_237_554_0, i_8_237_604_0, i_8_237_616_0, i_8_237_633_0,
    i_8_237_634_0, i_8_237_654_0, i_8_237_658_0, i_8_237_660_0,
    i_8_237_661_0, i_8_237_663_0, i_8_237_706_0, i_8_237_717_0,
    i_8_237_719_0, i_8_237_778_0, i_8_237_840_0, i_8_237_841_0,
    i_8_237_880_0, i_8_237_881_0, i_8_237_903_0, i_8_237_967_0,
    i_8_237_970_0, i_8_237_994_0, i_8_237_1024_0, i_8_237_1074_0,
    i_8_237_1081_0, i_8_237_1111_0, i_8_237_1121_0, i_8_237_1122_0,
    i_8_237_1129_0, i_8_237_1131_0, i_8_237_1198_0, i_8_237_1237_0,
    i_8_237_1249_0, i_8_237_1289_0, i_8_237_1292_0, i_8_237_1294_0,
    i_8_237_1321_0, i_8_237_1326_0, i_8_237_1357_0, i_8_237_1431_0,
    i_8_237_1434_0, i_8_237_1450_0, i_8_237_1471_0, i_8_237_1484_0,
    i_8_237_1489_0, i_8_237_1504_0, i_8_237_1519_0, i_8_237_1538_0,
    i_8_237_1542_0, i_8_237_1605_0, i_8_237_1625_0, i_8_237_1630_0,
    i_8_237_1632_0, i_8_237_1705_0, i_8_237_1743_0, i_8_237_1745_0,
    i_8_237_1749_0, i_8_237_1752_0, i_8_237_1753_0, i_8_237_1790_0,
    i_8_237_1804_0, i_8_237_1805_0, i_8_237_1813_0, i_8_237_1822_0,
    i_8_237_1823_0, i_8_237_1843_0, i_8_237_1849_0, i_8_237_1894_0,
    i_8_237_1922_0, i_8_237_1927_0, i_8_237_1947_0, i_8_237_1965_0,
    i_8_237_1992_0, i_8_237_2044_0, i_8_237_2093_0, i_8_237_2101_0,
    i_8_237_2146_0, i_8_237_2271_0, i_8_237_2289_0, i_8_237_2302_0;
  output o_8_237_0_0;
  assign o_8_237_0_0 = 0;
endmodule



// Benchmark "kernel_8_238" written by ABC on Sun Jul 19 10:07:12 2020

module kernel_8_238 ( 
    i_8_238_111_0, i_8_238_117_0, i_8_238_120_0, i_8_238_165_0,
    i_8_238_166_0, i_8_238_169_0, i_8_238_187_0, i_8_238_265_0,
    i_8_238_283_0, i_8_238_289_0, i_8_238_290_0, i_8_238_291_0,
    i_8_238_297_0, i_8_238_319_0, i_8_238_321_0, i_8_238_366_0,
    i_8_238_367_0, i_8_238_368_0, i_8_238_433_0, i_8_238_436_0,
    i_8_238_499_0, i_8_238_546_0, i_8_238_555_0, i_8_238_588_0,
    i_8_238_606_0, i_8_238_635_0, i_8_238_642_0, i_8_238_672_0,
    i_8_238_673_0, i_8_238_674_0, i_8_238_678_0, i_8_238_695_0,
    i_8_238_708_0, i_8_238_724_0, i_8_238_726_0, i_8_238_727_0,
    i_8_238_781_0, i_8_238_783_0, i_8_238_804_0, i_8_238_805_0,
    i_8_238_810_0, i_8_238_811_0, i_8_238_813_0, i_8_238_814_0,
    i_8_238_829_0, i_8_238_849_0, i_8_238_877_0, i_8_238_964_0,
    i_8_238_967_0, i_8_238_973_0, i_8_238_1011_0, i_8_238_1029_0,
    i_8_238_1030_0, i_8_238_1032_0, i_8_238_1119_0, i_8_238_1200_0,
    i_8_238_1239_0, i_8_238_1264_0, i_8_238_1299_0, i_8_238_1324_0,
    i_8_238_1345_0, i_8_238_1351_0, i_8_238_1441_0, i_8_238_1452_0,
    i_8_238_1491_0, i_8_238_1507_0, i_8_238_1533_0, i_8_238_1542_0,
    i_8_238_1546_0, i_8_238_1578_0, i_8_238_1587_0, i_8_238_1588_0,
    i_8_238_1623_0, i_8_238_1731_0, i_8_238_1749_0, i_8_238_1767_0,
    i_8_238_1770_0, i_8_238_1779_0, i_8_238_1782_0, i_8_238_1821_0,
    i_8_238_1824_0, i_8_238_1825_0, i_8_238_1846_0, i_8_238_1848_0,
    i_8_238_1851_0, i_8_238_1876_0, i_8_238_1903_0, i_8_238_1938_0,
    i_8_238_1993_0, i_8_238_1996_0, i_8_238_2029_0, i_8_238_2031_0,
    i_8_238_2037_0, i_8_238_2038_0, i_8_238_2074_0, i_8_238_2116_0,
    i_8_238_2128_0, i_8_238_2150_0, i_8_238_2190_0, i_8_238_2272_0,
    o_8_238_0_0  );
  input  i_8_238_111_0, i_8_238_117_0, i_8_238_120_0, i_8_238_165_0,
    i_8_238_166_0, i_8_238_169_0, i_8_238_187_0, i_8_238_265_0,
    i_8_238_283_0, i_8_238_289_0, i_8_238_290_0, i_8_238_291_0,
    i_8_238_297_0, i_8_238_319_0, i_8_238_321_0, i_8_238_366_0,
    i_8_238_367_0, i_8_238_368_0, i_8_238_433_0, i_8_238_436_0,
    i_8_238_499_0, i_8_238_546_0, i_8_238_555_0, i_8_238_588_0,
    i_8_238_606_0, i_8_238_635_0, i_8_238_642_0, i_8_238_672_0,
    i_8_238_673_0, i_8_238_674_0, i_8_238_678_0, i_8_238_695_0,
    i_8_238_708_0, i_8_238_724_0, i_8_238_726_0, i_8_238_727_0,
    i_8_238_781_0, i_8_238_783_0, i_8_238_804_0, i_8_238_805_0,
    i_8_238_810_0, i_8_238_811_0, i_8_238_813_0, i_8_238_814_0,
    i_8_238_829_0, i_8_238_849_0, i_8_238_877_0, i_8_238_964_0,
    i_8_238_967_0, i_8_238_973_0, i_8_238_1011_0, i_8_238_1029_0,
    i_8_238_1030_0, i_8_238_1032_0, i_8_238_1119_0, i_8_238_1200_0,
    i_8_238_1239_0, i_8_238_1264_0, i_8_238_1299_0, i_8_238_1324_0,
    i_8_238_1345_0, i_8_238_1351_0, i_8_238_1441_0, i_8_238_1452_0,
    i_8_238_1491_0, i_8_238_1507_0, i_8_238_1533_0, i_8_238_1542_0,
    i_8_238_1546_0, i_8_238_1578_0, i_8_238_1587_0, i_8_238_1588_0,
    i_8_238_1623_0, i_8_238_1731_0, i_8_238_1749_0, i_8_238_1767_0,
    i_8_238_1770_0, i_8_238_1779_0, i_8_238_1782_0, i_8_238_1821_0,
    i_8_238_1824_0, i_8_238_1825_0, i_8_238_1846_0, i_8_238_1848_0,
    i_8_238_1851_0, i_8_238_1876_0, i_8_238_1903_0, i_8_238_1938_0,
    i_8_238_1993_0, i_8_238_1996_0, i_8_238_2029_0, i_8_238_2031_0,
    i_8_238_2037_0, i_8_238_2038_0, i_8_238_2074_0, i_8_238_2116_0,
    i_8_238_2128_0, i_8_238_2150_0, i_8_238_2190_0, i_8_238_2272_0;
  output o_8_238_0_0;
  assign o_8_238_0_0 = 0;
endmodule



// Benchmark "kernel_8_239" written by ABC on Sun Jul 19 10:07:13 2020

module kernel_8_239 ( 
    i_8_239_23_0, i_8_239_31_0, i_8_239_32_0, i_8_239_34_0, i_8_239_165_0,
    i_8_239_201_0, i_8_239_225_0, i_8_239_263_0, i_8_239_265_0,
    i_8_239_279_0, i_8_239_318_0, i_8_239_335_0, i_8_239_365_0,
    i_8_239_368_0, i_8_239_417_0, i_8_239_443_0, i_8_239_447_0,
    i_8_239_451_0, i_8_239_452_0, i_8_239_483_0, i_8_239_525_0,
    i_8_239_530_0, i_8_239_533_0, i_8_239_615_0, i_8_239_616_0,
    i_8_239_631_0, i_8_239_688_0, i_8_239_689_0, i_8_239_704_0,
    i_8_239_717_0, i_8_239_772_0, i_8_239_831_0, i_8_239_842_0,
    i_8_239_874_0, i_8_239_875_0, i_8_239_938_0, i_8_239_970_0,
    i_8_239_1054_0, i_8_239_1057_0, i_8_239_1075_0, i_8_239_1077_0,
    i_8_239_1078_0, i_8_239_1099_0, i_8_239_1225_0, i_8_239_1228_0,
    i_8_239_1246_0, i_8_239_1247_0, i_8_239_1261_0, i_8_239_1282_0,
    i_8_239_1305_0, i_8_239_1309_0, i_8_239_1385_0, i_8_239_1407_0,
    i_8_239_1410_0, i_8_239_1423_0, i_8_239_1435_0, i_8_239_1436_0,
    i_8_239_1437_0, i_8_239_1469_0, i_8_239_1472_0, i_8_239_1536_0,
    i_8_239_1562_0, i_8_239_1567_0, i_8_239_1591_0, i_8_239_1598_0,
    i_8_239_1607_0, i_8_239_1622_0, i_8_239_1626_0, i_8_239_1654_0,
    i_8_239_1675_0, i_8_239_1684_0, i_8_239_1702_0, i_8_239_1722_0,
    i_8_239_1723_0, i_8_239_1752_0, i_8_239_1810_0, i_8_239_1825_0,
    i_8_239_1837_0, i_8_239_1838_0, i_8_239_1841_0, i_8_239_1868_0,
    i_8_239_1870_0, i_8_239_1901_0, i_8_239_1930_0, i_8_239_1967_0,
    i_8_239_2045_0, i_8_239_2117_0, i_8_239_2126_0, i_8_239_2129_0,
    i_8_239_2143_0, i_8_239_2144_0, i_8_239_2209_0, i_8_239_2212_0,
    i_8_239_2214_0, i_8_239_2242_0, i_8_239_2246_0, i_8_239_2257_0,
    i_8_239_2264_0, i_8_239_2292_0, i_8_239_2303_0,
    o_8_239_0_0  );
  input  i_8_239_23_0, i_8_239_31_0, i_8_239_32_0, i_8_239_34_0,
    i_8_239_165_0, i_8_239_201_0, i_8_239_225_0, i_8_239_263_0,
    i_8_239_265_0, i_8_239_279_0, i_8_239_318_0, i_8_239_335_0,
    i_8_239_365_0, i_8_239_368_0, i_8_239_417_0, i_8_239_443_0,
    i_8_239_447_0, i_8_239_451_0, i_8_239_452_0, i_8_239_483_0,
    i_8_239_525_0, i_8_239_530_0, i_8_239_533_0, i_8_239_615_0,
    i_8_239_616_0, i_8_239_631_0, i_8_239_688_0, i_8_239_689_0,
    i_8_239_704_0, i_8_239_717_0, i_8_239_772_0, i_8_239_831_0,
    i_8_239_842_0, i_8_239_874_0, i_8_239_875_0, i_8_239_938_0,
    i_8_239_970_0, i_8_239_1054_0, i_8_239_1057_0, i_8_239_1075_0,
    i_8_239_1077_0, i_8_239_1078_0, i_8_239_1099_0, i_8_239_1225_0,
    i_8_239_1228_0, i_8_239_1246_0, i_8_239_1247_0, i_8_239_1261_0,
    i_8_239_1282_0, i_8_239_1305_0, i_8_239_1309_0, i_8_239_1385_0,
    i_8_239_1407_0, i_8_239_1410_0, i_8_239_1423_0, i_8_239_1435_0,
    i_8_239_1436_0, i_8_239_1437_0, i_8_239_1469_0, i_8_239_1472_0,
    i_8_239_1536_0, i_8_239_1562_0, i_8_239_1567_0, i_8_239_1591_0,
    i_8_239_1598_0, i_8_239_1607_0, i_8_239_1622_0, i_8_239_1626_0,
    i_8_239_1654_0, i_8_239_1675_0, i_8_239_1684_0, i_8_239_1702_0,
    i_8_239_1722_0, i_8_239_1723_0, i_8_239_1752_0, i_8_239_1810_0,
    i_8_239_1825_0, i_8_239_1837_0, i_8_239_1838_0, i_8_239_1841_0,
    i_8_239_1868_0, i_8_239_1870_0, i_8_239_1901_0, i_8_239_1930_0,
    i_8_239_1967_0, i_8_239_2045_0, i_8_239_2117_0, i_8_239_2126_0,
    i_8_239_2129_0, i_8_239_2143_0, i_8_239_2144_0, i_8_239_2209_0,
    i_8_239_2212_0, i_8_239_2214_0, i_8_239_2242_0, i_8_239_2246_0,
    i_8_239_2257_0, i_8_239_2264_0, i_8_239_2292_0, i_8_239_2303_0;
  output o_8_239_0_0;
  assign o_8_239_0_0 = 0;
endmodule



// Benchmark "kernel_8_240" written by ABC on Sun Jul 19 10:07:14 2020

module kernel_8_240 ( 
    i_8_240_11_0, i_8_240_84_0, i_8_240_87_0, i_8_240_96_0, i_8_240_97_0,
    i_8_240_102_0, i_8_240_107_0, i_8_240_222_0, i_8_240_223_0,
    i_8_240_240_0, i_8_240_255_0, i_8_240_282_0, i_8_240_300_0,
    i_8_240_301_0, i_8_240_375_0, i_8_240_444_0, i_8_240_453_0,
    i_8_240_454_0, i_8_240_475_0, i_8_240_483_0, i_8_240_485_0,
    i_8_240_555_0, i_8_240_588_0, i_8_240_596_0, i_8_240_601_0,
    i_8_240_613_0, i_8_240_621_0, i_8_240_714_0, i_8_240_717_0,
    i_8_240_720_0, i_8_240_759_0, i_8_240_771_0, i_8_240_780_0,
    i_8_240_795_0, i_8_240_811_0, i_8_240_813_0, i_8_240_825_0,
    i_8_240_840_0, i_8_240_889_0, i_8_240_972_0, i_8_240_1014_0,
    i_8_240_1026_0, i_8_240_1029_0, i_8_240_1049_0, i_8_240_1111_0,
    i_8_240_1113_0, i_8_240_1135_0, i_8_240_1137_0, i_8_240_1233_0,
    i_8_240_1255_0, i_8_240_1257_0, i_8_240_1281_0, i_8_240_1313_0,
    i_8_240_1438_0, i_8_240_1443_0, i_8_240_1482_0, i_8_240_1533_0,
    i_8_240_1534_0, i_8_240_1541_0, i_8_240_1542_0, i_8_240_1548_0,
    i_8_240_1555_0, i_8_240_1587_0, i_8_240_1588_0, i_8_240_1590_0,
    i_8_240_1668_0, i_8_240_1677_0, i_8_240_1725_0, i_8_240_1753_0,
    i_8_240_1761_0, i_8_240_1762_0, i_8_240_1780_0, i_8_240_1785_0,
    i_8_240_1788_0, i_8_240_1812_0, i_8_240_1813_0, i_8_240_1840_0,
    i_8_240_1867_0, i_8_240_1893_0, i_8_240_1914_0, i_8_240_1918_0,
    i_8_240_1923_0, i_8_240_1968_0, i_8_240_1969_0, i_8_240_1974_0,
    i_8_240_1995_0, i_8_240_2001_0, i_8_240_2031_0, i_8_240_2046_0,
    i_8_240_2050_0, i_8_240_2054_0, i_8_240_2130_0, i_8_240_2136_0,
    i_8_240_2181_0, i_8_240_2214_0, i_8_240_2215_0, i_8_240_2263_0,
    i_8_240_2271_0, i_8_240_2272_0, i_8_240_2284_0,
    o_8_240_0_0  );
  input  i_8_240_11_0, i_8_240_84_0, i_8_240_87_0, i_8_240_96_0,
    i_8_240_97_0, i_8_240_102_0, i_8_240_107_0, i_8_240_222_0,
    i_8_240_223_0, i_8_240_240_0, i_8_240_255_0, i_8_240_282_0,
    i_8_240_300_0, i_8_240_301_0, i_8_240_375_0, i_8_240_444_0,
    i_8_240_453_0, i_8_240_454_0, i_8_240_475_0, i_8_240_483_0,
    i_8_240_485_0, i_8_240_555_0, i_8_240_588_0, i_8_240_596_0,
    i_8_240_601_0, i_8_240_613_0, i_8_240_621_0, i_8_240_714_0,
    i_8_240_717_0, i_8_240_720_0, i_8_240_759_0, i_8_240_771_0,
    i_8_240_780_0, i_8_240_795_0, i_8_240_811_0, i_8_240_813_0,
    i_8_240_825_0, i_8_240_840_0, i_8_240_889_0, i_8_240_972_0,
    i_8_240_1014_0, i_8_240_1026_0, i_8_240_1029_0, i_8_240_1049_0,
    i_8_240_1111_0, i_8_240_1113_0, i_8_240_1135_0, i_8_240_1137_0,
    i_8_240_1233_0, i_8_240_1255_0, i_8_240_1257_0, i_8_240_1281_0,
    i_8_240_1313_0, i_8_240_1438_0, i_8_240_1443_0, i_8_240_1482_0,
    i_8_240_1533_0, i_8_240_1534_0, i_8_240_1541_0, i_8_240_1542_0,
    i_8_240_1548_0, i_8_240_1555_0, i_8_240_1587_0, i_8_240_1588_0,
    i_8_240_1590_0, i_8_240_1668_0, i_8_240_1677_0, i_8_240_1725_0,
    i_8_240_1753_0, i_8_240_1761_0, i_8_240_1762_0, i_8_240_1780_0,
    i_8_240_1785_0, i_8_240_1788_0, i_8_240_1812_0, i_8_240_1813_0,
    i_8_240_1840_0, i_8_240_1867_0, i_8_240_1893_0, i_8_240_1914_0,
    i_8_240_1918_0, i_8_240_1923_0, i_8_240_1968_0, i_8_240_1969_0,
    i_8_240_1974_0, i_8_240_1995_0, i_8_240_2001_0, i_8_240_2031_0,
    i_8_240_2046_0, i_8_240_2050_0, i_8_240_2054_0, i_8_240_2130_0,
    i_8_240_2136_0, i_8_240_2181_0, i_8_240_2214_0, i_8_240_2215_0,
    i_8_240_2263_0, i_8_240_2271_0, i_8_240_2272_0, i_8_240_2284_0;
  output o_8_240_0_0;
  assign o_8_240_0_0 = 0;
endmodule



// Benchmark "kernel_8_241" written by ABC on Sun Jul 19 10:07:16 2020

module kernel_8_241 ( 
    i_8_241_36_0, i_8_241_63_0, i_8_241_189_0, i_8_241_190_0,
    i_8_241_191_0, i_8_241_192_0, i_8_241_193_0, i_8_241_194_0,
    i_8_241_223_0, i_8_241_237_0, i_8_241_238_0, i_8_241_258_0,
    i_8_241_300_0, i_8_241_325_0, i_8_241_327_0, i_8_241_328_0,
    i_8_241_360_0, i_8_241_393_0, i_8_241_529_0, i_8_241_615_0,
    i_8_241_618_0, i_8_241_624_0, i_8_241_628_0, i_8_241_665_0,
    i_8_241_689_0, i_8_241_696_0, i_8_241_716_0, i_8_241_781_0,
    i_8_241_837_0, i_8_241_842_0, i_8_241_844_0, i_8_241_849_0,
    i_8_241_853_0, i_8_241_861_0, i_8_241_862_0, i_8_241_874_0,
    i_8_241_875_0, i_8_241_877_0, i_8_241_878_0, i_8_241_937_0,
    i_8_241_939_0, i_8_241_970_0, i_8_241_996_0, i_8_241_1014_0,
    i_8_241_1015_0, i_8_241_1029_0, i_8_241_1030_0, i_8_241_1038_0,
    i_8_241_1050_0, i_8_241_1158_0, i_8_241_1231_0, i_8_241_1240_0,
    i_8_241_1263_0, i_8_241_1267_0, i_8_241_1269_0, i_8_241_1284_0,
    i_8_241_1285_0, i_8_241_1290_0, i_8_241_1291_0, i_8_241_1294_0,
    i_8_241_1315_0, i_8_241_1407_0, i_8_241_1408_0, i_8_241_1437_0,
    i_8_241_1444_0, i_8_241_1473_0, i_8_241_1492_0, i_8_241_1510_0,
    i_8_241_1530_0, i_8_241_1545_0, i_8_241_1546_0, i_8_241_1638_0,
    i_8_241_1647_0, i_8_241_1648_0, i_8_241_1651_0, i_8_241_1680_0,
    i_8_241_1700_0, i_8_241_1750_0, i_8_241_1768_0, i_8_241_1769_0,
    i_8_241_1779_0, i_8_241_1815_0, i_8_241_1822_0, i_8_241_1827_0,
    i_8_241_1830_0, i_8_241_1844_0, i_8_241_1881_0, i_8_241_1883_0,
    i_8_241_2037_0, i_8_241_2040_0, i_8_241_2070_0, i_8_241_2091_0,
    i_8_241_2156_0, i_8_241_2157_0, i_8_241_2158_0, i_8_241_2173_0,
    i_8_241_2218_0, i_8_241_2238_0, i_8_241_2239_0, i_8_241_2262_0,
    o_8_241_0_0  );
  input  i_8_241_36_0, i_8_241_63_0, i_8_241_189_0, i_8_241_190_0,
    i_8_241_191_0, i_8_241_192_0, i_8_241_193_0, i_8_241_194_0,
    i_8_241_223_0, i_8_241_237_0, i_8_241_238_0, i_8_241_258_0,
    i_8_241_300_0, i_8_241_325_0, i_8_241_327_0, i_8_241_328_0,
    i_8_241_360_0, i_8_241_393_0, i_8_241_529_0, i_8_241_615_0,
    i_8_241_618_0, i_8_241_624_0, i_8_241_628_0, i_8_241_665_0,
    i_8_241_689_0, i_8_241_696_0, i_8_241_716_0, i_8_241_781_0,
    i_8_241_837_0, i_8_241_842_0, i_8_241_844_0, i_8_241_849_0,
    i_8_241_853_0, i_8_241_861_0, i_8_241_862_0, i_8_241_874_0,
    i_8_241_875_0, i_8_241_877_0, i_8_241_878_0, i_8_241_937_0,
    i_8_241_939_0, i_8_241_970_0, i_8_241_996_0, i_8_241_1014_0,
    i_8_241_1015_0, i_8_241_1029_0, i_8_241_1030_0, i_8_241_1038_0,
    i_8_241_1050_0, i_8_241_1158_0, i_8_241_1231_0, i_8_241_1240_0,
    i_8_241_1263_0, i_8_241_1267_0, i_8_241_1269_0, i_8_241_1284_0,
    i_8_241_1285_0, i_8_241_1290_0, i_8_241_1291_0, i_8_241_1294_0,
    i_8_241_1315_0, i_8_241_1407_0, i_8_241_1408_0, i_8_241_1437_0,
    i_8_241_1444_0, i_8_241_1473_0, i_8_241_1492_0, i_8_241_1510_0,
    i_8_241_1530_0, i_8_241_1545_0, i_8_241_1546_0, i_8_241_1638_0,
    i_8_241_1647_0, i_8_241_1648_0, i_8_241_1651_0, i_8_241_1680_0,
    i_8_241_1700_0, i_8_241_1750_0, i_8_241_1768_0, i_8_241_1769_0,
    i_8_241_1779_0, i_8_241_1815_0, i_8_241_1822_0, i_8_241_1827_0,
    i_8_241_1830_0, i_8_241_1844_0, i_8_241_1881_0, i_8_241_1883_0,
    i_8_241_2037_0, i_8_241_2040_0, i_8_241_2070_0, i_8_241_2091_0,
    i_8_241_2156_0, i_8_241_2157_0, i_8_241_2158_0, i_8_241_2173_0,
    i_8_241_2218_0, i_8_241_2238_0, i_8_241_2239_0, i_8_241_2262_0;
  output o_8_241_0_0;
  assign o_8_241_0_0 = ~((~i_8_241_689_0 & ((~i_8_241_1648_0 & ((~i_8_241_36_0 & i_8_241_325_0 & ((~i_8_241_189_0 & ~i_8_241_191_0 & ~i_8_241_1473_0 & ~i_8_241_1647_0 & ~i_8_241_1750_0 & ~i_8_241_1815_0 & ~i_8_241_1883_0) | (~i_8_241_849_0 & ~i_8_241_937_0 & ~i_8_241_1231_0 & ~i_8_241_1881_0 & ~i_8_241_2040_0 & ~i_8_241_2070_0 & ~i_8_241_2158_0 & ~i_8_241_2173_0))) | (~i_8_241_615_0 & ((~i_8_241_190_0 & ~i_8_241_191_0 & ~i_8_241_258_0 & ~i_8_241_328_0 & i_8_241_970_0 & ~i_8_241_1240_0 & ~i_8_241_1267_0 & ~i_8_241_1285_0 & ~i_8_241_1680_0 & ~i_8_241_1750_0 & ~i_8_241_1815_0 & ~i_8_241_2156_0 & ~i_8_241_2157_0) | (~i_8_241_63_0 & ~i_8_241_842_0 & ~i_8_241_844_0 & i_8_241_874_0 & ~i_8_241_1269_0 & ~i_8_241_1822_0 & ~i_8_241_2070_0 & ~i_8_241_2158_0 & ~i_8_241_2218_0))) | (i_8_241_877_0 & ((~i_8_241_696_0 & i_8_241_875_0 & ~i_8_241_2157_0) | (~i_8_241_189_0 & ~i_8_241_192_0 & ~i_8_241_842_0 & ~i_8_241_1050_0 & ~i_8_241_1231_0 & ~i_8_241_1315_0 & ~i_8_241_1407_0 & ~i_8_241_1638_0 & ~i_8_241_1647_0 & ~i_8_241_1815_0 & ~i_8_241_2070_0 & ~i_8_241_2156_0 & ~i_8_241_2218_0 & ~i_8_241_2262_0))) | (~i_8_241_861_0 & i_8_241_1492_0 & i_8_241_1769_0 & ~i_8_241_2040_0))) | (~i_8_241_191_0 & ((~i_8_241_63_0 & ((~i_8_241_190_0 & ~i_8_241_237_0 & ~i_8_241_853_0 & ~i_8_241_1290_0 & ~i_8_241_1530_0 & ~i_8_241_1638_0 & i_8_241_1750_0 & ~i_8_241_1815_0 & i_8_241_1822_0 & ~i_8_241_2037_0) | (~i_8_241_696_0 & ~i_8_241_716_0 & ~i_8_241_861_0 & ~i_8_241_878_0 & ~i_8_241_939_0 & ~i_8_241_1285_0 & ~i_8_241_1291_0 & i_8_241_1651_0 & ~i_8_241_1779_0 & ~i_8_241_1883_0 & ~i_8_241_2040_0 & ~i_8_241_2070_0 & ~i_8_241_2157_0 & ~i_8_241_2262_0))) | (i_8_241_327_0 & i_8_241_393_0 & ~i_8_241_853_0 & ~i_8_241_1294_0 & ~i_8_241_1444_0 & ~i_8_241_1827_0 & ~i_8_241_1830_0) | (i_8_241_842_0 & ~i_8_241_844_0 & i_8_241_878_0 & ~i_8_241_937_0 & ~i_8_241_1408_0 & ~i_8_241_1473_0 & ~i_8_241_1638_0 & ~i_8_241_1883_0 & ~i_8_241_2218_0))) | (~i_8_241_2157_0 & ((~i_8_241_238_0 & ~i_8_241_1473_0 & ((~i_8_241_190_0 & ~i_8_241_849_0 & ~i_8_241_877_0 & i_8_241_1050_0 & ~i_8_241_1680_0 & ~i_8_241_1779_0 & ~i_8_241_2173_0) | (~i_8_241_189_0 & ~i_8_241_258_0 & ~i_8_241_878_0 & ~i_8_241_1240_0 & ~i_8_241_1285_0 & i_8_241_1510_0 & ~i_8_241_1883_0 & ~i_8_241_2040_0 & ~i_8_241_2239_0))) | (~i_8_241_192_0 & ~i_8_241_325_0 & ~i_8_241_1291_0 & ~i_8_241_1407_0 & ~i_8_241_1437_0 & ~i_8_241_1638_0 & ~i_8_241_1830_0 & ~i_8_241_2070_0 & i_8_241_2091_0 & ~i_8_241_2158_0) | (~i_8_241_237_0 & ~i_8_241_328_0 & i_8_241_781_0 & ~i_8_241_875_0 & ~i_8_241_1050_0 & ~i_8_241_1545_0 & ~i_8_241_1883_0 & ~i_8_241_2040_0 & ~i_8_241_2091_0 & ~i_8_241_2218_0))) | (~i_8_241_1437_0 & ~i_8_241_1881_0 & ((~i_8_241_327_0 & i_8_241_877_0 & ~i_8_241_878_0 & i_8_241_1285_0 & ~i_8_241_2158_0 & ~i_8_241_2238_0) | (~i_8_241_618_0 & i_8_241_837_0 & ~i_8_241_862_0 & ~i_8_241_937_0 & i_8_241_1038_0 & ~i_8_241_1827_0 & ~i_8_241_2262_0))) | (~i_8_241_258_0 & ~i_8_241_665_0 & ~i_8_241_696_0 & ~i_8_241_996_0 & ~i_8_241_1290_0 & ~i_8_241_1294_0 & ~i_8_241_1530_0 & ~i_8_241_1638_0 & ~i_8_241_1647_0 & i_8_241_1680_0 & ~i_8_241_1769_0 & ~i_8_241_1822_0 & ~i_8_241_1883_0 & ~i_8_241_2262_0))) | (~i_8_241_194_0 & ((~i_8_241_63_0 & ~i_8_241_874_0 & i_8_241_1029_0 & ~i_8_241_1231_0 & ~i_8_241_1648_0 & ~i_8_241_1815_0 & ~i_8_241_2173_0) | (~i_8_241_36_0 & ~i_8_241_191_0 & i_8_241_716_0 & ~i_8_241_875_0 & ~i_8_241_1291_0 & ~i_8_241_1294_0 & ~i_8_241_1315_0 & ~i_8_241_1651_0 & ~i_8_241_2218_0))) | (~i_8_241_237_0 & ((~i_8_241_258_0 & ~i_8_241_996_0 & i_8_241_1284_0 & i_8_241_1545_0 & ~i_8_241_1779_0 & ~i_8_241_1881_0) | (~i_8_241_300_0 & ~i_8_241_327_0 & ~i_8_241_328_0 & ~i_8_241_861_0 & i_8_241_1231_0 & i_8_241_1267_0 & ~i_8_241_1285_0 & ~i_8_241_1291_0 & ~i_8_241_1315_0 & ~i_8_241_1407_0 & ~i_8_241_1647_0 & ~i_8_241_2091_0))) | (i_8_241_325_0 & ((i_8_241_194_0 & ~i_8_241_696_0 & ~i_8_241_844_0 & i_8_241_1030_0 & ~i_8_241_1830_0) | (~i_8_241_63_0 & ~i_8_241_189_0 & i_8_241_874_0 & ~i_8_241_1290_0 & ~i_8_241_1648_0 & ~i_8_241_1651_0 & ~i_8_241_1827_0 & ~i_8_241_2037_0))) | (~i_8_241_1648_0 & ((~i_8_241_853_0 & ((~i_8_241_191_0 & ((i_8_241_194_0 & ~i_8_241_258_0 & ~i_8_241_615_0 & ~i_8_241_716_0 & ~i_8_241_1263_0 & ~i_8_241_1315_0 & ~i_8_241_1492_0 & ~i_8_241_1680_0) | (~i_8_241_665_0 & ~i_8_241_1408_0 & ~i_8_241_1750_0 & ~i_8_241_1822_0 & ~i_8_241_1883_0 & i_8_241_2156_0 & ~i_8_241_2238_0))) | (~i_8_241_63_0 & ~i_8_241_189_0 & i_8_241_300_0 & ~i_8_241_878_0 & ~i_8_241_939_0 & ~i_8_241_1290_0 & ~i_8_241_1294_0 & ~i_8_241_1779_0 & ~i_8_241_2037_0 & ~i_8_241_2040_0 & ~i_8_241_2173_0))) | (~i_8_241_615_0 & ~i_8_241_1291_0 & ((~i_8_241_996_0 & ~i_8_241_1029_0 & i_8_241_1510_0 & ~i_8_241_1680_0 & i_8_241_1750_0 & ~i_8_241_2040_0) | (~i_8_241_223_0 & ~i_8_241_327_0 & ~i_8_241_328_0 & i_8_241_1240_0 & ~i_8_241_1437_0 & ~i_8_241_1492_0 & ~i_8_241_1815_0 & i_8_241_2156_0))) | (i_8_241_842_0 & ~i_8_241_1285_0 & ((i_8_241_328_0 & ~i_8_241_665_0 & ~i_8_241_696_0 & ~i_8_241_1883_0) | (~i_8_241_190_0 & i_8_241_194_0 & ~i_8_241_300_0 & ~i_8_241_325_0 & ~i_8_241_2158_0 & ~i_8_241_2238_0 & ~i_8_241_844_0 & ~i_8_241_1284_0))) | (~i_8_241_696_0 & ((i_8_241_875_0 & ~i_8_241_1294_0 & ~i_8_241_1407_0 & i_8_241_1769_0) | (~i_8_241_878_0 & ~i_8_241_1029_0 & i_8_241_1030_0 & ~i_8_241_1263_0 & ~i_8_241_1315_0 & ~i_8_241_1822_0 & ~i_8_241_2173_0 & ~i_8_241_2239_0))) | (~i_8_241_1815_0 & ((i_8_241_223_0 & i_8_241_781_0 & ~i_8_241_844_0 & ~i_8_241_862_0 & ~i_8_241_1651_0 & ~i_8_241_1830_0 & ~i_8_241_2040_0) | (~i_8_241_36_0 & i_8_241_716_0 & i_8_241_875_0 & ~i_8_241_2239_0))))) | (~i_8_241_63_0 & ((i_8_241_300_0 & ((~i_8_241_937_0 & ~i_8_241_1240_0 & ~i_8_241_1290_0 & ~i_8_241_1408_0 & ~i_8_241_1437_0 & ~i_8_241_2070_0 & ~i_8_241_2218_0) | (~i_8_241_615_0 & ~i_8_241_696_0 & ~i_8_241_862_0 & i_8_241_877_0 & ~i_8_241_1267_0 & ~i_8_241_1315_0 & ~i_8_241_1815_0 & ~i_8_241_2262_0))) | (~i_8_241_937_0 & ((~i_8_241_1883_0 & ((~i_8_241_190_0 & ~i_8_241_191_0 & ~i_8_241_238_0 & i_8_241_327_0 & ~i_8_241_1231_0 & ~i_8_241_1290_0 & ~i_8_241_1294_0 & ~i_8_241_1815_0 & ~i_8_241_2070_0 & ~i_8_241_2238_0) | (i_8_241_716_0 & ~i_8_241_853_0 & ~i_8_241_1267_0 & ~i_8_241_1444_0 & ~i_8_241_2173_0 & ~i_8_241_2239_0 & ~i_8_241_2037_0 & ~i_8_241_2157_0))) | (i_8_241_193_0 & i_8_241_328_0 & ~i_8_241_665_0 & ~i_8_241_2157_0 & ~i_8_241_2262_0 & ~i_8_241_1263_0 & ~i_8_241_1530_0))) | (~i_8_241_189_0 & ~i_8_241_861_0 & i_8_241_1158_0 & ~i_8_241_1647_0 & i_8_241_1779_0 & ~i_8_241_2037_0 & ~i_8_241_2156_0 & ~i_8_241_2262_0))) | (i_8_241_878_0 & ((~i_8_241_238_0 & ((~i_8_241_862_0 & ~i_8_241_1263_0 & ~i_8_241_1407_0 & i_8_241_1768_0 & ~i_8_241_1822_0 & ~i_8_241_1881_0) | (~i_8_241_191_0 & ~i_8_241_327_0 & ~i_8_241_529_0 & i_8_241_877_0 & ~i_8_241_937_0 & ~i_8_241_1269_0 & ~i_8_241_1294_0 & ~i_8_241_1530_0 & ~i_8_241_1827_0 & ~i_8_241_1883_0 & ~i_8_241_2070_0 & ~i_8_241_2239_0 & ~i_8_241_2262_0))) | (i_8_241_223_0 & i_8_241_1050_0 & ~i_8_241_1408_0 & ~i_8_241_1815_0 & ~i_8_241_2040_0) | (~i_8_241_996_0 & ~i_8_241_1290_0 & ~i_8_241_190_0 & i_8_241_874_0 & ~i_8_241_1530_0 & ~i_8_241_1651_0 & ~i_8_241_2156_0 & ~i_8_241_2158_0))) | (~i_8_241_2158_0 & ((~i_8_241_36_0 & ~i_8_241_939_0 & ((~i_8_241_1290_0 & i_8_241_1768_0 & i_8_241_1769_0 & ~i_8_241_1883_0) | (i_8_241_193_0 & i_8_241_844_0 & ~i_8_241_937_0 & i_8_241_1050_0 & ~i_8_241_1510_0 & ~i_8_241_2238_0))) | (~i_8_241_190_0 & ~i_8_241_2037_0 & ((i_8_241_193_0 & ~i_8_241_258_0 & ~i_8_241_628_0 & ~i_8_241_696_0 & ~i_8_241_1267_0 & ~i_8_241_1408_0 & ~i_8_241_1530_0) | (~i_8_241_878_0 & ~i_8_241_996_0 & i_8_241_1015_0 & ~i_8_241_1444_0 & ~i_8_241_1750_0 & ~i_8_241_2157_0))) | (~i_8_241_193_0 & ~i_8_241_258_0 & ~i_8_241_861_0 & i_8_241_1240_0 & ~i_8_241_1291_0 & ~i_8_241_1294_0 & ~i_8_241_1315_0 & i_8_241_1510_0 & ~i_8_241_1700_0) | (i_8_241_223_0 & ~i_8_241_1050_0 & i_8_241_1267_0 & ~i_8_241_1492_0 & ~i_8_241_1769_0 & i_8_241_1822_0 & ~i_8_241_2173_0 & ~i_8_241_2238_0))) | (~i_8_241_2040_0 & ((~i_8_241_258_0 & ((i_8_241_327_0 & i_8_241_624_0 & ~i_8_241_1815_0 & ~i_8_241_1830_0) | (i_8_241_192_0 & i_8_241_193_0 & ~i_8_241_862_0 & ~i_8_241_1050_0 & ~i_8_241_1651_0 & ~i_8_241_1769_0 & ~i_8_241_2037_0))) | (~i_8_241_189_0 & i_8_241_328_0 & ~i_8_241_393_0 & ~i_8_241_1294_0 & ~i_8_241_1408_0 & i_8_241_1492_0 & ~i_8_241_1769_0 & ~i_8_241_2037_0 & ~i_8_241_2156_0))) | (~i_8_241_189_0 & ((~i_8_241_36_0 & ~i_8_241_191_0 & i_8_241_360_0 & ~i_8_241_1029_0 & ~i_8_241_1038_0 & ~i_8_241_1284_0 & ~i_8_241_1530_0 & ~i_8_241_1638_0 & ~i_8_241_1651_0 & ~i_8_241_1680_0 & ~i_8_241_2218_0) | (i_8_241_223_0 & ~i_8_241_696_0 & ~i_8_241_874_0 & i_8_241_1015_0 & ~i_8_241_1815_0 & ~i_8_241_2239_0))) | (~i_8_241_191_0 & ((i_8_241_223_0 & ((~i_8_241_1315_0 & i_8_241_1769_0 & i_8_241_1883_0) | (~i_8_241_618_0 & i_8_241_842_0 & ~i_8_241_853_0 & ~i_8_241_1883_0))) | (~i_8_241_1651_0 & ((i_8_241_328_0 & i_8_241_842_0 & i_8_241_1768_0 & ~i_8_241_1779_0) | (i_8_241_624_0 & ~i_8_241_696_0 & ~i_8_241_861_0 & ~i_8_241_1881_0 & ~i_8_241_2239_0))))) | (~i_8_241_2239_0 & ((~i_8_241_1647_0 & ((~i_8_241_1291_0 & ((i_8_241_393_0 & i_8_241_529_0 & ~i_8_241_1284_0 & ~i_8_241_1290_0 & ~i_8_241_1844_0) | (~i_8_241_696_0 & ~i_8_241_996_0 & ~i_8_241_1269_0 & ~i_8_241_1294_0 & ~i_8_241_1408_0 & i_8_241_1444_0 & ~i_8_241_1883_0))) | (~i_8_241_844_0 & ~i_8_241_1285_0 & ~i_8_241_1294_0 & i_8_241_1700_0 & ~i_8_241_1822_0))) | (~i_8_241_618_0 & ~i_8_241_1291_0 & ~i_8_241_1315_0 & i_8_241_1769_0 & ~i_8_241_1827_0 & ~i_8_241_1830_0 & ~i_8_241_1881_0 & ~i_8_241_1883_0 & ~i_8_241_2157_0))) | (i_8_241_327_0 & ~i_8_241_328_0 & ~i_8_241_615_0 & ~i_8_241_937_0 & ~i_8_241_1038_0 & ~i_8_241_1267_0 & i_8_241_1647_0 & i_8_241_1822_0));
endmodule



// Benchmark "kernel_8_242" written by ABC on Sun Jul 19 10:07:17 2020

module kernel_8_242 ( 
    i_8_242_67_0, i_8_242_75_0, i_8_242_76_0, i_8_242_120_0, i_8_242_125_0,
    i_8_242_138_0, i_8_242_169_0, i_8_242_192_0, i_8_242_195_0,
    i_8_242_196_0, i_8_242_198_0, i_8_242_225_0, i_8_242_228_0,
    i_8_242_229_0, i_8_242_261_0, i_8_242_301_0, i_8_242_312_0,
    i_8_242_324_0, i_8_242_354_0, i_8_242_355_0, i_8_242_402_0,
    i_8_242_417_0, i_8_242_433_0, i_8_242_522_0, i_8_242_556_0,
    i_8_242_571_0, i_8_242_586_0, i_8_242_588_0, i_8_242_634_0,
    i_8_242_657_0, i_8_242_660_0, i_8_242_671_0, i_8_242_672_0,
    i_8_242_697_0, i_8_242_709_0, i_8_242_732_0, i_8_242_747_0,
    i_8_242_753_0, i_8_242_782_0, i_8_242_831_0, i_8_242_835_0,
    i_8_242_837_0, i_8_242_838_0, i_8_242_840_0, i_8_242_858_0,
    i_8_242_925_0, i_8_242_943_0, i_8_242_969_0, i_8_242_970_0,
    i_8_242_971_0, i_8_242_973_0, i_8_242_983_0, i_8_242_985_0,
    i_8_242_990_0, i_8_242_993_0, i_8_242_1003_0, i_8_242_1038_0,
    i_8_242_1129_0, i_8_242_1138_0, i_8_242_1144_0, i_8_242_1266_0,
    i_8_242_1282_0, i_8_242_1293_0, i_8_242_1299_0, i_8_242_1300_0,
    i_8_242_1368_0, i_8_242_1390_0, i_8_242_1445_0, i_8_242_1452_0,
    i_8_242_1457_0, i_8_242_1470_0, i_8_242_1480_0, i_8_242_1486_0,
    i_8_242_1524_0, i_8_242_1549_0, i_8_242_1551_0, i_8_242_1573_0,
    i_8_242_1605_0, i_8_242_1633_0, i_8_242_1641_0, i_8_242_1651_0,
    i_8_242_1663_0, i_8_242_1849_0, i_8_242_1857_0, i_8_242_1922_0,
    i_8_242_1938_0, i_8_242_1946_0, i_8_242_1965_0, i_8_242_1968_0,
    i_8_242_1983_0, i_8_242_1995_0, i_8_242_2025_0, i_8_242_2053_0,
    i_8_242_2073_0, i_8_242_2082_0, i_8_242_2146_0, i_8_242_2191_0,
    i_8_242_2232_0, i_8_242_2233_0, i_8_242_2276_0,
    o_8_242_0_0  );
  input  i_8_242_67_0, i_8_242_75_0, i_8_242_76_0, i_8_242_120_0,
    i_8_242_125_0, i_8_242_138_0, i_8_242_169_0, i_8_242_192_0,
    i_8_242_195_0, i_8_242_196_0, i_8_242_198_0, i_8_242_225_0,
    i_8_242_228_0, i_8_242_229_0, i_8_242_261_0, i_8_242_301_0,
    i_8_242_312_0, i_8_242_324_0, i_8_242_354_0, i_8_242_355_0,
    i_8_242_402_0, i_8_242_417_0, i_8_242_433_0, i_8_242_522_0,
    i_8_242_556_0, i_8_242_571_0, i_8_242_586_0, i_8_242_588_0,
    i_8_242_634_0, i_8_242_657_0, i_8_242_660_0, i_8_242_671_0,
    i_8_242_672_0, i_8_242_697_0, i_8_242_709_0, i_8_242_732_0,
    i_8_242_747_0, i_8_242_753_0, i_8_242_782_0, i_8_242_831_0,
    i_8_242_835_0, i_8_242_837_0, i_8_242_838_0, i_8_242_840_0,
    i_8_242_858_0, i_8_242_925_0, i_8_242_943_0, i_8_242_969_0,
    i_8_242_970_0, i_8_242_971_0, i_8_242_973_0, i_8_242_983_0,
    i_8_242_985_0, i_8_242_990_0, i_8_242_993_0, i_8_242_1003_0,
    i_8_242_1038_0, i_8_242_1129_0, i_8_242_1138_0, i_8_242_1144_0,
    i_8_242_1266_0, i_8_242_1282_0, i_8_242_1293_0, i_8_242_1299_0,
    i_8_242_1300_0, i_8_242_1368_0, i_8_242_1390_0, i_8_242_1445_0,
    i_8_242_1452_0, i_8_242_1457_0, i_8_242_1470_0, i_8_242_1480_0,
    i_8_242_1486_0, i_8_242_1524_0, i_8_242_1549_0, i_8_242_1551_0,
    i_8_242_1573_0, i_8_242_1605_0, i_8_242_1633_0, i_8_242_1641_0,
    i_8_242_1651_0, i_8_242_1663_0, i_8_242_1849_0, i_8_242_1857_0,
    i_8_242_1922_0, i_8_242_1938_0, i_8_242_1946_0, i_8_242_1965_0,
    i_8_242_1968_0, i_8_242_1983_0, i_8_242_1995_0, i_8_242_2025_0,
    i_8_242_2053_0, i_8_242_2073_0, i_8_242_2082_0, i_8_242_2146_0,
    i_8_242_2191_0, i_8_242_2232_0, i_8_242_2233_0, i_8_242_2276_0;
  output o_8_242_0_0;
  assign o_8_242_0_0 = ~((~i_8_242_120_0 & ((~i_8_242_192_0 & ~i_8_242_1368_0 & ~i_8_242_1524_0) | (~i_8_242_198_0 & ~i_8_242_990_0 & ~i_8_242_1605_0 & ~i_8_242_2073_0))) | (~i_8_242_196_0 & ((~i_8_242_732_0 & ~i_8_242_925_0 & ~i_8_242_970_0 & ~i_8_242_1651_0 & ~i_8_242_1995_0) | (~i_8_242_634_0 & ~i_8_242_660_0 & ~i_8_242_1368_0 & ~i_8_242_1480_0 & ~i_8_242_1641_0 & ~i_8_242_2233_0))) | (~i_8_242_225_0 & ((~i_8_242_753_0 & i_8_242_837_0 & ~i_8_242_990_0) | (~i_8_242_76_0 & ~i_8_242_192_0 & ~i_8_242_198_0 & ~i_8_242_402_0 & ~i_8_242_586_0 & ~i_8_242_671_0 & i_8_242_1038_0 & ~i_8_242_1144_0 & ~i_8_242_1266_0 & ~i_8_242_1605_0))) | (~i_8_242_417_0 & ((i_8_242_75_0 & ~i_8_242_993_0) | (~i_8_242_195_0 & ~i_8_242_672_0 & ~i_8_242_985_0 & ~i_8_242_1144_0 & ~i_8_242_1368_0))) | (~i_8_242_312_0 & ((~i_8_242_671_0 & ((~i_8_242_831_0 & ~i_8_242_1452_0 & ~i_8_242_1965_0) | (~i_8_242_522_0 & ~i_8_242_586_0 & ~i_8_242_1549_0 & ~i_8_242_1651_0 & ~i_8_242_2082_0))) | (i_8_242_196_0 & ~i_8_242_969_0 & ~i_8_242_1129_0 & ~i_8_242_1983_0))) | (~i_8_242_1038_0 & (~i_8_242_1857_0 | (~i_8_242_747_0 & ~i_8_242_1486_0 & ~i_8_242_1524_0))) | (i_8_242_67_0 & i_8_242_971_0) | (~i_8_242_782_0 & ~i_8_242_835_0 & ~i_8_242_840_0 & ~i_8_242_1138_0 & i_8_242_1857_0 & ~i_8_242_1938_0 & i_8_242_1965_0) | (~i_8_242_1857_0 & ~i_8_242_1968_0 & ~i_8_242_1983_0) | (i_8_242_672_0 & i_8_242_1129_0 & ~i_8_242_2073_0));
endmodule



// Benchmark "kernel_8_243" written by ABC on Sun Jul 19 10:07:18 2020

module kernel_8_243 ( 
    i_8_243_39_0, i_8_243_42_0, i_8_243_49_0, i_8_243_58_0, i_8_243_82_0,
    i_8_243_115_0, i_8_243_117_0, i_8_243_148_0, i_8_243_151_0,
    i_8_243_166_0, i_8_243_221_0, i_8_243_241_0, i_8_243_273_0,
    i_8_243_275_0, i_8_243_343_0, i_8_243_356_0, i_8_243_370_0,
    i_8_243_432_0, i_8_243_444_0, i_8_243_453_0, i_8_243_461_0,
    i_8_243_476_0, i_8_243_477_0, i_8_243_517_0, i_8_243_523_0,
    i_8_243_524_0, i_8_243_545_0, i_8_243_621_0, i_8_243_667_0,
    i_8_243_668_0, i_8_243_712_0, i_8_243_760_0, i_8_243_769_0,
    i_8_243_776_0, i_8_243_790_0, i_8_243_805_0, i_8_243_813_0,
    i_8_243_861_0, i_8_243_868_0, i_8_243_923_0, i_8_243_944_0,
    i_8_243_993_0, i_8_243_1160_0, i_8_243_1184_0, i_8_243_1201_0,
    i_8_243_1254_0, i_8_243_1281_0, i_8_243_1282_0, i_8_243_1300_0,
    i_8_243_1301_0, i_8_243_1356_0, i_8_243_1382_0, i_8_243_1387_0,
    i_8_243_1435_0, i_8_243_1497_0, i_8_243_1498_0, i_8_243_1535_0,
    i_8_243_1542_0, i_8_243_1543_0, i_8_243_1585_0, i_8_243_1587_0,
    i_8_243_1588_0, i_8_243_1595_0, i_8_243_1604_0, i_8_243_1622_0,
    i_8_243_1650_0, i_8_243_1676_0, i_8_243_1681_0, i_8_243_1688_0,
    i_8_243_1720_0, i_8_243_1753_0, i_8_243_1759_0, i_8_243_1762_0,
    i_8_243_1808_0, i_8_243_1814_0, i_8_243_1848_0, i_8_243_1855_0,
    i_8_243_1872_0, i_8_243_1886_0, i_8_243_1945_0, i_8_243_1946_0,
    i_8_243_1982_0, i_8_243_1993_0, i_8_243_2001_0, i_8_243_2028_0,
    i_8_243_2041_0, i_8_243_2072_0, i_8_243_2073_0, i_8_243_2093_0,
    i_8_243_2107_0, i_8_243_2108_0, i_8_243_2122_0, i_8_243_2123_0,
    i_8_243_2126_0, i_8_243_2174_0, i_8_243_2245_0, i_8_243_2246_0,
    i_8_243_2271_0, i_8_243_2299_0, i_8_243_2300_0,
    o_8_243_0_0  );
  input  i_8_243_39_0, i_8_243_42_0, i_8_243_49_0, i_8_243_58_0,
    i_8_243_82_0, i_8_243_115_0, i_8_243_117_0, i_8_243_148_0,
    i_8_243_151_0, i_8_243_166_0, i_8_243_221_0, i_8_243_241_0,
    i_8_243_273_0, i_8_243_275_0, i_8_243_343_0, i_8_243_356_0,
    i_8_243_370_0, i_8_243_432_0, i_8_243_444_0, i_8_243_453_0,
    i_8_243_461_0, i_8_243_476_0, i_8_243_477_0, i_8_243_517_0,
    i_8_243_523_0, i_8_243_524_0, i_8_243_545_0, i_8_243_621_0,
    i_8_243_667_0, i_8_243_668_0, i_8_243_712_0, i_8_243_760_0,
    i_8_243_769_0, i_8_243_776_0, i_8_243_790_0, i_8_243_805_0,
    i_8_243_813_0, i_8_243_861_0, i_8_243_868_0, i_8_243_923_0,
    i_8_243_944_0, i_8_243_993_0, i_8_243_1160_0, i_8_243_1184_0,
    i_8_243_1201_0, i_8_243_1254_0, i_8_243_1281_0, i_8_243_1282_0,
    i_8_243_1300_0, i_8_243_1301_0, i_8_243_1356_0, i_8_243_1382_0,
    i_8_243_1387_0, i_8_243_1435_0, i_8_243_1497_0, i_8_243_1498_0,
    i_8_243_1535_0, i_8_243_1542_0, i_8_243_1543_0, i_8_243_1585_0,
    i_8_243_1587_0, i_8_243_1588_0, i_8_243_1595_0, i_8_243_1604_0,
    i_8_243_1622_0, i_8_243_1650_0, i_8_243_1676_0, i_8_243_1681_0,
    i_8_243_1688_0, i_8_243_1720_0, i_8_243_1753_0, i_8_243_1759_0,
    i_8_243_1762_0, i_8_243_1808_0, i_8_243_1814_0, i_8_243_1848_0,
    i_8_243_1855_0, i_8_243_1872_0, i_8_243_1886_0, i_8_243_1945_0,
    i_8_243_1946_0, i_8_243_1982_0, i_8_243_1993_0, i_8_243_2001_0,
    i_8_243_2028_0, i_8_243_2041_0, i_8_243_2072_0, i_8_243_2073_0,
    i_8_243_2093_0, i_8_243_2107_0, i_8_243_2108_0, i_8_243_2122_0,
    i_8_243_2123_0, i_8_243_2126_0, i_8_243_2174_0, i_8_243_2245_0,
    i_8_243_2246_0, i_8_243_2271_0, i_8_243_2299_0, i_8_243_2300_0;
  output o_8_243_0_0;
  assign o_8_243_0_0 = 0;
endmodule



// Benchmark "kernel_8_244" written by ABC on Sun Jul 19 10:07:19 2020

module kernel_8_244 ( 
    i_8_244_0_0, i_8_244_78_0, i_8_244_84_0, i_8_244_94_0, i_8_244_103_0,
    i_8_244_120_0, i_8_244_126_0, i_8_244_135_0, i_8_244_156_0,
    i_8_244_184_0, i_8_244_190_0, i_8_244_217_0, i_8_244_255_0,
    i_8_244_297_0, i_8_244_328_0, i_8_244_364_0, i_8_244_381_0,
    i_8_244_451_0, i_8_244_454_0, i_8_244_480_0, i_8_244_493_0,
    i_8_244_525_0, i_8_244_544_0, i_8_244_549_0, i_8_244_553_0,
    i_8_244_561_0, i_8_244_580_0, i_8_244_589_0, i_8_244_595_0,
    i_8_244_610_0, i_8_244_622_0, i_8_244_628_0, i_8_244_631_0,
    i_8_244_640_0, i_8_244_661_0, i_8_244_679_0, i_8_244_682_0,
    i_8_244_715_0, i_8_244_718_0, i_8_244_733_0, i_8_244_786_0,
    i_8_244_792_0, i_8_244_832_0, i_8_244_841_0, i_8_244_842_0,
    i_8_244_847_0, i_8_244_850_0, i_8_244_911_0, i_8_244_964_0,
    i_8_244_967_0, i_8_244_976_0, i_8_244_1071_0, i_8_244_1072_0,
    i_8_244_1108_0, i_8_244_1111_0, i_8_244_1210_0, i_8_244_1255_0,
    i_8_244_1257_0, i_8_244_1264_0, i_8_244_1266_0, i_8_244_1270_0,
    i_8_244_1279_0, i_8_244_1297_0, i_8_244_1321_0, i_8_244_1326_0,
    i_8_244_1416_0, i_8_244_1435_0, i_8_244_1437_0, i_8_244_1438_0,
    i_8_244_1450_0, i_8_244_1453_0, i_8_244_1465_0, i_8_244_1551_0,
    i_8_244_1563_0, i_8_244_1564_0, i_8_244_1593_0, i_8_244_1625_0,
    i_8_244_1680_0, i_8_244_1722_0, i_8_244_1759_0, i_8_244_1762_0,
    i_8_244_1764_0, i_8_244_1802_0, i_8_244_1805_0, i_8_244_1809_0,
    i_8_244_1995_0, i_8_244_2026_0, i_8_244_2053_0, i_8_244_2116_0,
    i_8_244_2119_0, i_8_244_2125_0, i_8_244_2128_0, i_8_244_2223_0,
    i_8_244_2233_0, i_8_244_2242_0, i_8_244_2275_0, i_8_244_2280_0,
    i_8_244_2283_0, i_8_244_2286_0, i_8_244_2290_0,
    o_8_244_0_0  );
  input  i_8_244_0_0, i_8_244_78_0, i_8_244_84_0, i_8_244_94_0,
    i_8_244_103_0, i_8_244_120_0, i_8_244_126_0, i_8_244_135_0,
    i_8_244_156_0, i_8_244_184_0, i_8_244_190_0, i_8_244_217_0,
    i_8_244_255_0, i_8_244_297_0, i_8_244_328_0, i_8_244_364_0,
    i_8_244_381_0, i_8_244_451_0, i_8_244_454_0, i_8_244_480_0,
    i_8_244_493_0, i_8_244_525_0, i_8_244_544_0, i_8_244_549_0,
    i_8_244_553_0, i_8_244_561_0, i_8_244_580_0, i_8_244_589_0,
    i_8_244_595_0, i_8_244_610_0, i_8_244_622_0, i_8_244_628_0,
    i_8_244_631_0, i_8_244_640_0, i_8_244_661_0, i_8_244_679_0,
    i_8_244_682_0, i_8_244_715_0, i_8_244_718_0, i_8_244_733_0,
    i_8_244_786_0, i_8_244_792_0, i_8_244_832_0, i_8_244_841_0,
    i_8_244_842_0, i_8_244_847_0, i_8_244_850_0, i_8_244_911_0,
    i_8_244_964_0, i_8_244_967_0, i_8_244_976_0, i_8_244_1071_0,
    i_8_244_1072_0, i_8_244_1108_0, i_8_244_1111_0, i_8_244_1210_0,
    i_8_244_1255_0, i_8_244_1257_0, i_8_244_1264_0, i_8_244_1266_0,
    i_8_244_1270_0, i_8_244_1279_0, i_8_244_1297_0, i_8_244_1321_0,
    i_8_244_1326_0, i_8_244_1416_0, i_8_244_1435_0, i_8_244_1437_0,
    i_8_244_1438_0, i_8_244_1450_0, i_8_244_1453_0, i_8_244_1465_0,
    i_8_244_1551_0, i_8_244_1563_0, i_8_244_1564_0, i_8_244_1593_0,
    i_8_244_1625_0, i_8_244_1680_0, i_8_244_1722_0, i_8_244_1759_0,
    i_8_244_1762_0, i_8_244_1764_0, i_8_244_1802_0, i_8_244_1805_0,
    i_8_244_1809_0, i_8_244_1995_0, i_8_244_2026_0, i_8_244_2053_0,
    i_8_244_2116_0, i_8_244_2119_0, i_8_244_2125_0, i_8_244_2128_0,
    i_8_244_2223_0, i_8_244_2233_0, i_8_244_2242_0, i_8_244_2275_0,
    i_8_244_2280_0, i_8_244_2283_0, i_8_244_2286_0, i_8_244_2290_0;
  output o_8_244_0_0;
  assign o_8_244_0_0 = 0;
endmodule



// Benchmark "kernel_8_245" written by ABC on Sun Jul 19 10:07:19 2020

module kernel_8_245 ( 
    i_8_245_32_0, i_8_245_76_0, i_8_245_167_0, i_8_245_173_0,
    i_8_245_209_0, i_8_245_256_0, i_8_245_262_0, i_8_245_326_0,
    i_8_245_344_0, i_8_245_362_0, i_8_245_364_0, i_8_245_365_0,
    i_8_245_425_0, i_8_245_434_0, i_8_245_454_0, i_8_245_482_0,
    i_8_245_491_0, i_8_245_553_0, i_8_245_590_0, i_8_245_626_0,
    i_8_245_634_0, i_8_245_641_0, i_8_245_703_0, i_8_245_706_0,
    i_8_245_707_0, i_8_245_738_0, i_8_245_767_0, i_8_245_795_0,
    i_8_245_837_0, i_8_245_839_0, i_8_245_842_0, i_8_245_845_0,
    i_8_245_919_0, i_8_245_920_0, i_8_245_929_0, i_8_245_956_0,
    i_8_245_1055_0, i_8_245_1061_0, i_8_245_1067_0, i_8_245_1100_0,
    i_8_245_1114_0, i_8_245_1171_0, i_8_245_1172_0, i_8_245_1235_0,
    i_8_245_1264_0, i_8_245_1278_0, i_8_245_1282_0, i_8_245_1283_0,
    i_8_245_1316_0, i_8_245_1372_0, i_8_245_1379_0, i_8_245_1382_0,
    i_8_245_1413_0, i_8_245_1433_0, i_8_245_1478_0, i_8_245_1544_0,
    i_8_245_1559_0, i_8_245_1562_0, i_8_245_1565_0, i_8_245_1571_0,
    i_8_245_1613_0, i_8_245_1625_0, i_8_245_1633_0, i_8_245_1643_0,
    i_8_245_1685_0, i_8_245_1688_0, i_8_245_1694_0, i_8_245_1702_0,
    i_8_245_1703_0, i_8_245_1706_0, i_8_245_1711_0, i_8_245_1721_0,
    i_8_245_1765_0, i_8_245_1774_0, i_8_245_1775_0, i_8_245_1820_0,
    i_8_245_1821_0, i_8_245_1822_0, i_8_245_1832_0, i_8_245_1859_0,
    i_8_245_1863_0, i_8_245_1867_0, i_8_245_1882_0, i_8_245_1883_0,
    i_8_245_1982_0, i_8_245_2009_0, i_8_245_2017_0, i_8_245_2018_0,
    i_8_245_2108_0, i_8_245_2111_0, i_8_245_2144_0, i_8_245_2146_0,
    i_8_245_2147_0, i_8_245_2170_0, i_8_245_2192_0, i_8_245_2197_0,
    i_8_245_2198_0, i_8_245_2206_0, i_8_245_2242_0, i_8_245_2243_0,
    o_8_245_0_0  );
  input  i_8_245_32_0, i_8_245_76_0, i_8_245_167_0, i_8_245_173_0,
    i_8_245_209_0, i_8_245_256_0, i_8_245_262_0, i_8_245_326_0,
    i_8_245_344_0, i_8_245_362_0, i_8_245_364_0, i_8_245_365_0,
    i_8_245_425_0, i_8_245_434_0, i_8_245_454_0, i_8_245_482_0,
    i_8_245_491_0, i_8_245_553_0, i_8_245_590_0, i_8_245_626_0,
    i_8_245_634_0, i_8_245_641_0, i_8_245_703_0, i_8_245_706_0,
    i_8_245_707_0, i_8_245_738_0, i_8_245_767_0, i_8_245_795_0,
    i_8_245_837_0, i_8_245_839_0, i_8_245_842_0, i_8_245_845_0,
    i_8_245_919_0, i_8_245_920_0, i_8_245_929_0, i_8_245_956_0,
    i_8_245_1055_0, i_8_245_1061_0, i_8_245_1067_0, i_8_245_1100_0,
    i_8_245_1114_0, i_8_245_1171_0, i_8_245_1172_0, i_8_245_1235_0,
    i_8_245_1264_0, i_8_245_1278_0, i_8_245_1282_0, i_8_245_1283_0,
    i_8_245_1316_0, i_8_245_1372_0, i_8_245_1379_0, i_8_245_1382_0,
    i_8_245_1413_0, i_8_245_1433_0, i_8_245_1478_0, i_8_245_1544_0,
    i_8_245_1559_0, i_8_245_1562_0, i_8_245_1565_0, i_8_245_1571_0,
    i_8_245_1613_0, i_8_245_1625_0, i_8_245_1633_0, i_8_245_1643_0,
    i_8_245_1685_0, i_8_245_1688_0, i_8_245_1694_0, i_8_245_1702_0,
    i_8_245_1703_0, i_8_245_1706_0, i_8_245_1711_0, i_8_245_1721_0,
    i_8_245_1765_0, i_8_245_1774_0, i_8_245_1775_0, i_8_245_1820_0,
    i_8_245_1821_0, i_8_245_1822_0, i_8_245_1832_0, i_8_245_1859_0,
    i_8_245_1863_0, i_8_245_1867_0, i_8_245_1882_0, i_8_245_1883_0,
    i_8_245_1982_0, i_8_245_2009_0, i_8_245_2017_0, i_8_245_2018_0,
    i_8_245_2108_0, i_8_245_2111_0, i_8_245_2144_0, i_8_245_2146_0,
    i_8_245_2147_0, i_8_245_2170_0, i_8_245_2192_0, i_8_245_2197_0,
    i_8_245_2198_0, i_8_245_2206_0, i_8_245_2242_0, i_8_245_2243_0;
  output o_8_245_0_0;
  assign o_8_245_0_0 = 0;
endmodule



// Benchmark "kernel_8_246" written by ABC on Sun Jul 19 10:07:21 2020

module kernel_8_246 ( 
    i_8_246_114_0, i_8_246_186_0, i_8_246_241_0, i_8_246_294_0,
    i_8_246_295_0, i_8_246_296_0, i_8_246_303_0, i_8_246_304_0,
    i_8_246_321_0, i_8_246_337_0, i_8_246_348_0, i_8_246_350_0,
    i_8_246_364_0, i_8_246_453_0, i_8_246_458_0, i_8_246_488_0,
    i_8_246_553_0, i_8_246_554_0, i_8_246_590_0, i_8_246_597_0,
    i_8_246_599_0, i_8_246_613_0, i_8_246_614_0, i_8_246_615_0,
    i_8_246_617_0, i_8_246_619_0, i_8_246_645_0, i_8_246_672_0,
    i_8_246_689_0, i_8_246_705_0, i_8_246_710_0, i_8_246_717_0,
    i_8_246_778_0, i_8_246_799_0, i_8_246_851_0, i_8_246_872_0,
    i_8_246_875_0, i_8_246_878_0, i_8_246_969_0, i_8_246_970_0,
    i_8_246_990_0, i_8_246_991_0, i_8_246_1031_0, i_8_246_1072_0,
    i_8_246_1074_0, i_8_246_1108_0, i_8_246_1112_0, i_8_246_1113_0,
    i_8_246_1119_0, i_8_246_1120_0, i_8_246_1121_0, i_8_246_1122_0,
    i_8_246_1123_0, i_8_246_1124_0, i_8_246_1229_0, i_8_246_1282_0,
    i_8_246_1306_0, i_8_246_1329_0, i_8_246_1330_0, i_8_246_1331_0,
    i_8_246_1407_0, i_8_246_1408_0, i_8_246_1411_0, i_8_246_1437_0,
    i_8_246_1489_0, i_8_246_1490_0, i_8_246_1509_0, i_8_246_1511_0,
    i_8_246_1545_0, i_8_246_1619_0, i_8_246_1650_0, i_8_246_1654_0,
    i_8_246_1672_0, i_8_246_1675_0, i_8_246_1677_0, i_8_246_1679_0,
    i_8_246_1790_0, i_8_246_1803_0, i_8_246_1806_0, i_8_246_1815_0,
    i_8_246_1823_0, i_8_246_1826_0, i_8_246_1866_0, i_8_246_1876_0,
    i_8_246_1884_0, i_8_246_1885_0, i_8_246_1983_0, i_8_246_1986_0,
    i_8_246_1988_0, i_8_246_2028_0, i_8_246_2056_0, i_8_246_2075_0,
    i_8_246_2090_0, i_8_246_2131_0, i_8_246_2193_0, i_8_246_2194_0,
    i_8_246_2219_0, i_8_246_2228_0, i_8_246_2249_0, i_8_246_2272_0,
    o_8_246_0_0  );
  input  i_8_246_114_0, i_8_246_186_0, i_8_246_241_0, i_8_246_294_0,
    i_8_246_295_0, i_8_246_296_0, i_8_246_303_0, i_8_246_304_0,
    i_8_246_321_0, i_8_246_337_0, i_8_246_348_0, i_8_246_350_0,
    i_8_246_364_0, i_8_246_453_0, i_8_246_458_0, i_8_246_488_0,
    i_8_246_553_0, i_8_246_554_0, i_8_246_590_0, i_8_246_597_0,
    i_8_246_599_0, i_8_246_613_0, i_8_246_614_0, i_8_246_615_0,
    i_8_246_617_0, i_8_246_619_0, i_8_246_645_0, i_8_246_672_0,
    i_8_246_689_0, i_8_246_705_0, i_8_246_710_0, i_8_246_717_0,
    i_8_246_778_0, i_8_246_799_0, i_8_246_851_0, i_8_246_872_0,
    i_8_246_875_0, i_8_246_878_0, i_8_246_969_0, i_8_246_970_0,
    i_8_246_990_0, i_8_246_991_0, i_8_246_1031_0, i_8_246_1072_0,
    i_8_246_1074_0, i_8_246_1108_0, i_8_246_1112_0, i_8_246_1113_0,
    i_8_246_1119_0, i_8_246_1120_0, i_8_246_1121_0, i_8_246_1122_0,
    i_8_246_1123_0, i_8_246_1124_0, i_8_246_1229_0, i_8_246_1282_0,
    i_8_246_1306_0, i_8_246_1329_0, i_8_246_1330_0, i_8_246_1331_0,
    i_8_246_1407_0, i_8_246_1408_0, i_8_246_1411_0, i_8_246_1437_0,
    i_8_246_1489_0, i_8_246_1490_0, i_8_246_1509_0, i_8_246_1511_0,
    i_8_246_1545_0, i_8_246_1619_0, i_8_246_1650_0, i_8_246_1654_0,
    i_8_246_1672_0, i_8_246_1675_0, i_8_246_1677_0, i_8_246_1679_0,
    i_8_246_1790_0, i_8_246_1803_0, i_8_246_1806_0, i_8_246_1815_0,
    i_8_246_1823_0, i_8_246_1826_0, i_8_246_1866_0, i_8_246_1876_0,
    i_8_246_1884_0, i_8_246_1885_0, i_8_246_1983_0, i_8_246_1986_0,
    i_8_246_1988_0, i_8_246_2028_0, i_8_246_2056_0, i_8_246_2075_0,
    i_8_246_2090_0, i_8_246_2131_0, i_8_246_2193_0, i_8_246_2194_0,
    i_8_246_2219_0, i_8_246_2228_0, i_8_246_2249_0, i_8_246_2272_0;
  output o_8_246_0_0;
  assign o_8_246_0_0 = ~((~i_8_246_114_0 & ((~i_8_246_186_0 & ~i_8_246_295_0 & ~i_8_246_453_0 & ~i_8_246_878_0 & ~i_8_246_990_0 & i_8_246_1407_0) | (~i_8_246_348_0 & i_8_246_619_0 & ~i_8_246_689_0 & ~i_8_246_1072_0 & ~i_8_246_1120_0 & ~i_8_246_1330_0 & ~i_8_246_1331_0 & ~i_8_246_2193_0))) | (~i_8_246_1545_0 & ((~i_8_246_304_0 & ((~i_8_246_645_0 & i_8_246_1113_0 & ~i_8_246_1120_0 & ~i_8_246_1122_0 & i_8_246_1437_0) | (~i_8_246_303_0 & ~i_8_246_851_0 & ~i_8_246_1119_0 & ~i_8_246_1790_0 & ~i_8_246_1876_0 & ~i_8_246_1885_0 & i_8_246_1986_0))) | (~i_8_246_2194_0 & ((i_8_246_364_0 & ~i_8_246_1408_0 & ((~i_8_246_689_0 & ~i_8_246_1123_0 & i_8_246_1803_0 & ~i_8_246_1815_0) | (~i_8_246_878_0 & ~i_8_246_990_0 & ~i_8_246_1072_0 & ~i_8_246_1511_0 & ~i_8_246_1803_0 & ~i_8_246_2028_0 & ~i_8_246_2090_0))) | (~i_8_246_295_0 & ~i_8_246_458_0 & ~i_8_246_969_0 & ~i_8_246_1306_0 & i_8_246_1411_0 & ~i_8_246_1677_0 & ~i_8_246_1986_0 & ~i_8_246_2219_0))) | (i_8_246_617_0 & ((~i_8_246_878_0 & ~i_8_246_1124_0 & ~i_8_246_1331_0) | (~i_8_246_645_0 & ~i_8_246_799_0 & ~i_8_246_1120_0 & ~i_8_246_1306_0 & ~i_8_246_2075_0 & ~i_8_246_2131_0))) | (~i_8_246_296_0 & ~i_8_246_590_0 & ~i_8_246_689_0 & ~i_8_246_872_0 & ~i_8_246_875_0 & ~i_8_246_990_0 & ~i_8_246_1122_0 & ~i_8_246_1124_0 & ~i_8_246_1229_0 & i_8_246_1282_0 & ~i_8_246_1511_0 & ~i_8_246_2090_0 & ~i_8_246_2131_0) | (~i_8_246_294_0 & i_8_246_348_0 & ~i_8_246_672_0 & i_8_246_1509_0 & i_8_246_1650_0 & ~i_8_246_2193_0) | (~i_8_246_453_0 & ~i_8_246_597_0 & ~i_8_246_799_0 & ~i_8_246_1108_0 & i_8_246_1654_0 & ~i_8_246_1677_0 & ~i_8_246_1679_0 & ~i_8_246_1823_0 & ~i_8_246_2219_0))) | (~i_8_246_458_0 & ((~i_8_246_294_0 & ((~i_8_246_296_0 & ((~i_8_246_321_0 & i_8_246_337_0 & ~i_8_246_348_0 & ~i_8_246_453_0 & ~i_8_246_597_0 & ~i_8_246_1072_0 & ~i_8_246_2028_0) | (~i_8_246_186_0 & ~i_8_246_304_0 & ~i_8_246_672_0 & i_8_246_1411_0 & ~i_8_246_1509_0 & ~i_8_246_1511_0 & ~i_8_246_2131_0))) | (~i_8_246_453_0 & ~i_8_246_1331_0 & ((~i_8_246_645_0 & ~i_8_246_1124_0 & ~i_8_246_1490_0 & ~i_8_246_1509_0 & i_8_246_1803_0 & ~i_8_246_1823_0) | (~i_8_246_241_0 & ~i_8_246_295_0 & ~i_8_246_590_0 & ~i_8_246_689_0 & ~i_8_246_799_0 & ~i_8_246_969_0 & ~i_8_246_990_0 & ~i_8_246_991_0 & ~i_8_246_1411_0 & ~i_8_246_2028_0 & ~i_8_246_2056_0 & ~i_8_246_2075_0 & i_8_246_2131_0))))) | (~i_8_246_2194_0 & ((~i_8_246_350_0 & ((~i_8_246_488_0 & ~i_8_246_990_0 & ~i_8_246_1072_0 & i_8_246_1112_0 & ~i_8_246_1120_0 & ~i_8_246_1329_0 & ~i_8_246_1331_0 & ~i_8_246_1408_0 & ~i_8_246_1489_0) | (~i_8_246_599_0 & ~i_8_246_1108_0 & i_8_246_1282_0 & i_8_246_2219_0))) | (~i_8_246_645_0 & ~i_8_246_717_0 & ~i_8_246_990_0 & ~i_8_246_1121_0 & ~i_8_246_1329_0 & i_8_246_1437_0 & ~i_8_246_1490_0 & ~i_8_246_1823_0 & ~i_8_246_1866_0))) | (~i_8_246_304_0 & ~i_8_246_590_0 & ~i_8_246_599_0 & i_8_246_1108_0 & ~i_8_246_1437_0 & ~i_8_246_1679_0 & ~i_8_246_1876_0 & ~i_8_246_2028_0 & ~i_8_246_2193_0))) | (~i_8_246_186_0 & ((~i_8_246_296_0 & ((~i_8_246_321_0 & ~i_8_246_851_0 & ~i_8_246_1122_0 & ~i_8_246_1123_0 & ~i_8_246_1509_0 & i_8_246_1885_0) | (~i_8_246_303_0 & ~i_8_246_348_0 & ~i_8_246_991_0 & i_8_246_1408_0 & ~i_8_246_1490_0 & ~i_8_246_1803_0 & ~i_8_246_1986_0 & ~i_8_246_2028_0 & ~i_8_246_2090_0 & ~i_8_246_2194_0))) | (~i_8_246_321_0 & ~i_8_246_597_0 & ~i_8_246_599_0 & i_8_246_705_0 & ~i_8_246_1074_0 & ~i_8_246_1306_0 & ~i_8_246_1866_0) | (~i_8_246_672_0 & ~i_8_246_1509_0 & ~i_8_246_1511_0 & i_8_246_1650_0 & ~i_8_246_1885_0 & ~i_8_246_2028_0))) | (~i_8_246_689_0 & ((~i_8_246_453_0 & ((~i_8_246_295_0 & ~i_8_246_645_0 & i_8_246_1074_0 & ~i_8_246_1330_0 & ~i_8_246_1866_0 & ~i_8_246_2249_0) | (~i_8_246_619_0 & i_8_246_1072_0 & ~i_8_246_1876_0 & ~i_8_246_2090_0 & ~i_8_246_2219_0 & ~i_8_246_2272_0))) | (~i_8_246_597_0 & ((~i_8_246_778_0 & ~i_8_246_875_0 & ~i_8_246_1074_0 & ~i_8_246_1123_0 & i_8_246_1489_0) | (~i_8_246_348_0 & ~i_8_246_990_0 & ~i_8_246_1437_0 & i_8_246_1675_0 & ~i_8_246_1876_0 & ~i_8_246_2028_0))) | (i_8_246_114_0 & ~i_8_246_615_0 & ~i_8_246_645_0 & ~i_8_246_672_0 & ~i_8_246_851_0 & ~i_8_246_872_0 & ~i_8_246_991_0 & ~i_8_246_1074_0 & ~i_8_246_1330_0 & ~i_8_246_1650_0) | (~i_8_246_303_0 & ~i_8_246_614_0 & i_8_246_710_0 & i_8_246_1112_0 & ~i_8_246_1121_0 & ~i_8_246_2075_0 & ~i_8_246_2194_0))) | (~i_8_246_303_0 & ((i_8_246_1408_0 & i_8_246_1650_0 & i_8_246_1884_0) | (~i_8_246_599_0 & ~i_8_246_1306_0 & ~i_8_246_1329_0 & i_8_246_1983_0 & ~i_8_246_2090_0 & ~i_8_246_2219_0))) | (~i_8_246_348_0 & ((~i_8_246_296_0 & ~i_8_246_599_0 & i_8_246_1112_0 & ~i_8_246_1331_0 & ~i_8_246_1437_0 & i_8_246_1823_0) | (i_8_246_1108_0 & ~i_8_246_1121_0 & i_8_246_1675_0 & ~i_8_246_2028_0 & ~i_8_246_2193_0))) | (i_8_246_590_0 & ((~i_8_246_488_0 & ~i_8_246_1121_0 & ~i_8_246_1306_0 & ~i_8_246_2090_0 & ~i_8_246_2131_0 & ~i_8_246_1511_0 & ~i_8_246_1790_0) | (i_8_246_613_0 & ~i_8_246_799_0 & i_8_246_1282_0 & ~i_8_246_2193_0))) | (~i_8_246_488_0 & ((~i_8_246_599_0 & ~i_8_246_1123_0 & i_8_246_1619_0) | (~i_8_246_295_0 & ~i_8_246_296_0 & ~i_8_246_590_0 & ~i_8_246_705_0 & ~i_8_246_875_0 & ~i_8_246_1306_0 & ~i_8_246_1329_0 & i_8_246_1679_0 & ~i_8_246_1815_0 & ~i_8_246_1823_0 & ~i_8_246_1884_0 & ~i_8_246_1885_0))) | (~i_8_246_295_0 & ~i_8_246_1876_0 & ((~i_8_246_296_0 & i_8_246_554_0 & ~i_8_246_799_0 & ~i_8_246_851_0 & ~i_8_246_878_0 & ~i_8_246_1122_0 & ~i_8_246_1675_0 & ~i_8_246_1885_0) | (~i_8_246_590_0 & ~i_8_246_970_0 & i_8_246_1031_0 & ~i_8_246_1677_0 & i_8_246_1679_0 & ~i_8_246_1790_0 & ~i_8_246_2090_0))) | (~i_8_246_645_0 & ((~i_8_246_717_0 & ~i_8_246_875_0 & ~i_8_246_1031_0 & i_8_246_1677_0 & i_8_246_1983_0 & ~i_8_246_2090_0) | (~i_8_246_294_0 & ~i_8_246_296_0 & ~i_8_246_350_0 & ~i_8_246_553_0 & ~i_8_246_597_0 & ~i_8_246_990_0 & ~i_8_246_1122_0 & ~i_8_246_1306_0 & i_8_246_1329_0 & ~i_8_246_2194_0))) | (~i_8_246_2028_0 & ((~i_8_246_294_0 & ((~i_8_246_296_0 & ~i_8_246_597_0 & ~i_8_246_991_0 & ~i_8_246_1074_0 & ~i_8_246_1121_0 & i_8_246_1677_0) | (i_8_246_553_0 & i_8_246_1986_0 & ~i_8_246_2249_0))) | (i_8_246_614_0 & ~i_8_246_851_0 & ~i_8_246_1122_0 & ~i_8_246_2090_0))) | (~i_8_246_717_0 & ((~i_8_246_296_0 & ~i_8_246_991_0 & ~i_8_246_1031_0 & ~i_8_246_1121_0 & ~i_8_246_1282_0 & ~i_8_246_1675_0 & i_8_246_1988_0) | (i_8_246_878_0 & ~i_8_246_1229_0 & ~i_8_246_1330_0 & ~i_8_246_2194_0 & ~i_8_246_2219_0 & i_8_246_2249_0))) | (i_8_246_1823_0 & ((~i_8_246_1031_0 & i_8_246_2075_0) | (~i_8_246_350_0 & ~i_8_246_991_0 & ~i_8_246_1112_0 & ~i_8_246_1120_0 & ~i_8_246_1123_0 & i_8_246_1229_0 & ~i_8_246_1619_0 & ~i_8_246_1679_0 & ~i_8_246_2219_0))) | (~i_8_246_350_0 & ((~i_8_246_590_0 & i_8_246_613_0 & ~i_8_246_1072_0 & ~i_8_246_1122_0) | (~i_8_246_597_0 & ~i_8_246_851_0 & ~i_8_246_990_0 & i_8_246_1490_0 & ~i_8_246_1806_0 & ~i_8_246_2090_0))) | (i_8_246_710_0 & ~i_8_246_1074_0 & ~i_8_246_1121_0 & ~i_8_246_1124_0 & ~i_8_246_1330_0 & i_8_246_1826_0) | (~i_8_246_1282_0 & ~i_8_246_1329_0 & i_8_246_1677_0 & i_8_246_1866_0 & ~i_8_246_2090_0) | (i_8_246_2056_0 & ~i_8_246_2131_0 & i_8_246_2194_0 & i_8_246_2272_0));
endmodule



// Benchmark "kernel_8_247" written by ABC on Sun Jul 19 10:07:22 2020

module kernel_8_247 ( 
    i_8_247_52_0, i_8_247_76_0, i_8_247_80_0, i_8_247_104_0, i_8_247_107_0,
    i_8_247_166_0, i_8_247_169_0, i_8_247_219_0, i_8_247_225_0,
    i_8_247_228_0, i_8_247_257_0, i_8_247_323_0, i_8_247_368_0,
    i_8_247_382_0, i_8_247_427_0, i_8_247_436_0, i_8_247_440_0,
    i_8_247_450_0, i_8_247_489_0, i_8_247_490_0, i_8_247_491_0,
    i_8_247_492_0, i_8_247_548_0, i_8_247_556_0, i_8_247_581_0,
    i_8_247_587_0, i_8_247_626_0, i_8_247_635_0, i_8_247_658_0,
    i_8_247_661_0, i_8_247_679_0, i_8_247_693_0, i_8_247_694_0,
    i_8_247_695_0, i_8_247_698_0, i_8_247_699_0, i_8_247_716_0,
    i_8_247_723_0, i_8_247_724_0, i_8_247_725_0, i_8_247_805_0,
    i_8_247_809_0, i_8_247_812_0, i_8_247_833_0, i_8_247_840_0,
    i_8_247_851_0, i_8_247_955_0, i_8_247_970_0, i_8_247_977_0,
    i_8_247_1031_0, i_8_247_1076_0, i_8_247_1111_0, i_8_247_1115_0,
    i_8_247_1184_0, i_8_247_1192_0, i_8_247_1210_0, i_8_247_1211_0,
    i_8_247_1226_0, i_8_247_1234_0, i_8_247_1255_0, i_8_247_1273_0,
    i_8_247_1280_0, i_8_247_1300_0, i_8_247_1301_0, i_8_247_1328_0,
    i_8_247_1360_0, i_8_247_1373_0, i_8_247_1391_0, i_8_247_1456_0,
    i_8_247_1471_0, i_8_247_1472_0, i_8_247_1577_0, i_8_247_1748_0,
    i_8_247_1773_0, i_8_247_1786_0, i_8_247_1789_0, i_8_247_1790_0,
    i_8_247_1818_0, i_8_247_1849_0, i_8_247_1850_0, i_8_247_1858_0,
    i_8_247_1867_0, i_8_247_1901_0, i_8_247_1904_0, i_8_247_1907_0,
    i_8_247_1979_0, i_8_247_1982_0, i_8_247_1996_0, i_8_247_2003_0,
    i_8_247_2029_0, i_8_247_2032_0, i_8_247_2038_0, i_8_247_2133_0,
    i_8_247_2134_0, i_8_247_2191_0, i_8_247_2200_0, i_8_247_2214_0,
    i_8_247_2223_0, i_8_247_2224_0, i_8_247_2273_0,
    o_8_247_0_0  );
  input  i_8_247_52_0, i_8_247_76_0, i_8_247_80_0, i_8_247_104_0,
    i_8_247_107_0, i_8_247_166_0, i_8_247_169_0, i_8_247_219_0,
    i_8_247_225_0, i_8_247_228_0, i_8_247_257_0, i_8_247_323_0,
    i_8_247_368_0, i_8_247_382_0, i_8_247_427_0, i_8_247_436_0,
    i_8_247_440_0, i_8_247_450_0, i_8_247_489_0, i_8_247_490_0,
    i_8_247_491_0, i_8_247_492_0, i_8_247_548_0, i_8_247_556_0,
    i_8_247_581_0, i_8_247_587_0, i_8_247_626_0, i_8_247_635_0,
    i_8_247_658_0, i_8_247_661_0, i_8_247_679_0, i_8_247_693_0,
    i_8_247_694_0, i_8_247_695_0, i_8_247_698_0, i_8_247_699_0,
    i_8_247_716_0, i_8_247_723_0, i_8_247_724_0, i_8_247_725_0,
    i_8_247_805_0, i_8_247_809_0, i_8_247_812_0, i_8_247_833_0,
    i_8_247_840_0, i_8_247_851_0, i_8_247_955_0, i_8_247_970_0,
    i_8_247_977_0, i_8_247_1031_0, i_8_247_1076_0, i_8_247_1111_0,
    i_8_247_1115_0, i_8_247_1184_0, i_8_247_1192_0, i_8_247_1210_0,
    i_8_247_1211_0, i_8_247_1226_0, i_8_247_1234_0, i_8_247_1255_0,
    i_8_247_1273_0, i_8_247_1280_0, i_8_247_1300_0, i_8_247_1301_0,
    i_8_247_1328_0, i_8_247_1360_0, i_8_247_1373_0, i_8_247_1391_0,
    i_8_247_1456_0, i_8_247_1471_0, i_8_247_1472_0, i_8_247_1577_0,
    i_8_247_1748_0, i_8_247_1773_0, i_8_247_1786_0, i_8_247_1789_0,
    i_8_247_1790_0, i_8_247_1818_0, i_8_247_1849_0, i_8_247_1850_0,
    i_8_247_1858_0, i_8_247_1867_0, i_8_247_1901_0, i_8_247_1904_0,
    i_8_247_1907_0, i_8_247_1979_0, i_8_247_1982_0, i_8_247_1996_0,
    i_8_247_2003_0, i_8_247_2029_0, i_8_247_2032_0, i_8_247_2038_0,
    i_8_247_2133_0, i_8_247_2134_0, i_8_247_2191_0, i_8_247_2200_0,
    i_8_247_2214_0, i_8_247_2223_0, i_8_247_2224_0, i_8_247_2273_0;
  output o_8_247_0_0;
  assign o_8_247_0_0 = 0;
endmodule



// Benchmark "kernel_8_248" written by ABC on Sun Jul 19 10:07:23 2020

module kernel_8_248 ( 
    i_8_248_31_0, i_8_248_39_0, i_8_248_42_0, i_8_248_51_0, i_8_248_55_0,
    i_8_248_96_0, i_8_248_97_0, i_8_248_169_0, i_8_248_256_0,
    i_8_248_258_0, i_8_248_300_0, i_8_248_307_0, i_8_248_319_0,
    i_8_248_331_0, i_8_248_334_0, i_8_248_360_0, i_8_248_363_0,
    i_8_248_417_0, i_8_248_418_0, i_8_248_421_0, i_8_248_440_0,
    i_8_248_481_0, i_8_248_483_0, i_8_248_484_0, i_8_248_529_0,
    i_8_248_587_0, i_8_248_588_0, i_8_248_601_0, i_8_248_628_0,
    i_8_248_653_0, i_8_248_661_0, i_8_248_669_0, i_8_248_680_0,
    i_8_248_691_0, i_8_248_707_0, i_8_248_747_0, i_8_248_748_0,
    i_8_248_786_0, i_8_248_789_0, i_8_248_823_0, i_8_248_839_0,
    i_8_248_842_0, i_8_248_844_0, i_8_248_845_0, i_8_248_868_0,
    i_8_248_894_0, i_8_248_993_0, i_8_248_994_0, i_8_248_996_0,
    i_8_248_1039_0, i_8_248_1050_0, i_8_248_1074_0, i_8_248_1075_0,
    i_8_248_1110_0, i_8_248_1112_0, i_8_248_1202_0, i_8_248_1227_0,
    i_8_248_1270_0, i_8_248_1274_0, i_8_248_1278_0, i_8_248_1282_0,
    i_8_248_1300_0, i_8_248_1307_0, i_8_248_1308_0, i_8_248_1359_0,
    i_8_248_1456_0, i_8_248_1462_0, i_8_248_1474_0, i_8_248_1507_0,
    i_8_248_1511_0, i_8_248_1516_0, i_8_248_1525_0, i_8_248_1540_0,
    i_8_248_1558_0, i_8_248_1561_0, i_8_248_1572_0, i_8_248_1633_0,
    i_8_248_1720_0, i_8_248_1726_0, i_8_248_1740_0, i_8_248_1749_0,
    i_8_248_1753_0, i_8_248_1775_0, i_8_248_1783_0, i_8_248_1796_0,
    i_8_248_1810_0, i_8_248_1828_0, i_8_248_1876_0, i_8_248_1906_0,
    i_8_248_1969_0, i_8_248_1991_0, i_8_248_2031_0, i_8_248_2136_0,
    i_8_248_2154_0, i_8_248_2191_0, i_8_248_2214_0, i_8_248_2218_0,
    i_8_248_2236_0, i_8_248_2243_0, i_8_248_2293_0,
    o_8_248_0_0  );
  input  i_8_248_31_0, i_8_248_39_0, i_8_248_42_0, i_8_248_51_0,
    i_8_248_55_0, i_8_248_96_0, i_8_248_97_0, i_8_248_169_0, i_8_248_256_0,
    i_8_248_258_0, i_8_248_300_0, i_8_248_307_0, i_8_248_319_0,
    i_8_248_331_0, i_8_248_334_0, i_8_248_360_0, i_8_248_363_0,
    i_8_248_417_0, i_8_248_418_0, i_8_248_421_0, i_8_248_440_0,
    i_8_248_481_0, i_8_248_483_0, i_8_248_484_0, i_8_248_529_0,
    i_8_248_587_0, i_8_248_588_0, i_8_248_601_0, i_8_248_628_0,
    i_8_248_653_0, i_8_248_661_0, i_8_248_669_0, i_8_248_680_0,
    i_8_248_691_0, i_8_248_707_0, i_8_248_747_0, i_8_248_748_0,
    i_8_248_786_0, i_8_248_789_0, i_8_248_823_0, i_8_248_839_0,
    i_8_248_842_0, i_8_248_844_0, i_8_248_845_0, i_8_248_868_0,
    i_8_248_894_0, i_8_248_993_0, i_8_248_994_0, i_8_248_996_0,
    i_8_248_1039_0, i_8_248_1050_0, i_8_248_1074_0, i_8_248_1075_0,
    i_8_248_1110_0, i_8_248_1112_0, i_8_248_1202_0, i_8_248_1227_0,
    i_8_248_1270_0, i_8_248_1274_0, i_8_248_1278_0, i_8_248_1282_0,
    i_8_248_1300_0, i_8_248_1307_0, i_8_248_1308_0, i_8_248_1359_0,
    i_8_248_1456_0, i_8_248_1462_0, i_8_248_1474_0, i_8_248_1507_0,
    i_8_248_1511_0, i_8_248_1516_0, i_8_248_1525_0, i_8_248_1540_0,
    i_8_248_1558_0, i_8_248_1561_0, i_8_248_1572_0, i_8_248_1633_0,
    i_8_248_1720_0, i_8_248_1726_0, i_8_248_1740_0, i_8_248_1749_0,
    i_8_248_1753_0, i_8_248_1775_0, i_8_248_1783_0, i_8_248_1796_0,
    i_8_248_1810_0, i_8_248_1828_0, i_8_248_1876_0, i_8_248_1906_0,
    i_8_248_1969_0, i_8_248_1991_0, i_8_248_2031_0, i_8_248_2136_0,
    i_8_248_2154_0, i_8_248_2191_0, i_8_248_2214_0, i_8_248_2218_0,
    i_8_248_2236_0, i_8_248_2243_0, i_8_248_2293_0;
  output o_8_248_0_0;
  assign o_8_248_0_0 = 0;
endmodule



// Benchmark "kernel_8_249" written by ABC on Sun Jul 19 10:07:25 2020

module kernel_8_249 ( 
    i_8_249_35_0, i_8_249_48_0, i_8_249_49_0, i_8_249_50_0, i_8_249_51_0,
    i_8_249_52_0, i_8_249_53_0, i_8_249_58_0, i_8_249_97_0, i_8_249_163_0,
    i_8_249_164_0, i_8_249_167_0, i_8_249_185_0, i_8_249_188_0,
    i_8_249_217_0, i_8_249_292_0, i_8_249_349_0, i_8_249_450_0,
    i_8_249_552_0, i_8_249_554_0, i_8_249_555_0, i_8_249_556_0,
    i_8_249_557_0, i_8_249_578_0, i_8_249_581_0, i_8_249_603_0,
    i_8_249_606_0, i_8_249_637_0, i_8_249_648_0, i_8_249_652_0,
    i_8_249_684_0, i_8_249_703_0, i_8_249_704_0, i_8_249_747_0,
    i_8_249_780_0, i_8_249_860_0, i_8_249_927_0, i_8_249_930_0,
    i_8_249_931_0, i_8_249_932_0, i_8_249_956_0, i_8_249_964_0,
    i_8_249_968_0, i_8_249_1050_0, i_8_249_1109_0, i_8_249_1110_0,
    i_8_249_1111_0, i_8_249_1112_0, i_8_249_1113_0, i_8_249_1114_0,
    i_8_249_1115_0, i_8_249_1125_0, i_8_249_1129_0, i_8_249_1256_0,
    i_8_249_1269_0, i_8_249_1270_0, i_8_249_1271_0, i_8_249_1335_0,
    i_8_249_1343_0, i_8_249_1388_0, i_8_249_1409_0, i_8_249_1437_0,
    i_8_249_1457_0, i_8_249_1533_0, i_8_249_1563_0, i_8_249_1564_0,
    i_8_249_1570_0, i_8_249_1651_0, i_8_249_1676_0, i_8_249_1678_0,
    i_8_249_1679_0, i_8_249_1682_0, i_8_249_1763_0, i_8_249_1773_0,
    i_8_249_1774_0, i_8_249_1775_0, i_8_249_1778_0, i_8_249_1819_0,
    i_8_249_1820_0, i_8_249_1917_0, i_8_249_1918_0, i_8_249_1947_0,
    i_8_249_1963_0, i_8_249_1964_0, i_8_249_1985_0, i_8_249_2004_0,
    i_8_249_2016_0, i_8_249_2046_0, i_8_249_2047_0, i_8_249_2049_0,
    i_8_249_2116_0, i_8_249_2153_0, i_8_249_2169_0, i_8_249_2171_0,
    i_8_249_2172_0, i_8_249_2173_0, i_8_249_2174_0, i_8_249_2247_0,
    i_8_249_2261_0, i_8_249_2291_0,
    o_8_249_0_0  );
  input  i_8_249_35_0, i_8_249_48_0, i_8_249_49_0, i_8_249_50_0,
    i_8_249_51_0, i_8_249_52_0, i_8_249_53_0, i_8_249_58_0, i_8_249_97_0,
    i_8_249_163_0, i_8_249_164_0, i_8_249_167_0, i_8_249_185_0,
    i_8_249_188_0, i_8_249_217_0, i_8_249_292_0, i_8_249_349_0,
    i_8_249_450_0, i_8_249_552_0, i_8_249_554_0, i_8_249_555_0,
    i_8_249_556_0, i_8_249_557_0, i_8_249_578_0, i_8_249_581_0,
    i_8_249_603_0, i_8_249_606_0, i_8_249_637_0, i_8_249_648_0,
    i_8_249_652_0, i_8_249_684_0, i_8_249_703_0, i_8_249_704_0,
    i_8_249_747_0, i_8_249_780_0, i_8_249_860_0, i_8_249_927_0,
    i_8_249_930_0, i_8_249_931_0, i_8_249_932_0, i_8_249_956_0,
    i_8_249_964_0, i_8_249_968_0, i_8_249_1050_0, i_8_249_1109_0,
    i_8_249_1110_0, i_8_249_1111_0, i_8_249_1112_0, i_8_249_1113_0,
    i_8_249_1114_0, i_8_249_1115_0, i_8_249_1125_0, i_8_249_1129_0,
    i_8_249_1256_0, i_8_249_1269_0, i_8_249_1270_0, i_8_249_1271_0,
    i_8_249_1335_0, i_8_249_1343_0, i_8_249_1388_0, i_8_249_1409_0,
    i_8_249_1437_0, i_8_249_1457_0, i_8_249_1533_0, i_8_249_1563_0,
    i_8_249_1564_0, i_8_249_1570_0, i_8_249_1651_0, i_8_249_1676_0,
    i_8_249_1678_0, i_8_249_1679_0, i_8_249_1682_0, i_8_249_1763_0,
    i_8_249_1773_0, i_8_249_1774_0, i_8_249_1775_0, i_8_249_1778_0,
    i_8_249_1819_0, i_8_249_1820_0, i_8_249_1917_0, i_8_249_1918_0,
    i_8_249_1947_0, i_8_249_1963_0, i_8_249_1964_0, i_8_249_1985_0,
    i_8_249_2004_0, i_8_249_2016_0, i_8_249_2046_0, i_8_249_2047_0,
    i_8_249_2049_0, i_8_249_2116_0, i_8_249_2153_0, i_8_249_2169_0,
    i_8_249_2171_0, i_8_249_2172_0, i_8_249_2173_0, i_8_249_2174_0,
    i_8_249_2247_0, i_8_249_2261_0, i_8_249_2291_0;
  output o_8_249_0_0;
  assign o_8_249_0_0 = ~((i_8_249_217_0 & ((~i_8_249_53_0 & ~i_8_249_684_0 & ~i_8_249_964_0 & ~i_8_249_968_0 & ~i_8_249_1437_0 & ~i_8_249_1679_0 & i_8_249_1917_0) | (i_8_249_58_0 & i_8_249_1109_0 & i_8_249_2291_0))) | (~i_8_249_217_0 & ((~i_8_249_167_0 & ~i_8_249_185_0 & ~i_8_249_581_0 & ~i_8_249_1270_0 & ~i_8_249_1343_0 & i_8_249_1819_0 & i_8_249_1985_0 & ~i_8_249_2171_0) | (~i_8_249_49_0 & i_8_249_349_0 & ~i_8_249_557_0 & i_8_249_1115_0 & ~i_8_249_1409_0 & ~i_8_249_1963_0 & ~i_8_249_2173_0))) | (~i_8_249_185_0 & ((~i_8_249_450_0 & i_8_249_606_0 & ~i_8_249_930_0 & ~i_8_249_1110_0 & i_8_249_1335_0 & ~i_8_249_1564_0) | (~i_8_249_964_0 & ~i_8_249_1271_0 & ~i_8_249_1682_0 & ~i_8_249_2116_0 & i_8_249_2171_0 & ~i_8_249_2291_0))) | (~i_8_249_1050_0 & ((~i_8_249_48_0 & ((~i_8_249_49_0 & ~i_8_249_51_0 & i_8_249_349_0 & ~i_8_249_450_0 & i_8_249_1113_0 & ~i_8_249_1256_0 & ~i_8_249_2173_0) | (~i_8_249_188_0 & i_8_249_557_0 & i_8_249_1115_0 & ~i_8_249_1564_0 & ~i_8_249_1947_0 & ~i_8_249_2261_0))) | (~i_8_249_52_0 & ~i_8_249_1682_0 & ((~i_8_249_53_0 & ~i_8_249_349_0 & i_8_249_1114_0 & ~i_8_249_1256_0 & ~i_8_249_1437_0 & ~i_8_249_1651_0 & ~i_8_249_1918_0) | (~i_8_249_552_0 & ~i_8_249_684_0 & i_8_249_780_0 & i_8_249_1437_0 & ~i_8_249_1678_0 & ~i_8_249_1947_0))) | (~i_8_249_2004_0 & ((~i_8_249_450_0 & ((~i_8_249_49_0 & i_8_249_1110_0 & ~i_8_249_1114_0 & ~i_8_249_1269_0 & ~i_8_249_1409_0 & ~i_8_249_1437_0 & ~i_8_249_1963_0) | (i_8_249_552_0 & i_8_249_1533_0 & ~i_8_249_2261_0))) | (~i_8_249_50_0 & i_8_249_556_0 & ~i_8_249_1113_0 & ~i_8_249_1256_0 & ~i_8_249_1335_0 & ~i_8_249_1457_0 & ~i_8_249_1570_0 & ~i_8_249_1678_0 & ~i_8_249_2247_0 & ~i_8_249_2291_0))) | (~i_8_249_58_0 & i_8_249_349_0 & ~i_8_249_930_0 & i_8_249_1335_0 & ~i_8_249_1563_0 & ~i_8_249_1651_0 & ~i_8_249_1985_0))) | (~i_8_249_164_0 & ((~i_8_249_50_0 & ~i_8_249_2153_0 & ((~i_8_249_97_0 & ~i_8_249_167_0 & ~i_8_249_450_0 & ~i_8_249_1270_0 & ~i_8_249_1437_0 & i_8_249_1679_0 & i_8_249_1778_0 & ~i_8_249_1963_0) | (~i_8_249_58_0 & ~i_8_249_188_0 & ~i_8_249_603_0 & i_8_249_1111_0 & ~i_8_249_1335_0 & i_8_249_1651_0 & ~i_8_249_1678_0 & ~i_8_249_2004_0 & ~i_8_249_2173_0))) | (~i_8_249_2016_0 & ((~i_8_249_58_0 & ~i_8_249_968_0 & i_8_249_1109_0 & i_8_249_1778_0) | (~i_8_249_49_0 & ~i_8_249_53_0 & ~i_8_249_603_0 & ~i_8_249_606_0 & ~i_8_249_1111_0 & ~i_8_249_1343_0 & ~i_8_249_1409_0 & ~i_8_249_1533_0 & i_8_249_1819_0 & i_8_249_1918_0 & ~i_8_249_2004_0) | (~i_8_249_52_0 & ~i_8_249_163_0 & ~i_8_249_450_0 & ~i_8_249_780_0 & ~i_8_249_964_0 & i_8_249_1676_0 & ~i_8_249_1820_0 & i_8_249_2153_0))) | (~i_8_249_578_0 & i_8_249_704_0 & ~i_8_249_1256_0 & i_8_249_2171_0 & ~i_8_249_2172_0 & ~i_8_249_2291_0))) | (~i_8_249_349_0 & ((i_8_249_552_0 & ((~i_8_249_931_0 & i_8_249_1113_0 & ~i_8_249_1682_0 & ~i_8_249_2016_0) | (~i_8_249_52_0 & ~i_8_249_450_0 & i_8_249_637_0 & ~i_8_249_684_0 & ~i_8_249_968_0 & ~i_8_249_1409_0 & ~i_8_249_2047_0))) | (~i_8_249_780_0 & ~i_8_249_932_0 & i_8_249_1774_0 & i_8_249_1820_0))) | (~i_8_249_637_0 & ((i_8_249_35_0 & ~i_8_249_50_0 & ~i_8_249_52_0 & ~i_8_249_167_0 & ~i_8_249_860_0 & ~i_8_249_1112_0 & ~i_8_249_1409_0 & ~i_8_249_1778_0) | (~i_8_249_48_0 & i_8_249_1125_0 & ~i_8_249_1563_0 & i_8_249_1918_0 & ~i_8_249_1947_0))) | (~i_8_249_48_0 & ((~i_8_249_50_0 & ((i_8_249_53_0 & i_8_249_1115_0 & ~i_8_249_1270_0 & ~i_8_249_1457_0 & ~i_8_249_1820_0) | (~i_8_249_53_0 & ~i_8_249_578_0 & i_8_249_1775_0 & ~i_8_249_2116_0))) | (~i_8_249_53_0 & i_8_249_637_0 & ~i_8_249_932_0 & i_8_249_1115_0 & ~i_8_249_1256_0 & ~i_8_249_1651_0) | (i_8_249_606_0 & ~i_8_249_684_0 & i_8_249_1773_0) | (~i_8_249_51_0 & ~i_8_249_652_0 & i_8_249_780_0 & i_8_249_1563_0 & ~i_8_249_1918_0) | (~i_8_249_52_0 & ~i_8_249_97_0 & i_8_249_1113_0 & i_8_249_1114_0 & ~i_8_249_2291_0))) | (i_8_249_1679_0 & ((~i_8_249_167_0 & ((~i_8_249_163_0 & i_8_249_1112_0 & ~i_8_249_1388_0 & i_8_249_1918_0 & i_8_249_1985_0) | (~i_8_249_52_0 & ~i_8_249_964_0 & i_8_249_1115_0 & ~i_8_249_2116_0))) | (~i_8_249_163_0 & ((~i_8_249_1271_0 & ~i_8_249_1409_0 & i_8_249_1533_0 & ~i_8_249_1775_0 & i_8_249_1778_0) | (~i_8_249_97_0 & i_8_249_1115_0 & i_8_249_1963_0))) | (~i_8_249_930_0 & ~i_8_249_932_0 & i_8_249_1113_0 & ~i_8_249_1388_0) | (~i_8_249_49_0 & ~i_8_249_51_0 & i_8_249_1343_0 & ~i_8_249_2153_0))) | (~i_8_249_52_0 & ((~i_8_249_930_0 & i_8_249_968_0 & i_8_249_1112_0 & i_8_249_1115_0 & ~i_8_249_1256_0) | (~i_8_249_450_0 & i_8_249_648_0 & i_8_249_747_0 & ~i_8_249_1343_0))) | (~i_8_249_97_0 & ((~i_8_249_188_0 & i_8_249_603_0 & i_8_249_1125_0) | (i_8_249_557_0 & i_8_249_1115_0 & ~i_8_249_1335_0 & ~i_8_249_1564_0 & ~i_8_249_1682_0 & ~i_8_249_1963_0 & ~i_8_249_2153_0))) | (i_8_249_557_0 & ((~i_8_249_53_0 & ~i_8_249_554_0 & ~i_8_249_930_0 & i_8_249_1437_0 & ~i_8_249_2049_0) | (i_8_249_1114_0 & i_8_249_1115_0 & ~i_8_249_1570_0 & ~i_8_249_2261_0))) | (i_8_249_606_0 & ((~i_8_249_49_0 & ~i_8_249_163_0 & ~i_8_249_450_0 & ~i_8_249_684_0 & ~i_8_249_964_0 & ~i_8_249_968_0 & ~i_8_249_1269_0 & ~i_8_249_1563_0 & ~i_8_249_1682_0 & ~i_8_249_1774_0 & ~i_8_249_1819_0 & ~i_8_249_2169_0) | (i_8_249_1774_0 & i_8_249_2172_0))) | (i_8_249_747_0 & ((i_8_249_648_0 & i_8_249_1773_0) | (~i_8_249_964_0 & i_8_249_1678_0 & i_8_249_1918_0))) | (i_8_249_648_0 & ((~i_8_249_450_0 & i_8_249_1773_0) | (~i_8_249_1269_0 & ~i_8_249_1437_0 & i_8_249_1678_0 & ~i_8_249_1819_0 & i_8_249_1918_0))) | (~i_8_249_450_0 & ((~i_8_249_684_0 & i_8_249_1774_0 & ~i_8_249_1947_0 & i_8_249_2169_0) | (~i_8_249_552_0 & i_8_249_556_0 & ~i_8_249_1111_0 & i_8_249_1113_0 & i_8_249_1437_0 & i_8_249_1678_0 & ~i_8_249_2004_0 & ~i_8_249_2049_0 & ~i_8_249_2172_0))) | (~i_8_249_51_0 & ((~i_8_249_188_0 & ((i_8_249_1110_0 & i_8_249_1112_0 & ~i_8_249_1570_0 & i_8_249_1651_0) | (i_8_249_1113_0 & i_8_249_2049_0 & ~i_8_249_2174_0))) | (i_8_249_556_0 & ((~i_8_249_1114_0 & i_8_249_1335_0 & i_8_249_1437_0) | (i_8_249_555_0 & i_8_249_2049_0))) | (~i_8_249_49_0 & ~i_8_249_964_0 & i_8_249_1112_0 & i_8_249_1437_0 & ~i_8_249_1564_0 & ~i_8_249_2153_0))) | (~i_8_249_49_0 & i_8_249_2174_0 & ((~i_8_249_53_0 & ~i_8_249_188_0 & ~i_8_249_704_0 & ~i_8_249_1271_0 & ~i_8_249_1679_0) | (~i_8_249_964_0 & i_8_249_1115_0 & ~i_8_249_1570_0 & ~i_8_249_1947_0))) | (~i_8_249_53_0 & i_8_249_1682_0 & ((~i_8_249_930_0 & ~i_8_249_956_0 & ~i_8_249_968_0 & ~i_8_249_1113_0 & ~i_8_249_1269_0 & ~i_8_249_1271_0 & ~i_8_249_1343_0 & i_8_249_1918_0 & ~i_8_249_1963_0) | (i_8_249_780_0 & ~i_8_249_964_0 & ~i_8_249_1651_0 & ~i_8_249_1679_0 & ~i_8_249_2174_0 & ~i_8_249_2261_0))) | (i_8_249_1110_0 & ((~i_8_249_747_0 & ~i_8_249_1457_0 & i_8_249_1773_0) | (i_8_249_1113_0 & i_8_249_1437_0 & i_8_249_1917_0))) | (~i_8_249_2116_0 & ((i_8_249_652_0 & i_8_249_780_0 & ~i_8_249_956_0 & i_8_249_1111_0) | (~i_8_249_1256_0 & ~i_8_249_1533_0 & i_8_249_1775_0 & i_8_249_1819_0 & ~i_8_249_2016_0))) | (i_8_249_1774_0 & ~i_8_249_2172_0 & i_8_249_2173_0) | (i_8_249_1050_0 & i_8_249_1113_0 & ~i_8_249_1269_0 & ~i_8_249_1335_0 & i_8_249_1533_0 & ~i_8_249_2291_0));
endmodule



// Benchmark "kernel_8_250" written by ABC on Sun Jul 19 10:07:26 2020

module kernel_8_250 ( 
    i_8_250_3_0, i_8_250_12_0, i_8_250_18_0, i_8_250_21_0, i_8_250_22_0,
    i_8_250_52_0, i_8_250_66_0, i_8_250_75_0, i_8_250_114_0, i_8_250_147_0,
    i_8_250_192_0, i_8_250_202_0, i_8_250_226_0, i_8_250_273_0,
    i_8_250_274_0, i_8_250_276_0, i_8_250_321_0, i_8_250_354_0,
    i_8_250_375_0, i_8_250_400_0, i_8_250_516_0, i_8_250_526_0,
    i_8_250_574_0, i_8_250_579_0, i_8_250_590_0, i_8_250_598_0,
    i_8_250_616_0, i_8_250_619_0, i_8_250_633_0, i_8_250_643_0,
    i_8_250_649_0, i_8_250_651_0, i_8_250_693_0, i_8_250_696_0,
    i_8_250_701_0, i_8_250_703_0, i_8_250_732_0, i_8_250_780_0,
    i_8_250_831_0, i_8_250_841_0, i_8_250_858_0, i_8_250_861_0,
    i_8_250_977_0, i_8_250_1200_0, i_8_250_1228_0, i_8_250_1236_0,
    i_8_250_1237_0, i_8_250_1270_0, i_8_250_1296_0, i_8_250_1302_0,
    i_8_250_1317_0, i_8_250_1318_0, i_8_250_1323_0, i_8_250_1350_0,
    i_8_250_1353_0, i_8_250_1356_0, i_8_250_1389_0, i_8_250_1398_0,
    i_8_250_1408_0, i_8_250_1410_0, i_8_250_1423_0, i_8_250_1436_0,
    i_8_250_1488_0, i_8_250_1497_0, i_8_250_1505_0, i_8_250_1516_0,
    i_8_250_1534_0, i_8_250_1551_0, i_8_250_1569_0, i_8_250_1573_0,
    i_8_250_1639_0, i_8_250_1647_0, i_8_250_1659_0, i_8_250_1677_0,
    i_8_250_1701_0, i_8_250_1746_0, i_8_250_1753_0, i_8_250_1782_0,
    i_8_250_1813_0, i_8_250_1824_0, i_8_250_1839_0, i_8_250_1843_0,
    i_8_250_1866_0, i_8_250_1881_0, i_8_250_1884_0, i_8_250_1911_0,
    i_8_250_1917_0, i_8_250_1939_0, i_8_250_1944_0, i_8_250_1992_0,
    i_8_250_1993_0, i_8_250_2008_0, i_8_250_2010_0, i_8_250_2013_0,
    i_8_250_2046_0, i_8_250_2062_0, i_8_250_2064_0, i_8_250_2184_0,
    i_8_250_2215_0, i_8_250_2248_0,
    o_8_250_0_0  );
  input  i_8_250_3_0, i_8_250_12_0, i_8_250_18_0, i_8_250_21_0,
    i_8_250_22_0, i_8_250_52_0, i_8_250_66_0, i_8_250_75_0, i_8_250_114_0,
    i_8_250_147_0, i_8_250_192_0, i_8_250_202_0, i_8_250_226_0,
    i_8_250_273_0, i_8_250_274_0, i_8_250_276_0, i_8_250_321_0,
    i_8_250_354_0, i_8_250_375_0, i_8_250_400_0, i_8_250_516_0,
    i_8_250_526_0, i_8_250_574_0, i_8_250_579_0, i_8_250_590_0,
    i_8_250_598_0, i_8_250_616_0, i_8_250_619_0, i_8_250_633_0,
    i_8_250_643_0, i_8_250_649_0, i_8_250_651_0, i_8_250_693_0,
    i_8_250_696_0, i_8_250_701_0, i_8_250_703_0, i_8_250_732_0,
    i_8_250_780_0, i_8_250_831_0, i_8_250_841_0, i_8_250_858_0,
    i_8_250_861_0, i_8_250_977_0, i_8_250_1200_0, i_8_250_1228_0,
    i_8_250_1236_0, i_8_250_1237_0, i_8_250_1270_0, i_8_250_1296_0,
    i_8_250_1302_0, i_8_250_1317_0, i_8_250_1318_0, i_8_250_1323_0,
    i_8_250_1350_0, i_8_250_1353_0, i_8_250_1356_0, i_8_250_1389_0,
    i_8_250_1398_0, i_8_250_1408_0, i_8_250_1410_0, i_8_250_1423_0,
    i_8_250_1436_0, i_8_250_1488_0, i_8_250_1497_0, i_8_250_1505_0,
    i_8_250_1516_0, i_8_250_1534_0, i_8_250_1551_0, i_8_250_1569_0,
    i_8_250_1573_0, i_8_250_1639_0, i_8_250_1647_0, i_8_250_1659_0,
    i_8_250_1677_0, i_8_250_1701_0, i_8_250_1746_0, i_8_250_1753_0,
    i_8_250_1782_0, i_8_250_1813_0, i_8_250_1824_0, i_8_250_1839_0,
    i_8_250_1843_0, i_8_250_1866_0, i_8_250_1881_0, i_8_250_1884_0,
    i_8_250_1911_0, i_8_250_1917_0, i_8_250_1939_0, i_8_250_1944_0,
    i_8_250_1992_0, i_8_250_1993_0, i_8_250_2008_0, i_8_250_2010_0,
    i_8_250_2013_0, i_8_250_2046_0, i_8_250_2062_0, i_8_250_2064_0,
    i_8_250_2184_0, i_8_250_2215_0, i_8_250_2248_0;
  output o_8_250_0_0;
  assign o_8_250_0_0 = ~((~i_8_250_202_0 & ((~i_8_250_354_0 & ~i_8_250_696_0 & i_8_250_1753_0) | (~i_8_250_274_0 & ~i_8_250_598_0 & ~i_8_250_619_0 & ~i_8_250_732_0 & ~i_8_250_1389_0 & ~i_8_250_1659_0 & ~i_8_250_1843_0 & ~i_8_250_2184_0))) | (~i_8_250_276_0 & ((i_8_250_114_0 & ~i_8_250_321_0 & i_8_250_703_0 & ~i_8_250_1551_0 & ~i_8_250_1843_0 & i_8_250_1884_0) | (~i_8_250_590_0 & ~i_8_250_649_0 & ~i_8_250_841_0 & ~i_8_250_1200_0 & ~i_8_250_1296_0 & ~i_8_250_1497_0 & ~i_8_250_1813_0 & ~i_8_250_1911_0 & ~i_8_250_1993_0 & ~i_8_250_2010_0))) | (~i_8_250_354_0 & ((~i_8_250_3_0 & ~i_8_250_858_0 & ~i_8_250_1398_0 & i_8_250_1881_0) | (~i_8_250_579_0 & ~i_8_250_590_0 & ~i_8_250_651_0 & ~i_8_250_831_0 & ~i_8_250_1534_0 & ~i_8_250_1569_0 & ~i_8_250_1911_0 & ~i_8_250_2008_0))) | (~i_8_250_3_0 & ((~i_8_250_18_0 & ~i_8_250_52_0 & i_8_250_192_0 & ~i_8_250_274_0 & ~i_8_250_643_0 & ~i_8_250_1436_0 & ~i_8_250_1866_0) | (~i_8_250_732_0 & ~i_8_250_1317_0 & ~i_8_250_1389_0 & ~i_8_250_1839_0 & ~i_8_250_2046_0 & ~i_8_250_2064_0))) | (~i_8_250_274_0 & ((~i_8_250_12_0 & i_8_250_598_0 & ~i_8_250_831_0 & ~i_8_250_1881_0 & ~i_8_250_1911_0) | (~i_8_250_21_0 & ~i_8_250_273_0 & ~i_8_250_616_0 & ~i_8_250_1408_0 & ~i_8_250_1569_0 & ~i_8_250_1639_0 & ~i_8_250_1659_0 & ~i_8_250_1813_0 & ~i_8_250_2008_0 & ~i_8_250_2062_0))) | (~i_8_250_21_0 & ((~i_8_250_590_0 & ~i_8_250_651_0 & i_8_250_1639_0 & ~i_8_250_2010_0) | (~i_8_250_18_0 & ~i_8_250_52_0 & ~i_8_250_400_0 & ~i_8_250_579_0 & ~i_8_250_1270_0 & i_8_250_1488_0 & ~i_8_250_1573_0 & ~i_8_250_1659_0 & ~i_8_250_1866_0 & ~i_8_250_2062_0))) | (~i_8_250_18_0 & ((~i_8_250_732_0 & ~i_8_250_1228_0 & ~i_8_250_1497_0 & ~i_8_250_1866_0) | (~i_8_250_400_0 & ~i_8_250_633_0 & ~i_8_250_696_0 & ~i_8_250_1782_0 & ~i_8_250_1911_0 & ~i_8_250_2064_0))) | (~i_8_250_52_0 & ((~i_8_250_226_0 & ~i_8_250_579_0 & ~i_8_250_1497_0 & ~i_8_250_1534_0 & i_8_250_2046_0 & ~i_8_250_2064_0) | (~i_8_250_147_0 & ~i_8_250_780_0 & i_8_250_1296_0 & ~i_8_250_1389_0 & i_8_250_1647_0 & ~i_8_250_1911_0 & ~i_8_250_2215_0))) | (~i_8_250_273_0 & ((~i_8_250_516_0 & ~i_8_250_598_0 & ~i_8_250_831_0 & ~i_8_250_1423_0 & ~i_8_250_1505_0 & ~i_8_250_2062_0 & ~i_8_250_2064_0) | (i_8_250_1677_0 & i_8_250_1839_0 & ~i_8_250_2215_0))) | (~i_8_250_516_0 & ((~i_8_250_192_0 & i_8_250_693_0 & i_8_250_1353_0 & ~i_8_250_1389_0 & ~i_8_250_1408_0 & ~i_8_250_1505_0) | (~i_8_250_75_0 & ~i_8_250_590_0 & ~i_8_250_1236_0 & i_8_250_1551_0 & ~i_8_250_1659_0 & ~i_8_250_1993_0))) | (~i_8_250_1866_0 & ((~i_8_250_75_0 & ~i_8_250_1236_0 & ~i_8_250_1497_0 & ~i_8_250_1505_0 & i_8_250_1677_0 & ~i_8_250_1992_0 & ~i_8_250_2046_0) | (i_8_250_1237_0 & ~i_8_250_1323_0 & ~i_8_250_1350_0 & ~i_8_250_1389_0 & i_8_250_1824_0 & ~i_8_250_2064_0))) | (~i_8_250_75_0 & ((i_8_250_274_0 & ~i_8_250_1423_0 & ~i_8_250_1782_0 & ~i_8_250_2010_0) | (~i_8_250_22_0 & ~i_8_250_66_0 & ~i_8_250_616_0 & ~i_8_250_2064_0))));
endmodule



// Benchmark "kernel_8_251" written by ABC on Sun Jul 19 10:07:27 2020

module kernel_8_251 ( 
    i_8_251_28_0, i_8_251_67_0, i_8_251_72_0, i_8_251_140_0, i_8_251_143_0,
    i_8_251_201_0, i_8_251_258_0, i_8_251_259_0, i_8_251_275_0,
    i_8_251_385_0, i_8_251_392_0, i_8_251_401_0, i_8_251_429_0,
    i_8_251_457_0, i_8_251_492_0, i_8_251_498_0, i_8_251_499_0,
    i_8_251_522_0, i_8_251_550_0, i_8_251_556_0, i_8_251_630_0,
    i_8_251_632_0, i_8_251_655_0, i_8_251_659_0, i_8_251_662_0,
    i_8_251_672_0, i_8_251_673_0, i_8_251_695_0, i_8_251_820_0,
    i_8_251_843_0, i_8_251_854_0, i_8_251_859_0, i_8_251_880_0,
    i_8_251_881_0, i_8_251_916_0, i_8_251_959_0, i_8_251_995_0,
    i_8_251_1075_0, i_8_251_1084_0, i_8_251_1087_0, i_8_251_1106_0,
    i_8_251_1108_0, i_8_251_1109_0, i_8_251_1113_0, i_8_251_1174_0,
    i_8_251_1201_0, i_8_251_1230_0, i_8_251_1238_0, i_8_251_1267_0,
    i_8_251_1273_0, i_8_251_1322_0, i_8_251_1330_0, i_8_251_1331_0,
    i_8_251_1333_0, i_8_251_1411_0, i_8_251_1426_0, i_8_251_1433_0,
    i_8_251_1471_0, i_8_251_1480_0, i_8_251_1484_0, i_8_251_1498_0,
    i_8_251_1528_0, i_8_251_1547_0, i_8_251_1561_0, i_8_251_1573_0,
    i_8_251_1598_0, i_8_251_1641_0, i_8_251_1653_0, i_8_251_1659_0,
    i_8_251_1705_0, i_8_251_1732_0, i_8_251_1748_0, i_8_251_1750_0,
    i_8_251_1753_0, i_8_251_1754_0, i_8_251_1762_0, i_8_251_1774_0,
    i_8_251_1816_0, i_8_251_1849_0, i_8_251_1852_0, i_8_251_1865_0,
    i_8_251_1867_0, i_8_251_1876_0, i_8_251_1882_0, i_8_251_1889_0,
    i_8_251_1895_0, i_8_251_1912_0, i_8_251_1921_0, i_8_251_1952_0,
    i_8_251_1966_0, i_8_251_1975_0, i_8_251_2048_0, i_8_251_2066_0,
    i_8_251_2092_0, i_8_251_2093_0, i_8_251_2119_0, i_8_251_2150_0,
    i_8_251_2229_0, i_8_251_2230_0, i_8_251_2299_0,
    o_8_251_0_0  );
  input  i_8_251_28_0, i_8_251_67_0, i_8_251_72_0, i_8_251_140_0,
    i_8_251_143_0, i_8_251_201_0, i_8_251_258_0, i_8_251_259_0,
    i_8_251_275_0, i_8_251_385_0, i_8_251_392_0, i_8_251_401_0,
    i_8_251_429_0, i_8_251_457_0, i_8_251_492_0, i_8_251_498_0,
    i_8_251_499_0, i_8_251_522_0, i_8_251_550_0, i_8_251_556_0,
    i_8_251_630_0, i_8_251_632_0, i_8_251_655_0, i_8_251_659_0,
    i_8_251_662_0, i_8_251_672_0, i_8_251_673_0, i_8_251_695_0,
    i_8_251_820_0, i_8_251_843_0, i_8_251_854_0, i_8_251_859_0,
    i_8_251_880_0, i_8_251_881_0, i_8_251_916_0, i_8_251_959_0,
    i_8_251_995_0, i_8_251_1075_0, i_8_251_1084_0, i_8_251_1087_0,
    i_8_251_1106_0, i_8_251_1108_0, i_8_251_1109_0, i_8_251_1113_0,
    i_8_251_1174_0, i_8_251_1201_0, i_8_251_1230_0, i_8_251_1238_0,
    i_8_251_1267_0, i_8_251_1273_0, i_8_251_1322_0, i_8_251_1330_0,
    i_8_251_1331_0, i_8_251_1333_0, i_8_251_1411_0, i_8_251_1426_0,
    i_8_251_1433_0, i_8_251_1471_0, i_8_251_1480_0, i_8_251_1484_0,
    i_8_251_1498_0, i_8_251_1528_0, i_8_251_1547_0, i_8_251_1561_0,
    i_8_251_1573_0, i_8_251_1598_0, i_8_251_1641_0, i_8_251_1653_0,
    i_8_251_1659_0, i_8_251_1705_0, i_8_251_1732_0, i_8_251_1748_0,
    i_8_251_1750_0, i_8_251_1753_0, i_8_251_1754_0, i_8_251_1762_0,
    i_8_251_1774_0, i_8_251_1816_0, i_8_251_1849_0, i_8_251_1852_0,
    i_8_251_1865_0, i_8_251_1867_0, i_8_251_1876_0, i_8_251_1882_0,
    i_8_251_1889_0, i_8_251_1895_0, i_8_251_1912_0, i_8_251_1921_0,
    i_8_251_1952_0, i_8_251_1966_0, i_8_251_1975_0, i_8_251_2048_0,
    i_8_251_2066_0, i_8_251_2092_0, i_8_251_2093_0, i_8_251_2119_0,
    i_8_251_2150_0, i_8_251_2229_0, i_8_251_2230_0, i_8_251_2299_0;
  output o_8_251_0_0;
  assign o_8_251_0_0 = 0;
endmodule



// Benchmark "kernel_8_252" written by ABC on Sun Jul 19 10:07:28 2020

module kernel_8_252 ( 
    i_8_252_3_0, i_8_252_8_0, i_8_252_22_0, i_8_252_50_0, i_8_252_78_0,
    i_8_252_80_0, i_8_252_114_0, i_8_252_125_0, i_8_252_177_0,
    i_8_252_185_0, i_8_252_192_0, i_8_252_204_0, i_8_252_223_0,
    i_8_252_224_0, i_8_252_232_0, i_8_252_292_0, i_8_252_420_0,
    i_8_252_456_0, i_8_252_457_0, i_8_252_462_0, i_8_252_480_0,
    i_8_252_483_0, i_8_252_517_0, i_8_252_535_0, i_8_252_555_0,
    i_8_252_557_0, i_8_252_591_0, i_8_252_592_0, i_8_252_593_0,
    i_8_252_608_0, i_8_252_690_0, i_8_252_715_0, i_8_252_727_0,
    i_8_252_756_0, i_8_252_815_0, i_8_252_850_0, i_8_252_853_0,
    i_8_252_951_0, i_8_252_995_0, i_8_252_1052_0, i_8_252_1142_0,
    i_8_252_1174_0, i_8_252_1179_0, i_8_252_1180_0, i_8_252_1228_0,
    i_8_252_1230_0, i_8_252_1237_0, i_8_252_1261_0, i_8_252_1283_0,
    i_8_252_1308_0, i_8_252_1311_0, i_8_252_1312_0, i_8_252_1314_0,
    i_8_252_1316_0, i_8_252_1325_0, i_8_252_1329_0, i_8_252_1330_0,
    i_8_252_1346_0, i_8_252_1364_0, i_8_252_1401_0, i_8_252_1448_0,
    i_8_252_1462_0, i_8_252_1492_0, i_8_252_1497_0, i_8_252_1504_0,
    i_8_252_1507_0, i_8_252_1508_0, i_8_252_1555_0, i_8_252_1629_0,
    i_8_252_1634_0, i_8_252_1647_0, i_8_252_1648_0, i_8_252_1654_0,
    i_8_252_1670_0, i_8_252_1678_0, i_8_252_1679_0, i_8_252_1682_0,
    i_8_252_1720_0, i_8_252_1751_0, i_8_252_1753_0, i_8_252_1754_0,
    i_8_252_1805_0, i_8_252_1812_0, i_8_252_1824_0, i_8_252_1947_0,
    i_8_252_1948_0, i_8_252_1949_0, i_8_252_1951_0, i_8_252_2005_0,
    i_8_252_2055_0, i_8_252_2077_0, i_8_252_2158_0, i_8_252_2185_0,
    i_8_252_2217_0, i_8_252_2235_0, i_8_252_2236_0, i_8_252_2253_0,
    i_8_252_2275_0, i_8_252_2278_0, i_8_252_2293_0,
    o_8_252_0_0  );
  input  i_8_252_3_0, i_8_252_8_0, i_8_252_22_0, i_8_252_50_0,
    i_8_252_78_0, i_8_252_80_0, i_8_252_114_0, i_8_252_125_0,
    i_8_252_177_0, i_8_252_185_0, i_8_252_192_0, i_8_252_204_0,
    i_8_252_223_0, i_8_252_224_0, i_8_252_232_0, i_8_252_292_0,
    i_8_252_420_0, i_8_252_456_0, i_8_252_457_0, i_8_252_462_0,
    i_8_252_480_0, i_8_252_483_0, i_8_252_517_0, i_8_252_535_0,
    i_8_252_555_0, i_8_252_557_0, i_8_252_591_0, i_8_252_592_0,
    i_8_252_593_0, i_8_252_608_0, i_8_252_690_0, i_8_252_715_0,
    i_8_252_727_0, i_8_252_756_0, i_8_252_815_0, i_8_252_850_0,
    i_8_252_853_0, i_8_252_951_0, i_8_252_995_0, i_8_252_1052_0,
    i_8_252_1142_0, i_8_252_1174_0, i_8_252_1179_0, i_8_252_1180_0,
    i_8_252_1228_0, i_8_252_1230_0, i_8_252_1237_0, i_8_252_1261_0,
    i_8_252_1283_0, i_8_252_1308_0, i_8_252_1311_0, i_8_252_1312_0,
    i_8_252_1314_0, i_8_252_1316_0, i_8_252_1325_0, i_8_252_1329_0,
    i_8_252_1330_0, i_8_252_1346_0, i_8_252_1364_0, i_8_252_1401_0,
    i_8_252_1448_0, i_8_252_1462_0, i_8_252_1492_0, i_8_252_1497_0,
    i_8_252_1504_0, i_8_252_1507_0, i_8_252_1508_0, i_8_252_1555_0,
    i_8_252_1629_0, i_8_252_1634_0, i_8_252_1647_0, i_8_252_1648_0,
    i_8_252_1654_0, i_8_252_1670_0, i_8_252_1678_0, i_8_252_1679_0,
    i_8_252_1682_0, i_8_252_1720_0, i_8_252_1751_0, i_8_252_1753_0,
    i_8_252_1754_0, i_8_252_1805_0, i_8_252_1812_0, i_8_252_1824_0,
    i_8_252_1947_0, i_8_252_1948_0, i_8_252_1949_0, i_8_252_1951_0,
    i_8_252_2005_0, i_8_252_2055_0, i_8_252_2077_0, i_8_252_2158_0,
    i_8_252_2185_0, i_8_252_2217_0, i_8_252_2235_0, i_8_252_2236_0,
    i_8_252_2253_0, i_8_252_2275_0, i_8_252_2278_0, i_8_252_2293_0;
  output o_8_252_0_0;
  assign o_8_252_0_0 = ~((~i_8_252_125_0 & ((~i_8_252_177_0 & i_8_252_192_0 & ~i_8_252_462_0 & ~i_8_252_1312_0 & ~i_8_252_1316_0 & ~i_8_252_1329_0 & ~i_8_252_1330_0 & ~i_8_252_1462_0 & i_8_252_1824_0 & ~i_8_252_2217_0) | (~i_8_252_517_0 & ~i_8_252_1401_0 & ~i_8_252_1654_0 & ~i_8_252_1812_0 & ~i_8_252_2253_0))) | (~i_8_252_420_0 & ((~i_8_252_3_0 & ~i_8_252_535_0 & ~i_8_252_591_0 & ~i_8_252_592_0 & ~i_8_252_593_0 & ~i_8_252_1261_0 & ~i_8_252_1329_0 & ~i_8_252_1629_0) | (~i_8_252_177_0 & ~i_8_252_483_0 & ~i_8_252_517_0 & ~i_8_252_557_0 & ~i_8_252_1174_0 & ~i_8_252_1647_0 & ~i_8_252_1948_0))) | (~i_8_252_727_0 & ((~i_8_252_3_0 & ((~i_8_252_517_0 & ~i_8_252_1497_0 & ~i_8_252_1812_0 & ~i_8_252_1948_0 & ~i_8_252_1949_0 & ~i_8_252_2236_0) | (~i_8_252_1179_0 & ~i_8_252_1316_0 & ~i_8_252_1346_0 & ~i_8_252_1492_0 & ~i_8_252_2235_0 & ~i_8_252_2278_0))) | (~i_8_252_1311_0 & ((~i_8_252_591_0 & ~i_8_252_1179_0 & ~i_8_252_1308_0 & ~i_8_252_1812_0) | (~i_8_252_517_0 & ~i_8_252_1312_0 & ~i_8_252_1497_0 & ~i_8_252_1629_0 & ~i_8_252_1679_0 & ~i_8_252_1754_0 & ~i_8_252_2185_0 & ~i_8_252_2293_0))))) | (~i_8_252_456_0 & ((~i_8_252_78_0 & ~i_8_252_80_0 & ~i_8_252_204_0 & ~i_8_252_462_0 & ~i_8_252_593_0 & ~i_8_252_1174_0 & ~i_8_252_1330_0 & ~i_8_252_1462_0) | (~i_8_252_995_0 & ~i_8_252_1228_0 & ~i_8_252_1448_0 & ~i_8_252_1648_0 & ~i_8_252_1824_0))) | (~i_8_252_1497_0 & ((~i_8_252_204_0 & ~i_8_252_2005_0 & ((~i_8_252_22_0 & ~i_8_252_462_0 & ~i_8_252_517_0 & ~i_8_252_715_0 & ~i_8_252_1947_0) | (~i_8_252_1308_0 & ~i_8_252_1311_0 & ~i_8_252_1462_0 & ~i_8_252_2275_0))) | (~i_8_252_850_0 & ~i_8_252_1462_0 & ~i_8_252_1648_0 & ~i_8_252_1812_0 & ~i_8_252_1951_0 & ~i_8_252_2236_0))) | (~i_8_252_483_0 & ~i_8_252_1174_0 & ~i_8_252_1949_0 & ((i_8_252_457_0 & ~i_8_252_555_0 & ~i_8_252_1142_0 & ~i_8_252_1462_0 & ~i_8_252_1555_0 & ~i_8_252_1654_0) | (~i_8_252_457_0 & ~i_8_252_1314_0 & ~i_8_252_1401_0 & ~i_8_252_2158_0 & ~i_8_252_2293_0))) | (~i_8_252_1401_0 & ((~i_8_252_462_0 & ~i_8_252_1230_0 & ~i_8_252_1824_0 & ~i_8_252_1947_0 & ~i_8_252_1951_0 & ~i_8_252_2055_0) | (~i_8_252_690_0 & ~i_8_252_853_0 & ~i_8_252_1311_0 & ~i_8_252_1948_0 & ~i_8_252_2236_0))) | (i_8_252_850_0 & i_8_252_1462_0 & ~i_8_252_2236_0));
endmodule



// Benchmark "kernel_8_253" written by ABC on Sun Jul 19 10:07:30 2020

module kernel_8_253 ( 
    i_8_253_23_0, i_8_253_33_0, i_8_253_75_0, i_8_253_76_0, i_8_253_77_0,
    i_8_253_85_0, i_8_253_114_0, i_8_253_139_0, i_8_253_193_0,
    i_8_253_231_0, i_8_253_322_0, i_8_253_364_0, i_8_253_424_0,
    i_8_253_428_0, i_8_253_429_0, i_8_253_507_0, i_8_253_509_0,
    i_8_253_510_0, i_8_253_526_0, i_8_253_527_0, i_8_253_589_0,
    i_8_253_604_0, i_8_253_606_0, i_8_253_655_0, i_8_253_660_0,
    i_8_253_678_0, i_8_253_703_0, i_8_253_808_0, i_8_253_823_0,
    i_8_253_832_0, i_8_253_838_0, i_8_253_878_0, i_8_253_896_0,
    i_8_253_969_0, i_8_253_992_0, i_8_253_1012_0, i_8_253_1101_0,
    i_8_253_1155_0, i_8_253_1183_0, i_8_253_1189_0, i_8_253_1191_0,
    i_8_253_1229_0, i_8_253_1264_0, i_8_253_1266_0, i_8_253_1267_0,
    i_8_253_1282_0, i_8_253_1299_0, i_8_253_1318_0, i_8_253_1335_0,
    i_8_253_1336_0, i_8_253_1337_0, i_8_253_1366_0, i_8_253_1393_0,
    i_8_253_1399_0, i_8_253_1434_0, i_8_253_1437_0, i_8_253_1463_0,
    i_8_253_1508_0, i_8_253_1517_0, i_8_253_1519_0, i_8_253_1534_0,
    i_8_253_1543_0, i_8_253_1550_0, i_8_253_1625_0, i_8_253_1642_0,
    i_8_253_1686_0, i_8_253_1687_0, i_8_253_1689_0, i_8_253_1722_0,
    i_8_253_1723_0, i_8_253_1768_0, i_8_253_1770_0, i_8_253_1773_0,
    i_8_253_1774_0, i_8_253_1781_0, i_8_253_1782_0, i_8_253_1786_0,
    i_8_253_1804_0, i_8_253_1819_0, i_8_253_1822_0, i_8_253_1837_0,
    i_8_253_1848_0, i_8_253_1857_0, i_8_253_1858_0, i_8_253_1861_0,
    i_8_253_1866_0, i_8_253_1903_0, i_8_253_1938_0, i_8_253_1939_0,
    i_8_253_1995_0, i_8_253_1996_0, i_8_253_2029_0, i_8_253_2048_0,
    i_8_253_2118_0, i_8_253_2134_0, i_8_253_2149_0, i_8_253_2226_0,
    i_8_253_2245_0, i_8_253_2246_0, i_8_253_2247_0,
    o_8_253_0_0  );
  input  i_8_253_23_0, i_8_253_33_0, i_8_253_75_0, i_8_253_76_0,
    i_8_253_77_0, i_8_253_85_0, i_8_253_114_0, i_8_253_139_0,
    i_8_253_193_0, i_8_253_231_0, i_8_253_322_0, i_8_253_364_0,
    i_8_253_424_0, i_8_253_428_0, i_8_253_429_0, i_8_253_507_0,
    i_8_253_509_0, i_8_253_510_0, i_8_253_526_0, i_8_253_527_0,
    i_8_253_589_0, i_8_253_604_0, i_8_253_606_0, i_8_253_655_0,
    i_8_253_660_0, i_8_253_678_0, i_8_253_703_0, i_8_253_808_0,
    i_8_253_823_0, i_8_253_832_0, i_8_253_838_0, i_8_253_878_0,
    i_8_253_896_0, i_8_253_969_0, i_8_253_992_0, i_8_253_1012_0,
    i_8_253_1101_0, i_8_253_1155_0, i_8_253_1183_0, i_8_253_1189_0,
    i_8_253_1191_0, i_8_253_1229_0, i_8_253_1264_0, i_8_253_1266_0,
    i_8_253_1267_0, i_8_253_1282_0, i_8_253_1299_0, i_8_253_1318_0,
    i_8_253_1335_0, i_8_253_1336_0, i_8_253_1337_0, i_8_253_1366_0,
    i_8_253_1393_0, i_8_253_1399_0, i_8_253_1434_0, i_8_253_1437_0,
    i_8_253_1463_0, i_8_253_1508_0, i_8_253_1517_0, i_8_253_1519_0,
    i_8_253_1534_0, i_8_253_1543_0, i_8_253_1550_0, i_8_253_1625_0,
    i_8_253_1642_0, i_8_253_1686_0, i_8_253_1687_0, i_8_253_1689_0,
    i_8_253_1722_0, i_8_253_1723_0, i_8_253_1768_0, i_8_253_1770_0,
    i_8_253_1773_0, i_8_253_1774_0, i_8_253_1781_0, i_8_253_1782_0,
    i_8_253_1786_0, i_8_253_1804_0, i_8_253_1819_0, i_8_253_1822_0,
    i_8_253_1837_0, i_8_253_1848_0, i_8_253_1857_0, i_8_253_1858_0,
    i_8_253_1861_0, i_8_253_1866_0, i_8_253_1903_0, i_8_253_1938_0,
    i_8_253_1939_0, i_8_253_1995_0, i_8_253_1996_0, i_8_253_2029_0,
    i_8_253_2048_0, i_8_253_2118_0, i_8_253_2134_0, i_8_253_2149_0,
    i_8_253_2226_0, i_8_253_2245_0, i_8_253_2246_0, i_8_253_2247_0;
  output o_8_253_0_0;
  assign o_8_253_0_0 = ~((~i_8_253_1689_0 & ((~i_8_253_23_0 & ~i_8_253_655_0 & ~i_8_253_1995_0 & ((~i_8_253_509_0 & ~i_8_253_589_0 & ~i_8_253_1012_0 & ~i_8_253_1264_0 & ~i_8_253_1543_0 & ~i_8_253_1861_0) | (~i_8_253_838_0 & ~i_8_253_1508_0 & ~i_8_253_1686_0 & ~i_8_253_1939_0 & ~i_8_253_2226_0 & ~i_8_253_2245_0))) | (~i_8_253_604_0 & ~i_8_253_1723_0 & ((~i_8_253_429_0 & ~i_8_253_510_0 & ~i_8_253_1101_0 & ~i_8_253_1336_0 & ~i_8_253_1337_0 & ~i_8_253_1463_0 & ~i_8_253_1782_0 & ~i_8_253_1837_0) | (~i_8_253_606_0 & i_8_253_1299_0 & ~i_8_253_1543_0 & ~i_8_253_1686_0 & ~i_8_253_1770_0 & ~i_8_253_2246_0))) | (~i_8_253_823_0 & ~i_8_253_878_0 & ~i_8_253_896_0 & ~i_8_253_1266_0 & ~i_8_253_1299_0 & ~i_8_253_1463_0 & ~i_8_253_1508_0 & ~i_8_253_1517_0 & ~i_8_253_1686_0 & ~i_8_253_2246_0 & ~i_8_253_2247_0))) | (~i_8_253_231_0 & ((~i_8_253_75_0 & ~i_8_253_139_0 & ~i_8_253_1336_0 & ~i_8_253_1437_0 & ~i_8_253_1774_0 & ~i_8_253_1786_0 & ~i_8_253_1995_0) | (~i_8_253_76_0 & ~i_8_253_77_0 & ~i_8_253_808_0 & ~i_8_253_969_0 & ~i_8_253_1155_0 & ~i_8_253_1337_0 & ~i_8_253_1517_0 & ~i_8_253_1782_0 & ~i_8_253_2247_0))) | (i_8_253_364_0 & ((i_8_253_832_0 & ~i_8_253_1299_0 & ~i_8_253_1337_0) | (~i_8_253_139_0 & ~i_8_253_589_0 & ~i_8_253_678_0 & ~i_8_253_823_0 & ~i_8_253_1012_0 & ~i_8_253_1189_0 & ~i_8_253_1267_0 & ~i_8_253_1366_0 & ~i_8_253_1463_0))) | (~i_8_253_139_0 & ((~i_8_253_678_0 & ~i_8_253_1267_0 & ~i_8_253_1282_0 & ~i_8_253_1335_0 & ~i_8_253_1337_0 & i_8_253_1786_0 & i_8_253_1822_0 & ~i_8_253_1939_0) | (~i_8_253_1782_0 & ~i_8_253_1786_0 & ~i_8_253_1819_0 & ~i_8_253_2245_0 & ~i_8_253_2246_0))) | (~i_8_253_424_0 & ((~i_8_253_823_0 & ~i_8_253_1336_0 & ~i_8_253_1366_0 & ~i_8_253_1517_0 & ~i_8_253_1768_0 & ~i_8_253_2134_0) | (~i_8_253_969_0 & ~i_8_253_1229_0 & ~i_8_253_1819_0 & ~i_8_253_1822_0 & ~i_8_253_1996_0 & ~i_8_253_2245_0))) | (~i_8_253_969_0 & ((~i_8_253_678_0 & ~i_8_253_1517_0 & ~i_8_253_1519_0 & ~i_8_253_1768_0 & ~i_8_253_1770_0 & ~i_8_253_1938_0 & ~i_8_253_2134_0 & ~i_8_253_2246_0) | (~i_8_253_77_0 & ~i_8_253_1266_0 & ~i_8_253_1282_0 & ~i_8_253_1686_0 & ~i_8_253_2245_0 & ~i_8_253_2247_0))) | (~i_8_253_77_0 & ((~i_8_253_1155_0 & ~i_8_253_1264_0 & ~i_8_253_1266_0 & ~i_8_253_1336_0 & ~i_8_253_1463_0 & ~i_8_253_1786_0) | (~i_8_253_1335_0 & ~i_8_253_1366_0 & ~i_8_253_2134_0 & ~i_8_253_2246_0 & ~i_8_253_2247_0))) | (~i_8_253_1508_0 & ((~i_8_253_606_0 & ~i_8_253_896_0 & ~i_8_253_1335_0 & ~i_8_253_1336_0 & ~i_8_253_1723_0 & ~i_8_253_1782_0 & i_8_253_1804_0) | (~i_8_253_604_0 & i_8_253_660_0 & i_8_253_1191_0 & ~i_8_253_1996_0))) | (~i_8_253_678_0 & ((~i_8_253_509_0 & ((~i_8_253_604_0 & ~i_8_253_1267_0 & ~i_8_253_1463_0 & ~i_8_253_1519_0 & ~i_8_253_1550_0 & ~i_8_253_1786_0) | (~i_8_253_76_0 & ~i_8_253_1366_0 & ~i_8_253_1773_0 & ~i_8_253_1781_0 & ~i_8_253_2246_0))) | (~i_8_253_604_0 & ~i_8_253_1282_0 & ~i_8_253_1463_0 & ~i_8_253_1722_0 & ~i_8_253_1770_0 & ~i_8_253_1822_0) | (~i_8_253_838_0 & ~i_8_253_896_0 & ~i_8_253_1434_0 & ~i_8_253_1687_0 & ~i_8_253_1768_0 & ~i_8_253_1819_0 & ~i_8_253_2245_0))) | (~i_8_253_76_0 & ~i_8_253_1822_0 & ((~i_8_253_364_0 & ~i_8_253_1723_0 & ~i_8_253_1938_0 & ~i_8_253_2029_0 & ~i_8_253_2134_0 & ~i_8_253_2246_0) | (~i_8_253_1782_0 & ~i_8_253_2247_0 & ~i_8_253_896_0 & ~i_8_253_1773_0))) | (i_8_253_1848_0 & i_8_253_1858_0) | (~i_8_253_509_0 & ~i_8_253_660_0 & ~i_8_253_1463_0 & i_8_253_1642_0 & ~i_8_253_1939_0));
endmodule



// Benchmark "kernel_8_254" written by ABC on Sun Jul 19 10:07:31 2020

module kernel_8_254 ( 
    i_8_254_22_0, i_8_254_88_0, i_8_254_141_0, i_8_254_203_0,
    i_8_254_206_0, i_8_254_229_0, i_8_254_240_0, i_8_254_257_0,
    i_8_254_265_0, i_8_254_310_0, i_8_254_328_0, i_8_254_337_0,
    i_8_254_345_0, i_8_254_355_0, i_8_254_373_0, i_8_254_382_0,
    i_8_254_426_0, i_8_254_427_0, i_8_254_430_0, i_8_254_455_0,
    i_8_254_457_0, i_8_254_490_0, i_8_254_505_0, i_8_254_524_0,
    i_8_254_554_0, i_8_254_556_0, i_8_254_565_0, i_8_254_569_0,
    i_8_254_604_0, i_8_254_626_0, i_8_254_627_0, i_8_254_676_0,
    i_8_254_710_0, i_8_254_752_0, i_8_254_761_0, i_8_254_770_0,
    i_8_254_778_0, i_8_254_836_0, i_8_254_938_0, i_8_254_951_0,
    i_8_254_1039_0, i_8_254_1088_0, i_8_254_1108_0, i_8_254_1112_0,
    i_8_254_1114_0, i_8_254_1115_0, i_8_254_1147_0, i_8_254_1264_0,
    i_8_254_1306_0, i_8_254_1329_0, i_8_254_1366_0, i_8_254_1369_0,
    i_8_254_1404_0, i_8_254_1407_0, i_8_254_1414_0, i_8_254_1433_0,
    i_8_254_1462_0, i_8_254_1480_0, i_8_254_1481_0, i_8_254_1490_0,
    i_8_254_1493_0, i_8_254_1543_0, i_8_254_1546_0, i_8_254_1552_0,
    i_8_254_1553_0, i_8_254_1562_0, i_8_254_1582_0, i_8_254_1651_0,
    i_8_254_1654_0, i_8_254_1677_0, i_8_254_1681_0, i_8_254_1706_0,
    i_8_254_1717_0, i_8_254_1723_0, i_8_254_1732_0, i_8_254_1733_0,
    i_8_254_1774_0, i_8_254_1778_0, i_8_254_1805_0, i_8_254_1814_0,
    i_8_254_1820_0, i_8_254_1821_0, i_8_254_1823_0, i_8_254_1826_0,
    i_8_254_1883_0, i_8_254_1888_0, i_8_254_1894_0, i_8_254_1903_0,
    i_8_254_1915_0, i_8_254_1957_0, i_8_254_1964_0, i_8_254_1984_0,
    i_8_254_1993_0, i_8_254_2105_0, i_8_254_2127_0, i_8_254_2150_0,
    i_8_254_2224_0, i_8_254_2266_0, i_8_254_2268_0, i_8_254_2290_0,
    o_8_254_0_0  );
  input  i_8_254_22_0, i_8_254_88_0, i_8_254_141_0, i_8_254_203_0,
    i_8_254_206_0, i_8_254_229_0, i_8_254_240_0, i_8_254_257_0,
    i_8_254_265_0, i_8_254_310_0, i_8_254_328_0, i_8_254_337_0,
    i_8_254_345_0, i_8_254_355_0, i_8_254_373_0, i_8_254_382_0,
    i_8_254_426_0, i_8_254_427_0, i_8_254_430_0, i_8_254_455_0,
    i_8_254_457_0, i_8_254_490_0, i_8_254_505_0, i_8_254_524_0,
    i_8_254_554_0, i_8_254_556_0, i_8_254_565_0, i_8_254_569_0,
    i_8_254_604_0, i_8_254_626_0, i_8_254_627_0, i_8_254_676_0,
    i_8_254_710_0, i_8_254_752_0, i_8_254_761_0, i_8_254_770_0,
    i_8_254_778_0, i_8_254_836_0, i_8_254_938_0, i_8_254_951_0,
    i_8_254_1039_0, i_8_254_1088_0, i_8_254_1108_0, i_8_254_1112_0,
    i_8_254_1114_0, i_8_254_1115_0, i_8_254_1147_0, i_8_254_1264_0,
    i_8_254_1306_0, i_8_254_1329_0, i_8_254_1366_0, i_8_254_1369_0,
    i_8_254_1404_0, i_8_254_1407_0, i_8_254_1414_0, i_8_254_1433_0,
    i_8_254_1462_0, i_8_254_1480_0, i_8_254_1481_0, i_8_254_1490_0,
    i_8_254_1493_0, i_8_254_1543_0, i_8_254_1546_0, i_8_254_1552_0,
    i_8_254_1553_0, i_8_254_1562_0, i_8_254_1582_0, i_8_254_1651_0,
    i_8_254_1654_0, i_8_254_1677_0, i_8_254_1681_0, i_8_254_1706_0,
    i_8_254_1717_0, i_8_254_1723_0, i_8_254_1732_0, i_8_254_1733_0,
    i_8_254_1774_0, i_8_254_1778_0, i_8_254_1805_0, i_8_254_1814_0,
    i_8_254_1820_0, i_8_254_1821_0, i_8_254_1823_0, i_8_254_1826_0,
    i_8_254_1883_0, i_8_254_1888_0, i_8_254_1894_0, i_8_254_1903_0,
    i_8_254_1915_0, i_8_254_1957_0, i_8_254_1964_0, i_8_254_1984_0,
    i_8_254_1993_0, i_8_254_2105_0, i_8_254_2127_0, i_8_254_2150_0,
    i_8_254_2224_0, i_8_254_2266_0, i_8_254_2268_0, i_8_254_2290_0;
  output o_8_254_0_0;
  assign o_8_254_0_0 = 0;
endmodule



// Benchmark "kernel_8_255" written by ABC on Sun Jul 19 10:07:32 2020

module kernel_8_255 ( 
    i_8_255_54_0, i_8_255_63_0, i_8_255_84_0, i_8_255_145_0, i_8_255_191_0,
    i_8_255_255_0, i_8_255_285_0, i_8_255_303_0, i_8_255_318_0,
    i_8_255_383_0, i_8_255_385_0, i_8_255_386_0, i_8_255_420_0,
    i_8_255_423_0, i_8_255_438_0, i_8_255_445_0, i_8_255_450_0,
    i_8_255_453_0, i_8_255_499_0, i_8_255_507_0, i_8_255_508_0,
    i_8_255_523_0, i_8_255_529_0, i_8_255_537_0, i_8_255_564_0,
    i_8_255_628_0, i_8_255_633_0, i_8_255_637_0, i_8_255_648_0,
    i_8_255_664_0, i_8_255_696_0, i_8_255_709_0, i_8_255_760_0,
    i_8_255_763_0, i_8_255_768_0, i_8_255_777_0, i_8_255_782_0,
    i_8_255_865_0, i_8_255_894_0, i_8_255_895_0, i_8_255_933_0,
    i_8_255_969_0, i_8_255_975_0, i_8_255_996_0, i_8_255_1095_0,
    i_8_255_1098_0, i_8_255_1108_0, i_8_255_1110_0, i_8_255_1111_0,
    i_8_255_1113_0, i_8_255_1119_0, i_8_255_1237_0, i_8_255_1264_0,
    i_8_255_1269_0, i_8_255_1314_0, i_8_255_1317_0, i_8_255_1324_0,
    i_8_255_1365_0, i_8_255_1401_0, i_8_255_1450_0, i_8_255_1506_0,
    i_8_255_1512_0, i_8_255_1515_0, i_8_255_1533_0, i_8_255_1561_0,
    i_8_255_1629_0, i_8_255_1635_0, i_8_255_1636_0, i_8_255_1670_0,
    i_8_255_1677_0, i_8_255_1678_0, i_8_255_1680_0, i_8_255_1681_0,
    i_8_255_1683_0, i_8_255_1686_0, i_8_255_1701_0, i_8_255_1704_0,
    i_8_255_1746_0, i_8_255_1753_0, i_8_255_1773_0, i_8_255_1780_0,
    i_8_255_1790_0, i_8_255_1791_0, i_8_255_1804_0, i_8_255_1818_0,
    i_8_255_1819_0, i_8_255_1822_0, i_8_255_1825_0, i_8_255_1845_0,
    i_8_255_1858_0, i_8_255_1867_0, i_8_255_1881_0, i_8_255_1885_0,
    i_8_255_1917_0, i_8_255_2044_0, i_8_255_2125_0, i_8_255_2142_0,
    i_8_255_2145_0, i_8_255_2232_0, i_8_255_2233_0,
    o_8_255_0_0  );
  input  i_8_255_54_0, i_8_255_63_0, i_8_255_84_0, i_8_255_145_0,
    i_8_255_191_0, i_8_255_255_0, i_8_255_285_0, i_8_255_303_0,
    i_8_255_318_0, i_8_255_383_0, i_8_255_385_0, i_8_255_386_0,
    i_8_255_420_0, i_8_255_423_0, i_8_255_438_0, i_8_255_445_0,
    i_8_255_450_0, i_8_255_453_0, i_8_255_499_0, i_8_255_507_0,
    i_8_255_508_0, i_8_255_523_0, i_8_255_529_0, i_8_255_537_0,
    i_8_255_564_0, i_8_255_628_0, i_8_255_633_0, i_8_255_637_0,
    i_8_255_648_0, i_8_255_664_0, i_8_255_696_0, i_8_255_709_0,
    i_8_255_760_0, i_8_255_763_0, i_8_255_768_0, i_8_255_777_0,
    i_8_255_782_0, i_8_255_865_0, i_8_255_894_0, i_8_255_895_0,
    i_8_255_933_0, i_8_255_969_0, i_8_255_975_0, i_8_255_996_0,
    i_8_255_1095_0, i_8_255_1098_0, i_8_255_1108_0, i_8_255_1110_0,
    i_8_255_1111_0, i_8_255_1113_0, i_8_255_1119_0, i_8_255_1237_0,
    i_8_255_1264_0, i_8_255_1269_0, i_8_255_1314_0, i_8_255_1317_0,
    i_8_255_1324_0, i_8_255_1365_0, i_8_255_1401_0, i_8_255_1450_0,
    i_8_255_1506_0, i_8_255_1512_0, i_8_255_1515_0, i_8_255_1533_0,
    i_8_255_1561_0, i_8_255_1629_0, i_8_255_1635_0, i_8_255_1636_0,
    i_8_255_1670_0, i_8_255_1677_0, i_8_255_1678_0, i_8_255_1680_0,
    i_8_255_1681_0, i_8_255_1683_0, i_8_255_1686_0, i_8_255_1701_0,
    i_8_255_1704_0, i_8_255_1746_0, i_8_255_1753_0, i_8_255_1773_0,
    i_8_255_1780_0, i_8_255_1790_0, i_8_255_1791_0, i_8_255_1804_0,
    i_8_255_1818_0, i_8_255_1819_0, i_8_255_1822_0, i_8_255_1825_0,
    i_8_255_1845_0, i_8_255_1858_0, i_8_255_1867_0, i_8_255_1881_0,
    i_8_255_1885_0, i_8_255_1917_0, i_8_255_2044_0, i_8_255_2125_0,
    i_8_255_2142_0, i_8_255_2145_0, i_8_255_2232_0, i_8_255_2233_0;
  output o_8_255_0_0;
  assign o_8_255_0_0 = 0;
endmodule



// Benchmark "kernel_8_256" written by ABC on Sun Jul 19 10:07:32 2020

module kernel_8_256 ( 
    i_8_256_22_0, i_8_256_37_0, i_8_256_40_0, i_8_256_49_0, i_8_256_94_0,
    i_8_256_124_0, i_8_256_157_0, i_8_256_165_0, i_8_256_166_0,
    i_8_256_213_0, i_8_256_256_0, i_8_256_287_0, i_8_256_292_0,
    i_8_256_328_0, i_8_256_337_0, i_8_256_361_0, i_8_256_363_0,
    i_8_256_427_0, i_8_256_453_0, i_8_256_492_0, i_8_256_571_0,
    i_8_256_583_0, i_8_256_599_0, i_8_256_627_0, i_8_256_682_0,
    i_8_256_703_0, i_8_256_706_0, i_8_256_744_0, i_8_256_759_0,
    i_8_256_772_0, i_8_256_773_0, i_8_256_787_0, i_8_256_805_0,
    i_8_256_823_0, i_8_256_842_0, i_8_256_876_0, i_8_256_880_0,
    i_8_256_955_0, i_8_256_967_0, i_8_256_979_0, i_8_256_1002_0,
    i_8_256_1040_0, i_8_256_1057_0, i_8_256_1066_0, i_8_256_1110_0,
    i_8_256_1111_0, i_8_256_1185_0, i_8_256_1227_0, i_8_256_1228_0,
    i_8_256_1229_0, i_8_256_1231_0, i_8_256_1249_0, i_8_256_1255_0,
    i_8_256_1257_0, i_8_256_1267_0, i_8_256_1279_0, i_8_256_1305_0,
    i_8_256_1327_0, i_8_256_1351_0, i_8_256_1357_0, i_8_256_1372_0,
    i_8_256_1375_0, i_8_256_1380_0, i_8_256_1381_0, i_8_256_1438_0,
    i_8_256_1447_0, i_8_256_1453_0, i_8_256_1455_0, i_8_256_1456_0,
    i_8_256_1467_0, i_8_256_1471_0, i_8_256_1578_0, i_8_256_1606_0,
    i_8_256_1614_0, i_8_256_1639_0, i_8_256_1651_0, i_8_256_1671_0,
    i_8_256_1696_0, i_8_256_1699_0, i_8_256_1701_0, i_8_256_1733_0,
    i_8_256_1749_0, i_8_256_1768_0, i_8_256_1821_0, i_8_256_1857_0,
    i_8_256_1939_0, i_8_256_1981_0, i_8_256_1992_0, i_8_256_2040_0,
    i_8_256_2055_0, i_8_256_2074_0, i_8_256_2164_0, i_8_256_2185_0,
    i_8_256_2200_0, i_8_256_2227_0, i_8_256_2238_0, i_8_256_2239_0,
    i_8_256_2259_0, i_8_256_2263_0, i_8_256_2284_0,
    o_8_256_0_0  );
  input  i_8_256_22_0, i_8_256_37_0, i_8_256_40_0, i_8_256_49_0,
    i_8_256_94_0, i_8_256_124_0, i_8_256_157_0, i_8_256_165_0,
    i_8_256_166_0, i_8_256_213_0, i_8_256_256_0, i_8_256_287_0,
    i_8_256_292_0, i_8_256_328_0, i_8_256_337_0, i_8_256_361_0,
    i_8_256_363_0, i_8_256_427_0, i_8_256_453_0, i_8_256_492_0,
    i_8_256_571_0, i_8_256_583_0, i_8_256_599_0, i_8_256_627_0,
    i_8_256_682_0, i_8_256_703_0, i_8_256_706_0, i_8_256_744_0,
    i_8_256_759_0, i_8_256_772_0, i_8_256_773_0, i_8_256_787_0,
    i_8_256_805_0, i_8_256_823_0, i_8_256_842_0, i_8_256_876_0,
    i_8_256_880_0, i_8_256_955_0, i_8_256_967_0, i_8_256_979_0,
    i_8_256_1002_0, i_8_256_1040_0, i_8_256_1057_0, i_8_256_1066_0,
    i_8_256_1110_0, i_8_256_1111_0, i_8_256_1185_0, i_8_256_1227_0,
    i_8_256_1228_0, i_8_256_1229_0, i_8_256_1231_0, i_8_256_1249_0,
    i_8_256_1255_0, i_8_256_1257_0, i_8_256_1267_0, i_8_256_1279_0,
    i_8_256_1305_0, i_8_256_1327_0, i_8_256_1351_0, i_8_256_1357_0,
    i_8_256_1372_0, i_8_256_1375_0, i_8_256_1380_0, i_8_256_1381_0,
    i_8_256_1438_0, i_8_256_1447_0, i_8_256_1453_0, i_8_256_1455_0,
    i_8_256_1456_0, i_8_256_1467_0, i_8_256_1471_0, i_8_256_1578_0,
    i_8_256_1606_0, i_8_256_1614_0, i_8_256_1639_0, i_8_256_1651_0,
    i_8_256_1671_0, i_8_256_1696_0, i_8_256_1699_0, i_8_256_1701_0,
    i_8_256_1733_0, i_8_256_1749_0, i_8_256_1768_0, i_8_256_1821_0,
    i_8_256_1857_0, i_8_256_1939_0, i_8_256_1981_0, i_8_256_1992_0,
    i_8_256_2040_0, i_8_256_2055_0, i_8_256_2074_0, i_8_256_2164_0,
    i_8_256_2185_0, i_8_256_2200_0, i_8_256_2227_0, i_8_256_2238_0,
    i_8_256_2239_0, i_8_256_2259_0, i_8_256_2263_0, i_8_256_2284_0;
  output o_8_256_0_0;
  assign o_8_256_0_0 = 0;
endmodule



// Benchmark "kernel_8_257" written by ABC on Sun Jul 19 10:07:33 2020

module kernel_8_257 ( 
    i_8_257_37_0, i_8_257_82_0, i_8_257_165_0, i_8_257_210_0,
    i_8_257_262_0, i_8_257_265_0, i_8_257_279_0, i_8_257_307_0,
    i_8_257_336_0, i_8_257_358_0, i_8_257_384_0, i_8_257_393_0,
    i_8_257_394_0, i_8_257_421_0, i_8_257_456_0, i_8_257_489_0,
    i_8_257_492_0, i_8_257_498_0, i_8_257_527_0, i_8_257_549_0,
    i_8_257_591_0, i_8_257_622_0, i_8_257_625_0, i_8_257_636_0,
    i_8_257_637_0, i_8_257_642_0, i_8_257_658_0, i_8_257_660_0,
    i_8_257_663_0, i_8_257_673_0, i_8_257_688_0, i_8_257_696_0,
    i_8_257_699_0, i_8_257_701_0, i_8_257_729_0, i_8_257_747_0,
    i_8_257_751_0, i_8_257_837_0, i_8_257_843_0, i_8_257_874_0,
    i_8_257_882_0, i_8_257_921_0, i_8_257_930_0, i_8_257_973_0,
    i_8_257_983_0, i_8_257_1009_0, i_8_257_1050_0, i_8_257_1056_0,
    i_8_257_1071_0, i_8_257_1075_0, i_8_257_1084_0, i_8_257_1129_0,
    i_8_257_1182_0, i_8_257_1228_0, i_8_257_1234_0, i_8_257_1263_0,
    i_8_257_1278_0, i_8_257_1291_0, i_8_257_1296_0, i_8_257_1306_0,
    i_8_257_1357_0, i_8_257_1362_0, i_8_257_1383_0, i_8_257_1390_0,
    i_8_257_1399_0, i_8_257_1410_0, i_8_257_1411_0, i_8_257_1435_0,
    i_8_257_1440_0, i_8_257_1441_0, i_8_257_1479_0, i_8_257_1507_0,
    i_8_257_1548_0, i_8_257_1551_0, i_8_257_1565_0, i_8_257_1608_0,
    i_8_257_1681_0, i_8_257_1683_0, i_8_257_1687_0, i_8_257_1720_0,
    i_8_257_1729_0, i_8_257_1731_0, i_8_257_1746_0, i_8_257_1747_0,
    i_8_257_1752_0, i_8_257_1768_0, i_8_257_1824_0, i_8_257_1855_0,
    i_8_257_1884_0, i_8_257_1887_0, i_8_257_1980_0, i_8_257_1989_0,
    i_8_257_2019_0, i_8_257_2052_0, i_8_257_2070_0, i_8_257_2118_0,
    i_8_257_2142_0, i_8_257_2148_0, i_8_257_2226_0, i_8_257_2286_0,
    o_8_257_0_0  );
  input  i_8_257_37_0, i_8_257_82_0, i_8_257_165_0, i_8_257_210_0,
    i_8_257_262_0, i_8_257_265_0, i_8_257_279_0, i_8_257_307_0,
    i_8_257_336_0, i_8_257_358_0, i_8_257_384_0, i_8_257_393_0,
    i_8_257_394_0, i_8_257_421_0, i_8_257_456_0, i_8_257_489_0,
    i_8_257_492_0, i_8_257_498_0, i_8_257_527_0, i_8_257_549_0,
    i_8_257_591_0, i_8_257_622_0, i_8_257_625_0, i_8_257_636_0,
    i_8_257_637_0, i_8_257_642_0, i_8_257_658_0, i_8_257_660_0,
    i_8_257_663_0, i_8_257_673_0, i_8_257_688_0, i_8_257_696_0,
    i_8_257_699_0, i_8_257_701_0, i_8_257_729_0, i_8_257_747_0,
    i_8_257_751_0, i_8_257_837_0, i_8_257_843_0, i_8_257_874_0,
    i_8_257_882_0, i_8_257_921_0, i_8_257_930_0, i_8_257_973_0,
    i_8_257_983_0, i_8_257_1009_0, i_8_257_1050_0, i_8_257_1056_0,
    i_8_257_1071_0, i_8_257_1075_0, i_8_257_1084_0, i_8_257_1129_0,
    i_8_257_1182_0, i_8_257_1228_0, i_8_257_1234_0, i_8_257_1263_0,
    i_8_257_1278_0, i_8_257_1291_0, i_8_257_1296_0, i_8_257_1306_0,
    i_8_257_1357_0, i_8_257_1362_0, i_8_257_1383_0, i_8_257_1390_0,
    i_8_257_1399_0, i_8_257_1410_0, i_8_257_1411_0, i_8_257_1435_0,
    i_8_257_1440_0, i_8_257_1441_0, i_8_257_1479_0, i_8_257_1507_0,
    i_8_257_1548_0, i_8_257_1551_0, i_8_257_1565_0, i_8_257_1608_0,
    i_8_257_1681_0, i_8_257_1683_0, i_8_257_1687_0, i_8_257_1720_0,
    i_8_257_1729_0, i_8_257_1731_0, i_8_257_1746_0, i_8_257_1747_0,
    i_8_257_1752_0, i_8_257_1768_0, i_8_257_1824_0, i_8_257_1855_0,
    i_8_257_1884_0, i_8_257_1887_0, i_8_257_1980_0, i_8_257_1989_0,
    i_8_257_2019_0, i_8_257_2052_0, i_8_257_2070_0, i_8_257_2118_0,
    i_8_257_2142_0, i_8_257_2148_0, i_8_257_2226_0, i_8_257_2286_0;
  output o_8_257_0_0;
  assign o_8_257_0_0 = 0;
endmodule



// Benchmark "kernel_8_258" written by ABC on Sun Jul 19 10:07:34 2020

module kernel_8_258 ( 
    i_8_258_1_0, i_8_258_22_0, i_8_258_57_0, i_8_258_85_0, i_8_258_96_0,
    i_8_258_103_0, i_8_258_104_0, i_8_258_105_0, i_8_258_165_0,
    i_8_258_168_0, i_8_258_202_0, i_8_258_210_0, i_8_258_211_0,
    i_8_258_214_0, i_8_258_219_0, i_8_258_220_0, i_8_258_223_0,
    i_8_258_256_0, i_8_258_292_0, i_8_258_333_0, i_8_258_345_0,
    i_8_258_361_0, i_8_258_415_0, i_8_258_445_0, i_8_258_448_0,
    i_8_258_475_0, i_8_258_501_0, i_8_258_589_0, i_8_258_596_0,
    i_8_258_606_0, i_8_258_627_0, i_8_258_658_0, i_8_258_669_0,
    i_8_258_670_0, i_8_258_716_0, i_8_258_768_0, i_8_258_786_0,
    i_8_258_888_0, i_8_258_949_0, i_8_258_977_0, i_8_258_984_0,
    i_8_258_985_0, i_8_258_991_0, i_8_258_992_0, i_8_258_1084_0,
    i_8_258_1110_0, i_8_258_1113_0, i_8_258_1155_0, i_8_258_1216_0,
    i_8_258_1222_0, i_8_258_1232_0, i_8_258_1248_0, i_8_258_1267_0,
    i_8_258_1272_0, i_8_258_1344_0, i_8_258_1347_0, i_8_258_1402_0,
    i_8_258_1419_0, i_8_258_1420_0, i_8_258_1423_0, i_8_258_1428_0,
    i_8_258_1437_0, i_8_258_1467_0, i_8_258_1477_0, i_8_258_1489_0,
    i_8_258_1518_0, i_8_258_1524_0, i_8_258_1544_0, i_8_258_1555_0,
    i_8_258_1588_0, i_8_258_1615_0, i_8_258_1618_0, i_8_258_1636_0,
    i_8_258_1677_0, i_8_258_1678_0, i_8_258_1680_0, i_8_258_1704_0,
    i_8_258_1720_0, i_8_258_1749_0, i_8_258_1780_0, i_8_258_1783_0,
    i_8_258_1785_0, i_8_258_1786_0, i_8_258_1825_0, i_8_258_1855_0,
    i_8_258_1861_0, i_8_258_1902_0, i_8_258_1963_0, i_8_258_2009_0,
    i_8_258_2026_0, i_8_258_2126_0, i_8_258_2128_0, i_8_258_2139_0,
    i_8_258_2140_0, i_8_258_2143_0, i_8_258_2150_0, i_8_258_2152_0,
    i_8_258_2236_0, i_8_258_2293_0, i_8_258_2294_0,
    o_8_258_0_0  );
  input  i_8_258_1_0, i_8_258_22_0, i_8_258_57_0, i_8_258_85_0,
    i_8_258_96_0, i_8_258_103_0, i_8_258_104_0, i_8_258_105_0,
    i_8_258_165_0, i_8_258_168_0, i_8_258_202_0, i_8_258_210_0,
    i_8_258_211_0, i_8_258_214_0, i_8_258_219_0, i_8_258_220_0,
    i_8_258_223_0, i_8_258_256_0, i_8_258_292_0, i_8_258_333_0,
    i_8_258_345_0, i_8_258_361_0, i_8_258_415_0, i_8_258_445_0,
    i_8_258_448_0, i_8_258_475_0, i_8_258_501_0, i_8_258_589_0,
    i_8_258_596_0, i_8_258_606_0, i_8_258_627_0, i_8_258_658_0,
    i_8_258_669_0, i_8_258_670_0, i_8_258_716_0, i_8_258_768_0,
    i_8_258_786_0, i_8_258_888_0, i_8_258_949_0, i_8_258_977_0,
    i_8_258_984_0, i_8_258_985_0, i_8_258_991_0, i_8_258_992_0,
    i_8_258_1084_0, i_8_258_1110_0, i_8_258_1113_0, i_8_258_1155_0,
    i_8_258_1216_0, i_8_258_1222_0, i_8_258_1232_0, i_8_258_1248_0,
    i_8_258_1267_0, i_8_258_1272_0, i_8_258_1344_0, i_8_258_1347_0,
    i_8_258_1402_0, i_8_258_1419_0, i_8_258_1420_0, i_8_258_1423_0,
    i_8_258_1428_0, i_8_258_1437_0, i_8_258_1467_0, i_8_258_1477_0,
    i_8_258_1489_0, i_8_258_1518_0, i_8_258_1524_0, i_8_258_1544_0,
    i_8_258_1555_0, i_8_258_1588_0, i_8_258_1615_0, i_8_258_1618_0,
    i_8_258_1636_0, i_8_258_1677_0, i_8_258_1678_0, i_8_258_1680_0,
    i_8_258_1704_0, i_8_258_1720_0, i_8_258_1749_0, i_8_258_1780_0,
    i_8_258_1783_0, i_8_258_1785_0, i_8_258_1786_0, i_8_258_1825_0,
    i_8_258_1855_0, i_8_258_1861_0, i_8_258_1902_0, i_8_258_1963_0,
    i_8_258_2009_0, i_8_258_2026_0, i_8_258_2126_0, i_8_258_2128_0,
    i_8_258_2139_0, i_8_258_2140_0, i_8_258_2143_0, i_8_258_2150_0,
    i_8_258_2152_0, i_8_258_2236_0, i_8_258_2293_0, i_8_258_2294_0;
  output o_8_258_0_0;
  assign o_8_258_0_0 = 0;
endmodule



// Benchmark "kernel_8_259" written by ABC on Sun Jul 19 10:07:35 2020

module kernel_8_259 ( 
    i_8_259_41_0, i_8_259_83_0, i_8_259_104_0, i_8_259_115_0,
    i_8_259_166_0, i_8_259_247_0, i_8_259_266_0, i_8_259_283_0,
    i_8_259_302_0, i_8_259_304_0, i_8_259_326_0, i_8_259_362_0,
    i_8_259_364_0, i_8_259_383_0, i_8_259_419_0, i_8_259_427_0,
    i_8_259_437_0, i_8_259_440_0, i_8_259_451_0, i_8_259_457_0,
    i_8_259_490_0, i_8_259_500_0, i_8_259_505_0, i_8_259_527_0,
    i_8_259_545_0, i_8_259_548_0, i_8_259_572_0, i_8_259_594_0,
    i_8_259_598_0, i_8_259_599_0, i_8_259_635_0, i_8_259_643_0,
    i_8_259_658_0, i_8_259_662_0, i_8_259_695_0, i_8_259_698_0,
    i_8_259_699_0, i_8_259_700_0, i_8_259_716_0, i_8_259_781_0,
    i_8_259_782_0, i_8_259_787_0, i_8_259_789_0, i_8_259_808_0,
    i_8_259_812_0, i_8_259_815_0, i_8_259_824_0, i_8_259_841_0,
    i_8_259_853_0, i_8_259_877_0, i_8_259_974_0, i_8_259_992_0,
    i_8_259_1061_0, i_8_259_1067_0, i_8_259_1211_0, i_8_259_1224_0,
    i_8_259_1228_0, i_8_259_1236_0, i_8_259_1253_0, i_8_259_1273_0,
    i_8_259_1296_0, i_8_259_1358_0, i_8_259_1365_0, i_8_259_1399_0,
    i_8_259_1426_0, i_8_259_1444_0, i_8_259_1471_0, i_8_259_1552_0,
    i_8_259_1589_0, i_8_259_1637_0, i_8_259_1697_0, i_8_259_1700_0,
    i_8_259_1705_0, i_8_259_1747_0, i_8_259_1768_0, i_8_259_1781_0,
    i_8_259_1783_0, i_8_259_1787_0, i_8_259_1805_0, i_8_259_1807_0,
    i_8_259_1851_0, i_8_259_1854_0, i_8_259_1855_0, i_8_259_1858_0,
    i_8_259_1859_0, i_8_259_1886_0, i_8_259_1949_0, i_8_259_1984_0,
    i_8_259_1993_0, i_8_259_1995_0, i_8_259_2029_0, i_8_259_2032_0,
    i_8_259_2090_0, i_8_259_2117_0, i_8_259_2134_0, i_8_259_2137_0,
    i_8_259_2155_0, i_8_259_2162_0, i_8_259_2191_0, i_8_259_2244_0,
    o_8_259_0_0  );
  input  i_8_259_41_0, i_8_259_83_0, i_8_259_104_0, i_8_259_115_0,
    i_8_259_166_0, i_8_259_247_0, i_8_259_266_0, i_8_259_283_0,
    i_8_259_302_0, i_8_259_304_0, i_8_259_326_0, i_8_259_362_0,
    i_8_259_364_0, i_8_259_383_0, i_8_259_419_0, i_8_259_427_0,
    i_8_259_437_0, i_8_259_440_0, i_8_259_451_0, i_8_259_457_0,
    i_8_259_490_0, i_8_259_500_0, i_8_259_505_0, i_8_259_527_0,
    i_8_259_545_0, i_8_259_548_0, i_8_259_572_0, i_8_259_594_0,
    i_8_259_598_0, i_8_259_599_0, i_8_259_635_0, i_8_259_643_0,
    i_8_259_658_0, i_8_259_662_0, i_8_259_695_0, i_8_259_698_0,
    i_8_259_699_0, i_8_259_700_0, i_8_259_716_0, i_8_259_781_0,
    i_8_259_782_0, i_8_259_787_0, i_8_259_789_0, i_8_259_808_0,
    i_8_259_812_0, i_8_259_815_0, i_8_259_824_0, i_8_259_841_0,
    i_8_259_853_0, i_8_259_877_0, i_8_259_974_0, i_8_259_992_0,
    i_8_259_1061_0, i_8_259_1067_0, i_8_259_1211_0, i_8_259_1224_0,
    i_8_259_1228_0, i_8_259_1236_0, i_8_259_1253_0, i_8_259_1273_0,
    i_8_259_1296_0, i_8_259_1358_0, i_8_259_1365_0, i_8_259_1399_0,
    i_8_259_1426_0, i_8_259_1444_0, i_8_259_1471_0, i_8_259_1552_0,
    i_8_259_1589_0, i_8_259_1637_0, i_8_259_1697_0, i_8_259_1700_0,
    i_8_259_1705_0, i_8_259_1747_0, i_8_259_1768_0, i_8_259_1781_0,
    i_8_259_1783_0, i_8_259_1787_0, i_8_259_1805_0, i_8_259_1807_0,
    i_8_259_1851_0, i_8_259_1854_0, i_8_259_1855_0, i_8_259_1858_0,
    i_8_259_1859_0, i_8_259_1886_0, i_8_259_1949_0, i_8_259_1984_0,
    i_8_259_1993_0, i_8_259_1995_0, i_8_259_2029_0, i_8_259_2032_0,
    i_8_259_2090_0, i_8_259_2117_0, i_8_259_2134_0, i_8_259_2137_0,
    i_8_259_2155_0, i_8_259_2162_0, i_8_259_2191_0, i_8_259_2244_0;
  output o_8_259_0_0;
  assign o_8_259_0_0 = 0;
endmodule



// Benchmark "kernel_8_260" written by ABC on Sun Jul 19 10:07:36 2020

module kernel_8_260 ( 
    i_8_260_6_0, i_8_260_14_0, i_8_260_44_0, i_8_260_106_0, i_8_260_140_0,
    i_8_260_196_0, i_8_260_197_0, i_8_260_214_0, i_8_260_222_0,
    i_8_260_228_0, i_8_260_241_0, i_8_260_311_0, i_8_260_322_0,
    i_8_260_323_0, i_8_260_328_0, i_8_260_364_0, i_8_260_367_0,
    i_8_260_368_0, i_8_260_436_0, i_8_260_439_0, i_8_260_574_0,
    i_8_260_606_0, i_8_260_628_0, i_8_260_633_0, i_8_260_646_0,
    i_8_260_665_0, i_8_260_672_0, i_8_260_674_0, i_8_260_682_0,
    i_8_260_701_0, i_8_260_707_0, i_8_260_709_0, i_8_260_710_0,
    i_8_260_735_0, i_8_260_804_0, i_8_260_823_0, i_8_260_834_0,
    i_8_260_886_0, i_8_260_957_0, i_8_260_979_0, i_8_260_985_0,
    i_8_260_1060_0, i_8_260_1074_0, i_8_260_1105_0, i_8_260_1132_0,
    i_8_260_1158_0, i_8_260_1185_0, i_8_260_1236_0, i_8_260_1239_0,
    i_8_260_1266_0, i_8_260_1284_0, i_8_260_1310_0, i_8_260_1352_0,
    i_8_260_1353_0, i_8_260_1354_0, i_8_260_1357_0, i_8_260_1365_0,
    i_8_260_1374_0, i_8_260_1375_0, i_8_260_1384_0, i_8_260_1405_0,
    i_8_260_1426_0, i_8_260_1429_0, i_8_260_1480_0, i_8_260_1590_0,
    i_8_260_1623_0, i_8_260_1624_0, i_8_260_1636_0, i_8_260_1649_0,
    i_8_260_1671_0, i_8_260_1672_0, i_8_260_1731_0, i_8_260_1749_0,
    i_8_260_1752_0, i_8_260_1770_0, i_8_260_1797_0, i_8_260_1824_0,
    i_8_260_1825_0, i_8_260_1903_0, i_8_260_1905_0, i_8_260_1914_0,
    i_8_260_1942_0, i_8_260_2031_0, i_8_260_2056_0, i_8_260_2082_0,
    i_8_260_2128_0, i_8_260_2136_0, i_8_260_2148_0, i_8_260_2193_0,
    i_8_260_2194_0, i_8_260_2217_0, i_8_260_2230_0, i_8_260_2263_0,
    i_8_260_2269_0, i_8_260_2272_0, i_8_260_2273_0, i_8_260_2274_0,
    i_8_260_2275_0, i_8_260_2276_0, i_8_260_2290_0,
    o_8_260_0_0  );
  input  i_8_260_6_0, i_8_260_14_0, i_8_260_44_0, i_8_260_106_0,
    i_8_260_140_0, i_8_260_196_0, i_8_260_197_0, i_8_260_214_0,
    i_8_260_222_0, i_8_260_228_0, i_8_260_241_0, i_8_260_311_0,
    i_8_260_322_0, i_8_260_323_0, i_8_260_328_0, i_8_260_364_0,
    i_8_260_367_0, i_8_260_368_0, i_8_260_436_0, i_8_260_439_0,
    i_8_260_574_0, i_8_260_606_0, i_8_260_628_0, i_8_260_633_0,
    i_8_260_646_0, i_8_260_665_0, i_8_260_672_0, i_8_260_674_0,
    i_8_260_682_0, i_8_260_701_0, i_8_260_707_0, i_8_260_709_0,
    i_8_260_710_0, i_8_260_735_0, i_8_260_804_0, i_8_260_823_0,
    i_8_260_834_0, i_8_260_886_0, i_8_260_957_0, i_8_260_979_0,
    i_8_260_985_0, i_8_260_1060_0, i_8_260_1074_0, i_8_260_1105_0,
    i_8_260_1132_0, i_8_260_1158_0, i_8_260_1185_0, i_8_260_1236_0,
    i_8_260_1239_0, i_8_260_1266_0, i_8_260_1284_0, i_8_260_1310_0,
    i_8_260_1352_0, i_8_260_1353_0, i_8_260_1354_0, i_8_260_1357_0,
    i_8_260_1365_0, i_8_260_1374_0, i_8_260_1375_0, i_8_260_1384_0,
    i_8_260_1405_0, i_8_260_1426_0, i_8_260_1429_0, i_8_260_1480_0,
    i_8_260_1590_0, i_8_260_1623_0, i_8_260_1624_0, i_8_260_1636_0,
    i_8_260_1649_0, i_8_260_1671_0, i_8_260_1672_0, i_8_260_1731_0,
    i_8_260_1749_0, i_8_260_1752_0, i_8_260_1770_0, i_8_260_1797_0,
    i_8_260_1824_0, i_8_260_1825_0, i_8_260_1903_0, i_8_260_1905_0,
    i_8_260_1914_0, i_8_260_1942_0, i_8_260_2031_0, i_8_260_2056_0,
    i_8_260_2082_0, i_8_260_2128_0, i_8_260_2136_0, i_8_260_2148_0,
    i_8_260_2193_0, i_8_260_2194_0, i_8_260_2217_0, i_8_260_2230_0,
    i_8_260_2263_0, i_8_260_2269_0, i_8_260_2272_0, i_8_260_2273_0,
    i_8_260_2274_0, i_8_260_2275_0, i_8_260_2276_0, i_8_260_2290_0;
  output o_8_260_0_0;
  assign o_8_260_0_0 = 0;
endmodule



// Benchmark "kernel_8_261" written by ABC on Sun Jul 19 10:07:36 2020

module kernel_8_261 ( 
    i_8_261_14_0, i_8_261_50_0, i_8_261_55_0, i_8_261_58_0, i_8_261_141_0,
    i_8_261_143_0, i_8_261_157_0, i_8_261_159_0, i_8_261_187_0,
    i_8_261_259_0, i_8_261_310_0, i_8_261_373_0, i_8_261_378_0,
    i_8_261_429_0, i_8_261_437_0, i_8_261_442_0, i_8_261_445_0,
    i_8_261_474_0, i_8_261_481_0, i_8_261_526_0, i_8_261_582_0,
    i_8_261_596_0, i_8_261_601_0, i_8_261_607_0, i_8_261_627_0,
    i_8_261_691_0, i_8_261_693_0, i_8_261_710_0, i_8_261_714_0,
    i_8_261_717_0, i_8_261_760_0, i_8_261_778_0, i_8_261_818_0,
    i_8_261_884_0, i_8_261_913_0, i_8_261_941_0, i_8_261_956_0,
    i_8_261_1012_0, i_8_261_1048_0, i_8_261_1050_0, i_8_261_1056_0,
    i_8_261_1071_0, i_8_261_1088_0, i_8_261_1090_0, i_8_261_1116_0,
    i_8_261_1123_0, i_8_261_1133_0, i_8_261_1189_0, i_8_261_1241_0,
    i_8_261_1264_0, i_8_261_1267_0, i_8_261_1273_0, i_8_261_1276_0,
    i_8_261_1287_0, i_8_261_1295_0, i_8_261_1324_0, i_8_261_1326_0,
    i_8_261_1327_0, i_8_261_1335_0, i_8_261_1390_0, i_8_261_1435_0,
    i_8_261_1467_0, i_8_261_1472_0, i_8_261_1507_0, i_8_261_1545_0,
    i_8_261_1588_0, i_8_261_1599_0, i_8_261_1605_0, i_8_261_1629_0,
    i_8_261_1632_0, i_8_261_1653_0, i_8_261_1668_0, i_8_261_1719_0,
    i_8_261_1723_0, i_8_261_1746_0, i_8_261_1772_0, i_8_261_1784_0,
    i_8_261_1790_0, i_8_261_1797_0, i_8_261_1830_0, i_8_261_1831_0,
    i_8_261_1839_0, i_8_261_1877_0, i_8_261_1900_0, i_8_261_1917_0,
    i_8_261_1918_0, i_8_261_1919_0, i_8_261_1930_0, i_8_261_1939_0,
    i_8_261_1989_0, i_8_261_2028_0, i_8_261_2101_0, i_8_261_2112_0,
    i_8_261_2133_0, i_8_261_2185_0, i_8_261_2211_0, i_8_261_2241_0,
    i_8_261_2245_0, i_8_261_2270_0, i_8_261_2293_0,
    o_8_261_0_0  );
  input  i_8_261_14_0, i_8_261_50_0, i_8_261_55_0, i_8_261_58_0,
    i_8_261_141_0, i_8_261_143_0, i_8_261_157_0, i_8_261_159_0,
    i_8_261_187_0, i_8_261_259_0, i_8_261_310_0, i_8_261_373_0,
    i_8_261_378_0, i_8_261_429_0, i_8_261_437_0, i_8_261_442_0,
    i_8_261_445_0, i_8_261_474_0, i_8_261_481_0, i_8_261_526_0,
    i_8_261_582_0, i_8_261_596_0, i_8_261_601_0, i_8_261_607_0,
    i_8_261_627_0, i_8_261_691_0, i_8_261_693_0, i_8_261_710_0,
    i_8_261_714_0, i_8_261_717_0, i_8_261_760_0, i_8_261_778_0,
    i_8_261_818_0, i_8_261_884_0, i_8_261_913_0, i_8_261_941_0,
    i_8_261_956_0, i_8_261_1012_0, i_8_261_1048_0, i_8_261_1050_0,
    i_8_261_1056_0, i_8_261_1071_0, i_8_261_1088_0, i_8_261_1090_0,
    i_8_261_1116_0, i_8_261_1123_0, i_8_261_1133_0, i_8_261_1189_0,
    i_8_261_1241_0, i_8_261_1264_0, i_8_261_1267_0, i_8_261_1273_0,
    i_8_261_1276_0, i_8_261_1287_0, i_8_261_1295_0, i_8_261_1324_0,
    i_8_261_1326_0, i_8_261_1327_0, i_8_261_1335_0, i_8_261_1390_0,
    i_8_261_1435_0, i_8_261_1467_0, i_8_261_1472_0, i_8_261_1507_0,
    i_8_261_1545_0, i_8_261_1588_0, i_8_261_1599_0, i_8_261_1605_0,
    i_8_261_1629_0, i_8_261_1632_0, i_8_261_1653_0, i_8_261_1668_0,
    i_8_261_1719_0, i_8_261_1723_0, i_8_261_1746_0, i_8_261_1772_0,
    i_8_261_1784_0, i_8_261_1790_0, i_8_261_1797_0, i_8_261_1830_0,
    i_8_261_1831_0, i_8_261_1839_0, i_8_261_1877_0, i_8_261_1900_0,
    i_8_261_1917_0, i_8_261_1918_0, i_8_261_1919_0, i_8_261_1930_0,
    i_8_261_1939_0, i_8_261_1989_0, i_8_261_2028_0, i_8_261_2101_0,
    i_8_261_2112_0, i_8_261_2133_0, i_8_261_2185_0, i_8_261_2211_0,
    i_8_261_2241_0, i_8_261_2245_0, i_8_261_2270_0, i_8_261_2293_0;
  output o_8_261_0_0;
  assign o_8_261_0_0 = 0;
endmodule



// Benchmark "kernel_8_262" written by ABC on Sun Jul 19 10:07:38 2020

module kernel_8_262 ( 
    i_8_262_31_0, i_8_262_49_0, i_8_262_54_0, i_8_262_56_0, i_8_262_81_0,
    i_8_262_85_0, i_8_262_86_0, i_8_262_103_0, i_8_262_219_0,
    i_8_262_229_0, i_8_262_237_0, i_8_262_297_0, i_8_262_300_0,
    i_8_262_301_0, i_8_262_346_0, i_8_262_361_0, i_8_262_362_0,
    i_8_262_366_0, i_8_262_442_0, i_8_262_486_0, i_8_262_522_0,
    i_8_262_523_0, i_8_262_524_0, i_8_262_580_0, i_8_262_585_0,
    i_8_262_586_0, i_8_262_590_0, i_8_262_603_0, i_8_262_622_0,
    i_8_262_630_0, i_8_262_657_0, i_8_262_662_0, i_8_262_667_0,
    i_8_262_675_0, i_8_262_676_0, i_8_262_677_0, i_8_262_833_0,
    i_8_262_839_0, i_8_262_850_0, i_8_262_876_0, i_8_262_877_0,
    i_8_262_1048_0, i_8_262_1071_0, i_8_262_1072_0, i_8_262_1108_0,
    i_8_262_1189_0, i_8_262_1190_0, i_8_262_1225_0, i_8_262_1263_0,
    i_8_262_1264_0, i_8_262_1270_0, i_8_262_1271_0, i_8_262_1282_0,
    i_8_262_1283_0, i_8_262_1286_0, i_8_262_1296_0, i_8_262_1333_0,
    i_8_262_1334_0, i_8_262_1337_0, i_8_262_1353_0, i_8_262_1408_0,
    i_8_262_1409_0, i_8_262_1534_0, i_8_262_1550_0, i_8_262_1561_0,
    i_8_262_1620_0, i_8_262_1629_0, i_8_262_1631_0, i_8_262_1638_0,
    i_8_262_1648_0, i_8_262_1680_0, i_8_262_1728_0, i_8_262_1732_0,
    i_8_262_1768_0, i_8_262_1773_0, i_8_262_1774_0, i_8_262_1782_0,
    i_8_262_1784_0, i_8_262_1811_0, i_8_262_1818_0, i_8_262_1819_0,
    i_8_262_1830_0, i_8_262_1848_0, i_8_262_1855_0, i_8_262_1856_0,
    i_8_262_1888_0, i_8_262_1903_0, i_8_262_1904_0, i_8_262_1962_0,
    i_8_262_1982_0, i_8_262_1985_0, i_8_262_2037_0, i_8_262_2038_0,
    i_8_262_2133_0, i_8_262_2134_0, i_8_262_2147_0, i_8_262_2155_0,
    i_8_262_2245_0, i_8_262_2270_0, i_8_262_2293_0,
    o_8_262_0_0  );
  input  i_8_262_31_0, i_8_262_49_0, i_8_262_54_0, i_8_262_56_0,
    i_8_262_81_0, i_8_262_85_0, i_8_262_86_0, i_8_262_103_0, i_8_262_219_0,
    i_8_262_229_0, i_8_262_237_0, i_8_262_297_0, i_8_262_300_0,
    i_8_262_301_0, i_8_262_346_0, i_8_262_361_0, i_8_262_362_0,
    i_8_262_366_0, i_8_262_442_0, i_8_262_486_0, i_8_262_522_0,
    i_8_262_523_0, i_8_262_524_0, i_8_262_580_0, i_8_262_585_0,
    i_8_262_586_0, i_8_262_590_0, i_8_262_603_0, i_8_262_622_0,
    i_8_262_630_0, i_8_262_657_0, i_8_262_662_0, i_8_262_667_0,
    i_8_262_675_0, i_8_262_676_0, i_8_262_677_0, i_8_262_833_0,
    i_8_262_839_0, i_8_262_850_0, i_8_262_876_0, i_8_262_877_0,
    i_8_262_1048_0, i_8_262_1071_0, i_8_262_1072_0, i_8_262_1108_0,
    i_8_262_1189_0, i_8_262_1190_0, i_8_262_1225_0, i_8_262_1263_0,
    i_8_262_1264_0, i_8_262_1270_0, i_8_262_1271_0, i_8_262_1282_0,
    i_8_262_1283_0, i_8_262_1286_0, i_8_262_1296_0, i_8_262_1333_0,
    i_8_262_1334_0, i_8_262_1337_0, i_8_262_1353_0, i_8_262_1408_0,
    i_8_262_1409_0, i_8_262_1534_0, i_8_262_1550_0, i_8_262_1561_0,
    i_8_262_1620_0, i_8_262_1629_0, i_8_262_1631_0, i_8_262_1638_0,
    i_8_262_1648_0, i_8_262_1680_0, i_8_262_1728_0, i_8_262_1732_0,
    i_8_262_1768_0, i_8_262_1773_0, i_8_262_1774_0, i_8_262_1782_0,
    i_8_262_1784_0, i_8_262_1811_0, i_8_262_1818_0, i_8_262_1819_0,
    i_8_262_1830_0, i_8_262_1848_0, i_8_262_1855_0, i_8_262_1856_0,
    i_8_262_1888_0, i_8_262_1903_0, i_8_262_1904_0, i_8_262_1962_0,
    i_8_262_1982_0, i_8_262_1985_0, i_8_262_2037_0, i_8_262_2038_0,
    i_8_262_2133_0, i_8_262_2134_0, i_8_262_2147_0, i_8_262_2155_0,
    i_8_262_2245_0, i_8_262_2270_0, i_8_262_2293_0;
  output o_8_262_0_0;
  assign o_8_262_0_0 = ~((~i_8_262_31_0 & ((~i_8_262_49_0 & ~i_8_262_586_0 & ~i_8_262_590_0 & ~i_8_262_676_0 & ~i_8_262_1264_0 & ~i_8_262_1296_0 & ~i_8_262_1631_0 & ~i_8_262_1811_0 & i_8_262_1818_0 & ~i_8_262_1856_0) | (~i_8_262_229_0 & ~i_8_262_297_0 & i_8_262_346_0 & ~i_8_262_486_0 & ~i_8_262_585_0 & i_8_262_850_0 & i_8_262_1264_0 & i_8_262_2147_0))) | (~i_8_262_1353_0 & ((~i_8_262_54_0 & ~i_8_262_1282_0 & ((~i_8_262_523_0 & ~i_8_262_524_0 & ~i_8_262_590_0 & ~i_8_262_662_0 & ~i_8_262_850_0 & ~i_8_262_1283_0 & ~i_8_262_1629_0) | (~i_8_262_300_0 & ~i_8_262_677_0 & ~i_8_262_876_0 & ~i_8_262_1225_0 & ~i_8_262_1784_0 & ~i_8_262_1903_0 & ~i_8_262_2155_0 & ~i_8_262_2293_0))) | (~i_8_262_366_0 & i_8_262_523_0 & ~i_8_262_676_0 & ~i_8_262_1048_0 & ~i_8_262_1732_0 & ~i_8_262_1811_0 & ~i_8_262_1819_0))) | (~i_8_262_229_0 & ((~i_8_262_442_0 & i_8_262_1225_0 & ~i_8_262_1334_0 & ~i_8_262_1409_0 & ~i_8_262_1631_0 & ~i_8_262_1648_0 & i_8_262_1768_0 & ~i_8_262_1773_0 & ~i_8_262_1830_0) | (~i_8_262_630_0 & i_8_262_833_0 & ~i_8_262_1190_0 & ~i_8_262_1534_0 & ~i_8_262_1550_0 & ~i_8_262_1774_0 & ~i_8_262_1962_0))) | (~i_8_262_300_0 & ((~i_8_262_585_0 & ~i_8_262_590_0 & ~i_8_262_675_0 & ~i_8_262_677_0 & ~i_8_262_876_0 & ~i_8_262_1333_0 & ~i_8_262_1337_0) | (~i_8_262_219_0 & ~i_8_262_301_0 & ~i_8_262_1108_0 & ~i_8_262_1190_0 & ~i_8_262_1264_0 & ~i_8_262_1334_0 & ~i_8_262_1629_0 & ~i_8_262_1631_0 & ~i_8_262_2155_0))) | (~i_8_262_219_0 & ((~i_8_262_603_0 & ~i_8_262_677_0 & ~i_8_262_1048_0 & ~i_8_262_1286_0 & ~i_8_262_1333_0 & ~i_8_262_1334_0 & ~i_8_262_1811_0 & ~i_8_262_1830_0 & ~i_8_262_1962_0) | (~i_8_262_49_0 & ~i_8_262_662_0 & i_8_262_667_0 & ~i_8_262_675_0 & ~i_8_262_1409_0 & ~i_8_262_2038_0))) | (~i_8_262_1337_0 & ((~i_8_262_301_0 & ~i_8_262_657_0 & ((~i_8_262_366_0 & ~i_8_262_676_0 & i_8_262_1048_0 & ~i_8_262_1631_0 & ~i_8_262_1728_0 & ~i_8_262_1819_0) | (~i_8_262_1263_0 & ~i_8_262_1286_0 & ~i_8_262_1409_0 & ~i_8_262_1629_0 & ~i_8_262_1784_0 & ~i_8_262_1982_0))) | (~i_8_262_585_0 & ~i_8_262_586_0 & ~i_8_262_675_0 & ~i_8_262_1333_0 & ~i_8_262_1334_0 & i_8_262_1409_0) | (~i_8_262_49_0 & i_8_262_86_0 & ~i_8_262_297_0 & ~i_8_262_2245_0) | (i_8_262_522_0 & ~i_8_262_676_0 & ~i_8_262_1550_0 & ~i_8_262_2293_0))) | (~i_8_262_590_0 & ((i_8_262_49_0 & ~i_8_262_1286_0 & ~i_8_262_1629_0 & ~i_8_262_1768_0 & ~i_8_262_1774_0) | (~i_8_262_677_0 & ~i_8_262_1263_0 & ~i_8_262_1334_0 & ~i_8_262_1773_0 & ~i_8_262_1818_0))) | (~i_8_262_603_0 & ((~i_8_262_676_0 & i_8_262_1071_0 & ~i_8_262_1680_0 & ~i_8_262_1768_0) | (~i_8_262_586_0 & ~i_8_262_675_0 & ~i_8_262_49_0 & ~i_8_262_362_0 & ~i_8_262_677_0 & ~i_8_262_839_0 & ~i_8_262_850_0 & ~i_8_262_1408_0 & ~i_8_262_1888_0))) | (~i_8_262_362_0 & ((~i_8_262_586_0 & ((~i_8_262_662_0 & i_8_262_877_0 & ~i_8_262_1409_0 & ~i_8_262_1773_0 & ~i_8_262_1774_0 & ~i_8_262_1782_0 & ~i_8_262_1888_0) | (~i_8_262_675_0 & ~i_8_262_1190_0 & ~i_8_262_1225_0 & ~i_8_262_1334_0 & i_8_262_2147_0))) | (~i_8_262_297_0 & i_8_262_301_0 & ~i_8_262_486_0 & ~i_8_262_876_0 & ~i_8_262_1108_0 & ~i_8_262_1334_0 & ~i_8_262_1561_0))) | (~i_8_262_297_0 & ((~i_8_262_49_0 & ~i_8_262_839_0 & ~i_8_262_1264_0 & ~i_8_262_1631_0 & ~i_8_262_1782_0 & ~i_8_262_1985_0) | (~i_8_262_675_0 & ~i_8_262_1550_0 & i_8_262_1888_0 & i_8_262_2245_0))) | (~i_8_262_49_0 & ((~i_8_262_662_0 & ~i_8_262_676_0 & i_8_262_1190_0) | (~i_8_262_675_0 & ~i_8_262_1334_0 & ~i_8_262_1561_0 & ~i_8_262_1768_0 & ~i_8_262_1818_0 & ~i_8_262_1985_0 & ~i_8_262_2293_0))) | (~i_8_262_675_0 & ((~i_8_262_833_0 & i_8_262_1271_0 & ~i_8_262_1768_0) | (~i_8_262_103_0 & ~i_8_262_676_0 & ~i_8_262_1283_0 & ~i_8_262_1286_0 & ~i_8_262_1773_0 & ~i_8_262_1818_0 & ~i_8_262_1819_0 & ~i_8_262_1982_0))) | (~i_8_262_1629_0 & ~i_8_262_1768_0 & ~i_8_262_2134_0 & ((~i_8_262_662_0 & i_8_262_1408_0 & ~i_8_262_1982_0) | (~i_8_262_1631_0 & i_8_262_1818_0 & ~i_8_262_1985_0 & ~i_8_262_2133_0))) | (i_8_262_486_0 & ~i_8_262_1333_0 & i_8_262_1648_0 & i_8_262_1728_0) | (~i_8_262_677_0 & i_8_262_1409_0 & i_8_262_1620_0 & ~i_8_262_1773_0) | (~i_8_262_56_0 & i_8_262_219_0 & i_8_262_523_0 & ~i_8_262_657_0 & ~i_8_262_676_0 & ~i_8_262_2155_0));
endmodule



// Benchmark "kernel_8_263" written by ABC on Sun Jul 19 10:07:39 2020

module kernel_8_263 ( 
    i_8_263_20_0, i_8_263_36_0, i_8_263_135_0, i_8_263_253_0,
    i_8_263_280_0, i_8_263_297_0, i_8_263_364_0, i_8_263_396_0,
    i_8_263_432_0, i_8_263_480_0, i_8_263_530_0, i_8_263_544_0,
    i_8_263_585_0, i_8_263_595_0, i_8_263_615_0, i_8_263_621_0,
    i_8_263_630_0, i_8_263_636_0, i_8_263_657_0, i_8_263_666_0,
    i_8_263_667_0, i_8_263_675_0, i_8_263_682_0, i_8_263_703_0,
    i_8_263_720_0, i_8_263_721_0, i_8_263_724_0, i_8_263_765_0,
    i_8_263_801_0, i_8_263_804_0, i_8_263_822_0, i_8_263_847_0,
    i_8_263_866_0, i_8_263_868_0, i_8_263_879_0, i_8_263_892_0,
    i_8_263_955_0, i_8_263_965_0, i_8_263_967_0, i_8_263_985_0,
    i_8_263_991_0, i_8_263_1050_0, i_8_263_1071_0, i_8_263_1111_0,
    i_8_263_1188_0, i_8_263_1189_0, i_8_263_1233_0, i_8_263_1251_0,
    i_8_263_1261_0, i_8_263_1292_0, i_8_263_1300_0, i_8_263_1351_0,
    i_8_263_1353_0, i_8_263_1359_0, i_8_263_1365_0, i_8_263_1366_0,
    i_8_263_1367_0, i_8_263_1374_0, i_8_263_1382_0, i_8_263_1450_0,
    i_8_263_1467_0, i_8_263_1531_0, i_8_263_1536_0, i_8_263_1537_0,
    i_8_263_1549_0, i_8_263_1559_0, i_8_263_1565_0, i_8_263_1575_0,
    i_8_263_1584_0, i_8_263_1586_0, i_8_263_1588_0, i_8_263_1622_0,
    i_8_263_1624_0, i_8_263_1629_0, i_8_263_1639_0, i_8_263_1674_0,
    i_8_263_1680_0, i_8_263_1681_0, i_8_263_1697_0, i_8_263_1747_0,
    i_8_263_1750_0, i_8_263_1756_0, i_8_263_1762_0, i_8_263_1815_0,
    i_8_263_1837_0, i_8_263_1908_0, i_8_263_1944_0, i_8_263_1947_0,
    i_8_263_1982_0, i_8_263_2004_0, i_8_263_2107_0, i_8_263_2116_0,
    i_8_263_2125_0, i_8_263_2139_0, i_8_263_2147_0, i_8_263_2187_0,
    i_8_263_2188_0, i_8_263_2191_0, i_8_263_2255_0, i_8_263_2259_0,
    o_8_263_0_0  );
  input  i_8_263_20_0, i_8_263_36_0, i_8_263_135_0, i_8_263_253_0,
    i_8_263_280_0, i_8_263_297_0, i_8_263_364_0, i_8_263_396_0,
    i_8_263_432_0, i_8_263_480_0, i_8_263_530_0, i_8_263_544_0,
    i_8_263_585_0, i_8_263_595_0, i_8_263_615_0, i_8_263_621_0,
    i_8_263_630_0, i_8_263_636_0, i_8_263_657_0, i_8_263_666_0,
    i_8_263_667_0, i_8_263_675_0, i_8_263_682_0, i_8_263_703_0,
    i_8_263_720_0, i_8_263_721_0, i_8_263_724_0, i_8_263_765_0,
    i_8_263_801_0, i_8_263_804_0, i_8_263_822_0, i_8_263_847_0,
    i_8_263_866_0, i_8_263_868_0, i_8_263_879_0, i_8_263_892_0,
    i_8_263_955_0, i_8_263_965_0, i_8_263_967_0, i_8_263_985_0,
    i_8_263_991_0, i_8_263_1050_0, i_8_263_1071_0, i_8_263_1111_0,
    i_8_263_1188_0, i_8_263_1189_0, i_8_263_1233_0, i_8_263_1251_0,
    i_8_263_1261_0, i_8_263_1292_0, i_8_263_1300_0, i_8_263_1351_0,
    i_8_263_1353_0, i_8_263_1359_0, i_8_263_1365_0, i_8_263_1366_0,
    i_8_263_1367_0, i_8_263_1374_0, i_8_263_1382_0, i_8_263_1450_0,
    i_8_263_1467_0, i_8_263_1531_0, i_8_263_1536_0, i_8_263_1537_0,
    i_8_263_1549_0, i_8_263_1559_0, i_8_263_1565_0, i_8_263_1575_0,
    i_8_263_1584_0, i_8_263_1586_0, i_8_263_1588_0, i_8_263_1622_0,
    i_8_263_1624_0, i_8_263_1629_0, i_8_263_1639_0, i_8_263_1674_0,
    i_8_263_1680_0, i_8_263_1681_0, i_8_263_1697_0, i_8_263_1747_0,
    i_8_263_1750_0, i_8_263_1756_0, i_8_263_1762_0, i_8_263_1815_0,
    i_8_263_1837_0, i_8_263_1908_0, i_8_263_1944_0, i_8_263_1947_0,
    i_8_263_1982_0, i_8_263_2004_0, i_8_263_2107_0, i_8_263_2116_0,
    i_8_263_2125_0, i_8_263_2139_0, i_8_263_2147_0, i_8_263_2187_0,
    i_8_263_2188_0, i_8_263_2191_0, i_8_263_2255_0, i_8_263_2259_0;
  output o_8_263_0_0;
  assign o_8_263_0_0 = 0;
endmodule



// Benchmark "kernel_8_264" written by ABC on Sun Jul 19 10:07:40 2020

module kernel_8_264 ( 
    i_8_264_6_0, i_8_264_41_0, i_8_264_60_0, i_8_264_115_0, i_8_264_118_0,
    i_8_264_179_0, i_8_264_202_0, i_8_264_256_0, i_8_264_258_0,
    i_8_264_292_0, i_8_264_363_0, i_8_264_364_0, i_8_264_381_0,
    i_8_264_392_0, i_8_264_401_0, i_8_264_419_0, i_8_264_422_0,
    i_8_264_462_0, i_8_264_475_0, i_8_264_509_0, i_8_264_525_0,
    i_8_264_529_0, i_8_264_572_0, i_8_264_581_0, i_8_264_589_0,
    i_8_264_592_0, i_8_264_606_0, i_8_264_607_0, i_8_264_618_0,
    i_8_264_633_0, i_8_264_708_0, i_8_264_714_0, i_8_264_769_0,
    i_8_264_795_0, i_8_264_796_0, i_8_264_818_0, i_8_264_824_0,
    i_8_264_835_0, i_8_264_858_0, i_8_264_895_0, i_8_264_896_0,
    i_8_264_897_0, i_8_264_992_0, i_8_264_1040_0, i_8_264_1131_0,
    i_8_264_1132_0, i_8_264_1192_0, i_8_264_1202_0, i_8_264_1267_0,
    i_8_264_1278_0, i_8_264_1282_0, i_8_264_1286_0, i_8_264_1319_0,
    i_8_264_1328_0, i_8_264_1334_0, i_8_264_1382_0, i_8_264_1407_0,
    i_8_264_1427_0, i_8_264_1443_0, i_8_264_1448_0, i_8_264_1455_0,
    i_8_264_1481_0, i_8_264_1489_0, i_8_264_1490_0, i_8_264_1508_0,
    i_8_264_1550_0, i_8_264_1553_0, i_8_264_1578_0, i_8_264_1589_0,
    i_8_264_1597_0, i_8_264_1614_0, i_8_264_1632_0, i_8_264_1697_0,
    i_8_264_1705_0, i_8_264_1706_0, i_8_264_1751_0, i_8_264_1760_0,
    i_8_264_1762_0, i_8_264_1807_0, i_8_264_1808_0, i_8_264_1837_0,
    i_8_264_1841_0, i_8_264_1885_0, i_8_264_1888_0, i_8_264_1963_0,
    i_8_264_1994_0, i_8_264_2002_0, i_8_264_2011_0, i_8_264_2090_0,
    i_8_264_2111_0, i_8_264_2113_0, i_8_264_2127_0, i_8_264_2176_0,
    i_8_264_2177_0, i_8_264_2184_0, i_8_264_2188_0, i_8_264_2211_0,
    i_8_264_2262_0, i_8_264_2273_0, i_8_264_2291_0,
    o_8_264_0_0  );
  input  i_8_264_6_0, i_8_264_41_0, i_8_264_60_0, i_8_264_115_0,
    i_8_264_118_0, i_8_264_179_0, i_8_264_202_0, i_8_264_256_0,
    i_8_264_258_0, i_8_264_292_0, i_8_264_363_0, i_8_264_364_0,
    i_8_264_381_0, i_8_264_392_0, i_8_264_401_0, i_8_264_419_0,
    i_8_264_422_0, i_8_264_462_0, i_8_264_475_0, i_8_264_509_0,
    i_8_264_525_0, i_8_264_529_0, i_8_264_572_0, i_8_264_581_0,
    i_8_264_589_0, i_8_264_592_0, i_8_264_606_0, i_8_264_607_0,
    i_8_264_618_0, i_8_264_633_0, i_8_264_708_0, i_8_264_714_0,
    i_8_264_769_0, i_8_264_795_0, i_8_264_796_0, i_8_264_818_0,
    i_8_264_824_0, i_8_264_835_0, i_8_264_858_0, i_8_264_895_0,
    i_8_264_896_0, i_8_264_897_0, i_8_264_992_0, i_8_264_1040_0,
    i_8_264_1131_0, i_8_264_1132_0, i_8_264_1192_0, i_8_264_1202_0,
    i_8_264_1267_0, i_8_264_1278_0, i_8_264_1282_0, i_8_264_1286_0,
    i_8_264_1319_0, i_8_264_1328_0, i_8_264_1334_0, i_8_264_1382_0,
    i_8_264_1407_0, i_8_264_1427_0, i_8_264_1443_0, i_8_264_1448_0,
    i_8_264_1455_0, i_8_264_1481_0, i_8_264_1489_0, i_8_264_1490_0,
    i_8_264_1508_0, i_8_264_1550_0, i_8_264_1553_0, i_8_264_1578_0,
    i_8_264_1589_0, i_8_264_1597_0, i_8_264_1614_0, i_8_264_1632_0,
    i_8_264_1697_0, i_8_264_1705_0, i_8_264_1706_0, i_8_264_1751_0,
    i_8_264_1760_0, i_8_264_1762_0, i_8_264_1807_0, i_8_264_1808_0,
    i_8_264_1837_0, i_8_264_1841_0, i_8_264_1885_0, i_8_264_1888_0,
    i_8_264_1963_0, i_8_264_1994_0, i_8_264_2002_0, i_8_264_2011_0,
    i_8_264_2090_0, i_8_264_2111_0, i_8_264_2113_0, i_8_264_2127_0,
    i_8_264_2176_0, i_8_264_2177_0, i_8_264_2184_0, i_8_264_2188_0,
    i_8_264_2211_0, i_8_264_2262_0, i_8_264_2273_0, i_8_264_2291_0;
  output o_8_264_0_0;
  assign o_8_264_0_0 = 0;
endmodule



// Benchmark "kernel_8_265" written by ABC on Sun Jul 19 10:07:41 2020

module kernel_8_265 ( 
    i_8_265_1_0, i_8_265_2_0, i_8_265_19_0, i_8_265_31_0, i_8_265_60_0,
    i_8_265_115_0, i_8_265_116_0, i_8_265_198_0, i_8_265_266_0,
    i_8_265_269_0, i_8_265_284_0, i_8_265_293_0, i_8_265_346_0,
    i_8_265_349_0, i_8_265_366_0, i_8_265_378_0, i_8_265_380_0,
    i_8_265_385_0, i_8_265_427_0, i_8_265_437_0, i_8_265_445_0,
    i_8_265_446_0, i_8_265_463_0, i_8_265_464_0, i_8_265_488_0,
    i_8_265_492_0, i_8_265_556_0, i_8_265_572_0, i_8_265_586_0,
    i_8_265_590_0, i_8_265_599_0, i_8_265_614_0, i_8_265_649_0,
    i_8_265_658_0, i_8_265_660_0, i_8_265_665_0, i_8_265_673_0,
    i_8_265_674_0, i_8_265_716_0, i_8_265_718_0, i_8_265_725_0,
    i_8_265_735_0, i_8_265_782_0, i_8_265_796_0, i_8_265_827_0,
    i_8_265_841_0, i_8_265_956_0, i_8_265_976_0, i_8_265_997_0,
    i_8_265_998_0, i_8_265_1004_0, i_8_265_1007_0, i_8_265_1039_0,
    i_8_265_1058_0, i_8_265_1074_0, i_8_265_1114_0, i_8_265_1130_0,
    i_8_265_1211_0, i_8_265_1237_0, i_8_265_1259_0, i_8_265_1274_0,
    i_8_265_1281_0, i_8_265_1302_0, i_8_265_1355_0, i_8_265_1437_0,
    i_8_265_1525_0, i_8_265_1542_0, i_8_265_1543_0, i_8_265_1544_0,
    i_8_265_1546_0, i_8_265_1547_0, i_8_265_1589_0, i_8_265_1592_0,
    i_8_265_1598_0, i_8_265_1618_0, i_8_265_1634_0, i_8_265_1655_0,
    i_8_265_1669_0, i_8_265_1677_0, i_8_265_1699_0, i_8_265_1714_0,
    i_8_265_1723_0, i_8_265_1724_0, i_8_265_1730_0, i_8_265_1753_0,
    i_8_265_1780_0, i_8_265_1919_0, i_8_265_1922_0, i_8_265_1967_0,
    i_8_265_1970_0, i_8_265_2114_0, i_8_265_2120_0, i_8_265_2129_0,
    i_8_265_2149_0, i_8_265_2192_0, i_8_265_2195_0, i_8_265_2242_0,
    i_8_265_2263_0, i_8_265_2275_0, i_8_265_2294_0,
    o_8_265_0_0  );
  input  i_8_265_1_0, i_8_265_2_0, i_8_265_19_0, i_8_265_31_0,
    i_8_265_60_0, i_8_265_115_0, i_8_265_116_0, i_8_265_198_0,
    i_8_265_266_0, i_8_265_269_0, i_8_265_284_0, i_8_265_293_0,
    i_8_265_346_0, i_8_265_349_0, i_8_265_366_0, i_8_265_378_0,
    i_8_265_380_0, i_8_265_385_0, i_8_265_427_0, i_8_265_437_0,
    i_8_265_445_0, i_8_265_446_0, i_8_265_463_0, i_8_265_464_0,
    i_8_265_488_0, i_8_265_492_0, i_8_265_556_0, i_8_265_572_0,
    i_8_265_586_0, i_8_265_590_0, i_8_265_599_0, i_8_265_614_0,
    i_8_265_649_0, i_8_265_658_0, i_8_265_660_0, i_8_265_665_0,
    i_8_265_673_0, i_8_265_674_0, i_8_265_716_0, i_8_265_718_0,
    i_8_265_725_0, i_8_265_735_0, i_8_265_782_0, i_8_265_796_0,
    i_8_265_827_0, i_8_265_841_0, i_8_265_956_0, i_8_265_976_0,
    i_8_265_997_0, i_8_265_998_0, i_8_265_1004_0, i_8_265_1007_0,
    i_8_265_1039_0, i_8_265_1058_0, i_8_265_1074_0, i_8_265_1114_0,
    i_8_265_1130_0, i_8_265_1211_0, i_8_265_1237_0, i_8_265_1259_0,
    i_8_265_1274_0, i_8_265_1281_0, i_8_265_1302_0, i_8_265_1355_0,
    i_8_265_1437_0, i_8_265_1525_0, i_8_265_1542_0, i_8_265_1543_0,
    i_8_265_1544_0, i_8_265_1546_0, i_8_265_1547_0, i_8_265_1589_0,
    i_8_265_1592_0, i_8_265_1598_0, i_8_265_1618_0, i_8_265_1634_0,
    i_8_265_1655_0, i_8_265_1669_0, i_8_265_1677_0, i_8_265_1699_0,
    i_8_265_1714_0, i_8_265_1723_0, i_8_265_1724_0, i_8_265_1730_0,
    i_8_265_1753_0, i_8_265_1780_0, i_8_265_1919_0, i_8_265_1922_0,
    i_8_265_1967_0, i_8_265_1970_0, i_8_265_2114_0, i_8_265_2120_0,
    i_8_265_2129_0, i_8_265_2149_0, i_8_265_2192_0, i_8_265_2195_0,
    i_8_265_2242_0, i_8_265_2263_0, i_8_265_2275_0, i_8_265_2294_0;
  output o_8_265_0_0;
  assign o_8_265_0_0 = ~((~i_8_265_266_0 & ((~i_8_265_293_0 & ~i_8_265_1058_0 & ~i_8_265_1274_0 & ~i_8_265_1437_0 & ~i_8_265_1598_0 & ~i_8_265_2114_0) | (~i_8_265_349_0 & ~i_8_265_782_0 & ~i_8_265_1543_0 & ~i_8_265_1547_0 & ~i_8_265_1618_0 & ~i_8_265_2195_0))) | (~i_8_265_464_0 & ((~i_8_265_599_0 & ~i_8_265_718_0 & ~i_8_265_956_0 & ~i_8_265_1259_0) | (~i_8_265_427_0 & ~i_8_265_673_0 & ~i_8_265_827_0 & ~i_8_265_2192_0))) | (~i_8_265_1259_0 & ((~i_8_265_1543_0 & ~i_8_265_1730_0 & ~i_8_265_1967_0 & ~i_8_265_2192_0) | (~i_8_265_2_0 & ~i_8_265_590_0 & ~i_8_265_673_0 & ~i_8_265_998_0 & ~i_8_265_1074_0 & ~i_8_265_2242_0))) | (~i_8_265_1074_0 & ((~i_8_265_366_0 & ~i_8_265_586_0 & ~i_8_265_1058_0 & ~i_8_265_1730_0 & i_8_265_1753_0 & ~i_8_265_2114_0 & ~i_8_265_2129_0) | (~i_8_265_346_0 & ~i_8_265_735_0 & ~i_8_265_956_0 & ~i_8_265_1274_0 & ~i_8_265_1753_0 & ~i_8_265_2195_0 & ~i_8_265_2242_0))) | (~i_8_265_2114_0 & ((~i_8_265_1007_0 & ~i_8_265_1355_0 & i_8_265_1437_0 & ~i_8_265_1592_0 & ~i_8_265_2120_0) | (~i_8_265_463_0 & ~i_8_265_556_0 & i_8_265_782_0 & ~i_8_265_1281_0 & ~i_8_265_1546_0 & ~i_8_265_1547_0 & ~i_8_265_1699_0 & ~i_8_265_2275_0))) | (~i_8_265_2120_0 & ((~i_8_265_614_0 & ~i_8_265_1004_0 & ~i_8_265_1542_0 & ~i_8_265_1724_0 & ~i_8_265_1780_0 & ~i_8_265_2129_0 & ~i_8_265_2192_0) | (~i_8_265_674_0 & ~i_8_265_716_0 & ~i_8_265_2275_0))) | (i_8_265_445_0 & i_8_265_976_0 & ~i_8_265_2129_0) | i_8_265_1525_0 | (~i_8_265_293_0 & ~i_8_265_437_0 & ~i_8_265_827_0 & ~i_8_265_1598_0));
endmodule



// Benchmark "kernel_8_266" written by ABC on Sun Jul 19 10:07:42 2020

module kernel_8_266 ( 
    i_8_266_39_0, i_8_266_40_0, i_8_266_49_0, i_8_266_82_0, i_8_266_90_0,
    i_8_266_120_0, i_8_266_192_0, i_8_266_300_0, i_8_266_318_0,
    i_8_266_321_0, i_8_266_322_0, i_8_266_391_0, i_8_266_399_0,
    i_8_266_415_0, i_8_266_418_0, i_8_266_428_0, i_8_266_453_0,
    i_8_266_507_0, i_8_266_532_0, i_8_266_552_0, i_8_266_571_0,
    i_8_266_572_0, i_8_266_574_0, i_8_266_595_0, i_8_266_606_0,
    i_8_266_639_0, i_8_266_651_0, i_8_266_657_0, i_8_266_660_0,
    i_8_266_678_0, i_8_266_706_0, i_8_266_829_0, i_8_266_831_0,
    i_8_266_840_0, i_8_266_925_0, i_8_266_964_0, i_8_266_967_0,
    i_8_266_969_0, i_8_266_972_0, i_8_266_975_0, i_8_266_984_0,
    i_8_266_993_0, i_8_266_1011_0, i_8_266_1039_0, i_8_266_1101_0,
    i_8_266_1104_0, i_8_266_1105_0, i_8_266_1111_0, i_8_266_1228_0,
    i_8_266_1239_0, i_8_266_1245_0, i_8_266_1257_0, i_8_266_1266_0,
    i_8_266_1397_0, i_8_266_1407_0, i_8_266_1435_0, i_8_266_1440_0,
    i_8_266_1452_0, i_8_266_1456_0, i_8_266_1461_0, i_8_266_1462_0,
    i_8_266_1464_0, i_8_266_1470_0, i_8_266_1474_0, i_8_266_1476_0,
    i_8_266_1479_0, i_8_266_1480_0, i_8_266_1488_0, i_8_266_1549_0,
    i_8_266_1551_0, i_8_266_1552_0, i_8_266_1624_0, i_8_266_1659_0,
    i_8_266_1704_0, i_8_266_1705_0, i_8_266_1719_0, i_8_266_1724_0,
    i_8_266_1731_0, i_8_266_1749_0, i_8_266_1767_0, i_8_266_1775_0,
    i_8_266_1779_0, i_8_266_1794_0, i_8_266_1795_0, i_8_266_1801_0,
    i_8_266_1820_0, i_8_266_1836_0, i_8_266_1839_0, i_8_266_1858_0,
    i_8_266_1859_0, i_8_266_1885_0, i_8_266_1911_0, i_8_266_1948_0,
    i_8_266_1956_0, i_8_266_2075_0, i_8_266_2173_0, i_8_266_2190_0,
    i_8_266_2226_0, i_8_266_2258_0, i_8_266_2278_0,
    o_8_266_0_0  );
  input  i_8_266_39_0, i_8_266_40_0, i_8_266_49_0, i_8_266_82_0,
    i_8_266_90_0, i_8_266_120_0, i_8_266_192_0, i_8_266_300_0,
    i_8_266_318_0, i_8_266_321_0, i_8_266_322_0, i_8_266_391_0,
    i_8_266_399_0, i_8_266_415_0, i_8_266_418_0, i_8_266_428_0,
    i_8_266_453_0, i_8_266_507_0, i_8_266_532_0, i_8_266_552_0,
    i_8_266_571_0, i_8_266_572_0, i_8_266_574_0, i_8_266_595_0,
    i_8_266_606_0, i_8_266_639_0, i_8_266_651_0, i_8_266_657_0,
    i_8_266_660_0, i_8_266_678_0, i_8_266_706_0, i_8_266_829_0,
    i_8_266_831_0, i_8_266_840_0, i_8_266_925_0, i_8_266_964_0,
    i_8_266_967_0, i_8_266_969_0, i_8_266_972_0, i_8_266_975_0,
    i_8_266_984_0, i_8_266_993_0, i_8_266_1011_0, i_8_266_1039_0,
    i_8_266_1101_0, i_8_266_1104_0, i_8_266_1105_0, i_8_266_1111_0,
    i_8_266_1228_0, i_8_266_1239_0, i_8_266_1245_0, i_8_266_1257_0,
    i_8_266_1266_0, i_8_266_1397_0, i_8_266_1407_0, i_8_266_1435_0,
    i_8_266_1440_0, i_8_266_1452_0, i_8_266_1456_0, i_8_266_1461_0,
    i_8_266_1462_0, i_8_266_1464_0, i_8_266_1470_0, i_8_266_1474_0,
    i_8_266_1476_0, i_8_266_1479_0, i_8_266_1480_0, i_8_266_1488_0,
    i_8_266_1549_0, i_8_266_1551_0, i_8_266_1552_0, i_8_266_1624_0,
    i_8_266_1659_0, i_8_266_1704_0, i_8_266_1705_0, i_8_266_1719_0,
    i_8_266_1724_0, i_8_266_1731_0, i_8_266_1749_0, i_8_266_1767_0,
    i_8_266_1775_0, i_8_266_1779_0, i_8_266_1794_0, i_8_266_1795_0,
    i_8_266_1801_0, i_8_266_1820_0, i_8_266_1836_0, i_8_266_1839_0,
    i_8_266_1858_0, i_8_266_1859_0, i_8_266_1885_0, i_8_266_1911_0,
    i_8_266_1948_0, i_8_266_1956_0, i_8_266_2075_0, i_8_266_2173_0,
    i_8_266_2190_0, i_8_266_2226_0, i_8_266_2258_0, i_8_266_2278_0;
  output o_8_266_0_0;
  assign o_8_266_0_0 = 0;
endmodule



// Benchmark "kernel_8_267" written by ABC on Sun Jul 19 10:07:43 2020

module kernel_8_267 ( 
    i_8_267_50_0, i_8_267_52_0, i_8_267_58_0, i_8_267_59_0, i_8_267_71_0,
    i_8_267_89_0, i_8_267_97_0, i_8_267_118_0, i_8_267_142_0,
    i_8_267_157_0, i_8_267_160_0, i_8_267_204_0, i_8_267_205_0,
    i_8_267_210_0, i_8_267_212_0, i_8_267_214_0, i_8_267_223_0,
    i_8_267_241_0, i_8_267_244_0, i_8_267_258_0, i_8_267_346_0,
    i_8_267_373_0, i_8_267_419_0, i_8_267_440_0, i_8_267_476_0,
    i_8_267_498_0, i_8_267_499_0, i_8_267_500_0, i_8_267_502_0,
    i_8_267_522_0, i_8_267_588_0, i_8_267_589_0, i_8_267_605_0,
    i_8_267_662_0, i_8_267_715_0, i_8_267_730_0, i_8_267_765_0,
    i_8_267_781_0, i_8_267_784_0, i_8_267_877_0, i_8_267_904_0,
    i_8_267_907_0, i_8_267_925_0, i_8_267_975_0, i_8_267_986_0,
    i_8_267_1027_0, i_8_267_1074_0, i_8_267_1110_0, i_8_267_1186_0,
    i_8_267_1249_0, i_8_267_1250_0, i_8_267_1255_0, i_8_267_1281_0,
    i_8_267_1284_0, i_8_267_1341_0, i_8_267_1342_0, i_8_267_1420_0,
    i_8_267_1426_0, i_8_267_1435_0, i_8_267_1443_0, i_8_267_1470_0,
    i_8_267_1472_0, i_8_267_1492_0, i_8_267_1528_0, i_8_267_1541_0,
    i_8_267_1555_0, i_8_267_1588_0, i_8_267_1589_0, i_8_267_1596_0,
    i_8_267_1597_0, i_8_267_1598_0, i_8_267_1634_0, i_8_267_1647_0,
    i_8_267_1678_0, i_8_267_1699_0, i_8_267_1706_0, i_8_267_1711_0,
    i_8_267_1737_0, i_8_267_1753_0, i_8_267_1782_0, i_8_267_1796_0,
    i_8_267_1818_0, i_8_267_1819_0, i_8_267_1834_0, i_8_267_1844_0,
    i_8_267_1855_0, i_8_267_1867_0, i_8_267_1870_0, i_8_267_1903_0,
    i_8_267_1975_0, i_8_267_2046_0, i_8_267_2109_0, i_8_267_2110_0,
    i_8_267_2111_0, i_8_267_2143_0, i_8_267_2183_0, i_8_267_2190_0,
    i_8_267_2224_0, i_8_267_2244_0, i_8_267_2272_0,
    o_8_267_0_0  );
  input  i_8_267_50_0, i_8_267_52_0, i_8_267_58_0, i_8_267_59_0,
    i_8_267_71_0, i_8_267_89_0, i_8_267_97_0, i_8_267_118_0, i_8_267_142_0,
    i_8_267_157_0, i_8_267_160_0, i_8_267_204_0, i_8_267_205_0,
    i_8_267_210_0, i_8_267_212_0, i_8_267_214_0, i_8_267_223_0,
    i_8_267_241_0, i_8_267_244_0, i_8_267_258_0, i_8_267_346_0,
    i_8_267_373_0, i_8_267_419_0, i_8_267_440_0, i_8_267_476_0,
    i_8_267_498_0, i_8_267_499_0, i_8_267_500_0, i_8_267_502_0,
    i_8_267_522_0, i_8_267_588_0, i_8_267_589_0, i_8_267_605_0,
    i_8_267_662_0, i_8_267_715_0, i_8_267_730_0, i_8_267_765_0,
    i_8_267_781_0, i_8_267_784_0, i_8_267_877_0, i_8_267_904_0,
    i_8_267_907_0, i_8_267_925_0, i_8_267_975_0, i_8_267_986_0,
    i_8_267_1027_0, i_8_267_1074_0, i_8_267_1110_0, i_8_267_1186_0,
    i_8_267_1249_0, i_8_267_1250_0, i_8_267_1255_0, i_8_267_1281_0,
    i_8_267_1284_0, i_8_267_1341_0, i_8_267_1342_0, i_8_267_1420_0,
    i_8_267_1426_0, i_8_267_1435_0, i_8_267_1443_0, i_8_267_1470_0,
    i_8_267_1472_0, i_8_267_1492_0, i_8_267_1528_0, i_8_267_1541_0,
    i_8_267_1555_0, i_8_267_1588_0, i_8_267_1589_0, i_8_267_1596_0,
    i_8_267_1597_0, i_8_267_1598_0, i_8_267_1634_0, i_8_267_1647_0,
    i_8_267_1678_0, i_8_267_1699_0, i_8_267_1706_0, i_8_267_1711_0,
    i_8_267_1737_0, i_8_267_1753_0, i_8_267_1782_0, i_8_267_1796_0,
    i_8_267_1818_0, i_8_267_1819_0, i_8_267_1834_0, i_8_267_1844_0,
    i_8_267_1855_0, i_8_267_1867_0, i_8_267_1870_0, i_8_267_1903_0,
    i_8_267_1975_0, i_8_267_2046_0, i_8_267_2109_0, i_8_267_2110_0,
    i_8_267_2111_0, i_8_267_2143_0, i_8_267_2183_0, i_8_267_2190_0,
    i_8_267_2224_0, i_8_267_2244_0, i_8_267_2272_0;
  output o_8_267_0_0;
  assign o_8_267_0_0 = 0;
endmodule



// Benchmark "kernel_8_268" written by ABC on Sun Jul 19 10:07:44 2020

module kernel_8_268 ( 
    i_8_268_9_0, i_8_268_72_0, i_8_268_108_0, i_8_268_111_0, i_8_268_135_0,
    i_8_268_162_0, i_8_268_183_0, i_8_268_228_0, i_8_268_234_0,
    i_8_268_262_0, i_8_268_361_0, i_8_268_363_0, i_8_268_396_0,
    i_8_268_477_0, i_8_268_479_0, i_8_268_480_0, i_8_268_481_0,
    i_8_268_498_0, i_8_268_522_0, i_8_268_543_0, i_8_268_549_0,
    i_8_268_567_0, i_8_268_568_0, i_8_268_570_0, i_8_268_571_0,
    i_8_268_603_0, i_8_268_633_0, i_8_268_636_0, i_8_268_652_0,
    i_8_268_675_0, i_8_268_676_0, i_8_268_677_0, i_8_268_684_0,
    i_8_268_748_0, i_8_268_759_0, i_8_268_793_0, i_8_268_855_0,
    i_8_268_936_0, i_8_268_966_0, i_8_268_999_0, i_8_268_1010_0,
    i_8_268_1036_0, i_8_268_1183_0, i_8_268_1188_0, i_8_268_1228_0,
    i_8_268_1236_0, i_8_268_1263_0, i_8_268_1272_0, i_8_268_1296_0,
    i_8_268_1315_0, i_8_268_1323_0, i_8_268_1332_0, i_8_268_1434_0,
    i_8_268_1459_0, i_8_268_1476_0, i_8_268_1485_0, i_8_268_1486_0,
    i_8_268_1512_0, i_8_268_1521_0, i_8_268_1522_0, i_8_268_1553_0,
    i_8_268_1585_0, i_8_268_1596_0, i_8_268_1647_0, i_8_268_1650_0,
    i_8_268_1683_0, i_8_268_1696_0, i_8_268_1704_0, i_8_268_1719_0,
    i_8_268_1728_0, i_8_268_1737_0, i_8_268_1752_0, i_8_268_1755_0,
    i_8_268_1773_0, i_8_268_1774_0, i_8_268_1776_0, i_8_268_1804_0,
    i_8_268_1818_0, i_8_268_1827_0, i_8_268_1836_0, i_8_268_1837_0,
    i_8_268_1838_0, i_8_268_1839_0, i_8_268_1840_0, i_8_268_1846_0,
    i_8_268_1854_0, i_8_268_1881_0, i_8_268_1993_0, i_8_268_2070_0,
    i_8_268_2118_0, i_8_268_2133_0, i_8_268_2145_0, i_8_268_2146_0,
    i_8_268_2188_0, i_8_268_2214_0, i_8_268_2223_0, i_8_268_2241_0,
    i_8_268_2242_0, i_8_268_2262_0, i_8_268_2295_0,
    o_8_268_0_0  );
  input  i_8_268_9_0, i_8_268_72_0, i_8_268_108_0, i_8_268_111_0,
    i_8_268_135_0, i_8_268_162_0, i_8_268_183_0, i_8_268_228_0,
    i_8_268_234_0, i_8_268_262_0, i_8_268_361_0, i_8_268_363_0,
    i_8_268_396_0, i_8_268_477_0, i_8_268_479_0, i_8_268_480_0,
    i_8_268_481_0, i_8_268_498_0, i_8_268_522_0, i_8_268_543_0,
    i_8_268_549_0, i_8_268_567_0, i_8_268_568_0, i_8_268_570_0,
    i_8_268_571_0, i_8_268_603_0, i_8_268_633_0, i_8_268_636_0,
    i_8_268_652_0, i_8_268_675_0, i_8_268_676_0, i_8_268_677_0,
    i_8_268_684_0, i_8_268_748_0, i_8_268_759_0, i_8_268_793_0,
    i_8_268_855_0, i_8_268_936_0, i_8_268_966_0, i_8_268_999_0,
    i_8_268_1010_0, i_8_268_1036_0, i_8_268_1183_0, i_8_268_1188_0,
    i_8_268_1228_0, i_8_268_1236_0, i_8_268_1263_0, i_8_268_1272_0,
    i_8_268_1296_0, i_8_268_1315_0, i_8_268_1323_0, i_8_268_1332_0,
    i_8_268_1434_0, i_8_268_1459_0, i_8_268_1476_0, i_8_268_1485_0,
    i_8_268_1486_0, i_8_268_1512_0, i_8_268_1521_0, i_8_268_1522_0,
    i_8_268_1553_0, i_8_268_1585_0, i_8_268_1596_0, i_8_268_1647_0,
    i_8_268_1650_0, i_8_268_1683_0, i_8_268_1696_0, i_8_268_1704_0,
    i_8_268_1719_0, i_8_268_1728_0, i_8_268_1737_0, i_8_268_1752_0,
    i_8_268_1755_0, i_8_268_1773_0, i_8_268_1774_0, i_8_268_1776_0,
    i_8_268_1804_0, i_8_268_1818_0, i_8_268_1827_0, i_8_268_1836_0,
    i_8_268_1837_0, i_8_268_1838_0, i_8_268_1839_0, i_8_268_1840_0,
    i_8_268_1846_0, i_8_268_1854_0, i_8_268_1881_0, i_8_268_1993_0,
    i_8_268_2070_0, i_8_268_2118_0, i_8_268_2133_0, i_8_268_2145_0,
    i_8_268_2146_0, i_8_268_2188_0, i_8_268_2214_0, i_8_268_2223_0,
    i_8_268_2241_0, i_8_268_2242_0, i_8_268_2262_0, i_8_268_2295_0;
  output o_8_268_0_0;
  assign o_8_268_0_0 = 0;
endmodule



// Benchmark "kernel_8_269" written by ABC on Sun Jul 19 10:07:45 2020

module kernel_8_269 ( 
    i_8_269_1_0, i_8_269_24_0, i_8_269_28_0, i_8_269_62_0, i_8_269_64_0,
    i_8_269_155_0, i_8_269_163_0, i_8_269_166_0, i_8_269_189_0,
    i_8_269_193_0, i_8_269_217_0, i_8_269_218_0, i_8_269_220_0,
    i_8_269_234_0, i_8_269_240_0, i_8_269_256_0, i_8_269_293_0,
    i_8_269_296_0, i_8_269_304_0, i_8_269_334_0, i_8_269_338_0,
    i_8_269_360_0, i_8_269_361_0, i_8_269_385_0, i_8_269_386_0,
    i_8_269_425_0, i_8_269_490_0, i_8_269_593_0, i_8_269_602_0,
    i_8_269_619_0, i_8_269_620_0, i_8_269_631_0, i_8_269_658_0,
    i_8_269_693_0, i_8_269_704_0, i_8_269_707_0, i_8_269_709_0,
    i_8_269_731_0, i_8_269_757_0, i_8_269_777_0, i_8_269_789_0,
    i_8_269_812_0, i_8_269_843_0, i_8_269_848_0, i_8_269_854_0,
    i_8_269_881_0, i_8_269_1123_0, i_8_269_1127_0, i_8_269_1154_0,
    i_8_269_1157_0, i_8_269_1179_0, i_8_269_1180_0, i_8_269_1181_0,
    i_8_269_1261_0, i_8_269_1271_0, i_8_269_1274_0, i_8_269_1277_0,
    i_8_269_1293_0, i_8_269_1302_0, i_8_269_1330_0, i_8_269_1341_0,
    i_8_269_1388_0, i_8_269_1391_0, i_8_269_1408_0, i_8_269_1410_0,
    i_8_269_1473_0, i_8_269_1474_0, i_8_269_1538_0, i_8_269_1545_0,
    i_8_269_1546_0, i_8_269_1548_0, i_8_269_1549_0, i_8_269_1586_0,
    i_8_269_1601_0, i_8_269_1604_0, i_8_269_1629_0, i_8_269_1654_0,
    i_8_269_1678_0, i_8_269_1720_0, i_8_269_1735_0, i_8_269_1776_0,
    i_8_269_1800_0, i_8_269_1818_0, i_8_269_1819_0, i_8_269_1846_0,
    i_8_269_1860_0, i_8_269_1887_0, i_8_269_2005_0, i_8_269_2051_0,
    i_8_269_2077_0, i_8_269_2116_0, i_8_269_2117_0, i_8_269_2150_0,
    i_8_269_2154_0, i_8_269_2155_0, i_8_269_2230_0, i_8_269_2269_0,
    i_8_269_2291_0, i_8_269_2295_0, i_8_269_2297_0,
    o_8_269_0_0  );
  input  i_8_269_1_0, i_8_269_24_0, i_8_269_28_0, i_8_269_62_0,
    i_8_269_64_0, i_8_269_155_0, i_8_269_163_0, i_8_269_166_0,
    i_8_269_189_0, i_8_269_193_0, i_8_269_217_0, i_8_269_218_0,
    i_8_269_220_0, i_8_269_234_0, i_8_269_240_0, i_8_269_256_0,
    i_8_269_293_0, i_8_269_296_0, i_8_269_304_0, i_8_269_334_0,
    i_8_269_338_0, i_8_269_360_0, i_8_269_361_0, i_8_269_385_0,
    i_8_269_386_0, i_8_269_425_0, i_8_269_490_0, i_8_269_593_0,
    i_8_269_602_0, i_8_269_619_0, i_8_269_620_0, i_8_269_631_0,
    i_8_269_658_0, i_8_269_693_0, i_8_269_704_0, i_8_269_707_0,
    i_8_269_709_0, i_8_269_731_0, i_8_269_757_0, i_8_269_777_0,
    i_8_269_789_0, i_8_269_812_0, i_8_269_843_0, i_8_269_848_0,
    i_8_269_854_0, i_8_269_881_0, i_8_269_1123_0, i_8_269_1127_0,
    i_8_269_1154_0, i_8_269_1157_0, i_8_269_1179_0, i_8_269_1180_0,
    i_8_269_1181_0, i_8_269_1261_0, i_8_269_1271_0, i_8_269_1274_0,
    i_8_269_1277_0, i_8_269_1293_0, i_8_269_1302_0, i_8_269_1330_0,
    i_8_269_1341_0, i_8_269_1388_0, i_8_269_1391_0, i_8_269_1408_0,
    i_8_269_1410_0, i_8_269_1473_0, i_8_269_1474_0, i_8_269_1538_0,
    i_8_269_1545_0, i_8_269_1546_0, i_8_269_1548_0, i_8_269_1549_0,
    i_8_269_1586_0, i_8_269_1601_0, i_8_269_1604_0, i_8_269_1629_0,
    i_8_269_1654_0, i_8_269_1678_0, i_8_269_1720_0, i_8_269_1735_0,
    i_8_269_1776_0, i_8_269_1800_0, i_8_269_1818_0, i_8_269_1819_0,
    i_8_269_1846_0, i_8_269_1860_0, i_8_269_1887_0, i_8_269_2005_0,
    i_8_269_2051_0, i_8_269_2077_0, i_8_269_2116_0, i_8_269_2117_0,
    i_8_269_2150_0, i_8_269_2154_0, i_8_269_2155_0, i_8_269_2230_0,
    i_8_269_2269_0, i_8_269_2291_0, i_8_269_2295_0, i_8_269_2297_0;
  output o_8_269_0_0;
  assign o_8_269_0_0 = ~((~i_8_269_1181_0 & ((~i_8_269_1_0 & ((~i_8_269_189_0 & i_8_269_338_0 & ~i_8_269_789_0 & ~i_8_269_881_0 & ~i_8_269_1388_0 & ~i_8_269_1720_0) | (~i_8_269_296_0 & ~i_8_269_386_0 & i_8_269_425_0 & ~i_8_269_619_0 & ~i_8_269_854_0 & ~i_8_269_1474_0 & ~i_8_269_2116_0))) | (~i_8_269_28_0 & ~i_8_269_1274_0 & ((~i_8_269_163_0 & ~i_8_269_293_0 & ~i_8_269_296_0 & ~i_8_269_1546_0 & ~i_8_269_1601_0 & i_8_269_1678_0) | (~i_8_269_166_0 & ~i_8_269_304_0 & ~i_8_269_385_0 & ~i_8_269_709_0 & ~i_8_269_789_0 & ~i_8_269_1157_0 & ~i_8_269_1277_0 & i_8_269_1549_0 & ~i_8_269_2116_0 & ~i_8_269_2117_0 & ~i_8_269_2155_0 & ~i_8_269_2295_0 & ~i_8_269_2297_0))) | (~i_8_269_62_0 & ~i_8_269_163_0 & ~i_8_269_293_0 & ~i_8_269_593_0 & ~i_8_269_602_0 & ~i_8_269_789_0 & ~i_8_269_812_0 & ~i_8_269_848_0 & ~i_8_269_854_0 & ~i_8_269_1261_0 & ~i_8_269_1473_0 & ~i_8_269_1538_0 & ~i_8_269_1545_0 & ~i_8_269_1601_0 & ~i_8_269_2116_0))) | (~i_8_269_602_0 & ((~i_8_269_1586_0 & ((~i_8_269_62_0 & ~i_8_269_1123_0 & ((~i_8_269_155_0 & i_8_269_620_0 & ~i_8_269_1388_0 & ~i_8_269_1601_0) | (~i_8_269_189_0 & ~i_8_269_709_0 & ~i_8_269_757_0 & ~i_8_269_1261_0 & ~i_8_269_2116_0 & ~i_8_269_2117_0 & i_8_269_2155_0))) | (~i_8_269_296_0 & ~i_8_269_1601_0 & ((~i_8_269_24_0 & ~i_8_269_217_0 & ~i_8_269_234_0 & ~i_8_269_293_0 & ~i_8_269_386_0 & ~i_8_269_731_0 & ~i_8_269_789_0 & ~i_8_269_854_0 & ~i_8_269_1271_0 & ~i_8_269_1274_0 & ~i_8_269_1720_0 & ~i_8_269_1887_0 & ~i_8_269_2295_0) | (i_8_269_304_0 & ~i_8_269_631_0 & ~i_8_269_1388_0 & ~i_8_269_1545_0 & ~i_8_269_1546_0 & ~i_8_269_1800_0 & ~i_8_269_2297_0))))) | (~i_8_269_189_0 & ~i_8_269_234_0 & ~i_8_269_256_0 & ~i_8_269_1846_0 & i_8_269_1860_0 & ~i_8_269_2051_0 & ~i_8_269_2150_0) | (~i_8_269_64_0 & ~i_8_269_166_0 & ~i_8_269_304_0 & ~i_8_269_425_0 & ~i_8_269_1302_0 & ~i_8_269_1391_0 & ~i_8_269_1474_0 & ~i_8_269_1549_0 & i_8_269_1678_0 & ~i_8_269_2295_0))) | (~i_8_269_293_0 & ((~i_8_269_24_0 & ((~i_8_269_28_0 & ~i_8_269_62_0 & ~i_8_269_163_0 & ~i_8_269_296_0 & ~i_8_269_757_0 & ~i_8_269_789_0 & ~i_8_269_854_0 & ~i_8_269_1179_0 & ~i_8_269_1408_0 & ~i_8_269_1473_0 & ~i_8_269_1538_0 & ~i_8_269_1548_0 & ~i_8_269_1549_0 & ~i_8_269_1586_0 & ~i_8_269_2117_0) | (i_8_269_361_0 & ~i_8_269_593_0 & ~i_8_269_812_0 & ~i_8_269_1388_0 & ~i_8_269_2297_0))) | (~i_8_269_2297_0 & ((~i_8_269_593_0 & ~i_8_269_1274_0 & ~i_8_269_1538_0 & i_8_269_1548_0 & ~i_8_269_1549_0) | (i_8_269_704_0 & ~i_8_269_731_0 & ~i_8_269_1179_0 & ~i_8_269_2051_0))) | (~i_8_269_28_0 & ~i_8_269_189_0 & i_8_269_361_0 & ~i_8_269_709_0 & i_8_269_881_0))) | (~i_8_269_163_0 & ((i_8_269_360_0 & ~i_8_269_731_0 & ~i_8_269_1601_0) | (~i_8_269_334_0 & ~i_8_269_386_0 & i_8_269_707_0 & ~i_8_269_1408_0 & ~i_8_269_1546_0 & ~i_8_269_1586_0 & ~i_8_269_2230_0 & ~i_8_269_2295_0))) | (~i_8_269_217_0 & ((~i_8_269_848_0 & ~i_8_269_1123_0 & ~i_8_269_1391_0 & ~i_8_269_1538_0 & i_8_269_2005_0) | (~i_8_269_220_0 & i_8_269_304_0 & ~i_8_269_593_0 & ~i_8_269_854_0 & ~i_8_269_1277_0 & ~i_8_269_1408_0 & ~i_8_269_1549_0 & ~i_8_269_1678_0 & ~i_8_269_2155_0 & ~i_8_269_2295_0))) | (i_8_269_620_0 & ((~i_8_269_296_0 & ~i_8_269_386_0 & ~i_8_269_881_0 & ~i_8_269_1545_0) | (i_8_269_709_0 & ~i_8_269_1474_0 & ~i_8_269_1720_0 & ~i_8_269_2291_0))) | (~i_8_269_1391_0 & ((~i_8_269_304_0 & ((~i_8_269_386_0 & ~i_8_269_789_0 & ~i_8_269_1388_0 & i_8_269_1735_0 & ~i_8_269_2155_0) | (i_8_269_217_0 & ~i_8_269_360_0 & ~i_8_269_881_0 & ~i_8_269_1546_0 & ~i_8_269_1846_0 & ~i_8_269_2117_0 & ~i_8_269_2297_0))) | (~i_8_269_693_0 & ~i_8_269_709_0 & ~i_8_269_1408_0 & ~i_8_269_1654_0 & ((~i_8_269_62_0 & ~i_8_269_334_0 & ~i_8_269_386_0 & ~i_8_269_490_0 & ~i_8_269_593_0 & ~i_8_269_619_0 & ~i_8_269_848_0 & ~i_8_269_1180_0 & ~i_8_269_1388_0 & ~i_8_269_1473_0 & ~i_8_269_2116_0) | (~i_8_269_189_0 & ~i_8_269_296_0 & ~i_8_269_757_0 & ~i_8_269_881_0 & ~i_8_269_1154_0 & ~i_8_269_1274_0 & ~i_8_269_1277_0 & ~i_8_269_1330_0 & ~i_8_269_1545_0 & ~i_8_269_2117_0 & ~i_8_269_2155_0))))) | (~i_8_269_296_0 & ((~i_8_269_386_0 & ~i_8_269_1546_0 & ~i_8_269_1586_0 & (i_8_269_1410_0 | (i_8_269_220_0 & ~i_8_269_709_0 & ~i_8_269_1261_0 & ~i_8_269_1277_0 & ~i_8_269_2230_0 & ~i_8_269_2295_0 & ~i_8_269_1388_0 & ~i_8_269_2150_0))) | (~i_8_269_843_0 & ~i_8_269_1545_0 & ((~i_8_269_593_0 & i_8_269_1887_0) | (i_8_269_2150_0 & ~i_8_269_2155_0 & i_8_269_2230_0 & ~i_8_269_2291_0))) | (~i_8_269_704_0 & ~i_8_269_854_0 & i_8_269_1157_0 & ~i_8_269_1274_0 & ~i_8_269_1408_0))) | (i_8_269_843_0 & ((i_8_269_709_0 & i_8_269_1887_0) | (~i_8_269_731_0 & ~i_8_269_1123_0 & ~i_8_269_1410_0 & ~i_8_269_1473_0 & ~i_8_269_1474_0 & ~i_8_269_1549_0 & ~i_8_269_1654_0 & ~i_8_269_2005_0 & ~i_8_269_2116_0))) | (~i_8_269_1123_0 & ~i_8_269_2117_0 & ((~i_8_269_28_0 & i_8_269_338_0 & ~i_8_269_385_0 & ~i_8_269_789_0 & ~i_8_269_812_0 & ~i_8_269_1545_0) | (~i_8_269_854_0 & ~i_8_269_1274_0 & ~i_8_269_1388_0 & ~i_8_269_1586_0 & i_8_269_2154_0))) | (i_8_269_218_0 & ~i_8_269_593_0 & ~i_8_269_1271_0 & ~i_8_269_1388_0 & i_8_269_1408_0) | (~i_8_269_304_0 & i_8_269_1293_0 & ~i_8_269_2077_0) | (i_8_269_1549_0 & i_8_269_1604_0 & ~i_8_269_1846_0 & ~i_8_269_2155_0));
endmodule



// Benchmark "kernel_8_270" written by ABC on Sun Jul 19 10:07:46 2020

module kernel_8_270 ( 
    i_8_270_35_0, i_8_270_169_0, i_8_270_339_0, i_8_270_447_0,
    i_8_270_453_0, i_8_270_456_0, i_8_270_483_0, i_8_270_492_0,
    i_8_270_502_0, i_8_270_510_0, i_8_270_527_0, i_8_270_574_0,
    i_8_270_627_0, i_8_270_655_0, i_8_270_696_0, i_8_270_699_0,
    i_8_270_705_0, i_8_270_708_0, i_8_270_762_0, i_8_270_780_0,
    i_8_270_808_0, i_8_270_834_0, i_8_270_840_0, i_8_270_843_0,
    i_8_270_886_0, i_8_270_941_0, i_8_270_943_0, i_8_270_946_0,
    i_8_270_947_0, i_8_270_958_0, i_8_270_967_0, i_8_270_969_0,
    i_8_270_987_0, i_8_270_993_0, i_8_270_996_0, i_8_270_1032_0,
    i_8_270_1050_0, i_8_270_1060_0, i_8_270_1069_0, i_8_270_1093_0,
    i_8_270_1129_0, i_8_270_1168_0, i_8_270_1185_0, i_8_270_1186_0,
    i_8_270_1187_0, i_8_270_1232_0, i_8_270_1258_0, i_8_270_1285_0,
    i_8_270_1286_0, i_8_270_1306_0, i_8_270_1307_0, i_8_270_1310_0,
    i_8_270_1312_0, i_8_270_1336_0, i_8_270_1402_0, i_8_270_1410_0,
    i_8_270_1411_0, i_8_270_1438_0, i_8_270_1474_0, i_8_270_1490_0,
    i_8_270_1492_0, i_8_270_1510_0, i_8_270_1537_0, i_8_270_1538_0,
    i_8_270_1545_0, i_8_270_1554_0, i_8_270_1591_0, i_8_270_1624_0,
    i_8_270_1654_0, i_8_270_1655_0, i_8_270_1671_0, i_8_270_1725_0,
    i_8_270_1732_0, i_8_270_1734_0, i_8_270_1741_0, i_8_270_1744_0,
    i_8_270_1745_0, i_8_270_1762_0, i_8_270_1770_0, i_8_270_1788_0,
    i_8_270_1888_0, i_8_270_1896_0, i_8_270_1906_0, i_8_270_1984_0,
    i_8_270_2041_0, i_8_270_2058_0, i_8_270_2059_0, i_8_270_2073_0,
    i_8_270_2076_0, i_8_270_2092_0, i_8_270_2094_0, i_8_270_2095_0,
    i_8_270_2122_0, i_8_270_2132_0, i_8_270_2146_0, i_8_270_2218_0,
    i_8_270_2230_0, i_8_270_2236_0, i_8_270_2247_0, i_8_270_2302_0,
    o_8_270_0_0  );
  input  i_8_270_35_0, i_8_270_169_0, i_8_270_339_0, i_8_270_447_0,
    i_8_270_453_0, i_8_270_456_0, i_8_270_483_0, i_8_270_492_0,
    i_8_270_502_0, i_8_270_510_0, i_8_270_527_0, i_8_270_574_0,
    i_8_270_627_0, i_8_270_655_0, i_8_270_696_0, i_8_270_699_0,
    i_8_270_705_0, i_8_270_708_0, i_8_270_762_0, i_8_270_780_0,
    i_8_270_808_0, i_8_270_834_0, i_8_270_840_0, i_8_270_843_0,
    i_8_270_886_0, i_8_270_941_0, i_8_270_943_0, i_8_270_946_0,
    i_8_270_947_0, i_8_270_958_0, i_8_270_967_0, i_8_270_969_0,
    i_8_270_987_0, i_8_270_993_0, i_8_270_996_0, i_8_270_1032_0,
    i_8_270_1050_0, i_8_270_1060_0, i_8_270_1069_0, i_8_270_1093_0,
    i_8_270_1129_0, i_8_270_1168_0, i_8_270_1185_0, i_8_270_1186_0,
    i_8_270_1187_0, i_8_270_1232_0, i_8_270_1258_0, i_8_270_1285_0,
    i_8_270_1286_0, i_8_270_1306_0, i_8_270_1307_0, i_8_270_1310_0,
    i_8_270_1312_0, i_8_270_1336_0, i_8_270_1402_0, i_8_270_1410_0,
    i_8_270_1411_0, i_8_270_1438_0, i_8_270_1474_0, i_8_270_1490_0,
    i_8_270_1492_0, i_8_270_1510_0, i_8_270_1537_0, i_8_270_1538_0,
    i_8_270_1545_0, i_8_270_1554_0, i_8_270_1591_0, i_8_270_1624_0,
    i_8_270_1654_0, i_8_270_1655_0, i_8_270_1671_0, i_8_270_1725_0,
    i_8_270_1732_0, i_8_270_1734_0, i_8_270_1741_0, i_8_270_1744_0,
    i_8_270_1745_0, i_8_270_1762_0, i_8_270_1770_0, i_8_270_1788_0,
    i_8_270_1888_0, i_8_270_1896_0, i_8_270_1906_0, i_8_270_1984_0,
    i_8_270_2041_0, i_8_270_2058_0, i_8_270_2059_0, i_8_270_2073_0,
    i_8_270_2076_0, i_8_270_2092_0, i_8_270_2094_0, i_8_270_2095_0,
    i_8_270_2122_0, i_8_270_2132_0, i_8_270_2146_0, i_8_270_2218_0,
    i_8_270_2230_0, i_8_270_2236_0, i_8_270_2247_0, i_8_270_2302_0;
  output o_8_270_0_0;
  assign o_8_270_0_0 = 0;
endmodule



// Benchmark "kernel_8_271" written by ABC on Sun Jul 19 10:07:47 2020

module kernel_8_271 ( 
    i_8_271_50_0, i_8_271_112_0, i_8_271_114_0, i_8_271_218_0,
    i_8_271_253_0, i_8_271_255_0, i_8_271_301_0, i_8_271_316_0,
    i_8_271_343_0, i_8_271_361_0, i_8_271_418_0, i_8_271_426_0,
    i_8_271_427_0, i_8_271_453_0, i_8_271_454_0, i_8_271_455_0,
    i_8_271_505_0, i_8_271_532_0, i_8_271_586_0, i_8_271_595_0,
    i_8_271_639_0, i_8_271_648_0, i_8_271_650_0, i_8_271_651_0,
    i_8_271_657_0, i_8_271_661_0, i_8_271_675_0, i_8_271_676_0,
    i_8_271_677_0, i_8_271_706_0, i_8_271_713_0, i_8_271_820_0,
    i_8_271_849_0, i_8_271_850_0, i_8_271_875_0, i_8_271_886_0,
    i_8_271_892_0, i_8_271_991_0, i_8_271_992_0, i_8_271_1035_0,
    i_8_271_1054_0, i_8_271_1055_0, i_8_271_1102_0, i_8_271_1127_0,
    i_8_271_1217_0, i_8_271_1226_0, i_8_271_1234_0, i_8_271_1264_0,
    i_8_271_1270_0, i_8_271_1325_0, i_8_271_1327_0, i_8_271_1336_0,
    i_8_271_1424_0, i_8_271_1439_0, i_8_271_1452_0, i_8_271_1459_0,
    i_8_271_1462_0, i_8_271_1486_0, i_8_271_1487_0, i_8_271_1522_0,
    i_8_271_1524_0, i_8_271_1549_0, i_8_271_1603_0, i_8_271_1611_0,
    i_8_271_1612_0, i_8_271_1615_0, i_8_271_1629_0, i_8_271_1676_0,
    i_8_271_1680_0, i_8_271_1682_0, i_8_271_1693_0, i_8_271_1705_0,
    i_8_271_1747_0, i_8_271_1749_0, i_8_271_1769_0, i_8_271_1791_0,
    i_8_271_1810_0, i_8_271_1811_0, i_8_271_1825_0, i_8_271_1837_0,
    i_8_271_1881_0, i_8_271_1945_0, i_8_271_1946_0, i_8_271_1954_0,
    i_8_271_1957_0, i_8_271_1963_0, i_8_271_1966_0, i_8_271_1972_0,
    i_8_271_1981_0, i_8_271_1984_0, i_8_271_1990_0, i_8_271_2029_0,
    i_8_271_2054_0, i_8_271_2126_0, i_8_271_2223_0, i_8_271_2244_0,
    i_8_271_2245_0, i_8_271_2246_0, i_8_271_2260_0, i_8_271_2263_0,
    o_8_271_0_0  );
  input  i_8_271_50_0, i_8_271_112_0, i_8_271_114_0, i_8_271_218_0,
    i_8_271_253_0, i_8_271_255_0, i_8_271_301_0, i_8_271_316_0,
    i_8_271_343_0, i_8_271_361_0, i_8_271_418_0, i_8_271_426_0,
    i_8_271_427_0, i_8_271_453_0, i_8_271_454_0, i_8_271_455_0,
    i_8_271_505_0, i_8_271_532_0, i_8_271_586_0, i_8_271_595_0,
    i_8_271_639_0, i_8_271_648_0, i_8_271_650_0, i_8_271_651_0,
    i_8_271_657_0, i_8_271_661_0, i_8_271_675_0, i_8_271_676_0,
    i_8_271_677_0, i_8_271_706_0, i_8_271_713_0, i_8_271_820_0,
    i_8_271_849_0, i_8_271_850_0, i_8_271_875_0, i_8_271_886_0,
    i_8_271_892_0, i_8_271_991_0, i_8_271_992_0, i_8_271_1035_0,
    i_8_271_1054_0, i_8_271_1055_0, i_8_271_1102_0, i_8_271_1127_0,
    i_8_271_1217_0, i_8_271_1226_0, i_8_271_1234_0, i_8_271_1264_0,
    i_8_271_1270_0, i_8_271_1325_0, i_8_271_1327_0, i_8_271_1336_0,
    i_8_271_1424_0, i_8_271_1439_0, i_8_271_1452_0, i_8_271_1459_0,
    i_8_271_1462_0, i_8_271_1486_0, i_8_271_1487_0, i_8_271_1522_0,
    i_8_271_1524_0, i_8_271_1549_0, i_8_271_1603_0, i_8_271_1611_0,
    i_8_271_1612_0, i_8_271_1615_0, i_8_271_1629_0, i_8_271_1676_0,
    i_8_271_1680_0, i_8_271_1682_0, i_8_271_1693_0, i_8_271_1705_0,
    i_8_271_1747_0, i_8_271_1749_0, i_8_271_1769_0, i_8_271_1791_0,
    i_8_271_1810_0, i_8_271_1811_0, i_8_271_1825_0, i_8_271_1837_0,
    i_8_271_1881_0, i_8_271_1945_0, i_8_271_1946_0, i_8_271_1954_0,
    i_8_271_1957_0, i_8_271_1963_0, i_8_271_1966_0, i_8_271_1972_0,
    i_8_271_1981_0, i_8_271_1984_0, i_8_271_1990_0, i_8_271_2029_0,
    i_8_271_2054_0, i_8_271_2126_0, i_8_271_2223_0, i_8_271_2244_0,
    i_8_271_2245_0, i_8_271_2246_0, i_8_271_2260_0, i_8_271_2263_0;
  output o_8_271_0_0;
  assign o_8_271_0_0 = 0;
endmodule



// Benchmark "kernel_8_272" written by ABC on Sun Jul 19 10:07:49 2020

module kernel_8_272 ( 
    i_8_272_25_0, i_8_272_70_0, i_8_272_94_0, i_8_272_96_0, i_8_272_185_0,
    i_8_272_215_0, i_8_272_229_0, i_8_272_301_0, i_8_272_328_0,
    i_8_272_329_0, i_8_272_345_0, i_8_272_373_0, i_8_272_374_0,
    i_8_272_379_0, i_8_272_383_0, i_8_272_423_0, i_8_272_462_0,
    i_8_272_592_0, i_8_272_593_0, i_8_272_606_0, i_8_272_608_0,
    i_8_272_612_0, i_8_272_621_0, i_8_272_622_0, i_8_272_623_0,
    i_8_272_625_0, i_8_272_626_0, i_8_272_638_0, i_8_272_702_0,
    i_8_272_703_0, i_8_272_704_0, i_8_272_705_0, i_8_272_713_0,
    i_8_272_720_0, i_8_272_723_0, i_8_272_778_0, i_8_272_779_0,
    i_8_272_854_0, i_8_272_934_0, i_8_272_973_0, i_8_272_984_0,
    i_8_272_985_0, i_8_272_986_0, i_8_272_987_0, i_8_272_988_0,
    i_8_272_989_0, i_8_272_996_0, i_8_272_997_0, i_8_272_1027_0,
    i_8_272_1123_0, i_8_272_1191_0, i_8_272_1272_0, i_8_272_1273_0,
    i_8_272_1297_0, i_8_272_1305_0, i_8_272_1307_0, i_8_272_1330_0,
    i_8_272_1402_0, i_8_272_1410_0, i_8_272_1470_0, i_8_272_1471_0,
    i_8_272_1473_0, i_8_272_1483_0, i_8_272_1526_0, i_8_272_1529_0,
    i_8_272_1621_0, i_8_272_1623_0, i_8_272_1625_0, i_8_272_1626_0,
    i_8_272_1651_0, i_8_272_1661_0, i_8_272_1731_0, i_8_272_1733_0,
    i_8_272_1734_0, i_8_272_1735_0, i_8_272_1736_0, i_8_272_1752_0,
    i_8_272_1776_0, i_8_272_1789_0, i_8_272_1790_0, i_8_272_1818_0,
    i_8_272_1841_0, i_8_272_1857_0, i_8_272_1860_0, i_8_272_1862_0,
    i_8_272_1902_0, i_8_272_1950_0, i_8_272_1965_0, i_8_272_1967_0,
    i_8_272_1980_0, i_8_272_2015_0, i_8_272_2025_0, i_8_272_2026_0,
    i_8_272_2058_0, i_8_272_2070_0, i_8_272_2076_0, i_8_272_2154_0,
    i_8_272_2156_0, i_8_272_2169_0, i_8_272_2237_0,
    o_8_272_0_0  );
  input  i_8_272_25_0, i_8_272_70_0, i_8_272_94_0, i_8_272_96_0,
    i_8_272_185_0, i_8_272_215_0, i_8_272_229_0, i_8_272_301_0,
    i_8_272_328_0, i_8_272_329_0, i_8_272_345_0, i_8_272_373_0,
    i_8_272_374_0, i_8_272_379_0, i_8_272_383_0, i_8_272_423_0,
    i_8_272_462_0, i_8_272_592_0, i_8_272_593_0, i_8_272_606_0,
    i_8_272_608_0, i_8_272_612_0, i_8_272_621_0, i_8_272_622_0,
    i_8_272_623_0, i_8_272_625_0, i_8_272_626_0, i_8_272_638_0,
    i_8_272_702_0, i_8_272_703_0, i_8_272_704_0, i_8_272_705_0,
    i_8_272_713_0, i_8_272_720_0, i_8_272_723_0, i_8_272_778_0,
    i_8_272_779_0, i_8_272_854_0, i_8_272_934_0, i_8_272_973_0,
    i_8_272_984_0, i_8_272_985_0, i_8_272_986_0, i_8_272_987_0,
    i_8_272_988_0, i_8_272_989_0, i_8_272_996_0, i_8_272_997_0,
    i_8_272_1027_0, i_8_272_1123_0, i_8_272_1191_0, i_8_272_1272_0,
    i_8_272_1273_0, i_8_272_1297_0, i_8_272_1305_0, i_8_272_1307_0,
    i_8_272_1330_0, i_8_272_1402_0, i_8_272_1410_0, i_8_272_1470_0,
    i_8_272_1471_0, i_8_272_1473_0, i_8_272_1483_0, i_8_272_1526_0,
    i_8_272_1529_0, i_8_272_1621_0, i_8_272_1623_0, i_8_272_1625_0,
    i_8_272_1626_0, i_8_272_1651_0, i_8_272_1661_0, i_8_272_1731_0,
    i_8_272_1733_0, i_8_272_1734_0, i_8_272_1735_0, i_8_272_1736_0,
    i_8_272_1752_0, i_8_272_1776_0, i_8_272_1789_0, i_8_272_1790_0,
    i_8_272_1818_0, i_8_272_1841_0, i_8_272_1857_0, i_8_272_1860_0,
    i_8_272_1862_0, i_8_272_1902_0, i_8_272_1950_0, i_8_272_1965_0,
    i_8_272_1967_0, i_8_272_1980_0, i_8_272_2015_0, i_8_272_2025_0,
    i_8_272_2026_0, i_8_272_2058_0, i_8_272_2070_0, i_8_272_2076_0,
    i_8_272_2154_0, i_8_272_2156_0, i_8_272_2169_0, i_8_272_2237_0;
  output o_8_272_0_0;
  assign o_8_272_0_0 = ~((~i_8_272_1734_0 & ((~i_8_272_96_0 & ~i_8_272_2076_0 & ((~i_8_272_301_0 & ~i_8_272_622_0 & ~i_8_272_1273_0 & ~i_8_272_1626_0 & ~i_8_272_1862_0 & ~i_8_272_2025_0 & i_8_272_2058_0) | (~i_8_272_328_0 & ~i_8_272_623_0 & ~i_8_272_705_0 & ~i_8_272_988_0 & ~i_8_272_996_0 & ~i_8_272_1410_0 & ~i_8_272_1731_0 & ~i_8_272_1736_0 & ~i_8_272_1857_0 & ~i_8_272_2026_0 & i_8_272_2154_0))) | (i_8_272_229_0 & ((~i_8_272_301_0 & ~i_8_272_329_0 & ~i_8_272_704_0 & ~i_8_272_1027_0 & ~i_8_272_1273_0 & ~i_8_272_1526_0 & ~i_8_272_1736_0 & ~i_8_272_1860_0 & ~i_8_272_2025_0) | (~i_8_272_70_0 & ~i_8_272_720_0 & ~i_8_272_973_0 & ~i_8_272_1529_0 & ~i_8_272_1661_0 & i_8_272_1789_0 & ~i_8_272_2058_0))) | (~i_8_272_1731_0 & ((~i_8_272_70_0 & ((~i_8_272_1123_0 & i_8_272_1473_0 & ~i_8_272_1860_0) | (i_8_272_592_0 & ~i_8_272_713_0 & ~i_8_272_778_0 & ~i_8_272_1623_0 & ~i_8_272_1736_0 & ~i_8_272_1902_0 & ~i_8_272_2058_0))) | (~i_8_272_997_0 & ((~i_8_272_623_0 & ~i_8_272_625_0 & ~i_8_272_713_0 & ~i_8_272_1027_0 & ~i_8_272_1623_0 & ~i_8_272_1736_0 & i_8_272_1965_0 & ~i_8_272_2026_0) | (~i_8_272_622_0 & ~i_8_272_1735_0 & i_8_272_1752_0 & ~i_8_272_2058_0))))) | (i_8_272_705_0 & ((~i_8_272_383_0 & i_8_272_702_0 & i_8_272_703_0 & ~i_8_272_997_0) | (~i_8_272_621_0 & ~i_8_272_720_0 & ~i_8_272_1272_0 & ~i_8_272_1410_0 & i_8_272_1818_0 & ~i_8_272_2025_0))) | (~i_8_272_1027_0 & ((~i_8_272_621_0 & ~i_8_272_1626_0 & ((i_8_272_345_0 & ~i_8_272_720_0 & ~i_8_272_1623_0 & ~i_8_272_1733_0 & ~i_8_272_1965_0) | (i_8_272_383_0 & ~i_8_272_986_0 & ~i_8_272_989_0 & ~i_8_272_1529_0 & ~i_8_272_1860_0 & i_8_272_2156_0))) | (~i_8_272_94_0 & ~i_8_272_713_0 & ~i_8_272_720_0 & ~i_8_272_779_0 & ~i_8_272_984_0 & i_8_272_1297_0 & ~i_8_272_1470_0 & ~i_8_272_2015_0 & ~i_8_272_2025_0 & ~i_8_272_2026_0))) | (~i_8_272_215_0 & i_8_272_301_0 & ~i_8_272_462_0 & ~i_8_272_623_0 & ~i_8_272_626_0 & ~i_8_272_705_0 & ~i_8_272_723_0 & ~i_8_272_778_0 & ~i_8_272_779_0 & ~i_8_272_996_0 & ~i_8_272_1529_0 & ~i_8_272_1621_0 & ~i_8_272_1860_0))) | (~i_8_272_1735_0 & ((~i_8_272_94_0 & ((i_8_272_612_0 & ~i_8_272_621_0 & ~i_8_272_622_0 & ~i_8_272_713_0 & ~i_8_272_1733_0 & ~i_8_272_1736_0 & ~i_8_272_1860_0 & ~i_8_272_1902_0) | (~i_8_272_301_0 & ~i_8_272_592_0 & ~i_8_272_779_0 & ~i_8_272_987_0 & i_8_272_1330_0 & ~i_8_272_1529_0 & ~i_8_272_1857_0 & ~i_8_272_2015_0 & ~i_8_272_2154_0 & ~i_8_272_2237_0))) | (i_8_272_383_0 & ((~i_8_272_301_0 & ~i_8_272_623_0 & ~i_8_272_779_0 & ~i_8_272_1471_0 & ~i_8_272_1626_0 & ~i_8_272_1731_0 & ~i_8_272_1733_0 & ~i_8_272_1789_0 & ~i_8_272_1862_0) | (~i_8_272_622_0 & i_8_272_854_0 & i_8_272_1967_0))) | (~i_8_272_2025_0 & ((~i_8_272_623_0 & ((~i_8_272_379_0 & i_8_272_423_0 & ~i_8_272_703_0 & ~i_8_272_988_0 & ~i_8_272_1305_0 & i_8_272_1818_0) | (~i_8_272_713_0 & ~i_8_272_985_0 & ~i_8_272_989_0 & i_8_272_1123_0 & ~i_8_272_1526_0 & ~i_8_272_1860_0))) | (i_8_272_593_0 & ~i_8_272_1626_0 & ~i_8_272_1736_0 & ~i_8_272_1857_0 & ~i_8_272_1862_0 & ~i_8_272_2026_0))) | (~i_8_272_713_0 & ((~i_8_272_379_0 & ((~i_8_272_96_0 & i_8_272_625_0 & ~i_8_272_720_0 & ~i_8_272_723_0 & ~i_8_272_996_0 & ~i_8_272_1027_0 & i_8_272_1776_0) | (~i_8_272_626_0 & i_8_272_704_0 & ~i_8_272_779_0 & ~i_8_272_986_0 & ~i_8_272_1862_0))) | (~i_8_272_1862_0 & ((~i_8_272_984_0 & ~i_8_272_997_0 & ~i_8_272_1027_0 & i_8_272_1483_0) | (~i_8_272_779_0 & ~i_8_272_1661_0 & i_8_272_2237_0))) | (~i_8_272_985_0 & i_8_272_1651_0 & i_8_272_2070_0))) | (~i_8_272_215_0 & ~i_8_272_229_0 & ~i_8_272_702_0 & ~i_8_272_1027_0 & ~i_8_272_1273_0 & i_8_272_1841_0 & ~i_8_272_2015_0))) | (~i_8_272_215_0 & ((~i_8_272_94_0 & i_8_272_374_0 & ~i_8_272_379_0 & ~i_8_272_621_0 & i_8_272_778_0 & ~i_8_272_1483_0 & ~i_8_272_1626_0 & ~i_8_272_1860_0) | (i_8_272_608_0 & ~i_8_272_713_0 & ~i_8_272_986_0 & ~i_8_272_1736_0 & ~i_8_272_1776_0 & ~i_8_272_2015_0 & ~i_8_272_2058_0))) | (~i_8_272_229_0 & ((i_8_272_373_0 & ~i_8_272_778_0 & ~i_8_272_1027_0 & ~i_8_272_1330_0 & ~i_8_272_1483_0 & ~i_8_272_1529_0 & ~i_8_272_1625_0 & ~i_8_272_1661_0 & ~i_8_272_1731_0 & ~i_8_272_1841_0) | (~i_8_272_329_0 & ~i_8_272_623_0 & ~i_8_272_626_0 & ~i_8_272_985_0 & ~i_8_272_988_0 & ~i_8_272_996_0 & ~i_8_272_1736_0 & ~i_8_272_2026_0 & i_8_272_2156_0))) | (~i_8_272_328_0 & ((~i_8_272_70_0 & ~i_8_272_713_0 & ~i_8_272_778_0 & ~i_8_272_986_0 & i_8_272_1307_0 & ~i_8_272_1733_0) | (~i_8_272_625_0 & i_8_272_704_0 & ~i_8_272_985_0 & ~i_8_272_1776_0 & i_8_272_1790_0))) | (~i_8_272_329_0 & ((~i_8_272_723_0 & ~i_8_272_778_0 & ~i_8_272_779_0 & ~i_8_272_70_0 & ~i_8_272_626_0 & ~i_8_272_987_0 & ~i_8_272_996_0 & ~i_8_272_1736_0 & i_8_272_1789_0 & ~i_8_272_2015_0 & ~i_8_272_2058_0) | (i_8_272_704_0 & ~i_8_272_1862_0 & i_8_272_2156_0 & ~i_8_272_2237_0))) | (~i_8_272_70_0 & ((~i_8_272_96_0 & i_8_272_592_0 & ~i_8_272_713_0 & ~i_8_272_984_0 & ~i_8_272_986_0 & ~i_8_272_1027_0 & ~i_8_272_1626_0 & i_8_272_1789_0) | (~i_8_272_621_0 & ~i_8_272_720_0 & ~i_8_272_987_0 & ~i_8_272_996_0 & ~i_8_272_1841_0 & i_8_272_2070_0))) | (~i_8_272_96_0 & ((~i_8_272_379_0 & ~i_8_272_988_0 & ~i_8_272_1027_0 & ~i_8_272_1483_0 & ~i_8_272_1626_0 & i_8_272_1651_0 & ~i_8_272_1661_0 & ~i_8_272_1857_0 & ~i_8_272_1860_0) | (i_8_272_25_0 & ~i_8_272_94_0 & ~i_8_272_622_0 & ~i_8_272_987_0 & ~i_8_272_997_0 & i_8_272_1410_0 & ~i_8_272_2026_0))) | (i_8_272_423_0 & ((~i_8_272_623_0 & ~i_8_272_987_0 & i_8_272_1651_0 & ~i_8_272_1736_0) | (~i_8_272_778_0 & ~i_8_272_989_0 & i_8_272_1305_0 & ~i_8_272_1626_0 & ~i_8_272_1661_0 & i_8_272_1776_0 & ~i_8_272_1790_0))) | (~i_8_272_2025_0 & ((~i_8_272_94_0 & ((~i_8_272_593_0 & ~i_8_272_779_0 & ~i_8_272_2058_0 & ((~i_8_272_988_0 & ~i_8_272_1818_0 & i_8_272_1980_0) | (~i_8_272_625_0 & ~i_8_272_638_0 & i_8_272_703_0 & ~i_8_272_713_0 & ~i_8_272_720_0 & ~i_8_272_985_0 & ~i_8_272_1902_0 & ~i_8_272_2015_0))) | (i_8_272_606_0 & ~i_8_272_713_0 & ~i_8_272_973_0 & ~i_8_272_984_0 & ~i_8_272_1626_0 & ~i_8_272_1651_0 & i_8_272_1965_0))) | (~i_8_272_713_0 & ((i_8_272_379_0 & ~i_8_272_621_0 & ~i_8_272_988_0 & ~i_8_272_1273_0 & ~i_8_272_1623_0 & ~i_8_272_1776_0 & ~i_8_272_1857_0 & i_8_272_1965_0) | (~i_8_272_703_0 & ~i_8_272_934_0 & ~i_8_272_989_0 & ~i_8_272_1330_0 & ~i_8_272_1483_0 & ~i_8_272_1733_0 & i_8_272_1967_0 & ~i_8_272_2026_0 & ~i_8_272_2058_0))) | (~i_8_272_345_0 & ~i_8_272_383_0 & ~i_8_272_626_0 & ~i_8_272_988_0 & i_8_272_1967_0 & i_8_272_2237_0))) | (~i_8_272_720_0 & ((i_8_272_606_0 & ~i_8_272_986_0 & ((i_8_272_626_0 & ~i_8_272_779_0 & ~i_8_272_996_0 & ~i_8_272_1731_0) | (~i_8_272_612_0 & ~i_8_272_1307_0 & ~i_8_272_1626_0 & ~i_8_272_1736_0 & i_8_272_1776_0 & ~i_8_272_1857_0 & ~i_8_272_1902_0))) | (~i_8_272_713_0 & ((i_8_272_345_0 & i_8_272_626_0 & ~i_8_272_985_0 & i_8_272_1470_0 & ~i_8_272_1736_0) | (~i_8_272_1483_0 & ~i_8_272_1529_0 & ~i_8_272_1623_0 & ~i_8_272_1626_0 & ~i_8_272_2015_0 & i_8_272_2154_0 & i_8_272_2156_0))) | (~i_8_272_625_0 & i_8_272_703_0 & ~i_8_272_985_0 & ~i_8_272_997_0 & i_8_272_1297_0))) | (~i_8_272_996_0 & ((~i_8_272_625_0 & ((~i_8_272_713_0 & ~i_8_272_934_0 & ~i_8_272_1027_0 & i_8_272_1307_0 & i_8_272_1651_0) | (~i_8_272_704_0 & ~i_8_272_973_0 & ~i_8_272_984_0 & ~i_8_272_1621_0 & ~i_8_272_1626_0 & i_8_272_1950_0 & ~i_8_272_2015_0 & ~i_8_272_2154_0))) | (i_8_272_593_0 & ~i_8_272_608_0 & ~i_8_272_623_0 & ~i_8_272_704_0 & ~i_8_272_713_0 & ~i_8_272_988_0 & ~i_8_272_1123_0 & ~i_8_272_1733_0 & ~i_8_272_1902_0) | (~i_8_272_1626_0 & ~i_8_272_1731_0 & i_8_272_1752_0 & ~i_8_272_1789_0 & ~i_8_272_1860_0 & ~i_8_272_1862_0 & ~i_8_272_2058_0 & ~i_8_272_2076_0))) | (~i_8_272_778_0 & ((~i_8_272_592_0 & ~i_8_272_1623_0 & ~i_8_272_1651_0 & i_8_272_1965_0 & i_8_272_2070_0) | (~i_8_272_623_0 & ~i_8_272_985_0 & ~i_8_272_1857_0 & i_8_272_1967_0 & i_8_272_2156_0))) | (~i_8_272_623_0 & ((~i_8_272_622_0 & ~i_8_272_1027_0 & i_8_272_1273_0 & ~i_8_272_1626_0 & ~i_8_272_1860_0 & i_8_272_1471_0 & ~i_8_272_1526_0) | (i_8_272_703_0 & i_8_272_704_0 & i_8_272_985_0 & ~i_8_272_1307_0 & ~i_8_272_2015_0))) | (~i_8_272_622_0 & ~i_8_272_987_0 & ((i_8_272_462_0 & ~i_8_272_723_0 & ~i_8_272_985_0 & ~i_8_272_986_0 & ~i_8_272_997_0 & ~i_8_272_1857_0) | (~i_8_272_94_0 & ~i_8_272_705_0 & ~i_8_272_1626_0 & ~i_8_272_1733_0 & ~i_8_272_1902_0 & i_8_272_2076_0))) | (~i_8_272_997_0 & ~i_8_272_1862_0 & i_8_272_1950_0 & ~i_8_272_2058_0 & i_8_272_2154_0) | (~i_8_272_1027_0 & ~i_8_272_1623_0 & ~i_8_272_1731_0 & i_8_272_1857_0 & i_8_272_2169_0));
endmodule



// Benchmark "kernel_8_273" written by ABC on Sun Jul 19 10:07:50 2020

module kernel_8_273 ( 
    i_8_273_4_0, i_8_273_23_0, i_8_273_64_0, i_8_273_75_0, i_8_273_85_0,
    i_8_273_131_0, i_8_273_176_0, i_8_273_193_0, i_8_273_233_0,
    i_8_273_235_0, i_8_273_247_0, i_8_273_248_0, i_8_273_301_0,
    i_8_273_302_0, i_8_273_310_0, i_8_273_362_0, i_8_273_374_0,
    i_8_273_426_0, i_8_273_428_0, i_8_273_489_0, i_8_273_493_0,
    i_8_273_497_0, i_8_273_536_0, i_8_273_581_0, i_8_273_596_0,
    i_8_273_651_0, i_8_273_655_0, i_8_273_671_0, i_8_273_703_0,
    i_8_273_706_0, i_8_273_803_0, i_8_273_832_0, i_8_273_860_0,
    i_8_273_911_0, i_8_273_914_0, i_8_273_956_0, i_8_273_967_0,
    i_8_273_991_0, i_8_273_1030_0, i_8_273_1048_0, i_8_273_1085_0,
    i_8_273_1095_0, i_8_273_1112_0, i_8_273_1132_0, i_8_273_1135_0,
    i_8_273_1164_0, i_8_273_1190_0, i_8_273_1228_0, i_8_273_1271_0,
    i_8_273_1308_0, i_8_273_1324_0, i_8_273_1355_0, i_8_273_1397_0,
    i_8_273_1400_0, i_8_273_1405_0, i_8_273_1407_0, i_8_273_1408_0,
    i_8_273_1428_0, i_8_273_1468_0, i_8_273_1492_0, i_8_273_1493_0,
    i_8_273_1498_0, i_8_273_1532_0, i_8_273_1534_0, i_8_273_1535_0,
    i_8_273_1549_0, i_8_273_1632_0, i_8_273_1636_0, i_8_273_1642_0,
    i_8_273_1688_0, i_8_273_1781_0, i_8_273_1795_0, i_8_273_1804_0,
    i_8_273_1805_0, i_8_273_1807_0, i_8_273_1819_0, i_8_273_1821_0,
    i_8_273_1855_0, i_8_273_1868_0, i_8_273_1885_0, i_8_273_1905_0,
    i_8_273_1913_0, i_8_273_1919_0, i_8_273_1949_0, i_8_273_1992_0,
    i_8_273_1994_0, i_8_273_1996_0, i_8_273_2011_0, i_8_273_2047_0,
    i_8_273_2048_0, i_8_273_2063_0, i_8_273_2066_0, i_8_273_2119_0,
    i_8_273_2144_0, i_8_273_2145_0, i_8_273_2147_0, i_8_273_2149_0,
    i_8_273_2216_0, i_8_273_2234_0, i_8_273_2275_0,
    o_8_273_0_0  );
  input  i_8_273_4_0, i_8_273_23_0, i_8_273_64_0, i_8_273_75_0,
    i_8_273_85_0, i_8_273_131_0, i_8_273_176_0, i_8_273_193_0,
    i_8_273_233_0, i_8_273_235_0, i_8_273_247_0, i_8_273_248_0,
    i_8_273_301_0, i_8_273_302_0, i_8_273_310_0, i_8_273_362_0,
    i_8_273_374_0, i_8_273_426_0, i_8_273_428_0, i_8_273_489_0,
    i_8_273_493_0, i_8_273_497_0, i_8_273_536_0, i_8_273_581_0,
    i_8_273_596_0, i_8_273_651_0, i_8_273_655_0, i_8_273_671_0,
    i_8_273_703_0, i_8_273_706_0, i_8_273_803_0, i_8_273_832_0,
    i_8_273_860_0, i_8_273_911_0, i_8_273_914_0, i_8_273_956_0,
    i_8_273_967_0, i_8_273_991_0, i_8_273_1030_0, i_8_273_1048_0,
    i_8_273_1085_0, i_8_273_1095_0, i_8_273_1112_0, i_8_273_1132_0,
    i_8_273_1135_0, i_8_273_1164_0, i_8_273_1190_0, i_8_273_1228_0,
    i_8_273_1271_0, i_8_273_1308_0, i_8_273_1324_0, i_8_273_1355_0,
    i_8_273_1397_0, i_8_273_1400_0, i_8_273_1405_0, i_8_273_1407_0,
    i_8_273_1408_0, i_8_273_1428_0, i_8_273_1468_0, i_8_273_1492_0,
    i_8_273_1493_0, i_8_273_1498_0, i_8_273_1532_0, i_8_273_1534_0,
    i_8_273_1535_0, i_8_273_1549_0, i_8_273_1632_0, i_8_273_1636_0,
    i_8_273_1642_0, i_8_273_1688_0, i_8_273_1781_0, i_8_273_1795_0,
    i_8_273_1804_0, i_8_273_1805_0, i_8_273_1807_0, i_8_273_1819_0,
    i_8_273_1821_0, i_8_273_1855_0, i_8_273_1868_0, i_8_273_1885_0,
    i_8_273_1905_0, i_8_273_1913_0, i_8_273_1919_0, i_8_273_1949_0,
    i_8_273_1992_0, i_8_273_1994_0, i_8_273_1996_0, i_8_273_2011_0,
    i_8_273_2047_0, i_8_273_2048_0, i_8_273_2063_0, i_8_273_2066_0,
    i_8_273_2119_0, i_8_273_2144_0, i_8_273_2145_0, i_8_273_2147_0,
    i_8_273_2149_0, i_8_273_2216_0, i_8_273_2234_0, i_8_273_2275_0;
  output o_8_273_0_0;
  assign o_8_273_0_0 = 0;
endmodule



// Benchmark "kernel_8_274" written by ABC on Sun Jul 19 10:07:50 2020

module kernel_8_274 ( 
    i_8_274_27_0, i_8_274_28_0, i_8_274_217_0, i_8_274_254_0,
    i_8_274_257_0, i_8_274_299_0, i_8_274_305_0, i_8_274_316_0,
    i_8_274_323_0, i_8_274_368_0, i_8_274_381_0, i_8_274_428_0,
    i_8_274_454_0, i_8_274_470_0, i_8_274_488_0, i_8_274_572_0,
    i_8_274_587_0, i_8_274_595_0, i_8_274_610_0, i_8_274_631_0,
    i_8_274_632_0, i_8_274_649_0, i_8_274_678_0, i_8_274_695_0,
    i_8_274_697_0, i_8_274_778_0, i_8_274_779_0, i_8_274_796_0,
    i_8_274_833_0, i_8_274_839_0, i_8_274_844_0, i_8_274_847_0,
    i_8_274_848_0, i_8_274_856_0, i_8_274_860_0, i_8_274_868_0,
    i_8_274_874_0, i_8_274_875_0, i_8_274_877_0, i_8_274_878_0,
    i_8_274_883_0, i_8_274_965_0, i_8_274_969_0, i_8_274_1136_0,
    i_8_274_1216_0, i_8_274_1226_0, i_8_274_1228_0, i_8_274_1255_0,
    i_8_274_1262_0, i_8_274_1281_0, i_8_274_1285_0, i_8_274_1298_0,
    i_8_274_1355_0, i_8_274_1410_0, i_8_274_1442_0, i_8_274_1449_0,
    i_8_274_1514_0, i_8_274_1516_0, i_8_274_1526_0, i_8_274_1543_0,
    i_8_274_1544_0, i_8_274_1547_0, i_8_274_1559_0, i_8_274_1561_0,
    i_8_274_1607_0, i_8_274_1615_0, i_8_274_1621_0, i_8_274_1630_0,
    i_8_274_1631_0, i_8_274_1634_0, i_8_274_1675_0, i_8_274_1703_0,
    i_8_274_1704_0, i_8_274_1714_0, i_8_274_1720_0, i_8_274_1756_0,
    i_8_274_1757_0, i_8_274_1759_0, i_8_274_1776_0, i_8_274_1810_0,
    i_8_274_1882_0, i_8_274_1972_0, i_8_274_1982_0, i_8_274_1990_0,
    i_8_274_1994_0, i_8_274_2054_0, i_8_274_2099_0, i_8_274_2102_0,
    i_8_274_2134_0, i_8_274_2136_0, i_8_274_2140_0, i_8_274_2156_0,
    i_8_274_2170_0, i_8_274_2225_0, i_8_274_2242_0, i_8_274_2243_0,
    i_8_274_2263_0, i_8_274_2264_0, i_8_274_2270_0, i_8_274_2291_0,
    o_8_274_0_0  );
  input  i_8_274_27_0, i_8_274_28_0, i_8_274_217_0, i_8_274_254_0,
    i_8_274_257_0, i_8_274_299_0, i_8_274_305_0, i_8_274_316_0,
    i_8_274_323_0, i_8_274_368_0, i_8_274_381_0, i_8_274_428_0,
    i_8_274_454_0, i_8_274_470_0, i_8_274_488_0, i_8_274_572_0,
    i_8_274_587_0, i_8_274_595_0, i_8_274_610_0, i_8_274_631_0,
    i_8_274_632_0, i_8_274_649_0, i_8_274_678_0, i_8_274_695_0,
    i_8_274_697_0, i_8_274_778_0, i_8_274_779_0, i_8_274_796_0,
    i_8_274_833_0, i_8_274_839_0, i_8_274_844_0, i_8_274_847_0,
    i_8_274_848_0, i_8_274_856_0, i_8_274_860_0, i_8_274_868_0,
    i_8_274_874_0, i_8_274_875_0, i_8_274_877_0, i_8_274_878_0,
    i_8_274_883_0, i_8_274_965_0, i_8_274_969_0, i_8_274_1136_0,
    i_8_274_1216_0, i_8_274_1226_0, i_8_274_1228_0, i_8_274_1255_0,
    i_8_274_1262_0, i_8_274_1281_0, i_8_274_1285_0, i_8_274_1298_0,
    i_8_274_1355_0, i_8_274_1410_0, i_8_274_1442_0, i_8_274_1449_0,
    i_8_274_1514_0, i_8_274_1516_0, i_8_274_1526_0, i_8_274_1543_0,
    i_8_274_1544_0, i_8_274_1547_0, i_8_274_1559_0, i_8_274_1561_0,
    i_8_274_1607_0, i_8_274_1615_0, i_8_274_1621_0, i_8_274_1630_0,
    i_8_274_1631_0, i_8_274_1634_0, i_8_274_1675_0, i_8_274_1703_0,
    i_8_274_1704_0, i_8_274_1714_0, i_8_274_1720_0, i_8_274_1756_0,
    i_8_274_1757_0, i_8_274_1759_0, i_8_274_1776_0, i_8_274_1810_0,
    i_8_274_1882_0, i_8_274_1972_0, i_8_274_1982_0, i_8_274_1990_0,
    i_8_274_1994_0, i_8_274_2054_0, i_8_274_2099_0, i_8_274_2102_0,
    i_8_274_2134_0, i_8_274_2136_0, i_8_274_2140_0, i_8_274_2156_0,
    i_8_274_2170_0, i_8_274_2225_0, i_8_274_2242_0, i_8_274_2243_0,
    i_8_274_2263_0, i_8_274_2264_0, i_8_274_2270_0, i_8_274_2291_0;
  output o_8_274_0_0;
  assign o_8_274_0_0 = 0;
endmodule



// Benchmark "kernel_8_275" written by ABC on Sun Jul 19 10:07:51 2020

module kernel_8_275 ( 
    i_8_275_20_0, i_8_275_38_0, i_8_275_47_0, i_8_275_50_0, i_8_275_55_0,
    i_8_275_56_0, i_8_275_65_0, i_8_275_92_0, i_8_275_115_0, i_8_275_173_0,
    i_8_275_189_0, i_8_275_236_0, i_8_275_299_0, i_8_275_304_0,
    i_8_275_308_0, i_8_275_335_0, i_8_275_352_0, i_8_275_362_0,
    i_8_275_379_0, i_8_275_380_0, i_8_275_387_0, i_8_275_418_0,
    i_8_275_425_0, i_8_275_452_0, i_8_275_524_0, i_8_275_530_0,
    i_8_275_578_0, i_8_275_586_0, i_8_275_587_0, i_8_275_658_0,
    i_8_275_666_0, i_8_275_704_0, i_8_275_779_0, i_8_275_793_0,
    i_8_275_801_0, i_8_275_803_0, i_8_275_829_0, i_8_275_848_0,
    i_8_275_880_0, i_8_275_883_0, i_8_275_884_0, i_8_275_919_0,
    i_8_275_927_0, i_8_275_928_0, i_8_275_992_0, i_8_275_994_0,
    i_8_275_1033_0, i_8_275_1054_0, i_8_275_1079_0, i_8_275_1091_0,
    i_8_275_1129_0, i_8_275_1145_0, i_8_275_1163_0, i_8_275_1226_0,
    i_8_275_1271_0, i_8_275_1283_0, i_8_275_1289_0, i_8_275_1297_0,
    i_8_275_1328_0, i_8_275_1333_0, i_8_275_1405_0, i_8_275_1406_0,
    i_8_275_1459_0, i_8_275_1505_0, i_8_275_1559_0, i_8_275_1603_0,
    i_8_275_1604_0, i_8_275_1747_0, i_8_275_1817_0, i_8_275_1823_0,
    i_8_275_1862_0, i_8_275_1864_0, i_8_275_1865_0, i_8_275_1883_0,
    i_8_275_1884_0, i_8_275_1886_0, i_8_275_1907_0, i_8_275_1918_0,
    i_8_275_1937_0, i_8_275_1992_0, i_8_275_1993_0, i_8_275_2008_0,
    i_8_275_2026_0, i_8_275_2030_0, i_8_275_2045_0, i_8_275_2052_0,
    i_8_275_2054_0, i_8_275_2096_0, i_8_275_2107_0, i_8_275_2132_0,
    i_8_275_2144_0, i_8_275_2152_0, i_8_275_2153_0, i_8_275_2180_0,
    i_8_275_2196_0, i_8_275_2197_0, i_8_275_2206_0, i_8_275_2210_0,
    i_8_275_2227_0, i_8_275_2287_0,
    o_8_275_0_0  );
  input  i_8_275_20_0, i_8_275_38_0, i_8_275_47_0, i_8_275_50_0,
    i_8_275_55_0, i_8_275_56_0, i_8_275_65_0, i_8_275_92_0, i_8_275_115_0,
    i_8_275_173_0, i_8_275_189_0, i_8_275_236_0, i_8_275_299_0,
    i_8_275_304_0, i_8_275_308_0, i_8_275_335_0, i_8_275_352_0,
    i_8_275_362_0, i_8_275_379_0, i_8_275_380_0, i_8_275_387_0,
    i_8_275_418_0, i_8_275_425_0, i_8_275_452_0, i_8_275_524_0,
    i_8_275_530_0, i_8_275_578_0, i_8_275_586_0, i_8_275_587_0,
    i_8_275_658_0, i_8_275_666_0, i_8_275_704_0, i_8_275_779_0,
    i_8_275_793_0, i_8_275_801_0, i_8_275_803_0, i_8_275_829_0,
    i_8_275_848_0, i_8_275_880_0, i_8_275_883_0, i_8_275_884_0,
    i_8_275_919_0, i_8_275_927_0, i_8_275_928_0, i_8_275_992_0,
    i_8_275_994_0, i_8_275_1033_0, i_8_275_1054_0, i_8_275_1079_0,
    i_8_275_1091_0, i_8_275_1129_0, i_8_275_1145_0, i_8_275_1163_0,
    i_8_275_1226_0, i_8_275_1271_0, i_8_275_1283_0, i_8_275_1289_0,
    i_8_275_1297_0, i_8_275_1328_0, i_8_275_1333_0, i_8_275_1405_0,
    i_8_275_1406_0, i_8_275_1459_0, i_8_275_1505_0, i_8_275_1559_0,
    i_8_275_1603_0, i_8_275_1604_0, i_8_275_1747_0, i_8_275_1817_0,
    i_8_275_1823_0, i_8_275_1862_0, i_8_275_1864_0, i_8_275_1865_0,
    i_8_275_1883_0, i_8_275_1884_0, i_8_275_1886_0, i_8_275_1907_0,
    i_8_275_1918_0, i_8_275_1937_0, i_8_275_1992_0, i_8_275_1993_0,
    i_8_275_2008_0, i_8_275_2026_0, i_8_275_2030_0, i_8_275_2045_0,
    i_8_275_2052_0, i_8_275_2054_0, i_8_275_2096_0, i_8_275_2107_0,
    i_8_275_2132_0, i_8_275_2144_0, i_8_275_2152_0, i_8_275_2153_0,
    i_8_275_2180_0, i_8_275_2196_0, i_8_275_2197_0, i_8_275_2206_0,
    i_8_275_2210_0, i_8_275_2227_0, i_8_275_2287_0;
  output o_8_275_0_0;
  assign o_8_275_0_0 = ~(~i_8_275_2180_0 | (~i_8_275_1907_0 & ~i_8_275_2287_0) | (~i_8_275_927_0 & ~i_8_275_1823_0) | (i_8_275_848_0 & i_8_275_1079_0) | (~i_8_275_793_0 & ~i_8_275_2052_0 & ~i_8_275_2206_0) | (~i_8_275_55_0 & ~i_8_275_173_0 & ~i_8_275_2132_0));
endmodule



// Benchmark "kernel_8_276" written by ABC on Sun Jul 19 10:07:52 2020

module kernel_8_276 ( 
    i_8_276_14_0, i_8_276_26_0, i_8_276_27_0, i_8_276_54_0, i_8_276_57_0,
    i_8_276_87_0, i_8_276_168_0, i_8_276_169_0, i_8_276_189_0,
    i_8_276_228_0, i_8_276_259_0, i_8_276_300_0, i_8_276_338_0,
    i_8_276_344_0, i_8_276_346_0, i_8_276_360_0, i_8_276_383_0,
    i_8_276_403_0, i_8_276_427_0, i_8_276_428_0, i_8_276_455_0,
    i_8_276_555_0, i_8_276_574_0, i_8_276_635_0, i_8_276_659_0,
    i_8_276_694_0, i_8_276_700_0, i_8_276_705_0, i_8_276_706_0,
    i_8_276_708_0, i_8_276_762_0, i_8_276_791_0, i_8_276_798_0,
    i_8_276_799_0, i_8_276_874_0, i_8_276_920_0, i_8_276_929_0,
    i_8_276_997_0, i_8_276_998_0, i_8_276_1077_0, i_8_276_1103_0,
    i_8_276_1105_0, i_8_276_1192_0, i_8_276_1195_0, i_8_276_1239_0,
    i_8_276_1260_0, i_8_276_1265_0, i_8_276_1276_0, i_8_276_1283_0,
    i_8_276_1288_0, i_8_276_1289_0, i_8_276_1299_0, i_8_276_1308_0,
    i_8_276_1309_0, i_8_276_1318_0, i_8_276_1321_0, i_8_276_1348_0,
    i_8_276_1382_0, i_8_276_1385_0, i_8_276_1393_0, i_8_276_1410_0,
    i_8_276_1436_0, i_8_276_1451_0, i_8_276_1470_0, i_8_276_1549_0,
    i_8_276_1590_0, i_8_276_1591_0, i_8_276_1592_0, i_8_276_1623_0,
    i_8_276_1625_0, i_8_276_1639_0, i_8_276_1642_0, i_8_276_1649_0,
    i_8_276_1690_0, i_8_276_1743_0, i_8_276_1762_0, i_8_276_1823_0,
    i_8_276_1826_0, i_8_276_1885_0, i_8_276_1888_0, i_8_276_1940_0,
    i_8_276_1986_0, i_8_276_1993_0, i_8_276_2040_0, i_8_276_2055_0,
    i_8_276_2056_0, i_8_276_2059_0, i_8_276_2077_0, i_8_276_2132_0,
    i_8_276_2147_0, i_8_276_2177_0, i_8_276_2200_0, i_8_276_2210_0,
    i_8_276_2213_0, i_8_276_2217_0, i_8_276_2219_0, i_8_276_2239_0,
    i_8_276_2240_0, i_8_276_2301_0, i_8_276_2302_0,
    o_8_276_0_0  );
  input  i_8_276_14_0, i_8_276_26_0, i_8_276_27_0, i_8_276_54_0,
    i_8_276_57_0, i_8_276_87_0, i_8_276_168_0, i_8_276_169_0,
    i_8_276_189_0, i_8_276_228_0, i_8_276_259_0, i_8_276_300_0,
    i_8_276_338_0, i_8_276_344_0, i_8_276_346_0, i_8_276_360_0,
    i_8_276_383_0, i_8_276_403_0, i_8_276_427_0, i_8_276_428_0,
    i_8_276_455_0, i_8_276_555_0, i_8_276_574_0, i_8_276_635_0,
    i_8_276_659_0, i_8_276_694_0, i_8_276_700_0, i_8_276_705_0,
    i_8_276_706_0, i_8_276_708_0, i_8_276_762_0, i_8_276_791_0,
    i_8_276_798_0, i_8_276_799_0, i_8_276_874_0, i_8_276_920_0,
    i_8_276_929_0, i_8_276_997_0, i_8_276_998_0, i_8_276_1077_0,
    i_8_276_1103_0, i_8_276_1105_0, i_8_276_1192_0, i_8_276_1195_0,
    i_8_276_1239_0, i_8_276_1260_0, i_8_276_1265_0, i_8_276_1276_0,
    i_8_276_1283_0, i_8_276_1288_0, i_8_276_1289_0, i_8_276_1299_0,
    i_8_276_1308_0, i_8_276_1309_0, i_8_276_1318_0, i_8_276_1321_0,
    i_8_276_1348_0, i_8_276_1382_0, i_8_276_1385_0, i_8_276_1393_0,
    i_8_276_1410_0, i_8_276_1436_0, i_8_276_1451_0, i_8_276_1470_0,
    i_8_276_1549_0, i_8_276_1590_0, i_8_276_1591_0, i_8_276_1592_0,
    i_8_276_1623_0, i_8_276_1625_0, i_8_276_1639_0, i_8_276_1642_0,
    i_8_276_1649_0, i_8_276_1690_0, i_8_276_1743_0, i_8_276_1762_0,
    i_8_276_1823_0, i_8_276_1826_0, i_8_276_1885_0, i_8_276_1888_0,
    i_8_276_1940_0, i_8_276_1986_0, i_8_276_1993_0, i_8_276_2040_0,
    i_8_276_2055_0, i_8_276_2056_0, i_8_276_2059_0, i_8_276_2077_0,
    i_8_276_2132_0, i_8_276_2147_0, i_8_276_2177_0, i_8_276_2200_0,
    i_8_276_2210_0, i_8_276_2213_0, i_8_276_2217_0, i_8_276_2219_0,
    i_8_276_2239_0, i_8_276_2240_0, i_8_276_2301_0, i_8_276_2302_0;
  output o_8_276_0_0;
  assign o_8_276_0_0 = 0;
endmodule



// Benchmark "kernel_8_277" written by ABC on Sun Jul 19 10:07:53 2020

module kernel_8_277 ( 
    i_8_277_13_0, i_8_277_74_0, i_8_277_79_0, i_8_277_103_0, i_8_277_114_0,
    i_8_277_115_0, i_8_277_116_0, i_8_277_137_0, i_8_277_184_0,
    i_8_277_190_0, i_8_277_196_0, i_8_277_233_0, i_8_277_284_0,
    i_8_277_301_0, i_8_277_319_0, i_8_277_320_0, i_8_277_326_0,
    i_8_277_343_0, i_8_277_366_0, i_8_277_427_0, i_8_277_434_0,
    i_8_277_450_0, i_8_277_493_0, i_8_277_525_0, i_8_277_526_0,
    i_8_277_544_0, i_8_277_640_0, i_8_277_660_0, i_8_277_665_0,
    i_8_277_703_0, i_8_277_748_0, i_8_277_782_0, i_8_277_799_0,
    i_8_277_800_0, i_8_277_854_0, i_8_277_880_0, i_8_277_946_0,
    i_8_277_965_0, i_8_277_971_0, i_8_277_977_0, i_8_277_992_0,
    i_8_277_1051_0, i_8_277_1061_0, i_8_277_1110_0, i_8_277_1114_0,
    i_8_277_1228_0, i_8_277_1236_0, i_8_277_1246_0, i_8_277_1263_0,
    i_8_277_1294_0, i_8_277_1295_0, i_8_277_1316_0, i_8_277_1325_0,
    i_8_277_1328_0, i_8_277_1354_0, i_8_277_1363_0, i_8_277_1364_0,
    i_8_277_1417_0, i_8_277_1424_0, i_8_277_1432_0, i_8_277_1441_0,
    i_8_277_1462_0, i_8_277_1463_0, i_8_277_1468_0, i_8_277_1517_0,
    i_8_277_1522_0, i_8_277_1538_0, i_8_277_1552_0, i_8_277_1561_0,
    i_8_277_1614_0, i_8_277_1624_0, i_8_277_1651_0, i_8_277_1678_0,
    i_8_277_1694_0, i_8_277_1702_0, i_8_277_1730_0, i_8_277_1746_0,
    i_8_277_1747_0, i_8_277_1819_0, i_8_277_1855_0, i_8_277_1859_0,
    i_8_277_1913_0, i_8_277_1930_0, i_8_277_1939_0, i_8_277_1964_0,
    i_8_277_1982_0, i_8_277_1995_0, i_8_277_2008_0, i_8_277_2047_0,
    i_8_277_2074_0, i_8_277_2143_0, i_8_277_2149_0, i_8_277_2153_0,
    i_8_277_2156_0, i_8_277_2161_0, i_8_277_2170_0, i_8_277_2225_0,
    i_8_277_2245_0, i_8_277_2247_0, i_8_277_2249_0,
    o_8_277_0_0  );
  input  i_8_277_13_0, i_8_277_74_0, i_8_277_79_0, i_8_277_103_0,
    i_8_277_114_0, i_8_277_115_0, i_8_277_116_0, i_8_277_137_0,
    i_8_277_184_0, i_8_277_190_0, i_8_277_196_0, i_8_277_233_0,
    i_8_277_284_0, i_8_277_301_0, i_8_277_319_0, i_8_277_320_0,
    i_8_277_326_0, i_8_277_343_0, i_8_277_366_0, i_8_277_427_0,
    i_8_277_434_0, i_8_277_450_0, i_8_277_493_0, i_8_277_525_0,
    i_8_277_526_0, i_8_277_544_0, i_8_277_640_0, i_8_277_660_0,
    i_8_277_665_0, i_8_277_703_0, i_8_277_748_0, i_8_277_782_0,
    i_8_277_799_0, i_8_277_800_0, i_8_277_854_0, i_8_277_880_0,
    i_8_277_946_0, i_8_277_965_0, i_8_277_971_0, i_8_277_977_0,
    i_8_277_992_0, i_8_277_1051_0, i_8_277_1061_0, i_8_277_1110_0,
    i_8_277_1114_0, i_8_277_1228_0, i_8_277_1236_0, i_8_277_1246_0,
    i_8_277_1263_0, i_8_277_1294_0, i_8_277_1295_0, i_8_277_1316_0,
    i_8_277_1325_0, i_8_277_1328_0, i_8_277_1354_0, i_8_277_1363_0,
    i_8_277_1364_0, i_8_277_1417_0, i_8_277_1424_0, i_8_277_1432_0,
    i_8_277_1441_0, i_8_277_1462_0, i_8_277_1463_0, i_8_277_1468_0,
    i_8_277_1517_0, i_8_277_1522_0, i_8_277_1538_0, i_8_277_1552_0,
    i_8_277_1561_0, i_8_277_1614_0, i_8_277_1624_0, i_8_277_1651_0,
    i_8_277_1678_0, i_8_277_1694_0, i_8_277_1702_0, i_8_277_1730_0,
    i_8_277_1746_0, i_8_277_1747_0, i_8_277_1819_0, i_8_277_1855_0,
    i_8_277_1859_0, i_8_277_1913_0, i_8_277_1930_0, i_8_277_1939_0,
    i_8_277_1964_0, i_8_277_1982_0, i_8_277_1995_0, i_8_277_2008_0,
    i_8_277_2047_0, i_8_277_2074_0, i_8_277_2143_0, i_8_277_2149_0,
    i_8_277_2153_0, i_8_277_2156_0, i_8_277_2161_0, i_8_277_2170_0,
    i_8_277_2225_0, i_8_277_2245_0, i_8_277_2247_0, i_8_277_2249_0;
  output o_8_277_0_0;
  assign o_8_277_0_0 = 0;
endmodule



// Benchmark "kernel_8_278" written by ABC on Sun Jul 19 10:07:54 2020

module kernel_8_278 ( 
    i_8_278_19_0, i_8_278_25_0, i_8_278_35_0, i_8_278_48_0, i_8_278_93_0,
    i_8_278_139_0, i_8_278_141_0, i_8_278_142_0, i_8_278_246_0,
    i_8_278_310_0, i_8_278_349_0, i_8_278_453_0, i_8_278_455_0,
    i_8_278_481_0, i_8_278_485_0, i_8_278_491_0, i_8_278_522_0,
    i_8_278_525_0, i_8_278_526_0, i_8_278_527_0, i_8_278_529_0,
    i_8_278_530_0, i_8_278_535_0, i_8_278_544_0, i_8_278_546_0,
    i_8_278_563_0, i_8_278_593_0, i_8_278_625_0, i_8_278_638_0,
    i_8_278_655_0, i_8_278_661_0, i_8_278_691_0, i_8_278_693_0,
    i_8_278_697_0, i_8_278_739_0, i_8_278_762_0, i_8_278_763_0,
    i_8_278_764_0, i_8_278_771_0, i_8_278_825_0, i_8_278_874_0,
    i_8_278_882_0, i_8_278_943_0, i_8_278_949_0, i_8_278_968_0,
    i_8_278_994_0, i_8_278_996_0, i_8_278_1056_0, i_8_278_1059_0,
    i_8_278_1063_0, i_8_278_1066_0, i_8_278_1067_0, i_8_278_1129_0,
    i_8_278_1135_0, i_8_278_1138_0, i_8_278_1180_0, i_8_278_1192_0,
    i_8_278_1219_0, i_8_278_1237_0, i_8_278_1260_0, i_8_278_1268_0,
    i_8_278_1305_0, i_8_278_1306_0, i_8_278_1307_0, i_8_278_1308_0,
    i_8_278_1315_0, i_8_278_1322_0, i_8_278_1323_0, i_8_278_1421_0,
    i_8_278_1431_0, i_8_278_1510_0, i_8_278_1547_0, i_8_278_1564_0,
    i_8_278_1574_0, i_8_278_1606_0, i_8_278_1651_0, i_8_278_1670_0,
    i_8_278_1682_0, i_8_278_1696_0, i_8_278_1723_0, i_8_278_1732_0,
    i_8_278_1751_0, i_8_278_1752_0, i_8_278_1762_0, i_8_278_1795_0,
    i_8_278_1807_0, i_8_278_1842_0, i_8_278_1848_0, i_8_278_1885_0,
    i_8_278_1918_0, i_8_278_1947_0, i_8_278_1980_0, i_8_278_1994_0,
    i_8_278_2014_0, i_8_278_2150_0, i_8_278_2177_0, i_8_278_2183_0,
    i_8_278_2214_0, i_8_278_2223_0, i_8_278_2263_0,
    o_8_278_0_0  );
  input  i_8_278_19_0, i_8_278_25_0, i_8_278_35_0, i_8_278_48_0,
    i_8_278_93_0, i_8_278_139_0, i_8_278_141_0, i_8_278_142_0,
    i_8_278_246_0, i_8_278_310_0, i_8_278_349_0, i_8_278_453_0,
    i_8_278_455_0, i_8_278_481_0, i_8_278_485_0, i_8_278_491_0,
    i_8_278_522_0, i_8_278_525_0, i_8_278_526_0, i_8_278_527_0,
    i_8_278_529_0, i_8_278_530_0, i_8_278_535_0, i_8_278_544_0,
    i_8_278_546_0, i_8_278_563_0, i_8_278_593_0, i_8_278_625_0,
    i_8_278_638_0, i_8_278_655_0, i_8_278_661_0, i_8_278_691_0,
    i_8_278_693_0, i_8_278_697_0, i_8_278_739_0, i_8_278_762_0,
    i_8_278_763_0, i_8_278_764_0, i_8_278_771_0, i_8_278_825_0,
    i_8_278_874_0, i_8_278_882_0, i_8_278_943_0, i_8_278_949_0,
    i_8_278_968_0, i_8_278_994_0, i_8_278_996_0, i_8_278_1056_0,
    i_8_278_1059_0, i_8_278_1063_0, i_8_278_1066_0, i_8_278_1067_0,
    i_8_278_1129_0, i_8_278_1135_0, i_8_278_1138_0, i_8_278_1180_0,
    i_8_278_1192_0, i_8_278_1219_0, i_8_278_1237_0, i_8_278_1260_0,
    i_8_278_1268_0, i_8_278_1305_0, i_8_278_1306_0, i_8_278_1307_0,
    i_8_278_1308_0, i_8_278_1315_0, i_8_278_1322_0, i_8_278_1323_0,
    i_8_278_1421_0, i_8_278_1431_0, i_8_278_1510_0, i_8_278_1547_0,
    i_8_278_1564_0, i_8_278_1574_0, i_8_278_1606_0, i_8_278_1651_0,
    i_8_278_1670_0, i_8_278_1682_0, i_8_278_1696_0, i_8_278_1723_0,
    i_8_278_1732_0, i_8_278_1751_0, i_8_278_1752_0, i_8_278_1762_0,
    i_8_278_1795_0, i_8_278_1807_0, i_8_278_1842_0, i_8_278_1848_0,
    i_8_278_1885_0, i_8_278_1918_0, i_8_278_1947_0, i_8_278_1980_0,
    i_8_278_1994_0, i_8_278_2014_0, i_8_278_2150_0, i_8_278_2177_0,
    i_8_278_2183_0, i_8_278_2214_0, i_8_278_2223_0, i_8_278_2263_0;
  output o_8_278_0_0;
  assign o_8_278_0_0 = 0;
endmodule



// Benchmark "kernel_8_279" written by ABC on Sun Jul 19 10:07:55 2020

module kernel_8_279 ( 
    i_8_279_22_0, i_8_279_95_0, i_8_279_135_0, i_8_279_140_0,
    i_8_279_208_0, i_8_279_325_0, i_8_279_337_0, i_8_279_426_0,
    i_8_279_450_0, i_8_279_459_0, i_8_279_484_0, i_8_279_496_0,
    i_8_279_497_0, i_8_279_500_0, i_8_279_525_0, i_8_279_528_0,
    i_8_279_539_0, i_8_279_544_0, i_8_279_545_0, i_8_279_551_0,
    i_8_279_557_0, i_8_279_649_0, i_8_279_658_0, i_8_279_668_0,
    i_8_279_669_0, i_8_279_675_0, i_8_279_708_0, i_8_279_720_0,
    i_8_279_760_0, i_8_279_762_0, i_8_279_779_0, i_8_279_820_0,
    i_8_279_842_0, i_8_279_846_0, i_8_279_867_0, i_8_279_875_0,
    i_8_279_956_0, i_8_279_989_0, i_8_279_1010_0, i_8_279_1028_0,
    i_8_279_1107_0, i_8_279_1108_0, i_8_279_1109_0, i_8_279_1112_0,
    i_8_279_1151_0, i_8_279_1180_0, i_8_279_1231_0, i_8_279_1260_0,
    i_8_279_1263_0, i_8_279_1270_0, i_8_279_1279_0, i_8_279_1304_0,
    i_8_279_1315_0, i_8_279_1316_0, i_8_279_1324_0, i_8_279_1338_0,
    i_8_279_1343_0, i_8_279_1432_0, i_8_279_1435_0, i_8_279_1526_0,
    i_8_279_1534_0, i_8_279_1536_0, i_8_279_1537_0, i_8_279_1549_0,
    i_8_279_1565_0, i_8_279_1579_0, i_8_279_1585_0, i_8_279_1618_0,
    i_8_279_1619_0, i_8_279_1630_0, i_8_279_1662_0, i_8_279_1665_0,
    i_8_279_1679_0, i_8_279_1682_0, i_8_279_1705_0, i_8_279_1732_0,
    i_8_279_1735_0, i_8_279_1747_0, i_8_279_1754_0, i_8_279_1787_0,
    i_8_279_1790_0, i_8_279_1805_0, i_8_279_1821_0, i_8_279_1867_0,
    i_8_279_1887_0, i_8_279_1888_0, i_8_279_1898_0, i_8_279_1920_0,
    i_8_279_2013_0, i_8_279_2047_0, i_8_279_2073_0, i_8_279_2086_0,
    i_8_279_2087_0, i_8_279_2105_0, i_8_279_2141_0, i_8_279_2146_0,
    i_8_279_2216_0, i_8_279_2266_0, i_8_279_2288_0, i_8_279_2302_0,
    o_8_279_0_0  );
  input  i_8_279_22_0, i_8_279_95_0, i_8_279_135_0, i_8_279_140_0,
    i_8_279_208_0, i_8_279_325_0, i_8_279_337_0, i_8_279_426_0,
    i_8_279_450_0, i_8_279_459_0, i_8_279_484_0, i_8_279_496_0,
    i_8_279_497_0, i_8_279_500_0, i_8_279_525_0, i_8_279_528_0,
    i_8_279_539_0, i_8_279_544_0, i_8_279_545_0, i_8_279_551_0,
    i_8_279_557_0, i_8_279_649_0, i_8_279_658_0, i_8_279_668_0,
    i_8_279_669_0, i_8_279_675_0, i_8_279_708_0, i_8_279_720_0,
    i_8_279_760_0, i_8_279_762_0, i_8_279_779_0, i_8_279_820_0,
    i_8_279_842_0, i_8_279_846_0, i_8_279_867_0, i_8_279_875_0,
    i_8_279_956_0, i_8_279_989_0, i_8_279_1010_0, i_8_279_1028_0,
    i_8_279_1107_0, i_8_279_1108_0, i_8_279_1109_0, i_8_279_1112_0,
    i_8_279_1151_0, i_8_279_1180_0, i_8_279_1231_0, i_8_279_1260_0,
    i_8_279_1263_0, i_8_279_1270_0, i_8_279_1279_0, i_8_279_1304_0,
    i_8_279_1315_0, i_8_279_1316_0, i_8_279_1324_0, i_8_279_1338_0,
    i_8_279_1343_0, i_8_279_1432_0, i_8_279_1435_0, i_8_279_1526_0,
    i_8_279_1534_0, i_8_279_1536_0, i_8_279_1537_0, i_8_279_1549_0,
    i_8_279_1565_0, i_8_279_1579_0, i_8_279_1585_0, i_8_279_1618_0,
    i_8_279_1619_0, i_8_279_1630_0, i_8_279_1662_0, i_8_279_1665_0,
    i_8_279_1679_0, i_8_279_1682_0, i_8_279_1705_0, i_8_279_1732_0,
    i_8_279_1735_0, i_8_279_1747_0, i_8_279_1754_0, i_8_279_1787_0,
    i_8_279_1790_0, i_8_279_1805_0, i_8_279_1821_0, i_8_279_1867_0,
    i_8_279_1887_0, i_8_279_1888_0, i_8_279_1898_0, i_8_279_1920_0,
    i_8_279_2013_0, i_8_279_2047_0, i_8_279_2073_0, i_8_279_2086_0,
    i_8_279_2087_0, i_8_279_2105_0, i_8_279_2141_0, i_8_279_2146_0,
    i_8_279_2216_0, i_8_279_2266_0, i_8_279_2288_0, i_8_279_2302_0;
  output o_8_279_0_0;
  assign o_8_279_0_0 = 0;
endmodule



// Benchmark "kernel_8_280" written by ABC on Sun Jul 19 10:07:56 2020

module kernel_8_280 ( 
    i_8_280_23_0, i_8_280_77_0, i_8_280_85_0, i_8_280_119_0, i_8_280_137_0,
    i_8_280_163_0, i_8_280_244_0, i_8_280_247_0, i_8_280_266_0,
    i_8_280_274_0, i_8_280_311_0, i_8_280_353_0, i_8_280_388_0,
    i_8_280_389_0, i_8_280_418_0, i_8_280_460_0, i_8_280_523_0,
    i_8_280_524_0, i_8_280_536_0, i_8_280_550_0, i_8_280_581_0,
    i_8_280_605_0, i_8_280_632_0, i_8_280_635_0, i_8_280_640_0,
    i_8_280_641_0, i_8_280_653_0, i_8_280_670_0, i_8_280_685_0,
    i_8_280_694_0, i_8_280_728_0, i_8_280_733_0, i_8_280_802_0,
    i_8_280_831_0, i_8_280_838_0, i_8_280_841_0, i_8_280_859_0,
    i_8_280_883_0, i_8_280_977_0, i_8_280_991_0, i_8_280_992_0,
    i_8_280_1054_0, i_8_280_1172_0, i_8_280_1199_0, i_8_280_1225_0,
    i_8_280_1243_0, i_8_280_1246_0, i_8_280_1247_0, i_8_280_1263_0,
    i_8_280_1279_0, i_8_280_1319_0, i_8_280_1354_0, i_8_280_1355_0,
    i_8_280_1388_0, i_8_280_1405_0, i_8_280_1408_0, i_8_280_1468_0,
    i_8_280_1486_0, i_8_280_1487_0, i_8_280_1496_0, i_8_280_1506_0,
    i_8_280_1507_0, i_8_280_1531_0, i_8_280_1542_0, i_8_280_1544_0,
    i_8_280_1595_0, i_8_280_1634_0, i_8_280_1648_0, i_8_280_1702_0,
    i_8_280_1748_0, i_8_280_1780_0, i_8_280_1801_0, i_8_280_1805_0,
    i_8_280_1818_0, i_8_280_1822_0, i_8_280_1847_0, i_8_280_1885_0,
    i_8_280_1913_0, i_8_280_1939_0, i_8_280_1940_0, i_8_280_1966_0,
    i_8_280_1980_0, i_8_280_1981_0, i_8_280_1993_0, i_8_280_2009_0,
    i_8_280_2038_0, i_8_280_2045_0, i_8_280_2052_0, i_8_280_2062_0,
    i_8_280_2065_0, i_8_280_2089_0, i_8_280_2122_0, i_8_280_2123_0,
    i_8_280_2149_0, i_8_280_2152_0, i_8_280_2227_0, i_8_280_2228_0,
    i_8_280_2241_0, i_8_280_2254_0, i_8_280_2256_0,
    o_8_280_0_0  );
  input  i_8_280_23_0, i_8_280_77_0, i_8_280_85_0, i_8_280_119_0,
    i_8_280_137_0, i_8_280_163_0, i_8_280_244_0, i_8_280_247_0,
    i_8_280_266_0, i_8_280_274_0, i_8_280_311_0, i_8_280_353_0,
    i_8_280_388_0, i_8_280_389_0, i_8_280_418_0, i_8_280_460_0,
    i_8_280_523_0, i_8_280_524_0, i_8_280_536_0, i_8_280_550_0,
    i_8_280_581_0, i_8_280_605_0, i_8_280_632_0, i_8_280_635_0,
    i_8_280_640_0, i_8_280_641_0, i_8_280_653_0, i_8_280_670_0,
    i_8_280_685_0, i_8_280_694_0, i_8_280_728_0, i_8_280_733_0,
    i_8_280_802_0, i_8_280_831_0, i_8_280_838_0, i_8_280_841_0,
    i_8_280_859_0, i_8_280_883_0, i_8_280_977_0, i_8_280_991_0,
    i_8_280_992_0, i_8_280_1054_0, i_8_280_1172_0, i_8_280_1199_0,
    i_8_280_1225_0, i_8_280_1243_0, i_8_280_1246_0, i_8_280_1247_0,
    i_8_280_1263_0, i_8_280_1279_0, i_8_280_1319_0, i_8_280_1354_0,
    i_8_280_1355_0, i_8_280_1388_0, i_8_280_1405_0, i_8_280_1408_0,
    i_8_280_1468_0, i_8_280_1486_0, i_8_280_1487_0, i_8_280_1496_0,
    i_8_280_1506_0, i_8_280_1507_0, i_8_280_1531_0, i_8_280_1542_0,
    i_8_280_1544_0, i_8_280_1595_0, i_8_280_1634_0, i_8_280_1648_0,
    i_8_280_1702_0, i_8_280_1748_0, i_8_280_1780_0, i_8_280_1801_0,
    i_8_280_1805_0, i_8_280_1818_0, i_8_280_1822_0, i_8_280_1847_0,
    i_8_280_1885_0, i_8_280_1913_0, i_8_280_1939_0, i_8_280_1940_0,
    i_8_280_1966_0, i_8_280_1980_0, i_8_280_1981_0, i_8_280_1993_0,
    i_8_280_2009_0, i_8_280_2038_0, i_8_280_2045_0, i_8_280_2052_0,
    i_8_280_2062_0, i_8_280_2065_0, i_8_280_2089_0, i_8_280_2122_0,
    i_8_280_2123_0, i_8_280_2149_0, i_8_280_2152_0, i_8_280_2227_0,
    i_8_280_2228_0, i_8_280_2241_0, i_8_280_2254_0, i_8_280_2256_0;
  output o_8_280_0_0;
  assign o_8_280_0_0 = 0;
endmodule



// Benchmark "kernel_8_281" written by ABC on Sun Jul 19 10:07:57 2020

module kernel_8_281 ( 
    i_8_281_24_0, i_8_281_25_0, i_8_281_52_0, i_8_281_62_0, i_8_281_76_0,
    i_8_281_169_0, i_8_281_204_0, i_8_281_223_0, i_8_281_328_0,
    i_8_281_333_0, i_8_281_348_0, i_8_281_376_0, i_8_281_384_0,
    i_8_281_400_0, i_8_281_429_0, i_8_281_455_0, i_8_281_490_0,
    i_8_281_494_0, i_8_281_503_0, i_8_281_522_0, i_8_281_526_0,
    i_8_281_574_0, i_8_281_583_0, i_8_281_588_0, i_8_281_592_0,
    i_8_281_608_0, i_8_281_613_0, i_8_281_616_0, i_8_281_642_0,
    i_8_281_661_0, i_8_281_750_0, i_8_281_754_0, i_8_281_759_0,
    i_8_281_771_0, i_8_281_773_0, i_8_281_789_0, i_8_281_845_0,
    i_8_281_854_0, i_8_281_895_0, i_8_281_941_0, i_8_281_944_0,
    i_8_281_966_0, i_8_281_998_0, i_8_281_1050_0, i_8_281_1086_0,
    i_8_281_1110_0, i_8_281_1111_0, i_8_281_1113_0, i_8_281_1114_0,
    i_8_281_1120_0, i_8_281_1123_0, i_8_281_1162_0, i_8_281_1265_0,
    i_8_281_1305_0, i_8_281_1308_0, i_8_281_1321_0, i_8_281_1331_0,
    i_8_281_1339_0, i_8_281_1348_0, i_8_281_1383_0, i_8_281_1399_0,
    i_8_281_1425_0, i_8_281_1426_0, i_8_281_1429_0, i_8_281_1471_0,
    i_8_281_1474_0, i_8_281_1509_0, i_8_281_1510_0, i_8_281_1527_0,
    i_8_281_1564_0, i_8_281_1565_0, i_8_281_1570_0, i_8_281_1588_0,
    i_8_281_1635_0, i_8_281_1636_0, i_8_281_1650_0, i_8_281_1651_0,
    i_8_281_1654_0, i_8_281_1689_0, i_8_281_1704_0, i_8_281_1752_0,
    i_8_281_1821_0, i_8_281_1822_0, i_8_281_1858_0, i_8_281_1860_0,
    i_8_281_1870_0, i_8_281_1876_0, i_8_281_1897_0, i_8_281_1906_0,
    i_8_281_1907_0, i_8_281_1978_0, i_8_281_1993_0, i_8_281_2041_0,
    i_8_281_2074_0, i_8_281_2091_0, i_8_281_2093_0, i_8_281_2215_0,
    i_8_281_2217_0, i_8_281_2227_0, i_8_281_2235_0,
    o_8_281_0_0  );
  input  i_8_281_24_0, i_8_281_25_0, i_8_281_52_0, i_8_281_62_0,
    i_8_281_76_0, i_8_281_169_0, i_8_281_204_0, i_8_281_223_0,
    i_8_281_328_0, i_8_281_333_0, i_8_281_348_0, i_8_281_376_0,
    i_8_281_384_0, i_8_281_400_0, i_8_281_429_0, i_8_281_455_0,
    i_8_281_490_0, i_8_281_494_0, i_8_281_503_0, i_8_281_522_0,
    i_8_281_526_0, i_8_281_574_0, i_8_281_583_0, i_8_281_588_0,
    i_8_281_592_0, i_8_281_608_0, i_8_281_613_0, i_8_281_616_0,
    i_8_281_642_0, i_8_281_661_0, i_8_281_750_0, i_8_281_754_0,
    i_8_281_759_0, i_8_281_771_0, i_8_281_773_0, i_8_281_789_0,
    i_8_281_845_0, i_8_281_854_0, i_8_281_895_0, i_8_281_941_0,
    i_8_281_944_0, i_8_281_966_0, i_8_281_998_0, i_8_281_1050_0,
    i_8_281_1086_0, i_8_281_1110_0, i_8_281_1111_0, i_8_281_1113_0,
    i_8_281_1114_0, i_8_281_1120_0, i_8_281_1123_0, i_8_281_1162_0,
    i_8_281_1265_0, i_8_281_1305_0, i_8_281_1308_0, i_8_281_1321_0,
    i_8_281_1331_0, i_8_281_1339_0, i_8_281_1348_0, i_8_281_1383_0,
    i_8_281_1399_0, i_8_281_1425_0, i_8_281_1426_0, i_8_281_1429_0,
    i_8_281_1471_0, i_8_281_1474_0, i_8_281_1509_0, i_8_281_1510_0,
    i_8_281_1527_0, i_8_281_1564_0, i_8_281_1565_0, i_8_281_1570_0,
    i_8_281_1588_0, i_8_281_1635_0, i_8_281_1636_0, i_8_281_1650_0,
    i_8_281_1651_0, i_8_281_1654_0, i_8_281_1689_0, i_8_281_1704_0,
    i_8_281_1752_0, i_8_281_1821_0, i_8_281_1822_0, i_8_281_1858_0,
    i_8_281_1860_0, i_8_281_1870_0, i_8_281_1876_0, i_8_281_1897_0,
    i_8_281_1906_0, i_8_281_1907_0, i_8_281_1978_0, i_8_281_1993_0,
    i_8_281_2041_0, i_8_281_2074_0, i_8_281_2091_0, i_8_281_2093_0,
    i_8_281_2215_0, i_8_281_2217_0, i_8_281_2227_0, i_8_281_2235_0;
  output o_8_281_0_0;
  assign o_8_281_0_0 = 0;
endmodule



// Benchmark "kernel_8_282" written by ABC on Sun Jul 19 10:07:58 2020

module kernel_8_282 ( 
    i_8_282_17_0, i_8_282_175_0, i_8_282_186_0, i_8_282_193_0,
    i_8_282_219_0, i_8_282_220_0, i_8_282_258_0, i_8_282_326_0,
    i_8_282_328_0, i_8_282_366_0, i_8_282_399_0, i_8_282_401_0,
    i_8_282_499_0, i_8_282_510_0, i_8_282_511_0, i_8_282_516_0,
    i_8_282_526_0, i_8_282_543_0, i_8_282_544_0, i_8_282_556_0,
    i_8_282_587_0, i_8_282_592_0, i_8_282_598_0, i_8_282_600_0,
    i_8_282_633_0, i_8_282_656_0, i_8_282_697_0, i_8_282_704_0,
    i_8_282_739_0, i_8_282_742_0, i_8_282_781_0, i_8_282_785_0,
    i_8_282_792_0, i_8_282_812_0, i_8_282_818_0, i_8_282_823_0,
    i_8_282_841_0, i_8_282_879_0, i_8_282_1014_0, i_8_282_1016_0,
    i_8_282_1051_0, i_8_282_1110_0, i_8_282_1123_0, i_8_282_1137_0,
    i_8_282_1155_0, i_8_282_1156_0, i_8_282_1158_0, i_8_282_1193_0,
    i_8_282_1236_0, i_8_282_1258_0, i_8_282_1274_0, i_8_282_1275_0,
    i_8_282_1279_0, i_8_282_1297_0, i_8_282_1302_0, i_8_282_1307_0,
    i_8_282_1314_0, i_8_282_1322_0, i_8_282_1330_0, i_8_282_1335_0,
    i_8_282_1338_0, i_8_282_1403_0, i_8_282_1462_0, i_8_282_1468_0,
    i_8_282_1472_0, i_8_282_1498_0, i_8_282_1560_0, i_8_282_1565_0,
    i_8_282_1608_0, i_8_282_1609_0, i_8_282_1636_0, i_8_282_1652_0,
    i_8_282_1653_0, i_8_282_1703_0, i_8_282_1706_0, i_8_282_1712_0,
    i_8_282_1749_0, i_8_282_1762_0, i_8_282_1774_0, i_8_282_1778_0,
    i_8_282_1833_0, i_8_282_1852_0, i_8_282_1886_0, i_8_282_1888_0,
    i_8_282_1950_0, i_8_282_1972_0, i_8_282_2055_0, i_8_282_2058_0,
    i_8_282_2113_0, i_8_282_2119_0, i_8_282_2157_0, i_8_282_2167_0,
    i_8_282_2170_0, i_8_282_2203_0, i_8_282_2211_0, i_8_282_2219_0,
    i_8_282_2230_0, i_8_282_2239_0, i_8_282_2244_0, i_8_282_2283_0,
    o_8_282_0_0  );
  input  i_8_282_17_0, i_8_282_175_0, i_8_282_186_0, i_8_282_193_0,
    i_8_282_219_0, i_8_282_220_0, i_8_282_258_0, i_8_282_326_0,
    i_8_282_328_0, i_8_282_366_0, i_8_282_399_0, i_8_282_401_0,
    i_8_282_499_0, i_8_282_510_0, i_8_282_511_0, i_8_282_516_0,
    i_8_282_526_0, i_8_282_543_0, i_8_282_544_0, i_8_282_556_0,
    i_8_282_587_0, i_8_282_592_0, i_8_282_598_0, i_8_282_600_0,
    i_8_282_633_0, i_8_282_656_0, i_8_282_697_0, i_8_282_704_0,
    i_8_282_739_0, i_8_282_742_0, i_8_282_781_0, i_8_282_785_0,
    i_8_282_792_0, i_8_282_812_0, i_8_282_818_0, i_8_282_823_0,
    i_8_282_841_0, i_8_282_879_0, i_8_282_1014_0, i_8_282_1016_0,
    i_8_282_1051_0, i_8_282_1110_0, i_8_282_1123_0, i_8_282_1137_0,
    i_8_282_1155_0, i_8_282_1156_0, i_8_282_1158_0, i_8_282_1193_0,
    i_8_282_1236_0, i_8_282_1258_0, i_8_282_1274_0, i_8_282_1275_0,
    i_8_282_1279_0, i_8_282_1297_0, i_8_282_1302_0, i_8_282_1307_0,
    i_8_282_1314_0, i_8_282_1322_0, i_8_282_1330_0, i_8_282_1335_0,
    i_8_282_1338_0, i_8_282_1403_0, i_8_282_1462_0, i_8_282_1468_0,
    i_8_282_1472_0, i_8_282_1498_0, i_8_282_1560_0, i_8_282_1565_0,
    i_8_282_1608_0, i_8_282_1609_0, i_8_282_1636_0, i_8_282_1652_0,
    i_8_282_1653_0, i_8_282_1703_0, i_8_282_1706_0, i_8_282_1712_0,
    i_8_282_1749_0, i_8_282_1762_0, i_8_282_1774_0, i_8_282_1778_0,
    i_8_282_1833_0, i_8_282_1852_0, i_8_282_1886_0, i_8_282_1888_0,
    i_8_282_1950_0, i_8_282_1972_0, i_8_282_2055_0, i_8_282_2058_0,
    i_8_282_2113_0, i_8_282_2119_0, i_8_282_2157_0, i_8_282_2167_0,
    i_8_282_2170_0, i_8_282_2203_0, i_8_282_2211_0, i_8_282_2219_0,
    i_8_282_2230_0, i_8_282_2239_0, i_8_282_2244_0, i_8_282_2283_0;
  output o_8_282_0_0;
  assign o_8_282_0_0 = 0;
endmodule



// Benchmark "kernel_8_283" written by ABC on Sun Jul 19 10:07:59 2020

module kernel_8_283 ( 
    i_8_283_20_0, i_8_283_27_0, i_8_283_56_0, i_8_283_58_0, i_8_283_59_0,
    i_8_283_112_0, i_8_283_113_0, i_8_283_137_0, i_8_283_142_0,
    i_8_283_143_0, i_8_283_184_0, i_8_283_221_0, i_8_283_226_0,
    i_8_283_254_0, i_8_283_257_0, i_8_283_299_0, i_8_283_301_0,
    i_8_283_304_0, i_8_283_320_0, i_8_283_329_0, i_8_283_425_0,
    i_8_283_451_0, i_8_283_452_0, i_8_283_454_0, i_8_283_478_0,
    i_8_283_479_0, i_8_283_524_0, i_8_283_554_0, i_8_283_586_0,
    i_8_283_605_0, i_8_283_632_0, i_8_283_634_0, i_8_283_640_0,
    i_8_283_649_0, i_8_283_662_0, i_8_283_680_0, i_8_283_706_0,
    i_8_283_713_0, i_8_283_779_0, i_8_283_830_0, i_8_283_838_0,
    i_8_283_848_0, i_8_283_883_0, i_8_283_929_0, i_8_283_965_0,
    i_8_283_968_0, i_8_283_1049_0, i_8_283_1064_0, i_8_283_1099_0,
    i_8_283_1135_0, i_8_283_1136_0, i_8_283_1138_0, i_8_283_1160_0,
    i_8_283_1220_0, i_8_283_1228_0, i_8_283_1264_0, i_8_283_1279_0,
    i_8_283_1315_0, i_8_283_1366_0, i_8_283_1404_0, i_8_283_1451_0,
    i_8_283_1467_0, i_8_283_1471_0, i_8_283_1475_0, i_8_283_1514_0,
    i_8_283_1544_0, i_8_283_1631_0, i_8_283_1633_0, i_8_283_1676_0,
    i_8_283_1678_0, i_8_283_1687_0, i_8_283_1703_0, i_8_283_1719_0,
    i_8_283_1759_0, i_8_283_1769_0, i_8_283_1774_0, i_8_283_1804_0,
    i_8_283_1820_0, i_8_283_1856_0, i_8_283_1858_0, i_8_283_1885_0,
    i_8_283_1964_0, i_8_283_1976_0, i_8_283_1981_0, i_8_283_1982_0,
    i_8_283_1990_0, i_8_283_1991_0, i_8_283_1993_0, i_8_283_1997_0,
    i_8_283_2047_0, i_8_283_2072_0, i_8_283_2074_0, i_8_283_2099_0,
    i_8_283_2142_0, i_8_283_2144_0, i_8_283_2147_0, i_8_283_2228_0,
    i_8_283_2245_0, i_8_283_2279_0, i_8_283_2290_0,
    o_8_283_0_0  );
  input  i_8_283_20_0, i_8_283_27_0, i_8_283_56_0, i_8_283_58_0,
    i_8_283_59_0, i_8_283_112_0, i_8_283_113_0, i_8_283_137_0,
    i_8_283_142_0, i_8_283_143_0, i_8_283_184_0, i_8_283_221_0,
    i_8_283_226_0, i_8_283_254_0, i_8_283_257_0, i_8_283_299_0,
    i_8_283_301_0, i_8_283_304_0, i_8_283_320_0, i_8_283_329_0,
    i_8_283_425_0, i_8_283_451_0, i_8_283_452_0, i_8_283_454_0,
    i_8_283_478_0, i_8_283_479_0, i_8_283_524_0, i_8_283_554_0,
    i_8_283_586_0, i_8_283_605_0, i_8_283_632_0, i_8_283_634_0,
    i_8_283_640_0, i_8_283_649_0, i_8_283_662_0, i_8_283_680_0,
    i_8_283_706_0, i_8_283_713_0, i_8_283_779_0, i_8_283_830_0,
    i_8_283_838_0, i_8_283_848_0, i_8_283_883_0, i_8_283_929_0,
    i_8_283_965_0, i_8_283_968_0, i_8_283_1049_0, i_8_283_1064_0,
    i_8_283_1099_0, i_8_283_1135_0, i_8_283_1136_0, i_8_283_1138_0,
    i_8_283_1160_0, i_8_283_1220_0, i_8_283_1228_0, i_8_283_1264_0,
    i_8_283_1279_0, i_8_283_1315_0, i_8_283_1366_0, i_8_283_1404_0,
    i_8_283_1451_0, i_8_283_1467_0, i_8_283_1471_0, i_8_283_1475_0,
    i_8_283_1514_0, i_8_283_1544_0, i_8_283_1631_0, i_8_283_1633_0,
    i_8_283_1676_0, i_8_283_1678_0, i_8_283_1687_0, i_8_283_1703_0,
    i_8_283_1719_0, i_8_283_1759_0, i_8_283_1769_0, i_8_283_1774_0,
    i_8_283_1804_0, i_8_283_1820_0, i_8_283_1856_0, i_8_283_1858_0,
    i_8_283_1885_0, i_8_283_1964_0, i_8_283_1976_0, i_8_283_1981_0,
    i_8_283_1982_0, i_8_283_1990_0, i_8_283_1991_0, i_8_283_1993_0,
    i_8_283_1997_0, i_8_283_2047_0, i_8_283_2072_0, i_8_283_2074_0,
    i_8_283_2099_0, i_8_283_2142_0, i_8_283_2144_0, i_8_283_2147_0,
    i_8_283_2228_0, i_8_283_2245_0, i_8_283_2279_0, i_8_283_2290_0;
  output o_8_283_0_0;
  assign o_8_283_0_0 = 0;
endmodule



// Benchmark "kernel_8_284" written by ABC on Sun Jul 19 10:08:00 2020

module kernel_8_284 ( 
    i_8_284_33_0, i_8_284_52_0, i_8_284_55_0, i_8_284_84_0, i_8_284_85_0,
    i_8_284_87_0, i_8_284_94_0, i_8_284_151_0, i_8_284_201_0,
    i_8_284_202_0, i_8_284_210_0, i_8_284_219_0, i_8_284_249_0,
    i_8_284_255_0, i_8_284_297_0, i_8_284_326_0, i_8_284_345_0,
    i_8_284_374_0, i_8_284_383_0, i_8_284_440_0, i_8_284_443_0,
    i_8_284_454_0, i_8_284_455_0, i_8_284_461_0, i_8_284_463_0,
    i_8_284_472_0, i_8_284_501_0, i_8_284_540_0, i_8_284_550_0,
    i_8_284_552_0, i_8_284_589_0, i_8_284_590_0, i_8_284_625_0,
    i_8_284_626_0, i_8_284_672_0, i_8_284_714_0, i_8_284_726_0,
    i_8_284_778_0, i_8_284_813_0, i_8_284_822_0, i_8_284_831_0,
    i_8_284_878_0, i_8_284_903_0, i_8_284_948_0, i_8_284_949_0,
    i_8_284_985_0, i_8_284_991_0, i_8_284_994_0, i_8_284_1029_0,
    i_8_284_1039_0, i_8_284_1053_0, i_8_284_1071_0, i_8_284_1083_0,
    i_8_284_1085_0, i_8_284_1112_0, i_8_284_1121_0, i_8_284_1138_0,
    i_8_284_1219_0, i_8_284_1240_0, i_8_284_1256_0, i_8_284_1259_0,
    i_8_284_1270_0, i_8_284_1274_0, i_8_284_1282_0, i_8_284_1283_0,
    i_8_284_1328_0, i_8_284_1395_0, i_8_284_1454_0, i_8_284_1472_0,
    i_8_284_1479_0, i_8_284_1480_0, i_8_284_1508_0, i_8_284_1509_0,
    i_8_284_1533_0, i_8_284_1541_0, i_8_284_1549_0, i_8_284_1555_0,
    i_8_284_1597_0, i_8_284_1607_0, i_8_284_1614_0, i_8_284_1615_0,
    i_8_284_1627_0, i_8_284_1738_0, i_8_284_1754_0, i_8_284_1759_0,
    i_8_284_1838_0, i_8_284_1841_0, i_8_284_1858_0, i_8_284_1864_0,
    i_8_284_1929_0, i_8_284_1975_0, i_8_284_2010_0, i_8_284_2047_0,
    i_8_284_2048_0, i_8_284_2049_0, i_8_284_2091_0, i_8_284_2109_0,
    i_8_284_2191_0, i_8_284_2223_0, i_8_284_2247_0,
    o_8_284_0_0  );
  input  i_8_284_33_0, i_8_284_52_0, i_8_284_55_0, i_8_284_84_0,
    i_8_284_85_0, i_8_284_87_0, i_8_284_94_0, i_8_284_151_0, i_8_284_201_0,
    i_8_284_202_0, i_8_284_210_0, i_8_284_219_0, i_8_284_249_0,
    i_8_284_255_0, i_8_284_297_0, i_8_284_326_0, i_8_284_345_0,
    i_8_284_374_0, i_8_284_383_0, i_8_284_440_0, i_8_284_443_0,
    i_8_284_454_0, i_8_284_455_0, i_8_284_461_0, i_8_284_463_0,
    i_8_284_472_0, i_8_284_501_0, i_8_284_540_0, i_8_284_550_0,
    i_8_284_552_0, i_8_284_589_0, i_8_284_590_0, i_8_284_625_0,
    i_8_284_626_0, i_8_284_672_0, i_8_284_714_0, i_8_284_726_0,
    i_8_284_778_0, i_8_284_813_0, i_8_284_822_0, i_8_284_831_0,
    i_8_284_878_0, i_8_284_903_0, i_8_284_948_0, i_8_284_949_0,
    i_8_284_985_0, i_8_284_991_0, i_8_284_994_0, i_8_284_1029_0,
    i_8_284_1039_0, i_8_284_1053_0, i_8_284_1071_0, i_8_284_1083_0,
    i_8_284_1085_0, i_8_284_1112_0, i_8_284_1121_0, i_8_284_1138_0,
    i_8_284_1219_0, i_8_284_1240_0, i_8_284_1256_0, i_8_284_1259_0,
    i_8_284_1270_0, i_8_284_1274_0, i_8_284_1282_0, i_8_284_1283_0,
    i_8_284_1328_0, i_8_284_1395_0, i_8_284_1454_0, i_8_284_1472_0,
    i_8_284_1479_0, i_8_284_1480_0, i_8_284_1508_0, i_8_284_1509_0,
    i_8_284_1533_0, i_8_284_1541_0, i_8_284_1549_0, i_8_284_1555_0,
    i_8_284_1597_0, i_8_284_1607_0, i_8_284_1614_0, i_8_284_1615_0,
    i_8_284_1627_0, i_8_284_1738_0, i_8_284_1754_0, i_8_284_1759_0,
    i_8_284_1838_0, i_8_284_1841_0, i_8_284_1858_0, i_8_284_1864_0,
    i_8_284_1929_0, i_8_284_1975_0, i_8_284_2010_0, i_8_284_2047_0,
    i_8_284_2048_0, i_8_284_2049_0, i_8_284_2091_0, i_8_284_2109_0,
    i_8_284_2191_0, i_8_284_2223_0, i_8_284_2247_0;
  output o_8_284_0_0;
  assign o_8_284_0_0 = 0;
endmodule



// Benchmark "kernel_8_285" written by ABC on Sun Jul 19 10:08:01 2020

module kernel_8_285 ( 
    i_8_285_17_0, i_8_285_48_0, i_8_285_49_0, i_8_285_51_0, i_8_285_85_0,
    i_8_285_93_0, i_8_285_96_0, i_8_285_114_0, i_8_285_139_0,
    i_8_285_142_0, i_8_285_143_0, i_8_285_177_0, i_8_285_183_0,
    i_8_285_186_0, i_8_285_193_0, i_8_285_196_0, i_8_285_231_0,
    i_8_285_257_0, i_8_285_344_0, i_8_285_345_0, i_8_285_348_0,
    i_8_285_354_0, i_8_285_357_0, i_8_285_361_0, i_8_285_433_0,
    i_8_285_444_0, i_8_285_456_0, i_8_285_494_0, i_8_285_573_0,
    i_8_285_582_0, i_8_285_601_0, i_8_285_654_0, i_8_285_660_0,
    i_8_285_703_0, i_8_285_748_0, i_8_285_768_0, i_8_285_774_0,
    i_8_285_825_0, i_8_285_843_0, i_8_285_924_0, i_8_285_933_0,
    i_8_285_958_0, i_8_285_966_0, i_8_285_967_0, i_8_285_969_0,
    i_8_285_1059_0, i_8_285_1071_0, i_8_285_1113_0, i_8_285_1119_0,
    i_8_285_1121_0, i_8_285_1126_0, i_8_285_1155_0, i_8_285_1166_0,
    i_8_285_1182_0, i_8_285_1183_0, i_8_285_1191_0, i_8_285_1232_0,
    i_8_285_1305_0, i_8_285_1307_0, i_8_285_1320_0, i_8_285_1329_0,
    i_8_285_1362_0, i_8_285_1366_0, i_8_285_1372_0, i_8_285_1407_0,
    i_8_285_1411_0, i_8_285_1470_0, i_8_285_1492_0, i_8_285_1560_0,
    i_8_285_1563_0, i_8_285_1564_0, i_8_285_1574_0, i_8_285_1641_0,
    i_8_285_1644_0, i_8_285_1648_0, i_8_285_1652_0, i_8_285_1655_0,
    i_8_285_1681_0, i_8_285_1689_0, i_8_285_1776_0, i_8_285_1833_0,
    i_8_285_1842_0, i_8_285_1877_0, i_8_285_1965_0, i_8_285_1996_0,
    i_8_285_2004_0, i_8_285_2073_0, i_8_285_2112_0, i_8_285_2143_0,
    i_8_285_2149_0, i_8_285_2157_0, i_8_285_2211_0, i_8_285_2214_0,
    i_8_285_2215_0, i_8_285_2216_0, i_8_285_2218_0, i_8_285_2229_0,
    i_8_285_2230_0, i_8_285_2232_0, i_8_285_2244_0,
    o_8_285_0_0  );
  input  i_8_285_17_0, i_8_285_48_0, i_8_285_49_0, i_8_285_51_0,
    i_8_285_85_0, i_8_285_93_0, i_8_285_96_0, i_8_285_114_0, i_8_285_139_0,
    i_8_285_142_0, i_8_285_143_0, i_8_285_177_0, i_8_285_183_0,
    i_8_285_186_0, i_8_285_193_0, i_8_285_196_0, i_8_285_231_0,
    i_8_285_257_0, i_8_285_344_0, i_8_285_345_0, i_8_285_348_0,
    i_8_285_354_0, i_8_285_357_0, i_8_285_361_0, i_8_285_433_0,
    i_8_285_444_0, i_8_285_456_0, i_8_285_494_0, i_8_285_573_0,
    i_8_285_582_0, i_8_285_601_0, i_8_285_654_0, i_8_285_660_0,
    i_8_285_703_0, i_8_285_748_0, i_8_285_768_0, i_8_285_774_0,
    i_8_285_825_0, i_8_285_843_0, i_8_285_924_0, i_8_285_933_0,
    i_8_285_958_0, i_8_285_966_0, i_8_285_967_0, i_8_285_969_0,
    i_8_285_1059_0, i_8_285_1071_0, i_8_285_1113_0, i_8_285_1119_0,
    i_8_285_1121_0, i_8_285_1126_0, i_8_285_1155_0, i_8_285_1166_0,
    i_8_285_1182_0, i_8_285_1183_0, i_8_285_1191_0, i_8_285_1232_0,
    i_8_285_1305_0, i_8_285_1307_0, i_8_285_1320_0, i_8_285_1329_0,
    i_8_285_1362_0, i_8_285_1366_0, i_8_285_1372_0, i_8_285_1407_0,
    i_8_285_1411_0, i_8_285_1470_0, i_8_285_1492_0, i_8_285_1560_0,
    i_8_285_1563_0, i_8_285_1564_0, i_8_285_1574_0, i_8_285_1641_0,
    i_8_285_1644_0, i_8_285_1648_0, i_8_285_1652_0, i_8_285_1655_0,
    i_8_285_1681_0, i_8_285_1689_0, i_8_285_1776_0, i_8_285_1833_0,
    i_8_285_1842_0, i_8_285_1877_0, i_8_285_1965_0, i_8_285_1996_0,
    i_8_285_2004_0, i_8_285_2073_0, i_8_285_2112_0, i_8_285_2143_0,
    i_8_285_2149_0, i_8_285_2157_0, i_8_285_2211_0, i_8_285_2214_0,
    i_8_285_2215_0, i_8_285_2216_0, i_8_285_2218_0, i_8_285_2229_0,
    i_8_285_2230_0, i_8_285_2232_0, i_8_285_2244_0;
  output o_8_285_0_0;
  assign o_8_285_0_0 = ~((~i_8_285_51_0 & ((~i_8_285_139_0 & ~i_8_285_361_0 & ~i_8_285_1155_0) | (~i_8_285_1119_0 & ~i_8_285_1305_0 & ~i_8_285_1470_0))) | (~i_8_285_231_0 & ((~i_8_285_17_0 & ~i_8_285_1307_0 & i_8_285_1648_0 & ~i_8_285_1842_0) | (~i_8_285_969_0 & i_8_285_1564_0 & ~i_8_285_2112_0 & ~i_8_285_2229_0))) | (~i_8_285_17_0 & ~i_8_285_774_0 & ((~i_8_285_93_0 & ~i_8_285_573_0 & ~i_8_285_1305_0 & ~i_8_285_1644_0 & ~i_8_285_2214_0) | (~i_8_285_494_0 & ~i_8_285_748_0 & ~i_8_285_1059_0 & ~i_8_285_1366_0 & ~i_8_285_2232_0))) | (~i_8_285_958_0 & ((~i_8_285_924_0 & ~i_8_285_1121_0 & i_8_285_2073_0) | (~i_8_285_582_0 & ~i_8_285_969_0 & ~i_8_285_1307_0 & ~i_8_285_1563_0 & ~i_8_285_2149_0))) | (~i_8_285_933_0 & ((~i_8_285_966_0 & ((~i_8_285_1126_0 & i_8_285_1329_0 & ~i_8_285_2004_0) | (~i_8_285_143_0 & ~i_8_285_257_0 & ~i_8_285_1833_0 & ~i_8_285_2218_0))) | (~i_8_285_49_0 & ~i_8_285_183_0 & ~i_8_285_967_0))) | (~i_8_285_924_0 & ((~i_8_285_143_0 & ((~i_8_285_433_0 & ~i_8_285_768_0 & ~i_8_285_1362_0 & ~i_8_285_1877_0 & ~i_8_285_2073_0) | (~i_8_285_139_0 & ~i_8_285_1320_0 & ~i_8_285_2112_0))) | (i_8_285_1182_0 & ~i_8_285_1470_0 & ~i_8_285_1877_0 & ~i_8_285_2211_0))) | (~i_8_285_354_0 & ~i_8_285_969_0 & i_8_285_1121_0 & ~i_8_285_1366_0 & ~i_8_285_1563_0 & i_8_285_1641_0) | (i_8_285_573_0 & i_8_285_2143_0) | (~i_8_285_177_0 & ~i_8_285_1372_0 & ~i_8_285_1641_0 & ~i_8_285_1877_0 & ~i_8_285_2211_0));
endmodule



// Benchmark "kernel_8_286" written by ABC on Sun Jul 19 10:08:02 2020

module kernel_8_286 ( 
    i_8_286_20_0, i_8_286_33_0, i_8_286_49_0, i_8_286_63_0, i_8_286_80_0,
    i_8_286_82_0, i_8_286_84_0, i_8_286_139_0, i_8_286_141_0,
    i_8_286_157_0, i_8_286_265_0, i_8_286_282_0, i_8_286_284_0,
    i_8_286_285_0, i_8_286_292_0, i_8_286_319_0, i_8_286_321_0,
    i_8_286_324_0, i_8_286_380_0, i_8_286_403_0, i_8_286_404_0,
    i_8_286_436_0, i_8_286_465_0, i_8_286_534_0, i_8_286_552_0,
    i_8_286_581_0, i_8_286_582_0, i_8_286_601_0, i_8_286_608_0,
    i_8_286_610_0, i_8_286_625_0, i_8_286_633_0, i_8_286_678_0,
    i_8_286_708_0, i_8_286_716_0, i_8_286_723_0, i_8_286_726_0,
    i_8_286_736_0, i_8_286_737_0, i_8_286_795_0, i_8_286_813_0,
    i_8_286_870_0, i_8_286_922_0, i_8_286_931_0, i_8_286_951_0,
    i_8_286_980_0, i_8_286_985_0, i_8_286_991_0, i_8_286_1012_0,
    i_8_286_1030_0, i_8_286_1032_0, i_8_286_1110_0, i_8_286_1112_0,
    i_8_286_1182_0, i_8_286_1185_0, i_8_286_1236_0, i_8_286_1239_0,
    i_8_286_1240_0, i_8_286_1260_0, i_8_286_1261_0, i_8_286_1285_0,
    i_8_286_1331_0, i_8_286_1383_0, i_8_286_1401_0, i_8_286_1436_0,
    i_8_286_1443_0, i_8_286_1570_0, i_8_286_1614_0, i_8_286_1623_0,
    i_8_286_1635_0, i_8_286_1649_0, i_8_286_1675_0, i_8_286_1680_0,
    i_8_286_1722_0, i_8_286_1734_0, i_8_286_1736_0, i_8_286_1749_0,
    i_8_286_1822_0, i_8_286_1848_0, i_8_286_1858_0, i_8_286_1863_0,
    i_8_286_1902_0, i_8_286_1903_0, i_8_286_1911_0, i_8_286_1915_0,
    i_8_286_1948_0, i_8_286_1957_0, i_8_286_1960_0, i_8_286_2014_0,
    i_8_286_2015_0, i_8_286_2029_0, i_8_286_2031_0, i_8_286_2058_0,
    i_8_286_2136_0, i_8_286_2152_0, i_8_286_2153_0, i_8_286_2163_0,
    i_8_286_2241_0, i_8_286_2262_0, i_8_286_2266_0,
    o_8_286_0_0  );
  input  i_8_286_20_0, i_8_286_33_0, i_8_286_49_0, i_8_286_63_0,
    i_8_286_80_0, i_8_286_82_0, i_8_286_84_0, i_8_286_139_0, i_8_286_141_0,
    i_8_286_157_0, i_8_286_265_0, i_8_286_282_0, i_8_286_284_0,
    i_8_286_285_0, i_8_286_292_0, i_8_286_319_0, i_8_286_321_0,
    i_8_286_324_0, i_8_286_380_0, i_8_286_403_0, i_8_286_404_0,
    i_8_286_436_0, i_8_286_465_0, i_8_286_534_0, i_8_286_552_0,
    i_8_286_581_0, i_8_286_582_0, i_8_286_601_0, i_8_286_608_0,
    i_8_286_610_0, i_8_286_625_0, i_8_286_633_0, i_8_286_678_0,
    i_8_286_708_0, i_8_286_716_0, i_8_286_723_0, i_8_286_726_0,
    i_8_286_736_0, i_8_286_737_0, i_8_286_795_0, i_8_286_813_0,
    i_8_286_870_0, i_8_286_922_0, i_8_286_931_0, i_8_286_951_0,
    i_8_286_980_0, i_8_286_985_0, i_8_286_991_0, i_8_286_1012_0,
    i_8_286_1030_0, i_8_286_1032_0, i_8_286_1110_0, i_8_286_1112_0,
    i_8_286_1182_0, i_8_286_1185_0, i_8_286_1236_0, i_8_286_1239_0,
    i_8_286_1240_0, i_8_286_1260_0, i_8_286_1261_0, i_8_286_1285_0,
    i_8_286_1331_0, i_8_286_1383_0, i_8_286_1401_0, i_8_286_1436_0,
    i_8_286_1443_0, i_8_286_1570_0, i_8_286_1614_0, i_8_286_1623_0,
    i_8_286_1635_0, i_8_286_1649_0, i_8_286_1675_0, i_8_286_1680_0,
    i_8_286_1722_0, i_8_286_1734_0, i_8_286_1736_0, i_8_286_1749_0,
    i_8_286_1822_0, i_8_286_1848_0, i_8_286_1858_0, i_8_286_1863_0,
    i_8_286_1902_0, i_8_286_1903_0, i_8_286_1911_0, i_8_286_1915_0,
    i_8_286_1948_0, i_8_286_1957_0, i_8_286_1960_0, i_8_286_2014_0,
    i_8_286_2015_0, i_8_286_2029_0, i_8_286_2031_0, i_8_286_2058_0,
    i_8_286_2136_0, i_8_286_2152_0, i_8_286_2153_0, i_8_286_2163_0,
    i_8_286_2241_0, i_8_286_2262_0, i_8_286_2266_0;
  output o_8_286_0_0;
  assign o_8_286_0_0 = 0;
endmodule



// Benchmark "kernel_8_287" written by ABC on Sun Jul 19 10:08:03 2020

module kernel_8_287 ( 
    i_8_287_41_0, i_8_287_77_0, i_8_287_80_0, i_8_287_194_0, i_8_287_202_0,
    i_8_287_203_0, i_8_287_247_0, i_8_287_278_0, i_8_287_301_0,
    i_8_287_356_0, i_8_287_358_0, i_8_287_364_0, i_8_287_367_0,
    i_8_287_391_0, i_8_287_392_0, i_8_287_424_0, i_8_287_460_0,
    i_8_287_499_0, i_8_287_527_0, i_8_287_529_0, i_8_287_536_0,
    i_8_287_593_0, i_8_287_607_0, i_8_287_608_0, i_8_287_610_0,
    i_8_287_612_0, i_8_287_614_0, i_8_287_635_0, i_8_287_638_0,
    i_8_287_642_0, i_8_287_648_0, i_8_287_656_0, i_8_287_664_0,
    i_8_287_679_0, i_8_287_703_0, i_8_287_704_0, i_8_287_706_0,
    i_8_287_710_0, i_8_287_812_0, i_8_287_832_0, i_8_287_833_0,
    i_8_287_835_0, i_8_287_840_0, i_8_287_842_0, i_8_287_857_0,
    i_8_287_869_0, i_8_287_873_0, i_8_287_875_0, i_8_287_956_0,
    i_8_287_967_0, i_8_287_970_0, i_8_287_1053_0, i_8_287_1133_0,
    i_8_287_1154_0, i_8_287_1174_0, i_8_287_1192_0, i_8_287_1228_0,
    i_8_287_1267_0, i_8_287_1285_0, i_8_287_1286_0, i_8_287_1315_0,
    i_8_287_1352_0, i_8_287_1382_0, i_8_287_1400_0, i_8_287_1404_0,
    i_8_287_1436_0, i_8_287_1438_0, i_8_287_1496_0, i_8_287_1508_0,
    i_8_287_1532_0, i_8_287_1551_0, i_8_287_1574_0, i_8_287_1607_0,
    i_8_287_1660_0, i_8_287_1670_0, i_8_287_1702_0, i_8_287_1703_0,
    i_8_287_1750_0, i_8_287_1751_0, i_8_287_1775_0, i_8_287_1803_0,
    i_8_287_1823_0, i_8_287_1825_0, i_8_287_1913_0, i_8_287_1951_0,
    i_8_287_1967_0, i_8_287_1996_0, i_8_287_2012_0, i_8_287_2052_0,
    i_8_287_2065_0, i_8_287_2107_0, i_8_287_2120_0, i_8_287_2129_0,
    i_8_287_2144_0, i_8_287_2145_0, i_8_287_2224_0, i_8_287_2247_0,
    i_8_287_2297_0, i_8_287_2299_0, i_8_287_2300_0,
    o_8_287_0_0  );
  input  i_8_287_41_0, i_8_287_77_0, i_8_287_80_0, i_8_287_194_0,
    i_8_287_202_0, i_8_287_203_0, i_8_287_247_0, i_8_287_278_0,
    i_8_287_301_0, i_8_287_356_0, i_8_287_358_0, i_8_287_364_0,
    i_8_287_367_0, i_8_287_391_0, i_8_287_392_0, i_8_287_424_0,
    i_8_287_460_0, i_8_287_499_0, i_8_287_527_0, i_8_287_529_0,
    i_8_287_536_0, i_8_287_593_0, i_8_287_607_0, i_8_287_608_0,
    i_8_287_610_0, i_8_287_612_0, i_8_287_614_0, i_8_287_635_0,
    i_8_287_638_0, i_8_287_642_0, i_8_287_648_0, i_8_287_656_0,
    i_8_287_664_0, i_8_287_679_0, i_8_287_703_0, i_8_287_704_0,
    i_8_287_706_0, i_8_287_710_0, i_8_287_812_0, i_8_287_832_0,
    i_8_287_833_0, i_8_287_835_0, i_8_287_840_0, i_8_287_842_0,
    i_8_287_857_0, i_8_287_869_0, i_8_287_873_0, i_8_287_875_0,
    i_8_287_956_0, i_8_287_967_0, i_8_287_970_0, i_8_287_1053_0,
    i_8_287_1133_0, i_8_287_1154_0, i_8_287_1174_0, i_8_287_1192_0,
    i_8_287_1228_0, i_8_287_1267_0, i_8_287_1285_0, i_8_287_1286_0,
    i_8_287_1315_0, i_8_287_1352_0, i_8_287_1382_0, i_8_287_1400_0,
    i_8_287_1404_0, i_8_287_1436_0, i_8_287_1438_0, i_8_287_1496_0,
    i_8_287_1508_0, i_8_287_1532_0, i_8_287_1551_0, i_8_287_1574_0,
    i_8_287_1607_0, i_8_287_1660_0, i_8_287_1670_0, i_8_287_1702_0,
    i_8_287_1703_0, i_8_287_1750_0, i_8_287_1751_0, i_8_287_1775_0,
    i_8_287_1803_0, i_8_287_1823_0, i_8_287_1825_0, i_8_287_1913_0,
    i_8_287_1951_0, i_8_287_1967_0, i_8_287_1996_0, i_8_287_2012_0,
    i_8_287_2052_0, i_8_287_2065_0, i_8_287_2107_0, i_8_287_2120_0,
    i_8_287_2129_0, i_8_287_2144_0, i_8_287_2145_0, i_8_287_2224_0,
    i_8_287_2247_0, i_8_287_2297_0, i_8_287_2299_0, i_8_287_2300_0;
  output o_8_287_0_0;
  assign o_8_287_0_0 = 0;
endmodule



// Benchmark "kernel_8_288" written by ABC on Sun Jul 19 10:08:05 2020

module kernel_8_288 ( 
    i_8_288_19_0, i_8_288_30_0, i_8_288_31_0, i_8_288_32_0, i_8_288_53_0,
    i_8_288_85_0, i_8_288_103_0, i_8_288_109_0, i_8_288_111_0,
    i_8_288_153_0, i_8_288_163_0, i_8_288_228_0, i_8_288_236_0,
    i_8_288_238_0, i_8_288_326_0, i_8_288_373_0, i_8_288_378_0,
    i_8_288_439_0, i_8_288_471_0, i_8_288_480_0, i_8_288_549_0,
    i_8_288_568_0, i_8_288_569_0, i_8_288_610_0, i_8_288_613_0,
    i_8_288_615_0, i_8_288_684_0, i_8_288_692_0, i_8_288_698_0,
    i_8_288_703_0, i_8_288_705_0, i_8_288_759_0, i_8_288_847_0,
    i_8_288_858_0, i_8_288_882_0, i_8_288_937_0, i_8_288_939_0,
    i_8_288_956_0, i_8_288_985_0, i_8_288_1008_0, i_8_288_1038_0,
    i_8_288_1039_0, i_8_288_1041_0, i_8_288_1042_0, i_8_288_1069_0,
    i_8_288_1118_0, i_8_288_1120_0, i_8_288_1183_0, i_8_288_1188_0,
    i_8_288_1260_0, i_8_288_1288_0, i_8_288_1291_0, i_8_288_1296_0,
    i_8_288_1306_0, i_8_288_1411_0, i_8_288_1432_0, i_8_288_1433_0,
    i_8_288_1435_0, i_8_288_1449_0, i_8_288_1454_0, i_8_288_1472_0,
    i_8_288_1532_0, i_8_288_1574_0, i_8_288_1622_0, i_8_288_1676_0,
    i_8_288_1696_0, i_8_288_1719_0, i_8_288_1720_0, i_8_288_1740_0,
    i_8_288_1746_0, i_8_288_1770_0, i_8_288_1808_0, i_8_288_1821_0,
    i_8_288_1828_0, i_8_288_1830_0, i_8_288_1854_0, i_8_288_1855_0,
    i_8_288_1881_0, i_8_288_1882_0, i_8_288_1884_0, i_8_288_1892_0,
    i_8_288_1901_0, i_8_288_1903_0, i_8_288_1962_0, i_8_288_1982_0,
    i_8_288_2044_0, i_8_288_2047_0, i_8_288_2074_0, i_8_288_2144_0,
    i_8_288_2147_0, i_8_288_2149_0, i_8_288_2170_0, i_8_288_2172_0,
    i_8_288_2190_0, i_8_288_2215_0, i_8_288_2229_0, i_8_288_2242_0,
    i_8_288_2272_0, i_8_288_2296_0, i_8_288_2297_0,
    o_8_288_0_0  );
  input  i_8_288_19_0, i_8_288_30_0, i_8_288_31_0, i_8_288_32_0,
    i_8_288_53_0, i_8_288_85_0, i_8_288_103_0, i_8_288_109_0,
    i_8_288_111_0, i_8_288_153_0, i_8_288_163_0, i_8_288_228_0,
    i_8_288_236_0, i_8_288_238_0, i_8_288_326_0, i_8_288_373_0,
    i_8_288_378_0, i_8_288_439_0, i_8_288_471_0, i_8_288_480_0,
    i_8_288_549_0, i_8_288_568_0, i_8_288_569_0, i_8_288_610_0,
    i_8_288_613_0, i_8_288_615_0, i_8_288_684_0, i_8_288_692_0,
    i_8_288_698_0, i_8_288_703_0, i_8_288_705_0, i_8_288_759_0,
    i_8_288_847_0, i_8_288_858_0, i_8_288_882_0, i_8_288_937_0,
    i_8_288_939_0, i_8_288_956_0, i_8_288_985_0, i_8_288_1008_0,
    i_8_288_1038_0, i_8_288_1039_0, i_8_288_1041_0, i_8_288_1042_0,
    i_8_288_1069_0, i_8_288_1118_0, i_8_288_1120_0, i_8_288_1183_0,
    i_8_288_1188_0, i_8_288_1260_0, i_8_288_1288_0, i_8_288_1291_0,
    i_8_288_1296_0, i_8_288_1306_0, i_8_288_1411_0, i_8_288_1432_0,
    i_8_288_1433_0, i_8_288_1435_0, i_8_288_1449_0, i_8_288_1454_0,
    i_8_288_1472_0, i_8_288_1532_0, i_8_288_1574_0, i_8_288_1622_0,
    i_8_288_1676_0, i_8_288_1696_0, i_8_288_1719_0, i_8_288_1720_0,
    i_8_288_1740_0, i_8_288_1746_0, i_8_288_1770_0, i_8_288_1808_0,
    i_8_288_1821_0, i_8_288_1828_0, i_8_288_1830_0, i_8_288_1854_0,
    i_8_288_1855_0, i_8_288_1881_0, i_8_288_1882_0, i_8_288_1884_0,
    i_8_288_1892_0, i_8_288_1901_0, i_8_288_1903_0, i_8_288_1962_0,
    i_8_288_1982_0, i_8_288_2044_0, i_8_288_2047_0, i_8_288_2074_0,
    i_8_288_2144_0, i_8_288_2147_0, i_8_288_2149_0, i_8_288_2170_0,
    i_8_288_2172_0, i_8_288_2190_0, i_8_288_2215_0, i_8_288_2229_0,
    i_8_288_2242_0, i_8_288_2272_0, i_8_288_2296_0, i_8_288_2297_0;
  output o_8_288_0_0;
  assign o_8_288_0_0 = ~((~i_8_288_2044_0 & ((~i_8_288_1676_0 & ((~i_8_288_30_0 & ~i_8_288_1855_0 & ((~i_8_288_103_0 & ~i_8_288_163_0 & ~i_8_288_569_0 & ~i_8_288_698_0 & ~i_8_288_847_0 & ~i_8_288_882_0 & ~i_8_288_937_0 & ~i_8_288_939_0 & ~i_8_288_985_0 & ~i_8_288_1288_0 & ~i_8_288_1982_0 & ~i_8_288_2170_0 & ~i_8_288_2172_0) | (~i_8_288_236_0 & ~i_8_288_326_0 & ~i_8_288_480_0 & ~i_8_288_1449_0 & ~i_8_288_1454_0 & ~i_8_288_1719_0 & ~i_8_288_1720_0 & ~i_8_288_1854_0 & ~i_8_288_2242_0))) | (~i_8_288_53_0 & ~i_8_288_109_0 & ~i_8_288_439_0 & ~i_8_288_568_0 & ~i_8_288_985_0 & ~i_8_288_1433_0 & ~i_8_288_1532_0 & i_8_288_1719_0) | (i_8_288_378_0 & ~i_8_288_569_0 & i_8_288_759_0 & ~i_8_288_939_0 & ~i_8_288_1296_0 & ~i_8_288_2297_0))) | (~i_8_288_480_0 & ((~i_8_288_32_0 & ((~i_8_288_847_0 & ~i_8_288_937_0 & i_8_288_956_0 & i_8_288_1454_0) | (~i_8_288_53_0 & i_8_288_103_0 & ~i_8_288_109_0 & ~i_8_288_238_0 & ~i_8_288_569_0 & ~i_8_288_939_0 & ~i_8_288_985_0 & ~i_8_288_1291_0 & ~i_8_288_2144_0))) | (~i_8_288_326_0 & ~i_8_288_610_0 & ~i_8_288_613_0 & ~i_8_288_847_0 & ~i_8_288_882_0 & ~i_8_288_1008_0 & ~i_8_288_1038_0 & ~i_8_288_1433_0 & ~i_8_288_2147_0))) | (~i_8_288_373_0 & ((~i_8_288_109_0 & i_8_288_613_0 & i_8_288_1676_0 & ~i_8_288_1720_0 & i_8_288_2144_0) | (~i_8_288_568_0 & ~i_8_288_703_0 & ~i_8_288_847_0 & ~i_8_288_937_0 & ~i_8_288_1118_0 & i_8_288_1183_0 & ~i_8_288_1188_0 & ~i_8_288_1719_0 & ~i_8_288_1808_0 & ~i_8_288_2229_0))) | (~i_8_288_1291_0 & ~i_8_288_1622_0 & ((~i_8_288_236_0 & ~i_8_288_549_0 & ~i_8_288_568_0 & ~i_8_288_610_0 & i_8_288_703_0 & ~i_8_288_858_0 & ~i_8_288_1039_0 & ~i_8_288_1454_0) | (i_8_288_378_0 & i_8_288_847_0 & ~i_8_288_939_0 & ~i_8_288_956_0 & ~i_8_288_1720_0 & ~i_8_288_1854_0 & ~i_8_288_1881_0 & ~i_8_288_2047_0))))) | (~i_8_288_1720_0 & ((~i_8_288_30_0 & ((~i_8_288_53_0 & ~i_8_288_1433_0 & ~i_8_288_1828_0 & ((~i_8_288_228_0 & ~i_8_288_373_0 & ~i_8_288_549_0 & ~i_8_288_1038_0 & ~i_8_288_1449_0 & ~i_8_288_1622_0 & ~i_8_288_1901_0 & ~i_8_288_1982_0 & ~i_8_288_2047_0) | (~i_8_288_85_0 & ~i_8_288_236_0 & ~i_8_288_439_0 & ~i_8_288_480_0 & ~i_8_288_684_0 & ~i_8_288_939_0 & ~i_8_288_1288_0 & ~i_8_288_1532_0 & ~i_8_288_1676_0 & ~i_8_288_1808_0 & ~i_8_288_2242_0))) | (~i_8_288_1719_0 & ((~i_8_288_109_0 & ~i_8_288_236_0 & ~i_8_288_326_0 & ~i_8_288_985_0 & ~i_8_288_1622_0 & ~i_8_288_1746_0 & ~i_8_288_2190_0) | (~i_8_288_19_0 & ~i_8_288_163_0 & ~i_8_288_698_0 & ~i_8_288_1260_0 & ~i_8_288_1454_0 & i_8_288_1696_0 & ~i_8_288_2170_0 & ~i_8_288_2242_0))))) | (~i_8_288_1719_0 & ((~i_8_288_103_0 & ~i_8_288_1982_0 & ((~i_8_288_163_0 & ~i_8_288_326_0 & ~i_8_288_613_0 & ~i_8_288_985_0 & ~i_8_288_1676_0 & ~i_8_288_1740_0 & ~i_8_288_1746_0 & ~i_8_288_1808_0) | (~i_8_288_549_0 & ~i_8_288_1039_0 & i_8_288_1962_0 & ~i_8_288_2147_0 & ~i_8_288_2172_0))) | (~i_8_288_236_0 & ~i_8_288_326_0 & ~i_8_288_471_0 & ~i_8_288_858_0 & ~i_8_288_939_0 & ~i_8_288_1260_0 & ~i_8_288_1622_0 & ~i_8_288_1854_0 & ~i_8_288_1882_0 & ~i_8_288_2144_0 & ~i_8_288_2170_0))) | (i_8_288_703_0 & ((~i_8_288_228_0 & i_8_288_705_0 & i_8_288_1882_0) | (~i_8_288_568_0 & ~i_8_288_1038_0 & ~i_8_288_1260_0 & ~i_8_288_1433_0 & ~i_8_288_1435_0 & ~i_8_288_2297_0))) | (~i_8_288_2144_0 & ((~i_8_288_549_0 & i_8_288_705_0 & ~i_8_288_1433_0 & ~i_8_288_1449_0 & ~i_8_288_1622_0) | (~i_8_288_480_0 & i_8_288_1306_0 & i_8_288_1432_0 & ~i_8_288_2297_0))) | (~i_8_288_326_0 & i_8_288_613_0 & ~i_8_288_759_0 & ~i_8_288_1260_0 & ~i_8_288_1432_0 & ~i_8_288_1903_0 & ~i_8_288_1982_0))) | (~i_8_288_85_0 & ((i_8_288_985_0 & ~i_8_288_1042_0 & ~i_8_288_1435_0 & i_8_288_1454_0 & ~i_8_288_1472_0 & ~i_8_288_2144_0 & ~i_8_288_2172_0) | (~i_8_288_471_0 & ~i_8_288_569_0 & ~i_8_288_692_0 & ~i_8_288_985_0 & i_8_288_1291_0 & ~i_8_288_2229_0 & ~i_8_288_2296_0))) | (~i_8_288_1008_0 & ((i_8_288_109_0 & ~i_8_288_1676_0 & ~i_8_288_1746_0 & ((~i_8_288_30_0 & ~i_8_288_163_0 & ~i_8_288_568_0 & ~i_8_288_985_0 & ~i_8_288_1042_0 & ~i_8_288_1288_0 & ~i_8_288_1855_0 & ~i_8_288_1901_0 & ~i_8_288_1982_0) | (~i_8_288_103_0 & ~i_8_288_1038_0 & ~i_8_288_1039_0 & ~i_8_288_1260_0 & ~i_8_288_1454_0 & ~i_8_288_1622_0 & ~i_8_288_1719_0 & ~i_8_288_1962_0 & ~i_8_288_2170_0))) | (~i_8_288_569_0 & i_8_288_705_0 & ~i_8_288_1449_0 & ~i_8_288_1454_0 & i_8_288_1821_0 & ~i_8_288_1854_0) | (~i_8_288_163_0 & ~i_8_288_326_0 & ~i_8_288_373_0 & ~i_8_288_684_0 & ~i_8_288_858_0 & ~i_8_288_937_0 & ~i_8_288_1039_0 & ~i_8_288_1901_0 & ~i_8_288_2047_0 & i_8_288_2144_0 & ~i_8_288_2297_0))) | (~i_8_288_326_0 & ((~i_8_288_30_0 & ~i_8_288_1532_0 & ((~i_8_288_1120_0 & ~i_8_288_1188_0 & ~i_8_288_1260_0 & i_8_288_1472_0 & ~i_8_288_1901_0) | (~i_8_288_103_0 & i_8_288_111_0 & ~i_8_288_163_0 & ~i_8_288_1296_0 & ~i_8_288_1746_0 & ~i_8_288_2190_0))) | (~i_8_288_1982_0 & ((~i_8_288_31_0 & ~i_8_288_1901_0 & ((~i_8_288_236_0 & ~i_8_288_568_0 & i_8_288_705_0 & ~i_8_288_1472_0 & ~i_8_288_1854_0) | (~i_8_288_103_0 & ~i_8_288_569_0 & i_8_288_703_0 & ~i_8_288_939_0 & i_8_288_2272_0))) | (~i_8_288_103_0 & ~i_8_288_568_0 & ~i_8_288_569_0 & ~i_8_288_937_0 & ~i_8_288_939_0 & ~i_8_288_985_0 & ~i_8_288_1039_0 & ~i_8_288_1296_0 & ~i_8_288_1433_0 & ~i_8_288_1719_0))) | (~i_8_288_939_0 & ~i_8_288_956_0 & ~i_8_288_153_0 & i_8_288_615_0 & ~i_8_288_1288_0 & ~i_8_288_1306_0 & i_8_288_1432_0 & ~i_8_288_2296_0 & ~i_8_288_2297_0))) | (~i_8_288_163_0 & ((~i_8_288_103_0 & ~i_8_288_698_0 & ~i_8_288_1830_0 & ((~i_8_288_238_0 & i_8_288_373_0 & ~i_8_288_549_0 & ~i_8_288_568_0 & ~i_8_288_939_0 & ~i_8_288_956_0 & ~i_8_288_1296_0 & ~i_8_288_1901_0) | (~i_8_288_236_0 & ~i_8_288_439_0 & ~i_8_288_569_0 & ~i_8_288_1038_0 & ~i_8_288_1118_0 & ~i_8_288_1183_0 & ~i_8_288_1454_0 & ~i_8_288_1828_0 & ~i_8_288_1854_0 & ~i_8_288_1881_0 & ~i_8_288_1982_0 & ~i_8_288_2144_0 & ~i_8_288_2296_0))) | (~i_8_288_236_0 & ((~i_8_288_31_0 & i_8_288_373_0 & i_8_288_1884_0) | (~i_8_288_684_0 & ~i_8_288_1188_0 & ~i_8_288_1432_0 & i_8_288_1454_0 & ~i_8_288_1532_0 & ~i_8_288_1828_0 & ~i_8_288_1901_0 & ~i_8_288_2047_0))) | (~i_8_288_985_0 & ((~i_8_288_684_0 & ~i_8_288_1432_0 & ~i_8_288_1622_0 & ~i_8_288_1982_0 & i_8_288_2147_0) | (~i_8_288_549_0 & ~i_8_288_569_0 & ~i_8_288_937_0 & ~i_8_288_1039_0 & ~i_8_288_1288_0 & ~i_8_288_1291_0 & ~i_8_288_1676_0 & i_8_288_2242_0))))) | (~i_8_288_985_0 & ~i_8_288_1306_0 & ((~i_8_288_684_0 & ~i_8_288_692_0 & ~i_8_288_698_0 & ~i_8_288_703_0 & i_8_288_1892_0 & ~i_8_288_2047_0) | (~i_8_288_569_0 & ~i_8_288_1432_0 & i_8_288_1454_0 & ~i_8_288_1903_0 & i_8_288_2147_0 & ~i_8_288_2297_0))) | (i_8_288_1962_0 & i_8_288_1982_0 & i_8_288_2147_0 & ~i_8_288_2242_0 & i_8_288_2272_0));
endmodule



// Benchmark "kernel_8_289" written by ABC on Sun Jul 19 10:08:05 2020

module kernel_8_289 ( 
    i_8_289_24_0, i_8_289_26_0, i_8_289_33_0, i_8_289_57_0, i_8_289_61_0,
    i_8_289_88_0, i_8_289_105_0, i_8_289_142_0, i_8_289_168_0,
    i_8_289_177_0, i_8_289_196_0, i_8_289_228_0, i_8_289_258_0,
    i_8_289_303_0, i_8_289_333_0, i_8_289_336_0, i_8_289_369_0,
    i_8_289_393_0, i_8_289_394_0, i_8_289_420_0, i_8_289_426_0,
    i_8_289_465_0, i_8_289_492_0, i_8_289_539_0, i_8_289_591_0,
    i_8_289_595_0, i_8_289_597_0, i_8_289_600_0, i_8_289_610_0,
    i_8_289_642_0, i_8_289_661_0, i_8_289_690_0, i_8_289_703_0,
    i_8_289_708_0, i_8_289_733_0, i_8_289_754_0, i_8_289_780_0,
    i_8_289_840_0, i_8_289_852_0, i_8_289_867_0, i_8_289_876_0,
    i_8_289_888_0, i_8_289_924_0, i_8_289_958_0, i_8_289_982_0,
    i_8_289_993_0, i_8_289_1041_0, i_8_289_1105_0, i_8_289_1132_0,
    i_8_289_1176_0, i_8_289_1203_0, i_8_289_1227_0, i_8_289_1230_0,
    i_8_289_1231_0, i_8_289_1262_0, i_8_289_1263_0, i_8_289_1264_0,
    i_8_289_1281_0, i_8_289_1284_0, i_8_289_1311_0, i_8_289_1326_0,
    i_8_289_1362_0, i_8_289_1366_0, i_8_289_1389_0, i_8_289_1398_0,
    i_8_289_1407_0, i_8_289_1437_0, i_8_289_1440_0, i_8_289_1473_0,
    i_8_289_1501_0, i_8_289_1626_0, i_8_289_1674_0, i_8_289_1707_0,
    i_8_289_1749_0, i_8_289_1753_0, i_8_289_1770_0, i_8_289_1779_0,
    i_8_289_1786_0, i_8_289_1789_0, i_8_289_1812_0, i_8_289_1869_0,
    i_8_289_1875_0, i_8_289_1914_0, i_8_289_1965_0, i_8_289_1981_0,
    i_8_289_1983_0, i_8_289_1995_0, i_8_289_2067_0, i_8_289_2103_0,
    i_8_289_2136_0, i_8_289_2145_0, i_8_289_2148_0, i_8_289_2149_0,
    i_8_289_2151_0, i_8_289_2152_0, i_8_289_2154_0, i_8_289_2230_0,
    i_8_289_2235_0, i_8_289_2262_0, i_8_289_2293_0,
    o_8_289_0_0  );
  input  i_8_289_24_0, i_8_289_26_0, i_8_289_33_0, i_8_289_57_0,
    i_8_289_61_0, i_8_289_88_0, i_8_289_105_0, i_8_289_142_0,
    i_8_289_168_0, i_8_289_177_0, i_8_289_196_0, i_8_289_228_0,
    i_8_289_258_0, i_8_289_303_0, i_8_289_333_0, i_8_289_336_0,
    i_8_289_369_0, i_8_289_393_0, i_8_289_394_0, i_8_289_420_0,
    i_8_289_426_0, i_8_289_465_0, i_8_289_492_0, i_8_289_539_0,
    i_8_289_591_0, i_8_289_595_0, i_8_289_597_0, i_8_289_600_0,
    i_8_289_610_0, i_8_289_642_0, i_8_289_661_0, i_8_289_690_0,
    i_8_289_703_0, i_8_289_708_0, i_8_289_733_0, i_8_289_754_0,
    i_8_289_780_0, i_8_289_840_0, i_8_289_852_0, i_8_289_867_0,
    i_8_289_876_0, i_8_289_888_0, i_8_289_924_0, i_8_289_958_0,
    i_8_289_982_0, i_8_289_993_0, i_8_289_1041_0, i_8_289_1105_0,
    i_8_289_1132_0, i_8_289_1176_0, i_8_289_1203_0, i_8_289_1227_0,
    i_8_289_1230_0, i_8_289_1231_0, i_8_289_1262_0, i_8_289_1263_0,
    i_8_289_1264_0, i_8_289_1281_0, i_8_289_1284_0, i_8_289_1311_0,
    i_8_289_1326_0, i_8_289_1362_0, i_8_289_1366_0, i_8_289_1389_0,
    i_8_289_1398_0, i_8_289_1407_0, i_8_289_1437_0, i_8_289_1440_0,
    i_8_289_1473_0, i_8_289_1501_0, i_8_289_1626_0, i_8_289_1674_0,
    i_8_289_1707_0, i_8_289_1749_0, i_8_289_1753_0, i_8_289_1770_0,
    i_8_289_1779_0, i_8_289_1786_0, i_8_289_1789_0, i_8_289_1812_0,
    i_8_289_1869_0, i_8_289_1875_0, i_8_289_1914_0, i_8_289_1965_0,
    i_8_289_1981_0, i_8_289_1983_0, i_8_289_1995_0, i_8_289_2067_0,
    i_8_289_2103_0, i_8_289_2136_0, i_8_289_2145_0, i_8_289_2148_0,
    i_8_289_2149_0, i_8_289_2151_0, i_8_289_2152_0, i_8_289_2154_0,
    i_8_289_2230_0, i_8_289_2235_0, i_8_289_2262_0, i_8_289_2293_0;
  output o_8_289_0_0;
  assign o_8_289_0_0 = 0;
endmodule



// Benchmark "kernel_8_290" written by ABC on Sun Jul 19 10:08:06 2020

module kernel_8_290 ( 
    i_8_290_9_0, i_8_290_135_0, i_8_290_138_0, i_8_290_139_0,
    i_8_290_151_0, i_8_290_173_0, i_8_290_181_0, i_8_290_233_0,
    i_8_290_302_0, i_8_290_392_0, i_8_290_394_0, i_8_290_398_0,
    i_8_290_401_0, i_8_290_423_0, i_8_290_424_0, i_8_290_463_0,
    i_8_290_476_0, i_8_290_506_0, i_8_290_528_0, i_8_290_532_0,
    i_8_290_538_0, i_8_290_554_0, i_8_290_568_0, i_8_290_576_0,
    i_8_290_657_0, i_8_290_670_0, i_8_290_702_0, i_8_290_748_0,
    i_8_290_815_0, i_8_290_829_0, i_8_290_833_0, i_8_290_839_0,
    i_8_290_842_0, i_8_290_890_0, i_8_290_936_0, i_8_290_964_0,
    i_8_290_968_0, i_8_290_970_0, i_8_290_1052_0, i_8_290_1197_0,
    i_8_290_1198_0, i_8_290_1199_0, i_8_290_1202_0, i_8_290_1228_0,
    i_8_290_1235_0, i_8_290_1253_0, i_8_290_1291_0, i_8_290_1296_0,
    i_8_290_1300_0, i_8_290_1314_0, i_8_290_1315_0, i_8_290_1382_0,
    i_8_290_1398_0, i_8_290_1400_0, i_8_290_1403_0, i_8_290_1404_0,
    i_8_290_1407_0, i_8_290_1436_0, i_8_290_1459_0, i_8_290_1460_0,
    i_8_290_1467_0, i_8_290_1486_0, i_8_290_1494_0, i_8_290_1512_0,
    i_8_290_1524_0, i_8_290_1525_0, i_8_290_1538_0, i_8_290_1539_0,
    i_8_290_1650_0, i_8_290_1684_0, i_8_290_1707_0, i_8_290_1708_0,
    i_8_290_1719_0, i_8_290_1720_0, i_8_290_1727_0, i_8_290_1745_0,
    i_8_290_1756_0, i_8_290_1786_0, i_8_290_1809_0, i_8_290_1825_0,
    i_8_290_1826_0, i_8_290_1840_0, i_8_290_1861_0, i_8_290_1882_0,
    i_8_290_1935_0, i_8_290_1952_0, i_8_290_1974_0, i_8_290_2012_0,
    i_8_290_2072_0, i_8_290_2096_0, i_8_290_2120_0, i_8_290_2126_0,
    i_8_290_2152_0, i_8_290_2170_0, i_8_290_2171_0, i_8_290_2177_0,
    i_8_290_2233_0, i_8_290_2253_0, i_8_290_2295_0, i_8_290_2297_0,
    o_8_290_0_0  );
  input  i_8_290_9_0, i_8_290_135_0, i_8_290_138_0, i_8_290_139_0,
    i_8_290_151_0, i_8_290_173_0, i_8_290_181_0, i_8_290_233_0,
    i_8_290_302_0, i_8_290_392_0, i_8_290_394_0, i_8_290_398_0,
    i_8_290_401_0, i_8_290_423_0, i_8_290_424_0, i_8_290_463_0,
    i_8_290_476_0, i_8_290_506_0, i_8_290_528_0, i_8_290_532_0,
    i_8_290_538_0, i_8_290_554_0, i_8_290_568_0, i_8_290_576_0,
    i_8_290_657_0, i_8_290_670_0, i_8_290_702_0, i_8_290_748_0,
    i_8_290_815_0, i_8_290_829_0, i_8_290_833_0, i_8_290_839_0,
    i_8_290_842_0, i_8_290_890_0, i_8_290_936_0, i_8_290_964_0,
    i_8_290_968_0, i_8_290_970_0, i_8_290_1052_0, i_8_290_1197_0,
    i_8_290_1198_0, i_8_290_1199_0, i_8_290_1202_0, i_8_290_1228_0,
    i_8_290_1235_0, i_8_290_1253_0, i_8_290_1291_0, i_8_290_1296_0,
    i_8_290_1300_0, i_8_290_1314_0, i_8_290_1315_0, i_8_290_1382_0,
    i_8_290_1398_0, i_8_290_1400_0, i_8_290_1403_0, i_8_290_1404_0,
    i_8_290_1407_0, i_8_290_1436_0, i_8_290_1459_0, i_8_290_1460_0,
    i_8_290_1467_0, i_8_290_1486_0, i_8_290_1494_0, i_8_290_1512_0,
    i_8_290_1524_0, i_8_290_1525_0, i_8_290_1538_0, i_8_290_1539_0,
    i_8_290_1650_0, i_8_290_1684_0, i_8_290_1707_0, i_8_290_1708_0,
    i_8_290_1719_0, i_8_290_1720_0, i_8_290_1727_0, i_8_290_1745_0,
    i_8_290_1756_0, i_8_290_1786_0, i_8_290_1809_0, i_8_290_1825_0,
    i_8_290_1826_0, i_8_290_1840_0, i_8_290_1861_0, i_8_290_1882_0,
    i_8_290_1935_0, i_8_290_1952_0, i_8_290_1974_0, i_8_290_2012_0,
    i_8_290_2072_0, i_8_290_2096_0, i_8_290_2120_0, i_8_290_2126_0,
    i_8_290_2152_0, i_8_290_2170_0, i_8_290_2171_0, i_8_290_2177_0,
    i_8_290_2233_0, i_8_290_2253_0, i_8_290_2295_0, i_8_290_2297_0;
  output o_8_290_0_0;
  assign o_8_290_0_0 = 0;
endmodule



// Benchmark "kernel_8_291" written by ABC on Sun Jul 19 10:08:08 2020

module kernel_8_291 ( 
    i_8_291_9_0, i_8_291_31_0, i_8_291_87_0, i_8_291_88_0, i_8_291_92_0,
    i_8_291_111_0, i_8_291_112_0, i_8_291_135_0, i_8_291_147_0,
    i_8_291_189_0, i_8_291_268_0, i_8_291_280_0, i_8_291_281_0,
    i_8_291_295_0, i_8_291_304_0, i_8_291_339_0, i_8_291_345_0,
    i_8_291_347_0, i_8_291_353_0, i_8_291_370_0, i_8_291_389_0,
    i_8_291_396_0, i_8_291_397_0, i_8_291_415_0, i_8_291_416_0,
    i_8_291_418_0, i_8_291_424_0, i_8_291_448_0, i_8_291_453_0,
    i_8_291_489_0, i_8_291_508_0, i_8_291_522_0, i_8_291_550_0,
    i_8_291_568_0, i_8_291_569_0, i_8_291_657_0, i_8_291_658_0,
    i_8_291_701_0, i_8_291_747_0, i_8_291_766_0, i_8_291_842_0,
    i_8_291_844_0, i_8_291_847_0, i_8_291_892_0, i_8_291_937_0,
    i_8_291_938_0, i_8_291_966_0, i_8_291_1009_0, i_8_291_1010_0,
    i_8_291_1033_0, i_8_291_1065_0, i_8_291_1098_0, i_8_291_1109_0,
    i_8_291_1142_0, i_8_291_1152_0, i_8_291_1198_0, i_8_291_1281_0,
    i_8_291_1294_0, i_8_291_1305_0, i_8_291_1352_0, i_8_291_1393_0,
    i_8_291_1404_0, i_8_291_1422_0, i_8_291_1423_0, i_8_291_1487_0,
    i_8_291_1521_0, i_8_291_1522_0, i_8_291_1523_0, i_8_291_1530_0,
    i_8_291_1543_0, i_8_291_1548_0, i_8_291_1549_0, i_8_291_1604_0,
    i_8_291_1634_0, i_8_291_1649_0, i_8_291_1669_0, i_8_291_1670_0,
    i_8_291_1683_0, i_8_291_1721_0, i_8_291_1757_0, i_8_291_1765_0,
    i_8_291_1773_0, i_8_291_1803_0, i_8_291_1855_0, i_8_291_1889_0,
    i_8_291_1935_0, i_8_291_1936_0, i_8_291_1954_0, i_8_291_1955_0,
    i_8_291_2017_0, i_8_291_2026_0, i_8_291_2039_0, i_8_291_2161_0,
    i_8_291_2173_0, i_8_291_2206_0, i_8_291_2226_0, i_8_291_2243_0,
    i_8_291_2256_0, i_8_291_2271_0, i_8_291_2297_0,
    o_8_291_0_0  );
  input  i_8_291_9_0, i_8_291_31_0, i_8_291_87_0, i_8_291_88_0,
    i_8_291_92_0, i_8_291_111_0, i_8_291_112_0, i_8_291_135_0,
    i_8_291_147_0, i_8_291_189_0, i_8_291_268_0, i_8_291_280_0,
    i_8_291_281_0, i_8_291_295_0, i_8_291_304_0, i_8_291_339_0,
    i_8_291_345_0, i_8_291_347_0, i_8_291_353_0, i_8_291_370_0,
    i_8_291_389_0, i_8_291_396_0, i_8_291_397_0, i_8_291_415_0,
    i_8_291_416_0, i_8_291_418_0, i_8_291_424_0, i_8_291_448_0,
    i_8_291_453_0, i_8_291_489_0, i_8_291_508_0, i_8_291_522_0,
    i_8_291_550_0, i_8_291_568_0, i_8_291_569_0, i_8_291_657_0,
    i_8_291_658_0, i_8_291_701_0, i_8_291_747_0, i_8_291_766_0,
    i_8_291_842_0, i_8_291_844_0, i_8_291_847_0, i_8_291_892_0,
    i_8_291_937_0, i_8_291_938_0, i_8_291_966_0, i_8_291_1009_0,
    i_8_291_1010_0, i_8_291_1033_0, i_8_291_1065_0, i_8_291_1098_0,
    i_8_291_1109_0, i_8_291_1142_0, i_8_291_1152_0, i_8_291_1198_0,
    i_8_291_1281_0, i_8_291_1294_0, i_8_291_1305_0, i_8_291_1352_0,
    i_8_291_1393_0, i_8_291_1404_0, i_8_291_1422_0, i_8_291_1423_0,
    i_8_291_1487_0, i_8_291_1521_0, i_8_291_1522_0, i_8_291_1523_0,
    i_8_291_1530_0, i_8_291_1543_0, i_8_291_1548_0, i_8_291_1549_0,
    i_8_291_1604_0, i_8_291_1634_0, i_8_291_1649_0, i_8_291_1669_0,
    i_8_291_1670_0, i_8_291_1683_0, i_8_291_1721_0, i_8_291_1757_0,
    i_8_291_1765_0, i_8_291_1773_0, i_8_291_1803_0, i_8_291_1855_0,
    i_8_291_1889_0, i_8_291_1935_0, i_8_291_1936_0, i_8_291_1954_0,
    i_8_291_1955_0, i_8_291_2017_0, i_8_291_2026_0, i_8_291_2039_0,
    i_8_291_2161_0, i_8_291_2173_0, i_8_291_2206_0, i_8_291_2226_0,
    i_8_291_2243_0, i_8_291_2256_0, i_8_291_2271_0, i_8_291_2297_0;
  output o_8_291_0_0;
  assign o_8_291_0_0 = 0;
endmodule



// Benchmark "kernel_8_292" written by ABC on Sun Jul 19 10:08:09 2020

module kernel_8_292 ( 
    i_8_292_3_0, i_8_292_35_0, i_8_292_42_0, i_8_292_43_0, i_8_292_44_0,
    i_8_292_66_0, i_8_292_79_0, i_8_292_129_0, i_8_292_138_0,
    i_8_292_141_0, i_8_292_150_0, i_8_292_190_0, i_8_292_202_0,
    i_8_292_355_0, i_8_292_384_0, i_8_292_421_0, i_8_292_498_0,
    i_8_292_499_0, i_8_292_500_0, i_8_292_507_0, i_8_292_553_0,
    i_8_292_554_0, i_8_292_594_0, i_8_292_607_0, i_8_292_624_0,
    i_8_292_642_0, i_8_292_643_0, i_8_292_656_0, i_8_292_789_0,
    i_8_292_811_0, i_8_292_828_0, i_8_292_831_0, i_8_292_840_0,
    i_8_292_876_0, i_8_292_877_0, i_8_292_880_0, i_8_292_958_0,
    i_8_292_1005_0, i_8_292_1039_0, i_8_292_1053_0, i_8_292_1083_0,
    i_8_292_1132_0, i_8_292_1155_0, i_8_292_1156_0, i_8_292_1200_0,
    i_8_292_1230_0, i_8_292_1272_0, i_8_292_1317_0, i_8_292_1318_0,
    i_8_292_1321_0, i_8_292_1326_0, i_8_292_1350_0, i_8_292_1372_0,
    i_8_292_1384_0, i_8_292_1385_0, i_8_292_1389_0, i_8_292_1390_0,
    i_8_292_1393_0, i_8_292_1399_0, i_8_292_1402_0, i_8_292_1449_0,
    i_8_292_1473_0, i_8_292_1483_0, i_8_292_1485_0, i_8_292_1486_0,
    i_8_292_1498_0, i_8_292_1503_0, i_8_292_1524_0, i_8_292_1533_0,
    i_8_292_1599_0, i_8_292_1615_0, i_8_292_1652_0, i_8_292_1654_0,
    i_8_292_1696_0, i_8_292_1753_0, i_8_292_1828_0, i_8_292_1876_0,
    i_8_292_1887_0, i_8_292_1897_0, i_8_292_1915_0, i_8_292_1950_0,
    i_8_292_1981_0, i_8_292_1996_0, i_8_292_2010_0, i_8_292_2011_0,
    i_8_292_2023_0, i_8_292_2035_0, i_8_292_2043_0, i_8_292_2053_0,
    i_8_292_2068_0, i_8_292_2082_0, i_8_292_2089_0, i_8_292_2093_0,
    i_8_292_2122_0, i_8_292_2150_0, i_8_292_2173_0, i_8_292_2185_0,
    i_8_292_2237_0, i_8_292_2249_0, i_8_292_2284_0,
    o_8_292_0_0  );
  input  i_8_292_3_0, i_8_292_35_0, i_8_292_42_0, i_8_292_43_0,
    i_8_292_44_0, i_8_292_66_0, i_8_292_79_0, i_8_292_129_0, i_8_292_138_0,
    i_8_292_141_0, i_8_292_150_0, i_8_292_190_0, i_8_292_202_0,
    i_8_292_355_0, i_8_292_384_0, i_8_292_421_0, i_8_292_498_0,
    i_8_292_499_0, i_8_292_500_0, i_8_292_507_0, i_8_292_553_0,
    i_8_292_554_0, i_8_292_594_0, i_8_292_607_0, i_8_292_624_0,
    i_8_292_642_0, i_8_292_643_0, i_8_292_656_0, i_8_292_789_0,
    i_8_292_811_0, i_8_292_828_0, i_8_292_831_0, i_8_292_840_0,
    i_8_292_876_0, i_8_292_877_0, i_8_292_880_0, i_8_292_958_0,
    i_8_292_1005_0, i_8_292_1039_0, i_8_292_1053_0, i_8_292_1083_0,
    i_8_292_1132_0, i_8_292_1155_0, i_8_292_1156_0, i_8_292_1200_0,
    i_8_292_1230_0, i_8_292_1272_0, i_8_292_1317_0, i_8_292_1318_0,
    i_8_292_1321_0, i_8_292_1326_0, i_8_292_1350_0, i_8_292_1372_0,
    i_8_292_1384_0, i_8_292_1385_0, i_8_292_1389_0, i_8_292_1390_0,
    i_8_292_1393_0, i_8_292_1399_0, i_8_292_1402_0, i_8_292_1449_0,
    i_8_292_1473_0, i_8_292_1483_0, i_8_292_1485_0, i_8_292_1486_0,
    i_8_292_1498_0, i_8_292_1503_0, i_8_292_1524_0, i_8_292_1533_0,
    i_8_292_1599_0, i_8_292_1615_0, i_8_292_1652_0, i_8_292_1654_0,
    i_8_292_1696_0, i_8_292_1753_0, i_8_292_1828_0, i_8_292_1876_0,
    i_8_292_1887_0, i_8_292_1897_0, i_8_292_1915_0, i_8_292_1950_0,
    i_8_292_1981_0, i_8_292_1996_0, i_8_292_2010_0, i_8_292_2011_0,
    i_8_292_2023_0, i_8_292_2035_0, i_8_292_2043_0, i_8_292_2053_0,
    i_8_292_2068_0, i_8_292_2082_0, i_8_292_2089_0, i_8_292_2093_0,
    i_8_292_2122_0, i_8_292_2150_0, i_8_292_2173_0, i_8_292_2185_0,
    i_8_292_2237_0, i_8_292_2249_0, i_8_292_2284_0;
  output o_8_292_0_0;
  assign o_8_292_0_0 = 0;
endmodule



// Benchmark "kernel_8_293" written by ABC on Sun Jul 19 10:08:10 2020

module kernel_8_293 ( 
    i_8_293_50_0, i_8_293_60_0, i_8_293_61_0, i_8_293_62_0, i_8_293_96_0,
    i_8_293_125_0, i_8_293_141_0, i_8_293_143_0, i_8_293_185_0,
    i_8_293_189_0, i_8_293_229_0, i_8_293_259_0, i_8_293_260_0,
    i_8_293_303_0, i_8_293_308_0, i_8_293_349_0, i_8_293_365_0,
    i_8_293_366_0, i_8_293_382_0, i_8_293_420_0, i_8_293_427_0,
    i_8_293_448_0, i_8_293_449_0, i_8_293_456_0, i_8_293_457_0,
    i_8_293_511_0, i_8_293_555_0, i_8_293_556_0, i_8_293_591_0,
    i_8_293_592_0, i_8_293_602_0, i_8_293_617_0, i_8_293_622_0,
    i_8_293_633_0, i_8_293_636_0, i_8_293_768_0, i_8_293_789_0,
    i_8_293_790_0, i_8_293_795_0, i_8_293_818_0, i_8_293_826_0,
    i_8_293_827_0, i_8_293_845_0, i_8_293_857_0, i_8_293_881_0,
    i_8_293_969_0, i_8_293_970_0, i_8_293_995_0, i_8_293_1051_0,
    i_8_293_1076_0, i_8_293_1124_0, i_8_293_1228_0, i_8_293_1237_0,
    i_8_293_1268_0, i_8_293_1282_0, i_8_293_1283_0, i_8_293_1284_0,
    i_8_293_1285_0, i_8_293_1286_0, i_8_293_1295_0, i_8_293_1314_0,
    i_8_293_1319_0, i_8_293_1331_0, i_8_293_1407_0, i_8_293_1408_0,
    i_8_293_1439_0, i_8_293_1473_0, i_8_293_1474_0, i_8_293_1484_0,
    i_8_293_1541_0, i_8_293_1547_0, i_8_293_1574_0, i_8_293_1601_0,
    i_8_293_1605_0, i_8_293_1626_0, i_8_293_1635_0, i_8_293_1648_0,
    i_8_293_1649_0, i_8_293_1653_0, i_8_293_1669_0, i_8_293_1679_0,
    i_8_293_1724_0, i_8_293_1736_0, i_8_293_1747_0, i_8_293_1773_0,
    i_8_293_1857_0, i_8_293_1948_0, i_8_293_2031_0, i_8_293_2033_0,
    i_8_293_2046_0, i_8_293_2095_0, i_8_293_2096_0, i_8_293_2151_0,
    i_8_293_2152_0, i_8_293_2217_0, i_8_293_2218_0, i_8_293_2219_0,
    i_8_293_2226_0, i_8_293_2243_0, i_8_293_2286_0,
    o_8_293_0_0  );
  input  i_8_293_50_0, i_8_293_60_0, i_8_293_61_0, i_8_293_62_0,
    i_8_293_96_0, i_8_293_125_0, i_8_293_141_0, i_8_293_143_0,
    i_8_293_185_0, i_8_293_189_0, i_8_293_229_0, i_8_293_259_0,
    i_8_293_260_0, i_8_293_303_0, i_8_293_308_0, i_8_293_349_0,
    i_8_293_365_0, i_8_293_366_0, i_8_293_382_0, i_8_293_420_0,
    i_8_293_427_0, i_8_293_448_0, i_8_293_449_0, i_8_293_456_0,
    i_8_293_457_0, i_8_293_511_0, i_8_293_555_0, i_8_293_556_0,
    i_8_293_591_0, i_8_293_592_0, i_8_293_602_0, i_8_293_617_0,
    i_8_293_622_0, i_8_293_633_0, i_8_293_636_0, i_8_293_768_0,
    i_8_293_789_0, i_8_293_790_0, i_8_293_795_0, i_8_293_818_0,
    i_8_293_826_0, i_8_293_827_0, i_8_293_845_0, i_8_293_857_0,
    i_8_293_881_0, i_8_293_969_0, i_8_293_970_0, i_8_293_995_0,
    i_8_293_1051_0, i_8_293_1076_0, i_8_293_1124_0, i_8_293_1228_0,
    i_8_293_1237_0, i_8_293_1268_0, i_8_293_1282_0, i_8_293_1283_0,
    i_8_293_1284_0, i_8_293_1285_0, i_8_293_1286_0, i_8_293_1295_0,
    i_8_293_1314_0, i_8_293_1319_0, i_8_293_1331_0, i_8_293_1407_0,
    i_8_293_1408_0, i_8_293_1439_0, i_8_293_1473_0, i_8_293_1474_0,
    i_8_293_1484_0, i_8_293_1541_0, i_8_293_1547_0, i_8_293_1574_0,
    i_8_293_1601_0, i_8_293_1605_0, i_8_293_1626_0, i_8_293_1635_0,
    i_8_293_1648_0, i_8_293_1649_0, i_8_293_1653_0, i_8_293_1669_0,
    i_8_293_1679_0, i_8_293_1724_0, i_8_293_1736_0, i_8_293_1747_0,
    i_8_293_1773_0, i_8_293_1857_0, i_8_293_1948_0, i_8_293_2031_0,
    i_8_293_2033_0, i_8_293_2046_0, i_8_293_2095_0, i_8_293_2096_0,
    i_8_293_2151_0, i_8_293_2152_0, i_8_293_2217_0, i_8_293_2218_0,
    i_8_293_2219_0, i_8_293_2226_0, i_8_293_2243_0, i_8_293_2286_0;
  output o_8_293_0_0;
  assign o_8_293_0_0 = ~((~i_8_293_60_0 & ((i_8_293_448_0 & ~i_8_293_881_0 & ~i_8_293_1547_0 & ~i_8_293_1724_0) | (~i_8_293_185_0 & ~i_8_293_1319_0 & ~i_8_293_1473_0 & ~i_8_293_1474_0 & ~i_8_293_2217_0))) | (~i_8_293_420_0 & ~i_8_293_818_0 & ((~i_8_293_365_0 & ~i_8_293_591_0 & ~i_8_293_790_0 & ~i_8_293_1124_0 & ~i_8_293_1574_0 & ~i_8_293_1649_0) | (~i_8_293_448_0 & ~i_8_293_1724_0 & ~i_8_293_2218_0))) | (~i_8_293_456_0 & ~i_8_293_1626_0 & ((~i_8_293_143_0 & ~i_8_293_457_0 & ~i_8_293_1076_0 & ~i_8_293_1228_0 & ~i_8_293_1286_0) | (~i_8_293_795_0 & ~i_8_293_881_0 & i_8_293_1484_0))) | (~i_8_293_1314_0 & ((~i_8_293_789_0 & i_8_293_969_0 & i_8_293_970_0 & ~i_8_293_2219_0) | (i_8_293_591_0 & i_8_293_1284_0 & ~i_8_293_2033_0 & ~i_8_293_2243_0))) | (~i_8_293_789_0 & (i_8_293_1286_0 | (~i_8_293_61_0 & ~i_8_293_349_0 & ~i_8_293_449_0 & ~i_8_293_2031_0))) | (~i_8_293_1474_0 & ((~i_8_293_427_0 & ~i_8_293_448_0 & ~i_8_293_511_0 & ~i_8_293_995_0) | (~i_8_293_96_0 & ~i_8_293_1407_0 & ~i_8_293_2031_0 & ~i_8_293_2033_0 & ~i_8_293_2096_0))) | (~i_8_293_1635_0 & ((~i_8_293_260_0 & ~i_8_293_2031_0 & ~i_8_293_2096_0) | (~i_8_293_50_0 & ~i_8_293_141_0 & ~i_8_293_366_0 & ~i_8_293_591_0 & ~i_8_293_1948_0 & ~i_8_293_2033_0 & ~i_8_293_2152_0))) | (~i_8_293_303_0 & i_8_293_826_0) | (i_8_293_555_0 & ~i_8_293_1574_0 & ~i_8_293_1649_0 & ~i_8_293_2151_0) | (i_8_293_1439_0 & i_8_293_2226_0));
endmodule



// Benchmark "kernel_8_294" written by ABC on Sun Jul 19 10:08:12 2020

module kernel_8_294 ( 
    i_8_294_13_0, i_8_294_63_0, i_8_294_66_0, i_8_294_75_0, i_8_294_129_0,
    i_8_294_183_0, i_8_294_204_0, i_8_294_237_0, i_8_294_309_0,
    i_8_294_336_0, i_8_294_345_0, i_8_294_354_0, i_8_294_450_0,
    i_8_294_453_0, i_8_294_475_0, i_8_294_489_0, i_8_294_490_0,
    i_8_294_504_0, i_8_294_552_0, i_8_294_555_0, i_8_294_591_0,
    i_8_294_597_0, i_8_294_608_0, i_8_294_637_0, i_8_294_658_0,
    i_8_294_662_0, i_8_294_664_0, i_8_294_682_0, i_8_294_690_0,
    i_8_294_697_0, i_8_294_728_0, i_8_294_765_0, i_8_294_768_0,
    i_8_294_769_0, i_8_294_771_0, i_8_294_795_0, i_8_294_804_0,
    i_8_294_825_0, i_8_294_921_0, i_8_294_930_0, i_8_294_933_0,
    i_8_294_970_0, i_8_294_1029_0, i_8_294_1056_0, i_8_294_1060_0,
    i_8_294_1072_0, i_8_294_1074_0, i_8_294_1089_0, i_8_294_1168_0,
    i_8_294_1173_0, i_8_294_1176_0, i_8_294_1254_0, i_8_294_1264_0,
    i_8_294_1266_0, i_8_294_1267_0, i_8_294_1275_0, i_8_294_1297_0,
    i_8_294_1305_0, i_8_294_1440_0, i_8_294_1470_0, i_8_294_1536_0,
    i_8_294_1554_0, i_8_294_1560_0, i_8_294_1563_0, i_8_294_1596_0,
    i_8_294_1605_0, i_8_294_1621_0, i_8_294_1641_0, i_8_294_1645_0,
    i_8_294_1668_0, i_8_294_1680_0, i_8_294_1704_0, i_8_294_1737_0,
    i_8_294_1747_0, i_8_294_1759_0, i_8_294_1767_0, i_8_294_1770_0,
    i_8_294_1778_0, i_8_294_1821_0, i_8_294_1830_0, i_8_294_1831_0,
    i_8_294_1857_0, i_8_294_1861_0, i_8_294_1875_0, i_8_294_1879_0,
    i_8_294_1885_0, i_8_294_1929_0, i_8_294_1965_0, i_8_294_2017_0,
    i_8_294_2019_0, i_8_294_2059_0, i_8_294_2119_0, i_8_294_2148_0,
    i_8_294_2169_0, i_8_294_2182_0, i_8_294_2184_0, i_8_294_2194_0,
    i_8_294_2211_0, i_8_294_2215_0, i_8_294_2291_0,
    o_8_294_0_0  );
  input  i_8_294_13_0, i_8_294_63_0, i_8_294_66_0, i_8_294_75_0,
    i_8_294_129_0, i_8_294_183_0, i_8_294_204_0, i_8_294_237_0,
    i_8_294_309_0, i_8_294_336_0, i_8_294_345_0, i_8_294_354_0,
    i_8_294_450_0, i_8_294_453_0, i_8_294_475_0, i_8_294_489_0,
    i_8_294_490_0, i_8_294_504_0, i_8_294_552_0, i_8_294_555_0,
    i_8_294_591_0, i_8_294_597_0, i_8_294_608_0, i_8_294_637_0,
    i_8_294_658_0, i_8_294_662_0, i_8_294_664_0, i_8_294_682_0,
    i_8_294_690_0, i_8_294_697_0, i_8_294_728_0, i_8_294_765_0,
    i_8_294_768_0, i_8_294_769_0, i_8_294_771_0, i_8_294_795_0,
    i_8_294_804_0, i_8_294_825_0, i_8_294_921_0, i_8_294_930_0,
    i_8_294_933_0, i_8_294_970_0, i_8_294_1029_0, i_8_294_1056_0,
    i_8_294_1060_0, i_8_294_1072_0, i_8_294_1074_0, i_8_294_1089_0,
    i_8_294_1168_0, i_8_294_1173_0, i_8_294_1176_0, i_8_294_1254_0,
    i_8_294_1264_0, i_8_294_1266_0, i_8_294_1267_0, i_8_294_1275_0,
    i_8_294_1297_0, i_8_294_1305_0, i_8_294_1440_0, i_8_294_1470_0,
    i_8_294_1536_0, i_8_294_1554_0, i_8_294_1560_0, i_8_294_1563_0,
    i_8_294_1596_0, i_8_294_1605_0, i_8_294_1621_0, i_8_294_1641_0,
    i_8_294_1645_0, i_8_294_1668_0, i_8_294_1680_0, i_8_294_1704_0,
    i_8_294_1737_0, i_8_294_1747_0, i_8_294_1759_0, i_8_294_1767_0,
    i_8_294_1770_0, i_8_294_1778_0, i_8_294_1821_0, i_8_294_1830_0,
    i_8_294_1831_0, i_8_294_1857_0, i_8_294_1861_0, i_8_294_1875_0,
    i_8_294_1879_0, i_8_294_1885_0, i_8_294_1929_0, i_8_294_1965_0,
    i_8_294_2017_0, i_8_294_2019_0, i_8_294_2059_0, i_8_294_2119_0,
    i_8_294_2148_0, i_8_294_2169_0, i_8_294_2182_0, i_8_294_2184_0,
    i_8_294_2194_0, i_8_294_2211_0, i_8_294_2215_0, i_8_294_2291_0;
  output o_8_294_0_0;
  assign o_8_294_0_0 = ~((~i_8_294_1875_0 & ((~i_8_294_66_0 & ((~i_8_294_63_0 & ~i_8_294_697_0 & ~i_8_294_1072_0 & ~i_8_294_1173_0 & ~i_8_294_1176_0 & ~i_8_294_1470_0) | (~i_8_294_309_0 & ~i_8_294_450_0 & ~i_8_294_804_0 & ~i_8_294_921_0 & ~i_8_294_2291_0))) | (~i_8_294_765_0 & ~i_8_294_771_0 & ~i_8_294_921_0 & i_8_294_1264_0) | (~i_8_294_336_0 & ~i_8_294_804_0 & ~i_8_294_1264_0 & ~i_8_294_1470_0 & ~i_8_294_1563_0) | (i_8_294_552_0 & i_8_294_1680_0 & ~i_8_294_1821_0))) | (~i_8_294_309_0 & ((~i_8_294_608_0 & ~i_8_294_795_0 & i_8_294_1297_0 & ~i_8_294_1605_0 & ~i_8_294_1645_0) | (i_8_294_475_0 & i_8_294_1759_0))) | (~i_8_294_795_0 & ((~i_8_294_354_0 & ((~i_8_294_768_0 & ~i_8_294_930_0 & ~i_8_294_1668_0 & i_8_294_1965_0 & ~i_8_294_2017_0 & ~i_8_294_2148_0) | (~i_8_294_552_0 & ~i_8_294_970_0 & ~i_8_294_1470_0 & ~i_8_294_1560_0 & ~i_8_294_1965_0 & ~i_8_294_2211_0))) | (~i_8_294_345_0 & ~i_8_294_504_0 & ~i_8_294_1305_0 & ~i_8_294_1645_0 & ~i_8_294_1857_0 & ~i_8_294_2211_0))) | (~i_8_294_453_0 & ~i_8_294_2184_0 & ((~i_8_294_765_0 & ~i_8_294_921_0 & ~i_8_294_1173_0 & ~i_8_294_1470_0) | (i_8_294_75_0 & ~i_8_294_1275_0 & ~i_8_294_1560_0 & ~i_8_294_1737_0 & ~i_8_294_2017_0))) | (~i_8_294_662_0 & ((~i_8_294_63_0 & i_8_294_66_0 & ~i_8_294_597_0 & ~i_8_294_765_0 & ~i_8_294_804_0 & ~i_8_294_1440_0 & ~i_8_294_1563_0) | (i_8_294_345_0 & ~i_8_294_591_0 & i_8_294_768_0 & ~i_8_294_771_0 & ~i_8_294_1254_0 & i_8_294_1560_0 & ~i_8_294_1621_0 & ~i_8_294_1857_0 & ~i_8_294_1879_0))) | (~i_8_294_690_0 & ~i_8_294_921_0 & ((~i_8_294_450_0 & ~i_8_294_765_0 & ~i_8_294_933_0 & ~i_8_294_1560_0 & ~i_8_294_1641_0 & ~i_8_294_1668_0) | (~i_8_294_13_0 & ~i_8_294_1254_0 & ~i_8_294_1305_0 & i_8_294_2148_0 & ~i_8_294_2169_0 & ~i_8_294_2215_0))) | (~i_8_294_930_0 & ((~i_8_294_1275_0 & i_8_294_1440_0 & ~i_8_294_1560_0 & ~i_8_294_1641_0) | (~i_8_294_63_0 & ~i_8_294_1056_0 & ~i_8_294_1074_0 & ~i_8_294_1264_0 & ~i_8_294_1554_0 & ~i_8_294_1621_0 & ~i_8_294_2017_0))) | (~i_8_294_1176_0 & ((~i_8_294_63_0 & ~i_8_294_1737_0 & ((~i_8_294_555_0 & ~i_8_294_1440_0 & ~i_8_294_1704_0 & i_8_294_1770_0) | (~i_8_294_765_0 & ~i_8_294_1060_0 & ~i_8_294_1254_0 & ~i_8_294_1297_0 & ~i_8_294_2017_0 & ~i_8_294_2215_0))) | (i_8_294_697_0 & ~i_8_294_765_0 & ~i_8_294_768_0 & ~i_8_294_1074_0 & ~i_8_294_1747_0 & ~i_8_294_2169_0))) | (~i_8_294_765_0 & ~i_8_294_933_0 & i_8_294_1072_0 & ~i_8_294_1254_0 & i_8_294_1470_0 & i_8_294_1645_0 & ~i_8_294_1680_0) | (~i_8_294_129_0 & ~i_8_294_1470_0 & ~i_8_294_1641_0 & ~i_8_294_1737_0 & ~i_8_294_2169_0));
endmodule



// Benchmark "kernel_8_295" written by ABC on Sun Jul 19 10:08:12 2020

module kernel_8_295 ( 
    i_8_295_1_0, i_8_295_22_0, i_8_295_73_0, i_8_295_75_0, i_8_295_115_0,
    i_8_295_137_0, i_8_295_148_0, i_8_295_226_0, i_8_295_229_0,
    i_8_295_302_0, i_8_295_319_0, i_8_295_364_0, i_8_295_380_0,
    i_8_295_388_0, i_8_295_400_0, i_8_295_425_0, i_8_295_454_0,
    i_8_295_490_0, i_8_295_497_0, i_8_295_508_0, i_8_295_528_0,
    i_8_295_552_0, i_8_295_599_0, i_8_295_602_0, i_8_295_605_0,
    i_8_295_607_0, i_8_295_635_0, i_8_295_641_0, i_8_295_659_0,
    i_8_295_660_0, i_8_295_676_0, i_8_295_680_0, i_8_295_695_0,
    i_8_295_696_0, i_8_295_706_0, i_8_295_710_0, i_8_295_757_0,
    i_8_295_814_0, i_8_295_815_0, i_8_295_860_0, i_8_295_968_0,
    i_8_295_1013_0, i_8_295_1103_0, i_8_295_1108_0, i_8_295_1111_0,
    i_8_295_1202_0, i_8_295_1228_0, i_8_295_1264_0, i_8_295_1273_0,
    i_8_295_1307_0, i_8_295_1311_0, i_8_295_1328_0, i_8_295_1358_0,
    i_8_295_1387_0, i_8_295_1388_0, i_8_295_1414_0, i_8_295_1424_0,
    i_8_295_1432_0, i_8_295_1462_0, i_8_295_1463_0, i_8_295_1466_0,
    i_8_295_1474_0, i_8_295_1478_0, i_8_295_1511_0, i_8_295_1517_0,
    i_8_295_1526_0, i_8_295_1557_0, i_8_295_1633_0, i_8_295_1648_0,
    i_8_295_1667_0, i_8_295_1678_0, i_8_295_1691_0, i_8_295_1697_0,
    i_8_295_1750_0, i_8_295_1766_0, i_8_295_1769_0, i_8_295_1772_0,
    i_8_295_1775_0, i_8_295_1787_0, i_8_295_1789_0, i_8_295_1792_0,
    i_8_295_1807_0, i_8_295_1811_0, i_8_295_1841_0, i_8_295_1846_0,
    i_8_295_1910_0, i_8_295_1927_0, i_8_295_1940_0, i_8_295_1958_0,
    i_8_295_1964_0, i_8_295_1972_0, i_8_295_1976_0, i_8_295_1981_0,
    i_8_295_1982_0, i_8_295_1997_0, i_8_295_2002_0, i_8_295_2020_0,
    i_8_295_2055_0, i_8_295_2119_0, i_8_295_2149_0,
    o_8_295_0_0  );
  input  i_8_295_1_0, i_8_295_22_0, i_8_295_73_0, i_8_295_75_0,
    i_8_295_115_0, i_8_295_137_0, i_8_295_148_0, i_8_295_226_0,
    i_8_295_229_0, i_8_295_302_0, i_8_295_319_0, i_8_295_364_0,
    i_8_295_380_0, i_8_295_388_0, i_8_295_400_0, i_8_295_425_0,
    i_8_295_454_0, i_8_295_490_0, i_8_295_497_0, i_8_295_508_0,
    i_8_295_528_0, i_8_295_552_0, i_8_295_599_0, i_8_295_602_0,
    i_8_295_605_0, i_8_295_607_0, i_8_295_635_0, i_8_295_641_0,
    i_8_295_659_0, i_8_295_660_0, i_8_295_676_0, i_8_295_680_0,
    i_8_295_695_0, i_8_295_696_0, i_8_295_706_0, i_8_295_710_0,
    i_8_295_757_0, i_8_295_814_0, i_8_295_815_0, i_8_295_860_0,
    i_8_295_968_0, i_8_295_1013_0, i_8_295_1103_0, i_8_295_1108_0,
    i_8_295_1111_0, i_8_295_1202_0, i_8_295_1228_0, i_8_295_1264_0,
    i_8_295_1273_0, i_8_295_1307_0, i_8_295_1311_0, i_8_295_1328_0,
    i_8_295_1358_0, i_8_295_1387_0, i_8_295_1388_0, i_8_295_1414_0,
    i_8_295_1424_0, i_8_295_1432_0, i_8_295_1462_0, i_8_295_1463_0,
    i_8_295_1466_0, i_8_295_1474_0, i_8_295_1478_0, i_8_295_1511_0,
    i_8_295_1517_0, i_8_295_1526_0, i_8_295_1557_0, i_8_295_1633_0,
    i_8_295_1648_0, i_8_295_1667_0, i_8_295_1678_0, i_8_295_1691_0,
    i_8_295_1697_0, i_8_295_1750_0, i_8_295_1766_0, i_8_295_1769_0,
    i_8_295_1772_0, i_8_295_1775_0, i_8_295_1787_0, i_8_295_1789_0,
    i_8_295_1792_0, i_8_295_1807_0, i_8_295_1811_0, i_8_295_1841_0,
    i_8_295_1846_0, i_8_295_1910_0, i_8_295_1927_0, i_8_295_1940_0,
    i_8_295_1958_0, i_8_295_1964_0, i_8_295_1972_0, i_8_295_1976_0,
    i_8_295_1981_0, i_8_295_1982_0, i_8_295_1997_0, i_8_295_2002_0,
    i_8_295_2020_0, i_8_295_2055_0, i_8_295_2119_0, i_8_295_2149_0;
  output o_8_295_0_0;
  assign o_8_295_0_0 = 0;
endmodule



// Benchmark "kernel_8_296" written by ABC on Sun Jul 19 10:08:14 2020

module kernel_8_296 ( 
    i_8_296_0_0, i_8_296_1_0, i_8_296_104_0, i_8_296_155_0, i_8_296_163_0,
    i_8_296_216_0, i_8_296_232_0, i_8_296_233_0, i_8_296_262_0,
    i_8_296_289_0, i_8_296_325_0, i_8_296_326_0, i_8_296_366_0,
    i_8_296_432_0, i_8_296_433_0, i_8_296_480_0, i_8_296_481_0,
    i_8_296_486_0, i_8_296_489_0, i_8_296_550_0, i_8_296_556_0,
    i_8_296_603_0, i_8_296_621_0, i_8_296_630_0, i_8_296_694_0,
    i_8_296_695_0, i_8_296_696_0, i_8_296_697_0, i_8_296_701_0,
    i_8_296_709_0, i_8_296_721_0, i_8_296_783_0, i_8_296_802_0,
    i_8_296_811_0, i_8_296_812_0, i_8_296_820_0, i_8_296_825_0,
    i_8_296_827_0, i_8_296_840_0, i_8_296_865_0, i_8_296_874_0,
    i_8_296_967_0, i_8_296_970_0, i_8_296_973_0, i_8_296_996_0,
    i_8_296_1071_0, i_8_296_1154_0, i_8_296_1180_0, i_8_296_1207_0,
    i_8_296_1208_0, i_8_296_1224_0, i_8_296_1233_0, i_8_296_1234_0,
    i_8_296_1260_0, i_8_296_1270_0, i_8_296_1352_0, i_8_296_1360_0,
    i_8_296_1367_0, i_8_296_1387_0, i_8_296_1399_0, i_8_296_1435_0,
    i_8_296_1452_0, i_8_296_1537_0, i_8_296_1542_0, i_8_296_1548_0,
    i_8_296_1571_0, i_8_296_1584_0, i_8_296_1585_0, i_8_296_1622_0,
    i_8_296_1624_0, i_8_296_1650_0, i_8_296_1651_0, i_8_296_1720_0,
    i_8_296_1747_0, i_8_296_1770_0, i_8_296_1774_0, i_8_296_1818_0,
    i_8_296_1864_0, i_8_296_1874_0, i_8_296_1989_0, i_8_296_2025_0,
    i_8_296_2026_0, i_8_296_2034_0, i_8_296_2035_0, i_8_296_2038_0,
    i_8_296_2088_0, i_8_296_2116_0, i_8_296_2144_0, i_8_296_2147_0,
    i_8_296_2152_0, i_8_296_2153_0, i_8_296_2155_0, i_8_296_2188_0,
    i_8_296_2269_0, i_8_296_2272_0, i_8_296_2279_0, i_8_296_2281_0,
    i_8_296_2286_0, i_8_296_2289_0, i_8_296_2297_0,
    o_8_296_0_0  );
  input  i_8_296_0_0, i_8_296_1_0, i_8_296_104_0, i_8_296_155_0,
    i_8_296_163_0, i_8_296_216_0, i_8_296_232_0, i_8_296_233_0,
    i_8_296_262_0, i_8_296_289_0, i_8_296_325_0, i_8_296_326_0,
    i_8_296_366_0, i_8_296_432_0, i_8_296_433_0, i_8_296_480_0,
    i_8_296_481_0, i_8_296_486_0, i_8_296_489_0, i_8_296_550_0,
    i_8_296_556_0, i_8_296_603_0, i_8_296_621_0, i_8_296_630_0,
    i_8_296_694_0, i_8_296_695_0, i_8_296_696_0, i_8_296_697_0,
    i_8_296_701_0, i_8_296_709_0, i_8_296_721_0, i_8_296_783_0,
    i_8_296_802_0, i_8_296_811_0, i_8_296_812_0, i_8_296_820_0,
    i_8_296_825_0, i_8_296_827_0, i_8_296_840_0, i_8_296_865_0,
    i_8_296_874_0, i_8_296_967_0, i_8_296_970_0, i_8_296_973_0,
    i_8_296_996_0, i_8_296_1071_0, i_8_296_1154_0, i_8_296_1180_0,
    i_8_296_1207_0, i_8_296_1208_0, i_8_296_1224_0, i_8_296_1233_0,
    i_8_296_1234_0, i_8_296_1260_0, i_8_296_1270_0, i_8_296_1352_0,
    i_8_296_1360_0, i_8_296_1367_0, i_8_296_1387_0, i_8_296_1399_0,
    i_8_296_1435_0, i_8_296_1452_0, i_8_296_1537_0, i_8_296_1542_0,
    i_8_296_1548_0, i_8_296_1571_0, i_8_296_1584_0, i_8_296_1585_0,
    i_8_296_1622_0, i_8_296_1624_0, i_8_296_1650_0, i_8_296_1651_0,
    i_8_296_1720_0, i_8_296_1747_0, i_8_296_1770_0, i_8_296_1774_0,
    i_8_296_1818_0, i_8_296_1864_0, i_8_296_1874_0, i_8_296_1989_0,
    i_8_296_2025_0, i_8_296_2026_0, i_8_296_2034_0, i_8_296_2035_0,
    i_8_296_2038_0, i_8_296_2088_0, i_8_296_2116_0, i_8_296_2144_0,
    i_8_296_2147_0, i_8_296_2152_0, i_8_296_2153_0, i_8_296_2155_0,
    i_8_296_2188_0, i_8_296_2269_0, i_8_296_2272_0, i_8_296_2279_0,
    i_8_296_2281_0, i_8_296_2286_0, i_8_296_2289_0, i_8_296_2297_0;
  output o_8_296_0_0;
  assign o_8_296_0_0 = ~((~i_8_296_1234_0 & ((~i_8_296_0_0 & ~i_8_296_2038_0 & ((~i_8_296_326_0 & ~i_8_296_481_0 & ~i_8_296_550_0 & ~i_8_296_802_0 & ~i_8_296_1154_0 & ~i_8_296_1270_0 & ~i_8_296_1387_0 & ~i_8_296_1399_0 & ~i_8_296_1770_0 & ~i_8_296_2279_0) | (~i_8_296_155_0 & ~i_8_296_163_0 & i_8_296_325_0 & ~i_8_296_865_0 & ~i_8_296_1435_0 & ~i_8_296_1864_0 & ~i_8_296_2035_0 & ~i_8_296_2155_0 & ~i_8_296_2286_0))) | (~i_8_296_2144_0 & ((~i_8_296_155_0 & ((i_8_296_289_0 & ~i_8_296_366_0 & ~i_8_296_2272_0 & ~i_8_296_2279_0) | (~i_8_296_216_0 & ~i_8_296_232_0 & ~i_8_296_550_0 & ~i_8_296_996_0 & ~i_8_296_1270_0 & ~i_8_296_1360_0 & ~i_8_296_1864_0 & ~i_8_296_2188_0 & ~i_8_296_2281_0 & ~i_8_296_2286_0))) | (~i_8_296_1154_0 & ((~i_8_296_289_0 & ~i_8_296_630_0 & ~i_8_296_1720_0 & ~i_8_296_2035_0 & ~i_8_296_2088_0 & ~i_8_296_2269_0 & ~i_8_296_2279_0) | (~i_8_296_1233_0 & i_8_296_1435_0 & ~i_8_296_1770_0 & ~i_8_296_1774_0 & ~i_8_296_2025_0 & ~i_8_296_2297_0))) | (~i_8_296_366_0 & ~i_8_296_812_0 & ~i_8_296_865_0 & i_8_296_874_0 & ~i_8_296_1542_0 & ~i_8_296_1584_0 & ~i_8_296_1585_0 & ~i_8_296_1624_0 & ~i_8_296_2025_0))) | (~i_8_296_603_0 & ~i_8_296_2297_0 & ((~i_8_296_155_0 & ~i_8_296_325_0 & ~i_8_296_721_0 & ~i_8_296_825_0 & ~i_8_296_1260_0 & ~i_8_296_1360_0 & ~i_8_296_1571_0 & ~i_8_296_1747_0 & ~i_8_296_1774_0 & ~i_8_296_1989_0 & ~i_8_296_2034_0 & ~i_8_296_2155_0) | (~i_8_296_694_0 & ~i_8_296_695_0 & ~i_8_296_820_0 & ~i_8_296_967_0 & ~i_8_296_996_0 & ~i_8_296_1542_0 & ~i_8_296_1864_0 & ~i_8_296_2025_0 & ~i_8_296_2035_0 & ~i_8_296_2279_0))) | (~i_8_296_802_0 & ((~i_8_296_1154_0 & ((~i_8_296_820_0 & ~i_8_296_1571_0 & ~i_8_296_1624_0 & ~i_8_296_1989_0 & i_8_296_2152_0) | (~i_8_296_233_0 & ~i_8_296_973_0 & ~i_8_296_1399_0 & ~i_8_296_1435_0 & ~i_8_296_1720_0 & ~i_8_296_1818_0 & ~i_8_296_2035_0 & ~i_8_296_2153_0 & ~i_8_296_2286_0))) | (~i_8_296_489_0 & ~i_8_296_694_0 & ~i_8_296_865_0 & ~i_8_296_996_0 & ~i_8_296_2116_0 & ~i_8_296_2152_0 & i_8_296_2155_0 & ~i_8_296_2269_0 & ~i_8_296_2289_0))) | (~i_8_296_1367_0 & ((i_8_296_480_0 & i_8_296_481_0 & ~i_8_296_721_0 & ~i_8_296_840_0 & ~i_8_296_1624_0 & ~i_8_296_2025_0 & ~i_8_296_2026_0 & ~i_8_296_2088_0 & ~i_8_296_2279_0) | (~i_8_296_326_0 & ~i_8_296_812_0 & ~i_8_296_1747_0 & ~i_8_296_1864_0 & i_8_296_2153_0 & ~i_8_296_2281_0))) | (i_8_296_696_0 & i_8_296_840_0 & ~i_8_296_1224_0 & ~i_8_296_1270_0 & ~i_8_296_1548_0 & ~i_8_296_1864_0 & ~i_8_296_2026_0))) | (~i_8_296_1154_0 & ((~i_8_296_432_0 & ((~i_8_296_104_0 & ((i_8_296_216_0 & ~i_8_296_486_0 & ~i_8_296_630_0 & ~i_8_296_802_0 & i_8_296_874_0 & ~i_8_296_1452_0 & ~i_8_296_2144_0 & ~i_8_296_2286_0) | (~i_8_296_1_0 & ~i_8_296_163_0 & ~i_8_296_366_0 & ~i_8_296_550_0 & ~i_8_296_812_0 & ~i_8_296_820_0 & ~i_8_296_973_0 & ~i_8_296_1387_0 & ~i_8_296_1584_0 & ~i_8_296_1864_0 & ~i_8_296_2025_0 & ~i_8_296_2147_0 & ~i_8_296_2153_0 & ~i_8_296_2279_0 & ~i_8_296_2289_0))) | (~i_8_296_163_0 & ~i_8_296_232_0 & ~i_8_296_556_0 & ~i_8_296_812_0 & ~i_8_296_820_0 & ~i_8_296_825_0 & ~i_8_296_865_0 & ~i_8_296_1270_0 & ~i_8_296_1360_0 & ~i_8_296_1747_0 & ~i_8_296_1774_0 & ~i_8_296_1864_0 & ~i_8_296_2155_0 & ~i_8_296_2279_0))) | (~i_8_296_1_0 & ~i_8_296_326_0 & ((~i_8_296_232_0 & ~i_8_296_289_0 & ~i_8_296_433_0 & ~i_8_296_696_0 & ~i_8_296_1360_0 & ~i_8_296_1537_0 & ~i_8_296_1571_0 & ~i_8_296_1989_0 & ~i_8_296_2026_0 & ~i_8_296_2034_0 & ~i_8_296_2035_0 & ~i_8_296_2144_0) | (~i_8_296_163_0 & i_8_296_216_0 & ~i_8_296_262_0 & ~i_8_296_489_0 & ~i_8_296_556_0 & i_8_296_840_0 & ~i_8_296_1071_0 & ~i_8_296_1387_0 & ~i_8_296_1622_0 & ~i_8_296_2088_0 & ~i_8_296_2279_0))) | (~i_8_296_697_0 & ((~i_8_296_233_0 & ~i_8_296_721_0 & ~i_8_296_802_0 & ~i_8_296_840_0 & ~i_8_296_1224_0 & ~i_8_296_1399_0 & ~i_8_296_1624_0 & ~i_8_296_1770_0 & ~i_8_296_2116_0 & ~i_8_296_2155_0 & i_8_296_2272_0) | (~i_8_296_481_0 & ~i_8_296_820_0 & ~i_8_296_973_0 & ~i_8_296_1387_0 & ~i_8_296_1542_0 & ~i_8_296_1571_0 & ~i_8_296_1747_0 & ~i_8_296_1774_0 & ~i_8_296_2025_0 & ~i_8_296_2035_0 & ~i_8_296_2147_0 & ~i_8_296_2289_0))) | (~i_8_296_802_0 & ~i_8_296_2026_0 & ~i_8_296_2279_0 & ((~i_8_296_216_0 & ~i_8_296_325_0 & ~i_8_296_550_0 & ~i_8_296_1270_0 & ~i_8_296_1367_0 & ~i_8_296_1650_0 & ~i_8_296_1818_0 & i_8_296_2147_0) | (~i_8_296_163_0 & ~i_8_296_1224_0 & i_8_296_1260_0 & ~i_8_296_1360_0 & ~i_8_296_2269_0))))) | (~i_8_296_104_0 & ~i_8_296_289_0 & ~i_8_296_697_0 & ((~i_8_296_432_0 & ~i_8_296_433_0 & ~i_8_296_486_0 & i_8_296_550_0 & ~i_8_296_1270_0 & ~i_8_296_1452_0 & ~i_8_296_1571_0 & ~i_8_296_1774_0 & ~i_8_296_2144_0 & ~i_8_296_2279_0) | (i_8_296_216_0 & i_8_296_481_0 & ~i_8_296_996_0 & ~i_8_296_1360_0 & ~i_8_296_1585_0 & ~i_8_296_1650_0 & ~i_8_296_1770_0 & ~i_8_296_1989_0 & ~i_8_296_2116_0 & ~i_8_296_2297_0))) | (~i_8_296_1270_0 & ((~i_8_296_163_0 & ~i_8_296_2289_0 & ((~i_8_296_433_0 & i_8_296_694_0 & ~i_8_296_802_0 & ~i_8_296_820_0 & ~i_8_296_996_0 & ~i_8_296_2026_0 & ~i_8_296_2035_0 & ~i_8_296_2144_0 & ~i_8_296_2188_0) | (~i_8_296_550_0 & ~i_8_296_973_0 & ~i_8_296_1352_0 & i_8_296_1399_0 & ~i_8_296_1571_0 & ~i_8_296_1584_0 & ~i_8_296_1624_0 & ~i_8_296_2038_0 & ~i_8_296_2297_0))) | (i_8_296_874_0 & ~i_8_296_1360_0 & ((~i_8_296_366_0 & ~i_8_296_432_0 & i_8_296_696_0 & ~i_8_296_721_0 & ~i_8_296_973_0 & ~i_8_296_1260_0 & ~i_8_296_1367_0 & ~i_8_296_2188_0) | (~i_8_296_696_0 & ~i_8_296_820_0 & ~i_8_296_1537_0 & ~i_8_296_2026_0 & ~i_8_296_2269_0 & ~i_8_296_2297_0))) | (~i_8_296_603_0 & ~i_8_296_701_0 & i_8_296_967_0 & ~i_8_296_970_0 & ~i_8_296_2035_0 & ~i_8_296_2144_0 & ~i_8_296_2269_0 & ~i_8_296_2297_0))) | (~i_8_296_233_0 & ~i_8_296_2035_0 & ~i_8_296_2147_0 & ((~i_8_296_1_0 & ~i_8_296_155_0 & ~i_8_296_325_0 & i_8_296_480_0 & ~i_8_296_694_0 & ~i_8_296_1180_0 & ~i_8_296_1367_0 & ~i_8_296_1624_0 & ~i_8_296_1818_0 & ~i_8_296_2188_0) | (~i_8_296_486_0 & ~i_8_296_630_0 & ~i_8_296_802_0 & ~i_8_296_820_0 & ~i_8_296_1233_0 & ~i_8_296_1387_0 & ~i_8_296_1864_0 & ~i_8_296_1989_0 & ~i_8_296_2026_0 & ~i_8_296_2144_0 & ~i_8_296_2279_0))) | (~i_8_296_820_0 & ((~i_8_296_550_0 & ~i_8_296_1774_0 & ~i_8_296_2279_0 & ((~i_8_296_802_0 & i_8_296_1770_0 & ~i_8_296_1864_0 & ~i_8_296_2144_0) | (~i_8_296_1360_0 & ~i_8_296_1537_0 & ~i_8_296_694_0 & ~i_8_296_811_0 & ~i_8_296_1720_0 & ~i_8_296_2025_0 & ~i_8_296_2026_0 & ~i_8_296_2088_0 & ~i_8_296_2269_0))) | (~i_8_296_366_0 & ~i_8_296_630_0 & ~i_8_296_694_0 & i_8_296_709_0 & ~i_8_296_1387_0 & ~i_8_296_1571_0 & ~i_8_296_1622_0 & ~i_8_296_2116_0 & ~i_8_296_2286_0))) | (~i_8_296_695_0 & ~i_8_296_802_0 & ((~i_8_296_550_0 & ~i_8_296_1352_0 & ~i_8_296_1747_0 & i_8_296_1774_0 & ~i_8_296_1989_0 & ~i_8_296_2026_0) | (~i_8_296_996_0 & ~i_8_296_1224_0 & ~i_8_296_1774_0 & ~i_8_296_1864_0 & ~i_8_296_2144_0 & i_8_296_2152_0 & ~i_8_296_2297_0))));
endmodule



// Benchmark "kernel_8_297" written by ABC on Sun Jul 19 10:08:15 2020

module kernel_8_297 ( 
    i_8_297_29_0, i_8_297_82_0, i_8_297_100_0, i_8_297_154_0,
    i_8_297_162_0, i_8_297_171_0, i_8_297_175_0, i_8_297_190_0,
    i_8_297_218_0, i_8_297_257_0, i_8_297_259_0, i_8_297_266_0,
    i_8_297_281_0, i_8_297_339_0, i_8_297_379_0, i_8_297_380_0,
    i_8_297_427_0, i_8_297_436_0, i_8_297_437_0, i_8_297_459_0,
    i_8_297_478_0, i_8_297_572_0, i_8_297_587_0, i_8_297_598_0,
    i_8_297_621_0, i_8_297_626_0, i_8_297_684_0, i_8_297_696_0,
    i_8_297_703_0, i_8_297_707_0, i_8_297_716_0, i_8_297_757_0,
    i_8_297_761_0, i_8_297_775_0, i_8_297_778_0, i_8_297_802_0,
    i_8_297_821_0, i_8_297_876_0, i_8_297_991_0, i_8_297_992_0,
    i_8_297_1108_0, i_8_297_1111_0, i_8_297_1135_0, i_8_297_1136_0,
    i_8_297_1153_0, i_8_297_1157_0, i_8_297_1170_0, i_8_297_1180_0,
    i_8_297_1261_0, i_8_297_1279_0, i_8_297_1283_0, i_8_297_1306_0,
    i_8_297_1325_0, i_8_297_1352_0, i_8_297_1370_0, i_8_297_1381_0,
    i_8_297_1405_0, i_8_297_1407_0, i_8_297_1418_0, i_8_297_1433_0,
    i_8_297_1460_0, i_8_297_1472_0, i_8_297_1481_0, i_8_297_1487_0,
    i_8_297_1551_0, i_8_297_1568_0, i_8_297_1603_0, i_8_297_1611_0,
    i_8_297_1625_0, i_8_297_1642_0, i_8_297_1669_0, i_8_297_1675_0,
    i_8_297_1697_0, i_8_297_1737_0, i_8_297_1753_0, i_8_297_1759_0,
    i_8_297_1773_0, i_8_297_1774_0, i_8_297_1801_0, i_8_297_1805_0,
    i_8_297_1811_0, i_8_297_1823_0, i_8_297_1928_0, i_8_297_1946_0,
    i_8_297_1981_0, i_8_297_1992_0, i_8_297_1994_0, i_8_297_2054_0,
    i_8_297_2107_0, i_8_297_2112_0, i_8_297_2150_0, i_8_297_2151_0,
    i_8_297_2152_0, i_8_297_2189_0, i_8_297_2225_0, i_8_297_2241_0,
    i_8_297_2259_0, i_8_297_2287_0, i_8_297_2288_0, i_8_297_2299_0,
    o_8_297_0_0  );
  input  i_8_297_29_0, i_8_297_82_0, i_8_297_100_0, i_8_297_154_0,
    i_8_297_162_0, i_8_297_171_0, i_8_297_175_0, i_8_297_190_0,
    i_8_297_218_0, i_8_297_257_0, i_8_297_259_0, i_8_297_266_0,
    i_8_297_281_0, i_8_297_339_0, i_8_297_379_0, i_8_297_380_0,
    i_8_297_427_0, i_8_297_436_0, i_8_297_437_0, i_8_297_459_0,
    i_8_297_478_0, i_8_297_572_0, i_8_297_587_0, i_8_297_598_0,
    i_8_297_621_0, i_8_297_626_0, i_8_297_684_0, i_8_297_696_0,
    i_8_297_703_0, i_8_297_707_0, i_8_297_716_0, i_8_297_757_0,
    i_8_297_761_0, i_8_297_775_0, i_8_297_778_0, i_8_297_802_0,
    i_8_297_821_0, i_8_297_876_0, i_8_297_991_0, i_8_297_992_0,
    i_8_297_1108_0, i_8_297_1111_0, i_8_297_1135_0, i_8_297_1136_0,
    i_8_297_1153_0, i_8_297_1157_0, i_8_297_1170_0, i_8_297_1180_0,
    i_8_297_1261_0, i_8_297_1279_0, i_8_297_1283_0, i_8_297_1306_0,
    i_8_297_1325_0, i_8_297_1352_0, i_8_297_1370_0, i_8_297_1381_0,
    i_8_297_1405_0, i_8_297_1407_0, i_8_297_1418_0, i_8_297_1433_0,
    i_8_297_1460_0, i_8_297_1472_0, i_8_297_1481_0, i_8_297_1487_0,
    i_8_297_1551_0, i_8_297_1568_0, i_8_297_1603_0, i_8_297_1611_0,
    i_8_297_1625_0, i_8_297_1642_0, i_8_297_1669_0, i_8_297_1675_0,
    i_8_297_1697_0, i_8_297_1737_0, i_8_297_1753_0, i_8_297_1759_0,
    i_8_297_1773_0, i_8_297_1774_0, i_8_297_1801_0, i_8_297_1805_0,
    i_8_297_1811_0, i_8_297_1823_0, i_8_297_1928_0, i_8_297_1946_0,
    i_8_297_1981_0, i_8_297_1992_0, i_8_297_1994_0, i_8_297_2054_0,
    i_8_297_2107_0, i_8_297_2112_0, i_8_297_2150_0, i_8_297_2151_0,
    i_8_297_2152_0, i_8_297_2189_0, i_8_297_2225_0, i_8_297_2241_0,
    i_8_297_2259_0, i_8_297_2287_0, i_8_297_2288_0, i_8_297_2299_0;
  output o_8_297_0_0;
  assign o_8_297_0_0 = 0;
endmodule



// Benchmark "kernel_8_298" written by ABC on Sun Jul 19 10:08:16 2020

module kernel_8_298 ( 
    i_8_298_0_0, i_8_298_1_0, i_8_298_40_0, i_8_298_79_0, i_8_298_83_0,
    i_8_298_104_0, i_8_298_112_0, i_8_298_143_0, i_8_298_166_0,
    i_8_298_167_0, i_8_298_190_0, i_8_298_208_0, i_8_298_259_0,
    i_8_298_265_0, i_8_298_280_0, i_8_298_281_0, i_8_298_289_0,
    i_8_298_290_0, i_8_298_299_0, i_8_298_308_0, i_8_298_310_0,
    i_8_298_317_0, i_8_298_319_0, i_8_298_418_0, i_8_298_424_0,
    i_8_298_437_0, i_8_298_451_0, i_8_298_488_0, i_8_298_585_0,
    i_8_298_589_0, i_8_298_641_0, i_8_298_651_0, i_8_298_670_0,
    i_8_298_693_0, i_8_298_701_0, i_8_298_703_0, i_8_298_704_0,
    i_8_298_710_0, i_8_298_730_0, i_8_298_767_0, i_8_298_778_0,
    i_8_298_779_0, i_8_298_824_0, i_8_298_847_0, i_8_298_929_0,
    i_8_298_967_0, i_8_298_976_0, i_8_298_991_0, i_8_298_992_0,
    i_8_298_1028_0, i_8_298_1180_0, i_8_298_1234_0, i_8_298_1235_0,
    i_8_298_1256_0, i_8_298_1262_0, i_8_298_1283_0, i_8_298_1300_0,
    i_8_298_1316_0, i_8_298_1330_0, i_8_298_1352_0, i_8_298_1360_0,
    i_8_298_1384_0, i_8_298_1405_0, i_8_298_1438_0, i_8_298_1441_0,
    i_8_298_1442_0, i_8_298_1459_0, i_8_298_1486_0, i_8_298_1507_0,
    i_8_298_1541_0, i_8_298_1558_0, i_8_298_1585_0, i_8_298_1586_0,
    i_8_298_1639_0, i_8_298_1651_0, i_8_298_1682_0, i_8_298_1765_0,
    i_8_298_1766_0, i_8_298_1811_0, i_8_298_1823_0, i_8_298_1824_0,
    i_8_298_1838_0, i_8_298_1846_0, i_8_298_1982_0, i_8_298_1993_0,
    i_8_298_1994_0, i_8_298_1999_0, i_8_298_2026_0, i_8_298_2053_0,
    i_8_298_2074_0, i_8_298_2125_0, i_8_298_2126_0, i_8_298_2147_0,
    i_8_298_2158_0, i_8_298_2188_0, i_8_298_2189_0, i_8_298_2196_0,
    i_8_298_2224_0, i_8_298_2233_0, i_8_298_2242_0,
    o_8_298_0_0  );
  input  i_8_298_0_0, i_8_298_1_0, i_8_298_40_0, i_8_298_79_0,
    i_8_298_83_0, i_8_298_104_0, i_8_298_112_0, i_8_298_143_0,
    i_8_298_166_0, i_8_298_167_0, i_8_298_190_0, i_8_298_208_0,
    i_8_298_259_0, i_8_298_265_0, i_8_298_280_0, i_8_298_281_0,
    i_8_298_289_0, i_8_298_290_0, i_8_298_299_0, i_8_298_308_0,
    i_8_298_310_0, i_8_298_317_0, i_8_298_319_0, i_8_298_418_0,
    i_8_298_424_0, i_8_298_437_0, i_8_298_451_0, i_8_298_488_0,
    i_8_298_585_0, i_8_298_589_0, i_8_298_641_0, i_8_298_651_0,
    i_8_298_670_0, i_8_298_693_0, i_8_298_701_0, i_8_298_703_0,
    i_8_298_704_0, i_8_298_710_0, i_8_298_730_0, i_8_298_767_0,
    i_8_298_778_0, i_8_298_779_0, i_8_298_824_0, i_8_298_847_0,
    i_8_298_929_0, i_8_298_967_0, i_8_298_976_0, i_8_298_991_0,
    i_8_298_992_0, i_8_298_1028_0, i_8_298_1180_0, i_8_298_1234_0,
    i_8_298_1235_0, i_8_298_1256_0, i_8_298_1262_0, i_8_298_1283_0,
    i_8_298_1300_0, i_8_298_1316_0, i_8_298_1330_0, i_8_298_1352_0,
    i_8_298_1360_0, i_8_298_1384_0, i_8_298_1405_0, i_8_298_1438_0,
    i_8_298_1441_0, i_8_298_1442_0, i_8_298_1459_0, i_8_298_1486_0,
    i_8_298_1507_0, i_8_298_1541_0, i_8_298_1558_0, i_8_298_1585_0,
    i_8_298_1586_0, i_8_298_1639_0, i_8_298_1651_0, i_8_298_1682_0,
    i_8_298_1765_0, i_8_298_1766_0, i_8_298_1811_0, i_8_298_1823_0,
    i_8_298_1824_0, i_8_298_1838_0, i_8_298_1846_0, i_8_298_1982_0,
    i_8_298_1993_0, i_8_298_1994_0, i_8_298_1999_0, i_8_298_2026_0,
    i_8_298_2053_0, i_8_298_2074_0, i_8_298_2125_0, i_8_298_2126_0,
    i_8_298_2147_0, i_8_298_2158_0, i_8_298_2188_0, i_8_298_2189_0,
    i_8_298_2196_0, i_8_298_2224_0, i_8_298_2233_0, i_8_298_2242_0;
  output o_8_298_0_0;
  assign o_8_298_0_0 = ~((~i_8_298_1838_0 & ((~i_8_298_166_0 & ((~i_8_298_280_0 & ~i_8_298_281_0 & ~i_8_298_693_0 & ~i_8_298_1235_0 & ~i_8_298_1459_0 & ~i_8_298_2126_0) | (~i_8_298_730_0 & ~i_8_298_1316_0 & ~i_8_298_1352_0 & ~i_8_298_1486_0 & ~i_8_298_1982_0 & ~i_8_298_1994_0 & ~i_8_298_2189_0))) | (~i_8_298_641_0 & i_8_298_991_0 & ~i_8_298_1262_0 & ~i_8_298_2188_0))) | (~i_8_298_1459_0 & ((~i_8_298_641_0 & ((~i_8_298_280_0 & ~i_8_298_1586_0 & ((~i_8_298_289_0 & ~i_8_298_317_0 & ~i_8_298_1234_0 & ~i_8_298_1846_0) | (~i_8_298_265_0 & ~i_8_298_281_0 & ~i_8_298_1441_0 & ~i_8_298_1442_0 & ~i_8_298_2188_0))) | (~i_8_298_585_0 & ~i_8_298_1028_0 & i_8_298_1405_0 & ~i_8_298_1765_0 & ~i_8_298_1766_0))) | (~i_8_298_208_0 & ~i_8_298_281_0 & ~i_8_298_290_0 & ~i_8_298_1360_0 & ~i_8_298_1442_0 & ~i_8_298_1811_0 & i_8_298_1994_0) | (~i_8_298_299_0 & ~i_8_298_1028_0 & ~i_8_298_1180_0 & ~i_8_298_1256_0 & ~i_8_298_2189_0))) | (~i_8_298_290_0 & ((~i_8_298_83_0 & ~i_8_298_289_0 & ~i_8_298_317_0 & ~i_8_298_730_0 & ~i_8_298_967_0 & ~i_8_298_1405_0) | (i_8_298_424_0 & ~i_8_298_1262_0 & ~i_8_298_2026_0 & ~i_8_298_2188_0 & ~i_8_298_2189_0))) | (~i_8_298_585_0 & ((i_8_298_710_0 & ~i_8_298_1180_0 & i_8_298_1300_0 & ~i_8_298_1541_0 & ~i_8_298_2158_0) | (~i_8_298_104_0 & ~i_8_298_589_0 & ~i_8_298_778_0 & ~i_8_298_1283_0 & ~i_8_298_1765_0 & ~i_8_298_2196_0))) | (~i_8_298_281_0 & ((~i_8_298_1585_0 & ((~i_8_298_778_0 & ~i_8_298_1316_0 & ~i_8_298_2026_0 & i_8_298_2147_0) | (~i_8_298_437_0 & ~i_8_298_1262_0 & ~i_8_298_1438_0 & ~i_8_298_1993_0 & ~i_8_298_2074_0 & ~i_8_298_2188_0))) | (~i_8_298_317_0 & ~i_8_298_824_0 & ~i_8_298_847_0 & ~i_8_298_1360_0 & ~i_8_298_1766_0 & ~i_8_298_2189_0))) | (~i_8_298_704_0 & ~i_8_298_779_0 & ~i_8_298_929_0 & ~i_8_298_1028_0 & ~i_8_298_1651_0 & ~i_8_298_1765_0 & ~i_8_298_2188_0) | (i_8_298_418_0 & i_8_298_2196_0));
endmodule



// Benchmark "kernel_8_299" written by ABC on Sun Jul 19 10:08:17 2020

module kernel_8_299 ( 
    i_8_299_31_0, i_8_299_89_0, i_8_299_96_0, i_8_299_98_0, i_8_299_196_0,
    i_8_299_237_0, i_8_299_240_0, i_8_299_241_0, i_8_299_295_0,
    i_8_299_296_0, i_8_299_312_0, i_8_299_324_0, i_8_299_349_0,
    i_8_299_372_0, i_8_299_424_0, i_8_299_480_0, i_8_299_528_0,
    i_8_299_529_0, i_8_299_556_0, i_8_299_605_0, i_8_299_733_0,
    i_8_299_735_0, i_8_299_736_0, i_8_299_763_0, i_8_299_778_0,
    i_8_299_779_0, i_8_299_781_0, i_8_299_789_0, i_8_299_797_0,
    i_8_299_815_0, i_8_299_837_0, i_8_299_862_0, i_8_299_940_0,
    i_8_299_941_0, i_8_299_943_0, i_8_299_947_0, i_8_299_996_0,
    i_8_299_1005_0, i_8_299_1012_0, i_8_299_1015_0, i_8_299_1060_0,
    i_8_299_1114_0, i_8_299_1115_0, i_8_299_1127_0, i_8_299_1130_0,
    i_8_299_1195_0, i_8_299_1219_0, i_8_299_1223_0, i_8_299_1292_0,
    i_8_299_1294_0, i_8_299_1306_0, i_8_299_1307_0, i_8_299_1310_0,
    i_8_299_1311_0, i_8_299_1314_0, i_8_299_1336_0, i_8_299_1410_0,
    i_8_299_1438_0, i_8_299_1472_0, i_8_299_1537_0, i_8_299_1538_0,
    i_8_299_1544_0, i_8_299_1597_0, i_8_299_1609_0, i_8_299_1632_0,
    i_8_299_1645_0, i_8_299_1649_0, i_8_299_1667_0, i_8_299_1668_0,
    i_8_299_1677_0, i_8_299_1707_0, i_8_299_1722_0, i_8_299_1723_0,
    i_8_299_1724_0, i_8_299_1743_0, i_8_299_1763_0, i_8_299_1814_0,
    i_8_299_1815_0, i_8_299_1816_0, i_8_299_1825_0, i_8_299_1831_0,
    i_8_299_1894_0, i_8_299_1907_0, i_8_299_1919_0, i_8_299_1970_0,
    i_8_299_2003_0, i_8_299_2041_0, i_8_299_2047_0, i_8_299_2109_0,
    i_8_299_2121_0, i_8_299_2174_0, i_8_299_2177_0, i_8_299_2202_0,
    i_8_299_2203_0, i_8_299_2212_0, i_8_299_2215_0, i_8_299_2256_0,
    i_8_299_2257_0, i_8_299_2274_0, i_8_299_2298_0,
    o_8_299_0_0  );
  input  i_8_299_31_0, i_8_299_89_0, i_8_299_96_0, i_8_299_98_0,
    i_8_299_196_0, i_8_299_237_0, i_8_299_240_0, i_8_299_241_0,
    i_8_299_295_0, i_8_299_296_0, i_8_299_312_0, i_8_299_324_0,
    i_8_299_349_0, i_8_299_372_0, i_8_299_424_0, i_8_299_480_0,
    i_8_299_528_0, i_8_299_529_0, i_8_299_556_0, i_8_299_605_0,
    i_8_299_733_0, i_8_299_735_0, i_8_299_736_0, i_8_299_763_0,
    i_8_299_778_0, i_8_299_779_0, i_8_299_781_0, i_8_299_789_0,
    i_8_299_797_0, i_8_299_815_0, i_8_299_837_0, i_8_299_862_0,
    i_8_299_940_0, i_8_299_941_0, i_8_299_943_0, i_8_299_947_0,
    i_8_299_996_0, i_8_299_1005_0, i_8_299_1012_0, i_8_299_1015_0,
    i_8_299_1060_0, i_8_299_1114_0, i_8_299_1115_0, i_8_299_1127_0,
    i_8_299_1130_0, i_8_299_1195_0, i_8_299_1219_0, i_8_299_1223_0,
    i_8_299_1292_0, i_8_299_1294_0, i_8_299_1306_0, i_8_299_1307_0,
    i_8_299_1310_0, i_8_299_1311_0, i_8_299_1314_0, i_8_299_1336_0,
    i_8_299_1410_0, i_8_299_1438_0, i_8_299_1472_0, i_8_299_1537_0,
    i_8_299_1538_0, i_8_299_1544_0, i_8_299_1597_0, i_8_299_1609_0,
    i_8_299_1632_0, i_8_299_1645_0, i_8_299_1649_0, i_8_299_1667_0,
    i_8_299_1668_0, i_8_299_1677_0, i_8_299_1707_0, i_8_299_1722_0,
    i_8_299_1723_0, i_8_299_1724_0, i_8_299_1743_0, i_8_299_1763_0,
    i_8_299_1814_0, i_8_299_1815_0, i_8_299_1816_0, i_8_299_1825_0,
    i_8_299_1831_0, i_8_299_1894_0, i_8_299_1907_0, i_8_299_1919_0,
    i_8_299_1970_0, i_8_299_2003_0, i_8_299_2041_0, i_8_299_2047_0,
    i_8_299_2109_0, i_8_299_2121_0, i_8_299_2174_0, i_8_299_2177_0,
    i_8_299_2202_0, i_8_299_2203_0, i_8_299_2212_0, i_8_299_2215_0,
    i_8_299_2256_0, i_8_299_2257_0, i_8_299_2274_0, i_8_299_2298_0;
  output o_8_299_0_0;
  assign o_8_299_0_0 = 0;
endmodule



// Benchmark "kernel_8_300" written by ABC on Sun Jul 19 10:08:18 2020

module kernel_8_300 ( 
    i_8_300_22_0, i_8_300_23_0, i_8_300_53_0, i_8_300_115_0, i_8_300_121_0,
    i_8_300_142_0, i_8_300_143_0, i_8_300_188_0, i_8_300_212_0,
    i_8_300_229_0, i_8_300_304_0, i_8_300_382_0, i_8_300_383_0,
    i_8_300_384_0, i_8_300_385_0, i_8_300_386_0, i_8_300_419_0,
    i_8_300_421_0, i_8_300_422_0, i_8_300_464_0, i_8_300_484_0,
    i_8_300_485_0, i_8_300_556_0, i_8_300_572_0, i_8_300_575_0,
    i_8_300_591_0, i_8_300_598_0, i_8_300_599_0, i_8_300_637_0,
    i_8_300_673_0, i_8_300_695_0, i_8_300_832_0, i_8_300_841_0,
    i_8_300_854_0, i_8_300_880_0, i_8_300_896_0, i_8_300_966_0,
    i_8_300_968_0, i_8_300_995_0, i_8_300_1015_0, i_8_300_1039_0,
    i_8_300_1040_0, i_8_300_1132_0, i_8_300_1225_0, i_8_300_1228_0,
    i_8_300_1232_0, i_8_300_1233_0, i_8_300_1255_0, i_8_300_1258_0,
    i_8_300_1259_0, i_8_300_1273_0, i_8_300_1277_0, i_8_300_1283_0,
    i_8_300_1284_0, i_8_300_1427_0, i_8_300_1438_0, i_8_300_1472_0,
    i_8_300_1474_0, i_8_300_1475_0, i_8_300_1481_0, i_8_300_1484_0,
    i_8_300_1490_0, i_8_300_1525_0, i_8_300_1526_0, i_8_300_1528_0,
    i_8_300_1529_0, i_8_300_1553_0, i_8_300_1556_0, i_8_300_1621_0,
    i_8_300_1643_0, i_8_300_1649_0, i_8_300_1655_0, i_8_300_1688_0,
    i_8_300_1696_0, i_8_300_1697_0, i_8_300_1723_0, i_8_300_1726_0,
    i_8_300_1727_0, i_8_300_1752_0, i_8_300_1771_0, i_8_300_1776_0,
    i_8_300_1795_0, i_8_300_1904_0, i_8_300_1944_0, i_8_300_1966_0,
    i_8_300_1973_0, i_8_300_2014_0, i_8_300_2038_0, i_8_300_2050_0,
    i_8_300_2093_0, i_8_300_2137_0, i_8_300_2150_0, i_8_300_2153_0,
    i_8_300_2155_0, i_8_300_2156_0, i_8_300_2158_0, i_8_300_2203_0,
    i_8_300_2233_0, i_8_300_2272_0, i_8_300_2275_0,
    o_8_300_0_0  );
  input  i_8_300_22_0, i_8_300_23_0, i_8_300_53_0, i_8_300_115_0,
    i_8_300_121_0, i_8_300_142_0, i_8_300_143_0, i_8_300_188_0,
    i_8_300_212_0, i_8_300_229_0, i_8_300_304_0, i_8_300_382_0,
    i_8_300_383_0, i_8_300_384_0, i_8_300_385_0, i_8_300_386_0,
    i_8_300_419_0, i_8_300_421_0, i_8_300_422_0, i_8_300_464_0,
    i_8_300_484_0, i_8_300_485_0, i_8_300_556_0, i_8_300_572_0,
    i_8_300_575_0, i_8_300_591_0, i_8_300_598_0, i_8_300_599_0,
    i_8_300_637_0, i_8_300_673_0, i_8_300_695_0, i_8_300_832_0,
    i_8_300_841_0, i_8_300_854_0, i_8_300_880_0, i_8_300_896_0,
    i_8_300_966_0, i_8_300_968_0, i_8_300_995_0, i_8_300_1015_0,
    i_8_300_1039_0, i_8_300_1040_0, i_8_300_1132_0, i_8_300_1225_0,
    i_8_300_1228_0, i_8_300_1232_0, i_8_300_1233_0, i_8_300_1255_0,
    i_8_300_1258_0, i_8_300_1259_0, i_8_300_1273_0, i_8_300_1277_0,
    i_8_300_1283_0, i_8_300_1284_0, i_8_300_1427_0, i_8_300_1438_0,
    i_8_300_1472_0, i_8_300_1474_0, i_8_300_1475_0, i_8_300_1481_0,
    i_8_300_1484_0, i_8_300_1490_0, i_8_300_1525_0, i_8_300_1526_0,
    i_8_300_1528_0, i_8_300_1529_0, i_8_300_1553_0, i_8_300_1556_0,
    i_8_300_1621_0, i_8_300_1643_0, i_8_300_1649_0, i_8_300_1655_0,
    i_8_300_1688_0, i_8_300_1696_0, i_8_300_1697_0, i_8_300_1723_0,
    i_8_300_1726_0, i_8_300_1727_0, i_8_300_1752_0, i_8_300_1771_0,
    i_8_300_1776_0, i_8_300_1795_0, i_8_300_1904_0, i_8_300_1944_0,
    i_8_300_1966_0, i_8_300_1973_0, i_8_300_2014_0, i_8_300_2038_0,
    i_8_300_2050_0, i_8_300_2093_0, i_8_300_2137_0, i_8_300_2150_0,
    i_8_300_2153_0, i_8_300_2155_0, i_8_300_2156_0, i_8_300_2158_0,
    i_8_300_2203_0, i_8_300_2233_0, i_8_300_2272_0, i_8_300_2275_0;
  output o_8_300_0_0;
  assign o_8_300_0_0 = ~((~i_8_300_1529_0 & ((~i_8_300_115_0 & ((~i_8_300_142_0 & ~i_8_300_896_0 & ~i_8_300_1481_0 & i_8_300_1484_0 & ~i_8_300_1795_0 & ~i_8_300_1966_0) | (~i_8_300_968_0 & i_8_300_995_0 & ~i_8_300_1015_0 & i_8_300_1472_0 & ~i_8_300_1649_0 & ~i_8_300_1726_0 & ~i_8_300_2156_0))) | (~i_8_300_2050_0 & ((~i_8_300_832_0 & ((~i_8_300_22_0 & ~i_8_300_53_0 & ~i_8_300_384_0 & i_8_300_966_0 & i_8_300_968_0 & ~i_8_300_1490_0 & ~i_8_300_1525_0 & ~i_8_300_1526_0 & ~i_8_300_1966_0 & ~i_8_300_2014_0) | (~i_8_300_421_0 & ~i_8_300_556_0 & ~i_8_300_896_0 & ~i_8_300_1039_0 & ~i_8_300_1427_0 & ~i_8_300_1481_0 & ~i_8_300_1697_0 & ~i_8_300_1727_0 & ~i_8_300_2150_0 & ~i_8_300_2203_0))) | (~i_8_300_143_0 & i_8_300_382_0 & ~i_8_300_995_0 & ~i_8_300_1475_0 & ~i_8_300_1481_0) | (~i_8_300_419_0 & ~i_8_300_422_0 & ~i_8_300_485_0 & ~i_8_300_575_0 & ~i_8_300_1040_0 & ~i_8_300_1132_0 & ~i_8_300_1490_0 & ~i_8_300_1696_0))) | (~i_8_300_1697_0 & ((~i_8_300_575_0 & ((~i_8_300_896_0 & ~i_8_300_995_0 & ~i_8_300_1277_0 & i_8_300_1284_0 & ~i_8_300_1475_0 & ~i_8_300_1525_0 & ~i_8_300_1688_0) | (~i_8_300_229_0 & ~i_8_300_572_0 & i_8_300_1283_0 & ~i_8_300_1481_0 & ~i_8_300_1526_0 & ~i_8_300_1771_0))) | (~i_8_300_484_0 & ~i_8_300_1132_0 & ~i_8_300_1490_0 & ~i_8_300_1525_0 & ~i_8_300_1526_0 & ~i_8_300_1649_0 & ~i_8_300_1655_0 & ~i_8_300_1726_0 & ~i_8_300_1727_0 & ~i_8_300_1904_0))) | (i_8_300_1277_0 & ~i_8_300_1438_0 & i_8_300_1475_0 & ~i_8_300_1481_0 & i_8_300_1966_0) | (~i_8_300_142_0 & ~i_8_300_995_0 & ~i_8_300_1015_0 & ~i_8_300_1225_0 & ~i_8_300_1273_0 & ~i_8_300_1427_0 & ~i_8_300_1526_0 & ~i_8_300_1723_0 & ~i_8_300_1726_0 & ~i_8_300_1795_0 & ~i_8_300_2093_0 & ~i_8_300_2153_0))) | (~i_8_300_53_0 & ~i_8_300_556_0 & ((~i_8_300_464_0 & ~i_8_300_484_0 & ~i_8_300_485_0 & ~i_8_300_575_0 & ~i_8_300_832_0 & ~i_8_300_968_0 & ~i_8_300_1039_0 & ~i_8_300_1040_0 & ~i_8_300_1688_0 & ~i_8_300_2150_0) | (i_8_300_386_0 & ~i_8_300_1427_0 & ~i_8_300_1474_0 & ~i_8_300_1655_0 & ~i_8_300_1696_0 & ~i_8_300_2203_0))) | (~i_8_300_143_0 & ((~i_8_300_142_0 & ~i_8_300_575_0 & ~i_8_300_880_0 & ~i_8_300_1427_0 & i_8_300_1472_0 & ~i_8_300_1697_0 & ~i_8_300_1723_0 & ~i_8_300_1727_0) | (~i_8_300_572_0 & ~i_8_300_841_0 & ~i_8_300_896_0 & ~i_8_300_966_0 & ~i_8_300_995_0 & ~i_8_300_1132_0 & ~i_8_300_1277_0 & ~i_8_300_1553_0 & ~i_8_300_1655_0 & ~i_8_300_1795_0 & ~i_8_300_2150_0))) | (~i_8_300_1528_0 & ((~i_8_300_188_0 & ~i_8_300_1427_0 & ((~i_8_300_419_0 & ~i_8_300_485_0 & ~i_8_300_896_0 & ~i_8_300_1233_0 & ~i_8_300_1526_0 & ~i_8_300_1621_0 & ~i_8_300_1643_0 & ~i_8_300_1723_0 & ~i_8_300_1776_0 & i_8_300_1966_0) | (~i_8_300_422_0 & ~i_8_300_464_0 & ~i_8_300_575_0 & i_8_300_598_0 & ~i_8_300_1015_0 & ~i_8_300_2014_0 & ~i_8_300_2153_0))) | (~i_8_300_575_0 & ((~i_8_300_422_0 & ~i_8_300_995_0 & i_8_300_1277_0 & ~i_8_300_1723_0) | (i_8_300_53_0 & ~i_8_300_419_0 & i_8_300_880_0 & ~i_8_300_1688_0 & ~i_8_300_2153_0))) | (~i_8_300_1039_0 & ~i_8_300_1526_0 & ~i_8_300_1621_0 & ~i_8_300_1727_0 & ~i_8_300_1904_0 & i_8_300_2155_0 & ~i_8_300_2275_0))) | (~i_8_300_421_0 & ((~i_8_300_1525_0 & ~i_8_300_1526_0 & ~i_8_300_422_0 & i_8_300_599_0 & ~i_8_300_1621_0 & ~i_8_300_1697_0 & ~i_8_300_1795_0 & ~i_8_300_2050_0) | (~i_8_300_229_0 & ~i_8_300_484_0 & ~i_8_300_575_0 & i_8_300_841_0 & ~i_8_300_896_0 & i_8_300_968_0 & ~i_8_300_995_0 & ~i_8_300_1727_0 & ~i_8_300_2272_0))) | (~i_8_300_1427_0 & ((~i_8_300_575_0 & ((~i_8_300_422_0 & ((~i_8_300_142_0 & ~i_8_300_896_0 & ~i_8_300_968_0 & ~i_8_300_1472_0 & i_8_300_1556_0 & ~i_8_300_1723_0 & ~i_8_300_1771_0) | (~i_8_300_121_0 & ~i_8_300_832_0 & ~i_8_300_1277_0 & ~i_8_300_1526_0 & ~i_8_300_1697_0 & ~i_8_300_1727_0 & ~i_8_300_1795_0 & i_8_300_1966_0))) | (~i_8_300_572_0 & ~i_8_300_695_0 & i_8_300_1273_0 & ~i_8_300_1525_0 & ~i_8_300_1655_0 & ~i_8_300_1771_0 & ~i_8_300_2014_0 & ~i_8_300_2203_0))) | (~i_8_300_121_0 & ~i_8_300_1040_0 & ((~i_8_300_485_0 & ~i_8_300_572_0 & ~i_8_300_1015_0 & ~i_8_300_1553_0 & ~i_8_300_1649_0 & ~i_8_300_1688_0 & ~i_8_300_1726_0 & ~i_8_300_2050_0) | (i_8_300_422_0 & i_8_300_599_0 & ~i_8_300_1284_0 & ~i_8_300_1752_0 & ~i_8_300_1904_0 & i_8_300_2093_0))) | (~i_8_300_142_0 & ~i_8_300_1526_0 & ((i_8_300_591_0 & ~i_8_300_854_0 & ~i_8_300_995_0 & ~i_8_300_1039_0 & ~i_8_300_1727_0) | (~i_8_300_896_0 & ~i_8_300_1273_0 & ~i_8_300_1643_0 & ~i_8_300_1752_0 & i_8_300_1776_0 & ~i_8_300_1904_0 & ~i_8_300_2014_0 & ~i_8_300_2050_0))))) | (~i_8_300_1726_0 & ((~i_8_300_121_0 & ((~i_8_300_142_0 & ~i_8_300_572_0 & ~i_8_300_968_0 & ~i_8_300_1228_0 & ~i_8_300_1484_0 & ~i_8_300_1655_0 & ~i_8_300_1697_0 & ~i_8_300_2050_0 & ~i_8_300_2137_0 & ~i_8_300_2150_0 & ~i_8_300_2155_0) | (~i_8_300_484_0 & ~i_8_300_485_0 & ~i_8_300_575_0 & ~i_8_300_1040_0 & ~i_8_300_1526_0 & ~i_8_300_1688_0 & ~i_8_300_1944_0 & ~i_8_300_2272_0 & ~i_8_300_2275_0))) | (~i_8_300_188_0 & ~i_8_300_212_0 & ~i_8_300_484_0 & ~i_8_300_995_0 & ~i_8_300_1525_0 & ~i_8_300_1688_0 & i_8_300_2275_0))) | (~i_8_300_1727_0 & ((~i_8_300_572_0 & ((i_8_300_464_0 & ~i_8_300_575_0 & ~i_8_300_896_0 & ~i_8_300_966_0 & ~i_8_300_1039_0 & ~i_8_300_1132_0 & ~i_8_300_1283_0 & ~i_8_300_1438_0 & ~i_8_300_1771_0 & ~i_8_300_2050_0 & i_8_300_2093_0) | (~i_8_300_1525_0 & ~i_8_300_1556_0 & ~i_8_300_1966_0 & i_8_300_2203_0))) | (i_8_300_1273_0 & ~i_8_300_1484_0 & ~i_8_300_1723_0 & i_8_300_2155_0))) | (i_8_300_382_0 & i_8_300_383_0 & ~i_8_300_995_0 & i_8_300_1277_0 & ~i_8_300_1655_0) | (i_8_300_695_0 & i_8_300_1225_0 & i_8_300_1649_0 & ~i_8_300_1697_0));
endmodule



// Benchmark "kernel_8_301" written by ABC on Sun Jul 19 10:08:19 2020

module kernel_8_301 ( 
    i_8_301_40_0, i_8_301_41_0, i_8_301_43_0, i_8_301_44_0, i_8_301_97_0,
    i_8_301_118_0, i_8_301_170_0, i_8_301_178_0, i_8_301_239_0,
    i_8_301_242_0, i_8_301_256_0, i_8_301_259_0, i_8_301_260_0,
    i_8_301_269_0, i_8_301_301_0, i_8_301_304_0, i_8_301_305_0,
    i_8_301_347_0, i_8_301_363_0, i_8_301_377_0, i_8_301_380_0,
    i_8_301_401_0, i_8_301_430_0, i_8_301_453_0, i_8_301_454_0,
    i_8_301_456_0, i_8_301_494_0, i_8_301_528_0, i_8_301_584_0,
    i_8_301_634_0, i_8_301_638_0, i_8_301_647_0, i_8_301_662_0,
    i_8_301_679_0, i_8_301_680_0, i_8_301_692_0, i_8_301_698_0,
    i_8_301_709_0, i_8_301_796_0, i_8_301_842_0, i_8_301_855_0,
    i_8_301_886_0, i_8_301_955_0, i_8_301_1060_0, i_8_301_1080_0,
    i_8_301_1125_0, i_8_301_1192_0, i_8_301_1228_0, i_8_301_1237_0,
    i_8_301_1261_0, i_8_301_1274_0, i_8_301_1282_0, i_8_301_1285_0,
    i_8_301_1295_0, i_8_301_1308_0, i_8_301_1310_0, i_8_301_1336_0,
    i_8_301_1352_0, i_8_301_1354_0, i_8_301_1373_0, i_8_301_1411_0,
    i_8_301_1416_0, i_8_301_1419_0, i_8_301_1456_0, i_8_301_1457_0,
    i_8_301_1610_0, i_8_301_1615_0, i_8_301_1642_0, i_8_301_1645_0,
    i_8_301_1673_0, i_8_301_1690_0, i_8_301_1691_0, i_8_301_1703_0,
    i_8_301_1787_0, i_8_301_1855_0, i_8_301_1857_0, i_8_301_1859_0,
    i_8_301_1886_0, i_8_301_1922_0, i_8_301_1940_0, i_8_301_1970_0,
    i_8_301_1982_0, i_8_301_1989_0, i_8_301_1993_0, i_8_301_2003_0,
    i_8_301_2005_0, i_8_301_2006_0, i_8_301_2056_0, i_8_301_2113_0,
    i_8_301_2114_0, i_8_301_2154_0, i_8_301_2156_0, i_8_301_2159_0,
    i_8_301_2201_0, i_8_301_2213_0, i_8_301_2223_0, i_8_301_2257_0,
    i_8_301_2261_0, i_8_301_2284_0, i_8_301_2285_0,
    o_8_301_0_0  );
  input  i_8_301_40_0, i_8_301_41_0, i_8_301_43_0, i_8_301_44_0,
    i_8_301_97_0, i_8_301_118_0, i_8_301_170_0, i_8_301_178_0,
    i_8_301_239_0, i_8_301_242_0, i_8_301_256_0, i_8_301_259_0,
    i_8_301_260_0, i_8_301_269_0, i_8_301_301_0, i_8_301_304_0,
    i_8_301_305_0, i_8_301_347_0, i_8_301_363_0, i_8_301_377_0,
    i_8_301_380_0, i_8_301_401_0, i_8_301_430_0, i_8_301_453_0,
    i_8_301_454_0, i_8_301_456_0, i_8_301_494_0, i_8_301_528_0,
    i_8_301_584_0, i_8_301_634_0, i_8_301_638_0, i_8_301_647_0,
    i_8_301_662_0, i_8_301_679_0, i_8_301_680_0, i_8_301_692_0,
    i_8_301_698_0, i_8_301_709_0, i_8_301_796_0, i_8_301_842_0,
    i_8_301_855_0, i_8_301_886_0, i_8_301_955_0, i_8_301_1060_0,
    i_8_301_1080_0, i_8_301_1125_0, i_8_301_1192_0, i_8_301_1228_0,
    i_8_301_1237_0, i_8_301_1261_0, i_8_301_1274_0, i_8_301_1282_0,
    i_8_301_1285_0, i_8_301_1295_0, i_8_301_1308_0, i_8_301_1310_0,
    i_8_301_1336_0, i_8_301_1352_0, i_8_301_1354_0, i_8_301_1373_0,
    i_8_301_1411_0, i_8_301_1416_0, i_8_301_1419_0, i_8_301_1456_0,
    i_8_301_1457_0, i_8_301_1610_0, i_8_301_1615_0, i_8_301_1642_0,
    i_8_301_1645_0, i_8_301_1673_0, i_8_301_1690_0, i_8_301_1691_0,
    i_8_301_1703_0, i_8_301_1787_0, i_8_301_1855_0, i_8_301_1857_0,
    i_8_301_1859_0, i_8_301_1886_0, i_8_301_1922_0, i_8_301_1940_0,
    i_8_301_1970_0, i_8_301_1982_0, i_8_301_1989_0, i_8_301_1993_0,
    i_8_301_2003_0, i_8_301_2005_0, i_8_301_2006_0, i_8_301_2056_0,
    i_8_301_2113_0, i_8_301_2114_0, i_8_301_2154_0, i_8_301_2156_0,
    i_8_301_2159_0, i_8_301_2201_0, i_8_301_2213_0, i_8_301_2223_0,
    i_8_301_2257_0, i_8_301_2261_0, i_8_301_2284_0, i_8_301_2285_0;
  output o_8_301_0_0;
  assign o_8_301_0_0 = 0;
endmodule



// Benchmark "kernel_8_302" written by ABC on Sun Jul 19 10:08:20 2020

module kernel_8_302 ( 
    i_8_302_28_0, i_8_302_40_0, i_8_302_227_0, i_8_302_259_0,
    i_8_302_275_0, i_8_302_318_0, i_8_302_335_0, i_8_302_348_0,
    i_8_302_390_0, i_8_302_398_0, i_8_302_401_0, i_8_302_418_0,
    i_8_302_422_0, i_8_302_427_0, i_8_302_451_0, i_8_302_506_0,
    i_8_302_508_0, i_8_302_509_0, i_8_302_552_0, i_8_302_553_0,
    i_8_302_554_0, i_8_302_572_0, i_8_302_603_0, i_8_302_604_0,
    i_8_302_631_0, i_8_302_638_0, i_8_302_651_0, i_8_302_705_0,
    i_8_302_707_0, i_8_302_710_0, i_8_302_749_0, i_8_302_884_0,
    i_8_302_895_0, i_8_302_896_0, i_8_302_1011_0, i_8_302_1040_0,
    i_8_302_1052_0, i_8_302_1058_0, i_8_302_1103_0, i_8_302_1106_0,
    i_8_302_1107_0, i_8_302_1112_0, i_8_302_1138_0, i_8_302_1139_0,
    i_8_302_1154_0, i_8_302_1180_0, i_8_302_1202_0, i_8_302_1235_0,
    i_8_302_1238_0, i_8_302_1244_0, i_8_302_1279_0, i_8_302_1305_0,
    i_8_302_1319_0, i_8_302_1362_0, i_8_302_1364_0, i_8_302_1422_0,
    i_8_302_1427_0, i_8_302_1429_0, i_8_302_1436_0, i_8_302_1458_0,
    i_8_302_1461_0, i_8_302_1462_0, i_8_302_1463_0, i_8_302_1471_0,
    i_8_302_1479_0, i_8_302_1480_0, i_8_302_1487_0, i_8_302_1508_0,
    i_8_302_1511_0, i_8_302_1512_0, i_8_302_1515_0, i_8_302_1524_0,
    i_8_302_1551_0, i_8_302_1569_0, i_8_302_1678_0, i_8_302_1702_0,
    i_8_302_1705_0, i_8_302_1706_0, i_8_302_1774_0, i_8_302_1776_0,
    i_8_302_1784_0, i_8_302_1795_0, i_8_302_1836_0, i_8_302_1839_0,
    i_8_302_1841_0, i_8_302_1892_0, i_8_302_1919_0, i_8_302_1955_0,
    i_8_302_1974_0, i_8_302_1997_0, i_8_302_2057_0, i_8_302_2075_0,
    i_8_302_2151_0, i_8_302_2155_0, i_8_302_2223_0, i_8_302_2224_0,
    i_8_302_2225_0, i_8_302_2245_0, i_8_302_2248_0, i_8_302_2249_0,
    o_8_302_0_0  );
  input  i_8_302_28_0, i_8_302_40_0, i_8_302_227_0, i_8_302_259_0,
    i_8_302_275_0, i_8_302_318_0, i_8_302_335_0, i_8_302_348_0,
    i_8_302_390_0, i_8_302_398_0, i_8_302_401_0, i_8_302_418_0,
    i_8_302_422_0, i_8_302_427_0, i_8_302_451_0, i_8_302_506_0,
    i_8_302_508_0, i_8_302_509_0, i_8_302_552_0, i_8_302_553_0,
    i_8_302_554_0, i_8_302_572_0, i_8_302_603_0, i_8_302_604_0,
    i_8_302_631_0, i_8_302_638_0, i_8_302_651_0, i_8_302_705_0,
    i_8_302_707_0, i_8_302_710_0, i_8_302_749_0, i_8_302_884_0,
    i_8_302_895_0, i_8_302_896_0, i_8_302_1011_0, i_8_302_1040_0,
    i_8_302_1052_0, i_8_302_1058_0, i_8_302_1103_0, i_8_302_1106_0,
    i_8_302_1107_0, i_8_302_1112_0, i_8_302_1138_0, i_8_302_1139_0,
    i_8_302_1154_0, i_8_302_1180_0, i_8_302_1202_0, i_8_302_1235_0,
    i_8_302_1238_0, i_8_302_1244_0, i_8_302_1279_0, i_8_302_1305_0,
    i_8_302_1319_0, i_8_302_1362_0, i_8_302_1364_0, i_8_302_1422_0,
    i_8_302_1427_0, i_8_302_1429_0, i_8_302_1436_0, i_8_302_1458_0,
    i_8_302_1461_0, i_8_302_1462_0, i_8_302_1463_0, i_8_302_1471_0,
    i_8_302_1479_0, i_8_302_1480_0, i_8_302_1487_0, i_8_302_1508_0,
    i_8_302_1511_0, i_8_302_1512_0, i_8_302_1515_0, i_8_302_1524_0,
    i_8_302_1551_0, i_8_302_1569_0, i_8_302_1678_0, i_8_302_1702_0,
    i_8_302_1705_0, i_8_302_1706_0, i_8_302_1774_0, i_8_302_1776_0,
    i_8_302_1784_0, i_8_302_1795_0, i_8_302_1836_0, i_8_302_1839_0,
    i_8_302_1841_0, i_8_302_1892_0, i_8_302_1919_0, i_8_302_1955_0,
    i_8_302_1974_0, i_8_302_1997_0, i_8_302_2057_0, i_8_302_2075_0,
    i_8_302_2151_0, i_8_302_2155_0, i_8_302_2223_0, i_8_302_2224_0,
    i_8_302_2225_0, i_8_302_2245_0, i_8_302_2248_0, i_8_302_2249_0;
  output o_8_302_0_0;
  assign o_8_302_0_0 = 0;
endmodule



// Benchmark "kernel_8_303" written by ABC on Sun Jul 19 10:08:21 2020

module kernel_8_303 ( 
    i_8_303_20_0, i_8_303_107_0, i_8_303_240_0, i_8_303_255_0,
    i_8_303_324_0, i_8_303_325_0, i_8_303_328_0, i_8_303_345_0,
    i_8_303_348_0, i_8_303_380_0, i_8_303_382_0, i_8_303_391_0,
    i_8_303_440_0, i_8_303_460_0, i_8_303_469_0, i_8_303_474_0,
    i_8_303_478_0, i_8_303_483_0, i_8_303_507_0, i_8_303_523_0,
    i_8_303_524_0, i_8_303_527_0, i_8_303_549_0, i_8_303_551_0,
    i_8_303_552_0, i_8_303_599_0, i_8_303_604_0, i_8_303_637_0,
    i_8_303_712_0, i_8_303_715_0, i_8_303_732_0, i_8_303_757_0,
    i_8_303_763_0, i_8_303_778_0, i_8_303_800_0, i_8_303_943_0,
    i_8_303_945_0, i_8_303_946_0, i_8_303_947_0, i_8_303_990_0,
    i_8_303_997_0, i_8_303_1050_0, i_8_303_1072_0, i_8_303_1075_0,
    i_8_303_1110_0, i_8_303_1114_0, i_8_303_1117_0, i_8_303_1130_0,
    i_8_303_1169_0, i_8_303_1176_0, i_8_303_1190_0, i_8_303_1238_0,
    i_8_303_1257_0, i_8_303_1273_0, i_8_303_1284_0, i_8_303_1315_0,
    i_8_303_1323_0, i_8_303_1324_0, i_8_303_1326_0, i_8_303_1347_0,
    i_8_303_1387_0, i_8_303_1417_0, i_8_303_1438_0, i_8_303_1441_0,
    i_8_303_1452_0, i_8_303_1506_0, i_8_303_1530_0, i_8_303_1534_0,
    i_8_303_1562_0, i_8_303_1649_0, i_8_303_1671_0, i_8_303_1681_0,
    i_8_303_1716_0, i_8_303_1722_0, i_8_303_1723_0, i_8_303_1726_0,
    i_8_303_1732_0, i_8_303_1746_0, i_8_303_1833_0, i_8_303_1841_0,
    i_8_303_1854_0, i_8_303_1864_0, i_8_303_1887_0, i_8_303_1894_0,
    i_8_303_1949_0, i_8_303_1965_0, i_8_303_1992_0, i_8_303_2002_0,
    i_8_303_2028_0, i_8_303_2031_0, i_8_303_2032_0, i_8_303_2051_0,
    i_8_303_2064_0, i_8_303_2092_0, i_8_303_2115_0, i_8_303_2175_0,
    i_8_303_2215_0, i_8_303_2216_0, i_8_303_2219_0, i_8_303_2283_0,
    o_8_303_0_0  );
  input  i_8_303_20_0, i_8_303_107_0, i_8_303_240_0, i_8_303_255_0,
    i_8_303_324_0, i_8_303_325_0, i_8_303_328_0, i_8_303_345_0,
    i_8_303_348_0, i_8_303_380_0, i_8_303_382_0, i_8_303_391_0,
    i_8_303_440_0, i_8_303_460_0, i_8_303_469_0, i_8_303_474_0,
    i_8_303_478_0, i_8_303_483_0, i_8_303_507_0, i_8_303_523_0,
    i_8_303_524_0, i_8_303_527_0, i_8_303_549_0, i_8_303_551_0,
    i_8_303_552_0, i_8_303_599_0, i_8_303_604_0, i_8_303_637_0,
    i_8_303_712_0, i_8_303_715_0, i_8_303_732_0, i_8_303_757_0,
    i_8_303_763_0, i_8_303_778_0, i_8_303_800_0, i_8_303_943_0,
    i_8_303_945_0, i_8_303_946_0, i_8_303_947_0, i_8_303_990_0,
    i_8_303_997_0, i_8_303_1050_0, i_8_303_1072_0, i_8_303_1075_0,
    i_8_303_1110_0, i_8_303_1114_0, i_8_303_1117_0, i_8_303_1130_0,
    i_8_303_1169_0, i_8_303_1176_0, i_8_303_1190_0, i_8_303_1238_0,
    i_8_303_1257_0, i_8_303_1273_0, i_8_303_1284_0, i_8_303_1315_0,
    i_8_303_1323_0, i_8_303_1324_0, i_8_303_1326_0, i_8_303_1347_0,
    i_8_303_1387_0, i_8_303_1417_0, i_8_303_1438_0, i_8_303_1441_0,
    i_8_303_1452_0, i_8_303_1506_0, i_8_303_1530_0, i_8_303_1534_0,
    i_8_303_1562_0, i_8_303_1649_0, i_8_303_1671_0, i_8_303_1681_0,
    i_8_303_1716_0, i_8_303_1722_0, i_8_303_1723_0, i_8_303_1726_0,
    i_8_303_1732_0, i_8_303_1746_0, i_8_303_1833_0, i_8_303_1841_0,
    i_8_303_1854_0, i_8_303_1864_0, i_8_303_1887_0, i_8_303_1894_0,
    i_8_303_1949_0, i_8_303_1965_0, i_8_303_1992_0, i_8_303_2002_0,
    i_8_303_2028_0, i_8_303_2031_0, i_8_303_2032_0, i_8_303_2051_0,
    i_8_303_2064_0, i_8_303_2092_0, i_8_303_2115_0, i_8_303_2175_0,
    i_8_303_2215_0, i_8_303_2216_0, i_8_303_2219_0, i_8_303_2283_0;
  output o_8_303_0_0;
  assign o_8_303_0_0 = 0;
endmodule



// Benchmark "kernel_8_304" written by ABC on Sun Jul 19 10:08:23 2020

module kernel_8_304 ( 
    i_8_304_19_0, i_8_304_39_0, i_8_304_87_0, i_8_304_111_0, i_8_304_112_0,
    i_8_304_113_0, i_8_304_219_0, i_8_304_245_0, i_8_304_266_0,
    i_8_304_269_0, i_8_304_286_0, i_8_304_287_0, i_8_304_295_0,
    i_8_304_296_0, i_8_304_304_0, i_8_304_305_0, i_8_304_381_0,
    i_8_304_383_0, i_8_304_427_0, i_8_304_428_0, i_8_304_429_0,
    i_8_304_430_0, i_8_304_431_0, i_8_304_504_0, i_8_304_524_0,
    i_8_304_567_0, i_8_304_568_0, i_8_304_569_0, i_8_304_577_0,
    i_8_304_578_0, i_8_304_606_0, i_8_304_607_0, i_8_304_635_0,
    i_8_304_705_0, i_8_304_708_0, i_8_304_709_0, i_8_304_710_0,
    i_8_304_713_0, i_8_304_715_0, i_8_304_726_0, i_8_304_816_0,
    i_8_304_817_0, i_8_304_838_0, i_8_304_846_0, i_8_304_847_0,
    i_8_304_878_0, i_8_304_1078_0, i_8_304_1179_0, i_8_304_1180_0,
    i_8_304_1181_0, i_8_304_1189_0, i_8_304_1266_0, i_8_304_1315_0,
    i_8_304_1329_0, i_8_304_1359_0, i_8_304_1365_0, i_8_304_1394_0,
    i_8_304_1399_0, i_8_304_1467_0, i_8_304_1468_0, i_8_304_1469_0,
    i_8_304_1470_0, i_8_304_1472_0, i_8_304_1522_0, i_8_304_1534_0,
    i_8_304_1565_0, i_8_304_1621_0, i_8_304_1683_0, i_8_304_1684_0,
    i_8_304_1693_0, i_8_304_1694_0, i_8_304_1730_0, i_8_304_1747_0,
    i_8_304_1749_0, i_8_304_1765_0, i_8_304_1777_0, i_8_304_1780_0,
    i_8_304_1784_0, i_8_304_1785_0, i_8_304_1786_0, i_8_304_1787_0,
    i_8_304_1825_0, i_8_304_1826_0, i_8_304_1854_0, i_8_304_1873_0,
    i_8_304_1874_0, i_8_304_1889_0, i_8_304_1920_0, i_8_304_1946_0,
    i_8_304_2060_0, i_8_304_2070_0, i_8_304_2071_0, i_8_304_2088_0,
    i_8_304_2138_0, i_8_304_2139_0, i_8_304_2226_0, i_8_304_2227_0,
    i_8_304_2233_0, i_8_304_2243_0, i_8_304_2274_0,
    o_8_304_0_0  );
  input  i_8_304_19_0, i_8_304_39_0, i_8_304_87_0, i_8_304_111_0,
    i_8_304_112_0, i_8_304_113_0, i_8_304_219_0, i_8_304_245_0,
    i_8_304_266_0, i_8_304_269_0, i_8_304_286_0, i_8_304_287_0,
    i_8_304_295_0, i_8_304_296_0, i_8_304_304_0, i_8_304_305_0,
    i_8_304_381_0, i_8_304_383_0, i_8_304_427_0, i_8_304_428_0,
    i_8_304_429_0, i_8_304_430_0, i_8_304_431_0, i_8_304_504_0,
    i_8_304_524_0, i_8_304_567_0, i_8_304_568_0, i_8_304_569_0,
    i_8_304_577_0, i_8_304_578_0, i_8_304_606_0, i_8_304_607_0,
    i_8_304_635_0, i_8_304_705_0, i_8_304_708_0, i_8_304_709_0,
    i_8_304_710_0, i_8_304_713_0, i_8_304_715_0, i_8_304_726_0,
    i_8_304_816_0, i_8_304_817_0, i_8_304_838_0, i_8_304_846_0,
    i_8_304_847_0, i_8_304_878_0, i_8_304_1078_0, i_8_304_1179_0,
    i_8_304_1180_0, i_8_304_1181_0, i_8_304_1189_0, i_8_304_1266_0,
    i_8_304_1315_0, i_8_304_1329_0, i_8_304_1359_0, i_8_304_1365_0,
    i_8_304_1394_0, i_8_304_1399_0, i_8_304_1467_0, i_8_304_1468_0,
    i_8_304_1469_0, i_8_304_1470_0, i_8_304_1472_0, i_8_304_1522_0,
    i_8_304_1534_0, i_8_304_1565_0, i_8_304_1621_0, i_8_304_1683_0,
    i_8_304_1684_0, i_8_304_1693_0, i_8_304_1694_0, i_8_304_1730_0,
    i_8_304_1747_0, i_8_304_1749_0, i_8_304_1765_0, i_8_304_1777_0,
    i_8_304_1780_0, i_8_304_1784_0, i_8_304_1785_0, i_8_304_1786_0,
    i_8_304_1787_0, i_8_304_1825_0, i_8_304_1826_0, i_8_304_1854_0,
    i_8_304_1873_0, i_8_304_1874_0, i_8_304_1889_0, i_8_304_1920_0,
    i_8_304_1946_0, i_8_304_2060_0, i_8_304_2070_0, i_8_304_2071_0,
    i_8_304_2088_0, i_8_304_2138_0, i_8_304_2139_0, i_8_304_2226_0,
    i_8_304_2227_0, i_8_304_2233_0, i_8_304_2243_0, i_8_304_2274_0;
  output o_8_304_0_0;
  assign o_8_304_0_0 = ~((i_8_304_39_0 & ((i_8_304_606_0 & ~i_8_304_1467_0 & i_8_304_1747_0 & ~i_8_304_1749_0) | (~i_8_304_567_0 & ~i_8_304_816_0 & ~i_8_304_1078_0 & ~i_8_304_1179_0 & ~i_8_304_1365_0 & ~i_8_304_1621_0 & ~i_8_304_1684_0 & i_8_304_2226_0))) | (~i_8_304_1181_0 & ((~i_8_304_569_0 & ((~i_8_304_1694_0 & ((~i_8_304_87_0 & ((~i_8_304_112_0 & ~i_8_304_245_0 & ~i_8_304_296_0 & ~i_8_304_567_0 & ~i_8_304_606_0 & i_8_304_607_0 & ~i_8_304_1394_0 & ~i_8_304_1467_0 & ~i_8_304_1621_0 & ~i_8_304_1730_0 & ~i_8_304_2060_0) | (~i_8_304_111_0 & ~i_8_304_304_0 & ~i_8_304_568_0 & ~i_8_304_635_0 & ~i_8_304_817_0 & ~i_8_304_1469_0 & ~i_8_304_1472_0 & i_8_304_1787_0 & ~i_8_304_2233_0 & ~i_8_304_2243_0))) | (~i_8_304_266_0 & ~i_8_304_428_0 & ~i_8_304_578_0 & ~i_8_304_1179_0 & i_8_304_1784_0 & ~i_8_304_1854_0 & ~i_8_304_2070_0))) | (~i_8_304_113_0 & ~i_8_304_568_0 & ~i_8_304_578_0 & i_8_304_606_0 & i_8_304_607_0 & ~i_8_304_816_0 & ~i_8_304_838_0 & ~i_8_304_1179_0 & ~i_8_304_1684_0 & ~i_8_304_1693_0 & ~i_8_304_1854_0 & ~i_8_304_2071_0))) | (~i_8_304_219_0 & ((~i_8_304_287_0 & ~i_8_304_304_0 & ~i_8_304_427_0 & ~i_8_304_708_0 & ~i_8_304_838_0 & ~i_8_304_878_0 & ~i_8_304_1394_0 & i_8_304_1826_0 & ~i_8_304_2139_0) | (~i_8_304_578_0 & ~i_8_304_1749_0 & i_8_304_1946_0 & i_8_304_2138_0 & ~i_8_304_2274_0))) | (~i_8_304_1854_0 & ((~i_8_304_113_0 & ~i_8_304_817_0 & ((~i_8_304_266_0 & ~i_8_304_296_0 & i_8_304_428_0 & ~i_8_304_577_0 & ~i_8_304_1078_0 & ~i_8_304_1189_0 & ~i_8_304_1469_0 & ~i_8_304_1621_0 & ~i_8_304_1730_0 & ~i_8_304_1786_0) | (~i_8_304_245_0 & ~i_8_304_305_0 & ~i_8_304_524_0 & ~i_8_304_705_0 & i_8_304_878_0 & ~i_8_304_1684_0 & ~i_8_304_1693_0 & ~i_8_304_1749_0 & ~i_8_304_2071_0 & ~i_8_304_2243_0))) | (i_8_304_428_0 & ~i_8_304_578_0 & i_8_304_1469_0 & ~i_8_304_1683_0 & ~i_8_304_1693_0 & ~i_8_304_1786_0) | (~i_8_304_266_0 & ~i_8_304_269_0 & ~i_8_304_295_0 & ~i_8_304_305_0 & i_8_304_383_0 & ~i_8_304_2071_0 & i_8_304_2138_0))) | (~i_8_304_1359_0 & ((~i_8_304_295_0 & ((~i_8_304_269_0 & i_8_304_305_0 & i_8_304_430_0 & ~i_8_304_578_0 & ~i_8_304_1180_0 & ~i_8_304_1468_0) | (~i_8_304_287_0 & ~i_8_304_304_0 & i_8_304_383_0 & ~i_8_304_817_0 & ~i_8_304_1315_0 & ~i_8_304_1394_0 & ~i_8_304_1469_0 & i_8_304_1534_0 & ~i_8_304_1747_0 & ~i_8_304_1889_0 & ~i_8_304_2070_0))) | (~i_8_304_113_0 & ~i_8_304_428_0 & ~i_8_304_577_0 & ~i_8_304_578_0 & i_8_304_713_0 & ~i_8_304_816_0 & ~i_8_304_1621_0 & i_8_304_1747_0 & ~i_8_304_1765_0))) | (~i_8_304_304_0 & i_8_304_430_0 & ~i_8_304_567_0 & i_8_304_710_0 & ~i_8_304_1470_0) | (i_8_304_19_0 & i_8_304_847_0 & ~i_8_304_1365_0 & ~i_8_304_1693_0 & i_8_304_1786_0))) | (~i_8_304_578_0 & ((~i_8_304_111_0 & ((~i_8_304_113_0 & ~i_8_304_266_0 & ~i_8_304_295_0 & i_8_304_524_0 & ~i_8_304_817_0 & ~i_8_304_1180_0 & ~i_8_304_1621_0 & ~i_8_304_1693_0 & ~i_8_304_1785_0 & i_8_304_1787_0) | (~i_8_304_112_0 & ~i_8_304_286_0 & ~i_8_304_635_0 & i_8_304_705_0 & ~i_8_304_715_0 & ~i_8_304_726_0 & ~i_8_304_1683_0 & ~i_8_304_1765_0 & ~i_8_304_1784_0 & ~i_8_304_1854_0 & ~i_8_304_2070_0))) | (~i_8_304_635_0 & ((~i_8_304_266_0 & ~i_8_304_269_0 & ~i_8_304_296_0 & i_8_304_710_0 & ~i_8_304_1365_0 & i_8_304_1826_0 & ~i_8_304_1854_0 & ~i_8_304_1874_0) | (~i_8_304_838_0 & ~i_8_304_878_0 & ~i_8_304_112_0 & ~i_8_304_427_0 & ~i_8_304_1180_0 & i_8_304_1469_0 & ~i_8_304_1565_0 & ~i_8_304_2088_0))) | (i_8_304_847_0 & ~i_8_304_2243_0 & ((~i_8_304_87_0 & i_8_304_504_0 & ~i_8_304_567_0 & ~i_8_304_1359_0 & ~i_8_304_1683_0 & ~i_8_304_1694_0) | (~i_8_304_1078_0 & ~i_8_304_1179_0 & ~i_8_304_286_0 & ~i_8_304_606_0 & ~i_8_304_1365_0 & ~i_8_304_1693_0 & ~i_8_304_1765_0 & ~i_8_304_1825_0 & ~i_8_304_2070_0))) | (~i_8_304_383_0 & i_8_304_713_0 & ~i_8_304_1365_0 & ~i_8_304_1565_0 & ~i_8_304_1684_0 & ~i_8_304_1694_0 & i_8_304_1787_0 & ~i_8_304_2070_0 & ~i_8_304_2071_0))) | (~i_8_304_427_0 & ((~i_8_304_87_0 & ~i_8_304_304_0 & i_8_304_708_0 & i_8_304_709_0 & ~i_8_304_1179_0 & ~i_8_304_1399_0 & ~i_8_304_1765_0) | (~i_8_304_305_0 & ~i_8_304_1078_0 & ~i_8_304_1469_0 & i_8_304_1472_0 & ~i_8_304_1534_0 & ~i_8_304_1730_0 & ~i_8_304_1920_0))) | (~i_8_304_305_0 & ((i_8_304_383_0 & ~i_8_304_817_0 & ~i_8_304_878_0 & ~i_8_304_1399_0 & ~i_8_304_1684_0 & ~i_8_304_1694_0 & ~i_8_304_1777_0 & i_8_304_1826_0) | (~i_8_304_87_0 & ~i_8_304_112_0 & ~i_8_304_113_0 & ~i_8_304_1078_0 & i_8_304_1889_0 & ~i_8_304_2071_0))) | (i_8_304_383_0 & ((~i_8_304_111_0 & i_8_304_112_0 & i_8_304_431_0 & ~i_8_304_817_0 & ~i_8_304_838_0 & ~i_8_304_1621_0) | (~i_8_304_219_0 & i_8_304_1399_0 & ~i_8_304_1920_0 & i_8_304_2060_0))) | (~i_8_304_219_0 & ((~i_8_304_112_0 & ~i_8_304_381_0 & ~i_8_304_1315_0 & ~i_8_304_1693_0 & ~i_8_304_2070_0 & i_8_304_2088_0) | (~i_8_304_87_0 & ~i_8_304_705_0 & ~i_8_304_715_0 & ~i_8_304_1920_0 & i_8_304_2274_0))) | (~i_8_304_1394_0 & ((~i_8_304_112_0 & ((~i_8_304_87_0 & ~i_8_304_381_0 & ~i_8_304_567_0 & ~i_8_304_607_0 & ~i_8_304_838_0 & ~i_8_304_1078_0 & ~i_8_304_1189_0 & ~i_8_304_1399_0 & ~i_8_304_1468_0 & ~i_8_304_1765_0 & ~i_8_304_1825_0 & i_8_304_1920_0) | (~i_8_304_19_0 & ~i_8_304_286_0 & ~i_8_304_287_0 & i_8_304_431_0 & ~i_8_304_817_0 & ~i_8_304_1179_0 & ~i_8_304_1694_0 & i_8_304_1787_0 & ~i_8_304_2274_0))) | (~i_8_304_286_0 & ~i_8_304_1694_0 & ~i_8_304_1784_0 & ((~i_8_304_295_0 & ~i_8_304_296_0 & ~i_8_304_383_0 & i_8_304_431_0 & ~i_8_304_569_0 & ~i_8_304_1359_0 & ~i_8_304_1365_0 & ~i_8_304_1693_0 & ~i_8_304_1777_0) | (~i_8_304_287_0 & ~i_8_304_577_0 & i_8_304_635_0 & ~i_8_304_1469_0 & ~i_8_304_1747_0 & ~i_8_304_1854_0 & i_8_304_2138_0))) | (~i_8_304_838_0 & ~i_8_304_1329_0 & ~i_8_304_1399_0 & ~i_8_304_1683_0 & ((~i_8_304_381_0 & ~i_8_304_816_0 & ~i_8_304_847_0 & ~i_8_304_1266_0 & ~i_8_304_1315_0 & i_8_304_1825_0) | (~i_8_304_383_0 & ~i_8_304_429_0 & ~i_8_304_715_0 & ~i_8_304_1179_0 & ~i_8_304_1522_0 & ~i_8_304_1621_0 & ~i_8_304_1693_0 & ~i_8_304_1730_0 & i_8_304_1785_0 & ~i_8_304_2139_0))) | (~i_8_304_295_0 & i_8_304_429_0 & ~i_8_304_726_0 & ~i_8_304_878_0 & ~i_8_304_1179_0 & ~i_8_304_1189_0 & ~i_8_304_1365_0 & i_8_304_1399_0 & ~i_8_304_1470_0))) | (~i_8_304_1683_0 & ((~i_8_304_87_0 & ((i_8_304_111_0 & i_8_304_705_0 & ~i_8_304_1749_0 & ~i_8_304_1786_0 & ~i_8_304_1825_0 & i_8_304_1920_0) | (i_8_304_219_0 & ~i_8_304_296_0 & ~i_8_304_726_0 & ~i_8_304_1359_0 & ~i_8_304_1399_0 & ~i_8_304_1470_0 & i_8_304_1889_0 & ~i_8_304_2060_0 & ~i_8_304_2227_0))) | (~i_8_304_113_0 & ((~i_8_304_295_0 & i_8_304_429_0 & i_8_304_430_0 & ~i_8_304_715_0 & ~i_8_304_726_0 & ~i_8_304_1180_0 & ~i_8_304_1399_0) | (i_8_304_606_0 & i_8_304_635_0 & ~i_8_304_838_0 & ~i_8_304_1179_0 & ~i_8_304_1359_0 & ~i_8_304_1730_0))) | (~i_8_304_568_0 & i_8_304_606_0 & ((~i_8_304_816_0 & i_8_304_846_0 & ~i_8_304_1621_0 & ~i_8_304_1854_0) | (~i_8_304_1359_0 & ~i_8_304_1522_0 & ~i_8_304_1693_0 & ~i_8_304_1694_0 & i_8_304_1777_0 & i_8_304_1786_0 & ~i_8_304_1873_0))) | (~i_8_304_1078_0 & ((~i_8_304_838_0 & ~i_8_304_1693_0 & i_8_304_2088_0 & i_8_304_2233_0) | (~i_8_304_295_0 & ~i_8_304_816_0 & ~i_8_304_1621_0 & ~i_8_304_1730_0 & ~i_8_304_1854_0 & ~i_8_304_2139_0 & i_8_304_2226_0 & ~i_8_304_2233_0))) | (~i_8_304_816_0 & ~i_8_304_1179_0 & ~i_8_304_1315_0 & ((i_8_304_429_0 & i_8_304_1780_0 & i_8_304_1785_0) | (~i_8_304_567_0 & ~i_8_304_635_0 & i_8_304_705_0 & ~i_8_304_1359_0 & ~i_8_304_1920_0))))) | (~i_8_304_295_0 & ((~i_8_304_111_0 & ((i_8_304_219_0 & ~i_8_304_287_0 & ~i_8_304_381_0 & ~i_8_304_577_0 & ~i_8_304_726_0 & ~i_8_304_1078_0 & ~i_8_304_1179_0 & ~i_8_304_1565_0 & i_8_304_1749_0 & ~i_8_304_1784_0 & ~i_8_304_2070_0) | (~i_8_304_286_0 & i_8_304_429_0 & ~i_8_304_1266_0 & ~i_8_304_2243_0 & i_8_304_2274_0))) | (~i_8_304_1359_0 & ((i_8_304_705_0 & ((~i_8_304_567_0 & i_8_304_606_0 & ~i_8_304_1180_0 & ~i_8_304_1470_0 & ~i_8_304_1522_0 & i_8_304_1747_0 & ~i_8_304_2139_0) | (i_8_304_708_0 & ~i_8_304_816_0 & ~i_8_304_1179_0 & ~i_8_304_1854_0 & ~i_8_304_2233_0 & i_8_304_2274_0))) | (~i_8_304_269_0 & ~i_8_304_296_0 & i_8_304_427_0 & ~i_8_304_568_0 & ~i_8_304_607_0 & ~i_8_304_726_0 & ~i_8_304_1565_0 & ~i_8_304_1621_0 & i_8_304_1825_0))) | (~i_8_304_2070_0 & ((~i_8_304_577_0 & ~i_8_304_816_0 & ~i_8_304_1179_0 & ~i_8_304_1180_0 & i_8_304_1467_0 & ~i_8_304_1522_0 & i_8_304_1747_0) | (i_8_304_219_0 & i_8_304_430_0 & ~i_8_304_606_0 & ~i_8_304_1078_0 & ~i_8_304_1621_0 & ~i_8_304_1749_0))))) | (~i_8_304_269_0 & ((~i_8_304_111_0 & i_8_304_428_0 & ~i_8_304_430_0 & ~i_8_304_1693_0 & ~i_8_304_1730_0 & i_8_304_1787_0 & ~i_8_304_1946_0 & ~i_8_304_2070_0 & i_8_304_2138_0) | (i_8_304_713_0 & ~i_8_304_838_0 & ~i_8_304_878_0 & ~i_8_304_1078_0 & ~i_8_304_1694_0 & ~i_8_304_1747_0 & ~i_8_304_1874_0 & ~i_8_304_2243_0))) | (~i_8_304_296_0 & ((~i_8_304_112_0 & ~i_8_304_838_0 & ~i_8_304_847_0 & ~i_8_304_1179_0 & ~i_8_304_1180_0 & ~i_8_304_1359_0 & ~i_8_304_1365_0 & ~i_8_304_1472_0 & i_8_304_1749_0 & i_8_304_1785_0) | (~i_8_304_635_0 & ~i_8_304_1266_0 & ~i_8_304_1693_0 & ~i_8_304_1730_0 & i_8_304_1874_0))) | (i_8_304_429_0 & ((i_8_304_381_0 & ~i_8_304_606_0 & ~i_8_304_1078_0 & ~i_8_304_1329_0 & i_8_304_1777_0) | (~i_8_304_111_0 & i_8_304_708_0 & ~i_8_304_816_0 & ~i_8_304_838_0 & ~i_8_304_2139_0))) | (~i_8_304_1359_0 & ((~i_8_304_304_0 & i_8_304_1749_0 & ((~i_8_304_577_0 & i_8_304_708_0 & ~i_8_304_1180_0 & i_8_304_1266_0 & ~i_8_304_1565_0 & ~i_8_304_1621_0) | (~i_8_304_567_0 & ~i_8_304_715_0 & ~i_8_304_1315_0 & ~i_8_304_1399_0 & ~i_8_304_1470_0 & ~i_8_304_1693_0 & i_8_304_1785_0 & ~i_8_304_1825_0 & ~i_8_304_2243_0))) | (~i_8_304_111_0 & ~i_8_304_381_0 & ~i_8_304_568_0 & ~i_8_304_577_0 & i_8_304_846_0 & ~i_8_304_1078_0 & ~i_8_304_1179_0 & ~i_8_304_1180_0 & ~i_8_304_1315_0 & ~i_8_304_1621_0 & ~i_8_304_2226_0))) | (~i_8_304_878_0 & ((~i_8_304_111_0 & ((i_8_304_606_0 & ~i_8_304_1621_0 & i_8_304_2227_0) | (~i_8_304_113_0 & ~i_8_304_304_0 & ~i_8_304_381_0 & ~i_8_304_383_0 & ~i_8_304_705_0 & ~i_8_304_1329_0 & ~i_8_304_1534_0 & ~i_8_304_1747_0 & ~i_8_304_1749_0 & i_8_304_1785_0 & ~i_8_304_1786_0 & ~i_8_304_2070_0 & ~i_8_304_2274_0))) | (i_8_304_715_0 & ((i_8_304_1399_0 & ~i_8_304_1777_0 & i_8_304_1786_0) | (~i_8_304_381_0 & ~i_8_304_705_0 & ~i_8_304_1749_0 & i_8_304_1777_0 & ~i_8_304_1786_0 & ~i_8_304_2227_0))) | (~i_8_304_715_0 & ~i_8_304_838_0 & ~i_8_304_1534_0 & i_8_304_1747_0 & ~i_8_304_1787_0 & ~i_8_304_1920_0 & ~i_8_304_2070_0 & ~i_8_304_2243_0))) | (i_8_304_430_0 & ~i_8_304_726_0 & ~i_8_304_1078_0 & ~i_8_304_1765_0 & i_8_304_1780_0 & i_8_304_1825_0 & ~i_8_304_2070_0));
endmodule



// Benchmark "kernel_8_305" written by ABC on Sun Jul 19 10:08:24 2020

module kernel_8_305 ( 
    i_8_305_21_0, i_8_305_30_0, i_8_305_31_0, i_8_305_35_0, i_8_305_53_0,
    i_8_305_57_0, i_8_305_114_0, i_8_305_116_0, i_8_305_142_0,
    i_8_305_143_0, i_8_305_171_0, i_8_305_188_0, i_8_305_192_0,
    i_8_305_225_0, i_8_305_238_0, i_8_305_246_0, i_8_305_395_0,
    i_8_305_415_0, i_8_305_422_0, i_8_305_446_0, i_8_305_585_0,
    i_8_305_598_0, i_8_305_599_0, i_8_305_611_0, i_8_305_698_0,
    i_8_305_701_0, i_8_305_716_0, i_8_305_759_0, i_8_305_780_0,
    i_8_305_781_0, i_8_305_815_0, i_8_305_818_0, i_8_305_823_0,
    i_8_305_841_0, i_8_305_845_0, i_8_305_849_0, i_8_305_853_0,
    i_8_305_888_0, i_8_305_959_0, i_8_305_964_0, i_8_305_1016_0,
    i_8_305_1030_0, i_8_305_1034_0, i_8_305_1050_0, i_8_305_1051_0,
    i_8_305_1060_0, i_8_305_1114_0, i_8_305_1121_0, i_8_305_1160_0,
    i_8_305_1182_0, i_8_305_1183_0, i_8_305_1281_0, i_8_305_1282_0,
    i_8_305_1283_0, i_8_305_1284_0, i_8_305_1291_0, i_8_305_1300_0,
    i_8_305_1305_0, i_8_305_1306_0, i_8_305_1307_0, i_8_305_1330_0,
    i_8_305_1344_0, i_8_305_1347_0, i_8_305_1390_0, i_8_305_1391_0,
    i_8_305_1410_0, i_8_305_1437_0, i_8_305_1438_0, i_8_305_1453_0,
    i_8_305_1470_0, i_8_305_1471_0, i_8_305_1552_0, i_8_305_1574_0,
    i_8_305_1652_0, i_8_305_1677_0, i_8_305_1683_0, i_8_305_1699_0,
    i_8_305_1754_0, i_8_305_1875_0, i_8_305_1876_0, i_8_305_1877_0,
    i_8_305_1984_0, i_8_305_1988_0, i_8_305_1991_0, i_8_305_1992_0,
    i_8_305_1995_0, i_8_305_2033_0, i_8_305_2071_0, i_8_305_2076_0,
    i_8_305_2093_0, i_8_305_2114_0, i_8_305_2132_0, i_8_305_2151_0,
    i_8_305_2214_0, i_8_305_2215_0, i_8_305_2216_0, i_8_305_2237_0,
    i_8_305_2245_0, i_8_305_2261_0, i_8_305_2290_0,
    o_8_305_0_0  );
  input  i_8_305_21_0, i_8_305_30_0, i_8_305_31_0, i_8_305_35_0,
    i_8_305_53_0, i_8_305_57_0, i_8_305_114_0, i_8_305_116_0,
    i_8_305_142_0, i_8_305_143_0, i_8_305_171_0, i_8_305_188_0,
    i_8_305_192_0, i_8_305_225_0, i_8_305_238_0, i_8_305_246_0,
    i_8_305_395_0, i_8_305_415_0, i_8_305_422_0, i_8_305_446_0,
    i_8_305_585_0, i_8_305_598_0, i_8_305_599_0, i_8_305_611_0,
    i_8_305_698_0, i_8_305_701_0, i_8_305_716_0, i_8_305_759_0,
    i_8_305_780_0, i_8_305_781_0, i_8_305_815_0, i_8_305_818_0,
    i_8_305_823_0, i_8_305_841_0, i_8_305_845_0, i_8_305_849_0,
    i_8_305_853_0, i_8_305_888_0, i_8_305_959_0, i_8_305_964_0,
    i_8_305_1016_0, i_8_305_1030_0, i_8_305_1034_0, i_8_305_1050_0,
    i_8_305_1051_0, i_8_305_1060_0, i_8_305_1114_0, i_8_305_1121_0,
    i_8_305_1160_0, i_8_305_1182_0, i_8_305_1183_0, i_8_305_1281_0,
    i_8_305_1282_0, i_8_305_1283_0, i_8_305_1284_0, i_8_305_1291_0,
    i_8_305_1300_0, i_8_305_1305_0, i_8_305_1306_0, i_8_305_1307_0,
    i_8_305_1330_0, i_8_305_1344_0, i_8_305_1347_0, i_8_305_1390_0,
    i_8_305_1391_0, i_8_305_1410_0, i_8_305_1437_0, i_8_305_1438_0,
    i_8_305_1453_0, i_8_305_1470_0, i_8_305_1471_0, i_8_305_1552_0,
    i_8_305_1574_0, i_8_305_1652_0, i_8_305_1677_0, i_8_305_1683_0,
    i_8_305_1699_0, i_8_305_1754_0, i_8_305_1875_0, i_8_305_1876_0,
    i_8_305_1877_0, i_8_305_1984_0, i_8_305_1988_0, i_8_305_1991_0,
    i_8_305_1992_0, i_8_305_1995_0, i_8_305_2033_0, i_8_305_2071_0,
    i_8_305_2076_0, i_8_305_2093_0, i_8_305_2114_0, i_8_305_2132_0,
    i_8_305_2151_0, i_8_305_2214_0, i_8_305_2215_0, i_8_305_2216_0,
    i_8_305_2237_0, i_8_305_2245_0, i_8_305_2261_0, i_8_305_2290_0;
  output o_8_305_0_0;
  assign o_8_305_0_0 = ~((~i_8_305_57_0 & ((~i_8_305_1281_0 & ~i_8_305_1300_0 & ~i_8_305_1347_0 & ~i_8_305_1390_0 & i_8_305_1410_0 & i_8_305_1552_0 & ~i_8_305_1699_0) | (~i_8_305_246_0 & ~i_8_305_422_0 & ~i_8_305_1305_0 & ~i_8_305_1876_0 & ~i_8_305_2093_0))) | (~i_8_305_142_0 & ((~i_8_305_21_0 & ~i_8_305_598_0 & ~i_8_305_959_0 & ~i_8_305_1391_0 & ~i_8_305_1471_0 & ~i_8_305_1683_0) | (~i_8_305_246_0 & ~i_8_305_599_0 & ~i_8_305_759_0 & ~i_8_305_1330_0 & ~i_8_305_1875_0 & i_8_305_2215_0 & ~i_8_305_2237_0))) | (~i_8_305_1470_0 & ((~i_8_305_21_0 & ~i_8_305_1330_0 & ((~i_8_305_598_0 & ~i_8_305_1051_0 & ~i_8_305_1574_0 & ~i_8_305_1875_0 & ~i_8_305_1991_0) | (~i_8_305_415_0 & ~i_8_305_1060_0 & ~i_8_305_1291_0 & ~i_8_305_1347_0 & ~i_8_305_1410_0 & ~i_8_305_1876_0 & ~i_8_305_2033_0))) | (~i_8_305_188_0 & ~i_8_305_759_0 & ~i_8_305_1114_0 & ~i_8_305_1306_0 & ~i_8_305_1471_0 & ~i_8_305_1754_0))) | (~i_8_305_192_0 & ~i_8_305_225_0 & ((~i_8_305_171_0 & i_8_305_1284_0 & ~i_8_305_1877_0) | (~i_8_305_611_0 & ~i_8_305_1060_0 & ~i_8_305_1410_0 & ~i_8_305_2214_0 & ~i_8_305_2215_0))) | (~i_8_305_246_0 & ~i_8_305_446_0 & ~i_8_305_716_0 & ((~i_8_305_585_0 & ~i_8_305_759_0 & ~i_8_305_818_0 & ~i_8_305_849_0 & ~i_8_305_1050_0 & ~i_8_305_1437_0) | (~i_8_305_888_0 & ~i_8_305_959_0 & ~i_8_305_1347_0 & ~i_8_305_1453_0 & ~i_8_305_1677_0 & ~i_8_305_1699_0 & ~i_8_305_1876_0 & i_8_305_1992_0 & ~i_8_305_2214_0))) | (~i_8_305_818_0 & ((~i_8_305_171_0 & ~i_8_305_1471_0 & i_8_305_1699_0) | (~i_8_305_845_0 & i_8_305_1284_0 & ~i_8_305_1875_0 & ~i_8_305_1877_0 & ~i_8_305_1988_0))) | (~i_8_305_171_0 & ((~i_8_305_422_0 & i_8_305_759_0 & ~i_8_305_888_0 & ~i_8_305_1300_0 & ~i_8_305_1875_0 & ~i_8_305_1991_0 & ~i_8_305_1992_0) | (~i_8_305_53_0 & ~i_8_305_841_0 & ~i_8_305_959_0 & i_8_305_1114_0 & ~i_8_305_1281_0 & ~i_8_305_1306_0 & ~i_8_305_2290_0))) | (~i_8_305_53_0 & ((~i_8_305_849_0 & ~i_8_305_853_0 & ~i_8_305_1114_0 & ~i_8_305_1391_0 & ~i_8_305_1875_0 & ~i_8_305_1992_0 & ~i_8_305_1995_0) | (~i_8_305_1051_0 & ~i_8_305_1183_0 & ~i_8_305_1305_0 & ~i_8_305_1306_0 & ~i_8_305_1877_0 & ~i_8_305_2214_0 & ~i_8_305_2261_0))) | (~i_8_305_1875_0 & ~i_8_305_2216_0 & ((~i_8_305_238_0 & ~i_8_305_759_0 & ~i_8_305_1307_0 & ~i_8_305_1390_0 & ~i_8_305_1877_0 & ~i_8_305_2215_0) | (~i_8_305_1121_0 & i_8_305_1438_0 & ~i_8_305_2261_0))) | (~i_8_305_1390_0 & ((~i_8_305_1050_0 & i_8_305_1282_0 & ~i_8_305_1652_0 & ~i_8_305_2033_0) | (~i_8_305_116_0 & ~i_8_305_143_0 & ~i_8_305_1305_0 & ~i_8_305_1410_0 & ~i_8_305_1992_0 & ~i_8_305_2114_0 & ~i_8_305_2214_0))) | i_8_305_1160_0 | (i_8_305_841_0 & i_8_305_853_0 & ~i_8_305_1552_0 & i_8_305_2093_0));
endmodule



// Benchmark "kernel_8_306" written by ABC on Sun Jul 19 10:08:25 2020

module kernel_8_306 ( 
    i_8_306_9_0, i_8_306_10_0, i_8_306_47_0, i_8_306_112_0, i_8_306_118_0,
    i_8_306_136_0, i_8_306_137_0, i_8_306_139_0, i_8_306_140_0,
    i_8_306_221_0, i_8_306_230_0, i_8_306_265_0, i_8_306_316_0,
    i_8_306_383_0, i_8_306_391_0, i_8_306_398_0, i_8_306_414_0,
    i_8_306_415_0, i_8_306_417_0, i_8_306_425_0, i_8_306_427_0,
    i_8_306_478_0, i_8_306_481_0, i_8_306_510_0, i_8_306_522_0,
    i_8_306_524_0, i_8_306_526_0, i_8_306_528_0, i_8_306_553_0,
    i_8_306_554_0, i_8_306_568_0, i_8_306_577_0, i_8_306_585_0,
    i_8_306_632_0, i_8_306_640_0, i_8_306_651_0, i_8_306_704_0,
    i_8_306_730_0, i_8_306_784_0, i_8_306_792_0, i_8_306_793_0,
    i_8_306_823_0, i_8_306_837_0, i_8_306_847_0, i_8_306_859_0,
    i_8_306_874_0, i_8_306_887_0, i_8_306_892_0, i_8_306_964_0,
    i_8_306_991_0, i_8_306_1036_0, i_8_306_1072_0, i_8_306_1111_0,
    i_8_306_1199_0, i_8_306_1237_0, i_8_306_1315_0, i_8_306_1324_0,
    i_8_306_1352_0, i_8_306_1354_0, i_8_306_1360_0, i_8_306_1372_0,
    i_8_306_1388_0, i_8_306_1396_0, i_8_306_1438_0, i_8_306_1458_0,
    i_8_306_1459_0, i_8_306_1470_0, i_8_306_1477_0, i_8_306_1513_0,
    i_8_306_1521_0, i_8_306_1540_0, i_8_306_1566_0, i_8_306_1567_0,
    i_8_306_1571_0, i_8_306_1603_0, i_8_306_1630_0, i_8_306_1684_0,
    i_8_306_1693_0, i_8_306_1720_0, i_8_306_1751_0, i_8_306_1776_0,
    i_8_306_1777_0, i_8_306_1778_0, i_8_306_1781_0, i_8_306_1786_0,
    i_8_306_1837_0, i_8_306_1864_0, i_8_306_1885_0, i_8_306_1900_0,
    i_8_306_1935_0, i_8_306_1936_0, i_8_306_1954_0, i_8_306_1972_0,
    i_8_306_1993_0, i_8_306_2026_0, i_8_306_2092_0, i_8_306_2138_0,
    i_8_306_2147_0, i_8_306_2170_0, i_8_306_2241_0,
    o_8_306_0_0  );
  input  i_8_306_9_0, i_8_306_10_0, i_8_306_47_0, i_8_306_112_0,
    i_8_306_118_0, i_8_306_136_0, i_8_306_137_0, i_8_306_139_0,
    i_8_306_140_0, i_8_306_221_0, i_8_306_230_0, i_8_306_265_0,
    i_8_306_316_0, i_8_306_383_0, i_8_306_391_0, i_8_306_398_0,
    i_8_306_414_0, i_8_306_415_0, i_8_306_417_0, i_8_306_425_0,
    i_8_306_427_0, i_8_306_478_0, i_8_306_481_0, i_8_306_510_0,
    i_8_306_522_0, i_8_306_524_0, i_8_306_526_0, i_8_306_528_0,
    i_8_306_553_0, i_8_306_554_0, i_8_306_568_0, i_8_306_577_0,
    i_8_306_585_0, i_8_306_632_0, i_8_306_640_0, i_8_306_651_0,
    i_8_306_704_0, i_8_306_730_0, i_8_306_784_0, i_8_306_792_0,
    i_8_306_793_0, i_8_306_823_0, i_8_306_837_0, i_8_306_847_0,
    i_8_306_859_0, i_8_306_874_0, i_8_306_887_0, i_8_306_892_0,
    i_8_306_964_0, i_8_306_991_0, i_8_306_1036_0, i_8_306_1072_0,
    i_8_306_1111_0, i_8_306_1199_0, i_8_306_1237_0, i_8_306_1315_0,
    i_8_306_1324_0, i_8_306_1352_0, i_8_306_1354_0, i_8_306_1360_0,
    i_8_306_1372_0, i_8_306_1388_0, i_8_306_1396_0, i_8_306_1438_0,
    i_8_306_1458_0, i_8_306_1459_0, i_8_306_1470_0, i_8_306_1477_0,
    i_8_306_1513_0, i_8_306_1521_0, i_8_306_1540_0, i_8_306_1566_0,
    i_8_306_1567_0, i_8_306_1571_0, i_8_306_1603_0, i_8_306_1630_0,
    i_8_306_1684_0, i_8_306_1693_0, i_8_306_1720_0, i_8_306_1751_0,
    i_8_306_1776_0, i_8_306_1777_0, i_8_306_1778_0, i_8_306_1781_0,
    i_8_306_1786_0, i_8_306_1837_0, i_8_306_1864_0, i_8_306_1885_0,
    i_8_306_1900_0, i_8_306_1935_0, i_8_306_1936_0, i_8_306_1954_0,
    i_8_306_1972_0, i_8_306_1993_0, i_8_306_2026_0, i_8_306_2092_0,
    i_8_306_2138_0, i_8_306_2147_0, i_8_306_2170_0, i_8_306_2241_0;
  output o_8_306_0_0;
  assign o_8_306_0_0 = 0;
endmodule



// Benchmark "kernel_8_307" written by ABC on Sun Jul 19 10:08:26 2020

module kernel_8_307 ( 
    i_8_307_85_0, i_8_307_88_0, i_8_307_91_0, i_8_307_181_0, i_8_307_189_0,
    i_8_307_190_0, i_8_307_220_0, i_8_307_292_0, i_8_307_305_0,
    i_8_307_370_0, i_8_307_372_0, i_8_307_417_0, i_8_307_418_0,
    i_8_307_476_0, i_8_307_481_0, i_8_307_483_0, i_8_307_546_0,
    i_8_307_556_0, i_8_307_595_0, i_8_307_634_0, i_8_307_648_0,
    i_8_307_672_0, i_8_307_703_0, i_8_307_705_0, i_8_307_728_0,
    i_8_307_759_0, i_8_307_764_0, i_8_307_797_0, i_8_307_811_0,
    i_8_307_855_0, i_8_307_872_0, i_8_307_898_0, i_8_307_899_0,
    i_8_307_966_0, i_8_307_991_0, i_8_307_1000_0, i_8_307_1030_0,
    i_8_307_1060_0, i_8_307_1061_0, i_8_307_1111_0, i_8_307_1121_0,
    i_8_307_1179_0, i_8_307_1191_0, i_8_307_1285_0, i_8_307_1291_0,
    i_8_307_1296_0, i_8_307_1297_0, i_8_307_1305_0, i_8_307_1316_0,
    i_8_307_1319_0, i_8_307_1323_0, i_8_307_1327_0, i_8_307_1455_0,
    i_8_307_1456_0, i_8_307_1469_0, i_8_307_1490_0, i_8_307_1509_0,
    i_8_307_1528_0, i_8_307_1529_0, i_8_307_1531_0, i_8_307_1544_0,
    i_8_307_1553_0, i_8_307_1561_0, i_8_307_1588_0, i_8_307_1603_0,
    i_8_307_1618_0, i_8_307_1669_0, i_8_307_1678_0, i_8_307_1718_0,
    i_8_307_1737_0, i_8_307_1738_0, i_8_307_1752_0, i_8_307_1753_0,
    i_8_307_1754_0, i_8_307_1761_0, i_8_307_1803_0, i_8_307_1805_0,
    i_8_307_1808_0, i_8_307_1839_0, i_8_307_1857_0, i_8_307_1867_0,
    i_8_307_1874_0, i_8_307_1904_0, i_8_307_1906_0, i_8_307_1911_0,
    i_8_307_1933_0, i_8_307_1981_0, i_8_307_2006_0, i_8_307_2032_0,
    i_8_307_2046_0, i_8_307_2047_0, i_8_307_2116_0, i_8_307_2142_0,
    i_8_307_2152_0, i_8_307_2153_0, i_8_307_2216_0, i_8_307_2218_0,
    i_8_307_2254_0, i_8_307_2290_0, i_8_307_2296_0,
    o_8_307_0_0  );
  input  i_8_307_85_0, i_8_307_88_0, i_8_307_91_0, i_8_307_181_0,
    i_8_307_189_0, i_8_307_190_0, i_8_307_220_0, i_8_307_292_0,
    i_8_307_305_0, i_8_307_370_0, i_8_307_372_0, i_8_307_417_0,
    i_8_307_418_0, i_8_307_476_0, i_8_307_481_0, i_8_307_483_0,
    i_8_307_546_0, i_8_307_556_0, i_8_307_595_0, i_8_307_634_0,
    i_8_307_648_0, i_8_307_672_0, i_8_307_703_0, i_8_307_705_0,
    i_8_307_728_0, i_8_307_759_0, i_8_307_764_0, i_8_307_797_0,
    i_8_307_811_0, i_8_307_855_0, i_8_307_872_0, i_8_307_898_0,
    i_8_307_899_0, i_8_307_966_0, i_8_307_991_0, i_8_307_1000_0,
    i_8_307_1030_0, i_8_307_1060_0, i_8_307_1061_0, i_8_307_1111_0,
    i_8_307_1121_0, i_8_307_1179_0, i_8_307_1191_0, i_8_307_1285_0,
    i_8_307_1291_0, i_8_307_1296_0, i_8_307_1297_0, i_8_307_1305_0,
    i_8_307_1316_0, i_8_307_1319_0, i_8_307_1323_0, i_8_307_1327_0,
    i_8_307_1455_0, i_8_307_1456_0, i_8_307_1469_0, i_8_307_1490_0,
    i_8_307_1509_0, i_8_307_1528_0, i_8_307_1529_0, i_8_307_1531_0,
    i_8_307_1544_0, i_8_307_1553_0, i_8_307_1561_0, i_8_307_1588_0,
    i_8_307_1603_0, i_8_307_1618_0, i_8_307_1669_0, i_8_307_1678_0,
    i_8_307_1718_0, i_8_307_1737_0, i_8_307_1738_0, i_8_307_1752_0,
    i_8_307_1753_0, i_8_307_1754_0, i_8_307_1761_0, i_8_307_1803_0,
    i_8_307_1805_0, i_8_307_1808_0, i_8_307_1839_0, i_8_307_1857_0,
    i_8_307_1867_0, i_8_307_1874_0, i_8_307_1904_0, i_8_307_1906_0,
    i_8_307_1911_0, i_8_307_1933_0, i_8_307_1981_0, i_8_307_2006_0,
    i_8_307_2032_0, i_8_307_2046_0, i_8_307_2047_0, i_8_307_2116_0,
    i_8_307_2142_0, i_8_307_2152_0, i_8_307_2153_0, i_8_307_2216_0,
    i_8_307_2218_0, i_8_307_2254_0, i_8_307_2290_0, i_8_307_2296_0;
  output o_8_307_0_0;
  assign o_8_307_0_0 = 0;
endmodule



// Benchmark "kernel_8_308" written by ABC on Sun Jul 19 10:08:26 2020

module kernel_8_308 ( 
    i_8_308_22_0, i_8_308_23_0, i_8_308_28_0, i_8_308_50_0, i_8_308_140_0,
    i_8_308_202_0, i_8_308_260_0, i_8_308_262_0, i_8_308_263_0,
    i_8_308_281_0, i_8_308_289_0, i_8_308_291_0, i_8_308_301_0,
    i_8_308_302_0, i_8_308_322_0, i_8_308_345_0, i_8_308_346_0,
    i_8_308_362_0, i_8_308_375_0, i_8_308_381_0, i_8_308_382_0,
    i_8_308_391_0, i_8_308_460_0, i_8_308_505_0, i_8_308_517_0,
    i_8_308_523_0, i_8_308_525_0, i_8_308_526_0, i_8_308_529_0,
    i_8_308_553_0, i_8_308_670_0, i_8_308_702_0, i_8_308_763_0,
    i_8_308_769_0, i_8_308_775_0, i_8_308_804_0, i_8_308_805_0,
    i_8_308_832_0, i_8_308_892_0, i_8_308_905_0, i_8_308_968_0,
    i_8_308_971_0, i_8_308_1067_0, i_8_308_1074_0, i_8_308_1138_0,
    i_8_308_1173_0, i_8_308_1182_0, i_8_308_1233_0, i_8_308_1254_0,
    i_8_308_1255_0, i_8_308_1260_0, i_8_308_1273_0, i_8_308_1279_0,
    i_8_308_1281_0, i_8_308_1282_0, i_8_308_1286_0, i_8_308_1300_0,
    i_8_308_1327_0, i_8_308_1384_0, i_8_308_1424_0, i_8_308_1435_0,
    i_8_308_1452_0, i_8_308_1467_0, i_8_308_1490_0, i_8_308_1498_0,
    i_8_308_1528_0, i_8_308_1533_0, i_8_308_1542_0, i_8_308_1555_0,
    i_8_308_1587_0, i_8_308_1597_0, i_8_308_1606_0, i_8_308_1630_0,
    i_8_308_1631_0, i_8_308_1632_0, i_8_308_1654_0, i_8_308_1660_0,
    i_8_308_1690_0, i_8_308_1696_0, i_8_308_1719_0, i_8_308_1720_0,
    i_8_308_1723_0, i_8_308_1724_0, i_8_308_1740_0, i_8_308_1762_0,
    i_8_308_1792_0, i_8_308_1808_0, i_8_308_1820_0, i_8_308_1837_0,
    i_8_308_1876_0, i_8_308_1990_0, i_8_308_2047_0, i_8_308_2089_0,
    i_8_308_2118_0, i_8_308_2126_0, i_8_308_2143_0, i_8_308_2154_0,
    i_8_308_2188_0, i_8_308_2234_0, i_8_308_2290_0,
    o_8_308_0_0  );
  input  i_8_308_22_0, i_8_308_23_0, i_8_308_28_0, i_8_308_50_0,
    i_8_308_140_0, i_8_308_202_0, i_8_308_260_0, i_8_308_262_0,
    i_8_308_263_0, i_8_308_281_0, i_8_308_289_0, i_8_308_291_0,
    i_8_308_301_0, i_8_308_302_0, i_8_308_322_0, i_8_308_345_0,
    i_8_308_346_0, i_8_308_362_0, i_8_308_375_0, i_8_308_381_0,
    i_8_308_382_0, i_8_308_391_0, i_8_308_460_0, i_8_308_505_0,
    i_8_308_517_0, i_8_308_523_0, i_8_308_525_0, i_8_308_526_0,
    i_8_308_529_0, i_8_308_553_0, i_8_308_670_0, i_8_308_702_0,
    i_8_308_763_0, i_8_308_769_0, i_8_308_775_0, i_8_308_804_0,
    i_8_308_805_0, i_8_308_832_0, i_8_308_892_0, i_8_308_905_0,
    i_8_308_968_0, i_8_308_971_0, i_8_308_1067_0, i_8_308_1074_0,
    i_8_308_1138_0, i_8_308_1173_0, i_8_308_1182_0, i_8_308_1233_0,
    i_8_308_1254_0, i_8_308_1255_0, i_8_308_1260_0, i_8_308_1273_0,
    i_8_308_1279_0, i_8_308_1281_0, i_8_308_1282_0, i_8_308_1286_0,
    i_8_308_1300_0, i_8_308_1327_0, i_8_308_1384_0, i_8_308_1424_0,
    i_8_308_1435_0, i_8_308_1452_0, i_8_308_1467_0, i_8_308_1490_0,
    i_8_308_1498_0, i_8_308_1528_0, i_8_308_1533_0, i_8_308_1542_0,
    i_8_308_1555_0, i_8_308_1587_0, i_8_308_1597_0, i_8_308_1606_0,
    i_8_308_1630_0, i_8_308_1631_0, i_8_308_1632_0, i_8_308_1654_0,
    i_8_308_1660_0, i_8_308_1690_0, i_8_308_1696_0, i_8_308_1719_0,
    i_8_308_1720_0, i_8_308_1723_0, i_8_308_1724_0, i_8_308_1740_0,
    i_8_308_1762_0, i_8_308_1792_0, i_8_308_1808_0, i_8_308_1820_0,
    i_8_308_1837_0, i_8_308_1876_0, i_8_308_1990_0, i_8_308_2047_0,
    i_8_308_2089_0, i_8_308_2118_0, i_8_308_2126_0, i_8_308_2143_0,
    i_8_308_2154_0, i_8_308_2188_0, i_8_308_2234_0, i_8_308_2290_0;
  output o_8_308_0_0;
  assign o_8_308_0_0 = 0;
endmodule



// Benchmark "kernel_8_309" written by ABC on Sun Jul 19 10:08:27 2020

module kernel_8_309 ( 
    i_8_309_46_0, i_8_309_52_0, i_8_309_87_0, i_8_309_142_0, i_8_309_171_0,
    i_8_309_172_0, i_8_309_210_0, i_8_309_259_0, i_8_309_294_0,
    i_8_309_334_0, i_8_309_364_0, i_8_309_376_0, i_8_309_381_0,
    i_8_309_383_0, i_8_309_390_0, i_8_309_436_0, i_8_309_487_0,
    i_8_309_489_0, i_8_309_492_0, i_8_309_532_0, i_8_309_534_0,
    i_8_309_550_0, i_8_309_551_0, i_8_309_576_0, i_8_309_581_0,
    i_8_309_585_0, i_8_309_609_0, i_8_309_630_0, i_8_309_676_0,
    i_8_309_684_0, i_8_309_699_0, i_8_309_736_0, i_8_309_765_0,
    i_8_309_766_0, i_8_309_769_0, i_8_309_792_0, i_8_309_795_0,
    i_8_309_839_0, i_8_309_841_0, i_8_309_879_0, i_8_309_880_0,
    i_8_309_919_0, i_8_309_927_0, i_8_309_930_0, i_8_309_965_0,
    i_8_309_966_0, i_8_309_991_0, i_8_309_1036_0, i_8_309_1053_0,
    i_8_309_1171_0, i_8_309_1233_0, i_8_309_1234_0, i_8_309_1255_0,
    i_8_309_1263_0, i_8_309_1266_0, i_8_309_1288_0, i_8_309_1308_0,
    i_8_309_1315_0, i_8_309_1316_0, i_8_309_1393_0, i_8_309_1455_0,
    i_8_309_1471_0, i_8_309_1544_0, i_8_309_1558_0, i_8_309_1642_0,
    i_8_309_1650_0, i_8_309_1668_0, i_8_309_1669_0, i_8_309_1683_0,
    i_8_309_1702_0, i_8_309_1729_0, i_8_309_1749_0, i_8_309_1777_0,
    i_8_309_1821_0, i_8_309_1828_0, i_8_309_1854_0, i_8_309_1857_0,
    i_8_309_1858_0, i_8_309_1861_0, i_8_309_1885_0, i_8_309_1938_0,
    i_8_309_1947_0, i_8_309_1950_0, i_8_309_1981_0, i_8_309_1989_0,
    i_8_309_2001_0, i_8_309_2016_0, i_8_309_2017_0, i_8_309_2056_0,
    i_8_309_2106_0, i_8_309_2139_0, i_8_309_2152_0, i_8_309_2155_0,
    i_8_309_2182_0, i_8_309_2196_0, i_8_309_2199_0, i_8_309_2205_0,
    i_8_309_2259_0, i_8_309_2272_0, i_8_309_2277_0,
    o_8_309_0_0  );
  input  i_8_309_46_0, i_8_309_52_0, i_8_309_87_0, i_8_309_142_0,
    i_8_309_171_0, i_8_309_172_0, i_8_309_210_0, i_8_309_259_0,
    i_8_309_294_0, i_8_309_334_0, i_8_309_364_0, i_8_309_376_0,
    i_8_309_381_0, i_8_309_383_0, i_8_309_390_0, i_8_309_436_0,
    i_8_309_487_0, i_8_309_489_0, i_8_309_492_0, i_8_309_532_0,
    i_8_309_534_0, i_8_309_550_0, i_8_309_551_0, i_8_309_576_0,
    i_8_309_581_0, i_8_309_585_0, i_8_309_609_0, i_8_309_630_0,
    i_8_309_676_0, i_8_309_684_0, i_8_309_699_0, i_8_309_736_0,
    i_8_309_765_0, i_8_309_766_0, i_8_309_769_0, i_8_309_792_0,
    i_8_309_795_0, i_8_309_839_0, i_8_309_841_0, i_8_309_879_0,
    i_8_309_880_0, i_8_309_919_0, i_8_309_927_0, i_8_309_930_0,
    i_8_309_965_0, i_8_309_966_0, i_8_309_991_0, i_8_309_1036_0,
    i_8_309_1053_0, i_8_309_1171_0, i_8_309_1233_0, i_8_309_1234_0,
    i_8_309_1255_0, i_8_309_1263_0, i_8_309_1266_0, i_8_309_1288_0,
    i_8_309_1308_0, i_8_309_1315_0, i_8_309_1316_0, i_8_309_1393_0,
    i_8_309_1455_0, i_8_309_1471_0, i_8_309_1544_0, i_8_309_1558_0,
    i_8_309_1642_0, i_8_309_1650_0, i_8_309_1668_0, i_8_309_1669_0,
    i_8_309_1683_0, i_8_309_1702_0, i_8_309_1729_0, i_8_309_1749_0,
    i_8_309_1777_0, i_8_309_1821_0, i_8_309_1828_0, i_8_309_1854_0,
    i_8_309_1857_0, i_8_309_1858_0, i_8_309_1861_0, i_8_309_1885_0,
    i_8_309_1938_0, i_8_309_1947_0, i_8_309_1950_0, i_8_309_1981_0,
    i_8_309_1989_0, i_8_309_2001_0, i_8_309_2016_0, i_8_309_2017_0,
    i_8_309_2056_0, i_8_309_2106_0, i_8_309_2139_0, i_8_309_2152_0,
    i_8_309_2155_0, i_8_309_2182_0, i_8_309_2196_0, i_8_309_2199_0,
    i_8_309_2205_0, i_8_309_2259_0, i_8_309_2272_0, i_8_309_2277_0;
  output o_8_309_0_0;
  assign o_8_309_0_0 = 0;
endmodule



// Benchmark "kernel_8_310" written by ABC on Sun Jul 19 10:08:28 2020

module kernel_8_310 ( 
    i_8_310_22_0, i_8_310_54_0, i_8_310_64_0, i_8_310_219_0, i_8_310_220_0,
    i_8_310_283_0, i_8_310_319_0, i_8_310_321_0, i_8_310_397_0,
    i_8_310_424_0, i_8_310_441_0, i_8_310_496_0, i_8_310_504_0,
    i_8_310_524_0, i_8_310_526_0, i_8_310_571_0, i_8_310_580_0,
    i_8_310_589_0, i_8_310_596_0, i_8_310_613_0, i_8_310_622_0,
    i_8_310_642_0, i_8_310_659_0, i_8_310_660_0, i_8_310_675_0,
    i_8_310_676_0, i_8_310_699_0, i_8_310_700_0, i_8_310_707_0,
    i_8_310_730_0, i_8_310_750_0, i_8_310_751_0, i_8_310_766_0,
    i_8_310_812_0, i_8_310_814_0, i_8_310_822_0, i_8_310_837_0,
    i_8_310_838_0, i_8_310_874_0, i_8_310_877_0, i_8_310_883_0,
    i_8_310_914_0, i_8_310_919_0, i_8_310_938_0, i_8_310_959_0,
    i_8_310_1036_0, i_8_310_1071_0, i_8_310_1072_0, i_8_310_1108_0,
    i_8_310_1129_0, i_8_310_1153_0, i_8_310_1198_0, i_8_310_1201_0,
    i_8_310_1237_0, i_8_310_1243_0, i_8_310_1260_0, i_8_310_1265_0,
    i_8_310_1266_0, i_8_310_1318_0, i_8_310_1327_0, i_8_310_1335_0,
    i_8_310_1338_0, i_8_310_1355_0, i_8_310_1381_0, i_8_310_1441_0,
    i_8_310_1462_0, i_8_310_1480_0, i_8_310_1524_0, i_8_310_1539_0,
    i_8_310_1544_0, i_8_310_1630_0, i_8_310_1646_0, i_8_310_1647_0,
    i_8_310_1651_0, i_8_310_1667_0, i_8_310_1676_0, i_8_310_1687_0,
    i_8_310_1701_0, i_8_310_1702_0, i_8_310_1707_0, i_8_310_1747_0,
    i_8_310_1749_0, i_8_310_1765_0, i_8_310_1796_0, i_8_310_1800_0,
    i_8_310_1855_0, i_8_310_1864_0, i_8_310_1868_0, i_8_310_1957_0,
    i_8_310_1989_0, i_8_310_1993_0, i_8_310_1996_0, i_8_310_2044_0,
    i_8_310_2106_0, i_8_310_2148_0, i_8_310_2154_0, i_8_310_2226_0,
    i_8_310_2245_0, i_8_310_2290_0, i_8_310_2298_0,
    o_8_310_0_0  );
  input  i_8_310_22_0, i_8_310_54_0, i_8_310_64_0, i_8_310_219_0,
    i_8_310_220_0, i_8_310_283_0, i_8_310_319_0, i_8_310_321_0,
    i_8_310_397_0, i_8_310_424_0, i_8_310_441_0, i_8_310_496_0,
    i_8_310_504_0, i_8_310_524_0, i_8_310_526_0, i_8_310_571_0,
    i_8_310_580_0, i_8_310_589_0, i_8_310_596_0, i_8_310_613_0,
    i_8_310_622_0, i_8_310_642_0, i_8_310_659_0, i_8_310_660_0,
    i_8_310_675_0, i_8_310_676_0, i_8_310_699_0, i_8_310_700_0,
    i_8_310_707_0, i_8_310_730_0, i_8_310_750_0, i_8_310_751_0,
    i_8_310_766_0, i_8_310_812_0, i_8_310_814_0, i_8_310_822_0,
    i_8_310_837_0, i_8_310_838_0, i_8_310_874_0, i_8_310_877_0,
    i_8_310_883_0, i_8_310_914_0, i_8_310_919_0, i_8_310_938_0,
    i_8_310_959_0, i_8_310_1036_0, i_8_310_1071_0, i_8_310_1072_0,
    i_8_310_1108_0, i_8_310_1129_0, i_8_310_1153_0, i_8_310_1198_0,
    i_8_310_1201_0, i_8_310_1237_0, i_8_310_1243_0, i_8_310_1260_0,
    i_8_310_1265_0, i_8_310_1266_0, i_8_310_1318_0, i_8_310_1327_0,
    i_8_310_1335_0, i_8_310_1338_0, i_8_310_1355_0, i_8_310_1381_0,
    i_8_310_1441_0, i_8_310_1462_0, i_8_310_1480_0, i_8_310_1524_0,
    i_8_310_1539_0, i_8_310_1544_0, i_8_310_1630_0, i_8_310_1646_0,
    i_8_310_1647_0, i_8_310_1651_0, i_8_310_1667_0, i_8_310_1676_0,
    i_8_310_1687_0, i_8_310_1701_0, i_8_310_1702_0, i_8_310_1707_0,
    i_8_310_1747_0, i_8_310_1749_0, i_8_310_1765_0, i_8_310_1796_0,
    i_8_310_1800_0, i_8_310_1855_0, i_8_310_1864_0, i_8_310_1868_0,
    i_8_310_1957_0, i_8_310_1989_0, i_8_310_1993_0, i_8_310_1996_0,
    i_8_310_2044_0, i_8_310_2106_0, i_8_310_2148_0, i_8_310_2154_0,
    i_8_310_2226_0, i_8_310_2245_0, i_8_310_2290_0, i_8_310_2298_0;
  output o_8_310_0_0;
  assign o_8_310_0_0 = 0;
endmodule



// Benchmark "kernel_8_311" written by ABC on Sun Jul 19 10:08:29 2020

module kernel_8_311 ( 
    i_8_311_4_0, i_8_311_76_0, i_8_311_77_0, i_8_311_104_0, i_8_311_121_0,
    i_8_311_130_0, i_8_311_263_0, i_8_311_356_0, i_8_311_360_0,
    i_8_311_427_0, i_8_311_445_0, i_8_311_455_0, i_8_311_496_0,
    i_8_311_497_0, i_8_311_517_0, i_8_311_526_0, i_8_311_551_0,
    i_8_311_554_0, i_8_311_572_0, i_8_311_597_0, i_8_311_609_0,
    i_8_311_611_0, i_8_311_612_0, i_8_311_647_0, i_8_311_656_0,
    i_8_311_661_0, i_8_311_680_0, i_8_311_707_0, i_8_311_749_0,
    i_8_311_751_0, i_8_311_828_0, i_8_311_832_0, i_8_311_836_0,
    i_8_311_837_0, i_8_311_840_0, i_8_311_845_0, i_8_311_850_0,
    i_8_311_913_0, i_8_311_958_0, i_8_311_963_0, i_8_311_1003_0,
    i_8_311_1108_0, i_8_311_1109_0, i_8_311_1111_0, i_8_311_1129_0,
    i_8_311_1130_0, i_8_311_1154_0, i_8_311_1156_0, i_8_311_1177_0,
    i_8_311_1229_0, i_8_311_1234_0, i_8_311_1270_0, i_8_311_1299_0,
    i_8_311_1318_0, i_8_311_1322_0, i_8_311_1325_0, i_8_311_1390_0,
    i_8_311_1391_0, i_8_311_1399_0, i_8_311_1455_0, i_8_311_1460_0,
    i_8_311_1470_0, i_8_311_1493_0, i_8_311_1498_0, i_8_311_1598_0,
    i_8_311_1634_0, i_8_311_1643_0, i_8_311_1652_0, i_8_311_1706_0,
    i_8_311_1747_0, i_8_311_1757_0, i_8_311_1784_0, i_8_311_1807_0,
    i_8_311_1818_0, i_8_311_1844_0, i_8_311_1846_0, i_8_311_1849_0,
    i_8_311_1930_0, i_8_311_1972_0, i_8_311_1992_0, i_8_311_1993_0,
    i_8_311_2040_0, i_8_311_2041_0, i_8_311_2044_0, i_8_311_2065_0,
    i_8_311_2123_0, i_8_311_2134_0, i_8_311_2141_0, i_8_311_2145_0,
    i_8_311_2147_0, i_8_311_2149_0, i_8_311_2150_0, i_8_311_2159_0,
    i_8_311_2174_0, i_8_311_2176_0, i_8_311_2183_0, i_8_311_2228_0,
    i_8_311_2231_0, i_8_311_2248_0, i_8_311_2273_0,
    o_8_311_0_0  );
  input  i_8_311_4_0, i_8_311_76_0, i_8_311_77_0, i_8_311_104_0,
    i_8_311_121_0, i_8_311_130_0, i_8_311_263_0, i_8_311_356_0,
    i_8_311_360_0, i_8_311_427_0, i_8_311_445_0, i_8_311_455_0,
    i_8_311_496_0, i_8_311_497_0, i_8_311_517_0, i_8_311_526_0,
    i_8_311_551_0, i_8_311_554_0, i_8_311_572_0, i_8_311_597_0,
    i_8_311_609_0, i_8_311_611_0, i_8_311_612_0, i_8_311_647_0,
    i_8_311_656_0, i_8_311_661_0, i_8_311_680_0, i_8_311_707_0,
    i_8_311_749_0, i_8_311_751_0, i_8_311_828_0, i_8_311_832_0,
    i_8_311_836_0, i_8_311_837_0, i_8_311_840_0, i_8_311_845_0,
    i_8_311_850_0, i_8_311_913_0, i_8_311_958_0, i_8_311_963_0,
    i_8_311_1003_0, i_8_311_1108_0, i_8_311_1109_0, i_8_311_1111_0,
    i_8_311_1129_0, i_8_311_1130_0, i_8_311_1154_0, i_8_311_1156_0,
    i_8_311_1177_0, i_8_311_1229_0, i_8_311_1234_0, i_8_311_1270_0,
    i_8_311_1299_0, i_8_311_1318_0, i_8_311_1322_0, i_8_311_1325_0,
    i_8_311_1390_0, i_8_311_1391_0, i_8_311_1399_0, i_8_311_1455_0,
    i_8_311_1460_0, i_8_311_1470_0, i_8_311_1493_0, i_8_311_1498_0,
    i_8_311_1598_0, i_8_311_1634_0, i_8_311_1643_0, i_8_311_1652_0,
    i_8_311_1706_0, i_8_311_1747_0, i_8_311_1757_0, i_8_311_1784_0,
    i_8_311_1807_0, i_8_311_1818_0, i_8_311_1844_0, i_8_311_1846_0,
    i_8_311_1849_0, i_8_311_1930_0, i_8_311_1972_0, i_8_311_1992_0,
    i_8_311_1993_0, i_8_311_2040_0, i_8_311_2041_0, i_8_311_2044_0,
    i_8_311_2065_0, i_8_311_2123_0, i_8_311_2134_0, i_8_311_2141_0,
    i_8_311_2145_0, i_8_311_2147_0, i_8_311_2149_0, i_8_311_2150_0,
    i_8_311_2159_0, i_8_311_2174_0, i_8_311_2176_0, i_8_311_2183_0,
    i_8_311_2228_0, i_8_311_2231_0, i_8_311_2248_0, i_8_311_2273_0;
  output o_8_311_0_0;
  assign o_8_311_0_0 = 0;
endmodule



// Benchmark "kernel_8_312" written by ABC on Sun Jul 19 10:08:30 2020

module kernel_8_312 ( 
    i_8_312_23_0, i_8_312_26_0, i_8_312_34_0, i_8_312_120_0, i_8_312_139_0,
    i_8_312_148_0, i_8_312_202_0, i_8_312_239_0, i_8_312_275_0,
    i_8_312_278_0, i_8_312_308_0, i_8_312_310_0, i_8_312_365_0,
    i_8_312_384_0, i_8_312_425_0, i_8_312_453_0, i_8_312_490_0,
    i_8_312_491_0, i_8_312_522_0, i_8_312_523_0, i_8_312_552_0,
    i_8_312_553_0, i_8_312_569_0, i_8_312_608_0, i_8_312_612_0,
    i_8_312_667_0, i_8_312_734_0, i_8_312_748_0, i_8_312_760_0,
    i_8_312_767_0, i_8_312_771_0, i_8_312_787_0, i_8_312_800_0,
    i_8_312_814_0, i_8_312_828_0, i_8_312_838_0, i_8_312_844_0,
    i_8_312_874_0, i_8_312_964_0, i_8_312_970_0, i_8_312_985_0,
    i_8_312_993_0, i_8_312_996_0, i_8_312_1021_0, i_8_312_1050_0,
    i_8_312_1067_0, i_8_312_1084_0, i_8_312_1102_0, i_8_312_1131_0,
    i_8_312_1135_0, i_8_312_1234_0, i_8_312_1238_0, i_8_312_1264_0,
    i_8_312_1267_0, i_8_312_1284_0, i_8_312_1305_0, i_8_312_1357_0,
    i_8_312_1381_0, i_8_312_1400_0, i_8_312_1408_0, i_8_312_1432_0,
    i_8_312_1437_0, i_8_312_1452_0, i_8_312_1508_0, i_8_312_1531_0,
    i_8_312_1544_0, i_8_312_1607_0, i_8_312_1643_0, i_8_312_1666_0,
    i_8_312_1667_0, i_8_312_1669_0, i_8_312_1671_0, i_8_312_1678_0,
    i_8_312_1747_0, i_8_312_1754_0, i_8_312_1757_0, i_8_312_1810_0,
    i_8_312_1822_0, i_8_312_1843_0, i_8_312_1883_0, i_8_312_1887_0,
    i_8_312_1927_0, i_8_312_1966_0, i_8_312_2000_0, i_8_312_2008_0,
    i_8_312_2009_0, i_8_312_2023_0, i_8_312_2070_0, i_8_312_2084_0,
    i_8_312_2143_0, i_8_312_2151_0, i_8_312_2153_0, i_8_312_2164_0,
    i_8_312_2165_0, i_8_312_2170_0, i_8_312_2176_0, i_8_312_2224_0,
    i_8_312_2245_0, i_8_312_2264_0, i_8_312_2273_0,
    o_8_312_0_0  );
  input  i_8_312_23_0, i_8_312_26_0, i_8_312_34_0, i_8_312_120_0,
    i_8_312_139_0, i_8_312_148_0, i_8_312_202_0, i_8_312_239_0,
    i_8_312_275_0, i_8_312_278_0, i_8_312_308_0, i_8_312_310_0,
    i_8_312_365_0, i_8_312_384_0, i_8_312_425_0, i_8_312_453_0,
    i_8_312_490_0, i_8_312_491_0, i_8_312_522_0, i_8_312_523_0,
    i_8_312_552_0, i_8_312_553_0, i_8_312_569_0, i_8_312_608_0,
    i_8_312_612_0, i_8_312_667_0, i_8_312_734_0, i_8_312_748_0,
    i_8_312_760_0, i_8_312_767_0, i_8_312_771_0, i_8_312_787_0,
    i_8_312_800_0, i_8_312_814_0, i_8_312_828_0, i_8_312_838_0,
    i_8_312_844_0, i_8_312_874_0, i_8_312_964_0, i_8_312_970_0,
    i_8_312_985_0, i_8_312_993_0, i_8_312_996_0, i_8_312_1021_0,
    i_8_312_1050_0, i_8_312_1067_0, i_8_312_1084_0, i_8_312_1102_0,
    i_8_312_1131_0, i_8_312_1135_0, i_8_312_1234_0, i_8_312_1238_0,
    i_8_312_1264_0, i_8_312_1267_0, i_8_312_1284_0, i_8_312_1305_0,
    i_8_312_1357_0, i_8_312_1381_0, i_8_312_1400_0, i_8_312_1408_0,
    i_8_312_1432_0, i_8_312_1437_0, i_8_312_1452_0, i_8_312_1508_0,
    i_8_312_1531_0, i_8_312_1544_0, i_8_312_1607_0, i_8_312_1643_0,
    i_8_312_1666_0, i_8_312_1667_0, i_8_312_1669_0, i_8_312_1671_0,
    i_8_312_1678_0, i_8_312_1747_0, i_8_312_1754_0, i_8_312_1757_0,
    i_8_312_1810_0, i_8_312_1822_0, i_8_312_1843_0, i_8_312_1883_0,
    i_8_312_1887_0, i_8_312_1927_0, i_8_312_1966_0, i_8_312_2000_0,
    i_8_312_2008_0, i_8_312_2009_0, i_8_312_2023_0, i_8_312_2070_0,
    i_8_312_2084_0, i_8_312_2143_0, i_8_312_2151_0, i_8_312_2153_0,
    i_8_312_2164_0, i_8_312_2165_0, i_8_312_2170_0, i_8_312_2176_0,
    i_8_312_2224_0, i_8_312_2245_0, i_8_312_2264_0, i_8_312_2273_0;
  output o_8_312_0_0;
  assign o_8_312_0_0 = 0;
endmodule



// Benchmark "kernel_8_313" written by ABC on Sun Jul 19 10:08:30 2020

module kernel_8_313 ( 
    i_8_313_18_0, i_8_313_41_0, i_8_313_59_0, i_8_313_88_0, i_8_313_115_0,
    i_8_313_143_0, i_8_313_188_0, i_8_313_234_0, i_8_313_266_0,
    i_8_313_283_0, i_8_313_284_0, i_8_313_361_0, i_8_313_362_0,
    i_8_313_379_0, i_8_313_383_0, i_8_313_481_0, i_8_313_493_0,
    i_8_313_524_0, i_8_313_525_0, i_8_313_554_0, i_8_313_569_0,
    i_8_313_610_0, i_8_313_635_0, i_8_313_679_0, i_8_313_682_0,
    i_8_313_693_0, i_8_313_698_0, i_8_313_704_0, i_8_313_709_0,
    i_8_313_724_0, i_8_313_735_0, i_8_313_754_0, i_8_313_762_0,
    i_8_313_771_0, i_8_313_773_0, i_8_313_787_0, i_8_313_789_0,
    i_8_313_799_0, i_8_313_841_0, i_8_313_958_0, i_8_313_964_0,
    i_8_313_970_0, i_8_313_1075_0, i_8_313_1106_0, i_8_313_1109_0,
    i_8_313_1256_0, i_8_313_1268_0, i_8_313_1301_0, i_8_313_1305_0,
    i_8_313_1351_0, i_8_313_1363_0, i_8_313_1399_0, i_8_313_1436_0,
    i_8_313_1455_0, i_8_313_1467_0, i_8_313_1471_0, i_8_313_1481_0,
    i_8_313_1489_0, i_8_313_1490_0, i_8_313_1529_0, i_8_313_1534_0,
    i_8_313_1606_0, i_8_313_1644_0, i_8_313_1649_0, i_8_313_1652_0,
    i_8_313_1670_0, i_8_313_1689_0, i_8_313_1703_0, i_8_313_1723_0,
    i_8_313_1725_0, i_8_313_1751_0, i_8_313_1752_0, i_8_313_1759_0,
    i_8_313_1765_0, i_8_313_1795_0, i_8_313_1804_0, i_8_313_1826_0,
    i_8_313_1838_0, i_8_313_1848_0, i_8_313_1849_0, i_8_313_1866_0,
    i_8_313_1867_0, i_8_313_1882_0, i_8_313_1886_0, i_8_313_1912_0,
    i_8_313_1919_0, i_8_313_1982_0, i_8_313_2001_0, i_8_313_2028_0,
    i_8_313_2075_0, i_8_313_2092_0, i_8_313_2142_0, i_8_313_2194_0,
    i_8_313_2224_0, i_8_313_2229_0, i_8_313_2230_0, i_8_313_2232_0,
    i_8_313_2242_0, i_8_313_2248_0, i_8_313_2264_0,
    o_8_313_0_0  );
  input  i_8_313_18_0, i_8_313_41_0, i_8_313_59_0, i_8_313_88_0,
    i_8_313_115_0, i_8_313_143_0, i_8_313_188_0, i_8_313_234_0,
    i_8_313_266_0, i_8_313_283_0, i_8_313_284_0, i_8_313_361_0,
    i_8_313_362_0, i_8_313_379_0, i_8_313_383_0, i_8_313_481_0,
    i_8_313_493_0, i_8_313_524_0, i_8_313_525_0, i_8_313_554_0,
    i_8_313_569_0, i_8_313_610_0, i_8_313_635_0, i_8_313_679_0,
    i_8_313_682_0, i_8_313_693_0, i_8_313_698_0, i_8_313_704_0,
    i_8_313_709_0, i_8_313_724_0, i_8_313_735_0, i_8_313_754_0,
    i_8_313_762_0, i_8_313_771_0, i_8_313_773_0, i_8_313_787_0,
    i_8_313_789_0, i_8_313_799_0, i_8_313_841_0, i_8_313_958_0,
    i_8_313_964_0, i_8_313_970_0, i_8_313_1075_0, i_8_313_1106_0,
    i_8_313_1109_0, i_8_313_1256_0, i_8_313_1268_0, i_8_313_1301_0,
    i_8_313_1305_0, i_8_313_1351_0, i_8_313_1363_0, i_8_313_1399_0,
    i_8_313_1436_0, i_8_313_1455_0, i_8_313_1467_0, i_8_313_1471_0,
    i_8_313_1481_0, i_8_313_1489_0, i_8_313_1490_0, i_8_313_1529_0,
    i_8_313_1534_0, i_8_313_1606_0, i_8_313_1644_0, i_8_313_1649_0,
    i_8_313_1652_0, i_8_313_1670_0, i_8_313_1689_0, i_8_313_1703_0,
    i_8_313_1723_0, i_8_313_1725_0, i_8_313_1751_0, i_8_313_1752_0,
    i_8_313_1759_0, i_8_313_1765_0, i_8_313_1795_0, i_8_313_1804_0,
    i_8_313_1826_0, i_8_313_1838_0, i_8_313_1848_0, i_8_313_1849_0,
    i_8_313_1866_0, i_8_313_1867_0, i_8_313_1882_0, i_8_313_1886_0,
    i_8_313_1912_0, i_8_313_1919_0, i_8_313_1982_0, i_8_313_2001_0,
    i_8_313_2028_0, i_8_313_2075_0, i_8_313_2092_0, i_8_313_2142_0,
    i_8_313_2194_0, i_8_313_2224_0, i_8_313_2229_0, i_8_313_2230_0,
    i_8_313_2232_0, i_8_313_2242_0, i_8_313_2248_0, i_8_313_2264_0;
  output o_8_313_0_0;
  assign o_8_313_0_0 = 0;
endmodule



// Benchmark "kernel_8_314" written by ABC on Sun Jul 19 10:08:31 2020

module kernel_8_314 ( 
    i_8_314_33_0, i_8_314_85_0, i_8_314_100_0, i_8_314_135_0,
    i_8_314_183_0, i_8_314_207_0, i_8_314_208_0, i_8_314_209_0,
    i_8_314_217_0, i_8_314_220_0, i_8_314_223_0, i_8_314_304_0,
    i_8_314_326_0, i_8_314_362_0, i_8_314_450_0, i_8_314_452_0,
    i_8_314_493_0, i_8_314_498_0, i_8_314_514_0, i_8_314_523_0,
    i_8_314_540_0, i_8_314_605_0, i_8_314_612_0, i_8_314_621_0,
    i_8_314_631_0, i_8_314_632_0, i_8_314_634_0, i_8_314_715_0,
    i_8_314_721_0, i_8_314_725_0, i_8_314_734_0, i_8_314_759_0,
    i_8_314_766_0, i_8_314_767_0, i_8_314_769_0, i_8_314_779_0,
    i_8_314_796_0, i_8_314_833_0, i_8_314_864_0, i_8_314_880_0,
    i_8_314_883_0, i_8_314_901_0, i_8_314_903_0, i_8_314_918_0,
    i_8_314_947_0, i_8_314_983_0, i_8_314_991_0, i_8_314_1031_0,
    i_8_314_1066_0, i_8_314_1072_0, i_8_314_1073_0, i_8_314_1172_0,
    i_8_314_1174_0, i_8_314_1246_0, i_8_314_1247_0, i_8_314_1256_0,
    i_8_314_1288_0, i_8_314_1324_0, i_8_314_1417_0, i_8_314_1538_0,
    i_8_314_1555_0, i_8_314_1556_0, i_8_314_1561_0, i_8_314_1565_0,
    i_8_314_1576_0, i_8_314_1606_0, i_8_314_1613_0, i_8_314_1665_0,
    i_8_314_1670_0, i_8_314_1675_0, i_8_314_1681_0, i_8_314_1684_0,
    i_8_314_1703_0, i_8_314_1710_0, i_8_314_1711_0, i_8_314_1712_0,
    i_8_314_1716_0, i_8_314_1721_0, i_8_314_1730_0, i_8_314_1746_0,
    i_8_314_1752_0, i_8_314_1783_0, i_8_314_1811_0, i_8_314_1819_0,
    i_8_314_1822_0, i_8_314_1823_0, i_8_314_1855_0, i_8_314_1963_0,
    i_8_314_1972_0, i_8_314_1999_0, i_8_314_2000_0, i_8_314_2107_0,
    i_8_314_2139_0, i_8_314_2144_0, i_8_314_2147_0, i_8_314_2215_0,
    i_8_314_2243_0, i_8_314_2255_0, i_8_314_2289_0, i_8_314_2293_0,
    o_8_314_0_0  );
  input  i_8_314_33_0, i_8_314_85_0, i_8_314_100_0, i_8_314_135_0,
    i_8_314_183_0, i_8_314_207_0, i_8_314_208_0, i_8_314_209_0,
    i_8_314_217_0, i_8_314_220_0, i_8_314_223_0, i_8_314_304_0,
    i_8_314_326_0, i_8_314_362_0, i_8_314_450_0, i_8_314_452_0,
    i_8_314_493_0, i_8_314_498_0, i_8_314_514_0, i_8_314_523_0,
    i_8_314_540_0, i_8_314_605_0, i_8_314_612_0, i_8_314_621_0,
    i_8_314_631_0, i_8_314_632_0, i_8_314_634_0, i_8_314_715_0,
    i_8_314_721_0, i_8_314_725_0, i_8_314_734_0, i_8_314_759_0,
    i_8_314_766_0, i_8_314_767_0, i_8_314_769_0, i_8_314_779_0,
    i_8_314_796_0, i_8_314_833_0, i_8_314_864_0, i_8_314_880_0,
    i_8_314_883_0, i_8_314_901_0, i_8_314_903_0, i_8_314_918_0,
    i_8_314_947_0, i_8_314_983_0, i_8_314_991_0, i_8_314_1031_0,
    i_8_314_1066_0, i_8_314_1072_0, i_8_314_1073_0, i_8_314_1172_0,
    i_8_314_1174_0, i_8_314_1246_0, i_8_314_1247_0, i_8_314_1256_0,
    i_8_314_1288_0, i_8_314_1324_0, i_8_314_1417_0, i_8_314_1538_0,
    i_8_314_1555_0, i_8_314_1556_0, i_8_314_1561_0, i_8_314_1565_0,
    i_8_314_1576_0, i_8_314_1606_0, i_8_314_1613_0, i_8_314_1665_0,
    i_8_314_1670_0, i_8_314_1675_0, i_8_314_1681_0, i_8_314_1684_0,
    i_8_314_1703_0, i_8_314_1710_0, i_8_314_1711_0, i_8_314_1712_0,
    i_8_314_1716_0, i_8_314_1721_0, i_8_314_1730_0, i_8_314_1746_0,
    i_8_314_1752_0, i_8_314_1783_0, i_8_314_1811_0, i_8_314_1819_0,
    i_8_314_1822_0, i_8_314_1823_0, i_8_314_1855_0, i_8_314_1963_0,
    i_8_314_1972_0, i_8_314_1999_0, i_8_314_2000_0, i_8_314_2107_0,
    i_8_314_2139_0, i_8_314_2144_0, i_8_314_2147_0, i_8_314_2215_0,
    i_8_314_2243_0, i_8_314_2255_0, i_8_314_2289_0, i_8_314_2293_0;
  output o_8_314_0_0;
  assign o_8_314_0_0 = 0;
endmodule



// Benchmark "kernel_8_315" written by ABC on Sun Jul 19 10:08:32 2020

module kernel_8_315 ( 
    i_8_315_10_0, i_8_315_38_0, i_8_315_49_0, i_8_315_82_0, i_8_315_93_0,
    i_8_315_111_0, i_8_315_181_0, i_8_315_216_0, i_8_315_217_0,
    i_8_315_315_0, i_8_315_316_0, i_8_315_317_0, i_8_315_324_0,
    i_8_315_325_0, i_8_315_360_0, i_8_315_397_0, i_8_315_416_0,
    i_8_315_505_0, i_8_315_522_0, i_8_315_523_0, i_8_315_550_0,
    i_8_315_576_0, i_8_315_577_0, i_8_315_595_0, i_8_315_603_0,
    i_8_315_604_0, i_8_315_640_0, i_8_315_653_0, i_8_315_659_0,
    i_8_315_667_0, i_8_315_706_0, i_8_315_730_0, i_8_315_731_0,
    i_8_315_748_0, i_8_315_799_0, i_8_315_841_0, i_8_315_874_0,
    i_8_315_1010_0, i_8_315_1036_0, i_8_315_1108_0, i_8_315_1135_0,
    i_8_315_1136_0, i_8_315_1153_0, i_8_315_1156_0, i_8_315_1233_0,
    i_8_315_1234_0, i_8_315_1243_0, i_8_315_1244_0, i_8_315_1260_0,
    i_8_315_1269_0, i_8_315_1278_0, i_8_315_1296_0, i_8_315_1297_0,
    i_8_315_1324_0, i_8_315_1333_0, i_8_315_1360_0, i_8_315_1363_0,
    i_8_315_1388_0, i_8_315_1407_0, i_8_315_1423_0, i_8_315_1431_0,
    i_8_315_1450_0, i_8_315_1455_0, i_8_315_1459_0, i_8_315_1462_0,
    i_8_315_1468_0, i_8_315_1470_0, i_8_315_1471_0, i_8_315_1476_0,
    i_8_315_1489_0, i_8_315_1512_0, i_8_315_1513_0, i_8_315_1522_0,
    i_8_315_1523_0, i_8_315_1544_0, i_8_315_1594_0, i_8_315_1604_0,
    i_8_315_1675_0, i_8_315_1684_0, i_8_315_1693_0, i_8_315_1710_0,
    i_8_315_1774_0, i_8_315_1822_0, i_8_315_1837_0, i_8_315_1881_0,
    i_8_315_1888_0, i_8_315_1936_0, i_8_315_1971_0, i_8_315_1972_0,
    i_8_315_1990_0, i_8_315_1992_0, i_8_315_2043_0, i_8_315_2104_0,
    i_8_315_2133_0, i_8_315_2169_0, i_8_315_2187_0, i_8_315_2259_0,
    i_8_315_2260_0, i_8_315_2287_0, i_8_315_2291_0,
    o_8_315_0_0  );
  input  i_8_315_10_0, i_8_315_38_0, i_8_315_49_0, i_8_315_82_0,
    i_8_315_93_0, i_8_315_111_0, i_8_315_181_0, i_8_315_216_0,
    i_8_315_217_0, i_8_315_315_0, i_8_315_316_0, i_8_315_317_0,
    i_8_315_324_0, i_8_315_325_0, i_8_315_360_0, i_8_315_397_0,
    i_8_315_416_0, i_8_315_505_0, i_8_315_522_0, i_8_315_523_0,
    i_8_315_550_0, i_8_315_576_0, i_8_315_577_0, i_8_315_595_0,
    i_8_315_603_0, i_8_315_604_0, i_8_315_640_0, i_8_315_653_0,
    i_8_315_659_0, i_8_315_667_0, i_8_315_706_0, i_8_315_730_0,
    i_8_315_731_0, i_8_315_748_0, i_8_315_799_0, i_8_315_841_0,
    i_8_315_874_0, i_8_315_1010_0, i_8_315_1036_0, i_8_315_1108_0,
    i_8_315_1135_0, i_8_315_1136_0, i_8_315_1153_0, i_8_315_1156_0,
    i_8_315_1233_0, i_8_315_1234_0, i_8_315_1243_0, i_8_315_1244_0,
    i_8_315_1260_0, i_8_315_1269_0, i_8_315_1278_0, i_8_315_1296_0,
    i_8_315_1297_0, i_8_315_1324_0, i_8_315_1333_0, i_8_315_1360_0,
    i_8_315_1363_0, i_8_315_1388_0, i_8_315_1407_0, i_8_315_1423_0,
    i_8_315_1431_0, i_8_315_1450_0, i_8_315_1455_0, i_8_315_1459_0,
    i_8_315_1462_0, i_8_315_1468_0, i_8_315_1470_0, i_8_315_1471_0,
    i_8_315_1476_0, i_8_315_1489_0, i_8_315_1512_0, i_8_315_1513_0,
    i_8_315_1522_0, i_8_315_1523_0, i_8_315_1544_0, i_8_315_1594_0,
    i_8_315_1604_0, i_8_315_1675_0, i_8_315_1684_0, i_8_315_1693_0,
    i_8_315_1710_0, i_8_315_1774_0, i_8_315_1822_0, i_8_315_1837_0,
    i_8_315_1881_0, i_8_315_1888_0, i_8_315_1936_0, i_8_315_1971_0,
    i_8_315_1972_0, i_8_315_1990_0, i_8_315_1992_0, i_8_315_2043_0,
    i_8_315_2104_0, i_8_315_2133_0, i_8_315_2169_0, i_8_315_2187_0,
    i_8_315_2259_0, i_8_315_2260_0, i_8_315_2287_0, i_8_315_2291_0;
  output o_8_315_0_0;
  assign o_8_315_0_0 = 0;
endmodule



// Benchmark "kernel_8_316" written by ABC on Sun Jul 19 10:08:33 2020

module kernel_8_316 ( 
    i_8_316_30_0, i_8_316_31_0, i_8_316_37_0, i_8_316_82_0, i_8_316_84_0,
    i_8_316_114_0, i_8_316_115_0, i_8_316_128_0, i_8_316_136_0,
    i_8_316_143_0, i_8_316_150_0, i_8_316_194_0, i_8_316_247_0,
    i_8_316_382_0, i_8_316_383_0, i_8_316_386_0, i_8_316_389_0,
    i_8_316_391_0, i_8_316_398_0, i_8_316_419_0, i_8_316_433_0,
    i_8_316_491_0, i_8_316_496_0, i_8_316_497_0, i_8_316_517_0,
    i_8_316_556_0, i_8_316_605_0, i_8_316_607_0, i_8_316_614_0,
    i_8_316_631_0, i_8_316_634_0, i_8_316_638_0, i_8_316_661_0,
    i_8_316_747_0, i_8_316_786_0, i_8_316_842_0, i_8_316_850_0,
    i_8_316_858_0, i_8_316_931_0, i_8_316_940_0, i_8_316_959_0,
    i_8_316_964_0, i_8_316_1072_0, i_8_316_1082_0, i_8_316_1125_0,
    i_8_316_1135_0, i_8_316_1228_0, i_8_316_1237_0, i_8_316_1262_0,
    i_8_316_1264_0, i_8_316_1274_0, i_8_316_1304_0, i_8_316_1309_0,
    i_8_316_1355_0, i_8_316_1388_0, i_8_316_1400_0, i_8_316_1434_0,
    i_8_316_1435_0, i_8_316_1462_0, i_8_316_1509_0, i_8_316_1522_0,
    i_8_316_1525_0, i_8_316_1531_0, i_8_316_1642_0, i_8_316_1647_0,
    i_8_316_1667_0, i_8_316_1675_0, i_8_316_1697_0, i_8_316_1702_0,
    i_8_316_1717_0, i_8_316_1747_0, i_8_316_1760_0, i_8_316_1766_0,
    i_8_316_1792_0, i_8_316_1805_0, i_8_316_1808_0, i_8_316_1823_0,
    i_8_316_1826_0, i_8_316_1865_0, i_8_316_1866_0, i_8_316_1918_0,
    i_8_316_1948_0, i_8_316_1972_0, i_8_316_1997_0, i_8_316_2060_0,
    i_8_316_2110_0, i_8_316_2134_0, i_8_316_2138_0, i_8_316_2141_0,
    i_8_316_2144_0, i_8_316_2154_0, i_8_316_2155_0, i_8_316_2170_0,
    i_8_316_2209_0, i_8_316_2215_0, i_8_316_2218_0, i_8_316_2255_0,
    i_8_316_2281_0, i_8_316_2286_0, i_8_316_2298_0,
    o_8_316_0_0  );
  input  i_8_316_30_0, i_8_316_31_0, i_8_316_37_0, i_8_316_82_0,
    i_8_316_84_0, i_8_316_114_0, i_8_316_115_0, i_8_316_128_0,
    i_8_316_136_0, i_8_316_143_0, i_8_316_150_0, i_8_316_194_0,
    i_8_316_247_0, i_8_316_382_0, i_8_316_383_0, i_8_316_386_0,
    i_8_316_389_0, i_8_316_391_0, i_8_316_398_0, i_8_316_419_0,
    i_8_316_433_0, i_8_316_491_0, i_8_316_496_0, i_8_316_497_0,
    i_8_316_517_0, i_8_316_556_0, i_8_316_605_0, i_8_316_607_0,
    i_8_316_614_0, i_8_316_631_0, i_8_316_634_0, i_8_316_638_0,
    i_8_316_661_0, i_8_316_747_0, i_8_316_786_0, i_8_316_842_0,
    i_8_316_850_0, i_8_316_858_0, i_8_316_931_0, i_8_316_940_0,
    i_8_316_959_0, i_8_316_964_0, i_8_316_1072_0, i_8_316_1082_0,
    i_8_316_1125_0, i_8_316_1135_0, i_8_316_1228_0, i_8_316_1237_0,
    i_8_316_1262_0, i_8_316_1264_0, i_8_316_1274_0, i_8_316_1304_0,
    i_8_316_1309_0, i_8_316_1355_0, i_8_316_1388_0, i_8_316_1400_0,
    i_8_316_1434_0, i_8_316_1435_0, i_8_316_1462_0, i_8_316_1509_0,
    i_8_316_1522_0, i_8_316_1525_0, i_8_316_1531_0, i_8_316_1642_0,
    i_8_316_1647_0, i_8_316_1667_0, i_8_316_1675_0, i_8_316_1697_0,
    i_8_316_1702_0, i_8_316_1717_0, i_8_316_1747_0, i_8_316_1760_0,
    i_8_316_1766_0, i_8_316_1792_0, i_8_316_1805_0, i_8_316_1808_0,
    i_8_316_1823_0, i_8_316_1826_0, i_8_316_1865_0, i_8_316_1866_0,
    i_8_316_1918_0, i_8_316_1948_0, i_8_316_1972_0, i_8_316_1997_0,
    i_8_316_2060_0, i_8_316_2110_0, i_8_316_2134_0, i_8_316_2138_0,
    i_8_316_2141_0, i_8_316_2144_0, i_8_316_2154_0, i_8_316_2155_0,
    i_8_316_2170_0, i_8_316_2209_0, i_8_316_2215_0, i_8_316_2218_0,
    i_8_316_2255_0, i_8_316_2281_0, i_8_316_2286_0, i_8_316_2298_0;
  output o_8_316_0_0;
  assign o_8_316_0_0 = 0;
endmodule



// Benchmark "kernel_8_317" written by ABC on Sun Jul 19 10:08:34 2020

module kernel_8_317 ( 
    i_8_317_22_0, i_8_317_165_0, i_8_317_208_0, i_8_317_262_0,
    i_8_317_264_0, i_8_317_265_0, i_8_317_279_0, i_8_317_282_0,
    i_8_317_285_0, i_8_317_292_0, i_8_317_295_0, i_8_317_310_0,
    i_8_317_319_0, i_8_317_321_0, i_8_317_397_0, i_8_317_436_0,
    i_8_317_439_0, i_8_317_450_0, i_8_317_525_0, i_8_317_526_0,
    i_8_317_639_0, i_8_317_706_0, i_8_317_727_0, i_8_317_747_0,
    i_8_317_807_0, i_8_317_808_0, i_8_317_883_0, i_8_317_966_0,
    i_8_317_969_0, i_8_317_1035_0, i_8_317_1182_0, i_8_317_1191_0,
    i_8_317_1198_0, i_8_317_1227_0, i_8_317_1236_0, i_8_317_1264_0,
    i_8_317_1267_0, i_8_317_1290_0, i_8_317_1305_0, i_8_317_1310_0,
    i_8_317_1351_0, i_8_317_1354_0, i_8_317_1357_0, i_8_317_1359_0,
    i_8_317_1362_0, i_8_317_1365_0, i_8_317_1398_0, i_8_317_1440_0,
    i_8_317_1446_0, i_8_317_1456_0, i_8_317_1468_0, i_8_317_1470_0,
    i_8_317_1474_0, i_8_317_1489_0, i_8_317_1491_0, i_8_317_1524_0,
    i_8_317_1533_0, i_8_317_1536_0, i_8_317_1547_0, i_8_317_1560_0,
    i_8_317_1570_0, i_8_317_1627_0, i_8_317_1641_0, i_8_317_1645_0,
    i_8_317_1649_0, i_8_317_1674_0, i_8_317_1677_0, i_8_317_1678_0,
    i_8_317_1695_0, i_8_317_1696_0, i_8_317_1704_0, i_8_317_1713_0,
    i_8_317_1767_0, i_8_317_1780_0, i_8_317_1789_0, i_8_317_1791_0,
    i_8_317_1820_0, i_8_317_1822_0, i_8_317_1826_0, i_8_317_1836_0,
    i_8_317_1861_0, i_8_317_1876_0, i_8_317_1956_0, i_8_317_1987_0,
    i_8_317_1995_0, i_8_317_2028_0, i_8_317_2056_0, i_8_317_2112_0,
    i_8_317_2133_0, i_8_317_2136_0, i_8_317_2149_0, i_8_317_2154_0,
    i_8_317_2164_0, i_8_317_2172_0, i_8_317_2190_0, i_8_317_2193_0,
    i_8_317_2194_0, i_8_317_2228_0, i_8_317_2248_0, i_8_317_2260_0,
    o_8_317_0_0  );
  input  i_8_317_22_0, i_8_317_165_0, i_8_317_208_0, i_8_317_262_0,
    i_8_317_264_0, i_8_317_265_0, i_8_317_279_0, i_8_317_282_0,
    i_8_317_285_0, i_8_317_292_0, i_8_317_295_0, i_8_317_310_0,
    i_8_317_319_0, i_8_317_321_0, i_8_317_397_0, i_8_317_436_0,
    i_8_317_439_0, i_8_317_450_0, i_8_317_525_0, i_8_317_526_0,
    i_8_317_639_0, i_8_317_706_0, i_8_317_727_0, i_8_317_747_0,
    i_8_317_807_0, i_8_317_808_0, i_8_317_883_0, i_8_317_966_0,
    i_8_317_969_0, i_8_317_1035_0, i_8_317_1182_0, i_8_317_1191_0,
    i_8_317_1198_0, i_8_317_1227_0, i_8_317_1236_0, i_8_317_1264_0,
    i_8_317_1267_0, i_8_317_1290_0, i_8_317_1305_0, i_8_317_1310_0,
    i_8_317_1351_0, i_8_317_1354_0, i_8_317_1357_0, i_8_317_1359_0,
    i_8_317_1362_0, i_8_317_1365_0, i_8_317_1398_0, i_8_317_1440_0,
    i_8_317_1446_0, i_8_317_1456_0, i_8_317_1468_0, i_8_317_1470_0,
    i_8_317_1474_0, i_8_317_1489_0, i_8_317_1491_0, i_8_317_1524_0,
    i_8_317_1533_0, i_8_317_1536_0, i_8_317_1547_0, i_8_317_1560_0,
    i_8_317_1570_0, i_8_317_1627_0, i_8_317_1641_0, i_8_317_1645_0,
    i_8_317_1649_0, i_8_317_1674_0, i_8_317_1677_0, i_8_317_1678_0,
    i_8_317_1695_0, i_8_317_1696_0, i_8_317_1704_0, i_8_317_1713_0,
    i_8_317_1767_0, i_8_317_1780_0, i_8_317_1789_0, i_8_317_1791_0,
    i_8_317_1820_0, i_8_317_1822_0, i_8_317_1826_0, i_8_317_1836_0,
    i_8_317_1861_0, i_8_317_1876_0, i_8_317_1956_0, i_8_317_1987_0,
    i_8_317_1995_0, i_8_317_2028_0, i_8_317_2056_0, i_8_317_2112_0,
    i_8_317_2133_0, i_8_317_2136_0, i_8_317_2149_0, i_8_317_2154_0,
    i_8_317_2164_0, i_8_317_2172_0, i_8_317_2190_0, i_8_317_2193_0,
    i_8_317_2194_0, i_8_317_2228_0, i_8_317_2248_0, i_8_317_2260_0;
  output o_8_317_0_0;
  assign o_8_317_0_0 = ~((~i_8_317_285_0 & ((~i_8_317_808_0 & ((~i_8_317_264_0 & ~i_8_317_1359_0 & ((~i_8_317_319_0 & ~i_8_317_747_0 & ~i_8_317_1362_0 & ~i_8_317_1446_0 & ~i_8_317_1570_0 & ~i_8_317_1695_0) | (~i_8_317_165_0 & ~i_8_317_265_0 & ~i_8_317_439_0 & ~i_8_317_1365_0 & ~i_8_317_1696_0))) | (i_8_317_525_0 & ~i_8_317_639_0 & ~i_8_317_1570_0))) | (~i_8_317_1440_0 & ((~i_8_317_265_0 & ~i_8_317_279_0 & ~i_8_317_282_0 & ~i_8_317_436_0 & ~i_8_317_439_0 & ~i_8_317_727_0 & ~i_8_317_807_0 & ~i_8_317_1198_0 & ~i_8_317_2194_0) | (~i_8_317_1035_0 & ~i_8_317_1357_0 & ~i_8_317_1696_0 & ~i_8_317_1956_0 & ~i_8_317_2190_0 & ~i_8_317_2193_0 & ~i_8_317_2248_0))))) | (~i_8_317_279_0 & ((~i_8_317_319_0 & i_8_317_706_0 & ~i_8_317_1236_0 & ~i_8_317_1305_0 & i_8_317_2133_0) | (~i_8_317_292_0 & ~i_8_317_397_0 & ~i_8_317_969_0 & ~i_8_317_1440_0 & ~i_8_317_1704_0 & ~i_8_317_1995_0 & ~i_8_317_2154_0))) | (~i_8_317_319_0 & ~i_8_317_1446_0 & ((~i_8_317_807_0 & ~i_8_317_883_0 & ~i_8_317_1035_0 & ~i_8_317_1649_0 & ~i_8_317_1713_0 & ~i_8_317_2028_0 & i_8_317_2172_0) | (~i_8_317_1359_0 & ~i_8_317_1456_0 & ~i_8_317_1627_0 & ~i_8_317_1695_0 & ~i_8_317_1696_0 & ~i_8_317_1704_0 & ~i_8_317_1791_0 & ~i_8_317_2248_0))) | (~i_8_317_321_0 & ((~i_8_317_727_0 & i_8_317_808_0 & ~i_8_317_1456_0 & ~i_8_317_1570_0 & ~i_8_317_1822_0 & ~i_8_317_2028_0 & ~i_8_317_2136_0) | (~i_8_317_397_0 & i_8_317_706_0 & ~i_8_317_1182_0 & ~i_8_317_1267_0 & ~i_8_317_1359_0 & ~i_8_317_1536_0 & ~i_8_317_1627_0 & ~i_8_317_2154_0))) | (~i_8_317_439_0 & ((~i_8_317_706_0 & ~i_8_317_883_0 & ~i_8_317_966_0 & ~i_8_317_1357_0) | (~i_8_317_1182_0 & ~i_8_317_1524_0 & ~i_8_317_1570_0 & i_8_317_1780_0 & ~i_8_317_2149_0 & ~i_8_317_2172_0))) | (~i_8_317_1357_0 & ~i_8_317_1820_0 & ((~i_8_317_208_0 & ~i_8_317_262_0 & ~i_8_317_969_0 & ~i_8_317_1362_0 & ~i_8_317_1791_0 & ~i_8_317_1995_0) | (~i_8_317_282_0 & i_8_317_1440_0 & ~i_8_317_1491_0 & ~i_8_317_1956_0 & ~i_8_317_2190_0 & ~i_8_317_1524_0 & ~i_8_317_1674_0))) | (~i_8_317_1696_0 & (i_8_317_1474_0 | (~i_8_317_292_0 & ~i_8_317_397_0 & i_8_317_706_0 & i_8_317_1267_0 & ~i_8_317_1956_0 & ~i_8_317_2194_0))) | (i_8_317_310_0 & ~i_8_317_2136_0 & ~i_8_317_2194_0) | (~i_8_317_264_0 & ~i_8_317_436_0 & ~i_8_317_727_0 & ~i_8_317_807_0 & ~i_8_317_1264_0 & ~i_8_317_1354_0 & ~i_8_317_1704_0 & ~i_8_317_2028_0 & ~i_8_317_2190_0));
endmodule



// Benchmark "kernel_8_318" written by ABC on Sun Jul 19 10:08:35 2020

module kernel_8_318 ( 
    i_8_318_27_0, i_8_318_33_0, i_8_318_34_0, i_8_318_54_0, i_8_318_84_0,
    i_8_318_96_0, i_8_318_106_0, i_8_318_156_0, i_8_318_157_0,
    i_8_318_201_0, i_8_318_202_0, i_8_318_219_0, i_8_318_246_0,
    i_8_318_265_0, i_8_318_274_0, i_8_318_292_0, i_8_318_324_0,
    i_8_318_325_0, i_8_318_360_0, i_8_318_383_0, i_8_318_440_0,
    i_8_318_445_0, i_8_318_475_0, i_8_318_484_0, i_8_318_498_0,
    i_8_318_508_0, i_8_318_523_0, i_8_318_546_0, i_8_318_552_0,
    i_8_318_556_0, i_8_318_591_0, i_8_318_606_0, i_8_318_625_0,
    i_8_318_627_0, i_8_318_657_0, i_8_318_658_0, i_8_318_660_0,
    i_8_318_661_0, i_8_318_676_0, i_8_318_714_0, i_8_318_723_0,
    i_8_318_757_0, i_8_318_759_0, i_8_318_760_0, i_8_318_768_0,
    i_8_318_795_0, i_8_318_822_0, i_8_318_823_0, i_8_318_837_0,
    i_8_318_840_0, i_8_318_895_0, i_8_318_949_0, i_8_318_1050_0,
    i_8_318_1087_0, i_8_318_1107_0, i_8_318_1113_0, i_8_318_1114_0,
    i_8_318_1130_0, i_8_318_1134_0, i_8_318_1135_0, i_8_318_1155_0,
    i_8_318_1267_0, i_8_318_1305_0, i_8_318_1320_0, i_8_318_1346_0,
    i_8_318_1387_0, i_8_318_1408_0, i_8_318_1420_0, i_8_318_1470_0,
    i_8_318_1480_0, i_8_318_1524_0, i_8_318_1525_0, i_8_318_1551_0,
    i_8_318_1579_0, i_8_318_1589_0, i_8_318_1606_0, i_8_318_1629_0,
    i_8_318_1705_0, i_8_318_1716_0, i_8_318_1746_0, i_8_318_1781_0,
    i_8_318_1805_0, i_8_318_1809_0, i_8_318_1839_0, i_8_318_1858_0,
    i_8_318_1859_0, i_8_318_1902_0, i_8_318_1966_0, i_8_318_2001_0,
    i_8_318_2011_0, i_8_318_2028_0, i_8_318_2031_0, i_8_318_2043_0,
    i_8_318_2049_0, i_8_318_2127_0, i_8_318_2146_0, i_8_318_2187_0,
    i_8_318_2188_0, i_8_318_2263_0, i_8_318_2286_0,
    o_8_318_0_0  );
  input  i_8_318_27_0, i_8_318_33_0, i_8_318_34_0, i_8_318_54_0,
    i_8_318_84_0, i_8_318_96_0, i_8_318_106_0, i_8_318_156_0,
    i_8_318_157_0, i_8_318_201_0, i_8_318_202_0, i_8_318_219_0,
    i_8_318_246_0, i_8_318_265_0, i_8_318_274_0, i_8_318_292_0,
    i_8_318_324_0, i_8_318_325_0, i_8_318_360_0, i_8_318_383_0,
    i_8_318_440_0, i_8_318_445_0, i_8_318_475_0, i_8_318_484_0,
    i_8_318_498_0, i_8_318_508_0, i_8_318_523_0, i_8_318_546_0,
    i_8_318_552_0, i_8_318_556_0, i_8_318_591_0, i_8_318_606_0,
    i_8_318_625_0, i_8_318_627_0, i_8_318_657_0, i_8_318_658_0,
    i_8_318_660_0, i_8_318_661_0, i_8_318_676_0, i_8_318_714_0,
    i_8_318_723_0, i_8_318_757_0, i_8_318_759_0, i_8_318_760_0,
    i_8_318_768_0, i_8_318_795_0, i_8_318_822_0, i_8_318_823_0,
    i_8_318_837_0, i_8_318_840_0, i_8_318_895_0, i_8_318_949_0,
    i_8_318_1050_0, i_8_318_1087_0, i_8_318_1107_0, i_8_318_1113_0,
    i_8_318_1114_0, i_8_318_1130_0, i_8_318_1134_0, i_8_318_1135_0,
    i_8_318_1155_0, i_8_318_1267_0, i_8_318_1305_0, i_8_318_1320_0,
    i_8_318_1346_0, i_8_318_1387_0, i_8_318_1408_0, i_8_318_1420_0,
    i_8_318_1470_0, i_8_318_1480_0, i_8_318_1524_0, i_8_318_1525_0,
    i_8_318_1551_0, i_8_318_1579_0, i_8_318_1589_0, i_8_318_1606_0,
    i_8_318_1629_0, i_8_318_1705_0, i_8_318_1716_0, i_8_318_1746_0,
    i_8_318_1781_0, i_8_318_1805_0, i_8_318_1809_0, i_8_318_1839_0,
    i_8_318_1858_0, i_8_318_1859_0, i_8_318_1902_0, i_8_318_1966_0,
    i_8_318_2001_0, i_8_318_2011_0, i_8_318_2028_0, i_8_318_2031_0,
    i_8_318_2043_0, i_8_318_2049_0, i_8_318_2127_0, i_8_318_2146_0,
    i_8_318_2187_0, i_8_318_2188_0, i_8_318_2263_0, i_8_318_2286_0;
  output o_8_318_0_0;
  assign o_8_318_0_0 = 0;
endmodule



// Benchmark "kernel_8_319" written by ABC on Sun Jul 19 10:08:36 2020

module kernel_8_319 ( 
    i_8_319_34_0, i_8_319_80_0, i_8_319_85_0, i_8_319_125_0, i_8_319_139_0,
    i_8_319_142_0, i_8_319_151_0, i_8_319_194_0, i_8_319_197_0,
    i_8_319_230_0, i_8_319_365_0, i_8_319_373_0, i_8_319_427_0,
    i_8_319_430_0, i_8_319_454_0, i_8_319_490_0, i_8_319_491_0,
    i_8_319_538_0, i_8_319_556_0, i_8_319_584_0, i_8_319_605_0,
    i_8_319_616_0, i_8_319_628_0, i_8_319_629_0, i_8_319_662_0,
    i_8_319_665_0, i_8_319_677_0, i_8_319_694_0, i_8_319_696_0,
    i_8_319_697_0, i_8_319_698_0, i_8_319_725_0, i_8_319_731_0,
    i_8_319_736_0, i_8_319_755_0, i_8_319_782_0, i_8_319_784_0,
    i_8_319_808_0, i_8_319_838_0, i_8_319_842_0, i_8_319_843_0,
    i_8_319_844_0, i_8_319_845_0, i_8_319_869_0, i_8_319_952_0,
    i_8_319_989_0, i_8_319_995_0, i_8_319_1139_0, i_8_319_1142_0,
    i_8_319_1151_0, i_8_319_1241_0, i_8_319_1260_0, i_8_319_1283_0,
    i_8_319_1301_0, i_8_319_1331_0, i_8_319_1355_0, i_8_319_1376_0,
    i_8_319_1388_0, i_8_319_1411_0, i_8_319_1412_0, i_8_319_1450_0,
    i_8_319_1472_0, i_8_319_1483_0, i_8_319_1484_0, i_8_319_1529_0,
    i_8_319_1615_0, i_8_319_1664_0, i_8_319_1691_0, i_8_319_1701_0,
    i_8_319_1709_0, i_8_319_1732_0, i_8_319_1751_0, i_8_319_1771_0,
    i_8_319_1823_0, i_8_319_1825_0, i_8_319_1846_0, i_8_319_1858_0,
    i_8_319_1859_0, i_8_319_1886_0, i_8_319_1904_0, i_8_319_1961_0,
    i_8_319_1966_0, i_8_319_1990_0, i_8_319_1997_0, i_8_319_2012_0,
    i_8_319_2015_0, i_8_319_2060_0, i_8_319_2075_0, i_8_319_2087_0,
    i_8_319_2096_0, i_8_319_2129_0, i_8_319_2148_0, i_8_319_2153_0,
    i_8_319_2174_0, i_8_319_2176_0, i_8_319_2177_0, i_8_319_2236_0,
    i_8_319_2263_0, i_8_319_2275_0, i_8_319_2289_0,
    o_8_319_0_0  );
  input  i_8_319_34_0, i_8_319_80_0, i_8_319_85_0, i_8_319_125_0,
    i_8_319_139_0, i_8_319_142_0, i_8_319_151_0, i_8_319_194_0,
    i_8_319_197_0, i_8_319_230_0, i_8_319_365_0, i_8_319_373_0,
    i_8_319_427_0, i_8_319_430_0, i_8_319_454_0, i_8_319_490_0,
    i_8_319_491_0, i_8_319_538_0, i_8_319_556_0, i_8_319_584_0,
    i_8_319_605_0, i_8_319_616_0, i_8_319_628_0, i_8_319_629_0,
    i_8_319_662_0, i_8_319_665_0, i_8_319_677_0, i_8_319_694_0,
    i_8_319_696_0, i_8_319_697_0, i_8_319_698_0, i_8_319_725_0,
    i_8_319_731_0, i_8_319_736_0, i_8_319_755_0, i_8_319_782_0,
    i_8_319_784_0, i_8_319_808_0, i_8_319_838_0, i_8_319_842_0,
    i_8_319_843_0, i_8_319_844_0, i_8_319_845_0, i_8_319_869_0,
    i_8_319_952_0, i_8_319_989_0, i_8_319_995_0, i_8_319_1139_0,
    i_8_319_1142_0, i_8_319_1151_0, i_8_319_1241_0, i_8_319_1260_0,
    i_8_319_1283_0, i_8_319_1301_0, i_8_319_1331_0, i_8_319_1355_0,
    i_8_319_1376_0, i_8_319_1388_0, i_8_319_1411_0, i_8_319_1412_0,
    i_8_319_1450_0, i_8_319_1472_0, i_8_319_1483_0, i_8_319_1484_0,
    i_8_319_1529_0, i_8_319_1615_0, i_8_319_1664_0, i_8_319_1691_0,
    i_8_319_1701_0, i_8_319_1709_0, i_8_319_1732_0, i_8_319_1751_0,
    i_8_319_1771_0, i_8_319_1823_0, i_8_319_1825_0, i_8_319_1846_0,
    i_8_319_1858_0, i_8_319_1859_0, i_8_319_1886_0, i_8_319_1904_0,
    i_8_319_1961_0, i_8_319_1966_0, i_8_319_1990_0, i_8_319_1997_0,
    i_8_319_2012_0, i_8_319_2015_0, i_8_319_2060_0, i_8_319_2075_0,
    i_8_319_2087_0, i_8_319_2096_0, i_8_319_2129_0, i_8_319_2148_0,
    i_8_319_2153_0, i_8_319_2174_0, i_8_319_2176_0, i_8_319_2177_0,
    i_8_319_2236_0, i_8_319_2263_0, i_8_319_2275_0, i_8_319_2289_0;
  output o_8_319_0_0;
  assign o_8_319_0_0 = 0;
endmodule



// Benchmark "kernel_8_320" written by ABC on Sun Jul 19 10:08:37 2020

module kernel_8_320 ( 
    i_8_320_31_0, i_8_320_50_0, i_8_320_57_0, i_8_320_60_0, i_8_320_75_0,
    i_8_320_101_0, i_8_320_131_0, i_8_320_168_0, i_8_320_190_0,
    i_8_320_301_0, i_8_320_311_0, i_8_320_322_0, i_8_320_356_0,
    i_8_320_361_0, i_8_320_371_0, i_8_320_384_0, i_8_320_427_0,
    i_8_320_455_0, i_8_320_461_0, i_8_320_538_0, i_8_320_539_0,
    i_8_320_548_0, i_8_320_553_0, i_8_320_581_0, i_8_320_582_0,
    i_8_320_608_0, i_8_320_613_0, i_8_320_638_0, i_8_320_644_0,
    i_8_320_653_0, i_8_320_655_0, i_8_320_664_0, i_8_320_683_0,
    i_8_320_695_0, i_8_320_701_0, i_8_320_745_0, i_8_320_752_0,
    i_8_320_755_0, i_8_320_779_0, i_8_320_781_0, i_8_320_820_0,
    i_8_320_827_0, i_8_320_884_0, i_8_320_886_0, i_8_320_944_0,
    i_8_320_955_0, i_8_320_1006_0, i_8_320_1039_0, i_8_320_1127_0,
    i_8_320_1226_0, i_8_320_1246_0, i_8_320_1247_0, i_8_320_1267_0,
    i_8_320_1268_0, i_8_320_1282_0, i_8_320_1283_0, i_8_320_1301_0,
    i_8_320_1302_0, i_8_320_1303_0, i_8_320_1339_0, i_8_320_1350_0,
    i_8_320_1353_0, i_8_320_1432_0, i_8_320_1455_0, i_8_320_1603_0,
    i_8_320_1607_0, i_8_320_1608_0, i_8_320_1633_0, i_8_320_1668_0,
    i_8_320_1699_0, i_8_320_1709_0, i_8_320_1718_0, i_8_320_1737_0,
    i_8_320_1759_0, i_8_320_1768_0, i_8_320_1777_0, i_8_320_1780_0,
    i_8_320_1789_0, i_8_320_1807_0, i_8_320_1810_0, i_8_320_1903_0,
    i_8_320_1904_0, i_8_320_1912_0, i_8_320_1939_0, i_8_320_1973_0,
    i_8_320_1981_0, i_8_320_1984_0, i_8_320_1992_0, i_8_320_2039_0,
    i_8_320_2048_0, i_8_320_2107_0, i_8_320_2145_0, i_8_320_2155_0,
    i_8_320_2156_0, i_8_320_2173_0, i_8_320_2195_0, i_8_320_2249_0,
    i_8_320_2270_0, i_8_320_2290_0, i_8_320_2294_0,
    o_8_320_0_0  );
  input  i_8_320_31_0, i_8_320_50_0, i_8_320_57_0, i_8_320_60_0,
    i_8_320_75_0, i_8_320_101_0, i_8_320_131_0, i_8_320_168_0,
    i_8_320_190_0, i_8_320_301_0, i_8_320_311_0, i_8_320_322_0,
    i_8_320_356_0, i_8_320_361_0, i_8_320_371_0, i_8_320_384_0,
    i_8_320_427_0, i_8_320_455_0, i_8_320_461_0, i_8_320_538_0,
    i_8_320_539_0, i_8_320_548_0, i_8_320_553_0, i_8_320_581_0,
    i_8_320_582_0, i_8_320_608_0, i_8_320_613_0, i_8_320_638_0,
    i_8_320_644_0, i_8_320_653_0, i_8_320_655_0, i_8_320_664_0,
    i_8_320_683_0, i_8_320_695_0, i_8_320_701_0, i_8_320_745_0,
    i_8_320_752_0, i_8_320_755_0, i_8_320_779_0, i_8_320_781_0,
    i_8_320_820_0, i_8_320_827_0, i_8_320_884_0, i_8_320_886_0,
    i_8_320_944_0, i_8_320_955_0, i_8_320_1006_0, i_8_320_1039_0,
    i_8_320_1127_0, i_8_320_1226_0, i_8_320_1246_0, i_8_320_1247_0,
    i_8_320_1267_0, i_8_320_1268_0, i_8_320_1282_0, i_8_320_1283_0,
    i_8_320_1301_0, i_8_320_1302_0, i_8_320_1303_0, i_8_320_1339_0,
    i_8_320_1350_0, i_8_320_1353_0, i_8_320_1432_0, i_8_320_1455_0,
    i_8_320_1603_0, i_8_320_1607_0, i_8_320_1608_0, i_8_320_1633_0,
    i_8_320_1668_0, i_8_320_1699_0, i_8_320_1709_0, i_8_320_1718_0,
    i_8_320_1737_0, i_8_320_1759_0, i_8_320_1768_0, i_8_320_1777_0,
    i_8_320_1780_0, i_8_320_1789_0, i_8_320_1807_0, i_8_320_1810_0,
    i_8_320_1903_0, i_8_320_1904_0, i_8_320_1912_0, i_8_320_1939_0,
    i_8_320_1973_0, i_8_320_1981_0, i_8_320_1984_0, i_8_320_1992_0,
    i_8_320_2039_0, i_8_320_2048_0, i_8_320_2107_0, i_8_320_2145_0,
    i_8_320_2155_0, i_8_320_2156_0, i_8_320_2173_0, i_8_320_2195_0,
    i_8_320_2249_0, i_8_320_2270_0, i_8_320_2290_0, i_8_320_2294_0;
  output o_8_320_0_0;
  assign o_8_320_0_0 = 0;
endmodule



// Benchmark "kernel_8_321" written by ABC on Sun Jul 19 10:08:38 2020

module kernel_8_321 ( 
    i_8_321_49_0, i_8_321_51_0, i_8_321_52_0, i_8_321_70_0, i_8_321_132_0,
    i_8_321_159_0, i_8_321_168_0, i_8_321_177_0, i_8_321_191_0,
    i_8_321_213_0, i_8_321_214_0, i_8_321_215_0, i_8_321_273_0,
    i_8_321_285_0, i_8_321_292_0, i_8_321_294_0, i_8_321_300_0,
    i_8_321_303_0, i_8_321_304_0, i_8_321_328_0, i_8_321_339_0,
    i_8_321_340_0, i_8_321_357_0, i_8_321_382_0, i_8_321_429_0,
    i_8_321_431_0, i_8_321_456_0, i_8_321_501_0, i_8_321_528_0,
    i_8_321_552_0, i_8_321_592_0, i_8_321_606_0, i_8_321_607_0,
    i_8_321_610_0, i_8_321_615_0, i_8_321_638_0, i_8_321_646_0,
    i_8_321_660_0, i_8_321_707_0, i_8_321_753_0, i_8_321_754_0,
    i_8_321_768_0, i_8_321_771_0, i_8_321_772_0, i_8_321_881_0,
    i_8_321_924_0, i_8_321_925_0, i_8_321_933_0, i_8_321_991_0,
    i_8_321_1093_0, i_8_321_1158_0, i_8_321_1159_0, i_8_321_1176_0,
    i_8_321_1195_0, i_8_321_1230_0, i_8_321_1267_0, i_8_321_1299_0,
    i_8_321_1313_0, i_8_321_1338_0, i_8_321_1347_0, i_8_321_1385_0,
    i_8_321_1410_0, i_8_321_1422_0, i_8_321_1489_0, i_8_321_1493_0,
    i_8_321_1528_0, i_8_321_1534_0, i_8_321_1553_0, i_8_321_1649_0,
    i_8_321_1671_0, i_8_321_1687_0, i_8_321_1731_0, i_8_321_1735_0,
    i_8_321_1770_0, i_8_321_1771_0, i_8_321_1818_0, i_8_321_1823_0,
    i_8_321_1824_0, i_8_321_1826_0, i_8_321_1831_0, i_8_321_1863_0,
    i_8_321_1885_0, i_8_321_1995_0, i_8_321_2004_0, i_8_321_2005_0,
    i_8_321_2022_0, i_8_321_2038_0, i_8_321_2074_0, i_8_321_2130_0,
    i_8_321_2153_0, i_8_321_2155_0, i_8_321_2157_0, i_8_321_2182_0,
    i_8_321_2184_0, i_8_321_2202_0, i_8_321_2211_0, i_8_321_2212_0,
    i_8_321_2229_0, i_8_321_2263_0, i_8_321_2292_0,
    o_8_321_0_0  );
  input  i_8_321_49_0, i_8_321_51_0, i_8_321_52_0, i_8_321_70_0,
    i_8_321_132_0, i_8_321_159_0, i_8_321_168_0, i_8_321_177_0,
    i_8_321_191_0, i_8_321_213_0, i_8_321_214_0, i_8_321_215_0,
    i_8_321_273_0, i_8_321_285_0, i_8_321_292_0, i_8_321_294_0,
    i_8_321_300_0, i_8_321_303_0, i_8_321_304_0, i_8_321_328_0,
    i_8_321_339_0, i_8_321_340_0, i_8_321_357_0, i_8_321_382_0,
    i_8_321_429_0, i_8_321_431_0, i_8_321_456_0, i_8_321_501_0,
    i_8_321_528_0, i_8_321_552_0, i_8_321_592_0, i_8_321_606_0,
    i_8_321_607_0, i_8_321_610_0, i_8_321_615_0, i_8_321_638_0,
    i_8_321_646_0, i_8_321_660_0, i_8_321_707_0, i_8_321_753_0,
    i_8_321_754_0, i_8_321_768_0, i_8_321_771_0, i_8_321_772_0,
    i_8_321_881_0, i_8_321_924_0, i_8_321_925_0, i_8_321_933_0,
    i_8_321_991_0, i_8_321_1093_0, i_8_321_1158_0, i_8_321_1159_0,
    i_8_321_1176_0, i_8_321_1195_0, i_8_321_1230_0, i_8_321_1267_0,
    i_8_321_1299_0, i_8_321_1313_0, i_8_321_1338_0, i_8_321_1347_0,
    i_8_321_1385_0, i_8_321_1410_0, i_8_321_1422_0, i_8_321_1489_0,
    i_8_321_1493_0, i_8_321_1528_0, i_8_321_1534_0, i_8_321_1553_0,
    i_8_321_1649_0, i_8_321_1671_0, i_8_321_1687_0, i_8_321_1731_0,
    i_8_321_1735_0, i_8_321_1770_0, i_8_321_1771_0, i_8_321_1818_0,
    i_8_321_1823_0, i_8_321_1824_0, i_8_321_1826_0, i_8_321_1831_0,
    i_8_321_1863_0, i_8_321_1885_0, i_8_321_1995_0, i_8_321_2004_0,
    i_8_321_2005_0, i_8_321_2022_0, i_8_321_2038_0, i_8_321_2074_0,
    i_8_321_2130_0, i_8_321_2153_0, i_8_321_2155_0, i_8_321_2157_0,
    i_8_321_2182_0, i_8_321_2184_0, i_8_321_2202_0, i_8_321_2211_0,
    i_8_321_2212_0, i_8_321_2229_0, i_8_321_2263_0, i_8_321_2292_0;
  output o_8_321_0_0;
  assign o_8_321_0_0 = ~((i_8_321_49_0 & ((i_8_321_610_0 & i_8_321_2130_0) | (~i_8_321_213_0 & ~i_8_321_528_0 & ~i_8_321_933_0 & ~i_8_321_1313_0 & ~i_8_321_2211_0 & i_8_321_2263_0))) | (~i_8_321_924_0 & ((~i_8_321_2212_0 & ((~i_8_321_51_0 & ((~i_8_321_660_0 & ~i_8_321_768_0 & ~i_8_321_933_0 & ~i_8_321_1176_0 & ~i_8_321_1528_0 & ~i_8_321_1735_0) | (~i_8_321_213_0 & i_8_321_2130_0))) | (~i_8_321_70_0 & ~i_8_321_177_0 & ~i_8_321_501_0 & ~i_8_321_772_0 & ~i_8_321_1649_0 & ~i_8_321_2202_0))) | (~i_8_321_215_0 & ((~i_8_321_768_0 & ~i_8_321_1176_0 & ~i_8_321_1195_0 & ~i_8_321_1528_0 & ~i_8_321_1771_0 & ~i_8_321_1885_0 & ~i_8_321_2004_0 & ~i_8_321_2202_0) | (~i_8_321_49_0 & ~i_8_321_159_0 & ~i_8_321_357_0 & ~i_8_321_933_0 & ~i_8_321_1230_0 & ~i_8_321_1313_0 & ~i_8_321_1347_0 & ~i_8_321_1671_0 & ~i_8_321_2263_0))) | (~i_8_321_177_0 & ~i_8_321_292_0 & ~i_8_321_772_0 & ~i_8_321_1176_0 & ~i_8_321_1771_0 & ~i_8_321_1885_0 & ~i_8_321_1995_0 & ~i_8_321_2263_0) | (~i_8_321_52_0 & ~i_8_321_456_0 & ~i_8_321_501_0 & ~i_8_321_925_0 & ~i_8_321_933_0 & ~i_8_321_1159_0 & ~i_8_321_2211_0 & ~i_8_321_2229_0))) | (~i_8_321_213_0 & ((~i_8_321_177_0 & ~i_8_321_501_0 & ~i_8_321_2004_0 & ~i_8_321_2005_0 & ~i_8_321_2202_0 & ~i_8_321_2211_0) | (~i_8_321_191_0 & ~i_8_321_456_0 & ~i_8_321_933_0 & ~i_8_321_1313_0 & ~i_8_321_1770_0 & ~i_8_321_2130_0 & ~i_8_321_2212_0 & ~i_8_321_2229_0))) | (~i_8_321_501_0 & ((i_8_321_615_0 & i_8_321_1267_0 & ~i_8_321_1649_0) | (i_8_321_328_0 & ~i_8_321_638_0 & ~i_8_321_1299_0 & ~i_8_321_1338_0 & ~i_8_321_1422_0 & ~i_8_321_2038_0 & ~i_8_321_2202_0))) | (~i_8_321_925_0 & ((~i_8_321_429_0 & ~i_8_321_754_0 & ~i_8_321_1410_0 & ~i_8_321_1649_0 & ~i_8_321_1671_0 & ~i_8_321_1771_0 & ~i_8_321_1824_0 & ~i_8_321_1826_0 & ~i_8_321_1885_0 & ~i_8_321_2074_0) | (~i_8_321_168_0 & ~i_8_321_1528_0 & i_8_321_1534_0 & ~i_8_321_2292_0))) | (~i_8_321_2212_0 & ((~i_8_321_340_0 & i_8_321_382_0 & ~i_8_321_552_0 & ~i_8_321_1176_0 & ~i_8_321_1195_0 & ~i_8_321_2038_0) | (i_8_321_303_0 & ~i_8_321_771_0 & ~i_8_321_2184_0))));
endmodule



// Benchmark "kernel_8_322" written by ABC on Sun Jul 19 10:08:39 2020

module kernel_8_322 ( 
    i_8_322_1_0, i_8_322_31_0, i_8_322_34_0, i_8_322_54_0, i_8_322_55_0,
    i_8_322_58_0, i_8_322_93_0, i_8_322_94_0, i_8_322_138_0, i_8_322_169_0,
    i_8_322_220_0, i_8_322_241_0, i_8_322_255_0, i_8_322_256_0,
    i_8_322_265_0, i_8_322_292_0, i_8_322_360_0, i_8_322_362_0,
    i_8_322_363_0, i_8_322_381_0, i_8_322_382_0, i_8_322_442_0,
    i_8_322_458_0, i_8_322_489_0, i_8_322_499_0, i_8_322_523_0,
    i_8_322_547_0, i_8_322_594_0, i_8_322_625_0, i_8_322_633_0,
    i_8_322_657_0, i_8_322_706_0, i_8_322_732_0, i_8_322_736_0,
    i_8_322_751_0, i_8_322_786_0, i_8_322_805_0, i_8_322_811_0,
    i_8_322_838_0, i_8_322_840_0, i_8_322_871_0, i_8_322_873_0,
    i_8_322_958_0, i_8_322_976_0, i_8_322_995_0, i_8_322_1071_0,
    i_8_322_1074_0, i_8_322_1182_0, i_8_322_1225_0, i_8_322_1240_0,
    i_8_322_1347_0, i_8_322_1360_0, i_8_322_1387_0, i_8_322_1403_0,
    i_8_322_1453_0, i_8_322_1471_0, i_8_322_1506_0, i_8_322_1524_0,
    i_8_322_1579_0, i_8_322_1615_0, i_8_322_1621_0, i_8_322_1630_0,
    i_8_322_1678_0, i_8_322_1681_0, i_8_322_1734_0, i_8_322_1743_0,
    i_8_322_1749_0, i_8_322_1750_0, i_8_322_1759_0, i_8_322_1760_0,
    i_8_322_1765_0, i_8_322_1768_0, i_8_322_1774_0, i_8_322_1777_0,
    i_8_322_1790_0, i_8_322_1821_0, i_8_322_1848_0, i_8_322_1849_0,
    i_8_322_1856_0, i_8_322_1857_0, i_8_322_1858_0, i_8_322_1902_0,
    i_8_322_1903_0, i_8_322_1946_0, i_8_322_1984_0, i_8_322_1995_0,
    i_8_322_2028_0, i_8_322_2029_0, i_8_322_2031_0, i_8_322_2092_0,
    i_8_322_2098_0, i_8_322_2119_0, i_8_322_2128_0, i_8_322_2129_0,
    i_8_322_2133_0, i_8_322_2134_0, i_8_322_2232_0, i_8_322_2245_0,
    i_8_322_2248_0, i_8_322_2259_0,
    o_8_322_0_0  );
  input  i_8_322_1_0, i_8_322_31_0, i_8_322_34_0, i_8_322_54_0,
    i_8_322_55_0, i_8_322_58_0, i_8_322_93_0, i_8_322_94_0, i_8_322_138_0,
    i_8_322_169_0, i_8_322_220_0, i_8_322_241_0, i_8_322_255_0,
    i_8_322_256_0, i_8_322_265_0, i_8_322_292_0, i_8_322_360_0,
    i_8_322_362_0, i_8_322_363_0, i_8_322_381_0, i_8_322_382_0,
    i_8_322_442_0, i_8_322_458_0, i_8_322_489_0, i_8_322_499_0,
    i_8_322_523_0, i_8_322_547_0, i_8_322_594_0, i_8_322_625_0,
    i_8_322_633_0, i_8_322_657_0, i_8_322_706_0, i_8_322_732_0,
    i_8_322_736_0, i_8_322_751_0, i_8_322_786_0, i_8_322_805_0,
    i_8_322_811_0, i_8_322_838_0, i_8_322_840_0, i_8_322_871_0,
    i_8_322_873_0, i_8_322_958_0, i_8_322_976_0, i_8_322_995_0,
    i_8_322_1071_0, i_8_322_1074_0, i_8_322_1182_0, i_8_322_1225_0,
    i_8_322_1240_0, i_8_322_1347_0, i_8_322_1360_0, i_8_322_1387_0,
    i_8_322_1403_0, i_8_322_1453_0, i_8_322_1471_0, i_8_322_1506_0,
    i_8_322_1524_0, i_8_322_1579_0, i_8_322_1615_0, i_8_322_1621_0,
    i_8_322_1630_0, i_8_322_1678_0, i_8_322_1681_0, i_8_322_1734_0,
    i_8_322_1743_0, i_8_322_1749_0, i_8_322_1750_0, i_8_322_1759_0,
    i_8_322_1760_0, i_8_322_1765_0, i_8_322_1768_0, i_8_322_1774_0,
    i_8_322_1777_0, i_8_322_1790_0, i_8_322_1821_0, i_8_322_1848_0,
    i_8_322_1849_0, i_8_322_1856_0, i_8_322_1857_0, i_8_322_1858_0,
    i_8_322_1902_0, i_8_322_1903_0, i_8_322_1946_0, i_8_322_1984_0,
    i_8_322_1995_0, i_8_322_2028_0, i_8_322_2029_0, i_8_322_2031_0,
    i_8_322_2092_0, i_8_322_2098_0, i_8_322_2119_0, i_8_322_2128_0,
    i_8_322_2129_0, i_8_322_2133_0, i_8_322_2134_0, i_8_322_2232_0,
    i_8_322_2245_0, i_8_322_2248_0, i_8_322_2259_0;
  output o_8_322_0_0;
  assign o_8_322_0_0 = 0;
endmodule



// Benchmark "kernel_8_323" written by ABC on Sun Jul 19 10:08:40 2020

module kernel_8_323 ( 
    i_8_323_85_0, i_8_323_88_0, i_8_323_121_0, i_8_323_193_0,
    i_8_323_222_0, i_8_323_223_0, i_8_323_266_0, i_8_323_272_0,
    i_8_323_288_0, i_8_323_345_0, i_8_323_348_0, i_8_323_374_0,
    i_8_323_391_0, i_8_323_419_0, i_8_323_424_0, i_8_323_426_0,
    i_8_323_427_0, i_8_323_444_0, i_8_323_451_0, i_8_323_457_0,
    i_8_323_491_0, i_8_323_526_0, i_8_323_589_0, i_8_323_590_0,
    i_8_323_595_0, i_8_323_599_0, i_8_323_625_0, i_8_323_649_0,
    i_8_323_652_0, i_8_323_666_0, i_8_323_679_0, i_8_323_685_0,
    i_8_323_709_0, i_8_323_715_0, i_8_323_761_0, i_8_323_798_0,
    i_8_323_815_0, i_8_323_820_0, i_8_323_838_0, i_8_323_847_0,
    i_8_323_909_0, i_8_323_996_0, i_8_323_1040_0, i_8_323_1047_0,
    i_8_323_1048_0, i_8_323_1084_0, i_8_323_1139_0, i_8_323_1141_0,
    i_8_323_1219_0, i_8_323_1228_0, i_8_323_1264_0, i_8_323_1269_0,
    i_8_323_1280_0, i_8_323_1309_0, i_8_323_1360_0, i_8_323_1373_0,
    i_8_323_1398_0, i_8_323_1407_0, i_8_323_1426_0, i_8_323_1440_0,
    i_8_323_1473_0, i_8_323_1498_0, i_8_323_1535_0, i_8_323_1544_0,
    i_8_323_1555_0, i_8_323_1638_0, i_8_323_1651_0, i_8_323_1680_0,
    i_8_323_1681_0, i_8_323_1731_0, i_8_323_1741_0, i_8_323_1761_0,
    i_8_323_1804_0, i_8_323_1810_0, i_8_323_1857_0, i_8_323_1883_0,
    i_8_323_1885_0, i_8_323_1930_0, i_8_323_1948_0, i_8_323_1959_0,
    i_8_323_1980_0, i_8_323_1993_0, i_8_323_2025_0, i_8_323_2059_0,
    i_8_323_2066_0, i_8_323_2106_0, i_8_323_2111_0, i_8_323_2134_0,
    i_8_323_2150_0, i_8_323_2152_0, i_8_323_2172_0, i_8_323_2221_0,
    i_8_323_2227_0, i_8_323_2235_0, i_8_323_2245_0, i_8_323_2258_0,
    i_8_323_2263_0, i_8_323_2273_0, i_8_323_2275_0, i_8_323_2281_0,
    o_8_323_0_0  );
  input  i_8_323_85_0, i_8_323_88_0, i_8_323_121_0, i_8_323_193_0,
    i_8_323_222_0, i_8_323_223_0, i_8_323_266_0, i_8_323_272_0,
    i_8_323_288_0, i_8_323_345_0, i_8_323_348_0, i_8_323_374_0,
    i_8_323_391_0, i_8_323_419_0, i_8_323_424_0, i_8_323_426_0,
    i_8_323_427_0, i_8_323_444_0, i_8_323_451_0, i_8_323_457_0,
    i_8_323_491_0, i_8_323_526_0, i_8_323_589_0, i_8_323_590_0,
    i_8_323_595_0, i_8_323_599_0, i_8_323_625_0, i_8_323_649_0,
    i_8_323_652_0, i_8_323_666_0, i_8_323_679_0, i_8_323_685_0,
    i_8_323_709_0, i_8_323_715_0, i_8_323_761_0, i_8_323_798_0,
    i_8_323_815_0, i_8_323_820_0, i_8_323_838_0, i_8_323_847_0,
    i_8_323_909_0, i_8_323_996_0, i_8_323_1040_0, i_8_323_1047_0,
    i_8_323_1048_0, i_8_323_1084_0, i_8_323_1139_0, i_8_323_1141_0,
    i_8_323_1219_0, i_8_323_1228_0, i_8_323_1264_0, i_8_323_1269_0,
    i_8_323_1280_0, i_8_323_1309_0, i_8_323_1360_0, i_8_323_1373_0,
    i_8_323_1398_0, i_8_323_1407_0, i_8_323_1426_0, i_8_323_1440_0,
    i_8_323_1473_0, i_8_323_1498_0, i_8_323_1535_0, i_8_323_1544_0,
    i_8_323_1555_0, i_8_323_1638_0, i_8_323_1651_0, i_8_323_1680_0,
    i_8_323_1681_0, i_8_323_1731_0, i_8_323_1741_0, i_8_323_1761_0,
    i_8_323_1804_0, i_8_323_1810_0, i_8_323_1857_0, i_8_323_1883_0,
    i_8_323_1885_0, i_8_323_1930_0, i_8_323_1948_0, i_8_323_1959_0,
    i_8_323_1980_0, i_8_323_1993_0, i_8_323_2025_0, i_8_323_2059_0,
    i_8_323_2066_0, i_8_323_2106_0, i_8_323_2111_0, i_8_323_2134_0,
    i_8_323_2150_0, i_8_323_2152_0, i_8_323_2172_0, i_8_323_2221_0,
    i_8_323_2227_0, i_8_323_2235_0, i_8_323_2245_0, i_8_323_2258_0,
    i_8_323_2263_0, i_8_323_2273_0, i_8_323_2275_0, i_8_323_2281_0;
  output o_8_323_0_0;
  assign o_8_323_0_0 = 0;
endmodule



// Benchmark "kernel_8_324" written by ABC on Sun Jul 19 10:08:40 2020

module kernel_8_324 ( 
    i_8_324_6_0, i_8_324_11_0, i_8_324_14_0, i_8_324_43_0, i_8_324_61_0,
    i_8_324_78_0, i_8_324_79_0, i_8_324_80_0, i_8_324_85_0, i_8_324_87_0,
    i_8_324_105_0, i_8_324_106_0, i_8_324_124_0, i_8_324_141_0,
    i_8_324_142_0, i_8_324_258_0, i_8_324_268_0, i_8_324_285_0,
    i_8_324_294_0, i_8_324_295_0, i_8_324_309_0, i_8_324_336_0,
    i_8_324_339_0, i_8_324_345_0, i_8_324_364_0, i_8_324_370_0,
    i_8_324_525_0, i_8_324_529_0, i_8_324_555_0, i_8_324_564_0,
    i_8_324_595_0, i_8_324_598_0, i_8_324_601_0, i_8_324_608_0,
    i_8_324_609_0, i_8_324_624_0, i_8_324_634_0, i_8_324_642_0,
    i_8_324_645_0, i_8_324_654_0, i_8_324_660_0, i_8_324_664_0,
    i_8_324_688_0, i_8_324_708_0, i_8_324_718_0, i_8_324_726_0,
    i_8_324_753_0, i_8_324_768_0, i_8_324_783_0, i_8_324_789_0,
    i_8_324_825_0, i_8_324_834_0, i_8_324_835_0, i_8_324_840_0,
    i_8_324_853_0, i_8_324_870_0, i_8_324_939_0, i_8_324_950_0,
    i_8_324_958_0, i_8_324_1012_0, i_8_324_1116_0, i_8_324_1164_0,
    i_8_324_1185_0, i_8_324_1213_0, i_8_324_1299_0, i_8_324_1309_0,
    i_8_324_1317_0, i_8_324_1330_0, i_8_324_1357_0, i_8_324_1375_0,
    i_8_324_1380_0, i_8_324_1409_0, i_8_324_1437_0, i_8_324_1438_0,
    i_8_324_1446_0, i_8_324_1473_0, i_8_324_1542_0, i_8_324_1546_0,
    i_8_324_1565_0, i_8_324_1588_0, i_8_324_1590_0, i_8_324_1600_0,
    i_8_324_1734_0, i_8_324_1779_0, i_8_324_1857_0, i_8_324_1861_0,
    i_8_324_1905_0, i_8_324_1906_0, i_8_324_2034_0, i_8_324_2037_0,
    i_8_324_2049_0, i_8_324_2073_0, i_8_324_2085_0, i_8_324_2090_0,
    i_8_324_2121_0, i_8_324_2172_0, i_8_324_2191_0, i_8_324_2193_0,
    i_8_324_2235_0, i_8_324_2268_0,
    o_8_324_0_0  );
  input  i_8_324_6_0, i_8_324_11_0, i_8_324_14_0, i_8_324_43_0,
    i_8_324_61_0, i_8_324_78_0, i_8_324_79_0, i_8_324_80_0, i_8_324_85_0,
    i_8_324_87_0, i_8_324_105_0, i_8_324_106_0, i_8_324_124_0,
    i_8_324_141_0, i_8_324_142_0, i_8_324_258_0, i_8_324_268_0,
    i_8_324_285_0, i_8_324_294_0, i_8_324_295_0, i_8_324_309_0,
    i_8_324_336_0, i_8_324_339_0, i_8_324_345_0, i_8_324_364_0,
    i_8_324_370_0, i_8_324_525_0, i_8_324_529_0, i_8_324_555_0,
    i_8_324_564_0, i_8_324_595_0, i_8_324_598_0, i_8_324_601_0,
    i_8_324_608_0, i_8_324_609_0, i_8_324_624_0, i_8_324_634_0,
    i_8_324_642_0, i_8_324_645_0, i_8_324_654_0, i_8_324_660_0,
    i_8_324_664_0, i_8_324_688_0, i_8_324_708_0, i_8_324_718_0,
    i_8_324_726_0, i_8_324_753_0, i_8_324_768_0, i_8_324_783_0,
    i_8_324_789_0, i_8_324_825_0, i_8_324_834_0, i_8_324_835_0,
    i_8_324_840_0, i_8_324_853_0, i_8_324_870_0, i_8_324_939_0,
    i_8_324_950_0, i_8_324_958_0, i_8_324_1012_0, i_8_324_1116_0,
    i_8_324_1164_0, i_8_324_1185_0, i_8_324_1213_0, i_8_324_1299_0,
    i_8_324_1309_0, i_8_324_1317_0, i_8_324_1330_0, i_8_324_1357_0,
    i_8_324_1375_0, i_8_324_1380_0, i_8_324_1409_0, i_8_324_1437_0,
    i_8_324_1438_0, i_8_324_1446_0, i_8_324_1473_0, i_8_324_1542_0,
    i_8_324_1546_0, i_8_324_1565_0, i_8_324_1588_0, i_8_324_1590_0,
    i_8_324_1600_0, i_8_324_1734_0, i_8_324_1779_0, i_8_324_1857_0,
    i_8_324_1861_0, i_8_324_1905_0, i_8_324_1906_0, i_8_324_2034_0,
    i_8_324_2037_0, i_8_324_2049_0, i_8_324_2073_0, i_8_324_2085_0,
    i_8_324_2090_0, i_8_324_2121_0, i_8_324_2172_0, i_8_324_2191_0,
    i_8_324_2193_0, i_8_324_2235_0, i_8_324_2268_0;
  output o_8_324_0_0;
  assign o_8_324_0_0 = 0;
endmodule



// Benchmark "kernel_8_325" written by ABC on Sun Jul 19 10:08:41 2020

module kernel_8_325 ( 
    i_8_325_41_0, i_8_325_65_0, i_8_325_82_0, i_8_325_91_0, i_8_325_92_0,
    i_8_325_128_0, i_8_325_131_0, i_8_325_136_0, i_8_325_137_0,
    i_8_325_140_0, i_8_325_142_0, i_8_325_163_0, i_8_325_181_0,
    i_8_325_189_0, i_8_325_212_0, i_8_325_236_0, i_8_325_282_0,
    i_8_325_307_0, i_8_325_308_0, i_8_325_316_0, i_8_325_335_0,
    i_8_325_344_0, i_8_325_380_0, i_8_325_446_0, i_8_325_451_0,
    i_8_325_452_0, i_8_325_486_0, i_8_325_491_0, i_8_325_527_0,
    i_8_325_542_0, i_8_325_553_0, i_8_325_554_0, i_8_325_595_0,
    i_8_325_604_0, i_8_325_614_0, i_8_325_622_0, i_8_325_652_0,
    i_8_325_661_0, i_8_325_686_0, i_8_325_696_0, i_8_325_700_0,
    i_8_325_703_0, i_8_325_730_0, i_8_325_731_0, i_8_325_792_0,
    i_8_325_837_0, i_8_325_838_0, i_8_325_841_0, i_8_325_852_0,
    i_8_325_878_0, i_8_325_929_0, i_8_325_932_0, i_8_325_956_0,
    i_8_325_965_0, i_8_325_973_0, i_8_325_1018_0, i_8_325_1035_0,
    i_8_325_1061_0, i_8_325_1115_0, i_8_325_1271_0, i_8_325_1283_0,
    i_8_325_1297_0, i_8_325_1315_0, i_8_325_1325_0, i_8_325_1328_0,
    i_8_325_1367_0, i_8_325_1373_0, i_8_325_1449_0, i_8_325_1621_0,
    i_8_325_1622_0, i_8_325_1639_0, i_8_325_1682_0, i_8_325_1686_0,
    i_8_325_1707_0, i_8_325_1715_0, i_8_325_1729_0, i_8_325_1733_0,
    i_8_325_1744_0, i_8_325_1760_0, i_8_325_1764_0, i_8_325_1828_0,
    i_8_325_1838_0, i_8_325_1882_0, i_8_325_1900_0, i_8_325_1937_0,
    i_8_325_1949_0, i_8_325_2017_0, i_8_325_2020_0, i_8_325_2108_0,
    i_8_325_2110_0, i_8_325_2144_0, i_8_325_2146_0, i_8_325_2153_0,
    i_8_325_2180_0, i_8_325_2198_0, i_8_325_2206_0, i_8_325_2212_0,
    i_8_325_2246_0, i_8_325_2264_0, i_8_325_2270_0,
    o_8_325_0_0  );
  input  i_8_325_41_0, i_8_325_65_0, i_8_325_82_0, i_8_325_91_0,
    i_8_325_92_0, i_8_325_128_0, i_8_325_131_0, i_8_325_136_0,
    i_8_325_137_0, i_8_325_140_0, i_8_325_142_0, i_8_325_163_0,
    i_8_325_181_0, i_8_325_189_0, i_8_325_212_0, i_8_325_236_0,
    i_8_325_282_0, i_8_325_307_0, i_8_325_308_0, i_8_325_316_0,
    i_8_325_335_0, i_8_325_344_0, i_8_325_380_0, i_8_325_446_0,
    i_8_325_451_0, i_8_325_452_0, i_8_325_486_0, i_8_325_491_0,
    i_8_325_527_0, i_8_325_542_0, i_8_325_553_0, i_8_325_554_0,
    i_8_325_595_0, i_8_325_604_0, i_8_325_614_0, i_8_325_622_0,
    i_8_325_652_0, i_8_325_661_0, i_8_325_686_0, i_8_325_696_0,
    i_8_325_700_0, i_8_325_703_0, i_8_325_730_0, i_8_325_731_0,
    i_8_325_792_0, i_8_325_837_0, i_8_325_838_0, i_8_325_841_0,
    i_8_325_852_0, i_8_325_878_0, i_8_325_929_0, i_8_325_932_0,
    i_8_325_956_0, i_8_325_965_0, i_8_325_973_0, i_8_325_1018_0,
    i_8_325_1035_0, i_8_325_1061_0, i_8_325_1115_0, i_8_325_1271_0,
    i_8_325_1283_0, i_8_325_1297_0, i_8_325_1315_0, i_8_325_1325_0,
    i_8_325_1328_0, i_8_325_1367_0, i_8_325_1373_0, i_8_325_1449_0,
    i_8_325_1621_0, i_8_325_1622_0, i_8_325_1639_0, i_8_325_1682_0,
    i_8_325_1686_0, i_8_325_1707_0, i_8_325_1715_0, i_8_325_1729_0,
    i_8_325_1733_0, i_8_325_1744_0, i_8_325_1760_0, i_8_325_1764_0,
    i_8_325_1828_0, i_8_325_1838_0, i_8_325_1882_0, i_8_325_1900_0,
    i_8_325_1937_0, i_8_325_1949_0, i_8_325_2017_0, i_8_325_2020_0,
    i_8_325_2108_0, i_8_325_2110_0, i_8_325_2144_0, i_8_325_2146_0,
    i_8_325_2153_0, i_8_325_2180_0, i_8_325_2198_0, i_8_325_2206_0,
    i_8_325_2212_0, i_8_325_2246_0, i_8_325_2264_0, i_8_325_2270_0;
  output o_8_325_0_0;
  assign o_8_325_0_0 = 0;
endmodule



// Benchmark "kernel_8_326" written by ABC on Sun Jul 19 10:08:42 2020

module kernel_8_326 ( 
    i_8_326_21_0, i_8_326_22_0, i_8_326_32_0, i_8_326_73_0, i_8_326_103_0,
    i_8_326_148_0, i_8_326_150_0, i_8_326_190_0, i_8_326_202_0,
    i_8_326_247_0, i_8_326_275_0, i_8_326_355_0, i_8_326_365_0,
    i_8_326_373_0, i_8_326_382_0, i_8_326_383_0, i_8_326_386_0,
    i_8_326_426_0, i_8_326_445_0, i_8_326_469_0, i_8_326_490_0,
    i_8_326_499_0, i_8_326_517_0, i_8_326_652_0, i_8_326_704_0,
    i_8_326_733_0, i_8_326_751_0, i_8_326_752_0, i_8_326_777_0,
    i_8_326_814_0, i_8_326_832_0, i_8_326_837_0, i_8_326_846_0,
    i_8_326_913_0, i_8_326_941_0, i_8_326_967_0, i_8_326_1069_0,
    i_8_326_1072_0, i_8_326_1112_0, i_8_326_1174_0, i_8_326_1202_0,
    i_8_326_1224_0, i_8_326_1233_0, i_8_326_1264_0, i_8_326_1284_0,
    i_8_326_1350_0, i_8_326_1394_0, i_8_326_1399_0, i_8_326_1404_0,
    i_8_326_1452_0, i_8_326_1479_0, i_8_326_1497_0, i_8_326_1531_0,
    i_8_326_1552_0, i_8_326_1597_0, i_8_326_1625_0, i_8_326_1648_0,
    i_8_326_1649_0, i_8_326_1657_0, i_8_326_1660_0, i_8_326_1676_0,
    i_8_326_1677_0, i_8_326_1705_0, i_8_326_1746_0, i_8_326_1792_0,
    i_8_326_1805_0, i_8_326_1806_0, i_8_326_1808_0, i_8_326_1812_0,
    i_8_326_1821_0, i_8_326_1840_0, i_8_326_1848_0, i_8_326_1849_0,
    i_8_326_1850_0, i_8_326_1864_0, i_8_326_1866_0, i_8_326_1890_0,
    i_8_326_1917_0, i_8_326_1928_0, i_8_326_1951_0, i_8_326_1952_0,
    i_8_326_1966_0, i_8_326_1972_0, i_8_326_1989_0, i_8_326_1997_0,
    i_8_326_2011_0, i_8_326_2038_0, i_8_326_2088_0, i_8_326_2089_0,
    i_8_326_2145_0, i_8_326_2146_0, i_8_326_2148_0, i_8_326_2149_0,
    i_8_326_2150_0, i_8_326_2155_0, i_8_326_2224_0, i_8_326_2233_0,
    i_8_326_2257_0, i_8_326_2273_0, i_8_326_2299_0,
    o_8_326_0_0  );
  input  i_8_326_21_0, i_8_326_22_0, i_8_326_32_0, i_8_326_73_0,
    i_8_326_103_0, i_8_326_148_0, i_8_326_150_0, i_8_326_190_0,
    i_8_326_202_0, i_8_326_247_0, i_8_326_275_0, i_8_326_355_0,
    i_8_326_365_0, i_8_326_373_0, i_8_326_382_0, i_8_326_383_0,
    i_8_326_386_0, i_8_326_426_0, i_8_326_445_0, i_8_326_469_0,
    i_8_326_490_0, i_8_326_499_0, i_8_326_517_0, i_8_326_652_0,
    i_8_326_704_0, i_8_326_733_0, i_8_326_751_0, i_8_326_752_0,
    i_8_326_777_0, i_8_326_814_0, i_8_326_832_0, i_8_326_837_0,
    i_8_326_846_0, i_8_326_913_0, i_8_326_941_0, i_8_326_967_0,
    i_8_326_1069_0, i_8_326_1072_0, i_8_326_1112_0, i_8_326_1174_0,
    i_8_326_1202_0, i_8_326_1224_0, i_8_326_1233_0, i_8_326_1264_0,
    i_8_326_1284_0, i_8_326_1350_0, i_8_326_1394_0, i_8_326_1399_0,
    i_8_326_1404_0, i_8_326_1452_0, i_8_326_1479_0, i_8_326_1497_0,
    i_8_326_1531_0, i_8_326_1552_0, i_8_326_1597_0, i_8_326_1625_0,
    i_8_326_1648_0, i_8_326_1649_0, i_8_326_1657_0, i_8_326_1660_0,
    i_8_326_1676_0, i_8_326_1677_0, i_8_326_1705_0, i_8_326_1746_0,
    i_8_326_1792_0, i_8_326_1805_0, i_8_326_1806_0, i_8_326_1808_0,
    i_8_326_1812_0, i_8_326_1821_0, i_8_326_1840_0, i_8_326_1848_0,
    i_8_326_1849_0, i_8_326_1850_0, i_8_326_1864_0, i_8_326_1866_0,
    i_8_326_1890_0, i_8_326_1917_0, i_8_326_1928_0, i_8_326_1951_0,
    i_8_326_1952_0, i_8_326_1966_0, i_8_326_1972_0, i_8_326_1989_0,
    i_8_326_1997_0, i_8_326_2011_0, i_8_326_2038_0, i_8_326_2088_0,
    i_8_326_2089_0, i_8_326_2145_0, i_8_326_2146_0, i_8_326_2148_0,
    i_8_326_2149_0, i_8_326_2150_0, i_8_326_2155_0, i_8_326_2224_0,
    i_8_326_2233_0, i_8_326_2257_0, i_8_326_2273_0, i_8_326_2299_0;
  output o_8_326_0_0;
  assign o_8_326_0_0 = 0;
endmodule



// Benchmark "kernel_8_327" written by ABC on Sun Jul 19 10:08:43 2020

module kernel_8_327 ( 
    i_8_327_34_0, i_8_327_54_0, i_8_327_55_0, i_8_327_86_0, i_8_327_87_0,
    i_8_327_96_0, i_8_327_103_0, i_8_327_142_0, i_8_327_167_0,
    i_8_327_201_0, i_8_327_202_0, i_8_327_223_0, i_8_327_255_0,
    i_8_327_369_0, i_8_327_415_0, i_8_327_421_0, i_8_327_441_0,
    i_8_327_456_0, i_8_327_471_0, i_8_327_479_0, i_8_327_500_0,
    i_8_327_526_0, i_8_327_528_0, i_8_327_530_0, i_8_327_552_0,
    i_8_327_553_0, i_8_327_601_0, i_8_327_625_0, i_8_327_660_0,
    i_8_327_714_0, i_8_327_772_0, i_8_327_795_0, i_8_327_815_0,
    i_8_327_827_0, i_8_327_868_0, i_8_327_888_0, i_8_327_895_0,
    i_8_327_1012_0, i_8_327_1028_0, i_8_327_1051_0, i_8_327_1059_0,
    i_8_327_1061_0, i_8_327_1084_0, i_8_327_1112_0, i_8_327_1156_0,
    i_8_327_1188_0, i_8_327_1198_0, i_8_327_1215_0, i_8_327_1249_0,
    i_8_327_1259_0, i_8_327_1266_0, i_8_327_1274_0, i_8_327_1277_0,
    i_8_327_1281_0, i_8_327_1325_0, i_8_327_1390_0, i_8_327_1417_0,
    i_8_327_1435_0, i_8_327_1438_0, i_8_327_1449_0, i_8_327_1471_0,
    i_8_327_1480_0, i_8_327_1536_0, i_8_327_1549_0, i_8_327_1551_0,
    i_8_327_1552_0, i_8_327_1579_0, i_8_327_1627_0, i_8_327_1629_0,
    i_8_327_1633_0, i_8_327_1668_0, i_8_327_1675_0, i_8_327_1681_0,
    i_8_327_1682_0, i_8_327_1707_0, i_8_327_1726_0, i_8_327_1731_0,
    i_8_327_1732_0, i_8_327_1744_0, i_8_327_1749_0, i_8_327_1753_0,
    i_8_327_1758_0, i_8_327_1813_0, i_8_327_1855_0, i_8_327_1858_0,
    i_8_327_1872_0, i_8_327_1873_0, i_8_327_1889_0, i_8_327_1894_0,
    i_8_327_1902_0, i_8_327_2002_0, i_8_327_2074_0, i_8_327_2136_0,
    i_8_327_2154_0, i_8_327_2191_0, i_8_327_2212_0, i_8_327_2228_0,
    i_8_327_2259_0, i_8_327_2271_0, i_8_327_2272_0,
    o_8_327_0_0  );
  input  i_8_327_34_0, i_8_327_54_0, i_8_327_55_0, i_8_327_86_0,
    i_8_327_87_0, i_8_327_96_0, i_8_327_103_0, i_8_327_142_0,
    i_8_327_167_0, i_8_327_201_0, i_8_327_202_0, i_8_327_223_0,
    i_8_327_255_0, i_8_327_369_0, i_8_327_415_0, i_8_327_421_0,
    i_8_327_441_0, i_8_327_456_0, i_8_327_471_0, i_8_327_479_0,
    i_8_327_500_0, i_8_327_526_0, i_8_327_528_0, i_8_327_530_0,
    i_8_327_552_0, i_8_327_553_0, i_8_327_601_0, i_8_327_625_0,
    i_8_327_660_0, i_8_327_714_0, i_8_327_772_0, i_8_327_795_0,
    i_8_327_815_0, i_8_327_827_0, i_8_327_868_0, i_8_327_888_0,
    i_8_327_895_0, i_8_327_1012_0, i_8_327_1028_0, i_8_327_1051_0,
    i_8_327_1059_0, i_8_327_1061_0, i_8_327_1084_0, i_8_327_1112_0,
    i_8_327_1156_0, i_8_327_1188_0, i_8_327_1198_0, i_8_327_1215_0,
    i_8_327_1249_0, i_8_327_1259_0, i_8_327_1266_0, i_8_327_1274_0,
    i_8_327_1277_0, i_8_327_1281_0, i_8_327_1325_0, i_8_327_1390_0,
    i_8_327_1417_0, i_8_327_1435_0, i_8_327_1438_0, i_8_327_1449_0,
    i_8_327_1471_0, i_8_327_1480_0, i_8_327_1536_0, i_8_327_1549_0,
    i_8_327_1551_0, i_8_327_1552_0, i_8_327_1579_0, i_8_327_1627_0,
    i_8_327_1629_0, i_8_327_1633_0, i_8_327_1668_0, i_8_327_1675_0,
    i_8_327_1681_0, i_8_327_1682_0, i_8_327_1707_0, i_8_327_1726_0,
    i_8_327_1731_0, i_8_327_1732_0, i_8_327_1744_0, i_8_327_1749_0,
    i_8_327_1753_0, i_8_327_1758_0, i_8_327_1813_0, i_8_327_1855_0,
    i_8_327_1858_0, i_8_327_1872_0, i_8_327_1873_0, i_8_327_1889_0,
    i_8_327_1894_0, i_8_327_1902_0, i_8_327_2002_0, i_8_327_2074_0,
    i_8_327_2136_0, i_8_327_2154_0, i_8_327_2191_0, i_8_327_2212_0,
    i_8_327_2228_0, i_8_327_2259_0, i_8_327_2271_0, i_8_327_2272_0;
  output o_8_327_0_0;
  assign o_8_327_0_0 = 0;
endmodule



// Benchmark "kernel_8_328" written by ABC on Sun Jul 19 10:08:44 2020

module kernel_8_328 ( 
    i_8_328_22_0, i_8_328_64_0, i_8_328_67_0, i_8_328_94_0, i_8_328_114_0,
    i_8_328_193_0, i_8_328_194_0, i_8_328_226_0, i_8_328_275_0,
    i_8_328_283_0, i_8_328_297_0, i_8_328_361_0, i_8_328_382_0,
    i_8_328_391_0, i_8_328_416_0, i_8_328_426_0, i_8_328_484_0,
    i_8_328_492_0, i_8_328_493_0, i_8_328_505_0, i_8_328_518_0,
    i_8_328_535_0, i_8_328_546_0, i_8_328_567_0, i_8_328_631_0,
    i_8_328_635_0, i_8_328_652_0, i_8_328_660_0, i_8_328_691_0,
    i_8_328_693_0, i_8_328_709_0, i_8_328_739_0, i_8_328_750_0,
    i_8_328_751_0, i_8_328_814_0, i_8_328_815_0, i_8_328_837_0,
    i_8_328_851_0, i_8_328_865_0, i_8_328_904_0, i_8_328_964_0,
    i_8_328_970_0, i_8_328_1012_0, i_8_328_1033_0, i_8_328_1072_0,
    i_8_328_1102_0, i_8_328_1134_0, i_8_328_1135_0, i_8_328_1171_0,
    i_8_328_1192_0, i_8_328_1202_0, i_8_328_1229_0, i_8_328_1249_0,
    i_8_328_1278_0, i_8_328_1282_0, i_8_328_1283_0, i_8_328_1286_0,
    i_8_328_1306_0, i_8_328_1391_0, i_8_328_1397_0, i_8_328_1439_0,
    i_8_328_1450_0, i_8_328_1477_0, i_8_328_1478_0, i_8_328_1489_0,
    i_8_328_1526_0, i_8_328_1546_0, i_8_328_1552_0, i_8_328_1582_0,
    i_8_328_1606_0, i_8_328_1640_0, i_8_328_1660_0, i_8_328_1673_0,
    i_8_328_1704_0, i_8_328_1769_0, i_8_328_1784_0, i_8_328_1819_0,
    i_8_328_1840_0, i_8_328_1849_0, i_8_328_1885_0, i_8_328_1902_0,
    i_8_328_1957_0, i_8_328_1981_0, i_8_328_1997_0, i_8_328_2011_0,
    i_8_328_2014_0, i_8_328_2145_0, i_8_328_2149_0, i_8_328_2171_0,
    i_8_328_2174_0, i_8_328_2214_0, i_8_328_2216_0, i_8_328_2242_0,
    i_8_328_2245_0, i_8_328_2255_0, i_8_328_2258_0, i_8_328_2262_0,
    i_8_328_2289_0, i_8_328_2300_0, i_8_328_2303_0,
    o_8_328_0_0  );
  input  i_8_328_22_0, i_8_328_64_0, i_8_328_67_0, i_8_328_94_0,
    i_8_328_114_0, i_8_328_193_0, i_8_328_194_0, i_8_328_226_0,
    i_8_328_275_0, i_8_328_283_0, i_8_328_297_0, i_8_328_361_0,
    i_8_328_382_0, i_8_328_391_0, i_8_328_416_0, i_8_328_426_0,
    i_8_328_484_0, i_8_328_492_0, i_8_328_493_0, i_8_328_505_0,
    i_8_328_518_0, i_8_328_535_0, i_8_328_546_0, i_8_328_567_0,
    i_8_328_631_0, i_8_328_635_0, i_8_328_652_0, i_8_328_660_0,
    i_8_328_691_0, i_8_328_693_0, i_8_328_709_0, i_8_328_739_0,
    i_8_328_750_0, i_8_328_751_0, i_8_328_814_0, i_8_328_815_0,
    i_8_328_837_0, i_8_328_851_0, i_8_328_865_0, i_8_328_904_0,
    i_8_328_964_0, i_8_328_970_0, i_8_328_1012_0, i_8_328_1033_0,
    i_8_328_1072_0, i_8_328_1102_0, i_8_328_1134_0, i_8_328_1135_0,
    i_8_328_1171_0, i_8_328_1192_0, i_8_328_1202_0, i_8_328_1229_0,
    i_8_328_1249_0, i_8_328_1278_0, i_8_328_1282_0, i_8_328_1283_0,
    i_8_328_1286_0, i_8_328_1306_0, i_8_328_1391_0, i_8_328_1397_0,
    i_8_328_1439_0, i_8_328_1450_0, i_8_328_1477_0, i_8_328_1478_0,
    i_8_328_1489_0, i_8_328_1526_0, i_8_328_1546_0, i_8_328_1552_0,
    i_8_328_1582_0, i_8_328_1606_0, i_8_328_1640_0, i_8_328_1660_0,
    i_8_328_1673_0, i_8_328_1704_0, i_8_328_1769_0, i_8_328_1784_0,
    i_8_328_1819_0, i_8_328_1840_0, i_8_328_1849_0, i_8_328_1885_0,
    i_8_328_1902_0, i_8_328_1957_0, i_8_328_1981_0, i_8_328_1997_0,
    i_8_328_2011_0, i_8_328_2014_0, i_8_328_2145_0, i_8_328_2149_0,
    i_8_328_2171_0, i_8_328_2174_0, i_8_328_2214_0, i_8_328_2216_0,
    i_8_328_2242_0, i_8_328_2245_0, i_8_328_2255_0, i_8_328_2258_0,
    i_8_328_2262_0, i_8_328_2289_0, i_8_328_2300_0, i_8_328_2303_0;
  output o_8_328_0_0;
  assign o_8_328_0_0 = 0;
endmodule



// Benchmark "kernel_8_329" written by ABC on Sun Jul 19 10:08:44 2020

module kernel_8_329 ( 
    i_8_329_22_0, i_8_329_23_0, i_8_329_28_0, i_8_329_29_0, i_8_329_56_0,
    i_8_329_67_0, i_8_329_74_0, i_8_329_79_0, i_8_329_162_0, i_8_329_172_0,
    i_8_329_181_0, i_8_329_191_0, i_8_329_193_0, i_8_329_198_0,
    i_8_329_218_0, i_8_329_226_0, i_8_329_227_0, i_8_329_229_0,
    i_8_329_231_0, i_8_329_299_0, i_8_329_302_0, i_8_329_370_0,
    i_8_329_379_0, i_8_329_383_0, i_8_329_414_0, i_8_329_415_0,
    i_8_329_424_0, i_8_329_434_0, i_8_329_463_0, i_8_329_488_0,
    i_8_329_492_0, i_8_329_493_0, i_8_329_592_0, i_8_329_604_0,
    i_8_329_605_0, i_8_329_658_0, i_8_329_679_0, i_8_329_823_0,
    i_8_329_837_0, i_8_329_838_0, i_8_329_839_0, i_8_329_842_0,
    i_8_329_859_0, i_8_329_869_0, i_8_329_873_0, i_8_329_883_0,
    i_8_329_955_0, i_8_329_965_0, i_8_329_971_0, i_8_329_1041_0,
    i_8_329_1104_0, i_8_329_1129_0, i_8_329_1175_0, i_8_329_1189_0,
    i_8_329_1237_0, i_8_329_1279_0, i_8_329_1297_0, i_8_329_1307_0,
    i_8_329_1328_0, i_8_329_1341_0, i_8_329_1360_0, i_8_329_1382_0,
    i_8_329_1441_0, i_8_329_1471_0, i_8_329_1472_0, i_8_329_1564_0,
    i_8_329_1573_0, i_8_329_1585_0, i_8_329_1603_0, i_8_329_1604_0,
    i_8_329_1622_0, i_8_329_1634_0, i_8_329_1652_0, i_8_329_1688_0,
    i_8_329_1756_0, i_8_329_1774_0, i_8_329_1775_0, i_8_329_1805_0,
    i_8_329_1809_0, i_8_329_1843_0, i_8_329_1873_0, i_8_329_1874_0,
    i_8_329_1882_0, i_8_329_1909_0, i_8_329_1982_0, i_8_329_1989_0,
    i_8_329_1991_0, i_8_329_1995_0, i_8_329_2052_0, i_8_329_2054_0,
    i_8_329_2065_0, i_8_329_2140_0, i_8_329_2145_0, i_8_329_2170_0,
    i_8_329_2171_0, i_8_329_2214_0, i_8_329_2215_0, i_8_329_2216_0,
    i_8_329_2233_0, i_8_329_2243_0,
    o_8_329_0_0  );
  input  i_8_329_22_0, i_8_329_23_0, i_8_329_28_0, i_8_329_29_0,
    i_8_329_56_0, i_8_329_67_0, i_8_329_74_0, i_8_329_79_0, i_8_329_162_0,
    i_8_329_172_0, i_8_329_181_0, i_8_329_191_0, i_8_329_193_0,
    i_8_329_198_0, i_8_329_218_0, i_8_329_226_0, i_8_329_227_0,
    i_8_329_229_0, i_8_329_231_0, i_8_329_299_0, i_8_329_302_0,
    i_8_329_370_0, i_8_329_379_0, i_8_329_383_0, i_8_329_414_0,
    i_8_329_415_0, i_8_329_424_0, i_8_329_434_0, i_8_329_463_0,
    i_8_329_488_0, i_8_329_492_0, i_8_329_493_0, i_8_329_592_0,
    i_8_329_604_0, i_8_329_605_0, i_8_329_658_0, i_8_329_679_0,
    i_8_329_823_0, i_8_329_837_0, i_8_329_838_0, i_8_329_839_0,
    i_8_329_842_0, i_8_329_859_0, i_8_329_869_0, i_8_329_873_0,
    i_8_329_883_0, i_8_329_955_0, i_8_329_965_0, i_8_329_971_0,
    i_8_329_1041_0, i_8_329_1104_0, i_8_329_1129_0, i_8_329_1175_0,
    i_8_329_1189_0, i_8_329_1237_0, i_8_329_1279_0, i_8_329_1297_0,
    i_8_329_1307_0, i_8_329_1328_0, i_8_329_1341_0, i_8_329_1360_0,
    i_8_329_1382_0, i_8_329_1441_0, i_8_329_1471_0, i_8_329_1472_0,
    i_8_329_1564_0, i_8_329_1573_0, i_8_329_1585_0, i_8_329_1603_0,
    i_8_329_1604_0, i_8_329_1622_0, i_8_329_1634_0, i_8_329_1652_0,
    i_8_329_1688_0, i_8_329_1756_0, i_8_329_1774_0, i_8_329_1775_0,
    i_8_329_1805_0, i_8_329_1809_0, i_8_329_1843_0, i_8_329_1873_0,
    i_8_329_1874_0, i_8_329_1882_0, i_8_329_1909_0, i_8_329_1982_0,
    i_8_329_1989_0, i_8_329_1991_0, i_8_329_1995_0, i_8_329_2052_0,
    i_8_329_2054_0, i_8_329_2065_0, i_8_329_2140_0, i_8_329_2145_0,
    i_8_329_2170_0, i_8_329_2171_0, i_8_329_2214_0, i_8_329_2215_0,
    i_8_329_2216_0, i_8_329_2233_0, i_8_329_2243_0;
  output o_8_329_0_0;
  assign o_8_329_0_0 = 0;
endmodule



// Benchmark "kernel_8_330" written by ABC on Sun Jul 19 10:08:46 2020

module kernel_8_330 ( 
    i_8_330_58_0, i_8_330_104_0, i_8_330_106_0, i_8_330_107_0,
    i_8_330_110_0, i_8_330_163_0, i_8_330_256_0, i_8_330_257_0,
    i_8_330_346_0, i_8_330_368_0, i_8_330_377_0, i_8_330_378_0,
    i_8_330_384_0, i_8_330_385_0, i_8_330_396_0, i_8_330_398_0,
    i_8_330_451_0, i_8_330_453_0, i_8_330_493_0, i_8_330_580_0,
    i_8_330_601_0, i_8_330_642_0, i_8_330_648_0, i_8_330_702_0,
    i_8_330_732_0, i_8_330_748_0, i_8_330_751_0, i_8_330_752_0,
    i_8_330_847_0, i_8_330_868_0, i_8_330_965_0, i_8_330_1058_0,
    i_8_330_1134_0, i_8_330_1135_0, i_8_330_1137_0, i_8_330_1138_0,
    i_8_330_1153_0, i_8_330_1192_0, i_8_330_1228_0, i_8_330_1233_0,
    i_8_330_1234_0, i_8_330_1273_0, i_8_330_1274_0, i_8_330_1314_0,
    i_8_330_1319_0, i_8_330_1324_0, i_8_330_1326_0, i_8_330_1328_0,
    i_8_330_1353_0, i_8_330_1408_0, i_8_330_1440_0, i_8_330_1486_0,
    i_8_330_1490_0, i_8_330_1506_0, i_8_330_1507_0, i_8_330_1533_0,
    i_8_330_1534_0, i_8_330_1551_0, i_8_330_1613_0, i_8_330_1614_0,
    i_8_330_1615_0, i_8_330_1616_0, i_8_330_1630_0, i_8_330_1652_0,
    i_8_330_1686_0, i_8_330_1688_0, i_8_330_1691_0, i_8_330_1710_0,
    i_8_330_1711_0, i_8_330_1712_0, i_8_330_1713_0, i_8_330_1714_0,
    i_8_330_1715_0, i_8_330_1810_0, i_8_330_1811_0, i_8_330_1812_0,
    i_8_330_1813_0, i_8_330_1831_0, i_8_330_1836_0, i_8_330_1837_0,
    i_8_330_1838_0, i_8_330_1839_0, i_8_330_1840_0, i_8_330_1841_0,
    i_8_330_1862_0, i_8_330_1885_0, i_8_330_1894_0, i_8_330_1895_0,
    i_8_330_1939_0, i_8_330_1986_0, i_8_330_2093_0, i_8_330_2099_0,
    i_8_330_2133_0, i_8_330_2134_0, i_8_330_2171_0, i_8_330_2260_0,
    i_8_330_2262_0, i_8_330_2263_0, i_8_330_2264_0, i_8_330_2298_0,
    o_8_330_0_0  );
  input  i_8_330_58_0, i_8_330_104_0, i_8_330_106_0, i_8_330_107_0,
    i_8_330_110_0, i_8_330_163_0, i_8_330_256_0, i_8_330_257_0,
    i_8_330_346_0, i_8_330_368_0, i_8_330_377_0, i_8_330_378_0,
    i_8_330_384_0, i_8_330_385_0, i_8_330_396_0, i_8_330_398_0,
    i_8_330_451_0, i_8_330_453_0, i_8_330_493_0, i_8_330_580_0,
    i_8_330_601_0, i_8_330_642_0, i_8_330_648_0, i_8_330_702_0,
    i_8_330_732_0, i_8_330_748_0, i_8_330_751_0, i_8_330_752_0,
    i_8_330_847_0, i_8_330_868_0, i_8_330_965_0, i_8_330_1058_0,
    i_8_330_1134_0, i_8_330_1135_0, i_8_330_1137_0, i_8_330_1138_0,
    i_8_330_1153_0, i_8_330_1192_0, i_8_330_1228_0, i_8_330_1233_0,
    i_8_330_1234_0, i_8_330_1273_0, i_8_330_1274_0, i_8_330_1314_0,
    i_8_330_1319_0, i_8_330_1324_0, i_8_330_1326_0, i_8_330_1328_0,
    i_8_330_1353_0, i_8_330_1408_0, i_8_330_1440_0, i_8_330_1486_0,
    i_8_330_1490_0, i_8_330_1506_0, i_8_330_1507_0, i_8_330_1533_0,
    i_8_330_1534_0, i_8_330_1551_0, i_8_330_1613_0, i_8_330_1614_0,
    i_8_330_1615_0, i_8_330_1616_0, i_8_330_1630_0, i_8_330_1652_0,
    i_8_330_1686_0, i_8_330_1688_0, i_8_330_1691_0, i_8_330_1710_0,
    i_8_330_1711_0, i_8_330_1712_0, i_8_330_1713_0, i_8_330_1714_0,
    i_8_330_1715_0, i_8_330_1810_0, i_8_330_1811_0, i_8_330_1812_0,
    i_8_330_1813_0, i_8_330_1831_0, i_8_330_1836_0, i_8_330_1837_0,
    i_8_330_1838_0, i_8_330_1839_0, i_8_330_1840_0, i_8_330_1841_0,
    i_8_330_1862_0, i_8_330_1885_0, i_8_330_1894_0, i_8_330_1895_0,
    i_8_330_1939_0, i_8_330_1986_0, i_8_330_2093_0, i_8_330_2099_0,
    i_8_330_2133_0, i_8_330_2134_0, i_8_330_2171_0, i_8_330_2260_0,
    i_8_330_2262_0, i_8_330_2263_0, i_8_330_2264_0, i_8_330_2298_0;
  output o_8_330_0_0;
  assign o_8_330_0_0 = ~((i_8_330_377_0 & ((~i_8_330_106_0 & ~i_8_330_1616_0 & i_8_330_1652_0) | (~i_8_330_257_0 & ~i_8_330_384_0 & i_8_330_751_0 & ~i_8_330_1137_0 & ~i_8_330_2134_0))) | (~i_8_330_1812_0 & ((~i_8_330_104_0 & ((~i_8_330_1135_0 & i_8_330_1506_0 & ~i_8_330_1551_0 & ~i_8_330_1810_0 & ~i_8_330_1813_0 & ~i_8_330_2133_0) | (~i_8_330_58_0 & ~i_8_330_385_0 & ~i_8_330_702_0 & i_8_330_1319_0 & ~i_8_330_1862_0 & ~i_8_330_2099_0 & ~i_8_330_2262_0))) | (~i_8_330_453_0 & ((~i_8_330_110_0 & ~i_8_330_1711_0 & ~i_8_330_1714_0 & ~i_8_330_1810_0 & i_8_330_1831_0 & ~i_8_330_2093_0) | (i_8_330_385_0 & i_8_330_493_0 & ~i_8_330_601_0 & i_8_330_1137_0 & ~i_8_330_1614_0 & ~i_8_330_2133_0))) | (~i_8_330_493_0 & ((~i_8_330_377_0 & i_8_330_1234_0 & ~i_8_330_1613_0 & ~i_8_330_1616_0 & ~i_8_330_1715_0 & ~i_8_330_1810_0 & ~i_8_330_1831_0 & i_8_330_1838_0) | (~i_8_330_106_0 & ~i_8_330_368_0 & ~i_8_330_1135_0 & ~i_8_330_1137_0 & ~i_8_330_1353_0 & ~i_8_330_1408_0 & ~i_8_330_1533_0 & i_8_330_1551_0 & ~i_8_330_1630_0 & ~i_8_330_1811_0 & ~i_8_330_2099_0 & ~i_8_330_2133_0 & ~i_8_330_2260_0))) | (~i_8_330_58_0 & ((~i_8_330_368_0 & ((~i_8_330_648_0 & i_8_330_1353_0 & i_8_330_1885_0 & ~i_8_330_1939_0) | (i_8_330_493_0 & ~i_8_330_1137_0 & i_8_330_1986_0 & ~i_8_330_2133_0))) | (~i_8_330_1138_0 & ~i_8_330_2099_0 & ((i_8_330_847_0 & i_8_330_1233_0 & i_8_330_1234_0 & ~i_8_330_1328_0 & ~i_8_330_1710_0 & ~i_8_330_1713_0) | (~i_8_330_256_0 & ~i_8_330_1058_0 & ~i_8_330_1135_0 & ~i_8_330_1314_0 & ~i_8_330_1615_0 & ~i_8_330_1630_0 & ~i_8_330_1714_0 & i_8_330_1810_0 & ~i_8_330_1862_0 & ~i_8_330_1939_0 & ~i_8_330_2262_0))))) | (~i_8_330_1551_0 & ((~i_8_330_748_0 & ((i_8_330_1233_0 & ~i_8_330_1353_0 & ~i_8_330_1614_0 & ~i_8_330_1712_0 & ~i_8_330_1810_0 & ~i_8_330_2099_0) | (~i_8_330_751_0 & i_8_330_1137_0 & i_8_330_1408_0 & ~i_8_330_2133_0))) | (~i_8_330_384_0 & ~i_8_330_847_0 & ~i_8_330_1228_0 & ~i_8_330_1274_0 & ~i_8_330_1534_0 & ~i_8_330_1714_0 & ~i_8_330_1715_0 & ~i_8_330_1811_0 & i_8_330_2093_0 & ~i_8_330_2264_0))) | (i_8_330_1058_0 & ((~i_8_330_1712_0 & ~i_8_330_1714_0 & i_8_330_1841_0) | (i_8_330_58_0 & ~i_8_330_1534_0 & ~i_8_330_1652_0 & ~i_8_330_1862_0 & ~i_8_330_2099_0 & ~i_8_330_2264_0))) | (~i_8_330_451_0 & ~i_8_330_648_0 & i_8_330_732_0 & ~i_8_330_1134_0 & i_8_330_1551_0 & ~i_8_330_2134_0) | (~i_8_330_1353_0 & ~i_8_330_1408_0 & ~i_8_330_107_0 & i_8_330_346_0 & i_8_330_1534_0 & ~i_8_330_1616_0 & ~i_8_330_1710_0 & ~i_8_330_2171_0) | (~i_8_330_601_0 & ~i_8_330_1810_0 & ~i_8_330_2260_0 & i_8_330_2298_0))) | (i_8_330_1058_0 & ((~i_8_330_1408_0 & i_8_330_1534_0 & ~i_8_330_1630_0 & ~i_8_330_1688_0 & ~i_8_330_1811_0 & ~i_8_330_2134_0) | (i_8_330_1353_0 & i_8_330_1652_0 & ~i_8_330_2171_0))) | (~i_8_330_1058_0 & ((~i_8_330_257_0 & ~i_8_330_368_0 & i_8_330_1233_0 & i_8_330_1314_0 & ~i_8_330_1710_0 & ~i_8_330_1811_0 & ~i_8_330_2171_0) | (~i_8_330_106_0 & ~i_8_330_384_0 & i_8_330_493_0 & ~i_8_330_1137_0 & i_8_330_1408_0 & ~i_8_330_1616_0 & ~i_8_330_1712_0 & ~i_8_330_1715_0 & ~i_8_330_2134_0 & ~i_8_330_2263_0))) | (~i_8_330_257_0 & ((~i_8_330_104_0 & ~i_8_330_1138_0 & i_8_330_1328_0 & ~i_8_330_1811_0 & ~i_8_330_1831_0 & ~i_8_330_1895_0) | (~i_8_330_107_0 & ~i_8_330_110_0 & ~i_8_330_453_0 & i_8_330_493_0 & ~i_8_330_732_0 & i_8_330_1353_0 & ~i_8_330_1614_0 & ~i_8_330_1616_0 & ~i_8_330_1986_0 & ~i_8_330_2099_0))) | (~i_8_330_1273_0 & ((~i_8_330_104_0 & i_8_330_110_0 & i_8_330_965_0 & i_8_330_1534_0 & ~i_8_330_2099_0) | (~i_8_330_107_0 & ~i_8_330_378_0 & ~i_8_330_752_0 & ~i_8_330_847_0 & ~i_8_330_965_0 & ~i_8_330_1192_0 & ~i_8_330_1228_0 & i_8_330_1507_0 & ~i_8_330_1614_0 & ~i_8_330_1630_0 & ~i_8_330_1688_0 & ~i_8_330_1714_0 & ~i_8_330_1840_0 & ~i_8_330_2133_0))) | (~i_8_330_378_0 & ((~i_8_330_451_0 & i_8_330_732_0 & i_8_330_1506_0 & ~i_8_330_1712_0) | (~i_8_330_107_0 & i_8_330_368_0 & i_8_330_493_0 & ~i_8_330_1353_0 & ~i_8_330_1616_0 & ~i_8_330_1813_0 & ~i_8_330_1986_0 & ~i_8_330_2099_0 & ~i_8_330_2264_0))) | (~i_8_330_385_0 & ((i_8_330_368_0 & ((~i_8_330_752_0 & i_8_330_1408_0 & i_8_330_1652_0 & ~i_8_330_2134_0) | (~i_8_330_107_0 & ~i_8_330_1613_0 & ~i_8_330_1691_0 & i_8_330_1862_0 & ~i_8_330_2263_0 & i_8_330_2264_0))) | (i_8_330_732_0 & ~i_8_330_1713_0 & ((~i_8_330_1134_0 & ~i_8_330_1135_0 & ~i_8_330_1615_0 & ~i_8_330_1710_0 & i_8_330_2133_0) | (~i_8_330_453_0 & ~i_8_330_601_0 & ~i_8_330_648_0 & ~i_8_330_847_0 & ~i_8_330_1712_0 & ~i_8_330_1714_0 & ~i_8_330_2171_0 & ~i_8_330_2262_0))) | (~i_8_330_1813_0 & ((~i_8_330_110_0 & ~i_8_330_384_0 & i_8_330_751_0 & ~i_8_330_1233_0 & ~i_8_330_1408_0 & ~i_8_330_1534_0 & ~i_8_330_1630_0 & ~i_8_330_2134_0) | (i_8_330_346_0 & ~i_8_330_748_0 & ~i_8_330_1134_0 & ~i_8_330_1507_0 & ~i_8_330_1533_0 & ~i_8_330_1712_0 & ~i_8_330_1836_0 & ~i_8_330_1862_0 & ~i_8_330_2262_0))) | (~i_8_330_1137_0 & ~i_8_330_1138_0 & i_8_330_1839_0 & ~i_8_330_2134_0))) | (~i_8_330_1813_0 & ((~i_8_330_58_0 & ~i_8_330_110_0 & ((~i_8_330_104_0 & ~i_8_330_451_0 & ~i_8_330_601_0 & i_8_330_1324_0 & ~i_8_330_1862_0 & ~i_8_330_2099_0 & ~i_8_330_2134_0) | (~i_8_330_1134_0 & i_8_330_1233_0 & ~i_8_330_1234_0 & i_8_330_1353_0 & ~i_8_330_1711_0 & ~i_8_330_2263_0))) | (~i_8_330_1810_0 & ((~i_8_330_107_0 & ((i_8_330_398_0 & ~i_8_330_1811_0) | (~i_8_330_104_0 & ~i_8_330_368_0 & ~i_8_330_748_0 & ~i_8_330_1234_0 & i_8_330_1274_0 & ~i_8_330_1408_0 & ~i_8_330_1712_0 & ~i_8_330_2133_0 & ~i_8_330_2263_0))) | (i_8_330_1274_0 & i_8_330_1507_0 & ~i_8_330_1986_0))) | (i_8_330_965_0 & ((i_8_330_163_0 & ~i_8_330_648_0 & ~i_8_330_1134_0 & ~i_8_330_1615_0 & ~i_8_330_1616_0 & ~i_8_330_2093_0) | (~i_8_330_106_0 & i_8_330_110_0 & ~i_8_330_1534_0 & ~i_8_330_1811_0 & ~i_8_330_2134_0))) | (i_8_330_346_0 & i_8_330_1506_0 & ~i_8_330_1713_0) | (~i_8_330_1811_0 & ~i_8_330_2099_0 & i_8_330_1234_0 & i_8_330_1324_0) | (~i_8_330_1134_0 & ~i_8_330_1137_0 & i_8_330_1408_0 & ~i_8_330_1486_0 & ~i_8_330_1862_0 & i_8_330_1885_0 & ~i_8_330_1986_0 & ~i_8_330_2133_0 & ~i_8_330_2262_0))) | (~i_8_330_107_0 & ((i_8_330_493_0 & i_8_330_1234_0 & ~i_8_330_1613_0 & ~i_8_330_1712_0 & ~i_8_330_2262_0) | (~i_8_330_965_0 & ~i_8_330_1534_0 & ~i_8_330_1616_0 & ~i_8_330_1652_0 & i_8_330_1688_0 & ~i_8_330_1715_0 & ~i_8_330_2171_0 & ~i_8_330_2264_0))) | (~i_8_330_1616_0 & ((~i_8_330_451_0 & ((~i_8_330_601_0 & ~i_8_330_648_0 & i_8_330_965_0 & i_8_330_1490_0) | (~i_8_330_368_0 & i_8_330_1326_0 & ~i_8_330_1534_0 & ~i_8_330_1630_0 & ~i_8_330_1839_0 & ~i_8_330_1885_0 & ~i_8_330_1894_0 & ~i_8_330_2263_0 & ~i_8_330_2264_0))) | (~i_8_330_702_0 & ((~i_8_330_104_0 & ~i_8_330_847_0 & ~i_8_330_965_0 & ~i_8_330_1135_0 & ~i_8_330_1274_0 & ~i_8_330_1614_0 & ~i_8_330_1712_0 & i_8_330_1837_0) | (i_8_330_1319_0 & i_8_330_1841_0 & ~i_8_330_2264_0))) | (~i_8_330_104_0 & ((~i_8_330_601_0 & ~i_8_330_868_0 & i_8_330_1192_0 & ~i_8_330_1314_0 & ~i_8_330_1711_0 & ~i_8_330_1811_0 & ~i_8_330_1895_0) | (~i_8_330_58_0 & ~i_8_330_398_0 & ~i_8_330_1137_0 & i_8_330_1273_0 & ~i_8_330_1353_0 & ~i_8_330_1712_0 & ~i_8_330_1714_0 & ~i_8_330_1715_0 & ~i_8_330_1837_0 & ~i_8_330_2171_0 & ~i_8_330_2262_0 & ~i_8_330_1838_0 & ~i_8_330_1986_0))))) | (~i_8_330_648_0 & ((~i_8_330_58_0 & ~i_8_330_1138_0 & ~i_8_330_1319_0 & ~i_8_330_1507_0 & ~i_8_330_1711_0 & i_8_330_1836_0 & ~i_8_330_2099_0) | (~i_8_330_106_0 & i_8_330_110_0 & ~i_8_330_384_0 & ~i_8_330_1811_0 & ~i_8_330_2134_0 & ~i_8_330_1234_0 & i_8_330_1551_0))) | (i_8_330_110_0 & i_8_330_1838_0 & ((~i_8_330_752_0 & i_8_330_1534_0) | (~i_8_330_368_0 & ~i_8_330_1486_0 & ~i_8_330_2099_0))) | (~i_8_330_2262_0 & ((~i_8_330_106_0 & i_8_330_1353_0 & ~i_8_330_1986_0 & ((~i_8_330_384_0 & ~i_8_330_453_0 & ~i_8_330_702_0 & ~i_8_330_847_0 & i_8_330_1408_0 & ~i_8_330_1715_0) | (~i_8_330_1615_0 & i_8_330_2298_0))) | (i_8_330_732_0 & ~i_8_330_1810_0 & ((i_8_330_702_0 & i_8_330_1233_0) | (~i_8_330_453_0 & ~i_8_330_847_0 & i_8_330_1533_0 & ~i_8_330_1614_0 & ~i_8_330_1712_0))) | (~i_8_330_256_0 & ~i_8_330_1137_0 & i_8_330_1506_0 & ~i_8_330_1534_0 & ~i_8_330_1713_0 & ~i_8_330_1811_0 & ~i_8_330_2133_0 & ~i_8_330_2134_0))) | (~i_8_330_106_0 & ((~i_8_330_601_0 & i_8_330_1326_0 & ~i_8_330_1710_0 & i_8_330_1839_0) | (~i_8_330_1490_0 & ~i_8_330_1862_0 & i_8_330_1895_0 & ~i_8_330_2099_0))) | (~i_8_330_1613_0 & ((~i_8_330_384_0 & ~i_8_330_1713_0 & ~i_8_330_1715_0 & ((~i_8_330_256_0 & i_8_330_752_0 & i_8_330_1551_0 & ~i_8_330_1615_0 & ~i_8_330_2133_0) | (~i_8_330_163_0 & ~i_8_330_453_0 & ~i_8_330_1135_0 & ~i_8_330_1137_0 & i_8_330_1234_0 & i_8_330_1353_0 & i_8_330_1486_0 & ~i_8_330_1490_0 & ~i_8_330_1839_0 & ~i_8_330_2298_0))) | (~i_8_330_256_0 & ~i_8_330_702_0 & ((~i_8_330_58_0 & ~i_8_330_396_0 & ~i_8_330_601_0 & ~i_8_330_748_0 & i_8_330_1233_0 & ~i_8_330_1328_0 & ~i_8_330_2260_0) | (~i_8_330_847_0 & ~i_8_330_1614_0 & i_8_330_1710_0 & i_8_330_2262_0))) | (i_8_330_1652_0 & ~i_8_330_1710_0 & ~i_8_330_1811_0 & i_8_330_1885_0))) | (~i_8_330_368_0 & ((~i_8_330_58_0 & ((i_8_330_1324_0 & ~i_8_330_1630_0 & i_8_330_2093_0) | (i_8_330_1652_0 & ~i_8_330_2171_0 & i_8_330_752_0 & ~i_8_330_1490_0))) | (i_8_330_346_0 & ~i_8_330_1134_0 & ~i_8_330_1234_0 & ~i_8_330_1551_0 & ~i_8_330_1811_0 & ~i_8_330_1986_0 & ~i_8_330_2093_0 & ~i_8_330_2099_0))) | (~i_8_330_868_0 & ((i_8_330_451_0 & ~i_8_330_1153_0 & i_8_330_1490_0 & ~i_8_330_1711_0 & ~i_8_330_1712_0) | (~i_8_330_748_0 & i_8_330_1319_0 & i_8_330_1652_0 & ~i_8_330_1715_0 & ~i_8_330_1810_0 & ~i_8_330_2093_0 & ~i_8_330_2298_0))) | (i_8_330_1652_0 & ((i_8_330_493_0 & i_8_330_748_0 & i_8_330_752_0 & ~i_8_330_1710_0 & ~i_8_330_1715_0) | (~i_8_330_601_0 & i_8_330_1840_0 & ~i_8_330_1862_0 & ~i_8_330_2134_0))) | (~i_8_330_1712_0 & ((i_8_330_1534_0 & ~i_8_330_1810_0 & i_8_330_1839_0) | (~i_8_330_346_0 & ~i_8_330_752_0 & ~i_8_330_1138_0 & i_8_330_1841_0 & ~i_8_330_2171_0))) | (i_8_330_1353_0 & i_8_330_1686_0 & i_8_330_1986_0) | (i_8_330_396_0 & ~i_8_330_1314_0 & ~i_8_330_1614_0 & ~i_8_330_1711_0 & ~i_8_330_2099_0));
endmodule



// Benchmark "kernel_8_331" written by ABC on Sun Jul 19 10:08:48 2020

module kernel_8_331 ( 
    i_8_331_48_0, i_8_331_63_0, i_8_331_64_0, i_8_331_121_0, i_8_331_152_0,
    i_8_331_171_0, i_8_331_219_0, i_8_331_226_0, i_8_331_294_0,
    i_8_331_295_0, i_8_331_304_0, i_8_331_324_0, i_8_331_340_0,
    i_8_331_354_0, i_8_331_374_0, i_8_331_382_0, i_8_331_384_0,
    i_8_331_385_0, i_8_331_430_0, i_8_331_489_0, i_8_331_492_0,
    i_8_331_552_0, i_8_331_554_0, i_8_331_583_0, i_8_331_591_0,
    i_8_331_592_0, i_8_331_600_0, i_8_331_642_0, i_8_331_655_0,
    i_8_331_661_0, i_8_331_662_0, i_8_331_687_0, i_8_331_710_0,
    i_8_331_733_0, i_8_331_750_0, i_8_331_795_0, i_8_331_798_0,
    i_8_331_879_0, i_8_331_881_0, i_8_331_926_0, i_8_331_935_0,
    i_8_331_990_0, i_8_331_1032_0, i_8_331_1110_0, i_8_331_1152_0,
    i_8_331_1170_0, i_8_331_1188_0, i_8_331_1224_0, i_8_331_1257_0,
    i_8_331_1258_0, i_8_331_1259_0, i_8_331_1266_0, i_8_331_1267_0,
    i_8_331_1272_0, i_8_331_1276_0, i_8_331_1284_0, i_8_331_1285_0,
    i_8_331_1286_0, i_8_331_1330_0, i_8_331_1371_0, i_8_331_1375_0,
    i_8_331_1389_0, i_8_331_1443_0, i_8_331_1455_0, i_8_331_1552_0,
    i_8_331_1554_0, i_8_331_1607_0, i_8_331_1633_0, i_8_331_1635_0,
    i_8_331_1647_0, i_8_331_1653_0, i_8_331_1678_0, i_8_331_1686_0,
    i_8_331_1723_0, i_8_331_1730_0, i_8_331_1736_0, i_8_331_1747_0,
    i_8_331_1751_0, i_8_331_1777_0, i_8_331_1778_0, i_8_331_1869_0,
    i_8_331_1950_0, i_8_331_2013_0, i_8_331_2048_0, i_8_331_2056_0,
    i_8_331_2078_0, i_8_331_2095_0, i_8_331_2097_0, i_8_331_2112_0,
    i_8_331_2114_0, i_8_331_2131_0, i_8_331_2142_0, i_8_331_2157_0,
    i_8_331_2176_0, i_8_331_2185_0, i_8_331_2194_0, i_8_331_2222_0,
    i_8_331_2223_0, i_8_331_2249_0, i_8_331_2266_0,
    o_8_331_0_0  );
  input  i_8_331_48_0, i_8_331_63_0, i_8_331_64_0, i_8_331_121_0,
    i_8_331_152_0, i_8_331_171_0, i_8_331_219_0, i_8_331_226_0,
    i_8_331_294_0, i_8_331_295_0, i_8_331_304_0, i_8_331_324_0,
    i_8_331_340_0, i_8_331_354_0, i_8_331_374_0, i_8_331_382_0,
    i_8_331_384_0, i_8_331_385_0, i_8_331_430_0, i_8_331_489_0,
    i_8_331_492_0, i_8_331_552_0, i_8_331_554_0, i_8_331_583_0,
    i_8_331_591_0, i_8_331_592_0, i_8_331_600_0, i_8_331_642_0,
    i_8_331_655_0, i_8_331_661_0, i_8_331_662_0, i_8_331_687_0,
    i_8_331_710_0, i_8_331_733_0, i_8_331_750_0, i_8_331_795_0,
    i_8_331_798_0, i_8_331_879_0, i_8_331_881_0, i_8_331_926_0,
    i_8_331_935_0, i_8_331_990_0, i_8_331_1032_0, i_8_331_1110_0,
    i_8_331_1152_0, i_8_331_1170_0, i_8_331_1188_0, i_8_331_1224_0,
    i_8_331_1257_0, i_8_331_1258_0, i_8_331_1259_0, i_8_331_1266_0,
    i_8_331_1267_0, i_8_331_1272_0, i_8_331_1276_0, i_8_331_1284_0,
    i_8_331_1285_0, i_8_331_1286_0, i_8_331_1330_0, i_8_331_1371_0,
    i_8_331_1375_0, i_8_331_1389_0, i_8_331_1443_0, i_8_331_1455_0,
    i_8_331_1552_0, i_8_331_1554_0, i_8_331_1607_0, i_8_331_1633_0,
    i_8_331_1635_0, i_8_331_1647_0, i_8_331_1653_0, i_8_331_1678_0,
    i_8_331_1686_0, i_8_331_1723_0, i_8_331_1730_0, i_8_331_1736_0,
    i_8_331_1747_0, i_8_331_1751_0, i_8_331_1777_0, i_8_331_1778_0,
    i_8_331_1869_0, i_8_331_1950_0, i_8_331_2013_0, i_8_331_2048_0,
    i_8_331_2056_0, i_8_331_2078_0, i_8_331_2095_0, i_8_331_2097_0,
    i_8_331_2112_0, i_8_331_2114_0, i_8_331_2131_0, i_8_331_2142_0,
    i_8_331_2157_0, i_8_331_2176_0, i_8_331_2185_0, i_8_331_2194_0,
    i_8_331_2222_0, i_8_331_2223_0, i_8_331_2249_0, i_8_331_2266_0;
  output o_8_331_0_0;
  assign o_8_331_0_0 = ~((~i_8_331_121_0 & ((~i_8_331_64_0 & i_8_331_382_0 & ~i_8_331_430_0 & ~i_8_331_687_0 & ~i_8_331_1257_0 & ~i_8_331_1258_0 & ~i_8_331_1276_0 & ~i_8_331_1686_0 & ~i_8_331_1730_0 & ~i_8_331_2112_0) | (~i_8_331_171_0 & ~i_8_331_226_0 & i_8_331_552_0 & ~i_8_331_1188_0 & ~i_8_331_1375_0 & ~i_8_331_1455_0 & ~i_8_331_2114_0 & ~i_8_331_2157_0 & ~i_8_331_2249_0))) | (~i_8_331_554_0 & ((~i_8_331_385_0 & i_8_331_489_0 & ~i_8_331_1284_0 & ~i_8_331_1371_0 & i_8_331_1552_0 & ~i_8_331_1723_0 & ~i_8_331_1747_0 & ~i_8_331_1751_0) | (~i_8_331_294_0 & ~i_8_331_583_0 & ~i_8_331_1257_0 & ~i_8_331_1286_0 & ~i_8_331_1389_0 & i_8_331_1554_0 & ~i_8_331_1778_0 & ~i_8_331_2056_0 & ~i_8_331_2078_0 & ~i_8_331_2194_0 & ~i_8_331_2223_0))) | (~i_8_331_294_0 & ((~i_8_331_63_0 & ~i_8_331_489_0 & ~i_8_331_592_0 & ~i_8_331_798_0 & ~i_8_331_1259_0 & ~i_8_331_1869_0 & ~i_8_331_2112_0) | (~i_8_331_384_0 & ~i_8_331_385_0 & ~i_8_331_430_0 & ~i_8_331_926_0 & ~i_8_331_935_0 & ~i_8_331_1170_0 & ~i_8_331_1257_0 & ~i_8_331_1258_0 & ~i_8_331_1371_0 & ~i_8_331_2056_0 & ~i_8_331_2142_0))) | (~i_8_331_1443_0 & ((~i_8_331_171_0 & ~i_8_331_1286_0 & ((i_8_331_226_0 & ~i_8_331_655_0 & ~i_8_331_662_0 & i_8_331_2142_0) | (~i_8_331_384_0 & ~i_8_331_795_0 & ~i_8_331_926_0 & ~i_8_331_1170_0 & ~i_8_331_1258_0 & ~i_8_331_1276_0 & ~i_8_331_1455_0 & ~i_8_331_1730_0 & ~i_8_331_2185_0))) | (~i_8_331_385_0 & ~i_8_331_881_0 & ((~i_8_331_382_0 & ~i_8_331_1224_0 & ~i_8_331_1276_0 & i_8_331_1285_0 & ~i_8_331_1455_0 & ~i_8_331_1751_0 & ~i_8_331_2114_0) | (~i_8_331_64_0 & ~i_8_331_384_0 & ~i_8_331_592_0 & ~i_8_331_655_0 & ~i_8_331_879_0 & ~i_8_331_1686_0 & ~i_8_331_2223_0 & ~i_8_331_2266_0))) | (~i_8_331_926_0 & ~i_8_331_1224_0 & ~i_8_331_1259_0 & i_8_331_1723_0))) | (~i_8_331_171_0 & ((~i_8_331_295_0 & i_8_331_661_0 & ~i_8_331_798_0 & ~i_8_331_935_0 & i_8_331_1266_0) | (i_8_331_219_0 & ~i_8_331_600_0 & ~i_8_331_687_0 & ~i_8_331_795_0 & ~i_8_331_926_0 & ~i_8_331_1032_0 & ~i_8_331_2185_0))) | (~i_8_331_1258_0 & ((~i_8_331_63_0 & ((~i_8_331_64_0 & ~i_8_331_1257_0 & ~i_8_331_1455_0 & i_8_331_1777_0 & ~i_8_331_2112_0) | (~i_8_331_385_0 & ~i_8_331_489_0 & ~i_8_331_583_0 & ~i_8_331_795_0 & ~i_8_331_935_0 & ~i_8_331_1032_0 & ~i_8_331_1647_0 & ~i_8_331_2114_0))) | (~i_8_331_64_0 & ((~i_8_331_935_0 & ((~i_8_331_304_0 & ~i_8_331_492_0 & ~i_8_331_591_0 & ~i_8_331_750_0 & ~i_8_331_1224_0 & ~i_8_331_2056_0 & ~i_8_331_2112_0) | (i_8_331_655_0 & ~i_8_331_1371_0 & ~i_8_331_1375_0 & ~i_8_331_1455_0 & ~i_8_331_2194_0 & ~i_8_331_2223_0))) | (~i_8_331_385_0 & ~i_8_331_430_0 & ~i_8_331_926_0 & ~i_8_331_1032_0 & ~i_8_331_1272_0 & ~i_8_331_1285_0 & ~i_8_331_1778_0 & ~i_8_331_2223_0))) | (~i_8_331_295_0 & ~i_8_331_662_0 & ~i_8_331_1224_0 & ~i_8_331_1389_0 & i_8_331_2078_0 & ~i_8_331_2194_0) | (~i_8_331_489_0 & ~i_8_331_733_0 & ~i_8_331_798_0 & ~i_8_331_879_0 & ~i_8_331_1170_0 & ~i_8_331_1259_0 & ~i_8_331_2131_0 & ~i_8_331_2222_0))) | (~i_8_331_492_0 & ((~i_8_331_63_0 & ~i_8_331_219_0 & ~i_8_331_295_0 & ~i_8_331_710_0 & ~i_8_331_926_0 & ~i_8_331_1032_0 & ~i_8_331_1170_0 & ~i_8_331_1259_0 & ~i_8_331_1375_0 & ~i_8_331_1869_0 & ~i_8_331_1950_0 & ~i_8_331_2176_0 & ~i_8_331_2223_0) | (~i_8_331_1224_0 & i_8_331_1267_0 & i_8_331_1950_0 & ~i_8_331_2249_0))) | (~i_8_331_583_0 & ((~i_8_331_600_0 & ((~i_8_331_64_0 & ~i_8_331_552_0 & ~i_8_331_591_0 & ~i_8_331_642_0 & ~i_8_331_926_0 & ~i_8_331_1170_0 & ~i_8_331_1276_0 & ~i_8_331_1284_0 & ~i_8_331_1285_0 & ~i_8_331_1950_0 & ~i_8_331_2114_0) | (i_8_331_340_0 & i_8_331_385_0 & i_8_331_1258_0 & i_8_331_1285_0 & ~i_8_331_1455_0 & ~i_8_331_1552_0 & ~i_8_331_1723_0 & ~i_8_331_2222_0))) | (~i_8_331_295_0 & ~i_8_331_1389_0 & i_8_331_1607_0 & ~i_8_331_1736_0 & ~i_8_331_1869_0 & ~i_8_331_2095_0 & ~i_8_331_2223_0))) | (~i_8_331_295_0 & ((~i_8_331_430_0 & ~i_8_331_1224_0 & i_8_331_1635_0) | (~i_8_331_661_0 & ~i_8_331_795_0 & ~i_8_331_1330_0 & i_8_331_1778_0 & ~i_8_331_1869_0 & ~i_8_331_2142_0))) | (~i_8_331_354_0 & ~i_8_331_1257_0 & ~i_8_331_1330_0 & i_8_331_1443_0 & i_8_331_1751_0 & ~i_8_331_2048_0 & ~i_8_331_2056_0) | (i_8_331_382_0 & ~i_8_331_1285_0 & i_8_331_2097_0 & i_8_331_2266_0));
endmodule



// Benchmark "kernel_8_332" written by ABC on Sun Jul 19 10:08:49 2020

module kernel_8_332 ( 
    i_8_332_12_0, i_8_332_30_0, i_8_332_72_0, i_8_332_82_0, i_8_332_83_0,
    i_8_332_119_0, i_8_332_135_0, i_8_332_139_0, i_8_332_153_0,
    i_8_332_156_0, i_8_332_201_0, i_8_332_202_0, i_8_332_207_0,
    i_8_332_216_0, i_8_332_219_0, i_8_332_220_0, i_8_332_267_0,
    i_8_332_282_0, i_8_332_324_0, i_8_332_333_0, i_8_332_343_0,
    i_8_332_373_0, i_8_332_384_0, i_8_332_432_0, i_8_332_495_0,
    i_8_332_498_0, i_8_332_533_0, i_8_332_550_0, i_8_332_552_0,
    i_8_332_585_0, i_8_332_595_0, i_8_332_609_0, i_8_332_612_0,
    i_8_332_621_0, i_8_332_636_0, i_8_332_637_0, i_8_332_669_0,
    i_8_332_720_0, i_8_332_774_0, i_8_332_775_0, i_8_332_777_0,
    i_8_332_804_0, i_8_332_821_0, i_8_332_823_0, i_8_332_847_0,
    i_8_332_867_0, i_8_332_875_0, i_8_332_876_0, i_8_332_891_0,
    i_8_332_932_0, i_8_332_963_0, i_8_332_965_0, i_8_332_972_0,
    i_8_332_981_0, i_8_332_991_0, i_8_332_994_0, i_8_332_1008_0,
    i_8_332_1009_0, i_8_332_1011_0, i_8_332_1083_0, i_8_332_1129_0,
    i_8_332_1145_0, i_8_332_1155_0, i_8_332_1171_0, i_8_332_1245_0,
    i_8_332_1255_0, i_8_332_1270_0, i_8_332_1275_0, i_8_332_1288_0,
    i_8_332_1296_0, i_8_332_1312_0, i_8_332_1341_0, i_8_332_1342_0,
    i_8_332_1428_0, i_8_332_1432_0, i_8_332_1443_0, i_8_332_1516_0,
    i_8_332_1521_0, i_8_332_1524_0, i_8_332_1548_0, i_8_332_1549_0,
    i_8_332_1611_0, i_8_332_1669_0, i_8_332_1675_0, i_8_332_1705_0,
    i_8_332_1775_0, i_8_332_1800_0, i_8_332_1801_0, i_8_332_1839_0,
    i_8_332_1919_0, i_8_332_1945_0, i_8_332_1999_0, i_8_332_2038_0,
    i_8_332_2107_0, i_8_332_2117_0, i_8_332_2146_0, i_8_332_2269_0,
    i_8_332_2281_0, i_8_332_2286_0, i_8_332_2291_0,
    o_8_332_0_0  );
  input  i_8_332_12_0, i_8_332_30_0, i_8_332_72_0, i_8_332_82_0,
    i_8_332_83_0, i_8_332_119_0, i_8_332_135_0, i_8_332_139_0,
    i_8_332_153_0, i_8_332_156_0, i_8_332_201_0, i_8_332_202_0,
    i_8_332_207_0, i_8_332_216_0, i_8_332_219_0, i_8_332_220_0,
    i_8_332_267_0, i_8_332_282_0, i_8_332_324_0, i_8_332_333_0,
    i_8_332_343_0, i_8_332_373_0, i_8_332_384_0, i_8_332_432_0,
    i_8_332_495_0, i_8_332_498_0, i_8_332_533_0, i_8_332_550_0,
    i_8_332_552_0, i_8_332_585_0, i_8_332_595_0, i_8_332_609_0,
    i_8_332_612_0, i_8_332_621_0, i_8_332_636_0, i_8_332_637_0,
    i_8_332_669_0, i_8_332_720_0, i_8_332_774_0, i_8_332_775_0,
    i_8_332_777_0, i_8_332_804_0, i_8_332_821_0, i_8_332_823_0,
    i_8_332_847_0, i_8_332_867_0, i_8_332_875_0, i_8_332_876_0,
    i_8_332_891_0, i_8_332_932_0, i_8_332_963_0, i_8_332_965_0,
    i_8_332_972_0, i_8_332_981_0, i_8_332_991_0, i_8_332_994_0,
    i_8_332_1008_0, i_8_332_1009_0, i_8_332_1011_0, i_8_332_1083_0,
    i_8_332_1129_0, i_8_332_1145_0, i_8_332_1155_0, i_8_332_1171_0,
    i_8_332_1245_0, i_8_332_1255_0, i_8_332_1270_0, i_8_332_1275_0,
    i_8_332_1288_0, i_8_332_1296_0, i_8_332_1312_0, i_8_332_1341_0,
    i_8_332_1342_0, i_8_332_1428_0, i_8_332_1432_0, i_8_332_1443_0,
    i_8_332_1516_0, i_8_332_1521_0, i_8_332_1524_0, i_8_332_1548_0,
    i_8_332_1549_0, i_8_332_1611_0, i_8_332_1669_0, i_8_332_1675_0,
    i_8_332_1705_0, i_8_332_1775_0, i_8_332_1800_0, i_8_332_1801_0,
    i_8_332_1839_0, i_8_332_1919_0, i_8_332_1945_0, i_8_332_1999_0,
    i_8_332_2038_0, i_8_332_2107_0, i_8_332_2117_0, i_8_332_2146_0,
    i_8_332_2269_0, i_8_332_2281_0, i_8_332_2286_0, i_8_332_2291_0;
  output o_8_332_0_0;
  assign o_8_332_0_0 = ~((~i_8_332_12_0 & ((~i_8_332_119_0 & ~i_8_332_201_0 & ~i_8_332_432_0 & ~i_8_332_495_0 & ~i_8_332_720_0 & ~i_8_332_821_0 & ~i_8_332_823_0 & ~i_8_332_1521_0 & ~i_8_332_1919_0 & ~i_8_332_1999_0) | (~i_8_332_83_0 & ~i_8_332_219_0 & ~i_8_332_891_0 & ~i_8_332_1129_0 & ~i_8_332_1145_0 & ~i_8_332_1288_0 & ~i_8_332_1516_0 & ~i_8_332_2286_0))) | (~i_8_332_202_0 & ((~i_8_332_201_0 & ((~i_8_332_207_0 & ~i_8_332_282_0 & ~i_8_332_495_0 & ~i_8_332_991_0 & ~i_8_332_1009_0 & ~i_8_332_1341_0) | (~i_8_332_875_0 & ~i_8_332_965_0 & ~i_8_332_1145_0 & ~i_8_332_1255_0 & ~i_8_332_1342_0 & i_8_332_2146_0))) | (~i_8_332_2286_0 & ((~i_8_332_219_0 & ~i_8_332_621_0 & ~i_8_332_875_0 & ~i_8_332_932_0 & ~i_8_332_1129_0 & ~i_8_332_1270_0) | (~i_8_332_153_0 & ~i_8_332_282_0 & ~i_8_332_1008_0 & ~i_8_332_1443_0 & ~i_8_332_2117_0 & ~i_8_332_2281_0))))) | (~i_8_332_153_0 & ~i_8_332_774_0 & ((~i_8_332_720_0 & ~i_8_332_991_0 & ~i_8_332_1009_0 & ~i_8_332_1521_0 & ~i_8_332_1675_0 & ~i_8_332_2107_0 & ~i_8_332_2117_0) | (~i_8_332_156_0 & ~i_8_332_282_0 & ~i_8_332_384_0 & ~i_8_332_550_0 & ~i_8_332_867_0 & ~i_8_332_891_0 & ~i_8_332_981_0 & ~i_8_332_1145_0 & ~i_8_332_1155_0 & ~i_8_332_1516_0 & ~i_8_332_1705_0 & ~i_8_332_2286_0))) | (~i_8_332_267_0 & ((~i_8_332_83_0 & ~i_8_332_432_0 & ~i_8_332_495_0 & ~i_8_332_804_0 & ~i_8_332_1011_0 & ~i_8_332_1083_0 & ~i_8_332_1270_0 & ~i_8_332_1705_0 & i_8_332_1999_0) | (~i_8_332_282_0 & ~i_8_332_621_0 & ~i_8_332_891_0 & i_8_332_1296_0 & ~i_8_332_1521_0 & i_8_332_2038_0 & i_8_332_2269_0))) | (~i_8_332_343_0 & ~i_8_332_932_0 & ((~i_8_332_156_0 & ~i_8_332_495_0 & ~i_8_332_994_0 & ~i_8_332_1275_0 & ~i_8_332_1775_0 & ~i_8_332_1801_0) | (~i_8_332_324_0 & ~i_8_332_981_0 & ~i_8_332_1008_0 & ~i_8_332_2269_0 & ~i_8_332_2286_0))) | (~i_8_332_156_0 & ((~i_8_332_621_0 & ~i_8_332_821_0 & ~i_8_332_1009_0 & ~i_8_332_1083_0 & ~i_8_332_1342_0) | (~i_8_332_82_0 & ~i_8_332_119_0 & ~i_8_332_333_0 & ~i_8_332_533_0 & ~i_8_332_720_0 & ~i_8_332_2269_0))) | (~i_8_332_495_0 & ((~i_8_332_550_0 & ~i_8_332_981_0 & ~i_8_332_1171_0 & ~i_8_332_1275_0 & i_8_332_1296_0) | (i_8_332_585_0 & ~i_8_332_775_0 & ~i_8_332_965_0 & ~i_8_332_1083_0 & ~i_8_332_2269_0))) | (~i_8_332_1342_0 & ((~i_8_332_135_0 & ~i_8_332_595_0 & ~i_8_332_609_0 & ~i_8_332_612_0 & ~i_8_332_669_0 & ~i_8_332_1083_0 & ~i_8_332_1312_0 & ~i_8_332_1443_0 & ~i_8_332_1611_0) | (~i_8_332_1516_0 & ~i_8_332_1800_0 & ~i_8_332_1801_0))) | (i_8_332_82_0 & i_8_332_774_0 & ~i_8_332_821_0 & ~i_8_332_963_0 & ~i_8_332_1341_0 & i_8_332_1800_0) | (i_8_332_432_0 & i_8_332_1171_0 & i_8_332_2107_0));
endmodule



// Benchmark "kernel_8_333" written by ABC on Sun Jul 19 10:08:50 2020

module kernel_8_333 ( 
    i_8_333_34_0, i_8_333_35_0, i_8_333_50_0, i_8_333_53_0, i_8_333_60_0,
    i_8_333_65_0, i_8_333_95_0, i_8_333_125_0, i_8_333_143_0,
    i_8_333_169_0, i_8_333_233_0, i_8_333_242_0, i_8_333_278_0,
    i_8_333_347_0, i_8_333_350_0, i_8_333_360_0, i_8_333_365_0,
    i_8_333_401_0, i_8_333_431_0, i_8_333_454_0, i_8_333_455_0,
    i_8_333_553_0, i_8_333_557_0, i_8_333_581_0, i_8_333_590_0,
    i_8_333_607_0, i_8_333_613_0, i_8_333_614_0, i_8_333_638_0,
    i_8_333_656_0, i_8_333_661_0, i_8_333_662_0, i_8_333_679_0,
    i_8_333_680_0, i_8_333_697_0, i_8_333_700_0, i_8_333_701_0,
    i_8_333_707_0, i_8_333_711_0, i_8_333_731_0, i_8_333_759_0,
    i_8_333_779_0, i_8_333_782_0, i_8_333_793_0, i_8_333_799_0,
    i_8_333_844_0, i_8_333_969_0, i_8_333_1030_0, i_8_333_1103_0,
    i_8_333_1129_0, i_8_333_1146_0, i_8_333_1154_0, i_8_333_1157_0,
    i_8_333_1172_0, i_8_333_1175_0, i_8_333_1264_0, i_8_333_1265_0,
    i_8_333_1274_0, i_8_333_1292_0, i_8_333_1305_0, i_8_333_1373_0,
    i_8_333_1411_0, i_8_333_1412_0, i_8_333_1472_0, i_8_333_1493_0,
    i_8_333_1508_0, i_8_333_1525_0, i_8_333_1562_0, i_8_333_1607_0,
    i_8_333_1609_0, i_8_333_1628_0, i_8_333_1648_0, i_8_333_1649_0,
    i_8_333_1655_0, i_8_333_1664_0, i_8_333_1679_0, i_8_333_1698_0,
    i_8_333_1778_0, i_8_333_1803_0, i_8_333_1819_0, i_8_333_1823_0,
    i_8_333_1832_0, i_8_333_1854_0, i_8_333_1859_0, i_8_333_1886_0,
    i_8_333_1906_0, i_8_333_1967_0, i_8_333_1984_0, i_8_333_1985_0,
    i_8_333_1996_0, i_8_333_2018_0, i_8_333_2096_0, i_8_333_2146_0,
    i_8_333_2156_0, i_8_333_2183_0, i_8_333_2210_0, i_8_333_2219_0,
    i_8_333_2227_0, i_8_333_2244_0, i_8_333_2276_0,
    o_8_333_0_0  );
  input  i_8_333_34_0, i_8_333_35_0, i_8_333_50_0, i_8_333_53_0,
    i_8_333_60_0, i_8_333_65_0, i_8_333_95_0, i_8_333_125_0, i_8_333_143_0,
    i_8_333_169_0, i_8_333_233_0, i_8_333_242_0, i_8_333_278_0,
    i_8_333_347_0, i_8_333_350_0, i_8_333_360_0, i_8_333_365_0,
    i_8_333_401_0, i_8_333_431_0, i_8_333_454_0, i_8_333_455_0,
    i_8_333_553_0, i_8_333_557_0, i_8_333_581_0, i_8_333_590_0,
    i_8_333_607_0, i_8_333_613_0, i_8_333_614_0, i_8_333_638_0,
    i_8_333_656_0, i_8_333_661_0, i_8_333_662_0, i_8_333_679_0,
    i_8_333_680_0, i_8_333_697_0, i_8_333_700_0, i_8_333_701_0,
    i_8_333_707_0, i_8_333_711_0, i_8_333_731_0, i_8_333_759_0,
    i_8_333_779_0, i_8_333_782_0, i_8_333_793_0, i_8_333_799_0,
    i_8_333_844_0, i_8_333_969_0, i_8_333_1030_0, i_8_333_1103_0,
    i_8_333_1129_0, i_8_333_1146_0, i_8_333_1154_0, i_8_333_1157_0,
    i_8_333_1172_0, i_8_333_1175_0, i_8_333_1264_0, i_8_333_1265_0,
    i_8_333_1274_0, i_8_333_1292_0, i_8_333_1305_0, i_8_333_1373_0,
    i_8_333_1411_0, i_8_333_1412_0, i_8_333_1472_0, i_8_333_1493_0,
    i_8_333_1508_0, i_8_333_1525_0, i_8_333_1562_0, i_8_333_1607_0,
    i_8_333_1609_0, i_8_333_1628_0, i_8_333_1648_0, i_8_333_1649_0,
    i_8_333_1655_0, i_8_333_1664_0, i_8_333_1679_0, i_8_333_1698_0,
    i_8_333_1778_0, i_8_333_1803_0, i_8_333_1819_0, i_8_333_1823_0,
    i_8_333_1832_0, i_8_333_1854_0, i_8_333_1859_0, i_8_333_1886_0,
    i_8_333_1906_0, i_8_333_1967_0, i_8_333_1984_0, i_8_333_1985_0,
    i_8_333_1996_0, i_8_333_2018_0, i_8_333_2096_0, i_8_333_2146_0,
    i_8_333_2156_0, i_8_333_2183_0, i_8_333_2210_0, i_8_333_2219_0,
    i_8_333_2227_0, i_8_333_2244_0, i_8_333_2276_0;
  output o_8_333_0_0;
  assign o_8_333_0_0 = 0;
endmodule



// Benchmark "kernel_8_334" written by ABC on Sun Jul 19 10:08:52 2020

module kernel_8_334 ( 
    i_8_334_53_0, i_8_334_86_0, i_8_334_87_0, i_8_334_97_0, i_8_334_139_0,
    i_8_334_230_0, i_8_334_255_0, i_8_334_258_0, i_8_334_260_0,
    i_8_334_327_0, i_8_334_328_0, i_8_334_329_0, i_8_334_362_0,
    i_8_334_363_0, i_8_334_457_0, i_8_334_462_0, i_8_334_463_0,
    i_8_334_464_0, i_8_334_466_0, i_8_334_474_0, i_8_334_476_0,
    i_8_334_500_0, i_8_334_523_0, i_8_334_526_0, i_8_334_528_0,
    i_8_334_530_0, i_8_334_555_0, i_8_334_617_0, i_8_334_660_0,
    i_8_334_661_0, i_8_334_663_0, i_8_334_672_0, i_8_334_674_0,
    i_8_334_682_0, i_8_334_732_0, i_8_334_762_0, i_8_334_763_0,
    i_8_334_840_0, i_8_334_841_0, i_8_334_842_0, i_8_334_845_0,
    i_8_334_958_0, i_8_334_977_0, i_8_334_996_0, i_8_334_997_0,
    i_8_334_1052_0, i_8_334_1086_0, i_8_334_1113_0, i_8_334_1114_0,
    i_8_334_1133_0, i_8_334_1139_0, i_8_334_1156_0, i_8_334_1326_0,
    i_8_334_1327_0, i_8_334_1410_0, i_8_334_1527_0, i_8_334_1528_0,
    i_8_334_1535_0, i_8_334_1596_0, i_8_334_1598_0, i_8_334_1599_0,
    i_8_334_1600_0, i_8_334_1645_0, i_8_334_1654_0, i_8_334_1669_0,
    i_8_334_1762_0, i_8_334_1768_0, i_8_334_1771_0, i_8_334_1788_0,
    i_8_334_1802_0, i_8_334_1806_0, i_8_334_1807_0, i_8_334_1808_0,
    i_8_334_1867_0, i_8_334_1868_0, i_8_334_1870_0, i_8_334_1902_0,
    i_8_334_1903_0, i_8_334_1904_0, i_8_334_1918_0, i_8_334_1919_0,
    i_8_334_1921_0, i_8_334_1922_0, i_8_334_1949_0, i_8_334_1950_0,
    i_8_334_1952_0, i_8_334_1965_0, i_8_334_1969_0, i_8_334_1980_0,
    i_8_334_1983_0, i_8_334_2064_0, i_8_334_2118_0, i_8_334_2120_0,
    i_8_334_2121_0, i_8_334_2214_0, i_8_334_2216_0, i_8_334_2218_0,
    i_8_334_2219_0, i_8_334_2245_0, i_8_334_2267_0,
    o_8_334_0_0  );
  input  i_8_334_53_0, i_8_334_86_0, i_8_334_87_0, i_8_334_97_0,
    i_8_334_139_0, i_8_334_230_0, i_8_334_255_0, i_8_334_258_0,
    i_8_334_260_0, i_8_334_327_0, i_8_334_328_0, i_8_334_329_0,
    i_8_334_362_0, i_8_334_363_0, i_8_334_457_0, i_8_334_462_0,
    i_8_334_463_0, i_8_334_464_0, i_8_334_466_0, i_8_334_474_0,
    i_8_334_476_0, i_8_334_500_0, i_8_334_523_0, i_8_334_526_0,
    i_8_334_528_0, i_8_334_530_0, i_8_334_555_0, i_8_334_617_0,
    i_8_334_660_0, i_8_334_661_0, i_8_334_663_0, i_8_334_672_0,
    i_8_334_674_0, i_8_334_682_0, i_8_334_732_0, i_8_334_762_0,
    i_8_334_763_0, i_8_334_840_0, i_8_334_841_0, i_8_334_842_0,
    i_8_334_845_0, i_8_334_958_0, i_8_334_977_0, i_8_334_996_0,
    i_8_334_997_0, i_8_334_1052_0, i_8_334_1086_0, i_8_334_1113_0,
    i_8_334_1114_0, i_8_334_1133_0, i_8_334_1139_0, i_8_334_1156_0,
    i_8_334_1326_0, i_8_334_1327_0, i_8_334_1410_0, i_8_334_1527_0,
    i_8_334_1528_0, i_8_334_1535_0, i_8_334_1596_0, i_8_334_1598_0,
    i_8_334_1599_0, i_8_334_1600_0, i_8_334_1645_0, i_8_334_1654_0,
    i_8_334_1669_0, i_8_334_1762_0, i_8_334_1768_0, i_8_334_1771_0,
    i_8_334_1788_0, i_8_334_1802_0, i_8_334_1806_0, i_8_334_1807_0,
    i_8_334_1808_0, i_8_334_1867_0, i_8_334_1868_0, i_8_334_1870_0,
    i_8_334_1902_0, i_8_334_1903_0, i_8_334_1904_0, i_8_334_1918_0,
    i_8_334_1919_0, i_8_334_1921_0, i_8_334_1922_0, i_8_334_1949_0,
    i_8_334_1950_0, i_8_334_1952_0, i_8_334_1965_0, i_8_334_1969_0,
    i_8_334_1980_0, i_8_334_1983_0, i_8_334_2064_0, i_8_334_2118_0,
    i_8_334_2120_0, i_8_334_2121_0, i_8_334_2214_0, i_8_334_2216_0,
    i_8_334_2218_0, i_8_334_2219_0, i_8_334_2245_0, i_8_334_2267_0;
  output o_8_334_0_0;
  assign o_8_334_0_0 = ~((~i_8_334_474_0 & ((~i_8_334_86_0 & ((~i_8_334_464_0 & ~i_8_334_1599_0 & i_8_334_1645_0 & ~i_8_334_1868_0 & ~i_8_334_1919_0 & ~i_8_334_1965_0) | (~i_8_334_230_0 & ~i_8_334_476_0 & ~i_8_334_500_0 & ~i_8_334_1326_0 & ~i_8_334_1535_0 & ~i_8_334_1600_0 & ~i_8_334_1950_0 & ~i_8_334_2064_0 & ~i_8_334_2121_0))) | (~i_8_334_462_0 & ~i_8_334_464_0 & ((~i_8_334_476_0 & i_8_334_1904_0) | (~i_8_334_1599_0 & ~i_8_334_1600_0 & ~i_8_334_1654_0 & ~i_8_334_1870_0 & ~i_8_334_1919_0 & ~i_8_334_2121_0 & ~i_8_334_2219_0))) | (~i_8_334_260_0 & ~i_8_334_660_0 & ~i_8_334_672_0 & ~i_8_334_841_0 & i_8_334_996_0 & ~i_8_334_1086_0 & ~i_8_334_1139_0 & ~i_8_334_1326_0 & ~i_8_334_2064_0) | (~i_8_334_230_0 & ~i_8_334_463_0 & ~i_8_334_1599_0 & ~i_8_334_1868_0 & ~i_8_334_1969_0 & ~i_8_334_2120_0 & ~i_8_334_2214_0 & ~i_8_334_2218_0))) | (~i_8_334_466_0 & ((~i_8_334_86_0 & ((~i_8_334_462_0 & ~i_8_334_463_0 & ~i_8_334_660_0 & ~i_8_334_762_0 & ~i_8_334_763_0 & ~i_8_334_977_0 & ~i_8_334_1535_0 & ~i_8_334_1868_0 & ~i_8_334_1950_0 & ~i_8_334_2118_0) | (~i_8_334_476_0 & ~i_8_334_528_0 & ~i_8_334_1965_0 & ~i_8_334_2216_0))) | (i_8_334_86_0 & ~i_8_334_363_0 & ~i_8_334_958_0 & ~i_8_334_996_0 & ~i_8_334_1139_0 & ~i_8_334_1918_0 & i_8_334_1922_0 & ~i_8_334_1965_0 & ~i_8_334_2245_0))) | (~i_8_334_1600_0 & ((~i_8_334_363_0 & ~i_8_334_1949_0 & ((~i_8_334_462_0 & i_8_334_977_0 & ~i_8_334_1952_0) | (i_8_334_526_0 & ~i_8_334_1052_0 & ~i_8_334_1596_0 & ~i_8_334_1645_0 & ~i_8_334_1654_0 & ~i_8_334_1950_0 & ~i_8_334_2216_0 & ~i_8_334_2245_0))) | (~i_8_334_462_0 & ~i_8_334_463_0 & ~i_8_334_526_0 & ~i_8_334_762_0 & i_8_334_841_0 & ~i_8_334_1086_0 & ~i_8_334_1771_0 & ~i_8_334_1950_0))) | (~i_8_334_528_0 & ((~i_8_334_526_0 & ~i_8_334_617_0 & i_8_334_1918_0 & ~i_8_334_1921_0 & i_8_334_1965_0) | (~i_8_334_464_0 & i_8_334_523_0 & ~i_8_334_674_0 & ~i_8_334_840_0 & ~i_8_334_1598_0 & ~i_8_334_1771_0 & ~i_8_334_1788_0 & ~i_8_334_1870_0 & ~i_8_334_1980_0 & ~i_8_334_2064_0))) | (~i_8_334_1870_0 & ((~i_8_334_530_0 & ~i_8_334_674_0 & ((~i_8_334_464_0 & ~i_8_334_762_0 & ~i_8_334_1596_0 & ~i_8_334_1598_0 & ~i_8_334_1599_0 & ~i_8_334_1867_0 & ~i_8_334_2118_0 & ~i_8_334_2120_0) | (~i_8_334_462_0 & ~i_8_334_555_0 & ~i_8_334_763_0 & ~i_8_334_1645_0 & i_8_334_1918_0 & ~i_8_334_2214_0 & ~i_8_334_2216_0))) | (~i_8_334_500_0 & ~i_8_334_526_0 & ~i_8_334_762_0 & ~i_8_334_763_0 & i_8_334_841_0 & ~i_8_334_1086_0 & ~i_8_334_2064_0))) | (~i_8_334_476_0 & ((~i_8_334_462_0 & ((~i_8_334_464_0 & ~i_8_334_555_0 & ~i_8_334_617_0 & ~i_8_334_1598_0 & ~i_8_334_1806_0 & ~i_8_334_1808_0) | (~i_8_334_526_0 & ~i_8_334_763_0 & ~i_8_334_1599_0 & ~i_8_334_1950_0 & ~i_8_334_2118_0 & ~i_8_334_1867_0 & ~i_8_334_1868_0))) | (~i_8_334_2121_0 & ((i_8_334_526_0 & ~i_8_334_763_0 & ~i_8_334_996_0 & ~i_8_334_1596_0 & ~i_8_334_1868_0 & ~i_8_334_1904_0 & ~i_8_334_1919_0 & ~i_8_334_2118_0) | (~i_8_334_555_0 & ~i_8_334_1598_0 & ~i_8_334_1918_0 & ~i_8_334_2120_0 & ~i_8_334_2218_0))))) | (i_8_334_997_0 & (i_8_334_258_0 | (~i_8_334_463_0 & ~i_8_334_1599_0 & ~i_8_334_1762_0 & ~i_8_334_1952_0 & ~i_8_334_2064_0))) | (~i_8_334_1950_0 & ((~i_8_334_463_0 & ((~i_8_334_674_0 & ~i_8_334_1535_0 & ~i_8_334_1599_0 & ~i_8_334_1762_0 & ~i_8_334_1788_0 & ~i_8_334_1918_0) | (i_8_334_1902_0 & ~i_8_334_2216_0))) | (~i_8_334_523_0 & ~i_8_334_526_0 & ~i_8_334_530_0 & ~i_8_334_763_0 & ~i_8_334_1598_0 & ~i_8_334_1654_0 & ~i_8_334_1949_0 & ~i_8_334_1952_0))) | (~i_8_334_674_0 & ~i_8_334_1918_0 & ((i_8_334_530_0 & ~i_8_334_958_0 & ~i_8_334_1596_0 & ~i_8_334_1807_0 & ~i_8_334_1868_0 & ~i_8_334_2214_0) | (~i_8_334_672_0 & ~i_8_334_763_0 & ~i_8_334_1598_0 & ~i_8_334_2121_0 & ~i_8_334_2219_0 & ~i_8_334_1904_0 & ~i_8_334_2120_0))) | (~i_8_334_464_0 & ~i_8_334_763_0 & ~i_8_334_1133_0 & ~i_8_334_1410_0 & i_8_334_1788_0 & ~i_8_334_1921_0 & ~i_8_334_2120_0) | (~i_8_334_87_0 & i_8_334_660_0 & ~i_8_334_1762_0 & ~i_8_334_2118_0) | (~i_8_334_841_0 & ~i_8_334_845_0 & ~i_8_334_1139_0 & ~i_8_334_1806_0 & ~i_8_334_1868_0 & ~i_8_334_1919_0 & ~i_8_334_1952_0 & ~i_8_334_2121_0 & ~i_8_334_2218_0));
endmodule



// Benchmark "kernel_8_335" written by ABC on Sun Jul 19 10:08:53 2020

module kernel_8_335 ( 
    i_8_335_34_0, i_8_335_53_0, i_8_335_80_0, i_8_335_115_0, i_8_335_143_0,
    i_8_335_189_0, i_8_335_190_0, i_8_335_191_0, i_8_335_193_0,
    i_8_335_252_0, i_8_335_292_0, i_8_335_301_0, i_8_335_302_0,
    i_8_335_305_0, i_8_335_345_0, i_8_335_346_0, i_8_335_362_0,
    i_8_335_378_0, i_8_335_379_0, i_8_335_380_0, i_8_335_381_0,
    i_8_335_383_0, i_8_335_463_0, i_8_335_468_0, i_8_335_469_0,
    i_8_335_492_0, i_8_335_522_0, i_8_335_550_0, i_8_335_591_0,
    i_8_335_606_0, i_8_335_607_0, i_8_335_608_0, i_8_335_610_0,
    i_8_335_611_0, i_8_335_627_0, i_8_335_663_0, i_8_335_664_0,
    i_8_335_689_0, i_8_335_712_0, i_8_335_726_0, i_8_335_735_0,
    i_8_335_764_0, i_8_335_834_0, i_8_335_989_0, i_8_335_997_0,
    i_8_335_998_0, i_8_335_1086_0, i_8_335_1111_0, i_8_335_1112_0,
    i_8_335_1125_0, i_8_335_1235_0, i_8_335_1261_0, i_8_335_1273_0,
    i_8_335_1274_0, i_8_335_1286_0, i_8_335_1306_0, i_8_335_1410_0,
    i_8_335_1435_0, i_8_335_1436_0, i_8_335_1470_0, i_8_335_1471_0,
    i_8_335_1528_0, i_8_335_1529_0, i_8_335_1533_0, i_8_335_1537_0,
    i_8_335_1605_0, i_8_335_1617_0, i_8_335_1624_0, i_8_335_1660_0,
    i_8_335_1680_0, i_8_335_1681_0, i_8_335_1751_0, i_8_335_1758_0,
    i_8_335_1803_0, i_8_335_1804_0, i_8_335_1824_0, i_8_335_1863_0,
    i_8_335_1865_0, i_8_335_1887_0, i_8_335_1984_0, i_8_335_1991_0,
    i_8_335_1992_0, i_8_335_1996_0, i_8_335_2034_0, i_8_335_2073_0,
    i_8_335_2109_0, i_8_335_2139_0, i_8_335_2140_0, i_8_335_2141_0,
    i_8_335_2149_0, i_8_335_2151_0, i_8_335_2153_0, i_8_335_2154_0,
    i_8_335_2155_0, i_8_335_2156_0, i_8_335_2157_0, i_8_335_2214_0,
    i_8_335_2215_0, i_8_335_2216_0, i_8_335_2275_0,
    o_8_335_0_0  );
  input  i_8_335_34_0, i_8_335_53_0, i_8_335_80_0, i_8_335_115_0,
    i_8_335_143_0, i_8_335_189_0, i_8_335_190_0, i_8_335_191_0,
    i_8_335_193_0, i_8_335_252_0, i_8_335_292_0, i_8_335_301_0,
    i_8_335_302_0, i_8_335_305_0, i_8_335_345_0, i_8_335_346_0,
    i_8_335_362_0, i_8_335_378_0, i_8_335_379_0, i_8_335_380_0,
    i_8_335_381_0, i_8_335_383_0, i_8_335_463_0, i_8_335_468_0,
    i_8_335_469_0, i_8_335_492_0, i_8_335_522_0, i_8_335_550_0,
    i_8_335_591_0, i_8_335_606_0, i_8_335_607_0, i_8_335_608_0,
    i_8_335_610_0, i_8_335_611_0, i_8_335_627_0, i_8_335_663_0,
    i_8_335_664_0, i_8_335_689_0, i_8_335_712_0, i_8_335_726_0,
    i_8_335_735_0, i_8_335_764_0, i_8_335_834_0, i_8_335_989_0,
    i_8_335_997_0, i_8_335_998_0, i_8_335_1086_0, i_8_335_1111_0,
    i_8_335_1112_0, i_8_335_1125_0, i_8_335_1235_0, i_8_335_1261_0,
    i_8_335_1273_0, i_8_335_1274_0, i_8_335_1286_0, i_8_335_1306_0,
    i_8_335_1410_0, i_8_335_1435_0, i_8_335_1436_0, i_8_335_1470_0,
    i_8_335_1471_0, i_8_335_1528_0, i_8_335_1529_0, i_8_335_1533_0,
    i_8_335_1537_0, i_8_335_1605_0, i_8_335_1617_0, i_8_335_1624_0,
    i_8_335_1660_0, i_8_335_1680_0, i_8_335_1681_0, i_8_335_1751_0,
    i_8_335_1758_0, i_8_335_1803_0, i_8_335_1804_0, i_8_335_1824_0,
    i_8_335_1863_0, i_8_335_1865_0, i_8_335_1887_0, i_8_335_1984_0,
    i_8_335_1991_0, i_8_335_1992_0, i_8_335_1996_0, i_8_335_2034_0,
    i_8_335_2073_0, i_8_335_2109_0, i_8_335_2139_0, i_8_335_2140_0,
    i_8_335_2141_0, i_8_335_2149_0, i_8_335_2151_0, i_8_335_2153_0,
    i_8_335_2154_0, i_8_335_2155_0, i_8_335_2156_0, i_8_335_2157_0,
    i_8_335_2214_0, i_8_335_2215_0, i_8_335_2216_0, i_8_335_2275_0;
  output o_8_335_0_0;
  assign o_8_335_0_0 = ~((~i_8_335_189_0 & ((~i_8_335_190_0 & ((~i_8_335_34_0 & ((~i_8_335_252_0 & ~i_8_335_302_0 & ~i_8_335_362_0 & ~i_8_335_383_0 & i_8_335_607_0 & ~i_8_335_712_0 & ~i_8_335_726_0 & ~i_8_335_989_0 & ~i_8_335_1235_0 & ~i_8_335_1617_0 & ~i_8_335_1680_0 & ~i_8_335_2034_0) | (i_8_335_383_0 & ~i_8_335_998_0 & ~i_8_335_2140_0 & ~i_8_335_2153_0 & i_8_335_2156_0))) | (i_8_335_345_0 & ~i_8_335_591_0 & ~i_8_335_610_0 & ~i_8_335_664_0 & ~i_8_335_735_0 & i_8_335_1470_0 & ~i_8_335_1992_0 & ~i_8_335_2153_0 & ~i_8_335_2216_0))) | (~i_8_335_989_0 & ((~i_8_335_53_0 & ~i_8_335_1235_0 & ((~i_8_335_362_0 & ~i_8_335_469_0 & i_8_335_607_0 & i_8_335_608_0) | (~i_8_335_143_0 & ~i_8_335_302_0 & ~i_8_335_591_0 & ~i_8_335_611_0 & ~i_8_335_735_0 & ~i_8_335_834_0 & ~i_8_335_1086_0 & ~i_8_335_1528_0 & i_8_335_1537_0 & ~i_8_335_2139_0 & ~i_8_335_2151_0 & ~i_8_335_2153_0 & ~i_8_335_2156_0))) | (~i_8_335_664_0 & ((i_8_335_115_0 & ~i_8_335_381_0 & ~i_8_335_383_0 & ~i_8_335_712_0 & ~i_8_335_1617_0 & i_8_335_1996_0 & i_8_335_2149_0 & ~i_8_335_2151_0) | (~i_8_335_305_0 & ~i_8_335_378_0 & ~i_8_335_2034_0 & i_8_335_2155_0 & i_8_335_2156_0))) | (~i_8_335_191_0 & i_8_335_301_0 & i_8_335_468_0 & ~i_8_335_1261_0 & i_8_335_1751_0 & ~i_8_335_2139_0))) | (~i_8_335_2141_0 & ((~i_8_335_305_0 & ((~i_8_335_143_0 & i_8_335_1274_0 & i_8_335_1436_0 & ~i_8_335_1660_0 & ~i_8_335_1863_0 & ~i_8_335_1991_0 & ~i_8_335_2151_0) | (~i_8_335_345_0 & ~i_8_335_381_0 & ~i_8_335_522_0 & ~i_8_335_663_0 & ~i_8_335_998_0 & ~i_8_335_1410_0 & ~i_8_335_1617_0 & i_8_335_1681_0 & ~i_8_335_1751_0 & ~i_8_335_1804_0 & ~i_8_335_1824_0 & ~i_8_335_1887_0 & ~i_8_335_2140_0 & ~i_8_335_2157_0))) | (~i_8_335_663_0 & ~i_8_335_1125_0 & ~i_8_335_1991_0 & ~i_8_335_2151_0 & ((i_8_335_115_0 & ~i_8_335_610_0 & ~i_8_335_611_0 & ~i_8_335_726_0 & ~i_8_335_764_0 & ~i_8_335_1261_0 & ~i_8_335_1410_0 & ~i_8_335_1803_0 & ~i_8_335_1887_0) | (~i_8_335_379_0 & ~i_8_335_380_0 & ~i_8_335_591_0 & ~i_8_335_712_0 & ~i_8_335_998_0 & ~i_8_335_1086_0 & ~i_8_335_2139_0 & ~i_8_335_2140_0 & i_8_335_2215_0))) | (~i_8_335_345_0 & ~i_8_335_627_0 & ~i_8_335_735_0 & ~i_8_335_997_0 & ~i_8_335_1261_0 & ~i_8_335_1681_0 & i_8_335_1758_0 & ~i_8_335_1863_0 & ~i_8_335_1865_0 & ~i_8_335_2157_0))) | (~i_8_335_379_0 & ((~i_8_335_468_0 & ~i_8_335_591_0 & ~i_8_335_735_0 & ~i_8_335_764_0 & ~i_8_335_1125_0 & ~i_8_335_1261_0 & ~i_8_335_1470_0 & ~i_8_335_1617_0 & i_8_335_2154_0) | (~i_8_335_346_0 & ~i_8_335_611_0 & ~i_8_335_998_0 & ~i_8_335_1112_0 & ~i_8_335_1529_0 & ~i_8_335_1991_0 & ~i_8_335_2034_0 & ~i_8_335_2157_0 & i_8_335_2216_0))) | (~i_8_335_735_0 & ~i_8_335_1865_0 & ((i_8_335_383_0 & ~i_8_335_764_0 & ~i_8_335_998_0 & ~i_8_335_1235_0 & i_8_335_1435_0 & i_8_335_1436_0 & ~i_8_335_1470_0 & ~i_8_335_1537_0) | (~i_8_335_193_0 & ~i_8_335_380_0 & ~i_8_335_1410_0 & i_8_335_1470_0 & ~i_8_335_1617_0 & ~i_8_335_2151_0 & i_8_335_2157_0) | (~i_8_335_191_0 & ~i_8_335_468_0 & ~i_8_335_469_0 & ~i_8_335_664_0 & ~i_8_335_1111_0 & ~i_8_335_2034_0 & ~i_8_335_2139_0 & ~i_8_335_2156_0 & i_8_335_2215_0 & ~i_8_335_2275_0))))) | (~i_8_335_1537_0 & ((~i_8_335_2214_0 & ((~i_8_335_53_0 & ((~i_8_335_191_0 & ~i_8_335_378_0 & ~i_8_335_380_0 & ~i_8_335_591_0 & ~i_8_335_627_0 & ~i_8_335_663_0 & ~i_8_335_764_0 & ~i_8_335_834_0 & ~i_8_335_989_0 & ~i_8_335_997_0 & ~i_8_335_1436_0 & ~i_8_335_1680_0 & ~i_8_335_1863_0 & i_8_335_2149_0) | (i_8_335_115_0 & ~i_8_335_305_0 & ~i_8_335_346_0 & ~i_8_335_550_0 & ~i_8_335_611_0 & ~i_8_335_735_0 & ~i_8_335_998_0 & ~i_8_335_1125_0 & ~i_8_335_1617_0 & ~i_8_335_1991_0 & ~i_8_335_1992_0 & ~i_8_335_2151_0))) | (~i_8_335_190_0 & ~i_8_335_292_0 & ~i_8_335_301_0 & ~i_8_335_550_0 & ~i_8_335_664_0 & ~i_8_335_1086_0 & i_8_335_1471_0 & ~i_8_335_1681_0 & ~i_8_335_1865_0 & ~i_8_335_1991_0 & ~i_8_335_2151_0))) | (~i_8_335_378_0 & ((~i_8_335_381_0 & ~i_8_335_550_0 & ~i_8_335_1086_0 & ~i_8_335_1261_0 & ~i_8_335_1617_0 & i_8_335_1824_0 & i_8_335_2073_0 & ~i_8_335_2141_0) | (~i_8_335_346_0 & i_8_335_606_0 & ~i_8_335_608_0 & ~i_8_335_1125_0 & ~i_8_335_2139_0 & ~i_8_335_2151_0 & ~i_8_335_1751_0 & ~i_8_335_2034_0))) | (~i_8_335_663_0 & ((~i_8_335_190_0 & ~i_8_335_252_0 & ~i_8_335_345_0 & ~i_8_335_550_0 & i_8_335_591_0 & ~i_8_335_664_0 & ~i_8_335_712_0 & ~i_8_335_998_0 & ~i_8_335_2140_0) | (~i_8_335_834_0 & i_8_335_1470_0 & ~i_8_335_1624_0 & i_8_335_2109_0 & ~i_8_335_2141_0 & i_8_335_2154_0))) | (~i_8_335_190_0 & ((~i_8_335_380_0 & i_8_335_1274_0 & i_8_335_1991_0) | (i_8_335_302_0 & ~i_8_335_712_0 & ~i_8_335_1261_0 & ~i_8_335_1865_0 & ~i_8_335_2109_0 & ~i_8_335_2139_0 & ~i_8_335_2141_0 & ~i_8_335_2151_0 & ~i_8_335_2153_0 & ~i_8_335_2156_0))) | (~i_8_335_1617_0 & i_8_335_1824_0 & ~i_8_335_606_0 & ~i_8_335_1471_0 & i_8_335_2141_0 & i_8_335_2149_0 & ~i_8_335_2155_0 & ~i_8_335_2157_0))) | (~i_8_335_193_0 & ((~i_8_335_379_0 & ~i_8_335_468_0 & i_8_335_522_0 & ~i_8_335_1863_0 & ~i_8_335_1865_0 & i_8_335_1984_0 & ~i_8_335_2140_0) | (~i_8_335_252_0 & i_8_335_301_0 & ~i_8_335_378_0 & ~i_8_335_1086_0 & ~i_8_335_1112_0 & ~i_8_335_1286_0 & ~i_8_335_1436_0 & ~i_8_335_1681_0 & ~i_8_335_1804_0 & ~i_8_335_1991_0 & ~i_8_335_2034_0 & ~i_8_335_2157_0))) | (~i_8_335_191_0 & ((~i_8_335_1617_0 & ((~i_8_335_34_0 & ~i_8_335_664_0 & ((~i_8_335_379_0 & i_8_335_383_0 & ~i_8_335_550_0 & i_8_335_1111_0 & ~i_8_335_1306_0 & ~i_8_335_2141_0) | (~i_8_335_190_0 & ~i_8_335_591_0 & ~i_8_335_611_0 & ~i_8_335_627_0 & ~i_8_335_712_0 & ~i_8_335_998_0 & ~i_8_335_1086_0 & ~i_8_335_1111_0 & ~i_8_335_1528_0 & ~i_8_335_1865_0 & i_8_335_2149_0))) | (~i_8_335_252_0 & i_8_335_302_0 & ~i_8_335_380_0 & ~i_8_335_550_0 & ~i_8_335_998_0 & ~i_8_335_1529_0 & ~i_8_335_1681_0 & ~i_8_335_2140_0))) | (~i_8_335_522_0 & ~i_8_335_989_0 & ((i_8_335_689_0 & i_8_335_764_0 & ~i_8_335_1528_0 & ~i_8_335_1824_0 & ~i_8_335_1996_0) | (~i_8_335_469_0 & ~i_8_335_550_0 & ~i_8_335_607_0 & ~i_8_335_764_0 & ~i_8_335_998_0 & ~i_8_335_1261_0 & ~i_8_335_1436_0 & ~i_8_335_1681_0 & i_8_335_1751_0 & ~i_8_335_1758_0 & ~i_8_335_2141_0))) | (i_8_335_143_0 & ~i_8_335_764_0 & ~i_8_335_997_0 & ~i_8_335_1804_0 & ~i_8_335_2034_0 & ~i_8_335_2141_0 & ~i_8_335_2151_0 & ~i_8_335_2157_0) | (~i_8_335_252_0 & ~i_8_335_379_0 & ~i_8_335_712_0 & ~i_8_335_1086_0 & ~i_8_335_1235_0 & ~i_8_335_1529_0 & ~i_8_335_1680_0 & ~i_8_335_1865_0 & i_8_335_2155_0 & ~i_8_335_2275_0))) | (i_8_335_301_0 & ((~i_8_335_463_0 & i_8_335_607_0 & i_8_335_1112_0 & ~i_8_335_2139_0 & ~i_8_335_2151_0 & ~i_8_335_1274_0 & ~i_8_335_1470_0) | (i_8_335_664_0 & ~i_8_335_2140_0 & i_8_335_2155_0))) | (i_8_335_346_0 & ~i_8_335_378_0 & ((i_8_335_193_0 & ~i_8_335_522_0 & ~i_8_335_712_0 & ~i_8_335_735_0 & ~i_8_335_1086_0 & ~i_8_335_1261_0 & ~i_8_335_1529_0 & ~i_8_335_1617_0) | (~i_8_335_190_0 & ~i_8_335_380_0 & ~i_8_335_492_0 & ~i_8_335_627_0 & ~i_8_335_664_0 & ~i_8_335_764_0 & ~i_8_335_1758_0 & ~i_8_335_2141_0 & ~i_8_335_2153_0 & ~i_8_335_2214_0))) | (~i_8_335_80_0 & ((i_8_335_193_0 & ((~i_8_335_190_0 & ~i_8_335_997_0 & i_8_335_1996_0 & ~i_8_335_2034_0 & ~i_8_335_2139_0 & ~i_8_335_2151_0) | (~i_8_335_34_0 & i_8_335_383_0 & ~i_8_335_1086_0 & i_8_335_2156_0 & ~i_8_335_2215_0))) | (~i_8_335_190_0 & ((~i_8_335_611_0 & ~i_8_335_627_0 & ~i_8_335_712_0 & ~i_8_335_468_0 & ~i_8_335_522_0 & ~i_8_335_1086_0 & ~i_8_335_1235_0 & ~i_8_335_1529_0 & i_8_335_1624_0 & ~i_8_335_2140_0) | (~i_8_335_115_0 & ~i_8_335_379_0 & ~i_8_335_380_0 & i_8_335_463_0 & ~i_8_335_2139_0 & ~i_8_335_2151_0 & ~i_8_335_997_0 & ~i_8_335_1261_0))) | (~i_8_335_305_0 & ~i_8_335_345_0 & ~i_8_335_469_0 & ~i_8_335_611_0 & ~i_8_335_997_0 & i_8_335_1286_0 & ~i_8_335_2034_0 & ~i_8_335_2140_0 & ~i_8_335_2141_0 & ~i_8_335_2215_0))) | (~i_8_335_34_0 & ~i_8_335_305_0 & ((~i_8_335_380_0 & i_8_335_383_0 & ~i_8_335_468_0 & ~i_8_335_764_0 & ~i_8_335_997_0 & ~i_8_335_1086_0 & ~i_8_335_1617_0 & ~i_8_335_1660_0 & i_8_335_1751_0 & ~i_8_335_1863_0) | (~i_8_335_379_0 & ~i_8_335_834_0 & i_8_335_1410_0 & ~i_8_335_1436_0 & ~i_8_335_1470_0 & ~i_8_335_1471_0 & ~i_8_335_1528_0 & ~i_8_335_1681_0 & ~i_8_335_2034_0))) | (i_8_335_2215_0 & ((~i_8_335_379_0 & ((i_8_335_381_0 & ~i_8_335_726_0 & ~i_8_335_997_0 & ~i_8_335_1086_0 & ~i_8_335_1111_0 & ~i_8_335_1471_0 & ~i_8_335_2073_0) | (~i_8_335_468_0 & ~i_8_335_1306_0 & ~i_8_335_1751_0 & ~i_8_335_2139_0 & i_8_335_2214_0))) | (~i_8_335_190_0 & i_8_335_522_0 & ~i_8_335_550_0 & ~i_8_335_607_0 & ~i_8_335_1111_0 & ~i_8_335_1261_0 & ~i_8_335_1680_0 & ~i_8_335_2141_0 & ~i_8_335_2157_0 & i_8_335_2214_0))) | (~i_8_335_190_0 & ((~i_8_335_380_0 & ~i_8_335_611_0 & ~i_8_335_997_0 & ~i_8_335_1086_0 & ~i_8_335_1125_0 & ~i_8_335_1435_0 & i_8_335_2155_0 & ~i_8_335_2157_0) | (~i_8_335_522_0 & ~i_8_335_550_0 & ~i_8_335_627_0 & ~i_8_335_1235_0 & ~i_8_335_1436_0 & ~i_8_335_1865_0 & i_8_335_1984_0 & ~i_8_335_1992_0 & ~i_8_335_2140_0 & ~i_8_335_2141_0 & ~i_8_335_2153_0 & ~i_8_335_2215_0))) | (i_8_335_383_0 & ((~i_8_335_143_0 & ~i_8_335_627_0 & ~i_8_335_1086_0 & ~i_8_335_1529_0 & ~i_8_335_1533_0 & i_8_335_1996_0 & ~i_8_335_2140_0 & ~i_8_335_2153_0) | (~i_8_335_469_0 & ~i_8_335_998_0 & i_8_335_1286_0 & ~i_8_335_1681_0 & ~i_8_335_1751_0 & ~i_8_335_1803_0 & ~i_8_335_2156_0))) | (i_8_335_606_0 & ~i_8_335_1863_0 & ((~i_8_335_383_0 & ~i_8_335_1235_0 & ~i_8_335_1887_0 & ~i_8_335_2151_0 & ~i_8_335_2153_0 & i_8_335_2154_0) | (~i_8_335_468_0 & ~i_8_335_1086_0 & ~i_8_335_1529_0 & ~i_8_335_1992_0 & i_8_335_2155_0))) | (i_8_335_2156_0 & ((~i_8_335_469_0 & ((i_8_335_362_0 & i_8_335_1865_0 & ~i_8_335_2140_0 & i_8_335_2153_0) | (i_8_335_608_0 & ~i_8_335_712_0 & ~i_8_335_997_0 & ~i_8_335_1086_0 & ~i_8_335_2275_0))) | (~i_8_335_463_0 & ~i_8_335_550_0 & ~i_8_335_611_0 & ~i_8_335_664_0 & ~i_8_335_1751_0 & ~i_8_335_1804_0 & ~i_8_335_712_0 & ~i_8_335_1235_0))) | (~i_8_335_1261_0 & ((i_8_335_302_0 & ~i_8_335_1112_0 & ~i_8_335_1436_0 & ~i_8_335_1529_0 & ~i_8_335_2140_0 & ~i_8_335_2153_0 & ~i_8_335_1758_0 & ~i_8_335_1865_0) | (~i_8_335_380_0 & ~i_8_335_469_0 & i_8_335_607_0 & ~i_8_335_998_0 & ~i_8_335_1125_0 & ~i_8_335_1804_0 & i_8_335_1984_0 & ~i_8_335_2214_0))) | (~i_8_335_1533_0 & ~i_8_335_1803_0 & i_8_335_1992_0 & i_8_335_2034_0 & i_8_335_2073_0 & i_8_335_2109_0));
endmodule



// Benchmark "kernel_8_336" written by ABC on Sun Jul 19 10:08:54 2020

module kernel_8_336 ( 
    i_8_336_11_0, i_8_336_19_0, i_8_336_27_0, i_8_336_34_0, i_8_336_73_0,
    i_8_336_74_0, i_8_336_83_0, i_8_336_101_0, i_8_336_141_0,
    i_8_336_298_0, i_8_336_325_0, i_8_336_326_0, i_8_336_364_0,
    i_8_336_367_0, i_8_336_450_0, i_8_336_486_0, i_8_336_562_0,
    i_8_336_577_0, i_8_336_579_0, i_8_336_589_0, i_8_336_611_0,
    i_8_336_639_0, i_8_336_640_0, i_8_336_657_0, i_8_336_663_0,
    i_8_336_676_0, i_8_336_684_0, i_8_336_694_0, i_8_336_707_0,
    i_8_336_708_0, i_8_336_712_0, i_8_336_713_0, i_8_336_721_0,
    i_8_336_729_0, i_8_336_733_0, i_8_336_791_0, i_8_336_822_0,
    i_8_336_837_0, i_8_336_844_0, i_8_336_855_0, i_8_336_967_0,
    i_8_336_996_0, i_8_336_1026_0, i_8_336_1129_0, i_8_336_1134_0,
    i_8_336_1179_0, i_8_336_1183_0, i_8_336_1206_0, i_8_336_1243_0,
    i_8_336_1252_0, i_8_336_1261_0, i_8_336_1285_0, i_8_336_1286_0,
    i_8_336_1296_0, i_8_336_1395_0, i_8_336_1398_0, i_8_336_1473_0,
    i_8_336_1480_0, i_8_336_1507_0, i_8_336_1513_0, i_8_336_1516_0,
    i_8_336_1530_0, i_8_336_1534_0, i_8_336_1555_0, i_8_336_1563_0,
    i_8_336_1595_0, i_8_336_1605_0, i_8_336_1625_0, i_8_336_1668_0,
    i_8_336_1675_0, i_8_336_1680_0, i_8_336_1707_0, i_8_336_1710_0,
    i_8_336_1711_0, i_8_336_1745_0, i_8_336_1754_0, i_8_336_1756_0,
    i_8_336_1757_0, i_8_336_1789_0, i_8_336_1802_0, i_8_336_1810_0,
    i_8_336_1819_0, i_8_336_1826_0, i_8_336_1854_0, i_8_336_1883_0,
    i_8_336_1900_0, i_8_336_1989_0, i_8_336_1990_0, i_8_336_2011_0,
    i_8_336_2017_0, i_8_336_2025_0, i_8_336_2088_0, i_8_336_2137_0,
    i_8_336_2147_0, i_8_336_2152_0, i_8_336_2206_0, i_8_336_2245_0,
    i_8_336_2246_0, i_8_336_2265_0, i_8_336_2292_0,
    o_8_336_0_0  );
  input  i_8_336_11_0, i_8_336_19_0, i_8_336_27_0, i_8_336_34_0,
    i_8_336_73_0, i_8_336_74_0, i_8_336_83_0, i_8_336_101_0, i_8_336_141_0,
    i_8_336_298_0, i_8_336_325_0, i_8_336_326_0, i_8_336_364_0,
    i_8_336_367_0, i_8_336_450_0, i_8_336_486_0, i_8_336_562_0,
    i_8_336_577_0, i_8_336_579_0, i_8_336_589_0, i_8_336_611_0,
    i_8_336_639_0, i_8_336_640_0, i_8_336_657_0, i_8_336_663_0,
    i_8_336_676_0, i_8_336_684_0, i_8_336_694_0, i_8_336_707_0,
    i_8_336_708_0, i_8_336_712_0, i_8_336_713_0, i_8_336_721_0,
    i_8_336_729_0, i_8_336_733_0, i_8_336_791_0, i_8_336_822_0,
    i_8_336_837_0, i_8_336_844_0, i_8_336_855_0, i_8_336_967_0,
    i_8_336_996_0, i_8_336_1026_0, i_8_336_1129_0, i_8_336_1134_0,
    i_8_336_1179_0, i_8_336_1183_0, i_8_336_1206_0, i_8_336_1243_0,
    i_8_336_1252_0, i_8_336_1261_0, i_8_336_1285_0, i_8_336_1286_0,
    i_8_336_1296_0, i_8_336_1395_0, i_8_336_1398_0, i_8_336_1473_0,
    i_8_336_1480_0, i_8_336_1507_0, i_8_336_1513_0, i_8_336_1516_0,
    i_8_336_1530_0, i_8_336_1534_0, i_8_336_1555_0, i_8_336_1563_0,
    i_8_336_1595_0, i_8_336_1605_0, i_8_336_1625_0, i_8_336_1668_0,
    i_8_336_1675_0, i_8_336_1680_0, i_8_336_1707_0, i_8_336_1710_0,
    i_8_336_1711_0, i_8_336_1745_0, i_8_336_1754_0, i_8_336_1756_0,
    i_8_336_1757_0, i_8_336_1789_0, i_8_336_1802_0, i_8_336_1810_0,
    i_8_336_1819_0, i_8_336_1826_0, i_8_336_1854_0, i_8_336_1883_0,
    i_8_336_1900_0, i_8_336_1989_0, i_8_336_1990_0, i_8_336_2011_0,
    i_8_336_2017_0, i_8_336_2025_0, i_8_336_2088_0, i_8_336_2137_0,
    i_8_336_2147_0, i_8_336_2152_0, i_8_336_2206_0, i_8_336_2245_0,
    i_8_336_2246_0, i_8_336_2265_0, i_8_336_2292_0;
  output o_8_336_0_0;
  assign o_8_336_0_0 = 0;
endmodule



// Benchmark "kernel_8_337" written by ABC on Sun Jul 19 10:08:55 2020

module kernel_8_337 ( 
    i_8_337_5_0, i_8_337_20_0, i_8_337_49_0, i_8_337_64_0, i_8_337_83_0,
    i_8_337_89_0, i_8_337_101_0, i_8_337_257_0, i_8_337_263_0,
    i_8_337_275_0, i_8_337_290_0, i_8_337_301_0, i_8_337_303_0,
    i_8_337_366_0, i_8_337_367_0, i_8_337_368_0, i_8_337_380_0,
    i_8_337_382_0, i_8_337_401_0, i_8_337_434_0, i_8_337_440_0,
    i_8_337_452_0, i_8_337_455_0, i_8_337_476_0, i_8_337_486_0,
    i_8_337_491_0, i_8_337_506_0, i_8_337_518_0, i_8_337_528_0,
    i_8_337_547_0, i_8_337_586_0, i_8_337_590_0, i_8_337_626_0,
    i_8_337_632_0, i_8_337_634_0, i_8_337_658_0, i_8_337_670_0,
    i_8_337_671_0, i_8_337_694_0, i_8_337_703_0, i_8_337_706_0,
    i_8_337_716_0, i_8_337_803_0, i_8_337_824_0, i_8_337_830_0,
    i_8_337_839_0, i_8_337_844_0, i_8_337_845_0, i_8_337_877_0,
    i_8_337_1012_0, i_8_337_1028_0, i_8_337_1130_0, i_8_337_1225_0,
    i_8_337_1256_0, i_8_337_1286_0, i_8_337_1350_0, i_8_337_1355_0,
    i_8_337_1388_0, i_8_337_1420_0, i_8_337_1442_0, i_8_337_1445_0,
    i_8_337_1456_0, i_8_337_1471_0, i_8_337_1531_0, i_8_337_1532_0,
    i_8_337_1536_0, i_8_337_1537_0, i_8_337_1544_0, i_8_337_1576_0,
    i_8_337_1585_0, i_8_337_1615_0, i_8_337_1621_0, i_8_337_1622_0,
    i_8_337_1747_0, i_8_337_1751_0, i_8_337_1753_0, i_8_337_1768_0,
    i_8_337_1782_0, i_8_337_1802_0, i_8_337_1819_0, i_8_337_1838_0,
    i_8_337_1846_0, i_8_337_1847_0, i_8_337_1850_0, i_8_337_1892_0,
    i_8_337_1895_0, i_8_337_1963_0, i_8_337_1964_0, i_8_337_1990_0,
    i_8_337_1993_0, i_8_337_2000_0, i_8_337_2012_0, i_8_337_2047_0,
    i_8_337_2063_0, i_8_337_2111_0, i_8_337_2117_0, i_8_337_2141_0,
    i_8_337_2170_0, i_8_337_2227_0, i_8_337_2237_0,
    o_8_337_0_0  );
  input  i_8_337_5_0, i_8_337_20_0, i_8_337_49_0, i_8_337_64_0,
    i_8_337_83_0, i_8_337_89_0, i_8_337_101_0, i_8_337_257_0,
    i_8_337_263_0, i_8_337_275_0, i_8_337_290_0, i_8_337_301_0,
    i_8_337_303_0, i_8_337_366_0, i_8_337_367_0, i_8_337_368_0,
    i_8_337_380_0, i_8_337_382_0, i_8_337_401_0, i_8_337_434_0,
    i_8_337_440_0, i_8_337_452_0, i_8_337_455_0, i_8_337_476_0,
    i_8_337_486_0, i_8_337_491_0, i_8_337_506_0, i_8_337_518_0,
    i_8_337_528_0, i_8_337_547_0, i_8_337_586_0, i_8_337_590_0,
    i_8_337_626_0, i_8_337_632_0, i_8_337_634_0, i_8_337_658_0,
    i_8_337_670_0, i_8_337_671_0, i_8_337_694_0, i_8_337_703_0,
    i_8_337_706_0, i_8_337_716_0, i_8_337_803_0, i_8_337_824_0,
    i_8_337_830_0, i_8_337_839_0, i_8_337_844_0, i_8_337_845_0,
    i_8_337_877_0, i_8_337_1012_0, i_8_337_1028_0, i_8_337_1130_0,
    i_8_337_1225_0, i_8_337_1256_0, i_8_337_1286_0, i_8_337_1350_0,
    i_8_337_1355_0, i_8_337_1388_0, i_8_337_1420_0, i_8_337_1442_0,
    i_8_337_1445_0, i_8_337_1456_0, i_8_337_1471_0, i_8_337_1531_0,
    i_8_337_1532_0, i_8_337_1536_0, i_8_337_1537_0, i_8_337_1544_0,
    i_8_337_1576_0, i_8_337_1585_0, i_8_337_1615_0, i_8_337_1621_0,
    i_8_337_1622_0, i_8_337_1747_0, i_8_337_1751_0, i_8_337_1753_0,
    i_8_337_1768_0, i_8_337_1782_0, i_8_337_1802_0, i_8_337_1819_0,
    i_8_337_1838_0, i_8_337_1846_0, i_8_337_1847_0, i_8_337_1850_0,
    i_8_337_1892_0, i_8_337_1895_0, i_8_337_1963_0, i_8_337_1964_0,
    i_8_337_1990_0, i_8_337_1993_0, i_8_337_2000_0, i_8_337_2012_0,
    i_8_337_2047_0, i_8_337_2063_0, i_8_337_2111_0, i_8_337_2117_0,
    i_8_337_2141_0, i_8_337_2170_0, i_8_337_2227_0, i_8_337_2237_0;
  output o_8_337_0_0;
  assign o_8_337_0_0 = 0;
endmodule



// Benchmark "kernel_8_338" written by ABC on Sun Jul 19 10:08:56 2020

module kernel_8_338 ( 
    i_8_338_19_0, i_8_338_37_0, i_8_338_47_0, i_8_338_67_0, i_8_338_72_0,
    i_8_338_73_0, i_8_338_83_0, i_8_338_119_0, i_8_338_163_0,
    i_8_338_208_0, i_8_338_209_0, i_8_338_253_0, i_8_338_307_0,
    i_8_338_362_0, i_8_338_398_0, i_8_338_424_0, i_8_338_487_0,
    i_8_338_489_0, i_8_338_497_0, i_8_338_500_0, i_8_338_524_0,
    i_8_338_526_0, i_8_338_612_0, i_8_338_625_0, i_8_338_662_0,
    i_8_338_685_0, i_8_338_688_0, i_8_338_694_0, i_8_338_695_0,
    i_8_338_729_0, i_8_338_752_0, i_8_338_760_0, i_8_338_767_0,
    i_8_338_777_0, i_8_338_796_0, i_8_338_829_0, i_8_338_830_0,
    i_8_338_833_0, i_8_338_837_0, i_8_338_839_0, i_8_338_865_0,
    i_8_338_878_0, i_8_338_956_0, i_8_338_965_0, i_8_338_970_0,
    i_8_338_971_0, i_8_338_974_0, i_8_338_998_0, i_8_338_1018_0,
    i_8_338_1057_0, i_8_338_1073_0, i_8_338_1102_0, i_8_338_1171_0,
    i_8_338_1172_0, i_8_338_1234_0, i_8_338_1235_0, i_8_338_1267_0,
    i_8_338_1288_0, i_8_338_1289_0, i_8_338_1294_0, i_8_338_1307_0,
    i_8_338_1378_0, i_8_338_1400_0, i_8_338_1405_0, i_8_338_1453_0,
    i_8_338_1468_0, i_8_338_1471_0, i_8_338_1555_0, i_8_338_1559_0,
    i_8_338_1620_0, i_8_338_1639_0, i_8_338_1647_0, i_8_338_1682_0,
    i_8_338_1712_0, i_8_338_1733_0, i_8_338_1754_0, i_8_338_1760_0,
    i_8_338_1762_0, i_8_338_1775_0, i_8_338_1792_0, i_8_338_1883_0,
    i_8_338_1885_0, i_8_338_1928_0, i_8_338_1989_0, i_8_338_1997_0,
    i_8_338_2053_0, i_8_338_2054_0, i_8_338_2055_0, i_8_338_2107_0,
    i_8_338_2146_0, i_8_338_2147_0, i_8_338_2148_0, i_8_338_2149_0,
    i_8_338_2155_0, i_8_338_2162_0, i_8_338_2180_0, i_8_338_2210_0,
    i_8_338_2224_0, i_8_338_2225_0, i_8_338_2288_0,
    o_8_338_0_0  );
  input  i_8_338_19_0, i_8_338_37_0, i_8_338_47_0, i_8_338_67_0,
    i_8_338_72_0, i_8_338_73_0, i_8_338_83_0, i_8_338_119_0, i_8_338_163_0,
    i_8_338_208_0, i_8_338_209_0, i_8_338_253_0, i_8_338_307_0,
    i_8_338_362_0, i_8_338_398_0, i_8_338_424_0, i_8_338_487_0,
    i_8_338_489_0, i_8_338_497_0, i_8_338_500_0, i_8_338_524_0,
    i_8_338_526_0, i_8_338_612_0, i_8_338_625_0, i_8_338_662_0,
    i_8_338_685_0, i_8_338_688_0, i_8_338_694_0, i_8_338_695_0,
    i_8_338_729_0, i_8_338_752_0, i_8_338_760_0, i_8_338_767_0,
    i_8_338_777_0, i_8_338_796_0, i_8_338_829_0, i_8_338_830_0,
    i_8_338_833_0, i_8_338_837_0, i_8_338_839_0, i_8_338_865_0,
    i_8_338_878_0, i_8_338_956_0, i_8_338_965_0, i_8_338_970_0,
    i_8_338_971_0, i_8_338_974_0, i_8_338_998_0, i_8_338_1018_0,
    i_8_338_1057_0, i_8_338_1073_0, i_8_338_1102_0, i_8_338_1171_0,
    i_8_338_1172_0, i_8_338_1234_0, i_8_338_1235_0, i_8_338_1267_0,
    i_8_338_1288_0, i_8_338_1289_0, i_8_338_1294_0, i_8_338_1307_0,
    i_8_338_1378_0, i_8_338_1400_0, i_8_338_1405_0, i_8_338_1453_0,
    i_8_338_1468_0, i_8_338_1471_0, i_8_338_1555_0, i_8_338_1559_0,
    i_8_338_1620_0, i_8_338_1639_0, i_8_338_1647_0, i_8_338_1682_0,
    i_8_338_1712_0, i_8_338_1733_0, i_8_338_1754_0, i_8_338_1760_0,
    i_8_338_1762_0, i_8_338_1775_0, i_8_338_1792_0, i_8_338_1883_0,
    i_8_338_1885_0, i_8_338_1928_0, i_8_338_1989_0, i_8_338_1997_0,
    i_8_338_2053_0, i_8_338_2054_0, i_8_338_2055_0, i_8_338_2107_0,
    i_8_338_2146_0, i_8_338_2147_0, i_8_338_2148_0, i_8_338_2149_0,
    i_8_338_2155_0, i_8_338_2162_0, i_8_338_2180_0, i_8_338_2210_0,
    i_8_338_2224_0, i_8_338_2225_0, i_8_338_2288_0;
  output o_8_338_0_0;
  assign o_8_338_0_0 = 0;
endmodule



// Benchmark "kernel_8_339" written by ABC on Sun Jul 19 10:08:57 2020

module kernel_8_339 ( 
    i_8_339_138_0, i_8_339_146_0, i_8_339_148_0, i_8_339_189_0,
    i_8_339_227_0, i_8_339_229_0, i_8_339_273_0, i_8_339_302_0,
    i_8_339_359_0, i_8_339_366_0, i_8_339_392_0, i_8_339_432_0,
    i_8_339_455_0, i_8_339_464_0, i_8_339_470_0, i_8_339_475_0,
    i_8_339_490_0, i_8_339_503_0, i_8_339_512_0, i_8_339_529_0,
    i_8_339_551_0, i_8_339_583_0, i_8_339_592_0, i_8_339_595_0,
    i_8_339_610_0, i_8_339_614_0, i_8_339_637_0, i_8_339_656_0,
    i_8_339_679_0, i_8_339_718_0, i_8_339_751_0, i_8_339_812_0,
    i_8_339_819_0, i_8_339_827_0, i_8_339_860_0, i_8_339_863_0,
    i_8_339_866_0, i_8_339_874_0, i_8_339_914_0, i_8_339_917_0,
    i_8_339_985_0, i_8_339_1046_0, i_8_339_1055_0, i_8_339_1058_0,
    i_8_339_1174_0, i_8_339_1181_0, i_8_339_1188_0, i_8_339_1205_0,
    i_8_339_1243_0, i_8_339_1298_0, i_8_339_1305_0, i_8_339_1306_0,
    i_8_339_1311_0, i_8_339_1329_0, i_8_339_1334_0, i_8_339_1343_0,
    i_8_339_1354_0, i_8_339_1391_0, i_8_339_1410_0, i_8_339_1420_0,
    i_8_339_1470_0, i_8_339_1471_0, i_8_339_1487_0, i_8_339_1498_0,
    i_8_339_1502_0, i_8_339_1541_0, i_8_339_1554_0, i_8_339_1559_0,
    i_8_339_1637_0, i_8_339_1642_0, i_8_339_1647_0, i_8_339_1667_0,
    i_8_339_1675_0, i_8_339_1676_0, i_8_339_1703_0, i_8_339_1750_0,
    i_8_339_1751_0, i_8_339_1766_0, i_8_339_1780_0, i_8_339_1784_0,
    i_8_339_1838_0, i_8_339_1844_0, i_8_339_1919_0, i_8_339_1930_0,
    i_8_339_1973_0, i_8_339_1989_0, i_8_339_1993_0, i_8_339_1997_0,
    i_8_339_2000_0, i_8_339_2042_0, i_8_339_2056_0, i_8_339_2065_0,
    i_8_339_2066_0, i_8_339_2147_0, i_8_339_2191_0, i_8_339_2234_0,
    i_8_339_2242_0, i_8_339_2248_0, i_8_339_2249_0, i_8_339_2268_0,
    o_8_339_0_0  );
  input  i_8_339_138_0, i_8_339_146_0, i_8_339_148_0, i_8_339_189_0,
    i_8_339_227_0, i_8_339_229_0, i_8_339_273_0, i_8_339_302_0,
    i_8_339_359_0, i_8_339_366_0, i_8_339_392_0, i_8_339_432_0,
    i_8_339_455_0, i_8_339_464_0, i_8_339_470_0, i_8_339_475_0,
    i_8_339_490_0, i_8_339_503_0, i_8_339_512_0, i_8_339_529_0,
    i_8_339_551_0, i_8_339_583_0, i_8_339_592_0, i_8_339_595_0,
    i_8_339_610_0, i_8_339_614_0, i_8_339_637_0, i_8_339_656_0,
    i_8_339_679_0, i_8_339_718_0, i_8_339_751_0, i_8_339_812_0,
    i_8_339_819_0, i_8_339_827_0, i_8_339_860_0, i_8_339_863_0,
    i_8_339_866_0, i_8_339_874_0, i_8_339_914_0, i_8_339_917_0,
    i_8_339_985_0, i_8_339_1046_0, i_8_339_1055_0, i_8_339_1058_0,
    i_8_339_1174_0, i_8_339_1181_0, i_8_339_1188_0, i_8_339_1205_0,
    i_8_339_1243_0, i_8_339_1298_0, i_8_339_1305_0, i_8_339_1306_0,
    i_8_339_1311_0, i_8_339_1329_0, i_8_339_1334_0, i_8_339_1343_0,
    i_8_339_1354_0, i_8_339_1391_0, i_8_339_1410_0, i_8_339_1420_0,
    i_8_339_1470_0, i_8_339_1471_0, i_8_339_1487_0, i_8_339_1498_0,
    i_8_339_1502_0, i_8_339_1541_0, i_8_339_1554_0, i_8_339_1559_0,
    i_8_339_1637_0, i_8_339_1642_0, i_8_339_1647_0, i_8_339_1667_0,
    i_8_339_1675_0, i_8_339_1676_0, i_8_339_1703_0, i_8_339_1750_0,
    i_8_339_1751_0, i_8_339_1766_0, i_8_339_1780_0, i_8_339_1784_0,
    i_8_339_1838_0, i_8_339_1844_0, i_8_339_1919_0, i_8_339_1930_0,
    i_8_339_1973_0, i_8_339_1989_0, i_8_339_1993_0, i_8_339_1997_0,
    i_8_339_2000_0, i_8_339_2042_0, i_8_339_2056_0, i_8_339_2065_0,
    i_8_339_2066_0, i_8_339_2147_0, i_8_339_2191_0, i_8_339_2234_0,
    i_8_339_2242_0, i_8_339_2248_0, i_8_339_2249_0, i_8_339_2268_0;
  output o_8_339_0_0;
  assign o_8_339_0_0 = 0;
endmodule



// Benchmark "kernel_8_340" written by ABC on Sun Jul 19 10:08:58 2020

module kernel_8_340 ( 
    i_8_340_10_0, i_8_340_18_0, i_8_340_28_0, i_8_340_49_0, i_8_340_73_0,
    i_8_340_135_0, i_8_340_156_0, i_8_340_183_0, i_8_340_229_0,
    i_8_340_252_0, i_8_340_265_0, i_8_340_288_0, i_8_340_370_0,
    i_8_340_387_0, i_8_340_421_0, i_8_340_435_0, i_8_340_472_0,
    i_8_340_473_0, i_8_340_493_0, i_8_340_507_0, i_8_340_543_0,
    i_8_340_546_0, i_8_340_550_0, i_8_340_595_0, i_8_340_608_0,
    i_8_340_611_0, i_8_340_625_0, i_8_340_633_0, i_8_340_660_0,
    i_8_340_661_0, i_8_340_663_0, i_8_340_684_0, i_8_340_687_0,
    i_8_340_690_0, i_8_340_711_0, i_8_340_756_0, i_8_340_765_0,
    i_8_340_769_0, i_8_340_781_0, i_8_340_783_0, i_8_340_786_0,
    i_8_340_806_0, i_8_340_819_0, i_8_340_820_0, i_8_340_822_0,
    i_8_340_847_0, i_8_340_865_0, i_8_340_873_0, i_8_340_891_0,
    i_8_340_892_0, i_8_340_946_0, i_8_340_975_0, i_8_340_984_0,
    i_8_340_1009_0, i_8_340_1065_0, i_8_340_1107_0, i_8_340_1126_0,
    i_8_340_1127_0, i_8_340_1144_0, i_8_340_1159_0, i_8_340_1215_0,
    i_8_340_1245_0, i_8_340_1260_0, i_8_340_1286_0, i_8_340_1305_0,
    i_8_340_1341_0, i_8_340_1416_0, i_8_340_1417_0, i_8_340_1440_0,
    i_8_340_1471_0, i_8_340_1549_0, i_8_340_1557_0, i_8_340_1565_0,
    i_8_340_1629_0, i_8_340_1633_0, i_8_340_1671_0, i_8_340_1674_0,
    i_8_340_1677_0, i_8_340_1682_0, i_8_340_1702_0, i_8_340_1710_0,
    i_8_340_1719_0, i_8_340_1737_0, i_8_340_1750_0, i_8_340_1758_0,
    i_8_340_1783_0, i_8_340_1788_0, i_8_340_1803_0, i_8_340_1808_0,
    i_8_340_1854_0, i_8_340_1857_0, i_8_340_1861_0, i_8_340_1893_0,
    i_8_340_1995_0, i_8_340_2025_0, i_8_340_2089_0, i_8_340_2110_0,
    i_8_340_2181_0, i_8_340_2298_0, i_8_340_2299_0,
    o_8_340_0_0  );
  input  i_8_340_10_0, i_8_340_18_0, i_8_340_28_0, i_8_340_49_0,
    i_8_340_73_0, i_8_340_135_0, i_8_340_156_0, i_8_340_183_0,
    i_8_340_229_0, i_8_340_252_0, i_8_340_265_0, i_8_340_288_0,
    i_8_340_370_0, i_8_340_387_0, i_8_340_421_0, i_8_340_435_0,
    i_8_340_472_0, i_8_340_473_0, i_8_340_493_0, i_8_340_507_0,
    i_8_340_543_0, i_8_340_546_0, i_8_340_550_0, i_8_340_595_0,
    i_8_340_608_0, i_8_340_611_0, i_8_340_625_0, i_8_340_633_0,
    i_8_340_660_0, i_8_340_661_0, i_8_340_663_0, i_8_340_684_0,
    i_8_340_687_0, i_8_340_690_0, i_8_340_711_0, i_8_340_756_0,
    i_8_340_765_0, i_8_340_769_0, i_8_340_781_0, i_8_340_783_0,
    i_8_340_786_0, i_8_340_806_0, i_8_340_819_0, i_8_340_820_0,
    i_8_340_822_0, i_8_340_847_0, i_8_340_865_0, i_8_340_873_0,
    i_8_340_891_0, i_8_340_892_0, i_8_340_946_0, i_8_340_975_0,
    i_8_340_984_0, i_8_340_1009_0, i_8_340_1065_0, i_8_340_1107_0,
    i_8_340_1126_0, i_8_340_1127_0, i_8_340_1144_0, i_8_340_1159_0,
    i_8_340_1215_0, i_8_340_1245_0, i_8_340_1260_0, i_8_340_1286_0,
    i_8_340_1305_0, i_8_340_1341_0, i_8_340_1416_0, i_8_340_1417_0,
    i_8_340_1440_0, i_8_340_1471_0, i_8_340_1549_0, i_8_340_1557_0,
    i_8_340_1565_0, i_8_340_1629_0, i_8_340_1633_0, i_8_340_1671_0,
    i_8_340_1674_0, i_8_340_1677_0, i_8_340_1682_0, i_8_340_1702_0,
    i_8_340_1710_0, i_8_340_1719_0, i_8_340_1737_0, i_8_340_1750_0,
    i_8_340_1758_0, i_8_340_1783_0, i_8_340_1788_0, i_8_340_1803_0,
    i_8_340_1808_0, i_8_340_1854_0, i_8_340_1857_0, i_8_340_1861_0,
    i_8_340_1893_0, i_8_340_1995_0, i_8_340_2025_0, i_8_340_2089_0,
    i_8_340_2110_0, i_8_340_2181_0, i_8_340_2298_0, i_8_340_2299_0;
  output o_8_340_0_0;
  assign o_8_340_0_0 = 0;
endmodule



// Benchmark "kernel_8_341" written by ABC on Sun Jul 19 10:09:00 2020

module kernel_8_341 ( 
    i_8_341_27_0, i_8_341_45_0, i_8_341_49_0, i_8_341_82_0, i_8_341_111_0,
    i_8_341_162_0, i_8_341_190_0, i_8_341_216_0, i_8_341_217_0,
    i_8_341_220_0, i_8_341_223_0, i_8_341_229_0, i_8_341_237_0,
    i_8_341_253_0, i_8_341_257_0, i_8_341_325_0, i_8_341_361_0,
    i_8_341_363_0, i_8_341_364_0, i_8_341_388_0, i_8_341_414_0,
    i_8_341_425_0, i_8_341_436_0, i_8_341_451_0, i_8_341_452_0,
    i_8_341_461_0, i_8_341_493_0, i_8_341_570_0, i_8_341_571_0,
    i_8_341_607_0, i_8_341_608_0, i_8_341_631_0, i_8_341_661_0,
    i_8_341_687_0, i_8_341_694_0, i_8_341_732_0, i_8_341_735_0,
    i_8_341_756_0, i_8_341_758_0, i_8_341_767_0, i_8_341_803_0,
    i_8_341_811_0, i_8_341_840_0, i_8_341_841_0, i_8_341_842_0,
    i_8_341_856_0, i_8_341_876_0, i_8_341_919_0, i_8_341_936_0,
    i_8_341_937_0, i_8_341_938_0, i_8_341_991_0, i_8_341_995_0,
    i_8_341_996_0, i_8_341_1008_0, i_8_341_1155_0, i_8_341_1179_0,
    i_8_341_1180_0, i_8_341_1181_0, i_8_341_1182_0, i_8_341_1189_0,
    i_8_341_1224_0, i_8_341_1234_0, i_8_341_1282_0, i_8_341_1305_0,
    i_8_341_1333_0, i_8_341_1335_0, i_8_341_1407_0, i_8_341_1467_0,
    i_8_341_1486_0, i_8_341_1492_0, i_8_341_1493_0, i_8_341_1549_0,
    i_8_341_1621_0, i_8_341_1631_0, i_8_341_1635_0, i_8_341_1649_0,
    i_8_341_1674_0, i_8_341_1692_0, i_8_341_1694_0, i_8_341_1730_0,
    i_8_341_1740_0, i_8_341_1748_0, i_8_341_1758_0, i_8_341_1759_0,
    i_8_341_1783_0, i_8_341_1797_0, i_8_341_1819_0, i_8_341_1821_0,
    i_8_341_1822_0, i_8_341_1993_0, i_8_341_2029_0, i_8_341_2054_0,
    i_8_341_2073_0, i_8_341_2187_0, i_8_341_2245_0, i_8_341_2271_0,
    i_8_341_2295_0, i_8_341_2296_0, i_8_341_2297_0,
    o_8_341_0_0  );
  input  i_8_341_27_0, i_8_341_45_0, i_8_341_49_0, i_8_341_82_0,
    i_8_341_111_0, i_8_341_162_0, i_8_341_190_0, i_8_341_216_0,
    i_8_341_217_0, i_8_341_220_0, i_8_341_223_0, i_8_341_229_0,
    i_8_341_237_0, i_8_341_253_0, i_8_341_257_0, i_8_341_325_0,
    i_8_341_361_0, i_8_341_363_0, i_8_341_364_0, i_8_341_388_0,
    i_8_341_414_0, i_8_341_425_0, i_8_341_436_0, i_8_341_451_0,
    i_8_341_452_0, i_8_341_461_0, i_8_341_493_0, i_8_341_570_0,
    i_8_341_571_0, i_8_341_607_0, i_8_341_608_0, i_8_341_631_0,
    i_8_341_661_0, i_8_341_687_0, i_8_341_694_0, i_8_341_732_0,
    i_8_341_735_0, i_8_341_756_0, i_8_341_758_0, i_8_341_767_0,
    i_8_341_803_0, i_8_341_811_0, i_8_341_840_0, i_8_341_841_0,
    i_8_341_842_0, i_8_341_856_0, i_8_341_876_0, i_8_341_919_0,
    i_8_341_936_0, i_8_341_937_0, i_8_341_938_0, i_8_341_991_0,
    i_8_341_995_0, i_8_341_996_0, i_8_341_1008_0, i_8_341_1155_0,
    i_8_341_1179_0, i_8_341_1180_0, i_8_341_1181_0, i_8_341_1182_0,
    i_8_341_1189_0, i_8_341_1224_0, i_8_341_1234_0, i_8_341_1282_0,
    i_8_341_1305_0, i_8_341_1333_0, i_8_341_1335_0, i_8_341_1407_0,
    i_8_341_1467_0, i_8_341_1486_0, i_8_341_1492_0, i_8_341_1493_0,
    i_8_341_1549_0, i_8_341_1621_0, i_8_341_1631_0, i_8_341_1635_0,
    i_8_341_1649_0, i_8_341_1674_0, i_8_341_1692_0, i_8_341_1694_0,
    i_8_341_1730_0, i_8_341_1740_0, i_8_341_1748_0, i_8_341_1758_0,
    i_8_341_1759_0, i_8_341_1783_0, i_8_341_1797_0, i_8_341_1819_0,
    i_8_341_1821_0, i_8_341_1822_0, i_8_341_1993_0, i_8_341_2029_0,
    i_8_341_2054_0, i_8_341_2073_0, i_8_341_2187_0, i_8_341_2245_0,
    i_8_341_2271_0, i_8_341_2295_0, i_8_341_2296_0, i_8_341_2297_0;
  output o_8_341_0_0;
  assign o_8_341_0_0 = ~((~i_8_341_27_0 & ((~i_8_341_162_0 & i_8_341_216_0 & ~i_8_341_571_0 & ~i_8_341_1181_0) | (~i_8_341_570_0 & i_8_341_661_0 & ~i_8_341_936_0 & ~i_8_341_1621_0 & ~i_8_341_2187_0))) | (~i_8_341_631_0 & ((~i_8_341_111_0 & ~i_8_341_856_0 & ~i_8_341_1182_0 & ~i_8_341_1282_0 & ~i_8_341_1692_0 & ~i_8_341_1694_0 & ~i_8_341_1759_0 & ~i_8_341_1783_0 & ~i_8_341_2054_0 & ~i_8_341_2245_0) | (~i_8_341_803_0 & ~i_8_341_1407_0 & i_8_341_1549_0 & ~i_8_341_1621_0 & ~i_8_341_2295_0 & ~i_8_341_2296_0))) | (~i_8_341_1181_0 & ((~i_8_341_111_0 & ((~i_8_341_694_0 & ~i_8_341_1234_0 & ~i_8_341_1333_0 & ~i_8_341_1740_0 & ~i_8_341_1758_0) | (~i_8_341_607_0 & ~i_8_341_936_0 & ~i_8_341_937_0 & ~i_8_341_991_0 & ~i_8_341_1649_0 & ~i_8_341_1674_0 & ~i_8_341_1694_0 & ~i_8_341_2073_0 & ~i_8_341_2245_0))) | (~i_8_341_229_0 & i_8_341_363_0) | (~i_8_341_493_0 & i_8_341_842_0 & ~i_8_341_1234_0 & i_8_341_1282_0 & ~i_8_341_2296_0))) | (~i_8_341_607_0 & ((~i_8_341_938_0 & ~i_8_341_991_0 & ~i_8_341_1748_0 & ~i_8_341_1759_0 & i_8_341_2054_0) | (i_8_341_220_0 & ~i_8_341_1182_0 & ~i_8_341_1224_0 & ~i_8_341_1282_0 & ~i_8_341_1635_0 & ~i_8_341_2054_0))) | (~i_8_341_937_0 & ((~i_8_341_687_0 & ((~i_8_341_49_0 & i_8_341_607_0 & ~i_8_341_758_0 & ~i_8_341_938_0 & ~i_8_341_2295_0) | (~i_8_341_661_0 & ~i_8_341_694_0 & ~i_8_341_842_0 & ~i_8_341_991_0 & ~i_8_341_1305_0 & ~i_8_341_1335_0 & ~i_8_341_1631_0 & ~i_8_341_1759_0 & ~i_8_341_2297_0))) | (~i_8_341_936_0 & ~i_8_341_1740_0 & i_8_341_1822_0) | (~i_8_341_570_0 & i_8_341_876_0 & ~i_8_341_1179_0 & ~i_8_341_1282_0 & ~i_8_341_2296_0))) | (~i_8_341_570_0 & ((~i_8_341_841_0 & ~i_8_341_938_0 & ~i_8_341_1335_0 & ~i_8_341_1407_0 & ~i_8_341_1621_0 & ~i_8_341_1649_0 & ~i_8_341_1692_0 & ~i_8_341_1758_0) | (~i_8_341_414_0 & i_8_341_451_0 & ~i_8_341_756_0 & i_8_341_1282_0 & ~i_8_341_2296_0 & ~i_8_341_758_0 & ~i_8_341_995_0))) | (~i_8_341_938_0 & ((~i_8_341_811_0 & ~i_8_341_991_0 & i_8_341_995_0 & ~i_8_341_1333_0) | (~i_8_341_936_0 & ~i_8_341_1179_0 & ~i_8_341_1407_0 & ~i_8_341_1621_0 & ~i_8_341_1730_0 & i_8_341_1783_0))) | (i_8_341_1492_0 & ((i_8_341_1493_0 & i_8_341_1740_0) | (~i_8_341_996_0 & ~i_8_341_1730_0 & ~i_8_341_1740_0))) | (~i_8_341_1674_0 & ((i_8_341_223_0 & ~i_8_341_363_0 & ~i_8_341_1180_0) | (~i_8_341_216_0 & ~i_8_341_1694_0 & i_8_341_1748_0 & ~i_8_341_1783_0))) | (i_8_341_436_0 & ~i_8_341_1335_0 & ~i_8_341_1621_0) | (i_8_341_1649_0 & i_8_341_1819_0) | (i_8_341_493_0 & ~i_8_341_2073_0) | (~i_8_341_856_0 & i_8_341_2271_0) | (i_8_341_237_0 & ~i_8_341_842_0 & ~i_8_341_1467_0 & ~i_8_341_1730_0 & i_8_341_1740_0 & ~i_8_341_1758_0 & ~i_8_341_2295_0));
endmodule



// Benchmark "kernel_8_342" written by ABC on Sun Jul 19 10:09:00 2020

module kernel_8_342 ( 
    i_8_342_25_0, i_8_342_34_0, i_8_342_81_0, i_8_342_87_0, i_8_342_89_0,
    i_8_342_93_0, i_8_342_106_0, i_8_342_160_0, i_8_342_183_0,
    i_8_342_262_0, i_8_342_291_0, i_8_342_307_0, i_8_342_328_0,
    i_8_342_378_0, i_8_342_403_0, i_8_342_433_0, i_8_342_462_0,
    i_8_342_503_0, i_8_342_523_0, i_8_342_554_0, i_8_342_572_0,
    i_8_342_595_0, i_8_342_621_0, i_8_342_624_0, i_8_342_633_0,
    i_8_342_634_0, i_8_342_637_0, i_8_342_669_0, i_8_342_670_0,
    i_8_342_690_0, i_8_342_707_0, i_8_342_712_0, i_8_342_756_0,
    i_8_342_762_0, i_8_342_767_0, i_8_342_777_0, i_8_342_778_0,
    i_8_342_783_0, i_8_342_803_0, i_8_342_823_0, i_8_342_873_0,
    i_8_342_971_0, i_8_342_973_0, i_8_342_987_0, i_8_342_1026_0,
    i_8_342_1029_0, i_8_342_1111_0, i_8_342_1119_0, i_8_342_1171_0,
    i_8_342_1172_0, i_8_342_1219_0, i_8_342_1236_0, i_8_342_1254_0,
    i_8_342_1282_0, i_8_342_1285_0, i_8_342_1305_0, i_8_342_1314_0,
    i_8_342_1317_0, i_8_342_1402_0, i_8_342_1424_0, i_8_342_1441_0,
    i_8_342_1474_0, i_8_342_1476_0, i_8_342_1482_0, i_8_342_1545_0,
    i_8_342_1547_0, i_8_342_1563_0, i_8_342_1579_0, i_8_342_1585_0,
    i_8_342_1587_0, i_8_342_1600_0, i_8_342_1651_0, i_8_342_1663_0,
    i_8_342_1668_0, i_8_342_1671_0, i_8_342_1680_0, i_8_342_1681_0,
    i_8_342_1695_0, i_8_342_1698_0, i_8_342_1708_0, i_8_342_1746_0,
    i_8_342_1751_0, i_8_342_1792_0, i_8_342_1804_0, i_8_342_1822_0,
    i_8_342_1841_0, i_8_342_1902_0, i_8_342_1912_0, i_8_342_1947_0,
    i_8_342_2107_0, i_8_342_2109_0, i_8_342_2128_0, i_8_342_2136_0,
    i_8_342_2146_0, i_8_342_2190_0, i_8_342_2226_0, i_8_342_2244_0,
    i_8_342_2291_0, i_8_342_2292_0, i_8_342_2295_0,
    o_8_342_0_0  );
  input  i_8_342_25_0, i_8_342_34_0, i_8_342_81_0, i_8_342_87_0,
    i_8_342_89_0, i_8_342_93_0, i_8_342_106_0, i_8_342_160_0,
    i_8_342_183_0, i_8_342_262_0, i_8_342_291_0, i_8_342_307_0,
    i_8_342_328_0, i_8_342_378_0, i_8_342_403_0, i_8_342_433_0,
    i_8_342_462_0, i_8_342_503_0, i_8_342_523_0, i_8_342_554_0,
    i_8_342_572_0, i_8_342_595_0, i_8_342_621_0, i_8_342_624_0,
    i_8_342_633_0, i_8_342_634_0, i_8_342_637_0, i_8_342_669_0,
    i_8_342_670_0, i_8_342_690_0, i_8_342_707_0, i_8_342_712_0,
    i_8_342_756_0, i_8_342_762_0, i_8_342_767_0, i_8_342_777_0,
    i_8_342_778_0, i_8_342_783_0, i_8_342_803_0, i_8_342_823_0,
    i_8_342_873_0, i_8_342_971_0, i_8_342_973_0, i_8_342_987_0,
    i_8_342_1026_0, i_8_342_1029_0, i_8_342_1111_0, i_8_342_1119_0,
    i_8_342_1171_0, i_8_342_1172_0, i_8_342_1219_0, i_8_342_1236_0,
    i_8_342_1254_0, i_8_342_1282_0, i_8_342_1285_0, i_8_342_1305_0,
    i_8_342_1314_0, i_8_342_1317_0, i_8_342_1402_0, i_8_342_1424_0,
    i_8_342_1441_0, i_8_342_1474_0, i_8_342_1476_0, i_8_342_1482_0,
    i_8_342_1545_0, i_8_342_1547_0, i_8_342_1563_0, i_8_342_1579_0,
    i_8_342_1585_0, i_8_342_1587_0, i_8_342_1600_0, i_8_342_1651_0,
    i_8_342_1663_0, i_8_342_1668_0, i_8_342_1671_0, i_8_342_1680_0,
    i_8_342_1681_0, i_8_342_1695_0, i_8_342_1698_0, i_8_342_1708_0,
    i_8_342_1746_0, i_8_342_1751_0, i_8_342_1792_0, i_8_342_1804_0,
    i_8_342_1822_0, i_8_342_1841_0, i_8_342_1902_0, i_8_342_1912_0,
    i_8_342_1947_0, i_8_342_2107_0, i_8_342_2109_0, i_8_342_2128_0,
    i_8_342_2136_0, i_8_342_2146_0, i_8_342_2190_0, i_8_342_2226_0,
    i_8_342_2244_0, i_8_342_2291_0, i_8_342_2292_0, i_8_342_2295_0;
  output o_8_342_0_0;
  assign o_8_342_0_0 = 0;
endmodule



// Benchmark "kernel_8_343" written by ABC on Sun Jul 19 10:09:01 2020

module kernel_8_343 ( 
    i_8_343_36_0, i_8_343_135_0, i_8_343_172_0, i_8_343_193_0,
    i_8_343_226_0, i_8_343_261_0, i_8_343_309_0, i_8_343_321_0,
    i_8_343_345_0, i_8_343_364_0, i_8_343_396_0, i_8_343_414_0,
    i_8_343_417_0, i_8_343_418_0, i_8_343_422_0, i_8_343_453_0,
    i_8_343_472_0, i_8_343_480_0, i_8_343_504_0, i_8_343_507_0,
    i_8_343_508_0, i_8_343_522_0, i_8_343_523_0, i_8_343_525_0,
    i_8_343_534_0, i_8_343_552_0, i_8_343_567_0, i_8_343_571_0,
    i_8_343_573_0, i_8_343_579_0, i_8_343_582_0, i_8_343_604_0,
    i_8_343_625_0, i_8_343_696_0, i_8_343_702_0, i_8_343_751_0,
    i_8_343_756_0, i_8_343_759_0, i_8_343_823_0, i_8_343_891_0,
    i_8_343_963_0, i_8_343_1009_0, i_8_343_1098_0, i_8_343_1103_0,
    i_8_343_1128_0, i_8_343_1134_0, i_8_343_1179_0, i_8_343_1197_0,
    i_8_343_1234_0, i_8_343_1263_0, i_8_343_1266_0, i_8_343_1314_0,
    i_8_343_1362_0, i_8_343_1422_0, i_8_343_1440_0, i_8_343_1461_0,
    i_8_343_1464_0, i_8_343_1465_0, i_8_343_1485_0, i_8_343_1512_0,
    i_8_343_1513_0, i_8_343_1521_0, i_8_343_1522_0, i_8_343_1540_0,
    i_8_343_1544_0, i_8_343_1569_0, i_8_343_1597_0, i_8_343_1606_0,
    i_8_343_1629_0, i_8_343_1665_0, i_8_343_1692_0, i_8_343_1693_0,
    i_8_343_1696_0, i_8_343_1723_0, i_8_343_1765_0, i_8_343_1784_0,
    i_8_343_1794_0, i_8_343_1803_0, i_8_343_1804_0, i_8_343_1830_0,
    i_8_343_1836_0, i_8_343_1840_0, i_8_343_1887_0, i_8_343_1899_0,
    i_8_343_1911_0, i_8_343_1927_0, i_8_343_1935_0, i_8_343_1938_0,
    i_8_343_1956_0, i_8_343_1974_0, i_8_343_1992_0, i_8_343_1993_0,
    i_8_343_2070_0, i_8_343_2079_0, i_8_343_2107_0, i_8_343_2141_0,
    i_8_343_2151_0, i_8_343_2163_0, i_8_343_2208_0, i_8_343_2232_0,
    o_8_343_0_0  );
  input  i_8_343_36_0, i_8_343_135_0, i_8_343_172_0, i_8_343_193_0,
    i_8_343_226_0, i_8_343_261_0, i_8_343_309_0, i_8_343_321_0,
    i_8_343_345_0, i_8_343_364_0, i_8_343_396_0, i_8_343_414_0,
    i_8_343_417_0, i_8_343_418_0, i_8_343_422_0, i_8_343_453_0,
    i_8_343_472_0, i_8_343_480_0, i_8_343_504_0, i_8_343_507_0,
    i_8_343_508_0, i_8_343_522_0, i_8_343_523_0, i_8_343_525_0,
    i_8_343_534_0, i_8_343_552_0, i_8_343_567_0, i_8_343_571_0,
    i_8_343_573_0, i_8_343_579_0, i_8_343_582_0, i_8_343_604_0,
    i_8_343_625_0, i_8_343_696_0, i_8_343_702_0, i_8_343_751_0,
    i_8_343_756_0, i_8_343_759_0, i_8_343_823_0, i_8_343_891_0,
    i_8_343_963_0, i_8_343_1009_0, i_8_343_1098_0, i_8_343_1103_0,
    i_8_343_1128_0, i_8_343_1134_0, i_8_343_1179_0, i_8_343_1197_0,
    i_8_343_1234_0, i_8_343_1263_0, i_8_343_1266_0, i_8_343_1314_0,
    i_8_343_1362_0, i_8_343_1422_0, i_8_343_1440_0, i_8_343_1461_0,
    i_8_343_1464_0, i_8_343_1465_0, i_8_343_1485_0, i_8_343_1512_0,
    i_8_343_1513_0, i_8_343_1521_0, i_8_343_1522_0, i_8_343_1540_0,
    i_8_343_1544_0, i_8_343_1569_0, i_8_343_1597_0, i_8_343_1606_0,
    i_8_343_1629_0, i_8_343_1665_0, i_8_343_1692_0, i_8_343_1693_0,
    i_8_343_1696_0, i_8_343_1723_0, i_8_343_1765_0, i_8_343_1784_0,
    i_8_343_1794_0, i_8_343_1803_0, i_8_343_1804_0, i_8_343_1830_0,
    i_8_343_1836_0, i_8_343_1840_0, i_8_343_1887_0, i_8_343_1899_0,
    i_8_343_1911_0, i_8_343_1927_0, i_8_343_1935_0, i_8_343_1938_0,
    i_8_343_1956_0, i_8_343_1974_0, i_8_343_1992_0, i_8_343_1993_0,
    i_8_343_2070_0, i_8_343_2079_0, i_8_343_2107_0, i_8_343_2141_0,
    i_8_343_2151_0, i_8_343_2163_0, i_8_343_2208_0, i_8_343_2232_0;
  output o_8_343_0_0;
  assign o_8_343_0_0 = ~(~i_8_343_1521_0 | ~i_8_343_1830_0 | ~i_8_343_1362_0 | ~i_8_343_261_0 | ~i_8_343_396_0);
endmodule



// Benchmark "kernel_8_344" written by ABC on Sun Jul 19 10:09:02 2020

module kernel_8_344 ( 
    i_8_344_34_0, i_8_344_76_0, i_8_344_103_0, i_8_344_115_0,
    i_8_344_119_0, i_8_344_121_0, i_8_344_166_0, i_8_344_167_0,
    i_8_344_220_0, i_8_344_229_0, i_8_344_245_0, i_8_344_281_0,
    i_8_344_301_0, i_8_344_320_0, i_8_344_323_0, i_8_344_324_0,
    i_8_344_326_0, i_8_344_338_0, i_8_344_371_0, i_8_344_437_0,
    i_8_344_504_0, i_8_344_523_0, i_8_344_525_0, i_8_344_527_0,
    i_8_344_529_0, i_8_344_543_0, i_8_344_562_0, i_8_344_563_0,
    i_8_344_566_0, i_8_344_583_0, i_8_344_604_0, i_8_344_605_0,
    i_8_344_626_0, i_8_344_679_0, i_8_344_722_0, i_8_344_729_0,
    i_8_344_760_0, i_8_344_761_0, i_8_344_785_0, i_8_344_795_0,
    i_8_344_796_0, i_8_344_806_0, i_8_344_832_0, i_8_344_840_0,
    i_8_344_932_0, i_8_344_1049_0, i_8_344_1072_0, i_8_344_1073_0,
    i_8_344_1109_0, i_8_344_1111_0, i_8_344_1127_0, i_8_344_1154_0,
    i_8_344_1180_0, i_8_344_1277_0, i_8_344_1282_0, i_8_344_1298_0,
    i_8_344_1334_0, i_8_344_1346_0, i_8_344_1360_0, i_8_344_1361_0,
    i_8_344_1364_0, i_8_344_1381_0, i_8_344_1450_0, i_8_344_1454_0,
    i_8_344_1469_0, i_8_344_1477_0, i_8_344_1478_0, i_8_344_1481_0,
    i_8_344_1543_0, i_8_344_1544_0, i_8_344_1552_0, i_8_344_1553_0,
    i_8_344_1684_0, i_8_344_1701_0, i_8_344_1711_0, i_8_344_1733_0,
    i_8_344_1747_0, i_8_344_1767_0, i_8_344_1768_0, i_8_344_1787_0,
    i_8_344_1822_0, i_8_344_1846_0, i_8_344_1856_0, i_8_344_1859_0,
    i_8_344_1864_0, i_8_344_1919_0, i_8_344_1943_0, i_8_344_1975_0,
    i_8_344_1996_0, i_8_344_2056_0, i_8_344_2074_0, i_8_344_2075_0,
    i_8_344_2133_0, i_8_344_2141_0, i_8_344_2156_0, i_8_344_2171_0,
    i_8_344_2192_0, i_8_344_2223_0, i_8_344_2282_0, i_8_344_2296_0,
    o_8_344_0_0  );
  input  i_8_344_34_0, i_8_344_76_0, i_8_344_103_0, i_8_344_115_0,
    i_8_344_119_0, i_8_344_121_0, i_8_344_166_0, i_8_344_167_0,
    i_8_344_220_0, i_8_344_229_0, i_8_344_245_0, i_8_344_281_0,
    i_8_344_301_0, i_8_344_320_0, i_8_344_323_0, i_8_344_324_0,
    i_8_344_326_0, i_8_344_338_0, i_8_344_371_0, i_8_344_437_0,
    i_8_344_504_0, i_8_344_523_0, i_8_344_525_0, i_8_344_527_0,
    i_8_344_529_0, i_8_344_543_0, i_8_344_562_0, i_8_344_563_0,
    i_8_344_566_0, i_8_344_583_0, i_8_344_604_0, i_8_344_605_0,
    i_8_344_626_0, i_8_344_679_0, i_8_344_722_0, i_8_344_729_0,
    i_8_344_760_0, i_8_344_761_0, i_8_344_785_0, i_8_344_795_0,
    i_8_344_796_0, i_8_344_806_0, i_8_344_832_0, i_8_344_840_0,
    i_8_344_932_0, i_8_344_1049_0, i_8_344_1072_0, i_8_344_1073_0,
    i_8_344_1109_0, i_8_344_1111_0, i_8_344_1127_0, i_8_344_1154_0,
    i_8_344_1180_0, i_8_344_1277_0, i_8_344_1282_0, i_8_344_1298_0,
    i_8_344_1334_0, i_8_344_1346_0, i_8_344_1360_0, i_8_344_1361_0,
    i_8_344_1364_0, i_8_344_1381_0, i_8_344_1450_0, i_8_344_1454_0,
    i_8_344_1469_0, i_8_344_1477_0, i_8_344_1478_0, i_8_344_1481_0,
    i_8_344_1543_0, i_8_344_1544_0, i_8_344_1552_0, i_8_344_1553_0,
    i_8_344_1684_0, i_8_344_1701_0, i_8_344_1711_0, i_8_344_1733_0,
    i_8_344_1747_0, i_8_344_1767_0, i_8_344_1768_0, i_8_344_1787_0,
    i_8_344_1822_0, i_8_344_1846_0, i_8_344_1856_0, i_8_344_1859_0,
    i_8_344_1864_0, i_8_344_1919_0, i_8_344_1943_0, i_8_344_1975_0,
    i_8_344_1996_0, i_8_344_2056_0, i_8_344_2074_0, i_8_344_2075_0,
    i_8_344_2133_0, i_8_344_2141_0, i_8_344_2156_0, i_8_344_2171_0,
    i_8_344_2192_0, i_8_344_2223_0, i_8_344_2282_0, i_8_344_2296_0;
  output o_8_344_0_0;
  assign o_8_344_0_0 = 0;
endmodule



// Benchmark "kernel_8_345" written by ABC on Sun Jul 19 10:09:03 2020

module kernel_8_345 ( 
    i_8_345_84_0, i_8_345_85_0, i_8_345_96_0, i_8_345_106_0, i_8_345_138_0,
    i_8_345_245_0, i_8_345_291_0, i_8_345_294_0, i_8_345_304_0,
    i_8_345_327_0, i_8_345_372_0, i_8_345_375_0, i_8_345_381_0,
    i_8_345_384_0, i_8_345_385_0, i_8_345_419_0, i_8_345_436_0,
    i_8_345_462_0, i_8_345_475_0, i_8_345_480_0, i_8_345_481_0,
    i_8_345_483_0, i_8_345_523_0, i_8_345_526_0, i_8_345_598_0,
    i_8_345_599_0, i_8_345_601_0, i_8_345_672_0, i_8_345_699_0,
    i_8_345_759_0, i_8_345_780_0, i_8_345_781_0, i_8_345_795_0,
    i_8_345_813_0, i_8_345_826_0, i_8_345_843_0, i_8_345_879_0,
    i_8_345_940_0, i_8_345_969_0, i_8_345_985_0, i_8_345_1014_0,
    i_8_345_1032_0, i_8_345_1086_0, i_8_345_1115_0, i_8_345_1119_0,
    i_8_345_1132_0, i_8_345_1159_0, i_8_345_1218_0, i_8_345_1225_0,
    i_8_345_1248_0, i_8_345_1257_0, i_8_345_1284_0, i_8_345_1315_0,
    i_8_345_1327_0, i_8_345_1344_0, i_8_345_1389_0, i_8_345_1506_0,
    i_8_345_1524_0, i_8_345_1537_0, i_8_345_1542_0, i_8_345_1543_0,
    i_8_345_1545_0, i_8_345_1551_0, i_8_345_1590_0, i_8_345_1597_0,
    i_8_345_1606_0, i_8_345_1627_0, i_8_345_1632_0, i_8_345_1633_0,
    i_8_345_1680_0, i_8_345_1690_0, i_8_345_1698_0, i_8_345_1719_0,
    i_8_345_1722_0, i_8_345_1741_0, i_8_345_1752_0, i_8_345_1761_0,
    i_8_345_1803_0, i_8_345_1812_0, i_8_345_1813_0, i_8_345_1840_0,
    i_8_345_1841_0, i_8_345_1857_0, i_8_345_1866_0, i_8_345_1872_0,
    i_8_345_1875_0, i_8_345_1921_0, i_8_345_1950_0, i_8_345_2092_0,
    i_8_345_2110_0, i_8_345_2112_0, i_8_345_2113_0, i_8_345_2127_0,
    i_8_345_2131_0, i_8_345_2184_0, i_8_345_2185_0, i_8_345_2190_0,
    i_8_345_2214_0, i_8_345_2215_0, i_8_345_2289_0,
    o_8_345_0_0  );
  input  i_8_345_84_0, i_8_345_85_0, i_8_345_96_0, i_8_345_106_0,
    i_8_345_138_0, i_8_345_245_0, i_8_345_291_0, i_8_345_294_0,
    i_8_345_304_0, i_8_345_327_0, i_8_345_372_0, i_8_345_375_0,
    i_8_345_381_0, i_8_345_384_0, i_8_345_385_0, i_8_345_419_0,
    i_8_345_436_0, i_8_345_462_0, i_8_345_475_0, i_8_345_480_0,
    i_8_345_481_0, i_8_345_483_0, i_8_345_523_0, i_8_345_526_0,
    i_8_345_598_0, i_8_345_599_0, i_8_345_601_0, i_8_345_672_0,
    i_8_345_699_0, i_8_345_759_0, i_8_345_780_0, i_8_345_781_0,
    i_8_345_795_0, i_8_345_813_0, i_8_345_826_0, i_8_345_843_0,
    i_8_345_879_0, i_8_345_940_0, i_8_345_969_0, i_8_345_985_0,
    i_8_345_1014_0, i_8_345_1032_0, i_8_345_1086_0, i_8_345_1115_0,
    i_8_345_1119_0, i_8_345_1132_0, i_8_345_1159_0, i_8_345_1218_0,
    i_8_345_1225_0, i_8_345_1248_0, i_8_345_1257_0, i_8_345_1284_0,
    i_8_345_1315_0, i_8_345_1327_0, i_8_345_1344_0, i_8_345_1389_0,
    i_8_345_1506_0, i_8_345_1524_0, i_8_345_1537_0, i_8_345_1542_0,
    i_8_345_1543_0, i_8_345_1545_0, i_8_345_1551_0, i_8_345_1590_0,
    i_8_345_1597_0, i_8_345_1606_0, i_8_345_1627_0, i_8_345_1632_0,
    i_8_345_1633_0, i_8_345_1680_0, i_8_345_1690_0, i_8_345_1698_0,
    i_8_345_1719_0, i_8_345_1722_0, i_8_345_1741_0, i_8_345_1752_0,
    i_8_345_1761_0, i_8_345_1803_0, i_8_345_1812_0, i_8_345_1813_0,
    i_8_345_1840_0, i_8_345_1841_0, i_8_345_1857_0, i_8_345_1866_0,
    i_8_345_1872_0, i_8_345_1875_0, i_8_345_1921_0, i_8_345_1950_0,
    i_8_345_2092_0, i_8_345_2110_0, i_8_345_2112_0, i_8_345_2113_0,
    i_8_345_2127_0, i_8_345_2131_0, i_8_345_2184_0, i_8_345_2185_0,
    i_8_345_2190_0, i_8_345_2214_0, i_8_345_2215_0, i_8_345_2289_0;
  output o_8_345_0_0;
  assign o_8_345_0_0 = 0;
endmodule



// Benchmark "kernel_8_346" written by ABC on Sun Jul 19 10:09:05 2020

module kernel_8_346 ( 
    i_8_346_9_0, i_8_346_27_0, i_8_346_37_0, i_8_346_81_0, i_8_346_102_0,
    i_8_346_104_0, i_8_346_111_0, i_8_346_136_0, i_8_346_147_0,
    i_8_346_180_0, i_8_346_189_0, i_8_346_219_0, i_8_346_243_0,
    i_8_346_262_0, i_8_346_315_0, i_8_346_337_0, i_8_346_366_0,
    i_8_346_378_0, i_8_346_381_0, i_8_346_398_0, i_8_346_467_0,
    i_8_346_505_0, i_8_346_510_0, i_8_346_531_0, i_8_346_567_0,
    i_8_346_570_0, i_8_346_588_0, i_8_346_596_0, i_8_346_603_0,
    i_8_346_604_0, i_8_346_639_0, i_8_346_649_0, i_8_346_662_0,
    i_8_346_707_0, i_8_346_731_0, i_8_346_822_0, i_8_346_841_0,
    i_8_346_877_0, i_8_346_879_0, i_8_346_880_0, i_8_346_884_0,
    i_8_346_891_0, i_8_346_966_0, i_8_346_998_0, i_8_346_1008_0,
    i_8_346_1049_0, i_8_346_1098_0, i_8_346_1108_0, i_8_346_1109_0,
    i_8_346_1127_0, i_8_346_1140_0, i_8_346_1154_0, i_8_346_1171_0,
    i_8_346_1231_0, i_8_346_1233_0, i_8_346_1234_0, i_8_346_1276_0,
    i_8_346_1323_0, i_8_346_1324_0, i_8_346_1351_0, i_8_346_1354_0,
    i_8_346_1359_0, i_8_346_1404_0, i_8_346_1436_0, i_8_346_1457_0,
    i_8_346_1458_0, i_8_346_1476_0, i_8_346_1480_0, i_8_346_1491_0,
    i_8_346_1503_0, i_8_346_1522_0, i_8_346_1567_0, i_8_346_1602_0,
    i_8_346_1630_0, i_8_346_1683_0, i_8_346_1686_0, i_8_346_1696_0,
    i_8_346_1758_0, i_8_346_1764_0, i_8_346_1800_0, i_8_346_1810_0,
    i_8_346_1836_0, i_8_346_1837_0, i_8_346_1882_0, i_8_346_1890_0,
    i_8_346_1908_0, i_8_346_1936_0, i_8_346_1990_0, i_8_346_1992_0,
    i_8_346_2037_0, i_8_346_2066_0, i_8_346_2070_0, i_8_346_2071_0,
    i_8_346_2124_0, i_8_346_2145_0, i_8_346_2234_0, i_8_346_2244_0,
    i_8_346_2247_0, i_8_346_2269_0, i_8_346_2271_0,
    o_8_346_0_0  );
  input  i_8_346_9_0, i_8_346_27_0, i_8_346_37_0, i_8_346_81_0,
    i_8_346_102_0, i_8_346_104_0, i_8_346_111_0, i_8_346_136_0,
    i_8_346_147_0, i_8_346_180_0, i_8_346_189_0, i_8_346_219_0,
    i_8_346_243_0, i_8_346_262_0, i_8_346_315_0, i_8_346_337_0,
    i_8_346_366_0, i_8_346_378_0, i_8_346_381_0, i_8_346_398_0,
    i_8_346_467_0, i_8_346_505_0, i_8_346_510_0, i_8_346_531_0,
    i_8_346_567_0, i_8_346_570_0, i_8_346_588_0, i_8_346_596_0,
    i_8_346_603_0, i_8_346_604_0, i_8_346_639_0, i_8_346_649_0,
    i_8_346_662_0, i_8_346_707_0, i_8_346_731_0, i_8_346_822_0,
    i_8_346_841_0, i_8_346_877_0, i_8_346_879_0, i_8_346_880_0,
    i_8_346_884_0, i_8_346_891_0, i_8_346_966_0, i_8_346_998_0,
    i_8_346_1008_0, i_8_346_1049_0, i_8_346_1098_0, i_8_346_1108_0,
    i_8_346_1109_0, i_8_346_1127_0, i_8_346_1140_0, i_8_346_1154_0,
    i_8_346_1171_0, i_8_346_1231_0, i_8_346_1233_0, i_8_346_1234_0,
    i_8_346_1276_0, i_8_346_1323_0, i_8_346_1324_0, i_8_346_1351_0,
    i_8_346_1354_0, i_8_346_1359_0, i_8_346_1404_0, i_8_346_1436_0,
    i_8_346_1457_0, i_8_346_1458_0, i_8_346_1476_0, i_8_346_1480_0,
    i_8_346_1491_0, i_8_346_1503_0, i_8_346_1522_0, i_8_346_1567_0,
    i_8_346_1602_0, i_8_346_1630_0, i_8_346_1683_0, i_8_346_1686_0,
    i_8_346_1696_0, i_8_346_1758_0, i_8_346_1764_0, i_8_346_1800_0,
    i_8_346_1810_0, i_8_346_1836_0, i_8_346_1837_0, i_8_346_1882_0,
    i_8_346_1890_0, i_8_346_1908_0, i_8_346_1936_0, i_8_346_1990_0,
    i_8_346_1992_0, i_8_346_2037_0, i_8_346_2066_0, i_8_346_2070_0,
    i_8_346_2071_0, i_8_346_2124_0, i_8_346_2145_0, i_8_346_2234_0,
    i_8_346_2244_0, i_8_346_2247_0, i_8_346_2269_0, i_8_346_2271_0;
  output o_8_346_0_0;
  assign o_8_346_0_0 = ~((~i_8_346_136_0 & ((~i_8_346_567_0 & ~i_8_346_2070_0 & ~i_8_346_2247_0 & i_8_346_2271_0) | (~i_8_346_262_0 & i_8_346_1990_0 & ~i_8_346_2234_0 & ~i_8_346_2271_0))) | (~i_8_346_180_0 & ((~i_8_346_639_0 & i_8_346_1234_0 & i_8_346_1354_0) | (i_8_346_588_0 & ~i_8_346_1233_0 & ~i_8_346_1882_0))) | (~i_8_346_1458_0 & ((~i_8_346_262_0 & ((~i_8_346_315_0 & ~i_8_346_822_0 & ~i_8_346_1008_0 & ~i_8_346_2124_0) | (~i_8_346_1503_0 & ~i_8_346_1764_0 & ~i_8_346_1810_0 & ~i_8_346_2247_0))) | (~i_8_346_147_0 & ~i_8_346_315_0 & ~i_8_346_567_0 & ~i_8_346_1758_0 & ~i_8_346_2269_0))) | (~i_8_346_1683_0 & ((~i_8_346_315_0 & ((~i_8_346_567_0 & ~i_8_346_1359_0) | (~i_8_346_366_0 & ~i_8_346_1810_0 & ~i_8_346_1908_0))) | (~i_8_346_1049_0 & ~i_8_346_1098_0 & ~i_8_346_1837_0))) | (~i_8_346_1098_0 & ((~i_8_346_570_0 & ~i_8_346_604_0 & ~i_8_346_998_0 & ~i_8_346_1476_0) | (~i_8_346_1503_0 & ~i_8_346_1686_0 & ~i_8_346_1696_0))) | (~i_8_346_189_0 & ~i_8_346_510_0 & ~i_8_346_588_0 & ~i_8_346_603_0 & ~i_8_346_639_0) | (i_8_346_337_0 & ~i_8_346_1602_0 & ~i_8_346_1764_0 & ~i_8_346_1908_0));
endmodule



// Benchmark "kernel_8_347" written by ABC on Sun Jul 19 10:09:07 2020

module kernel_8_347 ( 
    i_8_347_79_0, i_8_347_84_0, i_8_347_85_0, i_8_347_88_0, i_8_347_168_0,
    i_8_347_193_0, i_8_347_224_0, i_8_347_295_0, i_8_347_303_0,
    i_8_347_323_0, i_8_347_364_0, i_8_347_499_0, i_8_347_500_0,
    i_8_347_525_0, i_8_347_526_0, i_8_347_527_0, i_8_347_528_0,
    i_8_347_529_0, i_8_347_530_0, i_8_347_591_0, i_8_347_592_0,
    i_8_347_593_0, i_8_347_606_0, i_8_347_629_0, i_8_347_634_0,
    i_8_347_660_0, i_8_347_665_0, i_8_347_670_0, i_8_347_678_0,
    i_8_347_679_0, i_8_347_682_0, i_8_347_683_0, i_8_347_707_0,
    i_8_347_708_0, i_8_347_763_0, i_8_347_807_0, i_8_347_813_0,
    i_8_347_842_0, i_8_347_964_0, i_8_347_1057_0, i_8_347_1058_0,
    i_8_347_1076_0, i_8_347_1192_0, i_8_347_1193_0, i_8_347_1266_0,
    i_8_347_1268_0, i_8_347_1272_0, i_8_347_1274_0, i_8_347_1299_0,
    i_8_347_1309_0, i_8_347_1339_0, i_8_347_1340_0, i_8_347_1353_0,
    i_8_347_1354_0, i_8_347_1390_0, i_8_347_1433_0, i_8_347_1437_0,
    i_8_347_1455_0, i_8_347_1485_0, i_8_347_1534_0, i_8_347_1536_0,
    i_8_347_1627_0, i_8_347_1632_0, i_8_347_1633_0, i_8_347_1634_0,
    i_8_347_1642_0, i_8_347_1732_0, i_8_347_1750_0, i_8_347_1752_0,
    i_8_347_1770_0, i_8_347_1771_0, i_8_347_1778_0, i_8_347_1783_0,
    i_8_347_1784_0, i_8_347_1785_0, i_8_347_1787_0, i_8_347_1789_0,
    i_8_347_1790_0, i_8_347_1822_0, i_8_347_1858_0, i_8_347_1859_0,
    i_8_347_1860_0, i_8_347_1861_0, i_8_347_1862_0, i_8_347_1866_0,
    i_8_347_1869_0, i_8_347_1905_0, i_8_347_1906_0, i_8_347_1975_0,
    i_8_347_1978_0, i_8_347_1996_0, i_8_347_2041_0, i_8_347_2136_0,
    i_8_347_2137_0, i_8_347_2214_0, i_8_347_2215_0, i_8_347_2226_0,
    i_8_347_2248_0, i_8_347_2249_0, i_8_347_2284_0,
    o_8_347_0_0  );
  input  i_8_347_79_0, i_8_347_84_0, i_8_347_85_0, i_8_347_88_0,
    i_8_347_168_0, i_8_347_193_0, i_8_347_224_0, i_8_347_295_0,
    i_8_347_303_0, i_8_347_323_0, i_8_347_364_0, i_8_347_499_0,
    i_8_347_500_0, i_8_347_525_0, i_8_347_526_0, i_8_347_527_0,
    i_8_347_528_0, i_8_347_529_0, i_8_347_530_0, i_8_347_591_0,
    i_8_347_592_0, i_8_347_593_0, i_8_347_606_0, i_8_347_629_0,
    i_8_347_634_0, i_8_347_660_0, i_8_347_665_0, i_8_347_670_0,
    i_8_347_678_0, i_8_347_679_0, i_8_347_682_0, i_8_347_683_0,
    i_8_347_707_0, i_8_347_708_0, i_8_347_763_0, i_8_347_807_0,
    i_8_347_813_0, i_8_347_842_0, i_8_347_964_0, i_8_347_1057_0,
    i_8_347_1058_0, i_8_347_1076_0, i_8_347_1192_0, i_8_347_1193_0,
    i_8_347_1266_0, i_8_347_1268_0, i_8_347_1272_0, i_8_347_1274_0,
    i_8_347_1299_0, i_8_347_1309_0, i_8_347_1339_0, i_8_347_1340_0,
    i_8_347_1353_0, i_8_347_1354_0, i_8_347_1390_0, i_8_347_1433_0,
    i_8_347_1437_0, i_8_347_1455_0, i_8_347_1485_0, i_8_347_1534_0,
    i_8_347_1536_0, i_8_347_1627_0, i_8_347_1632_0, i_8_347_1633_0,
    i_8_347_1634_0, i_8_347_1642_0, i_8_347_1732_0, i_8_347_1750_0,
    i_8_347_1752_0, i_8_347_1770_0, i_8_347_1771_0, i_8_347_1778_0,
    i_8_347_1783_0, i_8_347_1784_0, i_8_347_1785_0, i_8_347_1787_0,
    i_8_347_1789_0, i_8_347_1790_0, i_8_347_1822_0, i_8_347_1858_0,
    i_8_347_1859_0, i_8_347_1860_0, i_8_347_1861_0, i_8_347_1862_0,
    i_8_347_1866_0, i_8_347_1869_0, i_8_347_1905_0, i_8_347_1906_0,
    i_8_347_1975_0, i_8_347_1978_0, i_8_347_1996_0, i_8_347_2041_0,
    i_8_347_2136_0, i_8_347_2137_0, i_8_347_2214_0, i_8_347_2215_0,
    i_8_347_2226_0, i_8_347_2248_0, i_8_347_2249_0, i_8_347_2284_0;
  output o_8_347_0_0;
  assign o_8_347_0_0 = ~((~i_8_347_634_0 & ((~i_8_347_79_0 & ((i_8_347_84_0 & i_8_347_499_0) | (i_8_347_193_0 & ~i_8_347_364_0 & ~i_8_347_1266_0 & ~i_8_347_1268_0 & ~i_8_347_1771_0 & ~i_8_347_1783_0 & ~i_8_347_1785_0 & ~i_8_347_1861_0))) | (~i_8_347_364_0 & ((~i_8_347_303_0 & ~i_8_347_591_0 & ~i_8_347_606_0 & i_8_347_964_0 & ~i_8_347_1634_0) | (~i_8_347_499_0 & ~i_8_347_593_0 & ~i_8_347_1437_0 & ~i_8_347_1750_0 & ~i_8_347_1789_0 & ~i_8_347_1790_0 & i_8_347_1822_0 & ~i_8_347_2136_0))) | (~i_8_347_682_0 & ((i_8_347_84_0 & ~i_8_347_1309_0 & ~i_8_347_1339_0 & i_8_347_2136_0) | (~i_8_347_591_0 & i_8_347_670_0 & ~i_8_347_842_0 & ~i_8_347_1272_0 & ~i_8_347_1485_0 & ~i_8_347_2136_0))) | (~i_8_347_707_0 & ((~i_8_347_593_0 & ~i_8_347_606_0 & ~i_8_347_660_0 & ~i_8_347_1785_0 & i_8_347_1858_0 & ~i_8_347_2137_0) | (~i_8_347_683_0 & ~i_8_347_1266_0 & ~i_8_347_1268_0 & ~i_8_347_1309_0 & ~i_8_347_1433_0 & ~i_8_347_1750_0 & ~i_8_347_1752_0 & ~i_8_347_1783_0 & ~i_8_347_1789_0 & ~i_8_347_1790_0 & ~i_8_347_1822_0 & ~i_8_347_1858_0 & ~i_8_347_2136_0 & ~i_8_347_2249_0))) | (~i_8_347_593_0 & ((i_8_347_964_0 & ~i_8_347_1771_0 & ~i_8_347_1862_0 & i_8_347_2215_0) | (i_8_347_500_0 & ~i_8_347_1274_0 & ~i_8_347_1354_0 & ~i_8_347_1632_0 & ~i_8_347_1822_0 & ~i_8_347_1996_0 & ~i_8_347_2136_0 & ~i_8_347_2226_0))) | (~i_8_347_660_0 & ((~i_8_347_193_0 & ~i_8_347_500_0 & ~i_8_347_665_0 & ~i_8_347_679_0 & i_8_347_842_0 & ~i_8_347_1193_0 & ~i_8_347_1309_0 & ~i_8_347_1340_0 & ~i_8_347_1433_0 & ~i_8_347_1750_0 & i_8_347_1778_0) | (~i_8_347_1299_0 & ~i_8_347_1485_0 & i_8_347_1534_0 & i_8_347_1750_0 & ~i_8_347_1778_0))) | (i_8_347_1353_0 & ((~i_8_347_592_0 & ~i_8_347_678_0 & ~i_8_347_1437_0 & ~i_8_347_1783_0 & ~i_8_347_1787_0 & ~i_8_347_1822_0 & ~i_8_347_1996_0 & ~i_8_347_2214_0) | (i_8_347_364_0 & ~i_8_347_1057_0 & i_8_347_1354_0 & ~i_8_347_1632_0 & ~i_8_347_1634_0 & ~i_8_347_2215_0))) | (~i_8_347_592_0 & ((i_8_347_1455_0 & ~i_8_347_1485_0 & ~i_8_347_1634_0 & ~i_8_347_1752_0) | (~i_8_347_1787_0 & i_8_347_1858_0 & ~i_8_347_2136_0 & i_8_347_2137_0 & ~i_8_347_2215_0))) | (i_8_347_526_0 & ~i_8_347_708_0 & ~i_8_347_842_0 & ~i_8_347_1770_0 & ~i_8_347_1784_0 & ~i_8_347_1822_0 & ~i_8_347_1858_0 & ~i_8_347_2249_0))) | (~i_8_347_85_0 & ((~i_8_347_707_0 & ~i_8_347_842_0 & ~i_8_347_1309_0 & i_8_347_1433_0 & ~i_8_347_1485_0 & i_8_347_1534_0 & ~i_8_347_1866_0 & ~i_8_347_1996_0) | (i_8_347_1272_0 & ~i_8_347_1534_0 & ~i_8_347_1632_0 & ~i_8_347_1633_0 & ~i_8_347_1787_0 & ~i_8_347_1822_0 & ~i_8_347_2248_0))) | (~i_8_347_1778_0 & ((~i_8_347_224_0 & ((~i_8_347_303_0 & i_8_347_526_0 & ~i_8_347_660_0 & ~i_8_347_1785_0) | (i_8_347_85_0 & ~i_8_347_528_0 & ~i_8_347_1455_0 & ~i_8_347_1783_0 & ~i_8_347_1859_0 & ~i_8_347_2137_0))) | (~i_8_347_660_0 & ~i_8_347_1787_0 & ((i_8_347_1057_0 & ~i_8_347_1266_0 & ~i_8_347_1822_0 & ~i_8_347_2214_0) | (~i_8_347_606_0 & ~i_8_347_665_0 & ~i_8_347_1353_0 & ~i_8_347_1354_0 & ~i_8_347_1433_0 & ~i_8_347_1485_0 & ~i_8_347_1534_0 & ~i_8_347_1771_0 & ~i_8_347_1785_0 & ~i_8_347_1789_0 & ~i_8_347_2136_0 & ~i_8_347_2137_0 & ~i_8_347_2226_0))) | (~i_8_347_1783_0 & ~i_8_347_1822_0 & ((i_8_347_964_0 & ~i_8_347_1771_0) | (~i_8_347_665_0 & ~i_8_347_678_0 & ~i_8_347_1268_0 & ~i_8_347_1309_0 & i_8_347_1354_0 & ~i_8_347_2226_0 & ~i_8_347_2249_0))) | (~i_8_347_303_0 & ~i_8_347_1339_0 & ~i_8_347_1632_0 & i_8_347_1732_0))) | (~i_8_347_1770_0 & ((i_8_347_85_0 & ((~i_8_347_323_0 & i_8_347_526_0 & ~i_8_347_660_0 & ~i_8_347_1905_0 & ~i_8_347_1996_0 & ~i_8_347_2226_0) | (i_8_347_364_0 & ~i_8_347_1642_0 & ~i_8_347_1906_0 & ~i_8_347_2249_0))) | (~i_8_347_1785_0 & ((~i_8_347_224_0 & i_8_347_526_0 & ~i_8_347_1076_0 & ~i_8_347_1783_0) | (~i_8_347_678_0 & ~i_8_347_1634_0 & i_8_347_2284_0))) | (~i_8_347_1268_0 & i_8_347_1783_0 & ~i_8_347_1784_0 & ~i_8_347_1789_0 & i_8_347_1862_0) | (~i_8_347_591_0 & ~i_8_347_679_0 & ~i_8_347_1433_0 & ~i_8_347_1771_0 & i_8_347_1860_0 & ~i_8_347_2248_0))) | (~i_8_347_1433_0 & ((~i_8_347_323_0 & ~i_8_347_1437_0 & ((i_8_347_530_0 & ~i_8_347_683_0 & ~i_8_347_1634_0) | (i_8_347_1058_0 & ~i_8_347_1353_0 & ~i_8_347_1752_0 & ~i_8_347_1783_0))) | (i_8_347_525_0 & ~i_8_347_682_0 & ~i_8_347_1353_0 & ~i_8_347_1455_0 & ~i_8_347_1536_0 & ~i_8_347_1627_0 & i_8_347_1790_0) | (~i_8_347_1193_0 & ~i_8_347_1485_0 & ~i_8_347_1783_0 & ~i_8_347_1787_0 & i_8_347_1861_0 & i_8_347_1862_0) | (~i_8_347_79_0 & ~i_8_347_683_0 & ~i_8_347_1340_0 & ~i_8_347_1785_0 & i_8_347_1859_0 & ~i_8_347_2137_0))) | (i_8_347_526_0 & ((i_8_347_499_0 & i_8_347_525_0 & ~i_8_347_682_0) | (~i_8_347_660_0 & ~i_8_347_683_0 & i_8_347_1193_0 & ~i_8_347_1536_0))) | (~i_8_347_2249_0 & ((~i_8_347_1783_0 & ((~i_8_347_79_0 & ~i_8_347_1299_0 & ~i_8_347_2137_0 & ((~i_8_347_593_0 & ~i_8_347_683_0 & i_8_347_842_0 & ~i_8_347_1340_0 & ~i_8_347_1485_0 & ~i_8_347_1642_0 & ~i_8_347_1750_0 & ~i_8_347_1784_0) | (~i_8_347_592_0 & ~i_8_347_1858_0 & i_8_347_1861_0 & ~i_8_347_2226_0 & ~i_8_347_2248_0))) | (~i_8_347_364_0 & ~i_8_347_606_0 & ~i_8_347_1354_0 & ~i_8_347_1784_0 & i_8_347_1858_0 & ~i_8_347_2136_0 & ~i_8_347_2214_0))) | (i_8_347_525_0 & ~i_8_347_1784_0 & ((~i_8_347_679_0 & i_8_347_1272_0) | (~i_8_347_606_0 & ~i_8_347_1787_0 & i_8_347_1822_0))) | (i_8_347_1076_0 & ((~i_8_347_364_0 & ~i_8_347_660_0 & i_8_347_1778_0 & ~i_8_347_1785_0 & i_8_347_1859_0) | (~i_8_347_1309_0 & ~i_8_347_1822_0 & ~i_8_347_1996_0 & ~i_8_347_2136_0))) | (i_8_347_88_0 & i_8_347_529_0 & ~i_8_347_606_0 & ~i_8_347_683_0))) | (~i_8_347_678_0 & ((~i_8_347_527_0 & ((~i_8_347_364_0 & i_8_347_634_0 & ~i_8_347_660_0 & ~i_8_347_679_0 & i_8_347_964_0 & ~i_8_347_1057_0 & i_8_347_1783_0 & i_8_347_1858_0) | (~i_8_347_295_0 & ~i_8_347_500_0 & ~i_8_347_526_0 & ~i_8_347_665_0 & ~i_8_347_682_0 & ~i_8_347_683_0 & ~i_8_347_807_0 & ~i_8_347_1274_0 & i_8_347_1536_0 & ~i_8_347_1634_0 & i_8_347_1860_0 & ~i_8_347_2136_0))) | (i_8_347_528_0 & ~i_8_347_682_0 & ~i_8_347_683_0 & ~i_8_347_707_0 & ~i_8_347_964_0 & ~i_8_347_1266_0 & ~i_8_347_1632_0 & ~i_8_347_1732_0) | (~i_8_347_606_0 & i_8_347_707_0 & ~i_8_347_842_0 & ~i_8_347_1354_0 & ~i_8_347_1634_0 & i_8_347_1750_0 & i_8_347_1787_0 & ~i_8_347_1996_0))) | (~i_8_347_500_0 & ((~i_8_347_679_0 & ~i_8_347_683_0 & i_8_347_1274_0 & ~i_8_347_1634_0 & ~i_8_347_1783_0) | (~i_8_347_224_0 & ~i_8_347_592_0 & ~i_8_347_660_0 & ~i_8_347_1266_0 & ~i_8_347_1339_0 & ~i_8_347_1455_0 & i_8_347_1642_0 & ~i_8_347_2136_0))) | (~i_8_347_660_0 & ((~i_8_347_1353_0 & ~i_8_347_1783_0 & ~i_8_347_2136_0 & i_8_347_2214_0 & ~i_8_347_2215_0) | (i_8_347_193_0 & i_8_347_1272_0 & ~i_8_347_2248_0))) | (~i_8_347_707_0 & ((~i_8_347_708_0 & ~i_8_347_1299_0 & i_8_347_1353_0 & i_8_347_1354_0 & ~i_8_347_1752_0 & ~i_8_347_1783_0 & ~i_8_347_1784_0) | (i_8_347_1534_0 & ~i_8_347_2136_0 & ~i_8_347_2137_0 & i_8_347_2214_0))) | (i_8_347_1192_0 & ((~i_8_347_88_0 & i_8_347_364_0 & ~i_8_347_964_0 & ~i_8_347_1634_0 & ~i_8_347_1869_0 & ~i_8_347_2136_0) | (i_8_347_1354_0 & ~i_8_347_1771_0 & ~i_8_347_2214_0))) | (~i_8_347_1299_0 & ((~i_8_347_629_0 & i_8_347_1274_0 & ~i_8_347_1534_0 & ~i_8_347_1789_0 & i_8_347_1859_0) | (~i_8_347_193_0 & ~i_8_347_683_0 & ~i_8_347_1632_0 & ~i_8_347_1783_0 & ~i_8_347_1784_0 & ~i_8_347_1785_0 & i_8_347_1860_0))) | (i_8_347_1354_0 & ((i_8_347_527_0 & ~i_8_347_842_0 & ~i_8_347_1268_0) | (~i_8_347_79_0 & i_8_347_500_0 & ~i_8_347_1632_0 & ~i_8_347_1750_0 & ~i_8_347_1790_0))) | (~i_8_347_1783_0 & ((i_8_347_530_0 & ~i_8_347_592_0 & ~i_8_347_1274_0 & ~i_8_347_1340_0) | (~i_8_347_679_0 & i_8_347_1309_0 & i_8_347_1536_0))) | (~i_8_347_1785_0 & ((i_8_347_1058_0 & i_8_347_1193_0) | (~i_8_347_665_0 & i_8_347_1770_0 & ~i_8_347_1784_0 & ~i_8_347_1789_0 & ~i_8_347_2136_0 & ~i_8_347_2248_0))));
endmodule



// Benchmark "kernel_8_348" written by ABC on Sun Jul 19 10:09:07 2020

module kernel_8_348 ( 
    i_8_348_32_0, i_8_348_58_0, i_8_348_84_0, i_8_348_85_0, i_8_348_92_0,
    i_8_348_94_0, i_8_348_101_0, i_8_348_103_0, i_8_348_140_0,
    i_8_348_155_0, i_8_348_185_0, i_8_348_299_0, i_8_348_372_0,
    i_8_348_373_0, i_8_348_380_0, i_8_348_419_0, i_8_348_437_0,
    i_8_348_441_0, i_8_348_460_0, i_8_348_461_0, i_8_348_482_0,
    i_8_348_522_0, i_8_348_529_0, i_8_348_572_0, i_8_348_587_0,
    i_8_348_613_0, i_8_348_622_0, i_8_348_623_0, i_8_348_667_0,
    i_8_348_668_0, i_8_348_697_0, i_8_348_713_0, i_8_348_715_0,
    i_8_348_716_0, i_8_348_722_0, i_8_348_731_0, i_8_348_756_0,
    i_8_348_757_0, i_8_348_767_0, i_8_348_779_0, i_8_348_793_0,
    i_8_348_821_0, i_8_348_842_0, i_8_348_866_0, i_8_348_1010_0,
    i_8_348_1028_0, i_8_348_1043_0, i_8_348_1135_0, i_8_348_1153_0,
    i_8_348_1154_0, i_8_348_1157_0, i_8_348_1253_0, i_8_348_1279_0,
    i_8_348_1280_0, i_8_348_1305_0, i_8_348_1306_0, i_8_348_1313_0,
    i_8_348_1323_0, i_8_348_1342_0, i_8_348_1343_0, i_8_348_1435_0,
    i_8_348_1436_0, i_8_348_1452_0, i_8_348_1504_0, i_8_348_1505_0,
    i_8_348_1542_0, i_8_348_1550_0, i_8_348_1562_0, i_8_348_1603_0,
    i_8_348_1613_0, i_8_348_1630_0, i_8_348_1676_0, i_8_348_1697_0,
    i_8_348_1711_0, i_8_348_1748_0, i_8_348_1749_0, i_8_348_1759_0,
    i_8_348_1802_0, i_8_348_1818_0, i_8_348_1856_0, i_8_348_1886_0,
    i_8_348_1892_0, i_8_348_1964_0, i_8_348_1973_0, i_8_348_1985_0,
    i_8_348_1994_0, i_8_348_2036_0, i_8_348_2075_0, i_8_348_2108_0,
    i_8_348_2134_0, i_8_348_2141_0, i_8_348_2143_0, i_8_348_2144_0,
    i_8_348_2145_0, i_8_348_2153_0, i_8_348_2171_0, i_8_348_2188_0,
    i_8_348_2246_0, i_8_348_2272_0, i_8_348_2288_0,
    o_8_348_0_0  );
  input  i_8_348_32_0, i_8_348_58_0, i_8_348_84_0, i_8_348_85_0,
    i_8_348_92_0, i_8_348_94_0, i_8_348_101_0, i_8_348_103_0,
    i_8_348_140_0, i_8_348_155_0, i_8_348_185_0, i_8_348_299_0,
    i_8_348_372_0, i_8_348_373_0, i_8_348_380_0, i_8_348_419_0,
    i_8_348_437_0, i_8_348_441_0, i_8_348_460_0, i_8_348_461_0,
    i_8_348_482_0, i_8_348_522_0, i_8_348_529_0, i_8_348_572_0,
    i_8_348_587_0, i_8_348_613_0, i_8_348_622_0, i_8_348_623_0,
    i_8_348_667_0, i_8_348_668_0, i_8_348_697_0, i_8_348_713_0,
    i_8_348_715_0, i_8_348_716_0, i_8_348_722_0, i_8_348_731_0,
    i_8_348_756_0, i_8_348_757_0, i_8_348_767_0, i_8_348_779_0,
    i_8_348_793_0, i_8_348_821_0, i_8_348_842_0, i_8_348_866_0,
    i_8_348_1010_0, i_8_348_1028_0, i_8_348_1043_0, i_8_348_1135_0,
    i_8_348_1153_0, i_8_348_1154_0, i_8_348_1157_0, i_8_348_1253_0,
    i_8_348_1279_0, i_8_348_1280_0, i_8_348_1305_0, i_8_348_1306_0,
    i_8_348_1313_0, i_8_348_1323_0, i_8_348_1342_0, i_8_348_1343_0,
    i_8_348_1435_0, i_8_348_1436_0, i_8_348_1452_0, i_8_348_1504_0,
    i_8_348_1505_0, i_8_348_1542_0, i_8_348_1550_0, i_8_348_1562_0,
    i_8_348_1603_0, i_8_348_1613_0, i_8_348_1630_0, i_8_348_1676_0,
    i_8_348_1697_0, i_8_348_1711_0, i_8_348_1748_0, i_8_348_1749_0,
    i_8_348_1759_0, i_8_348_1802_0, i_8_348_1818_0, i_8_348_1856_0,
    i_8_348_1886_0, i_8_348_1892_0, i_8_348_1964_0, i_8_348_1973_0,
    i_8_348_1985_0, i_8_348_1994_0, i_8_348_2036_0, i_8_348_2075_0,
    i_8_348_2108_0, i_8_348_2134_0, i_8_348_2141_0, i_8_348_2143_0,
    i_8_348_2144_0, i_8_348_2145_0, i_8_348_2153_0, i_8_348_2171_0,
    i_8_348_2188_0, i_8_348_2246_0, i_8_348_2272_0, i_8_348_2288_0;
  output o_8_348_0_0;
  assign o_8_348_0_0 = 0;
endmodule



// Benchmark "kernel_8_349" written by ABC on Sun Jul 19 10:09:08 2020

module kernel_8_349 ( 
    i_8_349_6_0, i_8_349_24_0, i_8_349_25_0, i_8_349_78_0, i_8_349_115_0,
    i_8_349_177_0, i_8_349_249_0, i_8_349_250_0, i_8_349_265_0,
    i_8_349_349_0, i_8_349_355_0, i_8_349_357_0, i_8_349_373_0,
    i_8_349_384_0, i_8_349_385_0, i_8_349_395_0, i_8_349_445_0,
    i_8_349_465_0, i_8_349_475_0, i_8_349_481_0, i_8_349_493_0,
    i_8_349_501_0, i_8_349_520_0, i_8_349_522_0, i_8_349_556_0,
    i_8_349_580_0, i_8_349_673_0, i_8_349_710_0, i_8_349_762_0,
    i_8_349_770_0, i_8_349_771_0, i_8_349_807_0, i_8_349_842_0,
    i_8_349_850_0, i_8_349_856_0, i_8_349_861_0, i_8_349_889_0,
    i_8_349_944_0, i_8_349_967_0, i_8_349_968_0, i_8_349_1057_0,
    i_8_349_1059_0, i_8_349_1060_0, i_8_349_1087_0, i_8_349_1194_0,
    i_8_349_1227_0, i_8_349_1230_0, i_8_349_1239_0, i_8_349_1266_0,
    i_8_349_1272_0, i_8_349_1275_0, i_8_349_1276_0, i_8_349_1285_0,
    i_8_349_1299_0, i_8_349_1307_0, i_8_349_1317_0, i_8_349_1393_0,
    i_8_349_1399_0, i_8_349_1402_0, i_8_349_1404_0, i_8_349_1419_0,
    i_8_349_1432_0, i_8_349_1472_0, i_8_349_1473_0, i_8_349_1536_0,
    i_8_349_1538_0, i_8_349_1553_0, i_8_349_1632_0, i_8_349_1636_0,
    i_8_349_1654_0, i_8_349_1663_0, i_8_349_1699_0, i_8_349_1704_0,
    i_8_349_1716_0, i_8_349_1749_0, i_8_349_1808_0, i_8_349_1860_0,
    i_8_349_1862_0, i_8_349_1868_0, i_8_349_1879_0, i_8_349_1885_0,
    i_8_349_1888_0, i_8_349_1921_0, i_8_349_1929_0, i_8_349_1960_0,
    i_8_349_1969_0, i_8_349_1975_0, i_8_349_1995_0, i_8_349_2047_0,
    i_8_349_2058_0, i_8_349_2059_0, i_8_349_2068_0, i_8_349_2073_0,
    i_8_349_2076_0, i_8_349_2145_0, i_8_349_2158_0, i_8_349_2176_0,
    i_8_349_2219_0, i_8_349_2299_0, i_8_349_2302_0,
    o_8_349_0_0  );
  input  i_8_349_6_0, i_8_349_24_0, i_8_349_25_0, i_8_349_78_0,
    i_8_349_115_0, i_8_349_177_0, i_8_349_249_0, i_8_349_250_0,
    i_8_349_265_0, i_8_349_349_0, i_8_349_355_0, i_8_349_357_0,
    i_8_349_373_0, i_8_349_384_0, i_8_349_385_0, i_8_349_395_0,
    i_8_349_445_0, i_8_349_465_0, i_8_349_475_0, i_8_349_481_0,
    i_8_349_493_0, i_8_349_501_0, i_8_349_520_0, i_8_349_522_0,
    i_8_349_556_0, i_8_349_580_0, i_8_349_673_0, i_8_349_710_0,
    i_8_349_762_0, i_8_349_770_0, i_8_349_771_0, i_8_349_807_0,
    i_8_349_842_0, i_8_349_850_0, i_8_349_856_0, i_8_349_861_0,
    i_8_349_889_0, i_8_349_944_0, i_8_349_967_0, i_8_349_968_0,
    i_8_349_1057_0, i_8_349_1059_0, i_8_349_1060_0, i_8_349_1087_0,
    i_8_349_1194_0, i_8_349_1227_0, i_8_349_1230_0, i_8_349_1239_0,
    i_8_349_1266_0, i_8_349_1272_0, i_8_349_1275_0, i_8_349_1276_0,
    i_8_349_1285_0, i_8_349_1299_0, i_8_349_1307_0, i_8_349_1317_0,
    i_8_349_1393_0, i_8_349_1399_0, i_8_349_1402_0, i_8_349_1404_0,
    i_8_349_1419_0, i_8_349_1432_0, i_8_349_1472_0, i_8_349_1473_0,
    i_8_349_1536_0, i_8_349_1538_0, i_8_349_1553_0, i_8_349_1632_0,
    i_8_349_1636_0, i_8_349_1654_0, i_8_349_1663_0, i_8_349_1699_0,
    i_8_349_1704_0, i_8_349_1716_0, i_8_349_1749_0, i_8_349_1808_0,
    i_8_349_1860_0, i_8_349_1862_0, i_8_349_1868_0, i_8_349_1879_0,
    i_8_349_1885_0, i_8_349_1888_0, i_8_349_1921_0, i_8_349_1929_0,
    i_8_349_1960_0, i_8_349_1969_0, i_8_349_1975_0, i_8_349_1995_0,
    i_8_349_2047_0, i_8_349_2058_0, i_8_349_2059_0, i_8_349_2068_0,
    i_8_349_2073_0, i_8_349_2076_0, i_8_349_2145_0, i_8_349_2158_0,
    i_8_349_2176_0, i_8_349_2219_0, i_8_349_2299_0, i_8_349_2302_0;
  output o_8_349_0_0;
  assign o_8_349_0_0 = 0;
endmodule



// Benchmark "kernel_8_350" written by ABC on Sun Jul 19 10:09:09 2020

module kernel_8_350 ( 
    i_8_350_10_0, i_8_350_13_0, i_8_350_38_0, i_8_350_40_0, i_8_350_41_0,
    i_8_350_47_0, i_8_350_50_0, i_8_350_73_0, i_8_350_91_0, i_8_350_136_0,
    i_8_350_143_0, i_8_350_182_0, i_8_350_193_0, i_8_350_239_0,
    i_8_350_254_0, i_8_350_334_0, i_8_350_344_0, i_8_350_362_0,
    i_8_350_364_0, i_8_350_397_0, i_8_350_398_0, i_8_350_423_0,
    i_8_350_425_0, i_8_350_427_0, i_8_350_428_0, i_8_350_451_0,
    i_8_350_452_0, i_8_350_490_0, i_8_350_491_0, i_8_350_532_0,
    i_8_350_533_0, i_8_350_578_0, i_8_350_595_0, i_8_350_608_0,
    i_8_350_612_0, i_8_350_613_0, i_8_350_640_0, i_8_350_641_0,
    i_8_350_675_0, i_8_350_676_0, i_8_350_677_0, i_8_350_694_0,
    i_8_350_695_0, i_8_350_699_0, i_8_350_700_0, i_8_350_748_0,
    i_8_350_775_0, i_8_350_782_0, i_8_350_796_0, i_8_350_839_0,
    i_8_350_844_0, i_8_350_856_0, i_8_350_857_0, i_8_350_858_0,
    i_8_350_878_0, i_8_350_973_0, i_8_350_1034_0, i_8_350_1036_0,
    i_8_350_1057_0, i_8_350_1154_0, i_8_350_1156_0, i_8_350_1226_0,
    i_8_350_1235_0, i_8_350_1236_0, i_8_350_1243_0, i_8_350_1292_0,
    i_8_350_1314_0, i_8_350_1315_0, i_8_350_1325_0, i_8_350_1411_0,
    i_8_350_1468_0, i_8_350_1489_0, i_8_350_1490_0, i_8_350_1564_0,
    i_8_350_1624_0, i_8_350_1632_0, i_8_350_1669_0, i_8_350_1694_0,
    i_8_350_1764_0, i_8_350_1765_0, i_8_350_1767_0, i_8_350_1783_0,
    i_8_350_1786_0, i_8_350_1818_0, i_8_350_1819_0, i_8_350_1830_0,
    i_8_350_1837_0, i_8_350_1885_0, i_8_350_1940_0, i_8_350_1969_0,
    i_8_350_2110_0, i_8_350_2111_0, i_8_350_2133_0, i_8_350_2147_0,
    i_8_350_2148_0, i_8_350_2152_0, i_8_350_2165_0, i_8_350_2225_0,
    i_8_350_2236_0, i_8_350_2263_0,
    o_8_350_0_0  );
  input  i_8_350_10_0, i_8_350_13_0, i_8_350_38_0, i_8_350_40_0,
    i_8_350_41_0, i_8_350_47_0, i_8_350_50_0, i_8_350_73_0, i_8_350_91_0,
    i_8_350_136_0, i_8_350_143_0, i_8_350_182_0, i_8_350_193_0,
    i_8_350_239_0, i_8_350_254_0, i_8_350_334_0, i_8_350_344_0,
    i_8_350_362_0, i_8_350_364_0, i_8_350_397_0, i_8_350_398_0,
    i_8_350_423_0, i_8_350_425_0, i_8_350_427_0, i_8_350_428_0,
    i_8_350_451_0, i_8_350_452_0, i_8_350_490_0, i_8_350_491_0,
    i_8_350_532_0, i_8_350_533_0, i_8_350_578_0, i_8_350_595_0,
    i_8_350_608_0, i_8_350_612_0, i_8_350_613_0, i_8_350_640_0,
    i_8_350_641_0, i_8_350_675_0, i_8_350_676_0, i_8_350_677_0,
    i_8_350_694_0, i_8_350_695_0, i_8_350_699_0, i_8_350_700_0,
    i_8_350_748_0, i_8_350_775_0, i_8_350_782_0, i_8_350_796_0,
    i_8_350_839_0, i_8_350_844_0, i_8_350_856_0, i_8_350_857_0,
    i_8_350_858_0, i_8_350_878_0, i_8_350_973_0, i_8_350_1034_0,
    i_8_350_1036_0, i_8_350_1057_0, i_8_350_1154_0, i_8_350_1156_0,
    i_8_350_1226_0, i_8_350_1235_0, i_8_350_1236_0, i_8_350_1243_0,
    i_8_350_1292_0, i_8_350_1314_0, i_8_350_1315_0, i_8_350_1325_0,
    i_8_350_1411_0, i_8_350_1468_0, i_8_350_1489_0, i_8_350_1490_0,
    i_8_350_1564_0, i_8_350_1624_0, i_8_350_1632_0, i_8_350_1669_0,
    i_8_350_1694_0, i_8_350_1764_0, i_8_350_1765_0, i_8_350_1767_0,
    i_8_350_1783_0, i_8_350_1786_0, i_8_350_1818_0, i_8_350_1819_0,
    i_8_350_1830_0, i_8_350_1837_0, i_8_350_1885_0, i_8_350_1940_0,
    i_8_350_1969_0, i_8_350_2110_0, i_8_350_2111_0, i_8_350_2133_0,
    i_8_350_2147_0, i_8_350_2148_0, i_8_350_2152_0, i_8_350_2165_0,
    i_8_350_2225_0, i_8_350_2236_0, i_8_350_2263_0;
  output o_8_350_0_0;
  assign o_8_350_0_0 = 0;
endmodule



// Benchmark "kernel_8_351" written by ABC on Sun Jul 19 10:09:10 2020

module kernel_8_351 ( 
    i_8_351_22_0, i_8_351_29_0, i_8_351_34_0, i_8_351_56_0, i_8_351_57_0,
    i_8_351_73_0, i_8_351_95_0, i_8_351_136_0, i_8_351_184_0,
    i_8_351_231_0, i_8_351_253_0, i_8_351_254_0, i_8_351_259_0,
    i_8_351_305_0, i_8_351_365_0, i_8_351_378_0, i_8_351_398_0,
    i_8_351_424_0, i_8_351_454_0, i_8_351_469_0, i_8_351_505_0,
    i_8_351_506_0, i_8_351_554_0, i_8_351_581_0, i_8_351_586_0,
    i_8_351_609_0, i_8_351_622_0, i_8_351_637_0, i_8_351_639_0,
    i_8_351_678_0, i_8_351_680_0, i_8_351_704_0, i_8_351_706_0,
    i_8_351_709_0, i_8_351_710_0, i_8_351_730_0, i_8_351_751_0,
    i_8_351_778_0, i_8_351_785_0, i_8_351_839_0, i_8_351_856_0,
    i_8_351_866_0, i_8_351_875_0, i_8_351_965_0, i_8_351_1063_0,
    i_8_351_1064_0, i_8_351_1099_0, i_8_351_1102_0, i_8_351_1103_0,
    i_8_351_1130_0, i_8_351_1145_0, i_8_351_1265_0, i_8_351_1283_0,
    i_8_351_1297_0, i_8_351_1298_0, i_8_351_1299_0, i_8_351_1355_0,
    i_8_351_1360_0, i_8_351_1366_0, i_8_351_1385_0, i_8_351_1393_0,
    i_8_351_1397_0, i_8_351_1402_0, i_8_351_1431_0, i_8_351_1434_0,
    i_8_351_1462_0, i_8_351_1463_0, i_8_351_1471_0, i_8_351_1548_0,
    i_8_351_1559_0, i_8_351_1632_0, i_8_351_1633_0, i_8_351_1688_0,
    i_8_351_1705_0, i_8_351_1786_0, i_8_351_1789_0, i_8_351_1795_0,
    i_8_351_1812_0, i_8_351_1821_0, i_8_351_1886_0, i_8_351_1888_0,
    i_8_351_1889_0, i_8_351_1891_0, i_8_351_1940_0, i_8_351_1963_0,
    i_8_351_1989_0, i_8_351_2056_0, i_8_351_2101_0, i_8_351_2107_0,
    i_8_351_2131_0, i_8_351_2132_0, i_8_351_2153_0, i_8_351_2170_0,
    i_8_351_2225_0, i_8_351_2234_0, i_8_351_2244_0, i_8_351_2246_0,
    i_8_351_2261_0, i_8_351_2263_0, i_8_351_2264_0,
    o_8_351_0_0  );
  input  i_8_351_22_0, i_8_351_29_0, i_8_351_34_0, i_8_351_56_0,
    i_8_351_57_0, i_8_351_73_0, i_8_351_95_0, i_8_351_136_0, i_8_351_184_0,
    i_8_351_231_0, i_8_351_253_0, i_8_351_254_0, i_8_351_259_0,
    i_8_351_305_0, i_8_351_365_0, i_8_351_378_0, i_8_351_398_0,
    i_8_351_424_0, i_8_351_454_0, i_8_351_469_0, i_8_351_505_0,
    i_8_351_506_0, i_8_351_554_0, i_8_351_581_0, i_8_351_586_0,
    i_8_351_609_0, i_8_351_622_0, i_8_351_637_0, i_8_351_639_0,
    i_8_351_678_0, i_8_351_680_0, i_8_351_704_0, i_8_351_706_0,
    i_8_351_709_0, i_8_351_710_0, i_8_351_730_0, i_8_351_751_0,
    i_8_351_778_0, i_8_351_785_0, i_8_351_839_0, i_8_351_856_0,
    i_8_351_866_0, i_8_351_875_0, i_8_351_965_0, i_8_351_1063_0,
    i_8_351_1064_0, i_8_351_1099_0, i_8_351_1102_0, i_8_351_1103_0,
    i_8_351_1130_0, i_8_351_1145_0, i_8_351_1265_0, i_8_351_1283_0,
    i_8_351_1297_0, i_8_351_1298_0, i_8_351_1299_0, i_8_351_1355_0,
    i_8_351_1360_0, i_8_351_1366_0, i_8_351_1385_0, i_8_351_1393_0,
    i_8_351_1397_0, i_8_351_1402_0, i_8_351_1431_0, i_8_351_1434_0,
    i_8_351_1462_0, i_8_351_1463_0, i_8_351_1471_0, i_8_351_1548_0,
    i_8_351_1559_0, i_8_351_1632_0, i_8_351_1633_0, i_8_351_1688_0,
    i_8_351_1705_0, i_8_351_1786_0, i_8_351_1789_0, i_8_351_1795_0,
    i_8_351_1812_0, i_8_351_1821_0, i_8_351_1886_0, i_8_351_1888_0,
    i_8_351_1889_0, i_8_351_1891_0, i_8_351_1940_0, i_8_351_1963_0,
    i_8_351_1989_0, i_8_351_2056_0, i_8_351_2101_0, i_8_351_2107_0,
    i_8_351_2131_0, i_8_351_2132_0, i_8_351_2153_0, i_8_351_2170_0,
    i_8_351_2225_0, i_8_351_2234_0, i_8_351_2244_0, i_8_351_2246_0,
    i_8_351_2261_0, i_8_351_2263_0, i_8_351_2264_0;
  output o_8_351_0_0;
  assign o_8_351_0_0 = 0;
endmodule



// Benchmark "kernel_8_352" written by ABC on Sun Jul 19 10:09:11 2020

module kernel_8_352 ( 
    i_8_352_18_0, i_8_352_21_0, i_8_352_33_0, i_8_352_34_0, i_8_352_52_0,
    i_8_352_105_0, i_8_352_114_0, i_8_352_173_0, i_8_352_203_0,
    i_8_352_223_0, i_8_352_300_0, i_8_352_307_0, i_8_352_319_0,
    i_8_352_356_0, i_8_352_372_0, i_8_352_374_0, i_8_352_381_0,
    i_8_352_391_0, i_8_352_392_0, i_8_352_497_0, i_8_352_518_0,
    i_8_352_594_0, i_8_352_597_0, i_8_352_600_0, i_8_352_604_0,
    i_8_352_608_0, i_8_352_610_0, i_8_352_640_0, i_8_352_657_0,
    i_8_352_661_0, i_8_352_668_0, i_8_352_675_0, i_8_352_678_0,
    i_8_352_681_0, i_8_352_748_0, i_8_352_776_0, i_8_352_850_0,
    i_8_352_860_0, i_8_352_867_0, i_8_352_870_0, i_8_352_871_0,
    i_8_352_878_0, i_8_352_896_0, i_8_352_974_0, i_8_352_986_0,
    i_8_352_1037_0, i_8_352_1085_0, i_8_352_1101_0, i_8_352_1102_0,
    i_8_352_1125_0, i_8_352_1126_0, i_8_352_1136_0, i_8_352_1140_0,
    i_8_352_1218_0, i_8_352_1228_0, i_8_352_1317_0, i_8_352_1362_0,
    i_8_352_1382_0, i_8_352_1443_0, i_8_352_1459_0, i_8_352_1462_0,
    i_8_352_1470_0, i_8_352_1499_0, i_8_352_1514_0, i_8_352_1517_0,
    i_8_352_1533_0, i_8_352_1557_0, i_8_352_1596_0, i_8_352_1605_0,
    i_8_352_1680_0, i_8_352_1688_0, i_8_352_1701_0, i_8_352_1702_0,
    i_8_352_1713_0, i_8_352_1733_0, i_8_352_1747_0, i_8_352_1748_0,
    i_8_352_1761_0, i_8_352_1762_0, i_8_352_1776_0, i_8_352_1782_0,
    i_8_352_1783_0, i_8_352_1810_0, i_8_352_1812_0, i_8_352_1817_0,
    i_8_352_1821_0, i_8_352_1890_0, i_8_352_1891_0, i_8_352_1903_0,
    i_8_352_1910_0, i_8_352_1947_0, i_8_352_1981_0, i_8_352_2056_0,
    i_8_352_2107_0, i_8_352_2129_0, i_8_352_2154_0, i_8_352_2201_0,
    i_8_352_2235_0, i_8_352_2241_0, i_8_352_2262_0,
    o_8_352_0_0  );
  input  i_8_352_18_0, i_8_352_21_0, i_8_352_33_0, i_8_352_34_0,
    i_8_352_52_0, i_8_352_105_0, i_8_352_114_0, i_8_352_173_0,
    i_8_352_203_0, i_8_352_223_0, i_8_352_300_0, i_8_352_307_0,
    i_8_352_319_0, i_8_352_356_0, i_8_352_372_0, i_8_352_374_0,
    i_8_352_381_0, i_8_352_391_0, i_8_352_392_0, i_8_352_497_0,
    i_8_352_518_0, i_8_352_594_0, i_8_352_597_0, i_8_352_600_0,
    i_8_352_604_0, i_8_352_608_0, i_8_352_610_0, i_8_352_640_0,
    i_8_352_657_0, i_8_352_661_0, i_8_352_668_0, i_8_352_675_0,
    i_8_352_678_0, i_8_352_681_0, i_8_352_748_0, i_8_352_776_0,
    i_8_352_850_0, i_8_352_860_0, i_8_352_867_0, i_8_352_870_0,
    i_8_352_871_0, i_8_352_878_0, i_8_352_896_0, i_8_352_974_0,
    i_8_352_986_0, i_8_352_1037_0, i_8_352_1085_0, i_8_352_1101_0,
    i_8_352_1102_0, i_8_352_1125_0, i_8_352_1126_0, i_8_352_1136_0,
    i_8_352_1140_0, i_8_352_1218_0, i_8_352_1228_0, i_8_352_1317_0,
    i_8_352_1362_0, i_8_352_1382_0, i_8_352_1443_0, i_8_352_1459_0,
    i_8_352_1462_0, i_8_352_1470_0, i_8_352_1499_0, i_8_352_1514_0,
    i_8_352_1517_0, i_8_352_1533_0, i_8_352_1557_0, i_8_352_1596_0,
    i_8_352_1605_0, i_8_352_1680_0, i_8_352_1688_0, i_8_352_1701_0,
    i_8_352_1702_0, i_8_352_1713_0, i_8_352_1733_0, i_8_352_1747_0,
    i_8_352_1748_0, i_8_352_1761_0, i_8_352_1762_0, i_8_352_1776_0,
    i_8_352_1782_0, i_8_352_1783_0, i_8_352_1810_0, i_8_352_1812_0,
    i_8_352_1817_0, i_8_352_1821_0, i_8_352_1890_0, i_8_352_1891_0,
    i_8_352_1903_0, i_8_352_1910_0, i_8_352_1947_0, i_8_352_1981_0,
    i_8_352_2056_0, i_8_352_2107_0, i_8_352_2129_0, i_8_352_2154_0,
    i_8_352_2201_0, i_8_352_2235_0, i_8_352_2241_0, i_8_352_2262_0;
  output o_8_352_0_0;
  assign o_8_352_0_0 = 0;
endmodule



// Benchmark "kernel_8_353" written by ABC on Sun Jul 19 10:09:12 2020

module kernel_8_353 ( 
    i_8_353_17_0, i_8_353_40_0, i_8_353_45_0, i_8_353_65_0, i_8_353_68_0,
    i_8_353_142_0, i_8_353_184_0, i_8_353_187_0, i_8_353_205_0,
    i_8_353_222_0, i_8_353_228_0, i_8_353_237_0, i_8_353_243_0,
    i_8_353_252_0, i_8_353_281_0, i_8_353_298_0, i_8_353_322_0,
    i_8_353_335_0, i_8_353_360_0, i_8_353_382_0, i_8_353_417_0,
    i_8_353_426_0, i_8_353_451_0, i_8_353_471_0, i_8_353_505_0,
    i_8_353_514_0, i_8_353_549_0, i_8_353_556_0, i_8_353_583_0,
    i_8_353_584_0, i_8_353_637_0, i_8_353_655_0, i_8_353_681_0,
    i_8_353_738_0, i_8_353_749_0, i_8_353_763_0, i_8_353_770_0,
    i_8_353_778_0, i_8_353_796_0, i_8_353_797_0, i_8_353_840_0,
    i_8_353_842_0, i_8_353_917_0, i_8_353_940_0, i_8_353_941_0,
    i_8_353_1053_0, i_8_353_1112_0, i_8_353_1137_0, i_8_353_1147_0,
    i_8_353_1155_0, i_8_353_1227_0, i_8_353_1234_0, i_8_353_1245_0,
    i_8_353_1246_0, i_8_353_1256_0, i_8_353_1280_0, i_8_353_1285_0,
    i_8_353_1286_0, i_8_353_1288_0, i_8_353_1296_0, i_8_353_1331_0,
    i_8_353_1332_0, i_8_353_1335_0, i_8_353_1336_0, i_8_353_1365_0,
    i_8_353_1367_0, i_8_353_1384_0, i_8_353_1400_0, i_8_353_1440_0,
    i_8_353_1464_0, i_8_353_1467_0, i_8_353_1528_0, i_8_353_1556_0,
    i_8_353_1606_0, i_8_353_1678_0, i_8_353_1689_0, i_8_353_1696_0,
    i_8_353_1702_0, i_8_353_1706_0, i_8_353_1714_0, i_8_353_1722_0,
    i_8_353_1745_0, i_8_353_1753_0, i_8_353_1754_0, i_8_353_1784_0,
    i_8_353_1787_0, i_8_353_1822_0, i_8_353_1883_0, i_8_353_1902_0,
    i_8_353_1963_0, i_8_353_1975_0, i_8_353_1996_0, i_8_353_2001_0,
    i_8_353_2073_0, i_8_353_2097_0, i_8_353_2106_0, i_8_353_2170_0,
    i_8_353_2224_0, i_8_353_2259_0, i_8_353_2280_0,
    o_8_353_0_0  );
  input  i_8_353_17_0, i_8_353_40_0, i_8_353_45_0, i_8_353_65_0,
    i_8_353_68_0, i_8_353_142_0, i_8_353_184_0, i_8_353_187_0,
    i_8_353_205_0, i_8_353_222_0, i_8_353_228_0, i_8_353_237_0,
    i_8_353_243_0, i_8_353_252_0, i_8_353_281_0, i_8_353_298_0,
    i_8_353_322_0, i_8_353_335_0, i_8_353_360_0, i_8_353_382_0,
    i_8_353_417_0, i_8_353_426_0, i_8_353_451_0, i_8_353_471_0,
    i_8_353_505_0, i_8_353_514_0, i_8_353_549_0, i_8_353_556_0,
    i_8_353_583_0, i_8_353_584_0, i_8_353_637_0, i_8_353_655_0,
    i_8_353_681_0, i_8_353_738_0, i_8_353_749_0, i_8_353_763_0,
    i_8_353_770_0, i_8_353_778_0, i_8_353_796_0, i_8_353_797_0,
    i_8_353_840_0, i_8_353_842_0, i_8_353_917_0, i_8_353_940_0,
    i_8_353_941_0, i_8_353_1053_0, i_8_353_1112_0, i_8_353_1137_0,
    i_8_353_1147_0, i_8_353_1155_0, i_8_353_1227_0, i_8_353_1234_0,
    i_8_353_1245_0, i_8_353_1246_0, i_8_353_1256_0, i_8_353_1280_0,
    i_8_353_1285_0, i_8_353_1286_0, i_8_353_1288_0, i_8_353_1296_0,
    i_8_353_1331_0, i_8_353_1332_0, i_8_353_1335_0, i_8_353_1336_0,
    i_8_353_1365_0, i_8_353_1367_0, i_8_353_1384_0, i_8_353_1400_0,
    i_8_353_1440_0, i_8_353_1464_0, i_8_353_1467_0, i_8_353_1528_0,
    i_8_353_1556_0, i_8_353_1606_0, i_8_353_1678_0, i_8_353_1689_0,
    i_8_353_1696_0, i_8_353_1702_0, i_8_353_1706_0, i_8_353_1714_0,
    i_8_353_1722_0, i_8_353_1745_0, i_8_353_1753_0, i_8_353_1754_0,
    i_8_353_1784_0, i_8_353_1787_0, i_8_353_1822_0, i_8_353_1883_0,
    i_8_353_1902_0, i_8_353_1963_0, i_8_353_1975_0, i_8_353_1996_0,
    i_8_353_2001_0, i_8_353_2073_0, i_8_353_2097_0, i_8_353_2106_0,
    i_8_353_2170_0, i_8_353_2224_0, i_8_353_2259_0, i_8_353_2280_0;
  output o_8_353_0_0;
  assign o_8_353_0_0 = 0;
endmodule



// Benchmark "kernel_8_354" written by ABC on Sun Jul 19 10:09:13 2020

module kernel_8_354 ( 
    i_8_354_16_0, i_8_354_34_0, i_8_354_185_0, i_8_354_257_0,
    i_8_354_281_0, i_8_354_283_0, i_8_354_338_0, i_8_354_383_0,
    i_8_354_391_0, i_8_354_392_0, i_8_354_400_0, i_8_354_418_0,
    i_8_354_450_0, i_8_354_451_0, i_8_354_509_0, i_8_354_554_0,
    i_8_354_557_0, i_8_354_563_0, i_8_354_569_0, i_8_354_583_0,
    i_8_354_633_0, i_8_354_644_0, i_8_354_652_0, i_8_354_653_0,
    i_8_354_663_0, i_8_354_700_0, i_8_354_703_0, i_8_354_704_0,
    i_8_354_751_0, i_8_354_769_0, i_8_354_782_0, i_8_354_785_0,
    i_8_354_823_0, i_8_354_827_0, i_8_354_842_0, i_8_354_866_0,
    i_8_354_874_0, i_8_354_895_0, i_8_354_958_0, i_8_354_969_0,
    i_8_354_1012_0, i_8_354_1013_0, i_8_354_1036_0, i_8_354_1109_0,
    i_8_354_1129_0, i_8_354_1132_0, i_8_354_1201_0, i_8_354_1285_0,
    i_8_354_1300_0, i_8_354_1303_0, i_8_354_1328_0, i_8_354_1357_0,
    i_8_354_1382_0, i_8_354_1411_0, i_8_354_1435_0, i_8_354_1436_0,
    i_8_354_1452_0, i_8_354_1468_0, i_8_354_1477_0, i_8_354_1478_0,
    i_8_354_1489_0, i_8_354_1511_0, i_8_354_1525_0, i_8_354_1526_0,
    i_8_354_1547_0, i_8_354_1553_0, i_8_354_1571_0, i_8_354_1603_0,
    i_8_354_1679_0, i_8_354_1696_0, i_8_354_1705_0, i_8_354_1706_0,
    i_8_354_1723_0, i_8_354_1750_0, i_8_354_1784_0, i_8_354_1794_0,
    i_8_354_1796_0, i_8_354_1807_0, i_8_354_1821_0, i_8_354_1822_0,
    i_8_354_1824_0, i_8_354_1840_0, i_8_354_1841_0, i_8_354_1868_0,
    i_8_354_1886_0, i_8_354_1894_0, i_8_354_1895_0, i_8_354_1912_0,
    i_8_354_1939_0, i_8_354_1976_0, i_8_354_1982_0, i_8_354_2074_0,
    i_8_354_2075_0, i_8_354_2154_0, i_8_354_2159_0, i_8_354_2182_0,
    i_8_354_2224_0, i_8_354_2227_0, i_8_354_2248_0, i_8_354_2276_0,
    o_8_354_0_0  );
  input  i_8_354_16_0, i_8_354_34_0, i_8_354_185_0, i_8_354_257_0,
    i_8_354_281_0, i_8_354_283_0, i_8_354_338_0, i_8_354_383_0,
    i_8_354_391_0, i_8_354_392_0, i_8_354_400_0, i_8_354_418_0,
    i_8_354_450_0, i_8_354_451_0, i_8_354_509_0, i_8_354_554_0,
    i_8_354_557_0, i_8_354_563_0, i_8_354_569_0, i_8_354_583_0,
    i_8_354_633_0, i_8_354_644_0, i_8_354_652_0, i_8_354_653_0,
    i_8_354_663_0, i_8_354_700_0, i_8_354_703_0, i_8_354_704_0,
    i_8_354_751_0, i_8_354_769_0, i_8_354_782_0, i_8_354_785_0,
    i_8_354_823_0, i_8_354_827_0, i_8_354_842_0, i_8_354_866_0,
    i_8_354_874_0, i_8_354_895_0, i_8_354_958_0, i_8_354_969_0,
    i_8_354_1012_0, i_8_354_1013_0, i_8_354_1036_0, i_8_354_1109_0,
    i_8_354_1129_0, i_8_354_1132_0, i_8_354_1201_0, i_8_354_1285_0,
    i_8_354_1300_0, i_8_354_1303_0, i_8_354_1328_0, i_8_354_1357_0,
    i_8_354_1382_0, i_8_354_1411_0, i_8_354_1435_0, i_8_354_1436_0,
    i_8_354_1452_0, i_8_354_1468_0, i_8_354_1477_0, i_8_354_1478_0,
    i_8_354_1489_0, i_8_354_1511_0, i_8_354_1525_0, i_8_354_1526_0,
    i_8_354_1547_0, i_8_354_1553_0, i_8_354_1571_0, i_8_354_1603_0,
    i_8_354_1679_0, i_8_354_1696_0, i_8_354_1705_0, i_8_354_1706_0,
    i_8_354_1723_0, i_8_354_1750_0, i_8_354_1784_0, i_8_354_1794_0,
    i_8_354_1796_0, i_8_354_1807_0, i_8_354_1821_0, i_8_354_1822_0,
    i_8_354_1824_0, i_8_354_1840_0, i_8_354_1841_0, i_8_354_1868_0,
    i_8_354_1886_0, i_8_354_1894_0, i_8_354_1895_0, i_8_354_1912_0,
    i_8_354_1939_0, i_8_354_1976_0, i_8_354_1982_0, i_8_354_2074_0,
    i_8_354_2075_0, i_8_354_2154_0, i_8_354_2159_0, i_8_354_2182_0,
    i_8_354_2224_0, i_8_354_2227_0, i_8_354_2248_0, i_8_354_2276_0;
  output o_8_354_0_0;
  assign o_8_354_0_0 = 0;
endmodule



// Benchmark "kernel_8_355" written by ABC on Sun Jul 19 10:09:14 2020

module kernel_8_355 ( 
    i_8_355_50_0, i_8_355_59_0, i_8_355_76_0, i_8_355_85_0, i_8_355_104_0,
    i_8_355_107_0, i_8_355_118_0, i_8_355_218_0, i_8_355_304_0,
    i_8_355_322_0, i_8_355_362_0, i_8_355_367_0, i_8_355_368_0,
    i_8_355_374_0, i_8_355_385_0, i_8_355_414_0, i_8_355_453_0,
    i_8_355_488_0, i_8_355_524_0, i_8_355_530_0, i_8_355_547_0,
    i_8_355_556_0, i_8_355_557_0, i_8_355_608_0, i_8_355_611_0,
    i_8_355_616_0, i_8_355_633_0, i_8_355_634_0, i_8_355_652_0,
    i_8_355_655_0, i_8_355_656_0, i_8_355_657_0, i_8_355_661_0,
    i_8_355_662_0, i_8_355_665_0, i_8_355_697_0, i_8_355_700_0,
    i_8_355_707_0, i_8_355_760_0, i_8_355_769_0, i_8_355_772_0,
    i_8_355_827_0, i_8_355_844_0, i_8_355_869_0, i_8_355_877_0,
    i_8_355_886_0, i_8_355_943_0, i_8_355_956_0, i_8_355_958_0,
    i_8_355_959_0, i_8_355_965_0, i_8_355_970_0, i_8_355_977_0,
    i_8_355_991_0, i_8_355_1039_0, i_8_355_1115_0, i_8_355_1138_0,
    i_8_355_1256_0, i_8_355_1267_0, i_8_355_1268_0, i_8_355_1319_0,
    i_8_355_1348_0, i_8_355_1439_0, i_8_355_1453_0, i_8_355_1474_0,
    i_8_355_1489_0, i_8_355_1516_0, i_8_355_1525_0, i_8_355_1544_0,
    i_8_355_1546_0, i_8_355_1555_0, i_8_355_1562_0, i_8_355_1673_0,
    i_8_355_1732_0, i_8_355_1765_0, i_8_355_1787_0, i_8_355_1795_0,
    i_8_355_1813_0, i_8_355_1822_0, i_8_355_1859_0, i_8_355_1877_0,
    i_8_355_1887_0, i_8_355_1909_0, i_8_355_1915_0, i_8_355_1993_0,
    i_8_355_1996_0, i_8_355_2056_0, i_8_355_2090_0, i_8_355_2092_0,
    i_8_355_2093_0, i_8_355_2102_0, i_8_355_2125_0, i_8_355_2129_0,
    i_8_355_2135_0, i_8_355_2149_0, i_8_355_2156_0, i_8_355_2173_0,
    i_8_355_2227_0, i_8_355_2233_0, i_8_355_2245_0,
    o_8_355_0_0  );
  input  i_8_355_50_0, i_8_355_59_0, i_8_355_76_0, i_8_355_85_0,
    i_8_355_104_0, i_8_355_107_0, i_8_355_118_0, i_8_355_218_0,
    i_8_355_304_0, i_8_355_322_0, i_8_355_362_0, i_8_355_367_0,
    i_8_355_368_0, i_8_355_374_0, i_8_355_385_0, i_8_355_414_0,
    i_8_355_453_0, i_8_355_488_0, i_8_355_524_0, i_8_355_530_0,
    i_8_355_547_0, i_8_355_556_0, i_8_355_557_0, i_8_355_608_0,
    i_8_355_611_0, i_8_355_616_0, i_8_355_633_0, i_8_355_634_0,
    i_8_355_652_0, i_8_355_655_0, i_8_355_656_0, i_8_355_657_0,
    i_8_355_661_0, i_8_355_662_0, i_8_355_665_0, i_8_355_697_0,
    i_8_355_700_0, i_8_355_707_0, i_8_355_760_0, i_8_355_769_0,
    i_8_355_772_0, i_8_355_827_0, i_8_355_844_0, i_8_355_869_0,
    i_8_355_877_0, i_8_355_886_0, i_8_355_943_0, i_8_355_956_0,
    i_8_355_958_0, i_8_355_959_0, i_8_355_965_0, i_8_355_970_0,
    i_8_355_977_0, i_8_355_991_0, i_8_355_1039_0, i_8_355_1115_0,
    i_8_355_1138_0, i_8_355_1256_0, i_8_355_1267_0, i_8_355_1268_0,
    i_8_355_1319_0, i_8_355_1348_0, i_8_355_1439_0, i_8_355_1453_0,
    i_8_355_1474_0, i_8_355_1489_0, i_8_355_1516_0, i_8_355_1525_0,
    i_8_355_1544_0, i_8_355_1546_0, i_8_355_1555_0, i_8_355_1562_0,
    i_8_355_1673_0, i_8_355_1732_0, i_8_355_1765_0, i_8_355_1787_0,
    i_8_355_1795_0, i_8_355_1813_0, i_8_355_1822_0, i_8_355_1859_0,
    i_8_355_1877_0, i_8_355_1887_0, i_8_355_1909_0, i_8_355_1915_0,
    i_8_355_1993_0, i_8_355_1996_0, i_8_355_2056_0, i_8_355_2090_0,
    i_8_355_2092_0, i_8_355_2093_0, i_8_355_2102_0, i_8_355_2125_0,
    i_8_355_2129_0, i_8_355_2135_0, i_8_355_2149_0, i_8_355_2156_0,
    i_8_355_2173_0, i_8_355_2227_0, i_8_355_2233_0, i_8_355_2245_0;
  output o_8_355_0_0;
  assign o_8_355_0_0 = 0;
endmodule



// Benchmark "kernel_8_356" written by ABC on Sun Jul 19 10:09:15 2020

module kernel_8_356 ( 
    i_8_356_39_0, i_8_356_88_0, i_8_356_136_0, i_8_356_159_0,
    i_8_356_183_0, i_8_356_187_0, i_8_356_265_0, i_8_356_285_0,
    i_8_356_295_0, i_8_356_300_0, i_8_356_322_0, i_8_356_331_0,
    i_8_356_363_0, i_8_356_364_0, i_8_356_368_0, i_8_356_393_0,
    i_8_356_399_0, i_8_356_420_0, i_8_356_426_0, i_8_356_459_0,
    i_8_356_510_0, i_8_356_565_0, i_8_356_591_0, i_8_356_592_0,
    i_8_356_594_0, i_8_356_598_0, i_8_356_608_0, i_8_356_612_0,
    i_8_356_660_0, i_8_356_673_0, i_8_356_681_0, i_8_356_683_0,
    i_8_356_703_0, i_8_356_707_0, i_8_356_736_0, i_8_356_750_0,
    i_8_356_809_0, i_8_356_826_0, i_8_356_832_0, i_8_356_835_0,
    i_8_356_838_0, i_8_356_841_0, i_8_356_843_0, i_8_356_850_0,
    i_8_356_927_0, i_8_356_1024_0, i_8_356_1050_0, i_8_356_1052_0,
    i_8_356_1055_0, i_8_356_1060_0, i_8_356_1132_0, i_8_356_1165_0,
    i_8_356_1200_0, i_8_356_1229_0, i_8_356_1231_0, i_8_356_1236_0,
    i_8_356_1240_0, i_8_356_1326_0, i_8_356_1375_0, i_8_356_1376_0,
    i_8_356_1381_0, i_8_356_1384_0, i_8_356_1402_0, i_8_356_1426_0,
    i_8_356_1456_0, i_8_356_1510_0, i_8_356_1524_0, i_8_356_1549_0,
    i_8_356_1552_0, i_8_356_1600_0, i_8_356_1635_0, i_8_356_1680_0,
    i_8_356_1686_0, i_8_356_1687_0, i_8_356_1704_0, i_8_356_1705_0,
    i_8_356_1796_0, i_8_356_1798_0, i_8_356_1819_0, i_8_356_1842_0,
    i_8_356_1884_0, i_8_356_1938_0, i_8_356_1939_0, i_8_356_1978_0,
    i_8_356_2048_0, i_8_356_2113_0, i_8_356_2121_0, i_8_356_2122_0,
    i_8_356_2131_0, i_8_356_2132_0, i_8_356_2140_0, i_8_356_2145_0,
    i_8_356_2147_0, i_8_356_2153_0, i_8_356_2172_0, i_8_356_2173_0,
    i_8_356_2224_0, i_8_356_2247_0, i_8_356_2256_0, i_8_356_2293_0,
    o_8_356_0_0  );
  input  i_8_356_39_0, i_8_356_88_0, i_8_356_136_0, i_8_356_159_0,
    i_8_356_183_0, i_8_356_187_0, i_8_356_265_0, i_8_356_285_0,
    i_8_356_295_0, i_8_356_300_0, i_8_356_322_0, i_8_356_331_0,
    i_8_356_363_0, i_8_356_364_0, i_8_356_368_0, i_8_356_393_0,
    i_8_356_399_0, i_8_356_420_0, i_8_356_426_0, i_8_356_459_0,
    i_8_356_510_0, i_8_356_565_0, i_8_356_591_0, i_8_356_592_0,
    i_8_356_594_0, i_8_356_598_0, i_8_356_608_0, i_8_356_612_0,
    i_8_356_660_0, i_8_356_673_0, i_8_356_681_0, i_8_356_683_0,
    i_8_356_703_0, i_8_356_707_0, i_8_356_736_0, i_8_356_750_0,
    i_8_356_809_0, i_8_356_826_0, i_8_356_832_0, i_8_356_835_0,
    i_8_356_838_0, i_8_356_841_0, i_8_356_843_0, i_8_356_850_0,
    i_8_356_927_0, i_8_356_1024_0, i_8_356_1050_0, i_8_356_1052_0,
    i_8_356_1055_0, i_8_356_1060_0, i_8_356_1132_0, i_8_356_1165_0,
    i_8_356_1200_0, i_8_356_1229_0, i_8_356_1231_0, i_8_356_1236_0,
    i_8_356_1240_0, i_8_356_1326_0, i_8_356_1375_0, i_8_356_1376_0,
    i_8_356_1381_0, i_8_356_1384_0, i_8_356_1402_0, i_8_356_1426_0,
    i_8_356_1456_0, i_8_356_1510_0, i_8_356_1524_0, i_8_356_1549_0,
    i_8_356_1552_0, i_8_356_1600_0, i_8_356_1635_0, i_8_356_1680_0,
    i_8_356_1686_0, i_8_356_1687_0, i_8_356_1704_0, i_8_356_1705_0,
    i_8_356_1796_0, i_8_356_1798_0, i_8_356_1819_0, i_8_356_1842_0,
    i_8_356_1884_0, i_8_356_1938_0, i_8_356_1939_0, i_8_356_1978_0,
    i_8_356_2048_0, i_8_356_2113_0, i_8_356_2121_0, i_8_356_2122_0,
    i_8_356_2131_0, i_8_356_2132_0, i_8_356_2140_0, i_8_356_2145_0,
    i_8_356_2147_0, i_8_356_2153_0, i_8_356_2172_0, i_8_356_2173_0,
    i_8_356_2224_0, i_8_356_2247_0, i_8_356_2256_0, i_8_356_2293_0;
  output o_8_356_0_0;
  assign o_8_356_0_0 = 0;
endmodule



// Benchmark "kernel_8_357" written by ABC on Sun Jul 19 10:09:16 2020

module kernel_8_357 ( 
    i_8_357_30_0, i_8_357_112_0, i_8_357_119_0, i_8_357_194_0,
    i_8_357_220_0, i_8_357_223_0, i_8_357_289_0, i_8_357_298_0,
    i_8_357_317_0, i_8_357_343_0, i_8_357_344_0, i_8_357_380_0,
    i_8_357_382_0, i_8_357_431_0, i_8_357_442_0, i_8_357_451_0,
    i_8_357_453_0, i_8_357_463_0, i_8_357_496_0, i_8_357_498_0,
    i_8_357_529_0, i_8_357_549_0, i_8_357_605_0, i_8_357_610_0,
    i_8_357_611_0, i_8_357_622_0, i_8_357_668_0, i_8_357_686_0,
    i_8_357_697_0, i_8_357_704_0, i_8_357_707_0, i_8_357_711_0,
    i_8_357_752_0, i_8_357_765_0, i_8_357_792_0, i_8_357_794_0,
    i_8_357_820_0, i_8_357_823_0, i_8_357_837_0, i_8_357_840_0,
    i_8_357_875_0, i_8_357_991_0, i_8_357_1004_0, i_8_357_1045_0,
    i_8_357_1046_0, i_8_357_1077_0, i_8_357_1103_0, i_8_357_1107_0,
    i_8_357_1111_0, i_8_357_1117_0, i_8_357_1139_0, i_8_357_1253_0,
    i_8_357_1271_0, i_8_357_1297_0, i_8_357_1324_0, i_8_357_1335_0,
    i_8_357_1355_0, i_8_357_1449_0, i_8_357_1451_0, i_8_357_1468_0,
    i_8_357_1478_0, i_8_357_1507_0, i_8_357_1536_0, i_8_357_1537_0,
    i_8_357_1541_0, i_8_357_1544_0, i_8_357_1549_0, i_8_357_1550_0,
    i_8_357_1594_0, i_8_357_1602_0, i_8_357_1620_0, i_8_357_1643_0,
    i_8_357_1649_0, i_8_357_1674_0, i_8_357_1749_0, i_8_357_1751_0,
    i_8_357_1801_0, i_8_357_1821_0, i_8_357_1856_0, i_8_357_1859_0,
    i_8_357_1863_0, i_8_357_1891_0, i_8_357_1901_0, i_8_357_1927_0,
    i_8_357_1962_0, i_8_357_2072_0, i_8_357_2089_0, i_8_357_2090_0,
    i_8_357_2107_0, i_8_357_2124_0, i_8_357_2125_0, i_8_357_2126_0,
    i_8_357_2132_0, i_8_357_2146_0, i_8_357_2242_0, i_8_357_2254_0,
    i_8_357_2268_0, i_8_357_2269_0, i_8_357_2270_0, i_8_357_2287_0,
    o_8_357_0_0  );
  input  i_8_357_30_0, i_8_357_112_0, i_8_357_119_0, i_8_357_194_0,
    i_8_357_220_0, i_8_357_223_0, i_8_357_289_0, i_8_357_298_0,
    i_8_357_317_0, i_8_357_343_0, i_8_357_344_0, i_8_357_380_0,
    i_8_357_382_0, i_8_357_431_0, i_8_357_442_0, i_8_357_451_0,
    i_8_357_453_0, i_8_357_463_0, i_8_357_496_0, i_8_357_498_0,
    i_8_357_529_0, i_8_357_549_0, i_8_357_605_0, i_8_357_610_0,
    i_8_357_611_0, i_8_357_622_0, i_8_357_668_0, i_8_357_686_0,
    i_8_357_697_0, i_8_357_704_0, i_8_357_707_0, i_8_357_711_0,
    i_8_357_752_0, i_8_357_765_0, i_8_357_792_0, i_8_357_794_0,
    i_8_357_820_0, i_8_357_823_0, i_8_357_837_0, i_8_357_840_0,
    i_8_357_875_0, i_8_357_991_0, i_8_357_1004_0, i_8_357_1045_0,
    i_8_357_1046_0, i_8_357_1077_0, i_8_357_1103_0, i_8_357_1107_0,
    i_8_357_1111_0, i_8_357_1117_0, i_8_357_1139_0, i_8_357_1253_0,
    i_8_357_1271_0, i_8_357_1297_0, i_8_357_1324_0, i_8_357_1335_0,
    i_8_357_1355_0, i_8_357_1449_0, i_8_357_1451_0, i_8_357_1468_0,
    i_8_357_1478_0, i_8_357_1507_0, i_8_357_1536_0, i_8_357_1537_0,
    i_8_357_1541_0, i_8_357_1544_0, i_8_357_1549_0, i_8_357_1550_0,
    i_8_357_1594_0, i_8_357_1602_0, i_8_357_1620_0, i_8_357_1643_0,
    i_8_357_1649_0, i_8_357_1674_0, i_8_357_1749_0, i_8_357_1751_0,
    i_8_357_1801_0, i_8_357_1821_0, i_8_357_1856_0, i_8_357_1859_0,
    i_8_357_1863_0, i_8_357_1891_0, i_8_357_1901_0, i_8_357_1927_0,
    i_8_357_1962_0, i_8_357_2072_0, i_8_357_2089_0, i_8_357_2090_0,
    i_8_357_2107_0, i_8_357_2124_0, i_8_357_2125_0, i_8_357_2126_0,
    i_8_357_2132_0, i_8_357_2146_0, i_8_357_2242_0, i_8_357_2254_0,
    i_8_357_2268_0, i_8_357_2269_0, i_8_357_2270_0, i_8_357_2287_0;
  output o_8_357_0_0;
  assign o_8_357_0_0 = 0;
endmodule



// Benchmark "kernel_8_358" written by ABC on Sun Jul 19 10:09:17 2020

module kernel_8_358 ( 
    i_8_358_104_0, i_8_358_153_0, i_8_358_154_0, i_8_358_155_0,
    i_8_358_158_0, i_8_358_160_0, i_8_358_205_0, i_8_358_206_0,
    i_8_358_221_0, i_8_358_435_0, i_8_358_471_0, i_8_358_480_0,
    i_8_358_489_0, i_8_358_499_0, i_8_358_500_0, i_8_358_572_0,
    i_8_358_592_0, i_8_358_606_0, i_8_358_610_0, i_8_358_624_0,
    i_8_358_684_0, i_8_358_688_0, i_8_358_699_0, i_8_358_714_0,
    i_8_358_716_0, i_8_358_717_0, i_8_358_729_0, i_8_358_778_0,
    i_8_358_779_0, i_8_358_780_0, i_8_358_782_0, i_8_358_787_0,
    i_8_358_837_0, i_8_358_838_0, i_8_358_867_0, i_8_358_869_0,
    i_8_358_871_0, i_8_358_879_0, i_8_358_881_0, i_8_358_998_0,
    i_8_358_1008_0, i_8_358_1012_0, i_8_358_1026_0, i_8_358_1027_0,
    i_8_358_1031_0, i_8_358_1044_0, i_8_358_1112_0, i_8_358_1135_0,
    i_8_358_1154_0, i_8_358_1155_0, i_8_358_1229_0, i_8_358_1297_0,
    i_8_358_1300_0, i_8_358_1305_0, i_8_358_1306_0, i_8_358_1314_0,
    i_8_358_1341_0, i_8_358_1342_0, i_8_358_1343_0, i_8_358_1345_0,
    i_8_358_1346_0, i_8_358_1349_0, i_8_358_1355_0, i_8_358_1407_0,
    i_8_358_1434_0, i_8_358_1435_0, i_8_358_1436_0, i_8_358_1455_0,
    i_8_358_1542_0, i_8_358_1545_0, i_8_358_1548_0, i_8_358_1550_0,
    i_8_358_1551_0, i_8_358_1624_0, i_8_358_1647_0, i_8_358_1651_0,
    i_8_358_1652_0, i_8_358_1677_0, i_8_358_1682_0, i_8_358_1741_0,
    i_8_358_1748_0, i_8_358_1779_0, i_8_358_1803_0, i_8_358_1866_0,
    i_8_358_1884_0, i_8_358_1925_0, i_8_358_1945_0, i_8_358_1962_0,
    i_8_358_1983_0, i_8_358_1992_0, i_8_358_1994_0, i_8_358_1996_0,
    i_8_358_2049_0, i_8_358_2051_0, i_8_358_2147_0, i_8_358_2245_0,
    i_8_358_2271_0, i_8_358_2286_0, i_8_358_2290_0, i_8_358_2291_0,
    o_8_358_0_0  );
  input  i_8_358_104_0, i_8_358_153_0, i_8_358_154_0, i_8_358_155_0,
    i_8_358_158_0, i_8_358_160_0, i_8_358_205_0, i_8_358_206_0,
    i_8_358_221_0, i_8_358_435_0, i_8_358_471_0, i_8_358_480_0,
    i_8_358_489_0, i_8_358_499_0, i_8_358_500_0, i_8_358_572_0,
    i_8_358_592_0, i_8_358_606_0, i_8_358_610_0, i_8_358_624_0,
    i_8_358_684_0, i_8_358_688_0, i_8_358_699_0, i_8_358_714_0,
    i_8_358_716_0, i_8_358_717_0, i_8_358_729_0, i_8_358_778_0,
    i_8_358_779_0, i_8_358_780_0, i_8_358_782_0, i_8_358_787_0,
    i_8_358_837_0, i_8_358_838_0, i_8_358_867_0, i_8_358_869_0,
    i_8_358_871_0, i_8_358_879_0, i_8_358_881_0, i_8_358_998_0,
    i_8_358_1008_0, i_8_358_1012_0, i_8_358_1026_0, i_8_358_1027_0,
    i_8_358_1031_0, i_8_358_1044_0, i_8_358_1112_0, i_8_358_1135_0,
    i_8_358_1154_0, i_8_358_1155_0, i_8_358_1229_0, i_8_358_1297_0,
    i_8_358_1300_0, i_8_358_1305_0, i_8_358_1306_0, i_8_358_1314_0,
    i_8_358_1341_0, i_8_358_1342_0, i_8_358_1343_0, i_8_358_1345_0,
    i_8_358_1346_0, i_8_358_1349_0, i_8_358_1355_0, i_8_358_1407_0,
    i_8_358_1434_0, i_8_358_1435_0, i_8_358_1436_0, i_8_358_1455_0,
    i_8_358_1542_0, i_8_358_1545_0, i_8_358_1548_0, i_8_358_1550_0,
    i_8_358_1551_0, i_8_358_1624_0, i_8_358_1647_0, i_8_358_1651_0,
    i_8_358_1652_0, i_8_358_1677_0, i_8_358_1682_0, i_8_358_1741_0,
    i_8_358_1748_0, i_8_358_1779_0, i_8_358_1803_0, i_8_358_1866_0,
    i_8_358_1884_0, i_8_358_1925_0, i_8_358_1945_0, i_8_358_1962_0,
    i_8_358_1983_0, i_8_358_1992_0, i_8_358_1994_0, i_8_358_1996_0,
    i_8_358_2049_0, i_8_358_2051_0, i_8_358_2147_0, i_8_358_2245_0,
    i_8_358_2271_0, i_8_358_2286_0, i_8_358_2290_0, i_8_358_2291_0;
  output o_8_358_0_0;
  assign o_8_358_0_0 = ~((~i_8_358_592_0 & ((~i_8_358_104_0 & ~i_8_358_435_0 & i_8_358_572_0 & ~i_8_358_606_0 & ~i_8_358_1342_0 & ~i_8_358_1349_0) | (~i_8_358_153_0 & ~i_8_358_221_0 & ~i_8_358_624_0 & ~i_8_358_717_0 & ~i_8_358_871_0 & ~i_8_358_1436_0 & i_8_358_2271_0))) | (i_8_358_838_0 & ((~i_8_358_153_0 & ~i_8_358_716_0 & ~i_8_358_782_0 & ~i_8_358_1548_0 & ~i_8_358_1550_0 & ~i_8_358_1866_0 & ~i_8_358_2271_0) | (~i_8_358_480_0 & ~i_8_358_500_0 & ~i_8_358_1012_0 & ~i_8_358_1349_0 & ~i_8_358_2290_0))) | (~i_8_358_2051_0 & ((~i_8_358_1803_0 & ((~i_8_358_104_0 & ((~i_8_358_154_0 & ~i_8_358_1154_0 & ~i_8_358_1407_0 & i_8_358_1435_0 & i_8_358_1925_0) | (~i_8_358_155_0 & ~i_8_358_471_0 & ~i_8_358_716_0 & ~i_8_358_1008_0 & ~i_8_358_1341_0 & ~i_8_358_1342_0 & ~i_8_358_1355_0 & ~i_8_358_2049_0 & ~i_8_358_2290_0))) | (~i_8_358_154_0 & ~i_8_358_205_0 & ~i_8_358_206_0 & ~i_8_358_499_0 & ~i_8_358_500_0 & ~i_8_358_624_0 & ~i_8_358_871_0 & ~i_8_358_1012_0 & ~i_8_358_1342_0 & ~i_8_358_1345_0 & ~i_8_358_1435_0 & ~i_8_358_1866_0 & ~i_8_358_1945_0))) | (~i_8_358_160_0 & ((~i_8_358_154_0 & ((~i_8_358_206_0 & ~i_8_358_499_0 & ~i_8_358_624_0 & ~i_8_358_1008_0 & ~i_8_358_1026_0 & ~i_8_358_1343_0 & ~i_8_358_1435_0 & ~i_8_358_1436_0 & ~i_8_358_2049_0) | (~i_8_358_158_0 & ~i_8_358_714_0 & ~i_8_358_998_0 & i_8_358_1994_0 & ~i_8_358_2286_0))) | (~i_8_358_155_0 & ~i_8_358_158_0 & ~i_8_358_780_0 & ~i_8_358_1044_0 & ~i_8_358_1341_0 & ~i_8_358_1342_0 & i_8_358_1435_0 & ~i_8_358_1925_0 & ~i_8_358_1945_0 & ~i_8_358_1983_0 & ~i_8_358_2245_0))) | (~i_8_358_206_0 & ((~i_8_358_205_0 & ~i_8_358_716_0 & i_8_358_1355_0 & ~i_8_358_1866_0 & ~i_8_358_1983_0) | (i_8_358_699_0 & ~i_8_358_714_0 & ~i_8_358_1031_0 & ~i_8_358_1346_0 & ~i_8_358_1748_0 & ~i_8_358_2290_0))) | (~i_8_358_205_0 & ~i_8_358_1155_0 & ((~i_8_358_500_0 & i_8_358_610_0 & ~i_8_358_1026_0 & ~i_8_358_1748_0 & i_8_358_1803_0 & ~i_8_358_1996_0) | (~i_8_358_221_0 & ~i_8_358_716_0 & ~i_8_358_869_0 & ~i_8_358_1300_0 & ~i_8_358_1342_0 & ~i_8_358_1343_0 & ~i_8_358_1548_0 & ~i_8_358_1647_0 & ~i_8_358_1677_0 & ~i_8_358_2049_0 & ~i_8_358_2147_0))) | (~i_8_358_480_0 & ~i_8_358_1748_0 & ~i_8_358_2049_0 & ((~i_8_358_155_0 & ~i_8_358_716_0 & ~i_8_358_717_0 & ~i_8_358_869_0 & ~i_8_358_1341_0 & ~i_8_358_1345_0 & ~i_8_358_1346_0 & ~i_8_358_1435_0 & ~i_8_358_1436_0 & ~i_8_358_1925_0) | (~i_8_358_153_0 & ~i_8_358_435_0 & ~i_8_358_1044_0 & ~i_8_358_1112_0 & ~i_8_358_1154_0 & i_8_358_1346_0 & ~i_8_358_1647_0 & ~i_8_358_1945_0))) | (~i_8_358_624_0 & ~i_8_358_780_0 & ~i_8_358_782_0 & ~i_8_358_871_0 & ~i_8_358_1026_0 & ~i_8_358_1031_0 & ~i_8_358_1341_0 & ~i_8_358_1436_0 & ~i_8_358_1550_0))) | (~i_8_358_1343_0 & ((~i_8_358_160_0 & ~i_8_358_471_0 & ~i_8_358_2290_0 & ((~i_8_358_153_0 & ~i_8_358_154_0 & ~i_8_358_155_0 & ~i_8_358_221_0 & ~i_8_358_782_0 & ~i_8_358_1345_0 & ~i_8_358_1455_0 & ~i_8_358_1677_0) | (i_8_358_592_0 & ~i_8_358_624_0 & ~i_8_358_716_0 & ~i_8_358_717_0 & ~i_8_358_779_0 & ~i_8_358_2049_0))) | (~i_8_358_153_0 & ~i_8_358_155_0 & ~i_8_358_206_0 & ((~i_8_358_158_0 & ~i_8_358_435_0 & ~i_8_358_480_0 & ~i_8_358_714_0 & ~i_8_358_869_0 & ~i_8_358_998_0 & ~i_8_358_1026_0 & ~i_8_358_1031_0 & ~i_8_358_1342_0 & ~i_8_358_2049_0) | (~i_8_358_154_0 & ~i_8_358_205_0 & ~i_8_358_624_0 & ~i_8_358_716_0 & ~i_8_358_780_0 & ~i_8_358_782_0 & ~i_8_358_1027_0 & ~i_8_358_1112_0 & ~i_8_358_1349_0 & ~i_8_358_1355_0 & ~i_8_358_1647_0 & ~i_8_358_2271_0))) | (~i_8_358_154_0 & ~i_8_358_221_0 & ~i_8_358_778_0 & ~i_8_358_782_0 & ~i_8_358_867_0 & ~i_8_358_1112_0 & ~i_8_358_1346_0 & ~i_8_358_1436_0 & ~i_8_358_1551_0 & ~i_8_358_1779_0 & ~i_8_358_1992_0 & ~i_8_358_2049_0))) | (~i_8_358_153_0 & ((~i_8_358_499_0 & ~i_8_358_716_0 & ~i_8_358_998_0 & ~i_8_358_1155_0 & ~i_8_358_1355_0 & i_8_358_1884_0) | (~i_8_358_158_0 & ~i_8_358_205_0 & ~i_8_358_480_0 & ~i_8_358_500_0 & ~i_8_358_1026_0 & i_8_358_1866_0 & ~i_8_358_2291_0))) | (~i_8_358_1435_0 & ((~i_8_358_155_0 & ~i_8_358_1434_0 & ((i_8_358_500_0 & i_8_358_1229_0 & ~i_8_358_2271_0) | (~i_8_358_154_0 & ~i_8_358_206_0 & ~i_8_358_779_0 & ~i_8_358_782_0 & ~i_8_358_1008_0 & ~i_8_358_1342_0 & ~i_8_358_1349_0 & ~i_8_358_2049_0 & ~i_8_358_2286_0))) | (~i_8_358_1803_0 & i_8_358_1994_0 & i_8_358_2051_0))) | (~i_8_358_154_0 & ((~i_8_358_871_0 & ~i_8_358_1027_0 & ~i_8_358_1551_0 & i_8_358_1652_0) | (~i_8_358_158_0 & ~i_8_358_480_0 & ~i_8_358_1306_0 & ~i_8_358_1345_0 & i_8_358_1992_0))) | (~i_8_358_480_0 & ~i_8_358_1008_0 & ((i_8_358_435_0 & i_8_358_780_0 & ~i_8_358_1407_0 & ~i_8_358_1548_0) | (~i_8_358_606_0 & ~i_8_358_714_0 & ~i_8_358_871_0 & ~i_8_358_1112_0 & ~i_8_358_1341_0 & ~i_8_358_1342_0 & ~i_8_358_1682_0 & ~i_8_358_1748_0 & ~i_8_358_1803_0))) | (~i_8_358_717_0 & ((~i_8_358_205_0 & ~i_8_358_435_0 & ~i_8_358_499_0 & i_8_358_881_0 & ~i_8_358_1027_0 & ~i_8_358_1135_0 & ~i_8_358_1154_0 & ~i_8_358_1341_0 & ~i_8_358_1346_0) | (i_8_358_489_0 & i_8_358_837_0 & ~i_8_358_1550_0))) | (~i_8_358_205_0 & ~i_8_358_1155_0 & ~i_8_358_1341_0 & ((~i_8_358_158_0 & ~i_8_358_206_0 & ~i_8_358_1026_0 & ~i_8_358_2049_0 & i_8_358_2147_0) | (~i_8_358_782_0 & i_8_358_1647_0 & ~i_8_358_1866_0 & ~i_8_358_2291_0))) | (~i_8_358_1866_0 & ((~i_8_358_104_0 & ~i_8_358_779_0 & ~i_8_358_998_0 & ~i_8_358_1026_0 & i_8_358_1297_0) | (~i_8_358_1027_0 & i_8_358_1314_0 & i_8_358_1647_0))));
endmodule



// Benchmark "kernel_8_359" written by ABC on Sun Jul 19 10:09:18 2020

module kernel_8_359 ( 
    i_8_359_10_0, i_8_359_20_0, i_8_359_35_0, i_8_359_65_0, i_8_359_73_0,
    i_8_359_74_0, i_8_359_77_0, i_8_359_106_0, i_8_359_113_0,
    i_8_359_124_0, i_8_359_266_0, i_8_359_302_0, i_8_359_322_0,
    i_8_359_323_0, i_8_359_361_0, i_8_359_362_0, i_8_359_364_0,
    i_8_359_365_0, i_8_359_368_0, i_8_359_392_0, i_8_359_398_0,
    i_8_359_428_0, i_8_359_445_0, i_8_359_487_0, i_8_359_505_0,
    i_8_359_506_0, i_8_359_509_0, i_8_359_578_0, i_8_359_590_0,
    i_8_359_604_0, i_8_359_605_0, i_8_359_607_0, i_8_359_608_0,
    i_8_359_641_0, i_8_359_661_0, i_8_359_671_0, i_8_359_677_0,
    i_8_359_680_0, i_8_359_727_0, i_8_359_758_0, i_8_359_781_0,
    i_8_359_817_0, i_8_359_824_0, i_8_359_826_0, i_8_359_955_0,
    i_8_359_974_0, i_8_359_1037_0, i_8_359_1040_0, i_8_359_1109_0,
    i_8_359_1114_0, i_8_359_1127_0, i_8_359_1181_0, i_8_359_1183_0,
    i_8_359_1199_0, i_8_359_1225_0, i_8_359_1229_0, i_8_359_1244_0,
    i_8_359_1264_0, i_8_359_1265_0, i_8_359_1280_0, i_8_359_1295_0,
    i_8_359_1307_0, i_8_359_1315_0, i_8_359_1316_0, i_8_359_1325_0,
    i_8_359_1361_0, i_8_359_1397_0, i_8_359_1424_0, i_8_359_1436_0,
    i_8_359_1438_0, i_8_359_1460_0, i_8_359_1463_0, i_8_359_1465_0,
    i_8_359_1492_0, i_8_359_1510_0, i_8_359_1514_0, i_8_359_1522_0,
    i_8_359_1525_0, i_8_359_1549_0, i_8_359_1550_0, i_8_359_1553_0,
    i_8_359_1630_0, i_8_359_1631_0, i_8_359_1634_0, i_8_359_1679_0,
    i_8_359_1702_0, i_8_359_1747_0, i_8_359_1748_0, i_8_359_1792_0,
    i_8_359_1805_0, i_8_359_1819_0, i_8_359_1822_0, i_8_359_1838_0,
    i_8_359_1883_0, i_8_359_1976_0, i_8_359_1982_0, i_8_359_1993_0,
    i_8_359_2135_0, i_8_359_2245_0, i_8_359_2246_0,
    o_8_359_0_0  );
  input  i_8_359_10_0, i_8_359_20_0, i_8_359_35_0, i_8_359_65_0,
    i_8_359_73_0, i_8_359_74_0, i_8_359_77_0, i_8_359_106_0, i_8_359_113_0,
    i_8_359_124_0, i_8_359_266_0, i_8_359_302_0, i_8_359_322_0,
    i_8_359_323_0, i_8_359_361_0, i_8_359_362_0, i_8_359_364_0,
    i_8_359_365_0, i_8_359_368_0, i_8_359_392_0, i_8_359_398_0,
    i_8_359_428_0, i_8_359_445_0, i_8_359_487_0, i_8_359_505_0,
    i_8_359_506_0, i_8_359_509_0, i_8_359_578_0, i_8_359_590_0,
    i_8_359_604_0, i_8_359_605_0, i_8_359_607_0, i_8_359_608_0,
    i_8_359_641_0, i_8_359_661_0, i_8_359_671_0, i_8_359_677_0,
    i_8_359_680_0, i_8_359_727_0, i_8_359_758_0, i_8_359_781_0,
    i_8_359_817_0, i_8_359_824_0, i_8_359_826_0, i_8_359_955_0,
    i_8_359_974_0, i_8_359_1037_0, i_8_359_1040_0, i_8_359_1109_0,
    i_8_359_1114_0, i_8_359_1127_0, i_8_359_1181_0, i_8_359_1183_0,
    i_8_359_1199_0, i_8_359_1225_0, i_8_359_1229_0, i_8_359_1244_0,
    i_8_359_1264_0, i_8_359_1265_0, i_8_359_1280_0, i_8_359_1295_0,
    i_8_359_1307_0, i_8_359_1315_0, i_8_359_1316_0, i_8_359_1325_0,
    i_8_359_1361_0, i_8_359_1397_0, i_8_359_1424_0, i_8_359_1436_0,
    i_8_359_1438_0, i_8_359_1460_0, i_8_359_1463_0, i_8_359_1465_0,
    i_8_359_1492_0, i_8_359_1510_0, i_8_359_1514_0, i_8_359_1522_0,
    i_8_359_1525_0, i_8_359_1549_0, i_8_359_1550_0, i_8_359_1553_0,
    i_8_359_1630_0, i_8_359_1631_0, i_8_359_1634_0, i_8_359_1679_0,
    i_8_359_1702_0, i_8_359_1747_0, i_8_359_1748_0, i_8_359_1792_0,
    i_8_359_1805_0, i_8_359_1819_0, i_8_359_1822_0, i_8_359_1838_0,
    i_8_359_1883_0, i_8_359_1976_0, i_8_359_1982_0, i_8_359_1993_0,
    i_8_359_2135_0, i_8_359_2245_0, i_8_359_2246_0;
  output o_8_359_0_0;
  assign o_8_359_0_0 = 0;
endmodule



// Benchmark "kernel_8_360" written by ABC on Sun Jul 19 10:09:19 2020

module kernel_8_360 ( 
    i_8_360_26_0, i_8_360_63_0, i_8_360_76_0, i_8_360_192_0, i_8_360_279_0,
    i_8_360_318_0, i_8_360_324_0, i_8_360_327_0, i_8_360_350_0,
    i_8_360_367_0, i_8_360_373_0, i_8_360_383_0, i_8_360_391_0,
    i_8_360_450_0, i_8_360_504_0, i_8_360_526_0, i_8_360_531_0,
    i_8_360_556_0, i_8_360_557_0, i_8_360_562_0, i_8_360_585_0,
    i_8_360_589_0, i_8_360_602_0, i_8_360_603_0, i_8_360_604_0,
    i_8_360_607_0, i_8_360_630_0, i_8_360_631_0, i_8_360_639_0,
    i_8_360_675_0, i_8_360_676_0, i_8_360_700_0, i_8_360_702_0,
    i_8_360_703_0, i_8_360_706_0, i_8_360_793_0, i_8_360_838_0,
    i_8_360_937_0, i_8_360_968_0, i_8_360_1008_0, i_8_360_1036_0,
    i_8_360_1047_0, i_8_360_1106_0, i_8_360_1179_0, i_8_360_1197_0,
    i_8_360_1200_0, i_8_360_1225_0, i_8_360_1246_0, i_8_360_1261_0,
    i_8_360_1264_0, i_8_360_1296_0, i_8_360_1298_0, i_8_360_1299_0,
    i_8_360_1315_0, i_8_360_1327_0, i_8_360_1341_0, i_8_360_1354_0,
    i_8_360_1359_0, i_8_360_1362_0, i_8_360_1422_0, i_8_360_1423_0,
    i_8_360_1433_0, i_8_360_1434_0, i_8_360_1440_0, i_8_360_1461_0,
    i_8_360_1476_0, i_8_360_1512_0, i_8_360_1513_0, i_8_360_1515_0,
    i_8_360_1522_0, i_8_360_1539_0, i_8_360_1543_0, i_8_360_1564_0,
    i_8_360_1632_0, i_8_360_1651_0, i_8_360_1682_0, i_8_360_1701_0,
    i_8_360_1747_0, i_8_360_1748_0, i_8_360_1773_0, i_8_360_1786_0,
    i_8_360_1791_0, i_8_360_1810_0, i_8_360_1829_0, i_8_360_1887_0,
    i_8_360_1953_0, i_8_360_1957_0, i_8_360_1989_0, i_8_360_2011_0,
    i_8_360_2072_0, i_8_360_2132_0, i_8_360_2140_0, i_8_360_2142_0,
    i_8_360_2144_0, i_8_360_2145_0, i_8_360_2146_0, i_8_360_2154_0,
    i_8_360_2223_0, i_8_360_2226_0, i_8_360_2227_0,
    o_8_360_0_0  );
  input  i_8_360_26_0, i_8_360_63_0, i_8_360_76_0, i_8_360_192_0,
    i_8_360_279_0, i_8_360_318_0, i_8_360_324_0, i_8_360_327_0,
    i_8_360_350_0, i_8_360_367_0, i_8_360_373_0, i_8_360_383_0,
    i_8_360_391_0, i_8_360_450_0, i_8_360_504_0, i_8_360_526_0,
    i_8_360_531_0, i_8_360_556_0, i_8_360_557_0, i_8_360_562_0,
    i_8_360_585_0, i_8_360_589_0, i_8_360_602_0, i_8_360_603_0,
    i_8_360_604_0, i_8_360_607_0, i_8_360_630_0, i_8_360_631_0,
    i_8_360_639_0, i_8_360_675_0, i_8_360_676_0, i_8_360_700_0,
    i_8_360_702_0, i_8_360_703_0, i_8_360_706_0, i_8_360_793_0,
    i_8_360_838_0, i_8_360_937_0, i_8_360_968_0, i_8_360_1008_0,
    i_8_360_1036_0, i_8_360_1047_0, i_8_360_1106_0, i_8_360_1179_0,
    i_8_360_1197_0, i_8_360_1200_0, i_8_360_1225_0, i_8_360_1246_0,
    i_8_360_1261_0, i_8_360_1264_0, i_8_360_1296_0, i_8_360_1298_0,
    i_8_360_1299_0, i_8_360_1315_0, i_8_360_1327_0, i_8_360_1341_0,
    i_8_360_1354_0, i_8_360_1359_0, i_8_360_1362_0, i_8_360_1422_0,
    i_8_360_1423_0, i_8_360_1433_0, i_8_360_1434_0, i_8_360_1440_0,
    i_8_360_1461_0, i_8_360_1476_0, i_8_360_1512_0, i_8_360_1513_0,
    i_8_360_1515_0, i_8_360_1522_0, i_8_360_1539_0, i_8_360_1543_0,
    i_8_360_1564_0, i_8_360_1632_0, i_8_360_1651_0, i_8_360_1682_0,
    i_8_360_1701_0, i_8_360_1747_0, i_8_360_1748_0, i_8_360_1773_0,
    i_8_360_1786_0, i_8_360_1791_0, i_8_360_1810_0, i_8_360_1829_0,
    i_8_360_1887_0, i_8_360_1953_0, i_8_360_1957_0, i_8_360_1989_0,
    i_8_360_2011_0, i_8_360_2072_0, i_8_360_2132_0, i_8_360_2140_0,
    i_8_360_2142_0, i_8_360_2144_0, i_8_360_2145_0, i_8_360_2146_0,
    i_8_360_2154_0, i_8_360_2223_0, i_8_360_2226_0, i_8_360_2227_0;
  output o_8_360_0_0;
  assign o_8_360_0_0 = 0;
endmodule



// Benchmark "kernel_8_361" written by ABC on Sun Jul 19 10:09:20 2020

module kernel_8_361 ( 
    i_8_361_0_0, i_8_361_63_0, i_8_361_84_0, i_8_361_139_0, i_8_361_283_0,
    i_8_361_381_0, i_8_361_383_0, i_8_361_423_0, i_8_361_482_0,
    i_8_361_499_0, i_8_361_516_0, i_8_361_520_0, i_8_361_525_0,
    i_8_361_526_0, i_8_361_527_0, i_8_361_528_0, i_8_361_549_0,
    i_8_361_579_0, i_8_361_609_0, i_8_361_700_0, i_8_361_704_0,
    i_8_361_705_0, i_8_361_751_0, i_8_361_777_0, i_8_361_778_0,
    i_8_361_850_0, i_8_361_937_0, i_8_361_968_0, i_8_361_970_0,
    i_8_361_1010_0, i_8_361_1047_0, i_8_361_1074_0, i_8_361_1117_0,
    i_8_361_1127_0, i_8_361_1128_0, i_8_361_1138_0, i_8_361_1180_0,
    i_8_361_1227_0, i_8_361_1263_0, i_8_361_1279_0, i_8_361_1283_0,
    i_8_361_1286_0, i_8_361_1294_0, i_8_361_1296_0, i_8_361_1297_0,
    i_8_361_1332_0, i_8_361_1359_0, i_8_361_1395_0, i_8_361_1434_0,
    i_8_361_1437_0, i_8_361_1438_0, i_8_361_1456_0, i_8_361_1457_0,
    i_8_361_1467_0, i_8_361_1469_0, i_8_361_1486_0, i_8_361_1489_0,
    i_8_361_1494_0, i_8_361_1531_0, i_8_361_1585_0, i_8_361_1600_0,
    i_8_361_1601_0, i_8_361_1602_0, i_8_361_1603_0, i_8_361_1620_0,
    i_8_361_1638_0, i_8_361_1664_0, i_8_361_1686_0, i_8_361_1728_0,
    i_8_361_1746_0, i_8_361_1748_0, i_8_361_1756_0, i_8_361_1758_0,
    i_8_361_1765_0, i_8_361_1768_0, i_8_361_1787_0, i_8_361_1789_0,
    i_8_361_1792_0, i_8_361_1804_0, i_8_361_1805_0, i_8_361_1807_0,
    i_8_361_1808_0, i_8_361_1873_0, i_8_361_1881_0, i_8_361_1948_0,
    i_8_361_1951_0, i_8_361_1963_0, i_8_361_1965_0, i_8_361_1966_0,
    i_8_361_1970_0, i_8_361_2047_0, i_8_361_2068_0, i_8_361_2101_0,
    i_8_361_2133_0, i_8_361_2136_0, i_8_361_2140_0, i_8_361_2149_0,
    i_8_361_2226_0, i_8_361_2273_0, i_8_361_2295_0,
    o_8_361_0_0  );
  input  i_8_361_0_0, i_8_361_63_0, i_8_361_84_0, i_8_361_139_0,
    i_8_361_283_0, i_8_361_381_0, i_8_361_383_0, i_8_361_423_0,
    i_8_361_482_0, i_8_361_499_0, i_8_361_516_0, i_8_361_520_0,
    i_8_361_525_0, i_8_361_526_0, i_8_361_527_0, i_8_361_528_0,
    i_8_361_549_0, i_8_361_579_0, i_8_361_609_0, i_8_361_700_0,
    i_8_361_704_0, i_8_361_705_0, i_8_361_751_0, i_8_361_777_0,
    i_8_361_778_0, i_8_361_850_0, i_8_361_937_0, i_8_361_968_0,
    i_8_361_970_0, i_8_361_1010_0, i_8_361_1047_0, i_8_361_1074_0,
    i_8_361_1117_0, i_8_361_1127_0, i_8_361_1128_0, i_8_361_1138_0,
    i_8_361_1180_0, i_8_361_1227_0, i_8_361_1263_0, i_8_361_1279_0,
    i_8_361_1283_0, i_8_361_1286_0, i_8_361_1294_0, i_8_361_1296_0,
    i_8_361_1297_0, i_8_361_1332_0, i_8_361_1359_0, i_8_361_1395_0,
    i_8_361_1434_0, i_8_361_1437_0, i_8_361_1438_0, i_8_361_1456_0,
    i_8_361_1457_0, i_8_361_1467_0, i_8_361_1469_0, i_8_361_1486_0,
    i_8_361_1489_0, i_8_361_1494_0, i_8_361_1531_0, i_8_361_1585_0,
    i_8_361_1600_0, i_8_361_1601_0, i_8_361_1602_0, i_8_361_1603_0,
    i_8_361_1620_0, i_8_361_1638_0, i_8_361_1664_0, i_8_361_1686_0,
    i_8_361_1728_0, i_8_361_1746_0, i_8_361_1748_0, i_8_361_1756_0,
    i_8_361_1758_0, i_8_361_1765_0, i_8_361_1768_0, i_8_361_1787_0,
    i_8_361_1789_0, i_8_361_1792_0, i_8_361_1804_0, i_8_361_1805_0,
    i_8_361_1807_0, i_8_361_1808_0, i_8_361_1873_0, i_8_361_1881_0,
    i_8_361_1948_0, i_8_361_1951_0, i_8_361_1963_0, i_8_361_1965_0,
    i_8_361_1966_0, i_8_361_1970_0, i_8_361_2047_0, i_8_361_2068_0,
    i_8_361_2101_0, i_8_361_2133_0, i_8_361_2136_0, i_8_361_2140_0,
    i_8_361_2149_0, i_8_361_2226_0, i_8_361_2273_0, i_8_361_2295_0;
  output o_8_361_0_0;
  assign o_8_361_0_0 = 0;
endmodule



// Benchmark "kernel_8_362" written by ABC on Sun Jul 19 10:09:21 2020

module kernel_8_362 ( 
    i_8_362_25_0, i_8_362_33_0, i_8_362_62_0, i_8_362_98_0, i_8_362_140_0,
    i_8_362_160_0, i_8_362_192_0, i_8_362_197_0, i_8_362_224_0,
    i_8_362_250_0, i_8_362_268_0, i_8_362_291_0, i_8_362_338_0,
    i_8_362_357_0, i_8_362_359_0, i_8_362_384_0, i_8_362_420_0,
    i_8_362_458_0, i_8_362_464_0, i_8_362_480_0, i_8_362_485_0,
    i_8_362_503_0, i_8_362_522_0, i_8_362_528_0, i_8_362_570_0,
    i_8_362_629_0, i_8_362_709_0, i_8_362_715_0, i_8_362_726_0,
    i_8_362_764_0, i_8_362_787_0, i_8_362_817_0, i_8_362_907_0,
    i_8_362_922_0, i_8_362_924_0, i_8_362_952_0, i_8_362_985_0,
    i_8_362_987_0, i_8_362_1075_0, i_8_362_1113_0, i_8_362_1124_0,
    i_8_362_1128_0, i_8_362_1132_0, i_8_362_1137_0, i_8_362_1138_0,
    i_8_362_1140_0, i_8_362_1194_0, i_8_362_1419_0, i_8_362_1420_0,
    i_8_362_1421_0, i_8_362_1429_0, i_8_362_1437_0, i_8_362_1455_0,
    i_8_362_1483_0, i_8_362_1527_0, i_8_362_1543_0, i_8_362_1545_0,
    i_8_362_1554_0, i_8_362_1601_0, i_8_362_1609_0, i_8_362_1617_0,
    i_8_362_1618_0, i_8_362_1635_0, i_8_362_1663_0, i_8_362_1671_0,
    i_8_362_1672_0, i_8_362_1717_0, i_8_362_1732_0, i_8_362_1733_0,
    i_8_362_1743_0, i_8_362_1744_0, i_8_362_1750_0, i_8_362_1762_0,
    i_8_362_1797_0, i_8_362_1808_0, i_8_362_1821_0, i_8_362_1839_0,
    i_8_362_1872_0, i_8_362_1875_0, i_8_362_1877_0, i_8_362_1880_0,
    i_8_362_1906_0, i_8_362_1921_0, i_8_362_1922_0, i_8_362_1929_0,
    i_8_362_1966_0, i_8_362_1967_0, i_8_362_1984_0, i_8_362_2031_0,
    i_8_362_2049_0, i_8_362_2055_0, i_8_362_2059_0, i_8_362_2096_0,
    i_8_362_2112_0, i_8_362_2120_0, i_8_362_2154_0, i_8_362_2218_0,
    i_8_362_2219_0, i_8_362_2229_0, i_8_362_2274_0,
    o_8_362_0_0  );
  input  i_8_362_25_0, i_8_362_33_0, i_8_362_62_0, i_8_362_98_0,
    i_8_362_140_0, i_8_362_160_0, i_8_362_192_0, i_8_362_197_0,
    i_8_362_224_0, i_8_362_250_0, i_8_362_268_0, i_8_362_291_0,
    i_8_362_338_0, i_8_362_357_0, i_8_362_359_0, i_8_362_384_0,
    i_8_362_420_0, i_8_362_458_0, i_8_362_464_0, i_8_362_480_0,
    i_8_362_485_0, i_8_362_503_0, i_8_362_522_0, i_8_362_528_0,
    i_8_362_570_0, i_8_362_629_0, i_8_362_709_0, i_8_362_715_0,
    i_8_362_726_0, i_8_362_764_0, i_8_362_787_0, i_8_362_817_0,
    i_8_362_907_0, i_8_362_922_0, i_8_362_924_0, i_8_362_952_0,
    i_8_362_985_0, i_8_362_987_0, i_8_362_1075_0, i_8_362_1113_0,
    i_8_362_1124_0, i_8_362_1128_0, i_8_362_1132_0, i_8_362_1137_0,
    i_8_362_1138_0, i_8_362_1140_0, i_8_362_1194_0, i_8_362_1419_0,
    i_8_362_1420_0, i_8_362_1421_0, i_8_362_1429_0, i_8_362_1437_0,
    i_8_362_1455_0, i_8_362_1483_0, i_8_362_1527_0, i_8_362_1543_0,
    i_8_362_1545_0, i_8_362_1554_0, i_8_362_1601_0, i_8_362_1609_0,
    i_8_362_1617_0, i_8_362_1618_0, i_8_362_1635_0, i_8_362_1663_0,
    i_8_362_1671_0, i_8_362_1672_0, i_8_362_1717_0, i_8_362_1732_0,
    i_8_362_1733_0, i_8_362_1743_0, i_8_362_1744_0, i_8_362_1750_0,
    i_8_362_1762_0, i_8_362_1797_0, i_8_362_1808_0, i_8_362_1821_0,
    i_8_362_1839_0, i_8_362_1872_0, i_8_362_1875_0, i_8_362_1877_0,
    i_8_362_1880_0, i_8_362_1906_0, i_8_362_1921_0, i_8_362_1922_0,
    i_8_362_1929_0, i_8_362_1966_0, i_8_362_1967_0, i_8_362_1984_0,
    i_8_362_2031_0, i_8_362_2049_0, i_8_362_2055_0, i_8_362_2059_0,
    i_8_362_2096_0, i_8_362_2112_0, i_8_362_2120_0, i_8_362_2154_0,
    i_8_362_2218_0, i_8_362_2219_0, i_8_362_2229_0, i_8_362_2274_0;
  output o_8_362_0_0;
  assign o_8_362_0_0 = 0;
endmodule



// Benchmark "kernel_8_363" written by ABC on Sun Jul 19 10:09:22 2020

module kernel_8_363 ( 
    i_8_363_31_0, i_8_363_38_0, i_8_363_83_0, i_8_363_139_0, i_8_363_217_0,
    i_8_363_229_0, i_8_363_281_0, i_8_363_304_0, i_8_363_379_0,
    i_8_363_388_0, i_8_363_416_0, i_8_363_425_0, i_8_363_439_0,
    i_8_363_442_0, i_8_363_443_0, i_8_363_453_0, i_8_363_473_0,
    i_8_363_550_0, i_8_363_571_0, i_8_363_585_0, i_8_363_586_0,
    i_8_363_587_0, i_8_363_604_0, i_8_363_605_0, i_8_363_608_0,
    i_8_363_611_0, i_8_363_622_0, i_8_363_631_0, i_8_363_638_0,
    i_8_363_667_0, i_8_363_669_0, i_8_363_677_0, i_8_363_685_0,
    i_8_363_704_0, i_8_363_736_0, i_8_363_749_0, i_8_363_821_0,
    i_8_363_830_0, i_8_363_839_0, i_8_363_864_0, i_8_363_967_0,
    i_8_363_968_0, i_8_363_1009_0, i_8_363_1031_0, i_8_363_1100_0,
    i_8_363_1118_0, i_8_363_1130_0, i_8_363_1154_0, i_8_363_1180_0,
    i_8_363_1181_0, i_8_363_1225_0, i_8_363_1226_0, i_8_363_1234_0,
    i_8_363_1235_0, i_8_363_1270_0, i_8_363_1280_0, i_8_363_1316_0,
    i_8_363_1327_0, i_8_363_1334_0, i_8_363_1406_0, i_8_363_1439_0,
    i_8_363_1460_0, i_8_363_1534_0, i_8_363_1536_0, i_8_363_1549_0,
    i_8_363_1555_0, i_8_363_1595_0, i_8_363_1658_0, i_8_363_1670_0,
    i_8_363_1681_0, i_8_363_1709_0, i_8_363_1745_0, i_8_363_1757_0,
    i_8_363_1758_0, i_8_363_1759_0, i_8_363_1774_0, i_8_363_1837_0,
    i_8_363_1838_0, i_8_363_1841_0, i_8_363_1891_0, i_8_363_1892_0,
    i_8_363_1895_0, i_8_363_1936_0, i_8_363_1963_0, i_8_363_1964_0,
    i_8_363_2008_0, i_8_363_2026_0, i_8_363_2037_0, i_8_363_2072_0,
    i_8_363_2108_0, i_8_363_2110_0, i_8_363_2140_0, i_8_363_2142_0,
    i_8_363_2143_0, i_8_363_2145_0, i_8_363_2152_0, i_8_363_2171_0,
    i_8_363_2188_0, i_8_363_2189_0, i_8_363_2191_0,
    o_8_363_0_0  );
  input  i_8_363_31_0, i_8_363_38_0, i_8_363_83_0, i_8_363_139_0,
    i_8_363_217_0, i_8_363_229_0, i_8_363_281_0, i_8_363_304_0,
    i_8_363_379_0, i_8_363_388_0, i_8_363_416_0, i_8_363_425_0,
    i_8_363_439_0, i_8_363_442_0, i_8_363_443_0, i_8_363_453_0,
    i_8_363_473_0, i_8_363_550_0, i_8_363_571_0, i_8_363_585_0,
    i_8_363_586_0, i_8_363_587_0, i_8_363_604_0, i_8_363_605_0,
    i_8_363_608_0, i_8_363_611_0, i_8_363_622_0, i_8_363_631_0,
    i_8_363_638_0, i_8_363_667_0, i_8_363_669_0, i_8_363_677_0,
    i_8_363_685_0, i_8_363_704_0, i_8_363_736_0, i_8_363_749_0,
    i_8_363_821_0, i_8_363_830_0, i_8_363_839_0, i_8_363_864_0,
    i_8_363_967_0, i_8_363_968_0, i_8_363_1009_0, i_8_363_1031_0,
    i_8_363_1100_0, i_8_363_1118_0, i_8_363_1130_0, i_8_363_1154_0,
    i_8_363_1180_0, i_8_363_1181_0, i_8_363_1225_0, i_8_363_1226_0,
    i_8_363_1234_0, i_8_363_1235_0, i_8_363_1270_0, i_8_363_1280_0,
    i_8_363_1316_0, i_8_363_1327_0, i_8_363_1334_0, i_8_363_1406_0,
    i_8_363_1439_0, i_8_363_1460_0, i_8_363_1534_0, i_8_363_1536_0,
    i_8_363_1549_0, i_8_363_1555_0, i_8_363_1595_0, i_8_363_1658_0,
    i_8_363_1670_0, i_8_363_1681_0, i_8_363_1709_0, i_8_363_1745_0,
    i_8_363_1757_0, i_8_363_1758_0, i_8_363_1759_0, i_8_363_1774_0,
    i_8_363_1837_0, i_8_363_1838_0, i_8_363_1841_0, i_8_363_1891_0,
    i_8_363_1892_0, i_8_363_1895_0, i_8_363_1936_0, i_8_363_1963_0,
    i_8_363_1964_0, i_8_363_2008_0, i_8_363_2026_0, i_8_363_2037_0,
    i_8_363_2072_0, i_8_363_2108_0, i_8_363_2110_0, i_8_363_2140_0,
    i_8_363_2142_0, i_8_363_2143_0, i_8_363_2145_0, i_8_363_2152_0,
    i_8_363_2171_0, i_8_363_2188_0, i_8_363_2189_0, i_8_363_2191_0;
  output o_8_363_0_0;
  assign o_8_363_0_0 = 0;
endmodule



// Benchmark "kernel_8_364" written by ABC on Sun Jul 19 10:09:23 2020

module kernel_8_364 ( 
    i_8_364_12_0, i_8_364_44_0, i_8_364_66_0, i_8_364_106_0, i_8_364_115_0,
    i_8_364_133_0, i_8_364_139_0, i_8_364_172_0, i_8_364_256_0,
    i_8_364_273_0, i_8_364_283_0, i_8_364_309_0, i_8_364_321_0,
    i_8_364_381_0, i_8_364_399_0, i_8_364_400_0, i_8_364_471_0,
    i_8_364_498_0, i_8_364_524_0, i_8_364_549_0, i_8_364_555_0,
    i_8_364_571_0, i_8_364_577_0, i_8_364_591_0, i_8_364_608_0,
    i_8_364_630_0, i_8_364_635_0, i_8_364_642_0, i_8_364_666_0,
    i_8_364_672_0, i_8_364_681_0, i_8_364_707_0, i_8_364_750_0,
    i_8_364_780_0, i_8_364_825_0, i_8_364_841_0, i_8_364_845_0,
    i_8_364_966_0, i_8_364_967_0, i_8_364_1035_0, i_8_364_1038_0,
    i_8_364_1039_0, i_8_364_1042_0, i_8_364_1072_0, i_8_364_1074_0,
    i_8_364_1225_0, i_8_364_1227_0, i_8_364_1236_0, i_8_364_1237_0,
    i_8_364_1246_0, i_8_364_1263_0, i_8_364_1270_0, i_8_364_1300_0,
    i_8_364_1314_0, i_8_364_1317_0, i_8_364_1318_0, i_8_364_1327_0,
    i_8_364_1330_0, i_8_364_1338_0, i_8_364_1362_0, i_8_364_1372_0,
    i_8_364_1390_0, i_8_364_1422_0, i_8_364_1437_0, i_8_364_1442_0,
    i_8_364_1464_0, i_8_364_1465_0, i_8_364_1506_0, i_8_364_1525_0,
    i_8_364_1527_0, i_8_364_1545_0, i_8_364_1564_0, i_8_364_1573_0,
    i_8_364_1623_0, i_8_364_1636_0, i_8_364_1641_0, i_8_364_1651_0,
    i_8_364_1678_0, i_8_364_1681_0, i_8_364_1698_0, i_8_364_1782_0,
    i_8_364_1787_0, i_8_364_1824_0, i_8_364_1893_0, i_8_364_1912_0,
    i_8_364_1938_0, i_8_364_1960_0, i_8_364_1969_0, i_8_364_1975_0,
    i_8_364_1977_0, i_8_364_1984_0, i_8_364_2071_0, i_8_364_2179_0,
    i_8_364_2208_0, i_8_364_2226_0, i_8_364_2231_0, i_8_364_2246_0,
    i_8_364_2247_0, i_8_364_2271_0, i_8_364_2298_0,
    o_8_364_0_0  );
  input  i_8_364_12_0, i_8_364_44_0, i_8_364_66_0, i_8_364_106_0,
    i_8_364_115_0, i_8_364_133_0, i_8_364_139_0, i_8_364_172_0,
    i_8_364_256_0, i_8_364_273_0, i_8_364_283_0, i_8_364_309_0,
    i_8_364_321_0, i_8_364_381_0, i_8_364_399_0, i_8_364_400_0,
    i_8_364_471_0, i_8_364_498_0, i_8_364_524_0, i_8_364_549_0,
    i_8_364_555_0, i_8_364_571_0, i_8_364_577_0, i_8_364_591_0,
    i_8_364_608_0, i_8_364_630_0, i_8_364_635_0, i_8_364_642_0,
    i_8_364_666_0, i_8_364_672_0, i_8_364_681_0, i_8_364_707_0,
    i_8_364_750_0, i_8_364_780_0, i_8_364_825_0, i_8_364_841_0,
    i_8_364_845_0, i_8_364_966_0, i_8_364_967_0, i_8_364_1035_0,
    i_8_364_1038_0, i_8_364_1039_0, i_8_364_1042_0, i_8_364_1072_0,
    i_8_364_1074_0, i_8_364_1225_0, i_8_364_1227_0, i_8_364_1236_0,
    i_8_364_1237_0, i_8_364_1246_0, i_8_364_1263_0, i_8_364_1270_0,
    i_8_364_1300_0, i_8_364_1314_0, i_8_364_1317_0, i_8_364_1318_0,
    i_8_364_1327_0, i_8_364_1330_0, i_8_364_1338_0, i_8_364_1362_0,
    i_8_364_1372_0, i_8_364_1390_0, i_8_364_1422_0, i_8_364_1437_0,
    i_8_364_1442_0, i_8_364_1464_0, i_8_364_1465_0, i_8_364_1506_0,
    i_8_364_1525_0, i_8_364_1527_0, i_8_364_1545_0, i_8_364_1564_0,
    i_8_364_1573_0, i_8_364_1623_0, i_8_364_1636_0, i_8_364_1641_0,
    i_8_364_1651_0, i_8_364_1678_0, i_8_364_1681_0, i_8_364_1698_0,
    i_8_364_1782_0, i_8_364_1787_0, i_8_364_1824_0, i_8_364_1893_0,
    i_8_364_1912_0, i_8_364_1938_0, i_8_364_1960_0, i_8_364_1969_0,
    i_8_364_1975_0, i_8_364_1977_0, i_8_364_1984_0, i_8_364_2071_0,
    i_8_364_2179_0, i_8_364_2208_0, i_8_364_2226_0, i_8_364_2231_0,
    i_8_364_2246_0, i_8_364_2247_0, i_8_364_2271_0, i_8_364_2298_0;
  output o_8_364_0_0;
  assign o_8_364_0_0 = 0;
endmodule



// Benchmark "kernel_8_365" written by ABC on Sun Jul 19 10:09:25 2020

module kernel_8_365 ( 
    i_8_365_18_0, i_8_365_19_0, i_8_365_47_0, i_8_365_51_0, i_8_365_54_0,
    i_8_365_55_0, i_8_365_58_0, i_8_365_138_0, i_8_365_216_0,
    i_8_365_228_0, i_8_365_229_0, i_8_365_252_0, i_8_365_272_0,
    i_8_365_292_0, i_8_365_350_0, i_8_365_363_0, i_8_365_399_0,
    i_8_365_427_0, i_8_365_433_0, i_8_365_436_0, i_8_365_457_0,
    i_8_365_552_0, i_8_365_597_0, i_8_365_615_0, i_8_365_621_0,
    i_8_365_631_0, i_8_365_657_0, i_8_365_664_0, i_8_365_665_0,
    i_8_365_689_0, i_8_365_697_0, i_8_365_699_0, i_8_365_709_0,
    i_8_365_716_0, i_8_365_729_0, i_8_365_730_0, i_8_365_759_0,
    i_8_365_783_0, i_8_365_792_0, i_8_365_847_0, i_8_365_880_0,
    i_8_365_990_0, i_8_365_998_0, i_8_365_1027_0, i_8_365_1045_0,
    i_8_365_1047_0, i_8_365_1077_0, i_8_365_1090_0, i_8_365_1109_0,
    i_8_365_1117_0, i_8_365_1129_0, i_8_365_1188_0, i_8_365_1233_0,
    i_8_365_1266_0, i_8_365_1270_0, i_8_365_1317_0, i_8_365_1369_0,
    i_8_365_1436_0, i_8_365_1441_0, i_8_365_1449_0, i_8_365_1452_0,
    i_8_365_1467_0, i_8_365_1468_0, i_8_365_1505_0, i_8_365_1534_0,
    i_8_365_1539_0, i_8_365_1546_0, i_8_365_1562_0, i_8_365_1591_0,
    i_8_365_1603_0, i_8_365_1611_0, i_8_365_1620_0, i_8_365_1629_0,
    i_8_365_1658_0, i_8_365_1666_0, i_8_365_1676_0, i_8_365_1678_0,
    i_8_365_1679_0, i_8_365_1681_0, i_8_365_1682_0, i_8_365_1740_0,
    i_8_365_1802_0, i_8_365_1855_0, i_8_365_1856_0, i_8_365_1873_0,
    i_8_365_1989_0, i_8_365_1991_0, i_8_365_2029_0, i_8_365_2035_0,
    i_8_365_2046_0, i_8_365_2053_0, i_8_365_2093_0, i_8_365_2125_0,
    i_8_365_2138_0, i_8_365_2139_0, i_8_365_2156_0, i_8_365_2232_0,
    i_8_365_2259_0, i_8_365_2261_0, i_8_365_2286_0,
    o_8_365_0_0  );
  input  i_8_365_18_0, i_8_365_19_0, i_8_365_47_0, i_8_365_51_0,
    i_8_365_54_0, i_8_365_55_0, i_8_365_58_0, i_8_365_138_0, i_8_365_216_0,
    i_8_365_228_0, i_8_365_229_0, i_8_365_252_0, i_8_365_272_0,
    i_8_365_292_0, i_8_365_350_0, i_8_365_363_0, i_8_365_399_0,
    i_8_365_427_0, i_8_365_433_0, i_8_365_436_0, i_8_365_457_0,
    i_8_365_552_0, i_8_365_597_0, i_8_365_615_0, i_8_365_621_0,
    i_8_365_631_0, i_8_365_657_0, i_8_365_664_0, i_8_365_665_0,
    i_8_365_689_0, i_8_365_697_0, i_8_365_699_0, i_8_365_709_0,
    i_8_365_716_0, i_8_365_729_0, i_8_365_730_0, i_8_365_759_0,
    i_8_365_783_0, i_8_365_792_0, i_8_365_847_0, i_8_365_880_0,
    i_8_365_990_0, i_8_365_998_0, i_8_365_1027_0, i_8_365_1045_0,
    i_8_365_1047_0, i_8_365_1077_0, i_8_365_1090_0, i_8_365_1109_0,
    i_8_365_1117_0, i_8_365_1129_0, i_8_365_1188_0, i_8_365_1233_0,
    i_8_365_1266_0, i_8_365_1270_0, i_8_365_1317_0, i_8_365_1369_0,
    i_8_365_1436_0, i_8_365_1441_0, i_8_365_1449_0, i_8_365_1452_0,
    i_8_365_1467_0, i_8_365_1468_0, i_8_365_1505_0, i_8_365_1534_0,
    i_8_365_1539_0, i_8_365_1546_0, i_8_365_1562_0, i_8_365_1591_0,
    i_8_365_1603_0, i_8_365_1611_0, i_8_365_1620_0, i_8_365_1629_0,
    i_8_365_1658_0, i_8_365_1666_0, i_8_365_1676_0, i_8_365_1678_0,
    i_8_365_1679_0, i_8_365_1681_0, i_8_365_1682_0, i_8_365_1740_0,
    i_8_365_1802_0, i_8_365_1855_0, i_8_365_1856_0, i_8_365_1873_0,
    i_8_365_1989_0, i_8_365_1991_0, i_8_365_2029_0, i_8_365_2035_0,
    i_8_365_2046_0, i_8_365_2053_0, i_8_365_2093_0, i_8_365_2125_0,
    i_8_365_2138_0, i_8_365_2139_0, i_8_365_2156_0, i_8_365_2232_0,
    i_8_365_2259_0, i_8_365_2261_0, i_8_365_2286_0;
  output o_8_365_0_0;
  assign o_8_365_0_0 = ~((~i_8_365_272_0 & ((~i_8_365_51_0 & ~i_8_365_54_0 & i_8_365_729_0 & ~i_8_365_1467_0 & ~i_8_365_1629_0) | (~i_8_365_47_0 & ~i_8_365_1129_0 & i_8_365_1188_0 & ~i_8_365_1562_0 & i_8_365_1620_0 & ~i_8_365_1681_0))) | (~i_8_365_292_0 & ((~i_8_365_18_0 & ~i_8_365_847_0 & ~i_8_365_880_0 & ~i_8_365_1045_0 & ~i_8_365_1117_0 & ~i_8_365_1441_0 & ~i_8_365_1629_0 & ~i_8_365_1856_0) | (~i_8_365_47_0 & ~i_8_365_51_0 & ~i_8_365_399_0 & ~i_8_365_457_0 & ~i_8_365_689_0 & ~i_8_365_990_0 & i_8_365_1270_0 & ~i_8_365_1989_0 & ~i_8_365_2093_0 & ~i_8_365_2138_0))) | (~i_8_365_51_0 & ((~i_8_365_47_0 & i_8_365_615_0 & ~i_8_365_1027_0 & ~i_8_365_1045_0 & i_8_365_1266_0 & ~i_8_365_1611_0 & ~i_8_365_2261_0) | (~i_8_365_54_0 & i_8_365_216_0 & ~i_8_365_665_0 & ~i_8_365_689_0 & ~i_8_365_847_0 & ~i_8_365_1467_0 & ~i_8_365_2035_0 & ~i_8_365_2259_0 & ~i_8_365_2286_0))) | (~i_8_365_783_0 & ((~i_8_365_54_0 & ((~i_8_365_47_0 & ~i_8_365_55_0 & ~i_8_365_597_0 & ~i_8_365_990_0 & ~i_8_365_1266_0 & ~i_8_365_1270_0 & ~i_8_365_1467_0 & i_8_365_1603_0) | (~i_8_365_252_0 & ~i_8_365_1117_0 & ~i_8_365_1436_0 & ~i_8_365_1505_0 & ~i_8_365_1534_0 & ~i_8_365_1603_0 & ~i_8_365_1611_0 & ~i_8_365_1678_0 & ~i_8_365_1855_0 & ~i_8_365_2156_0 & ~i_8_365_2259_0 & ~i_8_365_2261_0 & ~i_8_365_2286_0))) | (~i_8_365_55_0 & ((i_8_365_552_0 & ~i_8_365_631_0 & ~i_8_365_998_0 & ~i_8_365_1047_0 & ~i_8_365_2093_0) | (~i_8_365_1109_0 & ~i_8_365_1117_0 & ~i_8_365_1467_0 & ~i_8_365_1873_0 & ~i_8_365_1989_0 & ~i_8_365_2259_0))) | (~i_8_365_252_0 & i_8_365_631_0 & ~i_8_365_847_0 & ~i_8_365_2156_0 & ~i_8_365_2259_0 & ~i_8_365_1603_0 & ~i_8_365_2035_0) | (~i_8_365_228_0 & ~i_8_365_689_0 & ~i_8_365_709_0 & i_8_365_880_0 & ~i_8_365_1317_0 & ~i_8_365_1505_0 & ~i_8_365_1539_0 & ~i_8_365_1562_0 & ~i_8_365_2046_0 & ~i_8_365_2261_0 & ~i_8_365_2286_0))) | (~i_8_365_1989_0 & ((~i_8_365_1991_0 & ((~i_8_365_47_0 & ((~i_8_365_1270_0 & i_8_365_1562_0 & ~i_8_365_1658_0) | (~i_8_365_58_0 & ~i_8_365_228_0 & ~i_8_365_998_0 & ~i_8_365_1539_0 & ~i_8_365_1546_0 & ~i_8_365_1740_0 & ~i_8_365_2093_0 & ~i_8_365_2232_0))) | (i_8_365_1452_0 & i_8_365_1855_0))) | (~i_8_365_138_0 & ~i_8_365_350_0 & ~i_8_365_1562_0 & ((~i_8_365_730_0 & ~i_8_365_1045_0 & ~i_8_365_1109_0 & ~i_8_365_1534_0 & ~i_8_365_1629_0 & ~i_8_365_1682_0) | (~i_8_365_631_0 & ~i_8_365_709_0 & ~i_8_365_847_0 & ~i_8_365_1740_0 & ~i_8_365_1856_0 & ~i_8_365_2138_0 & ~i_8_365_2156_0 & ~i_8_365_2232_0))))) | (~i_8_365_58_0 & ((i_8_365_759_0 & ~i_8_365_1090_0 & ~i_8_365_1468_0 & ~i_8_365_1678_0 & ~i_8_365_1681_0 & ~i_8_365_2156_0) | (~i_8_365_55_0 & ~i_8_365_631_0 & ~i_8_365_699_0 & ~i_8_365_730_0 & ~i_8_365_759_0 & ~i_8_365_792_0 & ~i_8_365_1441_0 & ~i_8_365_1629_0 & ~i_8_365_1740_0 & ~i_8_365_2232_0 & ~i_8_365_2286_0))) | (~i_8_365_1562_0 & ((~i_8_365_55_0 & ((~i_8_365_138_0 & ~i_8_365_631_0 & ~i_8_365_689_0 & ~i_8_365_1117_0 & ~i_8_365_1233_0 & ~i_8_365_1467_0 & ~i_8_365_1629_0 & ~i_8_365_1740_0) | (~i_8_365_252_0 & i_8_365_427_0 & ~i_8_365_1047_0 & ~i_8_365_1468_0 & ~i_8_365_1873_0 & ~i_8_365_2232_0))) | (~i_8_365_1658_0 & ((i_8_365_363_0 & ~i_8_365_998_0 & ~i_8_365_1117_0 & ~i_8_365_1591_0 & i_8_365_1682_0 & ~i_8_365_1740_0 & ~i_8_365_2035_0) | (~i_8_365_138_0 & i_8_365_631_0 & ~i_8_365_792_0 & ~i_8_365_990_0 & ~i_8_365_1611_0 & i_8_365_2138_0 & ~i_8_365_2286_0))))) | (~i_8_365_1117_0 & ((~i_8_365_228_0 & ((~i_8_365_847_0 & i_8_365_1534_0 & i_8_365_1679_0 & ~i_8_365_2139_0) | (i_8_365_138_0 & ~i_8_365_729_0 & ~i_8_365_1045_0 & ~i_8_365_1188_0 & ~i_8_365_1629_0 & ~i_8_365_1991_0 & ~i_8_365_2232_0))) | (~i_8_365_1629_0 & ~i_8_365_1856_0 & ~i_8_365_363_0 & i_8_365_1436_0 & ~i_8_365_1873_0 & ~i_8_365_2035_0 & ~i_8_365_2139_0 & i_8_365_2156_0))) | (~i_8_365_657_0 & ((i_8_365_427_0 & ~i_8_365_990_0 & ~i_8_365_1109_0 & ~i_8_365_1467_0 & ~i_8_365_1991_0 & ~i_8_365_2029_0) | (~i_8_365_55_0 & ~i_8_365_1047_0 & ~i_8_365_1658_0 & i_8_365_2138_0 & ~i_8_365_2261_0))) | (~i_8_365_689_0 & ~i_8_365_1452_0 & ((i_8_365_597_0 & ~i_8_365_847_0 & ~i_8_365_1090_0 & ~i_8_365_1129_0 & ~i_8_365_1658_0 & ~i_8_365_1873_0) | (~i_8_365_252_0 & ~i_8_365_1047_0 & ~i_8_365_1270_0 & ~i_8_365_1317_0 & ~i_8_365_1441_0 & ~i_8_365_1467_0 & ~i_8_365_1468_0 & ~i_8_365_1620_0 & ~i_8_365_2053_0 & ~i_8_365_2093_0))) | (~i_8_365_1270_0 & ((~i_8_365_216_0 & ~i_8_365_697_0 & ~i_8_365_1045_0 & ~i_8_365_1188_0 & ~i_8_365_1317_0 & i_8_365_1678_0) | (~i_8_365_427_0 & i_8_365_716_0 & i_8_365_847_0 & ~i_8_365_1873_0 & ~i_8_365_2125_0))) | (~i_8_365_1188_0 & ((i_8_365_1233_0 & i_8_365_1369_0 & ~i_8_365_1539_0 & i_8_365_1611_0) | (~i_8_365_552_0 & i_8_365_1270_0 & ~i_8_365_1505_0 & i_8_365_2286_0))) | (i_8_365_664_0 & i_8_365_1666_0 & i_8_365_2138_0) | (i_8_365_436_0 & i_8_365_2046_0 & ~i_8_365_2139_0) | (~i_8_365_19_0 & ~i_8_365_1266_0 & ~i_8_365_1740_0 & i_8_365_1856_0 & ~i_8_365_2261_0));
endmodule



// Benchmark "kernel_8_366" written by ABC on Sun Jul 19 10:09:26 2020

module kernel_8_366 ( 
    i_8_366_30_0, i_8_366_33_0, i_8_366_53_0, i_8_366_79_0, i_8_366_84_0,
    i_8_366_118_0, i_8_366_138_0, i_8_366_165_0, i_8_366_184_0,
    i_8_366_187_0, i_8_366_192_0, i_8_366_210_0, i_8_366_240_0,
    i_8_366_241_0, i_8_366_301_0, i_8_366_336_0, i_8_366_369_0,
    i_8_366_381_0, i_8_366_382_0, i_8_366_439_0, i_8_366_472_0,
    i_8_366_522_0, i_8_366_543_0, i_8_366_573_0, i_8_366_608_0,
    i_8_366_638_0, i_8_366_760_0, i_8_366_771_0, i_8_366_774_0,
    i_8_366_810_0, i_8_366_811_0, i_8_366_858_0, i_8_366_861_0,
    i_8_366_878_0, i_8_366_879_0, i_8_366_939_0, i_8_366_940_0,
    i_8_366_968_0, i_8_366_984_0, i_8_366_1059_0, i_8_366_1060_0,
    i_8_366_1133_0, i_8_366_1138_0, i_8_366_1182_0, i_8_366_1188_0,
    i_8_366_1191_0, i_8_366_1264_0, i_8_366_1266_0, i_8_366_1269_0,
    i_8_366_1282_0, i_8_366_1287_0, i_8_366_1288_0, i_8_366_1291_0,
    i_8_366_1293_0, i_8_366_1305_0, i_8_366_1326_0, i_8_366_1333_0,
    i_8_366_1386_0, i_8_366_1387_0, i_8_366_1403_0, i_8_366_1407_0,
    i_8_366_1411_0, i_8_366_1489_0, i_8_366_1531_0, i_8_366_1545_0,
    i_8_366_1553_0, i_8_366_1600_0, i_8_366_1614_0, i_8_366_1633_0,
    i_8_366_1678_0, i_8_366_1681_0, i_8_366_1713_0, i_8_366_1719_0,
    i_8_366_1720_0, i_8_366_1731_0, i_8_366_1734_0, i_8_366_1747_0,
    i_8_366_1758_0, i_8_366_1759_0, i_8_366_1771_0, i_8_366_1783_0,
    i_8_366_1790_0, i_8_366_1796_0, i_8_366_1804_0, i_8_366_1822_0,
    i_8_366_1839_0, i_8_366_1857_0, i_8_366_1885_0, i_8_366_1918_0,
    i_8_366_1981_0, i_8_366_1998_0, i_8_366_2022_0, i_8_366_2047_0,
    i_8_366_2056_0, i_8_366_2124_0, i_8_366_2149_0, i_8_366_2169_0,
    i_8_366_2223_0, i_8_366_2235_0, i_8_366_2298_0,
    o_8_366_0_0  );
  input  i_8_366_30_0, i_8_366_33_0, i_8_366_53_0, i_8_366_79_0,
    i_8_366_84_0, i_8_366_118_0, i_8_366_138_0, i_8_366_165_0,
    i_8_366_184_0, i_8_366_187_0, i_8_366_192_0, i_8_366_210_0,
    i_8_366_240_0, i_8_366_241_0, i_8_366_301_0, i_8_366_336_0,
    i_8_366_369_0, i_8_366_381_0, i_8_366_382_0, i_8_366_439_0,
    i_8_366_472_0, i_8_366_522_0, i_8_366_543_0, i_8_366_573_0,
    i_8_366_608_0, i_8_366_638_0, i_8_366_760_0, i_8_366_771_0,
    i_8_366_774_0, i_8_366_810_0, i_8_366_811_0, i_8_366_858_0,
    i_8_366_861_0, i_8_366_878_0, i_8_366_879_0, i_8_366_939_0,
    i_8_366_940_0, i_8_366_968_0, i_8_366_984_0, i_8_366_1059_0,
    i_8_366_1060_0, i_8_366_1133_0, i_8_366_1138_0, i_8_366_1182_0,
    i_8_366_1188_0, i_8_366_1191_0, i_8_366_1264_0, i_8_366_1266_0,
    i_8_366_1269_0, i_8_366_1282_0, i_8_366_1287_0, i_8_366_1288_0,
    i_8_366_1291_0, i_8_366_1293_0, i_8_366_1305_0, i_8_366_1326_0,
    i_8_366_1333_0, i_8_366_1386_0, i_8_366_1387_0, i_8_366_1403_0,
    i_8_366_1407_0, i_8_366_1411_0, i_8_366_1489_0, i_8_366_1531_0,
    i_8_366_1545_0, i_8_366_1553_0, i_8_366_1600_0, i_8_366_1614_0,
    i_8_366_1633_0, i_8_366_1678_0, i_8_366_1681_0, i_8_366_1713_0,
    i_8_366_1719_0, i_8_366_1720_0, i_8_366_1731_0, i_8_366_1734_0,
    i_8_366_1747_0, i_8_366_1758_0, i_8_366_1759_0, i_8_366_1771_0,
    i_8_366_1783_0, i_8_366_1790_0, i_8_366_1796_0, i_8_366_1804_0,
    i_8_366_1822_0, i_8_366_1839_0, i_8_366_1857_0, i_8_366_1885_0,
    i_8_366_1918_0, i_8_366_1981_0, i_8_366_1998_0, i_8_366_2022_0,
    i_8_366_2047_0, i_8_366_2056_0, i_8_366_2124_0, i_8_366_2149_0,
    i_8_366_2169_0, i_8_366_2223_0, i_8_366_2235_0, i_8_366_2298_0;
  output o_8_366_0_0;
  assign o_8_366_0_0 = 0;
endmodule



// Benchmark "kernel_8_367" written by ABC on Sun Jul 19 10:09:27 2020

module kernel_8_367 ( 
    i_8_367_51_0, i_8_367_97_0, i_8_367_120_0, i_8_367_138_0,
    i_8_367_163_0, i_8_367_193_0, i_8_367_202_0, i_8_367_233_0,
    i_8_367_246_0, i_8_367_252_0, i_8_367_256_0, i_8_367_264_0,
    i_8_367_282_0, i_8_367_291_0, i_8_367_292_0, i_8_367_293_0,
    i_8_367_321_0, i_8_367_328_0, i_8_367_330_0, i_8_367_345_0,
    i_8_367_346_0, i_8_367_364_0, i_8_367_394_0, i_8_367_437_0,
    i_8_367_439_0, i_8_367_450_0, i_8_367_455_0, i_8_367_456_0,
    i_8_367_480_0, i_8_367_598_0, i_8_367_601_0, i_8_367_612_0,
    i_8_367_616_0, i_8_367_672_0, i_8_367_701_0, i_8_367_702_0,
    i_8_367_706_0, i_8_367_709_0, i_8_367_715_0, i_8_367_723_0,
    i_8_367_786_0, i_8_367_797_0, i_8_367_822_0, i_8_367_826_0,
    i_8_367_874_0, i_8_367_966_0, i_8_367_969_0, i_8_367_972_0,
    i_8_367_995_0, i_8_367_1050_0, i_8_367_1061_0, i_8_367_1074_0,
    i_8_367_1080_0, i_8_367_1081_0, i_8_367_1119_0, i_8_367_1182_0,
    i_8_367_1234_0, i_8_367_1237_0, i_8_367_1273_0, i_8_367_1347_0,
    i_8_367_1354_0, i_8_367_1389_0, i_8_367_1390_0, i_8_367_1408_0,
    i_8_367_1411_0, i_8_367_1437_0, i_8_367_1439_0, i_8_367_1452_0,
    i_8_367_1464_0, i_8_367_1527_0, i_8_367_1545_0, i_8_367_1546_0,
    i_8_367_1570_0, i_8_367_1573_0, i_8_367_1632_0, i_8_367_1681_0,
    i_8_367_1719_0, i_8_367_1746_0, i_8_367_1758_0, i_8_367_1759_0,
    i_8_367_1867_0, i_8_367_1884_0, i_8_367_1885_0, i_8_367_1887_0,
    i_8_367_1902_0, i_8_367_1948_0, i_8_367_1992_0, i_8_367_1995_0,
    i_8_367_2028_0, i_8_367_2031_0, i_8_367_2056_0, i_8_367_2058_0,
    i_8_367_2077_0, i_8_367_2128_0, i_8_367_2140_0, i_8_367_2156_0,
    i_8_367_2190_0, i_8_367_2215_0, i_8_367_2216_0, i_8_367_2270_0,
    o_8_367_0_0  );
  input  i_8_367_51_0, i_8_367_97_0, i_8_367_120_0, i_8_367_138_0,
    i_8_367_163_0, i_8_367_193_0, i_8_367_202_0, i_8_367_233_0,
    i_8_367_246_0, i_8_367_252_0, i_8_367_256_0, i_8_367_264_0,
    i_8_367_282_0, i_8_367_291_0, i_8_367_292_0, i_8_367_293_0,
    i_8_367_321_0, i_8_367_328_0, i_8_367_330_0, i_8_367_345_0,
    i_8_367_346_0, i_8_367_364_0, i_8_367_394_0, i_8_367_437_0,
    i_8_367_439_0, i_8_367_450_0, i_8_367_455_0, i_8_367_456_0,
    i_8_367_480_0, i_8_367_598_0, i_8_367_601_0, i_8_367_612_0,
    i_8_367_616_0, i_8_367_672_0, i_8_367_701_0, i_8_367_702_0,
    i_8_367_706_0, i_8_367_709_0, i_8_367_715_0, i_8_367_723_0,
    i_8_367_786_0, i_8_367_797_0, i_8_367_822_0, i_8_367_826_0,
    i_8_367_874_0, i_8_367_966_0, i_8_367_969_0, i_8_367_972_0,
    i_8_367_995_0, i_8_367_1050_0, i_8_367_1061_0, i_8_367_1074_0,
    i_8_367_1080_0, i_8_367_1081_0, i_8_367_1119_0, i_8_367_1182_0,
    i_8_367_1234_0, i_8_367_1237_0, i_8_367_1273_0, i_8_367_1347_0,
    i_8_367_1354_0, i_8_367_1389_0, i_8_367_1390_0, i_8_367_1408_0,
    i_8_367_1411_0, i_8_367_1437_0, i_8_367_1439_0, i_8_367_1452_0,
    i_8_367_1464_0, i_8_367_1527_0, i_8_367_1545_0, i_8_367_1546_0,
    i_8_367_1570_0, i_8_367_1573_0, i_8_367_1632_0, i_8_367_1681_0,
    i_8_367_1719_0, i_8_367_1746_0, i_8_367_1758_0, i_8_367_1759_0,
    i_8_367_1867_0, i_8_367_1884_0, i_8_367_1885_0, i_8_367_1887_0,
    i_8_367_1902_0, i_8_367_1948_0, i_8_367_1992_0, i_8_367_1995_0,
    i_8_367_2028_0, i_8_367_2031_0, i_8_367_2056_0, i_8_367_2058_0,
    i_8_367_2077_0, i_8_367_2128_0, i_8_367_2140_0, i_8_367_2156_0,
    i_8_367_2190_0, i_8_367_2215_0, i_8_367_2216_0, i_8_367_2270_0;
  output o_8_367_0_0;
  assign o_8_367_0_0 = ~((~i_8_367_2028_0 & ((~i_8_367_97_0 & ((~i_8_367_723_0 & ~i_8_367_874_0 & ~i_8_367_1050_0 & ~i_8_367_1545_0 & ~i_8_367_1573_0 & ~i_8_367_2031_0) | (~i_8_367_120_0 & ~i_8_367_264_0 & i_8_367_598_0 & ~i_8_367_715_0 & ~i_8_367_1408_0 & ~i_8_367_1464_0 & ~i_8_367_2216_0))) | (~i_8_367_291_0 & ~i_8_367_1746_0 & ((~i_8_367_233_0 & ~i_8_367_282_0 & ~i_8_367_439_0 & ~i_8_367_601_0 & ~i_8_367_723_0 & ~i_8_367_995_0 & ~i_8_367_1061_0 & ~i_8_367_1464_0) | (~i_8_367_51_0 & ~i_8_367_264_0 & ~i_8_367_1389_0 & i_8_367_1948_0 & ~i_8_367_2215_0))) | (~i_8_367_672_0 & ((~i_8_367_480_0 & ~i_8_367_701_0 & ~i_8_367_1237_0 & ~i_8_367_1354_0 & ~i_8_367_1390_0 & ~i_8_367_1545_0 & ~i_8_367_1885_0) | (~i_8_367_256_0 & ~i_8_367_328_0 & ~i_8_367_450_0 & ~i_8_367_874_0 & i_8_367_1632_0 & ~i_8_367_2270_0))))) | (~i_8_367_282_0 & ((~i_8_367_120_0 & ~i_8_367_330_0 & ~i_8_367_439_0 & ~i_8_367_601_0 & ~i_8_367_786_0 & ~i_8_367_1273_0 & ~i_8_367_1452_0) | (~i_8_367_51_0 & ~i_8_367_246_0 & ~i_8_367_264_0 & ~i_8_367_291_0 & ~i_8_367_598_0 & ~i_8_367_1182_0 & ~i_8_367_1902_0 & i_8_367_2140_0))) | (~i_8_367_723_0 & ((~i_8_367_246_0 & ((~i_8_367_786_0 & ~i_8_367_874_0 & ~i_8_367_1273_0 & ~i_8_367_1573_0 & ~i_8_367_2031_0 & ~i_8_367_1390_0 & ~i_8_367_1439_0) | (~i_8_367_292_0 & ~i_8_367_601_0 & ~i_8_367_672_0 & ~i_8_367_1995_0 & ~i_8_367_2190_0))) | (~i_8_367_439_0 & ((~i_8_367_120_0 & ~i_8_367_966_0 & ~i_8_367_995_0 & i_8_367_1050_0 & ~i_8_367_1074_0 & ~i_8_367_1867_0 & ~i_8_367_2031_0) | (~i_8_367_51_0 & ~i_8_367_321_0 & ~i_8_367_456_0 & i_8_367_480_0 & ~i_8_367_672_0 & ~i_8_367_969_0 & ~i_8_367_1545_0 & ~i_8_367_2216_0))) | (~i_8_367_598_0 & ~i_8_367_601_0 & i_8_367_1885_0))) | (~i_8_367_51_0 & ~i_8_367_455_0 & ((~i_8_367_480_0 & i_8_367_601_0 & ~i_8_367_612_0 & ~i_8_367_1050_0 & ~i_8_367_1390_0 & ~i_8_367_1437_0 & ~i_8_367_1546_0) | (~i_8_367_120_0 & ~i_8_367_291_0 & ~i_8_367_328_0 & i_8_367_1884_0 & ~i_8_367_2031_0))) | (~i_8_367_120_0 & ~i_8_367_1902_0 & ((~i_8_367_437_0 & ~i_8_367_1074_0 & ~i_8_367_1273_0 & ~i_8_367_1545_0 & ~i_8_367_1546_0 & i_8_367_1681_0) | (~i_8_367_346_0 & ~i_8_367_439_0 & ~i_8_367_450_0 & ~i_8_367_822_0 & ~i_8_367_969_0 & ~i_8_367_995_0 & ~i_8_367_1527_0 & ~i_8_367_2056_0 & ~i_8_367_2140_0))) | (~i_8_367_2031_0 & ((~i_8_367_321_0 & ~i_8_367_437_0 & ~i_8_367_439_0 & ~i_8_367_715_0 & ~i_8_367_786_0 & ~i_8_367_1182_0 & ~i_8_367_1390_0) | (~i_8_367_163_0 & ~i_8_367_291_0 & ~i_8_367_480_0 & ~i_8_367_672_0 & ~i_8_367_826_0 & ~i_8_367_1234_0 & ~i_8_367_1452_0 & ~i_8_367_1546_0 & ~i_8_367_1573_0))) | (~i_8_367_601_0 & i_8_367_1237_0 & i_8_367_1354_0 & i_8_367_1948_0));
endmodule



// Benchmark "kernel_8_368" written by ABC on Sun Jul 19 10:09:28 2020

module kernel_8_368 ( 
    i_8_368_13_0, i_8_368_50_0, i_8_368_139_0, i_8_368_170_0,
    i_8_368_188_0, i_8_368_192_0, i_8_368_226_0, i_8_368_229_0,
    i_8_368_257_0, i_8_368_263_0, i_8_368_277_0, i_8_368_278_0,
    i_8_368_283_0, i_8_368_365_0, i_8_368_383_0, i_8_368_385_0,
    i_8_368_425_0, i_8_368_449_0, i_8_368_454_0, i_8_368_457_0,
    i_8_368_490_0, i_8_368_493_0, i_8_368_526_0, i_8_368_528_0,
    i_8_368_530_0, i_8_368_544_0, i_8_368_606_0, i_8_368_613_0,
    i_8_368_617_0, i_8_368_631_0, i_8_368_632_0, i_8_368_655_0,
    i_8_368_656_0, i_8_368_661_0, i_8_368_703_0, i_8_368_709_0,
    i_8_368_710_0, i_8_368_785_0, i_8_368_798_0, i_8_368_854_0,
    i_8_368_866_0, i_8_368_892_0, i_8_368_935_0, i_8_368_977_0,
    i_8_368_1019_0, i_8_368_1023_0, i_8_368_1060_0, i_8_368_1075_0,
    i_8_368_1103_0, i_8_368_1163_0, i_8_368_1174_0, i_8_368_1228_0,
    i_8_368_1280_0, i_8_368_1282_0, i_8_368_1307_0, i_8_368_1334_0,
    i_8_368_1379_0, i_8_368_1414_0, i_8_368_1424_0, i_8_368_1471_0,
    i_8_368_1538_0, i_8_368_1558_0, i_8_368_1610_0, i_8_368_1642_0,
    i_8_368_1655_0, i_8_368_1685_0, i_8_368_1705_0, i_8_368_1750_0,
    i_8_368_1811_0, i_8_368_1849_0, i_8_368_1910_0, i_8_368_1913_0,
    i_8_368_1946_0, i_8_368_1952_0, i_8_368_1964_0, i_8_368_1973_0,
    i_8_368_1978_0, i_8_368_1982_0, i_8_368_1997_0, i_8_368_2006_0,
    i_8_368_2009_0, i_8_368_2038_0, i_8_368_2039_0, i_8_368_2091_0,
    i_8_368_2095_0, i_8_368_2126_0, i_8_368_2144_0, i_8_368_2146_0,
    i_8_368_2164_0, i_8_368_2168_0, i_8_368_2171_0, i_8_368_2173_0,
    i_8_368_2183_0, i_8_368_2186_0, i_8_368_2228_0, i_8_368_2239_0,
    i_8_368_2249_0, i_8_368_2259_0, i_8_368_2268_0, i_8_368_2293_0,
    o_8_368_0_0  );
  input  i_8_368_13_0, i_8_368_50_0, i_8_368_139_0, i_8_368_170_0,
    i_8_368_188_0, i_8_368_192_0, i_8_368_226_0, i_8_368_229_0,
    i_8_368_257_0, i_8_368_263_0, i_8_368_277_0, i_8_368_278_0,
    i_8_368_283_0, i_8_368_365_0, i_8_368_383_0, i_8_368_385_0,
    i_8_368_425_0, i_8_368_449_0, i_8_368_454_0, i_8_368_457_0,
    i_8_368_490_0, i_8_368_493_0, i_8_368_526_0, i_8_368_528_0,
    i_8_368_530_0, i_8_368_544_0, i_8_368_606_0, i_8_368_613_0,
    i_8_368_617_0, i_8_368_631_0, i_8_368_632_0, i_8_368_655_0,
    i_8_368_656_0, i_8_368_661_0, i_8_368_703_0, i_8_368_709_0,
    i_8_368_710_0, i_8_368_785_0, i_8_368_798_0, i_8_368_854_0,
    i_8_368_866_0, i_8_368_892_0, i_8_368_935_0, i_8_368_977_0,
    i_8_368_1019_0, i_8_368_1023_0, i_8_368_1060_0, i_8_368_1075_0,
    i_8_368_1103_0, i_8_368_1163_0, i_8_368_1174_0, i_8_368_1228_0,
    i_8_368_1280_0, i_8_368_1282_0, i_8_368_1307_0, i_8_368_1334_0,
    i_8_368_1379_0, i_8_368_1414_0, i_8_368_1424_0, i_8_368_1471_0,
    i_8_368_1538_0, i_8_368_1558_0, i_8_368_1610_0, i_8_368_1642_0,
    i_8_368_1655_0, i_8_368_1685_0, i_8_368_1705_0, i_8_368_1750_0,
    i_8_368_1811_0, i_8_368_1849_0, i_8_368_1910_0, i_8_368_1913_0,
    i_8_368_1946_0, i_8_368_1952_0, i_8_368_1964_0, i_8_368_1973_0,
    i_8_368_1978_0, i_8_368_1982_0, i_8_368_1997_0, i_8_368_2006_0,
    i_8_368_2009_0, i_8_368_2038_0, i_8_368_2039_0, i_8_368_2091_0,
    i_8_368_2095_0, i_8_368_2126_0, i_8_368_2144_0, i_8_368_2146_0,
    i_8_368_2164_0, i_8_368_2168_0, i_8_368_2171_0, i_8_368_2173_0,
    i_8_368_2183_0, i_8_368_2186_0, i_8_368_2228_0, i_8_368_2239_0,
    i_8_368_2249_0, i_8_368_2259_0, i_8_368_2268_0, i_8_368_2293_0;
  output o_8_368_0_0;
  assign o_8_368_0_0 = 0;
endmodule



// Benchmark "kernel_8_369" written by ABC on Sun Jul 19 10:09:30 2020

module kernel_8_369 ( 
    i_8_369_37_0, i_8_369_52_0, i_8_369_80_0, i_8_369_89_0, i_8_369_130_0,
    i_8_369_139_0, i_8_369_166_0, i_8_369_192_0, i_8_369_304_0,
    i_8_369_325_0, i_8_369_356_0, i_8_369_367_0, i_8_369_368_0,
    i_8_369_464_0, i_8_369_483_0, i_8_369_486_0, i_8_369_487_0,
    i_8_369_489_0, i_8_369_517_0, i_8_369_518_0, i_8_369_526_0,
    i_8_369_527_0, i_8_369_595_0, i_8_369_608_0, i_8_369_613_0,
    i_8_369_621_0, i_8_369_696_0, i_8_369_699_0, i_8_369_705_0,
    i_8_369_748_0, i_8_369_750_0, i_8_369_757_0, i_8_369_760_0,
    i_8_369_761_0, i_8_369_829_0, i_8_369_840_0, i_8_369_841_0,
    i_8_369_869_0, i_8_369_967_0, i_8_369_981_0, i_8_369_982_0,
    i_8_369_990_0, i_8_369_1074_0, i_8_369_1075_0, i_8_369_1076_0,
    i_8_369_1084_0, i_8_369_1128_0, i_8_369_1224_0, i_8_369_1234_0,
    i_8_369_1264_0, i_8_369_1265_0, i_8_369_1268_0, i_8_369_1273_0,
    i_8_369_1282_0, i_8_369_1305_0, i_8_369_1327_0, i_8_369_1331_0,
    i_8_369_1358_0, i_8_369_1408_0, i_8_369_1476_0, i_8_369_1481_0,
    i_8_369_1498_0, i_8_369_1499_0, i_8_369_1548_0, i_8_369_1557_0,
    i_8_369_1579_0, i_8_369_1613_0, i_8_369_1642_0, i_8_369_1648_0,
    i_8_369_1670_0, i_8_369_1710_0, i_8_369_1729_0, i_8_369_1746_0,
    i_8_369_1748_0, i_8_369_1753_0, i_8_369_1754_0, i_8_369_1779_0,
    i_8_369_1783_0, i_8_369_1787_0, i_8_369_1795_0, i_8_369_1800_0,
    i_8_369_1821_0, i_8_369_1858_0, i_8_369_1867_0, i_8_369_1877_0,
    i_8_369_1900_0, i_8_369_1999_0, i_8_369_2003_0, i_8_369_2008_0,
    i_8_369_2026_0, i_8_369_2047_0, i_8_369_2080_0, i_8_369_2154_0,
    i_8_369_2170_0, i_8_369_2174_0, i_8_369_2215_0, i_8_369_2216_0,
    i_8_369_2246_0, i_8_369_2253_0, i_8_369_2260_0,
    o_8_369_0_0  );
  input  i_8_369_37_0, i_8_369_52_0, i_8_369_80_0, i_8_369_89_0,
    i_8_369_130_0, i_8_369_139_0, i_8_369_166_0, i_8_369_192_0,
    i_8_369_304_0, i_8_369_325_0, i_8_369_356_0, i_8_369_367_0,
    i_8_369_368_0, i_8_369_464_0, i_8_369_483_0, i_8_369_486_0,
    i_8_369_487_0, i_8_369_489_0, i_8_369_517_0, i_8_369_518_0,
    i_8_369_526_0, i_8_369_527_0, i_8_369_595_0, i_8_369_608_0,
    i_8_369_613_0, i_8_369_621_0, i_8_369_696_0, i_8_369_699_0,
    i_8_369_705_0, i_8_369_748_0, i_8_369_750_0, i_8_369_757_0,
    i_8_369_760_0, i_8_369_761_0, i_8_369_829_0, i_8_369_840_0,
    i_8_369_841_0, i_8_369_869_0, i_8_369_967_0, i_8_369_981_0,
    i_8_369_982_0, i_8_369_990_0, i_8_369_1074_0, i_8_369_1075_0,
    i_8_369_1076_0, i_8_369_1084_0, i_8_369_1128_0, i_8_369_1224_0,
    i_8_369_1234_0, i_8_369_1264_0, i_8_369_1265_0, i_8_369_1268_0,
    i_8_369_1273_0, i_8_369_1282_0, i_8_369_1305_0, i_8_369_1327_0,
    i_8_369_1331_0, i_8_369_1358_0, i_8_369_1408_0, i_8_369_1476_0,
    i_8_369_1481_0, i_8_369_1498_0, i_8_369_1499_0, i_8_369_1548_0,
    i_8_369_1557_0, i_8_369_1579_0, i_8_369_1613_0, i_8_369_1642_0,
    i_8_369_1648_0, i_8_369_1670_0, i_8_369_1710_0, i_8_369_1729_0,
    i_8_369_1746_0, i_8_369_1748_0, i_8_369_1753_0, i_8_369_1754_0,
    i_8_369_1779_0, i_8_369_1783_0, i_8_369_1787_0, i_8_369_1795_0,
    i_8_369_1800_0, i_8_369_1821_0, i_8_369_1858_0, i_8_369_1867_0,
    i_8_369_1877_0, i_8_369_1900_0, i_8_369_1999_0, i_8_369_2003_0,
    i_8_369_2008_0, i_8_369_2026_0, i_8_369_2047_0, i_8_369_2080_0,
    i_8_369_2154_0, i_8_369_2170_0, i_8_369_2174_0, i_8_369_2215_0,
    i_8_369_2216_0, i_8_369_2246_0, i_8_369_2253_0, i_8_369_2260_0;
  output o_8_369_0_0;
  assign o_8_369_0_0 = ~((~i_8_369_2003_0 & ((~i_8_369_37_0 & ~i_8_369_1795_0 & ((~i_8_369_80_0 & ~i_8_369_705_0 & ~i_8_369_1224_0 & ~i_8_369_1557_0 & ~i_8_369_1729_0 & ~i_8_369_1821_0 & i_8_369_1858_0 & ~i_8_369_2080_0) | (~i_8_369_139_0 & ~i_8_369_518_0 & ~i_8_369_750_0 & ~i_8_369_761_0 & ~i_8_369_981_0 & ~i_8_369_982_0 & i_8_369_1264_0 & ~i_8_369_1481_0 & ~i_8_369_1779_0 & ~i_8_369_2008_0 & ~i_8_369_2215_0))) | (~i_8_369_518_0 & ((~i_8_369_52_0 & ~i_8_369_517_0 & ~i_8_369_829_0 & ~i_8_369_869_0 & ~i_8_369_1476_0 & ~i_8_369_1729_0 & ~i_8_369_1746_0 & ~i_8_369_2047_0 & ~i_8_369_2170_0 & ~i_8_369_2216_0) | (~i_8_369_304_0 & ~i_8_369_757_0 & ~i_8_369_967_0 & ~i_8_369_1265_0 & ~i_8_369_1498_0 & ~i_8_369_1710_0 & ~i_8_369_2008_0 & ~i_8_369_2026_0 & ~i_8_369_2253_0))) | (~i_8_369_608_0 & ((i_8_369_367_0 & ~i_8_369_464_0 & ~i_8_369_1076_0 & ~i_8_369_1858_0 & ~i_8_369_2008_0) | (~i_8_369_483_0 & ~i_8_369_829_0 & ~i_8_369_1498_0 & ~i_8_369_1499_0 & ~i_8_369_1783_0 & ~i_8_369_1999_0 & i_8_369_2215_0))) | (~i_8_369_981_0 & ((~i_8_369_517_0 & ((i_8_369_526_0 & ~i_8_369_705_0 & ~i_8_369_829_0 & ~i_8_369_967_0 & ~i_8_369_982_0 & ~i_8_369_1084_0 & ~i_8_369_1331_0 & ~i_8_369_1481_0 & ~i_8_369_1499_0 & ~i_8_369_1900_0 & ~i_8_369_1999_0) | (i_8_369_841_0 & ~i_8_369_1779_0 & ~i_8_369_2008_0 & ~i_8_369_2080_0))) | (~i_8_369_89_0 & ~i_8_369_487_0 & ~i_8_369_982_0 & ~i_8_369_1128_0 & ~i_8_369_1408_0 & ~i_8_369_1481_0 & i_8_369_1748_0 & ~i_8_369_1858_0 & ~i_8_369_1999_0))) | (~i_8_369_1265_0 & ~i_8_369_1282_0 & ~i_8_369_1746_0 & i_8_369_1753_0 & i_8_369_1754_0 & ~i_8_369_2047_0) | (~i_8_369_356_0 & ~i_8_369_517_0 & i_8_369_760_0 & ~i_8_369_2080_0 & i_8_369_2170_0 & ~i_8_369_2253_0))) | (~i_8_369_2080_0 & ((~i_8_369_325_0 & ~i_8_369_621_0 & ((~i_8_369_464_0 & ~i_8_369_1268_0 & i_8_369_1273_0 & ~i_8_369_1476_0 & ~i_8_369_1613_0 & ~i_8_369_1710_0) | (~i_8_369_356_0 & ~i_8_369_517_0 & ~i_8_369_518_0 & ~i_8_369_526_0 & ~i_8_369_981_0 & ~i_8_369_1076_0 & ~i_8_369_1900_0 & ~i_8_369_2008_0))) | (~i_8_369_518_0 & ~i_8_369_990_0 & ((~i_8_369_517_0 & ~i_8_369_982_0 & i_8_369_1224_0) | (~i_8_369_139_0 & i_8_369_748_0 & ~i_8_369_1084_0 & ~i_8_369_1481_0 & ~i_8_369_1900_0 & ~i_8_369_1999_0))) | (~i_8_369_517_0 & ~i_8_369_1476_0 & ((~i_8_369_192_0 & ~i_8_369_304_0 & ~i_8_369_613_0 & ~i_8_369_757_0 & ~i_8_369_760_0 & ~i_8_369_982_0 & ~i_8_369_1076_0 & ~i_8_369_1795_0 & ~i_8_369_1999_0) | (~i_8_369_89_0 & ~i_8_369_761_0 & ~i_8_369_1670_0 & ~i_8_369_2008_0 & i_8_369_2170_0))) | (~i_8_369_613_0 & ~i_8_369_967_0 & ~i_8_369_1999_0 & ((~i_8_369_841_0 & i_8_369_1265_0 & ~i_8_369_1795_0 & ~i_8_369_2253_0) | (~i_8_369_464_0 & ~i_8_369_981_0 & ~i_8_369_1613_0 & ~i_8_369_1710_0 & i_8_369_1753_0 & ~i_8_369_2174_0 & ~i_8_369_2260_0))) | (i_8_369_367_0 & ~i_8_369_760_0 & ~i_8_369_761_0 & ~i_8_369_869_0 & ~i_8_369_1557_0 & ~i_8_369_1746_0 & ~i_8_369_1783_0 & ~i_8_369_2047_0 & ~i_8_369_2246_0))) | (~i_8_369_1999_0 & ((~i_8_369_89_0 & ~i_8_369_757_0 & ((~i_8_369_621_0 & ~i_8_369_760_0 & ~i_8_369_982_0 & ~i_8_369_1075_0 & ~i_8_369_1498_0 & i_8_369_1783_0) | (~i_8_369_52_0 & ~i_8_369_192_0 & ~i_8_369_304_0 & ~i_8_369_1729_0 & ~i_8_369_2008_0 & i_8_369_2174_0 & ~i_8_369_2215_0))) | (~i_8_369_517_0 & ~i_8_369_982_0 & ((~i_8_369_356_0 & ~i_8_369_489_0 & i_8_369_1282_0 & ~i_8_369_1331_0 & ~i_8_369_1476_0 & ~i_8_369_1498_0 & ~i_8_369_1613_0 & ~i_8_369_1900_0) | (~i_8_369_192_0 & ~i_8_369_464_0 & ~i_8_369_696_0 & ~i_8_369_750_0 & ~i_8_369_841_0 & ~i_8_369_869_0 & ~i_8_369_1265_0 & ~i_8_369_1729_0 & ~i_8_369_2008_0 & ~i_8_369_2170_0 & ~i_8_369_2246_0 & ~i_8_369_2253_0))) | (~i_8_369_696_0 & i_8_369_750_0 & ~i_8_369_1327_0 & ~i_8_369_1476_0 & ~i_8_369_2026_0 & ~i_8_369_2047_0))) | (~i_8_369_139_0 & ((~i_8_369_829_0 & ~i_8_369_967_0 & ~i_8_369_1481_0 & ~i_8_369_1499_0 & i_8_369_1754_0 & ~i_8_369_2047_0) | (~i_8_369_487_0 & ~i_8_369_1268_0 & ~i_8_369_1498_0 & ~i_8_369_1858_0 & i_8_369_2246_0 & ~i_8_369_2253_0))) | (~i_8_369_304_0 & ((~i_8_369_613_0 & i_8_369_1265_0 & i_8_369_1358_0 & ~i_8_369_1642_0 & ~i_8_369_2170_0) | (~i_8_369_517_0 & ~i_8_369_608_0 & ~i_8_369_757_0 & ~i_8_369_982_0 & ~i_8_369_1084_0 & i_8_369_1282_0 & ~i_8_369_1648_0 & ~i_8_369_2216_0))) | (i_8_369_368_0 & ~i_8_369_2170_0 & ((~i_8_369_356_0 & ~i_8_369_483_0 & ~i_8_369_518_0 & ~i_8_369_760_0) | (i_8_369_80_0 & ~i_8_369_748_0 & ~i_8_369_829_0 & ~i_8_369_1084_0 & ~i_8_369_1548_0 & ~i_8_369_1779_0 & ~i_8_369_1783_0 & ~i_8_369_2246_0))) | (i_8_369_608_0 & ((~i_8_369_527_0 & i_8_369_757_0 & ~i_8_369_760_0 & ~i_8_369_1476_0 & ~i_8_369_2026_0) | (~i_8_369_192_0 & ~i_8_369_518_0 & ~i_8_369_705_0 & ~i_8_369_1084_0 & ~i_8_369_1234_0 & ~i_8_369_1710_0 & ~i_8_369_1877_0 & i_8_369_2215_0))) | (~i_8_369_518_0 & ((~i_8_369_621_0 & ~i_8_369_760_0 & ~i_8_369_981_0 & ~i_8_369_982_0 & ~i_8_369_1746_0 & i_8_369_1821_0) | (i_8_369_487_0 & ~i_8_369_517_0 & ~i_8_369_526_0 & ~i_8_369_748_0 & ~i_8_369_757_0 & ~i_8_369_1476_0 & ~i_8_369_1481_0 & ~i_8_369_2008_0))) | (i_8_369_517_0 & ~i_8_369_1074_0 & i_8_369_1264_0 & i_8_369_1800_0 & ~i_8_369_2026_0 & i_8_369_2154_0) | (i_8_369_699_0 & ~i_8_369_761_0 & ~i_8_369_1476_0 & ~i_8_369_1548_0 & ~i_8_369_2246_0));
endmodule



// Benchmark "kernel_8_370" written by ABC on Sun Jul 19 10:09:31 2020

module kernel_8_370 ( 
    i_8_370_4_0, i_8_370_18_0, i_8_370_20_0, i_8_370_35_0, i_8_370_40_0,
    i_8_370_41_0, i_8_370_88_0, i_8_370_114_0, i_8_370_115_0,
    i_8_370_166_0, i_8_370_184_0, i_8_370_275_0, i_8_370_307_0,
    i_8_370_319_0, i_8_370_320_0, i_8_370_335_0, i_8_370_343_0,
    i_8_370_364_0, i_8_370_418_0, i_8_370_419_0, i_8_370_427_0,
    i_8_370_453_0, i_8_370_454_0, i_8_370_508_0, i_8_370_526_0,
    i_8_370_554_0, i_8_370_572_0, i_8_370_590_0, i_8_370_599_0,
    i_8_370_613_0, i_8_370_614_0, i_8_370_635_0, i_8_370_638_0,
    i_8_370_640_0, i_8_370_671_0, i_8_370_695_0, i_8_370_769_0,
    i_8_370_882_0, i_8_370_893_0, i_8_370_991_0, i_8_370_1033_0,
    i_8_370_1040_0, i_8_370_1061_0, i_8_370_1084_0, i_8_370_1112_0,
    i_8_370_1115_0, i_8_370_1129_0, i_8_370_1130_0, i_8_370_1174_0,
    i_8_370_1226_0, i_8_370_1229_0, i_8_370_1240_0, i_8_370_1270_0,
    i_8_370_1298_0, i_8_370_1300_0, i_8_370_1396_0, i_8_370_1397_0,
    i_8_370_1408_0, i_8_370_1481_0, i_8_370_1498_0, i_8_370_1526_0,
    i_8_370_1532_0, i_8_370_1544_0, i_8_370_1546_0, i_8_370_1552_0,
    i_8_370_1630_0, i_8_370_1640_0, i_8_370_1642_0, i_8_370_1648_0,
    i_8_370_1651_0, i_8_370_1661_0, i_8_370_1663_0, i_8_370_1693_0,
    i_8_370_1694_0, i_8_370_1705_0, i_8_370_1707_0, i_8_370_1750_0,
    i_8_370_1754_0, i_8_370_1779_0, i_8_370_1807_0, i_8_370_1858_0,
    i_8_370_1883_0, i_8_370_1885_0, i_8_370_1886_0, i_8_370_1949_0,
    i_8_370_1966_0, i_8_370_1968_0, i_8_370_2000_0, i_8_370_2054_0,
    i_8_370_2093_0, i_8_370_2094_0, i_8_370_2135_0, i_8_370_2139_0,
    i_8_370_2140_0, i_8_370_2170_0, i_8_370_2171_0, i_8_370_2192_0,
    i_8_370_2233_0, i_8_370_2257_0, i_8_370_2258_0,
    o_8_370_0_0  );
  input  i_8_370_4_0, i_8_370_18_0, i_8_370_20_0, i_8_370_35_0,
    i_8_370_40_0, i_8_370_41_0, i_8_370_88_0, i_8_370_114_0, i_8_370_115_0,
    i_8_370_166_0, i_8_370_184_0, i_8_370_275_0, i_8_370_307_0,
    i_8_370_319_0, i_8_370_320_0, i_8_370_335_0, i_8_370_343_0,
    i_8_370_364_0, i_8_370_418_0, i_8_370_419_0, i_8_370_427_0,
    i_8_370_453_0, i_8_370_454_0, i_8_370_508_0, i_8_370_526_0,
    i_8_370_554_0, i_8_370_572_0, i_8_370_590_0, i_8_370_599_0,
    i_8_370_613_0, i_8_370_614_0, i_8_370_635_0, i_8_370_638_0,
    i_8_370_640_0, i_8_370_671_0, i_8_370_695_0, i_8_370_769_0,
    i_8_370_882_0, i_8_370_893_0, i_8_370_991_0, i_8_370_1033_0,
    i_8_370_1040_0, i_8_370_1061_0, i_8_370_1084_0, i_8_370_1112_0,
    i_8_370_1115_0, i_8_370_1129_0, i_8_370_1130_0, i_8_370_1174_0,
    i_8_370_1226_0, i_8_370_1229_0, i_8_370_1240_0, i_8_370_1270_0,
    i_8_370_1298_0, i_8_370_1300_0, i_8_370_1396_0, i_8_370_1397_0,
    i_8_370_1408_0, i_8_370_1481_0, i_8_370_1498_0, i_8_370_1526_0,
    i_8_370_1532_0, i_8_370_1544_0, i_8_370_1546_0, i_8_370_1552_0,
    i_8_370_1630_0, i_8_370_1640_0, i_8_370_1642_0, i_8_370_1648_0,
    i_8_370_1651_0, i_8_370_1661_0, i_8_370_1663_0, i_8_370_1693_0,
    i_8_370_1694_0, i_8_370_1705_0, i_8_370_1707_0, i_8_370_1750_0,
    i_8_370_1754_0, i_8_370_1779_0, i_8_370_1807_0, i_8_370_1858_0,
    i_8_370_1883_0, i_8_370_1885_0, i_8_370_1886_0, i_8_370_1949_0,
    i_8_370_1966_0, i_8_370_1968_0, i_8_370_2000_0, i_8_370_2054_0,
    i_8_370_2093_0, i_8_370_2094_0, i_8_370_2135_0, i_8_370_2139_0,
    i_8_370_2140_0, i_8_370_2170_0, i_8_370_2171_0, i_8_370_2192_0,
    i_8_370_2233_0, i_8_370_2257_0, i_8_370_2258_0;
  output o_8_370_0_0;
  assign o_8_370_0_0 = 0;
endmodule



// Benchmark "kernel_8_371" written by ABC on Sun Jul 19 10:09:32 2020

module kernel_8_371 ( 
    i_8_371_14_0, i_8_371_60_0, i_8_371_61_0, i_8_371_76_0, i_8_371_140_0,
    i_8_371_188_0, i_8_371_263_0, i_8_371_341_0, i_8_371_362_0,
    i_8_371_422_0, i_8_371_457_0, i_8_371_491_0, i_8_371_494_0,
    i_8_371_512_0, i_8_371_523_0, i_8_371_575_0, i_8_371_607_0,
    i_8_371_610_0, i_8_371_633_0, i_8_371_652_0, i_8_371_700_0,
    i_8_371_709_0, i_8_371_719_0, i_8_371_736_0, i_8_371_773_0,
    i_8_371_781_0, i_8_371_787_0, i_8_371_788_0, i_8_371_863_0,
    i_8_371_871_0, i_8_371_912_0, i_8_371_998_0, i_8_371_1075_0,
    i_8_371_1106_0, i_8_371_1111_0, i_8_371_1112_0, i_8_371_1114_0,
    i_8_371_1115_0, i_8_371_1157_0, i_8_371_1202_0, i_8_371_1204_0,
    i_8_371_1229_0, i_8_371_1231_0, i_8_371_1240_0, i_8_371_1247_0,
    i_8_371_1263_0, i_8_371_1300_0, i_8_371_1319_0, i_8_371_1322_0,
    i_8_371_1329_0, i_8_371_1331_0, i_8_371_1334_0, i_8_371_1397_0,
    i_8_371_1401_0, i_8_371_1402_0, i_8_371_1403_0, i_8_371_1435_0,
    i_8_371_1439_0, i_8_371_1445_0, i_8_371_1466_0, i_8_371_1490_0,
    i_8_371_1528_0, i_8_371_1552_0, i_8_371_1555_0, i_8_371_1597_0,
    i_8_371_1640_0, i_8_371_1645_0, i_8_371_1667_0, i_8_371_1679_0,
    i_8_371_1703_0, i_8_371_1717_0, i_8_371_1724_0, i_8_371_1748_0,
    i_8_371_1751_0, i_8_371_1762_0, i_8_371_1771_0, i_8_371_1778_0,
    i_8_371_1787_0, i_8_371_1808_0, i_8_371_1825_0, i_8_371_1835_0,
    i_8_371_1841_0, i_8_371_1848_0, i_8_371_1884_0, i_8_371_1888_0,
    i_8_371_1895_0, i_8_371_1948_0, i_8_371_1952_0, i_8_371_1966_0,
    i_8_371_1992_0, i_8_371_2012_0, i_8_371_2138_0, i_8_371_2140_0,
    i_8_371_2144_0, i_8_371_2147_0, i_8_371_2236_0, i_8_371_2237_0,
    i_8_371_2249_0, i_8_371_2264_0, i_8_371_2290_0,
    o_8_371_0_0  );
  input  i_8_371_14_0, i_8_371_60_0, i_8_371_61_0, i_8_371_76_0,
    i_8_371_140_0, i_8_371_188_0, i_8_371_263_0, i_8_371_341_0,
    i_8_371_362_0, i_8_371_422_0, i_8_371_457_0, i_8_371_491_0,
    i_8_371_494_0, i_8_371_512_0, i_8_371_523_0, i_8_371_575_0,
    i_8_371_607_0, i_8_371_610_0, i_8_371_633_0, i_8_371_652_0,
    i_8_371_700_0, i_8_371_709_0, i_8_371_719_0, i_8_371_736_0,
    i_8_371_773_0, i_8_371_781_0, i_8_371_787_0, i_8_371_788_0,
    i_8_371_863_0, i_8_371_871_0, i_8_371_912_0, i_8_371_998_0,
    i_8_371_1075_0, i_8_371_1106_0, i_8_371_1111_0, i_8_371_1112_0,
    i_8_371_1114_0, i_8_371_1115_0, i_8_371_1157_0, i_8_371_1202_0,
    i_8_371_1204_0, i_8_371_1229_0, i_8_371_1231_0, i_8_371_1240_0,
    i_8_371_1247_0, i_8_371_1263_0, i_8_371_1300_0, i_8_371_1319_0,
    i_8_371_1322_0, i_8_371_1329_0, i_8_371_1331_0, i_8_371_1334_0,
    i_8_371_1397_0, i_8_371_1401_0, i_8_371_1402_0, i_8_371_1403_0,
    i_8_371_1435_0, i_8_371_1439_0, i_8_371_1445_0, i_8_371_1466_0,
    i_8_371_1490_0, i_8_371_1528_0, i_8_371_1552_0, i_8_371_1555_0,
    i_8_371_1597_0, i_8_371_1640_0, i_8_371_1645_0, i_8_371_1667_0,
    i_8_371_1679_0, i_8_371_1703_0, i_8_371_1717_0, i_8_371_1724_0,
    i_8_371_1748_0, i_8_371_1751_0, i_8_371_1762_0, i_8_371_1771_0,
    i_8_371_1778_0, i_8_371_1787_0, i_8_371_1808_0, i_8_371_1825_0,
    i_8_371_1835_0, i_8_371_1841_0, i_8_371_1848_0, i_8_371_1884_0,
    i_8_371_1888_0, i_8_371_1895_0, i_8_371_1948_0, i_8_371_1952_0,
    i_8_371_1966_0, i_8_371_1992_0, i_8_371_2012_0, i_8_371_2138_0,
    i_8_371_2140_0, i_8_371_2144_0, i_8_371_2147_0, i_8_371_2236_0,
    i_8_371_2237_0, i_8_371_2249_0, i_8_371_2264_0, i_8_371_2290_0;
  output o_8_371_0_0;
  assign o_8_371_0_0 = 0;
endmodule



// Benchmark "kernel_8_372" written by ABC on Sun Jul 19 10:09:32 2020

module kernel_8_372 ( 
    i_8_372_34_0, i_8_372_88_0, i_8_372_96_0, i_8_372_143_0, i_8_372_258_0,
    i_8_372_330_0, i_8_372_331_0, i_8_372_332_0, i_8_372_349_0,
    i_8_372_363_0, i_8_372_366_0, i_8_372_385_0, i_8_372_448_0,
    i_8_372_449_0, i_8_372_466_0, i_8_372_485_0, i_8_372_502_0,
    i_8_372_522_0, i_8_372_523_0, i_8_372_524_0, i_8_372_527_0,
    i_8_372_553_0, i_8_372_556_0, i_8_372_557_0, i_8_372_599_0,
    i_8_372_601_0, i_8_372_663_0, i_8_372_871_0, i_8_372_898_0,
    i_8_372_926_0, i_8_372_988_0, i_8_372_989_0, i_8_372_993_0,
    i_8_372_994_0, i_8_372_996_0, i_8_372_1015_0, i_8_372_1016_0,
    i_8_372_1032_0, i_8_372_1069_0, i_8_372_1074_0, i_8_372_1087_0,
    i_8_372_1088_0, i_8_372_1112_0, i_8_372_1120_0, i_8_372_1138_0,
    i_8_372_1140_0, i_8_372_1195_0, i_8_372_1258_0, i_8_372_1264_0,
    i_8_372_1265_0, i_8_372_1282_0, i_8_372_1286_0, i_8_372_1307_0,
    i_8_372_1309_0, i_8_372_1456_0, i_8_372_1528_0, i_8_372_1536_0,
    i_8_372_1543_0, i_8_372_1552_0, i_8_372_1555_0, i_8_372_1556_0,
    i_8_372_1574_0, i_8_372_1610_0, i_8_372_1617_0, i_8_372_1628_0,
    i_8_372_1635_0, i_8_372_1636_0, i_8_372_1637_0, i_8_372_1651_0,
    i_8_372_1652_0, i_8_372_1671_0, i_8_372_1672_0, i_8_372_1673_0,
    i_8_372_1679_0, i_8_372_1699_0, i_8_372_1700_0, i_8_372_1704_0,
    i_8_372_1717_0, i_8_372_1735_0, i_8_372_1736_0, i_8_372_1750_0,
    i_8_372_1809_0, i_8_372_1810_0, i_8_372_1858_0, i_8_372_1861_0,
    i_8_372_1905_0, i_8_372_1906_0, i_8_372_1933_0, i_8_372_1934_0,
    i_8_372_1992_0, i_8_372_1994_0, i_8_372_1995_0, i_8_372_2005_0,
    i_8_372_2006_0, i_8_372_2015_0, i_8_372_2114_0, i_8_372_2146_0,
    i_8_372_2215_0, i_8_372_2266_0, i_8_372_2267_0,
    o_8_372_0_0  );
  input  i_8_372_34_0, i_8_372_88_0, i_8_372_96_0, i_8_372_143_0,
    i_8_372_258_0, i_8_372_330_0, i_8_372_331_0, i_8_372_332_0,
    i_8_372_349_0, i_8_372_363_0, i_8_372_366_0, i_8_372_385_0,
    i_8_372_448_0, i_8_372_449_0, i_8_372_466_0, i_8_372_485_0,
    i_8_372_502_0, i_8_372_522_0, i_8_372_523_0, i_8_372_524_0,
    i_8_372_527_0, i_8_372_553_0, i_8_372_556_0, i_8_372_557_0,
    i_8_372_599_0, i_8_372_601_0, i_8_372_663_0, i_8_372_871_0,
    i_8_372_898_0, i_8_372_926_0, i_8_372_988_0, i_8_372_989_0,
    i_8_372_993_0, i_8_372_994_0, i_8_372_996_0, i_8_372_1015_0,
    i_8_372_1016_0, i_8_372_1032_0, i_8_372_1069_0, i_8_372_1074_0,
    i_8_372_1087_0, i_8_372_1088_0, i_8_372_1112_0, i_8_372_1120_0,
    i_8_372_1138_0, i_8_372_1140_0, i_8_372_1195_0, i_8_372_1258_0,
    i_8_372_1264_0, i_8_372_1265_0, i_8_372_1282_0, i_8_372_1286_0,
    i_8_372_1307_0, i_8_372_1309_0, i_8_372_1456_0, i_8_372_1528_0,
    i_8_372_1536_0, i_8_372_1543_0, i_8_372_1552_0, i_8_372_1555_0,
    i_8_372_1556_0, i_8_372_1574_0, i_8_372_1610_0, i_8_372_1617_0,
    i_8_372_1628_0, i_8_372_1635_0, i_8_372_1636_0, i_8_372_1637_0,
    i_8_372_1651_0, i_8_372_1652_0, i_8_372_1671_0, i_8_372_1672_0,
    i_8_372_1673_0, i_8_372_1679_0, i_8_372_1699_0, i_8_372_1700_0,
    i_8_372_1704_0, i_8_372_1717_0, i_8_372_1735_0, i_8_372_1736_0,
    i_8_372_1750_0, i_8_372_1809_0, i_8_372_1810_0, i_8_372_1858_0,
    i_8_372_1861_0, i_8_372_1905_0, i_8_372_1906_0, i_8_372_1933_0,
    i_8_372_1934_0, i_8_372_1992_0, i_8_372_1994_0, i_8_372_1995_0,
    i_8_372_2005_0, i_8_372_2006_0, i_8_372_2015_0, i_8_372_2114_0,
    i_8_372_2146_0, i_8_372_2215_0, i_8_372_2266_0, i_8_372_2267_0;
  output o_8_372_0_0;
  assign o_8_372_0_0 = 0;
endmodule



// Benchmark "kernel_8_373" written by ABC on Sun Jul 19 10:09:34 2020

module kernel_8_373 ( 
    i_8_373_0_0, i_8_373_1_0, i_8_373_31_0, i_8_373_81_0, i_8_373_82_0,
    i_8_373_83_0, i_8_373_84_0, i_8_373_102_0, i_8_373_111_0,
    i_8_373_184_0, i_8_373_203_0, i_8_373_244_0, i_8_373_259_0,
    i_8_373_280_0, i_8_373_306_0, i_8_373_307_0, i_8_373_342_0,
    i_8_373_343_0, i_8_373_346_0, i_8_373_349_0, i_8_373_350_0,
    i_8_373_360_0, i_8_373_388_0, i_8_373_423_0, i_8_373_424_0,
    i_8_373_450_0, i_8_373_460_0, i_8_373_599_0, i_8_373_603_0,
    i_8_373_630_0, i_8_373_632_0, i_8_373_634_0, i_8_373_661_0,
    i_8_373_702_0, i_8_373_706_0, i_8_373_710_0, i_8_373_711_0,
    i_8_373_712_0, i_8_373_756_0, i_8_373_757_0, i_8_373_758_0,
    i_8_373_779_0, i_8_373_780_0, i_8_373_811_0, i_8_373_838_0,
    i_8_373_858_0, i_8_373_993_0, i_8_373_996_0, i_8_373_1035_0,
    i_8_373_1078_0, i_8_373_1093_0, i_8_373_1098_0, i_8_373_1099_0,
    i_8_373_1100_0, i_8_373_1101_0, i_8_373_1103_0, i_8_373_1110_0,
    i_8_373_1115_0, i_8_373_1260_0, i_8_373_1266_0, i_8_373_1314_0,
    i_8_373_1328_0, i_8_373_1331_0, i_8_373_1388_0, i_8_373_1438_0,
    i_8_373_1507_0, i_8_373_1516_0, i_8_373_1532_0, i_8_373_1533_0,
    i_8_373_1642_0, i_8_373_1678_0, i_8_373_1679_0, i_8_373_1683_0,
    i_8_373_1684_0, i_8_373_1685_0, i_8_373_1759_0, i_8_373_1763_0,
    i_8_373_1779_0, i_8_373_1804_0, i_8_373_1805_0, i_8_373_1826_0,
    i_8_373_1935_0, i_8_373_1936_0, i_8_373_1937_0, i_8_373_1938_0,
    i_8_373_1939_0, i_8_373_1964_0, i_8_373_1969_0, i_8_373_2026_0,
    i_8_373_2115_0, i_8_373_2116_0, i_8_373_2117_0, i_8_373_2136_0,
    i_8_373_2137_0, i_8_373_2138_0, i_8_373_2229_0, i_8_373_2245_0,
    i_8_373_2248_0, i_8_373_2260_0, i_8_373_2270_0,
    o_8_373_0_0  );
  input  i_8_373_0_0, i_8_373_1_0, i_8_373_31_0, i_8_373_81_0,
    i_8_373_82_0, i_8_373_83_0, i_8_373_84_0, i_8_373_102_0, i_8_373_111_0,
    i_8_373_184_0, i_8_373_203_0, i_8_373_244_0, i_8_373_259_0,
    i_8_373_280_0, i_8_373_306_0, i_8_373_307_0, i_8_373_342_0,
    i_8_373_343_0, i_8_373_346_0, i_8_373_349_0, i_8_373_350_0,
    i_8_373_360_0, i_8_373_388_0, i_8_373_423_0, i_8_373_424_0,
    i_8_373_450_0, i_8_373_460_0, i_8_373_599_0, i_8_373_603_0,
    i_8_373_630_0, i_8_373_632_0, i_8_373_634_0, i_8_373_661_0,
    i_8_373_702_0, i_8_373_706_0, i_8_373_710_0, i_8_373_711_0,
    i_8_373_712_0, i_8_373_756_0, i_8_373_757_0, i_8_373_758_0,
    i_8_373_779_0, i_8_373_780_0, i_8_373_811_0, i_8_373_838_0,
    i_8_373_858_0, i_8_373_993_0, i_8_373_996_0, i_8_373_1035_0,
    i_8_373_1078_0, i_8_373_1093_0, i_8_373_1098_0, i_8_373_1099_0,
    i_8_373_1100_0, i_8_373_1101_0, i_8_373_1103_0, i_8_373_1110_0,
    i_8_373_1115_0, i_8_373_1260_0, i_8_373_1266_0, i_8_373_1314_0,
    i_8_373_1328_0, i_8_373_1331_0, i_8_373_1388_0, i_8_373_1438_0,
    i_8_373_1507_0, i_8_373_1516_0, i_8_373_1532_0, i_8_373_1533_0,
    i_8_373_1642_0, i_8_373_1678_0, i_8_373_1679_0, i_8_373_1683_0,
    i_8_373_1684_0, i_8_373_1685_0, i_8_373_1759_0, i_8_373_1763_0,
    i_8_373_1779_0, i_8_373_1804_0, i_8_373_1805_0, i_8_373_1826_0,
    i_8_373_1935_0, i_8_373_1936_0, i_8_373_1937_0, i_8_373_1938_0,
    i_8_373_1939_0, i_8_373_1964_0, i_8_373_1969_0, i_8_373_2026_0,
    i_8_373_2115_0, i_8_373_2116_0, i_8_373_2117_0, i_8_373_2136_0,
    i_8_373_2137_0, i_8_373_2138_0, i_8_373_2229_0, i_8_373_2245_0,
    i_8_373_2248_0, i_8_373_2260_0, i_8_373_2270_0;
  output o_8_373_0_0;
  assign o_8_373_0_0 = ~((i_8_373_203_0 & ((i_8_373_1759_0 & i_8_373_1804_0 & ~i_8_373_1805_0) | (~i_8_373_1098_0 & ~i_8_373_1103_0 & i_8_373_1805_0 & ~i_8_373_1936_0))) | (~i_8_373_460_0 & ((~i_8_373_1098_0 & ~i_8_373_1100_0 & ~i_8_373_1101_0 & i_8_373_1115_0 & ~i_8_373_1679_0 & i_8_373_2137_0) | (~i_8_373_259_0 & ~i_8_373_423_0 & ~i_8_373_1093_0 & ~i_8_373_1099_0 & i_8_373_1266_0 & ~i_8_373_1678_0 & ~i_8_373_1683_0 & ~i_8_373_1937_0 & ~i_8_373_2260_0))) | (~i_8_373_388_0 & ((~i_8_373_259_0 & ~i_8_373_424_0 & ((~i_8_373_706_0 & i_8_373_711_0 & ~i_8_373_757_0 & ~i_8_373_1098_0 & ~i_8_373_1266_0) | (~i_8_373_84_0 & ~i_8_373_111_0 & ~i_8_373_306_0 & ~i_8_373_307_0 & ~i_8_373_360_0 & ~i_8_373_603_0 & ~i_8_373_630_0 & ~i_8_373_710_0 & ~i_8_373_712_0 & ~i_8_373_996_0 & ~i_8_373_1093_0 & ~i_8_373_1099_0 & ~i_8_373_1100_0 & ~i_8_373_1101_0 & ~i_8_373_1103_0 & ~i_8_373_1685_0 & ~i_8_373_1759_0 & ~i_8_373_1937_0 & ~i_8_373_1969_0 & ~i_8_373_2136_0 & ~i_8_373_2245_0))) | (~i_8_373_711_0 & ((~i_8_373_342_0 & ~i_8_373_780_0 & ~i_8_373_1093_0 & ~i_8_373_1100_0 & i_8_373_1110_0 & ~i_8_373_1266_0 & ~i_8_373_1507_0 & ~i_8_373_1642_0 & ~i_8_373_1804_0 & i_8_373_2245_0) | (~i_8_373_349_0 & i_8_373_706_0 & ~i_8_373_710_0 & ~i_8_373_1516_0 & i_8_373_1805_0 & ~i_8_373_2136_0 & ~i_8_373_2248_0))) | (~i_8_373_306_0 & ~i_8_373_423_0 & i_8_373_779_0 & i_8_373_1115_0 & ~i_8_373_1314_0 & ~i_8_373_1685_0) | (i_8_373_424_0 & ~i_8_373_603_0 & ~i_8_373_706_0 & ~i_8_373_1266_0 & ~i_8_373_1328_0 & ~i_8_373_1516_0 & ~i_8_373_1532_0 & i_8_373_1679_0 & ~i_8_373_1935_0))) | (i_8_373_757_0 & ((i_8_373_1679_0 & ~i_8_373_1826_0) | (~i_8_373_858_0 & ~i_8_373_1101_0 & ~i_8_373_1103_0 & ~i_8_373_1642_0 & ~i_8_373_1683_0 & ~i_8_373_1939_0))) | (i_8_373_858_0 & ((~i_8_373_342_0 & i_8_373_780_0) | (~i_8_373_349_0 & ~i_8_373_1098_0 & ~i_8_373_1507_0 & ~i_8_373_1683_0 & ~i_8_373_1935_0 & ~i_8_373_1939_0 & ~i_8_373_2026_0))) | (i_8_373_780_0 & ((~i_8_373_346_0 & ~i_8_373_1101_0 & ~i_8_373_1103_0 & i_8_373_1759_0) | (~i_8_373_350_0 & ~i_8_373_423_0 & ~i_8_373_838_0 & ~i_8_373_996_0 & ~i_8_373_1099_0 & ~i_8_373_2229_0))) | (~i_8_373_1939_0 & ((~i_8_373_1685_0 & ((i_8_373_350_0 & ((i_8_373_710_0 & ~i_8_373_1099_0 & i_8_373_1115_0 & ~i_8_373_1266_0 & ~i_8_373_1937_0) | (~i_8_373_423_0 & ~i_8_373_1098_0 & i_8_373_1438_0 & i_8_373_1826_0 & ~i_8_373_1969_0))) | (~i_8_373_424_0 & ~i_8_373_996_0 & ~i_8_373_1078_0 & ~i_8_373_1093_0 & ~i_8_373_1103_0 & i_8_373_1759_0 & ~i_8_373_2245_0))) | (~i_8_373_1099_0 & ((~i_8_373_1101_0 & ((~i_8_373_203_0 & ~i_8_373_1098_0 & i_8_373_1115_0 & i_8_373_1331_0 & ~i_8_373_1937_0) | (i_8_373_634_0 & ~i_8_373_1035_0 & i_8_373_2136_0 & i_8_373_2137_0))) | (i_8_373_84_0 & ~i_8_373_634_0 & ~i_8_373_1103_0 & ~i_8_373_1266_0 & ~i_8_373_1507_0 & ~i_8_373_1516_0 & ~i_8_373_1533_0 & ~i_8_373_1684_0 & ~i_8_373_1969_0 & ~i_8_373_2245_0))) | (i_8_373_1804_0 & i_8_373_1826_0 & ((~i_8_373_346_0 & i_8_373_1759_0) | (~i_8_373_111_0 & ~i_8_373_1100_0 & ~i_8_373_1103_0 & ~i_8_373_1516_0 & ~i_8_373_1533_0 & ~i_8_373_1938_0))))) | (~i_8_373_1103_0 & ((~i_8_373_1101_0 & ((~i_8_373_111_0 & ~i_8_373_450_0 & ~i_8_373_1936_0 & ((~i_8_373_346_0 & ~i_8_373_632_0 & ~i_8_373_838_0 & ~i_8_373_1683_0 & i_8_373_2229_0 & ~i_8_373_2245_0) | (~i_8_373_102_0 & ~i_8_373_307_0 & ~i_8_373_343_0 & ~i_8_373_350_0 & ~i_8_373_661_0 & ~i_8_373_706_0 & ~i_8_373_993_0 & ~i_8_373_996_0 & ~i_8_373_1078_0 & ~i_8_373_1098_0 & ~i_8_373_1100_0 & ~i_8_373_1507_0 & ~i_8_373_1685_0 & ~i_8_373_1937_0 & ~i_8_373_1969_0 & ~i_8_373_2260_0))) | (~i_8_373_184_0 & ~i_8_373_1098_0 & ((~i_8_373_259_0 & ~i_8_373_423_0 & ~i_8_373_632_0 & ~i_8_373_1093_0 & ~i_8_373_1100_0 & i_8_373_1438_0 & ~i_8_373_1532_0 & ~i_8_373_1533_0) | (i_8_373_349_0 & i_8_373_350_0 & ~i_8_373_1078_0 & ~i_8_373_1328_0 & ~i_8_373_1685_0 & ~i_8_373_2137_0 & ~i_8_373_2260_0))) | (~i_8_373_259_0 & ~i_8_373_424_0 & ~i_8_373_838_0 & ~i_8_373_1507_0 & ~i_8_373_1684_0 & i_8_373_2245_0))) | (~i_8_373_1804_0 & ((~i_8_373_423_0 & ((~i_8_373_838_0 & ~i_8_373_1093_0 & ~i_8_373_1507_0 & ~i_8_373_1533_0 & i_8_373_1779_0) | (~i_8_373_306_0 & ~i_8_373_350_0 & ~i_8_373_712_0 & ~i_8_373_1678_0 & i_8_373_1826_0 & ~i_8_373_2026_0 & ~i_8_373_2136_0))) | (~i_8_373_342_0 & ~i_8_373_343_0 & ~i_8_373_706_0 & ~i_8_373_996_0 & ~i_8_373_1098_0 & i_8_373_1110_0 & ~i_8_373_1507_0 & ~i_8_373_1533_0 & ~i_8_373_1969_0 & ~i_8_373_2229_0))) | (~i_8_373_702_0 & ((i_8_373_81_0 & ~i_8_373_1098_0 & i_8_373_1110_0 & ~i_8_373_1685_0 & ~i_8_373_1763_0) | (~i_8_373_630_0 & ~i_8_373_1035_0 & ~i_8_373_1093_0 & ~i_8_373_1438_0 & ~i_8_373_1507_0 & ~i_8_373_1935_0 & ~i_8_373_1936_0 & ~i_8_373_1938_0 & i_8_373_2136_0 & ~i_8_373_2260_0 & ~i_8_373_2270_0))) | (~i_8_373_838_0 & ~i_8_373_1093_0 & ((~i_8_373_424_0 & i_8_373_632_0 & ~i_8_373_634_0 & ~i_8_373_779_0 & ~i_8_373_1078_0) | (~i_8_373_1507_0 & ~i_8_373_1684_0 & ~i_8_373_1936_0 & ~i_8_373_1969_0 & i_8_373_2229_0))) | (~i_8_373_1328_0 & ~i_8_373_1969_0 & ((~i_8_373_1100_0 & ~i_8_373_1507_0 & ~i_8_373_1679_0 & i_8_373_1804_0 & i_8_373_1805_0) | (~i_8_373_349_0 & i_8_373_350_0 & i_8_373_710_0 & ~i_8_373_1642_0 & ~i_8_373_1937_0))) | (i_8_373_1388_0 & ~i_8_373_1507_0) | (~i_8_373_346_0 & ~i_8_373_996_0 & i_8_373_1759_0 & i_8_373_1804_0 & i_8_373_1969_0) | (~i_8_373_82_0 & ~i_8_373_280_0 & i_8_373_634_0 & ~i_8_373_1683_0 & ~i_8_373_1684_0 & i_8_373_2248_0))) | (~i_8_373_1684_0 & ((i_8_373_84_0 & ((i_8_373_423_0 & ~i_8_373_450_0 & ~i_8_373_811_0 & ~i_8_373_993_0 & ~i_8_373_1098_0 & ~i_8_373_2026_0) | (~i_8_373_306_0 & ~i_8_373_343_0 & ~i_8_373_706_0 & ~i_8_373_1100_0 & ~i_8_373_1101_0 & ~i_8_373_1260_0 & ~i_8_373_1314_0 & ~i_8_373_1516_0 & ~i_8_373_1683_0 & ~i_8_373_2260_0))) | (~i_8_373_184_0 & ~i_8_373_1093_0 & ~i_8_373_1331_0 & ((~i_8_373_306_0 & ~i_8_373_307_0 & ~i_8_373_343_0 & ~i_8_373_632_0 & ~i_8_373_996_0 & ~i_8_373_1098_0 & ~i_8_373_1101_0 & ~i_8_373_1328_0 & i_8_373_1678_0 & ~i_8_373_1683_0 & ~i_8_373_1685_0 & ~i_8_373_1935_0 & ~i_8_373_1937_0 & ~i_8_373_2026_0) | (i_8_373_710_0 & ~i_8_373_858_0 & ~i_8_373_993_0 & i_8_373_2138_0))) | (~i_8_373_996_0 & ((~i_8_373_0_0 & i_8_373_81_0 & ~i_8_373_342_0 & ~i_8_373_350_0 & ~i_8_373_1683_0 & ~i_8_373_1936_0) | (~i_8_373_346_0 & ~i_8_373_1098_0 & ~i_8_373_1260_0 & i_8_373_1679_0 & ~i_8_373_1685_0 & i_8_373_1804_0 & ~i_8_373_1938_0))) | (~i_8_373_1098_0 & ~i_8_373_1101_0 & ((~i_8_373_702_0 & ~i_8_373_706_0 & ~i_8_373_1516_0 & ~i_8_373_1678_0 & i_8_373_1679_0 & ~i_8_373_1937_0) | (~i_8_373_423_0 & ~i_8_373_424_0 & ~i_8_373_1110_0 & ~i_8_373_1328_0 & i_8_373_1779_0 & ~i_8_373_1826_0 & i_8_373_1969_0))) | (~i_8_373_423_0 & ((~i_8_373_343_0 & ~i_8_373_661_0 & ~i_8_373_706_0 & ~i_8_373_1779_0 & ~i_8_373_1935_0 & ~i_8_373_1969_0 & i_8_373_2136_0) | (~i_8_373_634_0 & ~i_8_373_1100_0 & ~i_8_373_1516_0 & ~i_8_373_1805_0 & i_8_373_1964_0 & ~i_8_373_2260_0))) | (~i_8_373_307_0 & ~i_8_373_632_0 & ~i_8_373_706_0 & ~i_8_373_838_0 & ~i_8_373_1100_0 & ~i_8_373_1507_0 & ~i_8_373_1678_0 & i_8_373_1685_0 & ~i_8_373_1804_0 & ~i_8_373_1805_0))) | (~i_8_373_259_0 & ((i_8_373_81_0 & ((i_8_373_811_0 & ~i_8_373_1683_0) | (~i_8_373_1093_0 & i_8_373_1260_0 & ~i_8_373_2136_0))) | (~i_8_373_349_0 & ~i_8_373_1078_0 & ~i_8_373_1100_0 & ~i_8_373_1110_0 & i_8_373_1115_0 & ~i_8_373_1685_0 & ~i_8_373_1804_0 & ~i_8_373_1826_0))) | (~i_8_373_360_0 & ((~i_8_373_184_0 & ~i_8_373_1100_0 & ((i_8_373_634_0 & ~i_8_373_702_0 & ~i_8_373_996_0 & ~i_8_373_1260_0 & ~i_8_373_1331_0 & ~i_8_373_1935_0 & ~i_8_373_1937_0) | (~i_8_373_343_0 & ~i_8_373_710_0 & ~i_8_373_1438_0 & ~i_8_373_1685_0 & ~i_8_373_1804_0 & ~i_8_373_2026_0 & i_8_373_2137_0 & ~i_8_373_2245_0 & ~i_8_373_2270_0))) | (~i_8_373_450_0 & ((~i_8_373_993_0 & ~i_8_373_996_0 & ~i_8_373_343_0 & ~i_8_373_349_0 & ~i_8_373_1035_0 & ~i_8_373_1078_0 & ~i_8_373_1260_0 & i_8_373_1266_0) | (i_8_373_111_0 & ~i_8_373_702_0 & i_8_373_2026_0))))) | (~i_8_373_424_0 & ((~i_8_373_423_0 & ((i_8_373_630_0 & ~i_8_373_1098_0 & ~i_8_373_1100_0 & ~i_8_373_1533_0) | (~i_8_373_603_0 & ~i_8_373_630_0 & i_8_373_712_0 & ~i_8_373_1078_0 & ~i_8_373_1099_0 & ~i_8_373_1331_0 & ~i_8_373_1935_0 & ~i_8_373_1937_0 & ~i_8_373_2115_0))) | (~i_8_373_661_0 & ((~i_8_373_630_0 & ~i_8_373_706_0 & ~i_8_373_1093_0 & ~i_8_373_1101_0 & i_8_373_1110_0 & ~i_8_373_1260_0 & ~i_8_373_1314_0 & ~i_8_373_2138_0) | (i_8_373_779_0 & ~i_8_373_1098_0 & ~i_8_373_1685_0 & ~i_8_373_1826_0 & ~i_8_373_1937_0 & ~i_8_373_2245_0))))) | (~i_8_373_1100_0 & ((~i_8_373_1093_0 & ((~i_8_373_423_0 & ((~i_8_373_702_0 & ~i_8_373_996_0 & ~i_8_373_349_0 & ~i_8_373_450_0 & ~i_8_373_1099_0 & i_8_373_1533_0 & ~i_8_373_1935_0 & ~i_8_373_2260_0) | (~i_8_373_306_0 & ~i_8_373_346_0 & ~i_8_373_634_0 & ~i_8_373_706_0 & ~i_8_373_1098_0 & ~i_8_373_1110_0 & i_8_373_1678_0 & ~i_8_373_1685_0 & ~i_8_373_2270_0))) | (~i_8_373_996_0 & ~i_8_373_1507_0 & ~i_8_373_1642_0 & i_8_373_1804_0 & i_8_373_1805_0))) | (~i_8_373_1438_0 & i_8_373_1763_0 & i_8_373_1969_0) | (~i_8_373_1314_0 & ~i_8_373_1533_0 & ~i_8_373_1937_0 & i_8_373_2117_0))) | (~i_8_373_993_0 & ((~i_8_373_632_0 & ~i_8_373_1098_0 & i_8_373_1763_0 & i_8_373_1804_0 & ~i_8_373_1938_0) | (~i_8_373_111_0 & ~i_8_373_342_0 & i_8_373_1533_0 & ~i_8_373_1685_0 & i_8_373_1779_0 & ~i_8_373_2260_0))) | (i_8_373_1115_0 & ((~i_8_373_996_0 & i_8_373_1078_0 & ~i_8_373_1093_0 & ~i_8_373_1099_0 & ~i_8_373_1507_0) | (~i_8_373_184_0 & ~i_8_373_599_0 & ~i_8_373_1098_0 & ~i_8_373_1328_0 & i_8_373_1826_0 & ~i_8_373_1937_0 & ~i_8_373_2137_0))) | (i_8_373_82_0 & i_8_373_83_0 & ~i_8_373_661_0 & ~i_8_373_1078_0 & ~i_8_373_1331_0) | (i_8_373_84_0 & i_8_373_102_0 & i_8_373_1759_0) | (i_8_373_758_0 & ~i_8_373_1507_0 & i_8_373_1969_0));
endmodule



// Benchmark "kernel_8_374" written by ABC on Sun Jul 19 10:09:35 2020

module kernel_8_374 ( 
    i_8_374_6_0, i_8_374_7_0, i_8_374_37_0, i_8_374_41_0, i_8_374_64_0,
    i_8_374_111_0, i_8_374_130_0, i_8_374_172_0, i_8_374_178_0,
    i_8_374_263_0, i_8_374_297_0, i_8_374_301_0, i_8_374_307_0,
    i_8_374_316_0, i_8_374_319_0, i_8_374_355_0, i_8_374_356_0,
    i_8_374_361_0, i_8_374_363_0, i_8_374_414_0, i_8_374_424_0,
    i_8_374_447_0, i_8_374_527_0, i_8_374_532_0, i_8_374_568_0,
    i_8_374_612_0, i_8_374_624_0, i_8_374_639_0, i_8_374_661_0,
    i_8_374_664_0, i_8_374_667_0, i_8_374_675_0, i_8_374_682_0,
    i_8_374_684_0, i_8_374_704_0, i_8_374_796_0, i_8_374_837_0,
    i_8_374_838_0, i_8_374_853_0, i_8_374_870_0, i_8_374_874_0,
    i_8_374_975_0, i_8_374_1008_0, i_8_374_1053_0, i_8_374_1099_0,
    i_8_374_1126_0, i_8_374_1145_0, i_8_374_1174_0, i_8_374_1225_0,
    i_8_374_1233_0, i_8_374_1241_0, i_8_374_1285_0, i_8_374_1296_0,
    i_8_374_1297_0, i_8_374_1331_0, i_8_374_1337_0, i_8_374_1350_0,
    i_8_374_1380_0, i_8_374_1383_0, i_8_374_1446_0, i_8_374_1467_0,
    i_8_374_1488_0, i_8_374_1510_0, i_8_374_1522_0, i_8_374_1614_0,
    i_8_374_1631_0, i_8_374_1638_0, i_8_374_1645_0, i_8_374_1705_0,
    i_8_374_1707_0, i_8_374_1750_0, i_8_374_1764_0, i_8_374_1768_0,
    i_8_374_1773_0, i_8_374_1781_0, i_8_374_1809_0, i_8_374_1819_0,
    i_8_374_1855_0, i_8_374_1887_0, i_8_374_1891_0, i_8_374_1929_0,
    i_8_374_1935_0, i_8_374_1948_0, i_8_374_1953_0, i_8_374_2012_0,
    i_8_374_2016_0, i_8_374_2044_0, i_8_374_2053_0, i_8_374_2061_0,
    i_8_374_2071_0, i_8_374_2079_0, i_8_374_2080_0, i_8_374_2134_0,
    i_8_374_2140_0, i_8_374_2167_0, i_8_374_2185_0, i_8_374_2216_0,
    i_8_374_2230_0, i_8_374_2236_0, i_8_374_2284_0,
    o_8_374_0_0  );
  input  i_8_374_6_0, i_8_374_7_0, i_8_374_37_0, i_8_374_41_0,
    i_8_374_64_0, i_8_374_111_0, i_8_374_130_0, i_8_374_172_0,
    i_8_374_178_0, i_8_374_263_0, i_8_374_297_0, i_8_374_301_0,
    i_8_374_307_0, i_8_374_316_0, i_8_374_319_0, i_8_374_355_0,
    i_8_374_356_0, i_8_374_361_0, i_8_374_363_0, i_8_374_414_0,
    i_8_374_424_0, i_8_374_447_0, i_8_374_527_0, i_8_374_532_0,
    i_8_374_568_0, i_8_374_612_0, i_8_374_624_0, i_8_374_639_0,
    i_8_374_661_0, i_8_374_664_0, i_8_374_667_0, i_8_374_675_0,
    i_8_374_682_0, i_8_374_684_0, i_8_374_704_0, i_8_374_796_0,
    i_8_374_837_0, i_8_374_838_0, i_8_374_853_0, i_8_374_870_0,
    i_8_374_874_0, i_8_374_975_0, i_8_374_1008_0, i_8_374_1053_0,
    i_8_374_1099_0, i_8_374_1126_0, i_8_374_1145_0, i_8_374_1174_0,
    i_8_374_1225_0, i_8_374_1233_0, i_8_374_1241_0, i_8_374_1285_0,
    i_8_374_1296_0, i_8_374_1297_0, i_8_374_1331_0, i_8_374_1337_0,
    i_8_374_1350_0, i_8_374_1380_0, i_8_374_1383_0, i_8_374_1446_0,
    i_8_374_1467_0, i_8_374_1488_0, i_8_374_1510_0, i_8_374_1522_0,
    i_8_374_1614_0, i_8_374_1631_0, i_8_374_1638_0, i_8_374_1645_0,
    i_8_374_1705_0, i_8_374_1707_0, i_8_374_1750_0, i_8_374_1764_0,
    i_8_374_1768_0, i_8_374_1773_0, i_8_374_1781_0, i_8_374_1809_0,
    i_8_374_1819_0, i_8_374_1855_0, i_8_374_1887_0, i_8_374_1891_0,
    i_8_374_1929_0, i_8_374_1935_0, i_8_374_1948_0, i_8_374_1953_0,
    i_8_374_2012_0, i_8_374_2016_0, i_8_374_2044_0, i_8_374_2053_0,
    i_8_374_2061_0, i_8_374_2071_0, i_8_374_2079_0, i_8_374_2080_0,
    i_8_374_2134_0, i_8_374_2140_0, i_8_374_2167_0, i_8_374_2185_0,
    i_8_374_2216_0, i_8_374_2230_0, i_8_374_2236_0, i_8_374_2284_0;
  output o_8_374_0_0;
  assign o_8_374_0_0 = 0;
endmodule



// Benchmark "kernel_8_375" written by ABC on Sun Jul 19 10:09:36 2020

module kernel_8_375 ( 
    i_8_375_21_0, i_8_375_45_0, i_8_375_73_0, i_8_375_129_0, i_8_375_130_0,
    i_8_375_147_0, i_8_375_150_0, i_8_375_192_0, i_8_375_193_0,
    i_8_375_222_0, i_8_375_329_0, i_8_375_355_0, i_8_375_378_0,
    i_8_375_385_0, i_8_375_462_0, i_8_375_472_0, i_8_375_493_0,
    i_8_375_516_0, i_8_375_517_0, i_8_375_519_0, i_8_375_525_0,
    i_8_375_549_0, i_8_375_606_0, i_8_375_613_0, i_8_375_624_0,
    i_8_375_631_0, i_8_375_652_0, i_8_375_658_0, i_8_375_659_0,
    i_8_375_661_0, i_8_375_694_0, i_8_375_703_0, i_8_375_705_0,
    i_8_375_715_0, i_8_375_733_0, i_8_375_831_0, i_8_375_832_0,
    i_8_375_876_0, i_8_375_879_0, i_8_375_925_0, i_8_375_963_0,
    i_8_375_1000_0, i_8_375_1003_0, i_8_375_1059_0, i_8_375_1086_0,
    i_8_375_1158_0, i_8_375_1164_0, i_8_375_1192_0, i_8_375_1224_0,
    i_8_375_1266_0, i_8_375_1281_0, i_8_375_1284_0, i_8_375_1302_0,
    i_8_375_1335_0, i_8_375_1336_0, i_8_375_1348_0, i_8_375_1354_0,
    i_8_375_1390_0, i_8_375_1435_0, i_8_375_1438_0, i_8_375_1455_0,
    i_8_375_1464_0, i_8_375_1489_0, i_8_375_1498_0, i_8_375_1539_0,
    i_8_375_1593_0, i_8_375_1596_0, i_8_375_1621_0, i_8_375_1641_0,
    i_8_375_1650_0, i_8_375_1659_0, i_8_375_1660_0, i_8_375_1662_0,
    i_8_375_1696_0, i_8_375_1704_0, i_8_375_1740_0, i_8_375_1743_0,
    i_8_375_1750_0, i_8_375_1875_0, i_8_375_1876_0, i_8_375_1881_0,
    i_8_375_1974_0, i_8_375_2010_0, i_8_375_2011_0, i_8_375_2046_0,
    i_8_375_2047_0, i_8_375_2057_0, i_8_375_2064_0, i_8_375_2092_0,
    i_8_375_2118_0, i_8_375_2146_0, i_8_375_2169_0, i_8_375_2172_0,
    i_8_375_2173_0, i_8_375_2185_0, i_8_375_2209_0, i_8_375_2253_0,
    i_8_375_2254_0, i_8_375_2256_0, i_8_375_2257_0,
    o_8_375_0_0  );
  input  i_8_375_21_0, i_8_375_45_0, i_8_375_73_0, i_8_375_129_0,
    i_8_375_130_0, i_8_375_147_0, i_8_375_150_0, i_8_375_192_0,
    i_8_375_193_0, i_8_375_222_0, i_8_375_329_0, i_8_375_355_0,
    i_8_375_378_0, i_8_375_385_0, i_8_375_462_0, i_8_375_472_0,
    i_8_375_493_0, i_8_375_516_0, i_8_375_517_0, i_8_375_519_0,
    i_8_375_525_0, i_8_375_549_0, i_8_375_606_0, i_8_375_613_0,
    i_8_375_624_0, i_8_375_631_0, i_8_375_652_0, i_8_375_658_0,
    i_8_375_659_0, i_8_375_661_0, i_8_375_694_0, i_8_375_703_0,
    i_8_375_705_0, i_8_375_715_0, i_8_375_733_0, i_8_375_831_0,
    i_8_375_832_0, i_8_375_876_0, i_8_375_879_0, i_8_375_925_0,
    i_8_375_963_0, i_8_375_1000_0, i_8_375_1003_0, i_8_375_1059_0,
    i_8_375_1086_0, i_8_375_1158_0, i_8_375_1164_0, i_8_375_1192_0,
    i_8_375_1224_0, i_8_375_1266_0, i_8_375_1281_0, i_8_375_1284_0,
    i_8_375_1302_0, i_8_375_1335_0, i_8_375_1336_0, i_8_375_1348_0,
    i_8_375_1354_0, i_8_375_1390_0, i_8_375_1435_0, i_8_375_1438_0,
    i_8_375_1455_0, i_8_375_1464_0, i_8_375_1489_0, i_8_375_1498_0,
    i_8_375_1539_0, i_8_375_1593_0, i_8_375_1596_0, i_8_375_1621_0,
    i_8_375_1641_0, i_8_375_1650_0, i_8_375_1659_0, i_8_375_1660_0,
    i_8_375_1662_0, i_8_375_1696_0, i_8_375_1704_0, i_8_375_1740_0,
    i_8_375_1743_0, i_8_375_1750_0, i_8_375_1875_0, i_8_375_1876_0,
    i_8_375_1881_0, i_8_375_1974_0, i_8_375_2010_0, i_8_375_2011_0,
    i_8_375_2046_0, i_8_375_2047_0, i_8_375_2057_0, i_8_375_2064_0,
    i_8_375_2092_0, i_8_375_2118_0, i_8_375_2146_0, i_8_375_2169_0,
    i_8_375_2172_0, i_8_375_2173_0, i_8_375_2185_0, i_8_375_2209_0,
    i_8_375_2253_0, i_8_375_2254_0, i_8_375_2256_0, i_8_375_2257_0;
  output o_8_375_0_0;
  assign o_8_375_0_0 = ~((~i_8_375_192_0 & ((~i_8_375_45_0 & ~i_8_375_516_0 & ~i_8_375_517_0 & ~i_8_375_1086_0 & ~i_8_375_1164_0 & ~i_8_375_1539_0) | (~i_8_375_1659_0 & ~i_8_375_2092_0 & ~i_8_375_2257_0))) | (~i_8_375_516_0 & ((~i_8_375_150_0 & ~i_8_375_525_0 & ~i_8_375_624_0 & ~i_8_375_2011_0 & ~i_8_375_2118_0) | (~i_8_375_715_0 & ~i_8_375_1539_0 & ~i_8_375_1662_0 & i_8_375_1750_0 & ~i_8_375_2256_0))) | (~i_8_375_832_0 & ((~i_8_375_21_0 & i_8_375_525_0 & ~i_8_375_606_0 & ~i_8_375_1335_0 & ~i_8_375_1650_0 & ~i_8_375_1704_0) | (~i_8_375_147_0 & ~i_8_375_831_0 & ~i_8_375_1158_0 & ~i_8_375_1660_0 & ~i_8_375_2256_0))) | (~i_8_375_147_0 & ((~i_8_375_1266_0 & ((~i_8_375_378_0 & ~i_8_375_879_0 & ~i_8_375_1621_0 & ~i_8_375_1650_0) | (i_8_375_493_0 & ~i_8_375_549_0 & i_8_375_705_0 & ~i_8_375_1348_0 & ~i_8_375_1539_0 & ~i_8_375_1875_0 & ~i_8_375_2057_0))) | (~i_8_375_1348_0 & ~i_8_375_1641_0 & ~i_8_375_2169_0 & ~i_8_375_2209_0 & ~i_8_375_2253_0))) | (~i_8_375_2011_0 & ~i_8_375_2118_0 & ((~i_8_375_658_0 & ~i_8_375_733_0 & ~i_8_375_1335_0 & ~i_8_375_1455_0 & ~i_8_375_1539_0 & ~i_8_375_2046_0 & ~i_8_375_2209_0) | (~i_8_375_193_0 & ~i_8_375_385_0 & ~i_8_375_694_0 & ~i_8_375_1498_0 & ~i_8_375_2256_0))) | (~i_8_375_130_0 & i_8_375_694_0 & ~i_8_375_1000_0 & ~i_8_375_1164_0 & ~i_8_375_1593_0) | (~i_8_375_659_0 & ~i_8_375_703_0 & ~i_8_375_1059_0 & ~i_8_375_1224_0 & ~i_8_375_1662_0 & ~i_8_375_1876_0 & ~i_8_375_1881_0) | (~i_8_375_517_0 & ~i_8_375_705_0 & ~i_8_375_2010_0 & ~i_8_375_2173_0));
endmodule



// Benchmark "kernel_8_376" written by ABC on Sun Jul 19 10:09:37 2020

module kernel_8_376 ( 
    i_8_376_11_0, i_8_376_27_0, i_8_376_32_0, i_8_376_51_0, i_8_376_97_0,
    i_8_376_141_0, i_8_376_142_0, i_8_376_169_0, i_8_376_223_0,
    i_8_376_224_0, i_8_376_230_0, i_8_376_259_0, i_8_376_260_0,
    i_8_376_346_0, i_8_376_372_0, i_8_376_418_0, i_8_376_440_0,
    i_8_376_480_0, i_8_376_501_0, i_8_376_505_0, i_8_376_507_0,
    i_8_376_523_0, i_8_376_524_0, i_8_376_555_0, i_8_376_556_0,
    i_8_376_591_0, i_8_376_598_0, i_8_376_602_0, i_8_376_617_0,
    i_8_376_649_0, i_8_376_687_0, i_8_376_692_0, i_8_376_702_0,
    i_8_376_705_0, i_8_376_750_0, i_8_376_760_0, i_8_376_762_0,
    i_8_376_763_0, i_8_376_838_0, i_8_376_843_0, i_8_376_844_0,
    i_8_376_850_0, i_8_376_886_0, i_8_376_958_0, i_8_376_969_0,
    i_8_376_994_0, i_8_376_1032_0, i_8_376_1051_0, i_8_376_1074_0,
    i_8_376_1075_0, i_8_376_1077_0, i_8_376_1094_0, i_8_376_1096_0,
    i_8_376_1123_0, i_8_376_1124_0, i_8_376_1191_0, i_8_376_1222_0,
    i_8_376_1282_0, i_8_376_1285_0, i_8_376_1305_0, i_8_376_1306_0,
    i_8_376_1316_0, i_8_376_1318_0, i_8_376_1330_0, i_8_376_1331_0,
    i_8_376_1386_0, i_8_376_1387_0, i_8_376_1390_0, i_8_376_1410_0,
    i_8_376_1411_0, i_8_376_1470_0, i_8_376_1471_0, i_8_376_1507_0,
    i_8_376_1509_0, i_8_376_1533_0, i_8_376_1548_0, i_8_376_1560_0,
    i_8_376_1564_0, i_8_376_1573_0, i_8_376_1574_0, i_8_376_1635_0,
    i_8_376_1655_0, i_8_376_1680_0, i_8_376_1681_0, i_8_376_1682_0,
    i_8_376_1704_0, i_8_376_1722_0, i_8_376_1723_0, i_8_376_1821_0,
    i_8_376_1834_0, i_8_376_1858_0, i_8_376_1906_0, i_8_376_2032_0,
    i_8_376_2119_0, i_8_376_2122_0, i_8_376_2145_0, i_8_376_2211_0,
    i_8_376_2214_0, i_8_376_2215_0, i_8_376_2216_0,
    o_8_376_0_0  );
  input  i_8_376_11_0, i_8_376_27_0, i_8_376_32_0, i_8_376_51_0,
    i_8_376_97_0, i_8_376_141_0, i_8_376_142_0, i_8_376_169_0,
    i_8_376_223_0, i_8_376_224_0, i_8_376_230_0, i_8_376_259_0,
    i_8_376_260_0, i_8_376_346_0, i_8_376_372_0, i_8_376_418_0,
    i_8_376_440_0, i_8_376_480_0, i_8_376_501_0, i_8_376_505_0,
    i_8_376_507_0, i_8_376_523_0, i_8_376_524_0, i_8_376_555_0,
    i_8_376_556_0, i_8_376_591_0, i_8_376_598_0, i_8_376_602_0,
    i_8_376_617_0, i_8_376_649_0, i_8_376_687_0, i_8_376_692_0,
    i_8_376_702_0, i_8_376_705_0, i_8_376_750_0, i_8_376_760_0,
    i_8_376_762_0, i_8_376_763_0, i_8_376_838_0, i_8_376_843_0,
    i_8_376_844_0, i_8_376_850_0, i_8_376_886_0, i_8_376_958_0,
    i_8_376_969_0, i_8_376_994_0, i_8_376_1032_0, i_8_376_1051_0,
    i_8_376_1074_0, i_8_376_1075_0, i_8_376_1077_0, i_8_376_1094_0,
    i_8_376_1096_0, i_8_376_1123_0, i_8_376_1124_0, i_8_376_1191_0,
    i_8_376_1222_0, i_8_376_1282_0, i_8_376_1285_0, i_8_376_1305_0,
    i_8_376_1306_0, i_8_376_1316_0, i_8_376_1318_0, i_8_376_1330_0,
    i_8_376_1331_0, i_8_376_1386_0, i_8_376_1387_0, i_8_376_1390_0,
    i_8_376_1410_0, i_8_376_1411_0, i_8_376_1470_0, i_8_376_1471_0,
    i_8_376_1507_0, i_8_376_1509_0, i_8_376_1533_0, i_8_376_1548_0,
    i_8_376_1560_0, i_8_376_1564_0, i_8_376_1573_0, i_8_376_1574_0,
    i_8_376_1635_0, i_8_376_1655_0, i_8_376_1680_0, i_8_376_1681_0,
    i_8_376_1682_0, i_8_376_1704_0, i_8_376_1722_0, i_8_376_1723_0,
    i_8_376_1821_0, i_8_376_1834_0, i_8_376_1858_0, i_8_376_1906_0,
    i_8_376_2032_0, i_8_376_2119_0, i_8_376_2122_0, i_8_376_2145_0,
    i_8_376_2211_0, i_8_376_2214_0, i_8_376_2215_0, i_8_376_2216_0;
  output o_8_376_0_0;
  assign o_8_376_0_0 = 0;
endmodule



// Benchmark "kernel_8_377" written by ABC on Sun Jul 19 10:09:39 2020

module kernel_8_377 ( 
    i_8_377_3_0, i_8_377_6_0, i_8_377_7_0, i_8_377_19_0, i_8_377_36_0,
    i_8_377_84_0, i_8_377_87_0, i_8_377_184_0, i_8_377_193_0,
    i_8_377_230_0, i_8_377_246_0, i_8_377_247_0, i_8_377_249_0,
    i_8_377_250_0, i_8_377_347_0, i_8_377_350_0, i_8_377_360_0,
    i_8_377_361_0, i_8_377_427_0, i_8_377_430_0, i_8_377_439_0,
    i_8_377_499_0, i_8_377_518_0, i_8_377_525_0, i_8_377_528_0,
    i_8_377_571_0, i_8_377_573_0, i_8_377_597_0, i_8_377_601_0,
    i_8_377_606_0, i_8_377_607_0, i_8_377_608_0, i_8_377_654_0,
    i_8_377_661_0, i_8_377_669_0, i_8_377_672_0, i_8_377_685_0,
    i_8_377_703_0, i_8_377_706_0, i_8_377_717_0, i_8_377_718_0,
    i_8_377_726_0, i_8_377_762_0, i_8_377_777_0, i_8_377_813_0,
    i_8_377_814_0, i_8_377_816_0, i_8_377_817_0, i_8_377_831_0,
    i_8_377_832_0, i_8_377_838_0, i_8_377_1071_0, i_8_377_1074_0,
    i_8_377_1084_0, i_8_377_1155_0, i_8_377_1159_0, i_8_377_1192_0,
    i_8_377_1285_0, i_8_377_1291_0, i_8_377_1295_0, i_8_377_1389_0,
    i_8_377_1392_0, i_8_377_1434_0, i_8_377_1497_0, i_8_377_1498_0,
    i_8_377_1542_0, i_8_377_1573_0, i_8_377_1658_0, i_8_377_1696_0,
    i_8_377_1749_0, i_8_377_1763_0, i_8_377_1819_0, i_8_377_1830_0,
    i_8_377_1833_0, i_8_377_1848_0, i_8_377_1851_0, i_8_377_1852_0,
    i_8_377_1866_0, i_8_377_1915_0, i_8_377_1938_0, i_8_377_1946_0,
    i_8_377_1947_0, i_8_377_1963_0, i_8_377_1974_0, i_8_377_1984_0,
    i_8_377_1985_0, i_8_377_2028_0, i_8_377_2031_0, i_8_377_2037_0,
    i_8_377_2047_0, i_8_377_2056_0, i_8_377_2064_0, i_8_377_2073_0,
    i_8_377_2076_0, i_8_377_2091_0, i_8_377_2095_0, i_8_377_2113_0,
    i_8_377_2118_0, i_8_377_2246_0, i_8_377_2281_0,
    o_8_377_0_0  );
  input  i_8_377_3_0, i_8_377_6_0, i_8_377_7_0, i_8_377_19_0,
    i_8_377_36_0, i_8_377_84_0, i_8_377_87_0, i_8_377_184_0, i_8_377_193_0,
    i_8_377_230_0, i_8_377_246_0, i_8_377_247_0, i_8_377_249_0,
    i_8_377_250_0, i_8_377_347_0, i_8_377_350_0, i_8_377_360_0,
    i_8_377_361_0, i_8_377_427_0, i_8_377_430_0, i_8_377_439_0,
    i_8_377_499_0, i_8_377_518_0, i_8_377_525_0, i_8_377_528_0,
    i_8_377_571_0, i_8_377_573_0, i_8_377_597_0, i_8_377_601_0,
    i_8_377_606_0, i_8_377_607_0, i_8_377_608_0, i_8_377_654_0,
    i_8_377_661_0, i_8_377_669_0, i_8_377_672_0, i_8_377_685_0,
    i_8_377_703_0, i_8_377_706_0, i_8_377_717_0, i_8_377_718_0,
    i_8_377_726_0, i_8_377_762_0, i_8_377_777_0, i_8_377_813_0,
    i_8_377_814_0, i_8_377_816_0, i_8_377_817_0, i_8_377_831_0,
    i_8_377_832_0, i_8_377_838_0, i_8_377_1071_0, i_8_377_1074_0,
    i_8_377_1084_0, i_8_377_1155_0, i_8_377_1159_0, i_8_377_1192_0,
    i_8_377_1285_0, i_8_377_1291_0, i_8_377_1295_0, i_8_377_1389_0,
    i_8_377_1392_0, i_8_377_1434_0, i_8_377_1497_0, i_8_377_1498_0,
    i_8_377_1542_0, i_8_377_1573_0, i_8_377_1658_0, i_8_377_1696_0,
    i_8_377_1749_0, i_8_377_1763_0, i_8_377_1819_0, i_8_377_1830_0,
    i_8_377_1833_0, i_8_377_1848_0, i_8_377_1851_0, i_8_377_1852_0,
    i_8_377_1866_0, i_8_377_1915_0, i_8_377_1938_0, i_8_377_1946_0,
    i_8_377_1947_0, i_8_377_1963_0, i_8_377_1974_0, i_8_377_1984_0,
    i_8_377_1985_0, i_8_377_2028_0, i_8_377_2031_0, i_8_377_2037_0,
    i_8_377_2047_0, i_8_377_2056_0, i_8_377_2064_0, i_8_377_2073_0,
    i_8_377_2076_0, i_8_377_2091_0, i_8_377_2095_0, i_8_377_2113_0,
    i_8_377_2118_0, i_8_377_2246_0, i_8_377_2281_0;
  output o_8_377_0_0;
  assign o_8_377_0_0 = ~((~i_8_377_1498_0 & ((~i_8_377_1389_0 & ((~i_8_377_3_0 & ~i_8_377_87_0 & ((~i_8_377_6_0 & ~i_8_377_246_0 & ~i_8_377_250_0 & ~i_8_377_597_0 & ~i_8_377_814_0 & i_8_377_838_0 & ~i_8_377_1573_0 & ~i_8_377_1749_0 & ~i_8_377_1833_0 & ~i_8_377_1851_0) | (~i_8_377_36_0 & ~i_8_377_230_0 & ~i_8_377_247_0 & ~i_8_377_717_0 & ~i_8_377_831_0 & ~i_8_377_1392_0 & i_8_377_1749_0 & ~i_8_377_1866_0 & ~i_8_377_2047_0))) | (~i_8_377_193_0 & ~i_8_377_246_0 & ~i_8_377_601_0 & ~i_8_377_817_0 & ~i_8_377_1392_0 & ((~i_8_377_84_0 & ~i_8_377_499_0 & ~i_8_377_718_0 & ~i_8_377_777_0 & ~i_8_377_1963_0 & ~i_8_377_2031_0 & ~i_8_377_2064_0) | (~i_8_377_247_0 & ~i_8_377_525_0 & ~i_8_377_597_0 & ~i_8_377_717_0 & ~i_8_377_832_0 & ~i_8_377_1573_0 & ~i_8_377_2047_0 & ~i_8_377_2118_0))))) | (~i_8_377_1392_0 & ((~i_8_377_832_0 & ((~i_8_377_817_0 & ((~i_8_377_84_0 & ~i_8_377_525_0 & ~i_8_377_2028_0 & ((~i_8_377_249_0 & ~i_8_377_439_0 & ~i_8_377_499_0 & ~i_8_377_1573_0 & i_8_377_2095_0) | (~i_8_377_19_0 & ~i_8_377_250_0 & ~i_8_377_654_0 & ~i_8_377_717_0 & ~i_8_377_718_0 & ~i_8_377_816_0 & ~i_8_377_831_0 & ~i_8_377_1084_0 & ~i_8_377_1749_0 & ~i_8_377_1866_0 & ~i_8_377_2031_0 & ~i_8_377_2037_0 & ~i_8_377_2095_0))) | (~i_8_377_193_0 & ~i_8_377_246_0 & ~i_8_377_439_0 & ~i_8_377_601_0 & ~i_8_377_669_0 & ~i_8_377_672_0 & ~i_8_377_838_0 & ~i_8_377_1192_0 & ~i_8_377_1763_0 & ~i_8_377_1852_0 & ~i_8_377_2037_0 & ~i_8_377_2047_0 & ~i_8_377_2118_0 & ~i_8_377_2246_0))) | (~i_8_377_6_0 & i_8_377_84_0 & ~i_8_377_246_0 & ~i_8_377_571_0 & ~i_8_377_762_0 & ~i_8_377_814_0 & ~i_8_377_816_0 & ~i_8_377_831_0 & ~i_8_377_1074_0 & ~i_8_377_1084_0 & ~i_8_377_1573_0 & ~i_8_377_1947_0))) | (~i_8_377_814_0 & ((i_8_377_606_0 & ~i_8_377_813_0 & ~i_8_377_1159_0 & i_8_377_1434_0 & ~i_8_377_1658_0) | (~i_8_377_250_0 & ~i_8_377_597_0 & ~i_8_377_661_0 & ~i_8_377_669_0 & i_8_377_718_0 & ~i_8_377_1573_0 & ~i_8_377_2037_0 & ~i_8_377_2091_0 & ~i_8_377_2095_0 & ~i_8_377_2281_0))))) | (~i_8_377_2281_0 & ((~i_8_377_246_0 & ~i_8_377_718_0 & i_8_377_777_0 & i_8_377_838_0 & ~i_8_377_2028_0) | (~i_8_377_661_0 & ~i_8_377_669_0 & ~i_8_377_1071_0 & ~i_8_377_1749_0 & i_8_377_1819_0 & ~i_8_377_1866_0 & ~i_8_377_1947_0 & ~i_8_377_2047_0))))) | (~i_8_377_7_0 & ((~i_8_377_84_0 & ~i_8_377_250_0 & i_8_377_361_0 & ~i_8_377_718_0 & ~i_8_377_814_0 & ~i_8_377_1830_0 & ~i_8_377_1946_0) | (~i_8_377_87_0 & ~i_8_377_247_0 & i_8_377_430_0 & ~i_8_377_525_0 & ~i_8_377_672_0 & ~i_8_377_717_0 & ~i_8_377_817_0 & ~i_8_377_831_0 & ~i_8_377_2028_0))) | (~i_8_377_2095_0 & ((~i_8_377_19_0 & ((~i_8_377_87_0 & ~i_8_377_230_0 & ~i_8_377_249_0 & ~i_8_377_601_0 & ~i_8_377_654_0 & i_8_377_661_0 & ~i_8_377_762_0 & ~i_8_377_816_0 & ~i_8_377_817_0 & ~i_8_377_1542_0 & ~i_8_377_1848_0 & ~i_8_377_1851_0 & ~i_8_377_1915_0 & ~i_8_377_1963_0 & ~i_8_377_2064_0) | (i_8_377_230_0 & ~i_8_377_718_0 & ~i_8_377_1071_0 & ~i_8_377_1159_0 & ~i_8_377_1573_0 & ~i_8_377_2091_0 & ~i_8_377_2113_0 & ~i_8_377_2118_0 & ~i_8_377_2281_0))) | (~i_8_377_499_0 & ~i_8_377_718_0 & ~i_8_377_832_0 & ((~i_8_377_528_0 & ~i_8_377_816_0 & ~i_8_377_1851_0 & ~i_8_377_2028_0 & i_8_377_2246_0) | (~i_8_377_250_0 & ~i_8_377_518_0 & ~i_8_377_601_0 & ~i_8_377_669_0 & ~i_8_377_1071_0 & ~i_8_377_1392_0 & ~i_8_377_1542_0 & ~i_8_377_1749_0 & ~i_8_377_1852_0 & ~i_8_377_1915_0 & ~i_8_377_2091_0 & ~i_8_377_2246_0))) | (~i_8_377_3_0 & i_8_377_427_0 & ~i_8_377_518_0 & ~i_8_377_528_0 & ~i_8_377_717_0 & ~i_8_377_762_0 & ~i_8_377_1497_0 & ~i_8_377_1866_0 & ~i_8_377_2064_0 & ~i_8_377_2091_0))) | (~i_8_377_1392_0 & ((~i_8_377_2064_0 & ((~i_8_377_87_0 & ~i_8_377_2047_0 & ((~i_8_377_246_0 & ~i_8_377_249_0 & ~i_8_377_528_0 & ~i_8_377_601_0 & ~i_8_377_669_0 & ~i_8_377_718_0 & ~i_8_377_814_0 & ~i_8_377_817_0 & ~i_8_377_1071_0 & ~i_8_377_1497_0 & ~i_8_377_1866_0 & ~i_8_377_2028_0) | (~i_8_377_250_0 & i_8_377_777_0 & ~i_8_377_813_0 & ~i_8_377_1285_0 & ~i_8_377_1295_0 & ~i_8_377_1389_0 & ~i_8_377_2037_0))) | (~i_8_377_84_0 & ~i_8_377_193_0 & ~i_8_377_246_0 & ~i_8_377_247_0 & i_8_377_525_0 & ~i_8_377_717_0 & ~i_8_377_718_0 & ~i_8_377_762_0 & ~i_8_377_1389_0 & ~i_8_377_1658_0 & ~i_8_377_2028_0))) | (~i_8_377_2031_0 & ((~i_8_377_350_0 & ~i_8_377_1295_0 & ~i_8_377_2091_0 & ((i_8_377_525_0 & ~i_8_377_717_0 & ~i_8_377_1071_0 & ~i_8_377_1084_0 & ~i_8_377_1573_0 & ~i_8_377_1848_0 & i_8_377_1947_0) | (~i_8_377_193_0 & ~i_8_377_518_0 & ~i_8_377_597_0 & ~i_8_377_601_0 & ~i_8_377_703_0 & ~i_8_377_1389_0 & i_8_377_2095_0 & ~i_8_377_2113_0))) | (~i_8_377_249_0 & i_8_377_350_0 & i_8_377_430_0 & ~i_8_377_685_0 & ~i_8_377_2118_0 & ~i_8_377_2281_0))))) | (~i_8_377_250_0 & ((i_8_377_525_0 & i_8_377_607_0 & ~i_8_377_817_0 & ~i_8_377_1074_0 & ~i_8_377_1084_0 & ~i_8_377_1573_0 & ~i_8_377_1696_0 & ~i_8_377_2064_0) | (~i_8_377_814_0 & i_8_377_1155_0 & ~i_8_377_1389_0 & ~i_8_377_2031_0 & i_8_377_2073_0))) | (~i_8_377_601_0 & ((~i_8_377_247_0 & ~i_8_377_427_0 & ~i_8_377_661_0 & ~i_8_377_813_0 & ~i_8_377_831_0 & i_8_377_838_0 & ~i_8_377_2047_0) | (i_8_377_193_0 & ~i_8_377_430_0 & ~i_8_377_669_0 & ~i_8_377_703_0 & ~i_8_377_717_0 & ~i_8_377_1497_0 & ~i_8_377_1542_0 & ~i_8_377_1851_0 & ~i_8_377_1947_0 & i_8_377_2091_0))) | (~i_8_377_1852_0 & ((~i_8_377_247_0 & ((~i_8_377_36_0 & ~i_8_377_246_0 & i_8_377_706_0 & ~i_8_377_718_0 & ~i_8_377_814_0 & ~i_8_377_1285_0 & ~i_8_377_1389_0 & ~i_8_377_1658_0 & ~i_8_377_2031_0) | (i_8_377_347_0 & ~i_8_377_669_0 & ~i_8_377_762_0 & ~i_8_377_813_0 & ~i_8_377_817_0 & ~i_8_377_1159_0 & ~i_8_377_1851_0 & ~i_8_377_2047_0 & ~i_8_377_2118_0))) | (i_8_377_247_0 & ~i_8_377_361_0 & ~i_8_377_518_0 & ~i_8_377_669_0 & ~i_8_377_814_0 & ~i_8_377_817_0 & ~i_8_377_1434_0 & ~i_8_377_2028_0 & ~i_8_377_2047_0 & ~i_8_377_2113_0))) | (~i_8_377_654_0 & ((i_8_377_607_0 & ~i_8_377_685_0 & i_8_377_1984_0) | (i_8_377_427_0 & ~i_8_377_816_0 & ~i_8_377_1497_0 & ~i_8_377_1573_0 & i_8_377_2246_0))) | (i_8_377_2076_0 & ((~i_8_377_672_0 & ~i_8_377_703_0 & ~i_8_377_718_0 & ~i_8_377_1573_0 & ~i_8_377_1947_0 & ~i_8_377_1389_0 & ~i_8_377_1497_0) | (~i_8_377_762_0 & i_8_377_816_0 & ~i_8_377_1848_0 & ~i_8_377_2281_0))));
endmodule



// Benchmark "kernel_8_378" written by ABC on Sun Jul 19 10:09:40 2020

module kernel_8_378 ( 
    i_8_378_33_0, i_8_378_96_0, i_8_378_97_0, i_8_378_114_0, i_8_378_211_0,
    i_8_378_258_0, i_8_378_259_0, i_8_378_294_0, i_8_378_297_0,
    i_8_378_298_0, i_8_378_330_0, i_8_378_367_0, i_8_378_421_0,
    i_8_378_442_0, i_8_378_444_0, i_8_378_445_0, i_8_378_457_0,
    i_8_378_476_0, i_8_378_483_0, i_8_378_484_0, i_8_378_525_0,
    i_8_378_555_0, i_8_378_568_0, i_8_378_602_0, i_8_378_607_0,
    i_8_378_609_0, i_8_378_660_0, i_8_378_661_0, i_8_378_662_0,
    i_8_378_705_0, i_8_378_706_0, i_8_378_780_0, i_8_378_781_0,
    i_8_378_834_0, i_8_378_840_0, i_8_378_867_0, i_8_378_877_0,
    i_8_378_886_0, i_8_378_990_0, i_8_378_993_0, i_8_378_1026_0,
    i_8_378_1060_0, i_8_378_1071_0, i_8_378_1072_0, i_8_378_1074_0,
    i_8_378_1084_0, i_8_378_1111_0, i_8_378_1113_0, i_8_378_1141_0,
    i_8_378_1239_0, i_8_378_1261_0, i_8_378_1274_0, i_8_378_1283_0,
    i_8_378_1284_0, i_8_378_1285_0, i_8_378_1327_0, i_8_378_1392_0,
    i_8_378_1393_0, i_8_378_1408_0, i_8_378_1435_0, i_8_378_1437_0,
    i_8_378_1438_0, i_8_378_1507_0, i_8_378_1538_0, i_8_378_1584_0,
    i_8_378_1587_0, i_8_378_1590_0, i_8_378_1591_0, i_8_378_1598_0,
    i_8_378_1632_0, i_8_378_1633_0, i_8_378_1679_0, i_8_378_1699_0,
    i_8_378_1741_0, i_8_378_1744_0, i_8_378_1759_0, i_8_378_1761_0,
    i_8_378_1762_0, i_8_378_1821_0, i_8_378_1824_0, i_8_378_1825_0,
    i_8_378_1862_0, i_8_378_1902_0, i_8_378_1918_0, i_8_378_1989_0,
    i_8_378_1996_0, i_8_378_2058_0, i_8_378_2076_0, i_8_378_2089_0,
    i_8_378_2111_0, i_8_378_2114_0, i_8_378_2125_0, i_8_378_2187_0,
    i_8_378_2214_0, i_8_378_2215_0, i_8_378_2248_0, i_8_378_2249_0,
    i_8_378_2262_0, i_8_378_2295_0, i_8_378_2303_0,
    o_8_378_0_0  );
  input  i_8_378_33_0, i_8_378_96_0, i_8_378_97_0, i_8_378_114_0,
    i_8_378_211_0, i_8_378_258_0, i_8_378_259_0, i_8_378_294_0,
    i_8_378_297_0, i_8_378_298_0, i_8_378_330_0, i_8_378_367_0,
    i_8_378_421_0, i_8_378_442_0, i_8_378_444_0, i_8_378_445_0,
    i_8_378_457_0, i_8_378_476_0, i_8_378_483_0, i_8_378_484_0,
    i_8_378_525_0, i_8_378_555_0, i_8_378_568_0, i_8_378_602_0,
    i_8_378_607_0, i_8_378_609_0, i_8_378_660_0, i_8_378_661_0,
    i_8_378_662_0, i_8_378_705_0, i_8_378_706_0, i_8_378_780_0,
    i_8_378_781_0, i_8_378_834_0, i_8_378_840_0, i_8_378_867_0,
    i_8_378_877_0, i_8_378_886_0, i_8_378_990_0, i_8_378_993_0,
    i_8_378_1026_0, i_8_378_1060_0, i_8_378_1071_0, i_8_378_1072_0,
    i_8_378_1074_0, i_8_378_1084_0, i_8_378_1111_0, i_8_378_1113_0,
    i_8_378_1141_0, i_8_378_1239_0, i_8_378_1261_0, i_8_378_1274_0,
    i_8_378_1283_0, i_8_378_1284_0, i_8_378_1285_0, i_8_378_1327_0,
    i_8_378_1392_0, i_8_378_1393_0, i_8_378_1408_0, i_8_378_1435_0,
    i_8_378_1437_0, i_8_378_1438_0, i_8_378_1507_0, i_8_378_1538_0,
    i_8_378_1584_0, i_8_378_1587_0, i_8_378_1590_0, i_8_378_1591_0,
    i_8_378_1598_0, i_8_378_1632_0, i_8_378_1633_0, i_8_378_1679_0,
    i_8_378_1699_0, i_8_378_1741_0, i_8_378_1744_0, i_8_378_1759_0,
    i_8_378_1761_0, i_8_378_1762_0, i_8_378_1821_0, i_8_378_1824_0,
    i_8_378_1825_0, i_8_378_1862_0, i_8_378_1902_0, i_8_378_1918_0,
    i_8_378_1989_0, i_8_378_1996_0, i_8_378_2058_0, i_8_378_2076_0,
    i_8_378_2089_0, i_8_378_2111_0, i_8_378_2114_0, i_8_378_2125_0,
    i_8_378_2187_0, i_8_378_2214_0, i_8_378_2215_0, i_8_378_2248_0,
    i_8_378_2249_0, i_8_378_2262_0, i_8_378_2295_0, i_8_378_2303_0;
  output o_8_378_0_0;
  assign o_8_378_0_0 = ~((i_8_378_662_0 & ((~i_8_378_781_0 & ~i_8_378_1111_0 & i_8_378_1435_0 & ~i_8_378_1538_0 & ~i_8_378_1590_0 & i_8_378_1918_0) | (~i_8_378_602_0 & ~i_8_378_705_0 & ~i_8_378_1283_0 & ~i_8_378_1284_0 & i_8_378_2089_0 & ~i_8_378_2214_0))) | (i_8_378_706_0 & ((~i_8_378_1274_0 & ~i_8_378_1283_0 & ~i_8_378_1327_0 & ~i_8_378_1587_0) | (~i_8_378_484_0 & ~i_8_378_602_0 & i_8_378_1435_0 & ~i_8_378_2089_0 & ~i_8_378_2187_0 & ~i_8_378_2215_0))) | (~i_8_378_297_0 & ((~i_8_378_780_0 & ((~i_8_378_484_0 & i_8_378_1072_0 & ~i_8_378_1285_0 & ~i_8_378_1759_0) | (~i_8_378_476_0 & ~i_8_378_1026_0 & ~i_8_378_1261_0 & ~i_8_378_1283_0 & ~i_8_378_1408_0 & ~i_8_378_1584_0 & ~i_8_378_1591_0 & ~i_8_378_1762_0 & ~i_8_378_1824_0 & ~i_8_378_2076_0 & ~i_8_378_2125_0))) | (~i_8_378_1283_0 & ~i_8_378_1862_0 & ((~i_8_378_114_0 & ~i_8_378_607_0 & ~i_8_378_662_0 & ~i_8_378_840_0 & ~i_8_378_1284_0 & ~i_8_378_1507_0 & ~i_8_378_1591_0 & ~i_8_378_1744_0 & ~i_8_378_2187_0 & ~i_8_378_2215_0) | (~i_8_378_781_0 & ~i_8_378_1261_0 & ~i_8_378_1285_0 & ~i_8_378_1435_0 & ~i_8_378_1587_0 & ~i_8_378_1759_0 & ~i_8_378_2076_0 & ~i_8_378_2125_0 & ~i_8_378_2249_0))) | (~i_8_378_555_0 & ~i_8_378_1591_0 & i_8_378_1825_0 & ~i_8_378_2125_0))) | (~i_8_378_484_0 & ((i_8_378_660_0 & ~i_8_378_834_0 & i_8_378_1435_0 & ~i_8_378_1598_0 & ~i_8_378_2111_0) | (~i_8_378_476_0 & ~i_8_378_483_0 & ~i_8_378_555_0 & ~i_8_378_662_0 & ~i_8_378_1283_0 & ~i_8_378_1327_0 & ~i_8_378_1435_0 & ~i_8_378_1587_0 & ~i_8_378_1989_0 & ~i_8_378_2125_0 & ~i_8_378_2187_0 & ~i_8_378_2303_0))) | (~i_8_378_298_0 & ((~i_8_378_476_0 & ((~i_8_378_294_0 & ~i_8_378_1507_0 & ((~i_8_378_607_0 & ~i_8_378_877_0 & i_8_378_1111_0 & ~i_8_378_1327_0 & i_8_378_1438_0 & ~i_8_378_1590_0) | (~i_8_378_555_0 & ~i_8_378_1274_0 & ~i_8_378_1587_0 & ~i_8_378_1591_0 & ~i_8_378_1598_0 & ~i_8_378_1741_0 & ~i_8_378_1762_0 & ~i_8_378_2058_0 & ~i_8_378_2125_0 & ~i_8_378_2187_0))) | (~i_8_378_1283_0 & ((~i_8_378_1584_0 & ~i_8_378_1762_0 & ((~i_8_378_1538_0 & ~i_8_378_1587_0 & ~i_8_378_1590_0 & ~i_8_378_2125_0 & ~i_8_378_2214_0) | (~i_8_378_602_0 & ~i_8_378_834_0 & ~i_8_378_1111_0 & ~i_8_378_1393_0 & i_8_378_1918_0 & ~i_8_378_2249_0))) | (~i_8_378_483_0 & ~i_8_378_1590_0 & ~i_8_378_1741_0 & ~i_8_378_1918_0 & ~i_8_378_2187_0 & ~i_8_378_2303_0))) | (~i_8_378_525_0 & ~i_8_378_555_0 & ~i_8_378_662_0 & ~i_8_378_781_0 & ~i_8_378_867_0 & ~i_8_378_993_0 & ~i_8_378_1261_0 & ~i_8_378_1285_0 & ~i_8_378_1587_0 & ~i_8_378_1679_0))) | (~i_8_378_2111_0 & ((~i_8_378_483_0 & ((~i_8_378_993_0 & ~i_8_378_1285_0 & ~i_8_378_1507_0 & ~i_8_378_1587_0 & ~i_8_378_1744_0 & ~i_8_378_1918_0 & ~i_8_378_2114_0 & ~i_8_378_2214_0) | (~i_8_378_886_0 & ~i_8_378_1283_0 & ~i_8_378_1408_0 & ~i_8_378_1590_0 & ~i_8_378_2125_0 & ~i_8_378_2187_0 & ~i_8_378_2303_0 & ~i_8_378_1598_0 & i_8_378_1918_0))) | (~i_8_378_1285_0 & ~i_8_378_2187_0 & ((~i_8_378_607_0 & i_8_378_1111_0 & ~i_8_378_1507_0 & ~i_8_378_1761_0 & ~i_8_378_2248_0) | (~i_8_378_114_0 & ~i_8_378_555_0 & ~i_8_378_781_0 & ~i_8_378_867_0 & ~i_8_378_1261_0 & ~i_8_378_1435_0 & ~i_8_378_1591_0 & ~i_8_378_1598_0 & ~i_8_378_1762_0 & ~i_8_378_2249_0))))))) | (~i_8_378_2125_0 & ((~i_8_378_114_0 & ~i_8_378_1507_0 & ((~i_8_378_330_0 & ~i_8_378_867_0 & ~i_8_378_1584_0 & i_8_378_1821_0) | (~i_8_378_33_0 & ~i_8_378_607_0 & ~i_8_378_877_0 & ~i_8_378_1060_0 & ~i_8_378_1284_0 & ~i_8_378_1598_0 & ~i_8_378_1761_0 & ~i_8_378_1862_0 & ~i_8_378_1918_0 & ~i_8_378_2058_0 & ~i_8_378_2248_0 & ~i_8_378_2249_0))) | (~i_8_378_2187_0 & ((~i_8_378_607_0 & ((~i_8_378_1590_0 & ~i_8_378_1741_0 & i_8_378_840_0 & ~i_8_378_886_0) | (~i_8_378_993_0 & ~i_8_378_1327_0 & ~i_8_378_1408_0 & ~i_8_378_1538_0 & ~i_8_378_1598_0 & ~i_8_378_1632_0 & ~i_8_378_1633_0 & ~i_8_378_2111_0 & i_8_378_2215_0 & ~i_8_378_2303_0))) | (~i_8_378_602_0 & ~i_8_378_834_0 & ~i_8_378_1026_0 & ~i_8_378_1408_0 & ~i_8_378_1591_0 & ~i_8_378_1598_0 & ~i_8_378_1679_0 & ~i_8_378_1761_0 & ~i_8_378_1918_0 & ~i_8_378_2076_0 & ~i_8_378_2248_0))) | (~i_8_378_662_0 & i_8_378_1071_0 & ~i_8_378_1435_0 & ~i_8_378_2114_0) | (i_8_378_607_0 & ~i_8_378_1072_0 & ~i_8_378_1113_0 & ~i_8_378_1538_0 & i_8_378_1759_0 & ~i_8_378_2249_0))) | (~i_8_378_662_0 & ((~i_8_378_555_0 & ~i_8_378_1590_0 & ~i_8_378_1699_0 & ~i_8_378_1918_0 & i_8_378_1996_0) | (~i_8_378_211_0 & i_8_378_877_0 & ~i_8_378_1026_0 & ~i_8_378_1261_0 & ~i_8_378_1285_0 & ~i_8_378_1591_0 & ~i_8_378_1598_0 & ~i_8_378_1761_0 & ~i_8_378_1762_0 & ~i_8_378_2187_0 & ~i_8_378_2248_0))) | (~i_8_378_1026_0 & ((~i_8_378_609_0 & i_8_378_661_0 & ~i_8_378_886_0 & ~i_8_378_1538_0 & ~i_8_378_1590_0 & ~i_8_378_2214_0) | (i_8_378_705_0 & ~i_8_378_1762_0 & ~i_8_378_1862_0 & ~i_8_378_2215_0))) | (~i_8_378_1762_0 & ((i_8_378_1285_0 & ((~i_8_378_1261_0 & ~i_8_378_1584_0 & ~i_8_378_1591_0 & ~i_8_378_1598_0 & ~i_8_378_1679_0 & ~i_8_378_1741_0 & ~i_8_378_2089_0) | (~i_8_378_1438_0 & ~i_8_378_1507_0 & ~i_8_378_1761_0 & i_8_378_2111_0))) | (i_8_378_445_0 & ~i_8_378_2215_0 & ~i_8_378_2249_0))) | (~i_8_378_1584_0 & ~i_8_378_1598_0 & ~i_8_378_1744_0 & ((~i_8_378_568_0 & ~i_8_378_602_0 & i_8_378_1408_0 & ~i_8_378_1587_0 & ~i_8_378_1590_0 & ~i_8_378_1759_0 & ~i_8_378_2215_0 & ~i_8_378_2248_0) | (~i_8_378_294_0 & i_8_378_993_0 & ~i_8_378_1072_0 & ~i_8_378_2187_0 & ~i_8_378_2303_0 & ~i_8_378_1239_0 & ~i_8_378_1507_0))) | (~i_8_378_2187_0 & ((i_8_378_258_0 & i_8_378_1392_0) | (~i_8_378_421_0 & i_8_378_834_0 & i_8_378_840_0 & ~i_8_378_1071_0 & ~i_8_378_1633_0))) | (i_8_378_442_0 & ~i_8_378_607_0 & ~i_8_378_1761_0) | (i_8_378_457_0 & i_8_378_525_0 & i_8_378_886_0 & ~i_8_378_2214_0) | (i_8_378_484_0 & ~i_8_378_1284_0 & i_8_378_1996_0 & ~i_8_378_2111_0 & ~i_8_378_2215_0) | (~i_8_378_1918_0 & i_8_378_2076_0 & ~i_8_378_2248_0 & i_8_378_2295_0));
endmodule



// Benchmark "kernel_8_379" written by ABC on Sun Jul 19 10:09:41 2020

module kernel_8_379 ( 
    i_8_379_3_0, i_8_379_4_0, i_8_379_39_0, i_8_379_67_0, i_8_379_147_0,
    i_8_379_192_0, i_8_379_201_0, i_8_379_228_0, i_8_379_244_0,
    i_8_379_246_0, i_8_379_247_0, i_8_379_307_0, i_8_379_378_0,
    i_8_379_379_0, i_8_379_390_0, i_8_379_418_0, i_8_379_427_0,
    i_8_379_469_0, i_8_379_472_0, i_8_379_481_0, i_8_379_495_0,
    i_8_379_507_0, i_8_379_516_0, i_8_379_555_0, i_8_379_571_0,
    i_8_379_594_0, i_8_379_598_0, i_8_379_634_0, i_8_379_659_0,
    i_8_379_707_0, i_8_379_748_0, i_8_379_753_0, i_8_379_759_0,
    i_8_379_762_0, i_8_379_813_0, i_8_379_840_0, i_8_379_858_0,
    i_8_379_867_0, i_8_379_913_0, i_8_379_954_0, i_8_379_955_0,
    i_8_379_963_0, i_8_379_967_0, i_8_379_1030_0, i_8_379_1036_0,
    i_8_379_1071_0, i_8_379_1173_0, i_8_379_1191_0, i_8_379_1200_0,
    i_8_379_1203_0, i_8_379_1236_0, i_8_379_1269_0, i_8_379_1270_0,
    i_8_379_1296_0, i_8_379_1336_0, i_8_379_1353_0, i_8_379_1354_0,
    i_8_379_1389_0, i_8_379_1390_0, i_8_379_1401_0, i_8_379_1407_0,
    i_8_379_1485_0, i_8_379_1489_0, i_8_379_1494_0, i_8_379_1495_0,
    i_8_379_1497_0, i_8_379_1534_0, i_8_379_1597_0, i_8_379_1641_0,
    i_8_379_1651_0, i_8_379_1659_0, i_8_379_1696_0, i_8_379_1748_0,
    i_8_379_1750_0, i_8_379_1777_0, i_8_379_1794_0, i_8_379_1836_0,
    i_8_379_1848_0, i_8_379_1849_0, i_8_379_1855_0, i_8_379_1863_0,
    i_8_379_1872_0, i_8_379_1873_0, i_8_379_1882_0, i_8_379_1888_0,
    i_8_379_1911_0, i_8_379_1948_0, i_8_379_1950_0, i_8_379_1965_0,
    i_8_379_1971_0, i_8_379_2010_0, i_8_379_2047_0, i_8_379_2065_0,
    i_8_379_2091_0, i_8_379_2119_0, i_8_379_2146_0, i_8_379_2149_0,
    i_8_379_2229_0, i_8_379_2233_0, i_8_379_2256_0,
    o_8_379_0_0  );
  input  i_8_379_3_0, i_8_379_4_0, i_8_379_39_0, i_8_379_67_0,
    i_8_379_147_0, i_8_379_192_0, i_8_379_201_0, i_8_379_228_0,
    i_8_379_244_0, i_8_379_246_0, i_8_379_247_0, i_8_379_307_0,
    i_8_379_378_0, i_8_379_379_0, i_8_379_390_0, i_8_379_418_0,
    i_8_379_427_0, i_8_379_469_0, i_8_379_472_0, i_8_379_481_0,
    i_8_379_495_0, i_8_379_507_0, i_8_379_516_0, i_8_379_555_0,
    i_8_379_571_0, i_8_379_594_0, i_8_379_598_0, i_8_379_634_0,
    i_8_379_659_0, i_8_379_707_0, i_8_379_748_0, i_8_379_753_0,
    i_8_379_759_0, i_8_379_762_0, i_8_379_813_0, i_8_379_840_0,
    i_8_379_858_0, i_8_379_867_0, i_8_379_913_0, i_8_379_954_0,
    i_8_379_955_0, i_8_379_963_0, i_8_379_967_0, i_8_379_1030_0,
    i_8_379_1036_0, i_8_379_1071_0, i_8_379_1173_0, i_8_379_1191_0,
    i_8_379_1200_0, i_8_379_1203_0, i_8_379_1236_0, i_8_379_1269_0,
    i_8_379_1270_0, i_8_379_1296_0, i_8_379_1336_0, i_8_379_1353_0,
    i_8_379_1354_0, i_8_379_1389_0, i_8_379_1390_0, i_8_379_1401_0,
    i_8_379_1407_0, i_8_379_1485_0, i_8_379_1489_0, i_8_379_1494_0,
    i_8_379_1495_0, i_8_379_1497_0, i_8_379_1534_0, i_8_379_1597_0,
    i_8_379_1641_0, i_8_379_1651_0, i_8_379_1659_0, i_8_379_1696_0,
    i_8_379_1748_0, i_8_379_1750_0, i_8_379_1777_0, i_8_379_1794_0,
    i_8_379_1836_0, i_8_379_1848_0, i_8_379_1849_0, i_8_379_1855_0,
    i_8_379_1863_0, i_8_379_1872_0, i_8_379_1873_0, i_8_379_1882_0,
    i_8_379_1888_0, i_8_379_1911_0, i_8_379_1948_0, i_8_379_1950_0,
    i_8_379_1965_0, i_8_379_1971_0, i_8_379_2010_0, i_8_379_2047_0,
    i_8_379_2065_0, i_8_379_2091_0, i_8_379_2119_0, i_8_379_2146_0,
    i_8_379_2149_0, i_8_379_2229_0, i_8_379_2233_0, i_8_379_2256_0;
  output o_8_379_0_0;
  assign o_8_379_0_0 = 0;
endmodule



// Benchmark "kernel_8_380" written by ABC on Sun Jul 19 10:09:42 2020

module kernel_8_380 ( 
    i_8_380_28_0, i_8_380_31_0, i_8_380_54_0, i_8_380_56_0, i_8_380_118_0,
    i_8_380_218_0, i_8_380_221_0, i_8_380_227_0, i_8_380_253_0,
    i_8_380_365_0, i_8_380_417_0, i_8_380_451_0, i_8_380_478_0,
    i_8_380_480_0, i_8_380_481_0, i_8_380_500_0, i_8_380_507_0,
    i_8_380_545_0, i_8_380_552_0, i_8_380_553_0, i_8_380_582_0,
    i_8_380_594_0, i_8_380_599_0, i_8_380_604_0, i_8_380_606_0,
    i_8_380_607_0, i_8_380_608_0, i_8_380_612_0, i_8_380_649_0,
    i_8_380_655_0, i_8_380_660_0, i_8_380_715_0, i_8_380_756_0,
    i_8_380_768_0, i_8_380_781_0, i_8_380_789_0, i_8_380_795_0,
    i_8_380_847_0, i_8_380_903_0, i_8_380_981_0, i_8_380_1008_0,
    i_8_380_1059_0, i_8_380_1060_0, i_8_380_1110_0, i_8_380_1111_0,
    i_8_380_1127_0, i_8_380_1130_0, i_8_380_1234_0, i_8_380_1260_0,
    i_8_380_1261_0, i_8_380_1292_0, i_8_380_1297_0, i_8_380_1307_0,
    i_8_380_1344_0, i_8_380_1345_0, i_8_380_1350_0, i_8_380_1379_0,
    i_8_380_1401_0, i_8_380_1416_0, i_8_380_1431_0, i_8_380_1443_0,
    i_8_380_1468_0, i_8_380_1541_0, i_8_380_1552_0, i_8_380_1555_0,
    i_8_380_1578_0, i_8_380_1588_0, i_8_380_1603_0, i_8_380_1680_0,
    i_8_380_1752_0, i_8_380_1753_0, i_8_380_1755_0, i_8_380_1756_0,
    i_8_380_1775_0, i_8_380_1783_0, i_8_380_1784_0, i_8_380_1788_0,
    i_8_380_1789_0, i_8_380_1801_0, i_8_380_1810_0, i_8_380_1822_0,
    i_8_380_1825_0, i_8_380_1837_0, i_8_380_1945_0, i_8_380_1946_0,
    i_8_380_1949_0, i_8_380_1973_0, i_8_380_1998_0, i_8_380_2050_0,
    i_8_380_2133_0, i_8_380_2142_0, i_8_380_2152_0, i_8_380_2153_0,
    i_8_380_2170_0, i_8_380_2214_0, i_8_380_2224_0, i_8_380_2227_0,
    i_8_380_2232_0, i_8_380_2287_0, i_8_380_2292_0,
    o_8_380_0_0  );
  input  i_8_380_28_0, i_8_380_31_0, i_8_380_54_0, i_8_380_56_0,
    i_8_380_118_0, i_8_380_218_0, i_8_380_221_0, i_8_380_227_0,
    i_8_380_253_0, i_8_380_365_0, i_8_380_417_0, i_8_380_451_0,
    i_8_380_478_0, i_8_380_480_0, i_8_380_481_0, i_8_380_500_0,
    i_8_380_507_0, i_8_380_545_0, i_8_380_552_0, i_8_380_553_0,
    i_8_380_582_0, i_8_380_594_0, i_8_380_599_0, i_8_380_604_0,
    i_8_380_606_0, i_8_380_607_0, i_8_380_608_0, i_8_380_612_0,
    i_8_380_649_0, i_8_380_655_0, i_8_380_660_0, i_8_380_715_0,
    i_8_380_756_0, i_8_380_768_0, i_8_380_781_0, i_8_380_789_0,
    i_8_380_795_0, i_8_380_847_0, i_8_380_903_0, i_8_380_981_0,
    i_8_380_1008_0, i_8_380_1059_0, i_8_380_1060_0, i_8_380_1110_0,
    i_8_380_1111_0, i_8_380_1127_0, i_8_380_1130_0, i_8_380_1234_0,
    i_8_380_1260_0, i_8_380_1261_0, i_8_380_1292_0, i_8_380_1297_0,
    i_8_380_1307_0, i_8_380_1344_0, i_8_380_1345_0, i_8_380_1350_0,
    i_8_380_1379_0, i_8_380_1401_0, i_8_380_1416_0, i_8_380_1431_0,
    i_8_380_1443_0, i_8_380_1468_0, i_8_380_1541_0, i_8_380_1552_0,
    i_8_380_1555_0, i_8_380_1578_0, i_8_380_1588_0, i_8_380_1603_0,
    i_8_380_1680_0, i_8_380_1752_0, i_8_380_1753_0, i_8_380_1755_0,
    i_8_380_1756_0, i_8_380_1775_0, i_8_380_1783_0, i_8_380_1784_0,
    i_8_380_1788_0, i_8_380_1789_0, i_8_380_1801_0, i_8_380_1810_0,
    i_8_380_1822_0, i_8_380_1825_0, i_8_380_1837_0, i_8_380_1945_0,
    i_8_380_1946_0, i_8_380_1949_0, i_8_380_1973_0, i_8_380_1998_0,
    i_8_380_2050_0, i_8_380_2133_0, i_8_380_2142_0, i_8_380_2152_0,
    i_8_380_2153_0, i_8_380_2170_0, i_8_380_2214_0, i_8_380_2224_0,
    i_8_380_2227_0, i_8_380_2232_0, i_8_380_2287_0, i_8_380_2292_0;
  output o_8_380_0_0;
  assign o_8_380_0_0 = 0;
endmodule



// Benchmark "kernel_8_381" written by ABC on Sun Jul 19 10:09:43 2020

module kernel_8_381 ( 
    i_8_381_32_0, i_8_381_51_0, i_8_381_95_0, i_8_381_97_0, i_8_381_114_0,
    i_8_381_115_0, i_8_381_141_0, i_8_381_258_0, i_8_381_331_0,
    i_8_381_332_0, i_8_381_377_0, i_8_381_383_0, i_8_381_421_0,
    i_8_381_457_0, i_8_381_462_0, i_8_381_463_0, i_8_381_476_0,
    i_8_381_479_0, i_8_381_482_0, i_8_381_527_0, i_8_381_553_0,
    i_8_381_556_0, i_8_381_606_0, i_8_381_608_0, i_8_381_661_0,
    i_8_381_662_0, i_8_381_663_0, i_8_381_682_0, i_8_381_782_0,
    i_8_381_817_0, i_8_381_818_0, i_8_381_840_0, i_8_381_841_0,
    i_8_381_847_0, i_8_381_851_0, i_8_381_1074_0, i_8_381_1077_0,
    i_8_381_1239_0, i_8_381_1240_0, i_8_381_1259_0, i_8_381_1283_0,
    i_8_381_1292_0, i_8_381_1307_0, i_8_381_1437_0, i_8_381_1438_0,
    i_8_381_1439_0, i_8_381_1534_0, i_8_381_1535_0, i_8_381_1540_0,
    i_8_381_1551_0, i_8_381_1588_0, i_8_381_1589_0, i_8_381_1590_0,
    i_8_381_1591_0, i_8_381_1592_0, i_8_381_1600_0, i_8_381_1615_0,
    i_8_381_1616_0, i_8_381_1633_0, i_8_381_1634_0, i_8_381_1636_0,
    i_8_381_1637_0, i_8_381_1671_0, i_8_381_1679_0, i_8_381_1680_0,
    i_8_381_1742_0, i_8_381_1744_0, i_8_381_1751_0, i_8_381_1760_0,
    i_8_381_1761_0, i_8_381_1762_0, i_8_381_1763_0, i_8_381_1825_0,
    i_8_381_1826_0, i_8_381_1834_0, i_8_381_1839_0, i_8_381_1843_0,
    i_8_381_1879_0, i_8_381_1904_0, i_8_381_1922_0, i_8_381_1967_0,
    i_8_381_1985_0, i_8_381_1993_0, i_8_381_1994_0, i_8_381_1997_0,
    i_8_381_2056_0, i_8_381_2059_0, i_8_381_2090_0, i_8_381_2107_0,
    i_8_381_2130_0, i_8_381_2149_0, i_8_381_2172_0, i_8_381_2190_0,
    i_8_381_2214_0, i_8_381_2215_0, i_8_381_2216_0, i_8_381_2219_0,
    i_8_381_2264_0, i_8_381_2296_0, i_8_381_2303_0,
    o_8_381_0_0  );
  input  i_8_381_32_0, i_8_381_51_0, i_8_381_95_0, i_8_381_97_0,
    i_8_381_114_0, i_8_381_115_0, i_8_381_141_0, i_8_381_258_0,
    i_8_381_331_0, i_8_381_332_0, i_8_381_377_0, i_8_381_383_0,
    i_8_381_421_0, i_8_381_457_0, i_8_381_462_0, i_8_381_463_0,
    i_8_381_476_0, i_8_381_479_0, i_8_381_482_0, i_8_381_527_0,
    i_8_381_553_0, i_8_381_556_0, i_8_381_606_0, i_8_381_608_0,
    i_8_381_661_0, i_8_381_662_0, i_8_381_663_0, i_8_381_682_0,
    i_8_381_782_0, i_8_381_817_0, i_8_381_818_0, i_8_381_840_0,
    i_8_381_841_0, i_8_381_847_0, i_8_381_851_0, i_8_381_1074_0,
    i_8_381_1077_0, i_8_381_1239_0, i_8_381_1240_0, i_8_381_1259_0,
    i_8_381_1283_0, i_8_381_1292_0, i_8_381_1307_0, i_8_381_1437_0,
    i_8_381_1438_0, i_8_381_1439_0, i_8_381_1534_0, i_8_381_1535_0,
    i_8_381_1540_0, i_8_381_1551_0, i_8_381_1588_0, i_8_381_1589_0,
    i_8_381_1590_0, i_8_381_1591_0, i_8_381_1592_0, i_8_381_1600_0,
    i_8_381_1615_0, i_8_381_1616_0, i_8_381_1633_0, i_8_381_1634_0,
    i_8_381_1636_0, i_8_381_1637_0, i_8_381_1671_0, i_8_381_1679_0,
    i_8_381_1680_0, i_8_381_1742_0, i_8_381_1744_0, i_8_381_1751_0,
    i_8_381_1760_0, i_8_381_1761_0, i_8_381_1762_0, i_8_381_1763_0,
    i_8_381_1825_0, i_8_381_1826_0, i_8_381_1834_0, i_8_381_1839_0,
    i_8_381_1843_0, i_8_381_1879_0, i_8_381_1904_0, i_8_381_1922_0,
    i_8_381_1967_0, i_8_381_1985_0, i_8_381_1993_0, i_8_381_1994_0,
    i_8_381_1997_0, i_8_381_2056_0, i_8_381_2059_0, i_8_381_2090_0,
    i_8_381_2107_0, i_8_381_2130_0, i_8_381_2149_0, i_8_381_2172_0,
    i_8_381_2190_0, i_8_381_2214_0, i_8_381_2215_0, i_8_381_2216_0,
    i_8_381_2219_0, i_8_381_2264_0, i_8_381_2296_0, i_8_381_2303_0;
  output o_8_381_0_0;
  assign o_8_381_0_0 = ~((~i_8_381_383_0 & ((~i_8_381_114_0 & ~i_8_381_377_0 & ~i_8_381_606_0 & ~i_8_381_1535_0 & ~i_8_381_2056_0 & ~i_8_381_2059_0 & ~i_8_381_2130_0) | (i_8_381_377_0 & ~i_8_381_1439_0 & ~i_8_381_1590_0 & ~i_8_381_2190_0))) | (~i_8_381_462_0 & ((~i_8_381_476_0 & ~i_8_381_1239_0 & ~i_8_381_1283_0 & ~i_8_381_1592_0 & ~i_8_381_1760_0 & ~i_8_381_1761_0 & ~i_8_381_1763_0 & ~i_8_381_1839_0) | (~i_8_381_527_0 & ~i_8_381_556_0 & ~i_8_381_1535_0 & ~i_8_381_1744_0 & ~i_8_381_1879_0 & ~i_8_381_2172_0))) | (~i_8_381_2059_0 & ((~i_8_381_482_0 & ((~i_8_381_476_0 & ~i_8_381_606_0 & ~i_8_381_1077_0 & ~i_8_381_1535_0 & ~i_8_381_1540_0 & ~i_8_381_1636_0 & ~i_8_381_1761_0) | (~i_8_381_661_0 & ~i_8_381_1259_0 & ~i_8_381_1590_0 & ~i_8_381_1762_0 & ~i_8_381_1763_0 & ~i_8_381_2214_0))) | (~i_8_381_608_0 & i_8_381_1240_0 & i_8_381_1438_0 & i_8_381_1439_0 & ~i_8_381_1540_0 & ~i_8_381_1834_0 & ~i_8_381_2172_0 & ~i_8_381_2215_0))) | (~i_8_381_1590_0 & ((~i_8_381_476_0 & ((~i_8_381_1615_0 & i_8_381_1634_0 & ~i_8_381_2090_0 & ~i_8_381_2130_0) | (i_8_381_482_0 & ~i_8_381_818_0 & ~i_8_381_1283_0 & ~i_8_381_1839_0 & ~i_8_381_1997_0 & ~i_8_381_2056_0 & ~i_8_381_2107_0 & ~i_8_381_2172_0))) | (i_8_381_1437_0 & ~i_8_381_1535_0 & ~i_8_381_1588_0 & ~i_8_381_1600_0 & ~i_8_381_1834_0 & ~i_8_381_2056_0 & ~i_8_381_2107_0) | (~i_8_381_608_0 & ~i_8_381_1437_0 & i_8_381_1993_0) | (~i_8_381_527_0 & i_8_381_661_0 & ~i_8_381_2190_0))) | (~i_8_381_463_0 & ((~i_8_381_606_0 & ((~i_8_381_1534_0 & ~i_8_381_1763_0 & i_8_381_1825_0) | (~i_8_381_1589_0 & ~i_8_381_1592_0 & ~i_8_381_1744_0 & ~i_8_381_1839_0 & ~i_8_381_1922_0 & ~i_8_381_2219_0 & ~i_8_381_2296_0))) | (~i_8_381_556_0 & ~i_8_381_1240_0 & ~i_8_381_1283_0 & ~i_8_381_1535_0 & ~i_8_381_2090_0 & ~i_8_381_2130_0 & ~i_8_381_1615_0 & ~i_8_381_1671_0) | (~i_8_381_32_0 & i_8_381_1438_0 & ~i_8_381_1600_0 & ~i_8_381_1744_0 & ~i_8_381_1760_0 & ~i_8_381_1879_0 & ~i_8_381_2149_0 & ~i_8_381_2190_0 & ~i_8_381_2219_0) | (~i_8_381_1534_0 & ~i_8_381_1540_0 & ~i_8_381_1592_0 & ~i_8_381_1680_0 & ~i_8_381_1834_0 & ~i_8_381_2215_0))) | (~i_8_381_1437_0 & ((~i_8_381_1259_0 & ~i_8_381_1540_0 & ~i_8_381_1588_0 & ~i_8_381_1839_0 & ~i_8_381_2219_0) | (~i_8_381_661_0 & ~i_8_381_1074_0 & ~i_8_381_1438_0 & ~i_8_381_1439_0 & ~i_8_381_1763_0 & ~i_8_381_1843_0 & ~i_8_381_1985_0 & ~i_8_381_2190_0 & ~i_8_381_2296_0))) | (~i_8_381_115_0 & ~i_8_381_421_0 & ~i_8_381_553_0 & ~i_8_381_1535_0 & ~i_8_381_1591_0 & ~i_8_381_1834_0 & ~i_8_381_2090_0) | (~i_8_381_1592_0 & ~i_8_381_1600_0 & ~i_8_381_1616_0 & ~i_8_381_1761_0 & ~i_8_381_1762_0 & ~i_8_381_2149_0 & ~i_8_381_2190_0 & ~i_8_381_2214_0 & ~i_8_381_2296_0));
endmodule



// Benchmark "kernel_8_382" written by ABC on Sun Jul 19 10:09:44 2020

module kernel_8_382 ( 
    i_8_382_28_0, i_8_382_57_0, i_8_382_87_0, i_8_382_143_0, i_8_382_214_0,
    i_8_382_264_0, i_8_382_268_0, i_8_382_269_0, i_8_382_328_0,
    i_8_382_349_0, i_8_382_360_0, i_8_382_376_0, i_8_382_378_0,
    i_8_382_379_0, i_8_382_381_0, i_8_382_384_0, i_8_382_417_0,
    i_8_382_463_0, i_8_382_481_0, i_8_382_490_0, i_8_382_500_0,
    i_8_382_529_0, i_8_382_589_0, i_8_382_590_0, i_8_382_592_0,
    i_8_382_599_0, i_8_382_608_0, i_8_382_611_0, i_8_382_615_0,
    i_8_382_616_0, i_8_382_628_0, i_8_382_633_0, i_8_382_637_0,
    i_8_382_638_0, i_8_382_661_0, i_8_382_664_0, i_8_382_670_0,
    i_8_382_682_0, i_8_382_715_0, i_8_382_716_0, i_8_382_760_0,
    i_8_382_769_0, i_8_382_778_0, i_8_382_823_0, i_8_382_843_0,
    i_8_382_870_0, i_8_382_871_0, i_8_382_898_0, i_8_382_899_0,
    i_8_382_984_0, i_8_382_985_0, i_8_382_1016_0, i_8_382_1079_0,
    i_8_382_1086_0, i_8_382_1110_0, i_8_382_1111_0, i_8_382_1114_0,
    i_8_382_1189_0, i_8_382_1236_0, i_8_382_1250_0, i_8_382_1281_0,
    i_8_382_1305_0, i_8_382_1307_0, i_8_382_1328_0, i_8_382_1345_0,
    i_8_382_1347_0, i_8_382_1449_0, i_8_382_1455_0, i_8_382_1456_0,
    i_8_382_1492_0, i_8_382_1534_0, i_8_382_1538_0, i_8_382_1579_0,
    i_8_382_1605_0, i_8_382_1606_0, i_8_382_1607_0, i_8_382_1608_0,
    i_8_382_1609_0, i_8_382_1644_0, i_8_382_1671_0, i_8_382_1706_0,
    i_8_382_1725_0, i_8_382_1726_0, i_8_382_1749_0, i_8_382_1763_0,
    i_8_382_1779_0, i_8_382_1823_0, i_8_382_1834_0, i_8_382_1870_0,
    i_8_382_1952_0, i_8_382_2012_0, i_8_382_2014_0, i_8_382_2050_0,
    i_8_382_2092_0, i_8_382_2129_0, i_8_382_2173_0, i_8_382_2199_0,
    i_8_382_2275_0, i_8_382_2293_0, i_8_382_2294_0,
    o_8_382_0_0  );
  input  i_8_382_28_0, i_8_382_57_0, i_8_382_87_0, i_8_382_143_0,
    i_8_382_214_0, i_8_382_264_0, i_8_382_268_0, i_8_382_269_0,
    i_8_382_328_0, i_8_382_349_0, i_8_382_360_0, i_8_382_376_0,
    i_8_382_378_0, i_8_382_379_0, i_8_382_381_0, i_8_382_384_0,
    i_8_382_417_0, i_8_382_463_0, i_8_382_481_0, i_8_382_490_0,
    i_8_382_500_0, i_8_382_529_0, i_8_382_589_0, i_8_382_590_0,
    i_8_382_592_0, i_8_382_599_0, i_8_382_608_0, i_8_382_611_0,
    i_8_382_615_0, i_8_382_616_0, i_8_382_628_0, i_8_382_633_0,
    i_8_382_637_0, i_8_382_638_0, i_8_382_661_0, i_8_382_664_0,
    i_8_382_670_0, i_8_382_682_0, i_8_382_715_0, i_8_382_716_0,
    i_8_382_760_0, i_8_382_769_0, i_8_382_778_0, i_8_382_823_0,
    i_8_382_843_0, i_8_382_870_0, i_8_382_871_0, i_8_382_898_0,
    i_8_382_899_0, i_8_382_984_0, i_8_382_985_0, i_8_382_1016_0,
    i_8_382_1079_0, i_8_382_1086_0, i_8_382_1110_0, i_8_382_1111_0,
    i_8_382_1114_0, i_8_382_1189_0, i_8_382_1236_0, i_8_382_1250_0,
    i_8_382_1281_0, i_8_382_1305_0, i_8_382_1307_0, i_8_382_1328_0,
    i_8_382_1345_0, i_8_382_1347_0, i_8_382_1449_0, i_8_382_1455_0,
    i_8_382_1456_0, i_8_382_1492_0, i_8_382_1534_0, i_8_382_1538_0,
    i_8_382_1579_0, i_8_382_1605_0, i_8_382_1606_0, i_8_382_1607_0,
    i_8_382_1608_0, i_8_382_1609_0, i_8_382_1644_0, i_8_382_1671_0,
    i_8_382_1706_0, i_8_382_1725_0, i_8_382_1726_0, i_8_382_1749_0,
    i_8_382_1763_0, i_8_382_1779_0, i_8_382_1823_0, i_8_382_1834_0,
    i_8_382_1870_0, i_8_382_1952_0, i_8_382_2012_0, i_8_382_2014_0,
    i_8_382_2050_0, i_8_382_2092_0, i_8_382_2129_0, i_8_382_2173_0,
    i_8_382_2199_0, i_8_382_2275_0, i_8_382_2293_0, i_8_382_2294_0;
  output o_8_382_0_0;
  assign o_8_382_0_0 = 0;
endmodule



// Benchmark "kernel_8_383" written by ABC on Sun Jul 19 10:09:45 2020

module kernel_8_383 ( 
    i_8_383_12_0, i_8_383_31_0, i_8_383_58_0, i_8_383_64_0, i_8_383_136_0,
    i_8_383_180_0, i_8_383_185_0, i_8_383_221_0, i_8_383_226_0,
    i_8_383_289_0, i_8_383_301_0, i_8_383_335_0, i_8_383_386_0,
    i_8_383_389_0, i_8_383_397_0, i_8_383_423_0, i_8_383_427_0,
    i_8_383_433_0, i_8_383_453_0, i_8_383_479_0, i_8_383_507_0,
    i_8_383_517_0, i_8_383_530_0, i_8_383_557_0, i_8_383_587_0,
    i_8_383_614_0, i_8_383_652_0, i_8_383_657_0, i_8_383_661_0,
    i_8_383_676_0, i_8_383_677_0, i_8_383_758_0, i_8_383_790_0,
    i_8_383_821_0, i_8_383_847_0, i_8_383_848_0, i_8_383_865_0,
    i_8_383_868_0, i_8_383_875_0, i_8_383_881_0, i_8_383_882_0,
    i_8_383_883_0, i_8_383_884_0, i_8_383_998_0, i_8_383_1049_0,
    i_8_383_1103_0, i_8_383_1106_0, i_8_383_1110_0, i_8_383_1115_0,
    i_8_383_1156_0, i_8_383_1199_0, i_8_383_1237_0, i_8_383_1255_0,
    i_8_383_1265_0, i_8_383_1286_0, i_8_383_1296_0, i_8_383_1298_0,
    i_8_383_1333_0, i_8_383_1340_0, i_8_383_1403_0, i_8_383_1408_0,
    i_8_383_1423_0, i_8_383_1435_0, i_8_383_1481_0, i_8_383_1507_0,
    i_8_383_1508_0, i_8_383_1539_0, i_8_383_1545_0, i_8_383_1558_0,
    i_8_383_1561_0, i_8_383_1581_0, i_8_383_1631_0, i_8_383_1642_0,
    i_8_383_1682_0, i_8_383_1683_0, i_8_383_1684_0, i_8_383_1737_0,
    i_8_383_1749_0, i_8_383_1750_0, i_8_383_1767_0, i_8_383_1771_0,
    i_8_383_1772_0, i_8_383_1778_0, i_8_383_1846_0, i_8_383_1881_0,
    i_8_383_1884_0, i_8_383_1885_0, i_8_383_1888_0, i_8_383_1947_0,
    i_8_383_1981_0, i_8_383_1992_0, i_8_383_2045_0, i_8_383_2098_0,
    i_8_383_2126_0, i_8_383_2170_0, i_8_383_2173_0, i_8_383_2268_0,
    i_8_383_2296_0, i_8_383_2297_0, i_8_383_2299_0,
    o_8_383_0_0  );
  input  i_8_383_12_0, i_8_383_31_0, i_8_383_58_0, i_8_383_64_0,
    i_8_383_136_0, i_8_383_180_0, i_8_383_185_0, i_8_383_221_0,
    i_8_383_226_0, i_8_383_289_0, i_8_383_301_0, i_8_383_335_0,
    i_8_383_386_0, i_8_383_389_0, i_8_383_397_0, i_8_383_423_0,
    i_8_383_427_0, i_8_383_433_0, i_8_383_453_0, i_8_383_479_0,
    i_8_383_507_0, i_8_383_517_0, i_8_383_530_0, i_8_383_557_0,
    i_8_383_587_0, i_8_383_614_0, i_8_383_652_0, i_8_383_657_0,
    i_8_383_661_0, i_8_383_676_0, i_8_383_677_0, i_8_383_758_0,
    i_8_383_790_0, i_8_383_821_0, i_8_383_847_0, i_8_383_848_0,
    i_8_383_865_0, i_8_383_868_0, i_8_383_875_0, i_8_383_881_0,
    i_8_383_882_0, i_8_383_883_0, i_8_383_884_0, i_8_383_998_0,
    i_8_383_1049_0, i_8_383_1103_0, i_8_383_1106_0, i_8_383_1110_0,
    i_8_383_1115_0, i_8_383_1156_0, i_8_383_1199_0, i_8_383_1237_0,
    i_8_383_1255_0, i_8_383_1265_0, i_8_383_1286_0, i_8_383_1296_0,
    i_8_383_1298_0, i_8_383_1333_0, i_8_383_1340_0, i_8_383_1403_0,
    i_8_383_1408_0, i_8_383_1423_0, i_8_383_1435_0, i_8_383_1481_0,
    i_8_383_1507_0, i_8_383_1508_0, i_8_383_1539_0, i_8_383_1545_0,
    i_8_383_1558_0, i_8_383_1561_0, i_8_383_1581_0, i_8_383_1631_0,
    i_8_383_1642_0, i_8_383_1682_0, i_8_383_1683_0, i_8_383_1684_0,
    i_8_383_1737_0, i_8_383_1749_0, i_8_383_1750_0, i_8_383_1767_0,
    i_8_383_1771_0, i_8_383_1772_0, i_8_383_1778_0, i_8_383_1846_0,
    i_8_383_1881_0, i_8_383_1884_0, i_8_383_1885_0, i_8_383_1888_0,
    i_8_383_1947_0, i_8_383_1981_0, i_8_383_1992_0, i_8_383_2045_0,
    i_8_383_2098_0, i_8_383_2126_0, i_8_383_2170_0, i_8_383_2173_0,
    i_8_383_2268_0, i_8_383_2296_0, i_8_383_2297_0, i_8_383_2299_0;
  output o_8_383_0_0;
  assign o_8_383_0_0 = 0;
endmodule



// Benchmark "kernel_8_384" written by ABC on Sun Jul 19 10:09:46 2020

module kernel_8_384 ( 
    i_8_384_11_0, i_8_384_80_0, i_8_384_85_0, i_8_384_120_0, i_8_384_121_0,
    i_8_384_143_0, i_8_384_147_0, i_8_384_184_0, i_8_384_191_0,
    i_8_384_316_0, i_8_384_317_0, i_8_384_360_0, i_8_384_361_0,
    i_8_384_366_0, i_8_384_368_0, i_8_384_386_0, i_8_384_435_0,
    i_8_384_500_0, i_8_384_508_0, i_8_384_532_0, i_8_384_533_0,
    i_8_384_535_0, i_8_384_580_0, i_8_384_604_0, i_8_384_633_0,
    i_8_384_644_0, i_8_384_653_0, i_8_384_656_0, i_8_384_662_0,
    i_8_384_732_0, i_8_384_733_0, i_8_384_748_0, i_8_384_749_0,
    i_8_384_787_0, i_8_384_826_0, i_8_384_829_0, i_8_384_831_0,
    i_8_384_850_0, i_8_384_872_0, i_8_384_873_0, i_8_384_893_0,
    i_8_384_1037_0, i_8_384_1103_0, i_8_384_1138_0, i_8_384_1153_0,
    i_8_384_1202_0, i_8_384_1227_0, i_8_384_1240_0, i_8_384_1241_0,
    i_8_384_1244_0, i_8_384_1256_0, i_8_384_1319_0, i_8_384_1327_0,
    i_8_384_1336_0, i_8_384_1354_0, i_8_384_1364_0, i_8_384_1424_0,
    i_8_384_1456_0, i_8_384_1457_0, i_8_384_1462_0, i_8_384_1463_0,
    i_8_384_1471_0, i_8_384_1478_0, i_8_384_1493_0, i_8_384_1514_0,
    i_8_384_1522_0, i_8_384_1526_0, i_8_384_1540_0, i_8_384_1544_0,
    i_8_384_1570_0, i_8_384_1571_0, i_8_384_1591_0, i_8_384_1675_0,
    i_8_384_1696_0, i_8_384_1702_0, i_8_384_1703_0, i_8_384_1748_0,
    i_8_384_1766_0, i_8_384_1781_0, i_8_384_1783_0, i_8_384_1821_0,
    i_8_384_1844_0, i_8_384_1858_0, i_8_384_1882_0, i_8_384_1883_0,
    i_8_384_1892_0, i_8_384_1936_0, i_8_384_1954_0, i_8_384_1958_0,
    i_8_384_1975_0, i_8_384_1976_0, i_8_384_1985_0, i_8_384_1992_0,
    i_8_384_2044_0, i_8_384_2146_0, i_8_384_2155_0, i_8_384_2227_0,
    i_8_384_2231_0, i_8_384_2246_0, i_8_384_2257_0,
    o_8_384_0_0  );
  input  i_8_384_11_0, i_8_384_80_0, i_8_384_85_0, i_8_384_120_0,
    i_8_384_121_0, i_8_384_143_0, i_8_384_147_0, i_8_384_184_0,
    i_8_384_191_0, i_8_384_316_0, i_8_384_317_0, i_8_384_360_0,
    i_8_384_361_0, i_8_384_366_0, i_8_384_368_0, i_8_384_386_0,
    i_8_384_435_0, i_8_384_500_0, i_8_384_508_0, i_8_384_532_0,
    i_8_384_533_0, i_8_384_535_0, i_8_384_580_0, i_8_384_604_0,
    i_8_384_633_0, i_8_384_644_0, i_8_384_653_0, i_8_384_656_0,
    i_8_384_662_0, i_8_384_732_0, i_8_384_733_0, i_8_384_748_0,
    i_8_384_749_0, i_8_384_787_0, i_8_384_826_0, i_8_384_829_0,
    i_8_384_831_0, i_8_384_850_0, i_8_384_872_0, i_8_384_873_0,
    i_8_384_893_0, i_8_384_1037_0, i_8_384_1103_0, i_8_384_1138_0,
    i_8_384_1153_0, i_8_384_1202_0, i_8_384_1227_0, i_8_384_1240_0,
    i_8_384_1241_0, i_8_384_1244_0, i_8_384_1256_0, i_8_384_1319_0,
    i_8_384_1327_0, i_8_384_1336_0, i_8_384_1354_0, i_8_384_1364_0,
    i_8_384_1424_0, i_8_384_1456_0, i_8_384_1457_0, i_8_384_1462_0,
    i_8_384_1463_0, i_8_384_1471_0, i_8_384_1478_0, i_8_384_1493_0,
    i_8_384_1514_0, i_8_384_1522_0, i_8_384_1526_0, i_8_384_1540_0,
    i_8_384_1544_0, i_8_384_1570_0, i_8_384_1571_0, i_8_384_1591_0,
    i_8_384_1675_0, i_8_384_1696_0, i_8_384_1702_0, i_8_384_1703_0,
    i_8_384_1748_0, i_8_384_1766_0, i_8_384_1781_0, i_8_384_1783_0,
    i_8_384_1821_0, i_8_384_1844_0, i_8_384_1858_0, i_8_384_1882_0,
    i_8_384_1883_0, i_8_384_1892_0, i_8_384_1936_0, i_8_384_1954_0,
    i_8_384_1958_0, i_8_384_1975_0, i_8_384_1976_0, i_8_384_1985_0,
    i_8_384_1992_0, i_8_384_2044_0, i_8_384_2146_0, i_8_384_2155_0,
    i_8_384_2227_0, i_8_384_2231_0, i_8_384_2246_0, i_8_384_2257_0;
  output o_8_384_0_0;
  assign o_8_384_0_0 = 0;
endmodule



// Benchmark "kernel_8_385" written by ABC on Sun Jul 19 10:09:47 2020

module kernel_8_385 ( 
    i_8_385_20_0, i_8_385_35_0, i_8_385_85_0, i_8_385_94_0, i_8_385_224_0,
    i_8_385_264_0, i_8_385_269_0, i_8_385_323_0, i_8_385_356_0,
    i_8_385_370_0, i_8_385_445_0, i_8_385_453_0, i_8_385_460_0,
    i_8_385_506_0, i_8_385_538_0, i_8_385_554_0, i_8_385_556_0,
    i_8_385_565_0, i_8_385_620_0, i_8_385_647_0, i_8_385_658_0,
    i_8_385_662_0, i_8_385_698_0, i_8_385_708_0, i_8_385_718_0,
    i_8_385_721_0, i_8_385_733_0, i_8_385_734_0, i_8_385_779_0,
    i_8_385_793_0, i_8_385_843_0, i_8_385_923_0, i_8_385_935_0,
    i_8_385_950_0, i_8_385_953_0, i_8_385_977_0, i_8_385_988_0,
    i_8_385_989_0, i_8_385_994_0, i_8_385_997_0, i_8_385_998_0,
    i_8_385_1060_0, i_8_385_1105_0, i_8_385_1139_0, i_8_385_1183_0,
    i_8_385_1203_0, i_8_385_1234_0, i_8_385_1259_0, i_8_385_1260_0,
    i_8_385_1261_0, i_8_385_1268_0, i_8_385_1282_0, i_8_385_1283_0,
    i_8_385_1286_0, i_8_385_1319_0, i_8_385_1321_0, i_8_385_1325_0,
    i_8_385_1327_0, i_8_385_1328_0, i_8_385_1332_0, i_8_385_1366_0,
    i_8_385_1416_0, i_8_385_1418_0, i_8_385_1450_0, i_8_385_1452_0,
    i_8_385_1470_0, i_8_385_1481_0, i_8_385_1526_0, i_8_385_1532_0,
    i_8_385_1538_0, i_8_385_1553_0, i_8_385_1603_0, i_8_385_1604_0,
    i_8_385_1723_0, i_8_385_1754_0, i_8_385_1770_0, i_8_385_1771_0,
    i_8_385_1772_0, i_8_385_1788_0, i_8_385_1796_0, i_8_385_1813_0,
    i_8_385_1823_0, i_8_385_1931_0, i_8_385_1964_0, i_8_385_1983_0,
    i_8_385_1988_0, i_8_385_1989_0, i_8_385_2042_0, i_8_385_2067_0,
    i_8_385_2069_0, i_8_385_2077_0, i_8_385_2078_0, i_8_385_2113_0,
    i_8_385_2114_0, i_8_385_2136_0, i_8_385_2218_0, i_8_385_2226_0,
    i_8_385_2264_0, i_8_385_2294_0, i_8_385_2299_0,
    o_8_385_0_0  );
  input  i_8_385_20_0, i_8_385_35_0, i_8_385_85_0, i_8_385_94_0,
    i_8_385_224_0, i_8_385_264_0, i_8_385_269_0, i_8_385_323_0,
    i_8_385_356_0, i_8_385_370_0, i_8_385_445_0, i_8_385_453_0,
    i_8_385_460_0, i_8_385_506_0, i_8_385_538_0, i_8_385_554_0,
    i_8_385_556_0, i_8_385_565_0, i_8_385_620_0, i_8_385_647_0,
    i_8_385_658_0, i_8_385_662_0, i_8_385_698_0, i_8_385_708_0,
    i_8_385_718_0, i_8_385_721_0, i_8_385_733_0, i_8_385_734_0,
    i_8_385_779_0, i_8_385_793_0, i_8_385_843_0, i_8_385_923_0,
    i_8_385_935_0, i_8_385_950_0, i_8_385_953_0, i_8_385_977_0,
    i_8_385_988_0, i_8_385_989_0, i_8_385_994_0, i_8_385_997_0,
    i_8_385_998_0, i_8_385_1060_0, i_8_385_1105_0, i_8_385_1139_0,
    i_8_385_1183_0, i_8_385_1203_0, i_8_385_1234_0, i_8_385_1259_0,
    i_8_385_1260_0, i_8_385_1261_0, i_8_385_1268_0, i_8_385_1282_0,
    i_8_385_1283_0, i_8_385_1286_0, i_8_385_1319_0, i_8_385_1321_0,
    i_8_385_1325_0, i_8_385_1327_0, i_8_385_1328_0, i_8_385_1332_0,
    i_8_385_1366_0, i_8_385_1416_0, i_8_385_1418_0, i_8_385_1450_0,
    i_8_385_1452_0, i_8_385_1470_0, i_8_385_1481_0, i_8_385_1526_0,
    i_8_385_1532_0, i_8_385_1538_0, i_8_385_1553_0, i_8_385_1603_0,
    i_8_385_1604_0, i_8_385_1723_0, i_8_385_1754_0, i_8_385_1770_0,
    i_8_385_1771_0, i_8_385_1772_0, i_8_385_1788_0, i_8_385_1796_0,
    i_8_385_1813_0, i_8_385_1823_0, i_8_385_1931_0, i_8_385_1964_0,
    i_8_385_1983_0, i_8_385_1988_0, i_8_385_1989_0, i_8_385_2042_0,
    i_8_385_2067_0, i_8_385_2069_0, i_8_385_2077_0, i_8_385_2078_0,
    i_8_385_2113_0, i_8_385_2114_0, i_8_385_2136_0, i_8_385_2218_0,
    i_8_385_2226_0, i_8_385_2264_0, i_8_385_2294_0, i_8_385_2299_0;
  output o_8_385_0_0;
  assign o_8_385_0_0 = 0;
endmodule



// Benchmark "kernel_8_386" written by ABC on Sun Jul 19 10:09:47 2020

module kernel_8_386 ( 
    i_8_386_19_0, i_8_386_31_0, i_8_386_32_0, i_8_386_54_0, i_8_386_55_0,
    i_8_386_81_0, i_8_386_84_0, i_8_386_100_0, i_8_386_107_0,
    i_8_386_117_0, i_8_386_205_0, i_8_386_255_0, i_8_386_256_0,
    i_8_386_297_0, i_8_386_304_0, i_8_386_423_0, i_8_386_495_0,
    i_8_386_502_0, i_8_386_530_0, i_8_386_549_0, i_8_386_554_0,
    i_8_386_576_0, i_8_386_586_0, i_8_386_589_0, i_8_386_603_0,
    i_8_386_606_0, i_8_386_607_0, i_8_386_627_0, i_8_386_628_0,
    i_8_386_631_0, i_8_386_632_0, i_8_386_677_0, i_8_386_703_0,
    i_8_386_730_0, i_8_386_735_0, i_8_386_764_0, i_8_386_823_0,
    i_8_386_846_0, i_8_386_855_0, i_8_386_864_0, i_8_386_865_0,
    i_8_386_882_0, i_8_386_883_0, i_8_386_945_0, i_8_386_948_0,
    i_8_386_1033_0, i_8_386_1034_0, i_8_386_1062_0, i_8_386_1063_0,
    i_8_386_1111_0, i_8_386_1125_0, i_8_386_1134_0, i_8_386_1143_0,
    i_8_386_1144_0, i_8_386_1152_0, i_8_386_1171_0, i_8_386_1226_0,
    i_8_386_1233_0, i_8_386_1297_0, i_8_386_1299_0, i_8_386_1305_0,
    i_8_386_1332_0, i_8_386_1333_0, i_8_386_1403_0, i_8_386_1431_0,
    i_8_386_1432_0, i_8_386_1436_0, i_8_386_1467_0, i_8_386_1530_0,
    i_8_386_1543_0, i_8_386_1602_0, i_8_386_1615_0, i_8_386_1623_0,
    i_8_386_1631_0, i_8_386_1650_0, i_8_386_1652_0, i_8_386_1660_0,
    i_8_386_1693_0, i_8_386_1702_0, i_8_386_1710_0, i_8_386_1747_0,
    i_8_386_1755_0, i_8_386_1756_0, i_8_386_1762_0, i_8_386_1774_0,
    i_8_386_1776_0, i_8_386_1793_0, i_8_386_1809_0, i_8_386_1815_0,
    i_8_386_1872_0, i_8_386_1963_0, i_8_386_1980_0, i_8_386_2137_0,
    i_8_386_2143_0, i_8_386_2151_0, i_8_386_2196_0, i_8_386_2224_0,
    i_8_386_2234_0, i_8_386_2242_0, i_8_386_2245_0,
    o_8_386_0_0  );
  input  i_8_386_19_0, i_8_386_31_0, i_8_386_32_0, i_8_386_54_0,
    i_8_386_55_0, i_8_386_81_0, i_8_386_84_0, i_8_386_100_0, i_8_386_107_0,
    i_8_386_117_0, i_8_386_205_0, i_8_386_255_0, i_8_386_256_0,
    i_8_386_297_0, i_8_386_304_0, i_8_386_423_0, i_8_386_495_0,
    i_8_386_502_0, i_8_386_530_0, i_8_386_549_0, i_8_386_554_0,
    i_8_386_576_0, i_8_386_586_0, i_8_386_589_0, i_8_386_603_0,
    i_8_386_606_0, i_8_386_607_0, i_8_386_627_0, i_8_386_628_0,
    i_8_386_631_0, i_8_386_632_0, i_8_386_677_0, i_8_386_703_0,
    i_8_386_730_0, i_8_386_735_0, i_8_386_764_0, i_8_386_823_0,
    i_8_386_846_0, i_8_386_855_0, i_8_386_864_0, i_8_386_865_0,
    i_8_386_882_0, i_8_386_883_0, i_8_386_945_0, i_8_386_948_0,
    i_8_386_1033_0, i_8_386_1034_0, i_8_386_1062_0, i_8_386_1063_0,
    i_8_386_1111_0, i_8_386_1125_0, i_8_386_1134_0, i_8_386_1143_0,
    i_8_386_1144_0, i_8_386_1152_0, i_8_386_1171_0, i_8_386_1226_0,
    i_8_386_1233_0, i_8_386_1297_0, i_8_386_1299_0, i_8_386_1305_0,
    i_8_386_1332_0, i_8_386_1333_0, i_8_386_1403_0, i_8_386_1431_0,
    i_8_386_1432_0, i_8_386_1436_0, i_8_386_1467_0, i_8_386_1530_0,
    i_8_386_1543_0, i_8_386_1602_0, i_8_386_1615_0, i_8_386_1623_0,
    i_8_386_1631_0, i_8_386_1650_0, i_8_386_1652_0, i_8_386_1660_0,
    i_8_386_1693_0, i_8_386_1702_0, i_8_386_1710_0, i_8_386_1747_0,
    i_8_386_1755_0, i_8_386_1756_0, i_8_386_1762_0, i_8_386_1774_0,
    i_8_386_1776_0, i_8_386_1793_0, i_8_386_1809_0, i_8_386_1815_0,
    i_8_386_1872_0, i_8_386_1963_0, i_8_386_1980_0, i_8_386_2137_0,
    i_8_386_2143_0, i_8_386_2151_0, i_8_386_2196_0, i_8_386_2224_0,
    i_8_386_2234_0, i_8_386_2242_0, i_8_386_2245_0;
  output o_8_386_0_0;
  assign o_8_386_0_0 = 0;
endmodule



// Benchmark "kernel_8_387" written by ABC on Sun Jul 19 10:09:48 2020

module kernel_8_387 ( 
    i_8_387_14_0, i_8_387_30_0, i_8_387_98_0, i_8_387_102_0, i_8_387_103_0,
    i_8_387_107_0, i_8_387_114_0, i_8_387_216_0, i_8_387_223_0,
    i_8_387_297_0, i_8_387_300_0, i_8_387_345_0, i_8_387_361_0,
    i_8_387_362_0, i_8_387_365_0, i_8_387_367_0, i_8_387_391_0,
    i_8_387_418_0, i_8_387_444_0, i_8_387_453_0, i_8_387_525_0,
    i_8_387_530_0, i_8_387_535_0, i_8_387_546_0, i_8_387_552_0,
    i_8_387_589_0, i_8_387_591_0, i_8_387_607_0, i_8_387_609_0,
    i_8_387_630_0, i_8_387_637_0, i_8_387_659_0, i_8_387_665_0,
    i_8_387_694_0, i_8_387_697_0, i_8_387_723_0, i_8_387_738_0,
    i_8_387_780_0, i_8_387_781_0, i_8_387_786_0, i_8_387_822_0,
    i_8_387_842_0, i_8_387_874_0, i_8_387_894_0, i_8_387_958_0,
    i_8_387_970_0, i_8_387_987_0, i_8_387_1071_0, i_8_387_1107_0,
    i_8_387_1138_0, i_8_387_1145_0, i_8_387_1159_0, i_8_387_1204_0,
    i_8_387_1227_0, i_8_387_1228_0, i_8_387_1264_0, i_8_387_1279_0,
    i_8_387_1282_0, i_8_387_1285_0, i_8_387_1344_0, i_8_387_1426_0,
    i_8_387_1437_0, i_8_387_1438_0, i_8_387_1461_0, i_8_387_1525_0,
    i_8_387_1542_0, i_8_387_1552_0, i_8_387_1563_0, i_8_387_1564_0,
    i_8_387_1614_0, i_8_387_1635_0, i_8_387_1668_0, i_8_387_1681_0,
    i_8_387_1701_0, i_8_387_1719_0, i_8_387_1749_0, i_8_387_1761_0,
    i_8_387_1765_0, i_8_387_1773_0, i_8_387_1780_0, i_8_387_1782_0,
    i_8_387_1785_0, i_8_387_1786_0, i_8_387_1815_0, i_8_387_1843_0,
    i_8_387_2109_0, i_8_387_2110_0, i_8_387_2134_0, i_8_387_2139_0,
    i_8_387_2147_0, i_8_387_2157_0, i_8_387_2158_0, i_8_387_2184_0,
    i_8_387_2190_0, i_8_387_2215_0, i_8_387_2226_0, i_8_387_2232_0,
    i_8_387_2233_0, i_8_387_2265_0, i_8_387_2287_0,
    o_8_387_0_0  );
  input  i_8_387_14_0, i_8_387_30_0, i_8_387_98_0, i_8_387_102_0,
    i_8_387_103_0, i_8_387_107_0, i_8_387_114_0, i_8_387_216_0,
    i_8_387_223_0, i_8_387_297_0, i_8_387_300_0, i_8_387_345_0,
    i_8_387_361_0, i_8_387_362_0, i_8_387_365_0, i_8_387_367_0,
    i_8_387_391_0, i_8_387_418_0, i_8_387_444_0, i_8_387_453_0,
    i_8_387_525_0, i_8_387_530_0, i_8_387_535_0, i_8_387_546_0,
    i_8_387_552_0, i_8_387_589_0, i_8_387_591_0, i_8_387_607_0,
    i_8_387_609_0, i_8_387_630_0, i_8_387_637_0, i_8_387_659_0,
    i_8_387_665_0, i_8_387_694_0, i_8_387_697_0, i_8_387_723_0,
    i_8_387_738_0, i_8_387_780_0, i_8_387_781_0, i_8_387_786_0,
    i_8_387_822_0, i_8_387_842_0, i_8_387_874_0, i_8_387_894_0,
    i_8_387_958_0, i_8_387_970_0, i_8_387_987_0, i_8_387_1071_0,
    i_8_387_1107_0, i_8_387_1138_0, i_8_387_1145_0, i_8_387_1159_0,
    i_8_387_1204_0, i_8_387_1227_0, i_8_387_1228_0, i_8_387_1264_0,
    i_8_387_1279_0, i_8_387_1282_0, i_8_387_1285_0, i_8_387_1344_0,
    i_8_387_1426_0, i_8_387_1437_0, i_8_387_1438_0, i_8_387_1461_0,
    i_8_387_1525_0, i_8_387_1542_0, i_8_387_1552_0, i_8_387_1563_0,
    i_8_387_1564_0, i_8_387_1614_0, i_8_387_1635_0, i_8_387_1668_0,
    i_8_387_1681_0, i_8_387_1701_0, i_8_387_1719_0, i_8_387_1749_0,
    i_8_387_1761_0, i_8_387_1765_0, i_8_387_1773_0, i_8_387_1780_0,
    i_8_387_1782_0, i_8_387_1785_0, i_8_387_1786_0, i_8_387_1815_0,
    i_8_387_1843_0, i_8_387_2109_0, i_8_387_2110_0, i_8_387_2134_0,
    i_8_387_2139_0, i_8_387_2147_0, i_8_387_2157_0, i_8_387_2158_0,
    i_8_387_2184_0, i_8_387_2190_0, i_8_387_2215_0, i_8_387_2226_0,
    i_8_387_2232_0, i_8_387_2233_0, i_8_387_2265_0, i_8_387_2287_0;
  output o_8_387_0_0;
  assign o_8_387_0_0 = 0;
endmodule



// Benchmark "kernel_8_388" written by ABC on Sun Jul 19 10:09:50 2020

module kernel_8_388 ( 
    i_8_388_4_0, i_8_388_7_0, i_8_388_86_0, i_8_388_89_0, i_8_388_121_0,
    i_8_388_151_0, i_8_388_197_0, i_8_388_202_0, i_8_388_214_0,
    i_8_388_220_0, i_8_388_247_0, i_8_388_248_0, i_8_388_301_0,
    i_8_388_342_0, i_8_388_346_0, i_8_388_367_0, i_8_388_376_0,
    i_8_388_400_0, i_8_388_401_0, i_8_388_440_0, i_8_388_455_0,
    i_8_388_516_0, i_8_388_517_0, i_8_388_527_0, i_8_388_529_0,
    i_8_388_530_0, i_8_388_571_0, i_8_388_659_0, i_8_388_683_0,
    i_8_388_688_0, i_8_388_699_0, i_8_388_701_0, i_8_388_727_0,
    i_8_388_728_0, i_8_388_763_0, i_8_388_781_0, i_8_388_815_0,
    i_8_388_818_0, i_8_388_835_0, i_8_388_862_0, i_8_388_982_0,
    i_8_388_985_0, i_8_388_1003_0, i_8_388_1004_0, i_8_388_1045_0,
    i_8_388_1114_0, i_8_388_1153_0, i_8_388_1155_0, i_8_388_1157_0,
    i_8_388_1186_0, i_8_388_1281_0, i_8_388_1328_0, i_8_388_1330_0,
    i_8_388_1331_0, i_8_388_1342_0, i_8_388_1344_0, i_8_388_1358_0,
    i_8_388_1365_0, i_8_388_1434_0, i_8_388_1473_0, i_8_388_1474_0,
    i_8_388_1490_0, i_8_388_1535_0, i_8_388_1565_0, i_8_388_1610_0,
    i_8_388_1634_0, i_8_388_1642_0, i_8_388_1661_0, i_8_388_1662_0,
    i_8_388_1732_0, i_8_388_1733_0, i_8_388_1750_0, i_8_388_1753_0,
    i_8_388_1786_0, i_8_388_1787_0, i_8_388_1804_0, i_8_388_1806_0,
    i_8_388_1807_0, i_8_388_1840_0, i_8_388_1858_0, i_8_388_1861_0,
    i_8_388_1885_0, i_8_388_1975_0, i_8_388_1997_0, i_8_388_2011_0,
    i_8_388_2012_0, i_8_388_2032_0, i_8_388_2113_0, i_8_388_2120_0,
    i_8_388_2122_0, i_8_388_2123_0, i_8_388_2159_0, i_8_388_2174_0,
    i_8_388_2200_0, i_8_388_2215_0, i_8_388_2216_0, i_8_388_2225_0,
    i_8_388_2254_0, i_8_388_2289_0, i_8_388_2294_0,
    o_8_388_0_0  );
  input  i_8_388_4_0, i_8_388_7_0, i_8_388_86_0, i_8_388_89_0,
    i_8_388_121_0, i_8_388_151_0, i_8_388_197_0, i_8_388_202_0,
    i_8_388_214_0, i_8_388_220_0, i_8_388_247_0, i_8_388_248_0,
    i_8_388_301_0, i_8_388_342_0, i_8_388_346_0, i_8_388_367_0,
    i_8_388_376_0, i_8_388_400_0, i_8_388_401_0, i_8_388_440_0,
    i_8_388_455_0, i_8_388_516_0, i_8_388_517_0, i_8_388_527_0,
    i_8_388_529_0, i_8_388_530_0, i_8_388_571_0, i_8_388_659_0,
    i_8_388_683_0, i_8_388_688_0, i_8_388_699_0, i_8_388_701_0,
    i_8_388_727_0, i_8_388_728_0, i_8_388_763_0, i_8_388_781_0,
    i_8_388_815_0, i_8_388_818_0, i_8_388_835_0, i_8_388_862_0,
    i_8_388_982_0, i_8_388_985_0, i_8_388_1003_0, i_8_388_1004_0,
    i_8_388_1045_0, i_8_388_1114_0, i_8_388_1153_0, i_8_388_1155_0,
    i_8_388_1157_0, i_8_388_1186_0, i_8_388_1281_0, i_8_388_1328_0,
    i_8_388_1330_0, i_8_388_1331_0, i_8_388_1342_0, i_8_388_1344_0,
    i_8_388_1358_0, i_8_388_1365_0, i_8_388_1434_0, i_8_388_1473_0,
    i_8_388_1474_0, i_8_388_1490_0, i_8_388_1535_0, i_8_388_1565_0,
    i_8_388_1610_0, i_8_388_1634_0, i_8_388_1642_0, i_8_388_1661_0,
    i_8_388_1662_0, i_8_388_1732_0, i_8_388_1733_0, i_8_388_1750_0,
    i_8_388_1753_0, i_8_388_1786_0, i_8_388_1787_0, i_8_388_1804_0,
    i_8_388_1806_0, i_8_388_1807_0, i_8_388_1840_0, i_8_388_1858_0,
    i_8_388_1861_0, i_8_388_1885_0, i_8_388_1975_0, i_8_388_1997_0,
    i_8_388_2011_0, i_8_388_2012_0, i_8_388_2032_0, i_8_388_2113_0,
    i_8_388_2120_0, i_8_388_2122_0, i_8_388_2123_0, i_8_388_2159_0,
    i_8_388_2174_0, i_8_388_2200_0, i_8_388_2215_0, i_8_388_2216_0,
    i_8_388_2225_0, i_8_388_2254_0, i_8_388_2289_0, i_8_388_2294_0;
  output o_8_388_0_0;
  assign o_8_388_0_0 = ~((~i_8_388_2120_0 & ((~i_8_388_728_0 & ((~i_8_388_121_0 & ~i_8_388_781_0 & ((~i_8_388_342_0 & ~i_8_388_367_0 & ~i_8_388_527_0 & ~i_8_388_815_0 & ~i_8_388_1330_0 & ~i_8_388_1661_0 & ~i_8_388_1885_0 & ~i_8_388_2032_0) | (~i_8_388_214_0 & ~i_8_388_247_0 & ~i_8_388_516_0 & ~i_8_388_517_0 & ~i_8_388_683_0 & ~i_8_388_701_0 & ~i_8_388_982_0 & ~i_8_388_1490_0 & ~i_8_388_1806_0 & ~i_8_388_2122_0 & ~i_8_388_2123_0 & ~i_8_388_2174_0 & ~i_8_388_2200_0))) | (~i_8_388_214_0 & i_8_388_376_0 & ~i_8_388_516_0 & ~i_8_388_530_0 & ~i_8_388_571_0 & ~i_8_388_688_0 & ~i_8_388_1045_0 & ~i_8_388_1661_0 & ~i_8_388_1732_0 & ~i_8_388_1733_0 & ~i_8_388_2122_0 & ~i_8_388_2123_0))) | (~i_8_388_151_0 & ((~i_8_388_202_0 & ~i_8_388_1733_0 & ((~i_8_388_455_0 & ~i_8_388_571_0 & ~i_8_388_699_0 & ~i_8_388_701_0 & ~i_8_388_727_0 & ~i_8_388_818_0 & ~i_8_388_1358_0 & ~i_8_388_1365_0 & ~i_8_388_2011_0 & ~i_8_388_2123_0) | (~i_8_388_197_0 & ~i_8_388_247_0 & i_8_388_529_0 & ~i_8_388_985_0 & ~i_8_388_1186_0 & ~i_8_388_1858_0 & ~i_8_388_2012_0 & ~i_8_388_2032_0 & ~i_8_388_2216_0 & ~i_8_388_2294_0))) | (~i_8_388_440_0 & ~i_8_388_985_0 & ((~i_8_388_248_0 & ~i_8_388_301_0 & ~i_8_388_517_0 & ~i_8_388_763_0 & ~i_8_388_835_0 & ~i_8_388_982_0 & ~i_8_388_1365_0 & ~i_8_388_1473_0 & ~i_8_388_1490_0 & ~i_8_388_1662_0 & ~i_8_388_1806_0 & ~i_8_388_1997_0) | (~i_8_388_214_0 & ~i_8_388_688_0 & ~i_8_388_727_0 & ~i_8_388_815_0 & ~i_8_388_1004_0 & ~i_8_388_2011_0 & ~i_8_388_2122_0 & ~i_8_388_2123_0 & ~i_8_388_2254_0))))) | (~i_8_388_2032_0 & ((~i_8_388_1733_0 & ((~i_8_388_7_0 & ~i_8_388_440_0 & ~i_8_388_699_0 & ~i_8_388_818_0 & ~i_8_388_1186_0 & ~i_8_388_1661_0 & ~i_8_388_1732_0 & ~i_8_388_1885_0 & ~i_8_388_2012_0) | (i_8_388_1434_0 & ~i_8_388_1610_0 & ~i_8_388_2122_0 & ~i_8_388_2254_0))) | (~i_8_388_248_0 & ~i_8_388_516_0 & ~i_8_388_571_0 & ~i_8_388_688_0 & ~i_8_388_985_0 & i_8_388_1114_0 & ~i_8_388_1662_0 & i_8_388_1753_0 & i_8_388_1804_0 & ~i_8_388_2012_0 & ~i_8_388_2123_0))))) | (~i_8_388_89_0 & ((~i_8_388_818_0 & ((~i_8_388_2012_0 & ((~i_8_388_4_0 & ~i_8_388_151_0 & ~i_8_388_2123_0 & ((~i_8_388_7_0 & ~i_8_388_516_0 & ~i_8_388_683_0 & ~i_8_388_701_0 & ~i_8_388_835_0 & ~i_8_388_1661_0 & ~i_8_388_1807_0 & ~i_8_388_1997_0 & ~i_8_388_2122_0 & ~i_8_388_2174_0) | (~i_8_388_727_0 & ~i_8_388_763_0 & ~i_8_388_862_0 & ~i_8_388_985_0 & ~i_8_388_1662_0 & ~i_8_388_1733_0 & ~i_8_388_2011_0 & ~i_8_388_2216_0))) | (~i_8_388_7_0 & ~i_8_388_121_0 & ~i_8_388_197_0 & ~i_8_388_214_0 & ~i_8_388_1342_0 & ~i_8_388_1358_0 & ~i_8_388_1490_0 & ~i_8_388_1662_0 & ~i_8_388_2122_0 & ~i_8_388_2216_0))) | (~i_8_388_376_0 & ~i_8_388_401_0 & ~i_8_388_527_0 & ~i_8_388_728_0 & ~i_8_388_835_0 & ~i_8_388_1806_0 & ~i_8_388_1858_0 & ~i_8_388_1861_0 & ~i_8_388_2011_0 & ~i_8_388_2294_0))) | (~i_8_388_121_0 & ~i_8_388_376_0 & ~i_8_388_571_0 & ~i_8_388_835_0 & ~i_8_388_1358_0 & ~i_8_388_1661_0 & ~i_8_388_1997_0 & ~i_8_388_2032_0 & ~i_8_388_2254_0))) | (~i_8_388_2011_0 & ((~i_8_388_4_0 & ~i_8_388_197_0 & ((~i_8_388_376_0 & ~i_8_388_530_0 & ~i_8_388_683_0 & ~i_8_388_763_0 & ~i_8_388_1358_0 & ~i_8_388_1365_0 & i_8_388_1804_0 & ~i_8_388_2122_0 & ~i_8_388_2174_0) | (~i_8_388_7_0 & ~i_8_388_248_0 & ~i_8_388_818_0 & ~i_8_388_1003_0 & i_8_388_1114_0 & ~i_8_388_2123_0 & ~i_8_388_2200_0))) | (~i_8_388_815_0 & ~i_8_388_2012_0 & ((~i_8_388_151_0 & ~i_8_388_220_0 & ~i_8_388_440_0 & ~i_8_388_517_0 & ~i_8_388_763_0 & ~i_8_388_1535_0 & ~i_8_388_1750_0 & ~i_8_388_1753_0 & ~i_8_388_1804_0 & ~i_8_388_2123_0 & ~i_8_388_2215_0) | (~i_8_388_247_0 & ~i_8_388_659_0 & ~i_8_388_835_0 & ~i_8_388_1186_0 & ~i_8_388_1885_0 & ~i_8_388_1997_0 & ~i_8_388_2032_0 & ~i_8_388_2122_0 & ~i_8_388_2159_0 & ~i_8_388_2225_0))) | (i_8_388_220_0 & ~i_8_388_248_0 & ~i_8_388_516_0 & ~i_8_388_1114_0 & ~i_8_388_2122_0 & ~i_8_388_2174_0 & ~i_8_388_1358_0 & ~i_8_388_1365_0))) | (~i_8_388_151_0 & ((~i_8_388_517_0 & ~i_8_388_818_0 & ~i_8_388_1003_0 & ~i_8_388_1186_0 & ~i_8_388_1662_0 & i_8_388_1786_0 & ~i_8_388_2174_0) | (~i_8_388_763_0 & i_8_388_1281_0 & ~i_8_388_1344_0 & ~i_8_388_1365_0 & ~i_8_388_2032_0 & ~i_8_388_2254_0 & ~i_8_388_1732_0 & ~i_8_388_1858_0))) | (~i_8_388_247_0 & ((~i_8_388_4_0 & ~i_8_388_376_0 & ~i_8_388_688_0 & ~i_8_388_699_0 & ~i_8_388_727_0 & ~i_8_388_728_0 & ~i_8_388_1045_0 & ~i_8_388_1610_0 & ~i_8_388_1642_0 & ~i_8_388_1661_0 & i_8_388_1753_0 & ~i_8_388_2032_0) | (~i_8_388_530_0 & ~i_8_388_763_0 & ~i_8_388_835_0 & ~i_8_388_2012_0 & ~i_8_388_2123_0 & ~i_8_388_1732_0 & i_8_388_1787_0))) | (~i_8_388_2012_0 & ((~i_8_388_86_0 & i_8_388_248_0 & ~i_8_388_1003_0 & i_8_388_1750_0) | (~i_8_388_248_0 & ~i_8_388_516_0 & ~i_8_388_530_0 & ~i_8_388_699_0 & ~i_8_388_818_0 & ~i_8_388_1490_0 & ~i_8_388_1661_0 & ~i_8_388_1806_0 & ~i_8_388_1885_0 & ~i_8_388_2113_0))) | (~i_8_388_86_0 & ((~i_8_388_220_0 & ~i_8_388_763_0 & i_8_388_1331_0 & ~i_8_388_1997_0) | (~i_8_388_835_0 & ~i_8_388_982_0 & i_8_388_1330_0 & ~i_8_388_2032_0 & ~i_8_388_2122_0 & ~i_8_388_2123_0))));
endmodule



// Benchmark "kernel_8_389" written by ABC on Sun Jul 19 10:09:51 2020

module kernel_8_389 ( 
    i_8_389_47_0, i_8_389_92_0, i_8_389_101_0, i_8_389_112_0,
    i_8_389_164_0, i_8_389_172_0, i_8_389_226_0, i_8_389_232_0,
    i_8_389_307_0, i_8_389_308_0, i_8_389_334_0, i_8_389_335_0,
    i_8_389_345_0, i_8_389_350_0, i_8_389_352_0, i_8_389_353_0,
    i_8_389_362_0, i_8_389_374_0, i_8_389_380_0, i_8_389_418_0,
    i_8_389_424_0, i_8_389_451_0, i_8_389_452_0, i_8_389_479_0,
    i_8_389_488_0, i_8_389_550_0, i_8_389_551_0, i_8_389_568_0,
    i_8_389_685_0, i_8_389_695_0, i_8_389_703_0, i_8_389_796_0,
    i_8_389_805_0, i_8_389_928_0, i_8_389_1018_0, i_8_389_1035_0,
    i_8_389_1054_0, i_8_389_1055_0, i_8_389_1057_0, i_8_389_1099_0,
    i_8_389_1100_0, i_8_389_1181_0, i_8_389_1229_0, i_8_389_1253_0,
    i_8_389_1274_0, i_8_389_1280_0, i_8_389_1289_0, i_8_389_1292_0,
    i_8_389_1297_0, i_8_389_1309_0, i_8_389_1315_0, i_8_389_1370_0,
    i_8_389_1378_0, i_8_389_1379_0, i_8_389_1381_0, i_8_389_1382_0,
    i_8_389_1408_0, i_8_389_1436_0, i_8_389_1443_0, i_8_389_1521_0,
    i_8_389_1549_0, i_8_389_1558_0, i_8_389_1559_0, i_8_389_1562_0,
    i_8_389_1603_0, i_8_389_1607_0, i_8_389_1624_0, i_8_389_1639_0,
    i_8_389_1640_0, i_8_389_1649_0, i_8_389_1650_0, i_8_389_1694_0,
    i_8_389_1702_0, i_8_389_1703_0, i_8_389_1752_0, i_8_389_1804_0,
    i_8_389_1820_0, i_8_389_1822_0, i_8_389_1829_0, i_8_389_1847_0,
    i_8_389_1855_0, i_8_389_1937_0, i_8_389_2002_0, i_8_389_2035_0,
    i_8_389_2036_0, i_8_389_2063_0, i_8_389_2072_0, i_8_389_2107_0,
    i_8_389_2143_0, i_8_389_2144_0, i_8_389_2152_0, i_8_389_2153_0,
    i_8_389_2197_0, i_8_389_2198_0, i_8_389_2207_0, i_8_389_2215_0,
    i_8_389_2225_0, i_8_389_2241_0, i_8_389_2245_0, i_8_389_2287_0,
    o_8_389_0_0  );
  input  i_8_389_47_0, i_8_389_92_0, i_8_389_101_0, i_8_389_112_0,
    i_8_389_164_0, i_8_389_172_0, i_8_389_226_0, i_8_389_232_0,
    i_8_389_307_0, i_8_389_308_0, i_8_389_334_0, i_8_389_335_0,
    i_8_389_345_0, i_8_389_350_0, i_8_389_352_0, i_8_389_353_0,
    i_8_389_362_0, i_8_389_374_0, i_8_389_380_0, i_8_389_418_0,
    i_8_389_424_0, i_8_389_451_0, i_8_389_452_0, i_8_389_479_0,
    i_8_389_488_0, i_8_389_550_0, i_8_389_551_0, i_8_389_568_0,
    i_8_389_685_0, i_8_389_695_0, i_8_389_703_0, i_8_389_796_0,
    i_8_389_805_0, i_8_389_928_0, i_8_389_1018_0, i_8_389_1035_0,
    i_8_389_1054_0, i_8_389_1055_0, i_8_389_1057_0, i_8_389_1099_0,
    i_8_389_1100_0, i_8_389_1181_0, i_8_389_1229_0, i_8_389_1253_0,
    i_8_389_1274_0, i_8_389_1280_0, i_8_389_1289_0, i_8_389_1292_0,
    i_8_389_1297_0, i_8_389_1309_0, i_8_389_1315_0, i_8_389_1370_0,
    i_8_389_1378_0, i_8_389_1379_0, i_8_389_1381_0, i_8_389_1382_0,
    i_8_389_1408_0, i_8_389_1436_0, i_8_389_1443_0, i_8_389_1521_0,
    i_8_389_1549_0, i_8_389_1558_0, i_8_389_1559_0, i_8_389_1562_0,
    i_8_389_1603_0, i_8_389_1607_0, i_8_389_1624_0, i_8_389_1639_0,
    i_8_389_1640_0, i_8_389_1649_0, i_8_389_1650_0, i_8_389_1694_0,
    i_8_389_1702_0, i_8_389_1703_0, i_8_389_1752_0, i_8_389_1804_0,
    i_8_389_1820_0, i_8_389_1822_0, i_8_389_1829_0, i_8_389_1847_0,
    i_8_389_1855_0, i_8_389_1937_0, i_8_389_2002_0, i_8_389_2035_0,
    i_8_389_2036_0, i_8_389_2063_0, i_8_389_2072_0, i_8_389_2107_0,
    i_8_389_2143_0, i_8_389_2144_0, i_8_389_2152_0, i_8_389_2153_0,
    i_8_389_2197_0, i_8_389_2198_0, i_8_389_2207_0, i_8_389_2215_0,
    i_8_389_2225_0, i_8_389_2241_0, i_8_389_2245_0, i_8_389_2287_0;
  output o_8_389_0_0;
  assign o_8_389_0_0 = 0;
endmodule



// Benchmark "kernel_8_390" written by ABC on Sun Jul 19 10:09:52 2020

module kernel_8_390 ( 
    i_8_390_53_0, i_8_390_193_0, i_8_390_238_0, i_8_390_255_0,
    i_8_390_256_0, i_8_390_258_0, i_8_390_259_0, i_8_390_260_0,
    i_8_390_289_0, i_8_390_299_0, i_8_390_364_0, i_8_390_366_0,
    i_8_390_367_0, i_8_390_379_0, i_8_390_380_0, i_8_390_382_0,
    i_8_390_393_0, i_8_390_394_0, i_8_390_395_0, i_8_390_446_0,
    i_8_390_457_0, i_8_390_465_0, i_8_390_475_0, i_8_390_555_0,
    i_8_390_585_0, i_8_390_587_0, i_8_390_606_0, i_8_390_612_0,
    i_8_390_613_0, i_8_390_614_0, i_8_390_615_0, i_8_390_616_0,
    i_8_390_658_0, i_8_390_660_0, i_8_390_661_0, i_8_390_697_0,
    i_8_390_702_0, i_8_390_711_0, i_8_390_712_0, i_8_390_813_0,
    i_8_390_814_0, i_8_390_815_0, i_8_390_816_0, i_8_390_817_0,
    i_8_390_820_0, i_8_390_955_0, i_8_390_990_0, i_8_390_992_0,
    i_8_390_1026_0, i_8_390_1072_0, i_8_390_1074_0, i_8_390_1076_0,
    i_8_390_1077_0, i_8_390_1111_0, i_8_390_1112_0, i_8_390_1159_0,
    i_8_390_1230_0, i_8_390_1232_0, i_8_390_1260_0, i_8_390_1264_0,
    i_8_390_1268_0, i_8_390_1299_0, i_8_390_1455_0, i_8_390_1457_0,
    i_8_390_1491_0, i_8_390_1492_0, i_8_390_1539_0, i_8_390_1542_0,
    i_8_390_1543_0, i_8_390_1554_0, i_8_390_1601_0, i_8_390_1637_0,
    i_8_390_1650_0, i_8_390_1651_0, i_8_390_1652_0, i_8_390_1685_0,
    i_8_390_1700_0, i_8_390_1735_0, i_8_390_1779_0, i_8_390_1780_0,
    i_8_390_1896_0, i_8_390_1897_0, i_8_390_1898_0, i_8_390_1904_0,
    i_8_390_1915_0, i_8_390_2008_0, i_8_390_2031_0, i_8_390_2053_0,
    i_8_390_2077_0, i_8_390_2111_0, i_8_390_2127_0, i_8_390_2128_0,
    i_8_390_2130_0, i_8_390_2171_0, i_8_390_2187_0, i_8_390_2188_0,
    i_8_390_2189_0, i_8_390_2264_0, i_8_390_2267_0, i_8_390_2291_0,
    o_8_390_0_0  );
  input  i_8_390_53_0, i_8_390_193_0, i_8_390_238_0, i_8_390_255_0,
    i_8_390_256_0, i_8_390_258_0, i_8_390_259_0, i_8_390_260_0,
    i_8_390_289_0, i_8_390_299_0, i_8_390_364_0, i_8_390_366_0,
    i_8_390_367_0, i_8_390_379_0, i_8_390_380_0, i_8_390_382_0,
    i_8_390_393_0, i_8_390_394_0, i_8_390_395_0, i_8_390_446_0,
    i_8_390_457_0, i_8_390_465_0, i_8_390_475_0, i_8_390_555_0,
    i_8_390_585_0, i_8_390_587_0, i_8_390_606_0, i_8_390_612_0,
    i_8_390_613_0, i_8_390_614_0, i_8_390_615_0, i_8_390_616_0,
    i_8_390_658_0, i_8_390_660_0, i_8_390_661_0, i_8_390_697_0,
    i_8_390_702_0, i_8_390_711_0, i_8_390_712_0, i_8_390_813_0,
    i_8_390_814_0, i_8_390_815_0, i_8_390_816_0, i_8_390_817_0,
    i_8_390_820_0, i_8_390_955_0, i_8_390_990_0, i_8_390_992_0,
    i_8_390_1026_0, i_8_390_1072_0, i_8_390_1074_0, i_8_390_1076_0,
    i_8_390_1077_0, i_8_390_1111_0, i_8_390_1112_0, i_8_390_1159_0,
    i_8_390_1230_0, i_8_390_1232_0, i_8_390_1260_0, i_8_390_1264_0,
    i_8_390_1268_0, i_8_390_1299_0, i_8_390_1455_0, i_8_390_1457_0,
    i_8_390_1491_0, i_8_390_1492_0, i_8_390_1539_0, i_8_390_1542_0,
    i_8_390_1543_0, i_8_390_1554_0, i_8_390_1601_0, i_8_390_1637_0,
    i_8_390_1650_0, i_8_390_1651_0, i_8_390_1652_0, i_8_390_1685_0,
    i_8_390_1700_0, i_8_390_1735_0, i_8_390_1779_0, i_8_390_1780_0,
    i_8_390_1896_0, i_8_390_1897_0, i_8_390_1898_0, i_8_390_1904_0,
    i_8_390_1915_0, i_8_390_2008_0, i_8_390_2031_0, i_8_390_2053_0,
    i_8_390_2077_0, i_8_390_2111_0, i_8_390_2127_0, i_8_390_2128_0,
    i_8_390_2130_0, i_8_390_2171_0, i_8_390_2187_0, i_8_390_2188_0,
    i_8_390_2189_0, i_8_390_2264_0, i_8_390_2267_0, i_8_390_2291_0;
  output o_8_390_0_0;
  assign o_8_390_0_0 = ~((i_8_390_255_0 & ((~i_8_390_382_0 & ~i_8_390_394_0 & ~i_8_390_1491_0 & ~i_8_390_1492_0 & ~i_8_390_1542_0 & ~i_8_390_2128_0) | (~i_8_390_289_0 & i_8_390_364_0 & ~i_8_390_395_0 & i_8_390_615_0 & ~i_8_390_2188_0))) | (~i_8_390_711_0 & ((~i_8_390_1111_0 & ((i_8_390_299_0 & ((~i_8_390_606_0 & ~i_8_390_614_0 & ~i_8_390_697_0 & i_8_390_992_0 & ~i_8_390_1554_0) | (~i_8_390_379_0 & ~i_8_390_587_0 & i_8_390_2171_0 & ~i_8_390_2291_0))) | (~i_8_390_299_0 & ~i_8_390_585_0 & i_8_390_614_0 & ~i_8_390_1542_0 & ~i_8_390_1735_0 & ~i_8_390_2188_0))) | (~i_8_390_380_0 & ~i_8_390_1542_0 & ((~i_8_390_379_0 & i_8_390_612_0 & ~i_8_390_697_0 & ~i_8_390_1026_0 & ~i_8_390_1112_0 & ~i_8_390_1492_0 & ~i_8_390_1896_0 & ~i_8_390_2008_0) | (~i_8_390_364_0 & ~i_8_390_382_0 & i_8_390_661_0 & ~i_8_390_1780_0 & ~i_8_390_2130_0 & ~i_8_390_2187_0))) | (~i_8_390_393_0 & ((~i_8_390_394_0 & ~i_8_390_395_0 & ((~i_8_390_299_0 & ~i_8_390_585_0 & i_8_390_661_0 & ~i_8_390_697_0 & ~i_8_390_1264_0 & ~i_8_390_1897_0 & ~i_8_390_2127_0) | (i_8_390_367_0 & ~i_8_390_612_0 & i_8_390_1264_0 & ~i_8_390_1491_0 & ~i_8_390_2008_0 & ~i_8_390_2187_0 & ~i_8_390_2189_0))) | (i_8_390_606_0 & ~i_8_390_820_0 & i_8_390_990_0 & ~i_8_390_992_0 & ~i_8_390_1650_0 & ~i_8_390_2291_0))) | (~i_8_390_299_0 & ((~i_8_390_587_0 & ~i_8_390_1112_0 & ~i_8_390_1260_0 & ((i_8_390_1264_0 & ~i_8_390_1455_0 & ~i_8_390_1491_0) | (~i_8_390_255_0 & ~i_8_390_394_0 & ~i_8_390_585_0 & ~i_8_390_697_0 & ~i_8_390_712_0 & ~i_8_390_1539_0 & ~i_8_390_1700_0 & ~i_8_390_2077_0 & i_8_390_2128_0))) | (~i_8_390_238_0 & ~i_8_390_1077_0 & ~i_8_390_1455_0 & ~i_8_390_1457_0 & i_8_390_1651_0 & ~i_8_390_1898_0 & ~i_8_390_2077_0 & ~i_8_390_2130_0 & ~i_8_390_2187_0))) | (~i_8_390_606_0 & ~i_8_390_616_0 & ~i_8_390_697_0 & ~i_8_390_712_0 & ~i_8_390_820_0 & i_8_390_1264_0 & ~i_8_390_1491_0 & ~i_8_390_1898_0 & ~i_8_390_2128_0 & ~i_8_390_2188_0))) | (~i_8_390_2128_0 & ((~i_8_390_238_0 & ((~i_8_390_393_0 & ~i_8_390_394_0 & ~i_8_390_616_0 & i_8_390_1230_0 & ~i_8_390_1457_0 & ~i_8_390_1897_0) | (~i_8_390_366_0 & ~i_8_390_382_0 & ~i_8_390_395_0 & ~i_8_390_585_0 & i_8_390_616_0 & ~i_8_390_661_0 & ~i_8_390_1542_0 & ~i_8_390_2111_0))) | (~i_8_390_2187_0 & ((~i_8_390_393_0 & ~i_8_390_1554_0 & ((~i_8_390_380_0 & ~i_8_390_616_0 & i_8_390_711_0 & ~i_8_390_813_0 & ~i_8_390_955_0 & ~i_8_390_1539_0) | (~i_8_390_394_0 & ~i_8_390_395_0 & ~i_8_390_606_0 & i_8_390_616_0 & ~i_8_390_820_0 & ~i_8_390_1457_0 & ~i_8_390_2189_0))) | (i_8_390_702_0 & ~i_8_390_1077_0 & ~i_8_390_1112_0 & ~i_8_390_1268_0 & ~i_8_390_1455_0 & ~i_8_390_1492_0 & ~i_8_390_1539_0) | (~i_8_390_379_0 & ~i_8_390_465_0 & ~i_8_390_587_0 & i_8_390_658_0 & ~i_8_390_1260_0 & ~i_8_390_1542_0 & ~i_8_390_1700_0 & ~i_8_390_1896_0 & ~i_8_390_1915_0) | (~i_8_390_258_0 & ~i_8_390_299_0 & ~i_8_390_394_0 & i_8_390_1076_0 & ~i_8_390_1898_0 & ~i_8_390_2127_0))) | (~i_8_390_382_0 & ~i_8_390_587_0 & ~i_8_390_1260_0 & ~i_8_390_1543_0 & ~i_8_390_1898_0 & i_8_390_2053_0 & ~i_8_390_2130_0) | (~i_8_390_289_0 & ~i_8_390_1026_0 & ~i_8_390_1601_0 & ~i_8_390_2111_0 & ~i_8_390_2188_0 & i_8_390_2264_0))) | (i_8_390_364_0 & ((~i_8_390_193_0 & ~i_8_390_289_0 & ~i_8_390_299_0 & ~i_8_390_585_0 & ~i_8_390_820_0 & ~i_8_390_1074_0 & ~i_8_390_1260_0 & ~i_8_390_1542_0 & ~i_8_390_1601_0 & ~i_8_390_1700_0 & ~i_8_390_1735_0 & ~i_8_390_1779_0) | (~i_8_390_379_0 & ~i_8_390_1111_0 & i_8_390_1260_0 & ~i_8_390_1539_0 & ~i_8_390_2130_0 & ~i_8_390_2187_0))) | (~i_8_390_1026_0 & ((~i_8_390_366_0 & ((i_8_390_616_0 & i_8_390_1264_0 & ~i_8_390_1491_0 & i_8_390_1651_0 & ~i_8_390_1779_0 & ~i_8_390_1896_0) | (~i_8_390_380_0 & ~i_8_390_394_0 & i_8_390_697_0 & ~i_8_390_992_0 & ~i_8_390_1111_0 & ~i_8_390_1539_0 & ~i_8_390_1543_0 & ~i_8_390_1780_0 & i_8_390_2128_0 & ~i_8_390_2187_0 & ~i_8_390_2189_0))) | (~i_8_390_585_0 & ((~i_8_390_393_0 & ((i_8_390_193_0 & i_8_390_382_0 & ~i_8_390_475_0 & ~i_8_390_606_0 & ~i_8_390_1112_0 & ~i_8_390_1455_0 & ~i_8_390_1896_0 & ~i_8_390_2187_0) | (~i_8_390_395_0 & ~i_8_390_555_0 & ~i_8_390_587_0 & ~i_8_390_992_0 & i_8_390_1299_0 & ~i_8_390_1650_0 & ~i_8_390_2188_0))) | (~i_8_390_299_0 & ~i_8_390_380_0 & ~i_8_390_395_0 & ~i_8_390_465_0 & ~i_8_390_658_0 & i_8_390_697_0 & ~i_8_390_1111_0 & ~i_8_390_1159_0 & ~i_8_390_1455_0 & ~i_8_390_1491_0 & ~i_8_390_1700_0 & ~i_8_390_2187_0 & ~i_8_390_2188_0 & ~i_8_390_2291_0))) | (~i_8_390_393_0 & ~i_8_390_587_0 & ((~i_8_390_992_0 & ((~i_8_390_395_0 & i_8_390_614_0 & ~i_8_390_660_0 & ~i_8_390_1074_0 & ~i_8_390_1542_0 & ~i_8_390_2171_0 & ~i_8_390_2188_0) | (i_8_390_615_0 & ~i_8_390_1077_0 & ~i_8_390_1457_0 & ~i_8_390_1539_0 & ~i_8_390_1637_0 & ~i_8_390_1897_0 & ~i_8_390_2127_0 & ~i_8_390_2189_0))) | (i_8_390_379_0 & i_8_390_457_0 & ~i_8_390_1542_0 & ~i_8_390_2171_0))))) | (~i_8_390_1457_0 & ((~i_8_390_193_0 & ~i_8_390_820_0 & ~i_8_390_2189_0 & ((~i_8_390_53_0 & ~i_8_390_364_0 & ~i_8_390_367_0 & ~i_8_390_555_0 & ~i_8_390_613_0 & ~i_8_390_1077_0 & i_8_390_1111_0 & ~i_8_390_1159_0 & ~i_8_390_1260_0 & i_8_390_1780_0) | (~i_8_390_299_0 & ~i_8_390_379_0 & ~i_8_390_395_0 & ~i_8_390_475_0 & ~i_8_390_712_0 & ~i_8_390_1111_0 & ~i_8_390_1264_0 & ~i_8_390_1543_0 & ~i_8_390_1779_0 & ~i_8_390_1898_0 & ~i_8_390_2130_0 & ~i_8_390_2187_0 & ~i_8_390_2077_0 & ~i_8_390_2127_0))) | (~i_8_390_393_0 & ~i_8_390_1539_0 & ((~i_8_390_367_0 & ~i_8_390_587_0 & ~i_8_390_613_0 & ~i_8_390_1159_0 & ~i_8_390_1637_0 & i_8_390_1651_0 & ~i_8_390_2008_0 & ~i_8_390_2130_0) | (~i_8_390_289_0 & i_8_390_702_0 & i_8_390_1264_0 & ~i_8_390_1455_0 & ~i_8_390_1542_0 & ~i_8_390_2264_0))) | (~i_8_390_380_0 & i_8_390_1074_0 & i_8_390_1077_0 & ~i_8_390_1685_0 & ~i_8_390_1896_0 & ~i_8_390_2127_0))) | (~i_8_390_380_0 & ((~i_8_390_1539_0 & ((~i_8_390_193_0 & ((i_8_390_367_0 & ~i_8_390_465_0 & ~i_8_390_475_0 & ~i_8_390_955_0 & ~i_8_390_1491_0 & ~i_8_390_1542_0 & ~i_8_390_1601_0 & ~i_8_390_1650_0 & ~i_8_390_1700_0 & ~i_8_390_1915_0 & ~i_8_390_2008_0 & ~i_8_390_2111_0) | (~i_8_390_364_0 & ~i_8_390_379_0 & ~i_8_390_661_0 & ~i_8_390_1260_0 & ~i_8_390_1264_0 & ~i_8_390_1779_0 & i_8_390_2127_0 & i_8_390_2128_0 & ~i_8_390_2291_0))) | (~i_8_390_697_0 & ~i_8_390_1076_0 & ~i_8_390_1111_0 & i_8_390_1268_0 & ~i_8_390_1492_0 & ~i_8_390_1601_0 & ~i_8_390_1651_0))) | (i_8_390_256_0 & i_8_390_382_0 & ~i_8_390_394_0 & ~i_8_390_1735_0 & ~i_8_390_1779_0) | (~i_8_390_712_0 & i_8_390_1111_0 & ~i_8_390_1159_0 & ~i_8_390_1230_0 & ~i_8_390_1260_0 & i_8_390_1268_0 & ~i_8_390_1601_0 & ~i_8_390_1700_0 & ~i_8_390_1898_0 & ~i_8_390_2077_0 & ~i_8_390_2187_0))) | (~i_8_390_382_0 & ((~i_8_390_379_0 & ~i_8_390_585_0 & i_8_390_702_0 & ~i_8_390_820_0 & i_8_390_1026_0 & ~i_8_390_1072_0 & ~i_8_390_1896_0) | (~i_8_390_364_0 & ~i_8_390_394_0 & i_8_390_1072_0 & ~i_8_390_1159_0 & ~i_8_390_1299_0 & ~i_8_390_1539_0 & ~i_8_390_1897_0 & ~i_8_390_1904_0 & ~i_8_390_2008_0 & ~i_8_390_2127_0 & ~i_8_390_2187_0))) | (~i_8_390_1554_0 & ((~i_8_390_364_0 & ((~i_8_390_1111_0 & ~i_8_390_1112_0 & i_8_390_1652_0 & ~i_8_390_1898_0 & ~i_8_390_1904_0) | (~i_8_390_289_0 & ~i_8_390_475_0 & ~i_8_390_587_0 & ~i_8_390_820_0 & ~i_8_390_992_0 & i_8_390_1074_0 & ~i_8_390_2187_0))) | (~i_8_390_712_0 & ~i_8_390_2111_0 & ((i_8_390_457_0 & ~i_8_390_1112_0 & ~i_8_390_2130_0) | (~i_8_390_1780_0 & i_8_390_1904_0 & ~i_8_390_2291_0))) | (i_8_390_613_0 & ~i_8_390_820_0 & i_8_390_1111_0 & ~i_8_390_1735_0 & ~i_8_390_1780_0 & ~i_8_390_2188_0))) | (~i_8_390_1601_0 & ((~i_8_390_393_0 & ~i_8_390_1898_0 & ((~i_8_390_299_0 & ~i_8_390_395_0 & ~i_8_390_555_0 & ~i_8_390_813_0 & i_8_390_992_0 & ~i_8_390_1539_0 & ~i_8_390_1896_0 & ~i_8_390_2077_0 & ~i_8_390_2187_0) | (~i_8_390_394_0 & i_8_390_1111_0 & i_8_390_1112_0 & ~i_8_390_1542_0 & ~i_8_390_1637_0 & i_8_390_1651_0 & ~i_8_390_2189_0 & ~i_8_390_2264_0 & ~i_8_390_2291_0))) | (i_8_390_193_0 & ~i_8_390_660_0 & ~i_8_390_712_0 & ~i_8_390_814_0 & i_8_390_1077_0 & ~i_8_390_1260_0 & ~i_8_390_1700_0 & ~i_8_390_2291_0) | (~i_8_390_289_0 & i_8_390_815_0 & ~i_8_390_1780_0 & ~i_8_390_1897_0 & ~i_8_390_2189_0) | (~i_8_390_555_0 & i_8_390_816_0 & ~i_8_390_1779_0 & ~i_8_390_2111_0))) | (~i_8_390_394_0 & ((i_8_390_193_0 & ((~i_8_390_289_0 & i_8_390_1652_0 & ~i_8_390_1915_0 & ~i_8_390_2111_0) | (~i_8_390_658_0 & ~i_8_390_697_0 & ~i_8_390_820_0 & ~i_8_390_1543_0 & ~i_8_390_1780_0 & ~i_8_390_2130_0))) | (~i_8_390_379_0 & ~i_8_390_395_0 & i_8_390_1232_0 & ~i_8_390_1915_0 & ~i_8_390_2130_0 & ~i_8_390_2189_0 & ~i_8_390_2264_0))) | (~i_8_390_299_0 & ((~i_8_390_393_0 & i_8_390_612_0 & ~i_8_390_820_0 & i_8_390_1299_0 & ~i_8_390_1542_0 & ~i_8_390_1897_0) | (~i_8_390_395_0 & ~i_8_390_587_0 & i_8_390_1651_0 & ~i_8_390_1779_0 & ~i_8_390_2077_0 & ~i_8_390_2187_0))) | (~i_8_390_379_0 & ((~i_8_390_395_0 & i_8_390_817_0 & ~i_8_390_1491_0 & ~i_8_390_1898_0 & ~i_8_390_2130_0) | (~i_8_390_587_0 & ~i_8_390_1232_0 & ~i_8_390_1543_0 & ~i_8_390_1915_0 & ~i_8_390_2187_0 & i_8_390_2264_0))) | (~i_8_390_395_0 & ~i_8_390_1543_0 & ~i_8_390_1685_0 & ((~i_8_390_612_0 & i_8_390_1264_0 & i_8_390_1268_0) | (~i_8_390_289_0 & ~i_8_390_712_0 & i_8_390_2053_0 & i_8_390_2171_0 & ~i_8_390_2189_0))) | (~i_8_390_1700_0 & ~i_8_390_2127_0 & ((i_8_390_238_0 & i_8_390_661_0 & ~i_8_390_1264_0 & ~i_8_390_2130_0 & ~i_8_390_2187_0) | (~i_8_390_712_0 & ~i_8_390_1268_0 & i_8_390_1685_0 & ~i_8_390_1780_0 & ~i_8_390_2189_0))) | (i_8_390_259_0 & i_8_390_457_0 & ~i_8_390_1896_0 & ~i_8_390_2171_0));
endmodule



// Benchmark "kernel_8_391" written by ABC on Sun Jul 19 10:09:53 2020

module kernel_8_391 ( 
    i_8_391_18_0, i_8_391_22_0, i_8_391_26_0, i_8_391_41_0, i_8_391_67_0,
    i_8_391_115_0, i_8_391_130_0, i_8_391_139_0, i_8_391_179_0,
    i_8_391_197_0, i_8_391_204_0, i_8_391_262_0, i_8_391_266_0,
    i_8_391_273_0, i_8_391_305_0, i_8_391_355_0, i_8_391_385_0,
    i_8_391_428_0, i_8_391_429_0, i_8_391_445_0, i_8_391_457_0,
    i_8_391_458_0, i_8_391_460_0, i_8_391_464_0, i_8_391_481_0,
    i_8_391_509_0, i_8_391_535_0, i_8_391_538_0, i_8_391_583_0,
    i_8_391_599_0, i_8_391_626_0, i_8_391_657_0, i_8_391_661_0,
    i_8_391_664_0, i_8_391_682_0, i_8_391_694_0, i_8_391_710_0,
    i_8_391_715_0, i_8_391_769_0, i_8_391_790_0, i_8_391_838_0,
    i_8_391_887_0, i_8_391_896_0, i_8_391_911_0, i_8_391_1041_0,
    i_8_391_1075_0, i_8_391_1076_0, i_8_391_1115_0, i_8_391_1133_0,
    i_8_391_1175_0, i_8_391_1192_0, i_8_391_1229_0, i_8_391_1232_0,
    i_8_391_1241_0, i_8_391_1296_0, i_8_391_1315_0, i_8_391_1318_0,
    i_8_391_1354_0, i_8_391_1386_0, i_8_391_1387_0, i_8_391_1395_0,
    i_8_391_1398_0, i_8_391_1399_0, i_8_391_1403_0, i_8_391_1407_0,
    i_8_391_1434_0, i_8_391_1436_0, i_8_391_1490_0, i_8_391_1494_0,
    i_8_391_1495_0, i_8_391_1498_0, i_8_391_1529_0, i_8_391_1634_0,
    i_8_391_1656_0, i_8_391_1702_0, i_8_391_1703_0, i_8_391_1706_0,
    i_8_391_1750_0, i_8_391_1768_0, i_8_391_1773_0, i_8_391_1795_0,
    i_8_391_1796_0, i_8_391_1819_0, i_8_391_1820_0, i_8_391_1826_0,
    i_8_391_1863_0, i_8_391_1919_0, i_8_391_1976_0, i_8_391_2007_0,
    i_8_391_2062_0, i_8_391_2138_0, i_8_391_2144_0, i_8_391_2147_0,
    i_8_391_2149_0, i_8_391_2216_0, i_8_391_2232_0, i_8_391_2237_0,
    i_8_391_2245_0, i_8_391_2246_0, i_8_391_2253_0,
    o_8_391_0_0  );
  input  i_8_391_18_0, i_8_391_22_0, i_8_391_26_0, i_8_391_41_0,
    i_8_391_67_0, i_8_391_115_0, i_8_391_130_0, i_8_391_139_0,
    i_8_391_179_0, i_8_391_197_0, i_8_391_204_0, i_8_391_262_0,
    i_8_391_266_0, i_8_391_273_0, i_8_391_305_0, i_8_391_355_0,
    i_8_391_385_0, i_8_391_428_0, i_8_391_429_0, i_8_391_445_0,
    i_8_391_457_0, i_8_391_458_0, i_8_391_460_0, i_8_391_464_0,
    i_8_391_481_0, i_8_391_509_0, i_8_391_535_0, i_8_391_538_0,
    i_8_391_583_0, i_8_391_599_0, i_8_391_626_0, i_8_391_657_0,
    i_8_391_661_0, i_8_391_664_0, i_8_391_682_0, i_8_391_694_0,
    i_8_391_710_0, i_8_391_715_0, i_8_391_769_0, i_8_391_790_0,
    i_8_391_838_0, i_8_391_887_0, i_8_391_896_0, i_8_391_911_0,
    i_8_391_1041_0, i_8_391_1075_0, i_8_391_1076_0, i_8_391_1115_0,
    i_8_391_1133_0, i_8_391_1175_0, i_8_391_1192_0, i_8_391_1229_0,
    i_8_391_1232_0, i_8_391_1241_0, i_8_391_1296_0, i_8_391_1315_0,
    i_8_391_1318_0, i_8_391_1354_0, i_8_391_1386_0, i_8_391_1387_0,
    i_8_391_1395_0, i_8_391_1398_0, i_8_391_1399_0, i_8_391_1403_0,
    i_8_391_1407_0, i_8_391_1434_0, i_8_391_1436_0, i_8_391_1490_0,
    i_8_391_1494_0, i_8_391_1495_0, i_8_391_1498_0, i_8_391_1529_0,
    i_8_391_1634_0, i_8_391_1656_0, i_8_391_1702_0, i_8_391_1703_0,
    i_8_391_1706_0, i_8_391_1750_0, i_8_391_1768_0, i_8_391_1773_0,
    i_8_391_1795_0, i_8_391_1796_0, i_8_391_1819_0, i_8_391_1820_0,
    i_8_391_1826_0, i_8_391_1863_0, i_8_391_1919_0, i_8_391_1976_0,
    i_8_391_2007_0, i_8_391_2062_0, i_8_391_2138_0, i_8_391_2144_0,
    i_8_391_2147_0, i_8_391_2149_0, i_8_391_2216_0, i_8_391_2232_0,
    i_8_391_2237_0, i_8_391_2245_0, i_8_391_2246_0, i_8_391_2253_0;
  output o_8_391_0_0;
  assign o_8_391_0_0 = 0;
endmodule



// Benchmark "kernel_8_392" written by ABC on Sun Jul 19 10:09:54 2020

module kernel_8_392 ( 
    i_8_392_4_0, i_8_392_67_0, i_8_392_140_0, i_8_392_148_0, i_8_392_169_0,
    i_8_392_202_0, i_8_392_203_0, i_8_392_248_0, i_8_392_274_0,
    i_8_392_334_0, i_8_392_362_0, i_8_392_364_0, i_8_392_373_0,
    i_8_392_422_0, i_8_392_445_0, i_8_392_454_0, i_8_392_464_0,
    i_8_392_473_0, i_8_392_493_0, i_8_392_529_0, i_8_392_535_0,
    i_8_392_547_0, i_8_392_553_0, i_8_392_608_0, i_8_392_634_0,
    i_8_392_706_0, i_8_392_707_0, i_8_392_736_0, i_8_392_739_0,
    i_8_392_760_0, i_8_392_790_0, i_8_392_814_0, i_8_392_835_0,
    i_8_392_860_0, i_8_392_873_0, i_8_392_916_0, i_8_392_971_0,
    i_8_392_1067_0, i_8_392_1103_0, i_8_392_1114_0, i_8_392_1115_0,
    i_8_392_1129_0, i_8_392_1130_0, i_8_392_1201_0, i_8_392_1267_0,
    i_8_392_1301_0, i_8_392_1305_0, i_8_392_1306_0, i_8_392_1357_0,
    i_8_392_1399_0, i_8_392_1400_0, i_8_392_1407_0, i_8_392_1419_0,
    i_8_392_1435_0, i_8_392_1468_0, i_8_392_1489_0, i_8_392_1490_0,
    i_8_392_1492_0, i_8_392_1499_0, i_8_392_1546_0, i_8_392_1564_0,
    i_8_392_1573_0, i_8_392_1580_0, i_8_392_1595_0, i_8_392_1606_0,
    i_8_392_1633_0, i_8_392_1634_0, i_8_392_1705_0, i_8_392_1706_0,
    i_8_392_1729_0, i_8_392_1733_0, i_8_392_1774_0, i_8_392_1778_0,
    i_8_392_1782_0, i_8_392_1805_0, i_8_392_1810_0, i_8_392_1822_0,
    i_8_392_1823_0, i_8_392_1825_0, i_8_392_1826_0, i_8_392_1885_0,
    i_8_392_1886_0, i_8_392_1888_0, i_8_392_1904_0, i_8_392_1939_0,
    i_8_392_1981_0, i_8_392_1982_0, i_8_392_1985_0, i_8_392_2135_0,
    i_8_392_2145_0, i_8_392_2147_0, i_8_392_2150_0, i_8_392_2233_0,
    i_8_392_2249_0, i_8_392_2254_0, i_8_392_2258_0, i_8_392_2263_0,
    i_8_392_2266_0, i_8_392_2293_0, i_8_392_2299_0,
    o_8_392_0_0  );
  input  i_8_392_4_0, i_8_392_67_0, i_8_392_140_0, i_8_392_148_0,
    i_8_392_169_0, i_8_392_202_0, i_8_392_203_0, i_8_392_248_0,
    i_8_392_274_0, i_8_392_334_0, i_8_392_362_0, i_8_392_364_0,
    i_8_392_373_0, i_8_392_422_0, i_8_392_445_0, i_8_392_454_0,
    i_8_392_464_0, i_8_392_473_0, i_8_392_493_0, i_8_392_529_0,
    i_8_392_535_0, i_8_392_547_0, i_8_392_553_0, i_8_392_608_0,
    i_8_392_634_0, i_8_392_706_0, i_8_392_707_0, i_8_392_736_0,
    i_8_392_739_0, i_8_392_760_0, i_8_392_790_0, i_8_392_814_0,
    i_8_392_835_0, i_8_392_860_0, i_8_392_873_0, i_8_392_916_0,
    i_8_392_971_0, i_8_392_1067_0, i_8_392_1103_0, i_8_392_1114_0,
    i_8_392_1115_0, i_8_392_1129_0, i_8_392_1130_0, i_8_392_1201_0,
    i_8_392_1267_0, i_8_392_1301_0, i_8_392_1305_0, i_8_392_1306_0,
    i_8_392_1357_0, i_8_392_1399_0, i_8_392_1400_0, i_8_392_1407_0,
    i_8_392_1419_0, i_8_392_1435_0, i_8_392_1468_0, i_8_392_1489_0,
    i_8_392_1490_0, i_8_392_1492_0, i_8_392_1499_0, i_8_392_1546_0,
    i_8_392_1564_0, i_8_392_1573_0, i_8_392_1580_0, i_8_392_1595_0,
    i_8_392_1606_0, i_8_392_1633_0, i_8_392_1634_0, i_8_392_1705_0,
    i_8_392_1706_0, i_8_392_1729_0, i_8_392_1733_0, i_8_392_1774_0,
    i_8_392_1778_0, i_8_392_1782_0, i_8_392_1805_0, i_8_392_1810_0,
    i_8_392_1822_0, i_8_392_1823_0, i_8_392_1825_0, i_8_392_1826_0,
    i_8_392_1885_0, i_8_392_1886_0, i_8_392_1888_0, i_8_392_1904_0,
    i_8_392_1939_0, i_8_392_1981_0, i_8_392_1982_0, i_8_392_1985_0,
    i_8_392_2135_0, i_8_392_2145_0, i_8_392_2147_0, i_8_392_2150_0,
    i_8_392_2233_0, i_8_392_2249_0, i_8_392_2254_0, i_8_392_2258_0,
    i_8_392_2263_0, i_8_392_2266_0, i_8_392_2293_0, i_8_392_2299_0;
  output o_8_392_0_0;
  assign o_8_392_0_0 = 0;
endmodule



// Benchmark "kernel_8_393" written by ABC on Sun Jul 19 10:09:55 2020

module kernel_8_393 ( 
    i_8_393_4_0, i_8_393_9_0, i_8_393_24_0, i_8_393_40_0, i_8_393_43_0,
    i_8_393_53_0, i_8_393_70_0, i_8_393_85_0, i_8_393_94_0, i_8_393_104_0,
    i_8_393_141_0, i_8_393_157_0, i_8_393_159_0, i_8_393_160_0,
    i_8_393_192_0, i_8_393_241_0, i_8_393_265_0, i_8_393_293_0,
    i_8_393_346_0, i_8_393_355_0, i_8_393_371_0, i_8_393_391_0,
    i_8_393_394_0, i_8_393_417_0, i_8_393_418_0, i_8_393_420_0,
    i_8_393_421_0, i_8_393_427_0, i_8_393_428_0, i_8_393_433_0,
    i_8_393_481_0, i_8_393_483_0, i_8_393_493_0, i_8_393_535_0,
    i_8_393_553_0, i_8_393_557_0, i_8_393_605_0, i_8_393_608_0,
    i_8_393_627_0, i_8_393_628_0, i_8_393_633_0, i_8_393_662_0,
    i_8_393_672_0, i_8_393_704_0, i_8_393_709_0, i_8_393_769_0,
    i_8_393_825_0, i_8_393_849_0, i_8_393_850_0, i_8_393_922_0,
    i_8_393_938_0, i_8_393_943_0, i_8_393_951_0, i_8_393_968_0,
    i_8_393_976_0, i_8_393_991_0, i_8_393_1030_0, i_8_393_1113_0,
    i_8_393_1158_0, i_8_393_1201_0, i_8_393_1203_0, i_8_393_1258_0,
    i_8_393_1305_0, i_8_393_1307_0, i_8_393_1471_0, i_8_393_1489_0,
    i_8_393_1490_0, i_8_393_1534_0, i_8_393_1639_0, i_8_393_1654_0,
    i_8_393_1659_0, i_8_393_1671_0, i_8_393_1700_0, i_8_393_1702_0,
    i_8_393_1703_0, i_8_393_1704_0, i_8_393_1708_0, i_8_393_1729_0,
    i_8_393_1750_0, i_8_393_1781_0, i_8_393_1808_0, i_8_393_1819_0,
    i_8_393_1822_0, i_8_393_1824_0, i_8_393_1826_0, i_8_393_1974_0,
    i_8_393_1997_0, i_8_393_2001_0, i_8_393_2029_0, i_8_393_2047_0,
    i_8_393_2092_0, i_8_393_2146_0, i_8_393_2170_0, i_8_393_2182_0,
    i_8_393_2183_0, i_8_393_2214_0, i_8_393_2215_0, i_8_393_2247_0,
    i_8_393_2258_0, i_8_393_2281_0,
    o_8_393_0_0  );
  input  i_8_393_4_0, i_8_393_9_0, i_8_393_24_0, i_8_393_40_0,
    i_8_393_43_0, i_8_393_53_0, i_8_393_70_0, i_8_393_85_0, i_8_393_94_0,
    i_8_393_104_0, i_8_393_141_0, i_8_393_157_0, i_8_393_159_0,
    i_8_393_160_0, i_8_393_192_0, i_8_393_241_0, i_8_393_265_0,
    i_8_393_293_0, i_8_393_346_0, i_8_393_355_0, i_8_393_371_0,
    i_8_393_391_0, i_8_393_394_0, i_8_393_417_0, i_8_393_418_0,
    i_8_393_420_0, i_8_393_421_0, i_8_393_427_0, i_8_393_428_0,
    i_8_393_433_0, i_8_393_481_0, i_8_393_483_0, i_8_393_493_0,
    i_8_393_535_0, i_8_393_553_0, i_8_393_557_0, i_8_393_605_0,
    i_8_393_608_0, i_8_393_627_0, i_8_393_628_0, i_8_393_633_0,
    i_8_393_662_0, i_8_393_672_0, i_8_393_704_0, i_8_393_709_0,
    i_8_393_769_0, i_8_393_825_0, i_8_393_849_0, i_8_393_850_0,
    i_8_393_922_0, i_8_393_938_0, i_8_393_943_0, i_8_393_951_0,
    i_8_393_968_0, i_8_393_976_0, i_8_393_991_0, i_8_393_1030_0,
    i_8_393_1113_0, i_8_393_1158_0, i_8_393_1201_0, i_8_393_1203_0,
    i_8_393_1258_0, i_8_393_1305_0, i_8_393_1307_0, i_8_393_1471_0,
    i_8_393_1489_0, i_8_393_1490_0, i_8_393_1534_0, i_8_393_1639_0,
    i_8_393_1654_0, i_8_393_1659_0, i_8_393_1671_0, i_8_393_1700_0,
    i_8_393_1702_0, i_8_393_1703_0, i_8_393_1704_0, i_8_393_1708_0,
    i_8_393_1729_0, i_8_393_1750_0, i_8_393_1781_0, i_8_393_1808_0,
    i_8_393_1819_0, i_8_393_1822_0, i_8_393_1824_0, i_8_393_1826_0,
    i_8_393_1974_0, i_8_393_1997_0, i_8_393_2001_0, i_8_393_2029_0,
    i_8_393_2047_0, i_8_393_2092_0, i_8_393_2146_0, i_8_393_2170_0,
    i_8_393_2182_0, i_8_393_2183_0, i_8_393_2214_0, i_8_393_2215_0,
    i_8_393_2247_0, i_8_393_2258_0, i_8_393_2281_0;
  output o_8_393_0_0;
  assign o_8_393_0_0 = 0;
endmodule



// Benchmark "kernel_8_394" written by ABC on Sun Jul 19 10:09:56 2020

module kernel_8_394 ( 
    i_8_394_15_0, i_8_394_23_0, i_8_394_43_0, i_8_394_66_0, i_8_394_79_0,
    i_8_394_98_0, i_8_394_118_0, i_8_394_169_0, i_8_394_191_0,
    i_8_394_257_0, i_8_394_265_0, i_8_394_266_0, i_8_394_268_0,
    i_8_394_282_0, i_8_394_283_0, i_8_394_287_0, i_8_394_296_0,
    i_8_394_299_0, i_8_394_338_0, i_8_394_340_0, i_8_394_382_0,
    i_8_394_430_0, i_8_394_454_0, i_8_394_456_0, i_8_394_491_0,
    i_8_394_492_0, i_8_394_493_0, i_8_394_502_0, i_8_394_529_0,
    i_8_394_530_0, i_8_394_583_0, i_8_394_588_0, i_8_394_592_0,
    i_8_394_615_0, i_8_394_628_0, i_8_394_672_0, i_8_394_673_0,
    i_8_394_690_0, i_8_394_693_0, i_8_394_711_0, i_8_394_716_0,
    i_8_394_718_0, i_8_394_719_0, i_8_394_750_0, i_8_394_769_0,
    i_8_394_770_0, i_8_394_772_0, i_8_394_789_0, i_8_394_795_0,
    i_8_394_822_0, i_8_394_842_0, i_8_394_843_0, i_8_394_845_0,
    i_8_394_880_0, i_8_394_894_0, i_8_394_954_0, i_8_394_1012_0,
    i_8_394_1021_0, i_8_394_1024_0, i_8_394_1033_0, i_8_394_1074_0,
    i_8_394_1078_0, i_8_394_1079_0, i_8_394_1087_0, i_8_394_1220_0,
    i_8_394_1242_0, i_8_394_1249_0, i_8_394_1254_0, i_8_394_1257_0,
    i_8_394_1258_0, i_8_394_1259_0, i_8_394_1267_0, i_8_394_1270_0,
    i_8_394_1295_0, i_8_394_1297_0, i_8_394_1310_0, i_8_394_1353_0,
    i_8_394_1417_0, i_8_394_1434_0, i_8_394_1457_0, i_8_394_1464_0,
    i_8_394_1617_0, i_8_394_1639_0, i_8_394_1650_0, i_8_394_1696_0,
    i_8_394_1704_0, i_8_394_1706_0, i_8_394_1728_0, i_8_394_1763_0,
    i_8_394_1927_0, i_8_394_1929_0, i_8_394_1936_0, i_8_394_2022_0,
    i_8_394_2023_0, i_8_394_2194_0, i_8_394_2195_0, i_8_394_2212_0,
    i_8_394_2262_0, i_8_394_2266_0, i_8_394_2281_0,
    o_8_394_0_0  );
  input  i_8_394_15_0, i_8_394_23_0, i_8_394_43_0, i_8_394_66_0,
    i_8_394_79_0, i_8_394_98_0, i_8_394_118_0, i_8_394_169_0,
    i_8_394_191_0, i_8_394_257_0, i_8_394_265_0, i_8_394_266_0,
    i_8_394_268_0, i_8_394_282_0, i_8_394_283_0, i_8_394_287_0,
    i_8_394_296_0, i_8_394_299_0, i_8_394_338_0, i_8_394_340_0,
    i_8_394_382_0, i_8_394_430_0, i_8_394_454_0, i_8_394_456_0,
    i_8_394_491_0, i_8_394_492_0, i_8_394_493_0, i_8_394_502_0,
    i_8_394_529_0, i_8_394_530_0, i_8_394_583_0, i_8_394_588_0,
    i_8_394_592_0, i_8_394_615_0, i_8_394_628_0, i_8_394_672_0,
    i_8_394_673_0, i_8_394_690_0, i_8_394_693_0, i_8_394_711_0,
    i_8_394_716_0, i_8_394_718_0, i_8_394_719_0, i_8_394_750_0,
    i_8_394_769_0, i_8_394_770_0, i_8_394_772_0, i_8_394_789_0,
    i_8_394_795_0, i_8_394_822_0, i_8_394_842_0, i_8_394_843_0,
    i_8_394_845_0, i_8_394_880_0, i_8_394_894_0, i_8_394_954_0,
    i_8_394_1012_0, i_8_394_1021_0, i_8_394_1024_0, i_8_394_1033_0,
    i_8_394_1074_0, i_8_394_1078_0, i_8_394_1079_0, i_8_394_1087_0,
    i_8_394_1220_0, i_8_394_1242_0, i_8_394_1249_0, i_8_394_1254_0,
    i_8_394_1257_0, i_8_394_1258_0, i_8_394_1259_0, i_8_394_1267_0,
    i_8_394_1270_0, i_8_394_1295_0, i_8_394_1297_0, i_8_394_1310_0,
    i_8_394_1353_0, i_8_394_1417_0, i_8_394_1434_0, i_8_394_1457_0,
    i_8_394_1464_0, i_8_394_1617_0, i_8_394_1639_0, i_8_394_1650_0,
    i_8_394_1696_0, i_8_394_1704_0, i_8_394_1706_0, i_8_394_1728_0,
    i_8_394_1763_0, i_8_394_1927_0, i_8_394_1929_0, i_8_394_1936_0,
    i_8_394_2022_0, i_8_394_2023_0, i_8_394_2194_0, i_8_394_2195_0,
    i_8_394_2212_0, i_8_394_2262_0, i_8_394_2266_0, i_8_394_2281_0;
  output o_8_394_0_0;
  assign o_8_394_0_0 = 0;
endmodule



// Benchmark "kernel_8_395" written by ABC on Sun Jul 19 10:09:57 2020

module kernel_8_395 ( 
    i_8_395_5_0, i_8_395_69_0, i_8_395_78_0, i_8_395_79_0, i_8_395_88_0,
    i_8_395_114_0, i_8_395_159_0, i_8_395_204_0, i_8_395_205_0,
    i_8_395_206_0, i_8_395_249_0, i_8_395_251_0, i_8_395_277_0,
    i_8_395_278_0, i_8_395_286_0, i_8_395_305_0, i_8_395_332_0,
    i_8_395_348_0, i_8_395_349_0, i_8_395_350_0, i_8_395_355_0,
    i_8_395_358_0, i_8_395_363_0, i_8_395_393_0, i_8_395_404_0,
    i_8_395_422_0, i_8_395_445_0, i_8_395_446_0, i_8_395_519_0,
    i_8_395_528_0, i_8_395_555_0, i_8_395_592_0, i_8_395_601_0,
    i_8_395_602_0, i_8_395_615_0, i_8_395_618_0, i_8_395_619_0,
    i_8_395_696_0, i_8_395_706_0, i_8_395_726_0, i_8_395_762_0,
    i_8_395_818_0, i_8_395_836_0, i_8_395_840_0, i_8_395_845_0,
    i_8_395_849_0, i_8_395_868_0, i_8_395_880_0, i_8_395_918_0,
    i_8_395_951_0, i_8_395_961_0, i_8_395_1015_0, i_8_395_1060_0,
    i_8_395_1075_0, i_8_395_1086_0, i_8_395_1087_0, i_8_395_1088_0,
    i_8_395_1115_0, i_8_395_1178_0, i_8_395_1203_0, i_8_395_1258_0,
    i_8_395_1284_0, i_8_395_1286_0, i_8_395_1328_0, i_8_395_1410_0,
    i_8_395_1438_0, i_8_395_1456_0, i_8_395_1457_0, i_8_395_1502_0,
    i_8_395_1543_0, i_8_395_1591_0, i_8_395_1592_0, i_8_395_1617_0,
    i_8_395_1661_0, i_8_395_1749_0, i_8_395_1752_0, i_8_395_1753_0,
    i_8_395_1772_0, i_8_395_1797_0, i_8_395_1799_0, i_8_395_1808_0,
    i_8_395_1815_0, i_8_395_1816_0, i_8_395_1835_0, i_8_395_1853_0,
    i_8_395_1896_0, i_8_395_1897_0, i_8_395_1941_0, i_8_395_1969_0,
    i_8_395_1978_0, i_8_395_2004_0, i_8_395_2013_0, i_8_395_2014_0,
    i_8_395_2058_0, i_8_395_2059_0, i_8_395_2069_0, i_8_395_2152_0,
    i_8_395_2193_0, i_8_395_2194_0, i_8_395_2218_0,
    o_8_395_0_0  );
  input  i_8_395_5_0, i_8_395_69_0, i_8_395_78_0, i_8_395_79_0,
    i_8_395_88_0, i_8_395_114_0, i_8_395_159_0, i_8_395_204_0,
    i_8_395_205_0, i_8_395_206_0, i_8_395_249_0, i_8_395_251_0,
    i_8_395_277_0, i_8_395_278_0, i_8_395_286_0, i_8_395_305_0,
    i_8_395_332_0, i_8_395_348_0, i_8_395_349_0, i_8_395_350_0,
    i_8_395_355_0, i_8_395_358_0, i_8_395_363_0, i_8_395_393_0,
    i_8_395_404_0, i_8_395_422_0, i_8_395_445_0, i_8_395_446_0,
    i_8_395_519_0, i_8_395_528_0, i_8_395_555_0, i_8_395_592_0,
    i_8_395_601_0, i_8_395_602_0, i_8_395_615_0, i_8_395_618_0,
    i_8_395_619_0, i_8_395_696_0, i_8_395_706_0, i_8_395_726_0,
    i_8_395_762_0, i_8_395_818_0, i_8_395_836_0, i_8_395_840_0,
    i_8_395_845_0, i_8_395_849_0, i_8_395_868_0, i_8_395_880_0,
    i_8_395_918_0, i_8_395_951_0, i_8_395_961_0, i_8_395_1015_0,
    i_8_395_1060_0, i_8_395_1075_0, i_8_395_1086_0, i_8_395_1087_0,
    i_8_395_1088_0, i_8_395_1115_0, i_8_395_1178_0, i_8_395_1203_0,
    i_8_395_1258_0, i_8_395_1284_0, i_8_395_1286_0, i_8_395_1328_0,
    i_8_395_1410_0, i_8_395_1438_0, i_8_395_1456_0, i_8_395_1457_0,
    i_8_395_1502_0, i_8_395_1543_0, i_8_395_1591_0, i_8_395_1592_0,
    i_8_395_1617_0, i_8_395_1661_0, i_8_395_1749_0, i_8_395_1752_0,
    i_8_395_1753_0, i_8_395_1772_0, i_8_395_1797_0, i_8_395_1799_0,
    i_8_395_1808_0, i_8_395_1815_0, i_8_395_1816_0, i_8_395_1835_0,
    i_8_395_1853_0, i_8_395_1896_0, i_8_395_1897_0, i_8_395_1941_0,
    i_8_395_1969_0, i_8_395_1978_0, i_8_395_2004_0, i_8_395_2013_0,
    i_8_395_2014_0, i_8_395_2058_0, i_8_395_2059_0, i_8_395_2069_0,
    i_8_395_2152_0, i_8_395_2193_0, i_8_395_2194_0, i_8_395_2218_0;
  output o_8_395_0_0;
  assign o_8_395_0_0 = ~((~i_8_395_1088_0 & ((~i_8_395_88_0 & ((~i_8_395_278_0 & ~i_8_395_555_0 & ~i_8_395_1502_0 & ~i_8_395_1797_0 & ~i_8_395_1816_0) | (~i_8_395_5_0 & ~i_8_395_249_0 & ~i_8_395_762_0 & ~i_8_395_1086_0 & ~i_8_395_1617_0 & ~i_8_395_1853_0 & ~i_8_395_2069_0 & ~i_8_395_2152_0))) | (~i_8_395_355_0 & ~i_8_395_696_0 & ~i_8_395_1075_0 & i_8_395_1438_0 & ~i_8_395_1896_0 & ~i_8_395_2013_0 & ~i_8_395_2059_0 & ~i_8_395_2069_0) | (i_8_395_88_0 & ~i_8_395_251_0 & ~i_8_395_445_0 & ~i_8_395_726_0 & ~i_8_395_918_0 & ~i_8_395_1815_0 & ~i_8_395_1816_0 & ~i_8_395_1941_0 & ~i_8_395_2004_0 & ~i_8_395_2152_0 & ~i_8_395_2194_0) | (~i_8_395_358_0 & ~i_8_395_615_0 & ~i_8_395_762_0 & ~i_8_395_1087_0 & ~i_8_395_1203_0 & ~i_8_395_1799_0 & ~i_8_395_2014_0 & ~i_8_395_2218_0))) | (~i_8_395_205_0 & ((~i_8_395_204_0 & ~i_8_395_1086_0 & ((~i_8_395_278_0 & ~i_8_395_618_0 & ~i_8_395_1178_0 & ~i_8_395_1502_0 & ~i_8_395_1799_0) | (~i_8_395_206_0 & ~i_8_395_393_0 & ~i_8_395_528_0 & ~i_8_395_961_0 & ~i_8_395_1853_0))) | (i_8_395_277_0 & ~i_8_395_1075_0 & ~i_8_395_1438_0 & ~i_8_395_1808_0 & ~i_8_395_1815_0 & ~i_8_395_1853_0))) | (~i_8_395_726_0 & ((~i_8_395_206_0 & ((~i_8_395_277_0 & ~i_8_395_358_0 & ~i_8_395_519_0 & ~i_8_395_1087_0 & ~i_8_395_1115_0 & ~i_8_395_1797_0) | (~i_8_395_602_0 & ~i_8_395_849_0 & ~i_8_395_1086_0 & ~i_8_395_1749_0 & ~i_8_395_1816_0 & ~i_8_395_2152_0 & ~i_8_395_2218_0))) | (~i_8_395_519_0 & ~i_8_395_528_0 & i_8_395_592_0 & ~i_8_395_762_0 & ~i_8_395_1115_0))) | (~i_8_395_355_0 & ((~i_8_395_249_0 & ((i_8_395_350_0 & ~i_8_395_836_0 & ~i_8_395_1328_0 & ~i_8_395_1456_0 & ~i_8_395_2013_0) | (~i_8_395_445_0 & ~i_8_395_615_0 & ~i_8_395_1410_0 & ~i_8_395_1502_0 & ~i_8_395_1799_0 & ~i_8_395_2014_0))) | (~i_8_395_159_0 & ~i_8_395_358_0 & ~i_8_395_422_0 & ~i_8_395_519_0 & ~i_8_395_762_0 & i_8_395_1438_0 & ~i_8_395_1502_0 & ~i_8_395_1543_0 & ~i_8_395_1661_0 & ~i_8_395_2013_0))) | (~i_8_395_818_0 & ((~i_8_395_78_0 & i_8_395_1286_0 & ~i_8_395_1799_0 & ~i_8_395_1816_0) | (~i_8_395_445_0 & ~i_8_395_706_0 & i_8_395_1015_0 & ~i_8_395_1087_0 & i_8_395_1456_0 & ~i_8_395_1853_0))) | (i_8_395_592_0 & i_8_395_845_0 & i_8_395_1543_0) | (~i_8_395_278_0 & ~i_8_395_446_0 & i_8_395_555_0 & ~i_8_395_1502_0 & ~i_8_395_1797_0 & ~i_8_395_1815_0 & ~i_8_395_1816_0));
endmodule



// Benchmark "kernel_8_396" written by ABC on Sun Jul 19 10:09:58 2020

module kernel_8_396 ( 
    i_8_396_43_0, i_8_396_55_0, i_8_396_61_0, i_8_396_96_0, i_8_396_106_0,
    i_8_396_121_0, i_8_396_142_0, i_8_396_249_0, i_8_396_255_0,
    i_8_396_295_0, i_8_396_300_0, i_8_396_301_0, i_8_396_321_0,
    i_8_396_328_0, i_8_396_330_0, i_8_396_340_0, i_8_396_367_0,
    i_8_396_429_0, i_8_396_436_0, i_8_396_439_0, i_8_396_440_0,
    i_8_396_457_0, i_8_396_460_0, i_8_396_484_0, i_8_396_486_0,
    i_8_396_489_0, i_8_396_492_0, i_8_396_588_0, i_8_396_593_0,
    i_8_396_618_0, i_8_396_624_0, i_8_396_627_0, i_8_396_635_0,
    i_8_396_661_0, i_8_396_664_0, i_8_396_672_0, i_8_396_708_0,
    i_8_396_717_0, i_8_396_736_0, i_8_396_768_0, i_8_396_807_0,
    i_8_396_808_0, i_8_396_835_0, i_8_396_840_0, i_8_396_845_0,
    i_8_396_873_0, i_8_396_970_0, i_8_396_979_0, i_8_396_993_0,
    i_8_396_1104_0, i_8_396_1105_0, i_8_396_1115_0, i_8_396_1152_0,
    i_8_396_1183_0, i_8_396_1228_0, i_8_396_1239_0, i_8_396_1258_0,
    i_8_396_1270_0, i_8_396_1354_0, i_8_396_1357_0, i_8_396_1393_0,
    i_8_396_1401_0, i_8_396_1428_0, i_8_396_1440_0, i_8_396_1447_0,
    i_8_396_1545_0, i_8_396_1588_0, i_8_396_1591_0, i_8_396_1681_0,
    i_8_396_1701_0, i_8_396_1705_0, i_8_396_1752_0, i_8_396_1754_0,
    i_8_396_1767_0, i_8_396_1768_0, i_8_396_1770_0, i_8_396_1777_0,
    i_8_396_1788_0, i_8_396_1789_0, i_8_396_1824_0, i_8_396_1825_0,
    i_8_396_1854_0, i_8_396_1857_0, i_8_396_1858_0, i_8_396_1861_0,
    i_8_396_1907_0, i_8_396_1942_0, i_8_396_1990_0, i_8_396_1995_0,
    i_8_396_2028_0, i_8_396_2031_0, i_8_396_2058_0, i_8_396_2091_0,
    i_8_396_2100_0, i_8_396_2109_0, i_8_396_2131_0, i_8_396_2133_0,
    i_8_396_2193_0, i_8_396_2194_0, i_8_396_2278_0,
    o_8_396_0_0  );
  input  i_8_396_43_0, i_8_396_55_0, i_8_396_61_0, i_8_396_96_0,
    i_8_396_106_0, i_8_396_121_0, i_8_396_142_0, i_8_396_249_0,
    i_8_396_255_0, i_8_396_295_0, i_8_396_300_0, i_8_396_301_0,
    i_8_396_321_0, i_8_396_328_0, i_8_396_330_0, i_8_396_340_0,
    i_8_396_367_0, i_8_396_429_0, i_8_396_436_0, i_8_396_439_0,
    i_8_396_440_0, i_8_396_457_0, i_8_396_460_0, i_8_396_484_0,
    i_8_396_486_0, i_8_396_489_0, i_8_396_492_0, i_8_396_588_0,
    i_8_396_593_0, i_8_396_618_0, i_8_396_624_0, i_8_396_627_0,
    i_8_396_635_0, i_8_396_661_0, i_8_396_664_0, i_8_396_672_0,
    i_8_396_708_0, i_8_396_717_0, i_8_396_736_0, i_8_396_768_0,
    i_8_396_807_0, i_8_396_808_0, i_8_396_835_0, i_8_396_840_0,
    i_8_396_845_0, i_8_396_873_0, i_8_396_970_0, i_8_396_979_0,
    i_8_396_993_0, i_8_396_1104_0, i_8_396_1105_0, i_8_396_1115_0,
    i_8_396_1152_0, i_8_396_1183_0, i_8_396_1228_0, i_8_396_1239_0,
    i_8_396_1258_0, i_8_396_1270_0, i_8_396_1354_0, i_8_396_1357_0,
    i_8_396_1393_0, i_8_396_1401_0, i_8_396_1428_0, i_8_396_1440_0,
    i_8_396_1447_0, i_8_396_1545_0, i_8_396_1588_0, i_8_396_1591_0,
    i_8_396_1681_0, i_8_396_1701_0, i_8_396_1705_0, i_8_396_1752_0,
    i_8_396_1754_0, i_8_396_1767_0, i_8_396_1768_0, i_8_396_1770_0,
    i_8_396_1777_0, i_8_396_1788_0, i_8_396_1789_0, i_8_396_1824_0,
    i_8_396_1825_0, i_8_396_1854_0, i_8_396_1857_0, i_8_396_1858_0,
    i_8_396_1861_0, i_8_396_1907_0, i_8_396_1942_0, i_8_396_1990_0,
    i_8_396_1995_0, i_8_396_2028_0, i_8_396_2031_0, i_8_396_2058_0,
    i_8_396_2091_0, i_8_396_2100_0, i_8_396_2109_0, i_8_396_2131_0,
    i_8_396_2133_0, i_8_396_2193_0, i_8_396_2194_0, i_8_396_2278_0;
  output o_8_396_0_0;
  assign o_8_396_0_0 = 0;
endmodule



// Benchmark "kernel_8_397" written by ABC on Sun Jul 19 10:10:00 2020

module kernel_8_397 ( 
    i_8_397_22_0, i_8_397_79_0, i_8_397_142_0, i_8_397_196_0,
    i_8_397_229_0, i_8_397_232_0, i_8_397_266_0, i_8_397_309_0,
    i_8_397_312_0, i_8_397_348_0, i_8_397_366_0, i_8_397_385_0,
    i_8_397_401_0, i_8_397_489_0, i_8_397_571_0, i_8_397_572_0,
    i_8_397_582_0, i_8_397_589_0, i_8_397_606_0, i_8_397_625_0,
    i_8_397_654_0, i_8_397_655_0, i_8_397_679_0, i_8_397_696_0,
    i_8_397_697_0, i_8_397_698_0, i_8_397_699_0, i_8_397_700_0,
    i_8_397_701_0, i_8_397_705_0, i_8_397_708_0, i_8_397_733_0,
    i_8_397_751_0, i_8_397_835_0, i_8_397_840_0, i_8_397_843_0,
    i_8_397_864_0, i_8_397_880_0, i_8_397_886_0, i_8_397_966_0,
    i_8_397_968_0, i_8_397_1041_0, i_8_397_1049_0, i_8_397_1093_0,
    i_8_397_1132_0, i_8_397_1147_0, i_8_397_1148_0, i_8_397_1168_0,
    i_8_397_1227_0, i_8_397_1230_0, i_8_397_1231_0, i_8_397_1267_0,
    i_8_397_1305_0, i_8_397_1317_0, i_8_397_1318_0, i_8_397_1357_0,
    i_8_397_1358_0, i_8_397_1373_0, i_8_397_1375_0, i_8_397_1390_0,
    i_8_397_1405_0, i_8_397_1449_0, i_8_397_1491_0, i_8_397_1492_0,
    i_8_397_1525_0, i_8_397_1543_0, i_8_397_1552_0, i_8_397_1599_0,
    i_8_397_1600_0, i_8_397_1624_0, i_8_397_1641_0, i_8_397_1642_0,
    i_8_397_1654_0, i_8_397_1655_0, i_8_397_1663_0, i_8_397_1751_0,
    i_8_397_1779_0, i_8_397_1780_0, i_8_397_1824_0, i_8_397_1825_0,
    i_8_397_1857_0, i_8_397_1860_0, i_8_397_1874_0, i_8_397_1904_0,
    i_8_397_1929_0, i_8_397_1939_0, i_8_397_1982_0, i_8_397_1992_0,
    i_8_397_2075_0, i_8_397_2086_0, i_8_397_2092_0, i_8_397_2093_0,
    i_8_397_2149_0, i_8_397_2152_0, i_8_397_2167_0, i_8_397_2174_0,
    i_8_397_2233_0, i_8_397_2244_0, i_8_397_2257_0, i_8_397_2273_0,
    o_8_397_0_0  );
  input  i_8_397_22_0, i_8_397_79_0, i_8_397_142_0, i_8_397_196_0,
    i_8_397_229_0, i_8_397_232_0, i_8_397_266_0, i_8_397_309_0,
    i_8_397_312_0, i_8_397_348_0, i_8_397_366_0, i_8_397_385_0,
    i_8_397_401_0, i_8_397_489_0, i_8_397_571_0, i_8_397_572_0,
    i_8_397_582_0, i_8_397_589_0, i_8_397_606_0, i_8_397_625_0,
    i_8_397_654_0, i_8_397_655_0, i_8_397_679_0, i_8_397_696_0,
    i_8_397_697_0, i_8_397_698_0, i_8_397_699_0, i_8_397_700_0,
    i_8_397_701_0, i_8_397_705_0, i_8_397_708_0, i_8_397_733_0,
    i_8_397_751_0, i_8_397_835_0, i_8_397_840_0, i_8_397_843_0,
    i_8_397_864_0, i_8_397_880_0, i_8_397_886_0, i_8_397_966_0,
    i_8_397_968_0, i_8_397_1041_0, i_8_397_1049_0, i_8_397_1093_0,
    i_8_397_1132_0, i_8_397_1147_0, i_8_397_1148_0, i_8_397_1168_0,
    i_8_397_1227_0, i_8_397_1230_0, i_8_397_1231_0, i_8_397_1267_0,
    i_8_397_1305_0, i_8_397_1317_0, i_8_397_1318_0, i_8_397_1357_0,
    i_8_397_1358_0, i_8_397_1373_0, i_8_397_1375_0, i_8_397_1390_0,
    i_8_397_1405_0, i_8_397_1449_0, i_8_397_1491_0, i_8_397_1492_0,
    i_8_397_1525_0, i_8_397_1543_0, i_8_397_1552_0, i_8_397_1599_0,
    i_8_397_1600_0, i_8_397_1624_0, i_8_397_1641_0, i_8_397_1642_0,
    i_8_397_1654_0, i_8_397_1655_0, i_8_397_1663_0, i_8_397_1751_0,
    i_8_397_1779_0, i_8_397_1780_0, i_8_397_1824_0, i_8_397_1825_0,
    i_8_397_1857_0, i_8_397_1860_0, i_8_397_1874_0, i_8_397_1904_0,
    i_8_397_1929_0, i_8_397_1939_0, i_8_397_1982_0, i_8_397_1992_0,
    i_8_397_2075_0, i_8_397_2086_0, i_8_397_2092_0, i_8_397_2093_0,
    i_8_397_2149_0, i_8_397_2152_0, i_8_397_2167_0, i_8_397_2174_0,
    i_8_397_2233_0, i_8_397_2244_0, i_8_397_2257_0, i_8_397_2273_0;
  output o_8_397_0_0;
  assign o_8_397_0_0 = 0;
endmodule



// Benchmark "kernel_8_398" written by ABC on Sun Jul 19 10:10:00 2020

module kernel_8_398 ( 
    i_8_398_19_0, i_8_398_109_0, i_8_398_139_0, i_8_398_238_0,
    i_8_398_300_0, i_8_398_310_0, i_8_398_372_0, i_8_398_373_0,
    i_8_398_375_0, i_8_398_381_0, i_8_398_383_0, i_8_398_419_0,
    i_8_398_431_0, i_8_398_460_0, i_8_398_463_0, i_8_398_479_0,
    i_8_398_480_0, i_8_398_506_0, i_8_398_510_0, i_8_398_529_0,
    i_8_398_549_0, i_8_398_552_0, i_8_398_553_0, i_8_398_590_0,
    i_8_398_603_0, i_8_398_606_0, i_8_398_613_0, i_8_398_706_0,
    i_8_398_796_0, i_8_398_858_0, i_8_398_867_0, i_8_398_868_0,
    i_8_398_878_0, i_8_398_976_0, i_8_398_991_0, i_8_398_1030_0,
    i_8_398_1084_0, i_8_398_1127_0, i_8_398_1130_0, i_8_398_1158_0,
    i_8_398_1188_0, i_8_398_1189_0, i_8_398_1192_0, i_8_398_1255_0,
    i_8_398_1279_0, i_8_398_1283_0, i_8_398_1325_0, i_8_398_1326_0,
    i_8_398_1327_0, i_8_398_1480_0, i_8_398_1507_0, i_8_398_1524_0,
    i_8_398_1533_0, i_8_398_1534_0, i_8_398_1535_0, i_8_398_1596_0,
    i_8_398_1597_0, i_8_398_1605_0, i_8_398_1606_0, i_8_398_1616_0,
    i_8_398_1660_0, i_8_398_1676_0, i_8_398_1681_0, i_8_398_1701_0,
    i_8_398_1733_0, i_8_398_1746_0, i_8_398_1779_0, i_8_398_1781_0,
    i_8_398_1782_0, i_8_398_1789_0, i_8_398_1790_0, i_8_398_1805_0,
    i_8_398_1806_0, i_8_398_1815_0, i_8_398_1821_0, i_8_398_1836_0,
    i_8_398_1837_0, i_8_398_1840_0, i_8_398_1844_0, i_8_398_1864_0,
    i_8_398_1891_0, i_8_398_1894_0, i_8_398_1901_0, i_8_398_1917_0,
    i_8_398_1919_0, i_8_398_1921_0, i_8_398_1951_0, i_8_398_1965_0,
    i_8_398_2053_0, i_8_398_2117_0, i_8_398_2127_0, i_8_398_2128_0,
    i_8_398_2169_0, i_8_398_2176_0, i_8_398_2179_0, i_8_398_2232_0,
    i_8_398_2244_0, i_8_398_2294_0, i_8_398_2297_0, i_8_398_2303_0,
    o_8_398_0_0  );
  input  i_8_398_19_0, i_8_398_109_0, i_8_398_139_0, i_8_398_238_0,
    i_8_398_300_0, i_8_398_310_0, i_8_398_372_0, i_8_398_373_0,
    i_8_398_375_0, i_8_398_381_0, i_8_398_383_0, i_8_398_419_0,
    i_8_398_431_0, i_8_398_460_0, i_8_398_463_0, i_8_398_479_0,
    i_8_398_480_0, i_8_398_506_0, i_8_398_510_0, i_8_398_529_0,
    i_8_398_549_0, i_8_398_552_0, i_8_398_553_0, i_8_398_590_0,
    i_8_398_603_0, i_8_398_606_0, i_8_398_613_0, i_8_398_706_0,
    i_8_398_796_0, i_8_398_858_0, i_8_398_867_0, i_8_398_868_0,
    i_8_398_878_0, i_8_398_976_0, i_8_398_991_0, i_8_398_1030_0,
    i_8_398_1084_0, i_8_398_1127_0, i_8_398_1130_0, i_8_398_1158_0,
    i_8_398_1188_0, i_8_398_1189_0, i_8_398_1192_0, i_8_398_1255_0,
    i_8_398_1279_0, i_8_398_1283_0, i_8_398_1325_0, i_8_398_1326_0,
    i_8_398_1327_0, i_8_398_1480_0, i_8_398_1507_0, i_8_398_1524_0,
    i_8_398_1533_0, i_8_398_1534_0, i_8_398_1535_0, i_8_398_1596_0,
    i_8_398_1597_0, i_8_398_1605_0, i_8_398_1606_0, i_8_398_1616_0,
    i_8_398_1660_0, i_8_398_1676_0, i_8_398_1681_0, i_8_398_1701_0,
    i_8_398_1733_0, i_8_398_1746_0, i_8_398_1779_0, i_8_398_1781_0,
    i_8_398_1782_0, i_8_398_1789_0, i_8_398_1790_0, i_8_398_1805_0,
    i_8_398_1806_0, i_8_398_1815_0, i_8_398_1821_0, i_8_398_1836_0,
    i_8_398_1837_0, i_8_398_1840_0, i_8_398_1844_0, i_8_398_1864_0,
    i_8_398_1891_0, i_8_398_1894_0, i_8_398_1901_0, i_8_398_1917_0,
    i_8_398_1919_0, i_8_398_1921_0, i_8_398_1951_0, i_8_398_1965_0,
    i_8_398_2053_0, i_8_398_2117_0, i_8_398_2127_0, i_8_398_2128_0,
    i_8_398_2169_0, i_8_398_2176_0, i_8_398_2179_0, i_8_398_2232_0,
    i_8_398_2244_0, i_8_398_2294_0, i_8_398_2297_0, i_8_398_2303_0;
  output o_8_398_0_0;
  assign o_8_398_0_0 = 0;
endmodule



// Benchmark "kernel_8_399" written by ABC on Sun Jul 19 10:10:02 2020

module kernel_8_399 ( 
    i_8_399_27_0, i_8_399_33_0, i_8_399_34_0, i_8_399_35_0, i_8_399_61_0,
    i_8_399_62_0, i_8_399_79_0, i_8_399_80_0, i_8_399_140_0, i_8_399_187_0,
    i_8_399_191_0, i_8_399_239_0, i_8_399_256_0, i_8_399_269_0,
    i_8_399_296_0, i_8_399_347_0, i_8_399_349_0, i_8_399_350_0,
    i_8_399_401_0, i_8_399_482_0, i_8_399_507_0, i_8_399_524_0,
    i_8_399_554_0, i_8_399_615_0, i_8_399_633_0, i_8_399_637_0,
    i_8_399_638_0, i_8_399_700_0, i_8_399_701_0, i_8_399_705_0,
    i_8_399_706_0, i_8_399_714_0, i_8_399_754_0, i_8_399_850_0,
    i_8_399_861_0, i_8_399_862_0, i_8_399_880_0, i_8_399_887_0,
    i_8_399_888_0, i_8_399_889_0, i_8_399_890_0, i_8_399_944_0,
    i_8_399_991_0, i_8_399_992_0, i_8_399_995_0, i_8_399_1016_0,
    i_8_399_1028_0, i_8_399_1050_0, i_8_399_1057_0, i_8_399_1060_0,
    i_8_399_1106_0, i_8_399_1131_0, i_8_399_1132_0, i_8_399_1157_0,
    i_8_399_1186_0, i_8_399_1187_0, i_8_399_1267_0, i_8_399_1268_0,
    i_8_399_1286_0, i_8_399_1297_0, i_8_399_1303_0, i_8_399_1322_0,
    i_8_399_1400_0, i_8_399_1483_0, i_8_399_1504_0, i_8_399_1505_0,
    i_8_399_1543_0, i_8_399_1545_0, i_8_399_1553_0, i_8_399_1556_0,
    i_8_399_1591_0, i_8_399_1648_0, i_8_399_1650_0, i_8_399_1690_0,
    i_8_399_1697_0, i_8_399_1751_0, i_8_399_1760_0, i_8_399_1762_0,
    i_8_399_1763_0, i_8_399_1857_0, i_8_399_1859_0, i_8_399_1886_0,
    i_8_399_1888_0, i_8_399_1898_0, i_8_399_1904_0, i_8_399_1949_0,
    i_8_399_1970_0, i_8_399_1985_0, i_8_399_1991_0, i_8_399_2015_0,
    i_8_399_2137_0, i_8_399_2146_0, i_8_399_2150_0, i_8_399_2159_0,
    i_8_399_2219_0, i_8_399_2241_0, i_8_399_2243_0, i_8_399_2248_0,
    i_8_399_2249_0, i_8_399_2263_0,
    o_8_399_0_0  );
  input  i_8_399_27_0, i_8_399_33_0, i_8_399_34_0, i_8_399_35_0,
    i_8_399_61_0, i_8_399_62_0, i_8_399_79_0, i_8_399_80_0, i_8_399_140_0,
    i_8_399_187_0, i_8_399_191_0, i_8_399_239_0, i_8_399_256_0,
    i_8_399_269_0, i_8_399_296_0, i_8_399_347_0, i_8_399_349_0,
    i_8_399_350_0, i_8_399_401_0, i_8_399_482_0, i_8_399_507_0,
    i_8_399_524_0, i_8_399_554_0, i_8_399_615_0, i_8_399_633_0,
    i_8_399_637_0, i_8_399_638_0, i_8_399_700_0, i_8_399_701_0,
    i_8_399_705_0, i_8_399_706_0, i_8_399_714_0, i_8_399_754_0,
    i_8_399_850_0, i_8_399_861_0, i_8_399_862_0, i_8_399_880_0,
    i_8_399_887_0, i_8_399_888_0, i_8_399_889_0, i_8_399_890_0,
    i_8_399_944_0, i_8_399_991_0, i_8_399_992_0, i_8_399_995_0,
    i_8_399_1016_0, i_8_399_1028_0, i_8_399_1050_0, i_8_399_1057_0,
    i_8_399_1060_0, i_8_399_1106_0, i_8_399_1131_0, i_8_399_1132_0,
    i_8_399_1157_0, i_8_399_1186_0, i_8_399_1187_0, i_8_399_1267_0,
    i_8_399_1268_0, i_8_399_1286_0, i_8_399_1297_0, i_8_399_1303_0,
    i_8_399_1322_0, i_8_399_1400_0, i_8_399_1483_0, i_8_399_1504_0,
    i_8_399_1505_0, i_8_399_1543_0, i_8_399_1545_0, i_8_399_1553_0,
    i_8_399_1556_0, i_8_399_1591_0, i_8_399_1648_0, i_8_399_1650_0,
    i_8_399_1690_0, i_8_399_1697_0, i_8_399_1751_0, i_8_399_1760_0,
    i_8_399_1762_0, i_8_399_1763_0, i_8_399_1857_0, i_8_399_1859_0,
    i_8_399_1886_0, i_8_399_1888_0, i_8_399_1898_0, i_8_399_1904_0,
    i_8_399_1949_0, i_8_399_1970_0, i_8_399_1985_0, i_8_399_1991_0,
    i_8_399_2015_0, i_8_399_2137_0, i_8_399_2146_0, i_8_399_2150_0,
    i_8_399_2159_0, i_8_399_2219_0, i_8_399_2241_0, i_8_399_2243_0,
    i_8_399_2248_0, i_8_399_2249_0, i_8_399_2263_0;
  output o_8_399_0_0;
  assign o_8_399_0_0 = ~((~i_8_399_1762_0 & ((~i_8_399_191_0 & ((i_8_399_700_0 & ~i_8_399_944_0 & ~i_8_399_1303_0 & ~i_8_399_1400_0 & i_8_399_1985_0) | (~i_8_399_296_0 & ~i_8_399_482_0 & ~i_8_399_861_0 & ~i_8_399_995_0 & i_8_399_1050_0 & ~i_8_399_1763_0 & ~i_8_399_1904_0 & ~i_8_399_2243_0))) | (~i_8_399_34_0 & ~i_8_399_35_0 & ~i_8_399_296_0 & i_8_399_554_0 & ~i_8_399_1186_0) | (~i_8_399_701_0 & ~i_8_399_861_0 & ~i_8_399_887_0 & ~i_8_399_1303_0 & ~i_8_399_1763_0 & ~i_8_399_2150_0 & ~i_8_399_2219_0 & ~i_8_399_2248_0))) | (~i_8_399_34_0 & ((~i_8_399_862_0 & i_8_399_1505_0 & ~i_8_399_2159_0) | (~i_8_399_33_0 & ~i_8_399_633_0 & ~i_8_399_1157_0 & i_8_399_1556_0 & ~i_8_399_1591_0 & ~i_8_399_2243_0))) | (~i_8_399_35_0 & ((~i_8_399_33_0 & i_8_399_706_0 & ~i_8_399_862_0 & ~i_8_399_1016_0 & ~i_8_399_1648_0 & ~i_8_399_1650_0 & ~i_8_399_1763_0) | (i_8_399_79_0 & i_8_399_350_0 & ~i_8_399_1591_0 & ~i_8_399_1949_0 & ~i_8_399_1985_0 & ~i_8_399_2263_0))) | (~i_8_399_701_0 & ((~i_8_399_191_0 & ((~i_8_399_700_0 & ~i_8_399_862_0 & i_8_399_1553_0) | (~i_8_399_861_0 & ~i_8_399_880_0 & ~i_8_399_1187_0 & ~i_8_399_1267_0 & ~i_8_399_1763_0 & ~i_8_399_1888_0 & ~i_8_399_2159_0))) | (~i_8_399_638_0 & ~i_8_399_700_0 & ~i_8_399_861_0 & ~i_8_399_1186_0 & ~i_8_399_2146_0 & ~i_8_399_2150_0 & ~i_8_399_2248_0))) | (~i_8_399_633_0 & ((~i_8_399_637_0 & i_8_399_1543_0 & ~i_8_399_1591_0) | (i_8_399_706_0 & ~i_8_399_1648_0 & i_8_399_1886_0))) | (~i_8_399_637_0 & ((~i_8_399_61_0 & ~i_8_399_62_0 & ~i_8_399_638_0 & ~i_8_399_888_0 & ~i_8_399_890_0 & ~i_8_399_1187_0) | (~i_8_399_80_0 & i_8_399_1016_0 & ~i_8_399_1050_0 & ~i_8_399_1400_0 & ~i_8_399_2241_0))) | (~i_8_399_2137_0 & ((~i_8_399_61_0 & ~i_8_399_62_0 & ((~i_8_399_80_0 & ~i_8_399_887_0 & ~i_8_399_888_0 & ~i_8_399_1186_0 & ~i_8_399_1751_0 & ~i_8_399_1760_0) | (i_8_399_637_0 & ~i_8_399_850_0 & ~i_8_399_889_0 & ~i_8_399_944_0 & ~i_8_399_2159_0))) | (~i_8_399_887_0 & ~i_8_399_888_0 & ~i_8_399_80_0 & ~i_8_399_482_0 & ~i_8_399_995_0 & ~i_8_399_1591_0 & ~i_8_399_1763_0 & ~i_8_399_1857_0 & ~i_8_399_1970_0))) | (i_8_399_754_0 & ((~i_8_399_62_0 & ~i_8_399_861_0 & ~i_8_399_889_0 & ~i_8_399_2243_0) | (~i_8_399_33_0 & i_8_399_861_0 & ~i_8_399_2248_0))) | (~i_8_399_62_0 & ((~i_8_399_862_0 & ~i_8_399_890_0 & ~i_8_399_1286_0 & ~i_8_399_1591_0 & i_8_399_2150_0) | (i_8_399_349_0 & ~i_8_399_1132_0 & i_8_399_1888_0 & ~i_8_399_2219_0 & ~i_8_399_2243_0))) | (~i_8_399_1050_0 & ~i_8_399_2263_0 & ((~i_8_399_33_0 & ~i_8_399_347_0 & ~i_8_399_714_0 & ~i_8_399_1268_0 & ~i_8_399_1763_0 & i_8_399_1888_0) | (~i_8_399_889_0 & ~i_8_399_1504_0 & i_8_399_2146_0 & ~i_8_399_2219_0 & ~i_8_399_2249_0))) | (~i_8_399_33_0 & ((i_8_399_524_0 & ~i_8_399_1763_0) | (~i_8_399_507_0 & i_8_399_633_0 & ~i_8_399_862_0 & ~i_8_399_1545_0 & ~i_8_399_1949_0 & ~i_8_399_2159_0) | (~i_8_399_61_0 & i_8_399_1057_0 & ~i_8_399_1187_0 & i_8_399_1591_0 & ~i_8_399_2249_0))) | (~i_8_399_700_0 & ~i_8_399_1060_0 & i_8_399_1131_0) | (~i_8_399_1057_0 & ~i_8_399_1286_0 & i_8_399_1504_0 & ~i_8_399_1543_0 & ~i_8_399_1857_0) | (i_8_399_1132_0 & i_8_399_1904_0));
endmodule



// Benchmark "kernel_8_400" written by ABC on Sun Jul 19 10:10:03 2020

module kernel_8_400 ( 
    i_8_400_9_0, i_8_400_12_0, i_8_400_20_0, i_8_400_50_0, i_8_400_74_0,
    i_8_400_101_0, i_8_400_140_0, i_8_400_149_0, i_8_400_165_0,
    i_8_400_254_0, i_8_400_290_0, i_8_400_299_0, i_8_400_304_0,
    i_8_400_362_0, i_8_400_364_0, i_8_400_379_0, i_8_400_380_0,
    i_8_400_423_0, i_8_400_424_0, i_8_400_490_0, i_8_400_554_0,
    i_8_400_578_0, i_8_400_582_0, i_8_400_583_0, i_8_400_598_0,
    i_8_400_605_0, i_8_400_640_0, i_8_400_650_0, i_8_400_653_0,
    i_8_400_677_0, i_8_400_679_0, i_8_400_695_0, i_8_400_697_0,
    i_8_400_731_0, i_8_400_775_0, i_8_400_776_0, i_8_400_787_0,
    i_8_400_794_0, i_8_400_803_0, i_8_400_842_0, i_8_400_850_0,
    i_8_400_878_0, i_8_400_883_0, i_8_400_936_0, i_8_400_965_0,
    i_8_400_971_0, i_8_400_1037_0, i_8_400_1199_0, i_8_400_1231_0,
    i_8_400_1255_0, i_8_400_1271_0, i_8_400_1282_0, i_8_400_1299_0,
    i_8_400_1313_0, i_8_400_1316_0, i_8_400_1339_0, i_8_400_1345_0,
    i_8_400_1378_0, i_8_400_1397_0, i_8_400_1433_0, i_8_400_1457_0,
    i_8_400_1471_0, i_8_400_1538_0, i_8_400_1557_0, i_8_400_1571_0,
    i_8_400_1607_0, i_8_400_1622_0, i_8_400_1629_0, i_8_400_1703_0,
    i_8_400_1715_0, i_8_400_1750_0, i_8_400_1755_0, i_8_400_1756_0,
    i_8_400_1768_0, i_8_400_1777_0, i_8_400_1791_0, i_8_400_1818_0,
    i_8_400_1819_0, i_8_400_1823_0, i_8_400_1832_0, i_8_400_1888_0,
    i_8_400_1973_0, i_8_400_1981_0, i_8_400_1993_0, i_8_400_2052_0,
    i_8_400_2054_0, i_8_400_2072_0, i_8_400_2099_0, i_8_400_2106_0,
    i_8_400_2108_0, i_8_400_2135_0, i_8_400_2143_0, i_8_400_2155_0,
    i_8_400_2170_0, i_8_400_2188_0, i_8_400_2230_0, i_8_400_2243_0,
    i_8_400_2264_0, i_8_400_2295_0, i_8_400_2298_0,
    o_8_400_0_0  );
  input  i_8_400_9_0, i_8_400_12_0, i_8_400_20_0, i_8_400_50_0,
    i_8_400_74_0, i_8_400_101_0, i_8_400_140_0, i_8_400_149_0,
    i_8_400_165_0, i_8_400_254_0, i_8_400_290_0, i_8_400_299_0,
    i_8_400_304_0, i_8_400_362_0, i_8_400_364_0, i_8_400_379_0,
    i_8_400_380_0, i_8_400_423_0, i_8_400_424_0, i_8_400_490_0,
    i_8_400_554_0, i_8_400_578_0, i_8_400_582_0, i_8_400_583_0,
    i_8_400_598_0, i_8_400_605_0, i_8_400_640_0, i_8_400_650_0,
    i_8_400_653_0, i_8_400_677_0, i_8_400_679_0, i_8_400_695_0,
    i_8_400_697_0, i_8_400_731_0, i_8_400_775_0, i_8_400_776_0,
    i_8_400_787_0, i_8_400_794_0, i_8_400_803_0, i_8_400_842_0,
    i_8_400_850_0, i_8_400_878_0, i_8_400_883_0, i_8_400_936_0,
    i_8_400_965_0, i_8_400_971_0, i_8_400_1037_0, i_8_400_1199_0,
    i_8_400_1231_0, i_8_400_1255_0, i_8_400_1271_0, i_8_400_1282_0,
    i_8_400_1299_0, i_8_400_1313_0, i_8_400_1316_0, i_8_400_1339_0,
    i_8_400_1345_0, i_8_400_1378_0, i_8_400_1397_0, i_8_400_1433_0,
    i_8_400_1457_0, i_8_400_1471_0, i_8_400_1538_0, i_8_400_1557_0,
    i_8_400_1571_0, i_8_400_1607_0, i_8_400_1622_0, i_8_400_1629_0,
    i_8_400_1703_0, i_8_400_1715_0, i_8_400_1750_0, i_8_400_1755_0,
    i_8_400_1756_0, i_8_400_1768_0, i_8_400_1777_0, i_8_400_1791_0,
    i_8_400_1818_0, i_8_400_1819_0, i_8_400_1823_0, i_8_400_1832_0,
    i_8_400_1888_0, i_8_400_1973_0, i_8_400_1981_0, i_8_400_1993_0,
    i_8_400_2052_0, i_8_400_2054_0, i_8_400_2072_0, i_8_400_2099_0,
    i_8_400_2106_0, i_8_400_2108_0, i_8_400_2135_0, i_8_400_2143_0,
    i_8_400_2155_0, i_8_400_2170_0, i_8_400_2188_0, i_8_400_2230_0,
    i_8_400_2243_0, i_8_400_2264_0, i_8_400_2295_0, i_8_400_2298_0;
  output o_8_400_0_0;
  assign o_8_400_0_0 = 0;
endmodule



// Benchmark "kernel_8_401" written by ABC on Sun Jul 19 10:10:04 2020

module kernel_8_401 ( 
    i_8_401_30_0, i_8_401_31_0, i_8_401_84_0, i_8_401_88_0, i_8_401_111_0,
    i_8_401_114_0, i_8_401_165_0, i_8_401_238_0, i_8_401_240_0,
    i_8_401_372_0, i_8_401_386_0, i_8_401_390_0, i_8_401_421_0,
    i_8_401_427_0, i_8_401_437_0, i_8_401_474_0, i_8_401_475_0,
    i_8_401_483_0, i_8_401_520_0, i_8_401_522_0, i_8_401_540_0,
    i_8_401_553_0, i_8_401_571_0, i_8_401_574_0, i_8_401_598_0,
    i_8_401_606_0, i_8_401_633_0, i_8_401_693_0, i_8_401_694_0,
    i_8_401_706_0, i_8_401_709_0, i_8_401_712_0, i_8_401_759_0,
    i_8_401_762_0, i_8_401_763_0, i_8_401_778_0, i_8_401_799_0,
    i_8_401_839_0, i_8_401_888_0, i_8_401_940_0, i_8_401_943_0,
    i_8_401_966_0, i_8_401_994_0, i_8_401_1056_0, i_8_401_1059_0,
    i_8_401_1090_0, i_8_401_1102_0, i_8_401_1182_0, i_8_401_1185_0,
    i_8_401_1281_0, i_8_401_1293_0, i_8_401_1300_0, i_8_401_1305_0,
    i_8_401_1309_0, i_8_401_1318_0, i_8_401_1345_0, i_8_401_1390_0,
    i_8_401_1438_0, i_8_401_1516_0, i_8_401_1533_0, i_8_401_1534_0,
    i_8_401_1563_0, i_8_401_1590_0, i_8_401_1603_0, i_8_401_1614_0,
    i_8_401_1624_0, i_8_401_1654_0, i_8_401_1686_0, i_8_401_1690_0,
    i_8_401_1731_0, i_8_401_1735_0, i_8_401_1747_0, i_8_401_1749_0,
    i_8_401_1751_0, i_8_401_1753_0, i_8_401_1762_0, i_8_401_1780_0,
    i_8_401_1789_0, i_8_401_1804_0, i_8_401_1824_0, i_8_401_1825_0,
    i_8_401_1831_0, i_8_401_1917_0, i_8_401_1929_0, i_8_401_1996_0,
    i_8_401_2019_0, i_8_401_2047_0, i_8_401_2058_0, i_8_401_2077_0,
    i_8_401_2118_0, i_8_401_2122_0, i_8_401_2124_0, i_8_401_2142_0,
    i_8_401_2150_0, i_8_401_2173_0, i_8_401_2224_0, i_8_401_2260_0,
    i_8_401_2290_0, i_8_401_2295_0, i_8_401_2299_0,
    o_8_401_0_0  );
  input  i_8_401_30_0, i_8_401_31_0, i_8_401_84_0, i_8_401_88_0,
    i_8_401_111_0, i_8_401_114_0, i_8_401_165_0, i_8_401_238_0,
    i_8_401_240_0, i_8_401_372_0, i_8_401_386_0, i_8_401_390_0,
    i_8_401_421_0, i_8_401_427_0, i_8_401_437_0, i_8_401_474_0,
    i_8_401_475_0, i_8_401_483_0, i_8_401_520_0, i_8_401_522_0,
    i_8_401_540_0, i_8_401_553_0, i_8_401_571_0, i_8_401_574_0,
    i_8_401_598_0, i_8_401_606_0, i_8_401_633_0, i_8_401_693_0,
    i_8_401_694_0, i_8_401_706_0, i_8_401_709_0, i_8_401_712_0,
    i_8_401_759_0, i_8_401_762_0, i_8_401_763_0, i_8_401_778_0,
    i_8_401_799_0, i_8_401_839_0, i_8_401_888_0, i_8_401_940_0,
    i_8_401_943_0, i_8_401_966_0, i_8_401_994_0, i_8_401_1056_0,
    i_8_401_1059_0, i_8_401_1090_0, i_8_401_1102_0, i_8_401_1182_0,
    i_8_401_1185_0, i_8_401_1281_0, i_8_401_1293_0, i_8_401_1300_0,
    i_8_401_1305_0, i_8_401_1309_0, i_8_401_1318_0, i_8_401_1345_0,
    i_8_401_1390_0, i_8_401_1438_0, i_8_401_1516_0, i_8_401_1533_0,
    i_8_401_1534_0, i_8_401_1563_0, i_8_401_1590_0, i_8_401_1603_0,
    i_8_401_1614_0, i_8_401_1624_0, i_8_401_1654_0, i_8_401_1686_0,
    i_8_401_1690_0, i_8_401_1731_0, i_8_401_1735_0, i_8_401_1747_0,
    i_8_401_1749_0, i_8_401_1751_0, i_8_401_1753_0, i_8_401_1762_0,
    i_8_401_1780_0, i_8_401_1789_0, i_8_401_1804_0, i_8_401_1824_0,
    i_8_401_1825_0, i_8_401_1831_0, i_8_401_1917_0, i_8_401_1929_0,
    i_8_401_1996_0, i_8_401_2019_0, i_8_401_2047_0, i_8_401_2058_0,
    i_8_401_2077_0, i_8_401_2118_0, i_8_401_2122_0, i_8_401_2124_0,
    i_8_401_2142_0, i_8_401_2150_0, i_8_401_2173_0, i_8_401_2224_0,
    i_8_401_2260_0, i_8_401_2290_0, i_8_401_2295_0, i_8_401_2299_0;
  output o_8_401_0_0;
  assign o_8_401_0_0 = 0;
endmodule



// Benchmark "kernel_8_402" written by ABC on Sun Jul 19 10:10:05 2020

module kernel_8_402 ( 
    i_8_402_55_0, i_8_402_78_0, i_8_402_95_0, i_8_402_97_0, i_8_402_105_0,
    i_8_402_106_0, i_8_402_107_0, i_8_402_141_0, i_8_402_220_0,
    i_8_402_223_0, i_8_402_228_0, i_8_402_229_0, i_8_402_256_0,
    i_8_402_276_0, i_8_402_379_0, i_8_402_492_0, i_8_402_573_0,
    i_8_402_580_0, i_8_402_583_0, i_8_402_597_0, i_8_402_636_0,
    i_8_402_658_0, i_8_402_661_0, i_8_402_663_0, i_8_402_664_0,
    i_8_402_672_0, i_8_402_700_0, i_8_402_704_0, i_8_402_733_0,
    i_8_402_763_0, i_8_402_781_0, i_8_402_822_0, i_8_402_858_0,
    i_8_402_861_0, i_8_402_871_0, i_8_402_894_0, i_8_402_925_0,
    i_8_402_969_0, i_8_402_975_0, i_8_402_976_0, i_8_402_1107_0,
    i_8_402_1108_0, i_8_402_1122_0, i_8_402_1228_0, i_8_402_1237_0,
    i_8_402_1272_0, i_8_402_1302_0, i_8_402_1322_0, i_8_402_1348_0,
    i_8_402_1393_0, i_8_402_1470_0, i_8_402_1473_0, i_8_402_1479_0,
    i_8_402_1483_0, i_8_402_1506_0, i_8_402_1509_0, i_8_402_1524_0,
    i_8_402_1561_0, i_8_402_1563_0, i_8_402_1606_0, i_8_402_1617_0,
    i_8_402_1618_0, i_8_402_1620_0, i_8_402_1677_0, i_8_402_1700_0,
    i_8_402_1702_0, i_8_402_1704_0, i_8_402_1750_0, i_8_402_1771_0,
    i_8_402_1785_0, i_8_402_1786_0, i_8_402_1810_0, i_8_402_1812_0,
    i_8_402_1833_0, i_8_402_1842_0, i_8_402_1866_0, i_8_402_1878_0,
    i_8_402_1885_0, i_8_402_1947_0, i_8_402_1949_0, i_8_402_1962_0,
    i_8_402_1965_0, i_8_402_1968_0, i_8_402_1974_0, i_8_402_1983_0,
    i_8_402_1986_0, i_8_402_1988_0, i_8_402_1992_0, i_8_402_2055_0,
    i_8_402_2112_0, i_8_402_2148_0, i_8_402_2154_0, i_8_402_2172_0,
    i_8_402_2175_0, i_8_402_2185_0, i_8_402_2188_0, i_8_402_2202_0,
    i_8_402_2229_0, i_8_402_2262_0, i_8_402_2278_0,
    o_8_402_0_0  );
  input  i_8_402_55_0, i_8_402_78_0, i_8_402_95_0, i_8_402_97_0,
    i_8_402_105_0, i_8_402_106_0, i_8_402_107_0, i_8_402_141_0,
    i_8_402_220_0, i_8_402_223_0, i_8_402_228_0, i_8_402_229_0,
    i_8_402_256_0, i_8_402_276_0, i_8_402_379_0, i_8_402_492_0,
    i_8_402_573_0, i_8_402_580_0, i_8_402_583_0, i_8_402_597_0,
    i_8_402_636_0, i_8_402_658_0, i_8_402_661_0, i_8_402_663_0,
    i_8_402_664_0, i_8_402_672_0, i_8_402_700_0, i_8_402_704_0,
    i_8_402_733_0, i_8_402_763_0, i_8_402_781_0, i_8_402_822_0,
    i_8_402_858_0, i_8_402_861_0, i_8_402_871_0, i_8_402_894_0,
    i_8_402_925_0, i_8_402_969_0, i_8_402_975_0, i_8_402_976_0,
    i_8_402_1107_0, i_8_402_1108_0, i_8_402_1122_0, i_8_402_1228_0,
    i_8_402_1237_0, i_8_402_1272_0, i_8_402_1302_0, i_8_402_1322_0,
    i_8_402_1348_0, i_8_402_1393_0, i_8_402_1470_0, i_8_402_1473_0,
    i_8_402_1479_0, i_8_402_1483_0, i_8_402_1506_0, i_8_402_1509_0,
    i_8_402_1524_0, i_8_402_1561_0, i_8_402_1563_0, i_8_402_1606_0,
    i_8_402_1617_0, i_8_402_1618_0, i_8_402_1620_0, i_8_402_1677_0,
    i_8_402_1700_0, i_8_402_1702_0, i_8_402_1704_0, i_8_402_1750_0,
    i_8_402_1771_0, i_8_402_1785_0, i_8_402_1786_0, i_8_402_1810_0,
    i_8_402_1812_0, i_8_402_1833_0, i_8_402_1842_0, i_8_402_1866_0,
    i_8_402_1878_0, i_8_402_1885_0, i_8_402_1947_0, i_8_402_1949_0,
    i_8_402_1962_0, i_8_402_1965_0, i_8_402_1968_0, i_8_402_1974_0,
    i_8_402_1983_0, i_8_402_1986_0, i_8_402_1988_0, i_8_402_1992_0,
    i_8_402_2055_0, i_8_402_2112_0, i_8_402_2148_0, i_8_402_2154_0,
    i_8_402_2172_0, i_8_402_2175_0, i_8_402_2185_0, i_8_402_2188_0,
    i_8_402_2202_0, i_8_402_2229_0, i_8_402_2262_0, i_8_402_2278_0;
  output o_8_402_0_0;
  assign o_8_402_0_0 = ~((~i_8_402_2188_0 & ((~i_8_402_106_0 & ((i_8_402_220_0 & ~i_8_402_663_0 & ((~i_8_402_78_0 & ~i_8_402_672_0 & i_8_402_1237_0 & ~i_8_402_1483_0 & ~i_8_402_1988_0) | (i_8_402_658_0 & ~i_8_402_1704_0 & ~i_8_402_1949_0 & ~i_8_402_1965_0 & ~i_8_402_2055_0))) | (~i_8_402_55_0 & ~i_8_402_573_0 & ~i_8_402_583_0 & ~i_8_402_672_0 & ~i_8_402_763_0 & ~i_8_402_858_0 & ~i_8_402_871_0 & ~i_8_402_1322_0 & ~i_8_402_1563_0 & ~i_8_402_1968_0 & i_8_402_1992_0))) | (~i_8_402_1563_0 & ((~i_8_402_276_0 & ((~i_8_402_105_0 & ~i_8_402_256_0 & ~i_8_402_658_0 & ~i_8_402_969_0 & ~i_8_402_1322_0 & ~i_8_402_1810_0 & ~i_8_402_1947_0 & ~i_8_402_1962_0 & ~i_8_402_1965_0 & ~i_8_402_1986_0) | (~i_8_402_573_0 & ~i_8_402_733_0 & ~i_8_402_1272_0 & ~i_8_402_1302_0 & ~i_8_402_1470_0 & ~i_8_402_1473_0 & ~i_8_402_1506_0 & ~i_8_402_1617_0 & ~i_8_402_1704_0 & ~i_8_402_2172_0 & ~i_8_402_2202_0 & ~i_8_402_2262_0))) | (~i_8_402_78_0 & i_8_402_223_0 & ~i_8_402_664_0 & ~i_8_402_1107_0 & ~i_8_402_1272_0 & ~i_8_402_1302_0 & i_8_402_1677_0 & ~i_8_402_1810_0 & ~i_8_402_2202_0))) | (~i_8_402_78_0 & ((~i_8_402_871_0 & ~i_8_402_2278_0 & ((i_8_402_492_0 & i_8_402_1108_0 & ~i_8_402_1470_0 & ~i_8_402_1524_0 & ~i_8_402_2175_0) | (~i_8_402_223_0 & ~i_8_402_858_0 & ~i_8_402_1122_0 & ~i_8_402_1479_0 & ~i_8_402_1509_0 & ~i_8_402_1812_0 & ~i_8_402_1866_0 & ~i_8_402_1878_0 & ~i_8_402_2112_0 & ~i_8_402_2154_0 & ~i_8_402_2262_0))) | (~i_8_402_1272_0 & ~i_8_402_1302_0 & ~i_8_402_228_0 & ~i_8_402_861_0 & ~i_8_402_1470_0 & ~i_8_402_1479_0 & ~i_8_402_1606_0 & ~i_8_402_1810_0 & ~i_8_402_1866_0))) | (i_8_402_661_0 & i_8_402_664_0 & ~i_8_402_1302_0 & ~i_8_402_1479_0 & ~i_8_402_1506_0 & ~i_8_402_1949_0 & ~i_8_402_2172_0))) | (~i_8_402_2172_0 & ((~i_8_402_1483_0 & ((~i_8_402_55_0 & ~i_8_402_106_0 & ~i_8_402_1810_0 & ((~i_8_402_105_0 & ~i_8_402_636_0 & ~i_8_402_700_0 & ~i_8_402_733_0 & ~i_8_402_822_0 & ~i_8_402_1107_0 & ~i_8_402_1322_0 & ~i_8_402_1620_0 & ~i_8_402_1949_0) | (~i_8_402_256_0 & ~i_8_402_597_0 & ~i_8_402_664_0 & ~i_8_402_858_0 & ~i_8_402_1122_0 & ~i_8_402_1618_0 & ~i_8_402_1771_0 & i_8_402_1785_0 & ~i_8_402_2112_0 & ~i_8_402_2229_0))) | (~i_8_402_223_0 & ~i_8_402_1509_0 & ~i_8_402_1606_0 & ~i_8_402_1866_0 & ~i_8_402_1965_0 & i_8_402_2148_0))) | (~i_8_402_1302_0 & ~i_8_402_1947_0 & ~i_8_402_2202_0 & ((~i_8_402_573_0 & i_8_402_597_0 & ~i_8_402_663_0 & ~i_8_402_1108_0 & ~i_8_402_1393_0 & ~i_8_402_1563_0 & ~i_8_402_1700_0) | (~i_8_402_858_0 & ~i_8_402_871_0 & ~i_8_402_894_0 & ~i_8_402_1506_0 & ~i_8_402_1785_0 & ~i_8_402_1866_0 & ~i_8_402_2175_0))) | (~i_8_402_78_0 & ~i_8_402_1322_0 & i_8_402_1885_0 & ~i_8_402_2055_0 & ~i_8_402_2278_0))) | (~i_8_402_105_0 & ((~i_8_402_228_0 & ~i_8_402_733_0 & ~i_8_402_822_0 & ~i_8_402_858_0 & ~i_8_402_871_0 & ~i_8_402_1302_0 & ~i_8_402_1470_0 & ~i_8_402_2154_0 & ~i_8_402_2229_0) | (i_8_402_223_0 & ~i_8_402_573_0 & ~i_8_402_763_0 & ~i_8_402_1108_0 & ~i_8_402_1563_0 & ~i_8_402_1618_0 & ~i_8_402_1842_0 & ~i_8_402_1878_0 & ~i_8_402_1965_0 & i_8_402_2148_0 & ~i_8_402_2262_0))) | (~i_8_402_228_0 & ((~i_8_402_78_0 & ~i_8_402_220_0 & i_8_402_1237_0 & ~i_8_402_1393_0 & ~i_8_402_1509_0) | (~i_8_402_636_0 & ~i_8_402_763_0 & ~i_8_402_861_0 & ~i_8_402_1228_0 & ~i_8_402_1470_0 & ~i_8_402_1524_0 & ~i_8_402_1561_0 & ~i_8_402_1606_0 & ~i_8_402_1878_0 & ~i_8_402_2154_0 & ~i_8_402_2278_0))) | (~i_8_402_858_0 & ((~i_8_402_55_0 & ~i_8_402_1833_0 & ((~i_8_402_78_0 & ~i_8_402_663_0 & ~i_8_402_871_0 & ~i_8_402_1617_0 & ~i_8_402_1618_0 & ~i_8_402_1704_0 & ~i_8_402_1750_0 & i_8_402_1786_0) | (~i_8_402_220_0 & ~i_8_402_573_0 & ~i_8_402_597_0 & ~i_8_402_636_0 & ~i_8_402_733_0 & ~i_8_402_1483_0 & ~i_8_402_1606_0 & ~i_8_402_2229_0))) | (~i_8_402_379_0 & ((i_8_402_106_0 & ~i_8_402_1237_0 & ~i_8_402_1947_0 & i_8_402_1968_0 & ~i_8_402_2112_0) | (~i_8_402_78_0 & ~i_8_402_220_0 & ~i_8_402_1302_0 & ~i_8_402_1618_0 & ~i_8_402_1810_0 & ~i_8_402_1988_0 & ~i_8_402_2055_0 & ~i_8_402_2202_0))) | (~i_8_402_733_0 & ((~i_8_402_861_0 & i_8_402_1509_0 & ~i_8_402_1866_0 & ~i_8_402_1947_0 & ~i_8_402_1949_0 & i_8_402_1986_0 & i_8_402_2175_0) | (~i_8_402_223_0 & ~i_8_402_672_0 & ~i_8_402_871_0 & ~i_8_402_1107_0 & ~i_8_402_1228_0 & ~i_8_402_1272_0 & ~i_8_402_1483_0 & ~i_8_402_1563_0 & ~i_8_402_1771_0 & ~i_8_402_1842_0 & ~i_8_402_2185_0 & ~i_8_402_2278_0))) | (~i_8_402_1771_0 & ((i_8_402_658_0 & ~i_8_402_781_0 & ~i_8_402_822_0 & ~i_8_402_1479_0 & ~i_8_402_1810_0 & ~i_8_402_1988_0) | (~i_8_402_95_0 & ~i_8_402_636_0 & ~i_8_402_894_0 & ~i_8_402_1302_0 & ~i_8_402_1606_0 & ~i_8_402_1677_0 & ~i_8_402_1785_0 & ~i_8_402_2154_0))))) | (~i_8_402_223_0 & ((~i_8_402_55_0 & ~i_8_402_276_0 & ~i_8_402_379_0 & ~i_8_402_733_0 & ~i_8_402_976_0 & ~i_8_402_1506_0 & ~i_8_402_1677_0 & ~i_8_402_1750_0 & ~i_8_402_2055_0) | (~i_8_402_78_0 & ~i_8_402_861_0 & ~i_8_402_975_0 & ~i_8_402_1108_0 & ~i_8_402_1122_0 & i_8_402_1506_0 & ~i_8_402_1704_0 & ~i_8_402_1810_0 & ~i_8_402_2278_0))) | (~i_8_402_861_0 & ~i_8_402_1108_0 & ~i_8_402_1878_0 & ((i_8_402_97_0 & ~i_8_402_925_0 & ~i_8_402_1302_0 & i_8_402_1750_0 & ~i_8_402_2148_0 & ~i_8_402_2154_0) | (~i_8_402_1750_0 & ~i_8_402_1771_0 & ~i_8_402_1947_0 & i_8_402_1983_0 & ~i_8_402_2175_0))) | (~i_8_402_1107_0 & ((~i_8_402_379_0 & ~i_8_402_597_0 & ~i_8_402_672_0 & ~i_8_402_1561_0 & ~i_8_402_1563_0 & ~i_8_402_1617_0 & ~i_8_402_1618_0 & ~i_8_402_1677_0 & i_8_402_1771_0 & ~i_8_402_2202_0) | (~i_8_402_781_0 & ~i_8_402_1302_0 & ~i_8_402_1322_0 & ~i_8_402_1348_0 & ~i_8_402_1470_0 & ~i_8_402_1750_0 & ~i_8_402_1947_0 & ~i_8_402_2229_0))) | (~i_8_402_1348_0 & ~i_8_402_1470_0 & ~i_8_402_1866_0 & ((~i_8_402_573_0 & ~i_8_402_733_0 & ~i_8_402_871_0 & ~i_8_402_1122_0 & ~i_8_402_1509_0 & ~i_8_402_1606_0 & i_8_402_1786_0 & ~i_8_402_2229_0) | (i_8_402_658_0 & i_8_402_1107_0 & i_8_402_1228_0 & ~i_8_402_1677_0 & ~i_8_402_2175_0 & ~i_8_402_2278_0))) | (i_8_402_379_0 & ~i_8_402_663_0 & ~i_8_402_763_0 & ~i_8_402_1393_0 & ~i_8_402_1473_0 & ~i_8_402_1479_0 & ~i_8_402_1506_0 & ~i_8_402_1606_0 & ~i_8_402_1704_0 & ~i_8_402_1750_0));
endmodule



// Benchmark "kernel_8_403" written by ABC on Sun Jul 19 10:10:07 2020

module kernel_8_403 ( 
    i_8_403_25_0, i_8_403_39_0, i_8_403_51_0, i_8_403_66_0, i_8_403_67_0,
    i_8_403_143_0, i_8_403_195_0, i_8_403_219_0, i_8_403_228_0,
    i_8_403_230_0, i_8_403_267_0, i_8_403_269_0, i_8_403_286_0,
    i_8_403_287_0, i_8_403_313_0, i_8_403_402_0, i_8_403_403_0,
    i_8_403_423_0, i_8_403_467_0, i_8_403_492_0, i_8_403_522_0,
    i_8_403_526_0, i_8_403_527_0, i_8_403_551_0, i_8_403_582_0,
    i_8_403_583_0, i_8_403_588_0, i_8_403_619_0, i_8_403_652_0,
    i_8_403_654_0, i_8_403_665_0, i_8_403_703_0, i_8_403_726_0,
    i_8_403_807_0, i_8_403_823_0, i_8_403_840_0, i_8_403_843_0,
    i_8_403_844_0, i_8_403_876_0, i_8_403_883_0, i_8_403_886_0,
    i_8_403_897_0, i_8_403_898_0, i_8_403_922_0, i_8_403_924_0,
    i_8_403_930_0, i_8_403_931_0, i_8_403_933_0, i_8_403_964_0,
    i_8_403_978_0, i_8_403_979_0, i_8_403_980_0, i_8_403_1030_0,
    i_8_403_1074_0, i_8_403_1276_0, i_8_403_1307_0, i_8_403_1428_0,
    i_8_403_1429_0, i_8_403_1438_0, i_8_403_1446_0, i_8_403_1447_0,
    i_8_403_1455_0, i_8_403_1534_0, i_8_403_1535_0, i_8_403_1599_0,
    i_8_403_1624_0, i_8_403_1632_0, i_8_403_1671_0, i_8_403_1672_0,
    i_8_403_1725_0, i_8_403_1733_0, i_8_403_1744_0, i_8_403_1748_0,
    i_8_403_1773_0, i_8_403_1774_0, i_8_403_1803_0, i_8_403_1857_0,
    i_8_403_1903_0, i_8_403_1941_0, i_8_403_1950_0, i_8_403_1962_0,
    i_8_403_1968_0, i_8_403_1969_0, i_8_403_2004_0, i_8_403_2100_0,
    i_8_403_2104_0, i_8_403_2143_0, i_8_403_2158_0, i_8_403_2172_0,
    i_8_403_2174_0, i_8_403_2175_0, i_8_403_2176_0, i_8_403_2177_0,
    i_8_403_2209_0, i_8_403_2233_0, i_8_403_2245_0, i_8_403_2262_0,
    i_8_403_2263_0, i_8_403_2265_0, i_8_403_2271_0,
    o_8_403_0_0  );
  input  i_8_403_25_0, i_8_403_39_0, i_8_403_51_0, i_8_403_66_0,
    i_8_403_67_0, i_8_403_143_0, i_8_403_195_0, i_8_403_219_0,
    i_8_403_228_0, i_8_403_230_0, i_8_403_267_0, i_8_403_269_0,
    i_8_403_286_0, i_8_403_287_0, i_8_403_313_0, i_8_403_402_0,
    i_8_403_403_0, i_8_403_423_0, i_8_403_467_0, i_8_403_492_0,
    i_8_403_522_0, i_8_403_526_0, i_8_403_527_0, i_8_403_551_0,
    i_8_403_582_0, i_8_403_583_0, i_8_403_588_0, i_8_403_619_0,
    i_8_403_652_0, i_8_403_654_0, i_8_403_665_0, i_8_403_703_0,
    i_8_403_726_0, i_8_403_807_0, i_8_403_823_0, i_8_403_840_0,
    i_8_403_843_0, i_8_403_844_0, i_8_403_876_0, i_8_403_883_0,
    i_8_403_886_0, i_8_403_897_0, i_8_403_898_0, i_8_403_922_0,
    i_8_403_924_0, i_8_403_930_0, i_8_403_931_0, i_8_403_933_0,
    i_8_403_964_0, i_8_403_978_0, i_8_403_979_0, i_8_403_980_0,
    i_8_403_1030_0, i_8_403_1074_0, i_8_403_1276_0, i_8_403_1307_0,
    i_8_403_1428_0, i_8_403_1429_0, i_8_403_1438_0, i_8_403_1446_0,
    i_8_403_1447_0, i_8_403_1455_0, i_8_403_1534_0, i_8_403_1535_0,
    i_8_403_1599_0, i_8_403_1624_0, i_8_403_1632_0, i_8_403_1671_0,
    i_8_403_1672_0, i_8_403_1725_0, i_8_403_1733_0, i_8_403_1744_0,
    i_8_403_1748_0, i_8_403_1773_0, i_8_403_1774_0, i_8_403_1803_0,
    i_8_403_1857_0, i_8_403_1903_0, i_8_403_1941_0, i_8_403_1950_0,
    i_8_403_1962_0, i_8_403_1968_0, i_8_403_1969_0, i_8_403_2004_0,
    i_8_403_2100_0, i_8_403_2104_0, i_8_403_2143_0, i_8_403_2158_0,
    i_8_403_2172_0, i_8_403_2174_0, i_8_403_2175_0, i_8_403_2176_0,
    i_8_403_2177_0, i_8_403_2209_0, i_8_403_2233_0, i_8_403_2245_0,
    i_8_403_2262_0, i_8_403_2263_0, i_8_403_2265_0, i_8_403_2271_0;
  output o_8_403_0_0;
  assign o_8_403_0_0 = ~((~i_8_403_467_0 & ((~i_8_403_313_0 & i_8_403_526_0 & ~i_8_403_844_0 & ~i_8_403_922_0 & ~i_8_403_1428_0 & ~i_8_403_1447_0 & ~i_8_403_1733_0 & ~i_8_403_1748_0 & ~i_8_403_2143_0 & ~i_8_403_2263_0) | (~i_8_403_143_0 & ~i_8_403_403_0 & i_8_403_619_0 & ~i_8_403_840_0 & ~i_8_403_931_0 & ~i_8_403_978_0 & ~i_8_403_980_0 & ~i_8_403_1429_0 & ~i_8_403_1857_0 & ~i_8_403_1950_0 & ~i_8_403_2004_0 & ~i_8_403_2158_0 & ~i_8_403_2265_0 & ~i_8_403_2271_0))) | (i_8_403_526_0 & ((~i_8_403_619_0 & ~i_8_403_1428_0 & ~i_8_403_1632_0 & i_8_403_1671_0 & ~i_8_403_1857_0) | (~i_8_403_287_0 & ~i_8_403_403_0 & ~i_8_403_930_0 & ~i_8_403_980_0 & ~i_8_403_1074_0 & ~i_8_403_1671_0 & ~i_8_403_1725_0 & ~i_8_403_1744_0 & ~i_8_403_1941_0 & ~i_8_403_2176_0 & ~i_8_403_2233_0 & ~i_8_403_2245_0))) | (~i_8_403_403_0 & ((~i_8_403_39_0 & ~i_8_403_269_0 & ~i_8_403_551_0 & ~i_8_403_582_0 & ~i_8_403_931_0 & ~i_8_403_1725_0 & i_8_403_2177_0) | (~i_8_403_67_0 & ~i_8_403_286_0 & ~i_8_403_823_0 & ~i_8_403_898_0 & ~i_8_403_924_0 & ~i_8_403_978_0 & ~i_8_403_1447_0 & ~i_8_403_1671_0 & ~i_8_403_1941_0 & i_8_403_2100_0 & ~i_8_403_2209_0))) | (~i_8_403_402_0 & ((~i_8_403_269_0 & ((~i_8_403_267_0 & ~i_8_403_619_0 & i_8_403_1030_0 & ~i_8_403_1624_0 & ~i_8_403_1671_0 & ~i_8_403_1903_0 & ~i_8_403_2143_0) | (~i_8_403_39_0 & ~i_8_403_287_0 & ~i_8_403_844_0 & ~i_8_403_883_0 & ~i_8_403_922_0 & ~i_8_403_1428_0 & ~i_8_403_1446_0 & i_8_403_2104_0 & ~i_8_403_2209_0))) | (~i_8_403_980_0 & ((i_8_403_219_0 & ((~i_8_403_67_0 & ~i_8_403_313_0 & ~i_8_403_933_0 & ~i_8_403_964_0 & ~i_8_403_978_0 & ~i_8_403_1307_0 & ~i_8_403_1428_0 & ~i_8_403_1447_0) | (~i_8_403_286_0 & ~i_8_403_583_0 & ~i_8_403_726_0 & ~i_8_403_843_0 & ~i_8_403_931_0 & ~i_8_403_1774_0 & ~i_8_403_2174_0 & ~i_8_403_2209_0 & ~i_8_403_2265_0))) | (~i_8_403_51_0 & ~i_8_403_286_0 & ~i_8_403_582_0 & ~i_8_403_897_0 & ~i_8_403_930_0 & ~i_8_403_1446_0 & i_8_403_2175_0 & ~i_8_403_2177_0 & ~i_8_403_2209_0 & ~i_8_403_2265_0))) | (~i_8_403_665_0 & ~i_8_403_1428_0 & ((~i_8_403_931_0 & ((i_8_403_219_0 & ~i_8_403_1429_0 & ~i_8_403_1455_0 & ~i_8_403_1733_0 & ~i_8_403_1941_0) | (~i_8_403_582_0 & ~i_8_403_979_0 & ~i_8_403_1748_0 & i_8_403_2177_0))) | (~i_8_403_287_0 & ~i_8_403_313_0 & ~i_8_403_619_0 & ~i_8_403_840_0 & ~i_8_403_844_0 & ~i_8_403_922_0 & ~i_8_403_1725_0 & ~i_8_403_1941_0))))) | (~i_8_403_1725_0 & ((~i_8_403_267_0 & ((~i_8_403_665_0 & ~i_8_403_1446_0 & ((~i_8_403_67_0 & ~i_8_403_1672_0 & ((~i_8_403_287_0 & ~i_8_403_551_0 & ~i_8_403_583_0 & ~i_8_403_843_0 & ~i_8_403_924_0 & ~i_8_403_931_0 & ~i_8_403_1074_0 & ~i_8_403_1624_0 & ~i_8_403_1671_0 & ~i_8_403_1857_0) | (~i_8_403_313_0 & ~i_8_403_492_0 & ~i_8_403_807_0 & ~i_8_403_897_0 & ~i_8_403_930_0 & ~i_8_403_980_0 & ~i_8_403_1438_0 & ~i_8_403_1733_0 & ~i_8_403_1744_0 & ~i_8_403_1803_0 & ~i_8_403_2143_0))) | (~i_8_403_143_0 & ~i_8_403_287_0 & ~i_8_403_313_0 & ~i_8_403_492_0 & ~i_8_403_619_0 & ~i_8_403_922_0 & ~i_8_403_933_0 & ~i_8_403_980_0 & ~i_8_403_1074_0 & ~i_8_403_1941_0 & ~i_8_403_2158_0))) | (~i_8_403_39_0 & ~i_8_403_898_0 & ~i_8_403_978_0 & ~i_8_403_1671_0 & ~i_8_403_1903_0 & i_8_403_2175_0))) | (~i_8_403_843_0 & i_8_403_844_0 & ~i_8_403_931_0 & ~i_8_403_1733_0 & i_8_403_2233_0) | (~i_8_403_51_0 & ~i_8_403_313_0 & i_8_403_423_0 & ~i_8_403_930_0 & ~i_8_403_1429_0 & ~i_8_403_1672_0 & ~i_8_403_2233_0 & ~i_8_403_2263_0))) | (~i_8_403_39_0 & ~i_8_403_980_0 & ((~i_8_403_143_0 & ~i_8_403_313_0 & ~i_8_403_619_0 & ~i_8_403_924_0 & ~i_8_403_978_0 & ~i_8_403_1733_0 & i_8_403_1968_0) | (~i_8_403_807_0 & ~i_8_403_898_0 & ~i_8_403_1671_0 & i_8_403_1748_0 & ~i_8_403_2004_0))) | (~i_8_403_978_0 & ((~i_8_403_51_0 & ~i_8_403_1447_0 & ((~i_8_403_143_0 & ~i_8_403_582_0 & ~i_8_403_898_0 & ~i_8_403_1446_0 & ~i_8_403_1773_0 & ~i_8_403_1857_0 & ~i_8_403_1941_0 & i_8_403_1969_0 & ~i_8_403_2100_0) | (~i_8_403_619_0 & i_8_403_823_0 & ~i_8_403_922_0 & ~i_8_403_1276_0 & ~i_8_403_1534_0 & ~i_8_403_1968_0 & ~i_8_403_2174_0 & ~i_8_403_2209_0))) | (~i_8_403_313_0 & ~i_8_403_492_0 & ~i_8_403_583_0 & i_8_403_654_0 & ~i_8_403_876_0 & ~i_8_403_1969_0) | (~i_8_403_219_0 & ~i_8_403_269_0 & ~i_8_403_1429_0 & ~i_8_403_2004_0 & i_8_403_2176_0 & ~i_8_403_2263_0))) | (~i_8_403_143_0 & ((~i_8_403_843_0 & ~i_8_403_922_0 & i_8_403_1535_0) | (~i_8_403_287_0 & ~i_8_403_619_0 & i_8_403_665_0 & ~i_8_403_840_0 & ~i_8_403_844_0 & ~i_8_403_979_0 & ~i_8_403_1857_0 & ~i_8_403_2104_0))) | (~i_8_403_582_0 & ((~i_8_403_66_0 & ~i_8_403_551_0 & ~i_8_403_665_0 & ~i_8_403_807_0 & ~i_8_403_823_0 & i_8_403_840_0 & ~i_8_403_924_0 & ~i_8_403_931_0 & ~i_8_403_1428_0 & ~i_8_403_1438_0 & ~i_8_403_1632_0 & ~i_8_403_1671_0) | (~i_8_403_898_0 & ~i_8_403_1624_0 & i_8_403_1773_0 & ~i_8_403_2209_0))) | (i_8_403_883_0 & ~i_8_403_898_0 & ~i_8_403_922_0 & ~i_8_403_930_0 & ~i_8_403_933_0) | (~i_8_403_840_0 & ~i_8_403_1438_0 & i_8_403_1969_0 & i_8_403_2143_0) | (i_8_403_66_0 & ~i_8_403_844_0 & i_8_403_1774_0 & ~i_8_403_2143_0) | (~i_8_403_287_0 & ~i_8_403_843_0 & ~i_8_403_979_0 & ~i_8_403_1857_0 & ~i_8_403_1903_0 & ~i_8_403_2104_0 & i_8_403_2174_0) | (i_8_403_195_0 & ~i_8_403_583_0 & ~i_8_403_897_0 & ~i_8_403_1733_0 & i_8_403_1803_0 & ~i_8_403_2262_0));
endmodule



// Benchmark "kernel_8_404" written by ABC on Sun Jul 19 10:10:08 2020

module kernel_8_404 ( 
    i_8_404_25_0, i_8_404_31_0, i_8_404_35_0, i_8_404_86_0, i_8_404_160_0,
    i_8_404_188_0, i_8_404_205_0, i_8_404_295_0, i_8_404_296_0,
    i_8_404_332_0, i_8_404_377_0, i_8_404_457_0, i_8_404_463_0,
    i_8_404_483_0, i_8_404_484_0, i_8_404_502_0, i_8_404_508_0,
    i_8_404_528_0, i_8_404_529_0, i_8_404_539_0, i_8_404_553_0,
    i_8_404_556_0, i_8_404_626_0, i_8_404_629_0, i_8_404_636_0,
    i_8_404_664_0, i_8_404_692_0, i_8_404_716_0, i_8_404_718_0,
    i_8_404_719_0, i_8_404_727_0, i_8_404_735_0, i_8_404_760_0,
    i_8_404_762_0, i_8_404_769_0, i_8_404_772_0, i_8_404_870_0,
    i_8_404_871_0, i_8_404_880_0, i_8_404_897_0, i_8_404_926_0,
    i_8_404_951_0, i_8_404_978_0, i_8_404_988_0, i_8_404_989_0,
    i_8_404_993_0, i_8_404_994_0, i_8_404_995_0, i_8_404_1032_0,
    i_8_404_1033_0, i_8_404_1034_0, i_8_404_1093_0, i_8_404_1113_0,
    i_8_404_1114_0, i_8_404_1203_0, i_8_404_1230_0, i_8_404_1239_0,
    i_8_404_1293_0, i_8_404_1330_0, i_8_404_1347_0, i_8_404_1407_0,
    i_8_404_1452_0, i_8_404_1482_0, i_8_404_1484_0, i_8_404_1509_0,
    i_8_404_1528_0, i_8_404_1529_0, i_8_404_1601_0, i_8_404_1618_0,
    i_8_404_1680_0, i_8_404_1705_0, i_8_404_1708_0, i_8_404_1716_0,
    i_8_404_1717_0, i_8_404_1718_0, i_8_404_1730_0, i_8_404_1735_0,
    i_8_404_1743_0, i_8_404_1762_0, i_8_404_1778_0, i_8_404_1784_0,
    i_8_404_1798_0, i_8_404_1808_0, i_8_404_1822_0, i_8_404_1905_0,
    i_8_404_1920_0, i_8_404_1929_0, i_8_404_1933_0, i_8_404_1969_0,
    i_8_404_1985_0, i_8_404_2013_0, i_8_404_2015_0, i_8_404_2029_0,
    i_8_404_2113_0, i_8_404_2140_0, i_8_404_2145_0, i_8_404_2146_0,
    i_8_404_2191_0, i_8_404_2230_0, i_8_404_2272_0,
    o_8_404_0_0  );
  input  i_8_404_25_0, i_8_404_31_0, i_8_404_35_0, i_8_404_86_0,
    i_8_404_160_0, i_8_404_188_0, i_8_404_205_0, i_8_404_295_0,
    i_8_404_296_0, i_8_404_332_0, i_8_404_377_0, i_8_404_457_0,
    i_8_404_463_0, i_8_404_483_0, i_8_404_484_0, i_8_404_502_0,
    i_8_404_508_0, i_8_404_528_0, i_8_404_529_0, i_8_404_539_0,
    i_8_404_553_0, i_8_404_556_0, i_8_404_626_0, i_8_404_629_0,
    i_8_404_636_0, i_8_404_664_0, i_8_404_692_0, i_8_404_716_0,
    i_8_404_718_0, i_8_404_719_0, i_8_404_727_0, i_8_404_735_0,
    i_8_404_760_0, i_8_404_762_0, i_8_404_769_0, i_8_404_772_0,
    i_8_404_870_0, i_8_404_871_0, i_8_404_880_0, i_8_404_897_0,
    i_8_404_926_0, i_8_404_951_0, i_8_404_978_0, i_8_404_988_0,
    i_8_404_989_0, i_8_404_993_0, i_8_404_994_0, i_8_404_995_0,
    i_8_404_1032_0, i_8_404_1033_0, i_8_404_1034_0, i_8_404_1093_0,
    i_8_404_1113_0, i_8_404_1114_0, i_8_404_1203_0, i_8_404_1230_0,
    i_8_404_1239_0, i_8_404_1293_0, i_8_404_1330_0, i_8_404_1347_0,
    i_8_404_1407_0, i_8_404_1452_0, i_8_404_1482_0, i_8_404_1484_0,
    i_8_404_1509_0, i_8_404_1528_0, i_8_404_1529_0, i_8_404_1601_0,
    i_8_404_1618_0, i_8_404_1680_0, i_8_404_1705_0, i_8_404_1708_0,
    i_8_404_1716_0, i_8_404_1717_0, i_8_404_1718_0, i_8_404_1730_0,
    i_8_404_1735_0, i_8_404_1743_0, i_8_404_1762_0, i_8_404_1778_0,
    i_8_404_1784_0, i_8_404_1798_0, i_8_404_1808_0, i_8_404_1822_0,
    i_8_404_1905_0, i_8_404_1920_0, i_8_404_1929_0, i_8_404_1933_0,
    i_8_404_1969_0, i_8_404_1985_0, i_8_404_2013_0, i_8_404_2015_0,
    i_8_404_2029_0, i_8_404_2113_0, i_8_404_2140_0, i_8_404_2145_0,
    i_8_404_2146_0, i_8_404_2191_0, i_8_404_2230_0, i_8_404_2272_0;
  output o_8_404_0_0;
  assign o_8_404_0_0 = 0;
endmodule



// Benchmark "kernel_8_405" written by ABC on Sun Jul 19 10:10:09 2020

module kernel_8_405 ( 
    i_8_405_1_0, i_8_405_2_0, i_8_405_82_0, i_8_405_83_0, i_8_405_95_0,
    i_8_405_101_0, i_8_405_104_0, i_8_405_154_0, i_8_405_221_0,
    i_8_405_244_0, i_8_405_281_0, i_8_405_289_0, i_8_405_290_0,
    i_8_405_292_0, i_8_405_293_0, i_8_405_326_0, i_8_405_342_0,
    i_8_405_343_0, i_8_405_363_0, i_8_405_382_0, i_8_405_401_0,
    i_8_405_419_0, i_8_405_434_0, i_8_405_437_0, i_8_405_440_0,
    i_8_405_454_0, i_8_405_478_0, i_8_405_479_0, i_8_405_545_0,
    i_8_405_585_0, i_8_405_607_0, i_8_405_608_0, i_8_405_613_0,
    i_8_405_622_0, i_8_405_623_0, i_8_405_625_0, i_8_405_631_0,
    i_8_405_659_0, i_8_405_666_0, i_8_405_667_0, i_8_405_682_0,
    i_8_405_703_0, i_8_405_704_0, i_8_405_713_0, i_8_405_721_0,
    i_8_405_722_0, i_8_405_776_0, i_8_405_784_0, i_8_405_796_0,
    i_8_405_823_0, i_8_405_830_0, i_8_405_832_0, i_8_405_833_0,
    i_8_405_838_0, i_8_405_843_0, i_8_405_868_0, i_8_405_968_0,
    i_8_405_974_0, i_8_405_977_0, i_8_405_1031_0, i_8_405_1040_0,
    i_8_405_1049_0, i_8_405_1112_0, i_8_405_1161_0, i_8_405_1180_0,
    i_8_405_1181_0, i_8_405_1208_0, i_8_405_1238_0, i_8_405_1265_0,
    i_8_405_1298_0, i_8_405_1355_0, i_8_405_1373_0, i_8_405_1388_0,
    i_8_405_1435_0, i_8_405_1547_0, i_8_405_1565_0, i_8_405_1576_0,
    i_8_405_1585_0, i_8_405_1586_0, i_8_405_1679_0, i_8_405_1750_0,
    i_8_405_1783_0, i_8_405_1801_0, i_8_405_1807_0, i_8_405_1855_0,
    i_8_405_1858_0, i_8_405_1876_0, i_8_405_1900_0, i_8_405_1904_0,
    i_8_405_1985_0, i_8_405_1991_0, i_8_405_1992_0, i_8_405_1994_0,
    i_8_405_2036_0, i_8_405_2093_0, i_8_405_2110_0, i_8_405_2143_0,
    i_8_405_2146_0, i_8_405_2182_0, i_8_405_2279_0,
    o_8_405_0_0  );
  input  i_8_405_1_0, i_8_405_2_0, i_8_405_82_0, i_8_405_83_0,
    i_8_405_95_0, i_8_405_101_0, i_8_405_104_0, i_8_405_154_0,
    i_8_405_221_0, i_8_405_244_0, i_8_405_281_0, i_8_405_289_0,
    i_8_405_290_0, i_8_405_292_0, i_8_405_293_0, i_8_405_326_0,
    i_8_405_342_0, i_8_405_343_0, i_8_405_363_0, i_8_405_382_0,
    i_8_405_401_0, i_8_405_419_0, i_8_405_434_0, i_8_405_437_0,
    i_8_405_440_0, i_8_405_454_0, i_8_405_478_0, i_8_405_479_0,
    i_8_405_545_0, i_8_405_585_0, i_8_405_607_0, i_8_405_608_0,
    i_8_405_613_0, i_8_405_622_0, i_8_405_623_0, i_8_405_625_0,
    i_8_405_631_0, i_8_405_659_0, i_8_405_666_0, i_8_405_667_0,
    i_8_405_682_0, i_8_405_703_0, i_8_405_704_0, i_8_405_713_0,
    i_8_405_721_0, i_8_405_722_0, i_8_405_776_0, i_8_405_784_0,
    i_8_405_796_0, i_8_405_823_0, i_8_405_830_0, i_8_405_832_0,
    i_8_405_833_0, i_8_405_838_0, i_8_405_843_0, i_8_405_868_0,
    i_8_405_968_0, i_8_405_974_0, i_8_405_977_0, i_8_405_1031_0,
    i_8_405_1040_0, i_8_405_1049_0, i_8_405_1112_0, i_8_405_1161_0,
    i_8_405_1180_0, i_8_405_1181_0, i_8_405_1208_0, i_8_405_1238_0,
    i_8_405_1265_0, i_8_405_1298_0, i_8_405_1355_0, i_8_405_1373_0,
    i_8_405_1388_0, i_8_405_1435_0, i_8_405_1547_0, i_8_405_1565_0,
    i_8_405_1576_0, i_8_405_1585_0, i_8_405_1586_0, i_8_405_1679_0,
    i_8_405_1750_0, i_8_405_1783_0, i_8_405_1801_0, i_8_405_1807_0,
    i_8_405_1855_0, i_8_405_1858_0, i_8_405_1876_0, i_8_405_1900_0,
    i_8_405_1904_0, i_8_405_1985_0, i_8_405_1991_0, i_8_405_1992_0,
    i_8_405_1994_0, i_8_405_2036_0, i_8_405_2093_0, i_8_405_2110_0,
    i_8_405_2143_0, i_8_405_2146_0, i_8_405_2182_0, i_8_405_2279_0;
  output o_8_405_0_0;
  assign o_8_405_0_0 = ~((~i_8_405_2_0 & ((~i_8_405_83_0 & ~i_8_405_437_0 & ~i_8_405_703_0 & ~i_8_405_713_0 & ~i_8_405_722_0 & ~i_8_405_868_0) | (~i_8_405_101_0 & ~i_8_405_154_0 & ~i_8_405_281_0 & ~i_8_405_292_0 & ~i_8_405_667_0 & ~i_8_405_776_0 & ~i_8_405_1161_0 & ~i_8_405_1180_0 & ~i_8_405_1181_0 & ~i_8_405_1238_0 & ~i_8_405_1435_0))) | (~i_8_405_104_0 & ((~i_8_405_1_0 & ~i_8_405_244_0 & ~i_8_405_326_0 & ~i_8_405_623_0 & ~i_8_405_784_0 & i_8_405_830_0 & ~i_8_405_974_0 & ~i_8_405_1565_0 & ~i_8_405_1807_0) | (~i_8_405_667_0 & ~i_8_405_721_0 & ~i_8_405_830_0 & i_8_405_1750_0 & ~i_8_405_2182_0))) | (~i_8_405_1_0 & ((i_8_405_703_0 & ~i_8_405_713_0 & ~i_8_405_833_0 & ~i_8_405_1876_0 & ~i_8_405_1900_0) | (~i_8_405_83_0 & ~i_8_405_281_0 & ~i_8_405_622_0 & ~i_8_405_784_0 & ~i_8_405_830_0 & ~i_8_405_2279_0))) | (~i_8_405_244_0 & ((i_8_405_289_0 & i_8_405_1031_0) | (~i_8_405_281_0 & ~i_8_405_401_0 & ~i_8_405_721_0 & ~i_8_405_1388_0 & ~i_8_405_1855_0 & ~i_8_405_1876_0 & i_8_405_1991_0))) | (~i_8_405_631_0 & ((~i_8_405_95_0 & ~i_8_405_221_0 & ~i_8_405_419_0 & ~i_8_405_722_0 & ~i_8_405_843_0 & ~i_8_405_968_0 & ~i_8_405_974_0 & ~i_8_405_1181_0) | (~i_8_405_281_0 & ~i_8_405_823_0 & i_8_405_968_0 & i_8_405_1238_0))) | (~i_8_405_290_0 & ((~i_8_405_281_0 & ((~i_8_405_342_0 & ~i_8_405_608_0 & ~i_8_405_622_0 & i_8_405_1238_0 & ~i_8_405_1855_0 & ~i_8_405_1904_0 & i_8_405_1994_0 & i_8_405_2093_0) | (~i_8_405_292_0 & ~i_8_405_437_0 & ~i_8_405_666_0 & ~i_8_405_721_0 & ~i_8_405_784_0 & ~i_8_405_832_0 & ~i_8_405_1181_0 & ~i_8_405_1298_0 & ~i_8_405_1783_0 & ~i_8_405_2143_0))) | (~i_8_405_667_0 & ((~i_8_405_833_0 & i_8_405_838_0 & ~i_8_405_1112_0 & ~i_8_405_1750_0) | (~i_8_405_382_0 & ~i_8_405_585_0 & ~i_8_405_830_0 & ~i_8_405_1040_0 & ~i_8_405_1180_0 & ~i_8_405_1586_0 & i_8_405_1679_0 & ~i_8_405_2146_0))) | (~i_8_405_434_0 & ~i_8_405_666_0 & ~i_8_405_830_0 & ~i_8_405_974_0 & ~i_8_405_1355_0 & ~i_8_405_1750_0) | (~i_8_405_293_0 & ~i_8_405_722_0 & ~i_8_405_776_0 & i_8_405_1783_0 & ~i_8_405_1855_0 & i_8_405_2143_0))) | (~i_8_405_434_0 & ((i_8_405_221_0 & ~i_8_405_722_0 & i_8_405_838_0 & i_8_405_1994_0) | (~i_8_405_363_0 & ~i_8_405_968_0 & ~i_8_405_1112_0 & ~i_8_405_1388_0 & ~i_8_405_1855_0 & ~i_8_405_2110_0))) | (~i_8_405_722_0 & ((~i_8_405_101_0 & ~i_8_405_721_0 & ~i_8_405_968_0 & ~i_8_405_1388_0 & i_8_405_1679_0 & ~i_8_405_1991_0) | (~i_8_405_326_0 & i_8_405_607_0 & ~i_8_405_843_0 & ~i_8_405_1049_0 & ~i_8_405_1876_0 & ~i_8_405_2110_0 & ~i_8_405_2279_0))) | (~i_8_405_721_0 & ~i_8_405_1904_0 & ((~i_8_405_343_0 & ~i_8_405_776_0 & ~i_8_405_968_0 & i_8_405_1858_0 & ~i_8_405_1994_0) | (~i_8_405_289_0 & ~i_8_405_830_0 & ~i_8_405_1388_0 & i_8_405_1435_0 & ~i_8_405_1679_0 & ~i_8_405_2093_0))) | (~i_8_405_713_0 & i_8_405_1904_0) | (i_8_405_977_0 & ~i_8_405_1181_0 & ~i_8_405_2036_0 & ~i_8_405_2182_0));
endmodule



// Benchmark "kernel_8_406" written by ABC on Sun Jul 19 10:10:11 2020

module kernel_8_406 ( 
    i_8_406_3_0, i_8_406_23_0, i_8_406_51_0, i_8_406_52_0, i_8_406_58_0,
    i_8_406_68_0, i_8_406_97_0, i_8_406_98_0, i_8_406_140_0, i_8_406_142_0,
    i_8_406_160_0, i_8_406_219_0, i_8_406_241_0, i_8_406_247_0,
    i_8_406_304_0, i_8_406_311_0, i_8_406_328_0, i_8_406_329_0,
    i_8_406_346_0, i_8_406_347_0, i_8_406_388_0, i_8_406_437_0,
    i_8_406_440_0, i_8_406_507_0, i_8_406_528_0, i_8_406_555_0,
    i_8_406_580_0, i_8_406_599_0, i_8_406_600_0, i_8_406_606_0,
    i_8_406_608_0, i_8_406_610_0, i_8_406_634_0, i_8_406_642_0,
    i_8_406_655_0, i_8_406_705_0, i_8_406_706_0, i_8_406_709_0,
    i_8_406_716_0, i_8_406_723_0, i_8_406_724_0, i_8_406_760_0,
    i_8_406_813_0, i_8_406_814_0, i_8_406_815_0, i_8_406_836_0,
    i_8_406_840_0, i_8_406_875_0, i_8_406_970_0, i_8_406_971_0,
    i_8_406_1034_0, i_8_406_1050_0, i_8_406_1051_0, i_8_406_1071_0,
    i_8_406_1114_0, i_8_406_1241_0, i_8_406_1281_0, i_8_406_1292_0,
    i_8_406_1305_0, i_8_406_1306_0, i_8_406_1316_0, i_8_406_1355_0,
    i_8_406_1389_0, i_8_406_1391_0, i_8_406_1407_0, i_8_406_1409_0,
    i_8_406_1410_0, i_8_406_1411_0, i_8_406_1471_0, i_8_406_1507_0,
    i_8_406_1531_0, i_8_406_1570_0, i_8_406_1573_0, i_8_406_1574_0,
    i_8_406_1642_0, i_8_406_1653_0, i_8_406_1664_0, i_8_406_1678_0,
    i_8_406_1679_0, i_8_406_1719_0, i_8_406_1731_0, i_8_406_1760_0,
    i_8_406_1784_0, i_8_406_1820_0, i_8_406_1887_0, i_8_406_1948_0,
    i_8_406_1963_0, i_8_406_1983_0, i_8_406_1997_0, i_8_406_2028_0,
    i_8_406_2031_0, i_8_406_2056_0, i_8_406_2057_0, i_8_406_2109_0,
    i_8_406_2151_0, i_8_406_2154_0, i_8_406_2156_0, i_8_406_2190_0,
    i_8_406_2216_0, i_8_406_2282_0,
    o_8_406_0_0  );
  input  i_8_406_3_0, i_8_406_23_0, i_8_406_51_0, i_8_406_52_0,
    i_8_406_58_0, i_8_406_68_0, i_8_406_97_0, i_8_406_98_0, i_8_406_140_0,
    i_8_406_142_0, i_8_406_160_0, i_8_406_219_0, i_8_406_241_0,
    i_8_406_247_0, i_8_406_304_0, i_8_406_311_0, i_8_406_328_0,
    i_8_406_329_0, i_8_406_346_0, i_8_406_347_0, i_8_406_388_0,
    i_8_406_437_0, i_8_406_440_0, i_8_406_507_0, i_8_406_528_0,
    i_8_406_555_0, i_8_406_580_0, i_8_406_599_0, i_8_406_600_0,
    i_8_406_606_0, i_8_406_608_0, i_8_406_610_0, i_8_406_634_0,
    i_8_406_642_0, i_8_406_655_0, i_8_406_705_0, i_8_406_706_0,
    i_8_406_709_0, i_8_406_716_0, i_8_406_723_0, i_8_406_724_0,
    i_8_406_760_0, i_8_406_813_0, i_8_406_814_0, i_8_406_815_0,
    i_8_406_836_0, i_8_406_840_0, i_8_406_875_0, i_8_406_970_0,
    i_8_406_971_0, i_8_406_1034_0, i_8_406_1050_0, i_8_406_1051_0,
    i_8_406_1071_0, i_8_406_1114_0, i_8_406_1241_0, i_8_406_1281_0,
    i_8_406_1292_0, i_8_406_1305_0, i_8_406_1306_0, i_8_406_1316_0,
    i_8_406_1355_0, i_8_406_1389_0, i_8_406_1391_0, i_8_406_1407_0,
    i_8_406_1409_0, i_8_406_1410_0, i_8_406_1411_0, i_8_406_1471_0,
    i_8_406_1507_0, i_8_406_1531_0, i_8_406_1570_0, i_8_406_1573_0,
    i_8_406_1574_0, i_8_406_1642_0, i_8_406_1653_0, i_8_406_1664_0,
    i_8_406_1678_0, i_8_406_1679_0, i_8_406_1719_0, i_8_406_1731_0,
    i_8_406_1760_0, i_8_406_1784_0, i_8_406_1820_0, i_8_406_1887_0,
    i_8_406_1948_0, i_8_406_1963_0, i_8_406_1983_0, i_8_406_1997_0,
    i_8_406_2028_0, i_8_406_2031_0, i_8_406_2056_0, i_8_406_2057_0,
    i_8_406_2109_0, i_8_406_2151_0, i_8_406_2154_0, i_8_406_2156_0,
    i_8_406_2190_0, i_8_406_2216_0, i_8_406_2282_0;
  output o_8_406_0_0;
  assign o_8_406_0_0 = ~((~i_8_406_329_0 & ((~i_8_406_52_0 & ~i_8_406_437_0 & ~i_8_406_507_0 & ~i_8_406_642_0 & ~i_8_406_723_0 & ~i_8_406_1389_0 & ~i_8_406_1391_0 & ~i_8_406_1573_0 & ~i_8_406_2031_0) | (~i_8_406_97_0 & ~i_8_406_98_0 & ~i_8_406_600_0 & i_8_406_705_0 & ~i_8_406_724_0 & ~i_8_406_1679_0 & ~i_8_406_2190_0))) | (~i_8_406_1573_0 & ((~i_8_406_388_0 & ((~i_8_406_437_0 & ~i_8_406_813_0 & ~i_8_406_815_0 & ~i_8_406_1306_0 & ~i_8_406_1389_0 & ~i_8_406_1391_0 & ~i_8_406_1997_0 & ~i_8_406_2028_0 & ~i_8_406_2031_0) | (~i_8_406_51_0 & ~i_8_406_52_0 & ~i_8_406_97_0 & ~i_8_406_142_0 & ~i_8_406_311_0 & ~i_8_406_971_0 & ~i_8_406_1071_0 & ~i_8_406_1574_0 & ~i_8_406_1719_0 & ~i_8_406_2282_0))) | (~i_8_406_440_0 & i_8_406_608_0 & ~i_8_406_1391_0 & ~i_8_406_1719_0))) | (~i_8_406_724_0 & ((~i_8_406_51_0 & ~i_8_406_1051_0 & ((~i_8_406_437_0 & i_8_406_528_0 & ~i_8_406_716_0 & ~i_8_406_1570_0 & ~i_8_406_1679_0 & ~i_8_406_2190_0 & ~i_8_406_2216_0) | (~i_8_406_58_0 & ~i_8_406_440_0 & ~i_8_406_599_0 & ~i_8_406_608_0 & ~i_8_406_1316_0 & ~i_8_406_1391_0 & ~i_8_406_1411_0 & ~i_8_406_1471_0 & ~i_8_406_1784_0 & ~i_8_406_1963_0 & ~i_8_406_2151_0 & ~i_8_406_2282_0))) | (~i_8_406_52_0 & ~i_8_406_247_0 & ((~i_8_406_440_0 & ~i_8_406_599_0 & ~i_8_406_97_0 & ~i_8_406_98_0 & ~i_8_406_2028_0 & ~i_8_406_2031_0 & ~i_8_406_642_0 & ~i_8_406_1306_0) | (~i_8_406_580_0 & ~i_8_406_655_0 & ~i_8_406_705_0 & ~i_8_406_836_0 & i_8_406_1114_0 & ~i_8_406_1355_0 & ~i_8_406_1389_0 & ~i_8_406_2056_0))) | (~i_8_406_98_0 & ~i_8_406_814_0 & ~i_8_406_1389_0 & ((~i_8_406_140_0 & ~i_8_406_304_0 & ~i_8_406_440_0 & ~i_8_406_600_0 & ~i_8_406_723_0 & ~i_8_406_1391_0 & ~i_8_406_1411_0 & ~i_8_406_1760_0) | (i_8_406_610_0 & ~i_8_406_716_0 & ~i_8_406_2028_0))) | (i_8_406_1292_0 & i_8_406_1409_0 & ~i_8_406_1410_0) | (i_8_406_1114_0 & i_8_406_1281_0 & ~i_8_406_1574_0 & ~i_8_406_2031_0 & ~i_8_406_2156_0))) | (~i_8_406_2028_0 & ((~i_8_406_52_0 & ((~i_8_406_51_0 & ~i_8_406_247_0 & ~i_8_406_437_0 & ~i_8_406_815_0 & i_8_406_1355_0) | (~i_8_406_97_0 & ~i_8_406_440_0 & ~i_8_406_600_0 & ~i_8_406_642_0 & ~i_8_406_814_0 & ~i_8_406_1034_0 & ~i_8_406_1389_0 & ~i_8_406_1574_0 & ~i_8_406_1678_0 & ~i_8_406_1760_0 & ~i_8_406_2154_0 & ~i_8_406_2216_0))) | (~i_8_406_98_0 & ~i_8_406_813_0 & ~i_8_406_970_0 & ~i_8_406_1050_0 & ~i_8_406_1391_0 & ~i_8_406_2031_0 & ~i_8_406_2190_0 & ~i_8_406_2282_0))) | (~i_8_406_51_0 & ((~i_8_406_440_0 & i_8_406_1407_0 & i_8_406_1409_0) | (~i_8_406_247_0 & ~i_8_406_760_0 & ~i_8_406_970_0 & i_8_406_2056_0))) | (~i_8_406_97_0 & ~i_8_406_723_0 & ((~i_8_406_241_0 & ~i_8_406_813_0 & ~i_8_406_971_0 & ~i_8_406_1306_0 & ~i_8_406_1389_0 & i_8_406_1678_0) | (~i_8_406_528_0 & ~i_8_406_642_0 & ~i_8_406_836_0 & ~i_8_406_875_0 & ~i_8_406_1574_0 & i_8_406_1963_0 & ~i_8_406_1997_0))) | (i_8_406_706_0 & ((i_8_406_606_0 & i_8_406_610_0) | (i_8_406_1305_0 & i_8_406_1679_0))) | (~i_8_406_1051_0 & ~i_8_406_1389_0 & ((~i_8_406_1391_0 & i_8_406_1411_0 & ~i_8_406_2151_0) | (~i_8_406_23_0 & ~i_8_406_160_0 & ~i_8_406_247_0 & ~i_8_406_437_0 & ~i_8_406_1241_0 & ~i_8_406_1355_0 & ~i_8_406_1507_0 & ~i_8_406_1731_0 & ~i_8_406_2282_0))) | (~i_8_406_3_0 & ~i_8_406_1292_0 & i_8_406_1410_0 & i_8_406_1411_0 & ~i_8_406_1574_0));
endmodule



// Benchmark "kernel_8_407" written by ABC on Sun Jul 19 10:10:12 2020

module kernel_8_407 ( 
    i_8_407_22_0, i_8_407_34_0, i_8_407_52_0, i_8_407_53_0, i_8_407_58_0,
    i_8_407_69_0, i_8_407_94_0, i_8_407_97_0, i_8_407_103_0, i_8_407_106_0,
    i_8_407_107_0, i_8_407_135_0, i_8_407_214_0, i_8_407_223_0,
    i_8_407_224_0, i_8_407_241_0, i_8_407_255_0, i_8_407_256_0,
    i_8_407_257_0, i_8_407_304_0, i_8_407_429_0, i_8_407_453_0,
    i_8_407_454_0, i_8_407_507_0, i_8_407_527_0, i_8_407_586_0,
    i_8_407_598_0, i_8_407_606_0, i_8_407_607_0, i_8_407_633_0,
    i_8_407_658_0, i_8_407_660_0, i_8_407_661_0, i_8_407_663_0,
    i_8_407_664_0, i_8_407_678_0, i_8_407_679_0, i_8_407_688_0,
    i_8_407_736_0, i_8_407_766_0, i_8_407_782_0, i_8_407_825_0,
    i_8_407_850_0, i_8_407_868_0, i_8_407_871_0, i_8_407_922_0,
    i_8_407_969_0, i_8_407_990_0, i_8_407_1051_0, i_8_407_1060_0,
    i_8_407_1066_0, i_8_407_1071_0, i_8_407_1137_0, i_8_407_1138_0,
    i_8_407_1268_0, i_8_407_1351_0, i_8_407_1431_0, i_8_407_1444_0,
    i_8_407_1453_0, i_8_407_1454_0, i_8_407_1490_0, i_8_407_1533_0,
    i_8_407_1535_0, i_8_407_1549_0, i_8_407_1561_0, i_8_407_1564_0,
    i_8_407_1596_0, i_8_407_1614_0, i_8_407_1618_0, i_8_407_1633_0,
    i_8_407_1713_0, i_8_407_1714_0, i_8_407_1742_0, i_8_407_1750_0,
    i_8_407_1813_0, i_8_407_1839_0, i_8_407_1840_0, i_8_407_1841_0,
    i_8_407_1860_0, i_8_407_1884_0, i_8_407_1887_0, i_8_407_1893_0,
    i_8_407_1894_0, i_8_407_1904_0, i_8_407_1969_0, i_8_407_1987_0,
    i_8_407_2002_0, i_8_407_2005_0, i_8_407_2077_0, i_8_407_2111_0,
    i_8_407_2127_0, i_8_407_2129_0, i_8_407_2131_0, i_8_407_2137_0,
    i_8_407_2200_0, i_8_407_2215_0, i_8_407_2227_0, i_8_407_2236_0,
    i_8_407_2260_0, i_8_407_2263_0,
    o_8_407_0_0  );
  input  i_8_407_22_0, i_8_407_34_0, i_8_407_52_0, i_8_407_53_0,
    i_8_407_58_0, i_8_407_69_0, i_8_407_94_0, i_8_407_97_0, i_8_407_103_0,
    i_8_407_106_0, i_8_407_107_0, i_8_407_135_0, i_8_407_214_0,
    i_8_407_223_0, i_8_407_224_0, i_8_407_241_0, i_8_407_255_0,
    i_8_407_256_0, i_8_407_257_0, i_8_407_304_0, i_8_407_429_0,
    i_8_407_453_0, i_8_407_454_0, i_8_407_507_0, i_8_407_527_0,
    i_8_407_586_0, i_8_407_598_0, i_8_407_606_0, i_8_407_607_0,
    i_8_407_633_0, i_8_407_658_0, i_8_407_660_0, i_8_407_661_0,
    i_8_407_663_0, i_8_407_664_0, i_8_407_678_0, i_8_407_679_0,
    i_8_407_688_0, i_8_407_736_0, i_8_407_766_0, i_8_407_782_0,
    i_8_407_825_0, i_8_407_850_0, i_8_407_868_0, i_8_407_871_0,
    i_8_407_922_0, i_8_407_969_0, i_8_407_990_0, i_8_407_1051_0,
    i_8_407_1060_0, i_8_407_1066_0, i_8_407_1071_0, i_8_407_1137_0,
    i_8_407_1138_0, i_8_407_1268_0, i_8_407_1351_0, i_8_407_1431_0,
    i_8_407_1444_0, i_8_407_1453_0, i_8_407_1454_0, i_8_407_1490_0,
    i_8_407_1533_0, i_8_407_1535_0, i_8_407_1549_0, i_8_407_1561_0,
    i_8_407_1564_0, i_8_407_1596_0, i_8_407_1614_0, i_8_407_1618_0,
    i_8_407_1633_0, i_8_407_1713_0, i_8_407_1714_0, i_8_407_1742_0,
    i_8_407_1750_0, i_8_407_1813_0, i_8_407_1839_0, i_8_407_1840_0,
    i_8_407_1841_0, i_8_407_1860_0, i_8_407_1884_0, i_8_407_1887_0,
    i_8_407_1893_0, i_8_407_1894_0, i_8_407_1904_0, i_8_407_1969_0,
    i_8_407_1987_0, i_8_407_2002_0, i_8_407_2005_0, i_8_407_2077_0,
    i_8_407_2111_0, i_8_407_2127_0, i_8_407_2129_0, i_8_407_2131_0,
    i_8_407_2137_0, i_8_407_2200_0, i_8_407_2215_0, i_8_407_2227_0,
    i_8_407_2236_0, i_8_407_2260_0, i_8_407_2263_0;
  output o_8_407_0_0;
  assign o_8_407_0_0 = ~((~i_8_407_1713_0 & ((~i_8_407_1071_0 & ((~i_8_407_22_0 & ~i_8_407_678_0 & ((~i_8_407_257_0 & ~i_8_407_453_0 & ~i_8_407_664_0 & ~i_8_407_679_0 & ~i_8_407_868_0 & ~i_8_407_1561_0 & ~i_8_407_1614_0 & ~i_8_407_1987_0 & ~i_8_407_2005_0) | (~i_8_407_52_0 & ~i_8_407_58_0 & ~i_8_407_97_0 & ~i_8_407_106_0 & ~i_8_407_107_0 & ~i_8_407_871_0 & ~i_8_407_990_0 & ~i_8_407_2263_0))) | (~i_8_407_53_0 & ~i_8_407_94_0 & ~i_8_407_107_0 & ~i_8_407_214_0 & ~i_8_407_660_0 & ~i_8_407_688_0 & ~i_8_407_782_0 & ~i_8_407_871_0 & ~i_8_407_990_0 & ~i_8_407_1549_0 & ~i_8_407_2263_0))) | (~i_8_407_214_0 & ((~i_8_407_34_0 & ~i_8_407_53_0 & ((~i_8_407_58_0 & ~i_8_407_256_0 & ~i_8_407_453_0 & ~i_8_407_679_0 & ~i_8_407_922_0 & ~i_8_407_1618_0 & ~i_8_407_1904_0 & ~i_8_407_2077_0) | (~i_8_407_97_0 & ~i_8_407_454_0 & ~i_8_407_688_0 & ~i_8_407_782_0 & ~i_8_407_1060_0 & ~i_8_407_1561_0 & ~i_8_407_1614_0 & ~i_8_407_2260_0))) | (~i_8_407_52_0 & ~i_8_407_94_0 & ~i_8_407_135_0 & ~i_8_407_664_0 & ~i_8_407_688_0 & ~i_8_407_1614_0 & ~i_8_407_1618_0 & ~i_8_407_1813_0 & ~i_8_407_2200_0 & ~i_8_407_2260_0 & ~i_8_407_2263_0))) | (~i_8_407_2005_0 & ((~i_8_407_106_0 & ~i_8_407_257_0 & ~i_8_407_1060_0 & ~i_8_407_1351_0 & ~i_8_407_1431_0 & ~i_8_407_1549_0 & ~i_8_407_1742_0 & ~i_8_407_1860_0 & ~i_8_407_2002_0) | (~i_8_407_223_0 & ~i_8_407_255_0 & ~i_8_407_850_0 & ~i_8_407_1137_0 & ~i_8_407_1138_0 & ~i_8_407_1564_0 & ~i_8_407_1633_0 & ~i_8_407_1714_0 & ~i_8_407_1813_0 & ~i_8_407_2227_0 & ~i_8_407_2260_0))))) | (~i_8_407_2263_0 & ((~i_8_407_214_0 & ((~i_8_407_34_0 & ~i_8_407_256_0 & ~i_8_407_850_0 & ((~i_8_407_135_0 & ~i_8_407_660_0 & ~i_8_407_661_0 & ~i_8_407_663_0 & ~i_8_407_679_0 & ~i_8_407_922_0 & ~i_8_407_1564_0 & ~i_8_407_1742_0 & ~i_8_407_1904_0) | (~i_8_407_69_0 & ~i_8_407_255_0 & ~i_8_407_1051_0 & ~i_8_407_1618_0 & ~i_8_407_1714_0 & ~i_8_407_2005_0 & ~i_8_407_2236_0))) | (~i_8_407_527_0 & ~i_8_407_660_0 & ~i_8_407_1071_0 & ~i_8_407_1268_0 & i_8_407_1840_0 & ~i_8_407_2077_0))) | (i_8_407_607_0 & ((~i_8_407_107_0 & i_8_407_224_0 & ~i_8_407_990_0 & ~i_8_407_1618_0 & ~i_8_407_1860_0) | (i_8_407_658_0 & ~i_8_407_782_0 & ~i_8_407_1138_0 & ~i_8_407_1614_0 & ~i_8_407_1904_0))) | (~i_8_407_1714_0 & ~i_8_407_2260_0 & ((~i_8_407_135_0 & ~i_8_407_664_0 & i_8_407_1060_0 & ~i_8_407_1840_0 & i_8_407_1841_0) | (~i_8_407_97_0 & ~i_8_407_663_0 & ~i_8_407_990_0 & ~i_8_407_1904_0 & i_8_407_1969_0 & ~i_8_407_1987_0))))) | (~i_8_407_214_0 & ((~i_8_407_34_0 & ~i_8_407_241_0 & ~i_8_407_2200_0 & ~i_8_407_2236_0 & ((~i_8_407_106_0 & ~i_8_407_224_0 & ~i_8_407_871_0 & ~i_8_407_922_0 & ~i_8_407_1051_0 & ~i_8_407_1887_0 & ~i_8_407_1987_0) | (~i_8_407_453_0 & ~i_8_407_598_0 & ~i_8_407_825_0 & ~i_8_407_850_0 & ~i_8_407_1431_0 & ~i_8_407_1813_0 & ~i_8_407_2215_0))) | (~i_8_407_97_0 & ((~i_8_407_52_0 & ~i_8_407_922_0 & ~i_8_407_2005_0 & ((~i_8_407_256_0 & ~i_8_407_257_0 & ~i_8_407_454_0 & ~i_8_407_598_0 & ~i_8_407_1614_0 & ~i_8_407_1618_0) | (~i_8_407_53_0 & ~i_8_407_106_0 & ~i_8_407_107_0 & ~i_8_407_255_0 & ~i_8_407_1714_0 & ~i_8_407_1987_0 & ~i_8_407_2131_0))) | (~i_8_407_58_0 & ~i_8_407_106_0 & ~i_8_407_107_0 & ~i_8_407_969_0 & ~i_8_407_1051_0 & ~i_8_407_1453_0 & ~i_8_407_1750_0 & ~i_8_407_2002_0))) | (~i_8_407_106_0 & ~i_8_407_223_0 & i_8_407_664_0 & ~i_8_407_825_0 & ~i_8_407_1561_0 & ~i_8_407_1614_0 & ~i_8_407_2077_0 & ~i_8_407_2215_0))) | (~i_8_407_58_0 & ((~i_8_407_94_0 & ~i_8_407_106_0 & ~i_8_407_586_0 & ~i_8_407_678_0 & i_8_407_1071_0 & ~i_8_407_1614_0 & ~i_8_407_1813_0) | (~i_8_407_454_0 & ~i_8_407_1071_0 & ~i_8_407_1564_0 & i_8_407_1887_0))) | (~i_8_407_94_0 & ((~i_8_407_97_0 & ~i_8_407_106_0 & ~i_8_407_255_0 & ~i_8_407_257_0 & ~i_8_407_453_0 & ~i_8_407_850_0 & ~i_8_407_1051_0 & ~i_8_407_1618_0) | (~i_8_407_107_0 & ~i_8_407_679_0 & ~i_8_407_922_0 & ~i_8_407_1714_0 & ~i_8_407_1813_0 & ~i_8_407_2200_0 & i_8_407_2227_0))) | (~i_8_407_922_0 & ~i_8_407_1137_0 & ((~i_8_407_34_0 & ~i_8_407_52_0 & ~i_8_407_850_0 & ~i_8_407_990_0 & ~i_8_407_1614_0 & i_8_407_1750_0 & ~i_8_407_1813_0) | (~i_8_407_453_0 & ~i_8_407_766_0 & i_8_407_1533_0 & ~i_8_407_1893_0 & ~i_8_407_2005_0))) | (~i_8_407_2200_0 & ((~i_8_407_103_0 & i_8_407_850_0 & i_8_407_1268_0 & i_8_407_1490_0 & ~i_8_407_2002_0) | (~i_8_407_1969_0 & ~i_8_407_1987_0 & i_8_407_2002_0 & i_8_407_2005_0 & i_8_407_2131_0))) | (~i_8_407_257_0 & ~i_8_407_454_0 & ~i_8_407_661_0 & i_8_407_1535_0));
endmodule



// Benchmark "kernel_8_408" written by ABC on Sun Jul 19 10:10:13 2020

module kernel_8_408 ( 
    i_8_408_21_0, i_8_408_76_0, i_8_408_84_0, i_8_408_91_0, i_8_408_159_0,
    i_8_408_224_0, i_8_408_325_0, i_8_408_329_0, i_8_408_345_0,
    i_8_408_367_0, i_8_408_381_0, i_8_408_382_0, i_8_408_384_0,
    i_8_408_390_0, i_8_408_391_0, i_8_408_399_0, i_8_408_462_0,
    i_8_408_463_0, i_8_408_478_0, i_8_408_483_0, i_8_408_484_0,
    i_8_408_501_0, i_8_408_525_0, i_8_408_526_0, i_8_408_529_0,
    i_8_408_621_0, i_8_408_669_0, i_8_408_673_0, i_8_408_685_0,
    i_8_408_753_0, i_8_408_759_0, i_8_408_760_0, i_8_408_768_0,
    i_8_408_823_0, i_8_408_827_0, i_8_408_840_0, i_8_408_841_0,
    i_8_408_892_0, i_8_408_992_0, i_8_408_1031_0, i_8_408_1075_0,
    i_8_408_1159_0, i_8_408_1191_0, i_8_408_1204_0, i_8_408_1218_0,
    i_8_408_1249_0, i_8_408_1254_0, i_8_408_1255_0, i_8_408_1272_0,
    i_8_408_1273_0, i_8_408_1274_0, i_8_408_1281_0, i_8_408_1303_0,
    i_8_408_1326_0, i_8_408_1358_0, i_8_408_1401_0, i_8_408_1402_0,
    i_8_408_1470_0, i_8_408_1506_0, i_8_408_1539_0, i_8_408_1542_0,
    i_8_408_1554_0, i_8_408_1587_0, i_8_408_1597_0, i_8_408_1600_0,
    i_8_408_1605_0, i_8_408_1633_0, i_8_408_1647_0, i_8_408_1680_0,
    i_8_408_1720_0, i_8_408_1741_0, i_8_408_1761_0, i_8_408_1762_0,
    i_8_408_1803_0, i_8_408_1807_0, i_8_408_1821_0, i_8_408_1839_0,
    i_8_408_1866_0, i_8_408_1867_0, i_8_408_1875_0, i_8_408_1893_0,
    i_8_408_1899_0, i_8_408_1917_0, i_8_408_1918_0, i_8_408_1921_0,
    i_8_408_1947_0, i_8_408_1950_0, i_8_408_1965_0, i_8_408_1967_0,
    i_8_408_2030_0, i_8_408_2033_0, i_8_408_2049_0, i_8_408_2088_0,
    i_8_408_2110_0, i_8_408_2150_0, i_8_408_2181_0, i_8_408_2190_0,
    i_8_408_2191_0, i_8_408_2215_0, i_8_408_2229_0,
    o_8_408_0_0  );
  input  i_8_408_21_0, i_8_408_76_0, i_8_408_84_0, i_8_408_91_0,
    i_8_408_159_0, i_8_408_224_0, i_8_408_325_0, i_8_408_329_0,
    i_8_408_345_0, i_8_408_367_0, i_8_408_381_0, i_8_408_382_0,
    i_8_408_384_0, i_8_408_390_0, i_8_408_391_0, i_8_408_399_0,
    i_8_408_462_0, i_8_408_463_0, i_8_408_478_0, i_8_408_483_0,
    i_8_408_484_0, i_8_408_501_0, i_8_408_525_0, i_8_408_526_0,
    i_8_408_529_0, i_8_408_621_0, i_8_408_669_0, i_8_408_673_0,
    i_8_408_685_0, i_8_408_753_0, i_8_408_759_0, i_8_408_760_0,
    i_8_408_768_0, i_8_408_823_0, i_8_408_827_0, i_8_408_840_0,
    i_8_408_841_0, i_8_408_892_0, i_8_408_992_0, i_8_408_1031_0,
    i_8_408_1075_0, i_8_408_1159_0, i_8_408_1191_0, i_8_408_1204_0,
    i_8_408_1218_0, i_8_408_1249_0, i_8_408_1254_0, i_8_408_1255_0,
    i_8_408_1272_0, i_8_408_1273_0, i_8_408_1274_0, i_8_408_1281_0,
    i_8_408_1303_0, i_8_408_1326_0, i_8_408_1358_0, i_8_408_1401_0,
    i_8_408_1402_0, i_8_408_1470_0, i_8_408_1506_0, i_8_408_1539_0,
    i_8_408_1542_0, i_8_408_1554_0, i_8_408_1587_0, i_8_408_1597_0,
    i_8_408_1600_0, i_8_408_1605_0, i_8_408_1633_0, i_8_408_1647_0,
    i_8_408_1680_0, i_8_408_1720_0, i_8_408_1741_0, i_8_408_1761_0,
    i_8_408_1762_0, i_8_408_1803_0, i_8_408_1807_0, i_8_408_1821_0,
    i_8_408_1839_0, i_8_408_1866_0, i_8_408_1867_0, i_8_408_1875_0,
    i_8_408_1893_0, i_8_408_1899_0, i_8_408_1917_0, i_8_408_1918_0,
    i_8_408_1921_0, i_8_408_1947_0, i_8_408_1950_0, i_8_408_1965_0,
    i_8_408_1967_0, i_8_408_2030_0, i_8_408_2033_0, i_8_408_2049_0,
    i_8_408_2088_0, i_8_408_2110_0, i_8_408_2150_0, i_8_408_2181_0,
    i_8_408_2190_0, i_8_408_2191_0, i_8_408_2215_0, i_8_408_2229_0;
  output o_8_408_0_0;
  assign o_8_408_0_0 = 0;
endmodule



// Benchmark "kernel_8_409" written by ABC on Sun Jul 19 10:10:14 2020

module kernel_8_409 ( 
    i_8_409_9_0, i_8_409_12_0, i_8_409_33_0, i_8_409_61_0, i_8_409_63_0,
    i_8_409_72_0, i_8_409_75_0, i_8_409_135_0, i_8_409_180_0,
    i_8_409_181_0, i_8_409_208_0, i_8_409_279_0, i_8_409_318_0,
    i_8_409_397_0, i_8_409_399_0, i_8_409_417_0, i_8_409_426_0,
    i_8_409_427_0, i_8_409_450_0, i_8_409_453_0, i_8_409_495_0,
    i_8_409_504_0, i_8_409_525_0, i_8_409_528_0, i_8_409_535_0,
    i_8_409_570_0, i_8_409_573_0, i_8_409_579_0, i_8_409_585_0,
    i_8_409_589_0, i_8_409_658_0, i_8_409_660_0, i_8_409_661_0,
    i_8_409_662_0, i_8_409_702_0, i_8_409_748_0, i_8_409_751_0,
    i_8_409_777_0, i_8_409_783_0, i_8_409_797_0, i_8_409_822_0,
    i_8_409_829_0, i_8_409_838_0, i_8_409_841_0, i_8_409_858_0,
    i_8_409_865_0, i_8_409_867_0, i_8_409_877_0, i_8_409_973_0,
    i_8_409_1101_0, i_8_409_1107_0, i_8_409_1152_0, i_8_409_1153_0,
    i_8_409_1198_0, i_8_409_1293_0, i_8_409_1294_0, i_8_409_1314_0,
    i_8_409_1326_0, i_8_409_1332_0, i_8_409_1354_0, i_8_409_1355_0,
    i_8_409_1363_0, i_8_409_1395_0, i_8_409_1398_0, i_8_409_1422_0,
    i_8_409_1425_0, i_8_409_1440_0, i_8_409_1467_0, i_8_409_1480_0,
    i_8_409_1515_0, i_8_409_1521_0, i_8_409_1522_0, i_8_409_1539_0,
    i_8_409_1551_0, i_8_409_1611_0, i_8_409_1629_0, i_8_409_1689_0,
    i_8_409_1701_0, i_8_409_1705_0, i_8_409_1746_0, i_8_409_1764_0,
    i_8_409_1791_0, i_8_409_1794_0, i_8_409_1803_0, i_8_409_1818_0,
    i_8_409_1822_0, i_8_409_1836_0, i_8_409_1837_0, i_8_409_1891_0,
    i_8_409_1956_0, i_8_409_1974_0, i_8_409_1992_0, i_8_409_1996_0,
    i_8_409_2008_0, i_8_409_2052_0, i_8_409_2133_0, i_8_409_2147_0,
    i_8_409_2223_0, i_8_409_2243_0, i_8_409_2273_0,
    o_8_409_0_0  );
  input  i_8_409_9_0, i_8_409_12_0, i_8_409_33_0, i_8_409_61_0,
    i_8_409_63_0, i_8_409_72_0, i_8_409_75_0, i_8_409_135_0, i_8_409_180_0,
    i_8_409_181_0, i_8_409_208_0, i_8_409_279_0, i_8_409_318_0,
    i_8_409_397_0, i_8_409_399_0, i_8_409_417_0, i_8_409_426_0,
    i_8_409_427_0, i_8_409_450_0, i_8_409_453_0, i_8_409_495_0,
    i_8_409_504_0, i_8_409_525_0, i_8_409_528_0, i_8_409_535_0,
    i_8_409_570_0, i_8_409_573_0, i_8_409_579_0, i_8_409_585_0,
    i_8_409_589_0, i_8_409_658_0, i_8_409_660_0, i_8_409_661_0,
    i_8_409_662_0, i_8_409_702_0, i_8_409_748_0, i_8_409_751_0,
    i_8_409_777_0, i_8_409_783_0, i_8_409_797_0, i_8_409_822_0,
    i_8_409_829_0, i_8_409_838_0, i_8_409_841_0, i_8_409_858_0,
    i_8_409_865_0, i_8_409_867_0, i_8_409_877_0, i_8_409_973_0,
    i_8_409_1101_0, i_8_409_1107_0, i_8_409_1152_0, i_8_409_1153_0,
    i_8_409_1198_0, i_8_409_1293_0, i_8_409_1294_0, i_8_409_1314_0,
    i_8_409_1326_0, i_8_409_1332_0, i_8_409_1354_0, i_8_409_1355_0,
    i_8_409_1363_0, i_8_409_1395_0, i_8_409_1398_0, i_8_409_1422_0,
    i_8_409_1425_0, i_8_409_1440_0, i_8_409_1467_0, i_8_409_1480_0,
    i_8_409_1515_0, i_8_409_1521_0, i_8_409_1522_0, i_8_409_1539_0,
    i_8_409_1551_0, i_8_409_1611_0, i_8_409_1629_0, i_8_409_1689_0,
    i_8_409_1701_0, i_8_409_1705_0, i_8_409_1746_0, i_8_409_1764_0,
    i_8_409_1791_0, i_8_409_1794_0, i_8_409_1803_0, i_8_409_1818_0,
    i_8_409_1822_0, i_8_409_1836_0, i_8_409_1837_0, i_8_409_1891_0,
    i_8_409_1956_0, i_8_409_1974_0, i_8_409_1992_0, i_8_409_1996_0,
    i_8_409_2008_0, i_8_409_2052_0, i_8_409_2133_0, i_8_409_2147_0,
    i_8_409_2223_0, i_8_409_2243_0, i_8_409_2273_0;
  output o_8_409_0_0;
  assign o_8_409_0_0 = 0;
endmodule



// Benchmark "kernel_8_410" written by ABC on Sun Jul 19 10:10:15 2020

module kernel_8_410 ( 
    i_8_410_4_0, i_8_410_21_0, i_8_410_24_0, i_8_410_53_0, i_8_410_89_0,
    i_8_410_115_0, i_8_410_175_0, i_8_410_188_0, i_8_410_193_0,
    i_8_410_255_0, i_8_410_256_0, i_8_410_277_0, i_8_410_310_0,
    i_8_410_313_0, i_8_410_336_0, i_8_410_355_0, i_8_410_356_0,
    i_8_410_364_0, i_8_410_463_0, i_8_410_516_0, i_8_410_517_0,
    i_8_410_571_0, i_8_410_580_0, i_8_410_604_0, i_8_410_615_0,
    i_8_410_616_0, i_8_410_617_0, i_8_410_652_0, i_8_410_669_0,
    i_8_410_671_0, i_8_410_678_0, i_8_410_697_0, i_8_410_708_0,
    i_8_410_815_0, i_8_410_831_0, i_8_410_832_0, i_8_410_840_0,
    i_8_410_842_0, i_8_410_846_0, i_8_410_991_0, i_8_410_1057_0,
    i_8_410_1126_0, i_8_410_1131_0, i_8_410_1156_0, i_8_410_1159_0,
    i_8_410_1173_0, i_8_410_1183_0, i_8_410_1201_0, i_8_410_1237_0,
    i_8_410_1273_0, i_8_410_1284_0, i_8_410_1285_0, i_8_410_1305_0,
    i_8_410_1306_0, i_8_410_1336_0, i_8_410_1353_0, i_8_410_1393_0,
    i_8_410_1470_0, i_8_410_1490_0, i_8_410_1498_0, i_8_410_1499_0,
    i_8_410_1525_0, i_8_410_1526_0, i_8_410_1534_0, i_8_410_1597_0,
    i_8_410_1629_0, i_8_410_1653_0, i_8_410_1659_0, i_8_410_1660_0,
    i_8_410_1696_0, i_8_410_1697_0, i_8_410_1724_0, i_8_410_1746_0,
    i_8_410_1771_0, i_8_410_1780_0, i_8_410_1802_0, i_8_410_1806_0,
    i_8_410_1807_0, i_8_410_1808_0, i_8_410_1825_0, i_8_410_1857_0,
    i_8_410_1858_0, i_8_410_1866_0, i_8_410_1876_0, i_8_410_1906_0,
    i_8_410_1919_0, i_8_410_1949_0, i_8_410_1969_0, i_8_410_1974_0,
    i_8_410_2038_0, i_8_410_2047_0, i_8_410_2048_0, i_8_410_2050_0,
    i_8_410_2066_0, i_8_410_2092_0, i_8_410_2108_0, i_8_410_2137_0,
    i_8_410_2147_0, i_8_410_2154_0, i_8_410_2257_0,
    o_8_410_0_0  );
  input  i_8_410_4_0, i_8_410_21_0, i_8_410_24_0, i_8_410_53_0,
    i_8_410_89_0, i_8_410_115_0, i_8_410_175_0, i_8_410_188_0,
    i_8_410_193_0, i_8_410_255_0, i_8_410_256_0, i_8_410_277_0,
    i_8_410_310_0, i_8_410_313_0, i_8_410_336_0, i_8_410_355_0,
    i_8_410_356_0, i_8_410_364_0, i_8_410_463_0, i_8_410_516_0,
    i_8_410_517_0, i_8_410_571_0, i_8_410_580_0, i_8_410_604_0,
    i_8_410_615_0, i_8_410_616_0, i_8_410_617_0, i_8_410_652_0,
    i_8_410_669_0, i_8_410_671_0, i_8_410_678_0, i_8_410_697_0,
    i_8_410_708_0, i_8_410_815_0, i_8_410_831_0, i_8_410_832_0,
    i_8_410_840_0, i_8_410_842_0, i_8_410_846_0, i_8_410_991_0,
    i_8_410_1057_0, i_8_410_1126_0, i_8_410_1131_0, i_8_410_1156_0,
    i_8_410_1159_0, i_8_410_1173_0, i_8_410_1183_0, i_8_410_1201_0,
    i_8_410_1237_0, i_8_410_1273_0, i_8_410_1284_0, i_8_410_1285_0,
    i_8_410_1305_0, i_8_410_1306_0, i_8_410_1336_0, i_8_410_1353_0,
    i_8_410_1393_0, i_8_410_1470_0, i_8_410_1490_0, i_8_410_1498_0,
    i_8_410_1499_0, i_8_410_1525_0, i_8_410_1526_0, i_8_410_1534_0,
    i_8_410_1597_0, i_8_410_1629_0, i_8_410_1653_0, i_8_410_1659_0,
    i_8_410_1660_0, i_8_410_1696_0, i_8_410_1697_0, i_8_410_1724_0,
    i_8_410_1746_0, i_8_410_1771_0, i_8_410_1780_0, i_8_410_1802_0,
    i_8_410_1806_0, i_8_410_1807_0, i_8_410_1808_0, i_8_410_1825_0,
    i_8_410_1857_0, i_8_410_1858_0, i_8_410_1866_0, i_8_410_1876_0,
    i_8_410_1906_0, i_8_410_1919_0, i_8_410_1949_0, i_8_410_1969_0,
    i_8_410_1974_0, i_8_410_2038_0, i_8_410_2047_0, i_8_410_2048_0,
    i_8_410_2050_0, i_8_410_2066_0, i_8_410_2092_0, i_8_410_2108_0,
    i_8_410_2137_0, i_8_410_2147_0, i_8_410_2154_0, i_8_410_2257_0;
  output o_8_410_0_0;
  assign o_8_410_0_0 = ~((~i_8_410_356_0 & ((~i_8_410_175_0 & ~i_8_410_188_0 & i_8_410_336_0 & ~i_8_410_516_0 & ~i_8_410_652_0 & ~i_8_410_1353_0 & ~i_8_410_1597_0 & ~i_8_410_1825_0 & ~i_8_410_1949_0) | (~i_8_410_21_0 & ~i_8_410_89_0 & ~i_8_410_463_0 & ~i_8_410_708_0 & ~i_8_410_1057_0 & ~i_8_410_1393_0 & ~i_8_410_1659_0 & ~i_8_410_1746_0 & ~i_8_410_2050_0))) | (~i_8_410_832_0 & ((~i_8_410_188_0 & ((~i_8_410_24_0 & ~i_8_410_313_0 & ~i_8_410_516_0 & ~i_8_410_517_0 & ~i_8_410_1159_0 & ~i_8_410_1808_0 & ~i_8_410_1866_0 & ~i_8_410_2066_0) | (~i_8_410_256_0 & ~i_8_410_697_0 & ~i_8_410_831_0 & ~i_8_410_1273_0 & ~i_8_410_1353_0 & ~i_8_410_1393_0 & ~i_8_410_1499_0 & ~i_8_410_1876_0 & ~i_8_410_2047_0 & ~i_8_410_2147_0))) | (~i_8_410_89_0 & ~i_8_410_516_0 & ~i_8_410_1131_0 & ~i_8_410_1534_0 & ~i_8_410_1825_0 & ~i_8_410_1876_0 & ~i_8_410_1969_0 & ~i_8_410_2038_0))) | (i_8_410_364_0 & ((~i_8_410_516_0 & ~i_8_410_517_0 & ~i_8_410_831_0 & ~i_8_410_1806_0 & ~i_8_410_1807_0 & ~i_8_410_1949_0) | (i_8_410_193_0 & ~i_8_410_463_0 & ~i_8_410_617_0 & ~i_8_410_846_0 & ~i_8_410_1173_0 & ~i_8_410_1866_0 & ~i_8_410_2038_0))) | (~i_8_410_193_0 & ((~i_8_410_463_0 & ((~i_8_410_21_0 & ~i_8_410_24_0 & ~i_8_410_516_0 & i_8_410_697_0 & ~i_8_410_815_0 & ~i_8_410_1131_0 & ~i_8_410_1526_0) | (~i_8_410_571_0 & ~i_8_410_671_0 & ~i_8_410_1470_0 & ~i_8_410_1653_0 & ~i_8_410_1825_0 & ~i_8_410_1857_0 & ~i_8_410_1969_0 & ~i_8_410_2092_0))) | (~i_8_410_1393_0 & ~i_8_410_2066_0 & ((~i_8_410_1159_0 & ~i_8_410_1499_0 & ~i_8_410_1659_0 & ~i_8_410_1746_0 & ~i_8_410_1780_0 & ~i_8_410_1806_0) | (~i_8_410_89_0 & ~i_8_410_652_0 & i_8_410_1057_0 & ~i_8_410_1597_0 & ~i_8_410_2257_0))) | (~i_8_410_571_0 & i_8_410_840_0 & ~i_8_410_1173_0 & ~i_8_410_1201_0 & ~i_8_410_1490_0 & ~i_8_410_2050_0))) | (~i_8_410_463_0 & ((~i_8_410_89_0 & i_8_410_571_0 & ~i_8_410_1201_0 & i_8_410_1780_0 & ~i_8_410_1866_0 & ~i_8_410_2048_0 & ~i_8_410_2137_0) | (~i_8_410_1131_0 & ~i_8_410_1499_0 & ~i_8_410_1659_0 & ~i_8_410_1660_0 & ~i_8_410_1807_0 & ~i_8_410_2066_0 & ~i_8_410_2257_0))) | (~i_8_410_1597_0 & ((~i_8_410_89_0 & ((i_8_410_842_0 & ~i_8_410_1131_0 & ~i_8_410_1771_0 & i_8_410_1825_0 & ~i_8_410_2137_0) | (~i_8_410_21_0 & ~i_8_410_617_0 & ~i_8_410_1173_0 & ~i_8_410_1806_0 & ~i_8_410_1866_0 & ~i_8_410_2047_0 & ~i_8_410_2257_0))) | (~i_8_410_4_0 & ~i_8_410_355_0 & ~i_8_410_517_0 & ~i_8_410_1653_0 & ~i_8_410_1659_0 & ~i_8_410_1807_0 & ~i_8_410_1808_0 & ~i_8_410_2257_0))) | (~i_8_410_21_0 & ~i_8_410_671_0 & ((~i_8_410_516_0 & ~i_8_410_1393_0 & ~i_8_410_1470_0 & ~i_8_410_1825_0 & ~i_8_410_1949_0 & ~i_8_410_1490_0 & ~i_8_410_1660_0) | (~i_8_410_517_0 & ~i_8_410_1806_0 & ~i_8_410_1906_0 & i_8_410_1969_0 & ~i_8_410_2050_0 & i_8_410_2092_0))) | (~i_8_410_516_0 & ((~i_8_410_1306_0 & ((~i_8_410_24_0 & ~i_8_410_517_0 & ~i_8_410_1393_0 & ~i_8_410_1949_0 & ~i_8_410_2092_0 & i_8_410_2137_0) | (~i_8_410_1499_0 & ~i_8_410_1659_0 & ~i_8_410_1808_0 & ~i_8_410_1969_0 & ~i_8_410_2048_0 & ~i_8_410_2147_0 & ~i_8_410_2257_0))) | (~i_8_410_604_0 & i_8_410_1353_0 & ~i_8_410_1393_0 & ~i_8_410_1534_0 & ~i_8_410_1659_0 & ~i_8_410_1807_0 & ~i_8_410_1866_0))) | (~i_8_410_24_0 & ((~i_8_410_669_0 & ~i_8_410_697_0 & i_8_410_1285_0 & ~i_8_410_1806_0 & ~i_8_410_1949_0 & ~i_8_410_2066_0) | (~i_8_410_277_0 & ~i_8_410_336_0 & ~i_8_410_617_0 & ~i_8_410_1057_0 & ~i_8_410_1173_0 & ~i_8_410_1305_0 & ~i_8_410_1490_0 & ~i_8_410_1653_0 & ~i_8_410_1919_0 & ~i_8_410_2092_0))) | (~i_8_410_1499_0 & ((~i_8_410_1393_0 & ~i_8_410_1498_0 & i_8_410_1724_0 & ~i_8_410_1866_0) | (i_8_410_671_0 & ~i_8_410_815_0 & ~i_8_410_1131_0 & ~i_8_410_1746_0 & ~i_8_410_1876_0 & i_8_410_1919_0))) | (i_8_410_89_0 & i_8_410_1525_0 & ~i_8_410_1857_0 & ~i_8_410_2257_0));
endmodule



// Benchmark "kernel_8_411" written by ABC on Sun Jul 19 10:10:16 2020

module kernel_8_411 ( 
    i_8_411_18_0, i_8_411_96_0, i_8_411_106_0, i_8_411_196_0,
    i_8_411_222_0, i_8_411_225_0, i_8_411_258_0, i_8_411_348_0,
    i_8_411_364_0, i_8_411_365_0, i_8_411_421_0, i_8_411_439_0,
    i_8_411_486_0, i_8_411_610_0, i_8_411_627_0, i_8_411_635_0,
    i_8_411_648_0, i_8_411_651_0, i_8_411_654_0, i_8_411_664_0,
    i_8_411_682_0, i_8_411_693_0, i_8_411_697_0, i_8_411_700_0,
    i_8_411_706_0, i_8_411_708_0, i_8_411_726_0, i_8_411_729_0,
    i_8_411_732_0, i_8_411_733_0, i_8_411_747_0, i_8_411_751_0,
    i_8_411_769_0, i_8_411_777_0, i_8_411_842_0, i_8_411_874_0,
    i_8_411_876_0, i_8_411_877_0, i_8_411_880_0, i_8_411_882_0,
    i_8_411_967_0, i_8_411_969_0, i_8_411_981_0, i_8_411_984_0,
    i_8_411_990_0, i_8_411_996_0, i_8_411_1030_0, i_8_411_1128_0,
    i_8_411_1173_0, i_8_411_1174_0, i_8_411_1224_0, i_8_411_1372_0,
    i_8_411_1410_0, i_8_411_1470_0, i_8_411_1483_0, i_8_411_1527_0,
    i_8_411_1530_0, i_8_411_1533_0, i_8_411_1540_0, i_8_411_1542_0,
    i_8_411_1546_0, i_8_411_1548_0, i_8_411_1555_0, i_8_411_1624_0,
    i_8_411_1642_0, i_8_411_1659_0, i_8_411_1663_0, i_8_411_1683_0,
    i_8_411_1686_0, i_8_411_1691_0, i_8_411_1696_0, i_8_411_1701_0,
    i_8_411_1705_0, i_8_411_1725_0, i_8_411_1734_0, i_8_411_1759_0,
    i_8_411_1767_0, i_8_411_1809_0, i_8_411_1812_0, i_8_411_1824_0,
    i_8_411_1855_0, i_8_411_1885_0, i_8_411_1962_0, i_8_411_1965_0,
    i_8_411_1986_0, i_8_411_1995_0, i_8_411_2007_0, i_8_411_2070_0,
    i_8_411_2083_0, i_8_411_2088_0, i_8_411_2091_0, i_8_411_2104_0,
    i_8_411_2146_0, i_8_411_2223_0, i_8_411_2236_0, i_8_411_2242_0,
    i_8_411_2247_0, i_8_411_2253_0, i_8_411_2254_0, i_8_411_2262_0,
    o_8_411_0_0  );
  input  i_8_411_18_0, i_8_411_96_0, i_8_411_106_0, i_8_411_196_0,
    i_8_411_222_0, i_8_411_225_0, i_8_411_258_0, i_8_411_348_0,
    i_8_411_364_0, i_8_411_365_0, i_8_411_421_0, i_8_411_439_0,
    i_8_411_486_0, i_8_411_610_0, i_8_411_627_0, i_8_411_635_0,
    i_8_411_648_0, i_8_411_651_0, i_8_411_654_0, i_8_411_664_0,
    i_8_411_682_0, i_8_411_693_0, i_8_411_697_0, i_8_411_700_0,
    i_8_411_706_0, i_8_411_708_0, i_8_411_726_0, i_8_411_729_0,
    i_8_411_732_0, i_8_411_733_0, i_8_411_747_0, i_8_411_751_0,
    i_8_411_769_0, i_8_411_777_0, i_8_411_842_0, i_8_411_874_0,
    i_8_411_876_0, i_8_411_877_0, i_8_411_880_0, i_8_411_882_0,
    i_8_411_967_0, i_8_411_969_0, i_8_411_981_0, i_8_411_984_0,
    i_8_411_990_0, i_8_411_996_0, i_8_411_1030_0, i_8_411_1128_0,
    i_8_411_1173_0, i_8_411_1174_0, i_8_411_1224_0, i_8_411_1372_0,
    i_8_411_1410_0, i_8_411_1470_0, i_8_411_1483_0, i_8_411_1527_0,
    i_8_411_1530_0, i_8_411_1533_0, i_8_411_1540_0, i_8_411_1542_0,
    i_8_411_1546_0, i_8_411_1548_0, i_8_411_1555_0, i_8_411_1624_0,
    i_8_411_1642_0, i_8_411_1659_0, i_8_411_1663_0, i_8_411_1683_0,
    i_8_411_1686_0, i_8_411_1691_0, i_8_411_1696_0, i_8_411_1701_0,
    i_8_411_1705_0, i_8_411_1725_0, i_8_411_1734_0, i_8_411_1759_0,
    i_8_411_1767_0, i_8_411_1809_0, i_8_411_1812_0, i_8_411_1824_0,
    i_8_411_1855_0, i_8_411_1885_0, i_8_411_1962_0, i_8_411_1965_0,
    i_8_411_1986_0, i_8_411_1995_0, i_8_411_2007_0, i_8_411_2070_0,
    i_8_411_2083_0, i_8_411_2088_0, i_8_411_2091_0, i_8_411_2104_0,
    i_8_411_2146_0, i_8_411_2223_0, i_8_411_2236_0, i_8_411_2242_0,
    i_8_411_2247_0, i_8_411_2253_0, i_8_411_2254_0, i_8_411_2262_0;
  output o_8_411_0_0;
  assign o_8_411_0_0 = 0;
endmodule



// Benchmark "kernel_8_412" written by ABC on Sun Jul 19 10:10:18 2020

module kernel_8_412 ( 
    i_8_412_59_0, i_8_412_60_0, i_8_412_105_0, i_8_412_107_0,
    i_8_412_108_0, i_8_412_184_0, i_8_412_225_0, i_8_412_226_0,
    i_8_412_228_0, i_8_412_229_0, i_8_412_258_0, i_8_412_285_0,
    i_8_412_337_0, i_8_412_349_0, i_8_412_367_0, i_8_412_393_0,
    i_8_412_484_0, i_8_412_485_0, i_8_412_504_0, i_8_412_505_0,
    i_8_412_526_0, i_8_412_592_0, i_8_412_600_0, i_8_412_602_0,
    i_8_412_630_0, i_8_412_701_0, i_8_412_750_0, i_8_412_780_0,
    i_8_412_850_0, i_8_412_851_0, i_8_412_876_0, i_8_412_879_0,
    i_8_412_882_0, i_8_412_1013_0, i_8_412_1016_0, i_8_412_1032_0,
    i_8_412_1102_0, i_8_412_1138_0, i_8_412_1155_0, i_8_412_1203_0,
    i_8_412_1231_0, i_8_412_1237_0, i_8_412_1238_0, i_8_412_1240_0,
    i_8_412_1241_0, i_8_412_1261_0, i_8_412_1274_0, i_8_412_1311_0,
    i_8_412_1314_0, i_8_412_1315_0, i_8_412_1317_0, i_8_412_1322_0,
    i_8_412_1326_0, i_8_412_1331_0, i_8_412_1353_0, i_8_412_1354_0,
    i_8_412_1361_0, i_8_412_1479_0, i_8_412_1484_0, i_8_412_1490_0,
    i_8_412_1542_0, i_8_412_1548_0, i_8_412_1551_0, i_8_412_1552_0,
    i_8_412_1553_0, i_8_412_1556_0, i_8_412_1653_0, i_8_412_1689_0,
    i_8_412_1691_0, i_8_412_1697_0, i_8_412_1701_0, i_8_412_1708_0,
    i_8_412_1713_0, i_8_412_1715_0, i_8_412_1716_0, i_8_412_1717_0,
    i_8_412_1726_0, i_8_412_1813_0, i_8_412_1814_0, i_8_412_1816_0,
    i_8_412_1825_0, i_8_412_1859_0, i_8_412_1884_0, i_8_412_1885_0,
    i_8_412_1887_0, i_8_412_1888_0, i_8_412_1938_0, i_8_412_1939_0,
    i_8_412_1940_0, i_8_412_1941_0, i_8_412_1980_0, i_8_412_1995_0,
    i_8_412_2053_0, i_8_412_2115_0, i_8_412_2140_0, i_8_412_2169_0,
    i_8_412_2170_0, i_8_412_2287_0, i_8_412_2290_0, i_8_412_2301_0,
    o_8_412_0_0  );
  input  i_8_412_59_0, i_8_412_60_0, i_8_412_105_0, i_8_412_107_0,
    i_8_412_108_0, i_8_412_184_0, i_8_412_225_0, i_8_412_226_0,
    i_8_412_228_0, i_8_412_229_0, i_8_412_258_0, i_8_412_285_0,
    i_8_412_337_0, i_8_412_349_0, i_8_412_367_0, i_8_412_393_0,
    i_8_412_484_0, i_8_412_485_0, i_8_412_504_0, i_8_412_505_0,
    i_8_412_526_0, i_8_412_592_0, i_8_412_600_0, i_8_412_602_0,
    i_8_412_630_0, i_8_412_701_0, i_8_412_750_0, i_8_412_780_0,
    i_8_412_850_0, i_8_412_851_0, i_8_412_876_0, i_8_412_879_0,
    i_8_412_882_0, i_8_412_1013_0, i_8_412_1016_0, i_8_412_1032_0,
    i_8_412_1102_0, i_8_412_1138_0, i_8_412_1155_0, i_8_412_1203_0,
    i_8_412_1231_0, i_8_412_1237_0, i_8_412_1238_0, i_8_412_1240_0,
    i_8_412_1241_0, i_8_412_1261_0, i_8_412_1274_0, i_8_412_1311_0,
    i_8_412_1314_0, i_8_412_1315_0, i_8_412_1317_0, i_8_412_1322_0,
    i_8_412_1326_0, i_8_412_1331_0, i_8_412_1353_0, i_8_412_1354_0,
    i_8_412_1361_0, i_8_412_1479_0, i_8_412_1484_0, i_8_412_1490_0,
    i_8_412_1542_0, i_8_412_1548_0, i_8_412_1551_0, i_8_412_1552_0,
    i_8_412_1553_0, i_8_412_1556_0, i_8_412_1653_0, i_8_412_1689_0,
    i_8_412_1691_0, i_8_412_1697_0, i_8_412_1701_0, i_8_412_1708_0,
    i_8_412_1713_0, i_8_412_1715_0, i_8_412_1716_0, i_8_412_1717_0,
    i_8_412_1726_0, i_8_412_1813_0, i_8_412_1814_0, i_8_412_1816_0,
    i_8_412_1825_0, i_8_412_1859_0, i_8_412_1884_0, i_8_412_1885_0,
    i_8_412_1887_0, i_8_412_1888_0, i_8_412_1938_0, i_8_412_1939_0,
    i_8_412_1940_0, i_8_412_1941_0, i_8_412_1980_0, i_8_412_1995_0,
    i_8_412_2053_0, i_8_412_2115_0, i_8_412_2140_0, i_8_412_2169_0,
    i_8_412_2170_0, i_8_412_2287_0, i_8_412_2290_0, i_8_412_2301_0;
  output o_8_412_0_0;
  assign o_8_412_0_0 = ~((~i_8_412_882_0 & ((~i_8_412_60_0 & ((~i_8_412_105_0 & ~i_8_412_226_0 & i_8_412_349_0 & ~i_8_412_750_0 & i_8_412_1552_0 & ~i_8_412_1814_0) | (~i_8_412_59_0 & i_8_412_1326_0 & i_8_412_1884_0))) | (~i_8_412_105_0 & ((~i_8_412_107_0 & ~i_8_412_2140_0 & ((i_8_412_108_0 & ~i_8_412_393_0 & ~i_8_412_1713_0 & i_8_412_1885_0) | (~i_8_412_876_0 & ~i_8_412_1102_0 & i_8_412_1353_0 & i_8_412_1551_0 & ~i_8_412_1825_0 & ~i_8_412_2115_0 & ~i_8_412_2170_0))) | (~i_8_412_602_0 & ~i_8_412_851_0 & ~i_8_412_1542_0 & i_8_412_1940_0))) | (~i_8_412_226_0 & ((~i_8_412_701_0 & ~i_8_412_850_0 & ~i_8_412_879_0 & ~i_8_412_1032_0 & i_8_412_1315_0) | (~i_8_412_592_0 & ~i_8_412_750_0 & ~i_8_412_780_0 & ~i_8_412_851_0 & i_8_412_1261_0 & ~i_8_412_1995_0 & i_8_412_2053_0 & ~i_8_412_2115_0 & ~i_8_412_2170_0))) | (~i_8_412_630_0 & ((~i_8_412_229_0 & ((i_8_412_337_0 & ~i_8_412_592_0 & ~i_8_412_1354_0 & i_8_412_1548_0) | (i_8_412_1314_0 & ~i_8_412_1713_0))) | (~i_8_412_258_0 & ~i_8_412_780_0 & i_8_412_1311_0 & i_8_412_1353_0 & ~i_8_412_1995_0))) | (~i_8_412_367_0 & ((~i_8_412_258_0 & ~i_8_412_592_0 & ~i_8_412_701_0 & i_8_412_1708_0) | (i_8_412_108_0 & ~i_8_412_850_0 & ~i_8_412_879_0 & ~i_8_412_1311_0 & ~i_8_412_1980_0 & ~i_8_412_2287_0 & ~i_8_412_2290_0))) | (~i_8_412_879_0 & i_8_412_1885_0 & ((~i_8_412_600_0 & ~i_8_412_876_0 & ~i_8_412_1240_0 & ~i_8_412_1354_0) | (~i_8_412_59_0 & ~i_8_412_1274_0 & ~i_8_412_1314_0 & i_8_412_1553_0))) | (~i_8_412_59_0 & ((~i_8_412_850_0 & ~i_8_412_851_0 & ~i_8_412_1813_0 & ~i_8_412_1814_0 & i_8_412_1859_0) | (~i_8_412_1032_0 & ~i_8_412_1825_0 & ~i_8_412_2053_0 & ~i_8_412_2115_0 & i_8_412_2287_0))) | (~i_8_412_393_0 & i_8_412_484_0 & i_8_412_485_0 & i_8_412_526_0 & ~i_8_412_1013_0 & ~i_8_412_1016_0 & ~i_8_412_1361_0 & ~i_8_412_1717_0 & ~i_8_412_1813_0 & ~i_8_412_2290_0))) | (~i_8_412_1980_0 & ((~i_8_412_1138_0 & ((~i_8_412_105_0 & ((~i_8_412_59_0 & ~i_8_412_229_0 & ~i_8_412_349_0 & i_8_412_526_0 & ~i_8_412_602_0 & ~i_8_412_780_0 & ~i_8_412_1238_0 & ~i_8_412_1240_0 & ~i_8_412_1542_0 & ~i_8_412_1653_0 & ~i_8_412_1713_0 & ~i_8_412_1813_0 & ~i_8_412_1885_0 & ~i_8_412_1995_0) | (i_8_412_349_0 & ~i_8_412_393_0 & ~i_8_412_485_0 & ~i_8_412_1231_0 & ~i_8_412_1241_0 & ~i_8_412_1331_0 & ~i_8_412_1717_0 & ~i_8_412_2140_0))) | (~i_8_412_1713_0 & i_8_412_1885_0 & i_8_412_229_0 & i_8_412_1240_0))) | (~i_8_412_600_0 & ((~i_8_412_59_0 & ((~i_8_412_1353_0 & i_8_412_1553_0 & ~i_8_412_1813_0 & i_8_412_1825_0) | (~i_8_412_367_0 & ~i_8_412_850_0 & ~i_8_412_876_0 & ~i_8_412_2287_0 & i_8_412_2290_0))) | (~i_8_412_505_0 & i_8_412_526_0 & ~i_8_412_1240_0 & ~i_8_412_1315_0 & i_8_412_1885_0))) | (~i_8_412_226_0 & ((~i_8_412_1354_0 & i_8_412_1552_0 & i_8_412_1553_0 & ~i_8_412_1556_0 & ~i_8_412_1813_0) | (~i_8_412_349_0 & ~i_8_412_485_0 & i_8_412_1155_0 & ~i_8_412_1353_0 & ~i_8_412_1717_0 & ~i_8_412_1888_0 & ~i_8_412_1940_0 & ~i_8_412_2115_0))) | (~i_8_412_2115_0 & ((~i_8_412_1274_0 & ((~i_8_412_367_0 & i_8_412_1553_0 & i_8_412_1859_0) | (i_8_412_228_0 & i_8_412_229_0 & ~i_8_412_485_0 & ~i_8_412_1032_0 & ~i_8_412_1231_0 & ~i_8_412_1713_0 & ~i_8_412_1884_0))) | (~i_8_412_228_0 & ~i_8_412_630_0 & ~i_8_412_780_0 & ~i_8_412_850_0 & ~i_8_412_1237_0 & ~i_8_412_1240_0 & ~i_8_412_1551_0 & ~i_8_412_1716_0 & ~i_8_412_1859_0 & ~i_8_412_2140_0 & i_8_412_2290_0))) | (~i_8_412_602_0 & ~i_8_412_1016_0 & i_8_412_1274_0 & ~i_8_412_1322_0 & ~i_8_412_1701_0 & ~i_8_412_1813_0 & i_8_412_1859_0))) | (~i_8_412_505_0 & ((~i_8_412_59_0 & ~i_8_412_60_0 & ~i_8_412_105_0 & ~i_8_412_107_0 & ~i_8_412_228_0 & ~i_8_412_337_0 & ~i_8_412_367_0 & ~i_8_412_484_0 & ~i_8_412_504_0 & i_8_412_526_0 & ~i_8_412_600_0 & ~i_8_412_630_0 & ~i_8_412_851_0 & ~i_8_412_1032_0 & ~i_8_412_1653_0 & ~i_8_412_1715_0 & ~i_8_412_1717_0 & ~i_8_412_1885_0) | (~i_8_412_526_0 & i_8_412_1274_0 & i_8_412_1551_0 & ~i_8_412_1816_0 & ~i_8_412_2287_0))) | (~i_8_412_504_0 & ((~i_8_412_60_0 & ~i_8_412_630_0 & i_8_412_1032_0 & ~i_8_412_1261_0 & i_8_412_1653_0) | (i_8_412_505_0 & ~i_8_412_850_0 & i_8_412_1553_0 & ~i_8_412_2053_0))) | (~i_8_412_851_0 & ((~i_8_412_107_0 & ((i_8_412_701_0 & i_8_412_1016_0 & ~i_8_412_1231_0 & ~i_8_412_1552_0) | (~i_8_412_879_0 & ~i_8_412_1102_0 & i_8_412_1322_0 & ~i_8_412_1556_0))) | (~i_8_412_526_0 & ((i_8_412_1238_0 & i_8_412_1552_0 & i_8_412_1556_0) | (~i_8_412_225_0 & i_8_412_505_0 & ~i_8_412_780_0 & ~i_8_412_879_0 & ~i_8_412_1237_0 & ~i_8_412_1274_0 & ~i_8_412_1542_0 & ~i_8_412_1708_0 & ~i_8_412_2169_0 & ~i_8_412_2170_0))) | (~i_8_412_876_0 & ((~i_8_412_1138_0 & i_8_412_1241_0 & i_8_412_1331_0 & ~i_8_412_1717_0) | (~i_8_412_108_0 & ~i_8_412_226_0 & ~i_8_412_600_0 & ~i_8_412_1237_0 & ~i_8_412_1238_0 & i_8_412_1261_0 & ~i_8_412_1888_0 & ~i_8_412_2140_0 & ~i_8_412_2170_0 & ~i_8_412_2287_0))) | (~i_8_412_367_0 & i_8_412_701_0 & ~i_8_412_1315_0 & i_8_412_1552_0 & i_8_412_1556_0) | (~i_8_412_337_0 & ~i_8_412_592_0 & i_8_412_1490_0 & ~i_8_412_1697_0) | (~i_8_412_105_0 & ~i_8_412_228_0 & ~i_8_412_1542_0 & i_8_412_1887_0 & ~i_8_412_2170_0) | (~i_8_412_879_0 & i_8_412_1238_0 & i_8_412_1354_0 & ~i_8_412_1552_0 & ~i_8_412_1814_0 & ~i_8_412_2053_0 & ~i_8_412_2140_0) | (i_8_412_1013_0 & ~i_8_412_1314_0 & i_8_412_1553_0 & ~i_8_412_1995_0 & ~i_8_412_2115_0))) | (~i_8_412_592_0 & ((~i_8_412_59_0 & ((~i_8_412_225_0 & i_8_412_1490_0 & i_8_412_1553_0 & ~i_8_412_1689_0 & ~i_8_412_2053_0) | (~i_8_412_701_0 & ~i_8_412_1353_0 & i_8_412_1354_0 & i_8_412_1556_0 & ~i_8_412_2140_0 & ~i_8_412_2169_0))) | (~i_8_412_107_0 & ((~i_8_412_602_0 & i_8_412_1238_0 & i_8_412_1241_0 & i_8_412_1354_0 & ~i_8_412_1825_0) | (~i_8_412_108_0 & ~i_8_412_1354_0 & i_8_412_1490_0 & ~i_8_412_1995_0 & ~i_8_412_2115_0))) | (i_8_412_226_0 & ~i_8_412_337_0 & ~i_8_412_850_0 & ~i_8_412_1361_0 & ~i_8_412_1552_0 & i_8_412_2053_0 & ~i_8_412_2115_0 & ~i_8_412_2169_0))) | (~i_8_412_850_0 & ((~i_8_412_59_0 & ((~i_8_412_630_0 & i_8_412_1691_0 & ~i_8_412_1814_0 & ~i_8_412_1887_0) | (~i_8_412_225_0 & ~i_8_412_258_0 & ~i_8_412_337_0 & ~i_8_412_526_0 & ~i_8_412_600_0 & ~i_8_412_701_0 & ~i_8_412_876_0 & ~i_8_412_1238_0 & ~i_8_412_1241_0 & ~i_8_412_1311_0 & ~i_8_412_1354_0 & ~i_8_412_1552_0 & ~i_8_412_1553_0 & ~i_8_412_1653_0 & ~i_8_412_1813_0 & ~i_8_412_1816_0 & ~i_8_412_1825_0 & ~i_8_412_1859_0 & ~i_8_412_2115_0 & ~i_8_412_2169_0 & ~i_8_412_2170_0 & ~i_8_412_2290_0))) | (i_8_412_1552_0 & ((~i_8_412_226_0 & ~i_8_412_1813_0 & ((~i_8_412_1138_0 & ~i_8_412_1261_0 & i_8_412_1354_0 & i_8_412_1553_0) | (~i_8_412_105_0 & i_8_412_337_0 & i_8_412_1237_0 & ~i_8_412_2053_0))) | (~i_8_412_225_0 & ~i_8_412_750_0 & ~i_8_412_1155_0 & ~i_8_412_1551_0 & i_8_412_1980_0 & ~i_8_412_1995_0 & ~i_8_412_2170_0))) | (~i_8_412_229_0 & ((~i_8_412_879_0 & ~i_8_412_1231_0 & i_8_412_1726_0 & ~i_8_412_1814_0 & ~i_8_412_1941_0) | (~i_8_412_337_0 & i_8_412_592_0 & ~i_8_412_630_0 & ~i_8_412_780_0 & i_8_412_879_0 & ~i_8_412_1816_0 & ~i_8_412_1825_0 & ~i_8_412_1885_0 & ~i_8_412_1995_0 & ~i_8_412_2169_0 & ~i_8_412_2287_0))) | (i_8_412_526_0 & ((~i_8_412_701_0 & ~i_8_412_879_0 & ~i_8_412_1032_0 & ~i_8_412_1354_0 & ~i_8_412_1479_0 & ~i_8_412_1552_0 & ~i_8_412_1715_0 & ~i_8_412_1884_0 & ~i_8_412_1887_0 & ~i_8_412_1939_0 & ~i_8_412_2169_0) | (~i_8_412_1102_0 & ~i_8_412_1825_0 & ~i_8_412_2115_0 & i_8_412_2290_0))) | (~i_8_412_2170_0 & ((~i_8_412_630_0 & ((~i_8_412_1353_0 & i_8_412_1361_0 & ~i_8_412_1715_0 & ~i_8_412_1717_0) | (~i_8_412_600_0 & i_8_412_750_0 & ~i_8_412_1716_0 & ~i_8_412_1816_0 & i_8_412_1995_0))) | (~i_8_412_285_0 & ~i_8_412_367_0 & ~i_8_412_876_0 & ~i_8_412_1013_0 & i_8_412_1203_0 & ~i_8_412_1314_0 & ~i_8_412_1479_0))) | (~i_8_412_258_0 & ~i_8_412_876_0 & ~i_8_412_1032_0 & ~i_8_412_1887_0 & ~i_8_412_2115_0 & i_8_412_2301_0))) | (~i_8_412_229_0 & ((~i_8_412_367_0 & i_8_412_485_0 & ~i_8_412_602_0 & ~i_8_412_1713_0 & ~i_8_412_1813_0 & ~i_8_412_1814_0) | (~i_8_412_225_0 & i_8_412_505_0 & i_8_412_1490_0 & ~i_8_412_1708_0 & ~i_8_412_1716_0 & ~i_8_412_1816_0 & ~i_8_412_2053_0 & i_8_412_2170_0))) | (i_8_412_1551_0 & ((~i_8_412_225_0 & ((i_8_412_876_0 & ~i_8_412_879_0 & i_8_412_1548_0) | (~i_8_412_600_0 & i_8_412_1261_0 & i_8_412_1552_0 & ~i_8_412_1859_0 & ~i_8_412_2169_0))) | (~i_8_412_876_0 & i_8_412_1653_0 & ~i_8_412_2115_0))) | (~i_8_412_367_0 & ((i_8_412_505_0 & ~i_8_412_876_0 & ~i_8_412_1138_0 & i_8_412_1261_0 & i_8_412_1315_0 & ~i_8_412_1691_0 & ~i_8_412_1715_0) | (~i_8_412_105_0 & ~i_8_412_630_0 & ~i_8_412_1237_0 & i_8_412_1548_0 & ~i_8_412_1825_0 & i_8_412_2287_0))) | (i_8_412_485_0 & ((~i_8_412_60_0 & i_8_412_602_0 & ~i_8_412_1102_0 & ~i_8_412_1556_0 & ~i_8_412_1813_0 & ~i_8_412_1326_0 & ~i_8_412_1552_0) | (~i_8_412_59_0 & ~i_8_412_750_0 & i_8_412_1013_0 & ~i_8_412_1689_0 & ~i_8_412_1887_0 & ~i_8_412_2115_0))) | (~i_8_412_59_0 & ((~i_8_412_1032_0 & ((~i_8_412_60_0 & ((~i_8_412_1013_0 & ~i_8_412_1713_0 & i_8_412_1887_0) | (i_8_412_1238_0 & ~i_8_412_1552_0 & i_8_412_1556_0 & ~i_8_412_1717_0 & ~i_8_412_1816_0 & ~i_8_412_2170_0))) | (~i_8_412_226_0 & ~i_8_412_600_0 & i_8_412_1013_0 & ~i_8_412_1240_0 & ~i_8_412_1717_0 & ~i_8_412_1940_0))) | (~i_8_412_228_0 & i_8_412_504_0 & i_8_412_1314_0 & i_8_412_1548_0) | (i_8_412_258_0 & i_8_412_526_0 & i_8_412_600_0 & ~i_8_412_1138_0 & ~i_8_412_1708_0 & ~i_8_412_1717_0 & ~i_8_412_1816_0 & ~i_8_412_1884_0) | (~i_8_412_105_0 & i_8_412_184_0 & i_8_412_1317_0 & i_8_412_1885_0) | (~i_8_412_184_0 & ~i_8_412_600_0 & ~i_8_412_780_0 & i_8_412_1240_0 & i_8_412_1888_0 & ~i_8_412_2170_0))) | (~i_8_412_105_0 & ((i_8_412_1653_0 & ~i_8_412_1713_0 & i_8_412_1887_0) | (~i_8_412_108_0 & ~i_8_412_228_0 & i_8_412_850_0 & ~i_8_412_1155_0 & ~i_8_412_1331_0 & ~i_8_412_1354_0 & i_8_412_1552_0 & ~i_8_412_1814_0 & ~i_8_412_2170_0))) | (~i_8_412_226_0 & ~i_8_412_2169_0 & ((~i_8_412_780_0 & ~i_8_412_1231_0 & ~i_8_412_1237_0 & i_8_412_1553_0 & i_8_412_1556_0 & ~i_8_412_1715_0) | (~i_8_412_258_0 & ~i_8_412_602_0 & ~i_8_412_750_0 & ~i_8_412_879_0 & ~i_8_412_1032_0 & ~i_8_412_1331_0 & ~i_8_412_1552_0 & ~i_8_412_1556_0 & ~i_8_412_1814_0 & ~i_8_412_1816_0 & i_8_412_2140_0))) | (~i_8_412_228_0 & i_8_412_1552_0 & ((~i_8_412_780_0 & i_8_412_1155_0 & ~i_8_412_1353_0 & ~i_8_412_2053_0) | (~i_8_412_750_0 & i_8_412_882_0 & ~i_8_412_1261_0 & ~i_8_412_2170_0 & i_8_412_2290_0))) | (~i_8_412_750_0 & ((~i_8_412_526_0 & ~i_8_412_780_0 & i_8_412_1553_0 & i_8_412_1701_0) | (~i_8_412_701_0 & ~i_8_412_876_0 & i_8_412_1689_0 & ~i_8_412_1717_0 & i_8_412_2140_0))) | (~i_8_412_349_0 & ~i_8_412_602_0 & ~i_8_412_1231_0 & i_8_412_1484_0 & ~i_8_412_1490_0 & i_8_412_1556_0) | (~i_8_412_60_0 & i_8_412_393_0 & ~i_8_412_1138_0 & ~i_8_412_1237_0 & ~i_8_412_1354_0 & ~i_8_412_1708_0 & ~i_8_412_1716_0 & ~i_8_412_1825_0 & ~i_8_412_1941_0));
endmodule



// Benchmark "kernel_8_413" written by ABC on Sun Jul 19 10:10:19 2020

module kernel_8_413 ( 
    i_8_413_17_0, i_8_413_20_0, i_8_413_41_0, i_8_413_89_0, i_8_413_113_0,
    i_8_413_167_0, i_8_413_197_0, i_8_413_201_0, i_8_413_233_0,
    i_8_413_242_0, i_8_413_248_0, i_8_413_347_0, i_8_413_352_0,
    i_8_413_361_0, i_8_413_362_0, i_8_413_365_0, i_8_413_374_0,
    i_8_413_386_0, i_8_413_427_0, i_8_413_441_0, i_8_413_454_0,
    i_8_413_488_0, i_8_413_524_0, i_8_413_527_0, i_8_413_581_0,
    i_8_413_595_0, i_8_413_609_0, i_8_413_652_0, i_8_413_657_0,
    i_8_413_659_0, i_8_413_676_0, i_8_413_677_0, i_8_413_693_0,
    i_8_413_698_0, i_8_413_703_0, i_8_413_709_0, i_8_413_729_0,
    i_8_413_734_0, i_8_413_761_0, i_8_413_764_0, i_8_413_778_0,
    i_8_413_833_0, i_8_413_835_0, i_8_413_838_0, i_8_413_839_0,
    i_8_413_848_0, i_8_413_850_0, i_8_413_862_0, i_8_413_869_0,
    i_8_413_878_0, i_8_413_881_0, i_8_413_887_0, i_8_413_941_0,
    i_8_413_959_0, i_8_413_1075_0, i_8_413_1076_0, i_8_413_1118_0,
    i_8_413_1136_0, i_8_413_1193_0, i_8_413_1237_0, i_8_413_1262_0,
    i_8_413_1283_0, i_8_413_1325_0, i_8_413_1342_0, i_8_413_1357_0,
    i_8_413_1411_0, i_8_413_1414_0, i_8_413_1474_0, i_8_413_1477_0,
    i_8_413_1478_0, i_8_413_1526_0, i_8_413_1534_0, i_8_413_1543_0,
    i_8_413_1552_0, i_8_413_1589_0, i_8_413_1603_0, i_8_413_1612_0,
    i_8_413_1625_0, i_8_413_1631_0, i_8_413_1697_0, i_8_413_1712_0,
    i_8_413_1736_0, i_8_413_1741_0, i_8_413_1742_0, i_8_413_1863_0,
    i_8_413_1886_0, i_8_413_1889_0, i_8_413_1895_0, i_8_413_1901_0,
    i_8_413_1964_0, i_8_413_1982_0, i_8_413_1985_0, i_8_413_2007_0,
    i_8_413_2011_0, i_8_413_2075_0, i_8_413_2077_0, i_8_413_2134_0,
    i_8_413_2147_0, i_8_413_2150_0, i_8_413_2156_0,
    o_8_413_0_0  );
  input  i_8_413_17_0, i_8_413_20_0, i_8_413_41_0, i_8_413_89_0,
    i_8_413_113_0, i_8_413_167_0, i_8_413_197_0, i_8_413_201_0,
    i_8_413_233_0, i_8_413_242_0, i_8_413_248_0, i_8_413_347_0,
    i_8_413_352_0, i_8_413_361_0, i_8_413_362_0, i_8_413_365_0,
    i_8_413_374_0, i_8_413_386_0, i_8_413_427_0, i_8_413_441_0,
    i_8_413_454_0, i_8_413_488_0, i_8_413_524_0, i_8_413_527_0,
    i_8_413_581_0, i_8_413_595_0, i_8_413_609_0, i_8_413_652_0,
    i_8_413_657_0, i_8_413_659_0, i_8_413_676_0, i_8_413_677_0,
    i_8_413_693_0, i_8_413_698_0, i_8_413_703_0, i_8_413_709_0,
    i_8_413_729_0, i_8_413_734_0, i_8_413_761_0, i_8_413_764_0,
    i_8_413_778_0, i_8_413_833_0, i_8_413_835_0, i_8_413_838_0,
    i_8_413_839_0, i_8_413_848_0, i_8_413_850_0, i_8_413_862_0,
    i_8_413_869_0, i_8_413_878_0, i_8_413_881_0, i_8_413_887_0,
    i_8_413_941_0, i_8_413_959_0, i_8_413_1075_0, i_8_413_1076_0,
    i_8_413_1118_0, i_8_413_1136_0, i_8_413_1193_0, i_8_413_1237_0,
    i_8_413_1262_0, i_8_413_1283_0, i_8_413_1325_0, i_8_413_1342_0,
    i_8_413_1357_0, i_8_413_1411_0, i_8_413_1414_0, i_8_413_1474_0,
    i_8_413_1477_0, i_8_413_1478_0, i_8_413_1526_0, i_8_413_1534_0,
    i_8_413_1543_0, i_8_413_1552_0, i_8_413_1589_0, i_8_413_1603_0,
    i_8_413_1612_0, i_8_413_1625_0, i_8_413_1631_0, i_8_413_1697_0,
    i_8_413_1712_0, i_8_413_1736_0, i_8_413_1741_0, i_8_413_1742_0,
    i_8_413_1863_0, i_8_413_1886_0, i_8_413_1889_0, i_8_413_1895_0,
    i_8_413_1901_0, i_8_413_1964_0, i_8_413_1982_0, i_8_413_1985_0,
    i_8_413_2007_0, i_8_413_2011_0, i_8_413_2075_0, i_8_413_2077_0,
    i_8_413_2134_0, i_8_413_2147_0, i_8_413_2150_0, i_8_413_2156_0;
  output o_8_413_0_0;
  assign o_8_413_0_0 = 0;
endmodule



// Benchmark "kernel_8_414" written by ABC on Sun Jul 19 10:10:19 2020

module kernel_8_414 ( 
    i_8_414_3_0, i_8_414_4_0, i_8_414_27_0, i_8_414_44_0, i_8_414_51_0,
    i_8_414_57_0, i_8_414_75_0, i_8_414_117_0, i_8_414_165_0,
    i_8_414_168_0, i_8_414_192_0, i_8_414_193_0, i_8_414_221_0,
    i_8_414_255_0, i_8_414_265_0, i_8_414_282_0, i_8_414_292_0,
    i_8_414_300_0, i_8_414_337_0, i_8_414_339_0, i_8_414_346_0,
    i_8_414_363_0, i_8_414_364_0, i_8_414_366_0, i_8_414_368_0,
    i_8_414_381_0, i_8_414_382_0, i_8_414_417_0, i_8_414_436_0,
    i_8_414_439_0, i_8_414_455_0, i_8_414_479_0, i_8_414_480_0,
    i_8_414_523_0, i_8_414_525_0, i_8_414_526_0, i_8_414_528_0,
    i_8_414_595_0, i_8_414_615_0, i_8_414_624_0, i_8_414_633_0,
    i_8_414_642_0, i_8_414_661_0, i_8_414_665_0, i_8_414_672_0,
    i_8_414_678_0, i_8_414_694_0, i_8_414_705_0, i_8_414_715_0,
    i_8_414_723_0, i_8_414_759_0, i_8_414_804_0, i_8_414_837_0,
    i_8_414_840_0, i_8_414_841_0, i_8_414_844_0, i_8_414_876_0,
    i_8_414_966_0, i_8_414_969_0, i_8_414_971_0, i_8_414_1072_0,
    i_8_414_1074_0, i_8_414_1182_0, i_8_414_1199_0, i_8_414_1227_0,
    i_8_414_1231_0, i_8_414_1254_0, i_8_414_1263_0, i_8_414_1301_0,
    i_8_414_1305_0, i_8_414_1336_0, i_8_414_1357_0, i_8_414_1551_0,
    i_8_414_1570_0, i_8_414_1574_0, i_8_414_1587_0, i_8_414_1623_0,
    i_8_414_1624_0, i_8_414_1641_0, i_8_414_1644_0, i_8_414_1677_0,
    i_8_414_1717_0, i_8_414_1731_0, i_8_414_1749_0, i_8_414_1807_0,
    i_8_414_1830_0, i_8_414_1857_0, i_8_414_1866_0, i_8_414_1903_0,
    i_8_414_1992_0, i_8_414_1995_0, i_8_414_2028_0, i_8_414_2036_0,
    i_8_414_2056_0, i_8_414_2090_0, i_8_414_2133_0, i_8_414_2190_0,
    i_8_414_2194_0, i_8_414_2293_0, i_8_414_2301_0,
    o_8_414_0_0  );
  input  i_8_414_3_0, i_8_414_4_0, i_8_414_27_0, i_8_414_44_0,
    i_8_414_51_0, i_8_414_57_0, i_8_414_75_0, i_8_414_117_0, i_8_414_165_0,
    i_8_414_168_0, i_8_414_192_0, i_8_414_193_0, i_8_414_221_0,
    i_8_414_255_0, i_8_414_265_0, i_8_414_282_0, i_8_414_292_0,
    i_8_414_300_0, i_8_414_337_0, i_8_414_339_0, i_8_414_346_0,
    i_8_414_363_0, i_8_414_364_0, i_8_414_366_0, i_8_414_368_0,
    i_8_414_381_0, i_8_414_382_0, i_8_414_417_0, i_8_414_436_0,
    i_8_414_439_0, i_8_414_455_0, i_8_414_479_0, i_8_414_480_0,
    i_8_414_523_0, i_8_414_525_0, i_8_414_526_0, i_8_414_528_0,
    i_8_414_595_0, i_8_414_615_0, i_8_414_624_0, i_8_414_633_0,
    i_8_414_642_0, i_8_414_661_0, i_8_414_665_0, i_8_414_672_0,
    i_8_414_678_0, i_8_414_694_0, i_8_414_705_0, i_8_414_715_0,
    i_8_414_723_0, i_8_414_759_0, i_8_414_804_0, i_8_414_837_0,
    i_8_414_840_0, i_8_414_841_0, i_8_414_844_0, i_8_414_876_0,
    i_8_414_966_0, i_8_414_969_0, i_8_414_971_0, i_8_414_1072_0,
    i_8_414_1074_0, i_8_414_1182_0, i_8_414_1199_0, i_8_414_1227_0,
    i_8_414_1231_0, i_8_414_1254_0, i_8_414_1263_0, i_8_414_1301_0,
    i_8_414_1305_0, i_8_414_1336_0, i_8_414_1357_0, i_8_414_1551_0,
    i_8_414_1570_0, i_8_414_1574_0, i_8_414_1587_0, i_8_414_1623_0,
    i_8_414_1624_0, i_8_414_1641_0, i_8_414_1644_0, i_8_414_1677_0,
    i_8_414_1717_0, i_8_414_1731_0, i_8_414_1749_0, i_8_414_1807_0,
    i_8_414_1830_0, i_8_414_1857_0, i_8_414_1866_0, i_8_414_1903_0,
    i_8_414_1992_0, i_8_414_1995_0, i_8_414_2028_0, i_8_414_2036_0,
    i_8_414_2056_0, i_8_414_2090_0, i_8_414_2133_0, i_8_414_2190_0,
    i_8_414_2194_0, i_8_414_2293_0, i_8_414_2301_0;
  output o_8_414_0_0;
  assign o_8_414_0_0 = 0;
endmodule



// Benchmark "kernel_8_415" written by ABC on Sun Jul 19 10:10:20 2020

module kernel_8_415 ( 
    i_8_415_13_0, i_8_415_38_0, i_8_415_40_0, i_8_415_75_0, i_8_415_113_0,
    i_8_415_135_0, i_8_415_193_0, i_8_415_226_0, i_8_415_262_0,
    i_8_415_264_0, i_8_415_308_0, i_8_415_320_0, i_8_415_361_0,
    i_8_415_362_0, i_8_415_422_0, i_8_415_490_0, i_8_415_509_0,
    i_8_415_514_0, i_8_415_520_0, i_8_415_535_0, i_8_415_543_0,
    i_8_415_544_0, i_8_415_580_0, i_8_415_604_0, i_8_415_612_0,
    i_8_415_613_0, i_8_415_634_0, i_8_415_653_0, i_8_415_656_0,
    i_8_415_748_0, i_8_415_751_0, i_8_415_756_0, i_8_415_766_0,
    i_8_415_800_0, i_8_415_802_0, i_8_415_815_0, i_8_415_837_0,
    i_8_415_881_0, i_8_415_896_0, i_8_415_937_0, i_8_415_967_0,
    i_8_415_968_0, i_8_415_974_0, i_8_415_1071_0, i_8_415_1085_0,
    i_8_415_1102_0, i_8_415_1117_0, i_8_415_1163_0, i_8_415_1228_0,
    i_8_415_1253_0, i_8_415_1260_0, i_8_415_1262_0, i_8_415_1270_0,
    i_8_415_1273_0, i_8_415_1295_0, i_8_415_1432_0, i_8_415_1463_0,
    i_8_415_1495_0, i_8_415_1496_0, i_8_415_1498_0, i_8_415_1514_0,
    i_8_415_1516_0, i_8_415_1519_0, i_8_415_1526_0, i_8_415_1531_0,
    i_8_415_1596_0, i_8_415_1638_0, i_8_415_1651_0, i_8_415_1676_0,
    i_8_415_1682_0, i_8_415_1688_0, i_8_415_1694_0, i_8_415_1702_0,
    i_8_415_1729_0, i_8_415_1747_0, i_8_415_1760_0, i_8_415_1769_0,
    i_8_415_1773_0, i_8_415_1784_0, i_8_415_1819_0, i_8_415_1822_0,
    i_8_415_1837_0, i_8_415_1873_0, i_8_415_1881_0, i_8_415_1884_0,
    i_8_415_1891_0, i_8_415_1912_0, i_8_415_1927_0, i_8_415_1939_0,
    i_8_415_1965_0, i_8_415_1971_0, i_8_415_1980_0, i_8_415_2017_0,
    i_8_415_2054_0, i_8_415_2072_0, i_8_415_2146_0, i_8_415_2152_0,
    i_8_415_2244_0, i_8_415_2246_0, i_8_415_2270_0,
    o_8_415_0_0  );
  input  i_8_415_13_0, i_8_415_38_0, i_8_415_40_0, i_8_415_75_0,
    i_8_415_113_0, i_8_415_135_0, i_8_415_193_0, i_8_415_226_0,
    i_8_415_262_0, i_8_415_264_0, i_8_415_308_0, i_8_415_320_0,
    i_8_415_361_0, i_8_415_362_0, i_8_415_422_0, i_8_415_490_0,
    i_8_415_509_0, i_8_415_514_0, i_8_415_520_0, i_8_415_535_0,
    i_8_415_543_0, i_8_415_544_0, i_8_415_580_0, i_8_415_604_0,
    i_8_415_612_0, i_8_415_613_0, i_8_415_634_0, i_8_415_653_0,
    i_8_415_656_0, i_8_415_748_0, i_8_415_751_0, i_8_415_756_0,
    i_8_415_766_0, i_8_415_800_0, i_8_415_802_0, i_8_415_815_0,
    i_8_415_837_0, i_8_415_881_0, i_8_415_896_0, i_8_415_937_0,
    i_8_415_967_0, i_8_415_968_0, i_8_415_974_0, i_8_415_1071_0,
    i_8_415_1085_0, i_8_415_1102_0, i_8_415_1117_0, i_8_415_1163_0,
    i_8_415_1228_0, i_8_415_1253_0, i_8_415_1260_0, i_8_415_1262_0,
    i_8_415_1270_0, i_8_415_1273_0, i_8_415_1295_0, i_8_415_1432_0,
    i_8_415_1463_0, i_8_415_1495_0, i_8_415_1496_0, i_8_415_1498_0,
    i_8_415_1514_0, i_8_415_1516_0, i_8_415_1519_0, i_8_415_1526_0,
    i_8_415_1531_0, i_8_415_1596_0, i_8_415_1638_0, i_8_415_1651_0,
    i_8_415_1676_0, i_8_415_1682_0, i_8_415_1688_0, i_8_415_1694_0,
    i_8_415_1702_0, i_8_415_1729_0, i_8_415_1747_0, i_8_415_1760_0,
    i_8_415_1769_0, i_8_415_1773_0, i_8_415_1784_0, i_8_415_1819_0,
    i_8_415_1822_0, i_8_415_1837_0, i_8_415_1873_0, i_8_415_1881_0,
    i_8_415_1884_0, i_8_415_1891_0, i_8_415_1912_0, i_8_415_1927_0,
    i_8_415_1939_0, i_8_415_1965_0, i_8_415_1971_0, i_8_415_1980_0,
    i_8_415_2017_0, i_8_415_2054_0, i_8_415_2072_0, i_8_415_2146_0,
    i_8_415_2152_0, i_8_415_2244_0, i_8_415_2246_0, i_8_415_2270_0;
  output o_8_415_0_0;
  assign o_8_415_0_0 = 0;
endmodule



// Benchmark "kernel_8_416" written by ABC on Sun Jul 19 10:10:21 2020

module kernel_8_416 ( 
    i_8_416_27_0, i_8_416_31_0, i_8_416_34_0, i_8_416_96_0, i_8_416_97_0,
    i_8_416_114_0, i_8_416_115_0, i_8_416_116_0, i_8_416_166_0,
    i_8_416_184_0, i_8_416_224_0, i_8_416_241_0, i_8_416_300_0,
    i_8_416_303_0, i_8_416_367_0, i_8_416_369_0, i_8_416_381_0,
    i_8_416_382_0, i_8_416_421_0, i_8_416_492_0, i_8_416_508_0,
    i_8_416_525_0, i_8_416_572_0, i_8_416_588_0, i_8_416_616_0,
    i_8_416_633_0, i_8_416_634_0, i_8_416_662_0, i_8_416_701_0,
    i_8_416_703_0, i_8_416_704_0, i_8_416_706_0, i_8_416_707_0,
    i_8_416_714_0, i_8_416_754_0, i_8_416_778_0, i_8_416_859_0,
    i_8_416_887_0, i_8_416_940_0, i_8_416_941_0, i_8_416_994_0,
    i_8_416_1030_0, i_8_416_1096_0, i_8_416_1113_0, i_8_416_1114_0,
    i_8_416_1120_0, i_8_416_1159_0, i_8_416_1182_0, i_8_416_1183_0,
    i_8_416_1186_0, i_8_416_1188_0, i_8_416_1197_0, i_8_416_1284_0,
    i_8_416_1292_0, i_8_416_1299_0, i_8_416_1307_0, i_8_416_1308_0,
    i_8_416_1330_0, i_8_416_1411_0, i_8_416_1412_0, i_8_416_1437_0,
    i_8_416_1535_0, i_8_416_1545_0, i_8_416_1551_0, i_8_416_1591_0,
    i_8_416_1635_0, i_8_416_1642_0, i_8_416_1654_0, i_8_416_1678_0,
    i_8_416_1684_0, i_8_416_1696_0, i_8_416_1731_0, i_8_416_1741_0,
    i_8_416_1742_0, i_8_416_1744_0, i_8_416_1751_0, i_8_416_1762_0,
    i_8_416_1785_0, i_8_416_1821_0, i_8_416_1825_0, i_8_416_1831_0,
    i_8_416_1858_0, i_8_416_1939_0, i_8_416_2047_0, i_8_416_2050_0,
    i_8_416_2075_0, i_8_416_2119_0, i_8_416_2122_0, i_8_416_2123_0,
    i_8_416_2153_0, i_8_416_2157_0, i_8_416_2172_0, i_8_416_2189_0,
    i_8_416_2214_0, i_8_416_2215_0, i_8_416_2217_0, i_8_416_2218_0,
    i_8_416_2245_0, i_8_416_2248_0, i_8_416_2303_0,
    o_8_416_0_0  );
  input  i_8_416_27_0, i_8_416_31_0, i_8_416_34_0, i_8_416_96_0,
    i_8_416_97_0, i_8_416_114_0, i_8_416_115_0, i_8_416_116_0,
    i_8_416_166_0, i_8_416_184_0, i_8_416_224_0, i_8_416_241_0,
    i_8_416_300_0, i_8_416_303_0, i_8_416_367_0, i_8_416_369_0,
    i_8_416_381_0, i_8_416_382_0, i_8_416_421_0, i_8_416_492_0,
    i_8_416_508_0, i_8_416_525_0, i_8_416_572_0, i_8_416_588_0,
    i_8_416_616_0, i_8_416_633_0, i_8_416_634_0, i_8_416_662_0,
    i_8_416_701_0, i_8_416_703_0, i_8_416_704_0, i_8_416_706_0,
    i_8_416_707_0, i_8_416_714_0, i_8_416_754_0, i_8_416_778_0,
    i_8_416_859_0, i_8_416_887_0, i_8_416_940_0, i_8_416_941_0,
    i_8_416_994_0, i_8_416_1030_0, i_8_416_1096_0, i_8_416_1113_0,
    i_8_416_1114_0, i_8_416_1120_0, i_8_416_1159_0, i_8_416_1182_0,
    i_8_416_1183_0, i_8_416_1186_0, i_8_416_1188_0, i_8_416_1197_0,
    i_8_416_1284_0, i_8_416_1292_0, i_8_416_1299_0, i_8_416_1307_0,
    i_8_416_1308_0, i_8_416_1330_0, i_8_416_1411_0, i_8_416_1412_0,
    i_8_416_1437_0, i_8_416_1535_0, i_8_416_1545_0, i_8_416_1551_0,
    i_8_416_1591_0, i_8_416_1635_0, i_8_416_1642_0, i_8_416_1654_0,
    i_8_416_1678_0, i_8_416_1684_0, i_8_416_1696_0, i_8_416_1731_0,
    i_8_416_1741_0, i_8_416_1742_0, i_8_416_1744_0, i_8_416_1751_0,
    i_8_416_1762_0, i_8_416_1785_0, i_8_416_1821_0, i_8_416_1825_0,
    i_8_416_1831_0, i_8_416_1858_0, i_8_416_1939_0, i_8_416_2047_0,
    i_8_416_2050_0, i_8_416_2075_0, i_8_416_2119_0, i_8_416_2122_0,
    i_8_416_2123_0, i_8_416_2153_0, i_8_416_2157_0, i_8_416_2172_0,
    i_8_416_2189_0, i_8_416_2214_0, i_8_416_2215_0, i_8_416_2217_0,
    i_8_416_2218_0, i_8_416_2245_0, i_8_416_2248_0, i_8_416_2303_0;
  output o_8_416_0_0;
  assign o_8_416_0_0 = ~((~i_8_416_31_0 & ((~i_8_416_34_0 & i_8_416_706_0 & ~i_8_416_1182_0 & ~i_8_416_1183_0 & ~i_8_416_1742_0) | (~i_8_416_572_0 & ~i_8_416_778_0 & ~i_8_416_994_0 & ~i_8_416_1696_0 & ~i_8_416_2245_0))) | (i_8_416_616_0 & ((i_8_416_34_0 & ~i_8_416_941_0 & ~i_8_416_1307_0 & ~i_8_416_1535_0 & ~i_8_416_1642_0 & ~i_8_416_1654_0 & i_8_416_1858_0) | (~i_8_416_114_0 & ~i_8_416_1762_0 & ~i_8_416_1858_0 & ~i_8_416_2075_0 & ~i_8_416_2217_0))) | (~i_8_416_1182_0 & ((~i_8_416_940_0 & ((~i_8_416_369_0 & ~i_8_416_572_0 & ~i_8_416_887_0 & ~i_8_416_1183_0 & ~i_8_416_1197_0 & ~i_8_416_2248_0) | (~i_8_416_1535_0 & ~i_8_416_2047_0 & ~i_8_416_2172_0 & ~i_8_416_2303_0))) | (i_8_416_707_0 & ~i_8_416_1742_0 & ~i_8_416_2217_0) | (~i_8_416_27_0 & ~i_8_416_116_0 & ~i_8_416_166_0 & ~i_8_416_754_0 & ~i_8_416_1183_0 & ~i_8_416_1535_0 & ~i_8_416_1591_0 & ~i_8_416_2245_0))) | (~i_8_416_166_0 & ((~i_8_416_859_0 & ~i_8_416_1307_0 & ~i_8_416_2119_0 & ~i_8_416_2123_0) | (~i_8_416_1186_0 & ~i_8_416_1437_0 & ~i_8_416_2172_0 & ~i_8_416_2215_0))) | (~i_8_416_1831_0 & ((~i_8_416_616_0 & ~i_8_416_634_0 & ~i_8_416_1299_0) | (~i_8_416_701_0 & ~i_8_416_940_0 & ~i_8_416_1696_0 & ~i_8_416_1858_0 & ~i_8_416_2050_0))) | (~i_8_416_34_0 & i_8_416_367_0 & ~i_8_416_994_0 & ~i_8_416_1684_0) | (~i_8_416_941_0 & ~i_8_416_2047_0 & ~i_8_416_2050_0 & ~i_8_416_2123_0 & ~i_8_416_2214_0) | (i_8_416_1821_0 & ~i_8_416_2215_0) | (i_8_416_701_0 & ~i_8_416_1188_0 & ~i_8_416_1292_0 & ~i_8_416_1437_0 & ~i_8_416_2218_0));
endmodule



// Benchmark "kernel_8_417" written by ABC on Sun Jul 19 10:10:23 2020

module kernel_8_417 ( 
    i_8_417_12_0, i_8_417_52_0, i_8_417_114_0, i_8_417_193_0,
    i_8_417_220_0, i_8_417_226_0, i_8_417_279_0, i_8_417_318_0,
    i_8_417_319_0, i_8_417_321_0, i_8_417_365_0, i_8_417_397_0,
    i_8_417_399_0, i_8_417_400_0, i_8_417_402_0, i_8_417_427_0,
    i_8_417_428_0, i_8_417_440_0, i_8_417_471_0, i_8_417_490_0,
    i_8_417_492_0, i_8_417_525_0, i_8_417_582_0, i_8_417_583_0,
    i_8_417_584_0, i_8_417_612_0, i_8_417_639_0, i_8_417_642_0,
    i_8_417_645_0, i_8_417_646_0, i_8_417_660_0, i_8_417_748_0,
    i_8_417_759_0, i_8_417_762_0, i_8_417_799_0, i_8_417_808_0,
    i_8_417_843_0, i_8_417_844_0, i_8_417_852_0, i_8_417_855_0,
    i_8_417_877_0, i_8_417_933_0, i_8_417_934_0, i_8_417_966_0,
    i_8_417_967_0, i_8_417_1179_0, i_8_417_1228_0, i_8_417_1240_0,
    i_8_417_1257_0, i_8_417_1263_0, i_8_417_1281_0, i_8_417_1284_0,
    i_8_417_1285_0, i_8_417_1303_0, i_8_417_1307_0, i_8_417_1318_0,
    i_8_417_1330_0, i_8_417_1359_0, i_8_417_1366_0, i_8_417_1435_0,
    i_8_417_1438_0, i_8_417_1440_0, i_8_417_1443_0, i_8_417_1456_0,
    i_8_417_1461_0, i_8_417_1464_0, i_8_417_1470_0, i_8_417_1493_0,
    i_8_417_1559_0, i_8_417_1564_0, i_8_417_1662_0, i_8_417_1677_0,
    i_8_417_1713_0, i_8_417_1717_0, i_8_417_1756_0, i_8_417_1876_0,
    i_8_417_1893_0, i_8_417_1935_0, i_8_417_1939_0, i_8_417_1966_0,
    i_8_417_1997_0, i_8_417_2041_0, i_8_417_2057_0, i_8_417_2091_0,
    i_8_417_2134_0, i_8_417_2146_0, i_8_417_2147_0, i_8_417_2149_0,
    i_8_417_2154_0, i_8_417_2170_0, i_8_417_2171_0, i_8_417_2173_0,
    i_8_417_2174_0, i_8_417_2175_0, i_8_417_2177_0, i_8_417_2185_0,
    i_8_417_2193_0, i_8_417_2194_0, i_8_417_2216_0, i_8_417_2232_0,
    o_8_417_0_0  );
  input  i_8_417_12_0, i_8_417_52_0, i_8_417_114_0, i_8_417_193_0,
    i_8_417_220_0, i_8_417_226_0, i_8_417_279_0, i_8_417_318_0,
    i_8_417_319_0, i_8_417_321_0, i_8_417_365_0, i_8_417_397_0,
    i_8_417_399_0, i_8_417_400_0, i_8_417_402_0, i_8_417_427_0,
    i_8_417_428_0, i_8_417_440_0, i_8_417_471_0, i_8_417_490_0,
    i_8_417_492_0, i_8_417_525_0, i_8_417_582_0, i_8_417_583_0,
    i_8_417_584_0, i_8_417_612_0, i_8_417_639_0, i_8_417_642_0,
    i_8_417_645_0, i_8_417_646_0, i_8_417_660_0, i_8_417_748_0,
    i_8_417_759_0, i_8_417_762_0, i_8_417_799_0, i_8_417_808_0,
    i_8_417_843_0, i_8_417_844_0, i_8_417_852_0, i_8_417_855_0,
    i_8_417_877_0, i_8_417_933_0, i_8_417_934_0, i_8_417_966_0,
    i_8_417_967_0, i_8_417_1179_0, i_8_417_1228_0, i_8_417_1240_0,
    i_8_417_1257_0, i_8_417_1263_0, i_8_417_1281_0, i_8_417_1284_0,
    i_8_417_1285_0, i_8_417_1303_0, i_8_417_1307_0, i_8_417_1318_0,
    i_8_417_1330_0, i_8_417_1359_0, i_8_417_1366_0, i_8_417_1435_0,
    i_8_417_1438_0, i_8_417_1440_0, i_8_417_1443_0, i_8_417_1456_0,
    i_8_417_1461_0, i_8_417_1464_0, i_8_417_1470_0, i_8_417_1493_0,
    i_8_417_1559_0, i_8_417_1564_0, i_8_417_1662_0, i_8_417_1677_0,
    i_8_417_1713_0, i_8_417_1717_0, i_8_417_1756_0, i_8_417_1876_0,
    i_8_417_1893_0, i_8_417_1935_0, i_8_417_1939_0, i_8_417_1966_0,
    i_8_417_1997_0, i_8_417_2041_0, i_8_417_2057_0, i_8_417_2091_0,
    i_8_417_2134_0, i_8_417_2146_0, i_8_417_2147_0, i_8_417_2149_0,
    i_8_417_2154_0, i_8_417_2170_0, i_8_417_2171_0, i_8_417_2173_0,
    i_8_417_2174_0, i_8_417_2175_0, i_8_417_2177_0, i_8_417_2185_0,
    i_8_417_2193_0, i_8_417_2194_0, i_8_417_2216_0, i_8_417_2232_0;
  output o_8_417_0_0;
  assign o_8_417_0_0 = ~((~i_8_417_748_0 & ((~i_8_417_114_0 & ((~i_8_417_52_0 & i_8_417_220_0 & ~i_8_417_427_0 & ~i_8_417_428_0 & ~i_8_417_855_0 & ~i_8_417_1179_0 & ~i_8_417_1330_0 & ~i_8_417_2041_0) | (~i_8_417_220_0 & ~i_8_417_321_0 & ~i_8_417_583_0 & ~i_8_417_584_0 & ~i_8_417_808_0 & ~i_8_417_933_0 & ~i_8_417_1228_0 & ~i_8_417_1359_0 & i_8_417_1435_0 & ~i_8_417_1493_0 & ~i_8_417_1662_0 & ~i_8_417_2091_0))) | (~i_8_417_319_0 & ~i_8_417_583_0 & ~i_8_417_808_0 & ~i_8_417_1240_0 & ~i_8_417_1366_0 & i_8_417_2057_0))) | (~i_8_417_52_0 & ((~i_8_417_12_0 & ~i_8_417_400_0 & i_8_417_428_0 & ~i_8_417_639_0 & ~i_8_417_1438_0 & ~i_8_417_1443_0) | (~i_8_417_279_0 & ~i_8_417_321_0 & ~i_8_417_397_0 & ~i_8_417_399_0 & ~i_8_417_646_0 & ~i_8_417_1240_0 & ~i_8_417_1257_0 & ~i_8_417_1281_0 & ~i_8_417_1359_0 & ~i_8_417_1470_0 & ~i_8_417_2193_0 & ~i_8_417_2194_0))) | (~i_8_417_646_0 & ((~i_8_417_12_0 & ((~i_8_417_397_0 & ~i_8_417_399_0 & ~i_8_417_402_0 & i_8_417_525_0 & ~i_8_417_584_0 & ~i_8_417_645_0 & ~i_8_417_1263_0) | (~i_8_417_639_0 & ~i_8_417_933_0 & ~i_8_417_934_0 & ~i_8_417_1461_0 & i_8_417_1677_0 & ~i_8_417_1939_0))) | (~i_8_417_397_0 & ((~i_8_417_400_0 & ((~i_8_417_321_0 & ((~i_8_417_402_0 & ~i_8_417_427_0 & ~i_8_417_582_0 & ~i_8_417_843_0 & ~i_8_417_933_0 & ~i_8_417_1179_0 & ~i_8_417_1366_0 & ~i_8_417_1440_0 & ~i_8_417_1456_0 & ~i_8_417_1461_0 & ~i_8_417_1564_0 & ~i_8_417_1935_0) | (~i_8_417_279_0 & ~i_8_417_440_0 & ~i_8_417_583_0 & ~i_8_417_584_0 & ~i_8_417_660_0 & i_8_417_843_0 & ~i_8_417_934_0 & ~i_8_417_1228_0 & ~i_8_417_1263_0 & ~i_8_417_1717_0 & ~i_8_417_2170_0 & ~i_8_417_2216_0))) | (~i_8_417_399_0 & ~i_8_417_440_0 & ~i_8_417_582_0 & ~i_8_417_583_0 & ~i_8_417_639_0 & ~i_8_417_843_0 & ~i_8_417_1257_0 & ~i_8_417_1440_0 & ~i_8_417_1564_0 & ~i_8_417_1893_0 & ~i_8_417_2149_0 & ~i_8_417_2194_0))) | (~i_8_417_402_0 & ~i_8_417_799_0 & ~i_8_417_843_0 & ~i_8_417_1228_0 & ~i_8_417_1257_0 & ~i_8_417_1359_0 & ~i_8_417_1440_0 & ~i_8_417_1893_0 & ~i_8_417_2041_0 & ~i_8_417_2091_0 & ~i_8_417_2134_0) | (~i_8_417_525_0 & ~i_8_417_584_0 & ~i_8_417_642_0 & ~i_8_417_808_0 & ~i_8_417_966_0 & i_8_417_2149_0 & i_8_417_2185_0 & ~i_8_417_2194_0))) | (~i_8_417_1330_0 & ~i_8_417_1935_0 & ((~i_8_417_318_0 & ~i_8_417_492_0 & ~i_8_417_639_0 & ~i_8_417_660_0 & ~i_8_417_808_0 & ~i_8_417_1440_0 & ~i_8_417_2147_0) | (~i_8_417_399_0 & ~i_8_417_400_0 & ~i_8_417_428_0 & ~i_8_417_582_0 & ~i_8_417_584_0 & ~i_8_417_799_0 & ~i_8_417_933_0 & ~i_8_417_966_0 & ~i_8_417_1179_0 & ~i_8_417_1359_0 & ~i_8_417_1564_0 & ~i_8_417_2041_0 & ~i_8_417_2175_0 & ~i_8_417_2177_0 & ~i_8_417_2194_0))))) | (~i_8_417_934_0 & ((~i_8_417_397_0 & ((~i_8_417_319_0 & ~i_8_417_1359_0 & ((~i_8_417_399_0 & ~i_8_417_583_0 & ~i_8_417_639_0 & ~i_8_417_808_0 & ~i_8_417_933_0 & ~i_8_417_1284_0 & ~i_8_417_1366_0 & ~i_8_417_1435_0 & ~i_8_417_1564_0 & ~i_8_417_2057_0) | (~i_8_417_428_0 & ~i_8_417_582_0 & ~i_8_417_844_0 & ~i_8_417_1228_0 & ~i_8_417_1257_0 & ~i_8_417_1443_0 & ~i_8_417_1713_0 & ~i_8_417_1893_0 & ~i_8_417_2175_0 & ~i_8_417_2185_0))) | (~i_8_417_321_0 & ~i_8_417_400_0 & ~i_8_417_402_0 & ~i_8_417_645_0 & ~i_8_417_1179_0 & i_8_417_1470_0 & ~i_8_417_1662_0 & ~i_8_417_1756_0 & ~i_8_417_1876_0 & ~i_8_417_1939_0))) | (~i_8_417_321_0 & i_8_417_471_0 & ~i_8_417_799_0 & ~i_8_417_1257_0 & ~i_8_417_1359_0 & ~i_8_417_1443_0 & ~i_8_417_1893_0 & ~i_8_417_1939_0))) | (~i_8_417_967_0 & ~i_8_417_2185_0 & ((~i_8_417_397_0 & ~i_8_417_1359_0 & ~i_8_417_1440_0 & ((~i_8_417_399_0 & ~i_8_417_402_0 & ~i_8_417_583_0 & ~i_8_417_584_0 & ~i_8_417_645_0 & ~i_8_417_1318_0 & ~i_8_417_1366_0) | (~i_8_417_400_0 & ~i_8_417_492_0 & ~i_8_417_808_0 & ~i_8_417_1284_0 & ~i_8_417_2154_0))) | (i_8_417_226_0 & ~i_8_417_583_0 & i_8_417_612_0 & ~i_8_417_843_0 & ~i_8_417_1997_0))) | (~i_8_417_583_0 & ((~i_8_417_319_0 & ~i_8_417_1440_0 & i_8_417_2174_0) | (~i_8_417_318_0 & ~i_8_417_400_0 & i_8_417_525_0 & ~i_8_417_1438_0 & ~i_8_417_2193_0))) | (i_8_417_1461_0 & i_8_417_1876_0) | (~i_8_417_440_0 & ~i_8_417_1359_0 & i_8_417_1559_0 & ~i_8_417_1939_0) | (i_8_417_492_0 & ~i_8_417_582_0 & i_8_417_966_0 & ~i_8_417_1257_0 & ~i_8_417_1366_0 & ~i_8_417_1443_0 & i_8_417_1966_0));
endmodule



// Benchmark "kernel_8_418" written by ABC on Sun Jul 19 10:10:24 2020

module kernel_8_418 ( 
    i_8_418_21_0, i_8_418_30_0, i_8_418_139_0, i_8_418_140_0,
    i_8_418_184_0, i_8_418_193_0, i_8_418_229_0, i_8_418_246_0,
    i_8_418_247_0, i_8_418_262_0, i_8_418_274_0, i_8_418_292_0,
    i_8_418_356_0, i_8_418_373_0, i_8_418_417_0, i_8_418_420_0,
    i_8_418_430_0, i_8_418_461_0, i_8_418_462_0, i_8_418_463_0,
    i_8_418_474_0, i_8_418_517_0, i_8_418_529_0, i_8_418_557_0,
    i_8_418_571_0, i_8_418_612_0, i_8_418_615_0, i_8_418_634_0,
    i_8_418_671_0, i_8_418_678_0, i_8_418_681_0, i_8_418_703_0,
    i_8_418_715_0, i_8_418_730_0, i_8_418_761_0, i_8_418_792_0,
    i_8_418_793_0, i_8_418_795_0, i_8_418_837_0, i_8_418_849_0,
    i_8_418_880_0, i_8_418_959_0, i_8_418_993_0, i_8_418_996_0,
    i_8_418_997_0, i_8_418_1081_0, i_8_418_1114_0, i_8_418_1157_0,
    i_8_418_1159_0, i_8_418_1192_0, i_8_418_1236_0, i_8_418_1237_0,
    i_8_418_1259_0, i_8_418_1270_0, i_8_418_1274_0, i_8_418_1281_0,
    i_8_418_1283_0, i_8_418_1284_0, i_8_418_1300_0, i_8_418_1307_0,
    i_8_418_1326_0, i_8_418_1387_0, i_8_418_1468_0, i_8_418_1483_0,
    i_8_418_1493_0, i_8_418_1539_0, i_8_418_1542_0, i_8_418_1546_0,
    i_8_418_1597_0, i_8_418_1598_0, i_8_418_1659_0, i_8_418_1731_0,
    i_8_418_1752_0, i_8_418_1776_0, i_8_418_1785_0, i_8_418_1803_0,
    i_8_418_1804_0, i_8_418_1812_0, i_8_418_1818_0, i_8_418_1820_0,
    i_8_418_1855_0, i_8_418_1867_0, i_8_418_1874_0, i_8_418_1876_0,
    i_8_418_1894_0, i_8_418_1912_0, i_8_418_1918_0, i_8_418_1919_0,
    i_8_418_1997_0, i_8_418_2007_0, i_8_418_2045_0, i_8_418_2065_0,
    i_8_418_2093_0, i_8_418_2109_0, i_8_418_2137_0, i_8_418_2158_0,
    i_8_418_2192_0, i_8_418_2254_0, i_8_418_2257_0, i_8_418_2291_0,
    o_8_418_0_0  );
  input  i_8_418_21_0, i_8_418_30_0, i_8_418_139_0, i_8_418_140_0,
    i_8_418_184_0, i_8_418_193_0, i_8_418_229_0, i_8_418_246_0,
    i_8_418_247_0, i_8_418_262_0, i_8_418_274_0, i_8_418_292_0,
    i_8_418_356_0, i_8_418_373_0, i_8_418_417_0, i_8_418_420_0,
    i_8_418_430_0, i_8_418_461_0, i_8_418_462_0, i_8_418_463_0,
    i_8_418_474_0, i_8_418_517_0, i_8_418_529_0, i_8_418_557_0,
    i_8_418_571_0, i_8_418_612_0, i_8_418_615_0, i_8_418_634_0,
    i_8_418_671_0, i_8_418_678_0, i_8_418_681_0, i_8_418_703_0,
    i_8_418_715_0, i_8_418_730_0, i_8_418_761_0, i_8_418_792_0,
    i_8_418_793_0, i_8_418_795_0, i_8_418_837_0, i_8_418_849_0,
    i_8_418_880_0, i_8_418_959_0, i_8_418_993_0, i_8_418_996_0,
    i_8_418_997_0, i_8_418_1081_0, i_8_418_1114_0, i_8_418_1157_0,
    i_8_418_1159_0, i_8_418_1192_0, i_8_418_1236_0, i_8_418_1237_0,
    i_8_418_1259_0, i_8_418_1270_0, i_8_418_1274_0, i_8_418_1281_0,
    i_8_418_1283_0, i_8_418_1284_0, i_8_418_1300_0, i_8_418_1307_0,
    i_8_418_1326_0, i_8_418_1387_0, i_8_418_1468_0, i_8_418_1483_0,
    i_8_418_1493_0, i_8_418_1539_0, i_8_418_1542_0, i_8_418_1546_0,
    i_8_418_1597_0, i_8_418_1598_0, i_8_418_1659_0, i_8_418_1731_0,
    i_8_418_1752_0, i_8_418_1776_0, i_8_418_1785_0, i_8_418_1803_0,
    i_8_418_1804_0, i_8_418_1812_0, i_8_418_1818_0, i_8_418_1820_0,
    i_8_418_1855_0, i_8_418_1867_0, i_8_418_1874_0, i_8_418_1876_0,
    i_8_418_1894_0, i_8_418_1912_0, i_8_418_1918_0, i_8_418_1919_0,
    i_8_418_1997_0, i_8_418_2007_0, i_8_418_2045_0, i_8_418_2065_0,
    i_8_418_2093_0, i_8_418_2109_0, i_8_418_2137_0, i_8_418_2158_0,
    i_8_418_2192_0, i_8_418_2254_0, i_8_418_2257_0, i_8_418_2291_0;
  output o_8_418_0_0;
  assign o_8_418_0_0 = 0;
endmodule



// Benchmark "kernel_8_419" written by ABC on Sun Jul 19 10:10:26 2020

module kernel_8_419 ( 
    i_8_419_44_0, i_8_419_93_0, i_8_419_95_0, i_8_419_131_0, i_8_419_174_0,
    i_8_419_175_0, i_8_419_185_0, i_8_419_223_0, i_8_419_241_0,
    i_8_419_264_0, i_8_419_276_0, i_8_419_282_0, i_8_419_302_0,
    i_8_419_309_0, i_8_419_310_0, i_8_419_312_0, i_8_419_314_0,
    i_8_419_338_0, i_8_419_391_0, i_8_419_430_0, i_8_419_527_0,
    i_8_419_591_0, i_8_419_592_0, i_8_419_593_0, i_8_419_607_0,
    i_8_419_617_0, i_8_419_626_0, i_8_419_655_0, i_8_419_661_0,
    i_8_419_663_0, i_8_419_664_0, i_8_419_692_0, i_8_419_822_0,
    i_8_419_826_0, i_8_419_827_0, i_8_419_838_0, i_8_419_955_0,
    i_8_419_959_0, i_8_419_969_0, i_8_419_970_0, i_8_419_996_0,
    i_8_419_1003_0, i_8_419_1047_0, i_8_419_1049_0, i_8_419_1060_0,
    i_8_419_1061_0, i_8_419_1092_0, i_8_419_1110_0, i_8_419_1159_0,
    i_8_419_1191_0, i_8_419_1192_0, i_8_419_1193_0, i_8_419_1236_0,
    i_8_419_1263_0, i_8_419_1264_0, i_8_419_1265_0, i_8_419_1278_0,
    i_8_419_1279_0, i_8_419_1280_0, i_8_419_1282_0, i_8_419_1300_0,
    i_8_419_1306_0, i_8_419_1308_0, i_8_419_1366_0, i_8_419_1410_0,
    i_8_419_1411_0, i_8_419_1412_0, i_8_419_1434_0, i_8_419_1435_0,
    i_8_419_1436_0, i_8_419_1471_0, i_8_419_1641_0, i_8_419_1643_0,
    i_8_419_1644_0, i_8_419_1645_0, i_8_419_1646_0, i_8_419_1653_0,
    i_8_419_1655_0, i_8_419_1662_0, i_8_419_1663_0, i_8_419_1664_0,
    i_8_419_1715_0, i_8_419_1819_0, i_8_419_1877_0, i_8_419_1899_0,
    i_8_419_1964_0, i_8_419_2073_0, i_8_419_2093_0, i_8_419_2135_0,
    i_8_419_2136_0, i_8_419_2141_0, i_8_419_2164_0, i_8_419_2175_0,
    i_8_419_2193_0, i_8_419_2215_0, i_8_419_2216_0, i_8_419_2219_0,
    i_8_419_2263_0, i_8_419_2264_0, i_8_419_2290_0,
    o_8_419_0_0  );
  input  i_8_419_44_0, i_8_419_93_0, i_8_419_95_0, i_8_419_131_0,
    i_8_419_174_0, i_8_419_175_0, i_8_419_185_0, i_8_419_223_0,
    i_8_419_241_0, i_8_419_264_0, i_8_419_276_0, i_8_419_282_0,
    i_8_419_302_0, i_8_419_309_0, i_8_419_310_0, i_8_419_312_0,
    i_8_419_314_0, i_8_419_338_0, i_8_419_391_0, i_8_419_430_0,
    i_8_419_527_0, i_8_419_591_0, i_8_419_592_0, i_8_419_593_0,
    i_8_419_607_0, i_8_419_617_0, i_8_419_626_0, i_8_419_655_0,
    i_8_419_661_0, i_8_419_663_0, i_8_419_664_0, i_8_419_692_0,
    i_8_419_822_0, i_8_419_826_0, i_8_419_827_0, i_8_419_838_0,
    i_8_419_955_0, i_8_419_959_0, i_8_419_969_0, i_8_419_970_0,
    i_8_419_996_0, i_8_419_1003_0, i_8_419_1047_0, i_8_419_1049_0,
    i_8_419_1060_0, i_8_419_1061_0, i_8_419_1092_0, i_8_419_1110_0,
    i_8_419_1159_0, i_8_419_1191_0, i_8_419_1192_0, i_8_419_1193_0,
    i_8_419_1236_0, i_8_419_1263_0, i_8_419_1264_0, i_8_419_1265_0,
    i_8_419_1278_0, i_8_419_1279_0, i_8_419_1280_0, i_8_419_1282_0,
    i_8_419_1300_0, i_8_419_1306_0, i_8_419_1308_0, i_8_419_1366_0,
    i_8_419_1410_0, i_8_419_1411_0, i_8_419_1412_0, i_8_419_1434_0,
    i_8_419_1435_0, i_8_419_1436_0, i_8_419_1471_0, i_8_419_1641_0,
    i_8_419_1643_0, i_8_419_1644_0, i_8_419_1645_0, i_8_419_1646_0,
    i_8_419_1653_0, i_8_419_1655_0, i_8_419_1662_0, i_8_419_1663_0,
    i_8_419_1664_0, i_8_419_1715_0, i_8_419_1819_0, i_8_419_1877_0,
    i_8_419_1899_0, i_8_419_1964_0, i_8_419_2073_0, i_8_419_2093_0,
    i_8_419_2135_0, i_8_419_2136_0, i_8_419_2141_0, i_8_419_2164_0,
    i_8_419_2175_0, i_8_419_2193_0, i_8_419_2215_0, i_8_419_2216_0,
    i_8_419_2219_0, i_8_419_2263_0, i_8_419_2264_0, i_8_419_2290_0;
  output o_8_419_0_0;
  assign o_8_419_0_0 = ~((~i_8_419_1662_0 & ((~i_8_419_2263_0 & ((~i_8_419_44_0 & ~i_8_419_1049_0 & ((~i_8_419_276_0 & ~i_8_419_310_0 & ~i_8_419_430_0 & ~i_8_419_617_0 & ~i_8_419_692_0 & ~i_8_419_1060_0 & ~i_8_419_1191_0 & ~i_8_419_1192_0 & ~i_8_419_1282_0 & ~i_8_419_1410_0 & ~i_8_419_1645_0 & ~i_8_419_1663_0 & ~i_8_419_1715_0 & ~i_8_419_1964_0) | (~i_8_419_174_0 & ~i_8_419_309_0 & ~i_8_419_312_0 & ~i_8_419_314_0 & ~i_8_419_955_0 & ~i_8_419_969_0 & ~i_8_419_1061_0 & ~i_8_419_1308_0 & ~i_8_419_1641_0 & ~i_8_419_2073_0 & ~i_8_419_2093_0 & ~i_8_419_2141_0))) | (~i_8_419_314_0 & ~i_8_419_1646_0 & ((~i_8_419_310_0 & ~i_8_419_593_0 & ~i_8_419_692_0 & ~i_8_419_838_0 & ~i_8_419_996_0 & ~i_8_419_1003_0 & ~i_8_419_1047_0 & ~i_8_419_1060_0 & ~i_8_419_1641_0) | (~i_8_419_276_0 & ~i_8_419_309_0 & ~i_8_419_391_0 & ~i_8_419_1191_0 & ~i_8_419_1193_0 & ~i_8_419_1263_0 & ~i_8_419_1308_0 & ~i_8_419_1645_0 & ~i_8_419_1877_0 & ~i_8_419_1899_0 & ~i_8_419_2093_0))))) | (~i_8_419_95_0 & ((~i_8_419_131_0 & ~i_8_419_174_0 & ~i_8_419_1003_0 & ((~i_8_419_185_0 & ~i_8_419_312_0 & ~i_8_419_1193_0 & ~i_8_419_1308_0 & ~i_8_419_1641_0 & ~i_8_419_1644_0 & ~i_8_419_1646_0 & ~i_8_419_1655_0) | (~i_8_419_692_0 & ~i_8_419_955_0 & ~i_8_419_969_0 & ~i_8_419_1061_0 & ~i_8_419_1306_0 & ~i_8_419_1410_0 & ~i_8_419_1411_0 & ~i_8_419_1645_0 & ~i_8_419_1715_0 & ~i_8_419_2164_0))) | (~i_8_419_93_0 & ~i_8_419_312_0 & ~i_8_419_338_0 & ~i_8_419_663_0 & ~i_8_419_1061_0 & ~i_8_419_1191_0 & ~i_8_419_1192_0 & ~i_8_419_1193_0 & ~i_8_419_1663_0 & ~i_8_419_1664_0 & ~i_8_419_1877_0 & ~i_8_419_2135_0 & ~i_8_419_2215_0 & ~i_8_419_2216_0 & ~i_8_419_2219_0))) | (i_8_419_223_0 & ~i_8_419_276_0 & ~i_8_419_959_0 & ~i_8_419_1061_0 & ~i_8_419_1308_0 & ~i_8_419_1643_0 & i_8_419_1655_0) | (~i_8_419_131_0 & ~i_8_419_312_0 & ~i_8_419_592_0 & i_8_419_822_0 & ~i_8_419_1265_0 & ~i_8_419_1471_0 & ~i_8_419_1715_0 & ~i_8_419_2264_0))) | (~i_8_419_310_0 & ((~i_8_419_95_0 & ((~i_8_419_591_0 & ~i_8_419_617_0 & ~i_8_419_1412_0 & i_8_419_1435_0 & i_8_419_1436_0) | (~i_8_419_175_0 & ~i_8_419_185_0 & ~i_8_419_314_0 & ~i_8_419_527_0 & ~i_8_419_1092_0 & ~i_8_419_1411_0 & ~i_8_419_1643_0 & ~i_8_419_1644_0 & ~i_8_419_1655_0 & ~i_8_419_1663_0 & ~i_8_419_1899_0 & ~i_8_419_2263_0 & ~i_8_419_2290_0))) | (~i_8_419_309_0 & ~i_8_419_527_0 & ~i_8_419_617_0 & ~i_8_419_1061_0 & ~i_8_419_1471_0 & ~i_8_419_1641_0 & ~i_8_419_1644_0 & ~i_8_419_1645_0 & ~i_8_419_1653_0 & ~i_8_419_1655_0 & ~i_8_419_1877_0) | (~i_8_419_174_0 & ~i_8_419_264_0 & ~i_8_419_314_0 & ~i_8_419_692_0 & ~i_8_419_1192_0 & i_8_419_1264_0 & ~i_8_419_1308_0 & ~i_8_419_2093_0))) | (~i_8_419_1060_0 & ((~i_8_419_1646_0 & ((~i_8_419_131_0 & ((~i_8_419_312_0 & ~i_8_419_338_0 & ~i_8_419_175_0 & ~i_8_419_241_0 & ~i_8_419_1049_0 & ~i_8_419_1306_0 & ~i_8_419_1641_0 & ~i_8_419_1653_0) | (~i_8_419_655_0 & ~i_8_419_970_0 & ~i_8_419_1092_0 & ~i_8_419_1191_0 & ~i_8_419_1192_0 & ~i_8_419_1193_0 & ~i_8_419_1236_0 & ~i_8_419_1663_0 & ~i_8_419_1664_0 & ~i_8_419_1899_0 & ~i_8_419_2175_0 & ~i_8_419_2215_0))) | (~i_8_419_655_0 & ~i_8_419_838_0 & ~i_8_419_955_0 & ~i_8_419_959_0 & ~i_8_419_1049_0 & ~i_8_419_1192_0 & ~i_8_419_1236_0 & ~i_8_419_1410_0 & ~i_8_419_1411_0 & ~i_8_419_1412_0 & ~i_8_419_1899_0 & ~i_8_419_2175_0))) | (~i_8_419_1653_0 & ((i_8_419_241_0 & i_8_419_822_0 & ~i_8_419_1300_0 & ~i_8_419_1664_0) | (~i_8_419_314_0 & ~i_8_419_338_0 & ~i_8_419_838_0 & ~i_8_419_955_0 & ~i_8_419_1047_0 & ~i_8_419_1092_0 & ~i_8_419_1410_0 & ~i_8_419_1643_0 & ~i_8_419_1644_0 & ~i_8_419_1655_0 & ~i_8_419_1877_0) | (~i_8_419_93_0 & ~i_8_419_309_0 & i_8_419_1644_0 & ~i_8_419_2073_0 & ~i_8_419_2093_0 & i_8_419_2215_0))))) | (~i_8_419_93_0 & ((~i_8_419_276_0 & i_8_419_617_0 & ~i_8_419_1061_0 & i_8_419_1265_0 & ~i_8_419_1411_0 & i_8_419_1436_0 & ~i_8_419_1644_0 & ~i_8_419_1663_0) | (~i_8_419_607_0 & i_8_419_838_0 & ~i_8_419_996_0 & ~i_8_419_1308_0 & ~i_8_419_1643_0 & ~i_8_419_1645_0 & i_8_419_1819_0 & ~i_8_419_2216_0))) | (~i_8_419_175_0 & ((~i_8_419_241_0 & i_8_419_338_0 & ~i_8_419_593_0 & ~i_8_419_692_0 & ~i_8_419_1061_0 & ~i_8_419_1643_0 & ~i_8_419_1653_0 & ~i_8_419_1655_0 & ~i_8_419_1819_0) | (~i_8_419_309_0 & ~i_8_419_314_0 & ~i_8_419_527_0 & i_8_419_607_0 & ~i_8_419_959_0 & ~i_8_419_1192_0 & ~i_8_419_1664_0 & ~i_8_419_2215_0))) | (~i_8_419_1643_0 & ((~i_8_419_185_0 & ~i_8_419_1644_0 & ((~i_8_419_661_0 & ~i_8_419_959_0 & ~i_8_419_1047_0 & ~i_8_419_1410_0 & ~i_8_419_1646_0 & ~i_8_419_1655_0 & ~i_8_419_1663_0 & i_8_419_2216_0) | (~i_8_419_309_0 & ~i_8_419_314_0 & ~i_8_419_1061_0 & ~i_8_419_1191_0 & ~i_8_419_1192_0 & ~i_8_419_2093_0 & ~i_8_419_2175_0 & ~i_8_419_2219_0))) | (~i_8_419_1191_0 & ((i_8_419_827_0 & ~i_8_419_1047_0 & ~i_8_419_1641_0 & ~i_8_419_1646_0 & ~i_8_419_1653_0 & ~i_8_419_2073_0) | (~i_8_419_174_0 & i_8_419_592_0 & ~i_8_419_692_0 & ~i_8_419_1193_0 & ~i_8_419_1645_0 & ~i_8_419_1663_0 & ~i_8_419_1664_0 & ~i_8_419_2164_0 & ~i_8_419_2215_0))))) | (~i_8_419_1877_0 & ((~i_8_419_314_0 & ((i_8_419_592_0 & ~i_8_419_1191_0 & ~i_8_419_1641_0 & ~i_8_419_1645_0 & ~i_8_419_1653_0 & ~i_8_419_1663_0 & ~i_8_419_2093_0 & ~i_8_419_2215_0) | (~i_8_419_276_0 & ~i_8_419_309_0 & ~i_8_419_970_0 & ~i_8_419_1192_0 & ~i_8_419_1646_0 & i_8_419_2136_0 & ~i_8_419_2216_0))) | (~i_8_419_338_0 & ~i_8_419_592_0 & ~i_8_419_996_0 & ~i_8_419_1047_0 & ~i_8_419_1049_0 & ~i_8_419_1061_0 & ~i_8_419_1308_0 & ~i_8_419_1411_0 & ~i_8_419_1434_0 & ~i_8_419_1653_0 & ~i_8_419_1663_0 & ~i_8_419_2263_0))) | (i_8_419_1366_0 & ~i_8_419_1645_0 & ~i_8_419_2175_0 & i_8_419_2219_0));
endmodule



// Benchmark "kernel_8_420" written by ABC on Sun Jul 19 10:10:27 2020

module kernel_8_420 ( 
    i_8_420_22_0, i_8_420_34_0, i_8_420_47_0, i_8_420_50_0, i_8_420_61_0,
    i_8_420_154_0, i_8_420_161_0, i_8_420_208_0, i_8_420_211_0,
    i_8_420_212_0, i_8_420_214_0, i_8_420_290_0, i_8_420_293_0,
    i_8_420_296_0, i_8_420_335_0, i_8_420_391_0, i_8_420_424_0,
    i_8_420_425_0, i_8_420_451_0, i_8_420_452_0, i_8_420_463_0,
    i_8_420_658_0, i_8_420_662_0, i_8_420_673_0, i_8_420_704_0,
    i_8_420_749_0, i_8_420_828_0, i_8_420_829_0, i_8_420_923_0,
    i_8_420_952_0, i_8_420_955_0, i_8_420_1027_0, i_8_420_1036_0,
    i_8_420_1135_0, i_8_420_1136_0, i_8_420_1138_0, i_8_420_1139_0,
    i_8_420_1225_0, i_8_420_1233_0, i_8_420_1272_0, i_8_420_1276_0,
    i_8_420_1286_0, i_8_420_1351_0, i_8_420_1354_0, i_8_420_1355_0,
    i_8_420_1357_0, i_8_420_1358_0, i_8_420_1361_0, i_8_420_1469_0,
    i_8_420_1486_0, i_8_420_1487_0, i_8_420_1506_0, i_8_420_1532_0,
    i_8_420_1533_0, i_8_420_1535_0, i_8_420_1544_0, i_8_420_1550_0,
    i_8_420_1558_0, i_8_420_1559_0, i_8_420_1603_0, i_8_420_1604_0,
    i_8_420_1702_0, i_8_420_1711_0, i_8_420_1714_0, i_8_420_1715_0,
    i_8_420_1719_0, i_8_420_1720_0, i_8_420_1821_0, i_8_420_1861_0,
    i_8_420_1881_0, i_8_420_1886_0, i_8_420_1895_0, i_8_420_1944_0,
    i_8_420_1985_0, i_8_420_1993_0, i_8_420_2002_0, i_8_420_2003_0,
    i_8_420_2005_0, i_8_420_2006_0, i_8_420_2045_0, i_8_420_2053_0,
    i_8_420_2117_0, i_8_420_2129_0, i_8_420_2142_0, i_8_420_2146_0,
    i_8_420_2153_0, i_8_420_2154_0, i_8_420_2179_0, i_8_420_2188_0,
    i_8_420_2191_0, i_8_420_2200_0, i_8_420_2210_0, i_8_420_2225_0,
    i_8_420_2227_0, i_8_420_2246_0, i_8_420_2260_0, i_8_420_2261_0,
    i_8_420_2263_0, i_8_420_2264_0, i_8_420_2273_0,
    o_8_420_0_0  );
  input  i_8_420_22_0, i_8_420_34_0, i_8_420_47_0, i_8_420_50_0,
    i_8_420_61_0, i_8_420_154_0, i_8_420_161_0, i_8_420_208_0,
    i_8_420_211_0, i_8_420_212_0, i_8_420_214_0, i_8_420_290_0,
    i_8_420_293_0, i_8_420_296_0, i_8_420_335_0, i_8_420_391_0,
    i_8_420_424_0, i_8_420_425_0, i_8_420_451_0, i_8_420_452_0,
    i_8_420_463_0, i_8_420_658_0, i_8_420_662_0, i_8_420_673_0,
    i_8_420_704_0, i_8_420_749_0, i_8_420_828_0, i_8_420_829_0,
    i_8_420_923_0, i_8_420_952_0, i_8_420_955_0, i_8_420_1027_0,
    i_8_420_1036_0, i_8_420_1135_0, i_8_420_1136_0, i_8_420_1138_0,
    i_8_420_1139_0, i_8_420_1225_0, i_8_420_1233_0, i_8_420_1272_0,
    i_8_420_1276_0, i_8_420_1286_0, i_8_420_1351_0, i_8_420_1354_0,
    i_8_420_1355_0, i_8_420_1357_0, i_8_420_1358_0, i_8_420_1361_0,
    i_8_420_1469_0, i_8_420_1486_0, i_8_420_1487_0, i_8_420_1506_0,
    i_8_420_1532_0, i_8_420_1533_0, i_8_420_1535_0, i_8_420_1544_0,
    i_8_420_1550_0, i_8_420_1558_0, i_8_420_1559_0, i_8_420_1603_0,
    i_8_420_1604_0, i_8_420_1702_0, i_8_420_1711_0, i_8_420_1714_0,
    i_8_420_1715_0, i_8_420_1719_0, i_8_420_1720_0, i_8_420_1821_0,
    i_8_420_1861_0, i_8_420_1881_0, i_8_420_1886_0, i_8_420_1895_0,
    i_8_420_1944_0, i_8_420_1985_0, i_8_420_1993_0, i_8_420_2002_0,
    i_8_420_2003_0, i_8_420_2005_0, i_8_420_2006_0, i_8_420_2045_0,
    i_8_420_2053_0, i_8_420_2117_0, i_8_420_2129_0, i_8_420_2142_0,
    i_8_420_2146_0, i_8_420_2153_0, i_8_420_2154_0, i_8_420_2179_0,
    i_8_420_2188_0, i_8_420_2191_0, i_8_420_2200_0, i_8_420_2210_0,
    i_8_420_2225_0, i_8_420_2227_0, i_8_420_2246_0, i_8_420_2260_0,
    i_8_420_2261_0, i_8_420_2263_0, i_8_420_2264_0, i_8_420_2273_0;
  output o_8_420_0_0;
  assign o_8_420_0_0 = ~((~i_8_420_452_0 & ((~i_8_420_22_0 & ((~i_8_420_208_0 & ~i_8_420_212_0 & ~i_8_420_1559_0 & ~i_8_420_1714_0 & i_8_420_1886_0 & ~i_8_420_2006_0 & ~i_8_420_2053_0 & ~i_8_420_2200_0 & ~i_8_420_2246_0 & ~i_8_420_2261_0) | (~i_8_420_34_0 & ~i_8_420_154_0 & ~i_8_420_214_0 & ~i_8_420_704_0 & ~i_8_420_1135_0 & ~i_8_420_1139_0 & ~i_8_420_1355_0 & ~i_8_420_1535_0 & ~i_8_420_1711_0 & ~i_8_420_1720_0 & ~i_8_420_2002_0 & ~i_8_420_2003_0 & ~i_8_420_2005_0 & ~i_8_420_2264_0))) | (~i_8_420_2002_0 & ((~i_8_420_50_0 & ~i_8_420_451_0 & ((~i_8_420_34_0 & ~i_8_420_161_0 & ~i_8_420_463_0 & ~i_8_420_1533_0 & ~i_8_420_1544_0 & ~i_8_420_1702_0 & ~i_8_420_1861_0 & i_8_420_2146_0) | (~i_8_420_658_0 & ~i_8_420_1136_0 & ~i_8_420_1138_0 & ~i_8_420_1559_0 & ~i_8_420_1821_0 & ~i_8_420_1993_0 & ~i_8_420_2003_0 & ~i_8_420_2005_0 & ~i_8_420_2006_0 & ~i_8_420_2263_0))) | (~i_8_420_424_0 & ~i_8_420_923_0 & ~i_8_420_1139_0 & ~i_8_420_1286_0 & ~i_8_420_1985_0 & ~i_8_420_2005_0 & ~i_8_420_2006_0 & ~i_8_420_2200_0))) | (~i_8_420_2260_0 & ((~i_8_420_212_0 & ~i_8_420_662_0 & ~i_8_420_1533_0 & i_8_420_1535_0 & ~i_8_420_1604_0 & i_8_420_1985_0 & ~i_8_420_2005_0) | (~i_8_420_47_0 & ~i_8_420_214_0 & ~i_8_420_1286_0 & ~i_8_420_1558_0 & ~i_8_420_1714_0 & i_8_420_1821_0 & i_8_420_2146_0 & ~i_8_420_2263_0))))) | (~i_8_420_1138_0 & ((~i_8_420_2006_0 & ((~i_8_420_47_0 & ((~i_8_420_34_0 & ~i_8_420_1135_0 & ~i_8_420_1139_0 & ~i_8_420_1711_0 & ~i_8_420_1861_0 & i_8_420_2154_0 & ~i_8_420_2200_0 & ~i_8_420_2227_0) | (~i_8_420_50_0 & i_8_420_662_0 & ~i_8_420_673_0 & ~i_8_420_1233_0 & ~i_8_420_1355_0 & ~i_8_420_1532_0 & ~i_8_420_1881_0 & ~i_8_420_1944_0 & ~i_8_420_2179_0 & ~i_8_420_2261_0 & ~i_8_420_2264_0))) | (~i_8_420_154_0 & ~i_8_420_214_0 & ~i_8_420_1136_0 & ~i_8_420_1272_0 & i_8_420_1354_0 & ~i_8_420_1559_0 & ~i_8_420_2002_0 & ~i_8_420_2153_0 & ~i_8_420_2200_0 & ~i_8_420_2260_0 & ~i_8_420_2261_0))) | (~i_8_420_34_0 & ((~i_8_420_61_0 & ~i_8_420_214_0 & ~i_8_420_1136_0 & ~i_8_420_1276_0 & ~i_8_420_1506_0 & ~i_8_420_1714_0 & i_8_420_1895_0) | (~i_8_420_161_0 & ~i_8_420_658_0 & ~i_8_420_1233_0 & ~i_8_420_1469_0 & i_8_420_1535_0 & ~i_8_420_1559_0 & ~i_8_420_2003_0 & ~i_8_420_2273_0))) | (~i_8_420_161_0 & ((~i_8_420_50_0 & ~i_8_420_335_0 & i_8_420_1233_0 & ~i_8_420_1603_0 & i_8_420_2153_0) | (i_8_420_1533_0 & ~i_8_420_1559_0 & ~i_8_420_1711_0 & ~i_8_420_1719_0 & ~i_8_420_2003_0 & ~i_8_420_2225_0 & ~i_8_420_2261_0))) | (~i_8_420_425_0 & ~i_8_420_1533_0 & ~i_8_420_1993_0 & ~i_8_420_2003_0 & i_8_420_2142_0 & i_8_420_2260_0))) | (~i_8_420_214_0 & ((~i_8_420_34_0 & ((~i_8_420_161_0 & ~i_8_420_1135_0 & ~i_8_420_1351_0 & i_8_420_1354_0 & ~i_8_420_1544_0 & ~i_8_420_1603_0 & ~i_8_420_1604_0 & ~i_8_420_2003_0 & ~i_8_420_2154_0) | (i_8_420_50_0 & ~i_8_420_425_0 & ~i_8_420_923_0 & ~i_8_420_1136_0 & ~i_8_420_1225_0 & ~i_8_420_1354_0 & ~i_8_420_1357_0 & ~i_8_420_1711_0 & ~i_8_420_1985_0 & ~i_8_420_2002_0 & ~i_8_420_2179_0 & ~i_8_420_2260_0))) | (~i_8_420_1139_0 & ((~i_8_420_658_0 & i_8_420_749_0 & ~i_8_420_1469_0 & ~i_8_420_2003_0 & ~i_8_420_2142_0 & ~i_8_420_2200_0) | (~i_8_420_61_0 & i_8_420_1355_0 & ~i_8_420_1558_0 & ~i_8_420_1559_0 & ~i_8_420_2002_0 & ~i_8_420_2006_0 & ~i_8_420_2210_0 & ~i_8_420_2263_0))) | (~i_8_420_2261_0 & ((i_8_420_1355_0 & ~i_8_420_2005_0 & ((~i_8_420_1027_0 & ~i_8_420_1486_0 & ~i_8_420_1559_0 & ~i_8_420_1603_0 & ~i_8_420_1711_0 & ~i_8_420_1715_0 & ~i_8_420_2154_0 & ~i_8_420_2210_0 & ~i_8_420_2227_0) | (~i_8_420_1604_0 & ~i_8_420_2153_0 & i_8_420_2246_0 & ~i_8_420_2260_0))) | (~i_8_420_923_0 & ~i_8_420_1355_0 & i_8_420_1506_0 & ~i_8_420_2246_0 & ~i_8_420_2260_0))) | (~i_8_420_1558_0 & ((~i_8_420_2006_0 & ((i_8_420_1233_0 & ~i_8_420_1604_0 & ~i_8_420_1714_0 & ~i_8_420_1985_0) | (~i_8_420_211_0 & ~i_8_420_335_0 & ~i_8_420_1136_0 & ~i_8_420_1711_0 & i_8_420_2129_0 & ~i_8_420_2225_0 & ~i_8_420_2263_0 & ~i_8_420_2264_0))) | (~i_8_420_212_0 & i_8_420_1719_0 & ~i_8_420_2200_0 & ~i_8_420_2263_0))) | (~i_8_420_955_0 & i_8_420_1272_0 & ~i_8_420_1821_0 & ~i_8_420_2053_0 & ~i_8_420_2179_0))) | (~i_8_420_61_0 & ((~i_8_420_47_0 & i_8_420_425_0 & ~i_8_420_1286_0 & ~i_8_420_1559_0 & ~i_8_420_1944_0 & i_8_420_1993_0 & ~i_8_420_2005_0 & ~i_8_420_2261_0) | (~i_8_420_211_0 & ~i_8_420_662_0 & i_8_420_673_0 & ~i_8_420_1233_0 & ~i_8_420_2002_0 & ~i_8_420_2154_0 & ~i_8_420_2263_0))) | (~i_8_420_47_0 & ((~i_8_420_290_0 & ~i_8_420_391_0 & ~i_8_420_662_0 & ~i_8_420_704_0 & ~i_8_420_829_0 & ~i_8_420_1135_0 & ~i_8_420_1225_0 & ~i_8_420_1286_0 & ~i_8_420_1354_0 & ~i_8_420_1604_0 & ~i_8_420_1861_0 & ~i_8_420_1895_0 & ~i_8_420_2005_0 & ~i_8_420_2006_0 & ~i_8_420_2142_0) | (~i_8_420_212_0 & ~i_8_420_425_0 & i_8_420_463_0 & ~i_8_420_2210_0 & ~i_8_420_2263_0 & ~i_8_420_1136_0 & ~i_8_420_2003_0))) | (~i_8_420_211_0 & ~i_8_420_1881_0 & ((~i_8_420_425_0 & i_8_420_1351_0 & ~i_8_420_1559_0 & ~i_8_420_2200_0 & ~i_8_420_2227_0 & ~i_8_420_1603_0 & ~i_8_420_2006_0) | (~i_8_420_424_0 & i_8_420_658_0 & ~i_8_420_1604_0 & ~i_8_420_1702_0 & ~i_8_420_1714_0 & ~i_8_420_1944_0 & i_8_420_2273_0))) | (~i_8_420_2200_0 & ((~i_8_420_212_0 & ((~i_8_420_424_0 & i_8_420_452_0 & ~i_8_420_1351_0 & ~i_8_420_1357_0 & ~i_8_420_1558_0 & ~i_8_420_1559_0 & ~i_8_420_1886_0 & ~i_8_420_2003_0 & ~i_8_420_2006_0 & ~i_8_420_2053_0) | (~i_8_420_1135_0 & i_8_420_1361_0 & ~i_8_420_1711_0 & ~i_8_420_1715_0 & ~i_8_420_2002_0 & ~i_8_420_2179_0))) | (~i_8_420_1276_0 & i_8_420_1354_0 & i_8_420_1506_0 & ~i_8_420_1711_0 & ~i_8_420_2006_0 & ~i_8_420_2264_0))) | (~i_8_420_2002_0 & ~i_8_420_2003_0 & ~i_8_420_2153_0 & ((~i_8_420_1139_0 & ~i_8_420_1225_0 & ~i_8_420_1702_0 & i_8_420_1711_0) | (~i_8_420_658_0 & ~i_8_420_1135_0 & i_8_420_1469_0 & ~i_8_420_2263_0 & ~i_8_420_2264_0 & ~i_8_420_1985_0 & ~i_8_420_2225_0))) | (~i_8_420_2264_0 & ((~i_8_420_2179_0 & ~i_8_420_2225_0 & ~i_8_420_2246_0 & ~i_8_420_2260_0 & i_8_420_2261_0 & i_8_420_2263_0) | (~i_8_420_293_0 & ~i_8_420_424_0 & ~i_8_420_1603_0 & ~i_8_420_1711_0 & ~i_8_420_1715_0 & i_8_420_1720_0 & ~i_8_420_1821_0 & ~i_8_420_2263_0))) | (~i_8_420_425_0 & ~i_8_420_923_0 & ~i_8_420_1286_0 & i_8_420_1357_0 & ~i_8_420_1558_0 & ~i_8_420_1895_0 & ~i_8_420_2005_0 & ~i_8_420_2129_0));
endmodule



// Benchmark "kernel_8_421" written by ABC on Sun Jul 19 10:10:28 2020

module kernel_8_421 ( 
    i_8_421_34_0, i_8_421_76_0, i_8_421_91_0, i_8_421_95_0, i_8_421_154_0,
    i_8_421_234_0, i_8_421_252_0, i_8_421_305_0, i_8_421_334_0,
    i_8_421_337_0, i_8_421_352_0, i_8_421_353_0, i_8_421_365_0,
    i_8_421_371_0, i_8_421_443_0, i_8_421_469_0, i_8_421_492_0,
    i_8_421_496_0, i_8_421_497_0, i_8_421_499_0, i_8_421_526_0,
    i_8_421_527_0, i_8_421_557_0, i_8_421_586_0, i_8_421_589_0,
    i_8_421_602_0, i_8_421_609_0, i_8_421_613_0, i_8_421_614_0,
    i_8_421_631_0, i_8_421_634_0, i_8_421_659_0, i_8_421_691_0,
    i_8_421_703_0, i_8_421_706_0, i_8_421_760_0, i_8_421_775_0,
    i_8_421_799_0, i_8_421_812_0, i_8_421_833_0, i_8_421_836_0,
    i_8_421_841_0, i_8_421_842_0, i_8_421_844_0, i_8_421_866_0,
    i_8_421_896_0, i_8_421_902_0, i_8_421_932_0, i_8_421_946_0,
    i_8_421_947_0, i_8_421_958_0, i_8_421_967_0, i_8_421_982_0,
    i_8_421_1057_0, i_8_421_1058_0, i_8_421_1225_0, i_8_421_1229_0,
    i_8_421_1247_0, i_8_421_1292_0, i_8_421_1318_0, i_8_421_1322_0,
    i_8_421_1349_0, i_8_421_1435_0, i_8_421_1436_0, i_8_421_1468_0,
    i_8_421_1485_0, i_8_421_1525_0, i_8_421_1538_0, i_8_421_1543_0,
    i_8_421_1553_0, i_8_421_1654_0, i_8_421_1655_0, i_8_421_1682_0,
    i_8_421_1723_0, i_8_421_1729_0, i_8_421_1733_0, i_8_421_1753_0,
    i_8_421_1784_0, i_8_421_1786_0, i_8_421_1787_0, i_8_421_1822_0,
    i_8_421_1871_0, i_8_421_1886_0, i_8_421_1972_0, i_8_421_1984_0,
    i_8_421_1992_0, i_8_421_1993_0, i_8_421_2005_0, i_8_421_2044_0,
    i_8_421_2125_0, i_8_421_2143_0, i_8_421_2144_0, i_8_421_2146_0,
    i_8_421_2147_0, i_8_421_2155_0, i_8_421_2200_0, i_8_421_2224_0,
    i_8_421_2245_0, i_8_421_2289_0, i_8_421_2294_0,
    o_8_421_0_0  );
  input  i_8_421_34_0, i_8_421_76_0, i_8_421_91_0, i_8_421_95_0,
    i_8_421_154_0, i_8_421_234_0, i_8_421_252_0, i_8_421_305_0,
    i_8_421_334_0, i_8_421_337_0, i_8_421_352_0, i_8_421_353_0,
    i_8_421_365_0, i_8_421_371_0, i_8_421_443_0, i_8_421_469_0,
    i_8_421_492_0, i_8_421_496_0, i_8_421_497_0, i_8_421_499_0,
    i_8_421_526_0, i_8_421_527_0, i_8_421_557_0, i_8_421_586_0,
    i_8_421_589_0, i_8_421_602_0, i_8_421_609_0, i_8_421_613_0,
    i_8_421_614_0, i_8_421_631_0, i_8_421_634_0, i_8_421_659_0,
    i_8_421_691_0, i_8_421_703_0, i_8_421_706_0, i_8_421_760_0,
    i_8_421_775_0, i_8_421_799_0, i_8_421_812_0, i_8_421_833_0,
    i_8_421_836_0, i_8_421_841_0, i_8_421_842_0, i_8_421_844_0,
    i_8_421_866_0, i_8_421_896_0, i_8_421_902_0, i_8_421_932_0,
    i_8_421_946_0, i_8_421_947_0, i_8_421_958_0, i_8_421_967_0,
    i_8_421_982_0, i_8_421_1057_0, i_8_421_1058_0, i_8_421_1225_0,
    i_8_421_1229_0, i_8_421_1247_0, i_8_421_1292_0, i_8_421_1318_0,
    i_8_421_1322_0, i_8_421_1349_0, i_8_421_1435_0, i_8_421_1436_0,
    i_8_421_1468_0, i_8_421_1485_0, i_8_421_1525_0, i_8_421_1538_0,
    i_8_421_1543_0, i_8_421_1553_0, i_8_421_1654_0, i_8_421_1655_0,
    i_8_421_1682_0, i_8_421_1723_0, i_8_421_1729_0, i_8_421_1733_0,
    i_8_421_1753_0, i_8_421_1784_0, i_8_421_1786_0, i_8_421_1787_0,
    i_8_421_1822_0, i_8_421_1871_0, i_8_421_1886_0, i_8_421_1972_0,
    i_8_421_1984_0, i_8_421_1992_0, i_8_421_1993_0, i_8_421_2005_0,
    i_8_421_2044_0, i_8_421_2125_0, i_8_421_2143_0, i_8_421_2144_0,
    i_8_421_2146_0, i_8_421_2147_0, i_8_421_2155_0, i_8_421_2200_0,
    i_8_421_2224_0, i_8_421_2245_0, i_8_421_2289_0, i_8_421_2294_0;
  output o_8_421_0_0;
  assign o_8_421_0_0 = 0;
endmodule



// Benchmark "kernel_8_422" written by ABC on Sun Jul 19 10:10:29 2020

module kernel_8_422 ( 
    i_8_422_38_0, i_8_422_47_0, i_8_422_55_0, i_8_422_64_0, i_8_422_65_0,
    i_8_422_73_0, i_8_422_77_0, i_8_422_107_0, i_8_422_127_0,
    i_8_422_140_0, i_8_422_236_0, i_8_422_262_0, i_8_422_263_0,
    i_8_422_309_0, i_8_422_312_0, i_8_422_319_0, i_8_422_344_0,
    i_8_422_360_0, i_8_422_371_0, i_8_422_373_0, i_8_422_374_0,
    i_8_422_388_0, i_8_422_389_0, i_8_422_398_0, i_8_422_416_0,
    i_8_422_419_0, i_8_422_424_0, i_8_422_451_0, i_8_422_457_0,
    i_8_422_529_0, i_8_422_533_0, i_8_422_545_0, i_8_422_559_0,
    i_8_422_577_0, i_8_422_580_0, i_8_422_589_0, i_8_422_610_0,
    i_8_422_632_0, i_8_422_693_0, i_8_422_694_0, i_8_422_698_0,
    i_8_422_702_0, i_8_422_721_0, i_8_422_749_0, i_8_422_782_0,
    i_8_422_838_0, i_8_422_866_0, i_8_422_929_0, i_8_422_967_0,
    i_8_422_968_0, i_8_422_973_0, i_8_422_978_0, i_8_422_1081_0,
    i_8_422_1127_0, i_8_422_1153_0, i_8_422_1172_0, i_8_422_1198_0,
    i_8_422_1234_0, i_8_422_1235_0, i_8_422_1279_0, i_8_422_1298_0,
    i_8_422_1315_0, i_8_422_1336_0, i_8_422_1351_0, i_8_422_1366_0,
    i_8_422_1379_0, i_8_422_1398_0, i_8_422_1406_0, i_8_422_1414_0,
    i_8_422_1442_0, i_8_422_1462_0, i_8_422_1468_0, i_8_422_1469_0,
    i_8_422_1487_0, i_8_422_1514_0, i_8_422_1605_0, i_8_422_1669_0,
    i_8_422_1684_0, i_8_422_1685_0, i_8_422_1688_0, i_8_422_1712_0,
    i_8_422_1777_0, i_8_422_1793_0, i_8_422_1801_0, i_8_422_1819_0,
    i_8_422_1820_0, i_8_422_1821_0, i_8_422_1837_0, i_8_422_1883_0,
    i_8_422_1910_0, i_8_422_1936_0, i_8_422_1939_0, i_8_422_1990_0,
    i_8_422_2005_0, i_8_422_2032_0, i_8_422_2059_0, i_8_422_2072_0,
    i_8_422_2189_0, i_8_422_2265_0, i_8_422_2296_0,
    o_8_422_0_0  );
  input  i_8_422_38_0, i_8_422_47_0, i_8_422_55_0, i_8_422_64_0,
    i_8_422_65_0, i_8_422_73_0, i_8_422_77_0, i_8_422_107_0, i_8_422_127_0,
    i_8_422_140_0, i_8_422_236_0, i_8_422_262_0, i_8_422_263_0,
    i_8_422_309_0, i_8_422_312_0, i_8_422_319_0, i_8_422_344_0,
    i_8_422_360_0, i_8_422_371_0, i_8_422_373_0, i_8_422_374_0,
    i_8_422_388_0, i_8_422_389_0, i_8_422_398_0, i_8_422_416_0,
    i_8_422_419_0, i_8_422_424_0, i_8_422_451_0, i_8_422_457_0,
    i_8_422_529_0, i_8_422_533_0, i_8_422_545_0, i_8_422_559_0,
    i_8_422_577_0, i_8_422_580_0, i_8_422_589_0, i_8_422_610_0,
    i_8_422_632_0, i_8_422_693_0, i_8_422_694_0, i_8_422_698_0,
    i_8_422_702_0, i_8_422_721_0, i_8_422_749_0, i_8_422_782_0,
    i_8_422_838_0, i_8_422_866_0, i_8_422_929_0, i_8_422_967_0,
    i_8_422_968_0, i_8_422_973_0, i_8_422_978_0, i_8_422_1081_0,
    i_8_422_1127_0, i_8_422_1153_0, i_8_422_1172_0, i_8_422_1198_0,
    i_8_422_1234_0, i_8_422_1235_0, i_8_422_1279_0, i_8_422_1298_0,
    i_8_422_1315_0, i_8_422_1336_0, i_8_422_1351_0, i_8_422_1366_0,
    i_8_422_1379_0, i_8_422_1398_0, i_8_422_1406_0, i_8_422_1414_0,
    i_8_422_1442_0, i_8_422_1462_0, i_8_422_1468_0, i_8_422_1469_0,
    i_8_422_1487_0, i_8_422_1514_0, i_8_422_1605_0, i_8_422_1669_0,
    i_8_422_1684_0, i_8_422_1685_0, i_8_422_1688_0, i_8_422_1712_0,
    i_8_422_1777_0, i_8_422_1793_0, i_8_422_1801_0, i_8_422_1819_0,
    i_8_422_1820_0, i_8_422_1821_0, i_8_422_1837_0, i_8_422_1883_0,
    i_8_422_1910_0, i_8_422_1936_0, i_8_422_1939_0, i_8_422_1990_0,
    i_8_422_2005_0, i_8_422_2032_0, i_8_422_2059_0, i_8_422_2072_0,
    i_8_422_2189_0, i_8_422_2265_0, i_8_422_2296_0;
  output o_8_422_0_0;
  assign o_8_422_0_0 = 0;
endmodule



// Benchmark "kernel_8_423" written by ABC on Sun Jul 19 10:10:31 2020

module kernel_8_423 ( 
    i_8_423_89_0, i_8_423_166_0, i_8_423_194_0, i_8_423_195_0,
    i_8_423_197_0, i_8_423_260_0, i_8_423_314_0, i_8_423_381_0,
    i_8_423_384_0, i_8_423_385_0, i_8_423_386_0, i_8_423_451_0,
    i_8_423_458_0, i_8_423_485_0, i_8_423_539_0, i_8_423_556_0,
    i_8_423_575_0, i_8_423_598_0, i_8_423_602_0, i_8_423_607_0,
    i_8_423_611_0, i_8_423_619_0, i_8_423_633_0, i_8_423_635_0,
    i_8_423_662_0, i_8_423_670_0, i_8_423_716_0, i_8_423_736_0,
    i_8_423_751_0, i_8_423_754_0, i_8_423_835_0, i_8_423_841_0,
    i_8_423_844_0, i_8_423_863_0, i_8_423_877_0, i_8_423_986_0,
    i_8_423_994_0, i_8_423_1039_0, i_8_423_1040_0, i_8_423_1042_0,
    i_8_423_1043_0, i_8_423_1051_0, i_8_423_1052_0, i_8_423_1074_0,
    i_8_423_1079_0, i_8_423_1106_0, i_8_423_1177_0, i_8_423_1227_0,
    i_8_423_1229_0, i_8_423_1231_0, i_8_423_1236_0, i_8_423_1262_0,
    i_8_423_1263_0, i_8_423_1264_0, i_8_423_1284_0, i_8_423_1294_0,
    i_8_423_1302_0, i_8_423_1402_0, i_8_423_1412_0, i_8_423_1475_0,
    i_8_423_1484_0, i_8_423_1493_0, i_8_423_1528_0, i_8_423_1529_0,
    i_8_423_1561_0, i_8_423_1562_0, i_8_423_1655_0, i_8_423_1663_0,
    i_8_423_1677_0, i_8_423_1679_0, i_8_423_1682_0, i_8_423_1689_0,
    i_8_423_1700_0, i_8_423_1724_0, i_8_423_1727_0, i_8_423_1751_0,
    i_8_423_1752_0, i_8_423_1771_0, i_8_423_1790_0, i_8_423_1807_0,
    i_8_423_1816_0, i_8_423_1825_0, i_8_423_1867_0, i_8_423_1871_0,
    i_8_423_1880_0, i_8_423_1888_0, i_8_423_1889_0, i_8_423_1967_0,
    i_8_423_1995_0, i_8_423_2014_0, i_8_423_2074_0, i_8_423_2075_0,
    i_8_423_2129_0, i_8_423_2132_0, i_8_423_2143_0, i_8_423_2195_0,
    i_8_423_2210_0, i_8_423_2239_0, i_8_423_2248_0, i_8_423_2249_0,
    o_8_423_0_0  );
  input  i_8_423_89_0, i_8_423_166_0, i_8_423_194_0, i_8_423_195_0,
    i_8_423_197_0, i_8_423_260_0, i_8_423_314_0, i_8_423_381_0,
    i_8_423_384_0, i_8_423_385_0, i_8_423_386_0, i_8_423_451_0,
    i_8_423_458_0, i_8_423_485_0, i_8_423_539_0, i_8_423_556_0,
    i_8_423_575_0, i_8_423_598_0, i_8_423_602_0, i_8_423_607_0,
    i_8_423_611_0, i_8_423_619_0, i_8_423_633_0, i_8_423_635_0,
    i_8_423_662_0, i_8_423_670_0, i_8_423_716_0, i_8_423_736_0,
    i_8_423_751_0, i_8_423_754_0, i_8_423_835_0, i_8_423_841_0,
    i_8_423_844_0, i_8_423_863_0, i_8_423_877_0, i_8_423_986_0,
    i_8_423_994_0, i_8_423_1039_0, i_8_423_1040_0, i_8_423_1042_0,
    i_8_423_1043_0, i_8_423_1051_0, i_8_423_1052_0, i_8_423_1074_0,
    i_8_423_1079_0, i_8_423_1106_0, i_8_423_1177_0, i_8_423_1227_0,
    i_8_423_1229_0, i_8_423_1231_0, i_8_423_1236_0, i_8_423_1262_0,
    i_8_423_1263_0, i_8_423_1264_0, i_8_423_1284_0, i_8_423_1294_0,
    i_8_423_1302_0, i_8_423_1402_0, i_8_423_1412_0, i_8_423_1475_0,
    i_8_423_1484_0, i_8_423_1493_0, i_8_423_1528_0, i_8_423_1529_0,
    i_8_423_1561_0, i_8_423_1562_0, i_8_423_1655_0, i_8_423_1663_0,
    i_8_423_1677_0, i_8_423_1679_0, i_8_423_1682_0, i_8_423_1689_0,
    i_8_423_1700_0, i_8_423_1724_0, i_8_423_1727_0, i_8_423_1751_0,
    i_8_423_1752_0, i_8_423_1771_0, i_8_423_1790_0, i_8_423_1807_0,
    i_8_423_1816_0, i_8_423_1825_0, i_8_423_1867_0, i_8_423_1871_0,
    i_8_423_1880_0, i_8_423_1888_0, i_8_423_1889_0, i_8_423_1967_0,
    i_8_423_1995_0, i_8_423_2014_0, i_8_423_2074_0, i_8_423_2075_0,
    i_8_423_2129_0, i_8_423_2132_0, i_8_423_2143_0, i_8_423_2195_0,
    i_8_423_2210_0, i_8_423_2239_0, i_8_423_2248_0, i_8_423_2249_0;
  output o_8_423_0_0;
  assign o_8_423_0_0 = ~((i_8_423_89_0 & ((i_8_423_451_0 & ~i_8_423_1727_0) | (~i_8_423_1051_0 & ~i_8_423_1889_0 & ~i_8_423_2075_0))) | (~i_8_423_1106_0 & ((~i_8_423_197_0 & ((~i_8_423_195_0 & ~i_8_423_575_0 & ~i_8_423_716_0 & ~i_8_423_835_0 & i_8_423_841_0 & ~i_8_423_1562_0 & ~i_8_423_1700_0 & ~i_8_423_1807_0 & ~i_8_423_1888_0 & ~i_8_423_2014_0) | (i_8_423_619_0 & ~i_8_423_1043_0 & ~i_8_423_1529_0 & ~i_8_423_1689_0 & ~i_8_423_2075_0))) | (~i_8_423_1529_0 & ((~i_8_423_598_0 & i_8_423_635_0 & ~i_8_423_1051_0 & ~i_8_423_1484_0) | (i_8_423_197_0 & ~i_8_423_877_0 & ~i_8_423_986_0 & ~i_8_423_1727_0 & ~i_8_423_1771_0) | (~i_8_423_386_0 & ~i_8_423_751_0 & ~i_8_423_994_0 & ~i_8_423_1229_0 & ~i_8_423_1262_0 & ~i_8_423_1528_0 & ~i_8_423_1663_0 & ~i_8_423_1679_0 & ~i_8_423_1724_0 & ~i_8_423_1967_0 & ~i_8_423_2014_0 & ~i_8_423_2129_0))))) | (~i_8_423_575_0 & ((~i_8_423_195_0 & ((~i_8_423_386_0 & ~i_8_423_607_0 & i_8_423_751_0 & ~i_8_423_1039_0 & ~i_8_423_1043_0) | (~i_8_423_539_0 & ~i_8_423_754_0 & ~i_8_423_1042_0 & ~i_8_423_1889_0 & ~i_8_423_2075_0))) | (~i_8_423_485_0 & ((~i_8_423_986_0 & ~i_8_423_1079_0 & i_8_423_1236_0 & ~i_8_423_1663_0 & ~i_8_423_1727_0) | (~i_8_423_598_0 & ~i_8_423_736_0 & ~i_8_423_1039_0 & ~i_8_423_1528_0 & ~i_8_423_1679_0 & i_8_423_1790_0))) | (~i_8_423_716_0 & ~i_8_423_1880_0 & ((~i_8_423_835_0 & ~i_8_423_844_0 & ~i_8_423_1655_0 & ~i_8_423_1679_0 & ~i_8_423_1682_0 & ~i_8_423_1700_0 & ~i_8_423_1771_0) | (~i_8_423_314_0 & i_8_423_386_0 & ~i_8_423_1294_0 & ~i_8_423_1484_0 & ~i_8_423_1528_0 & ~i_8_423_1562_0 & ~i_8_423_2014_0))) | (~i_8_423_1040_0 & ~i_8_423_1663_0 & i_8_423_1682_0 & ~i_8_423_1771_0) | (~i_8_423_89_0 & ~i_8_423_1051_0 & ~i_8_423_1727_0 & i_8_423_1751_0 & ~i_8_423_1825_0))) | (~i_8_423_635_0 & ((~i_8_423_194_0 & ~i_8_423_539_0 & ~i_8_423_736_0 & ~i_8_423_754_0 & ~i_8_423_841_0 & ~i_8_423_1493_0 & ~i_8_423_1677_0) | (~i_8_423_314_0 & i_8_423_1227_0 & ~i_8_423_1679_0 & ~i_8_423_1727_0 & ~i_8_423_2195_0))) | (~i_8_423_194_0 & ((~i_8_423_751_0 & ~i_8_423_986_0 & ~i_8_423_1051_0 & ~i_8_423_1052_0 & ~i_8_423_1529_0 & ~i_8_423_1727_0 & ~i_8_423_1995_0) | (i_8_423_385_0 & ~i_8_423_994_0 & ~i_8_423_1294_0 & ~i_8_423_1484_0 & ~i_8_423_1677_0 & ~i_8_423_1880_0 & ~i_8_423_2195_0))) | (~i_8_423_314_0 & ((~i_8_423_458_0 & ~i_8_423_602_0 & ~i_8_423_751_0 & ~i_8_423_1529_0 & ~i_8_423_1727_0 & ~i_8_423_1752_0 & ~i_8_423_1807_0 & ~i_8_423_1880_0 & ~i_8_423_1995_0 & ~i_8_423_2075_0 & ~i_8_423_2248_0) | (~i_8_423_539_0 & ~i_8_423_611_0 & ~i_8_423_662_0 & ~i_8_423_841_0 & ~i_8_423_1227_0 & ~i_8_423_1888_0 & ~i_8_423_2014_0 & ~i_8_423_2249_0))) | (~i_8_423_1039_0 & ((~i_8_423_751_0 & ~i_8_423_1040_0 & ((~i_8_423_539_0 & i_8_423_611_0 & ~i_8_423_1229_0 & ~i_8_423_1484_0 & ~i_8_423_1880_0) | (~i_8_423_835_0 & ~i_8_423_1700_0 & ~i_8_423_2132_0))) | (~i_8_423_986_0 & ~i_8_423_994_0 & ~i_8_423_1262_0 & ~i_8_423_1493_0 & ~i_8_423_1655_0 & ~i_8_423_1663_0 & ~i_8_423_1700_0 & ~i_8_423_1727_0 & ~i_8_423_1888_0 & ~i_8_423_1967_0))) | (~i_8_423_1689_0 & ((i_8_423_633_0 & ~i_8_423_1727_0 & ~i_8_423_1771_0 & ~i_8_423_2074_0) | (i_8_423_736_0 & ~i_8_423_994_0 & ~i_8_423_1562_0 & ~i_8_423_1679_0 & ~i_8_423_1700_0 & i_8_423_1888_0 & ~i_8_423_2195_0))) | (~i_8_423_1880_0 & ((~i_8_423_1724_0 & ~i_8_423_1727_0 & ((i_8_423_877_0 & i_8_423_1264_0) | (~i_8_423_662_0 & ~i_8_423_841_0 & ~i_8_423_1051_0 & ~i_8_423_1529_0 & ~i_8_423_1751_0 & ~i_8_423_2075_0))) | (~i_8_423_607_0 & ~i_8_423_844_0 & ~i_8_423_1052_0 & i_8_423_1682_0 & ~i_8_423_1889_0))) | (~i_8_423_835_0 & i_8_423_1677_0 & ~i_8_423_1771_0 & ~i_8_423_1995_0) | (i_8_423_260_0 & i_8_423_458_0 & ~i_8_423_2129_0));
endmodule



// Benchmark "kernel_8_424" written by ABC on Sun Jul 19 10:10:32 2020

module kernel_8_424 ( 
    i_8_424_36_0, i_8_424_41_0, i_8_424_67_0, i_8_424_72_0, i_8_424_73_0,
    i_8_424_74_0, i_8_424_76_0, i_8_424_104_0, i_8_424_136_0,
    i_8_424_173_0, i_8_424_220_0, i_8_424_244_0, i_8_424_304_0,
    i_8_424_352_0, i_8_424_353_0, i_8_424_356_0, i_8_424_361_0,
    i_8_424_365_0, i_8_424_389_0, i_8_424_426_0, i_8_424_427_0,
    i_8_424_470_0, i_8_424_490_0, i_8_424_505_0, i_8_424_514_0,
    i_8_424_515_0, i_8_424_526_0, i_8_424_527_0, i_8_424_569_0,
    i_8_424_582_0, i_8_424_587_0, i_8_424_596_0, i_8_424_603_0,
    i_8_424_611_0, i_8_424_623_0, i_8_424_676_0, i_8_424_679_0,
    i_8_424_748_0, i_8_424_757_0, i_8_424_793_0, i_8_424_826_0,
    i_8_424_829_0, i_8_424_847_0, i_8_424_866_0, i_8_424_911_0,
    i_8_424_1127_0, i_8_424_1161_0, i_8_424_1172_0, i_8_424_1199_0,
    i_8_424_1250_0, i_8_424_1316_0, i_8_424_1378_0, i_8_424_1397_0,
    i_8_424_1404_0, i_8_424_1468_0, i_8_424_1495_0, i_8_424_1531_0,
    i_8_424_1533_0, i_8_424_1534_0, i_8_424_1537_0, i_8_424_1538_0,
    i_8_424_1595_0, i_8_424_1639_0, i_8_424_1648_0, i_8_424_1657_0,
    i_8_424_1682_0, i_8_424_1694_0, i_8_424_1701_0, i_8_424_1706_0,
    i_8_424_1743_0, i_8_424_1754_0, i_8_424_1764_0, i_8_424_1802_0,
    i_8_424_1810_0, i_8_424_1838_0, i_8_424_1843_0, i_8_424_1846_0,
    i_8_424_1886_0, i_8_424_1909_0, i_8_424_1910_0, i_8_424_1948_0,
    i_8_424_1970_0, i_8_424_1972_0, i_8_424_1991_0, i_8_424_2063_0,
    i_8_424_2064_0, i_8_424_2093_0, i_8_424_2142_0, i_8_424_2144_0,
    i_8_424_2147_0, i_8_424_2150_0, i_8_424_2206_0, i_8_424_2242_0,
    i_8_424_2254_0, i_8_424_2255_0, i_8_424_2256_0, i_8_424_2273_0,
    i_8_424_2282_0, i_8_424_2293_0, i_8_424_2296_0,
    o_8_424_0_0  );
  input  i_8_424_36_0, i_8_424_41_0, i_8_424_67_0, i_8_424_72_0,
    i_8_424_73_0, i_8_424_74_0, i_8_424_76_0, i_8_424_104_0, i_8_424_136_0,
    i_8_424_173_0, i_8_424_220_0, i_8_424_244_0, i_8_424_304_0,
    i_8_424_352_0, i_8_424_353_0, i_8_424_356_0, i_8_424_361_0,
    i_8_424_365_0, i_8_424_389_0, i_8_424_426_0, i_8_424_427_0,
    i_8_424_470_0, i_8_424_490_0, i_8_424_505_0, i_8_424_514_0,
    i_8_424_515_0, i_8_424_526_0, i_8_424_527_0, i_8_424_569_0,
    i_8_424_582_0, i_8_424_587_0, i_8_424_596_0, i_8_424_603_0,
    i_8_424_611_0, i_8_424_623_0, i_8_424_676_0, i_8_424_679_0,
    i_8_424_748_0, i_8_424_757_0, i_8_424_793_0, i_8_424_826_0,
    i_8_424_829_0, i_8_424_847_0, i_8_424_866_0, i_8_424_911_0,
    i_8_424_1127_0, i_8_424_1161_0, i_8_424_1172_0, i_8_424_1199_0,
    i_8_424_1250_0, i_8_424_1316_0, i_8_424_1378_0, i_8_424_1397_0,
    i_8_424_1404_0, i_8_424_1468_0, i_8_424_1495_0, i_8_424_1531_0,
    i_8_424_1533_0, i_8_424_1534_0, i_8_424_1537_0, i_8_424_1538_0,
    i_8_424_1595_0, i_8_424_1639_0, i_8_424_1648_0, i_8_424_1657_0,
    i_8_424_1682_0, i_8_424_1694_0, i_8_424_1701_0, i_8_424_1706_0,
    i_8_424_1743_0, i_8_424_1754_0, i_8_424_1764_0, i_8_424_1802_0,
    i_8_424_1810_0, i_8_424_1838_0, i_8_424_1843_0, i_8_424_1846_0,
    i_8_424_1886_0, i_8_424_1909_0, i_8_424_1910_0, i_8_424_1948_0,
    i_8_424_1970_0, i_8_424_1972_0, i_8_424_1991_0, i_8_424_2063_0,
    i_8_424_2064_0, i_8_424_2093_0, i_8_424_2142_0, i_8_424_2144_0,
    i_8_424_2147_0, i_8_424_2150_0, i_8_424_2206_0, i_8_424_2242_0,
    i_8_424_2254_0, i_8_424_2255_0, i_8_424_2256_0, i_8_424_2273_0,
    i_8_424_2282_0, i_8_424_2293_0, i_8_424_2296_0;
  output o_8_424_0_0;
  assign o_8_424_0_0 = 0;
endmodule



// Benchmark "kernel_8_425" written by ABC on Sun Jul 19 10:10:32 2020

module kernel_8_425 ( 
    i_8_425_7_0, i_8_425_8_0, i_8_425_11_0, i_8_425_76_0, i_8_425_79_0,
    i_8_425_89_0, i_8_425_121_0, i_8_425_169_0, i_8_425_227_0,
    i_8_425_269_0, i_8_425_296_0, i_8_425_322_0, i_8_425_332_0,
    i_8_425_364_0, i_8_425_365_0, i_8_425_366_0, i_8_425_368_0,
    i_8_425_379_0, i_8_425_383_0, i_8_425_421_0, i_8_425_429_0,
    i_8_425_448_0, i_8_425_455_0, i_8_425_484_0, i_8_425_491_0,
    i_8_425_492_0, i_8_425_493_0, i_8_425_599_0, i_8_425_605_0,
    i_8_425_629_0, i_8_425_647_0, i_8_425_658_0, i_8_425_661_0,
    i_8_425_664_0, i_8_425_670_0, i_8_425_683_0, i_8_425_696_0,
    i_8_425_698_0, i_8_425_719_0, i_8_425_727_0, i_8_425_748_0,
    i_8_425_771_0, i_8_425_815_0, i_8_425_818_0, i_8_425_827_0,
    i_8_425_893_0, i_8_425_977_0, i_8_425_996_0, i_8_425_998_0,
    i_8_425_1025_0, i_8_425_1078_0, i_8_425_1126_0, i_8_425_1127_0,
    i_8_425_1186_0, i_8_425_1214_0, i_8_425_1241_0, i_8_425_1294_0,
    i_8_425_1301_0, i_8_425_1309_0, i_8_425_1318_0, i_8_425_1325_0,
    i_8_425_1358_0, i_8_425_1366_0, i_8_425_1388_0, i_8_425_1391_0,
    i_8_425_1394_0, i_8_425_1410_0, i_8_425_1411_0, i_8_425_1430_0,
    i_8_425_1591_0, i_8_425_1627_0, i_8_425_1628_0, i_8_425_1649_0,
    i_8_425_1655_0, i_8_425_1675_0, i_8_425_1679_0, i_8_425_1689_0,
    i_8_425_1699_0, i_8_425_1771_0, i_8_425_1779_0, i_8_425_1784_0,
    i_8_425_1807_0, i_8_425_1852_0, i_8_425_1862_0, i_8_425_1907_0,
    i_8_425_1954_0, i_8_425_1988_0, i_8_425_2032_0, i_8_425_2060_0,
    i_8_425_2089_0, i_8_425_2092_0, i_8_425_2122_0, i_8_425_2146_0,
    i_8_425_2149_0, i_8_425_2152_0, i_8_425_2153_0, i_8_425_2175_0,
    i_8_425_2180_0, i_8_425_2195_0, i_8_425_2219_0,
    o_8_425_0_0  );
  input  i_8_425_7_0, i_8_425_8_0, i_8_425_11_0, i_8_425_76_0,
    i_8_425_79_0, i_8_425_89_0, i_8_425_121_0, i_8_425_169_0,
    i_8_425_227_0, i_8_425_269_0, i_8_425_296_0, i_8_425_322_0,
    i_8_425_332_0, i_8_425_364_0, i_8_425_365_0, i_8_425_366_0,
    i_8_425_368_0, i_8_425_379_0, i_8_425_383_0, i_8_425_421_0,
    i_8_425_429_0, i_8_425_448_0, i_8_425_455_0, i_8_425_484_0,
    i_8_425_491_0, i_8_425_492_0, i_8_425_493_0, i_8_425_599_0,
    i_8_425_605_0, i_8_425_629_0, i_8_425_647_0, i_8_425_658_0,
    i_8_425_661_0, i_8_425_664_0, i_8_425_670_0, i_8_425_683_0,
    i_8_425_696_0, i_8_425_698_0, i_8_425_719_0, i_8_425_727_0,
    i_8_425_748_0, i_8_425_771_0, i_8_425_815_0, i_8_425_818_0,
    i_8_425_827_0, i_8_425_893_0, i_8_425_977_0, i_8_425_996_0,
    i_8_425_998_0, i_8_425_1025_0, i_8_425_1078_0, i_8_425_1126_0,
    i_8_425_1127_0, i_8_425_1186_0, i_8_425_1214_0, i_8_425_1241_0,
    i_8_425_1294_0, i_8_425_1301_0, i_8_425_1309_0, i_8_425_1318_0,
    i_8_425_1325_0, i_8_425_1358_0, i_8_425_1366_0, i_8_425_1388_0,
    i_8_425_1391_0, i_8_425_1394_0, i_8_425_1410_0, i_8_425_1411_0,
    i_8_425_1430_0, i_8_425_1591_0, i_8_425_1627_0, i_8_425_1628_0,
    i_8_425_1649_0, i_8_425_1655_0, i_8_425_1675_0, i_8_425_1679_0,
    i_8_425_1689_0, i_8_425_1699_0, i_8_425_1771_0, i_8_425_1779_0,
    i_8_425_1784_0, i_8_425_1807_0, i_8_425_1852_0, i_8_425_1862_0,
    i_8_425_1907_0, i_8_425_1954_0, i_8_425_1988_0, i_8_425_2032_0,
    i_8_425_2060_0, i_8_425_2089_0, i_8_425_2092_0, i_8_425_2122_0,
    i_8_425_2146_0, i_8_425_2149_0, i_8_425_2152_0, i_8_425_2153_0,
    i_8_425_2175_0, i_8_425_2180_0, i_8_425_2195_0, i_8_425_2219_0;
  output o_8_425_0_0;
  assign o_8_425_0_0 = 0;
endmodule



// Benchmark "kernel_8_426" written by ABC on Sun Jul 19 10:10:33 2020

module kernel_8_426 ( 
    i_8_426_21_0, i_8_426_48_0, i_8_426_78_0, i_8_426_106_0, i_8_426_114_0,
    i_8_426_115_0, i_8_426_143_0, i_8_426_157_0, i_8_426_190_0,
    i_8_426_265_0, i_8_426_288_0, i_8_426_366_0, i_8_426_381_0,
    i_8_426_400_0, i_8_426_452_0, i_8_426_454_0, i_8_426_469_0,
    i_8_426_508_0, i_8_426_527_0, i_8_426_550_0, i_8_426_554_0,
    i_8_426_557_0, i_8_426_579_0, i_8_426_581_0, i_8_426_583_0,
    i_8_426_584_0, i_8_426_601_0, i_8_426_633_0, i_8_426_634_0,
    i_8_426_642_0, i_8_426_643_0, i_8_426_653_0, i_8_426_660_0,
    i_8_426_662_0, i_8_426_679_0, i_8_426_680_0, i_8_426_683_0,
    i_8_426_702_0, i_8_426_710_0, i_8_426_720_0, i_8_426_751_0,
    i_8_426_754_0, i_8_426_819_0, i_8_426_826_0, i_8_426_827_0,
    i_8_426_851_0, i_8_426_868_0, i_8_426_895_0, i_8_426_940_0,
    i_8_426_961_0, i_8_426_971_0, i_8_426_993_0, i_8_426_1013_0,
    i_8_426_1039_0, i_8_426_1041_0, i_8_426_1115_0, i_8_426_1137_0,
    i_8_426_1146_0, i_8_426_1149_0, i_8_426_1198_0, i_8_426_1229_0,
    i_8_426_1236_0, i_8_426_1263_0, i_8_426_1267_0, i_8_426_1295_0,
    i_8_426_1300_0, i_8_426_1398_0, i_8_426_1431_0, i_8_426_1435_0,
    i_8_426_1436_0, i_8_426_1437_0, i_8_426_1463_0, i_8_426_1465_0,
    i_8_426_1470_0, i_8_426_1489_0, i_8_426_1491_0, i_8_426_1560_0,
    i_8_426_1679_0, i_8_426_1702_0, i_8_426_1750_0, i_8_426_1759_0,
    i_8_426_1767_0, i_8_426_1769_0, i_8_426_1774_0, i_8_426_1783_0,
    i_8_426_1795_0, i_8_426_1829_0, i_8_426_1837_0, i_8_426_1939_0,
    i_8_426_1947_0, i_8_426_1957_0, i_8_426_1983_0, i_8_426_2036_0,
    i_8_426_2055_0, i_8_426_2110_0, i_8_426_2134_0, i_8_426_2226_0,
    i_8_426_2235_0, i_8_426_2246_0, i_8_426_2263_0,
    o_8_426_0_0  );
  input  i_8_426_21_0, i_8_426_48_0, i_8_426_78_0, i_8_426_106_0,
    i_8_426_114_0, i_8_426_115_0, i_8_426_143_0, i_8_426_157_0,
    i_8_426_190_0, i_8_426_265_0, i_8_426_288_0, i_8_426_366_0,
    i_8_426_381_0, i_8_426_400_0, i_8_426_452_0, i_8_426_454_0,
    i_8_426_469_0, i_8_426_508_0, i_8_426_527_0, i_8_426_550_0,
    i_8_426_554_0, i_8_426_557_0, i_8_426_579_0, i_8_426_581_0,
    i_8_426_583_0, i_8_426_584_0, i_8_426_601_0, i_8_426_633_0,
    i_8_426_634_0, i_8_426_642_0, i_8_426_643_0, i_8_426_653_0,
    i_8_426_660_0, i_8_426_662_0, i_8_426_679_0, i_8_426_680_0,
    i_8_426_683_0, i_8_426_702_0, i_8_426_710_0, i_8_426_720_0,
    i_8_426_751_0, i_8_426_754_0, i_8_426_819_0, i_8_426_826_0,
    i_8_426_827_0, i_8_426_851_0, i_8_426_868_0, i_8_426_895_0,
    i_8_426_940_0, i_8_426_961_0, i_8_426_971_0, i_8_426_993_0,
    i_8_426_1013_0, i_8_426_1039_0, i_8_426_1041_0, i_8_426_1115_0,
    i_8_426_1137_0, i_8_426_1146_0, i_8_426_1149_0, i_8_426_1198_0,
    i_8_426_1229_0, i_8_426_1236_0, i_8_426_1263_0, i_8_426_1267_0,
    i_8_426_1295_0, i_8_426_1300_0, i_8_426_1398_0, i_8_426_1431_0,
    i_8_426_1435_0, i_8_426_1436_0, i_8_426_1437_0, i_8_426_1463_0,
    i_8_426_1465_0, i_8_426_1470_0, i_8_426_1489_0, i_8_426_1491_0,
    i_8_426_1560_0, i_8_426_1679_0, i_8_426_1702_0, i_8_426_1750_0,
    i_8_426_1759_0, i_8_426_1767_0, i_8_426_1769_0, i_8_426_1774_0,
    i_8_426_1783_0, i_8_426_1795_0, i_8_426_1829_0, i_8_426_1837_0,
    i_8_426_1939_0, i_8_426_1947_0, i_8_426_1957_0, i_8_426_1983_0,
    i_8_426_2036_0, i_8_426_2055_0, i_8_426_2110_0, i_8_426_2134_0,
    i_8_426_2226_0, i_8_426_2235_0, i_8_426_2246_0, i_8_426_2263_0;
  output o_8_426_0_0;
  assign o_8_426_0_0 = 0;
endmodule



// Benchmark "kernel_8_427" written by ABC on Sun Jul 19 10:10:34 2020

module kernel_8_427 ( 
    i_8_427_8_0, i_8_427_29_0, i_8_427_34_0, i_8_427_44_0, i_8_427_94_0,
    i_8_427_115_0, i_8_427_130_0, i_8_427_190_0, i_8_427_194_0,
    i_8_427_203_0, i_8_427_206_0, i_8_427_230_0, i_8_427_247_0,
    i_8_427_259_0, i_8_427_262_0, i_8_427_275_0, i_8_427_278_0,
    i_8_427_292_0, i_8_427_311_0, i_8_427_325_0, i_8_427_429_0,
    i_8_427_430_0, i_8_427_445_0, i_8_427_453_0, i_8_427_454_0,
    i_8_427_462_0, i_8_427_475_0, i_8_427_528_0, i_8_427_552_0,
    i_8_427_588_0, i_8_427_607_0, i_8_427_608_0, i_8_427_661_0,
    i_8_427_664_0, i_8_427_673_0, i_8_427_681_0, i_8_427_704_0,
    i_8_427_761_0, i_8_427_792_0, i_8_427_844_0, i_8_427_959_0,
    i_8_427_968_0, i_8_427_972_0, i_8_427_1087_0, i_8_427_1102_0,
    i_8_427_1112_0, i_8_427_1131_0, i_8_427_1132_0, i_8_427_1134_0,
    i_8_427_1159_0, i_8_427_1175_0, i_8_427_1231_0, i_8_427_1274_0,
    i_8_427_1312_0, i_8_427_1346_0, i_8_427_1370_0, i_8_427_1383_0,
    i_8_427_1385_0, i_8_427_1392_0, i_8_427_1407_0, i_8_427_1426_0,
    i_8_427_1482_0, i_8_427_1498_0, i_8_427_1534_0, i_8_427_1537_0,
    i_8_427_1553_0, i_8_427_1597_0, i_8_427_1598_0, i_8_427_1601_0,
    i_8_427_1615_0, i_8_427_1642_0, i_8_427_1645_0, i_8_427_1687_0,
    i_8_427_1748_0, i_8_427_1769_0, i_8_427_1770_0, i_8_427_1777_0,
    i_8_427_1779_0, i_8_427_1836_0, i_8_427_1842_0, i_8_427_1849_0,
    i_8_427_1852_0, i_8_427_1873_0, i_8_427_1877_0, i_8_427_1886_0,
    i_8_427_1887_0, i_8_427_1894_0, i_8_427_1919_0, i_8_427_1969_0,
    i_8_427_1983_0, i_8_427_1985_0, i_8_427_2024_0, i_8_427_2069_0,
    i_8_427_2084_0, i_8_427_2174_0, i_8_427_2177_0, i_8_427_2183_0,
    i_8_427_2191_0, i_8_427_2258_0, i_8_427_2275_0,
    o_8_427_0_0  );
  input  i_8_427_8_0, i_8_427_29_0, i_8_427_34_0, i_8_427_44_0,
    i_8_427_94_0, i_8_427_115_0, i_8_427_130_0, i_8_427_190_0,
    i_8_427_194_0, i_8_427_203_0, i_8_427_206_0, i_8_427_230_0,
    i_8_427_247_0, i_8_427_259_0, i_8_427_262_0, i_8_427_275_0,
    i_8_427_278_0, i_8_427_292_0, i_8_427_311_0, i_8_427_325_0,
    i_8_427_429_0, i_8_427_430_0, i_8_427_445_0, i_8_427_453_0,
    i_8_427_454_0, i_8_427_462_0, i_8_427_475_0, i_8_427_528_0,
    i_8_427_552_0, i_8_427_588_0, i_8_427_607_0, i_8_427_608_0,
    i_8_427_661_0, i_8_427_664_0, i_8_427_673_0, i_8_427_681_0,
    i_8_427_704_0, i_8_427_761_0, i_8_427_792_0, i_8_427_844_0,
    i_8_427_959_0, i_8_427_968_0, i_8_427_972_0, i_8_427_1087_0,
    i_8_427_1102_0, i_8_427_1112_0, i_8_427_1131_0, i_8_427_1132_0,
    i_8_427_1134_0, i_8_427_1159_0, i_8_427_1175_0, i_8_427_1231_0,
    i_8_427_1274_0, i_8_427_1312_0, i_8_427_1346_0, i_8_427_1370_0,
    i_8_427_1383_0, i_8_427_1385_0, i_8_427_1392_0, i_8_427_1407_0,
    i_8_427_1426_0, i_8_427_1482_0, i_8_427_1498_0, i_8_427_1534_0,
    i_8_427_1537_0, i_8_427_1553_0, i_8_427_1597_0, i_8_427_1598_0,
    i_8_427_1601_0, i_8_427_1615_0, i_8_427_1642_0, i_8_427_1645_0,
    i_8_427_1687_0, i_8_427_1748_0, i_8_427_1769_0, i_8_427_1770_0,
    i_8_427_1777_0, i_8_427_1779_0, i_8_427_1836_0, i_8_427_1842_0,
    i_8_427_1849_0, i_8_427_1852_0, i_8_427_1873_0, i_8_427_1877_0,
    i_8_427_1886_0, i_8_427_1887_0, i_8_427_1894_0, i_8_427_1919_0,
    i_8_427_1969_0, i_8_427_1983_0, i_8_427_1985_0, i_8_427_2024_0,
    i_8_427_2069_0, i_8_427_2084_0, i_8_427_2174_0, i_8_427_2177_0,
    i_8_427_2183_0, i_8_427_2191_0, i_8_427_2258_0, i_8_427_2275_0;
  output o_8_427_0_0;
  assign o_8_427_0_0 = 0;
endmodule



// Benchmark "kernel_8_428" written by ABC on Sun Jul 19 10:10:35 2020

module kernel_8_428 ( 
    i_8_428_20_0, i_8_428_22_0, i_8_428_23_0, i_8_428_24_0, i_8_428_40_0,
    i_8_428_52_0, i_8_428_67_0, i_8_428_91_0, i_8_428_114_0, i_8_428_142_0,
    i_8_428_175_0, i_8_428_193_0, i_8_428_200_0, i_8_428_244_0,
    i_8_428_273_0, i_8_428_274_0, i_8_428_356_0, i_8_428_365_0,
    i_8_428_368_0, i_8_428_382_0, i_8_428_385_0, i_8_428_430_0,
    i_8_428_468_0, i_8_428_469_0, i_8_428_571_0, i_8_428_599_0,
    i_8_428_651_0, i_8_428_703_0, i_8_428_706_0, i_8_428_707_0,
    i_8_428_730_0, i_8_428_751_0, i_8_428_814_0, i_8_428_853_0,
    i_8_428_856_0, i_8_428_883_0, i_8_428_955_0, i_8_428_1053_0,
    i_8_428_1066_0, i_8_428_1102_0, i_8_428_1105_0, i_8_428_1111_0,
    i_8_428_1123_0, i_8_428_1182_0, i_8_428_1228_0, i_8_428_1303_0,
    i_8_428_1343_0, i_8_428_1351_0, i_8_428_1390_0, i_8_428_1391_0,
    i_8_428_1400_0, i_8_428_1414_0, i_8_428_1453_0, i_8_428_1470_0,
    i_8_428_1473_0, i_8_428_1510_0, i_8_428_1542_0, i_8_428_1606_0,
    i_8_428_1633_0, i_8_428_1638_0, i_8_428_1642_0, i_8_428_1650_0,
    i_8_428_1653_0, i_8_428_1687_0, i_8_428_1694_0, i_8_428_1705_0,
    i_8_428_1732_0, i_8_428_1764_0, i_8_428_1771_0, i_8_428_1807_0,
    i_8_428_1808_0, i_8_428_1821_0, i_8_428_1873_0, i_8_428_1881_0,
    i_8_428_1882_0, i_8_428_1906_0, i_8_428_1913_0, i_8_428_1918_0,
    i_8_428_1939_0, i_8_428_1942_0, i_8_428_1949_0, i_8_428_1990_0,
    i_8_428_1991_0, i_8_428_2011_0, i_8_428_2065_0, i_8_428_2088_0,
    i_8_428_2091_0, i_8_428_2112_0, i_8_428_2120_0, i_8_428_2149_0,
    i_8_428_2153_0, i_8_428_2182_0, i_8_428_2183_0, i_8_428_2206_0,
    i_8_428_2207_0, i_8_428_2223_0, i_8_428_2233_0, i_8_428_2244_0,
    i_8_428_2272_0, i_8_428_2302_0,
    o_8_428_0_0  );
  input  i_8_428_20_0, i_8_428_22_0, i_8_428_23_0, i_8_428_24_0,
    i_8_428_40_0, i_8_428_52_0, i_8_428_67_0, i_8_428_91_0, i_8_428_114_0,
    i_8_428_142_0, i_8_428_175_0, i_8_428_193_0, i_8_428_200_0,
    i_8_428_244_0, i_8_428_273_0, i_8_428_274_0, i_8_428_356_0,
    i_8_428_365_0, i_8_428_368_0, i_8_428_382_0, i_8_428_385_0,
    i_8_428_430_0, i_8_428_468_0, i_8_428_469_0, i_8_428_571_0,
    i_8_428_599_0, i_8_428_651_0, i_8_428_703_0, i_8_428_706_0,
    i_8_428_707_0, i_8_428_730_0, i_8_428_751_0, i_8_428_814_0,
    i_8_428_853_0, i_8_428_856_0, i_8_428_883_0, i_8_428_955_0,
    i_8_428_1053_0, i_8_428_1066_0, i_8_428_1102_0, i_8_428_1105_0,
    i_8_428_1111_0, i_8_428_1123_0, i_8_428_1182_0, i_8_428_1228_0,
    i_8_428_1303_0, i_8_428_1343_0, i_8_428_1351_0, i_8_428_1390_0,
    i_8_428_1391_0, i_8_428_1400_0, i_8_428_1414_0, i_8_428_1453_0,
    i_8_428_1470_0, i_8_428_1473_0, i_8_428_1510_0, i_8_428_1542_0,
    i_8_428_1606_0, i_8_428_1633_0, i_8_428_1638_0, i_8_428_1642_0,
    i_8_428_1650_0, i_8_428_1653_0, i_8_428_1687_0, i_8_428_1694_0,
    i_8_428_1705_0, i_8_428_1732_0, i_8_428_1764_0, i_8_428_1771_0,
    i_8_428_1807_0, i_8_428_1808_0, i_8_428_1821_0, i_8_428_1873_0,
    i_8_428_1881_0, i_8_428_1882_0, i_8_428_1906_0, i_8_428_1913_0,
    i_8_428_1918_0, i_8_428_1939_0, i_8_428_1942_0, i_8_428_1949_0,
    i_8_428_1990_0, i_8_428_1991_0, i_8_428_2011_0, i_8_428_2065_0,
    i_8_428_2088_0, i_8_428_2091_0, i_8_428_2112_0, i_8_428_2120_0,
    i_8_428_2149_0, i_8_428_2153_0, i_8_428_2182_0, i_8_428_2183_0,
    i_8_428_2206_0, i_8_428_2207_0, i_8_428_2223_0, i_8_428_2233_0,
    i_8_428_2244_0, i_8_428_2272_0, i_8_428_2302_0;
  output o_8_428_0_0;
  assign o_8_428_0_0 = 0;
endmodule



// Benchmark "kernel_8_429" written by ABC on Sun Jul 19 10:10:36 2020

module kernel_8_429 ( 
    i_8_429_30_0, i_8_429_33_0, i_8_429_34_0, i_8_429_36_0, i_8_429_39_0,
    i_8_429_63_0, i_8_429_75_0, i_8_429_87_0, i_8_429_126_0, i_8_429_172_0,
    i_8_429_175_0, i_8_429_180_0, i_8_429_210_0, i_8_429_220_0,
    i_8_429_227_0, i_8_429_237_0, i_8_429_256_0, i_8_429_301_0,
    i_8_429_306_0, i_8_429_309_0, i_8_429_328_0, i_8_429_336_0,
    i_8_429_351_0, i_8_429_378_0, i_8_429_451_0, i_8_429_472_0,
    i_8_429_489_0, i_8_429_490_0, i_8_429_525_0, i_8_429_550_0,
    i_8_429_579_0, i_8_429_589_0, i_8_429_606_0, i_8_429_607_0,
    i_8_429_610_0, i_8_429_624_0, i_8_429_634_0, i_8_429_660_0,
    i_8_429_664_0, i_8_429_694_0, i_8_429_705_0, i_8_429_760_0,
    i_8_429_768_0, i_8_429_843_0, i_8_429_883_0, i_8_429_886_0,
    i_8_429_921_0, i_8_429_924_0, i_8_429_954_0, i_8_429_967_0,
    i_8_429_970_0, i_8_429_985_0, i_8_429_990_0, i_8_429_1026_0,
    i_8_429_1032_0, i_8_429_1056_0, i_8_429_1089_0, i_8_429_1170_0,
    i_8_429_1188_0, i_8_429_1227_0, i_8_429_1228_0, i_8_429_1233_0,
    i_8_429_1254_0, i_8_429_1275_0, i_8_429_1301_0, i_8_429_1329_0,
    i_8_429_1345_0, i_8_429_1371_0, i_8_429_1380_0, i_8_429_1461_0,
    i_8_429_1541_0, i_8_429_1557_0, i_8_429_1560_0, i_8_429_1638_0,
    i_8_429_1650_0, i_8_429_1671_0, i_8_429_1677_0, i_8_429_1701_0,
    i_8_429_1704_0, i_8_429_1749_0, i_8_429_1751_0, i_8_429_1768_0,
    i_8_429_1774_0, i_8_429_1780_0, i_8_429_1803_0, i_8_429_1827_0,
    i_8_429_1863_0, i_8_429_1888_0, i_8_429_1905_0, i_8_429_1906_0,
    i_8_429_2108_0, i_8_429_2133_0, i_8_429_2154_0, i_8_429_2158_0,
    i_8_429_2163_0, i_8_429_2178_0, i_8_429_2181_0, i_8_429_2245_0,
    i_8_429_2272_0, i_8_429_2289_0,
    o_8_429_0_0  );
  input  i_8_429_30_0, i_8_429_33_0, i_8_429_34_0, i_8_429_36_0,
    i_8_429_39_0, i_8_429_63_0, i_8_429_75_0, i_8_429_87_0, i_8_429_126_0,
    i_8_429_172_0, i_8_429_175_0, i_8_429_180_0, i_8_429_210_0,
    i_8_429_220_0, i_8_429_227_0, i_8_429_237_0, i_8_429_256_0,
    i_8_429_301_0, i_8_429_306_0, i_8_429_309_0, i_8_429_328_0,
    i_8_429_336_0, i_8_429_351_0, i_8_429_378_0, i_8_429_451_0,
    i_8_429_472_0, i_8_429_489_0, i_8_429_490_0, i_8_429_525_0,
    i_8_429_550_0, i_8_429_579_0, i_8_429_589_0, i_8_429_606_0,
    i_8_429_607_0, i_8_429_610_0, i_8_429_624_0, i_8_429_634_0,
    i_8_429_660_0, i_8_429_664_0, i_8_429_694_0, i_8_429_705_0,
    i_8_429_760_0, i_8_429_768_0, i_8_429_843_0, i_8_429_883_0,
    i_8_429_886_0, i_8_429_921_0, i_8_429_924_0, i_8_429_954_0,
    i_8_429_967_0, i_8_429_970_0, i_8_429_985_0, i_8_429_990_0,
    i_8_429_1026_0, i_8_429_1032_0, i_8_429_1056_0, i_8_429_1089_0,
    i_8_429_1170_0, i_8_429_1188_0, i_8_429_1227_0, i_8_429_1228_0,
    i_8_429_1233_0, i_8_429_1254_0, i_8_429_1275_0, i_8_429_1301_0,
    i_8_429_1329_0, i_8_429_1345_0, i_8_429_1371_0, i_8_429_1380_0,
    i_8_429_1461_0, i_8_429_1541_0, i_8_429_1557_0, i_8_429_1560_0,
    i_8_429_1638_0, i_8_429_1650_0, i_8_429_1671_0, i_8_429_1677_0,
    i_8_429_1701_0, i_8_429_1704_0, i_8_429_1749_0, i_8_429_1751_0,
    i_8_429_1768_0, i_8_429_1774_0, i_8_429_1780_0, i_8_429_1803_0,
    i_8_429_1827_0, i_8_429_1863_0, i_8_429_1888_0, i_8_429_1905_0,
    i_8_429_1906_0, i_8_429_2108_0, i_8_429_2133_0, i_8_429_2154_0,
    i_8_429_2158_0, i_8_429_2163_0, i_8_429_2178_0, i_8_429_2181_0,
    i_8_429_2245_0, i_8_429_2272_0, i_8_429_2289_0;
  output o_8_429_0_0;
  assign o_8_429_0_0 = ~((~i_8_429_39_0 & ((~i_8_429_172_0 & ~i_8_429_351_0 & ~i_8_429_705_0 & ~i_8_429_1461_0 & ~i_8_429_1638_0 & ~i_8_429_1751_0 & ~i_8_429_2181_0) | (~i_8_429_63_0 & ~i_8_429_306_0 & ~i_8_429_954_0 & ~i_8_429_1677_0 & ~i_8_429_1701_0 & ~i_8_429_2272_0))) | (~i_8_429_1704_0 & ((~i_8_429_172_0 & ((i_8_429_607_0 & ~i_8_429_1188_0 & ~i_8_429_1371_0) | (~i_8_429_924_0 & ~i_8_429_1827_0 & ~i_8_429_1863_0 & ~i_8_429_2178_0 & ~i_8_429_2181_0 & i_8_429_2272_0 & ~i_8_429_2289_0))) | (~i_8_429_126_0 & ~i_8_429_490_0 & ~i_8_429_607_0 & ~i_8_429_768_0 & ~i_8_429_921_0 & ~i_8_429_1780_0 & ~i_8_429_1888_0 & i_8_429_2181_0))) | (~i_8_429_694_0 & ((~i_8_429_210_0 & ((~i_8_429_306_0 & ~i_8_429_1461_0 & i_8_429_1888_0 & ~i_8_429_2181_0) | (~i_8_429_63_0 & ~i_8_429_301_0 & ~i_8_429_1170_0 & ~i_8_429_1380_0 & ~i_8_429_1560_0 & ~i_8_429_1803_0 & ~i_8_429_2133_0 & ~i_8_429_2245_0))) | (~i_8_429_351_0 & ~i_8_429_579_0 & ~i_8_429_924_0 & ~i_8_429_954_0 & ~i_8_429_1026_0 & ~i_8_429_1275_0 & i_8_429_1560_0 & ~i_8_429_2133_0 & ~i_8_429_2289_0))) | (i_8_429_220_0 & ((~i_8_429_336_0 & ~i_8_429_954_0 & ~i_8_429_1032_0 & ~i_8_429_1557_0 & ~i_8_429_1638_0 & ~i_8_429_2154_0) | (~i_8_429_30_0 & ~i_8_429_63_0 & i_8_429_489_0 & ~i_8_429_1329_0 & ~i_8_429_2133_0 & ~i_8_429_2245_0))) | (~i_8_429_1701_0 & ((~i_8_429_306_0 & ((~i_8_429_351_0 & ~i_8_429_579_0 & ~i_8_429_660_0 & ~i_8_429_954_0 & i_8_429_1774_0) | (~i_8_429_227_0 & i_8_429_489_0 & ~i_8_429_634_0 & ~i_8_429_1380_0 & ~i_8_429_1650_0 & ~i_8_429_2178_0 & ~i_8_429_2245_0))) | (~i_8_429_36_0 & ~i_8_429_579_0 & ~i_8_429_768_0 & ~i_8_429_1371_0 & ~i_8_429_1671_0 & ~i_8_429_1827_0 & ~i_8_429_2181_0))) | (~i_8_429_63_0 & ((~i_8_429_36_0 & ((~i_8_429_75_0 & ~i_8_429_180_0 & ~i_8_429_921_0 & ~i_8_429_954_0 & ~i_8_429_1254_0 & ~i_8_429_1380_0 & ~i_8_429_1638_0) | (~i_8_429_843_0 & ~i_8_429_1228_0 & ~i_8_429_1233_0 & ~i_8_429_1905_0 & ~i_8_429_2181_0))) | (~i_8_429_175_0 & i_8_429_301_0 & ~i_8_429_309_0 & ~i_8_429_351_0 & ~i_8_429_2163_0) | (~i_8_429_610_0 & ~i_8_429_768_0 & ~i_8_429_1056_0 & ~i_8_429_1170_0 & ~i_8_429_1275_0 & ~i_8_429_1560_0 & ~i_8_429_1671_0 & ~i_8_429_1905_0 & ~i_8_429_2178_0))) | (i_8_429_525_0 & ((i_8_429_1026_0 & i_8_429_1032_0) | (~i_8_429_1170_0 & ~i_8_429_1227_0 & i_8_429_1677_0 & i_8_429_1749_0))) | (~i_8_429_1560_0 & ((~i_8_429_378_0 & i_8_429_606_0 & ~i_8_429_921_0 & ~i_8_429_1170_0 & i_8_429_1677_0) | (~i_8_429_705_0 & i_8_429_990_0 & ~i_8_429_1905_0))) | (i_8_429_36_0 & ~i_8_429_336_0 & ~i_8_429_607_0 & ~i_8_429_886_0 & ~i_8_429_1671_0 & i_8_429_1774_0 & ~i_8_429_2163_0 & ~i_8_429_2178_0 & ~i_8_429_2181_0) | (~i_8_429_489_0 & ~i_8_429_1227_0 & ~i_8_429_1557_0 & i_8_429_1751_0 & ~i_8_429_2245_0));
endmodule



// Benchmark "kernel_8_430" written by ABC on Sun Jul 19 10:10:37 2020

module kernel_8_430 ( 
    i_8_430_3_0, i_8_430_28_0, i_8_430_33_0, i_8_430_36_0, i_8_430_57_0,
    i_8_430_94_0, i_8_430_106_0, i_8_430_168_0, i_8_430_224_0,
    i_8_430_259_0, i_8_430_323_0, i_8_430_361_0, i_8_430_390_0,
    i_8_430_470_0, i_8_430_498_0, i_8_430_507_0, i_8_430_523_0,
    i_8_430_582_0, i_8_430_597_0, i_8_430_607_0, i_8_430_642_0,
    i_8_430_651_0, i_8_430_654_0, i_8_430_659_0, i_8_430_678_0,
    i_8_430_681_0, i_8_430_751_0, i_8_430_786_0, i_8_430_845_0,
    i_8_430_861_0, i_8_430_870_0, i_8_430_871_0, i_8_430_885_0,
    i_8_430_940_0, i_8_430_1013_0, i_8_430_1038_0, i_8_430_1039_0,
    i_8_430_1084_0, i_8_430_1111_0, i_8_430_1114_0, i_8_430_1128_0,
    i_8_430_1129_0, i_8_430_1159_0, i_8_430_1182_0, i_8_430_1194_0,
    i_8_430_1258_0, i_8_430_1266_0, i_8_430_1272_0, i_8_430_1317_0,
    i_8_430_1338_0, i_8_430_1395_0, i_8_430_1410_0, i_8_430_1425_0,
    i_8_430_1434_0, i_8_430_1437_0, i_8_430_1438_0, i_8_430_1448_0,
    i_8_430_1464_0, i_8_430_1471_0, i_8_430_1483_0, i_8_430_1489_0,
    i_8_430_1492_0, i_8_430_1515_0, i_8_430_1516_0, i_8_430_1548_0,
    i_8_430_1551_0, i_8_430_1605_0, i_8_430_1623_0, i_8_430_1633_0,
    i_8_430_1683_0, i_8_430_1716_0, i_8_430_1722_0, i_8_430_1752_0,
    i_8_430_1759_0, i_8_430_1768_0, i_8_430_1794_0, i_8_430_1803_0,
    i_8_430_1812_0, i_8_430_1822_0, i_8_430_1824_0, i_8_430_1839_0,
    i_8_430_1840_0, i_8_430_1855_0, i_8_430_1881_0, i_8_430_1888_0,
    i_8_430_1938_0, i_8_430_1947_0, i_8_430_1965_0, i_8_430_1984_0,
    i_8_430_1987_0, i_8_430_2133_0, i_8_430_2147_0, i_8_430_2148_0,
    i_8_430_2154_0, i_8_430_2157_0, i_8_430_2158_0, i_8_430_2229_0,
    i_8_430_2233_0, i_8_430_2246_0, i_8_430_2248_0,
    o_8_430_0_0  );
  input  i_8_430_3_0, i_8_430_28_0, i_8_430_33_0, i_8_430_36_0,
    i_8_430_57_0, i_8_430_94_0, i_8_430_106_0, i_8_430_168_0,
    i_8_430_224_0, i_8_430_259_0, i_8_430_323_0, i_8_430_361_0,
    i_8_430_390_0, i_8_430_470_0, i_8_430_498_0, i_8_430_507_0,
    i_8_430_523_0, i_8_430_582_0, i_8_430_597_0, i_8_430_607_0,
    i_8_430_642_0, i_8_430_651_0, i_8_430_654_0, i_8_430_659_0,
    i_8_430_678_0, i_8_430_681_0, i_8_430_751_0, i_8_430_786_0,
    i_8_430_845_0, i_8_430_861_0, i_8_430_870_0, i_8_430_871_0,
    i_8_430_885_0, i_8_430_940_0, i_8_430_1013_0, i_8_430_1038_0,
    i_8_430_1039_0, i_8_430_1084_0, i_8_430_1111_0, i_8_430_1114_0,
    i_8_430_1128_0, i_8_430_1129_0, i_8_430_1159_0, i_8_430_1182_0,
    i_8_430_1194_0, i_8_430_1258_0, i_8_430_1266_0, i_8_430_1272_0,
    i_8_430_1317_0, i_8_430_1338_0, i_8_430_1395_0, i_8_430_1410_0,
    i_8_430_1425_0, i_8_430_1434_0, i_8_430_1437_0, i_8_430_1438_0,
    i_8_430_1448_0, i_8_430_1464_0, i_8_430_1471_0, i_8_430_1483_0,
    i_8_430_1489_0, i_8_430_1492_0, i_8_430_1515_0, i_8_430_1516_0,
    i_8_430_1548_0, i_8_430_1551_0, i_8_430_1605_0, i_8_430_1623_0,
    i_8_430_1633_0, i_8_430_1683_0, i_8_430_1716_0, i_8_430_1722_0,
    i_8_430_1752_0, i_8_430_1759_0, i_8_430_1768_0, i_8_430_1794_0,
    i_8_430_1803_0, i_8_430_1812_0, i_8_430_1822_0, i_8_430_1824_0,
    i_8_430_1839_0, i_8_430_1840_0, i_8_430_1855_0, i_8_430_1881_0,
    i_8_430_1888_0, i_8_430_1938_0, i_8_430_1947_0, i_8_430_1965_0,
    i_8_430_1984_0, i_8_430_1987_0, i_8_430_2133_0, i_8_430_2147_0,
    i_8_430_2148_0, i_8_430_2154_0, i_8_430_2157_0, i_8_430_2158_0,
    i_8_430_2229_0, i_8_430_2233_0, i_8_430_2246_0, i_8_430_2248_0;
  output o_8_430_0_0;
  assign o_8_430_0_0 = 0;
endmodule



// Benchmark "kernel_8_431" written by ABC on Sun Jul 19 10:10:38 2020

module kernel_8_431 ( 
    i_8_431_115_0, i_8_431_143_0, i_8_431_169_0, i_8_431_191_0,
    i_8_431_260_0, i_8_431_296_0, i_8_431_311_0, i_8_431_316_0,
    i_8_431_395_0, i_8_431_459_0, i_8_431_466_0, i_8_431_467_0,
    i_8_431_484_0, i_8_431_485_0, i_8_431_494_0, i_8_431_511_0,
    i_8_431_520_0, i_8_431_523_0, i_8_431_526_0, i_8_431_527_0,
    i_8_431_528_0, i_8_431_529_0, i_8_431_537_0, i_8_431_557_0,
    i_8_431_664_0, i_8_431_715_0, i_8_431_718_0, i_8_431_719_0,
    i_8_431_763_0, i_8_431_764_0, i_8_431_771_0, i_8_431_772_0,
    i_8_431_782_0, i_8_431_835_0, i_8_431_844_0, i_8_431_869_0,
    i_8_431_915_0, i_8_431_949_0, i_8_431_959_0, i_8_431_967_0,
    i_8_431_1040_0, i_8_431_1050_0, i_8_431_1114_0, i_8_431_1124_0,
    i_8_431_1223_0, i_8_431_1267_0, i_8_431_1277_0, i_8_431_1283_0,
    i_8_431_1308_0, i_8_431_1309_0, i_8_431_1319_0, i_8_431_1328_0,
    i_8_431_1330_0, i_8_431_1331_0, i_8_431_1346_0, i_8_431_1392_0,
    i_8_431_1402_0, i_8_431_1439_0, i_8_431_1447_0, i_8_431_1493_0,
    i_8_431_1501_0, i_8_431_1534_0, i_8_431_1537_0, i_8_431_1538_0,
    i_8_431_1555_0, i_8_431_1600_0, i_8_431_1601_0, i_8_431_1633_0,
    i_8_431_1651_0, i_8_431_1681_0, i_8_431_1682_0, i_8_431_1723_0,
    i_8_431_1732_0, i_8_431_1735_0, i_8_431_1768_0, i_8_431_1771_0,
    i_8_431_1796_0, i_8_431_1799_0, i_8_431_1825_0, i_8_431_1843_0,
    i_8_431_1871_0, i_8_431_1886_0, i_8_431_1916_0, i_8_431_1920_0,
    i_8_431_1921_0, i_8_431_1950_0, i_8_431_1979_0, i_8_431_1995_0,
    i_8_431_2014_0, i_8_431_2015_0, i_8_431_2032_0, i_8_431_2068_0,
    i_8_431_2095_0, i_8_431_2114_0, i_8_431_2122_0, i_8_431_2185_0,
    i_8_431_2218_0, i_8_431_2240_0, i_8_431_2247_0, i_8_431_2302_0,
    o_8_431_0_0  );
  input  i_8_431_115_0, i_8_431_143_0, i_8_431_169_0, i_8_431_191_0,
    i_8_431_260_0, i_8_431_296_0, i_8_431_311_0, i_8_431_316_0,
    i_8_431_395_0, i_8_431_459_0, i_8_431_466_0, i_8_431_467_0,
    i_8_431_484_0, i_8_431_485_0, i_8_431_494_0, i_8_431_511_0,
    i_8_431_520_0, i_8_431_523_0, i_8_431_526_0, i_8_431_527_0,
    i_8_431_528_0, i_8_431_529_0, i_8_431_537_0, i_8_431_557_0,
    i_8_431_664_0, i_8_431_715_0, i_8_431_718_0, i_8_431_719_0,
    i_8_431_763_0, i_8_431_764_0, i_8_431_771_0, i_8_431_772_0,
    i_8_431_782_0, i_8_431_835_0, i_8_431_844_0, i_8_431_869_0,
    i_8_431_915_0, i_8_431_949_0, i_8_431_959_0, i_8_431_967_0,
    i_8_431_1040_0, i_8_431_1050_0, i_8_431_1114_0, i_8_431_1124_0,
    i_8_431_1223_0, i_8_431_1267_0, i_8_431_1277_0, i_8_431_1283_0,
    i_8_431_1308_0, i_8_431_1309_0, i_8_431_1319_0, i_8_431_1328_0,
    i_8_431_1330_0, i_8_431_1331_0, i_8_431_1346_0, i_8_431_1392_0,
    i_8_431_1402_0, i_8_431_1439_0, i_8_431_1447_0, i_8_431_1493_0,
    i_8_431_1501_0, i_8_431_1534_0, i_8_431_1537_0, i_8_431_1538_0,
    i_8_431_1555_0, i_8_431_1600_0, i_8_431_1601_0, i_8_431_1633_0,
    i_8_431_1651_0, i_8_431_1681_0, i_8_431_1682_0, i_8_431_1723_0,
    i_8_431_1732_0, i_8_431_1735_0, i_8_431_1768_0, i_8_431_1771_0,
    i_8_431_1796_0, i_8_431_1799_0, i_8_431_1825_0, i_8_431_1843_0,
    i_8_431_1871_0, i_8_431_1886_0, i_8_431_1916_0, i_8_431_1920_0,
    i_8_431_1921_0, i_8_431_1950_0, i_8_431_1979_0, i_8_431_1995_0,
    i_8_431_2014_0, i_8_431_2015_0, i_8_431_2032_0, i_8_431_2068_0,
    i_8_431_2095_0, i_8_431_2114_0, i_8_431_2122_0, i_8_431_2185_0,
    i_8_431_2218_0, i_8_431_2240_0, i_8_431_2247_0, i_8_431_2302_0;
  output o_8_431_0_0;
  assign o_8_431_0_0 = 0;
endmodule



// Benchmark "kernel_8_432" written by ABC on Sun Jul 19 10:10:39 2020

module kernel_8_432 ( 
    i_8_432_52_0, i_8_432_57_0, i_8_432_84_0, i_8_432_141_0, i_8_432_142_0,
    i_8_432_143_0, i_8_432_192_0, i_8_432_225_0, i_8_432_255_0,
    i_8_432_328_0, i_8_432_370_0, i_8_432_373_0, i_8_432_382_0,
    i_8_432_417_0, i_8_432_480_0, i_8_432_481_0, i_8_432_483_0,
    i_8_432_484_0, i_8_432_500_0, i_8_432_507_0, i_8_432_510_0,
    i_8_432_522_0, i_8_432_526_0, i_8_432_528_0, i_8_432_530_0,
    i_8_432_544_0, i_8_432_596_0, i_8_432_602_0, i_8_432_610_0,
    i_8_432_651_0, i_8_432_656_0, i_8_432_661_0, i_8_432_702_0,
    i_8_432_759_0, i_8_432_760_0, i_8_432_763_0, i_8_432_777_0,
    i_8_432_778_0, i_8_432_789_0, i_8_432_796_0, i_8_432_813_0,
    i_8_432_814_0, i_8_432_836_0, i_8_432_842_0, i_8_432_871_0,
    i_8_432_879_0, i_8_432_904_0, i_8_432_949_0, i_8_432_993_0,
    i_8_432_1011_0, i_8_432_1016_0, i_8_432_1050_0, i_8_432_1074_0,
    i_8_432_1135_0, i_8_432_1177_0, i_8_432_1272_0, i_8_432_1284_0,
    i_8_432_1305_0, i_8_432_1306_0, i_8_432_1344_0, i_8_432_1348_0,
    i_8_432_1349_0, i_8_432_1357_0, i_8_432_1419_0, i_8_432_1437_0,
    i_8_432_1506_0, i_8_432_1527_0, i_8_432_1544_0, i_8_432_1545_0,
    i_8_432_1547_0, i_8_432_1573_0, i_8_432_1630_0, i_8_432_1633_0,
    i_8_432_1644_0, i_8_432_1668_0, i_8_432_1677_0, i_8_432_1679_0,
    i_8_432_1682_0, i_8_432_1710_0, i_8_432_1714_0, i_8_432_1717_0,
    i_8_432_1718_0, i_8_432_1722_0, i_8_432_1726_0, i_8_432_1732_0,
    i_8_432_1753_0, i_8_432_1867_0, i_8_432_1868_0, i_8_432_1906_0,
    i_8_432_1950_0, i_8_432_1997_0, i_8_432_2028_0, i_8_432_2101_0,
    i_8_432_2104_0, i_8_432_2128_0, i_8_432_2130_0, i_8_432_2131_0,
    i_8_432_2214_0, i_8_432_2215_0, i_8_432_2216_0,
    o_8_432_0_0  );
  input  i_8_432_52_0, i_8_432_57_0, i_8_432_84_0, i_8_432_141_0,
    i_8_432_142_0, i_8_432_143_0, i_8_432_192_0, i_8_432_225_0,
    i_8_432_255_0, i_8_432_328_0, i_8_432_370_0, i_8_432_373_0,
    i_8_432_382_0, i_8_432_417_0, i_8_432_480_0, i_8_432_481_0,
    i_8_432_483_0, i_8_432_484_0, i_8_432_500_0, i_8_432_507_0,
    i_8_432_510_0, i_8_432_522_0, i_8_432_526_0, i_8_432_528_0,
    i_8_432_530_0, i_8_432_544_0, i_8_432_596_0, i_8_432_602_0,
    i_8_432_610_0, i_8_432_651_0, i_8_432_656_0, i_8_432_661_0,
    i_8_432_702_0, i_8_432_759_0, i_8_432_760_0, i_8_432_763_0,
    i_8_432_777_0, i_8_432_778_0, i_8_432_789_0, i_8_432_796_0,
    i_8_432_813_0, i_8_432_814_0, i_8_432_836_0, i_8_432_842_0,
    i_8_432_871_0, i_8_432_879_0, i_8_432_904_0, i_8_432_949_0,
    i_8_432_993_0, i_8_432_1011_0, i_8_432_1016_0, i_8_432_1050_0,
    i_8_432_1074_0, i_8_432_1135_0, i_8_432_1177_0, i_8_432_1272_0,
    i_8_432_1284_0, i_8_432_1305_0, i_8_432_1306_0, i_8_432_1344_0,
    i_8_432_1348_0, i_8_432_1349_0, i_8_432_1357_0, i_8_432_1419_0,
    i_8_432_1437_0, i_8_432_1506_0, i_8_432_1527_0, i_8_432_1544_0,
    i_8_432_1545_0, i_8_432_1547_0, i_8_432_1573_0, i_8_432_1630_0,
    i_8_432_1633_0, i_8_432_1644_0, i_8_432_1668_0, i_8_432_1677_0,
    i_8_432_1679_0, i_8_432_1682_0, i_8_432_1710_0, i_8_432_1714_0,
    i_8_432_1717_0, i_8_432_1718_0, i_8_432_1722_0, i_8_432_1726_0,
    i_8_432_1732_0, i_8_432_1753_0, i_8_432_1867_0, i_8_432_1868_0,
    i_8_432_1906_0, i_8_432_1950_0, i_8_432_1997_0, i_8_432_2028_0,
    i_8_432_2101_0, i_8_432_2104_0, i_8_432_2128_0, i_8_432_2130_0,
    i_8_432_2131_0, i_8_432_2214_0, i_8_432_2215_0, i_8_432_2216_0;
  output o_8_432_0_0;
  assign o_8_432_0_0 = 0;
endmodule



// Benchmark "kernel_8_433" written by ABC on Sun Jul 19 10:10:40 2020

module kernel_8_433 ( 
    i_8_433_30_0, i_8_433_49_0, i_8_433_81_0, i_8_433_106_0, i_8_433_138_0,
    i_8_433_141_0, i_8_433_142_0, i_8_433_183_0, i_8_433_255_0,
    i_8_433_256_0, i_8_433_328_0, i_8_433_352_0, i_8_433_355_0,
    i_8_433_374_0, i_8_433_418_0, i_8_433_442_0, i_8_433_445_0,
    i_8_433_450_0, i_8_433_453_0, i_8_433_481_0, i_8_433_494_0,
    i_8_433_497_0, i_8_433_547_0, i_8_433_616_0, i_8_433_663_0,
    i_8_433_691_0, i_8_433_702_0, i_8_433_703_0, i_8_433_706_0,
    i_8_433_736_0, i_8_433_765_0, i_8_433_786_0, i_8_433_811_0,
    i_8_433_814_0, i_8_433_815_0, i_8_433_819_0, i_8_433_828_0,
    i_8_433_848_0, i_8_433_867_0, i_8_433_868_0, i_8_433_869_0,
    i_8_433_895_0, i_8_433_922_0, i_8_433_949_0, i_8_433_950_0,
    i_8_433_953_0, i_8_433_969_0, i_8_433_972_0, i_8_433_973_0,
    i_8_433_976_0, i_8_433_982_0, i_8_433_984_0, i_8_433_994_0,
    i_8_433_1011_0, i_8_433_1027_0, i_8_433_1074_0, i_8_433_1134_0,
    i_8_433_1155_0, i_8_433_1267_0, i_8_433_1273_0, i_8_433_1305_0,
    i_8_433_1325_0, i_8_433_1336_0, i_8_433_1342_0, i_8_433_1442_0,
    i_8_433_1468_0, i_8_433_1525_0, i_8_433_1559_0, i_8_433_1564_0,
    i_8_433_1617_0, i_8_433_1713_0, i_8_433_1714_0, i_8_433_1717_0,
    i_8_433_1726_0, i_8_433_1731_0, i_8_433_1732_0, i_8_433_1750_0,
    i_8_433_1753_0, i_8_433_1754_0, i_8_433_1786_0, i_8_433_1789_0,
    i_8_433_1802_0, i_8_433_1812_0, i_8_433_1813_0, i_8_433_1864_0,
    i_8_433_1903_0, i_8_433_1904_0, i_8_433_1930_0, i_8_433_1952_0,
    i_8_433_2007_0, i_8_433_2010_0, i_8_433_2011_0, i_8_433_2068_0,
    i_8_433_2069_0, i_8_433_2093_0, i_8_433_2131_0, i_8_433_2136_0,
    i_8_433_2214_0, i_8_433_2215_0, i_8_433_2244_0,
    o_8_433_0_0  );
  input  i_8_433_30_0, i_8_433_49_0, i_8_433_81_0, i_8_433_106_0,
    i_8_433_138_0, i_8_433_141_0, i_8_433_142_0, i_8_433_183_0,
    i_8_433_255_0, i_8_433_256_0, i_8_433_328_0, i_8_433_352_0,
    i_8_433_355_0, i_8_433_374_0, i_8_433_418_0, i_8_433_442_0,
    i_8_433_445_0, i_8_433_450_0, i_8_433_453_0, i_8_433_481_0,
    i_8_433_494_0, i_8_433_497_0, i_8_433_547_0, i_8_433_616_0,
    i_8_433_663_0, i_8_433_691_0, i_8_433_702_0, i_8_433_703_0,
    i_8_433_706_0, i_8_433_736_0, i_8_433_765_0, i_8_433_786_0,
    i_8_433_811_0, i_8_433_814_0, i_8_433_815_0, i_8_433_819_0,
    i_8_433_828_0, i_8_433_848_0, i_8_433_867_0, i_8_433_868_0,
    i_8_433_869_0, i_8_433_895_0, i_8_433_922_0, i_8_433_949_0,
    i_8_433_950_0, i_8_433_953_0, i_8_433_969_0, i_8_433_972_0,
    i_8_433_973_0, i_8_433_976_0, i_8_433_982_0, i_8_433_984_0,
    i_8_433_994_0, i_8_433_1011_0, i_8_433_1027_0, i_8_433_1074_0,
    i_8_433_1134_0, i_8_433_1155_0, i_8_433_1267_0, i_8_433_1273_0,
    i_8_433_1305_0, i_8_433_1325_0, i_8_433_1336_0, i_8_433_1342_0,
    i_8_433_1442_0, i_8_433_1468_0, i_8_433_1525_0, i_8_433_1559_0,
    i_8_433_1564_0, i_8_433_1617_0, i_8_433_1713_0, i_8_433_1714_0,
    i_8_433_1717_0, i_8_433_1726_0, i_8_433_1731_0, i_8_433_1732_0,
    i_8_433_1750_0, i_8_433_1753_0, i_8_433_1754_0, i_8_433_1786_0,
    i_8_433_1789_0, i_8_433_1802_0, i_8_433_1812_0, i_8_433_1813_0,
    i_8_433_1864_0, i_8_433_1903_0, i_8_433_1904_0, i_8_433_1930_0,
    i_8_433_1952_0, i_8_433_2007_0, i_8_433_2010_0, i_8_433_2011_0,
    i_8_433_2068_0, i_8_433_2069_0, i_8_433_2093_0, i_8_433_2131_0,
    i_8_433_2136_0, i_8_433_2214_0, i_8_433_2215_0, i_8_433_2244_0;
  output o_8_433_0_0;
  assign o_8_433_0_0 = 0;
endmodule



// Benchmark "kernel_8_434" written by ABC on Sun Jul 19 10:10:41 2020

module kernel_8_434 ( 
    i_8_434_48_0, i_8_434_49_0, i_8_434_66_0, i_8_434_67_0, i_8_434_72_0,
    i_8_434_78_0, i_8_434_93_0, i_8_434_107_0, i_8_434_114_0,
    i_8_434_130_0, i_8_434_138_0, i_8_434_166_0, i_8_434_174_0,
    i_8_434_178_0, i_8_434_183_0, i_8_434_191_0, i_8_434_237_0,
    i_8_434_304_0, i_8_434_321_0, i_8_434_334_0, i_8_434_336_0,
    i_8_434_337_0, i_8_434_361_0, i_8_434_381_0, i_8_434_382_0,
    i_8_434_399_0, i_8_434_400_0, i_8_434_579_0, i_8_434_607_0,
    i_8_434_608_0, i_8_434_642_0, i_8_434_651_0, i_8_434_693_0,
    i_8_434_694_0, i_8_434_705_0, i_8_434_729_0, i_8_434_795_0,
    i_8_434_831_0, i_8_434_864_0, i_8_434_882_0, i_8_434_930_0,
    i_8_434_954_0, i_8_434_969_0, i_8_434_1020_0, i_8_434_1092_0,
    i_8_434_1093_0, i_8_434_1128_0, i_8_434_1255_0, i_8_434_1263_0,
    i_8_434_1287_0, i_8_434_1300_0, i_8_434_1306_0, i_8_434_1311_0,
    i_8_434_1314_0, i_8_434_1317_0, i_8_434_1354_0, i_8_434_1388_0,
    i_8_434_1400_0, i_8_434_1448_0, i_8_434_1469_0, i_8_434_1493_0,
    i_8_434_1524_0, i_8_434_1527_0, i_8_434_1545_0, i_8_434_1560_0,
    i_8_434_1686_0, i_8_434_1687_0, i_8_434_1704_0, i_8_434_1706_0,
    i_8_434_1749_0, i_8_434_1821_0, i_8_434_1825_0, i_8_434_1830_0,
    i_8_434_1840_0, i_8_434_1846_0, i_8_434_1848_0, i_8_434_1851_0,
    i_8_434_1855_0, i_8_434_1869_0, i_8_434_1893_0, i_8_434_1938_0,
    i_8_434_1993_0, i_8_434_1995_0, i_8_434_2038_0, i_8_434_2040_0,
    i_8_434_2041_0, i_8_434_2056_0, i_8_434_2077_0, i_8_434_2145_0,
    i_8_434_2154_0, i_8_434_2155_0, i_8_434_2157_0, i_8_434_2181_0,
    i_8_434_2199_0, i_8_434_2200_0, i_8_434_2202_0, i_8_434_2220_0,
    i_8_434_2246_0, i_8_434_2275_0, i_8_434_2299_0,
    o_8_434_0_0  );
  input  i_8_434_48_0, i_8_434_49_0, i_8_434_66_0, i_8_434_67_0,
    i_8_434_72_0, i_8_434_78_0, i_8_434_93_0, i_8_434_107_0, i_8_434_114_0,
    i_8_434_130_0, i_8_434_138_0, i_8_434_166_0, i_8_434_174_0,
    i_8_434_178_0, i_8_434_183_0, i_8_434_191_0, i_8_434_237_0,
    i_8_434_304_0, i_8_434_321_0, i_8_434_334_0, i_8_434_336_0,
    i_8_434_337_0, i_8_434_361_0, i_8_434_381_0, i_8_434_382_0,
    i_8_434_399_0, i_8_434_400_0, i_8_434_579_0, i_8_434_607_0,
    i_8_434_608_0, i_8_434_642_0, i_8_434_651_0, i_8_434_693_0,
    i_8_434_694_0, i_8_434_705_0, i_8_434_729_0, i_8_434_795_0,
    i_8_434_831_0, i_8_434_864_0, i_8_434_882_0, i_8_434_930_0,
    i_8_434_954_0, i_8_434_969_0, i_8_434_1020_0, i_8_434_1092_0,
    i_8_434_1093_0, i_8_434_1128_0, i_8_434_1255_0, i_8_434_1263_0,
    i_8_434_1287_0, i_8_434_1300_0, i_8_434_1306_0, i_8_434_1311_0,
    i_8_434_1314_0, i_8_434_1317_0, i_8_434_1354_0, i_8_434_1388_0,
    i_8_434_1400_0, i_8_434_1448_0, i_8_434_1469_0, i_8_434_1493_0,
    i_8_434_1524_0, i_8_434_1527_0, i_8_434_1545_0, i_8_434_1560_0,
    i_8_434_1686_0, i_8_434_1687_0, i_8_434_1704_0, i_8_434_1706_0,
    i_8_434_1749_0, i_8_434_1821_0, i_8_434_1825_0, i_8_434_1830_0,
    i_8_434_1840_0, i_8_434_1846_0, i_8_434_1848_0, i_8_434_1851_0,
    i_8_434_1855_0, i_8_434_1869_0, i_8_434_1893_0, i_8_434_1938_0,
    i_8_434_1993_0, i_8_434_1995_0, i_8_434_2038_0, i_8_434_2040_0,
    i_8_434_2041_0, i_8_434_2056_0, i_8_434_2077_0, i_8_434_2145_0,
    i_8_434_2154_0, i_8_434_2155_0, i_8_434_2157_0, i_8_434_2181_0,
    i_8_434_2199_0, i_8_434_2200_0, i_8_434_2202_0, i_8_434_2220_0,
    i_8_434_2246_0, i_8_434_2275_0, i_8_434_2299_0;
  output o_8_434_0_0;
  assign o_8_434_0_0 = 0;
endmodule



// Benchmark "kernel_8_435" written by ABC on Sun Jul 19 10:10:42 2020

module kernel_8_435 ( 
    i_8_435_18_0, i_8_435_31_0, i_8_435_32_0, i_8_435_154_0, i_8_435_208_0,
    i_8_435_220_0, i_8_435_289_0, i_8_435_326_0, i_8_435_370_0,
    i_8_435_371_0, i_8_435_373_0, i_8_435_374_0, i_8_435_426_0,
    i_8_435_445_0, i_8_435_473_0, i_8_435_478_0, i_8_435_485_0,
    i_8_435_496_0, i_8_435_522_0, i_8_435_524_0, i_8_435_578_0,
    i_8_435_586_0, i_8_435_604_0, i_8_435_610_0, i_8_435_611_0,
    i_8_435_625_0, i_8_435_631_0, i_8_435_657_0, i_8_435_667_0,
    i_8_435_668_0, i_8_435_671_0, i_8_435_711_0, i_8_435_712_0,
    i_8_435_713_0, i_8_435_757_0, i_8_435_776_0, i_8_435_783_0,
    i_8_435_787_0, i_8_435_792_0, i_8_435_793_0, i_8_435_821_0,
    i_8_435_855_0, i_8_435_892_0, i_8_435_938_0, i_8_435_947_0,
    i_8_435_1112_0, i_8_435_1127_0, i_8_435_1130_0, i_8_435_1216_0,
    i_8_435_1225_0, i_8_435_1246_0, i_8_435_1247_0, i_8_435_1252_0,
    i_8_435_1260_0, i_8_435_1264_0, i_8_435_1279_0, i_8_435_1280_0,
    i_8_435_1297_0, i_8_435_1317_0, i_8_435_1318_0, i_8_435_1323_0,
    i_8_435_1431_0, i_8_435_1434_0, i_8_435_1450_0, i_8_435_1451_0,
    i_8_435_1503_0, i_8_435_1504_0, i_8_435_1505_0, i_8_435_1522_0,
    i_8_435_1585_0, i_8_435_1586_0, i_8_435_1595_0, i_8_435_1631_0,
    i_8_435_1634_0, i_8_435_1666_0, i_8_435_1681_0, i_8_435_1696_0,
    i_8_435_1713_0, i_8_435_1739_0, i_8_435_1752_0, i_8_435_1753_0,
    i_8_435_1759_0, i_8_435_1776_0, i_8_435_1802_0, i_8_435_1824_0,
    i_8_435_1837_0, i_8_435_1854_0, i_8_435_1856_0, i_8_435_1890_0,
    i_8_435_1891_0, i_8_435_1948_0, i_8_435_1965_0, i_8_435_2047_0,
    i_8_435_2125_0, i_8_435_2126_0, i_8_435_2147_0, i_8_435_2189_0,
    i_8_435_2245_0, i_8_435_2270_0, i_8_435_2286_0,
    o_8_435_0_0  );
  input  i_8_435_18_0, i_8_435_31_0, i_8_435_32_0, i_8_435_154_0,
    i_8_435_208_0, i_8_435_220_0, i_8_435_289_0, i_8_435_326_0,
    i_8_435_370_0, i_8_435_371_0, i_8_435_373_0, i_8_435_374_0,
    i_8_435_426_0, i_8_435_445_0, i_8_435_473_0, i_8_435_478_0,
    i_8_435_485_0, i_8_435_496_0, i_8_435_522_0, i_8_435_524_0,
    i_8_435_578_0, i_8_435_586_0, i_8_435_604_0, i_8_435_610_0,
    i_8_435_611_0, i_8_435_625_0, i_8_435_631_0, i_8_435_657_0,
    i_8_435_667_0, i_8_435_668_0, i_8_435_671_0, i_8_435_711_0,
    i_8_435_712_0, i_8_435_713_0, i_8_435_757_0, i_8_435_776_0,
    i_8_435_783_0, i_8_435_787_0, i_8_435_792_0, i_8_435_793_0,
    i_8_435_821_0, i_8_435_855_0, i_8_435_892_0, i_8_435_938_0,
    i_8_435_947_0, i_8_435_1112_0, i_8_435_1127_0, i_8_435_1130_0,
    i_8_435_1216_0, i_8_435_1225_0, i_8_435_1246_0, i_8_435_1247_0,
    i_8_435_1252_0, i_8_435_1260_0, i_8_435_1264_0, i_8_435_1279_0,
    i_8_435_1280_0, i_8_435_1297_0, i_8_435_1317_0, i_8_435_1318_0,
    i_8_435_1323_0, i_8_435_1431_0, i_8_435_1434_0, i_8_435_1450_0,
    i_8_435_1451_0, i_8_435_1503_0, i_8_435_1504_0, i_8_435_1505_0,
    i_8_435_1522_0, i_8_435_1585_0, i_8_435_1586_0, i_8_435_1595_0,
    i_8_435_1631_0, i_8_435_1634_0, i_8_435_1666_0, i_8_435_1681_0,
    i_8_435_1696_0, i_8_435_1713_0, i_8_435_1739_0, i_8_435_1752_0,
    i_8_435_1753_0, i_8_435_1759_0, i_8_435_1776_0, i_8_435_1802_0,
    i_8_435_1824_0, i_8_435_1837_0, i_8_435_1854_0, i_8_435_1856_0,
    i_8_435_1890_0, i_8_435_1891_0, i_8_435_1948_0, i_8_435_1965_0,
    i_8_435_2047_0, i_8_435_2125_0, i_8_435_2126_0, i_8_435_2147_0,
    i_8_435_2189_0, i_8_435_2245_0, i_8_435_2270_0, i_8_435_2286_0;
  output o_8_435_0_0;
  assign o_8_435_0_0 = 0;
endmodule



// Benchmark "kernel_8_436" written by ABC on Sun Jul 19 10:10:43 2020

module kernel_8_436 ( 
    i_8_436_18_0, i_8_436_48_0, i_8_436_78_0, i_8_436_117_0, i_8_436_141_0,
    i_8_436_142_0, i_8_436_219_0, i_8_436_259_0, i_8_436_310_0,
    i_8_436_322_0, i_8_436_336_0, i_8_436_345_0, i_8_436_346_0,
    i_8_436_348_0, i_8_436_360_0, i_8_436_363_0, i_8_436_367_0,
    i_8_436_378_0, i_8_436_381_0, i_8_436_400_0, i_8_436_402_0,
    i_8_436_417_0, i_8_436_427_0, i_8_436_454_0, i_8_436_493_0,
    i_8_436_499_0, i_8_436_579_0, i_8_436_603_0, i_8_436_615_0,
    i_8_436_643_0, i_8_436_654_0, i_8_436_658_0, i_8_436_660_0,
    i_8_436_675_0, i_8_436_696_0, i_8_436_702_0, i_8_436_750_0,
    i_8_436_795_0, i_8_436_799_0, i_8_436_849_0, i_8_436_873_0,
    i_8_436_889_0, i_8_436_991_0, i_8_436_1020_0, i_8_436_1056_0,
    i_8_436_1059_0, i_8_436_1092_0, i_8_436_1104_0, i_8_436_1115_0,
    i_8_436_1146_0, i_8_436_1152_0, i_8_436_1158_0, i_8_436_1266_0,
    i_8_436_1283_0, i_8_436_1284_0, i_8_436_1291_0, i_8_436_1314_0,
    i_8_436_1323_0, i_8_436_1383_0, i_8_436_1426_0, i_8_436_1439_0,
    i_8_436_1440_0, i_8_436_1444_0, i_8_436_1473_0, i_8_436_1597_0,
    i_8_436_1602_0, i_8_436_1633_0, i_8_436_1644_0, i_8_436_1671_0,
    i_8_436_1688_0, i_8_436_1699_0, i_8_436_1702_0, i_8_436_1704_0,
    i_8_436_1723_0, i_8_436_1749_0, i_8_436_1753_0, i_8_436_1803_0,
    i_8_436_1818_0, i_8_436_1830_0, i_8_436_1836_0, i_8_436_1840_0,
    i_8_436_1857_0, i_8_436_1885_0, i_8_436_1887_0, i_8_436_1899_0,
    i_8_436_1944_0, i_8_436_1947_0, i_8_436_1980_0, i_8_436_1981_0,
    i_8_436_2004_0, i_8_436_2184_0, i_8_436_2223_0, i_8_436_2227_0,
    i_8_436_2229_0, i_8_436_2238_0, i_8_436_2247_0, i_8_436_2248_0,
    i_8_436_2271_0, i_8_436_2277_0, i_8_436_2287_0,
    o_8_436_0_0  );
  input  i_8_436_18_0, i_8_436_48_0, i_8_436_78_0, i_8_436_117_0,
    i_8_436_141_0, i_8_436_142_0, i_8_436_219_0, i_8_436_259_0,
    i_8_436_310_0, i_8_436_322_0, i_8_436_336_0, i_8_436_345_0,
    i_8_436_346_0, i_8_436_348_0, i_8_436_360_0, i_8_436_363_0,
    i_8_436_367_0, i_8_436_378_0, i_8_436_381_0, i_8_436_400_0,
    i_8_436_402_0, i_8_436_417_0, i_8_436_427_0, i_8_436_454_0,
    i_8_436_493_0, i_8_436_499_0, i_8_436_579_0, i_8_436_603_0,
    i_8_436_615_0, i_8_436_643_0, i_8_436_654_0, i_8_436_658_0,
    i_8_436_660_0, i_8_436_675_0, i_8_436_696_0, i_8_436_702_0,
    i_8_436_750_0, i_8_436_795_0, i_8_436_799_0, i_8_436_849_0,
    i_8_436_873_0, i_8_436_889_0, i_8_436_991_0, i_8_436_1020_0,
    i_8_436_1056_0, i_8_436_1059_0, i_8_436_1092_0, i_8_436_1104_0,
    i_8_436_1115_0, i_8_436_1146_0, i_8_436_1152_0, i_8_436_1158_0,
    i_8_436_1266_0, i_8_436_1283_0, i_8_436_1284_0, i_8_436_1291_0,
    i_8_436_1314_0, i_8_436_1323_0, i_8_436_1383_0, i_8_436_1426_0,
    i_8_436_1439_0, i_8_436_1440_0, i_8_436_1444_0, i_8_436_1473_0,
    i_8_436_1597_0, i_8_436_1602_0, i_8_436_1633_0, i_8_436_1644_0,
    i_8_436_1671_0, i_8_436_1688_0, i_8_436_1699_0, i_8_436_1702_0,
    i_8_436_1704_0, i_8_436_1723_0, i_8_436_1749_0, i_8_436_1753_0,
    i_8_436_1803_0, i_8_436_1818_0, i_8_436_1830_0, i_8_436_1836_0,
    i_8_436_1840_0, i_8_436_1857_0, i_8_436_1885_0, i_8_436_1887_0,
    i_8_436_1899_0, i_8_436_1944_0, i_8_436_1947_0, i_8_436_1980_0,
    i_8_436_1981_0, i_8_436_2004_0, i_8_436_2184_0, i_8_436_2223_0,
    i_8_436_2227_0, i_8_436_2229_0, i_8_436_2238_0, i_8_436_2247_0,
    i_8_436_2248_0, i_8_436_2271_0, i_8_436_2277_0, i_8_436_2287_0;
  output o_8_436_0_0;
  assign o_8_436_0_0 = 0;
endmodule



// Benchmark "kernel_8_437" written by ABC on Sun Jul 19 10:10:44 2020

module kernel_8_437 ( 
    i_8_437_9_0, i_8_437_58_0, i_8_437_86_0, i_8_437_136_0, i_8_437_138_0,
    i_8_437_139_0, i_8_437_165_0, i_8_437_223_0, i_8_437_363_0,
    i_8_437_370_0, i_8_437_374_0, i_8_437_375_0, i_8_437_385_0,
    i_8_437_417_0, i_8_437_468_0, i_8_437_480_0, i_8_437_499_0,
    i_8_437_507_0, i_8_437_527_0, i_8_437_529_0, i_8_437_547_0,
    i_8_437_554_0, i_8_437_597_0, i_8_437_624_0, i_8_437_625_0,
    i_8_437_715_0, i_8_437_716_0, i_8_437_760_0, i_8_437_761_0,
    i_8_437_762_0, i_8_437_769_0, i_8_437_868_0, i_8_437_873_0,
    i_8_437_906_0, i_8_437_912_0, i_8_437_935_0, i_8_437_938_0,
    i_8_437_945_0, i_8_437_966_0, i_8_437_1029_0, i_8_437_1046_0,
    i_8_437_1050_0, i_8_437_1052_0, i_8_437_1074_0, i_8_437_1104_0,
    i_8_437_1111_0, i_8_437_1114_0, i_8_437_1128_0, i_8_437_1129_0,
    i_8_437_1222_0, i_8_437_1317_0, i_8_437_1323_0, i_8_437_1330_0,
    i_8_437_1346_0, i_8_437_1348_0, i_8_437_1378_0, i_8_437_1380_0,
    i_8_437_1438_0, i_8_437_1456_0, i_8_437_1459_0, i_8_437_1490_0,
    i_8_437_1506_0, i_8_437_1539_0, i_8_437_1542_0, i_8_437_1556_0,
    i_8_437_1560_0, i_8_437_1637_0, i_8_437_1667_0, i_8_437_1669_0,
    i_8_437_1678_0, i_8_437_1682_0, i_8_437_1704_0, i_8_437_1707_0,
    i_8_437_1722_0, i_8_437_1726_0, i_8_437_1753_0, i_8_437_1762_0,
    i_8_437_1785_0, i_8_437_1799_0, i_8_437_1863_0, i_8_437_1918_0,
    i_8_437_1919_0, i_8_437_1934_0, i_8_437_1977_0, i_8_437_1996_0,
    i_8_437_2006_0, i_8_437_2028_0, i_8_437_2101_0, i_8_437_2112_0,
    i_8_437_2119_0, i_8_437_2129_0, i_8_437_2141_0, i_8_437_2190_0,
    i_8_437_2209_0, i_8_437_2211_0, i_8_437_2217_0, i_8_437_2276_0,
    i_8_437_2290_0, i_8_437_2293_0, i_8_437_2294_0,
    o_8_437_0_0  );
  input  i_8_437_9_0, i_8_437_58_0, i_8_437_86_0, i_8_437_136_0,
    i_8_437_138_0, i_8_437_139_0, i_8_437_165_0, i_8_437_223_0,
    i_8_437_363_0, i_8_437_370_0, i_8_437_374_0, i_8_437_375_0,
    i_8_437_385_0, i_8_437_417_0, i_8_437_468_0, i_8_437_480_0,
    i_8_437_499_0, i_8_437_507_0, i_8_437_527_0, i_8_437_529_0,
    i_8_437_547_0, i_8_437_554_0, i_8_437_597_0, i_8_437_624_0,
    i_8_437_625_0, i_8_437_715_0, i_8_437_716_0, i_8_437_760_0,
    i_8_437_761_0, i_8_437_762_0, i_8_437_769_0, i_8_437_868_0,
    i_8_437_873_0, i_8_437_906_0, i_8_437_912_0, i_8_437_935_0,
    i_8_437_938_0, i_8_437_945_0, i_8_437_966_0, i_8_437_1029_0,
    i_8_437_1046_0, i_8_437_1050_0, i_8_437_1052_0, i_8_437_1074_0,
    i_8_437_1104_0, i_8_437_1111_0, i_8_437_1114_0, i_8_437_1128_0,
    i_8_437_1129_0, i_8_437_1222_0, i_8_437_1317_0, i_8_437_1323_0,
    i_8_437_1330_0, i_8_437_1346_0, i_8_437_1348_0, i_8_437_1378_0,
    i_8_437_1380_0, i_8_437_1438_0, i_8_437_1456_0, i_8_437_1459_0,
    i_8_437_1490_0, i_8_437_1506_0, i_8_437_1539_0, i_8_437_1542_0,
    i_8_437_1556_0, i_8_437_1560_0, i_8_437_1637_0, i_8_437_1667_0,
    i_8_437_1669_0, i_8_437_1678_0, i_8_437_1682_0, i_8_437_1704_0,
    i_8_437_1707_0, i_8_437_1722_0, i_8_437_1726_0, i_8_437_1753_0,
    i_8_437_1762_0, i_8_437_1785_0, i_8_437_1799_0, i_8_437_1863_0,
    i_8_437_1918_0, i_8_437_1919_0, i_8_437_1934_0, i_8_437_1977_0,
    i_8_437_1996_0, i_8_437_2006_0, i_8_437_2028_0, i_8_437_2101_0,
    i_8_437_2112_0, i_8_437_2119_0, i_8_437_2129_0, i_8_437_2141_0,
    i_8_437_2190_0, i_8_437_2209_0, i_8_437_2211_0, i_8_437_2217_0,
    i_8_437_2276_0, i_8_437_2290_0, i_8_437_2293_0, i_8_437_2294_0;
  output o_8_437_0_0;
  assign o_8_437_0_0 = 0;
endmodule



// Benchmark "kernel_8_438" written by ABC on Sun Jul 19 10:10:45 2020

module kernel_8_438 ( 
    i_8_438_6_0, i_8_438_21_0, i_8_438_25_0, i_8_438_35_0, i_8_438_78_0,
    i_8_438_79_0, i_8_438_87_0, i_8_438_120_0, i_8_438_121_0,
    i_8_438_123_0, i_8_438_141_0, i_8_438_171_0, i_8_438_193_0,
    i_8_438_195_0, i_8_438_214_0, i_8_438_264_0, i_8_438_268_0,
    i_8_438_286_0, i_8_438_321_0, i_8_438_489_0, i_8_438_492_0,
    i_8_438_582_0, i_8_438_591_0, i_8_438_601_0, i_8_438_627_0,
    i_8_438_628_0, i_8_438_636_0, i_8_438_645_0, i_8_438_672_0,
    i_8_438_693_0, i_8_438_703_0, i_8_438_706_0, i_8_438_735_0,
    i_8_438_813_0, i_8_438_825_0, i_8_438_834_0, i_8_438_835_0,
    i_8_438_860_0, i_8_438_876_0, i_8_438_888_0, i_8_438_969_0,
    i_8_438_978_0, i_8_438_979_0, i_8_438_994_0, i_8_438_1032_0,
    i_8_438_1033_0, i_8_438_1131_0, i_8_438_1167_0, i_8_438_1185_0,
    i_8_438_1187_0, i_8_438_1191_0, i_8_438_1213_0, i_8_438_1230_0,
    i_8_438_1257_0, i_8_438_1264_0, i_8_438_1275_0, i_8_438_1276_0,
    i_8_438_1281_0, i_8_438_1329_0, i_8_438_1330_0, i_8_438_1349_0,
    i_8_438_1362_0, i_8_438_1365_0, i_8_438_1404_0, i_8_438_1407_0,
    i_8_438_1452_0, i_8_438_1455_0, i_8_438_1474_0, i_8_438_1489_0,
    i_8_438_1491_0, i_8_438_1554_0, i_8_438_1573_0, i_8_438_1578_0,
    i_8_438_1582_0, i_8_438_1590_0, i_8_438_1651_0, i_8_438_1668_0,
    i_8_438_1689_0, i_8_438_1749_0, i_8_438_1786_0, i_8_438_1822_0,
    i_8_438_1858_0, i_8_438_1860_0, i_8_438_1861_0, i_8_438_1907_0,
    i_8_438_1965_0, i_8_438_1995_0, i_8_438_2013_0, i_8_438_2058_0,
    i_8_438_2096_0, i_8_438_2140_0, i_8_438_2145_0, i_8_438_2151_0,
    i_8_438_2152_0, i_8_438_2155_0, i_8_438_2172_0, i_8_438_2193_0,
    i_8_438_2194_0, i_8_438_2202_0, i_8_438_2247_0,
    o_8_438_0_0  );
  input  i_8_438_6_0, i_8_438_21_0, i_8_438_25_0, i_8_438_35_0,
    i_8_438_78_0, i_8_438_79_0, i_8_438_87_0, i_8_438_120_0, i_8_438_121_0,
    i_8_438_123_0, i_8_438_141_0, i_8_438_171_0, i_8_438_193_0,
    i_8_438_195_0, i_8_438_214_0, i_8_438_264_0, i_8_438_268_0,
    i_8_438_286_0, i_8_438_321_0, i_8_438_489_0, i_8_438_492_0,
    i_8_438_582_0, i_8_438_591_0, i_8_438_601_0, i_8_438_627_0,
    i_8_438_628_0, i_8_438_636_0, i_8_438_645_0, i_8_438_672_0,
    i_8_438_693_0, i_8_438_703_0, i_8_438_706_0, i_8_438_735_0,
    i_8_438_813_0, i_8_438_825_0, i_8_438_834_0, i_8_438_835_0,
    i_8_438_860_0, i_8_438_876_0, i_8_438_888_0, i_8_438_969_0,
    i_8_438_978_0, i_8_438_979_0, i_8_438_994_0, i_8_438_1032_0,
    i_8_438_1033_0, i_8_438_1131_0, i_8_438_1167_0, i_8_438_1185_0,
    i_8_438_1187_0, i_8_438_1191_0, i_8_438_1213_0, i_8_438_1230_0,
    i_8_438_1257_0, i_8_438_1264_0, i_8_438_1275_0, i_8_438_1276_0,
    i_8_438_1281_0, i_8_438_1329_0, i_8_438_1330_0, i_8_438_1349_0,
    i_8_438_1362_0, i_8_438_1365_0, i_8_438_1404_0, i_8_438_1407_0,
    i_8_438_1452_0, i_8_438_1455_0, i_8_438_1474_0, i_8_438_1489_0,
    i_8_438_1491_0, i_8_438_1554_0, i_8_438_1573_0, i_8_438_1578_0,
    i_8_438_1582_0, i_8_438_1590_0, i_8_438_1651_0, i_8_438_1668_0,
    i_8_438_1689_0, i_8_438_1749_0, i_8_438_1786_0, i_8_438_1822_0,
    i_8_438_1858_0, i_8_438_1860_0, i_8_438_1861_0, i_8_438_1907_0,
    i_8_438_1965_0, i_8_438_1995_0, i_8_438_2013_0, i_8_438_2058_0,
    i_8_438_2096_0, i_8_438_2140_0, i_8_438_2145_0, i_8_438_2151_0,
    i_8_438_2152_0, i_8_438_2155_0, i_8_438_2172_0, i_8_438_2193_0,
    i_8_438_2194_0, i_8_438_2202_0, i_8_438_2247_0;
  output o_8_438_0_0;
  assign o_8_438_0_0 = 0;
endmodule



// Benchmark "kernel_8_439" written by ABC on Sun Jul 19 10:10:47 2020

module kernel_8_439 ( 
    i_8_439_51_0, i_8_439_52_0, i_8_439_57_0, i_8_439_60_0, i_8_439_61_0,
    i_8_439_62_0, i_8_439_85_0, i_8_439_142_0, i_8_439_216_0,
    i_8_439_226_0, i_8_439_229_0, i_8_439_230_0, i_8_439_255_0,
    i_8_439_257_0, i_8_439_258_0, i_8_439_259_0, i_8_439_260_0,
    i_8_439_301_0, i_8_439_329_0, i_8_439_379_0, i_8_439_389_0,
    i_8_439_426_0, i_8_439_453_0, i_8_439_485_0, i_8_439_554_0,
    i_8_439_556_0, i_8_439_557_0, i_8_439_597_0, i_8_439_602_0,
    i_8_439_678_0, i_8_439_786_0, i_8_439_851_0, i_8_439_852_0,
    i_8_439_853_0, i_8_439_877_0, i_8_439_971_0, i_8_439_991_0,
    i_8_439_992_0, i_8_439_1013_0, i_8_439_1050_0, i_8_439_1052_0,
    i_8_439_1112_0, i_8_439_1120_0, i_8_439_1124_0, i_8_439_1129_0,
    i_8_439_1137_0, i_8_439_1159_0, i_8_439_1238_0, i_8_439_1261_0,
    i_8_439_1281_0, i_8_439_1286_0, i_8_439_1315_0, i_8_439_1316_0,
    i_8_439_1342_0, i_8_439_1407_0, i_8_439_1410_0, i_8_439_1411_0,
    i_8_439_1449_0, i_8_439_1489_0, i_8_439_1490_0, i_8_439_1535_0,
    i_8_439_1537_0, i_8_439_1545_0, i_8_439_1549_0, i_8_439_1551_0,
    i_8_439_1552_0, i_8_439_1553_0, i_8_439_1561_0, i_8_439_1564_0,
    i_8_439_1615_0, i_8_439_1625_0, i_8_439_1632_0, i_8_439_1633_0,
    i_8_439_1652_0, i_8_439_1653_0, i_8_439_1655_0, i_8_439_1696_0,
    i_8_439_1782_0, i_8_439_1789_0, i_8_439_1805_0, i_8_439_1813_0,
    i_8_439_1855_0, i_8_439_1858_0, i_8_439_1884_0, i_8_439_1885_0,
    i_8_439_1887_0, i_8_439_1888_0, i_8_439_1889_0, i_8_439_1944_0,
    i_8_439_1996_0, i_8_439_2028_0, i_8_439_2032_0, i_8_439_2048_0,
    i_8_439_2073_0, i_8_439_2139_0, i_8_439_2143_0, i_8_439_2147_0,
    i_8_439_2216_0, i_8_439_2236_0, i_8_439_2273_0,
    o_8_439_0_0  );
  input  i_8_439_51_0, i_8_439_52_0, i_8_439_57_0, i_8_439_60_0,
    i_8_439_61_0, i_8_439_62_0, i_8_439_85_0, i_8_439_142_0, i_8_439_216_0,
    i_8_439_226_0, i_8_439_229_0, i_8_439_230_0, i_8_439_255_0,
    i_8_439_257_0, i_8_439_258_0, i_8_439_259_0, i_8_439_260_0,
    i_8_439_301_0, i_8_439_329_0, i_8_439_379_0, i_8_439_389_0,
    i_8_439_426_0, i_8_439_453_0, i_8_439_485_0, i_8_439_554_0,
    i_8_439_556_0, i_8_439_557_0, i_8_439_597_0, i_8_439_602_0,
    i_8_439_678_0, i_8_439_786_0, i_8_439_851_0, i_8_439_852_0,
    i_8_439_853_0, i_8_439_877_0, i_8_439_971_0, i_8_439_991_0,
    i_8_439_992_0, i_8_439_1013_0, i_8_439_1050_0, i_8_439_1052_0,
    i_8_439_1112_0, i_8_439_1120_0, i_8_439_1124_0, i_8_439_1129_0,
    i_8_439_1137_0, i_8_439_1159_0, i_8_439_1238_0, i_8_439_1261_0,
    i_8_439_1281_0, i_8_439_1286_0, i_8_439_1315_0, i_8_439_1316_0,
    i_8_439_1342_0, i_8_439_1407_0, i_8_439_1410_0, i_8_439_1411_0,
    i_8_439_1449_0, i_8_439_1489_0, i_8_439_1490_0, i_8_439_1535_0,
    i_8_439_1537_0, i_8_439_1545_0, i_8_439_1549_0, i_8_439_1551_0,
    i_8_439_1552_0, i_8_439_1553_0, i_8_439_1561_0, i_8_439_1564_0,
    i_8_439_1615_0, i_8_439_1625_0, i_8_439_1632_0, i_8_439_1633_0,
    i_8_439_1652_0, i_8_439_1653_0, i_8_439_1655_0, i_8_439_1696_0,
    i_8_439_1782_0, i_8_439_1789_0, i_8_439_1805_0, i_8_439_1813_0,
    i_8_439_1855_0, i_8_439_1858_0, i_8_439_1884_0, i_8_439_1885_0,
    i_8_439_1887_0, i_8_439_1888_0, i_8_439_1889_0, i_8_439_1944_0,
    i_8_439_1996_0, i_8_439_2028_0, i_8_439_2032_0, i_8_439_2048_0,
    i_8_439_2073_0, i_8_439_2139_0, i_8_439_2143_0, i_8_439_2147_0,
    i_8_439_2216_0, i_8_439_2236_0, i_8_439_2273_0;
  output o_8_439_0_0;
  assign o_8_439_0_0 = ~((~i_8_439_229_0 & ((~i_8_439_52_0 & i_8_439_257_0 & ~i_8_439_1137_0 & ~i_8_439_1410_0 & ~i_8_439_1564_0 & i_8_439_1805_0) | (~i_8_439_57_0 & ~i_8_439_142_0 & ~i_8_439_230_0 & ~i_8_439_877_0 & ~i_8_439_1281_0 & ~i_8_439_1315_0 & ~i_8_439_1944_0 & ~i_8_439_2032_0 & i_8_439_2236_0))) | (~i_8_439_1789_0 & ((~i_8_439_60_0 & ~i_8_439_1315_0 & ((~i_8_439_301_0 & ~i_8_439_426_0 & ~i_8_439_786_0 & ~i_8_439_852_0 & ~i_8_439_1052_0 & i_8_439_1411_0) | (~i_8_439_52_0 & i_8_439_216_0 & ~i_8_439_226_0 & ~i_8_439_255_0 & ~i_8_439_992_0 & ~i_8_439_1615_0 & ~i_8_439_1632_0 & ~i_8_439_1652_0 & ~i_8_439_2028_0 & ~i_8_439_2236_0))) | (~i_8_439_142_0 & ((i_8_439_329_0 & i_8_439_992_0 & ~i_8_439_1782_0 & ~i_8_439_1813_0) | (~i_8_439_62_0 & ~i_8_439_257_0 & ~i_8_439_329_0 & i_8_439_1286_0 & ~i_8_439_1633_0 & ~i_8_439_1858_0 & ~i_8_439_2236_0))) | (~i_8_439_1052_0 & ((~i_8_439_485_0 & ((~i_8_439_57_0 & i_8_439_61_0 & ~i_8_439_678_0 & ~i_8_439_786_0 & ~i_8_439_1286_0 & ~i_8_439_1805_0 & ~i_8_439_2032_0) | (~i_8_439_85_0 & ~i_8_439_226_0 & ~i_8_439_260_0 & ~i_8_439_389_0 & ~i_8_439_453_0 & ~i_8_439_597_0 & ~i_8_439_852_0 & i_8_439_877_0 & ~i_8_439_971_0 & ~i_8_439_1281_0 & ~i_8_439_1316_0 & ~i_8_439_2139_0))) | (~i_8_439_51_0 & ~i_8_439_255_0 & ~i_8_439_678_0 & ~i_8_439_991_0 & i_8_439_1551_0 & ~i_8_439_1564_0 & ~i_8_439_1813_0 & ~i_8_439_1944_0 & ~i_8_439_2028_0))) | (~i_8_439_602_0 & ~i_8_439_851_0 & i_8_439_2147_0 & ~i_8_439_2236_0))) | (~i_8_439_453_0 & ((~i_8_439_226_0 & ((~i_8_439_142_0 & i_8_439_301_0 & ~i_8_439_1050_0 & ~i_8_439_1159_0 & i_8_439_1652_0) | (~i_8_439_60_0 & ~i_8_439_597_0 & ~i_8_439_1052_0 & ~i_8_439_1315_0 & ~i_8_439_1535_0 & ~i_8_439_1549_0 & i_8_439_1551_0 & ~i_8_439_1813_0 & ~i_8_439_1944_0))) | (~i_8_439_61_0 & ~i_8_439_259_0 & ~i_8_439_329_0 & ~i_8_439_678_0 & ~i_8_439_1050_0 & i_8_439_1112_0 & ~i_8_439_1124_0 & ~i_8_439_1996_0 & ~i_8_439_2032_0) | (~i_8_439_51_0 & ~i_8_439_52_0 & ~i_8_439_57_0 & ~i_8_439_230_0 & ~i_8_439_1052_0 & ~i_8_439_1535_0 & i_8_439_1549_0 & ~i_8_439_1625_0 & ~i_8_439_1858_0 & ~i_8_439_2048_0) | (~i_8_439_62_0 & ~i_8_439_852_0 & ~i_8_439_853_0 & ~i_8_439_971_0 & ~i_8_439_1889_0 & i_8_439_2273_0))) | (~i_8_439_230_0 & ((~i_8_439_52_0 & ~i_8_439_852_0 & ~i_8_439_971_0 & i_8_439_1553_0 & ~i_8_439_1561_0 & ~i_8_439_1782_0 & ~i_8_439_1813_0 & ~i_8_439_2032_0) | (i_8_439_257_0 & ~i_8_439_329_0 & ~i_8_439_678_0 & ~i_8_439_1238_0 & i_8_439_2216_0))) | (~i_8_439_853_0 & ((~i_8_439_57_0 & (i_8_439_1653_0 | (~i_8_439_51_0 & ~i_8_439_329_0 & i_8_439_556_0 & ~i_8_439_971_0 & ~i_8_439_1120_0 & ~i_8_439_1782_0))) | (~i_8_439_60_0 & ~i_8_439_786_0 & ((~i_8_439_62_0 & ~i_8_439_597_0 & ~i_8_439_1813_0 & i_8_439_1885_0 & ~i_8_439_1996_0) | (~i_8_439_61_0 & i_8_439_301_0 & ~i_8_439_556_0 & ~i_8_439_851_0 & ~i_8_439_991_0 & ~i_8_439_1137_0 & i_8_439_1281_0 & ~i_8_439_1315_0 & ~i_8_439_1615_0 & ~i_8_439_2032_0 & ~i_8_439_2048_0))) | (~i_8_439_260_0 & ((~i_8_439_61_0 & ~i_8_439_62_0 & i_8_439_379_0 & ~i_8_439_426_0 & ~i_8_439_597_0 & ~i_8_439_678_0 & ~i_8_439_971_0 & ~i_8_439_1449_0 & ~i_8_439_1564_0 & ~i_8_439_1632_0) | (i_8_439_971_0 & ~i_8_439_1561_0 & i_8_439_1888_0))) | (~i_8_439_142_0 & ~i_8_439_877_0 & ~i_8_439_1052_0 & ~i_8_439_1286_0 & ~i_8_439_1633_0 & ~i_8_439_1652_0 & ~i_8_439_1782_0 & i_8_439_1889_0 & ~i_8_439_1996_0))) | (~i_8_439_379_0 & ((~i_8_439_57_0 & ~i_8_439_301_0 & ~i_8_439_1052_0 & ~i_8_439_1615_0 & i_8_439_1655_0 & ~i_8_439_1858_0) | (i_8_439_1013_0 & i_8_439_1052_0 & ~i_8_439_1281_0 & i_8_439_1286_0 & ~i_8_439_2032_0))) | (~i_8_439_1561_0 & ((~i_8_439_51_0 & ~i_8_439_62_0 & ((~i_8_439_61_0 & ~i_8_439_257_0 & ~i_8_439_301_0 & ~i_8_439_597_0 & ~i_8_439_678_0 & ~i_8_439_851_0 & ~i_8_439_971_0 & ~i_8_439_1238_0 & ~i_8_439_1316_0 & ~i_8_439_1944_0 & ~i_8_439_2028_0 & ~i_8_439_1535_0 & i_8_439_1552_0) | (~i_8_439_1013_0 & i_8_439_1884_0 & i_8_439_2139_0))) | (~i_8_439_52_0 & ~i_8_439_57_0 & ~i_8_439_786_0 & ((~i_8_439_301_0 & ~i_8_439_1545_0 & i_8_439_1888_0 & ~i_8_439_1889_0) | (~i_8_439_258_0 & i_8_439_453_0 & ~i_8_439_992_0 & ~i_8_439_1316_0 & ~i_8_439_1410_0 & ~i_8_439_1535_0 & ~i_8_439_1551_0 & ~i_8_439_1632_0 & ~i_8_439_2032_0 & ~i_8_439_2236_0))))) | (~i_8_439_51_0 & ((~i_8_439_257_0 & ~i_8_439_258_0 & ~i_8_439_597_0 & ~i_8_439_786_0 & ~i_8_439_1052_0 & i_8_439_1537_0 & ~i_8_439_1552_0 & ~i_8_439_1633_0 & ~i_8_439_1944_0 & ~i_8_439_2216_0) | (~i_8_439_142_0 & i_8_439_329_0 & i_8_439_851_0 & ~i_8_439_1013_0 & ~i_8_439_1782_0 & i_8_439_1996_0 & ~i_8_439_2139_0 & ~i_8_439_2236_0))) | (~i_8_439_258_0 & ((i_8_439_1653_0 & i_8_439_1887_0) | (~i_8_439_57_0 & ~i_8_439_60_0 & ~i_8_439_851_0 & ~i_8_439_852_0 & ~i_8_439_971_0 & ~i_8_439_1137_0 & i_8_439_1888_0))) | (~i_8_439_62_0 & ((~i_8_439_57_0 & ~i_8_439_257_0 & i_8_439_1652_0 & ((~i_8_439_61_0 & i_8_439_554_0) | (~i_8_439_142_0 & ~i_8_439_602_0 & ~i_8_439_786_0 & ~i_8_439_852_0))) | (~i_8_439_52_0 & ~i_8_439_485_0 & ~i_8_439_678_0 & i_8_439_1052_0 & i_8_439_1655_0) | (i_8_439_1411_0 & i_8_439_1889_0))) | (~i_8_439_52_0 & ((~i_8_439_786_0 & ~i_8_439_1052_0 & i_8_439_1112_0 & i_8_439_1238_0 & ~i_8_439_1615_0 & ~i_8_439_1633_0) | (~i_8_439_61_0 & ~i_8_439_971_0 & ~i_8_439_1159_0 & i_8_439_1552_0 & i_8_439_1858_0))) | (~i_8_439_61_0 & ((~i_8_439_329_0 & ~i_8_439_971_0 & ~i_8_439_991_0 & ~i_8_439_992_0 & i_8_439_1286_0 & ~i_8_439_1316_0 & ~i_8_439_1625_0 & ~i_8_439_1655_0 & ~i_8_439_1805_0 & ~i_8_439_1885_0 & ~i_8_439_1887_0) | (~i_8_439_60_0 & ~i_8_439_142_0 & i_8_439_453_0 & ~i_8_439_786_0 & i_8_439_1050_0 & ~i_8_439_1052_0 & ~i_8_439_1137_0 & ~i_8_439_1782_0 & ~i_8_439_2216_0))) | (~i_8_439_60_0 & ((~i_8_439_142_0 & i_8_439_554_0 & ~i_8_439_851_0 & i_8_439_1805_0) | (~i_8_439_597_0 & ~i_8_439_877_0 & i_8_439_1884_0))) | (~i_8_439_786_0 & ((~i_8_439_678_0 & ~i_8_439_2073_0 & ((i_8_439_229_0 & ~i_8_439_1120_0 & i_8_439_1632_0 & ~i_8_439_1696_0 & ~i_8_439_2139_0 & ~i_8_439_2216_0) | (~i_8_439_257_0 & ~i_8_439_485_0 & ~i_8_439_602_0 & ~i_8_439_1124_0 & ~i_8_439_2032_0 & i_8_439_2143_0 & ~i_8_439_2273_0))) | (~i_8_439_851_0 & ~i_8_439_1552_0 & ~i_8_439_1632_0 & ~i_8_439_1813_0 & i_8_439_1858_0))) | (~i_8_439_2032_0 & ((~i_8_439_554_0 & ~i_8_439_851_0 & ~i_8_439_1050_0 & ~i_8_439_1535_0 & ~i_8_439_1549_0 & ~i_8_439_1124_0 & i_8_439_1238_0) | (~i_8_439_259_0 & i_8_439_597_0 & ~i_8_439_991_0 & ~i_8_439_1112_0 & ~i_8_439_1615_0 & i_8_439_1944_0 & ~i_8_439_1996_0))) | (~i_8_439_2139_0 & ((i_8_439_557_0 & ~i_8_439_1261_0 & i_8_439_1553_0 & ~i_8_439_2073_0) | (~i_8_439_142_0 & ~i_8_439_877_0 & ~i_8_439_1315_0 & i_8_439_1696_0 & ~i_8_439_1889_0 & ~i_8_439_2216_0))) | (i_8_439_1888_0 & i_8_439_2048_0));
endmodule



// Benchmark "kernel_8_440" written by ABC on Sun Jul 19 10:10:48 2020

module kernel_8_440 ( 
    i_8_440_13_0, i_8_440_77_0, i_8_440_80_0, i_8_440_140_0, i_8_440_167_0,
    i_8_440_184_0, i_8_440_221_0, i_8_440_233_0, i_8_440_253_0,
    i_8_440_254_0, i_8_440_259_0, i_8_440_263_0, i_8_440_281_0,
    i_8_440_284_0, i_8_440_302_0, i_8_440_304_0, i_8_440_322_0,
    i_8_440_335_0, i_8_440_364_0, i_8_440_376_0, i_8_440_400_0,
    i_8_440_437_0, i_8_440_439_0, i_8_440_440_0, i_8_440_488_0,
    i_8_440_494_0, i_8_440_578_0, i_8_440_580_0, i_8_440_590_0,
    i_8_440_619_0, i_8_440_625_0, i_8_440_626_0, i_8_440_643_0,
    i_8_440_662_0, i_8_440_664_0, i_8_440_698_0, i_8_440_702_0,
    i_8_440_707_0, i_8_440_712_0, i_8_440_716_0, i_8_440_725_0,
    i_8_440_732_0, i_8_440_808_0, i_8_440_812_0, i_8_440_853_0,
    i_8_440_869_0, i_8_440_878_0, i_8_440_942_0, i_8_440_968_0,
    i_8_440_1027_0, i_8_440_1057_0, i_8_440_1067_0, i_8_440_1075_0,
    i_8_440_1143_0, i_8_440_1192_0, i_8_440_1211_0, i_8_440_1220_0,
    i_8_440_1241_0, i_8_440_1277_0, i_8_440_1282_0, i_8_440_1323_0,
    i_8_440_1370_0, i_8_440_1411_0, i_8_440_1436_0, i_8_440_1453_0,
    i_8_440_1480_0, i_8_440_1489_0, i_8_440_1552_0, i_8_440_1561_0,
    i_8_440_1618_0, i_8_440_1625_0, i_8_440_1697_0, i_8_440_1716_0,
    i_8_440_1723_0, i_8_440_1729_0, i_8_440_1769_0, i_8_440_1779_0,
    i_8_440_1780_0, i_8_440_1801_0, i_8_440_1808_0, i_8_440_1825_0,
    i_8_440_1849_0, i_8_440_1855_0, i_8_440_1904_0, i_8_440_1945_0,
    i_8_440_1970_0, i_8_440_1993_0, i_8_440_2039_0, i_8_440_2083_0,
    i_8_440_2111_0, i_8_440_2129_0, i_8_440_2191_0, i_8_440_2192_0,
    i_8_440_2228_0, i_8_440_2245_0, i_8_440_2247_0, i_8_440_2248_0,
    i_8_440_2261_0, i_8_440_2282_0, i_8_440_2301_0,
    o_8_440_0_0  );
  input  i_8_440_13_0, i_8_440_77_0, i_8_440_80_0, i_8_440_140_0,
    i_8_440_167_0, i_8_440_184_0, i_8_440_221_0, i_8_440_233_0,
    i_8_440_253_0, i_8_440_254_0, i_8_440_259_0, i_8_440_263_0,
    i_8_440_281_0, i_8_440_284_0, i_8_440_302_0, i_8_440_304_0,
    i_8_440_322_0, i_8_440_335_0, i_8_440_364_0, i_8_440_376_0,
    i_8_440_400_0, i_8_440_437_0, i_8_440_439_0, i_8_440_440_0,
    i_8_440_488_0, i_8_440_494_0, i_8_440_578_0, i_8_440_580_0,
    i_8_440_590_0, i_8_440_619_0, i_8_440_625_0, i_8_440_626_0,
    i_8_440_643_0, i_8_440_662_0, i_8_440_664_0, i_8_440_698_0,
    i_8_440_702_0, i_8_440_707_0, i_8_440_712_0, i_8_440_716_0,
    i_8_440_725_0, i_8_440_732_0, i_8_440_808_0, i_8_440_812_0,
    i_8_440_853_0, i_8_440_869_0, i_8_440_878_0, i_8_440_942_0,
    i_8_440_968_0, i_8_440_1027_0, i_8_440_1057_0, i_8_440_1067_0,
    i_8_440_1075_0, i_8_440_1143_0, i_8_440_1192_0, i_8_440_1211_0,
    i_8_440_1220_0, i_8_440_1241_0, i_8_440_1277_0, i_8_440_1282_0,
    i_8_440_1323_0, i_8_440_1370_0, i_8_440_1411_0, i_8_440_1436_0,
    i_8_440_1453_0, i_8_440_1480_0, i_8_440_1489_0, i_8_440_1552_0,
    i_8_440_1561_0, i_8_440_1618_0, i_8_440_1625_0, i_8_440_1697_0,
    i_8_440_1716_0, i_8_440_1723_0, i_8_440_1729_0, i_8_440_1769_0,
    i_8_440_1779_0, i_8_440_1780_0, i_8_440_1801_0, i_8_440_1808_0,
    i_8_440_1825_0, i_8_440_1849_0, i_8_440_1855_0, i_8_440_1904_0,
    i_8_440_1945_0, i_8_440_1970_0, i_8_440_1993_0, i_8_440_2039_0,
    i_8_440_2083_0, i_8_440_2111_0, i_8_440_2129_0, i_8_440_2191_0,
    i_8_440_2192_0, i_8_440_2228_0, i_8_440_2245_0, i_8_440_2247_0,
    i_8_440_2248_0, i_8_440_2261_0, i_8_440_2282_0, i_8_440_2301_0;
  output o_8_440_0_0;
  assign o_8_440_0_0 = 0;
endmodule



// Benchmark "kernel_8_441" written by ABC on Sun Jul 19 10:10:49 2020

module kernel_8_441 ( 
    i_8_441_19_0, i_8_441_22_0, i_8_441_23_0, i_8_441_107_0, i_8_441_125_0,
    i_8_441_144_0, i_8_441_176_0, i_8_441_221_0, i_8_441_223_0,
    i_8_441_224_0, i_8_441_266_0, i_8_441_281_0, i_8_441_296_0,
    i_8_441_329_0, i_8_441_349_0, i_8_441_418_0, i_8_441_428_0,
    i_8_441_437_0, i_8_441_439_0, i_8_441_440_0, i_8_441_490_0,
    i_8_441_491_0, i_8_441_492_0, i_8_441_493_0, i_8_441_499_0,
    i_8_441_527_0, i_8_441_530_0, i_8_441_611_0, i_8_441_632_0,
    i_8_441_671_0, i_8_441_698_0, i_8_441_700_0, i_8_441_702_0,
    i_8_441_703_0, i_8_441_704_0, i_8_441_705_0, i_8_441_706_0,
    i_8_441_707_0, i_8_441_710_0, i_8_441_728_0, i_8_441_736_0,
    i_8_441_809_0, i_8_441_827_0, i_8_441_836_0, i_8_441_841_0,
    i_8_441_842_0, i_8_441_844_0, i_8_441_845_0, i_8_441_964_0,
    i_8_441_971_0, i_8_441_1047_0, i_8_441_1073_0, i_8_441_1103_0,
    i_8_441_1157_0, i_8_441_1183_0, i_8_441_1184_0, i_8_441_1300_0,
    i_8_441_1310_0, i_8_441_1358_0, i_8_441_1363_0, i_8_441_1390_0,
    i_8_441_1405_0, i_8_441_1411_0, i_8_441_1434_0, i_8_441_1442_0,
    i_8_441_1471_0, i_8_441_1473_0, i_8_441_1546_0, i_8_441_1565_0,
    i_8_441_1589_0, i_8_441_1592_0, i_8_441_1607_0, i_8_441_1628_0,
    i_8_441_1633_0, i_8_441_1643_0, i_8_441_1650_0, i_8_441_1681_0,
    i_8_441_1694_0, i_8_441_1733_0, i_8_441_1751_0, i_8_441_1771_0,
    i_8_441_1778_0, i_8_441_1817_0, i_8_441_1850_0, i_8_441_1862_0,
    i_8_441_1867_0, i_8_441_1871_0, i_8_441_1991_0, i_8_441_2026_0,
    i_8_441_2028_0, i_8_441_2030_0, i_8_441_2032_0, i_8_441_2074_0,
    i_8_441_2111_0, i_8_441_2120_0, i_8_441_2140_0, i_8_441_2189_0,
    i_8_441_2191_0, i_8_441_2192_0, i_8_441_2243_0,
    o_8_441_0_0  );
  input  i_8_441_19_0, i_8_441_22_0, i_8_441_23_0, i_8_441_107_0,
    i_8_441_125_0, i_8_441_144_0, i_8_441_176_0, i_8_441_221_0,
    i_8_441_223_0, i_8_441_224_0, i_8_441_266_0, i_8_441_281_0,
    i_8_441_296_0, i_8_441_329_0, i_8_441_349_0, i_8_441_418_0,
    i_8_441_428_0, i_8_441_437_0, i_8_441_439_0, i_8_441_440_0,
    i_8_441_490_0, i_8_441_491_0, i_8_441_492_0, i_8_441_493_0,
    i_8_441_499_0, i_8_441_527_0, i_8_441_530_0, i_8_441_611_0,
    i_8_441_632_0, i_8_441_671_0, i_8_441_698_0, i_8_441_700_0,
    i_8_441_702_0, i_8_441_703_0, i_8_441_704_0, i_8_441_705_0,
    i_8_441_706_0, i_8_441_707_0, i_8_441_710_0, i_8_441_728_0,
    i_8_441_736_0, i_8_441_809_0, i_8_441_827_0, i_8_441_836_0,
    i_8_441_841_0, i_8_441_842_0, i_8_441_844_0, i_8_441_845_0,
    i_8_441_964_0, i_8_441_971_0, i_8_441_1047_0, i_8_441_1073_0,
    i_8_441_1103_0, i_8_441_1157_0, i_8_441_1183_0, i_8_441_1184_0,
    i_8_441_1300_0, i_8_441_1310_0, i_8_441_1358_0, i_8_441_1363_0,
    i_8_441_1390_0, i_8_441_1405_0, i_8_441_1411_0, i_8_441_1434_0,
    i_8_441_1442_0, i_8_441_1471_0, i_8_441_1473_0, i_8_441_1546_0,
    i_8_441_1565_0, i_8_441_1589_0, i_8_441_1592_0, i_8_441_1607_0,
    i_8_441_1628_0, i_8_441_1633_0, i_8_441_1643_0, i_8_441_1650_0,
    i_8_441_1681_0, i_8_441_1694_0, i_8_441_1733_0, i_8_441_1751_0,
    i_8_441_1771_0, i_8_441_1778_0, i_8_441_1817_0, i_8_441_1850_0,
    i_8_441_1862_0, i_8_441_1867_0, i_8_441_1871_0, i_8_441_1991_0,
    i_8_441_2026_0, i_8_441_2028_0, i_8_441_2030_0, i_8_441_2032_0,
    i_8_441_2074_0, i_8_441_2111_0, i_8_441_2120_0, i_8_441_2140_0,
    i_8_441_2189_0, i_8_441_2191_0, i_8_441_2192_0, i_8_441_2243_0;
  output o_8_441_0_0;
  assign o_8_441_0_0 = ~((~i_8_441_266_0 & ((~i_8_441_704_0 & ~i_8_441_710_0 & ~i_8_441_736_0 & i_8_441_1681_0) | (~i_8_441_107_0 & ~i_8_441_223_0 & ~i_8_441_1073_0 & ~i_8_441_1358_0 & ~i_8_441_1442_0 & ~i_8_441_1771_0 & ~i_8_441_2028_0 & ~i_8_441_2140_0))) | (~i_8_441_296_0 & ((i_8_441_224_0 & ~i_8_441_703_0 & ~i_8_441_1183_0 & ~i_8_441_1184_0 & ~i_8_441_1628_0) | (i_8_441_428_0 & ~i_8_441_439_0 & ~i_8_441_1991_0))) | (i_8_441_527_0 & ((~i_8_441_841_0 & ~i_8_441_845_0) | (~i_8_441_698_0 & ~i_8_441_1592_0))) | (~i_8_441_728_0 & ((i_8_441_223_0 & i_8_441_493_0 & ~i_8_441_1681_0 & ~i_8_441_1862_0 & ~i_8_441_2028_0 & ~i_8_441_2120_0) | (~i_8_441_281_0 & ~i_8_441_439_0 & ~i_8_441_971_0 & ~i_8_441_1047_0 & ~i_8_441_1358_0 & ~i_8_441_1628_0 & ~i_8_441_1771_0 & ~i_8_441_2140_0))) | (~i_8_441_809_0 & ((~i_8_441_493_0 & ~i_8_441_844_0 & ~i_8_441_1442_0 & ~i_8_441_1589_0 & ~i_8_441_1817_0) | (~i_8_441_1363_0 & i_8_441_1778_0 & ~i_8_441_2030_0))) | (~i_8_441_836_0 & ((i_8_441_710_0 & ~i_8_441_1363_0 & ~i_8_441_1546_0 & ~i_8_441_1589_0) | (~i_8_441_439_0 & i_8_441_491_0 & ~i_8_441_827_0 & ~i_8_441_1157_0 & ~i_8_441_1411_0 & ~i_8_441_1442_0 & ~i_8_441_2032_0 & ~i_8_441_2192_0))) | (~i_8_441_1358_0 & ((~i_8_441_439_0 & ~i_8_441_698_0 & ~i_8_441_736_0 & ~i_8_441_2032_0) | (~i_8_441_700_0 & ~i_8_441_971_0 & ~i_8_441_1073_0 & ~i_8_441_1771_0 & ~i_8_441_2030_0 & ~i_8_441_2189_0))) | (~i_8_441_439_0 & ((~i_8_441_329_0 & ~i_8_441_490_0 & i_8_441_736_0 & ~i_8_441_1310_0 & ~i_8_441_1442_0) | (~i_8_441_611_0 & ~i_8_441_703_0 & ~i_8_441_1183_0 & ~i_8_441_1434_0 & ~i_8_441_1589_0 & ~i_8_441_1592_0 & ~i_8_441_1694_0 & ~i_8_441_1817_0 & ~i_8_441_2189_0))) | (~i_8_441_971_0 & ~i_8_441_2028_0 & ((~i_8_441_437_0 & ~i_8_441_440_0 & ~i_8_441_1589_0 & i_8_441_1681_0) | (~i_8_441_842_0 & ~i_8_441_1363_0 & ~i_8_441_1434_0 & ~i_8_441_1817_0 & ~i_8_441_1850_0 & ~i_8_441_2030_0))) | (~i_8_441_440_0 & (i_8_441_705_0 | (~i_8_441_671_0 & i_8_441_1778_0))) | (i_8_441_1300_0 & i_8_441_2192_0) | (i_8_441_703_0 & ~i_8_441_1733_0 & ~i_8_441_2192_0));
endmodule



// Benchmark "kernel_8_442" written by ABC on Sun Jul 19 10:10:50 2020

module kernel_8_442 ( 
    i_8_442_7_0, i_8_442_29_0, i_8_442_49_0, i_8_442_58_0, i_8_442_89_0,
    i_8_442_96_0, i_8_442_97_0, i_8_442_113_0, i_8_442_169_0,
    i_8_442_174_0, i_8_442_184_0, i_8_442_232_0, i_8_442_239_0,
    i_8_442_254_0, i_8_442_259_0, i_8_442_268_0, i_8_442_292_0,
    i_8_442_297_0, i_8_442_329_0, i_8_442_335_0, i_8_442_371_0,
    i_8_442_374_0, i_8_442_418_0, i_8_442_432_0, i_8_442_443_0,
    i_8_442_468_0, i_8_442_479_0, i_8_442_481_0, i_8_442_500_0,
    i_8_442_508_0, i_8_442_510_0, i_8_442_524_0, i_8_442_525_0,
    i_8_442_528_0, i_8_442_529_0, i_8_442_556_0, i_8_442_572_0,
    i_8_442_595_0, i_8_442_600_0, i_8_442_636_0, i_8_442_659_0,
    i_8_442_665_0, i_8_442_690_0, i_8_442_705_0, i_8_442_735_0,
    i_8_442_770_0, i_8_442_789_0, i_8_442_849_0, i_8_442_857_0,
    i_8_442_875_0, i_8_442_1039_0, i_8_442_1075_0, i_8_442_1093_0,
    i_8_442_1189_0, i_8_442_1190_0, i_8_442_1200_0, i_8_442_1219_0,
    i_8_442_1277_0, i_8_442_1293_0, i_8_442_1297_0, i_8_442_1307_0,
    i_8_442_1348_0, i_8_442_1408_0, i_8_442_1410_0, i_8_442_1437_0,
    i_8_442_1471_0, i_8_442_1487_0, i_8_442_1531_0, i_8_442_1536_0,
    i_8_442_1545_0, i_8_442_1586_0, i_8_442_1624_0, i_8_442_1633_0,
    i_8_442_1634_0, i_8_442_1669_0, i_8_442_1696_0, i_8_442_1704_0,
    i_8_442_1724_0, i_8_442_1739_0, i_8_442_1742_0, i_8_442_1768_0,
    i_8_442_1779_0, i_8_442_1794_0, i_8_442_1795_0, i_8_442_1799_0,
    i_8_442_1874_0, i_8_442_1906_0, i_8_442_1918_0, i_8_442_1957_0,
    i_8_442_1958_0, i_8_442_1965_0, i_8_442_1969_0, i_8_442_1981_0,
    i_8_442_2019_0, i_8_442_2032_0, i_8_442_2116_0, i_8_442_2122_0,
    i_8_442_2149_0, i_8_442_2236_0, i_8_442_2246_0,
    o_8_442_0_0  );
  input  i_8_442_7_0, i_8_442_29_0, i_8_442_49_0, i_8_442_58_0,
    i_8_442_89_0, i_8_442_96_0, i_8_442_97_0, i_8_442_113_0, i_8_442_169_0,
    i_8_442_174_0, i_8_442_184_0, i_8_442_232_0, i_8_442_239_0,
    i_8_442_254_0, i_8_442_259_0, i_8_442_268_0, i_8_442_292_0,
    i_8_442_297_0, i_8_442_329_0, i_8_442_335_0, i_8_442_371_0,
    i_8_442_374_0, i_8_442_418_0, i_8_442_432_0, i_8_442_443_0,
    i_8_442_468_0, i_8_442_479_0, i_8_442_481_0, i_8_442_500_0,
    i_8_442_508_0, i_8_442_510_0, i_8_442_524_0, i_8_442_525_0,
    i_8_442_528_0, i_8_442_529_0, i_8_442_556_0, i_8_442_572_0,
    i_8_442_595_0, i_8_442_600_0, i_8_442_636_0, i_8_442_659_0,
    i_8_442_665_0, i_8_442_690_0, i_8_442_705_0, i_8_442_735_0,
    i_8_442_770_0, i_8_442_789_0, i_8_442_849_0, i_8_442_857_0,
    i_8_442_875_0, i_8_442_1039_0, i_8_442_1075_0, i_8_442_1093_0,
    i_8_442_1189_0, i_8_442_1190_0, i_8_442_1200_0, i_8_442_1219_0,
    i_8_442_1277_0, i_8_442_1293_0, i_8_442_1297_0, i_8_442_1307_0,
    i_8_442_1348_0, i_8_442_1408_0, i_8_442_1410_0, i_8_442_1437_0,
    i_8_442_1471_0, i_8_442_1487_0, i_8_442_1531_0, i_8_442_1536_0,
    i_8_442_1545_0, i_8_442_1586_0, i_8_442_1624_0, i_8_442_1633_0,
    i_8_442_1634_0, i_8_442_1669_0, i_8_442_1696_0, i_8_442_1704_0,
    i_8_442_1724_0, i_8_442_1739_0, i_8_442_1742_0, i_8_442_1768_0,
    i_8_442_1779_0, i_8_442_1794_0, i_8_442_1795_0, i_8_442_1799_0,
    i_8_442_1874_0, i_8_442_1906_0, i_8_442_1918_0, i_8_442_1957_0,
    i_8_442_1958_0, i_8_442_1965_0, i_8_442_1969_0, i_8_442_1981_0,
    i_8_442_2019_0, i_8_442_2032_0, i_8_442_2116_0, i_8_442_2122_0,
    i_8_442_2149_0, i_8_442_2236_0, i_8_442_2246_0;
  output o_8_442_0_0;
  assign o_8_442_0_0 = 0;
endmodule



// Benchmark "kernel_8_443" written by ABC on Sun Jul 19 10:10:51 2020

module kernel_8_443 ( 
    i_8_443_11_0, i_8_443_48_0, i_8_443_103_0, i_8_443_112_0,
    i_8_443_125_0, i_8_443_134_0, i_8_443_280_0, i_8_443_301_0,
    i_8_443_335_0, i_8_443_349_0, i_8_443_367_0, i_8_443_377_0,
    i_8_443_385_0, i_8_443_390_0, i_8_443_399_0, i_8_443_428_0,
    i_8_443_430_0, i_8_443_454_0, i_8_443_458_0, i_8_443_569_0,
    i_8_443_576_0, i_8_443_588_0, i_8_443_589_0, i_8_443_604_0,
    i_8_443_628_0, i_8_443_653_0, i_8_443_655_0, i_8_443_658_0,
    i_8_443_736_0, i_8_443_819_0, i_8_443_893_0, i_8_443_934_0,
    i_8_443_985_0, i_8_443_988_0, i_8_443_995_0, i_8_443_1033_0,
    i_8_443_1036_0, i_8_443_1043_0, i_8_443_1078_0, i_8_443_1093_0,
    i_8_443_1108_0, i_8_443_1109_0, i_8_443_1180_0, i_8_443_1229_0,
    i_8_443_1232_0, i_8_443_1265_0, i_8_443_1284_0, i_8_443_1285_0,
    i_8_443_1286_0, i_8_443_1315_0, i_8_443_1319_0, i_8_443_1331_0,
    i_8_443_1356_0, i_8_443_1363_0, i_8_443_1399_0, i_8_443_1432_0,
    i_8_443_1459_0, i_8_443_1484_0, i_8_443_1486_0, i_8_443_1514_0,
    i_8_443_1527_0, i_8_443_1528_0, i_8_443_1548_0, i_8_443_1558_0,
    i_8_443_1624_0, i_8_443_1638_0, i_8_443_1652_0, i_8_443_1654_0,
    i_8_443_1658_0, i_8_443_1676_0, i_8_443_1687_0, i_8_443_1706_0,
    i_8_443_1748_0, i_8_443_1749_0, i_8_443_1765_0, i_8_443_1825_0,
    i_8_443_1834_0, i_8_443_1836_0, i_8_443_1837_0, i_8_443_1855_0,
    i_8_443_1860_0, i_8_443_1861_0, i_8_443_1888_0, i_8_443_1902_0,
    i_8_443_1909_0, i_8_443_1980_0, i_8_443_1992_0, i_8_443_2013_0,
    i_8_443_2087_0, i_8_443_2093_0, i_8_443_2101_0, i_8_443_2106_0,
    i_8_443_2132_0, i_8_443_2144_0, i_8_443_2146_0, i_8_443_2147_0,
    i_8_443_2150_0, i_8_443_2224_0, i_8_443_2245_0, i_8_443_2275_0,
    o_8_443_0_0  );
  input  i_8_443_11_0, i_8_443_48_0, i_8_443_103_0, i_8_443_112_0,
    i_8_443_125_0, i_8_443_134_0, i_8_443_280_0, i_8_443_301_0,
    i_8_443_335_0, i_8_443_349_0, i_8_443_367_0, i_8_443_377_0,
    i_8_443_385_0, i_8_443_390_0, i_8_443_399_0, i_8_443_428_0,
    i_8_443_430_0, i_8_443_454_0, i_8_443_458_0, i_8_443_569_0,
    i_8_443_576_0, i_8_443_588_0, i_8_443_589_0, i_8_443_604_0,
    i_8_443_628_0, i_8_443_653_0, i_8_443_655_0, i_8_443_658_0,
    i_8_443_736_0, i_8_443_819_0, i_8_443_893_0, i_8_443_934_0,
    i_8_443_985_0, i_8_443_988_0, i_8_443_995_0, i_8_443_1033_0,
    i_8_443_1036_0, i_8_443_1043_0, i_8_443_1078_0, i_8_443_1093_0,
    i_8_443_1108_0, i_8_443_1109_0, i_8_443_1180_0, i_8_443_1229_0,
    i_8_443_1232_0, i_8_443_1265_0, i_8_443_1284_0, i_8_443_1285_0,
    i_8_443_1286_0, i_8_443_1315_0, i_8_443_1319_0, i_8_443_1331_0,
    i_8_443_1356_0, i_8_443_1363_0, i_8_443_1399_0, i_8_443_1432_0,
    i_8_443_1459_0, i_8_443_1484_0, i_8_443_1486_0, i_8_443_1514_0,
    i_8_443_1527_0, i_8_443_1528_0, i_8_443_1548_0, i_8_443_1558_0,
    i_8_443_1624_0, i_8_443_1638_0, i_8_443_1652_0, i_8_443_1654_0,
    i_8_443_1658_0, i_8_443_1676_0, i_8_443_1687_0, i_8_443_1706_0,
    i_8_443_1748_0, i_8_443_1749_0, i_8_443_1765_0, i_8_443_1825_0,
    i_8_443_1834_0, i_8_443_1836_0, i_8_443_1837_0, i_8_443_1855_0,
    i_8_443_1860_0, i_8_443_1861_0, i_8_443_1888_0, i_8_443_1902_0,
    i_8_443_1909_0, i_8_443_1980_0, i_8_443_1992_0, i_8_443_2013_0,
    i_8_443_2087_0, i_8_443_2093_0, i_8_443_2101_0, i_8_443_2106_0,
    i_8_443_2132_0, i_8_443_2144_0, i_8_443_2146_0, i_8_443_2147_0,
    i_8_443_2150_0, i_8_443_2224_0, i_8_443_2245_0, i_8_443_2275_0;
  output o_8_443_0_0;
  assign o_8_443_0_0 = 0;
endmodule



// Benchmark "kernel_8_444" written by ABC on Sun Jul 19 10:10:52 2020

module kernel_8_444 ( 
    i_8_444_31_0, i_8_444_70_0, i_8_444_89_0, i_8_444_96_0, i_8_444_191_0,
    i_8_444_194_0, i_8_444_204_0, i_8_444_205_0, i_8_444_292_0,
    i_8_444_293_0, i_8_444_311_0, i_8_444_328_0, i_8_444_343_0,
    i_8_444_358_0, i_8_444_376_0, i_8_444_383_0, i_8_444_422_0,
    i_8_444_456_0, i_8_444_477_0, i_8_444_552_0, i_8_444_587_0,
    i_8_444_596_0, i_8_444_601_0, i_8_444_609_0, i_8_444_610_0,
    i_8_444_613_0, i_8_444_619_0, i_8_444_672_0, i_8_444_760_0,
    i_8_444_772_0, i_8_444_780_0, i_8_444_818_0, i_8_444_874_0,
    i_8_444_875_0, i_8_444_877_0, i_8_444_898_0, i_8_444_899_0,
    i_8_444_916_0, i_8_444_946_0, i_8_444_951_0, i_8_444_976_0,
    i_8_444_985_0, i_8_444_987_0, i_8_444_989_0, i_8_444_1030_0,
    i_8_444_1108_0, i_8_444_1110_0, i_8_444_1132_0, i_8_444_1141_0,
    i_8_444_1194_0, i_8_444_1223_0, i_8_444_1256_0, i_8_444_1257_0,
    i_8_444_1259_0, i_8_444_1262_0, i_8_444_1277_0, i_8_444_1281_0,
    i_8_444_1284_0, i_8_444_1430_0, i_8_444_1438_0, i_8_444_1455_0,
    i_8_444_1471_0, i_8_444_1483_0, i_8_444_1484_0, i_8_444_1527_0,
    i_8_444_1552_0, i_8_444_1553_0, i_8_444_1558_0, i_8_444_1582_0,
    i_8_444_1603_0, i_8_444_1606_0, i_8_444_1637_0, i_8_444_1672_0,
    i_8_444_1680_0, i_8_444_1699_0, i_8_444_1734_0, i_8_444_1735_0,
    i_8_444_1743_0, i_8_444_1745_0, i_8_444_1775_0, i_8_444_1779_0,
    i_8_444_1784_0, i_8_444_1788_0, i_8_444_1797_0, i_8_444_1815_0,
    i_8_444_1821_0, i_8_444_1822_0, i_8_444_1823_0, i_8_444_1839_0,
    i_8_444_1855_0, i_8_444_1867_0, i_8_444_1964_0, i_8_444_1982_0,
    i_8_444_2013_0, i_8_444_2014_0, i_8_444_2050_0, i_8_444_2108_0,
    i_8_444_2130_0, i_8_444_2193_0, i_8_444_2290_0,
    o_8_444_0_0  );
  input  i_8_444_31_0, i_8_444_70_0, i_8_444_89_0, i_8_444_96_0,
    i_8_444_191_0, i_8_444_194_0, i_8_444_204_0, i_8_444_205_0,
    i_8_444_292_0, i_8_444_293_0, i_8_444_311_0, i_8_444_328_0,
    i_8_444_343_0, i_8_444_358_0, i_8_444_376_0, i_8_444_383_0,
    i_8_444_422_0, i_8_444_456_0, i_8_444_477_0, i_8_444_552_0,
    i_8_444_587_0, i_8_444_596_0, i_8_444_601_0, i_8_444_609_0,
    i_8_444_610_0, i_8_444_613_0, i_8_444_619_0, i_8_444_672_0,
    i_8_444_760_0, i_8_444_772_0, i_8_444_780_0, i_8_444_818_0,
    i_8_444_874_0, i_8_444_875_0, i_8_444_877_0, i_8_444_898_0,
    i_8_444_899_0, i_8_444_916_0, i_8_444_946_0, i_8_444_951_0,
    i_8_444_976_0, i_8_444_985_0, i_8_444_987_0, i_8_444_989_0,
    i_8_444_1030_0, i_8_444_1108_0, i_8_444_1110_0, i_8_444_1132_0,
    i_8_444_1141_0, i_8_444_1194_0, i_8_444_1223_0, i_8_444_1256_0,
    i_8_444_1257_0, i_8_444_1259_0, i_8_444_1262_0, i_8_444_1277_0,
    i_8_444_1281_0, i_8_444_1284_0, i_8_444_1430_0, i_8_444_1438_0,
    i_8_444_1455_0, i_8_444_1471_0, i_8_444_1483_0, i_8_444_1484_0,
    i_8_444_1527_0, i_8_444_1552_0, i_8_444_1553_0, i_8_444_1558_0,
    i_8_444_1582_0, i_8_444_1603_0, i_8_444_1606_0, i_8_444_1637_0,
    i_8_444_1672_0, i_8_444_1680_0, i_8_444_1699_0, i_8_444_1734_0,
    i_8_444_1735_0, i_8_444_1743_0, i_8_444_1745_0, i_8_444_1775_0,
    i_8_444_1779_0, i_8_444_1784_0, i_8_444_1788_0, i_8_444_1797_0,
    i_8_444_1815_0, i_8_444_1821_0, i_8_444_1822_0, i_8_444_1823_0,
    i_8_444_1839_0, i_8_444_1855_0, i_8_444_1867_0, i_8_444_1964_0,
    i_8_444_1982_0, i_8_444_2013_0, i_8_444_2014_0, i_8_444_2050_0,
    i_8_444_2108_0, i_8_444_2130_0, i_8_444_2193_0, i_8_444_2290_0;
  output o_8_444_0_0;
  assign o_8_444_0_0 = 0;
endmodule



// Benchmark "kernel_8_445" written by ABC on Sun Jul 19 10:10:54 2020

module kernel_8_445 ( 
    i_8_445_7_0, i_8_445_18_0, i_8_445_59_0, i_8_445_112_0, i_8_445_136_0,
    i_8_445_142_0, i_8_445_154_0, i_8_445_162_0, i_8_445_163_0,
    i_8_445_220_0, i_8_445_222_0, i_8_445_225_0, i_8_445_300_0,
    i_8_445_330_0, i_8_445_378_0, i_8_445_382_0, i_8_445_493_0,
    i_8_445_516_0, i_8_445_522_0, i_8_445_530_0, i_8_445_576_0,
    i_8_445_580_0, i_8_445_589_0, i_8_445_590_0, i_8_445_600_0,
    i_8_445_628_0, i_8_445_631_0, i_8_445_639_0, i_8_445_640_0,
    i_8_445_648_0, i_8_445_649_0, i_8_445_658_0, i_8_445_675_0,
    i_8_445_693_0, i_8_445_694_0, i_8_445_703_0, i_8_445_708_0,
    i_8_445_729_0, i_8_445_747_0, i_8_445_748_0, i_8_445_820_0,
    i_8_445_829_0, i_8_445_877_0, i_8_445_886_0, i_8_445_956_0,
    i_8_445_973_0, i_8_445_990_0, i_8_445_993_0, i_8_445_999_0,
    i_8_445_1034_0, i_8_445_1107_0, i_8_445_1108_0, i_8_445_1125_0,
    i_8_445_1152_0, i_8_445_1156_0, i_8_445_1161_0, i_8_445_1162_0,
    i_8_445_1261_0, i_8_445_1275_0, i_8_445_1327_0, i_8_445_1335_0,
    i_8_445_1352_0, i_8_445_1355_0, i_8_445_1407_0, i_8_445_1433_0,
    i_8_445_1485_0, i_8_445_1486_0, i_8_445_1530_0, i_8_445_1593_0,
    i_8_445_1596_0, i_8_445_1609_0, i_8_445_1656_0, i_8_445_1659_0,
    i_8_445_1680_0, i_8_445_1681_0, i_8_445_1753_0, i_8_445_1773_0,
    i_8_445_1784_0, i_8_445_1804_0, i_8_445_1818_0, i_8_445_1819_0,
    i_8_445_1852_0, i_8_445_1853_0, i_8_445_1971_0, i_8_445_1972_0,
    i_8_445_1992_0, i_8_445_2007_0, i_8_445_2008_0, i_8_445_2043_0,
    i_8_445_2088_0, i_8_445_2089_0, i_8_445_2093_0, i_8_445_2098_0,
    i_8_445_2123_0, i_8_445_2145_0, i_8_445_2170_0, i_8_445_2206_0,
    i_8_445_2226_0, i_8_445_2253_0, i_8_445_2254_0,
    o_8_445_0_0  );
  input  i_8_445_7_0, i_8_445_18_0, i_8_445_59_0, i_8_445_112_0,
    i_8_445_136_0, i_8_445_142_0, i_8_445_154_0, i_8_445_162_0,
    i_8_445_163_0, i_8_445_220_0, i_8_445_222_0, i_8_445_225_0,
    i_8_445_300_0, i_8_445_330_0, i_8_445_378_0, i_8_445_382_0,
    i_8_445_493_0, i_8_445_516_0, i_8_445_522_0, i_8_445_530_0,
    i_8_445_576_0, i_8_445_580_0, i_8_445_589_0, i_8_445_590_0,
    i_8_445_600_0, i_8_445_628_0, i_8_445_631_0, i_8_445_639_0,
    i_8_445_640_0, i_8_445_648_0, i_8_445_649_0, i_8_445_658_0,
    i_8_445_675_0, i_8_445_693_0, i_8_445_694_0, i_8_445_703_0,
    i_8_445_708_0, i_8_445_729_0, i_8_445_747_0, i_8_445_748_0,
    i_8_445_820_0, i_8_445_829_0, i_8_445_877_0, i_8_445_886_0,
    i_8_445_956_0, i_8_445_973_0, i_8_445_990_0, i_8_445_993_0,
    i_8_445_999_0, i_8_445_1034_0, i_8_445_1107_0, i_8_445_1108_0,
    i_8_445_1125_0, i_8_445_1152_0, i_8_445_1156_0, i_8_445_1161_0,
    i_8_445_1162_0, i_8_445_1261_0, i_8_445_1275_0, i_8_445_1327_0,
    i_8_445_1335_0, i_8_445_1352_0, i_8_445_1355_0, i_8_445_1407_0,
    i_8_445_1433_0, i_8_445_1485_0, i_8_445_1486_0, i_8_445_1530_0,
    i_8_445_1593_0, i_8_445_1596_0, i_8_445_1609_0, i_8_445_1656_0,
    i_8_445_1659_0, i_8_445_1680_0, i_8_445_1681_0, i_8_445_1753_0,
    i_8_445_1773_0, i_8_445_1784_0, i_8_445_1804_0, i_8_445_1818_0,
    i_8_445_1819_0, i_8_445_1852_0, i_8_445_1853_0, i_8_445_1971_0,
    i_8_445_1972_0, i_8_445_1992_0, i_8_445_2007_0, i_8_445_2008_0,
    i_8_445_2043_0, i_8_445_2088_0, i_8_445_2089_0, i_8_445_2093_0,
    i_8_445_2098_0, i_8_445_2123_0, i_8_445_2145_0, i_8_445_2170_0,
    i_8_445_2206_0, i_8_445_2226_0, i_8_445_2253_0, i_8_445_2254_0;
  output o_8_445_0_0;
  assign o_8_445_0_0 = ~((~i_8_445_516_0 & ((~i_8_445_112_0 & ((~i_8_445_225_0 & ~i_8_445_628_0 & ~i_8_445_829_0 & ~i_8_445_2007_0 & ~i_8_445_2008_0 & ~i_8_445_2088_0 & ~i_8_445_2123_0) | (~i_8_445_648_0 & ~i_8_445_703_0 & ~i_8_445_1596_0 & ~i_8_445_1656_0 & ~i_8_445_1819_0 & ~i_8_445_2170_0 & ~i_8_445_2253_0))) | (~i_8_445_162_0 & ~i_8_445_747_0 & ~i_8_445_990_0 & ~i_8_445_1407_0 & ~i_8_445_1659_0 & i_8_445_1818_0))) | (~i_8_445_493_0 & ((~i_8_445_631_0 & ~i_8_445_729_0 & ~i_8_445_973_0 & ~i_8_445_1161_0 & ~i_8_445_1162_0 & ~i_8_445_1355_0 & ~i_8_445_1593_0 & ~i_8_445_1596_0 & ~i_8_445_1609_0 & ~i_8_445_2007_0) | (~i_8_445_300_0 & ~i_8_445_829_0 & ~i_8_445_877_0 & i_8_445_1125_0 & ~i_8_445_1275_0 & ~i_8_445_1352_0 & ~i_8_445_1784_0 & i_8_445_2089_0 & ~i_8_445_2253_0))) | (~i_8_445_1162_0 & ((~i_8_445_649_0 & ((~i_8_445_648_0 & ~i_8_445_1593_0 & ~i_8_445_1753_0 & ~i_8_445_1992_0 & ~i_8_445_2089_0) | (~i_8_445_1161_0 & ~i_8_445_1609_0 & ~i_8_445_1659_0 & ~i_8_445_2007_0 & ~i_8_445_2226_0 & ~i_8_445_2254_0))) | (~i_8_445_7_0 & ~i_8_445_136_0 & ~i_8_445_382_0 & i_8_445_522_0 & ~i_8_445_693_0 & ~i_8_445_729_0 & ~i_8_445_1355_0 & ~i_8_445_1593_0 & ~i_8_445_1773_0) | (i_8_445_820_0 & i_8_445_877_0 & ~i_8_445_1609_0 & ~i_8_445_2088_0) | (~i_8_445_163_0 & i_8_445_222_0 & ~i_8_445_1656_0 & ~i_8_445_2123_0 & ~i_8_445_2145_0))) | (~i_8_445_747_0 & ((~i_8_445_829_0 & ((~i_8_445_530_0 & ~i_8_445_631_0 & ~i_8_445_1355_0 & ~i_8_445_1656_0 & i_8_445_1753_0) | (~i_8_445_877_0 & ~i_8_445_1659_0 & i_8_445_1818_0 & ~i_8_445_1853_0 & ~i_8_445_2008_0 & ~i_8_445_2253_0))) | (~i_8_445_1992_0 & ((i_8_445_649_0 & ~i_8_445_675_0 & i_8_445_1261_0 & ~i_8_445_1275_0 & ~i_8_445_2088_0) | (~i_8_445_330_0 & ~i_8_445_658_0 & ~i_8_445_820_0 & ~i_8_445_877_0 & ~i_8_445_956_0 & i_8_445_1853_0 & i_8_445_2098_0))) | (~i_8_445_154_0 & i_8_445_589_0 & ~i_8_445_693_0 & ~i_8_445_729_0 & ~i_8_445_1107_0 & ~i_8_445_2123_0))) | (~i_8_445_693_0 & ~i_8_445_2253_0 & ((i_8_445_154_0 & ~i_8_445_703_0 & ~i_8_445_729_0 & ~i_8_445_1355_0) | (~i_8_445_1486_0 & ~i_8_445_1530_0 & ~i_8_445_1593_0 & ~i_8_445_1853_0 & ~i_8_445_2089_0))) | (~i_8_445_829_0 & ~i_8_445_2254_0 & ((~i_8_445_225_0 & i_8_445_648_0 & ~i_8_445_1161_0 & ~i_8_445_1530_0) | (~i_8_445_18_0 & ~i_8_445_729_0 & ~i_8_445_990_0 & ~i_8_445_1656_0 & ~i_8_445_1680_0 & ~i_8_445_2008_0))) | (~i_8_445_1161_0 & ((~i_8_445_220_0 & ~i_8_445_1125_0 & ~i_8_445_1596_0 & ~i_8_445_1659_0 & ~i_8_445_1773_0 & ~i_8_445_1819_0 & ~i_8_445_1992_0 & ~i_8_445_2093_0) | (~i_8_445_600_0 & ~i_8_445_694_0 & ~i_8_445_1034_0 & ~i_8_445_1485_0 & ~i_8_445_1486_0 & ~i_8_445_1530_0 & ~i_8_445_1681_0 & ~i_8_445_1753_0 & ~i_8_445_1852_0 & ~i_8_445_2170_0))) | (~i_8_445_1656_0 & i_8_445_1992_0 & ~i_8_445_2008_0 & ((i_8_445_300_0 & ~i_8_445_1804_0 & ~i_8_445_2089_0) | (~i_8_445_1593_0 & ~i_8_445_1596_0 & ~i_8_445_1659_0 & ~i_8_445_2007_0 & ~i_8_445_2093_0 & i_8_445_2145_0))) | (i_8_445_576_0 & i_8_445_1275_0) | (~i_8_445_748_0 & ~i_8_445_1659_0 & i_8_445_1681_0 & ~i_8_445_1773_0 & ~i_8_445_2145_0));
endmodule



// Benchmark "kernel_8_446" written by ABC on Sun Jul 19 10:10:55 2020

module kernel_8_446 ( 
    i_8_446_10_0, i_8_446_114_0, i_8_446_115_0, i_8_446_120_0,
    i_8_446_121_0, i_8_446_125_0, i_8_446_171_0, i_8_446_193_0,
    i_8_446_196_0, i_8_446_223_0, i_8_446_232_0, i_8_446_292_0,
    i_8_446_349_0, i_8_446_365_0, i_8_446_422_0, i_8_446_426_0,
    i_8_446_472_0, i_8_446_475_0, i_8_446_507_0, i_8_446_556_0,
    i_8_446_572_0, i_8_446_602_0, i_8_446_625_0, i_8_446_679_0,
    i_8_446_696_0, i_8_446_698_0, i_8_446_724_0, i_8_446_732_0,
    i_8_446_784_0, i_8_446_787_0, i_8_446_814_0, i_8_446_832_0,
    i_8_446_843_0, i_8_446_862_0, i_8_446_877_0, i_8_446_885_0,
    i_8_446_930_0, i_8_446_967_0, i_8_446_976_0, i_8_446_984_0,
    i_8_446_994_0, i_8_446_995_0, i_8_446_1003_0, i_8_446_1030_0,
    i_8_446_1040_0, i_8_446_1047_0, i_8_446_1057_0, i_8_446_1126_0,
    i_8_446_1179_0, i_8_446_1281_0, i_8_446_1315_0, i_8_446_1355_0,
    i_8_446_1372_0, i_8_446_1436_0, i_8_446_1453_0, i_8_446_1456_0,
    i_8_446_1484_0, i_8_446_1551_0, i_8_446_1553_0, i_8_446_1623_0,
    i_8_446_1624_0, i_8_446_1642_0, i_8_446_1650_0, i_8_446_1651_0,
    i_8_446_1652_0, i_8_446_1653_0, i_8_446_1655_0, i_8_446_1663_0,
    i_8_446_1696_0, i_8_446_1697_0, i_8_446_1699_0, i_8_446_1747_0,
    i_8_446_1767_0, i_8_446_1771_0, i_8_446_1804_0, i_8_446_1808_0,
    i_8_446_1821_0, i_8_446_1823_0, i_8_446_1826_0, i_8_446_1839_0,
    i_8_446_1867_0, i_8_446_1893_0, i_8_446_1967_0, i_8_446_1992_0,
    i_8_446_2073_0, i_8_446_2096_0, i_8_446_2100_0, i_8_446_2101_0,
    i_8_446_2109_0, i_8_446_2119_0, i_8_446_2126_0, i_8_446_2128_0,
    i_8_446_2134_0, i_8_446_2172_0, i_8_446_2173_0, i_8_446_2176_0,
    i_8_446_2230_0, i_8_446_2244_0, i_8_446_2245_0, i_8_446_2258_0,
    o_8_446_0_0  );
  input  i_8_446_10_0, i_8_446_114_0, i_8_446_115_0, i_8_446_120_0,
    i_8_446_121_0, i_8_446_125_0, i_8_446_171_0, i_8_446_193_0,
    i_8_446_196_0, i_8_446_223_0, i_8_446_232_0, i_8_446_292_0,
    i_8_446_349_0, i_8_446_365_0, i_8_446_422_0, i_8_446_426_0,
    i_8_446_472_0, i_8_446_475_0, i_8_446_507_0, i_8_446_556_0,
    i_8_446_572_0, i_8_446_602_0, i_8_446_625_0, i_8_446_679_0,
    i_8_446_696_0, i_8_446_698_0, i_8_446_724_0, i_8_446_732_0,
    i_8_446_784_0, i_8_446_787_0, i_8_446_814_0, i_8_446_832_0,
    i_8_446_843_0, i_8_446_862_0, i_8_446_877_0, i_8_446_885_0,
    i_8_446_930_0, i_8_446_967_0, i_8_446_976_0, i_8_446_984_0,
    i_8_446_994_0, i_8_446_995_0, i_8_446_1003_0, i_8_446_1030_0,
    i_8_446_1040_0, i_8_446_1047_0, i_8_446_1057_0, i_8_446_1126_0,
    i_8_446_1179_0, i_8_446_1281_0, i_8_446_1315_0, i_8_446_1355_0,
    i_8_446_1372_0, i_8_446_1436_0, i_8_446_1453_0, i_8_446_1456_0,
    i_8_446_1484_0, i_8_446_1551_0, i_8_446_1553_0, i_8_446_1623_0,
    i_8_446_1624_0, i_8_446_1642_0, i_8_446_1650_0, i_8_446_1651_0,
    i_8_446_1652_0, i_8_446_1653_0, i_8_446_1655_0, i_8_446_1663_0,
    i_8_446_1696_0, i_8_446_1697_0, i_8_446_1699_0, i_8_446_1747_0,
    i_8_446_1767_0, i_8_446_1771_0, i_8_446_1804_0, i_8_446_1808_0,
    i_8_446_1821_0, i_8_446_1823_0, i_8_446_1826_0, i_8_446_1839_0,
    i_8_446_1867_0, i_8_446_1893_0, i_8_446_1967_0, i_8_446_1992_0,
    i_8_446_2073_0, i_8_446_2096_0, i_8_446_2100_0, i_8_446_2101_0,
    i_8_446_2109_0, i_8_446_2119_0, i_8_446_2126_0, i_8_446_2128_0,
    i_8_446_2134_0, i_8_446_2172_0, i_8_446_2173_0, i_8_446_2176_0,
    i_8_446_2230_0, i_8_446_2244_0, i_8_446_2245_0, i_8_446_2258_0;
  output o_8_446_0_0;
  assign o_8_446_0_0 = 0;
endmodule



// Benchmark "kernel_8_447" written by ABC on Sun Jul 19 10:10:56 2020

module kernel_8_447 ( 
    i_8_447_138_0, i_8_447_232_0, i_8_447_233_0, i_8_447_360_0,
    i_8_447_361_0, i_8_447_365_0, i_8_447_366_0, i_8_447_368_0,
    i_8_447_372_0, i_8_447_378_0, i_8_447_382_0, i_8_447_422_0,
    i_8_447_426_0, i_8_447_427_0, i_8_447_428_0, i_8_447_474_0,
    i_8_447_477_0, i_8_447_478_0, i_8_447_479_0, i_8_447_480_0,
    i_8_447_482_0, i_8_447_492_0, i_8_447_493_0, i_8_447_592_0,
    i_8_447_612_0, i_8_447_670_0, i_8_447_671_0, i_8_447_673_0,
    i_8_447_674_0, i_8_447_684_0, i_8_447_687_0, i_8_447_689_0,
    i_8_447_691_0, i_8_447_695_0, i_8_447_696_0, i_8_447_697_0,
    i_8_447_703_0, i_8_447_704_0, i_8_447_757_0, i_8_447_758_0,
    i_8_447_763_0, i_8_447_837_0, i_8_447_838_0, i_8_447_839_0,
    i_8_447_878_0, i_8_447_955_0, i_8_447_1060_0, i_8_447_1079_0,
    i_8_447_1129_0, i_8_447_1132_0, i_8_447_1159_0, i_8_447_1185_0,
    i_8_447_1224_0, i_8_447_1226_0, i_8_447_1231_0, i_8_447_1273_0,
    i_8_447_1282_0, i_8_447_1303_0, i_8_447_1305_0, i_8_447_1306_0,
    i_8_447_1307_0, i_8_447_1332_0, i_8_447_1352_0, i_8_447_1456_0,
    i_8_447_1477_0, i_8_447_1552_0, i_8_447_1587_0, i_8_447_1719_0,
    i_8_447_1720_0, i_8_447_1722_0, i_8_447_1737_0, i_8_447_1740_0,
    i_8_447_1746_0, i_8_447_1807_0, i_8_447_1808_0, i_8_447_1818_0,
    i_8_447_1820_0, i_8_447_1821_0, i_8_447_1824_0, i_8_447_1832_0,
    i_8_447_1902_0, i_8_447_1951_0, i_8_447_1967_0, i_8_447_1981_0,
    i_8_447_1985_0, i_8_447_2143_0, i_8_447_2149_0, i_8_447_2150_0,
    i_8_447_2223_0, i_8_447_2226_0, i_8_447_2229_0, i_8_447_2272_0,
    i_8_447_2275_0, i_8_447_2276_0, i_8_447_2289_0, i_8_447_2290_0,
    i_8_447_2299_0, i_8_447_2300_0, i_8_447_2301_0, i_8_447_2303_0,
    o_8_447_0_0  );
  input  i_8_447_138_0, i_8_447_232_0, i_8_447_233_0, i_8_447_360_0,
    i_8_447_361_0, i_8_447_365_0, i_8_447_366_0, i_8_447_368_0,
    i_8_447_372_0, i_8_447_378_0, i_8_447_382_0, i_8_447_422_0,
    i_8_447_426_0, i_8_447_427_0, i_8_447_428_0, i_8_447_474_0,
    i_8_447_477_0, i_8_447_478_0, i_8_447_479_0, i_8_447_480_0,
    i_8_447_482_0, i_8_447_492_0, i_8_447_493_0, i_8_447_592_0,
    i_8_447_612_0, i_8_447_670_0, i_8_447_671_0, i_8_447_673_0,
    i_8_447_674_0, i_8_447_684_0, i_8_447_687_0, i_8_447_689_0,
    i_8_447_691_0, i_8_447_695_0, i_8_447_696_0, i_8_447_697_0,
    i_8_447_703_0, i_8_447_704_0, i_8_447_757_0, i_8_447_758_0,
    i_8_447_763_0, i_8_447_837_0, i_8_447_838_0, i_8_447_839_0,
    i_8_447_878_0, i_8_447_955_0, i_8_447_1060_0, i_8_447_1079_0,
    i_8_447_1129_0, i_8_447_1132_0, i_8_447_1159_0, i_8_447_1185_0,
    i_8_447_1224_0, i_8_447_1226_0, i_8_447_1231_0, i_8_447_1273_0,
    i_8_447_1282_0, i_8_447_1303_0, i_8_447_1305_0, i_8_447_1306_0,
    i_8_447_1307_0, i_8_447_1332_0, i_8_447_1352_0, i_8_447_1456_0,
    i_8_447_1477_0, i_8_447_1552_0, i_8_447_1587_0, i_8_447_1719_0,
    i_8_447_1720_0, i_8_447_1722_0, i_8_447_1737_0, i_8_447_1740_0,
    i_8_447_1746_0, i_8_447_1807_0, i_8_447_1808_0, i_8_447_1818_0,
    i_8_447_1820_0, i_8_447_1821_0, i_8_447_1824_0, i_8_447_1832_0,
    i_8_447_1902_0, i_8_447_1951_0, i_8_447_1967_0, i_8_447_1981_0,
    i_8_447_1985_0, i_8_447_2143_0, i_8_447_2149_0, i_8_447_2150_0,
    i_8_447_2223_0, i_8_447_2226_0, i_8_447_2229_0, i_8_447_2272_0,
    i_8_447_2275_0, i_8_447_2276_0, i_8_447_2289_0, i_8_447_2290_0,
    i_8_447_2299_0, i_8_447_2300_0, i_8_447_2301_0, i_8_447_2303_0;
  output o_8_447_0_0;
  assign o_8_447_0_0 = ~((i_8_447_361_0 & ((~i_8_447_684_0 & ~i_8_447_687_0 & ~i_8_447_1719_0 & ~i_8_447_1722_0 & ~i_8_447_1832_0 & i_8_447_2143_0) | (~i_8_447_480_0 & ~i_8_447_757_0 & ~i_8_447_1737_0 & ~i_8_447_1985_0 & ~i_8_447_2300_0))) | (~i_8_447_138_0 & ((~i_8_447_372_0 & ((~i_8_447_378_0 & ~i_8_447_477_0 & ~i_8_447_479_0 & ~i_8_447_687_0 & ~i_8_447_697_0 & ~i_8_447_763_0 & ~i_8_447_1746_0 & ~i_8_447_1818_0 & ~i_8_447_1985_0 & i_8_447_2290_0) | (~i_8_447_428_0 & ~i_8_447_1552_0 & i_8_447_2150_0 & ~i_8_447_2276_0 & ~i_8_447_2299_0 & ~i_8_447_2301_0 & ~i_8_447_2303_0))) | (~i_8_447_689_0 & ((~i_8_447_684_0 & ~i_8_447_878_0 & ~i_8_447_1746_0 & i_8_447_1820_0 & ~i_8_447_1824_0) | (~i_8_447_479_0 & i_8_447_839_0 & ~i_8_447_1332_0 & ~i_8_447_1720_0 & ~i_8_447_1820_0 & ~i_8_447_1967_0 & ~i_8_447_2303_0))) | (~i_8_447_482_0 & ((~i_8_447_479_0 & ~i_8_447_691_0 & ((~i_8_447_360_0 & ~i_8_447_422_0 & ~i_8_447_478_0 & ~i_8_447_684_0 & ~i_8_447_1282_0 & i_8_447_1552_0 & ~i_8_447_1587_0 & ~i_8_447_1985_0) | (~i_8_447_757_0 & ~i_8_447_1273_0 & i_8_447_2143_0 & ~i_8_447_2223_0))) | (~i_8_447_474_0 & ~i_8_447_684_0 & i_8_447_696_0 & ~i_8_447_1282_0 & ~i_8_447_1332_0 & ~i_8_447_1981_0 & ~i_8_447_2301_0))) | (~i_8_447_1303_0 & ((i_8_447_366_0 & ~i_8_447_382_0 & ~i_8_447_1719_0 & ~i_8_447_1740_0 & ~i_8_447_1951_0) | (~i_8_447_368_0 & i_8_447_427_0 & ~i_8_447_757_0 & ~i_8_447_1552_0 & ~i_8_447_1587_0 & ~i_8_447_2303_0))))) | (i_8_447_378_0 & ((~i_8_447_474_0 & i_8_447_696_0 & ~i_8_447_1740_0 & ~i_8_447_1981_0 & ~i_8_447_2149_0) | (~i_8_447_689_0 & ~i_8_447_1079_0 & i_8_447_1129_0 & ~i_8_447_1307_0 & ~i_8_447_1818_0 & ~i_8_447_2299_0 & ~i_8_447_2301_0))) | (~i_8_447_2299_0 & ((i_8_447_478_0 & ((~i_8_447_480_0 & ~i_8_447_763_0 & i_8_447_1129_0 & ~i_8_447_1720_0) | (~i_8_447_479_0 & ~i_8_447_673_0 & ~i_8_447_1306_0 & ~i_8_447_1818_0 & ~i_8_447_1902_0 & i_8_447_2226_0 & ~i_8_447_2301_0))) | (~i_8_447_233_0 & ~i_8_447_382_0 & ~i_8_447_427_0 & ~i_8_447_428_0 & ~i_8_447_493_0 & ~i_8_447_691_0 & i_8_447_697_0 & ~i_8_447_1720_0 & ~i_8_447_1737_0 & ~i_8_447_1807_0 & ~i_8_447_1967_0 & ~i_8_447_1985_0 & ~i_8_447_2149_0) | (~i_8_447_763_0 & ~i_8_447_1456_0 & i_8_447_2275_0))) | (~i_8_447_479_0 & ((~i_8_447_233_0 & ((i_8_447_382_0 & ~i_8_447_477_0 & ~i_8_447_492_0 & ~i_8_447_687_0 & ~i_8_447_691_0 & ~i_8_447_697_0 & ~i_8_447_1129_0 & ~i_8_447_1273_0 & i_8_447_1282_0 & ~i_8_447_1303_0) | (i_8_447_365_0 & ~i_8_447_838_0 & ~i_8_447_1079_0 & ~i_8_447_1456_0 & ~i_8_447_1720_0 & ~i_8_447_1722_0 & ~i_8_447_1746_0 & ~i_8_447_2300_0))) | (~i_8_447_478_0 & ((~i_8_447_477_0 & ~i_8_447_1332_0 & ((~i_8_447_360_0 & ~i_8_447_687_0 & ~i_8_447_689_0 & i_8_447_838_0 & ~i_8_447_1185_0 & ~i_8_447_1737_0) | (~i_8_447_592_0 & ~i_8_447_696_0 & ~i_8_447_1722_0 & i_8_447_1818_0))) | (i_8_447_1224_0 & ~i_8_447_1740_0) | (~i_8_447_382_0 & i_8_447_592_0 & ~i_8_447_689_0 & ~i_8_447_691_0 & ~i_8_447_1587_0 & ~i_8_447_1746_0 & ~i_8_447_1967_0 & ~i_8_447_2300_0))) | (~i_8_447_757_0 & ((~i_8_447_482_0 & ~i_8_447_689_0 & ((i_8_447_428_0 & ~i_8_447_763_0 & ~i_8_447_1552_0 & ~i_8_447_1807_0 & ~i_8_447_2275_0) | (i_8_447_426_0 & ~i_8_447_474_0 & ~i_8_447_492_0 & ~i_8_447_687_0 & ~i_8_447_691_0 & ~i_8_447_839_0 & ~i_8_447_1722_0 & ~i_8_447_2226_0 & ~i_8_447_2301_0))) | (~i_8_447_378_0 & ~i_8_447_422_0 & ~i_8_447_480_0 & i_8_447_592_0 & ~i_8_447_691_0 & ~i_8_447_1079_0 & ~i_8_447_1719_0 & ~i_8_447_1832_0 & ~i_8_447_1967_0 & ~i_8_447_2290_0))) | (i_8_447_427_0 & ~i_8_447_758_0 & ~i_8_447_1282_0 & i_8_447_1552_0 & ~i_8_447_1746_0 & ~i_8_447_2303_0))) | (~i_8_447_360_0 & ((~i_8_447_592_0 & ~i_8_447_687_0 & ~i_8_447_763_0 & ~i_8_447_1060_0 & i_8_447_1824_0 & ~i_8_447_1902_0) | (i_8_447_382_0 & ~i_8_447_478_0 & ~i_8_447_758_0 & ~i_8_447_1306_0 & ~i_8_447_1820_0 & i_8_447_1967_0 & ~i_8_447_2300_0 & ~i_8_447_2301_0))) | (i_8_447_365_0 & ((i_8_447_838_0 & ~i_8_447_1587_0 & i_8_447_1820_0) | (~i_8_447_482_0 & ~i_8_447_757_0 & ~i_8_447_1967_0 & i_8_447_1985_0 & ~i_8_447_2149_0))) | (~i_8_447_691_0 & ((i_8_447_426_0 & ((~i_8_447_478_0 & ~i_8_447_1231_0 & ~i_8_447_1477_0 & i_8_447_1587_0 & ~i_8_447_1722_0) | (~i_8_447_670_0 & ~i_8_447_1352_0 & ~i_8_447_1587_0 & ~i_8_447_1737_0 & ~i_8_447_1740_0 & i_8_447_1824_0))) | (~i_8_447_477_0 & ((~i_8_447_482_0 & i_8_447_839_0 & i_8_447_1552_0 & i_8_447_1967_0) | (i_8_447_763_0 & ~i_8_447_1719_0 & i_8_447_2276_0))) | (~i_8_447_366_0 & i_8_447_493_0 & ~i_8_447_1332_0 & i_8_447_1552_0 & ~i_8_447_1740_0 & ~i_8_447_1832_0))) | (i_8_447_366_0 & ((~i_8_447_474_0 & ((~i_8_447_670_0 & ~i_8_447_684_0 & i_8_447_691_0 & ~i_8_447_878_0 & ~i_8_447_1746_0 & ~i_8_447_2229_0) | (~i_8_447_592_0 & i_8_447_670_0 & ~i_8_447_687_0 & ~i_8_447_1303_0 & ~i_8_447_1902_0 & ~i_8_447_2301_0))) | (i_8_447_480_0 & ~i_8_447_612_0 & i_8_447_1552_0 & ~i_8_447_1720_0 & ~i_8_447_1824_0))) | (i_8_447_493_0 & ((~i_8_447_482_0 & i_8_447_2276_0) | (~i_8_447_480_0 & ~i_8_447_670_0 & ~i_8_447_1306_0 & ~i_8_447_1722_0 & i_8_447_2290_0))) | (~i_8_447_482_0 & ((i_8_447_382_0 & i_8_447_671_0 & i_8_447_691_0 & ~i_8_447_1060_0) | (~i_8_447_878_0 & ~i_8_447_1185_0 & ~i_8_447_1282_0 & i_8_447_1807_0 & ~i_8_447_2290_0 & ~i_8_447_2301_0))) | (~i_8_447_689_0 & ((~i_8_447_480_0 & ~i_8_447_1060_0 & ~i_8_447_1185_0 & ~i_8_447_1307_0 & ~i_8_447_1985_0 & i_8_447_2149_0 & i_8_447_2150_0) | (~i_8_447_757_0 & ~i_8_447_1303_0 & i_8_447_2276_0))) | (i_8_447_695_0 & ((i_8_447_704_0 & i_8_447_1820_0) | (~i_8_447_480_0 & i_8_447_1352_0 & ~i_8_447_1720_0 & ~i_8_447_1832_0 & ~i_8_447_1951_0))) | (~i_8_447_480_0 & ((~i_8_447_232_0 & i_8_447_674_0 & ~i_8_447_1060_0 & ~i_8_447_1808_0) | (~i_8_447_671_0 & ~i_8_447_1720_0 & i_8_447_2275_0 & ~i_8_447_2301_0))) | (~i_8_447_763_0 & ((i_8_447_492_0 & ~i_8_447_1185_0 & ~i_8_447_1722_0 & ~i_8_447_1737_0 & i_8_447_1821_0) | (~i_8_447_612_0 & ~i_8_447_684_0 & ~i_8_447_757_0 & ~i_8_447_1282_0 & i_8_447_2289_0))) | (~i_8_447_684_0 & ((i_8_447_360_0 & ~i_8_447_1587_0 & ~i_8_447_1719_0 & ~i_8_447_1720_0 & i_8_447_1821_0) | (i_8_447_612_0 & ~i_8_447_757_0 & i_8_447_1224_0 & ~i_8_447_1273_0 & ~i_8_447_1456_0 & ~i_8_447_1967_0 & ~i_8_447_1985_0))) | (i_8_447_1231_0 & ((~i_8_447_1720_0 & i_8_447_1807_0) | (i_8_447_592_0 & i_8_447_2149_0 & ~i_8_447_2301_0))) | (i_8_447_1808_0 & ((~i_8_447_757_0 & i_8_447_1951_0 & ~i_8_447_2300_0) | (~i_8_447_382_0 & i_8_447_670_0 & ~i_8_447_1807_0 & ~i_8_447_2303_0))) | (i_8_447_1818_0 & (i_8_447_2272_0 | (i_8_447_1282_0 & ~i_8_447_1737_0 & i_8_447_2290_0))) | (i_8_447_368_0 & ~i_8_447_704_0 & ~i_8_447_1129_0 & ~i_8_447_1185_0 & i_8_447_1456_0 & ~i_8_447_2303_0));
endmodule



// Benchmark "kernel_8_448" written by ABC on Sun Jul 19 10:10:57 2020

module kernel_8_448 ( 
    i_8_448_19_0, i_8_448_31_0, i_8_448_37_0, i_8_448_46_0, i_8_448_50_0,
    i_8_448_60_0, i_8_448_114_0, i_8_448_172_0, i_8_448_175_0,
    i_8_448_238_0, i_8_448_271_0, i_8_448_307_0, i_8_448_311_0,
    i_8_448_334_0, i_8_448_343_0, i_8_448_365_0, i_8_448_379_0,
    i_8_448_397_0, i_8_448_417_0, i_8_448_418_0, i_8_448_424_0,
    i_8_448_439_0, i_8_448_443_0, i_8_448_526_0, i_8_448_527_0,
    i_8_448_550_0, i_8_448_571_0, i_8_448_572_0, i_8_448_592_0,
    i_8_448_611_0, i_8_448_630_0, i_8_448_661_0, i_8_448_664_0,
    i_8_448_680_0, i_8_448_688_0, i_8_448_695_0, i_8_448_700_0,
    i_8_448_705_0, i_8_448_707_0, i_8_448_736_0, i_8_448_760_0,
    i_8_448_796_0, i_8_448_797_0, i_8_448_805_0, i_8_448_839_0,
    i_8_448_841_0, i_8_448_842_0, i_8_448_861_0, i_8_448_863_0,
    i_8_448_886_0, i_8_448_941_0, i_8_448_955_0, i_8_448_956_0,
    i_8_448_963_0, i_8_448_964_0, i_8_448_1018_0, i_8_448_1059_0,
    i_8_448_1066_0, i_8_448_1071_0, i_8_448_1090_0, i_8_448_1101_0,
    i_8_448_1179_0, i_8_448_1183_0, i_8_448_1226_0, i_8_448_1282_0,
    i_8_448_1291_0, i_8_448_1305_0, i_8_448_1336_0, i_8_448_1407_0,
    i_8_448_1408_0, i_8_448_1435_0, i_8_448_1542_0, i_8_448_1545_0,
    i_8_448_1561_0, i_8_448_1562_0, i_8_448_1587_0, i_8_448_1588_0,
    i_8_448_1610_0, i_8_448_1618_0, i_8_448_1634_0, i_8_448_1679_0,
    i_8_448_1697_0, i_8_448_1731_0, i_8_448_1733_0, i_8_448_1765_0,
    i_8_448_1818_0, i_8_448_1859_0, i_8_448_1888_0, i_8_448_1992_0,
    i_8_448_1996_0, i_8_448_2017_0, i_8_448_2056_0, i_8_448_2075_0,
    i_8_448_2145_0, i_8_448_2149_0, i_8_448_2152_0, i_8_448_2155_0,
    i_8_448_2156_0, i_8_448_2197_0, i_8_448_2209_0,
    o_8_448_0_0  );
  input  i_8_448_19_0, i_8_448_31_0, i_8_448_37_0, i_8_448_46_0,
    i_8_448_50_0, i_8_448_60_0, i_8_448_114_0, i_8_448_172_0,
    i_8_448_175_0, i_8_448_238_0, i_8_448_271_0, i_8_448_307_0,
    i_8_448_311_0, i_8_448_334_0, i_8_448_343_0, i_8_448_365_0,
    i_8_448_379_0, i_8_448_397_0, i_8_448_417_0, i_8_448_418_0,
    i_8_448_424_0, i_8_448_439_0, i_8_448_443_0, i_8_448_526_0,
    i_8_448_527_0, i_8_448_550_0, i_8_448_571_0, i_8_448_572_0,
    i_8_448_592_0, i_8_448_611_0, i_8_448_630_0, i_8_448_661_0,
    i_8_448_664_0, i_8_448_680_0, i_8_448_688_0, i_8_448_695_0,
    i_8_448_700_0, i_8_448_705_0, i_8_448_707_0, i_8_448_736_0,
    i_8_448_760_0, i_8_448_796_0, i_8_448_797_0, i_8_448_805_0,
    i_8_448_839_0, i_8_448_841_0, i_8_448_842_0, i_8_448_861_0,
    i_8_448_863_0, i_8_448_886_0, i_8_448_941_0, i_8_448_955_0,
    i_8_448_956_0, i_8_448_963_0, i_8_448_964_0, i_8_448_1018_0,
    i_8_448_1059_0, i_8_448_1066_0, i_8_448_1071_0, i_8_448_1090_0,
    i_8_448_1101_0, i_8_448_1179_0, i_8_448_1183_0, i_8_448_1226_0,
    i_8_448_1282_0, i_8_448_1291_0, i_8_448_1305_0, i_8_448_1336_0,
    i_8_448_1407_0, i_8_448_1408_0, i_8_448_1435_0, i_8_448_1542_0,
    i_8_448_1545_0, i_8_448_1561_0, i_8_448_1562_0, i_8_448_1587_0,
    i_8_448_1588_0, i_8_448_1610_0, i_8_448_1618_0, i_8_448_1634_0,
    i_8_448_1679_0, i_8_448_1697_0, i_8_448_1731_0, i_8_448_1733_0,
    i_8_448_1765_0, i_8_448_1818_0, i_8_448_1859_0, i_8_448_1888_0,
    i_8_448_1992_0, i_8_448_1996_0, i_8_448_2017_0, i_8_448_2056_0,
    i_8_448_2075_0, i_8_448_2145_0, i_8_448_2149_0, i_8_448_2152_0,
    i_8_448_2155_0, i_8_448_2156_0, i_8_448_2197_0, i_8_448_2209_0;
  output o_8_448_0_0;
  assign o_8_448_0_0 = 0;
endmodule



// Benchmark "kernel_8_449" written by ABC on Sun Jul 19 10:10:59 2020

module kernel_8_449 ( 
    i_8_449_28_0, i_8_449_38_0, i_8_449_107_0, i_8_449_142_0,
    i_8_449_171_0, i_8_449_213_0, i_8_449_214_0, i_8_449_272_0,
    i_8_449_292_0, i_8_449_295_0, i_8_449_298_0, i_8_449_300_0,
    i_8_449_301_0, i_8_449_302_0, i_8_449_307_0, i_8_449_308_0,
    i_8_449_310_0, i_8_449_314_0, i_8_449_338_0, i_8_449_351_0,
    i_8_449_420_0, i_8_449_421_0, i_8_449_430_0, i_8_449_483_0,
    i_8_449_489_0, i_8_449_492_0, i_8_449_496_0, i_8_449_498_0,
    i_8_449_528_0, i_8_449_589_0, i_8_449_591_0, i_8_449_592_0,
    i_8_449_605_0, i_8_449_606_0, i_8_449_631_0, i_8_449_633_0,
    i_8_449_635_0, i_8_449_677_0, i_8_449_679_0, i_8_449_689_0,
    i_8_449_706_0, i_8_449_709_0, i_8_449_766_0, i_8_449_780_0,
    i_8_449_830_0, i_8_449_849_0, i_8_449_925_0, i_8_449_954_0,
    i_8_449_985_0, i_8_449_1033_0, i_8_449_1138_0, i_8_449_1156_0,
    i_8_449_1263_0, i_8_449_1264_0, i_8_449_1267_0, i_8_449_1274_0,
    i_8_449_1283_0, i_8_449_1286_0, i_8_449_1332_0, i_8_449_1333_0,
    i_8_449_1335_0, i_8_449_1551_0, i_8_449_1558_0, i_8_449_1561_0,
    i_8_449_1595_0, i_8_449_1650_0, i_8_449_1651_0, i_8_449_1657_0,
    i_8_449_1658_0, i_8_449_1659_0, i_8_449_1671_0, i_8_449_1719_0,
    i_8_449_1740_0, i_8_449_1763_0, i_8_449_1779_0, i_8_449_1789_0,
    i_8_449_1801_0, i_8_449_1803_0, i_8_449_1805_0, i_8_449_1826_0,
    i_8_449_1861_0, i_8_449_1863_0, i_8_449_1989_0, i_8_449_1994_0,
    i_8_449_2004_0, i_8_449_2007_0, i_8_449_2010_0, i_8_449_2013_0,
    i_8_449_2150_0, i_8_449_2155_0, i_8_449_2164_0, i_8_449_2165_0,
    i_8_449_2253_0, i_8_449_2255_0, i_8_449_2256_0, i_8_449_2268_0,
    i_8_449_2272_0, i_8_449_2273_0, i_8_449_2275_0, i_8_449_2286_0,
    o_8_449_0_0  );
  input  i_8_449_28_0, i_8_449_38_0, i_8_449_107_0, i_8_449_142_0,
    i_8_449_171_0, i_8_449_213_0, i_8_449_214_0, i_8_449_272_0,
    i_8_449_292_0, i_8_449_295_0, i_8_449_298_0, i_8_449_300_0,
    i_8_449_301_0, i_8_449_302_0, i_8_449_307_0, i_8_449_308_0,
    i_8_449_310_0, i_8_449_314_0, i_8_449_338_0, i_8_449_351_0,
    i_8_449_420_0, i_8_449_421_0, i_8_449_430_0, i_8_449_483_0,
    i_8_449_489_0, i_8_449_492_0, i_8_449_496_0, i_8_449_498_0,
    i_8_449_528_0, i_8_449_589_0, i_8_449_591_0, i_8_449_592_0,
    i_8_449_605_0, i_8_449_606_0, i_8_449_631_0, i_8_449_633_0,
    i_8_449_635_0, i_8_449_677_0, i_8_449_679_0, i_8_449_689_0,
    i_8_449_706_0, i_8_449_709_0, i_8_449_766_0, i_8_449_780_0,
    i_8_449_830_0, i_8_449_849_0, i_8_449_925_0, i_8_449_954_0,
    i_8_449_985_0, i_8_449_1033_0, i_8_449_1138_0, i_8_449_1156_0,
    i_8_449_1263_0, i_8_449_1264_0, i_8_449_1267_0, i_8_449_1274_0,
    i_8_449_1283_0, i_8_449_1286_0, i_8_449_1332_0, i_8_449_1333_0,
    i_8_449_1335_0, i_8_449_1551_0, i_8_449_1558_0, i_8_449_1561_0,
    i_8_449_1595_0, i_8_449_1650_0, i_8_449_1651_0, i_8_449_1657_0,
    i_8_449_1658_0, i_8_449_1659_0, i_8_449_1671_0, i_8_449_1719_0,
    i_8_449_1740_0, i_8_449_1763_0, i_8_449_1779_0, i_8_449_1789_0,
    i_8_449_1801_0, i_8_449_1803_0, i_8_449_1805_0, i_8_449_1826_0,
    i_8_449_1861_0, i_8_449_1863_0, i_8_449_1989_0, i_8_449_1994_0,
    i_8_449_2004_0, i_8_449_2007_0, i_8_449_2010_0, i_8_449_2013_0,
    i_8_449_2150_0, i_8_449_2155_0, i_8_449_2164_0, i_8_449_2165_0,
    i_8_449_2253_0, i_8_449_2255_0, i_8_449_2256_0, i_8_449_2268_0,
    i_8_449_2272_0, i_8_449_2273_0, i_8_449_2275_0, i_8_449_2286_0;
  output o_8_449_0_0;
  assign o_8_449_0_0 = ~((~i_8_449_985_0 & ((i_8_449_300_0 & ((~i_8_449_213_0 & i_8_449_589_0 & ~i_8_449_954_0 & ~i_8_449_1805_0 & ~i_8_449_2007_0) | (~i_8_449_351_0 & ~i_8_449_766_0 & i_8_449_1156_0 & i_8_449_1267_0 & ~i_8_449_2010_0))) | (~i_8_449_351_0 & ((i_8_449_489_0 & i_8_449_606_0 & ~i_8_449_1803_0 & i_8_449_2268_0 & ~i_8_449_2272_0) | (~i_8_449_213_0 & ~i_8_449_308_0 & ~i_8_449_310_0 & ~i_8_449_314_0 & ~i_8_449_496_0 & ~i_8_449_780_0 & ~i_8_449_830_0 & ~i_8_449_954_0 & ~i_8_449_1650_0 & ~i_8_449_1651_0 & ~i_8_449_1763_0 & ~i_8_449_1801_0 & ~i_8_449_1863_0 & ~i_8_449_2004_0 & ~i_8_449_2007_0 & ~i_8_449_2013_0 & ~i_8_449_2253_0 & ~i_8_449_2273_0 & ~i_8_449_2275_0))) | (~i_8_449_492_0 & ((~i_8_449_308_0 & ~i_8_449_766_0 & ((~i_8_449_292_0 & i_8_449_298_0 & ~i_8_449_483_0 & ~i_8_449_1138_0 & ~i_8_449_1650_0 & ~i_8_449_1826_0 & ~i_8_449_2164_0 & ~i_8_449_2255_0 & ~i_8_449_2275_0) | (~i_8_449_38_0 & ~i_8_449_171_0 & ~i_8_449_213_0 & ~i_8_449_272_0 & ~i_8_449_310_0 & ~i_8_449_314_0 & ~i_8_449_498_0 & ~i_8_449_605_0 & ~i_8_449_1551_0 & ~i_8_449_1561_0 & ~i_8_449_1595_0 & ~i_8_449_1658_0 & ~i_8_449_1659_0 & ~i_8_449_1863_0 & ~i_8_449_2004_0 & ~i_8_449_2007_0 & ~i_8_449_2013_0 & ~i_8_449_2253_0 & ~i_8_449_2273_0 & ~i_8_449_2286_0))) | (~i_8_449_496_0 & ~i_8_449_780_0 & i_8_449_302_0 & ~i_8_449_314_0 & ~i_8_449_1138_0 & ~i_8_449_2253_0 & ~i_8_449_2255_0 & ~i_8_449_2268_0))) | (~i_8_449_2013_0 & ((~i_8_449_213_0 & ~i_8_449_421_0 & ~i_8_449_1658_0 & ~i_8_449_2256_0 & ~i_8_449_2286_0 & ((~i_8_449_308_0 & i_8_449_592_0 & ~i_8_449_633_0 & ~i_8_449_2268_0 & i_8_449_2275_0) | (~i_8_449_310_0 & ~i_8_449_338_0 & ~i_8_449_591_0 & ~i_8_449_631_0 & ~i_8_449_679_0 & ~i_8_449_709_0 & ~i_8_449_1551_0 & ~i_8_449_1657_0 & ~i_8_449_1671_0 & ~i_8_449_1805_0 & ~i_8_449_1826_0 & ~i_8_449_1861_0 & ~i_8_449_2255_0 & ~i_8_449_2275_0 & ~i_8_449_2010_0 & ~i_8_449_2253_0))) | (i_8_449_295_0 & ~i_8_449_307_0 & ~i_8_449_310_0 & ~i_8_449_1659_0 & ~i_8_449_1671_0))))) | (~i_8_449_2165_0 & ((~i_8_449_213_0 & ((~i_8_449_308_0 & ~i_8_449_351_0 & i_8_449_528_0 & ~i_8_449_633_0 & ~i_8_449_1156_0 & ~i_8_449_1658_0 & ~i_8_449_1826_0 & ~i_8_449_1863_0 & ~i_8_449_2010_0 & ~i_8_449_2013_0 & ~i_8_449_2253_0) | (i_8_449_301_0 & ~i_8_449_307_0 & ~i_8_449_605_0 & ~i_8_449_631_0 & ~i_8_449_709_0 & ~i_8_449_849_0 & ~i_8_449_1138_0 & ~i_8_449_1671_0 & ~i_8_449_2268_0 & ~i_8_449_2273_0))) | (~i_8_449_214_0 & ~i_8_449_272_0 & ((~i_8_449_307_0 & ~i_8_449_589_0 & ~i_8_449_766_0 & ~i_8_449_1138_0 & ~i_8_449_1551_0 & ~i_8_449_1763_0 & i_8_449_1994_0 & ~i_8_449_2255_0 & ~i_8_449_2268_0 & ~i_8_449_2272_0 & ~i_8_449_2275_0) | (~i_8_449_528_0 & ~i_8_449_633_0 & i_8_449_1283_0 & ~i_8_449_1558_0 & ~i_8_449_1657_0 & ~i_8_449_1658_0 & ~i_8_449_1805_0 & ~i_8_449_2273_0 & ~i_8_449_2286_0))) | (~i_8_449_314_0 & ~i_8_449_496_0 & ((i_8_449_301_0 & ~i_8_449_498_0 & ~i_8_449_1651_0 & ~i_8_449_1658_0 & ~i_8_449_1659_0 & ~i_8_449_1671_0 & ~i_8_449_2004_0 & ~i_8_449_2007_0 & ~i_8_449_2253_0) | (~i_8_449_307_0 & i_8_449_635_0 & ~i_8_449_679_0 & ~i_8_449_1263_0 & ~i_8_449_1335_0 & ~i_8_449_1803_0 & ~i_8_449_1989_0 & ~i_8_449_2272_0))) | (~i_8_449_1805_0 & ((i_8_449_1763_0 & ~i_8_449_2273_0 & ~i_8_449_2275_0) | (~i_8_449_38_0 & i_8_449_338_0 & ~i_8_449_706_0 & ~i_8_449_954_0 & ~i_8_449_1138_0 & ~i_8_449_1651_0 & ~i_8_449_1803_0 & ~i_8_449_2286_0))))) | (~i_8_449_498_0 & ((~i_8_449_214_0 & ~i_8_449_351_0 & ((~i_8_449_28_0 & ~i_8_449_171_0 & ~i_8_449_272_0 & ~i_8_449_307_0 & ~i_8_449_310_0 & ~i_8_449_420_0 & ~i_8_449_830_0 & ~i_8_449_1033_0 & i_8_449_1264_0 & ~i_8_449_1657_0 & ~i_8_449_1658_0 & ~i_8_449_1805_0 & ~i_8_449_2007_0 & ~i_8_449_2164_0) | (~i_8_449_308_0 & ~i_8_449_314_0 & ~i_8_449_489_0 & ~i_8_449_677_0 & ~i_8_449_706_0 & ~i_8_449_1719_0 & ~i_8_449_1994_0 & ~i_8_449_2004_0 & ~i_8_449_2010_0 & i_8_449_2155_0 & ~i_8_449_2253_0))) | (~i_8_449_307_0 & ((~i_8_449_338_0 & ~i_8_449_709_0 & i_8_449_1263_0 & ~i_8_449_1558_0 & ~i_8_449_1595_0 & ~i_8_449_1651_0 & ~i_8_449_1740_0 & ~i_8_449_1803_0 & ~i_8_449_2155_0 & ~i_8_449_2273_0) | (~i_8_449_213_0 & ~i_8_449_925_0 & i_8_449_1740_0 & ~i_8_449_1801_0 & ~i_8_449_2013_0 & ~i_8_449_2275_0))) | (~i_8_449_338_0 & ~i_8_449_421_0 & ~i_8_449_430_0 & ~i_8_449_489_0 & ~i_8_449_954_0 & ~i_8_449_1033_0 & ~i_8_449_1551_0 & ~i_8_449_1657_0 & ~i_8_449_1801_0 & ~i_8_449_1803_0 & ~i_8_449_1826_0 & ~i_8_449_1994_0 & ~i_8_449_2150_0 & ~i_8_449_2155_0))) | (~i_8_449_2164_0 & ((~i_8_449_28_0 & ((~i_8_449_107_0 & ~i_8_449_295_0 & ~i_8_449_633_0 & ~i_8_449_679_0 & ~i_8_449_706_0 & ~i_8_449_709_0 & i_8_449_1789_0 & ~i_8_449_2155_0 & ~i_8_449_2255_0 & ~i_8_449_2268_0 & ~i_8_449_2272_0) | (~i_8_449_171_0 & ~i_8_449_300_0 & ~i_8_449_351_0 & ~i_8_449_925_0 & i_8_449_1333_0 & ~i_8_449_1561_0 & ~i_8_449_1658_0 & ~i_8_449_1659_0 & ~i_8_449_1805_0 & ~i_8_449_2275_0))) | (~i_8_449_308_0 & ~i_8_449_1595_0 & ~i_8_449_2256_0 & ((~i_8_449_38_0 & i_8_449_302_0 & ~i_8_449_421_0 & ~i_8_449_496_0 & ~i_8_449_925_0 & ~i_8_449_1651_0 & ~i_8_449_1657_0 & ~i_8_449_1789_0 & ~i_8_449_2013_0) | (~i_8_449_213_0 & ~i_8_449_307_0 & ~i_8_449_314_0 & ~i_8_449_351_0 & ~i_8_449_430_0 & ~i_8_449_492_0 & ~i_8_449_954_0 & i_8_449_1551_0 & ~i_8_449_1658_0 & ~i_8_449_1861_0 & ~i_8_449_2010_0 & ~i_8_449_2268_0 & ~i_8_449_2273_0 & ~i_8_449_2275_0 & ~i_8_449_2286_0))) | (~i_8_449_310_0 & ~i_8_449_528_0 & i_8_449_633_0 & ~i_8_449_1671_0 & i_8_449_1779_0 & ~i_8_449_2268_0))) | (~i_8_449_214_0 & ((~i_8_449_38_0 & ((~i_8_449_709_0 & ~i_8_449_766_0 & ~i_8_449_830_0 & i_8_449_1286_0 & i_8_449_1789_0 & ~i_8_449_1861_0 & ~i_8_449_2004_0 & ~i_8_449_2010_0) | (~i_8_449_213_0 & ~i_8_449_925_0 & ~i_8_449_1033_0 & ~i_8_449_2272_0 & ~i_8_449_2275_0 & i_8_449_1335_0 & ~i_8_449_1863_0))) | (~i_8_449_308_0 & ~i_8_449_421_0 & ~i_8_449_528_0 & i_8_449_591_0 & ~i_8_449_605_0 & ~i_8_449_689_0 & ~i_8_449_925_0 & ~i_8_449_1561_0 & ~i_8_449_1657_0 & ~i_8_449_1659_0 & ~i_8_449_2013_0 & ~i_8_449_2253_0 & ~i_8_449_2256_0 & ~i_8_449_2268_0))) | (~i_8_449_308_0 & ((~i_8_449_272_0 & ((~i_8_449_314_0 & ~i_8_449_496_0 & ~i_8_449_605_0 & ~i_8_449_1138_0 & ~i_8_449_2272_0 & ~i_8_449_2275_0 & i_8_449_1286_0 & ~i_8_449_1863_0) | (~i_8_449_171_0 & ~i_8_449_310_0 & i_8_449_1558_0 & ~i_8_449_1657_0 & ~i_8_449_1803_0 & i_8_449_1989_0 & ~i_8_449_2286_0))) | (~i_8_449_307_0 & i_8_449_1274_0 & ~i_8_449_1595_0 & ~i_8_449_1651_0 & ~i_8_449_1658_0 & ~i_8_449_1805_0))) | (~i_8_449_307_0 & ((~i_8_449_314_0 & ~i_8_449_2268_0 & ((~i_8_449_351_0 & ~i_8_449_492_0 & ~i_8_449_496_0 & ~i_8_449_709_0 & ~i_8_449_766_0 & ~i_8_449_830_0 & ~i_8_449_954_0 & ~i_8_449_1283_0 & ~i_8_449_1650_0 & ~i_8_449_1803_0 & ~i_8_449_1805_0 & ~i_8_449_1861_0 & ~i_8_449_2255_0) | (~i_8_449_2004_0 & ~i_8_449_2010_0 & i_8_449_1779_0 & i_8_449_1789_0 & ~i_8_449_2273_0 & ~i_8_449_2286_0 & ~i_8_449_2155_0 & ~i_8_449_2253_0))) | (~i_8_449_1826_0 & ~i_8_449_1863_0 & ~i_8_449_1994_0 & ((~i_8_449_489_0 & i_8_449_606_0 & ~i_8_449_766_0 & ~i_8_449_780_0 & ~i_8_449_954_0 & ~i_8_449_1595_0 & ~i_8_449_1659_0 & ~i_8_449_2010_0) | (~i_8_449_1156_0 & ~i_8_449_1264_0 & i_8_449_1283_0 & ~i_8_449_1551_0 & ~i_8_449_1789_0 & ~i_8_449_2275_0))))) | (~i_8_449_213_0 & ~i_8_449_310_0 & i_8_449_780_0 & ~i_8_449_1033_0 & ~i_8_449_1558_0 & ~i_8_449_1671_0 & ~i_8_449_1861_0 & ~i_8_449_2004_0 & ~i_8_449_2007_0 & ~i_8_449_2255_0 & ~i_8_449_2256_0 & ~i_8_449_2273_0) | (i_8_449_605_0 & i_8_449_677_0 & ~i_8_449_1595_0 & ~i_8_449_2272_0));
endmodule



// Benchmark "kernel_8_450" written by ABC on Sun Jul 19 10:11:00 2020

module kernel_8_450 ( 
    i_8_450_35_0, i_8_450_43_0, i_8_450_88_0, i_8_450_114_0, i_8_450_115_0,
    i_8_450_124_0, i_8_450_130_0, i_8_450_148_0, i_8_450_193_0,
    i_8_450_194_0, i_8_450_338_0, i_8_450_363_0, i_8_450_371_0,
    i_8_450_377_0, i_8_450_421_0, i_8_450_455_0, i_8_450_494_0,
    i_8_450_509_0, i_8_450_534_0, i_8_450_553_0, i_8_450_556_0,
    i_8_450_616_0, i_8_450_637_0, i_8_450_653_0, i_8_450_656_0,
    i_8_450_694_0, i_8_450_697_0, i_8_450_833_0, i_8_450_959_0,
    i_8_450_992_0, i_8_450_1027_0, i_8_450_1037_0, i_8_450_1110_0,
    i_8_450_1111_0, i_8_450_1127_0, i_8_450_1130_0, i_8_450_1132_0,
    i_8_450_1202_0, i_8_450_1204_0, i_8_450_1224_0, i_8_450_1226_0,
    i_8_450_1306_0, i_8_450_1307_0, i_8_450_1310_0, i_8_450_1312_0,
    i_8_450_1399_0, i_8_450_1400_0, i_8_450_1444_0, i_8_450_1455_0,
    i_8_450_1462_0, i_8_450_1471_0, i_8_450_1472_0, i_8_450_1486_0,
    i_8_450_1490_0, i_8_450_1524_0, i_8_450_1547_0, i_8_450_1549_0,
    i_8_450_1550_0, i_8_450_1552_0, i_8_450_1562_0, i_8_450_1634_0,
    i_8_450_1641_0, i_8_450_1660_0, i_8_450_1669_0, i_8_450_1748_0,
    i_8_450_1750_0, i_8_450_1771_0, i_8_450_1795_0, i_8_450_1805_0,
    i_8_450_1810_0, i_8_450_1823_0, i_8_450_1824_0, i_8_450_1825_0,
    i_8_450_1881_0, i_8_450_1886_0, i_8_450_1895_0, i_8_450_1939_0,
    i_8_450_1951_0, i_8_450_1973_0, i_8_450_1976_0, i_8_450_2009_0,
    i_8_450_2011_0, i_8_450_2012_0, i_8_450_2045_0, i_8_450_2090_0,
    i_8_450_2098_0, i_8_450_2101_0, i_8_450_2122_0, i_8_450_2137_0,
    i_8_450_2143_0, i_8_450_2146_0, i_8_450_2150_0, i_8_450_2167_0,
    i_8_450_2170_0, i_8_450_2171_0, i_8_450_2194_0, i_8_450_2201_0,
    i_8_450_2236_0, i_8_450_2242_0, i_8_450_2245_0,
    o_8_450_0_0  );
  input  i_8_450_35_0, i_8_450_43_0, i_8_450_88_0, i_8_450_114_0,
    i_8_450_115_0, i_8_450_124_0, i_8_450_130_0, i_8_450_148_0,
    i_8_450_193_0, i_8_450_194_0, i_8_450_338_0, i_8_450_363_0,
    i_8_450_371_0, i_8_450_377_0, i_8_450_421_0, i_8_450_455_0,
    i_8_450_494_0, i_8_450_509_0, i_8_450_534_0, i_8_450_553_0,
    i_8_450_556_0, i_8_450_616_0, i_8_450_637_0, i_8_450_653_0,
    i_8_450_656_0, i_8_450_694_0, i_8_450_697_0, i_8_450_833_0,
    i_8_450_959_0, i_8_450_992_0, i_8_450_1027_0, i_8_450_1037_0,
    i_8_450_1110_0, i_8_450_1111_0, i_8_450_1127_0, i_8_450_1130_0,
    i_8_450_1132_0, i_8_450_1202_0, i_8_450_1204_0, i_8_450_1224_0,
    i_8_450_1226_0, i_8_450_1306_0, i_8_450_1307_0, i_8_450_1310_0,
    i_8_450_1312_0, i_8_450_1399_0, i_8_450_1400_0, i_8_450_1444_0,
    i_8_450_1455_0, i_8_450_1462_0, i_8_450_1471_0, i_8_450_1472_0,
    i_8_450_1486_0, i_8_450_1490_0, i_8_450_1524_0, i_8_450_1547_0,
    i_8_450_1549_0, i_8_450_1550_0, i_8_450_1552_0, i_8_450_1562_0,
    i_8_450_1634_0, i_8_450_1641_0, i_8_450_1660_0, i_8_450_1669_0,
    i_8_450_1748_0, i_8_450_1750_0, i_8_450_1771_0, i_8_450_1795_0,
    i_8_450_1805_0, i_8_450_1810_0, i_8_450_1823_0, i_8_450_1824_0,
    i_8_450_1825_0, i_8_450_1881_0, i_8_450_1886_0, i_8_450_1895_0,
    i_8_450_1939_0, i_8_450_1951_0, i_8_450_1973_0, i_8_450_1976_0,
    i_8_450_2009_0, i_8_450_2011_0, i_8_450_2012_0, i_8_450_2045_0,
    i_8_450_2090_0, i_8_450_2098_0, i_8_450_2101_0, i_8_450_2122_0,
    i_8_450_2137_0, i_8_450_2143_0, i_8_450_2146_0, i_8_450_2150_0,
    i_8_450_2167_0, i_8_450_2170_0, i_8_450_2171_0, i_8_450_2194_0,
    i_8_450_2201_0, i_8_450_2236_0, i_8_450_2242_0, i_8_450_2245_0;
  output o_8_450_0_0;
  assign o_8_450_0_0 = 0;
endmodule



// Benchmark "kernel_8_451" written by ABC on Sun Jul 19 10:11:01 2020

module kernel_8_451 ( 
    i_8_451_18_0, i_8_451_27_0, i_8_451_40_0, i_8_451_46_0, i_8_451_90_0,
    i_8_451_166_0, i_8_451_171_0, i_8_451_173_0, i_8_451_191_0,
    i_8_451_207_0, i_8_451_227_0, i_8_451_288_0, i_8_451_343_0,
    i_8_451_361_0, i_8_451_378_0, i_8_451_396_0, i_8_451_397_0,
    i_8_451_415_0, i_8_451_423_0, i_8_451_490_0, i_8_451_498_0,
    i_8_451_522_0, i_8_451_523_0, i_8_451_594_0, i_8_451_608_0,
    i_8_451_612_0, i_8_451_615_0, i_8_451_648_0, i_8_451_684_0,
    i_8_451_690_0, i_8_451_694_0, i_8_451_703_0, i_8_451_766_0,
    i_8_451_795_0, i_8_451_810_0, i_8_451_827_0, i_8_451_829_0,
    i_8_451_838_0, i_8_451_858_0, i_8_451_883_0, i_8_451_927_0,
    i_8_451_954_0, i_8_451_963_0, i_8_451_965_0, i_8_451_993_0,
    i_8_451_1017_0, i_8_451_1053_0, i_8_451_1054_0, i_8_451_1107_0,
    i_8_451_1143_0, i_8_451_1171_0, i_8_451_1224_0, i_8_451_1225_0,
    i_8_451_1261_0, i_8_451_1269_0, i_8_451_1278_0, i_8_451_1279_0,
    i_8_451_1287_0, i_8_451_1288_0, i_8_451_1297_0, i_8_451_1377_0,
    i_8_451_1380_0, i_8_451_1435_0, i_8_451_1467_0, i_8_451_1489_0,
    i_8_451_1548_0, i_8_451_1603_0, i_8_451_1629_0, i_8_451_1638_0,
    i_8_451_1641_0, i_8_451_1693_0, i_8_451_1720_0, i_8_451_1722_0,
    i_8_451_1729_0, i_8_451_1737_0, i_8_451_1740_0, i_8_451_1741_0,
    i_8_451_1869_0, i_8_451_1884_0, i_8_451_1936_0, i_8_451_1993_0,
    i_8_451_1994_0, i_8_451_1998_0, i_8_451_2034_0, i_8_451_2052_0,
    i_8_451_2053_0, i_8_451_2055_0, i_8_451_2089_0, i_8_451_2101_0,
    i_8_451_2102_0, i_8_451_2106_0, i_8_451_2140_0, i_8_451_2169_0,
    i_8_451_2172_0, i_8_451_2178_0, i_8_451_2196_0, i_8_451_2223_0,
    i_8_451_2225_0, i_8_451_2226_0, i_8_451_2296_0,
    o_8_451_0_0  );
  input  i_8_451_18_0, i_8_451_27_0, i_8_451_40_0, i_8_451_46_0,
    i_8_451_90_0, i_8_451_166_0, i_8_451_171_0, i_8_451_173_0,
    i_8_451_191_0, i_8_451_207_0, i_8_451_227_0, i_8_451_288_0,
    i_8_451_343_0, i_8_451_361_0, i_8_451_378_0, i_8_451_396_0,
    i_8_451_397_0, i_8_451_415_0, i_8_451_423_0, i_8_451_490_0,
    i_8_451_498_0, i_8_451_522_0, i_8_451_523_0, i_8_451_594_0,
    i_8_451_608_0, i_8_451_612_0, i_8_451_615_0, i_8_451_648_0,
    i_8_451_684_0, i_8_451_690_0, i_8_451_694_0, i_8_451_703_0,
    i_8_451_766_0, i_8_451_795_0, i_8_451_810_0, i_8_451_827_0,
    i_8_451_829_0, i_8_451_838_0, i_8_451_858_0, i_8_451_883_0,
    i_8_451_927_0, i_8_451_954_0, i_8_451_963_0, i_8_451_965_0,
    i_8_451_993_0, i_8_451_1017_0, i_8_451_1053_0, i_8_451_1054_0,
    i_8_451_1107_0, i_8_451_1143_0, i_8_451_1171_0, i_8_451_1224_0,
    i_8_451_1225_0, i_8_451_1261_0, i_8_451_1269_0, i_8_451_1278_0,
    i_8_451_1279_0, i_8_451_1287_0, i_8_451_1288_0, i_8_451_1297_0,
    i_8_451_1377_0, i_8_451_1380_0, i_8_451_1435_0, i_8_451_1467_0,
    i_8_451_1489_0, i_8_451_1548_0, i_8_451_1603_0, i_8_451_1629_0,
    i_8_451_1638_0, i_8_451_1641_0, i_8_451_1693_0, i_8_451_1720_0,
    i_8_451_1722_0, i_8_451_1729_0, i_8_451_1737_0, i_8_451_1740_0,
    i_8_451_1741_0, i_8_451_1869_0, i_8_451_1884_0, i_8_451_1936_0,
    i_8_451_1993_0, i_8_451_1994_0, i_8_451_1998_0, i_8_451_2034_0,
    i_8_451_2052_0, i_8_451_2053_0, i_8_451_2055_0, i_8_451_2089_0,
    i_8_451_2101_0, i_8_451_2102_0, i_8_451_2106_0, i_8_451_2140_0,
    i_8_451_2169_0, i_8_451_2172_0, i_8_451_2178_0, i_8_451_2196_0,
    i_8_451_2223_0, i_8_451_2225_0, i_8_451_2226_0, i_8_451_2296_0;
  output o_8_451_0_0;
  assign o_8_451_0_0 = 0;
endmodule



// Benchmark "kernel_8_452" written by ABC on Sun Jul 19 10:11:02 2020

module kernel_8_452 ( 
    i_8_452_44_0, i_8_452_45_0, i_8_452_60_0, i_8_452_69_0, i_8_452_70_0,
    i_8_452_90_0, i_8_452_106_0, i_8_452_166_0, i_8_452_194_0,
    i_8_452_224_0, i_8_452_225_0, i_8_452_226_0, i_8_452_227_0,
    i_8_452_241_0, i_8_452_301_0, i_8_452_340_0, i_8_452_341_0,
    i_8_452_348_0, i_8_452_362_0, i_8_452_402_0, i_8_452_528_0,
    i_8_452_529_0, i_8_452_601_0, i_8_452_602_0, i_8_452_628_0,
    i_8_452_630_0, i_8_452_631_0, i_8_452_632_0, i_8_452_651_0,
    i_8_452_652_0, i_8_452_653_0, i_8_452_654_0, i_8_452_660_0,
    i_8_452_665_0, i_8_452_672_0, i_8_452_691_0, i_8_452_717_0,
    i_8_452_719_0, i_8_452_765_0, i_8_452_768_0, i_8_452_795_0,
    i_8_452_836_0, i_8_452_839_0, i_8_452_844_0, i_8_452_853_0,
    i_8_452_857_0, i_8_452_877_0, i_8_452_880_0, i_8_452_881_0,
    i_8_452_1033_0, i_8_452_1042_0, i_8_452_1105_0, i_8_452_1132_0,
    i_8_452_1155_0, i_8_452_1156_0, i_8_452_1295_0, i_8_452_1314_0,
    i_8_452_1321_0, i_8_452_1322_0, i_8_452_1329_0, i_8_452_1330_0,
    i_8_452_1331_0, i_8_452_1338_0, i_8_452_1339_0, i_8_452_1356_0,
    i_8_452_1383_0, i_8_452_1384_0, i_8_452_1389_0, i_8_452_1407_0,
    i_8_452_1410_0, i_8_452_1435_0, i_8_452_1625_0, i_8_452_1673_0,
    i_8_452_1705_0, i_8_452_1708_0, i_8_452_1776_0, i_8_452_1818_0,
    i_8_452_1819_0, i_8_452_1821_0, i_8_452_1830_0, i_8_452_1834_0,
    i_8_452_1835_0, i_8_452_1844_0, i_8_452_1862_0, i_8_452_1942_0,
    i_8_452_1987_0, i_8_452_1995_0, i_8_452_1996_0, i_8_452_2016_0,
    i_8_452_2022_0, i_8_452_2095_0, i_8_452_2096_0, i_8_452_2109_0,
    i_8_452_2112_0, i_8_452_2113_0, i_8_452_2151_0, i_8_452_2171_0,
    i_8_452_2178_0, i_8_452_2227_0, i_8_452_2244_0,
    o_8_452_0_0  );
  input  i_8_452_44_0, i_8_452_45_0, i_8_452_60_0, i_8_452_69_0,
    i_8_452_70_0, i_8_452_90_0, i_8_452_106_0, i_8_452_166_0,
    i_8_452_194_0, i_8_452_224_0, i_8_452_225_0, i_8_452_226_0,
    i_8_452_227_0, i_8_452_241_0, i_8_452_301_0, i_8_452_340_0,
    i_8_452_341_0, i_8_452_348_0, i_8_452_362_0, i_8_452_402_0,
    i_8_452_528_0, i_8_452_529_0, i_8_452_601_0, i_8_452_602_0,
    i_8_452_628_0, i_8_452_630_0, i_8_452_631_0, i_8_452_632_0,
    i_8_452_651_0, i_8_452_652_0, i_8_452_653_0, i_8_452_654_0,
    i_8_452_660_0, i_8_452_665_0, i_8_452_672_0, i_8_452_691_0,
    i_8_452_717_0, i_8_452_719_0, i_8_452_765_0, i_8_452_768_0,
    i_8_452_795_0, i_8_452_836_0, i_8_452_839_0, i_8_452_844_0,
    i_8_452_853_0, i_8_452_857_0, i_8_452_877_0, i_8_452_880_0,
    i_8_452_881_0, i_8_452_1033_0, i_8_452_1042_0, i_8_452_1105_0,
    i_8_452_1132_0, i_8_452_1155_0, i_8_452_1156_0, i_8_452_1295_0,
    i_8_452_1314_0, i_8_452_1321_0, i_8_452_1322_0, i_8_452_1329_0,
    i_8_452_1330_0, i_8_452_1331_0, i_8_452_1338_0, i_8_452_1339_0,
    i_8_452_1356_0, i_8_452_1383_0, i_8_452_1384_0, i_8_452_1389_0,
    i_8_452_1407_0, i_8_452_1410_0, i_8_452_1435_0, i_8_452_1625_0,
    i_8_452_1673_0, i_8_452_1705_0, i_8_452_1708_0, i_8_452_1776_0,
    i_8_452_1818_0, i_8_452_1819_0, i_8_452_1821_0, i_8_452_1830_0,
    i_8_452_1834_0, i_8_452_1835_0, i_8_452_1844_0, i_8_452_1862_0,
    i_8_452_1942_0, i_8_452_1987_0, i_8_452_1995_0, i_8_452_1996_0,
    i_8_452_2016_0, i_8_452_2022_0, i_8_452_2095_0, i_8_452_2096_0,
    i_8_452_2109_0, i_8_452_2112_0, i_8_452_2113_0, i_8_452_2151_0,
    i_8_452_2171_0, i_8_452_2178_0, i_8_452_2227_0, i_8_452_2244_0;
  output o_8_452_0_0;
  assign o_8_452_0_0 = ~((~i_8_452_348_0 & ((i_8_452_225_0 & ~i_8_452_795_0 & i_8_452_1776_0 & ~i_8_452_1818_0) | (~i_8_452_45_0 & ~i_8_452_194_0 & ~i_8_452_765_0 & ~i_8_452_768_0 & i_8_452_877_0 & ~i_8_452_1156_0 & ~i_8_452_1322_0 & ~i_8_452_1410_0 & ~i_8_452_1435_0 & ~i_8_452_1705_0 & ~i_8_452_1821_0 & ~i_8_452_1987_0 & ~i_8_452_2151_0))) | (~i_8_452_1830_0 & ((~i_8_452_1987_0 & ((~i_8_452_44_0 & ~i_8_452_1155_0 & ~i_8_452_2178_0 & ((~i_8_452_529_0 & ~i_8_452_665_0 & ~i_8_452_765_0 & ~i_8_452_768_0 & ~i_8_452_877_0 & ~i_8_452_1156_0 & ~i_8_452_1295_0 & ~i_8_452_1321_0 & ~i_8_452_1329_0 & ~i_8_452_1330_0 & ~i_8_452_1383_0 & ~i_8_452_1407_0 & ~i_8_452_1625_0 & ~i_8_452_1705_0 & ~i_8_452_1818_0 & ~i_8_452_1942_0 & ~i_8_452_2016_0 & ~i_8_452_2113_0) | (~i_8_452_69_0 & ~i_8_452_691_0 & i_8_452_844_0 & ~i_8_452_1339_0 & ~i_8_452_1708_0 & ~i_8_452_1821_0 & ~i_8_452_1835_0 & ~i_8_452_1844_0 & ~i_8_452_1995_0 & ~i_8_452_2022_0 & ~i_8_452_2151_0 & ~i_8_452_2244_0))) | (~i_8_452_69_0 & i_8_452_630_0 & ~i_8_452_795_0 & ~i_8_452_1033_0 & ~i_8_452_1156_0 & ~i_8_452_1322_0))) | (~i_8_452_2227_0 & ((~i_8_452_765_0 & ((~i_8_452_44_0 & ~i_8_452_1295_0 & ~i_8_452_1708_0 & ((~i_8_452_45_0 & ~i_8_452_631_0 & ~i_8_452_717_0 & ~i_8_452_768_0 & i_8_452_880_0 & ~i_8_452_1339_0 & ~i_8_452_1942_0 & ~i_8_452_2022_0 & ~i_8_452_2113_0) | (i_8_452_301_0 & ~i_8_452_795_0 & ~i_8_452_1156_0 & ~i_8_452_1407_0 & ~i_8_452_1410_0 & ~i_8_452_1705_0 & ~i_8_452_1776_0 & ~i_8_452_1835_0 & ~i_8_452_2016_0 & ~i_8_452_2109_0 & ~i_8_452_2112_0 & ~i_8_452_2151_0))) | (~i_8_452_528_0 & ~i_8_452_665_0 & ~i_8_452_691_0 & i_8_452_844_0 & ~i_8_452_853_0 & ~i_8_452_880_0 & ~i_8_452_1322_0 & ~i_8_452_1821_0 & ~i_8_452_1834_0 & ~i_8_452_1996_0 & ~i_8_452_2112_0))) | (i_8_452_225_0 & ((~i_8_452_45_0 & ~i_8_452_853_0 & ~i_8_452_1322_0 & ~i_8_452_1339_0 & ~i_8_452_1942_0) | (~i_8_452_1155_0 & ~i_8_452_2109_0 & ~i_8_452_2178_0))))) | (i_8_452_628_0 & ((~i_8_452_90_0 & i_8_452_106_0 & ~i_8_452_402_0 & ~i_8_452_672_0 & ~i_8_452_1295_0 & ~i_8_452_1818_0) | (~i_8_452_765_0 & i_8_452_880_0 & ~i_8_452_1339_0 & ~i_8_452_1435_0 & ~i_8_452_2016_0 & ~i_8_452_2022_0 & ~i_8_452_2109_0))) | (~i_8_452_90_0 & ((~i_8_452_402_0 & i_8_452_631_0 & ~i_8_452_765_0 & ~i_8_452_1835_0 & ~i_8_452_1844_0) | (~i_8_452_660_0 & ~i_8_452_1321_0 & ~i_8_452_1330_0 & ~i_8_452_1384_0 & i_8_452_1819_0 & ~i_8_452_1834_0 & ~i_8_452_1996_0 & ~i_8_452_2016_0 & ~i_8_452_2178_0))) | (~i_8_452_1835_0 & ((~i_8_452_402_0 & ((~i_8_452_765_0 & ~i_8_452_768_0 & ~i_8_452_836_0 & i_8_452_839_0 & ~i_8_452_881_0 & ~i_8_452_1156_0 & ~i_8_452_1339_0 & ~i_8_452_1834_0 & ~i_8_452_1844_0 & ~i_8_452_1942_0 & ~i_8_452_2016_0) | (~i_8_452_224_0 & i_8_452_529_0 & ~i_8_452_691_0 & ~i_8_452_844_0 & ~i_8_452_1331_0 & ~i_8_452_1705_0 & ~i_8_452_2022_0 & ~i_8_452_2151_0))) | (~i_8_452_341_0 & ((~i_8_452_1156_0 & ~i_8_452_1383_0 & ((~i_8_452_166_0 & ~i_8_452_194_0 & ~i_8_452_630_0 & i_8_452_881_0 & ~i_8_452_1322_0 & ~i_8_452_1338_0 & ~i_8_452_1384_0) | (~i_8_452_45_0 & ~i_8_452_340_0 & ~i_8_452_665_0 & ~i_8_452_765_0 & ~i_8_452_768_0 & ~i_8_452_1329_0 & ~i_8_452_1330_0 & ~i_8_452_1410_0 & ~i_8_452_1435_0 & ~i_8_452_1625_0 & ~i_8_452_1708_0 & ~i_8_452_1844_0 & ~i_8_452_2178_0))) | (~i_8_452_44_0 & i_8_452_665_0 & i_8_452_1322_0 & ~i_8_452_1996_0 & ~i_8_452_2022_0))))) | (~i_8_452_839_0 & i_8_452_857_0 & ~i_8_452_1155_0 & ~i_8_452_1156_0 & ~i_8_452_1295_0 & ~i_8_452_1384_0 & ~i_8_452_1942_0))) | (~i_8_452_1155_0 & ((~i_8_452_69_0 & ~i_8_452_1384_0 & ((~i_8_452_340_0 & ~i_8_452_341_0 & ~i_8_452_628_0 & ~i_8_452_1105_0 & i_8_452_1410_0 & ~i_8_452_1818_0 & ~i_8_452_1834_0 & ~i_8_452_2112_0) | (i_8_452_226_0 & ~i_8_452_1295_0 & ~i_8_452_1330_0 & ~i_8_452_2178_0))) | (~i_8_452_70_0 & ((~i_8_452_241_0 & ~i_8_452_301_0 & ~i_8_452_844_0 & ~i_8_452_877_0 & ~i_8_452_1156_0 & ~i_8_452_1322_0 & ~i_8_452_1834_0 & i_8_452_1995_0) | (~i_8_452_90_0 & ~i_8_452_341_0 & ~i_8_452_628_0 & ~i_8_452_654_0 & ~i_8_452_672_0 & ~i_8_452_768_0 & ~i_8_452_1314_0 & ~i_8_452_1330_0 & i_8_452_1821_0 & ~i_8_452_1942_0 & ~i_8_452_2016_0 & ~i_8_452_2244_0))) | (~i_8_452_765_0 & ((~i_8_452_631_0 & ((~i_8_452_44_0 & ~i_8_452_90_0 & ~i_8_452_241_0 & ~i_8_452_402_0 & i_8_452_652_0 & ~i_8_452_1383_0 & ~i_8_452_1708_0) | (~i_8_452_691_0 & ~i_8_452_768_0 & ~i_8_452_795_0 & ~i_8_452_839_0 & ~i_8_452_1844_0 & ~i_8_452_2178_0 & ~i_8_452_1338_0 & i_8_452_1776_0))) | (~i_8_452_45_0 & ~i_8_452_166_0 & i_8_452_362_0 & ~i_8_452_1410_0 & ~i_8_452_1835_0 & ~i_8_452_2227_0))) | (i_8_452_839_0 & i_8_452_877_0 & i_8_452_1156_0 & i_8_452_1776_0) | (~i_8_452_194_0 & i_8_452_602_0 & ~i_8_452_1330_0 & ~i_8_452_1673_0 & ~i_8_452_1705_0 & ~i_8_452_1835_0 & ~i_8_452_1987_0) | (i_8_452_194_0 & i_8_452_301_0 & ~i_8_452_528_0 & ~i_8_452_1329_0 & ~i_8_452_1356_0 & ~i_8_452_1410_0 & ~i_8_452_1844_0 & ~i_8_452_1862_0 & ~i_8_452_2112_0))) | (i_8_452_194_0 & ((~i_8_452_340_0 & i_8_452_853_0 & ~i_8_452_1819_0) | (~i_8_452_90_0 & ~i_8_452_691_0 & ~i_8_452_765_0 & i_8_452_877_0 & ~i_8_452_1295_0 & ~i_8_452_1384_0 & ~i_8_452_1407_0 & ~i_8_452_2022_0))) | (~i_8_452_1295_0 & ((~i_8_452_194_0 & ((~i_8_452_60_0 & ~i_8_452_301_0 & ~i_8_452_340_0 & i_8_452_529_0 & i_8_452_691_0 & ~i_8_452_1321_0 & ~i_8_452_1625_0) | (~i_8_452_44_0 & ~i_8_452_166_0 & i_8_452_301_0 & ~i_8_452_768_0 & i_8_452_853_0 & ~i_8_452_1156_0 & ~i_8_452_1673_0 & ~i_8_452_2016_0))) | (~i_8_452_839_0 & ~i_8_452_853_0 & ~i_8_452_1435_0 & i_8_452_1673_0 & ~i_8_452_1844_0 & ~i_8_452_2227_0))) | (~i_8_452_765_0 & ((~i_8_452_45_0 & i_8_452_301_0 & ~i_8_452_1330_0 & ~i_8_452_1384_0 & ((~i_8_452_529_0 & ~i_8_452_768_0 & ~i_8_452_795_0 & i_8_452_877_0 & ~i_8_452_1862_0) | (~i_8_452_402_0 & ~i_8_452_660_0 & ~i_8_452_665_0 & ~i_8_452_844_0 & ~i_8_452_857_0 & ~i_8_452_1105_0 & ~i_8_452_1708_0 & ~i_8_452_1834_0 & ~i_8_452_2022_0 & ~i_8_452_2112_0 & ~i_8_452_2178_0 & ~i_8_452_2227_0))) | (i_8_452_528_0 & ((~i_8_452_44_0 & i_8_452_529_0 & i_8_452_717_0 & i_8_452_1033_0) | (i_8_452_654_0 & ~i_8_452_691_0 & ~i_8_452_1834_0))) | (~i_8_452_44_0 & ((~i_8_452_528_0 & ~i_8_452_651_0 & i_8_452_665_0 & ~i_8_452_1132_0 & ~i_8_452_1331_0 & ~i_8_452_1407_0 & i_8_452_1435_0 & ~i_8_452_1708_0 & ~i_8_452_1818_0 & ~i_8_452_2112_0) | (~i_8_452_341_0 & i_8_452_601_0 & ~i_8_452_1329_0 & ~i_8_452_1835_0 & ~i_8_452_1995_0 & ~i_8_452_2244_0))) | (~i_8_452_665_0 & ((~i_8_452_90_0 & ~i_8_452_651_0 & ~i_8_452_691_0 & i_8_452_719_0 & ~i_8_452_1338_0 & ~i_8_452_1705_0 & ~i_8_452_1942_0) | (~i_8_452_340_0 & i_8_452_717_0 & ~i_8_452_2109_0))) | (~i_8_452_90_0 & ((i_8_452_45_0 & i_8_452_877_0 & ~i_8_452_1407_0 & ~i_8_452_1435_0 & i_8_452_1818_0 & ~i_8_452_1819_0) | (~i_8_452_660_0 & ~i_8_452_877_0 & ~i_8_452_1339_0 & i_8_452_1776_0 & ~i_8_452_1821_0 & ~i_8_452_2109_0))))) | (~i_8_452_1383_0 & ((~i_8_452_90_0 & ~i_8_452_2178_0 & ((~i_8_452_44_0 & ~i_8_452_691_0 & i_8_452_1033_0 & ~i_8_452_1330_0 & ~i_8_452_2022_0) | (~i_8_452_529_0 & i_8_452_651_0 & ~i_8_452_1156_0 & ~i_8_452_1314_0 & ~i_8_452_1322_0 & ~i_8_452_1329_0 & ~i_8_452_1834_0 & ~i_8_452_2016_0 & ~i_8_452_2227_0))) | (~i_8_452_340_0 & ~i_8_452_1407_0 & ((~i_8_452_70_0 & i_8_452_224_0 & ~i_8_452_857_0 & i_8_452_881_0 & ~i_8_452_2022_0) | (~i_8_452_301_0 & ~i_8_452_880_0 & ~i_8_452_1435_0 & ~i_8_452_1818_0 & i_8_452_2244_0))) | (~i_8_452_654_0 & ~i_8_452_665_0 & i_8_452_717_0 & ~i_8_452_836_0 & ~i_8_452_844_0 & ~i_8_452_1384_0 & ~i_8_452_1834_0 & ~i_8_452_1942_0 & ~i_8_452_2016_0))) | (~i_8_452_839_0 & ((~i_8_452_227_0 & ~i_8_452_341_0 & i_8_452_836_0 & ~i_8_452_1331_0 & ~i_8_452_1834_0 & ~i_8_452_2151_0) | (i_8_452_362_0 & ~i_8_452_857_0 & ~i_8_452_1156_0 & ~i_8_452_1835_0 & ~i_8_452_2227_0))) | (~i_8_452_1105_0 & ((~i_8_452_241_0 & ~i_8_452_672_0 & ~i_8_452_1321_0 & ~i_8_452_1339_0 & ~i_8_452_1835_0 & ~i_8_452_2022_0 & i_8_452_2096_0 & ~i_8_452_2171_0) | (i_8_452_653_0 & ~i_8_452_665_0 & ~i_8_452_1331_0 & ~i_8_452_1834_0 & ~i_8_452_2178_0))) | (~i_8_452_2178_0 & ((~i_8_452_301_0 & i_8_452_628_0 & ~i_8_452_691_0 & ~i_8_452_857_0 & ~i_8_452_2022_0 & ~i_8_452_2109_0 & ~i_8_452_1384_0 & i_8_452_1776_0) | (~i_8_452_402_0 & i_8_452_719_0 & ~i_8_452_1625_0 & i_8_452_2096_0 & ~i_8_452_2151_0))) | (~i_8_452_45_0 & ~i_8_452_795_0 & ~i_8_452_853_0 & ~i_8_452_877_0 & ~i_8_452_1321_0 & ~i_8_452_1329_0 & i_8_452_1818_0 & i_8_452_1821_0) | (~i_8_452_340_0 & i_8_452_529_0 & i_8_452_665_0 & ~i_8_452_1331_0 & i_8_452_1844_0) | (i_8_452_839_0 & ~i_8_452_880_0 & ~i_8_452_1835_0 & i_8_452_1862_0 & ~i_8_452_1987_0));
endmodule



// Benchmark "kernel_8_453" written by ABC on Sun Jul 19 10:11:03 2020

module kernel_8_453 ( 
    i_8_453_21_0, i_8_453_24_0, i_8_453_30_0, i_8_453_39_0, i_8_453_43_0,
    i_8_453_115_0, i_8_453_120_0, i_8_453_121_0, i_8_453_124_0,
    i_8_453_129_0, i_8_453_140_0, i_8_453_150_0, i_8_453_160_0,
    i_8_453_175_0, i_8_453_273_0, i_8_453_276_0, i_8_453_309_0,
    i_8_453_310_0, i_8_453_324_0, i_8_453_345_0, i_8_453_348_0,
    i_8_453_351_0, i_8_453_354_0, i_8_453_365_0, i_8_453_378_0,
    i_8_453_387_0, i_8_453_426_0, i_8_453_529_0, i_8_453_553_0,
    i_8_453_555_0, i_8_453_624_0, i_8_453_625_0, i_8_453_643_0,
    i_8_453_652_0, i_8_453_654_0, i_8_453_672_0, i_8_453_673_0,
    i_8_453_697_0, i_8_453_741_0, i_8_453_762_0, i_8_453_768_0,
    i_8_453_829_0, i_8_453_833_0, i_8_453_841_0, i_8_453_848_0,
    i_8_453_854_0, i_8_453_877_0, i_8_453_881_0, i_8_453_915_0,
    i_8_453_943_0, i_8_453_944_0, i_8_453_951_0, i_8_453_954_0,
    i_8_453_969_0, i_8_453_987_0, i_8_453_1012_0, i_8_453_1203_0,
    i_8_453_1270_0, i_8_453_1271_0, i_8_453_1285_0, i_8_453_1324_0,
    i_8_453_1410_0, i_8_453_1432_0, i_8_453_1474_0, i_8_453_1479_0,
    i_8_453_1482_0, i_8_453_1492_0, i_8_453_1545_0, i_8_453_1546_0,
    i_8_453_1571_0, i_8_453_1580_0, i_8_453_1605_0, i_8_453_1606_0,
    i_8_453_1623_0, i_8_453_1641_0, i_8_453_1644_0, i_8_453_1660_0,
    i_8_453_1705_0, i_8_453_1749_0, i_8_453_1765_0, i_8_453_1806_0,
    i_8_453_1821_0, i_8_453_1848_0, i_8_453_1912_0, i_8_453_1951_0,
    i_8_453_1962_0, i_8_453_1969_0, i_8_453_1971_0, i_8_453_2011_0,
    i_8_453_2046_0, i_8_453_2064_0, i_8_453_2086_0, i_8_453_2094_0,
    i_8_453_2104_0, i_8_453_2215_0, i_8_453_2224_0, i_8_453_2245_0,
    i_8_453_2257_0, i_8_453_2272_0, i_8_453_2298_0,
    o_8_453_0_0  );
  input  i_8_453_21_0, i_8_453_24_0, i_8_453_30_0, i_8_453_39_0,
    i_8_453_43_0, i_8_453_115_0, i_8_453_120_0, i_8_453_121_0,
    i_8_453_124_0, i_8_453_129_0, i_8_453_140_0, i_8_453_150_0,
    i_8_453_160_0, i_8_453_175_0, i_8_453_273_0, i_8_453_276_0,
    i_8_453_309_0, i_8_453_310_0, i_8_453_324_0, i_8_453_345_0,
    i_8_453_348_0, i_8_453_351_0, i_8_453_354_0, i_8_453_365_0,
    i_8_453_378_0, i_8_453_387_0, i_8_453_426_0, i_8_453_529_0,
    i_8_453_553_0, i_8_453_555_0, i_8_453_624_0, i_8_453_625_0,
    i_8_453_643_0, i_8_453_652_0, i_8_453_654_0, i_8_453_672_0,
    i_8_453_673_0, i_8_453_697_0, i_8_453_741_0, i_8_453_762_0,
    i_8_453_768_0, i_8_453_829_0, i_8_453_833_0, i_8_453_841_0,
    i_8_453_848_0, i_8_453_854_0, i_8_453_877_0, i_8_453_881_0,
    i_8_453_915_0, i_8_453_943_0, i_8_453_944_0, i_8_453_951_0,
    i_8_453_954_0, i_8_453_969_0, i_8_453_987_0, i_8_453_1012_0,
    i_8_453_1203_0, i_8_453_1270_0, i_8_453_1271_0, i_8_453_1285_0,
    i_8_453_1324_0, i_8_453_1410_0, i_8_453_1432_0, i_8_453_1474_0,
    i_8_453_1479_0, i_8_453_1482_0, i_8_453_1492_0, i_8_453_1545_0,
    i_8_453_1546_0, i_8_453_1571_0, i_8_453_1580_0, i_8_453_1605_0,
    i_8_453_1606_0, i_8_453_1623_0, i_8_453_1641_0, i_8_453_1644_0,
    i_8_453_1660_0, i_8_453_1705_0, i_8_453_1749_0, i_8_453_1765_0,
    i_8_453_1806_0, i_8_453_1821_0, i_8_453_1848_0, i_8_453_1912_0,
    i_8_453_1951_0, i_8_453_1962_0, i_8_453_1969_0, i_8_453_1971_0,
    i_8_453_2011_0, i_8_453_2046_0, i_8_453_2064_0, i_8_453_2086_0,
    i_8_453_2094_0, i_8_453_2104_0, i_8_453_2215_0, i_8_453_2224_0,
    i_8_453_2245_0, i_8_453_2257_0, i_8_453_2272_0, i_8_453_2298_0;
  output o_8_453_0_0;
  assign o_8_453_0_0 = 0;
endmodule



// Benchmark "kernel_8_454" written by ABC on Sun Jul 19 10:11:05 2020

module kernel_8_454 ( 
    i_8_454_37_0, i_8_454_38_0, i_8_454_59_0, i_8_454_64_0, i_8_454_65_0,
    i_8_454_172_0, i_8_454_173_0, i_8_454_182_0, i_8_454_225_0,
    i_8_454_227_0, i_8_454_319_0, i_8_454_325_0, i_8_454_353_0,
    i_8_454_379_0, i_8_454_380_0, i_8_454_401_0, i_8_454_493_0,
    i_8_454_584_0, i_8_454_617_0, i_8_454_620_0, i_8_454_657_0,
    i_8_454_665_0, i_8_454_703_0, i_8_454_704_0, i_8_454_707_0,
    i_8_454_765_0, i_8_454_777_0, i_8_454_840_0, i_8_454_842_0,
    i_8_454_873_0, i_8_454_875_0, i_8_454_877_0, i_8_454_882_0,
    i_8_454_884_0, i_8_454_932_0, i_8_454_956_0, i_8_454_965_0,
    i_8_454_991_0, i_8_454_993_0, i_8_454_995_0, i_8_454_1026_0,
    i_8_454_1028_0, i_8_454_1031_0, i_8_454_1073_0, i_8_454_1103_0,
    i_8_454_1171_0, i_8_454_1172_0, i_8_454_1175_0, i_8_454_1199_0,
    i_8_454_1225_0, i_8_454_1234_0, i_8_454_1238_0, i_8_454_1315_0,
    i_8_454_1354_0, i_8_454_1381_0, i_8_454_1382_0, i_8_454_1397_0,
    i_8_454_1434_0, i_8_454_1439_0, i_8_454_1460_0, i_8_454_1468_0,
    i_8_454_1469_0, i_8_454_1489_0, i_8_454_1505_0, i_8_454_1543_0,
    i_8_454_1544_0, i_8_454_1552_0, i_8_454_1648_0, i_8_454_1654_0,
    i_8_454_1675_0, i_8_454_1676_0, i_8_454_1678_0, i_8_454_1679_0,
    i_8_454_1702_0, i_8_454_1703_0, i_8_454_1706_0, i_8_454_1746_0,
    i_8_454_1749_0, i_8_454_1777_0, i_8_454_1778_0, i_8_454_1792_0,
    i_8_454_1804_0, i_8_454_1819_0, i_8_454_1820_0, i_8_454_1823_0,
    i_8_454_1855_0, i_8_454_1910_0, i_8_454_1913_0, i_8_454_1918_0,
    i_8_454_1936_0, i_8_454_1943_0, i_8_454_2053_0, i_8_454_2099_0,
    i_8_454_2143_0, i_8_454_2144_0, i_8_454_2147_0, i_8_454_2168_0,
    i_8_454_2183_0, i_8_454_2210_0, i_8_454_2287_0,
    o_8_454_0_0  );
  input  i_8_454_37_0, i_8_454_38_0, i_8_454_59_0, i_8_454_64_0,
    i_8_454_65_0, i_8_454_172_0, i_8_454_173_0, i_8_454_182_0,
    i_8_454_225_0, i_8_454_227_0, i_8_454_319_0, i_8_454_325_0,
    i_8_454_353_0, i_8_454_379_0, i_8_454_380_0, i_8_454_401_0,
    i_8_454_493_0, i_8_454_584_0, i_8_454_617_0, i_8_454_620_0,
    i_8_454_657_0, i_8_454_665_0, i_8_454_703_0, i_8_454_704_0,
    i_8_454_707_0, i_8_454_765_0, i_8_454_777_0, i_8_454_840_0,
    i_8_454_842_0, i_8_454_873_0, i_8_454_875_0, i_8_454_877_0,
    i_8_454_882_0, i_8_454_884_0, i_8_454_932_0, i_8_454_956_0,
    i_8_454_965_0, i_8_454_991_0, i_8_454_993_0, i_8_454_995_0,
    i_8_454_1026_0, i_8_454_1028_0, i_8_454_1031_0, i_8_454_1073_0,
    i_8_454_1103_0, i_8_454_1171_0, i_8_454_1172_0, i_8_454_1175_0,
    i_8_454_1199_0, i_8_454_1225_0, i_8_454_1234_0, i_8_454_1238_0,
    i_8_454_1315_0, i_8_454_1354_0, i_8_454_1381_0, i_8_454_1382_0,
    i_8_454_1397_0, i_8_454_1434_0, i_8_454_1439_0, i_8_454_1460_0,
    i_8_454_1468_0, i_8_454_1469_0, i_8_454_1489_0, i_8_454_1505_0,
    i_8_454_1543_0, i_8_454_1544_0, i_8_454_1552_0, i_8_454_1648_0,
    i_8_454_1654_0, i_8_454_1675_0, i_8_454_1676_0, i_8_454_1678_0,
    i_8_454_1679_0, i_8_454_1702_0, i_8_454_1703_0, i_8_454_1706_0,
    i_8_454_1746_0, i_8_454_1749_0, i_8_454_1777_0, i_8_454_1778_0,
    i_8_454_1792_0, i_8_454_1804_0, i_8_454_1819_0, i_8_454_1820_0,
    i_8_454_1823_0, i_8_454_1855_0, i_8_454_1910_0, i_8_454_1913_0,
    i_8_454_1918_0, i_8_454_1936_0, i_8_454_1943_0, i_8_454_2053_0,
    i_8_454_2099_0, i_8_454_2143_0, i_8_454_2144_0, i_8_454_2147_0,
    i_8_454_2168_0, i_8_454_2183_0, i_8_454_2210_0, i_8_454_2287_0;
  output o_8_454_0_0;
  assign o_8_454_0_0 = ~((~i_8_454_840_0 & ((~i_8_454_319_0 & ~i_8_454_842_0 & ((i_8_454_617_0 & ~i_8_454_995_0 & ~i_8_454_1172_0 & ~i_8_454_1225_0 & ~i_8_454_1505_0 & ~i_8_454_1703_0 & ~i_8_454_1910_0 & i_8_454_1918_0 & ~i_8_454_1943_0) | (~i_8_454_173_0 & ~i_8_454_182_0 & ~i_8_454_379_0 & ~i_8_454_380_0 & ~i_8_454_956_0 & ~i_8_454_993_0 & ~i_8_454_1028_0 & ~i_8_454_1103_0 & ~i_8_454_1439_0 & ~i_8_454_1460_0 & ~i_8_454_1792_0 & ~i_8_454_2168_0))) | (~i_8_454_704_0 & ~i_8_454_1382_0 & ~i_8_454_1397_0 & ~i_8_454_1706_0 & i_8_454_1778_0 & i_8_454_1804_0 & ~i_8_454_2210_0))) | (~i_8_454_1382_0 & ((~i_8_454_64_0 & ((~i_8_454_38_0 & ~i_8_454_173_0 & ~i_8_454_182_0 & i_8_454_877_0 & ~i_8_454_1175_0 & ~i_8_454_1238_0 & ~i_8_454_1460_0 & ~i_8_454_1792_0) | (~i_8_454_37_0 & ~i_8_454_617_0 & ~i_8_454_665_0 & ~i_8_454_956_0 & ~i_8_454_1026_0 & ~i_8_454_1103_0 & ~i_8_454_1552_0 & ~i_8_454_1703_0 & ~i_8_454_1804_0 & ~i_8_454_1910_0))) | (~i_8_454_1792_0 & ((~i_8_454_1913_0 & ((~i_8_454_37_0 & ~i_8_454_2183_0 & ((~i_8_454_173_0 & ~i_8_454_765_0 & i_8_454_840_0 & ~i_8_454_1238_0) | (~i_8_454_38_0 & ~i_8_454_182_0 & ~i_8_454_584_0 & ~i_8_454_932_0 & ~i_8_454_1031_0 & ~i_8_454_1073_0 & ~i_8_454_1171_0 & ~i_8_454_1910_0 & ~i_8_454_1943_0))) | (~i_8_454_1943_0 & ((~i_8_454_173_0 & ~i_8_454_401_0 & ~i_8_454_965_0 & ~i_8_454_1028_0 & ~i_8_454_1315_0 & ~i_8_454_1648_0 & i_8_454_1778_0 & ~i_8_454_1910_0) | (~i_8_454_38_0 & i_8_454_703_0 & ~i_8_454_1225_0 & ~i_8_454_2210_0))))) | (~i_8_454_37_0 & ~i_8_454_65_0 & i_8_454_1552_0 & ~i_8_454_1703_0 & i_8_454_1777_0 & ~i_8_454_2168_0 & ~i_8_454_2210_0))) | (~i_8_454_65_0 & ~i_8_454_584_0 & ~i_8_454_1702_0 & ((~i_8_454_932_0 & ~i_8_454_1703_0 & i_8_454_1820_0 & ~i_8_454_2144_0) | (~i_8_454_37_0 & ~i_8_454_704_0 & ~i_8_454_1238_0 & ~i_8_454_1381_0 & ~i_8_454_2147_0))))) | (~i_8_454_64_0 & ((~i_8_454_37_0 & ((~i_8_454_873_0 & i_8_454_875_0 & ~i_8_454_965_0 & ~i_8_454_1439_0 & i_8_454_1823_0) | (~i_8_454_65_0 & ~i_8_454_932_0 & i_8_454_1679_0 & ~i_8_454_1913_0 & ~i_8_454_2147_0))) | (i_8_454_1749_0 & ~i_8_454_2147_0))) | (~i_8_454_65_0 & ~i_8_454_620_0 & ((~i_8_454_173_0 & ~i_8_454_493_0 & ~i_8_454_584_0 & ~i_8_454_1172_0 & ~i_8_454_1175_0 & ~i_8_454_1654_0 & ~i_8_454_1819_0 & ~i_8_454_1820_0 & ~i_8_454_1936_0 & ~i_8_454_2144_0) | (~i_8_454_379_0 & ~i_8_454_617_0 & ~i_8_454_1234_0 & ~i_8_454_1469_0 & ~i_8_454_1648_0 & ~i_8_454_1706_0 & i_8_454_1823_0 & ~i_8_454_1943_0 & i_8_454_2147_0))) | (~i_8_454_401_0 & ((~i_8_454_665_0 & ~i_8_454_956_0 & ~i_8_454_1397_0 & i_8_454_1678_0 & ~i_8_454_1702_0 & ~i_8_454_1703_0 & ~i_8_454_1910_0) | (i_8_454_620_0 & ~i_8_454_1073_0 & ~i_8_454_1238_0 & ~i_8_454_1706_0 & ~i_8_454_1819_0 & i_8_454_1823_0 & ~i_8_454_1913_0))) | (~i_8_454_2183_0 & ((~i_8_454_493_0 & ~i_8_454_932_0 & ((~i_8_454_173_0 & ~i_8_454_584_0 & ~i_8_454_657_0 & ~i_8_454_1175_0 & ~i_8_454_1439_0 & ~i_8_454_1469_0 & ~i_8_454_1489_0 & ~i_8_454_1505_0 & ~i_8_454_1552_0 & ~i_8_454_1648_0 & ~i_8_454_1706_0) | (~i_8_454_617_0 & ~i_8_454_704_0 & ~i_8_454_965_0 & ~i_8_454_995_0 & ~i_8_454_1172_0 & ~i_8_454_1702_0 & ~i_8_454_1943_0))) | (~i_8_454_1172_0 & ~i_8_454_1175_0 & ~i_8_454_1234_0 & i_8_454_1552_0 & ~i_8_454_1703_0 & ~i_8_454_1823_0 & ~i_8_454_1910_0 & ~i_8_454_2168_0))) | (~i_8_454_1910_0 & ((~i_8_454_173_0 & ((~i_8_454_584_0 & ~i_8_454_707_0 & i_8_454_995_0 & ~i_8_454_1172_0) | (~i_8_454_703_0 & ~i_8_454_1073_0 & i_8_454_1234_0 & ~i_8_454_1354_0 & ~i_8_454_1489_0 & ~i_8_454_1823_0))) | (i_8_454_379_0 & ~i_8_454_1381_0 & ~i_8_454_1544_0 & ~i_8_454_1702_0 & ~i_8_454_1820_0 & ~i_8_454_1913_0 & ~i_8_454_2210_0))) | (~i_8_454_1103_0 & ~i_8_454_1354_0 & ~i_8_454_1468_0 & i_8_454_1505_0 & i_8_454_1679_0 & ~i_8_454_1703_0));
endmodule



// Benchmark "kernel_8_455" written by ABC on Sun Jul 19 10:11:05 2020

module kernel_8_455 ( 
    i_8_455_7_0, i_8_455_26_0, i_8_455_79_0, i_8_455_86_0, i_8_455_134_0,
    i_8_455_140_0, i_8_455_184_0, i_8_455_206_0, i_8_455_250_0,
    i_8_455_314_0, i_8_455_359_0, i_8_455_366_0, i_8_455_401_0,
    i_8_455_499_0, i_8_455_521_0, i_8_455_529_0, i_8_455_539_0,
    i_8_455_556_0, i_8_455_575_0, i_8_455_583_0, i_8_455_601_0,
    i_8_455_611_0, i_8_455_652_0, i_8_455_656_0, i_8_455_664_0,
    i_8_455_665_0, i_8_455_719_0, i_8_455_737_0, i_8_455_754_0,
    i_8_455_763_0, i_8_455_781_0, i_8_455_789_0, i_8_455_844_0,
    i_8_455_886_0, i_8_455_896_0, i_8_455_917_0, i_8_455_923_0,
    i_8_455_959_0, i_8_455_962_0, i_8_455_968_0, i_8_455_1015_0,
    i_8_455_1075_0, i_8_455_1078_0, i_8_455_1088_0, i_8_455_1195_0,
    i_8_455_1196_0, i_8_455_1201_0, i_8_455_1205_0, i_8_455_1230_0,
    i_8_455_1339_0, i_8_455_1384_0, i_8_455_1385_0, i_8_455_1393_0,
    i_8_455_1394_0, i_8_455_1403_0, i_8_455_1410_0, i_8_455_1466_0,
    i_8_455_1484_0, i_8_455_1492_0, i_8_455_1502_0, i_8_455_1517_0,
    i_8_455_1528_0, i_8_455_1573_0, i_8_455_1601_0, i_8_455_1636_0,
    i_8_455_1646_0, i_8_455_1652_0, i_8_455_1663_0, i_8_455_1664_0,
    i_8_455_1700_0, i_8_455_1717_0, i_8_455_1718_0, i_8_455_1727_0,
    i_8_455_1753_0, i_8_455_1781_0, i_8_455_1826_0, i_8_455_1844_0,
    i_8_455_1852_0, i_8_455_1879_0, i_8_455_1880_0, i_8_455_1885_0,
    i_8_455_1922_0, i_8_455_1929_0, i_8_455_1939_0, i_8_455_1979_0,
    i_8_455_2015_0, i_8_455_2060_0, i_8_455_2065_0, i_8_455_2094_0,
    i_8_455_2146_0, i_8_455_2149_0, i_8_455_2150_0, i_8_455_2174_0,
    i_8_455_2177_0, i_8_455_2185_0, i_8_455_2214_0, i_8_455_2217_0,
    i_8_455_2218_0, i_8_455_2231_0, i_8_455_2240_0,
    o_8_455_0_0  );
  input  i_8_455_7_0, i_8_455_26_0, i_8_455_79_0, i_8_455_86_0,
    i_8_455_134_0, i_8_455_140_0, i_8_455_184_0, i_8_455_206_0,
    i_8_455_250_0, i_8_455_314_0, i_8_455_359_0, i_8_455_366_0,
    i_8_455_401_0, i_8_455_499_0, i_8_455_521_0, i_8_455_529_0,
    i_8_455_539_0, i_8_455_556_0, i_8_455_575_0, i_8_455_583_0,
    i_8_455_601_0, i_8_455_611_0, i_8_455_652_0, i_8_455_656_0,
    i_8_455_664_0, i_8_455_665_0, i_8_455_719_0, i_8_455_737_0,
    i_8_455_754_0, i_8_455_763_0, i_8_455_781_0, i_8_455_789_0,
    i_8_455_844_0, i_8_455_886_0, i_8_455_896_0, i_8_455_917_0,
    i_8_455_923_0, i_8_455_959_0, i_8_455_962_0, i_8_455_968_0,
    i_8_455_1015_0, i_8_455_1075_0, i_8_455_1078_0, i_8_455_1088_0,
    i_8_455_1195_0, i_8_455_1196_0, i_8_455_1201_0, i_8_455_1205_0,
    i_8_455_1230_0, i_8_455_1339_0, i_8_455_1384_0, i_8_455_1385_0,
    i_8_455_1393_0, i_8_455_1394_0, i_8_455_1403_0, i_8_455_1410_0,
    i_8_455_1466_0, i_8_455_1484_0, i_8_455_1492_0, i_8_455_1502_0,
    i_8_455_1517_0, i_8_455_1528_0, i_8_455_1573_0, i_8_455_1601_0,
    i_8_455_1636_0, i_8_455_1646_0, i_8_455_1652_0, i_8_455_1663_0,
    i_8_455_1664_0, i_8_455_1700_0, i_8_455_1717_0, i_8_455_1718_0,
    i_8_455_1727_0, i_8_455_1753_0, i_8_455_1781_0, i_8_455_1826_0,
    i_8_455_1844_0, i_8_455_1852_0, i_8_455_1879_0, i_8_455_1880_0,
    i_8_455_1885_0, i_8_455_1922_0, i_8_455_1929_0, i_8_455_1939_0,
    i_8_455_1979_0, i_8_455_2015_0, i_8_455_2060_0, i_8_455_2065_0,
    i_8_455_2094_0, i_8_455_2146_0, i_8_455_2149_0, i_8_455_2150_0,
    i_8_455_2174_0, i_8_455_2177_0, i_8_455_2185_0, i_8_455_2214_0,
    i_8_455_2217_0, i_8_455_2218_0, i_8_455_2231_0, i_8_455_2240_0;
  output o_8_455_0_0;
  assign o_8_455_0_0 = 0;
endmodule



// Benchmark "kernel_8_456" written by ABC on Sun Jul 19 10:11:06 2020

module kernel_8_456 ( 
    i_8_456_12_0, i_8_456_22_0, i_8_456_28_0, i_8_456_31_0, i_8_456_33_0,
    i_8_456_50_0, i_8_456_54_0, i_8_456_55_0, i_8_456_56_0, i_8_456_76_0,
    i_8_456_103_0, i_8_456_105_0, i_8_456_136_0, i_8_456_139_0,
    i_8_456_195_0, i_8_456_299_0, i_8_456_430_0, i_8_456_441_0,
    i_8_456_523_0, i_8_456_529_0, i_8_456_543_0, i_8_456_552_0,
    i_8_456_606_0, i_8_456_608_0, i_8_456_610_0, i_8_456_615_0,
    i_8_456_631_0, i_8_456_652_0, i_8_456_678_0, i_8_456_708_0,
    i_8_456_729_0, i_8_456_750_0, i_8_456_751_0, i_8_456_760_0,
    i_8_456_762_0, i_8_456_783_0, i_8_456_811_0, i_8_456_814_0,
    i_8_456_840_0, i_8_456_860_0, i_8_456_876_0, i_8_456_891_0,
    i_8_456_940_0, i_8_456_1050_0, i_8_456_1090_0, i_8_456_1104_0,
    i_8_456_1108_0, i_8_456_1111_0, i_8_456_1112_0, i_8_456_1139_0,
    i_8_456_1246_0, i_8_456_1254_0, i_8_456_1255_0, i_8_456_1294_0,
    i_8_456_1308_0, i_8_456_1309_0, i_8_456_1314_0, i_8_456_1324_0,
    i_8_456_1331_0, i_8_456_1334_0, i_8_456_1337_0, i_8_456_1362_0,
    i_8_456_1399_0, i_8_456_1422_0, i_8_456_1435_0, i_8_456_1441_0,
    i_8_456_1477_0, i_8_456_1480_0, i_8_456_1512_0, i_8_456_1513_0,
    i_8_456_1615_0, i_8_456_1632_0, i_8_456_1634_0, i_8_456_1635_0,
    i_8_456_1680_0, i_8_456_1682_0, i_8_456_1705_0, i_8_456_1714_0,
    i_8_456_1746_0, i_8_456_1756_0, i_8_456_1757_0, i_8_456_1784_0,
    i_8_456_1857_0, i_8_456_1885_0, i_8_456_1902_0, i_8_456_1904_0,
    i_8_456_1912_0, i_8_456_1926_0, i_8_456_1948_0, i_8_456_1975_0,
    i_8_456_1981_0, i_8_456_1993_0, i_8_456_2029_0, i_8_456_2053_0,
    i_8_456_2098_0, i_8_456_2149_0, i_8_456_2236_0, i_8_456_2273_0,
    i_8_456_2286_0, i_8_456_2295_0,
    o_8_456_0_0  );
  input  i_8_456_12_0, i_8_456_22_0, i_8_456_28_0, i_8_456_31_0,
    i_8_456_33_0, i_8_456_50_0, i_8_456_54_0, i_8_456_55_0, i_8_456_56_0,
    i_8_456_76_0, i_8_456_103_0, i_8_456_105_0, i_8_456_136_0,
    i_8_456_139_0, i_8_456_195_0, i_8_456_299_0, i_8_456_430_0,
    i_8_456_441_0, i_8_456_523_0, i_8_456_529_0, i_8_456_543_0,
    i_8_456_552_0, i_8_456_606_0, i_8_456_608_0, i_8_456_610_0,
    i_8_456_615_0, i_8_456_631_0, i_8_456_652_0, i_8_456_678_0,
    i_8_456_708_0, i_8_456_729_0, i_8_456_750_0, i_8_456_751_0,
    i_8_456_760_0, i_8_456_762_0, i_8_456_783_0, i_8_456_811_0,
    i_8_456_814_0, i_8_456_840_0, i_8_456_860_0, i_8_456_876_0,
    i_8_456_891_0, i_8_456_940_0, i_8_456_1050_0, i_8_456_1090_0,
    i_8_456_1104_0, i_8_456_1108_0, i_8_456_1111_0, i_8_456_1112_0,
    i_8_456_1139_0, i_8_456_1246_0, i_8_456_1254_0, i_8_456_1255_0,
    i_8_456_1294_0, i_8_456_1308_0, i_8_456_1309_0, i_8_456_1314_0,
    i_8_456_1324_0, i_8_456_1331_0, i_8_456_1334_0, i_8_456_1337_0,
    i_8_456_1362_0, i_8_456_1399_0, i_8_456_1422_0, i_8_456_1435_0,
    i_8_456_1441_0, i_8_456_1477_0, i_8_456_1480_0, i_8_456_1512_0,
    i_8_456_1513_0, i_8_456_1615_0, i_8_456_1632_0, i_8_456_1634_0,
    i_8_456_1635_0, i_8_456_1680_0, i_8_456_1682_0, i_8_456_1705_0,
    i_8_456_1714_0, i_8_456_1746_0, i_8_456_1756_0, i_8_456_1757_0,
    i_8_456_1784_0, i_8_456_1857_0, i_8_456_1885_0, i_8_456_1902_0,
    i_8_456_1904_0, i_8_456_1912_0, i_8_456_1926_0, i_8_456_1948_0,
    i_8_456_1975_0, i_8_456_1981_0, i_8_456_1993_0, i_8_456_2029_0,
    i_8_456_2053_0, i_8_456_2098_0, i_8_456_2149_0, i_8_456_2236_0,
    i_8_456_2273_0, i_8_456_2286_0, i_8_456_2295_0;
  output o_8_456_0_0;
  assign o_8_456_0_0 = 0;
endmodule



// Benchmark "kernel_8_457" written by ABC on Sun Jul 19 10:11:08 2020

module kernel_8_457 ( 
    i_8_457_19_0, i_8_457_46_0, i_8_457_67_0, i_8_457_70_0, i_8_457_88_0,
    i_8_457_136_0, i_8_457_232_0, i_8_457_252_0, i_8_457_255_0,
    i_8_457_343_0, i_8_457_350_0, i_8_457_378_0, i_8_457_379_0,
    i_8_457_429_0, i_8_457_430_0, i_8_457_450_0, i_8_457_454_0,
    i_8_457_484_0, i_8_457_496_0, i_8_457_507_0, i_8_457_556_0,
    i_8_457_585_0, i_8_457_586_0, i_8_457_610_0, i_8_457_634_0,
    i_8_457_655_0, i_8_457_699_0, i_8_457_702_0, i_8_457_703_0,
    i_8_457_708_0, i_8_457_709_0, i_8_457_718_0, i_8_457_733_0,
    i_8_457_814_0, i_8_457_841_0, i_8_457_879_0, i_8_457_880_0,
    i_8_457_889_0, i_8_457_978_0, i_8_457_979_0, i_8_457_996_0,
    i_8_457_1032_0, i_8_457_1078_0, i_8_457_1140_0, i_8_457_1141_0,
    i_8_457_1144_0, i_8_457_1149_0, i_8_457_1150_0, i_8_457_1168_0,
    i_8_457_1171_0, i_8_457_1227_0, i_8_457_1239_0, i_8_457_1240_0,
    i_8_457_1251_0, i_8_457_1264_0, i_8_457_1273_0, i_8_457_1275_0,
    i_8_457_1278_0, i_8_457_1356_0, i_8_457_1357_0, i_8_457_1359_0,
    i_8_457_1410_0, i_8_457_1412_0, i_8_457_1547_0, i_8_457_1602_0,
    i_8_457_1603_0, i_8_457_1604_0, i_8_457_1632_0, i_8_457_1637_0,
    i_8_457_1779_0, i_8_457_1803_0, i_8_457_1819_0, i_8_457_1824_0,
    i_8_457_1869_0, i_8_457_1986_0, i_8_457_1996_0, i_8_457_2058_0,
    i_8_457_2059_0, i_8_457_2107_0, i_8_457_2146_0, i_8_457_2148_0,
    i_8_457_2149_0, i_8_457_2150_0, i_8_457_2152_0, i_8_457_2157_0,
    i_8_457_2175_0, i_8_457_2176_0, i_8_457_2233_0, i_8_457_2238_0,
    i_8_457_2241_0, i_8_457_2242_0, i_8_457_2243_0, i_8_457_2244_0,
    i_8_457_2248_0, i_8_457_2260_0, i_8_457_2263_0, i_8_457_2272_0,
    i_8_457_2273_0, i_8_457_2301_0, i_8_457_2302_0,
    o_8_457_0_0  );
  input  i_8_457_19_0, i_8_457_46_0, i_8_457_67_0, i_8_457_70_0,
    i_8_457_88_0, i_8_457_136_0, i_8_457_232_0, i_8_457_252_0,
    i_8_457_255_0, i_8_457_343_0, i_8_457_350_0, i_8_457_378_0,
    i_8_457_379_0, i_8_457_429_0, i_8_457_430_0, i_8_457_450_0,
    i_8_457_454_0, i_8_457_484_0, i_8_457_496_0, i_8_457_507_0,
    i_8_457_556_0, i_8_457_585_0, i_8_457_586_0, i_8_457_610_0,
    i_8_457_634_0, i_8_457_655_0, i_8_457_699_0, i_8_457_702_0,
    i_8_457_703_0, i_8_457_708_0, i_8_457_709_0, i_8_457_718_0,
    i_8_457_733_0, i_8_457_814_0, i_8_457_841_0, i_8_457_879_0,
    i_8_457_880_0, i_8_457_889_0, i_8_457_978_0, i_8_457_979_0,
    i_8_457_996_0, i_8_457_1032_0, i_8_457_1078_0, i_8_457_1140_0,
    i_8_457_1141_0, i_8_457_1144_0, i_8_457_1149_0, i_8_457_1150_0,
    i_8_457_1168_0, i_8_457_1171_0, i_8_457_1227_0, i_8_457_1239_0,
    i_8_457_1240_0, i_8_457_1251_0, i_8_457_1264_0, i_8_457_1273_0,
    i_8_457_1275_0, i_8_457_1278_0, i_8_457_1356_0, i_8_457_1357_0,
    i_8_457_1359_0, i_8_457_1410_0, i_8_457_1412_0, i_8_457_1547_0,
    i_8_457_1602_0, i_8_457_1603_0, i_8_457_1604_0, i_8_457_1632_0,
    i_8_457_1637_0, i_8_457_1779_0, i_8_457_1803_0, i_8_457_1819_0,
    i_8_457_1824_0, i_8_457_1869_0, i_8_457_1986_0, i_8_457_1996_0,
    i_8_457_2058_0, i_8_457_2059_0, i_8_457_2107_0, i_8_457_2146_0,
    i_8_457_2148_0, i_8_457_2149_0, i_8_457_2150_0, i_8_457_2152_0,
    i_8_457_2157_0, i_8_457_2175_0, i_8_457_2176_0, i_8_457_2233_0,
    i_8_457_2238_0, i_8_457_2241_0, i_8_457_2242_0, i_8_457_2243_0,
    i_8_457_2244_0, i_8_457_2248_0, i_8_457_2260_0, i_8_457_2263_0,
    i_8_457_2272_0, i_8_457_2273_0, i_8_457_2301_0, i_8_457_2302_0;
  output o_8_457_0_0;
  assign o_8_457_0_0 = ~((i_8_457_88_0 & ((~i_8_457_19_0 & ~i_8_457_136_0 & i_8_457_484_0) | (~i_8_457_350_0 & ~i_8_457_496_0 & ~i_8_457_709_0 & ~i_8_457_1150_0 & ~i_8_457_2272_0))) | (~i_8_457_379_0 & ((i_8_457_70_0 & ~i_8_457_232_0 & ~i_8_457_343_0 & ~i_8_457_978_0 & ~i_8_457_1251_0 & ~i_8_457_1603_0 & ~i_8_457_1604_0 & ~i_8_457_2263_0) | (~i_8_457_378_0 & ~i_8_457_430_0 & ~i_8_457_879_0 & ~i_8_457_1141_0 & ~i_8_457_1168_0 & ~i_8_457_2238_0 & ~i_8_457_2272_0 & ~i_8_457_2273_0))) | (~i_8_457_46_0 & ((~i_8_457_1140_0 & ((~i_8_457_430_0 & ((~i_8_457_585_0 & ~i_8_457_634_0 & ~i_8_457_655_0 & ~i_8_457_1278_0 & ~i_8_457_2059_0 & ~i_8_457_2152_0 & ~i_8_457_2238_0 & ~i_8_457_2241_0 & ~i_8_457_2243_0 & ~i_8_457_2248_0 & i_8_457_2272_0) | (i_8_457_343_0 & ~i_8_457_378_0 & ~i_8_457_1150_0 & ~i_8_457_1273_0 & ~i_8_457_2058_0 & ~i_8_457_2260_0 & ~i_8_457_2273_0 & ~i_8_457_2302_0))) | (~i_8_457_484_0 & ~i_8_457_496_0 & ~i_8_457_585_0 & i_8_457_841_0 & ~i_8_457_889_0 & ~i_8_457_1547_0 & ~i_8_457_1604_0 & i_8_457_2152_0))) | (~i_8_457_1149_0 & ~i_8_457_1251_0 & ((~i_8_457_232_0 & ~i_8_457_1078_0 & i_8_457_1264_0 & ~i_8_457_1637_0 & i_8_457_2243_0) | (~i_8_457_350_0 & ~i_8_457_718_0 & i_8_457_2146_0 & ~i_8_457_2157_0 & i_8_457_2233_0 & i_8_457_2273_0))) | (~i_8_457_429_0 & i_8_457_430_0 & ~i_8_457_496_0 & ~i_8_457_879_0 & ~i_8_457_889_0 & ~i_8_457_1141_0 & ~i_8_457_1603_0) | (~i_8_457_484_0 & ~i_8_457_996_0 & ~i_8_457_1168_0 & i_8_457_1227_0 & i_8_457_1803_0 & ~i_8_457_1986_0) | (~i_8_457_19_0 & ~i_8_457_880_0 & ~i_8_457_2238_0 & i_8_457_2260_0))) | (~i_8_457_1144_0 & ((~i_8_457_350_0 & ~i_8_457_718_0 & ((~i_8_457_655_0 & ~i_8_457_709_0 & ~i_8_457_1140_0 & ~i_8_457_1603_0 & ~i_8_457_2107_0 & ~i_8_457_2157_0) | (~i_8_457_70_0 & ~i_8_457_343_0 & ~i_8_457_378_0 & ~i_8_457_1168_0 & ~i_8_457_1547_0 & ~i_8_457_1602_0 & ~i_8_457_1604_0 & ~i_8_457_1637_0 & ~i_8_457_1869_0 & ~i_8_457_2149_0 & ~i_8_457_2150_0 & ~i_8_457_2175_0 & ~i_8_457_2238_0))) | (~i_8_457_429_0 & ((~i_8_457_19_0 & ((~i_8_457_586_0 & ~i_8_457_610_0 & ~i_8_457_889_0 & ~i_8_457_1150_0 & ~i_8_457_2175_0) | (~i_8_457_343_0 & ~i_8_457_430_0 & ~i_8_457_709_0 & ~i_8_457_1278_0 & ~i_8_457_1603_0 & ~i_8_457_2176_0 & ~i_8_457_2260_0))) | (~i_8_457_232_0 & ~i_8_457_343_0 & ~i_8_457_450_0 & ~i_8_457_996_0 & ~i_8_457_1547_0 & ~i_8_457_1604_0 & ~i_8_457_2107_0 & ~i_8_457_2176_0 & ~i_8_457_2238_0))) | (~i_8_457_19_0 & ~i_8_457_879_0 & ~i_8_457_1168_0 & ~i_8_457_2107_0 & i_8_457_2148_0 & ~i_8_457_2152_0 & ~i_8_457_2248_0) | (~i_8_457_1032_0 & ~i_8_457_1149_0 & ~i_8_457_1603_0 & i_8_457_2157_0 & i_8_457_2272_0))) | (i_8_457_2149_0 & ((~i_8_457_450_0 & ((~i_8_457_232_0 & ~i_8_457_343_0 & ~i_8_457_1171_0 & ~i_8_457_1986_0 & ~i_8_457_2059_0 & ~i_8_457_2157_0) | (~i_8_457_996_0 & ~i_8_457_1140_0 & ~i_8_457_1547_0 & i_8_457_2058_0 & i_8_457_2176_0))) | (~i_8_457_610_0 & ~i_8_457_1032_0 & ~i_8_457_1168_0 & ~i_8_457_1410_0 & ~i_8_457_1603_0 & ~i_8_457_2175_0))) | (i_8_457_586_0 & ((~i_8_457_1140_0 & i_8_457_1264_0 & ~i_8_457_2152_0 & ~i_8_457_2233_0 & ~i_8_457_2243_0) | (~i_8_457_496_0 & ~i_8_457_708_0 & ~i_8_457_1168_0 & i_8_457_1278_0 & ~i_8_457_2149_0 & ~i_8_457_2238_0 & ~i_8_457_2301_0))) | (~i_8_457_1150_0 & ((~i_8_457_496_0 & ((~i_8_457_88_0 & i_8_457_702_0 & i_8_457_703_0 & ~i_8_457_841_0 & ~i_8_457_978_0 & ~i_8_457_1140_0 & ~i_8_457_1171_0) | (~i_8_457_343_0 & ~i_8_457_880_0 & ~i_8_457_1141_0 & ~i_8_457_1149_0 & ~i_8_457_1168_0 & ~i_8_457_1251_0 & ~i_8_457_2058_0 & ~i_8_457_2107_0))) | (~i_8_457_1140_0 & ((i_8_457_484_0 & ~i_8_457_610_0 & ~i_8_457_841_0 & ~i_8_457_1603_0) | (~i_8_457_586_0 & ~i_8_457_879_0 & ~i_8_457_1141_0 & ~i_8_457_1171_0 & ~i_8_457_2152_0 & ~i_8_457_2175_0 & ~i_8_457_2176_0 & ~i_8_457_2273_0))))) | (~i_8_457_343_0 & ((~i_8_457_1032_0 & ~i_8_457_1168_0 & i_8_457_1239_0 & ~i_8_457_1604_0 & ~i_8_457_2058_0) | (~i_8_457_19_0 & ~i_8_457_586_0 & ~i_8_457_1240_0 & i_8_457_1278_0 & ~i_8_457_1603_0 & ~i_8_457_1632_0 & ~i_8_457_1819_0 & ~i_8_457_2148_0 & ~i_8_457_2273_0))) | (~i_8_457_19_0 & ~i_8_457_1227_0 & ((~i_8_457_136_0 & ~i_8_457_1171_0 & ~i_8_457_1278_0 & ~i_8_457_1602_0 & ~i_8_457_2059_0 & ~i_8_457_2157_0 & i_8_457_2233_0) | (~i_8_457_889_0 & i_8_457_1078_0 & ~i_8_457_1604_0 & ~i_8_457_1824_0 & ~i_8_457_2301_0))) | (~i_8_457_586_0 & ~i_8_457_1602_0 & ((i_8_457_699_0 & i_8_457_1227_0 & i_8_457_2146_0) | (~i_8_457_232_0 & ~i_8_457_1251_0 & ~i_8_457_1603_0 & ~i_8_457_1803_0 & i_8_457_1986_0 & ~i_8_457_2059_0 & ~i_8_457_2176_0 & ~i_8_457_2238_0 & ~i_8_457_2263_0))) | (~i_8_457_232_0 & ~i_8_457_1171_0 & ((i_8_457_136_0 & ~i_8_457_255_0 & ~i_8_457_1251_0 & ~i_8_457_1547_0 & ~i_8_457_1603_0 & ~i_8_457_2058_0 & ~i_8_457_2059_0) | (~i_8_457_610_0 & ~i_8_457_709_0 & i_8_457_841_0 & ~i_8_457_889_0 & ~i_8_457_978_0 & ~i_8_457_1869_0 & ~i_8_457_2107_0 & ~i_8_457_2175_0 & ~i_8_457_2238_0 & ~i_8_457_2260_0))) | (~i_8_457_1140_0 & ~i_8_457_2107_0 & ~i_8_457_2176_0 & ((~i_8_457_378_0 & ~i_8_457_1356_0 & ~i_8_457_1412_0 & i_8_457_1547_0 & ~i_8_457_2148_0) | (~i_8_457_879_0 & ~i_8_457_1141_0 & ~i_8_457_1168_0 & ~i_8_457_1603_0 & ~i_8_457_1604_0 & ~i_8_457_1986_0 & ~i_8_457_2152_0 & ~i_8_457_2238_0))) | (~i_8_457_1547_0 & ((i_8_457_19_0 & i_8_457_634_0 & i_8_457_703_0 & ~i_8_457_1141_0 & ~i_8_457_1149_0) | (i_8_457_1275_0 & i_8_457_1410_0))) | (~i_8_457_1141_0 & ~i_8_457_2260_0 & ((i_8_457_1264_0 & ~i_8_457_1803_0 & i_8_457_2058_0) | (i_8_457_507_0 & ~i_8_457_634_0 & ~i_8_457_699_0 & ~i_8_457_1149_0 & ~i_8_457_1410_0 & ~i_8_457_2273_0))) | (i_8_457_1078_0 & i_8_457_1637_0) | (i_8_457_841_0 & i_8_457_889_0 & ~i_8_457_1149_0 & ~i_8_457_1168_0 & ~i_8_457_1412_0 & ~i_8_457_1604_0 & ~i_8_457_2058_0 & ~i_8_457_2157_0));
endmodule



// Benchmark "kernel_8_458" written by ABC on Sun Jul 19 10:11:09 2020

module kernel_8_458 ( 
    i_8_458_87_0, i_8_458_88_0, i_8_458_93_0, i_8_458_157_0, i_8_458_187_0,
    i_8_458_192_0, i_8_458_206_0, i_8_458_221_0, i_8_458_255_0,
    i_8_458_259_0, i_8_458_263_0, i_8_458_275_0, i_8_458_295_0,
    i_8_458_304_0, i_8_458_322_0, i_8_458_363_0, i_8_458_367_0,
    i_8_458_392_0, i_8_458_414_0, i_8_458_415_0, i_8_458_445_0,
    i_8_458_456_0, i_8_458_464_0, i_8_458_466_0, i_8_458_483_0,
    i_8_458_525_0, i_8_458_528_0, i_8_458_556_0, i_8_458_602_0,
    i_8_458_606_0, i_8_458_625_0, i_8_458_627_0, i_8_458_652_0,
    i_8_458_663_0, i_8_458_673_0, i_8_458_718_0, i_8_458_769_0,
    i_8_458_795_0, i_8_458_798_0, i_8_458_799_0, i_8_458_840_0,
    i_8_458_854_0, i_8_458_855_0, i_8_458_876_0, i_8_458_879_0,
    i_8_458_881_0, i_8_458_895_0, i_8_458_990_0, i_8_458_993_0,
    i_8_458_1033_0, i_8_458_1113_0, i_8_458_1114_0, i_8_458_1159_0,
    i_8_458_1216_0, i_8_458_1218_0, i_8_458_1263_0, i_8_458_1322_0,
    i_8_458_1325_0, i_8_458_1331_0, i_8_458_1349_0, i_8_458_1438_0,
    i_8_458_1443_0, i_8_458_1444_0, i_8_458_1447_0, i_8_458_1524_0,
    i_8_458_1528_0, i_8_458_1543_0, i_8_458_1555_0, i_8_458_1571_0,
    i_8_458_1587_0, i_8_458_1590_0, i_8_458_1600_0, i_8_458_1617_0,
    i_8_458_1648_0, i_8_458_1736_0, i_8_458_1744_0, i_8_458_1786_0,
    i_8_458_1807_0, i_8_458_1843_0, i_8_458_1844_0, i_8_458_1930_0,
    i_8_458_1951_0, i_8_458_1989_0, i_8_458_2025_0, i_8_458_2028_0,
    i_8_458_2050_0, i_8_458_2109_0, i_8_458_2110_0, i_8_458_2131_0,
    i_8_458_2184_0, i_8_458_2185_0, i_8_458_2186_0, i_8_458_2193_0,
    i_8_458_2214_0, i_8_458_2215_0, i_8_458_2217_0, i_8_458_2224_0,
    i_8_458_2235_0, i_8_458_2239_0, i_8_458_2293_0,
    o_8_458_0_0  );
  input  i_8_458_87_0, i_8_458_88_0, i_8_458_93_0, i_8_458_157_0,
    i_8_458_187_0, i_8_458_192_0, i_8_458_206_0, i_8_458_221_0,
    i_8_458_255_0, i_8_458_259_0, i_8_458_263_0, i_8_458_275_0,
    i_8_458_295_0, i_8_458_304_0, i_8_458_322_0, i_8_458_363_0,
    i_8_458_367_0, i_8_458_392_0, i_8_458_414_0, i_8_458_415_0,
    i_8_458_445_0, i_8_458_456_0, i_8_458_464_0, i_8_458_466_0,
    i_8_458_483_0, i_8_458_525_0, i_8_458_528_0, i_8_458_556_0,
    i_8_458_602_0, i_8_458_606_0, i_8_458_625_0, i_8_458_627_0,
    i_8_458_652_0, i_8_458_663_0, i_8_458_673_0, i_8_458_718_0,
    i_8_458_769_0, i_8_458_795_0, i_8_458_798_0, i_8_458_799_0,
    i_8_458_840_0, i_8_458_854_0, i_8_458_855_0, i_8_458_876_0,
    i_8_458_879_0, i_8_458_881_0, i_8_458_895_0, i_8_458_990_0,
    i_8_458_993_0, i_8_458_1033_0, i_8_458_1113_0, i_8_458_1114_0,
    i_8_458_1159_0, i_8_458_1216_0, i_8_458_1218_0, i_8_458_1263_0,
    i_8_458_1322_0, i_8_458_1325_0, i_8_458_1331_0, i_8_458_1349_0,
    i_8_458_1438_0, i_8_458_1443_0, i_8_458_1444_0, i_8_458_1447_0,
    i_8_458_1524_0, i_8_458_1528_0, i_8_458_1543_0, i_8_458_1555_0,
    i_8_458_1571_0, i_8_458_1587_0, i_8_458_1590_0, i_8_458_1600_0,
    i_8_458_1617_0, i_8_458_1648_0, i_8_458_1736_0, i_8_458_1744_0,
    i_8_458_1786_0, i_8_458_1807_0, i_8_458_1843_0, i_8_458_1844_0,
    i_8_458_1930_0, i_8_458_1951_0, i_8_458_1989_0, i_8_458_2025_0,
    i_8_458_2028_0, i_8_458_2050_0, i_8_458_2109_0, i_8_458_2110_0,
    i_8_458_2131_0, i_8_458_2184_0, i_8_458_2185_0, i_8_458_2186_0,
    i_8_458_2193_0, i_8_458_2214_0, i_8_458_2215_0, i_8_458_2217_0,
    i_8_458_2224_0, i_8_458_2235_0, i_8_458_2239_0, i_8_458_2293_0;
  output o_8_458_0_0;
  assign o_8_458_0_0 = 0;
endmodule



// Benchmark "kernel_8_459" written by ABC on Sun Jul 19 10:11:10 2020

module kernel_8_459 ( 
    i_8_459_86_0, i_8_459_148_0, i_8_459_157_0, i_8_459_201_0,
    i_8_459_203_0, i_8_459_207_0, i_8_459_221_0, i_8_459_231_0,
    i_8_459_232_0, i_8_459_298_0, i_8_459_300_0, i_8_459_340_0,
    i_8_459_342_0, i_8_459_350_0, i_8_459_370_0, i_8_459_388_0,
    i_8_459_454_0, i_8_459_473_0, i_8_459_479_0, i_8_459_484_0,
    i_8_459_485_0, i_8_459_498_0, i_8_459_525_0, i_8_459_543_0,
    i_8_459_552_0, i_8_459_574_0, i_8_459_625_0, i_8_459_659_0,
    i_8_459_663_0, i_8_459_666_0, i_8_459_667_0, i_8_459_678_0,
    i_8_459_704_0, i_8_459_708_0, i_8_459_762_0, i_8_459_768_0,
    i_8_459_778_0, i_8_459_779_0, i_8_459_829_0, i_8_459_867_0,
    i_8_459_949_0, i_8_459_984_0, i_8_459_991_0, i_8_459_1003_0,
    i_8_459_1013_0, i_8_459_1030_0, i_8_459_1031_0, i_8_459_1090_0,
    i_8_459_1104_0, i_8_459_1106_0, i_8_459_1108_0, i_8_459_1117_0,
    i_8_459_1129_0, i_8_459_1204_0, i_8_459_1217_0, i_8_459_1219_0,
    i_8_459_1220_0, i_8_459_1327_0, i_8_459_1345_0, i_8_459_1346_0,
    i_8_459_1358_0, i_8_459_1402_0, i_8_459_1417_0, i_8_459_1443_0,
    i_8_459_1514_0, i_8_459_1544_0, i_8_459_1563_0, i_8_459_1564_0,
    i_8_459_1578_0, i_8_459_1594_0, i_8_459_1597_0, i_8_459_1611_0,
    i_8_459_1613_0, i_8_459_1630_0, i_8_459_1669_0, i_8_459_1677_0,
    i_8_459_1707_0, i_8_459_1710_0, i_8_459_1713_0, i_8_459_1722_0,
    i_8_459_1735_0, i_8_459_1774_0, i_8_459_1798_0, i_8_459_1802_0,
    i_8_459_1826_0, i_8_459_1867_0, i_8_459_1872_0, i_8_459_1899_0,
    i_8_459_2047_0, i_8_459_2048_0, i_8_459_2049_0, i_8_459_2055_0,
    i_8_459_2070_0, i_8_459_2074_0, i_8_459_2088_0, i_8_459_2106_0,
    i_8_459_2227_0, i_8_459_2260_0, i_8_459_2286_0, i_8_459_2299_0,
    o_8_459_0_0  );
  input  i_8_459_86_0, i_8_459_148_0, i_8_459_157_0, i_8_459_201_0,
    i_8_459_203_0, i_8_459_207_0, i_8_459_221_0, i_8_459_231_0,
    i_8_459_232_0, i_8_459_298_0, i_8_459_300_0, i_8_459_340_0,
    i_8_459_342_0, i_8_459_350_0, i_8_459_370_0, i_8_459_388_0,
    i_8_459_454_0, i_8_459_473_0, i_8_459_479_0, i_8_459_484_0,
    i_8_459_485_0, i_8_459_498_0, i_8_459_525_0, i_8_459_543_0,
    i_8_459_552_0, i_8_459_574_0, i_8_459_625_0, i_8_459_659_0,
    i_8_459_663_0, i_8_459_666_0, i_8_459_667_0, i_8_459_678_0,
    i_8_459_704_0, i_8_459_708_0, i_8_459_762_0, i_8_459_768_0,
    i_8_459_778_0, i_8_459_779_0, i_8_459_829_0, i_8_459_867_0,
    i_8_459_949_0, i_8_459_984_0, i_8_459_991_0, i_8_459_1003_0,
    i_8_459_1013_0, i_8_459_1030_0, i_8_459_1031_0, i_8_459_1090_0,
    i_8_459_1104_0, i_8_459_1106_0, i_8_459_1108_0, i_8_459_1117_0,
    i_8_459_1129_0, i_8_459_1204_0, i_8_459_1217_0, i_8_459_1219_0,
    i_8_459_1220_0, i_8_459_1327_0, i_8_459_1345_0, i_8_459_1346_0,
    i_8_459_1358_0, i_8_459_1402_0, i_8_459_1417_0, i_8_459_1443_0,
    i_8_459_1514_0, i_8_459_1544_0, i_8_459_1563_0, i_8_459_1564_0,
    i_8_459_1578_0, i_8_459_1594_0, i_8_459_1597_0, i_8_459_1611_0,
    i_8_459_1613_0, i_8_459_1630_0, i_8_459_1669_0, i_8_459_1677_0,
    i_8_459_1707_0, i_8_459_1710_0, i_8_459_1713_0, i_8_459_1722_0,
    i_8_459_1735_0, i_8_459_1774_0, i_8_459_1798_0, i_8_459_1802_0,
    i_8_459_1826_0, i_8_459_1867_0, i_8_459_1872_0, i_8_459_1899_0,
    i_8_459_2047_0, i_8_459_2048_0, i_8_459_2049_0, i_8_459_2055_0,
    i_8_459_2070_0, i_8_459_2074_0, i_8_459_2088_0, i_8_459_2106_0,
    i_8_459_2227_0, i_8_459_2260_0, i_8_459_2286_0, i_8_459_2299_0;
  output o_8_459_0_0;
  assign o_8_459_0_0 = 0;
endmodule



// Benchmark "kernel_8_460" written by ABC on Sun Jul 19 10:11:11 2020

module kernel_8_460 ( 
    i_8_460_23_0, i_8_460_41_0, i_8_460_73_0, i_8_460_106_0, i_8_460_187_0,
    i_8_460_189_0, i_8_460_193_0, i_8_460_217_0, i_8_460_243_0,
    i_8_460_364_0, i_8_460_390_0, i_8_460_411_0, i_8_460_423_0,
    i_8_460_424_0, i_8_460_425_0, i_8_460_426_0, i_8_460_454_0,
    i_8_460_468_0, i_8_460_472_0, i_8_460_490_0, i_8_460_572_0,
    i_8_460_583_0, i_8_460_610_0, i_8_460_652_0, i_8_460_665_0,
    i_8_460_676_0, i_8_460_679_0, i_8_460_705_0, i_8_460_738_0,
    i_8_460_752_0, i_8_460_775_0, i_8_460_808_0, i_8_460_837_0,
    i_8_460_856_0, i_8_460_867_0, i_8_460_876_0, i_8_460_882_0,
    i_8_460_883_0, i_8_460_931_0, i_8_460_984_0, i_8_460_994_0,
    i_8_460_1039_0, i_8_460_1040_0, i_8_460_1048_0, i_8_460_1057_0,
    i_8_460_1123_0, i_8_460_1126_0, i_8_460_1138_0, i_8_460_1162_0,
    i_8_460_1174_0, i_8_460_1200_0, i_8_460_1223_0, i_8_460_1226_0,
    i_8_460_1239_0, i_8_460_1242_0, i_8_460_1245_0, i_8_460_1286_0,
    i_8_460_1294_0, i_8_460_1311_0, i_8_460_1348_0, i_8_460_1362_0,
    i_8_460_1363_0, i_8_460_1396_0, i_8_460_1431_0, i_8_460_1456_0,
    i_8_460_1539_0, i_8_460_1546_0, i_8_460_1547_0, i_8_460_1563_0,
    i_8_460_1564_0, i_8_460_1574_0, i_8_460_1601_0, i_8_460_1624_0,
    i_8_460_1639_0, i_8_460_1642_0, i_8_460_1655_0, i_8_460_1659_0,
    i_8_460_1679_0, i_8_460_1702_0, i_8_460_1713_0, i_8_460_1746_0,
    i_8_460_1783_0, i_8_460_1802_0, i_8_460_1861_0, i_8_460_1885_0,
    i_8_460_1920_0, i_8_460_1974_0, i_8_460_1981_0, i_8_460_1984_0,
    i_8_460_1992_0, i_8_460_2031_0, i_8_460_2083_0, i_8_460_2091_0,
    i_8_460_2137_0, i_8_460_2155_0, i_8_460_2164_0, i_8_460_2246_0,
    i_8_460_2247_0, i_8_460_2272_0, i_8_460_2275_0,
    o_8_460_0_0  );
  input  i_8_460_23_0, i_8_460_41_0, i_8_460_73_0, i_8_460_106_0,
    i_8_460_187_0, i_8_460_189_0, i_8_460_193_0, i_8_460_217_0,
    i_8_460_243_0, i_8_460_364_0, i_8_460_390_0, i_8_460_411_0,
    i_8_460_423_0, i_8_460_424_0, i_8_460_425_0, i_8_460_426_0,
    i_8_460_454_0, i_8_460_468_0, i_8_460_472_0, i_8_460_490_0,
    i_8_460_572_0, i_8_460_583_0, i_8_460_610_0, i_8_460_652_0,
    i_8_460_665_0, i_8_460_676_0, i_8_460_679_0, i_8_460_705_0,
    i_8_460_738_0, i_8_460_752_0, i_8_460_775_0, i_8_460_808_0,
    i_8_460_837_0, i_8_460_856_0, i_8_460_867_0, i_8_460_876_0,
    i_8_460_882_0, i_8_460_883_0, i_8_460_931_0, i_8_460_984_0,
    i_8_460_994_0, i_8_460_1039_0, i_8_460_1040_0, i_8_460_1048_0,
    i_8_460_1057_0, i_8_460_1123_0, i_8_460_1126_0, i_8_460_1138_0,
    i_8_460_1162_0, i_8_460_1174_0, i_8_460_1200_0, i_8_460_1223_0,
    i_8_460_1226_0, i_8_460_1239_0, i_8_460_1242_0, i_8_460_1245_0,
    i_8_460_1286_0, i_8_460_1294_0, i_8_460_1311_0, i_8_460_1348_0,
    i_8_460_1362_0, i_8_460_1363_0, i_8_460_1396_0, i_8_460_1431_0,
    i_8_460_1456_0, i_8_460_1539_0, i_8_460_1546_0, i_8_460_1547_0,
    i_8_460_1563_0, i_8_460_1564_0, i_8_460_1574_0, i_8_460_1601_0,
    i_8_460_1624_0, i_8_460_1639_0, i_8_460_1642_0, i_8_460_1655_0,
    i_8_460_1659_0, i_8_460_1679_0, i_8_460_1702_0, i_8_460_1713_0,
    i_8_460_1746_0, i_8_460_1783_0, i_8_460_1802_0, i_8_460_1861_0,
    i_8_460_1885_0, i_8_460_1920_0, i_8_460_1974_0, i_8_460_1981_0,
    i_8_460_1984_0, i_8_460_1992_0, i_8_460_2031_0, i_8_460_2083_0,
    i_8_460_2091_0, i_8_460_2137_0, i_8_460_2155_0, i_8_460_2164_0,
    i_8_460_2246_0, i_8_460_2247_0, i_8_460_2272_0, i_8_460_2275_0;
  output o_8_460_0_0;
  assign o_8_460_0_0 = 0;
endmodule



// Benchmark "kernel_8_461" written by ABC on Sun Jul 19 10:11:12 2020

module kernel_8_461 ( 
    i_8_461_30_0, i_8_461_143_0, i_8_461_214_0, i_8_461_215_0,
    i_8_461_219_0, i_8_461_259_0, i_8_461_268_0, i_8_461_347_0,
    i_8_461_350_0, i_8_461_377_0, i_8_461_378_0, i_8_461_383_0,
    i_8_461_385_0, i_8_461_430_0, i_8_461_456_0, i_8_461_468_0,
    i_8_461_469_0, i_8_461_556_0, i_8_461_557_0, i_8_461_606_0,
    i_8_461_615_0, i_8_461_618_0, i_8_461_627_0, i_8_461_646_0,
    i_8_461_663_0, i_8_461_772_0, i_8_461_780_0, i_8_461_796_0,
    i_8_461_871_0, i_8_461_881_0, i_8_461_898_0, i_8_461_899_0,
    i_8_461_921_0, i_8_461_952_0, i_8_461_953_0, i_8_461_975_0,
    i_8_461_978_0, i_8_461_979_0, i_8_461_1015_0, i_8_461_1027_0,
    i_8_461_1045_0, i_8_461_1051_0, i_8_461_1057_0, i_8_461_1140_0,
    i_8_461_1159_0, i_8_461_1185_0, i_8_461_1194_0, i_8_461_1204_0,
    i_8_461_1237_0, i_8_461_1239_0, i_8_461_1272_0, i_8_461_1282_0,
    i_8_461_1285_0, i_8_461_1286_0, i_8_461_1339_0, i_8_461_1429_0,
    i_8_461_1435_0, i_8_461_1438_0, i_8_461_1446_0, i_8_461_1447_0,
    i_8_461_1474_0, i_8_461_1506_0, i_8_461_1507_0, i_8_461_1527_0,
    i_8_461_1528_0, i_8_461_1529_0, i_8_461_1534_0, i_8_461_1538_0,
    i_8_461_1545_0, i_8_461_1555_0, i_8_461_1635_0, i_8_461_1645_0,
    i_8_461_1652_0, i_8_461_1671_0, i_8_461_1672_0, i_8_461_1735_0,
    i_8_461_1753_0, i_8_461_1779_0, i_8_461_1786_0, i_8_461_1798_0,
    i_8_461_1807_0, i_8_461_1840_0, i_8_461_1860_0, i_8_461_1867_0,
    i_8_461_1941_0, i_8_461_1942_0, i_8_461_1969_0, i_8_461_1987_0,
    i_8_461_2002_0, i_8_461_2004_0, i_8_461_2014_0, i_8_461_2113_0,
    i_8_461_2139_0, i_8_461_2151_0, i_8_461_2158_0, i_8_461_2219_0,
    i_8_461_2264_0, i_8_461_2267_0, i_8_461_2274_0, i_8_461_2293_0,
    o_8_461_0_0  );
  input  i_8_461_30_0, i_8_461_143_0, i_8_461_214_0, i_8_461_215_0,
    i_8_461_219_0, i_8_461_259_0, i_8_461_268_0, i_8_461_347_0,
    i_8_461_350_0, i_8_461_377_0, i_8_461_378_0, i_8_461_383_0,
    i_8_461_385_0, i_8_461_430_0, i_8_461_456_0, i_8_461_468_0,
    i_8_461_469_0, i_8_461_556_0, i_8_461_557_0, i_8_461_606_0,
    i_8_461_615_0, i_8_461_618_0, i_8_461_627_0, i_8_461_646_0,
    i_8_461_663_0, i_8_461_772_0, i_8_461_780_0, i_8_461_796_0,
    i_8_461_871_0, i_8_461_881_0, i_8_461_898_0, i_8_461_899_0,
    i_8_461_921_0, i_8_461_952_0, i_8_461_953_0, i_8_461_975_0,
    i_8_461_978_0, i_8_461_979_0, i_8_461_1015_0, i_8_461_1027_0,
    i_8_461_1045_0, i_8_461_1051_0, i_8_461_1057_0, i_8_461_1140_0,
    i_8_461_1159_0, i_8_461_1185_0, i_8_461_1194_0, i_8_461_1204_0,
    i_8_461_1237_0, i_8_461_1239_0, i_8_461_1272_0, i_8_461_1282_0,
    i_8_461_1285_0, i_8_461_1286_0, i_8_461_1339_0, i_8_461_1429_0,
    i_8_461_1435_0, i_8_461_1438_0, i_8_461_1446_0, i_8_461_1447_0,
    i_8_461_1474_0, i_8_461_1506_0, i_8_461_1507_0, i_8_461_1527_0,
    i_8_461_1528_0, i_8_461_1529_0, i_8_461_1534_0, i_8_461_1538_0,
    i_8_461_1545_0, i_8_461_1555_0, i_8_461_1635_0, i_8_461_1645_0,
    i_8_461_1652_0, i_8_461_1671_0, i_8_461_1672_0, i_8_461_1735_0,
    i_8_461_1753_0, i_8_461_1779_0, i_8_461_1786_0, i_8_461_1798_0,
    i_8_461_1807_0, i_8_461_1840_0, i_8_461_1860_0, i_8_461_1867_0,
    i_8_461_1941_0, i_8_461_1942_0, i_8_461_1969_0, i_8_461_1987_0,
    i_8_461_2002_0, i_8_461_2004_0, i_8_461_2014_0, i_8_461_2113_0,
    i_8_461_2139_0, i_8_461_2151_0, i_8_461_2158_0, i_8_461_2219_0,
    i_8_461_2264_0, i_8_461_2267_0, i_8_461_2274_0, i_8_461_2293_0;
  output o_8_461_0_0;
  assign o_8_461_0_0 = ~((~i_8_461_627_0 & ((~i_8_461_268_0 & ~i_8_461_898_0 & ~i_8_461_1527_0 & ~i_8_461_1529_0 & ~i_8_461_1941_0 & ~i_8_461_2219_0) | (~i_8_461_606_0 & ~i_8_461_978_0 & ~i_8_461_1435_0 & ~i_8_461_2113_0 & ~i_8_461_2293_0))) | (~i_8_461_268_0 & ((~i_8_461_456_0 & ~i_8_461_1045_0 & i_8_461_1506_0 & i_8_461_1672_0) | (~i_8_461_898_0 & ~i_8_461_921_0 & ~i_8_461_1140_0 & ~i_8_461_1671_0 & i_8_461_2219_0))) | (~i_8_461_646_0 & ((~i_8_461_215_0 & ~i_8_461_556_0 & ~i_8_461_1204_0 & ~i_8_461_1446_0) | (~i_8_461_780_0 & ~i_8_461_1429_0 & ~i_8_461_2139_0 & ~i_8_461_2267_0))) | (~i_8_461_898_0 & i_8_461_1051_0 & ((~i_8_461_618_0 & ~i_8_461_1529_0) | (~i_8_461_378_0 & ~i_8_461_1969_0 & ~i_8_461_2014_0 & ~i_8_461_2267_0))) | (~i_8_461_1051_0 & ~i_8_461_1942_0 & ~i_8_461_2267_0 & ((~i_8_461_468_0 & i_8_461_556_0 & ~i_8_461_1447_0 & ~i_8_461_1528_0 & i_8_461_1779_0) | (~i_8_461_871_0 & ~i_8_461_921_0 & ~i_8_461_1140_0 & i_8_461_1635_0 & i_8_461_1753_0 & ~i_8_461_1860_0 & ~i_8_461_1987_0))) | (~i_8_461_921_0 & ((~i_8_461_979_0 & ~i_8_461_1474_0 & ~i_8_461_1798_0 & ~i_8_461_1941_0 & ~i_8_461_2004_0 & ~i_8_461_2264_0) | (~i_8_461_978_0 & ~i_8_461_1204_0 & ~i_8_461_1429_0 & ~i_8_461_2293_0))) | (~i_8_461_2219_0 & ((~i_8_461_663_0 & ~i_8_461_772_0 & ~i_8_461_1446_0 & ~i_8_461_1527_0) | (~i_8_461_615_0 & ~i_8_461_1672_0 & i_8_461_2158_0))) | (i_8_461_1045_0 & i_8_461_1286_0) | (i_8_461_1474_0 & ~i_8_461_1528_0 & ~i_8_461_1635_0 & ~i_8_461_1798_0));
endmodule



// Benchmark "kernel_8_462" written by ABC on Sun Jul 19 10:11:13 2020

module kernel_8_462 ( 
    i_8_462_21_0, i_8_462_30_0, i_8_462_86_0, i_8_462_87_0, i_8_462_142_0,
    i_8_462_169_0, i_8_462_185_0, i_8_462_187_0, i_8_462_193_0,
    i_8_462_213_0, i_8_462_233_0, i_8_462_255_0, i_8_462_256_0,
    i_8_462_260_0, i_8_462_292_0, i_8_462_295_0, i_8_462_346_0,
    i_8_462_376_0, i_8_462_417_0, i_8_462_418_0, i_8_462_445_0,
    i_8_462_453_0, i_8_462_456_0, i_8_462_464_0, i_8_462_481_0,
    i_8_462_485_0, i_8_462_503_0, i_8_462_510_0, i_8_462_522_0,
    i_8_462_525_0, i_8_462_526_0, i_8_462_530_0, i_8_462_556_0,
    i_8_462_592_0, i_8_462_601_0, i_8_462_704_0, i_8_462_705_0,
    i_8_462_717_0, i_8_462_761_0, i_8_462_763_0, i_8_462_764_0,
    i_8_462_789_0, i_8_462_798_0, i_8_462_894_0, i_8_462_952_0,
    i_8_462_993_0, i_8_462_996_0, i_8_462_998_0, i_8_462_1050_0,
    i_8_462_1074_0, i_8_462_1078_0, i_8_462_1121_0, i_8_462_1123_0,
    i_8_462_1124_0, i_8_462_1159_0, i_8_462_1191_0, i_8_462_1305_0,
    i_8_462_1306_0, i_8_462_1307_0, i_8_462_1308_0, i_8_462_1310_0,
    i_8_462_1328_0, i_8_462_1411_0, i_8_462_1419_0, i_8_462_1444_0,
    i_8_462_1447_0, i_8_462_1471_0, i_8_462_1510_0, i_8_462_1543_0,
    i_8_462_1544_0, i_8_462_1545_0, i_8_462_1578_0, i_8_462_1633_0,
    i_8_462_1642_0, i_8_462_1707_0, i_8_462_1723_0, i_8_462_1730_0,
    i_8_462_1733_0, i_8_462_1741_0, i_8_462_1752_0, i_8_462_1779_0,
    i_8_462_1790_0, i_8_462_1805_0, i_8_462_1812_0, i_8_462_1813_0,
    i_8_462_1889_0, i_8_462_1906_0, i_8_462_1960_0, i_8_462_1993_0,
    i_8_462_2049_0, i_8_462_2104_0, i_8_462_2144_0, i_8_462_2218_0,
    i_8_462_2222_0, i_8_462_2236_0, i_8_462_2247_0, i_8_462_2263_0,
    i_8_462_2275_0, i_8_462_2292_0, i_8_462_2294_0,
    o_8_462_0_0  );
  input  i_8_462_21_0, i_8_462_30_0, i_8_462_86_0, i_8_462_87_0,
    i_8_462_142_0, i_8_462_169_0, i_8_462_185_0, i_8_462_187_0,
    i_8_462_193_0, i_8_462_213_0, i_8_462_233_0, i_8_462_255_0,
    i_8_462_256_0, i_8_462_260_0, i_8_462_292_0, i_8_462_295_0,
    i_8_462_346_0, i_8_462_376_0, i_8_462_417_0, i_8_462_418_0,
    i_8_462_445_0, i_8_462_453_0, i_8_462_456_0, i_8_462_464_0,
    i_8_462_481_0, i_8_462_485_0, i_8_462_503_0, i_8_462_510_0,
    i_8_462_522_0, i_8_462_525_0, i_8_462_526_0, i_8_462_530_0,
    i_8_462_556_0, i_8_462_592_0, i_8_462_601_0, i_8_462_704_0,
    i_8_462_705_0, i_8_462_717_0, i_8_462_761_0, i_8_462_763_0,
    i_8_462_764_0, i_8_462_789_0, i_8_462_798_0, i_8_462_894_0,
    i_8_462_952_0, i_8_462_993_0, i_8_462_996_0, i_8_462_998_0,
    i_8_462_1050_0, i_8_462_1074_0, i_8_462_1078_0, i_8_462_1121_0,
    i_8_462_1123_0, i_8_462_1124_0, i_8_462_1159_0, i_8_462_1191_0,
    i_8_462_1305_0, i_8_462_1306_0, i_8_462_1307_0, i_8_462_1308_0,
    i_8_462_1310_0, i_8_462_1328_0, i_8_462_1411_0, i_8_462_1419_0,
    i_8_462_1444_0, i_8_462_1447_0, i_8_462_1471_0, i_8_462_1510_0,
    i_8_462_1543_0, i_8_462_1544_0, i_8_462_1545_0, i_8_462_1578_0,
    i_8_462_1633_0, i_8_462_1642_0, i_8_462_1707_0, i_8_462_1723_0,
    i_8_462_1730_0, i_8_462_1733_0, i_8_462_1741_0, i_8_462_1752_0,
    i_8_462_1779_0, i_8_462_1790_0, i_8_462_1805_0, i_8_462_1812_0,
    i_8_462_1813_0, i_8_462_1889_0, i_8_462_1906_0, i_8_462_1960_0,
    i_8_462_1993_0, i_8_462_2049_0, i_8_462_2104_0, i_8_462_2144_0,
    i_8_462_2218_0, i_8_462_2222_0, i_8_462_2236_0, i_8_462_2247_0,
    i_8_462_2263_0, i_8_462_2275_0, i_8_462_2292_0, i_8_462_2294_0;
  output o_8_462_0_0;
  assign o_8_462_0_0 = 0;
endmodule



// Benchmark "kernel_8_463" written by ABC on Sun Jul 19 10:11:14 2020

module kernel_8_463 ( 
    i_8_463_3_0, i_8_463_48_0, i_8_463_53_0, i_8_463_106_0, i_8_463_120_0,
    i_8_463_156_0, i_8_463_197_0, i_8_463_258_0, i_8_463_265_0,
    i_8_463_282_0, i_8_463_285_0, i_8_463_376_0, i_8_463_397_0,
    i_8_463_409_0, i_8_463_412_0, i_8_463_439_0, i_8_463_454_0,
    i_8_463_456_0, i_8_463_488_0, i_8_463_490_0, i_8_463_534_0,
    i_8_463_546_0, i_8_463_588_0, i_8_463_591_0, i_8_463_621_0,
    i_8_463_624_0, i_8_463_625_0, i_8_463_628_0, i_8_463_654_0,
    i_8_463_658_0, i_8_463_661_0, i_8_463_663_0, i_8_463_664_0,
    i_8_463_673_0, i_8_463_675_0, i_8_463_682_0, i_8_463_693_0,
    i_8_463_703_0, i_8_463_732_0, i_8_463_735_0, i_8_463_742_0,
    i_8_463_780_0, i_8_463_835_0, i_8_463_841_0, i_8_463_879_0,
    i_8_463_943_0, i_8_463_971_0, i_8_463_985_0, i_8_463_991_0,
    i_8_463_1019_0, i_8_463_1025_0, i_8_463_1029_0, i_8_463_1066_0,
    i_8_463_1110_0, i_8_463_1213_0, i_8_463_1257_0, i_8_463_1281_0,
    i_8_463_1292_0, i_8_463_1362_0, i_8_463_1371_0, i_8_463_1380_0,
    i_8_463_1451_0, i_8_463_1488_0, i_8_463_1543_0, i_8_463_1544_0,
    i_8_463_1547_0, i_8_463_1561_0, i_8_463_1675_0, i_8_463_1689_0,
    i_8_463_1699_0, i_8_463_1704_0, i_8_463_1705_0, i_8_463_1753_0,
    i_8_463_1770_0, i_8_463_1776_0, i_8_463_1806_0, i_8_463_1807_0,
    i_8_463_1815_0, i_8_463_1821_0, i_8_463_1830_0, i_8_463_1848_0,
    i_8_463_1849_0, i_8_463_1857_0, i_8_463_1858_0, i_8_463_1866_0,
    i_8_463_1911_0, i_8_463_1951_0, i_8_463_1995_0, i_8_463_2010_0,
    i_8_463_2037_0, i_8_463_2041_0, i_8_463_2082_0, i_8_463_2112_0,
    i_8_463_2149_0, i_8_463_2193_0, i_8_463_2233_0, i_8_463_2235_0,
    i_8_463_2236_0, i_8_463_2242_0, i_8_463_2272_0,
    o_8_463_0_0  );
  input  i_8_463_3_0, i_8_463_48_0, i_8_463_53_0, i_8_463_106_0,
    i_8_463_120_0, i_8_463_156_0, i_8_463_197_0, i_8_463_258_0,
    i_8_463_265_0, i_8_463_282_0, i_8_463_285_0, i_8_463_376_0,
    i_8_463_397_0, i_8_463_409_0, i_8_463_412_0, i_8_463_439_0,
    i_8_463_454_0, i_8_463_456_0, i_8_463_488_0, i_8_463_490_0,
    i_8_463_534_0, i_8_463_546_0, i_8_463_588_0, i_8_463_591_0,
    i_8_463_621_0, i_8_463_624_0, i_8_463_625_0, i_8_463_628_0,
    i_8_463_654_0, i_8_463_658_0, i_8_463_661_0, i_8_463_663_0,
    i_8_463_664_0, i_8_463_673_0, i_8_463_675_0, i_8_463_682_0,
    i_8_463_693_0, i_8_463_703_0, i_8_463_732_0, i_8_463_735_0,
    i_8_463_742_0, i_8_463_780_0, i_8_463_835_0, i_8_463_841_0,
    i_8_463_879_0, i_8_463_943_0, i_8_463_971_0, i_8_463_985_0,
    i_8_463_991_0, i_8_463_1019_0, i_8_463_1025_0, i_8_463_1029_0,
    i_8_463_1066_0, i_8_463_1110_0, i_8_463_1213_0, i_8_463_1257_0,
    i_8_463_1281_0, i_8_463_1292_0, i_8_463_1362_0, i_8_463_1371_0,
    i_8_463_1380_0, i_8_463_1451_0, i_8_463_1488_0, i_8_463_1543_0,
    i_8_463_1544_0, i_8_463_1547_0, i_8_463_1561_0, i_8_463_1675_0,
    i_8_463_1689_0, i_8_463_1699_0, i_8_463_1704_0, i_8_463_1705_0,
    i_8_463_1753_0, i_8_463_1770_0, i_8_463_1776_0, i_8_463_1806_0,
    i_8_463_1807_0, i_8_463_1815_0, i_8_463_1821_0, i_8_463_1830_0,
    i_8_463_1848_0, i_8_463_1849_0, i_8_463_1857_0, i_8_463_1858_0,
    i_8_463_1866_0, i_8_463_1911_0, i_8_463_1951_0, i_8_463_1995_0,
    i_8_463_2010_0, i_8_463_2037_0, i_8_463_2041_0, i_8_463_2082_0,
    i_8_463_2112_0, i_8_463_2149_0, i_8_463_2193_0, i_8_463_2233_0,
    i_8_463_2235_0, i_8_463_2236_0, i_8_463_2242_0, i_8_463_2272_0;
  output o_8_463_0_0;
  assign o_8_463_0_0 = 0;
endmodule



// Benchmark "kernel_8_464" written by ABC on Sun Jul 19 10:11:15 2020

module kernel_8_464 ( 
    i_8_464_33_0, i_8_464_34_0, i_8_464_70_0, i_8_464_76_0, i_8_464_77_0,
    i_8_464_141_0, i_8_464_187_0, i_8_464_191_0, i_8_464_205_0,
    i_8_464_214_0, i_8_464_215_0, i_8_464_224_0, i_8_464_267_0,
    i_8_464_268_0, i_8_464_292_0, i_8_464_330_0, i_8_464_332_0,
    i_8_464_340_0, i_8_464_358_0, i_8_464_446_0, i_8_464_448_0,
    i_8_464_456_0, i_8_464_457_0, i_8_464_463_0, i_8_464_468_0,
    i_8_464_486_0, i_8_464_557_0, i_8_464_603_0, i_8_464_618_0,
    i_8_464_619_0, i_8_464_627_0, i_8_464_637_0, i_8_464_661_0,
    i_8_464_664_0, i_8_464_719_0, i_8_464_772_0, i_8_464_787_0,
    i_8_464_825_0, i_8_464_855_0, i_8_464_879_0, i_8_464_898_0,
    i_8_464_899_0, i_8_464_925_0, i_8_464_952_0, i_8_464_953_0,
    i_8_464_987_0, i_8_464_988_0, i_8_464_998_0, i_8_464_1014_0,
    i_8_464_1015_0, i_8_464_1016_0, i_8_464_1113_0, i_8_464_1114_0,
    i_8_464_1128_0, i_8_464_1131_0, i_8_464_1132_0, i_8_464_1141_0,
    i_8_464_1186_0, i_8_464_1195_0, i_8_464_1429_0, i_8_464_1430_0,
    i_8_464_1441_0, i_8_464_1455_0, i_8_464_1510_0, i_8_464_1516_0,
    i_8_464_1537_0, i_8_464_1556_0, i_8_464_1601_0, i_8_464_1618_0,
    i_8_464_1648_0, i_8_464_1672_0, i_8_464_1673_0, i_8_464_1699_0,
    i_8_464_1734_0, i_8_464_1741_0, i_8_464_1745_0, i_8_464_1780_0,
    i_8_464_1781_0, i_8_464_1817_0, i_8_464_1857_0, i_8_464_1907_0,
    i_8_464_1933_0, i_8_464_1934_0, i_8_464_1951_0, i_8_464_2005_0,
    i_8_464_2006_0, i_8_464_2013_0, i_8_464_2014_0, i_8_464_2015_0,
    i_8_464_2050_0, i_8_464_2051_0, i_8_464_2096_0, i_8_464_2130_0,
    i_8_464_2131_0, i_8_464_2132_0, i_8_464_2139_0, i_8_464_2152_0,
    i_8_464_2263_0, i_8_464_2274_0, i_8_464_2293_0,
    o_8_464_0_0  );
  input  i_8_464_33_0, i_8_464_34_0, i_8_464_70_0, i_8_464_76_0,
    i_8_464_77_0, i_8_464_141_0, i_8_464_187_0, i_8_464_191_0,
    i_8_464_205_0, i_8_464_214_0, i_8_464_215_0, i_8_464_224_0,
    i_8_464_267_0, i_8_464_268_0, i_8_464_292_0, i_8_464_330_0,
    i_8_464_332_0, i_8_464_340_0, i_8_464_358_0, i_8_464_446_0,
    i_8_464_448_0, i_8_464_456_0, i_8_464_457_0, i_8_464_463_0,
    i_8_464_468_0, i_8_464_486_0, i_8_464_557_0, i_8_464_603_0,
    i_8_464_618_0, i_8_464_619_0, i_8_464_627_0, i_8_464_637_0,
    i_8_464_661_0, i_8_464_664_0, i_8_464_719_0, i_8_464_772_0,
    i_8_464_787_0, i_8_464_825_0, i_8_464_855_0, i_8_464_879_0,
    i_8_464_898_0, i_8_464_899_0, i_8_464_925_0, i_8_464_952_0,
    i_8_464_953_0, i_8_464_987_0, i_8_464_988_0, i_8_464_998_0,
    i_8_464_1014_0, i_8_464_1015_0, i_8_464_1016_0, i_8_464_1113_0,
    i_8_464_1114_0, i_8_464_1128_0, i_8_464_1131_0, i_8_464_1132_0,
    i_8_464_1141_0, i_8_464_1186_0, i_8_464_1195_0, i_8_464_1429_0,
    i_8_464_1430_0, i_8_464_1441_0, i_8_464_1455_0, i_8_464_1510_0,
    i_8_464_1516_0, i_8_464_1537_0, i_8_464_1556_0, i_8_464_1601_0,
    i_8_464_1618_0, i_8_464_1648_0, i_8_464_1672_0, i_8_464_1673_0,
    i_8_464_1699_0, i_8_464_1734_0, i_8_464_1741_0, i_8_464_1745_0,
    i_8_464_1780_0, i_8_464_1781_0, i_8_464_1817_0, i_8_464_1857_0,
    i_8_464_1907_0, i_8_464_1933_0, i_8_464_1934_0, i_8_464_1951_0,
    i_8_464_2005_0, i_8_464_2006_0, i_8_464_2013_0, i_8_464_2014_0,
    i_8_464_2015_0, i_8_464_2050_0, i_8_464_2051_0, i_8_464_2096_0,
    i_8_464_2130_0, i_8_464_2131_0, i_8_464_2132_0, i_8_464_2139_0,
    i_8_464_2152_0, i_8_464_2263_0, i_8_464_2274_0, i_8_464_2293_0;
  output o_8_464_0_0;
  assign o_8_464_0_0 = 0;
endmodule



// Benchmark "kernel_8_465" written by ABC on Sun Jul 19 10:11:15 2020

module kernel_8_465 ( 
    i_8_465_25_0, i_8_465_76_0, i_8_465_77_0, i_8_465_79_0, i_8_465_185_0,
    i_8_465_211_0, i_8_465_259_0, i_8_465_349_0, i_8_465_362_0,
    i_8_465_365_0, i_8_465_367_0, i_8_465_368_0, i_8_465_401_0,
    i_8_465_458_0, i_8_465_484_0, i_8_465_532_0, i_8_465_539_0,
    i_8_465_572_0, i_8_465_589_0, i_8_465_598_0, i_8_465_608_0,
    i_8_465_628_0, i_8_465_643_0, i_8_465_647_0, i_8_465_653_0,
    i_8_465_656_0, i_8_465_679_0, i_8_465_697_0, i_8_465_778_0,
    i_8_465_781_0, i_8_465_782_0, i_8_465_784_0, i_8_465_796_0,
    i_8_465_815_0, i_8_465_817_0, i_8_465_833_0, i_8_465_838_0,
    i_8_465_839_0, i_8_465_851_0, i_8_465_853_0, i_8_465_862_0,
    i_8_465_878_0, i_8_465_959_0, i_8_465_1067_0, i_8_465_1070_0,
    i_8_465_1075_0, i_8_465_1134_0, i_8_465_1222_0, i_8_465_1254_0,
    i_8_465_1264_0, i_8_465_1282_0, i_8_465_1283_0, i_8_465_1286_0,
    i_8_465_1304_0, i_8_465_1305_0, i_8_465_1327_0, i_8_465_1337_0,
    i_8_465_1379_0, i_8_465_1391_0, i_8_465_1423_0, i_8_465_1427_0,
    i_8_465_1436_0, i_8_465_1444_0, i_8_465_1463_0, i_8_465_1466_0,
    i_8_465_1484_0, i_8_465_1514_0, i_8_465_1549_0, i_8_465_1613_0,
    i_8_465_1619_0, i_8_465_1630_0, i_8_465_1633_0, i_8_465_1688_0,
    i_8_465_1706_0, i_8_465_1721_0, i_8_465_1750_0, i_8_465_1751_0,
    i_8_465_1799_0, i_8_465_1803_0, i_8_465_1807_0, i_8_465_1877_0,
    i_8_465_1883_0, i_8_465_1898_0, i_8_465_1927_0, i_8_465_1951_0,
    i_8_465_1988_0, i_8_465_1993_0, i_8_465_1994_0, i_8_465_2006_0,
    i_8_465_2024_0, i_8_465_2093_0, i_8_465_2140_0, i_8_465_2144_0,
    i_8_465_2147_0, i_8_465_2158_0, i_8_465_2159_0, i_8_465_2229_0,
    i_8_465_2261_0, i_8_465_2263_0, i_8_465_2267_0,
    o_8_465_0_0  );
  input  i_8_465_25_0, i_8_465_76_0, i_8_465_77_0, i_8_465_79_0,
    i_8_465_185_0, i_8_465_211_0, i_8_465_259_0, i_8_465_349_0,
    i_8_465_362_0, i_8_465_365_0, i_8_465_367_0, i_8_465_368_0,
    i_8_465_401_0, i_8_465_458_0, i_8_465_484_0, i_8_465_532_0,
    i_8_465_539_0, i_8_465_572_0, i_8_465_589_0, i_8_465_598_0,
    i_8_465_608_0, i_8_465_628_0, i_8_465_643_0, i_8_465_647_0,
    i_8_465_653_0, i_8_465_656_0, i_8_465_679_0, i_8_465_697_0,
    i_8_465_778_0, i_8_465_781_0, i_8_465_782_0, i_8_465_784_0,
    i_8_465_796_0, i_8_465_815_0, i_8_465_817_0, i_8_465_833_0,
    i_8_465_838_0, i_8_465_839_0, i_8_465_851_0, i_8_465_853_0,
    i_8_465_862_0, i_8_465_878_0, i_8_465_959_0, i_8_465_1067_0,
    i_8_465_1070_0, i_8_465_1075_0, i_8_465_1134_0, i_8_465_1222_0,
    i_8_465_1254_0, i_8_465_1264_0, i_8_465_1282_0, i_8_465_1283_0,
    i_8_465_1286_0, i_8_465_1304_0, i_8_465_1305_0, i_8_465_1327_0,
    i_8_465_1337_0, i_8_465_1379_0, i_8_465_1391_0, i_8_465_1423_0,
    i_8_465_1427_0, i_8_465_1436_0, i_8_465_1444_0, i_8_465_1463_0,
    i_8_465_1466_0, i_8_465_1484_0, i_8_465_1514_0, i_8_465_1549_0,
    i_8_465_1613_0, i_8_465_1619_0, i_8_465_1630_0, i_8_465_1633_0,
    i_8_465_1688_0, i_8_465_1706_0, i_8_465_1721_0, i_8_465_1750_0,
    i_8_465_1751_0, i_8_465_1799_0, i_8_465_1803_0, i_8_465_1807_0,
    i_8_465_1877_0, i_8_465_1883_0, i_8_465_1898_0, i_8_465_1927_0,
    i_8_465_1951_0, i_8_465_1988_0, i_8_465_1993_0, i_8_465_1994_0,
    i_8_465_2006_0, i_8_465_2024_0, i_8_465_2093_0, i_8_465_2140_0,
    i_8_465_2144_0, i_8_465_2147_0, i_8_465_2158_0, i_8_465_2159_0,
    i_8_465_2229_0, i_8_465_2261_0, i_8_465_2263_0, i_8_465_2267_0;
  output o_8_465_0_0;
  assign o_8_465_0_0 = 0;
endmodule



// Benchmark "kernel_8_466" written by ABC on Sun Jul 19 10:11:17 2020

module kernel_8_466 ( 
    i_8_466_39_0, i_8_466_52_0, i_8_466_66_0, i_8_466_69_0, i_8_466_139_0,
    i_8_466_169_0, i_8_466_174_0, i_8_466_183_0, i_8_466_192_0,
    i_8_466_210_0, i_8_466_232_0, i_8_466_264_0, i_8_466_270_0,
    i_8_466_291_0, i_8_466_295_0, i_8_466_327_0, i_8_466_345_0,
    i_8_466_348_0, i_8_466_366_0, i_8_466_384_0, i_8_466_445_0,
    i_8_466_462_0, i_8_466_466_0, i_8_466_528_0, i_8_466_552_0,
    i_8_466_554_0, i_8_466_598_0, i_8_466_633_0, i_8_466_662_0,
    i_8_466_664_0, i_8_466_674_0, i_8_466_687_0, i_8_466_699_0,
    i_8_466_704_0, i_8_466_768_0, i_8_466_770_0, i_8_466_777_0,
    i_8_466_843_0, i_8_466_858_0, i_8_466_877_0, i_8_466_880_0,
    i_8_466_990_0, i_8_466_993_0, i_8_466_1056_0, i_8_466_1107_0,
    i_8_466_1113_0, i_8_466_1119_0, i_8_466_1155_0, i_8_466_1156_0,
    i_8_466_1158_0, i_8_466_1159_0, i_8_466_1173_0, i_8_466_1185_0,
    i_8_466_1191_0, i_8_466_1230_0, i_8_466_1231_0, i_8_466_1233_0,
    i_8_466_1237_0, i_8_466_1272_0, i_8_466_1302_0, i_8_466_1317_0,
    i_8_466_1324_0, i_8_466_1380_0, i_8_466_1452_0, i_8_466_1470_0,
    i_8_466_1509_0, i_8_466_1540_0, i_8_466_1542_0, i_8_466_1596_0,
    i_8_466_1600_0, i_8_466_1633_0, i_8_466_1704_0, i_8_466_1731_0,
    i_8_466_1740_0, i_8_466_1753_0, i_8_466_1806_0, i_8_466_1816_0,
    i_8_466_1830_0, i_8_466_1843_0, i_8_466_1879_0, i_8_466_1906_0,
    i_8_466_1948_0, i_8_466_1966_0, i_8_466_1969_0, i_8_466_1975_0,
    i_8_466_1989_0, i_8_466_1995_0, i_8_466_2109_0, i_8_466_2112_0,
    i_8_466_2114_0, i_8_466_2145_0, i_8_466_2152_0, i_8_466_2155_0,
    i_8_466_2158_0, i_8_466_2181_0, i_8_466_2182_0, i_8_466_2190_0,
    i_8_466_2211_0, i_8_466_2226_0, i_8_466_2275_0,
    o_8_466_0_0  );
  input  i_8_466_39_0, i_8_466_52_0, i_8_466_66_0, i_8_466_69_0,
    i_8_466_139_0, i_8_466_169_0, i_8_466_174_0, i_8_466_183_0,
    i_8_466_192_0, i_8_466_210_0, i_8_466_232_0, i_8_466_264_0,
    i_8_466_270_0, i_8_466_291_0, i_8_466_295_0, i_8_466_327_0,
    i_8_466_345_0, i_8_466_348_0, i_8_466_366_0, i_8_466_384_0,
    i_8_466_445_0, i_8_466_462_0, i_8_466_466_0, i_8_466_528_0,
    i_8_466_552_0, i_8_466_554_0, i_8_466_598_0, i_8_466_633_0,
    i_8_466_662_0, i_8_466_664_0, i_8_466_674_0, i_8_466_687_0,
    i_8_466_699_0, i_8_466_704_0, i_8_466_768_0, i_8_466_770_0,
    i_8_466_777_0, i_8_466_843_0, i_8_466_858_0, i_8_466_877_0,
    i_8_466_880_0, i_8_466_990_0, i_8_466_993_0, i_8_466_1056_0,
    i_8_466_1107_0, i_8_466_1113_0, i_8_466_1119_0, i_8_466_1155_0,
    i_8_466_1156_0, i_8_466_1158_0, i_8_466_1159_0, i_8_466_1173_0,
    i_8_466_1185_0, i_8_466_1191_0, i_8_466_1230_0, i_8_466_1231_0,
    i_8_466_1233_0, i_8_466_1237_0, i_8_466_1272_0, i_8_466_1302_0,
    i_8_466_1317_0, i_8_466_1324_0, i_8_466_1380_0, i_8_466_1452_0,
    i_8_466_1470_0, i_8_466_1509_0, i_8_466_1540_0, i_8_466_1542_0,
    i_8_466_1596_0, i_8_466_1600_0, i_8_466_1633_0, i_8_466_1704_0,
    i_8_466_1731_0, i_8_466_1740_0, i_8_466_1753_0, i_8_466_1806_0,
    i_8_466_1816_0, i_8_466_1830_0, i_8_466_1843_0, i_8_466_1879_0,
    i_8_466_1906_0, i_8_466_1948_0, i_8_466_1966_0, i_8_466_1969_0,
    i_8_466_1975_0, i_8_466_1989_0, i_8_466_1995_0, i_8_466_2109_0,
    i_8_466_2112_0, i_8_466_2114_0, i_8_466_2145_0, i_8_466_2152_0,
    i_8_466_2155_0, i_8_466_2158_0, i_8_466_2181_0, i_8_466_2182_0,
    i_8_466_2190_0, i_8_466_2211_0, i_8_466_2226_0, i_8_466_2275_0;
  output o_8_466_0_0;
  assign o_8_466_0_0 = ~((~i_8_466_139_0 & ((~i_8_466_52_0 & i_8_466_1107_0 & ~i_8_466_1185_0 & ~i_8_466_1452_0 & ~i_8_466_1542_0 & ~i_8_466_1806_0 & ~i_8_466_2112_0) | (~i_8_466_39_0 & ~i_8_466_1237_0 & ~i_8_466_1830_0 & ~i_8_466_2181_0 & ~i_8_466_2190_0))) | (~i_8_466_52_0 & ((~i_8_466_993_0 & ~i_8_466_1230_0 & i_8_466_1233_0 & ~i_8_466_2109_0 & ~i_8_466_2112_0 & ~i_8_466_2181_0) | (~i_8_466_264_0 & i_8_466_598_0 & ~i_8_466_1056_0 & i_8_466_1113_0 & ~i_8_466_1324_0 & ~i_8_466_1600_0 & ~i_8_466_1989_0 & ~i_8_466_2211_0))) | (~i_8_466_210_0 & ((~i_8_466_552_0 & ~i_8_466_768_0 & ~i_8_466_1113_0 & ~i_8_466_1173_0 & ~i_8_466_1324_0 & ~i_8_466_1704_0 & ~i_8_466_1740_0) | (~i_8_466_39_0 & ~i_8_466_264_0 & ~i_8_466_366_0 & ~i_8_466_633_0 & ~i_8_466_1155_0 & ~i_8_466_1596_0 & ~i_8_466_2275_0))) | (~i_8_466_345_0 & ~i_8_466_1272_0 & ((~i_8_466_291_0 & ~i_8_466_843_0 & ~i_8_466_1119_0 & ~i_8_466_1542_0) | (~i_8_466_348_0 & ~i_8_466_1830_0 & ~i_8_466_2182_0))) | (~i_8_466_990_0 & ~i_8_466_1740_0 & ((i_8_466_1113_0 & ~i_8_466_1155_0 & ~i_8_466_1158_0 & i_8_466_1302_0 & ~i_8_466_1906_0) | (~i_8_466_327_0 & ~i_8_466_384_0 & ~i_8_466_770_0 & ~i_8_466_1119_0 & ~i_8_466_1542_0 & ~i_8_466_2190_0 & ~i_8_466_2275_0))) | (~i_8_466_1380_0 & ((~i_8_466_39_0 & i_8_466_1155_0 & i_8_466_1158_0 & ~i_8_466_1540_0 & ~i_8_466_1596_0) | (~i_8_466_169_0 & ~i_8_466_174_0 & ~i_8_466_264_0 & ~i_8_466_768_0 & ~i_8_466_1158_0 & ~i_8_466_2182_0))) | (~i_8_466_39_0 & ((~i_8_466_192_0 & ~i_8_466_462_0 & ~i_8_466_843_0 & i_8_466_877_0 & ~i_8_466_1185_0 & ~i_8_466_1237_0) | (~i_8_466_183_0 & ~i_8_466_1107_0 & ~i_8_466_1470_0 & ~i_8_466_2155_0 & ~i_8_466_2226_0))) | (~i_8_466_291_0 & ((~i_8_466_183_0 & ((i_8_466_39_0 & ~i_8_466_687_0 & ~i_8_466_1509_0 & ~i_8_466_1542_0 & ~i_8_466_1633_0 & ~i_8_466_1969_0) | (~i_8_466_662_0 & ~i_8_466_1155_0 & ~i_8_466_1540_0 & ~i_8_466_1989_0 & ~i_8_466_2182_0 & ~i_8_466_2211_0))) | (~i_8_466_1119_0 & ~i_8_466_1231_0 & ~i_8_466_1324_0 & ~i_8_466_1989_0 & ~i_8_466_2181_0 & ~i_8_466_2226_0))) | (~i_8_466_66_0 & ~i_8_466_183_0 & ~i_8_466_528_0 & ~i_8_466_1830_0 & ~i_8_466_2190_0));
endmodule



// Benchmark "kernel_8_467" written by ABC on Sun Jul 19 10:11:17 2020

module kernel_8_467 ( 
    i_8_467_32_0, i_8_467_34_0, i_8_467_87_0, i_8_467_107_0, i_8_467_160_0,
    i_8_467_213_0, i_8_467_220_0, i_8_467_224_0, i_8_467_256_0,
    i_8_467_302_0, i_8_467_327_0, i_8_467_328_0, i_8_467_383_0,
    i_8_467_418_0, i_8_467_421_0, i_8_467_440_0, i_8_467_442_0,
    i_8_467_463_0, i_8_467_472_0, i_8_467_485_0, i_8_467_502_0,
    i_8_467_510_0, i_8_467_526_0, i_8_467_547_0, i_8_467_599_0,
    i_8_467_616_0, i_8_467_625_0, i_8_467_627_0, i_8_467_637_0,
    i_8_467_658_0, i_8_467_716_0, i_8_467_723_0, i_8_467_726_0,
    i_8_467_759_0, i_8_467_760_0, i_8_467_769_0, i_8_467_773_0,
    i_8_467_781_0, i_8_467_782_0, i_8_467_795_0, i_8_467_814_0,
    i_8_467_850_0, i_8_467_880_0, i_8_467_881_0, i_8_467_895_0,
    i_8_467_896_0, i_8_467_898_0, i_8_467_1012_0, i_8_467_1013_0,
    i_8_467_1029_0, i_8_467_1109_0, i_8_467_1115_0, i_8_467_1156_0,
    i_8_467_1159_0, i_8_467_1318_0, i_8_467_1345_0, i_8_467_1347_0,
    i_8_467_1348_0, i_8_467_1452_0, i_8_467_1453_0, i_8_467_1471_0,
    i_8_467_1472_0, i_8_467_1537_0, i_8_467_1544_0, i_8_467_1552_0,
    i_8_467_1579_0, i_8_467_1599_0, i_8_467_1603_0, i_8_467_1615_0,
    i_8_467_1633_0, i_8_467_1670_0, i_8_467_1681_0, i_8_467_1714_0,
    i_8_467_1715_0, i_8_467_1717_0, i_8_467_1726_0, i_8_467_1727_0,
    i_8_467_1748_0, i_8_467_1759_0, i_8_467_1762_0, i_8_467_1805_0,
    i_8_467_1860_0, i_8_467_1883_0, i_8_467_1895_0, i_8_467_1903_0,
    i_8_467_1931_0, i_8_467_1965_0, i_8_467_1995_0, i_8_467_2002_0,
    i_8_467_2012_0, i_8_467_2031_0, i_8_467_2049_0, i_8_467_2050_0,
    i_8_467_2110_0, i_8_467_2111_0, i_8_467_2136_0, i_8_467_2145_0,
    i_8_467_2146_0, i_8_467_2149_0, i_8_467_2215_0,
    o_8_467_0_0  );
  input  i_8_467_32_0, i_8_467_34_0, i_8_467_87_0, i_8_467_107_0,
    i_8_467_160_0, i_8_467_213_0, i_8_467_220_0, i_8_467_224_0,
    i_8_467_256_0, i_8_467_302_0, i_8_467_327_0, i_8_467_328_0,
    i_8_467_383_0, i_8_467_418_0, i_8_467_421_0, i_8_467_440_0,
    i_8_467_442_0, i_8_467_463_0, i_8_467_472_0, i_8_467_485_0,
    i_8_467_502_0, i_8_467_510_0, i_8_467_526_0, i_8_467_547_0,
    i_8_467_599_0, i_8_467_616_0, i_8_467_625_0, i_8_467_627_0,
    i_8_467_637_0, i_8_467_658_0, i_8_467_716_0, i_8_467_723_0,
    i_8_467_726_0, i_8_467_759_0, i_8_467_760_0, i_8_467_769_0,
    i_8_467_773_0, i_8_467_781_0, i_8_467_782_0, i_8_467_795_0,
    i_8_467_814_0, i_8_467_850_0, i_8_467_880_0, i_8_467_881_0,
    i_8_467_895_0, i_8_467_896_0, i_8_467_898_0, i_8_467_1012_0,
    i_8_467_1013_0, i_8_467_1029_0, i_8_467_1109_0, i_8_467_1115_0,
    i_8_467_1156_0, i_8_467_1159_0, i_8_467_1318_0, i_8_467_1345_0,
    i_8_467_1347_0, i_8_467_1348_0, i_8_467_1452_0, i_8_467_1453_0,
    i_8_467_1471_0, i_8_467_1472_0, i_8_467_1537_0, i_8_467_1544_0,
    i_8_467_1552_0, i_8_467_1579_0, i_8_467_1599_0, i_8_467_1603_0,
    i_8_467_1615_0, i_8_467_1633_0, i_8_467_1670_0, i_8_467_1681_0,
    i_8_467_1714_0, i_8_467_1715_0, i_8_467_1717_0, i_8_467_1726_0,
    i_8_467_1727_0, i_8_467_1748_0, i_8_467_1759_0, i_8_467_1762_0,
    i_8_467_1805_0, i_8_467_1860_0, i_8_467_1883_0, i_8_467_1895_0,
    i_8_467_1903_0, i_8_467_1931_0, i_8_467_1965_0, i_8_467_1995_0,
    i_8_467_2002_0, i_8_467_2012_0, i_8_467_2031_0, i_8_467_2049_0,
    i_8_467_2050_0, i_8_467_2110_0, i_8_467_2111_0, i_8_467_2136_0,
    i_8_467_2145_0, i_8_467_2146_0, i_8_467_2149_0, i_8_467_2215_0;
  output o_8_467_0_0;
  assign o_8_467_0_0 = 0;
endmodule



// Benchmark "kernel_8_468" written by ABC on Sun Jul 19 10:11:18 2020

module kernel_8_468 ( 
    i_8_468_13_0, i_8_468_35_0, i_8_468_41_0, i_8_468_87_0, i_8_468_142_0,
    i_8_468_187_0, i_8_468_189_0, i_8_468_190_0, i_8_468_214_0,
    i_8_468_224_0, i_8_468_228_0, i_8_468_300_0, i_8_468_347_0,
    i_8_468_368_0, i_8_468_377_0, i_8_468_381_0, i_8_468_383_0,
    i_8_468_429_0, i_8_468_431_0, i_8_468_444_0, i_8_468_454_0,
    i_8_468_457_0, i_8_468_488_0, i_8_468_505_0, i_8_468_510_0,
    i_8_468_511_0, i_8_468_557_0, i_8_468_605_0, i_8_468_629_0,
    i_8_468_661_0, i_8_468_682_0, i_8_468_688_0, i_8_468_696_0,
    i_8_468_699_0, i_8_468_700_0, i_8_468_707_0, i_8_468_710_0,
    i_8_468_719_0, i_8_468_743_0, i_8_468_764_0, i_8_468_815_0,
    i_8_468_845_0, i_8_468_868_0, i_8_468_869_0, i_8_468_877_0,
    i_8_468_951_0, i_8_468_971_0, i_8_468_977_0, i_8_468_980_0,
    i_8_468_1065_0, i_8_468_1106_0, i_8_468_1112_0, i_8_468_1132_0,
    i_8_468_1184_0, i_8_468_1193_0, i_8_468_1225_0, i_8_468_1232_0,
    i_8_468_1240_0, i_8_468_1249_0, i_8_468_1268_0, i_8_468_1344_0,
    i_8_468_1353_0, i_8_468_1417_0, i_8_468_1433_0, i_8_468_1519_0,
    i_8_468_1537_0, i_8_468_1544_0, i_8_468_1564_0, i_8_468_1581_0,
    i_8_468_1637_0, i_8_468_1650_0, i_8_468_1654_0, i_8_468_1673_0,
    i_8_468_1707_0, i_8_468_1717_0, i_8_468_1732_0, i_8_468_1792_0,
    i_8_468_1808_0, i_8_468_1815_0, i_8_468_1822_0, i_8_468_1861_0,
    i_8_468_1888_0, i_8_468_1922_0, i_8_468_1933_0, i_8_468_1947_0,
    i_8_468_2046_0, i_8_468_2056_0, i_8_468_2092_0, i_8_468_2111_0,
    i_8_468_2112_0, i_8_468_2131_0, i_8_468_2136_0, i_8_468_2137_0,
    i_8_468_2147_0, i_8_468_2214_0, i_8_468_2218_0, i_8_468_2219_0,
    i_8_468_2231_0, i_8_468_2244_0, i_8_468_2247_0,
    o_8_468_0_0  );
  input  i_8_468_13_0, i_8_468_35_0, i_8_468_41_0, i_8_468_87_0,
    i_8_468_142_0, i_8_468_187_0, i_8_468_189_0, i_8_468_190_0,
    i_8_468_214_0, i_8_468_224_0, i_8_468_228_0, i_8_468_300_0,
    i_8_468_347_0, i_8_468_368_0, i_8_468_377_0, i_8_468_381_0,
    i_8_468_383_0, i_8_468_429_0, i_8_468_431_0, i_8_468_444_0,
    i_8_468_454_0, i_8_468_457_0, i_8_468_488_0, i_8_468_505_0,
    i_8_468_510_0, i_8_468_511_0, i_8_468_557_0, i_8_468_605_0,
    i_8_468_629_0, i_8_468_661_0, i_8_468_682_0, i_8_468_688_0,
    i_8_468_696_0, i_8_468_699_0, i_8_468_700_0, i_8_468_707_0,
    i_8_468_710_0, i_8_468_719_0, i_8_468_743_0, i_8_468_764_0,
    i_8_468_815_0, i_8_468_845_0, i_8_468_868_0, i_8_468_869_0,
    i_8_468_877_0, i_8_468_951_0, i_8_468_971_0, i_8_468_977_0,
    i_8_468_980_0, i_8_468_1065_0, i_8_468_1106_0, i_8_468_1112_0,
    i_8_468_1132_0, i_8_468_1184_0, i_8_468_1193_0, i_8_468_1225_0,
    i_8_468_1232_0, i_8_468_1240_0, i_8_468_1249_0, i_8_468_1268_0,
    i_8_468_1344_0, i_8_468_1353_0, i_8_468_1417_0, i_8_468_1433_0,
    i_8_468_1519_0, i_8_468_1537_0, i_8_468_1544_0, i_8_468_1564_0,
    i_8_468_1581_0, i_8_468_1637_0, i_8_468_1650_0, i_8_468_1654_0,
    i_8_468_1673_0, i_8_468_1707_0, i_8_468_1717_0, i_8_468_1732_0,
    i_8_468_1792_0, i_8_468_1808_0, i_8_468_1815_0, i_8_468_1822_0,
    i_8_468_1861_0, i_8_468_1888_0, i_8_468_1922_0, i_8_468_1933_0,
    i_8_468_1947_0, i_8_468_2046_0, i_8_468_2056_0, i_8_468_2092_0,
    i_8_468_2111_0, i_8_468_2112_0, i_8_468_2131_0, i_8_468_2136_0,
    i_8_468_2137_0, i_8_468_2147_0, i_8_468_2214_0, i_8_468_2218_0,
    i_8_468_2219_0, i_8_468_2231_0, i_8_468_2244_0, i_8_468_2247_0;
  output o_8_468_0_0;
  assign o_8_468_0_0 = 0;
endmodule



// Benchmark "kernel_8_469" written by ABC on Sun Jul 19 10:11:19 2020

module kernel_8_469 ( 
    i_8_469_11_0, i_8_469_26_0, i_8_469_51_0, i_8_469_77_0, i_8_469_86_0,
    i_8_469_107_0, i_8_469_165_0, i_8_469_246_0, i_8_469_255_0,
    i_8_469_256_0, i_8_469_262_0, i_8_469_303_0, i_8_469_310_0,
    i_8_469_318_0, i_8_469_321_0, i_8_469_361_0, i_8_469_368_0,
    i_8_469_436_0, i_8_469_492_0, i_8_469_535_0, i_8_469_552_0,
    i_8_469_579_0, i_8_469_580_0, i_8_469_595_0, i_8_469_598_0,
    i_8_469_609_0, i_8_469_624_0, i_8_469_625_0, i_8_469_636_0,
    i_8_469_639_0, i_8_469_657_0, i_8_469_660_0, i_8_469_661_0,
    i_8_469_675_0, i_8_469_678_0, i_8_469_696_0, i_8_469_705_0,
    i_8_469_715_0, i_8_469_778_0, i_8_469_786_0, i_8_469_791_0,
    i_8_469_823_0, i_8_469_843_0, i_8_469_844_0, i_8_469_846_0,
    i_8_469_847_0, i_8_469_850_0, i_8_469_968_0, i_8_469_1040_0,
    i_8_469_1061_0, i_8_469_1074_0, i_8_469_1139_0, i_8_469_1146_0,
    i_8_469_1229_0, i_8_469_1233_0, i_8_469_1246_0, i_8_469_1255_0,
    i_8_469_1273_0, i_8_469_1284_0, i_8_469_1303_0, i_8_469_1317_0,
    i_8_469_1336_0, i_8_469_1359_0, i_8_469_1362_0, i_8_469_1387_0,
    i_8_469_1396_0, i_8_469_1455_0, i_8_469_1458_0, i_8_469_1470_0,
    i_8_469_1471_0, i_8_469_1489_0, i_8_469_1543_0, i_8_469_1545_0,
    i_8_469_1547_0, i_8_469_1570_0, i_8_469_1696_0, i_8_469_1697_0,
    i_8_469_1702_0, i_8_469_1733_0, i_8_469_1767_0, i_8_469_1804_0,
    i_8_469_1819_0, i_8_469_1839_0, i_8_469_1884_0, i_8_469_1885_0,
    i_8_469_1902_0, i_8_469_1911_0, i_8_469_1912_0, i_8_469_1997_0,
    i_8_469_2028_0, i_8_469_2095_0, i_8_469_2096_0, i_8_469_2129_0,
    i_8_469_2133_0, i_8_469_2140_0, i_8_469_2173_0, i_8_469_2191_0,
    i_8_469_2194_0, i_8_469_2284_0, i_8_469_2289_0,
    o_8_469_0_0  );
  input  i_8_469_11_0, i_8_469_26_0, i_8_469_51_0, i_8_469_77_0,
    i_8_469_86_0, i_8_469_107_0, i_8_469_165_0, i_8_469_246_0,
    i_8_469_255_0, i_8_469_256_0, i_8_469_262_0, i_8_469_303_0,
    i_8_469_310_0, i_8_469_318_0, i_8_469_321_0, i_8_469_361_0,
    i_8_469_368_0, i_8_469_436_0, i_8_469_492_0, i_8_469_535_0,
    i_8_469_552_0, i_8_469_579_0, i_8_469_580_0, i_8_469_595_0,
    i_8_469_598_0, i_8_469_609_0, i_8_469_624_0, i_8_469_625_0,
    i_8_469_636_0, i_8_469_639_0, i_8_469_657_0, i_8_469_660_0,
    i_8_469_661_0, i_8_469_675_0, i_8_469_678_0, i_8_469_696_0,
    i_8_469_705_0, i_8_469_715_0, i_8_469_778_0, i_8_469_786_0,
    i_8_469_791_0, i_8_469_823_0, i_8_469_843_0, i_8_469_844_0,
    i_8_469_846_0, i_8_469_847_0, i_8_469_850_0, i_8_469_968_0,
    i_8_469_1040_0, i_8_469_1061_0, i_8_469_1074_0, i_8_469_1139_0,
    i_8_469_1146_0, i_8_469_1229_0, i_8_469_1233_0, i_8_469_1246_0,
    i_8_469_1255_0, i_8_469_1273_0, i_8_469_1284_0, i_8_469_1303_0,
    i_8_469_1317_0, i_8_469_1336_0, i_8_469_1359_0, i_8_469_1362_0,
    i_8_469_1387_0, i_8_469_1396_0, i_8_469_1455_0, i_8_469_1458_0,
    i_8_469_1470_0, i_8_469_1471_0, i_8_469_1489_0, i_8_469_1543_0,
    i_8_469_1545_0, i_8_469_1547_0, i_8_469_1570_0, i_8_469_1696_0,
    i_8_469_1697_0, i_8_469_1702_0, i_8_469_1733_0, i_8_469_1767_0,
    i_8_469_1804_0, i_8_469_1819_0, i_8_469_1839_0, i_8_469_1884_0,
    i_8_469_1885_0, i_8_469_1902_0, i_8_469_1911_0, i_8_469_1912_0,
    i_8_469_1997_0, i_8_469_2028_0, i_8_469_2095_0, i_8_469_2096_0,
    i_8_469_2129_0, i_8_469_2133_0, i_8_469_2140_0, i_8_469_2173_0,
    i_8_469_2191_0, i_8_469_2194_0, i_8_469_2284_0, i_8_469_2289_0;
  output o_8_469_0_0;
  assign o_8_469_0_0 = 0;
endmodule



// Benchmark "kernel_8_470" written by ABC on Sun Jul 19 10:11:20 2020

module kernel_8_470 ( 
    i_8_470_19_0, i_8_470_21_0, i_8_470_28_0, i_8_470_30_0, i_8_470_34_0,
    i_8_470_37_0, i_8_470_229_0, i_8_470_340_0, i_8_470_364_0,
    i_8_470_365_0, i_8_470_366_0, i_8_470_468_0, i_8_470_469_0,
    i_8_470_478_0, i_8_470_480_0, i_8_470_487_0, i_8_470_490_0,
    i_8_470_528_0, i_8_470_540_0, i_8_470_567_0, i_8_470_568_0,
    i_8_470_611_0, i_8_470_612_0, i_8_470_622_0, i_8_470_652_0,
    i_8_470_656_0, i_8_470_685_0, i_8_470_709_0, i_8_470_755_0,
    i_8_470_766_0, i_8_470_789_0, i_8_470_844_0, i_8_470_875_0,
    i_8_470_928_0, i_8_470_983_0, i_8_470_992_0, i_8_470_997_0,
    i_8_470_999_0, i_8_470_1029_0, i_8_470_1042_0, i_8_470_1099_0,
    i_8_470_1127_0, i_8_470_1225_0, i_8_470_1226_0, i_8_470_1261_0,
    i_8_470_1262_0, i_8_470_1271_0, i_8_470_1277_0, i_8_470_1280_0,
    i_8_470_1283_0, i_8_470_1288_0, i_8_470_1297_0, i_8_470_1324_0,
    i_8_470_1325_0, i_8_470_1378_0, i_8_470_1379_0, i_8_470_1407_0,
    i_8_470_1468_0, i_8_470_1486_0, i_8_470_1495_0, i_8_470_1536_0,
    i_8_470_1538_0, i_8_470_1541_0, i_8_470_1549_0, i_8_470_1675_0,
    i_8_470_1681_0, i_8_470_1682_0, i_8_470_1696_0, i_8_470_1741_0,
    i_8_470_1752_0, i_8_470_1765_0, i_8_470_1772_0, i_8_470_1817_0,
    i_8_470_1820_0, i_8_470_1825_0, i_8_470_1827_0, i_8_470_1867_0,
    i_8_470_1888_0, i_8_470_1889_0, i_8_470_1900_0, i_8_470_1946_0,
    i_8_470_1971_0, i_8_470_1975_0, i_8_470_2000_0, i_8_470_2015_0,
    i_8_470_2052_0, i_8_470_2053_0, i_8_470_2130_0, i_8_470_2132_0,
    i_8_470_2133_0, i_8_470_2139_0, i_8_470_2145_0, i_8_470_2152_0,
    i_8_470_2224_0, i_8_470_2230_0, i_8_470_2242_0, i_8_470_2243_0,
    i_8_470_2246_0, i_8_470_2270_0, i_8_470_2273_0,
    o_8_470_0_0  );
  input  i_8_470_19_0, i_8_470_21_0, i_8_470_28_0, i_8_470_30_0,
    i_8_470_34_0, i_8_470_37_0, i_8_470_229_0, i_8_470_340_0,
    i_8_470_364_0, i_8_470_365_0, i_8_470_366_0, i_8_470_468_0,
    i_8_470_469_0, i_8_470_478_0, i_8_470_480_0, i_8_470_487_0,
    i_8_470_490_0, i_8_470_528_0, i_8_470_540_0, i_8_470_567_0,
    i_8_470_568_0, i_8_470_611_0, i_8_470_612_0, i_8_470_622_0,
    i_8_470_652_0, i_8_470_656_0, i_8_470_685_0, i_8_470_709_0,
    i_8_470_755_0, i_8_470_766_0, i_8_470_789_0, i_8_470_844_0,
    i_8_470_875_0, i_8_470_928_0, i_8_470_983_0, i_8_470_992_0,
    i_8_470_997_0, i_8_470_999_0, i_8_470_1029_0, i_8_470_1042_0,
    i_8_470_1099_0, i_8_470_1127_0, i_8_470_1225_0, i_8_470_1226_0,
    i_8_470_1261_0, i_8_470_1262_0, i_8_470_1271_0, i_8_470_1277_0,
    i_8_470_1280_0, i_8_470_1283_0, i_8_470_1288_0, i_8_470_1297_0,
    i_8_470_1324_0, i_8_470_1325_0, i_8_470_1378_0, i_8_470_1379_0,
    i_8_470_1407_0, i_8_470_1468_0, i_8_470_1486_0, i_8_470_1495_0,
    i_8_470_1536_0, i_8_470_1538_0, i_8_470_1541_0, i_8_470_1549_0,
    i_8_470_1675_0, i_8_470_1681_0, i_8_470_1682_0, i_8_470_1696_0,
    i_8_470_1741_0, i_8_470_1752_0, i_8_470_1765_0, i_8_470_1772_0,
    i_8_470_1817_0, i_8_470_1820_0, i_8_470_1825_0, i_8_470_1827_0,
    i_8_470_1867_0, i_8_470_1888_0, i_8_470_1889_0, i_8_470_1900_0,
    i_8_470_1946_0, i_8_470_1971_0, i_8_470_1975_0, i_8_470_2000_0,
    i_8_470_2015_0, i_8_470_2052_0, i_8_470_2053_0, i_8_470_2130_0,
    i_8_470_2132_0, i_8_470_2133_0, i_8_470_2139_0, i_8_470_2145_0,
    i_8_470_2152_0, i_8_470_2224_0, i_8_470_2230_0, i_8_470_2242_0,
    i_8_470_2243_0, i_8_470_2246_0, i_8_470_2270_0, i_8_470_2273_0;
  output o_8_470_0_0;
  assign o_8_470_0_0 = 0;
endmodule



// Benchmark "kernel_8_471" written by ABC on Sun Jul 19 10:11:21 2020

module kernel_8_471 ( 
    i_8_471_64_0, i_8_471_141_0, i_8_471_165_0, i_8_471_238_0,
    i_8_471_265_0, i_8_471_297_0, i_8_471_334_0, i_8_471_352_0,
    i_8_471_361_0, i_8_471_379_0, i_8_471_399_0, i_8_471_400_0,
    i_8_471_418_0, i_8_471_453_0, i_8_471_481_0, i_8_471_493_0,
    i_8_471_524_0, i_8_471_525_0, i_8_471_526_0, i_8_471_541_0,
    i_8_471_550_0, i_8_471_552_0, i_8_471_553_0, i_8_471_570_0,
    i_8_471_571_0, i_8_471_580_0, i_8_471_589_0, i_8_471_606_0,
    i_8_471_659_0, i_8_471_661_0, i_8_471_662_0, i_8_471_687_0,
    i_8_471_688_0, i_8_471_708_0, i_8_471_760_0, i_8_471_804_0,
    i_8_471_837_0, i_8_471_840_0, i_8_471_874_0, i_8_471_990_0,
    i_8_471_1057_0, i_8_471_1058_0, i_8_471_1111_0, i_8_471_1183_0,
    i_8_471_1200_0, i_8_471_1238_0, i_8_471_1266_0, i_8_471_1267_0,
    i_8_471_1271_0, i_8_471_1288_0, i_8_471_1291_0, i_8_471_1308_0,
    i_8_471_1399_0, i_8_471_1411_0, i_8_471_1416_0, i_8_471_1432_0,
    i_8_471_1437_0, i_8_471_1441_0, i_8_471_1462_0, i_8_471_1515_0,
    i_8_471_1544_0, i_8_471_1546_0, i_8_471_1547_0, i_8_471_1555_0,
    i_8_471_1561_0, i_8_471_1564_0, i_8_471_1602_0, i_8_471_1605_0,
    i_8_471_1611_0, i_8_471_1612_0, i_8_471_1641_0, i_8_471_1679_0,
    i_8_471_1692_0, i_8_471_1696_0, i_8_471_1714_0, i_8_471_1730_0,
    i_8_471_1732_0, i_8_471_1786_0, i_8_471_1790_0, i_8_471_1805_0,
    i_8_471_1809_0, i_8_471_1820_0, i_8_471_1830_0, i_8_471_1938_0,
    i_8_471_1948_0, i_8_471_1981_0, i_8_471_1992_0, i_8_471_1995_0,
    i_8_471_2071_0, i_8_471_2073_0, i_8_471_2092_0, i_8_471_2135_0,
    i_8_471_2142_0, i_8_471_2145_0, i_8_471_2216_0, i_8_471_2223_0,
    i_8_471_2234_0, i_8_471_2242_0, i_8_471_2244_0, i_8_471_2286_0,
    o_8_471_0_0  );
  input  i_8_471_64_0, i_8_471_141_0, i_8_471_165_0, i_8_471_238_0,
    i_8_471_265_0, i_8_471_297_0, i_8_471_334_0, i_8_471_352_0,
    i_8_471_361_0, i_8_471_379_0, i_8_471_399_0, i_8_471_400_0,
    i_8_471_418_0, i_8_471_453_0, i_8_471_481_0, i_8_471_493_0,
    i_8_471_524_0, i_8_471_525_0, i_8_471_526_0, i_8_471_541_0,
    i_8_471_550_0, i_8_471_552_0, i_8_471_553_0, i_8_471_570_0,
    i_8_471_571_0, i_8_471_580_0, i_8_471_589_0, i_8_471_606_0,
    i_8_471_659_0, i_8_471_661_0, i_8_471_662_0, i_8_471_687_0,
    i_8_471_688_0, i_8_471_708_0, i_8_471_760_0, i_8_471_804_0,
    i_8_471_837_0, i_8_471_840_0, i_8_471_874_0, i_8_471_990_0,
    i_8_471_1057_0, i_8_471_1058_0, i_8_471_1111_0, i_8_471_1183_0,
    i_8_471_1200_0, i_8_471_1238_0, i_8_471_1266_0, i_8_471_1267_0,
    i_8_471_1271_0, i_8_471_1288_0, i_8_471_1291_0, i_8_471_1308_0,
    i_8_471_1399_0, i_8_471_1411_0, i_8_471_1416_0, i_8_471_1432_0,
    i_8_471_1437_0, i_8_471_1441_0, i_8_471_1462_0, i_8_471_1515_0,
    i_8_471_1544_0, i_8_471_1546_0, i_8_471_1547_0, i_8_471_1555_0,
    i_8_471_1561_0, i_8_471_1564_0, i_8_471_1602_0, i_8_471_1605_0,
    i_8_471_1611_0, i_8_471_1612_0, i_8_471_1641_0, i_8_471_1679_0,
    i_8_471_1692_0, i_8_471_1696_0, i_8_471_1714_0, i_8_471_1730_0,
    i_8_471_1732_0, i_8_471_1786_0, i_8_471_1790_0, i_8_471_1805_0,
    i_8_471_1809_0, i_8_471_1820_0, i_8_471_1830_0, i_8_471_1938_0,
    i_8_471_1948_0, i_8_471_1981_0, i_8_471_1992_0, i_8_471_1995_0,
    i_8_471_2071_0, i_8_471_2073_0, i_8_471_2092_0, i_8_471_2135_0,
    i_8_471_2142_0, i_8_471_2145_0, i_8_471_2216_0, i_8_471_2223_0,
    i_8_471_2234_0, i_8_471_2242_0, i_8_471_2244_0, i_8_471_2286_0;
  output o_8_471_0_0;
  assign o_8_471_0_0 = 0;
endmodule



// Benchmark "kernel_8_472" written by ABC on Sun Jul 19 10:11:23 2020

module kernel_8_472 ( 
    i_8_472_96_0, i_8_472_111_0, i_8_472_114_0, i_8_472_137_0,
    i_8_472_189_0, i_8_472_190_0, i_8_472_193_0, i_8_472_204_0,
    i_8_472_211_0, i_8_472_220_0, i_8_472_258_0, i_8_472_259_0,
    i_8_472_330_0, i_8_472_363_0, i_8_472_382_0, i_8_472_393_0,
    i_8_472_394_0, i_8_472_427_0, i_8_472_440_0, i_8_472_447_0,
    i_8_472_456_0, i_8_472_492_0, i_8_472_495_0, i_8_472_510_0,
    i_8_472_511_0, i_8_472_556_0, i_8_472_601_0, i_8_472_609_0,
    i_8_472_610_0, i_8_472_631_0, i_8_472_659_0, i_8_472_673_0,
    i_8_472_706_0, i_8_472_726_0, i_8_472_750_0, i_8_472_789_0,
    i_8_472_813_0, i_8_472_856_0, i_8_472_876_0, i_8_472_889_0,
    i_8_472_933_0, i_8_472_934_0, i_8_472_958_0, i_8_472_987_0,
    i_8_472_994_0, i_8_472_1029_0, i_8_472_1052_0, i_8_472_1074_0,
    i_8_472_1087_0, i_8_472_1113_0, i_8_472_1114_0, i_8_472_1124_0,
    i_8_472_1221_0, i_8_472_1273_0, i_8_472_1281_0, i_8_472_1282_0,
    i_8_472_1285_0, i_8_472_1301_0, i_8_472_1305_0, i_8_472_1308_0,
    i_8_472_1331_0, i_8_472_1390_0, i_8_472_1410_0, i_8_472_1435_0,
    i_8_472_1439_0, i_8_472_1473_0, i_8_472_1493_0, i_8_472_1536_0,
    i_8_472_1542_0, i_8_472_1573_0, i_8_472_1599_0, i_8_472_1617_0,
    i_8_472_1635_0, i_8_472_1651_0, i_8_472_1653_0, i_8_472_1669_0,
    i_8_472_1678_0, i_8_472_1679_0, i_8_472_1681_0, i_8_472_1698_0,
    i_8_472_1710_0, i_8_472_1725_0, i_8_472_1740_0, i_8_472_1763_0,
    i_8_472_1851_0, i_8_472_1857_0, i_8_472_1879_0, i_8_472_1905_0,
    i_8_472_1906_0, i_8_472_1986_0, i_8_472_1987_0, i_8_472_1996_0,
    i_8_472_2031_0, i_8_472_2037_0, i_8_472_2058_0, i_8_472_2059_0,
    i_8_472_2107_0, i_8_472_2155_0, i_8_472_2217_0, i_8_472_2283_0,
    o_8_472_0_0  );
  input  i_8_472_96_0, i_8_472_111_0, i_8_472_114_0, i_8_472_137_0,
    i_8_472_189_0, i_8_472_190_0, i_8_472_193_0, i_8_472_204_0,
    i_8_472_211_0, i_8_472_220_0, i_8_472_258_0, i_8_472_259_0,
    i_8_472_330_0, i_8_472_363_0, i_8_472_382_0, i_8_472_393_0,
    i_8_472_394_0, i_8_472_427_0, i_8_472_440_0, i_8_472_447_0,
    i_8_472_456_0, i_8_472_492_0, i_8_472_495_0, i_8_472_510_0,
    i_8_472_511_0, i_8_472_556_0, i_8_472_601_0, i_8_472_609_0,
    i_8_472_610_0, i_8_472_631_0, i_8_472_659_0, i_8_472_673_0,
    i_8_472_706_0, i_8_472_726_0, i_8_472_750_0, i_8_472_789_0,
    i_8_472_813_0, i_8_472_856_0, i_8_472_876_0, i_8_472_889_0,
    i_8_472_933_0, i_8_472_934_0, i_8_472_958_0, i_8_472_987_0,
    i_8_472_994_0, i_8_472_1029_0, i_8_472_1052_0, i_8_472_1074_0,
    i_8_472_1087_0, i_8_472_1113_0, i_8_472_1114_0, i_8_472_1124_0,
    i_8_472_1221_0, i_8_472_1273_0, i_8_472_1281_0, i_8_472_1282_0,
    i_8_472_1285_0, i_8_472_1301_0, i_8_472_1305_0, i_8_472_1308_0,
    i_8_472_1331_0, i_8_472_1390_0, i_8_472_1410_0, i_8_472_1435_0,
    i_8_472_1439_0, i_8_472_1473_0, i_8_472_1493_0, i_8_472_1536_0,
    i_8_472_1542_0, i_8_472_1573_0, i_8_472_1599_0, i_8_472_1617_0,
    i_8_472_1635_0, i_8_472_1651_0, i_8_472_1653_0, i_8_472_1669_0,
    i_8_472_1678_0, i_8_472_1679_0, i_8_472_1681_0, i_8_472_1698_0,
    i_8_472_1710_0, i_8_472_1725_0, i_8_472_1740_0, i_8_472_1763_0,
    i_8_472_1851_0, i_8_472_1857_0, i_8_472_1879_0, i_8_472_1905_0,
    i_8_472_1906_0, i_8_472_1986_0, i_8_472_1987_0, i_8_472_1996_0,
    i_8_472_2031_0, i_8_472_2037_0, i_8_472_2058_0, i_8_472_2059_0,
    i_8_472_2107_0, i_8_472_2155_0, i_8_472_2217_0, i_8_472_2283_0;
  output o_8_472_0_0;
  assign o_8_472_0_0 = ~((~i_8_472_440_0 & ((~i_8_472_111_0 & ((i_8_472_114_0 & ~i_8_472_190_0 & ~i_8_472_789_0 & ~i_8_472_1087_0 & ~i_8_472_1473_0 & ~i_8_472_1740_0) | (~i_8_472_259_0 & ~i_8_472_726_0 & ~i_8_472_876_0 & ~i_8_472_987_0 & ~i_8_472_1273_0 & ~i_8_472_1635_0 & ~i_8_472_1906_0 & ~i_8_472_2283_0))) | (~i_8_472_1635_0 & ((~i_8_472_726_0 & ((~i_8_472_96_0 & i_8_472_456_0 & ~i_8_472_789_0 & ~i_8_472_1281_0 & ~i_8_472_1331_0 & ~i_8_472_1879_0 & ~i_8_472_2031_0) | (~i_8_472_259_0 & ~i_8_472_813_0 & ~i_8_472_994_0 & ~i_8_472_1435_0 & ~i_8_472_1573_0 & ~i_8_472_1725_0 & ~i_8_472_1763_0 & ~i_8_472_2283_0))) | (~i_8_472_258_0 & i_8_472_1679_0) | (~i_8_472_789_0 & ~i_8_472_813_0 & ~i_8_472_1124_0 & ~i_8_472_1308_0 & ~i_8_472_1435_0 & ~i_8_472_1573_0 & ~i_8_472_1599_0 & ~i_8_472_1617_0 & ~i_8_472_1905_0 & ~i_8_472_2031_0))) | (~i_8_472_813_0 & ((~i_8_472_2031_0 & ((~i_8_472_190_0 & ~i_8_472_193_0 & ~i_8_472_456_0 & ~i_8_472_1124_0 & ~i_8_472_1331_0 & ~i_8_472_1390_0 & ~i_8_472_1573_0 & ~i_8_472_1698_0) | (i_8_472_1281_0 & ~i_8_472_1617_0 & ~i_8_472_2283_0))) | (~i_8_472_394_0 & ~i_8_472_447_0 & ~i_8_472_934_0 & ~i_8_472_987_0 & ~i_8_472_1029_0 & ~i_8_472_1087_0 & ~i_8_472_1599_0 & ~i_8_472_1851_0 & ~i_8_472_1879_0 & ~i_8_472_1905_0 & ~i_8_472_2217_0))))) | (~i_8_472_789_0 & ((~i_8_472_259_0 & ((~i_8_472_96_0 & ~i_8_472_189_0 & ~i_8_472_750_0 & ~i_8_472_1074_0 & ~i_8_472_1542_0 & ~i_8_472_1573_0 & ~i_8_472_1617_0 & ~i_8_472_1635_0 & ~i_8_472_1905_0 & ~i_8_472_1996_0) | (i_8_472_427_0 & ~i_8_472_510_0 & ~i_8_472_2031_0))) | (~i_8_472_1573_0 & ((i_8_472_363_0 & ~i_8_472_447_0 & ~i_8_472_726_0 & ~i_8_472_1074_0) | (~i_8_472_456_0 & ~i_8_472_934_0 & ~i_8_472_1725_0 & i_8_472_1857_0 & ~i_8_472_2031_0 & ~i_8_472_2059_0 & ~i_8_472_2107_0))) | (~i_8_472_601_0 & i_8_472_1282_0 & ~i_8_472_1905_0 & ~i_8_472_1906_0 & ~i_8_472_2107_0))) | (~i_8_472_96_0 & i_8_472_1114_0 & ((~i_8_472_933_0 & ~i_8_472_1390_0 & ~i_8_472_1879_0 & ~i_8_472_1905_0 & ~i_8_472_1906_0 & ~i_8_472_2037_0) | (~i_8_472_1435_0 & ~i_8_472_1857_0 & i_8_472_1996_0 & ~i_8_472_2031_0 & ~i_8_472_2217_0))) | (~i_8_472_189_0 & ((~i_8_472_934_0 & ~i_8_472_987_0 & ~i_8_472_1052_0 & ~i_8_472_1273_0 & i_8_472_1410_0 & ~i_8_472_1536_0) | (~i_8_472_211_0 & ~i_8_472_456_0 & ~i_8_472_726_0 & ~i_8_472_933_0 & ~i_8_472_994_0 & i_8_472_1536_0 & ~i_8_472_1879_0))) | (i_8_472_427_0 & ((i_8_472_447_0 & ~i_8_472_726_0 & ~i_8_472_856_0 & ~i_8_472_1281_0 & ~i_8_472_1573_0 & i_8_472_1635_0 & ~i_8_472_1710_0 & ~i_8_472_1740_0) | (~i_8_472_204_0 & ~i_8_472_601_0 & ~i_8_472_631_0 & i_8_472_706_0 & ~i_8_472_889_0 & ~i_8_472_1681_0 & ~i_8_472_2217_0))) | (~i_8_472_933_0 & ((~i_8_472_673_0 & ((i_8_472_556_0 & ~i_8_472_601_0 & ~i_8_472_726_0 & ~i_8_472_2031_0) | (~i_8_472_1698_0 & ~i_8_472_1725_0 & ~i_8_472_1851_0 & i_8_472_2058_0))) | (~i_8_472_510_0 & ~i_8_472_726_0 & i_8_472_889_0 & ~i_8_472_994_0 & ~i_8_472_1087_0 & ~i_8_472_1617_0))) | (~i_8_472_258_0 & ~i_8_472_447_0 & ~i_8_472_726_0 & ~i_8_472_813_0 & ~i_8_472_934_0 & i_8_472_1435_0 & ~i_8_472_1599_0 & ~i_8_472_1906_0) | (~i_8_472_456_0 & ~i_8_472_958_0 & ~i_8_472_1635_0 & i_8_472_1986_0 & ~i_8_472_2107_0) | (i_8_472_220_0 & ~i_8_472_393_0 & ~i_8_472_659_0 & ~i_8_472_994_0 & ~i_8_472_1029_0 & ~i_8_472_1439_0 & ~i_8_472_1678_0 & ~i_8_472_1725_0 & ~i_8_472_1740_0 & i_8_472_1996_0 & ~i_8_472_2217_0));
endmodule



// Benchmark "kernel_8_473" written by ABC on Sun Jul 19 10:11:23 2020

module kernel_8_473 ( 
    i_8_473_86_0, i_8_473_88_0, i_8_473_143_0, i_8_473_160_0,
    i_8_473_169_0, i_8_473_170_0, i_8_473_212_0, i_8_473_221_0,
    i_8_473_266_0, i_8_473_269_0, i_8_473_296_0, i_8_473_311_0,
    i_8_473_329_0, i_8_473_440_0, i_8_473_454_0, i_8_473_455_0,
    i_8_473_464_0, i_8_473_481_0, i_8_473_485_0, i_8_473_493_0,
    i_8_473_494_0, i_8_473_502_0, i_8_473_553_0, i_8_473_554_0,
    i_8_473_593_0, i_8_473_606_0, i_8_473_625_0, i_8_473_626_0,
    i_8_473_637_0, i_8_473_661_0, i_8_473_714_0, i_8_473_716_0,
    i_8_473_727_0, i_8_473_769_0, i_8_473_781_0, i_8_473_782_0,
    i_8_473_787_0, i_8_473_833_0, i_8_473_836_0, i_8_473_844_0,
    i_8_473_854_0, i_8_473_872_0, i_8_473_881_0, i_8_473_896_0,
    i_8_473_949_0, i_8_473_977_0, i_8_473_995_0, i_8_473_1013_0,
    i_8_473_1067_0, i_8_473_1087_0, i_8_473_1112_0, i_8_473_1114_0,
    i_8_473_1159_0, i_8_473_1160_0, i_8_473_1228_0, i_8_473_1229_0,
    i_8_473_1250_0, i_8_473_1336_0, i_8_473_1346_0, i_8_473_1358_0,
    i_8_473_1401_0, i_8_473_1421_0, i_8_473_1439_0, i_8_473_1444_0,
    i_8_473_1451_0, i_8_473_1526_0, i_8_473_1546_0, i_8_473_1563_0,
    i_8_473_1579_0, i_8_473_1580_0, i_8_473_1598_0, i_8_473_1616_0,
    i_8_473_1625_0, i_8_473_1637_0, i_8_473_1670_0, i_8_473_1679_0,
    i_8_473_1700_0, i_8_473_1732_0, i_8_473_1750_0, i_8_473_1762_0,
    i_8_473_1805_0, i_8_473_1825_0, i_8_473_1840_0, i_8_473_1859_0,
    i_8_473_1862_0, i_8_473_1868_0, i_8_473_1965_0, i_8_473_2002_0,
    i_8_473_2003_0, i_8_473_2030_0, i_8_473_2032_0, i_8_473_2051_0,
    i_8_473_2132_0, i_8_473_2141_0, i_8_473_2148_0, i_8_473_2150_0,
    i_8_473_2151_0, i_8_473_2170_0, i_8_473_2223_0, i_8_473_2290_0,
    o_8_473_0_0  );
  input  i_8_473_86_0, i_8_473_88_0, i_8_473_143_0, i_8_473_160_0,
    i_8_473_169_0, i_8_473_170_0, i_8_473_212_0, i_8_473_221_0,
    i_8_473_266_0, i_8_473_269_0, i_8_473_296_0, i_8_473_311_0,
    i_8_473_329_0, i_8_473_440_0, i_8_473_454_0, i_8_473_455_0,
    i_8_473_464_0, i_8_473_481_0, i_8_473_485_0, i_8_473_493_0,
    i_8_473_494_0, i_8_473_502_0, i_8_473_553_0, i_8_473_554_0,
    i_8_473_593_0, i_8_473_606_0, i_8_473_625_0, i_8_473_626_0,
    i_8_473_637_0, i_8_473_661_0, i_8_473_714_0, i_8_473_716_0,
    i_8_473_727_0, i_8_473_769_0, i_8_473_781_0, i_8_473_782_0,
    i_8_473_787_0, i_8_473_833_0, i_8_473_836_0, i_8_473_844_0,
    i_8_473_854_0, i_8_473_872_0, i_8_473_881_0, i_8_473_896_0,
    i_8_473_949_0, i_8_473_977_0, i_8_473_995_0, i_8_473_1013_0,
    i_8_473_1067_0, i_8_473_1087_0, i_8_473_1112_0, i_8_473_1114_0,
    i_8_473_1159_0, i_8_473_1160_0, i_8_473_1228_0, i_8_473_1229_0,
    i_8_473_1250_0, i_8_473_1336_0, i_8_473_1346_0, i_8_473_1358_0,
    i_8_473_1401_0, i_8_473_1421_0, i_8_473_1439_0, i_8_473_1444_0,
    i_8_473_1451_0, i_8_473_1526_0, i_8_473_1546_0, i_8_473_1563_0,
    i_8_473_1579_0, i_8_473_1580_0, i_8_473_1598_0, i_8_473_1616_0,
    i_8_473_1625_0, i_8_473_1637_0, i_8_473_1670_0, i_8_473_1679_0,
    i_8_473_1700_0, i_8_473_1732_0, i_8_473_1750_0, i_8_473_1762_0,
    i_8_473_1805_0, i_8_473_1825_0, i_8_473_1840_0, i_8_473_1859_0,
    i_8_473_1862_0, i_8_473_1868_0, i_8_473_1965_0, i_8_473_2002_0,
    i_8_473_2003_0, i_8_473_2030_0, i_8_473_2032_0, i_8_473_2051_0,
    i_8_473_2132_0, i_8_473_2141_0, i_8_473_2148_0, i_8_473_2150_0,
    i_8_473_2151_0, i_8_473_2170_0, i_8_473_2223_0, i_8_473_2290_0;
  output o_8_473_0_0;
  assign o_8_473_0_0 = 0;
endmodule



// Benchmark "kernel_8_474" written by ABC on Sun Jul 19 10:11:24 2020

module kernel_8_474 ( 
    i_8_474_30_0, i_8_474_72_0, i_8_474_82_0, i_8_474_84_0, i_8_474_104_0,
    i_8_474_147_0, i_8_474_190_0, i_8_474_219_0, i_8_474_368_0,
    i_8_474_382_0, i_8_474_427_0, i_8_474_440_0, i_8_474_441_0,
    i_8_474_550_0, i_8_474_568_0, i_8_474_586_0, i_8_474_606_0,
    i_8_474_641_0, i_8_474_664_0, i_8_474_688_0, i_8_474_692_0,
    i_8_474_700_0, i_8_474_729_0, i_8_474_730_0, i_8_474_732_0,
    i_8_474_749_0, i_8_474_752_0, i_8_474_778_0, i_8_474_794_0,
    i_8_474_802_0, i_8_474_803_0, i_8_474_817_0, i_8_474_823_0,
    i_8_474_829_0, i_8_474_840_0, i_8_474_842_0, i_8_474_864_0,
    i_8_474_896_0, i_8_474_965_0, i_8_474_994_0, i_8_474_1003_0,
    i_8_474_1009_0, i_8_474_1128_0, i_8_474_1129_0, i_8_474_1156_0,
    i_8_474_1190_0, i_8_474_1198_0, i_8_474_1229_0, i_8_474_1233_0,
    i_8_474_1237_0, i_8_474_1261_0, i_8_474_1283_0, i_8_474_1285_0,
    i_8_474_1295_0, i_8_474_1296_0, i_8_474_1327_0, i_8_474_1351_0,
    i_8_474_1359_0, i_8_474_1360_0, i_8_474_1362_0, i_8_474_1397_0,
    i_8_474_1423_0, i_8_474_1432_0, i_8_474_1456_0, i_8_474_1469_0,
    i_8_474_1481_0, i_8_474_1503_0, i_8_474_1506_0, i_8_474_1513_0,
    i_8_474_1526_0, i_8_474_1534_0, i_8_474_1548_0, i_8_474_1550_0,
    i_8_474_1582_0, i_8_474_1672_0, i_8_474_1679_0, i_8_474_1705_0,
    i_8_474_1721_0, i_8_474_1745_0, i_8_474_1765_0, i_8_474_1804_0,
    i_8_474_1819_0, i_8_474_1838_0, i_8_474_1877_0, i_8_474_1894_0,
    i_8_474_1909_0, i_8_474_1910_0, i_8_474_1936_0, i_8_474_1962_0,
    i_8_474_1972_0, i_8_474_1973_0, i_8_474_1992_0, i_8_474_2072_0,
    i_8_474_2147_0, i_8_474_2149_0, i_8_474_2224_0, i_8_474_2225_0,
    i_8_474_2226_0, i_8_474_2273_0, i_8_474_2287_0,
    o_8_474_0_0  );
  input  i_8_474_30_0, i_8_474_72_0, i_8_474_82_0, i_8_474_84_0,
    i_8_474_104_0, i_8_474_147_0, i_8_474_190_0, i_8_474_219_0,
    i_8_474_368_0, i_8_474_382_0, i_8_474_427_0, i_8_474_440_0,
    i_8_474_441_0, i_8_474_550_0, i_8_474_568_0, i_8_474_586_0,
    i_8_474_606_0, i_8_474_641_0, i_8_474_664_0, i_8_474_688_0,
    i_8_474_692_0, i_8_474_700_0, i_8_474_729_0, i_8_474_730_0,
    i_8_474_732_0, i_8_474_749_0, i_8_474_752_0, i_8_474_778_0,
    i_8_474_794_0, i_8_474_802_0, i_8_474_803_0, i_8_474_817_0,
    i_8_474_823_0, i_8_474_829_0, i_8_474_840_0, i_8_474_842_0,
    i_8_474_864_0, i_8_474_896_0, i_8_474_965_0, i_8_474_994_0,
    i_8_474_1003_0, i_8_474_1009_0, i_8_474_1128_0, i_8_474_1129_0,
    i_8_474_1156_0, i_8_474_1190_0, i_8_474_1198_0, i_8_474_1229_0,
    i_8_474_1233_0, i_8_474_1237_0, i_8_474_1261_0, i_8_474_1283_0,
    i_8_474_1285_0, i_8_474_1295_0, i_8_474_1296_0, i_8_474_1327_0,
    i_8_474_1351_0, i_8_474_1359_0, i_8_474_1360_0, i_8_474_1362_0,
    i_8_474_1397_0, i_8_474_1423_0, i_8_474_1432_0, i_8_474_1456_0,
    i_8_474_1469_0, i_8_474_1481_0, i_8_474_1503_0, i_8_474_1506_0,
    i_8_474_1513_0, i_8_474_1526_0, i_8_474_1534_0, i_8_474_1548_0,
    i_8_474_1550_0, i_8_474_1582_0, i_8_474_1672_0, i_8_474_1679_0,
    i_8_474_1705_0, i_8_474_1721_0, i_8_474_1745_0, i_8_474_1765_0,
    i_8_474_1804_0, i_8_474_1819_0, i_8_474_1838_0, i_8_474_1877_0,
    i_8_474_1894_0, i_8_474_1909_0, i_8_474_1910_0, i_8_474_1936_0,
    i_8_474_1962_0, i_8_474_1972_0, i_8_474_1973_0, i_8_474_1992_0,
    i_8_474_2072_0, i_8_474_2147_0, i_8_474_2149_0, i_8_474_2224_0,
    i_8_474_2225_0, i_8_474_2226_0, i_8_474_2273_0, i_8_474_2287_0;
  output o_8_474_0_0;
  assign o_8_474_0_0 = 0;
endmodule



// Benchmark "kernel_8_475" written by ABC on Sun Jul 19 10:11:25 2020

module kernel_8_475 ( 
    i_8_475_31_0, i_8_475_49_0, i_8_475_56_0, i_8_475_104_0, i_8_475_117_0,
    i_8_475_125_0, i_8_475_169_0, i_8_475_188_0, i_8_475_198_0,
    i_8_475_230_0, i_8_475_418_0, i_8_475_423_0, i_8_475_490_0,
    i_8_475_496_0, i_8_475_511_0, i_8_475_523_0, i_8_475_524_0,
    i_8_475_527_0, i_8_475_556_0, i_8_475_590_0, i_8_475_608_0,
    i_8_475_610_0, i_8_475_625_0, i_8_475_631_0, i_8_475_637_0,
    i_8_475_659_0, i_8_475_664_0, i_8_475_698_0, i_8_475_699_0,
    i_8_475_710_0, i_8_475_742_0, i_8_475_747_0, i_8_475_772_0,
    i_8_475_786_0, i_8_475_789_0, i_8_475_790_0, i_8_475_850_0,
    i_8_475_857_0, i_8_475_963_0, i_8_475_966_0, i_8_475_971_0,
    i_8_475_1043_0, i_8_475_1059_0, i_8_475_1067_0, i_8_475_1078_0,
    i_8_475_1139_0, i_8_475_1148_0, i_8_475_1160_0, i_8_475_1197_0,
    i_8_475_1214_0, i_8_475_1233_0, i_8_475_1250_0, i_8_475_1251_0,
    i_8_475_1279_0, i_8_475_1306_0, i_8_475_1328_0, i_8_475_1354_0,
    i_8_475_1358_0, i_8_475_1359_0, i_8_475_1426_0, i_8_475_1432_0,
    i_8_475_1485_0, i_8_475_1490_0, i_8_475_1525_0, i_8_475_1543_0,
    i_8_475_1544_0, i_8_475_1547_0, i_8_475_1552_0, i_8_475_1630_0,
    i_8_475_1636_0, i_8_475_1669_0, i_8_475_1674_0, i_8_475_1680_0,
    i_8_475_1681_0, i_8_475_1682_0, i_8_475_1753_0, i_8_475_1764_0,
    i_8_475_1778_0, i_8_475_1790_0, i_8_475_1795_0, i_8_475_1801_0,
    i_8_475_1818_0, i_8_475_1822_0, i_8_475_1837_0, i_8_475_1849_0,
    i_8_475_1851_0, i_8_475_1888_0, i_8_475_1960_0, i_8_475_2057_0,
    i_8_475_2105_0, i_8_475_2125_0, i_8_475_2149_0, i_8_475_2150_0,
    i_8_475_2161_0, i_8_475_2227_0, i_8_475_2229_0, i_8_475_2242_0,
    i_8_475_2246_0, i_8_475_2254_0, i_8_475_2278_0,
    o_8_475_0_0  );
  input  i_8_475_31_0, i_8_475_49_0, i_8_475_56_0, i_8_475_104_0,
    i_8_475_117_0, i_8_475_125_0, i_8_475_169_0, i_8_475_188_0,
    i_8_475_198_0, i_8_475_230_0, i_8_475_418_0, i_8_475_423_0,
    i_8_475_490_0, i_8_475_496_0, i_8_475_511_0, i_8_475_523_0,
    i_8_475_524_0, i_8_475_527_0, i_8_475_556_0, i_8_475_590_0,
    i_8_475_608_0, i_8_475_610_0, i_8_475_625_0, i_8_475_631_0,
    i_8_475_637_0, i_8_475_659_0, i_8_475_664_0, i_8_475_698_0,
    i_8_475_699_0, i_8_475_710_0, i_8_475_742_0, i_8_475_747_0,
    i_8_475_772_0, i_8_475_786_0, i_8_475_789_0, i_8_475_790_0,
    i_8_475_850_0, i_8_475_857_0, i_8_475_963_0, i_8_475_966_0,
    i_8_475_971_0, i_8_475_1043_0, i_8_475_1059_0, i_8_475_1067_0,
    i_8_475_1078_0, i_8_475_1139_0, i_8_475_1148_0, i_8_475_1160_0,
    i_8_475_1197_0, i_8_475_1214_0, i_8_475_1233_0, i_8_475_1250_0,
    i_8_475_1251_0, i_8_475_1279_0, i_8_475_1306_0, i_8_475_1328_0,
    i_8_475_1354_0, i_8_475_1358_0, i_8_475_1359_0, i_8_475_1426_0,
    i_8_475_1432_0, i_8_475_1485_0, i_8_475_1490_0, i_8_475_1525_0,
    i_8_475_1543_0, i_8_475_1544_0, i_8_475_1547_0, i_8_475_1552_0,
    i_8_475_1630_0, i_8_475_1636_0, i_8_475_1669_0, i_8_475_1674_0,
    i_8_475_1680_0, i_8_475_1681_0, i_8_475_1682_0, i_8_475_1753_0,
    i_8_475_1764_0, i_8_475_1778_0, i_8_475_1790_0, i_8_475_1795_0,
    i_8_475_1801_0, i_8_475_1818_0, i_8_475_1822_0, i_8_475_1837_0,
    i_8_475_1849_0, i_8_475_1851_0, i_8_475_1888_0, i_8_475_1960_0,
    i_8_475_2057_0, i_8_475_2105_0, i_8_475_2125_0, i_8_475_2149_0,
    i_8_475_2150_0, i_8_475_2161_0, i_8_475_2227_0, i_8_475_2229_0,
    i_8_475_2242_0, i_8_475_2246_0, i_8_475_2254_0, i_8_475_2278_0;
  output o_8_475_0_0;
  assign o_8_475_0_0 = 0;
endmodule



// Benchmark "kernel_8_476" written by ABC on Sun Jul 19 10:11:27 2020

module kernel_8_476 ( 
    i_8_476_16_0, i_8_476_24_0, i_8_476_25_0, i_8_476_26_0, i_8_476_43_0,
    i_8_476_52_0, i_8_476_77_0, i_8_476_88_0, i_8_476_176_0, i_8_476_177_0,
    i_8_476_178_0, i_8_476_204_0, i_8_476_276_0, i_8_476_277_0,
    i_8_476_286_0, i_8_476_303_0, i_8_476_314_0, i_8_476_328_0,
    i_8_476_329_0, i_8_476_339_0, i_8_476_348_0, i_8_476_354_0,
    i_8_476_357_0, i_8_476_358_0, i_8_476_359_0, i_8_476_363_0,
    i_8_476_368_0, i_8_476_370_0, i_8_476_384_0, i_8_476_385_0,
    i_8_476_458_0, i_8_476_484_0, i_8_476_492_0, i_8_476_499_0,
    i_8_476_519_0, i_8_476_574_0, i_8_476_575_0, i_8_476_601_0,
    i_8_476_611_0, i_8_476_618_0, i_8_476_628_0, i_8_476_629_0,
    i_8_476_699_0, i_8_476_701_0, i_8_476_708_0, i_8_476_709_0,
    i_8_476_856_0, i_8_476_863_0, i_8_476_958_0, i_8_476_961_0,
    i_8_476_1015_0, i_8_476_1033_0, i_8_476_1040_0, i_8_476_1042_0,
    i_8_476_1096_0, i_8_476_1112_0, i_8_476_1176_0, i_8_476_1177_0,
    i_8_476_1178_0, i_8_476_1195_0, i_8_476_1231_0, i_8_476_1232_0,
    i_8_476_1274_0, i_8_476_1293_0, i_8_476_1294_0, i_8_476_1295_0,
    i_8_476_1309_0, i_8_476_1363_0, i_8_476_1365_0, i_8_476_1366_0,
    i_8_476_1367_0, i_8_476_1457_0, i_8_476_1474_0, i_8_476_1475_0,
    i_8_476_1564_0, i_8_476_1565_0, i_8_476_1590_0, i_8_476_1603_0,
    i_8_476_1709_0, i_8_476_1725_0, i_8_476_1726_0, i_8_476_1727_0,
    i_8_476_1761_0, i_8_476_1770_0, i_8_476_1771_0, i_8_476_1776_0,
    i_8_476_1825_0, i_8_476_1861_0, i_8_476_1921_0, i_8_476_2052_0,
    i_8_476_2067_0, i_8_476_2113_0, i_8_476_2157_0, i_8_476_2158_0,
    i_8_476_2194_0, i_8_476_2213_0, i_8_476_2219_0, i_8_476_2229_0,
    i_8_476_2239_0, i_8_476_2245_0,
    o_8_476_0_0  );
  input  i_8_476_16_0, i_8_476_24_0, i_8_476_25_0, i_8_476_26_0,
    i_8_476_43_0, i_8_476_52_0, i_8_476_77_0, i_8_476_88_0, i_8_476_176_0,
    i_8_476_177_0, i_8_476_178_0, i_8_476_204_0, i_8_476_276_0,
    i_8_476_277_0, i_8_476_286_0, i_8_476_303_0, i_8_476_314_0,
    i_8_476_328_0, i_8_476_329_0, i_8_476_339_0, i_8_476_348_0,
    i_8_476_354_0, i_8_476_357_0, i_8_476_358_0, i_8_476_359_0,
    i_8_476_363_0, i_8_476_368_0, i_8_476_370_0, i_8_476_384_0,
    i_8_476_385_0, i_8_476_458_0, i_8_476_484_0, i_8_476_492_0,
    i_8_476_499_0, i_8_476_519_0, i_8_476_574_0, i_8_476_575_0,
    i_8_476_601_0, i_8_476_611_0, i_8_476_618_0, i_8_476_628_0,
    i_8_476_629_0, i_8_476_699_0, i_8_476_701_0, i_8_476_708_0,
    i_8_476_709_0, i_8_476_856_0, i_8_476_863_0, i_8_476_958_0,
    i_8_476_961_0, i_8_476_1015_0, i_8_476_1033_0, i_8_476_1040_0,
    i_8_476_1042_0, i_8_476_1096_0, i_8_476_1112_0, i_8_476_1176_0,
    i_8_476_1177_0, i_8_476_1178_0, i_8_476_1195_0, i_8_476_1231_0,
    i_8_476_1232_0, i_8_476_1274_0, i_8_476_1293_0, i_8_476_1294_0,
    i_8_476_1295_0, i_8_476_1309_0, i_8_476_1363_0, i_8_476_1365_0,
    i_8_476_1366_0, i_8_476_1367_0, i_8_476_1457_0, i_8_476_1474_0,
    i_8_476_1475_0, i_8_476_1564_0, i_8_476_1565_0, i_8_476_1590_0,
    i_8_476_1603_0, i_8_476_1709_0, i_8_476_1725_0, i_8_476_1726_0,
    i_8_476_1727_0, i_8_476_1761_0, i_8_476_1770_0, i_8_476_1771_0,
    i_8_476_1776_0, i_8_476_1825_0, i_8_476_1861_0, i_8_476_1921_0,
    i_8_476_2052_0, i_8_476_2067_0, i_8_476_2113_0, i_8_476_2157_0,
    i_8_476_2158_0, i_8_476_2194_0, i_8_476_2213_0, i_8_476_2219_0,
    i_8_476_2229_0, i_8_476_2239_0, i_8_476_2245_0;
  output o_8_476_0_0;
  assign o_8_476_0_0 = ~((~i_8_476_24_0 & ((~i_8_476_354_0 & ~i_8_476_1096_0 & ~i_8_476_1195_0 & ~i_8_476_1295_0 & ~i_8_476_1309_0 & ~i_8_476_2067_0 & ~i_8_476_2113_0 & ~i_8_476_2158_0) | (~i_8_476_52_0 & i_8_476_77_0 & ~i_8_476_176_0 & ~i_8_476_958_0 & i_8_476_1112_0 & ~i_8_476_1177_0 & ~i_8_476_1274_0 & ~i_8_476_1457_0 & ~i_8_476_2213_0))) | (~i_8_476_25_0 & ((~i_8_476_26_0 & ~i_8_476_519_0 & i_8_476_601_0 & ~i_8_476_1176_0 & ~i_8_476_1295_0 & ~i_8_476_2113_0 & ~i_8_476_2219_0) | (i_8_476_1015_0 & ~i_8_476_1474_0 & ~i_8_476_1564_0 & ~i_8_476_2239_0))) | (~i_8_476_26_0 & ((~i_8_476_178_0 & ((~i_8_476_384_0 & ~i_8_476_499_0 & ~i_8_476_1015_0 & ~i_8_476_1096_0 & ~i_8_476_1274_0 & ~i_8_476_1293_0 & ~i_8_476_1295_0 & ~i_8_476_1709_0 & ~i_8_476_2158_0) | (i_8_476_328_0 & ~i_8_476_357_0 & i_8_476_385_0 & ~i_8_476_1294_0 & ~i_8_476_1366_0 & ~i_8_476_2219_0))) | (~i_8_476_204_0 & ~i_8_476_2113_0 & ((~i_8_476_314_0 & i_8_476_458_0) | (~i_8_476_77_0 & ~i_8_476_177_0 & ~i_8_476_359_0 & ~i_8_476_629_0 & ~i_8_476_961_0 & ~i_8_476_1195_0 & ~i_8_476_1294_0))) | (~i_8_476_385_0 & ~i_8_476_458_0 & ~i_8_476_699_0 & ~i_8_476_863_0 & ~i_8_476_1564_0 & ~i_8_476_1825_0 & ~i_8_476_2158_0 & ~i_8_476_2239_0))) | (~i_8_476_176_0 & ((~i_8_476_277_0 & ((~i_8_476_43_0 & ~i_8_476_314_0 & ~i_8_476_708_0 & ~i_8_476_1294_0 & ~i_8_476_1921_0) | (~i_8_476_177_0 & ~i_8_476_178_0 & ~i_8_476_357_0 & ~i_8_476_358_0 & ~i_8_476_384_0 & ~i_8_476_863_0 & ~i_8_476_1176_0 & ~i_8_476_1232_0 & i_8_476_2113_0))) | (~i_8_476_16_0 & ~i_8_476_276_0 & i_8_476_368_0 & ~i_8_476_575_0 & ~i_8_476_1177_0 & ~i_8_476_1474_0 & ~i_8_476_1475_0 & ~i_8_476_1603_0 & ~i_8_476_1776_0 & ~i_8_476_2052_0))) | (~i_8_476_177_0 & ~i_8_476_178_0 & ((~i_8_476_43_0 & ~i_8_476_357_0 & i_8_476_363_0 & ~i_8_476_368_0 & ~i_8_476_519_0) | (~i_8_476_499_0 & ~i_8_476_708_0 & ~i_8_476_863_0 & ~i_8_476_958_0 & ~i_8_476_1295_0 & ~i_8_476_2157_0 & ~i_8_476_2219_0 & ~i_8_476_2239_0))) | (~i_8_476_1178_0 & ((~i_8_476_1176_0 & ((~i_8_476_43_0 & ((~i_8_476_314_0 & ~i_8_476_575_0 & ~i_8_476_1294_0 & i_8_476_1474_0 & ~i_8_476_1564_0 & ~i_8_476_1761_0 & ~i_8_476_1861_0) | (~i_8_476_492_0 & ~i_8_476_1231_0 & ~i_8_476_1232_0 & ~i_8_476_2113_0 & ~i_8_476_2229_0))) | (~i_8_476_88_0 & ~i_8_476_276_0 & ~i_8_476_358_0 & ~i_8_476_1177_0 & ~i_8_476_2113_0 & ~i_8_476_2229_0 & ~i_8_476_1294_0 & ~i_8_476_1474_0))) | (i_8_476_303_0 & ~i_8_476_699_0 & ~i_8_476_701_0) | (~i_8_476_618_0 & ~i_8_476_1177_0 & ~i_8_476_1232_0 & ~i_8_476_1293_0 & ~i_8_476_1474_0 & ~i_8_476_2239_0))) | (~i_8_476_359_0 & ((i_8_476_368_0 & ~i_8_476_958_0 & ~i_8_476_1112_0 & i_8_476_1232_0 & ~i_8_476_1475_0 & i_8_476_1825_0) | (~i_8_476_276_0 & ~i_8_476_709_0 & ~i_8_476_1232_0 & ~i_8_476_1825_0 & ~i_8_476_2239_0))) | (i_8_476_88_0 & i_8_476_1727_0 & i_8_476_1861_0) | (~i_8_476_492_0 & i_8_476_701_0 & ~i_8_476_1112_0 & ~i_8_476_1231_0 & ~i_8_476_1603_0 & ~i_8_476_1709_0 & ~i_8_476_1921_0));
endmodule



// Benchmark "kernel_8_477" written by ABC on Sun Jul 19 10:11:28 2020

module kernel_8_477 ( 
    i_8_477_10_0, i_8_477_18_0, i_8_477_31_0, i_8_477_64_0, i_8_477_65_0,
    i_8_477_68_0, i_8_477_112_0, i_8_477_117_0, i_8_477_118_0,
    i_8_477_195_0, i_8_477_221_0, i_8_477_224_0, i_8_477_227_0,
    i_8_477_307_0, i_8_477_317_0, i_8_477_320_0, i_8_477_346_0,
    i_8_477_362_0, i_8_477_364_0, i_8_477_373_0, i_8_477_418_0,
    i_8_477_419_0, i_8_477_505_0, i_8_477_506_0, i_8_477_551_0,
    i_8_477_590_0, i_8_477_605_0, i_8_477_632_0, i_8_477_635_0,
    i_8_477_640_0, i_8_477_641_0, i_8_477_649_0, i_8_477_707_0,
    i_8_477_735_0, i_8_477_749_0, i_8_477_811_0, i_8_477_829_0,
    i_8_477_838_0, i_8_477_839_0, i_8_477_841_0, i_8_477_846_0,
    i_8_477_847_0, i_8_477_974_0, i_8_477_991_0, i_8_477_1035_0,
    i_8_477_1048_0, i_8_477_1071_0, i_8_477_1081_0, i_8_477_1109_0,
    i_8_477_1134_0, i_8_477_1135_0, i_8_477_1161_0, i_8_477_1215_0,
    i_8_477_1229_0, i_8_477_1296_0, i_8_477_1325_0, i_8_477_1360_0,
    i_8_477_1382_0, i_8_477_1387_0, i_8_477_1423_0, i_8_477_1424_0,
    i_8_477_1436_0, i_8_477_1460_0, i_8_477_1462_0, i_8_477_1463_0,
    i_8_477_1471_0, i_8_477_1507_0, i_8_477_1514_0, i_8_477_1522_0,
    i_8_477_1539_0, i_8_477_1570_0, i_8_477_1571_0, i_8_477_1634_0,
    i_8_477_1694_0, i_8_477_1703_0, i_8_477_1775_0, i_8_477_1781_0,
    i_8_477_1838_0, i_8_477_1886_0, i_8_477_1887_0, i_8_477_1888_0,
    i_8_477_1955_0, i_8_477_1957_0, i_8_477_1970_0, i_8_477_1973_0,
    i_8_477_1976_0, i_8_477_1982_0, i_8_477_1991_0, i_8_477_2011_0,
    i_8_477_2052_0, i_8_477_2089_0, i_8_477_2090_0, i_8_477_2097_0,
    i_8_477_2098_0, i_8_477_2135_0, i_8_477_2188_0, i_8_477_2224_0,
    i_8_477_2252_0, i_8_477_2255_0, i_8_477_2269_0,
    o_8_477_0_0  );
  input  i_8_477_10_0, i_8_477_18_0, i_8_477_31_0, i_8_477_64_0,
    i_8_477_65_0, i_8_477_68_0, i_8_477_112_0, i_8_477_117_0,
    i_8_477_118_0, i_8_477_195_0, i_8_477_221_0, i_8_477_224_0,
    i_8_477_227_0, i_8_477_307_0, i_8_477_317_0, i_8_477_320_0,
    i_8_477_346_0, i_8_477_362_0, i_8_477_364_0, i_8_477_373_0,
    i_8_477_418_0, i_8_477_419_0, i_8_477_505_0, i_8_477_506_0,
    i_8_477_551_0, i_8_477_590_0, i_8_477_605_0, i_8_477_632_0,
    i_8_477_635_0, i_8_477_640_0, i_8_477_641_0, i_8_477_649_0,
    i_8_477_707_0, i_8_477_735_0, i_8_477_749_0, i_8_477_811_0,
    i_8_477_829_0, i_8_477_838_0, i_8_477_839_0, i_8_477_841_0,
    i_8_477_846_0, i_8_477_847_0, i_8_477_974_0, i_8_477_991_0,
    i_8_477_1035_0, i_8_477_1048_0, i_8_477_1071_0, i_8_477_1081_0,
    i_8_477_1109_0, i_8_477_1134_0, i_8_477_1135_0, i_8_477_1161_0,
    i_8_477_1215_0, i_8_477_1229_0, i_8_477_1296_0, i_8_477_1325_0,
    i_8_477_1360_0, i_8_477_1382_0, i_8_477_1387_0, i_8_477_1423_0,
    i_8_477_1424_0, i_8_477_1436_0, i_8_477_1460_0, i_8_477_1462_0,
    i_8_477_1463_0, i_8_477_1471_0, i_8_477_1507_0, i_8_477_1514_0,
    i_8_477_1522_0, i_8_477_1539_0, i_8_477_1570_0, i_8_477_1571_0,
    i_8_477_1634_0, i_8_477_1694_0, i_8_477_1703_0, i_8_477_1775_0,
    i_8_477_1781_0, i_8_477_1838_0, i_8_477_1886_0, i_8_477_1887_0,
    i_8_477_1888_0, i_8_477_1955_0, i_8_477_1957_0, i_8_477_1970_0,
    i_8_477_1973_0, i_8_477_1976_0, i_8_477_1982_0, i_8_477_1991_0,
    i_8_477_2011_0, i_8_477_2052_0, i_8_477_2089_0, i_8_477_2090_0,
    i_8_477_2097_0, i_8_477_2098_0, i_8_477_2135_0, i_8_477_2188_0,
    i_8_477_2224_0, i_8_477_2252_0, i_8_477_2255_0, i_8_477_2269_0;
  output o_8_477_0_0;
  assign o_8_477_0_0 = 0;
endmodule



// Benchmark "kernel_8_478" written by ABC on Sun Jul 19 10:11:29 2020

module kernel_8_478 ( 
    i_8_478_18_0, i_8_478_21_0, i_8_478_22_0, i_8_478_27_0, i_8_478_30_0,
    i_8_478_31_0, i_8_478_32_0, i_8_478_54_0, i_8_478_57_0, i_8_478_99_0,
    i_8_478_100_0, i_8_478_141_0, i_8_478_201_0, i_8_478_202_0,
    i_8_478_216_0, i_8_478_255_0, i_8_478_262_0, i_8_478_298_0,
    i_8_478_300_0, i_8_478_318_0, i_8_478_319_0, i_8_478_379_0,
    i_8_478_417_0, i_8_478_418_0, i_8_478_426_0, i_8_478_543_0,
    i_8_478_544_0, i_8_478_555_0, i_8_478_572_0, i_8_478_580_0,
    i_8_478_604_0, i_8_478_630_0, i_8_478_640_0, i_8_478_652_0,
    i_8_478_702_0, i_8_478_707_0, i_8_478_747_0, i_8_478_792_0,
    i_8_478_858_0, i_8_478_859_0, i_8_478_882_0, i_8_478_900_0,
    i_8_478_936_0, i_8_478_937_0, i_8_478_963_0, i_8_478_966_0,
    i_8_478_1035_0, i_8_478_1065_0, i_8_478_1076_0, i_8_478_1161_0,
    i_8_478_1240_0, i_8_478_1315_0, i_8_478_1319_0, i_8_478_1332_0,
    i_8_478_1358_0, i_8_478_1359_0, i_8_478_1360_0, i_8_478_1362_0,
    i_8_478_1395_0, i_8_478_1398_0, i_8_478_1416_0, i_8_478_1462_0,
    i_8_478_1463_0, i_8_478_1467_0, i_8_478_1472_0, i_8_478_1521_0,
    i_8_478_1629_0, i_8_478_1630_0, i_8_478_1674_0, i_8_478_1675_0,
    i_8_478_1676_0, i_8_478_1677_0, i_8_478_1683_0, i_8_478_1710_0,
    i_8_478_1711_0, i_8_478_1713_0, i_8_478_1812_0, i_8_478_1836_0,
    i_8_478_1839_0, i_8_478_1926_0, i_8_478_1927_0, i_8_478_1944_0,
    i_8_478_1945_0, i_8_478_1947_0, i_8_478_1951_0, i_8_478_1962_0,
    i_8_478_1983_0, i_8_478_2008_0, i_8_478_2119_0, i_8_478_2133_0,
    i_8_478_2144_0, i_8_478_2154_0, i_8_478_2157_0, i_8_478_2169_0,
    i_8_478_2196_0, i_8_478_2224_0, i_8_478_2226_0, i_8_478_2232_0,
    i_8_478_2233_0, i_8_478_2259_0,
    o_8_478_0_0  );
  input  i_8_478_18_0, i_8_478_21_0, i_8_478_22_0, i_8_478_27_0,
    i_8_478_30_0, i_8_478_31_0, i_8_478_32_0, i_8_478_54_0, i_8_478_57_0,
    i_8_478_99_0, i_8_478_100_0, i_8_478_141_0, i_8_478_201_0,
    i_8_478_202_0, i_8_478_216_0, i_8_478_255_0, i_8_478_262_0,
    i_8_478_298_0, i_8_478_300_0, i_8_478_318_0, i_8_478_319_0,
    i_8_478_379_0, i_8_478_417_0, i_8_478_418_0, i_8_478_426_0,
    i_8_478_543_0, i_8_478_544_0, i_8_478_555_0, i_8_478_572_0,
    i_8_478_580_0, i_8_478_604_0, i_8_478_630_0, i_8_478_640_0,
    i_8_478_652_0, i_8_478_702_0, i_8_478_707_0, i_8_478_747_0,
    i_8_478_792_0, i_8_478_858_0, i_8_478_859_0, i_8_478_882_0,
    i_8_478_900_0, i_8_478_936_0, i_8_478_937_0, i_8_478_963_0,
    i_8_478_966_0, i_8_478_1035_0, i_8_478_1065_0, i_8_478_1076_0,
    i_8_478_1161_0, i_8_478_1240_0, i_8_478_1315_0, i_8_478_1319_0,
    i_8_478_1332_0, i_8_478_1358_0, i_8_478_1359_0, i_8_478_1360_0,
    i_8_478_1362_0, i_8_478_1395_0, i_8_478_1398_0, i_8_478_1416_0,
    i_8_478_1462_0, i_8_478_1463_0, i_8_478_1467_0, i_8_478_1472_0,
    i_8_478_1521_0, i_8_478_1629_0, i_8_478_1630_0, i_8_478_1674_0,
    i_8_478_1675_0, i_8_478_1676_0, i_8_478_1677_0, i_8_478_1683_0,
    i_8_478_1710_0, i_8_478_1711_0, i_8_478_1713_0, i_8_478_1812_0,
    i_8_478_1836_0, i_8_478_1839_0, i_8_478_1926_0, i_8_478_1927_0,
    i_8_478_1944_0, i_8_478_1945_0, i_8_478_1947_0, i_8_478_1951_0,
    i_8_478_1962_0, i_8_478_1983_0, i_8_478_2008_0, i_8_478_2119_0,
    i_8_478_2133_0, i_8_478_2144_0, i_8_478_2154_0, i_8_478_2157_0,
    i_8_478_2169_0, i_8_478_2196_0, i_8_478_2224_0, i_8_478_2226_0,
    i_8_478_2232_0, i_8_478_2233_0, i_8_478_2259_0;
  output o_8_478_0_0;
  assign o_8_478_0_0 = 0;
endmodule



// Benchmark "kernel_8_479" written by ABC on Sun Jul 19 10:11:29 2020

module kernel_8_479 ( 
    i_8_479_35_0, i_8_479_74_0, i_8_479_89_0, i_8_479_107_0, i_8_479_142_0,
    i_8_479_189_0, i_8_479_190_0, i_8_479_222_0, i_8_479_259_0,
    i_8_479_331_0, i_8_479_379_0, i_8_479_386_0, i_8_479_392_0,
    i_8_479_445_0, i_8_479_457_0, i_8_479_481_0, i_8_479_502_0,
    i_8_479_522_0, i_8_479_555_0, i_8_479_556_0, i_8_479_597_0,
    i_8_479_634_0, i_8_479_645_0, i_8_479_664_0, i_8_479_696_0,
    i_8_479_699_0, i_8_479_706_0, i_8_479_762_0, i_8_479_817_0,
    i_8_479_818_0, i_8_479_826_0, i_8_479_897_0, i_8_479_906_0,
    i_8_479_925_0, i_8_479_943_0, i_8_479_951_0, i_8_479_979_0,
    i_8_479_980_0, i_8_479_987_0, i_8_479_988_0, i_8_479_997_0,
    i_8_479_1012_0, i_8_479_1014_0, i_8_479_1015_0, i_8_479_1029_0,
    i_8_479_1113_0, i_8_479_1122_0, i_8_479_1131_0, i_8_479_1140_0,
    i_8_479_1186_0, i_8_479_1303_0, i_8_479_1308_0, i_8_479_1327_0,
    i_8_479_1330_0, i_8_479_1338_0, i_8_479_1348_0, i_8_479_1350_0,
    i_8_479_1453_0, i_8_479_1455_0, i_8_479_1489_0, i_8_479_1510_0,
    i_8_479_1527_0, i_8_479_1599_0, i_8_479_1608_0, i_8_479_1617_0,
    i_8_479_1618_0, i_8_479_1632_0, i_8_479_1651_0, i_8_479_1673_0,
    i_8_479_1681_0, i_8_479_1686_0, i_8_479_1704_0, i_8_479_1708_0,
    i_8_479_1716_0, i_8_479_1717_0, i_8_479_1732_0, i_8_479_1750_0,
    i_8_479_1812_0, i_8_479_1861_0, i_8_479_1862_0, i_8_479_1869_0,
    i_8_479_1870_0, i_8_479_1876_0, i_8_479_1904_0, i_8_479_1918_0,
    i_8_479_1949_0, i_8_479_1950_0, i_8_479_1981_0, i_8_479_1993_0,
    i_8_479_2001_0, i_8_479_2005_0, i_8_479_2049_0, i_8_479_2090_0,
    i_8_479_2093_0, i_8_479_2107_0, i_8_479_2139_0, i_8_479_2140_0,
    i_8_479_2184_0, i_8_479_2193_0, i_8_479_2265_0,
    o_8_479_0_0  );
  input  i_8_479_35_0, i_8_479_74_0, i_8_479_89_0, i_8_479_107_0,
    i_8_479_142_0, i_8_479_189_0, i_8_479_190_0, i_8_479_222_0,
    i_8_479_259_0, i_8_479_331_0, i_8_479_379_0, i_8_479_386_0,
    i_8_479_392_0, i_8_479_445_0, i_8_479_457_0, i_8_479_481_0,
    i_8_479_502_0, i_8_479_522_0, i_8_479_555_0, i_8_479_556_0,
    i_8_479_597_0, i_8_479_634_0, i_8_479_645_0, i_8_479_664_0,
    i_8_479_696_0, i_8_479_699_0, i_8_479_706_0, i_8_479_762_0,
    i_8_479_817_0, i_8_479_818_0, i_8_479_826_0, i_8_479_897_0,
    i_8_479_906_0, i_8_479_925_0, i_8_479_943_0, i_8_479_951_0,
    i_8_479_979_0, i_8_479_980_0, i_8_479_987_0, i_8_479_988_0,
    i_8_479_997_0, i_8_479_1012_0, i_8_479_1014_0, i_8_479_1015_0,
    i_8_479_1029_0, i_8_479_1113_0, i_8_479_1122_0, i_8_479_1131_0,
    i_8_479_1140_0, i_8_479_1186_0, i_8_479_1303_0, i_8_479_1308_0,
    i_8_479_1327_0, i_8_479_1330_0, i_8_479_1338_0, i_8_479_1348_0,
    i_8_479_1350_0, i_8_479_1453_0, i_8_479_1455_0, i_8_479_1489_0,
    i_8_479_1510_0, i_8_479_1527_0, i_8_479_1599_0, i_8_479_1608_0,
    i_8_479_1617_0, i_8_479_1618_0, i_8_479_1632_0, i_8_479_1651_0,
    i_8_479_1673_0, i_8_479_1681_0, i_8_479_1686_0, i_8_479_1704_0,
    i_8_479_1708_0, i_8_479_1716_0, i_8_479_1717_0, i_8_479_1732_0,
    i_8_479_1750_0, i_8_479_1812_0, i_8_479_1861_0, i_8_479_1862_0,
    i_8_479_1869_0, i_8_479_1870_0, i_8_479_1876_0, i_8_479_1904_0,
    i_8_479_1918_0, i_8_479_1949_0, i_8_479_1950_0, i_8_479_1981_0,
    i_8_479_1993_0, i_8_479_2001_0, i_8_479_2005_0, i_8_479_2049_0,
    i_8_479_2090_0, i_8_479_2093_0, i_8_479_2107_0, i_8_479_2139_0,
    i_8_479_2140_0, i_8_479_2184_0, i_8_479_2193_0, i_8_479_2265_0;
  output o_8_479_0_0;
  assign o_8_479_0_0 = 0;
endmodule



// Benchmark "kernel_8_480" written by ABC on Sun Jul 19 10:11:31 2020

module kernel_8_480 ( 
    i_8_480_13_0, i_8_480_21_0, i_8_480_22_0, i_8_480_58_0, i_8_480_66_0,
    i_8_480_109_0, i_8_480_114_0, i_8_480_138_0, i_8_480_194_0,
    i_8_480_219_0, i_8_480_220_0, i_8_480_279_0, i_8_480_285_0,
    i_8_480_321_0, i_8_480_325_0, i_8_480_328_0, i_8_480_345_0,
    i_8_480_364_0, i_8_480_384_0, i_8_480_396_0, i_8_480_400_0,
    i_8_480_486_0, i_8_480_492_0, i_8_480_527_0, i_8_480_530_0,
    i_8_480_552_0, i_8_480_555_0, i_8_480_573_0, i_8_480_589_0,
    i_8_480_594_0, i_8_480_595_0, i_8_480_606_0, i_8_480_608_0,
    i_8_480_615_0, i_8_480_696_0, i_8_480_777_0, i_8_480_822_0,
    i_8_480_838_0, i_8_480_874_0, i_8_480_877_0, i_8_480_880_0,
    i_8_480_883_0, i_8_480_891_0, i_8_480_894_0, i_8_480_969_0,
    i_8_480_970_0, i_8_480_972_0, i_8_480_1029_0, i_8_480_1036_0,
    i_8_480_1092_0, i_8_480_1111_0, i_8_480_1137_0, i_8_480_1146_0,
    i_8_480_1152_0, i_8_480_1155_0, i_8_480_1197_0, i_8_480_1255_0,
    i_8_480_1263_0, i_8_480_1317_0, i_8_480_1324_0, i_8_480_1336_0,
    i_8_480_1396_0, i_8_480_1400_0, i_8_480_1422_0, i_8_480_1423_0,
    i_8_480_1425_0, i_8_480_1440_0, i_8_480_1443_0, i_8_480_1461_0,
    i_8_480_1462_0, i_8_480_1481_0, i_8_480_1518_0, i_8_480_1524_0,
    i_8_480_1525_0, i_8_480_1548_0, i_8_480_1549_0, i_8_480_1587_0,
    i_8_480_1605_0, i_8_480_1638_0, i_8_480_1639_0, i_8_480_1695_0,
    i_8_480_1722_0, i_8_480_1724_0, i_8_480_1746_0, i_8_480_1783_0,
    i_8_480_1813_0, i_8_480_1839_0, i_8_480_1935_0, i_8_480_1967_0,
    i_8_480_1974_0, i_8_480_1995_0, i_8_480_2011_0, i_8_480_2053_0,
    i_8_480_2060_0, i_8_480_2110_0, i_8_480_2111_0, i_8_480_2232_0,
    i_8_480_2233_0, i_8_480_2247_0, i_8_480_2298_0,
    o_8_480_0_0  );
  input  i_8_480_13_0, i_8_480_21_0, i_8_480_22_0, i_8_480_58_0,
    i_8_480_66_0, i_8_480_109_0, i_8_480_114_0, i_8_480_138_0,
    i_8_480_194_0, i_8_480_219_0, i_8_480_220_0, i_8_480_279_0,
    i_8_480_285_0, i_8_480_321_0, i_8_480_325_0, i_8_480_328_0,
    i_8_480_345_0, i_8_480_364_0, i_8_480_384_0, i_8_480_396_0,
    i_8_480_400_0, i_8_480_486_0, i_8_480_492_0, i_8_480_527_0,
    i_8_480_530_0, i_8_480_552_0, i_8_480_555_0, i_8_480_573_0,
    i_8_480_589_0, i_8_480_594_0, i_8_480_595_0, i_8_480_606_0,
    i_8_480_608_0, i_8_480_615_0, i_8_480_696_0, i_8_480_777_0,
    i_8_480_822_0, i_8_480_838_0, i_8_480_874_0, i_8_480_877_0,
    i_8_480_880_0, i_8_480_883_0, i_8_480_891_0, i_8_480_894_0,
    i_8_480_969_0, i_8_480_970_0, i_8_480_972_0, i_8_480_1029_0,
    i_8_480_1036_0, i_8_480_1092_0, i_8_480_1111_0, i_8_480_1137_0,
    i_8_480_1146_0, i_8_480_1152_0, i_8_480_1155_0, i_8_480_1197_0,
    i_8_480_1255_0, i_8_480_1263_0, i_8_480_1317_0, i_8_480_1324_0,
    i_8_480_1336_0, i_8_480_1396_0, i_8_480_1400_0, i_8_480_1422_0,
    i_8_480_1423_0, i_8_480_1425_0, i_8_480_1440_0, i_8_480_1443_0,
    i_8_480_1461_0, i_8_480_1462_0, i_8_480_1481_0, i_8_480_1518_0,
    i_8_480_1524_0, i_8_480_1525_0, i_8_480_1548_0, i_8_480_1549_0,
    i_8_480_1587_0, i_8_480_1605_0, i_8_480_1638_0, i_8_480_1639_0,
    i_8_480_1695_0, i_8_480_1722_0, i_8_480_1724_0, i_8_480_1746_0,
    i_8_480_1783_0, i_8_480_1813_0, i_8_480_1839_0, i_8_480_1935_0,
    i_8_480_1967_0, i_8_480_1974_0, i_8_480_1995_0, i_8_480_2011_0,
    i_8_480_2053_0, i_8_480_2060_0, i_8_480_2110_0, i_8_480_2111_0,
    i_8_480_2232_0, i_8_480_2233_0, i_8_480_2247_0, i_8_480_2298_0;
  output o_8_480_0_0;
  assign o_8_480_0_0 = ~((~i_8_480_552_0 & ((~i_8_480_1425_0 & ((~i_8_480_109_0 & ((~i_8_480_13_0 & ~i_8_480_345_0 & ~i_8_480_486_0 & ~i_8_480_530_0 & ~i_8_480_894_0 & ~i_8_480_1336_0 & ~i_8_480_1524_0 & ~i_8_480_1839_0 & ~i_8_480_2060_0) | (i_8_480_970_0 & ~i_8_480_1324_0 & ~i_8_480_1462_0 & ~i_8_480_1548_0 & ~i_8_480_1695_0 & ~i_8_480_2298_0))) | (~i_8_480_114_0 & ~i_8_480_530_0 & i_8_480_696_0 & ~i_8_480_891_0 & ~i_8_480_894_0 & ~i_8_480_1155_0 & ~i_8_480_1461_0 & ~i_8_480_1525_0 & ~i_8_480_1935_0))) | (~i_8_480_285_0 & ~i_8_480_1422_0 & ((~i_8_480_138_0 & ~i_8_480_555_0 & ~i_8_480_777_0 & ~i_8_480_1036_0 & ~i_8_480_1152_0) | (~i_8_480_66_0 & i_8_480_877_0 & ~i_8_480_1423_0 & ~i_8_480_1440_0 & ~i_8_480_1443_0 & ~i_8_480_1695_0))) | (i_8_480_838_0 & i_8_480_2110_0) | (i_8_480_696_0 & ~i_8_480_969_0 & ~i_8_480_1461_0 & i_8_480_2232_0) | (~i_8_480_279_0 & ~i_8_480_400_0 & ~i_8_480_573_0 & ~i_8_480_970_0 & ~i_8_480_1152_0 & ~i_8_480_1155_0 & ~i_8_480_1518_0 & ~i_8_480_1549_0 & ~i_8_480_2011_0 & ~i_8_480_2298_0))) | (~i_8_480_894_0 & ((~i_8_480_13_0 & ~i_8_480_2247_0 & ((i_8_480_345_0 & ~i_8_480_492_0 & ~i_8_480_883_0 & ~i_8_480_1036_0 & ~i_8_480_1440_0 & ~i_8_480_1461_0 & ~i_8_480_1605_0 & ~i_8_480_1724_0) | (~i_8_480_321_0 & ~i_8_480_573_0 & ~i_8_480_838_0 & ~i_8_480_891_0 & ~i_8_480_1423_0 & ~i_8_480_1695_0 & ~i_8_480_1839_0))) | (~i_8_480_220_0 & ~i_8_480_1524_0 & ((~i_8_480_22_0 & ~i_8_480_279_0 & ~i_8_480_555_0 & ~i_8_480_573_0 & ~i_8_480_874_0 & ~i_8_480_969_0 & ~i_8_480_1137_0 & ~i_8_480_1155_0 & ~i_8_480_1440_0 & ~i_8_480_1462_0) | (~i_8_480_321_0 & ~i_8_480_589_0 & ~i_8_480_970_0 & ~i_8_480_1423_0 & ~i_8_480_1461_0 & ~i_8_480_1518_0 & ~i_8_480_1525_0 & ~i_8_480_1548_0 & ~i_8_480_1638_0))) | (~i_8_480_573_0 & ~i_8_480_822_0 & ~i_8_480_1092_0 & i_8_480_1111_0 & ~i_8_480_1152_0 & ~i_8_480_1197_0 & ~i_8_480_1423_0 & ~i_8_480_1481_0 & ~i_8_480_1548_0) | (~i_8_480_589_0 & ~i_8_480_606_0 & ~i_8_480_970_0 & ~i_8_480_1036_0 & ~i_8_480_1155_0 & ~i_8_480_1317_0 & ~i_8_480_1336_0 & ~i_8_480_1422_0 & ~i_8_480_1443_0 & ~i_8_480_1587_0 & ~i_8_480_1967_0))) | (~i_8_480_219_0 & ((i_8_480_492_0 & i_8_480_696_0 & ~i_8_480_1443_0 & ~i_8_480_1461_0) | (~i_8_480_321_0 & ~i_8_480_573_0 & ~i_8_480_589_0 & ~i_8_480_594_0 & ~i_8_480_891_0 & ~i_8_480_1111_0 & ~i_8_480_1524_0 & ~i_8_480_1695_0 & ~i_8_480_2298_0))) | (~i_8_480_1462_0 & ((~i_8_480_396_0 & ((i_8_480_220_0 & ~i_8_480_1036_0 & i_8_480_1111_0 & ~i_8_480_1155_0 & ~i_8_480_1422_0 & ~i_8_480_1443_0 & ~i_8_480_1525_0) | (i_8_480_384_0 & i_8_480_696_0 & ~i_8_480_1524_0 & ~i_8_480_1746_0))) | (i_8_480_21_0 & ~i_8_480_138_0 & ~i_8_480_883_0 & ~i_8_480_1324_0 & ~i_8_480_1461_0 & ~i_8_480_2298_0))) | (~i_8_480_138_0 & ~i_8_480_1443_0 & ((i_8_480_1029_0 & ~i_8_480_1422_0 & ~i_8_480_1839_0) | (~i_8_480_321_0 & ~i_8_480_530_0 & ~i_8_480_573_0 & ~i_8_480_589_0 & ~i_8_480_838_0 & ~i_8_480_972_0 & ~i_8_480_1155_0 & ~i_8_480_1461_0 & ~i_8_480_1524_0 & ~i_8_480_2060_0))) | (i_8_480_527_0 & ((~i_8_480_220_0 & ~i_8_480_1425_0) | (~i_8_480_615_0 & ~i_8_480_1440_0 & ~i_8_480_1461_0 & ~i_8_480_1481_0 & ~i_8_480_1524_0 & ~i_8_480_1549_0))) | (i_8_480_552_0 & ~i_8_480_1518_0 & ((i_8_480_364_0 & ~i_8_480_1152_0 & ~i_8_480_1197_0 & ~i_8_480_1317_0 & ~i_8_480_1422_0 & ~i_8_480_1461_0 & ~i_8_480_2247_0) | (i_8_480_345_0 & ~i_8_480_891_0 & ~i_8_480_1639_0 & ~i_8_480_1722_0 & ~i_8_480_1935_0 & ~i_8_480_2298_0))) | (~i_8_480_1152_0 & ((~i_8_480_970_0 & ~i_8_480_1440_0 & ((~i_8_480_1461_0 & i_8_480_2232_0) | (i_8_480_138_0 & ~i_8_480_1036_0 & ~i_8_480_1137_0 & ~i_8_480_1336_0 & ~i_8_480_1722_0 & ~i_8_480_1783_0 & ~i_8_480_2298_0))) | (~i_8_480_606_0 & ~i_8_480_608_0 & ~i_8_480_822_0 & ~i_8_480_891_0 & ~i_8_480_969_0 & ~i_8_480_1155_0 & ~i_8_480_1746_0 & ~i_8_480_1995_0 & ~i_8_480_2298_0))) | (~i_8_480_1722_0 & ((i_8_480_877_0 & i_8_480_1255_0) | (~i_8_480_279_0 & ~i_8_480_555_0 & ~i_8_480_1036_0 & ~i_8_480_1423_0 & ~i_8_480_1695_0 & ~i_8_480_1839_0 & i_8_480_1995_0 & ~i_8_480_2298_0))) | (~i_8_480_285_0 & i_8_480_589_0 & ~i_8_480_1197_0 & ~i_8_480_1524_0 & ~i_8_480_1783_0 & i_8_480_1813_0));
endmodule



// Benchmark "kernel_8_481" written by ABC on Sun Jul 19 10:11:32 2020

module kernel_8_481 ( 
    i_8_481_31_0, i_8_481_70_0, i_8_481_187_0, i_8_481_188_0,
    i_8_481_259_0, i_8_481_301_0, i_8_481_305_0, i_8_481_367_0,
    i_8_481_368_0, i_8_481_430_0, i_8_481_454_0, i_8_481_493_0,
    i_8_481_505_0, i_8_481_512_0, i_8_481_556_0, i_8_481_565_0,
    i_8_481_584_0, i_8_481_593_0, i_8_481_596_0, i_8_481_599_0,
    i_8_481_607_0, i_8_481_610_0, i_8_481_627_0, i_8_481_630_0,
    i_8_481_631_0, i_8_481_634_0, i_8_481_643_0, i_8_481_654_0,
    i_8_481_682_0, i_8_481_707_0, i_8_481_778_0, i_8_481_781_0,
    i_8_481_782_0, i_8_481_796_0, i_8_481_842_0, i_8_481_844_0,
    i_8_481_865_0, i_8_481_890_0, i_8_481_965_0, i_8_481_976_0,
    i_8_481_977_0, i_8_481_1042_0, i_8_481_1069_0, i_8_481_1105_0,
    i_8_481_1167_0, i_8_481_1183_0, i_8_481_1201_0, i_8_481_1222_0,
    i_8_481_1228_0, i_8_481_1244_0, i_8_481_1246_0, i_8_481_1262_0,
    i_8_481_1264_0, i_8_481_1297_0, i_8_481_1300_0, i_8_481_1313_0,
    i_8_481_1318_0, i_8_481_1331_0, i_8_481_1427_0, i_8_481_1465_0,
    i_8_481_1468_0, i_8_481_1471_0, i_8_481_1474_0, i_8_481_1483_0,
    i_8_481_1516_0, i_8_481_1525_0, i_8_481_1543_0, i_8_481_1552_0,
    i_8_481_1675_0, i_8_481_1688_0, i_8_481_1694_0, i_8_481_1705_0,
    i_8_481_1750_0, i_8_481_1752_0, i_8_481_1771_0, i_8_481_1772_0,
    i_8_481_1783_0, i_8_481_1792_0, i_8_481_1795_0, i_8_481_1821_0,
    i_8_481_1837_0, i_8_481_1843_0, i_8_481_1888_0, i_8_481_1912_0,
    i_8_481_1937_0, i_8_481_1943_0, i_8_481_1959_0, i_8_481_1996_0,
    i_8_481_2047_0, i_8_481_2063_0, i_8_481_2077_0, i_8_481_2132_0,
    i_8_481_2139_0, i_8_481_2149_0, i_8_481_2155_0, i_8_481_2165_0,
    i_8_481_2223_0, i_8_481_2227_0, i_8_481_2233_0, i_8_481_2248_0,
    o_8_481_0_0  );
  input  i_8_481_31_0, i_8_481_70_0, i_8_481_187_0, i_8_481_188_0,
    i_8_481_259_0, i_8_481_301_0, i_8_481_305_0, i_8_481_367_0,
    i_8_481_368_0, i_8_481_430_0, i_8_481_454_0, i_8_481_493_0,
    i_8_481_505_0, i_8_481_512_0, i_8_481_556_0, i_8_481_565_0,
    i_8_481_584_0, i_8_481_593_0, i_8_481_596_0, i_8_481_599_0,
    i_8_481_607_0, i_8_481_610_0, i_8_481_627_0, i_8_481_630_0,
    i_8_481_631_0, i_8_481_634_0, i_8_481_643_0, i_8_481_654_0,
    i_8_481_682_0, i_8_481_707_0, i_8_481_778_0, i_8_481_781_0,
    i_8_481_782_0, i_8_481_796_0, i_8_481_842_0, i_8_481_844_0,
    i_8_481_865_0, i_8_481_890_0, i_8_481_965_0, i_8_481_976_0,
    i_8_481_977_0, i_8_481_1042_0, i_8_481_1069_0, i_8_481_1105_0,
    i_8_481_1167_0, i_8_481_1183_0, i_8_481_1201_0, i_8_481_1222_0,
    i_8_481_1228_0, i_8_481_1244_0, i_8_481_1246_0, i_8_481_1262_0,
    i_8_481_1264_0, i_8_481_1297_0, i_8_481_1300_0, i_8_481_1313_0,
    i_8_481_1318_0, i_8_481_1331_0, i_8_481_1427_0, i_8_481_1465_0,
    i_8_481_1468_0, i_8_481_1471_0, i_8_481_1474_0, i_8_481_1483_0,
    i_8_481_1516_0, i_8_481_1525_0, i_8_481_1543_0, i_8_481_1552_0,
    i_8_481_1675_0, i_8_481_1688_0, i_8_481_1694_0, i_8_481_1705_0,
    i_8_481_1750_0, i_8_481_1752_0, i_8_481_1771_0, i_8_481_1772_0,
    i_8_481_1783_0, i_8_481_1792_0, i_8_481_1795_0, i_8_481_1821_0,
    i_8_481_1837_0, i_8_481_1843_0, i_8_481_1888_0, i_8_481_1912_0,
    i_8_481_1937_0, i_8_481_1943_0, i_8_481_1959_0, i_8_481_1996_0,
    i_8_481_2047_0, i_8_481_2063_0, i_8_481_2077_0, i_8_481_2132_0,
    i_8_481_2139_0, i_8_481_2149_0, i_8_481_2155_0, i_8_481_2165_0,
    i_8_481_2223_0, i_8_481_2227_0, i_8_481_2233_0, i_8_481_2248_0;
  output o_8_481_0_0;
  assign o_8_481_0_0 = 0;
endmodule



// Benchmark "kernel_8_482" written by ABC on Sun Jul 19 10:11:33 2020

module kernel_8_482 ( 
    i_8_482_49_0, i_8_482_65_0, i_8_482_114_0, i_8_482_168_0,
    i_8_482_211_0, i_8_482_212_0, i_8_482_219_0, i_8_482_223_0,
    i_8_482_227_0, i_8_482_252_0, i_8_482_353_0, i_8_482_372_0,
    i_8_482_422_0, i_8_482_453_0, i_8_482_456_0, i_8_482_472_0,
    i_8_482_481_0, i_8_482_483_0, i_8_482_496_0, i_8_482_526_0,
    i_8_482_552_0, i_8_482_555_0, i_8_482_573_0, i_8_482_628_0,
    i_8_482_636_0, i_8_482_661_0, i_8_482_698_0, i_8_482_708_0,
    i_8_482_807_0, i_8_482_840_0, i_8_482_861_0, i_8_482_888_0,
    i_8_482_923_0, i_8_482_929_0, i_8_482_942_0, i_8_482_993_0,
    i_8_482_996_0, i_8_482_1102_0, i_8_482_1113_0, i_8_482_1114_0,
    i_8_482_1123_0, i_8_482_1171_0, i_8_482_1172_0, i_8_482_1185_0,
    i_8_482_1215_0, i_8_482_1224_0, i_8_482_1225_0, i_8_482_1260_0,
    i_8_482_1261_0, i_8_482_1263_0, i_8_482_1281_0, i_8_482_1282_0,
    i_8_482_1284_0, i_8_482_1287_0, i_8_482_1288_0, i_8_482_1293_0,
    i_8_482_1299_0, i_8_482_1308_0, i_8_482_1318_0, i_8_482_1324_0,
    i_8_482_1338_0, i_8_482_1386_0, i_8_482_1389_0, i_8_482_1395_0,
    i_8_482_1534_0, i_8_482_1542_0, i_8_482_1590_0, i_8_482_1591_0,
    i_8_482_1623_0, i_8_482_1626_0, i_8_482_1645_0, i_8_482_1653_0,
    i_8_482_1677_0, i_8_482_1680_0, i_8_482_1686_0, i_8_482_1689_0,
    i_8_482_1690_0, i_8_482_1698_0, i_8_482_1722_0, i_8_482_1735_0,
    i_8_482_1740_0, i_8_482_1741_0, i_8_482_1820_0, i_8_482_1822_0,
    i_8_482_1887_0, i_8_482_1914_0, i_8_482_1969_0, i_8_482_1996_0,
    i_8_482_2016_0, i_8_482_2018_0, i_8_482_2077_0, i_8_482_2121_0,
    i_8_482_2146_0, i_8_482_2155_0, i_8_482_2175_0, i_8_482_2244_0,
    i_8_482_2247_0, i_8_482_2259_0, i_8_482_2266_0, i_8_482_2287_0,
    o_8_482_0_0  );
  input  i_8_482_49_0, i_8_482_65_0, i_8_482_114_0, i_8_482_168_0,
    i_8_482_211_0, i_8_482_212_0, i_8_482_219_0, i_8_482_223_0,
    i_8_482_227_0, i_8_482_252_0, i_8_482_353_0, i_8_482_372_0,
    i_8_482_422_0, i_8_482_453_0, i_8_482_456_0, i_8_482_472_0,
    i_8_482_481_0, i_8_482_483_0, i_8_482_496_0, i_8_482_526_0,
    i_8_482_552_0, i_8_482_555_0, i_8_482_573_0, i_8_482_628_0,
    i_8_482_636_0, i_8_482_661_0, i_8_482_698_0, i_8_482_708_0,
    i_8_482_807_0, i_8_482_840_0, i_8_482_861_0, i_8_482_888_0,
    i_8_482_923_0, i_8_482_929_0, i_8_482_942_0, i_8_482_993_0,
    i_8_482_996_0, i_8_482_1102_0, i_8_482_1113_0, i_8_482_1114_0,
    i_8_482_1123_0, i_8_482_1171_0, i_8_482_1172_0, i_8_482_1185_0,
    i_8_482_1215_0, i_8_482_1224_0, i_8_482_1225_0, i_8_482_1260_0,
    i_8_482_1261_0, i_8_482_1263_0, i_8_482_1281_0, i_8_482_1282_0,
    i_8_482_1284_0, i_8_482_1287_0, i_8_482_1288_0, i_8_482_1293_0,
    i_8_482_1299_0, i_8_482_1308_0, i_8_482_1318_0, i_8_482_1324_0,
    i_8_482_1338_0, i_8_482_1386_0, i_8_482_1389_0, i_8_482_1395_0,
    i_8_482_1534_0, i_8_482_1542_0, i_8_482_1590_0, i_8_482_1591_0,
    i_8_482_1623_0, i_8_482_1626_0, i_8_482_1645_0, i_8_482_1653_0,
    i_8_482_1677_0, i_8_482_1680_0, i_8_482_1686_0, i_8_482_1689_0,
    i_8_482_1690_0, i_8_482_1698_0, i_8_482_1722_0, i_8_482_1735_0,
    i_8_482_1740_0, i_8_482_1741_0, i_8_482_1820_0, i_8_482_1822_0,
    i_8_482_1887_0, i_8_482_1914_0, i_8_482_1969_0, i_8_482_1996_0,
    i_8_482_2016_0, i_8_482_2018_0, i_8_482_2077_0, i_8_482_2121_0,
    i_8_482_2146_0, i_8_482_2155_0, i_8_482_2175_0, i_8_482_2244_0,
    i_8_482_2247_0, i_8_482_2259_0, i_8_482_2266_0, i_8_482_2287_0;
  output o_8_482_0_0;
  assign o_8_482_0_0 = 0;
endmodule



// Benchmark "kernel_8_483" written by ABC on Sun Jul 19 10:11:34 2020

module kernel_8_483 ( 
    i_8_483_19_0, i_8_483_77_0, i_8_483_116_0, i_8_483_143_0,
    i_8_483_151_0, i_8_483_189_0, i_8_483_247_0, i_8_483_302_0,
    i_8_483_310_0, i_8_483_319_0, i_8_483_322_0, i_8_483_323_0,
    i_8_483_346_0, i_8_483_361_0, i_8_483_427_0, i_8_483_481_0,
    i_8_483_489_0, i_8_483_492_0, i_8_483_498_0, i_8_483_508_0,
    i_8_483_523_0, i_8_483_536_0, i_8_483_553_0, i_8_483_556_0,
    i_8_483_572_0, i_8_483_575_0, i_8_483_580_0, i_8_483_584_0,
    i_8_483_607_0, i_8_483_636_0, i_8_483_637_0, i_8_483_643_0,
    i_8_483_644_0, i_8_483_650_0, i_8_483_682_0, i_8_483_703_0,
    i_8_483_705_0, i_8_483_751_0, i_8_483_841_0, i_8_483_928_0,
    i_8_483_941_0, i_8_483_973_0, i_8_483_1015_0, i_8_483_1083_0,
    i_8_483_1115_0, i_8_483_1237_0, i_8_483_1282_0, i_8_483_1315_0,
    i_8_483_1328_0, i_8_483_1339_0, i_8_483_1382_0, i_8_483_1403_0,
    i_8_483_1436_0, i_8_483_1445_0, i_8_483_1462_0, i_8_483_1463_0,
    i_8_483_1477_0, i_8_483_1507_0, i_8_483_1508_0, i_8_483_1510_0,
    i_8_483_1511_0, i_8_483_1520_0, i_8_483_1535_0, i_8_483_1552_0,
    i_8_483_1555_0, i_8_483_1628_0, i_8_483_1633_0, i_8_483_1648_0,
    i_8_483_1690_0, i_8_483_1691_0, i_8_483_1694_0, i_8_483_1700_0,
    i_8_483_1750_0, i_8_483_1751_0, i_8_483_1753_0, i_8_483_1754_0,
    i_8_483_1771_0, i_8_483_1772_0, i_8_483_1822_0, i_8_483_1840_0,
    i_8_483_1841_0, i_8_483_1864_0, i_8_483_1894_0, i_8_483_1912_0,
    i_8_483_1940_0, i_8_483_1952_0, i_8_483_1974_0, i_8_483_1983_0,
    i_8_483_1997_0, i_8_483_2075_0, i_8_483_2104_0, i_8_483_2137_0,
    i_8_483_2138_0, i_8_483_2140_0, i_8_483_2147_0, i_8_483_2153_0,
    i_8_483_2158_0, i_8_483_2216_0, i_8_483_2230_0, i_8_483_2289_0,
    o_8_483_0_0  );
  input  i_8_483_19_0, i_8_483_77_0, i_8_483_116_0, i_8_483_143_0,
    i_8_483_151_0, i_8_483_189_0, i_8_483_247_0, i_8_483_302_0,
    i_8_483_310_0, i_8_483_319_0, i_8_483_322_0, i_8_483_323_0,
    i_8_483_346_0, i_8_483_361_0, i_8_483_427_0, i_8_483_481_0,
    i_8_483_489_0, i_8_483_492_0, i_8_483_498_0, i_8_483_508_0,
    i_8_483_523_0, i_8_483_536_0, i_8_483_553_0, i_8_483_556_0,
    i_8_483_572_0, i_8_483_575_0, i_8_483_580_0, i_8_483_584_0,
    i_8_483_607_0, i_8_483_636_0, i_8_483_637_0, i_8_483_643_0,
    i_8_483_644_0, i_8_483_650_0, i_8_483_682_0, i_8_483_703_0,
    i_8_483_705_0, i_8_483_751_0, i_8_483_841_0, i_8_483_928_0,
    i_8_483_941_0, i_8_483_973_0, i_8_483_1015_0, i_8_483_1083_0,
    i_8_483_1115_0, i_8_483_1237_0, i_8_483_1282_0, i_8_483_1315_0,
    i_8_483_1328_0, i_8_483_1339_0, i_8_483_1382_0, i_8_483_1403_0,
    i_8_483_1436_0, i_8_483_1445_0, i_8_483_1462_0, i_8_483_1463_0,
    i_8_483_1477_0, i_8_483_1507_0, i_8_483_1508_0, i_8_483_1510_0,
    i_8_483_1511_0, i_8_483_1520_0, i_8_483_1535_0, i_8_483_1552_0,
    i_8_483_1555_0, i_8_483_1628_0, i_8_483_1633_0, i_8_483_1648_0,
    i_8_483_1690_0, i_8_483_1691_0, i_8_483_1694_0, i_8_483_1700_0,
    i_8_483_1750_0, i_8_483_1751_0, i_8_483_1753_0, i_8_483_1754_0,
    i_8_483_1771_0, i_8_483_1772_0, i_8_483_1822_0, i_8_483_1840_0,
    i_8_483_1841_0, i_8_483_1864_0, i_8_483_1894_0, i_8_483_1912_0,
    i_8_483_1940_0, i_8_483_1952_0, i_8_483_1974_0, i_8_483_1983_0,
    i_8_483_1997_0, i_8_483_2075_0, i_8_483_2104_0, i_8_483_2137_0,
    i_8_483_2138_0, i_8_483_2140_0, i_8_483_2147_0, i_8_483_2153_0,
    i_8_483_2158_0, i_8_483_2216_0, i_8_483_2230_0, i_8_483_2289_0;
  output o_8_483_0_0;
  assign o_8_483_0_0 = 0;
endmodule



// Benchmark "kernel_8_484" written by ABC on Sun Jul 19 10:11:35 2020

module kernel_8_484 ( 
    i_8_484_104_0, i_8_484_127_0, i_8_484_145_0, i_8_484_176_0,
    i_8_484_190_0, i_8_484_217_0, i_8_484_219_0, i_8_484_274_0,
    i_8_484_305_0, i_8_484_334_0, i_8_484_352_0, i_8_484_360_0,
    i_8_484_370_0, i_8_484_417_0, i_8_484_427_0, i_8_484_481_0,
    i_8_484_490_0, i_8_484_495_0, i_8_484_496_0, i_8_484_514_0,
    i_8_484_522_0, i_8_484_523_0, i_8_484_552_0, i_8_484_595_0,
    i_8_484_604_0, i_8_484_607_0, i_8_484_658_0, i_8_484_667_0,
    i_8_484_669_0, i_8_484_712_0, i_8_484_828_0, i_8_484_831_0,
    i_8_484_849_0, i_8_484_855_0, i_8_484_878_0, i_8_484_1027_0,
    i_8_484_1041_0, i_8_484_1071_0, i_8_484_1126_0, i_8_484_1129_0,
    i_8_484_1156_0, i_8_484_1174_0, i_8_484_1197_0, i_8_484_1225_0,
    i_8_484_1260_0, i_8_484_1282_0, i_8_484_1296_0, i_8_484_1297_0,
    i_8_484_1354_0, i_8_484_1387_0, i_8_484_1396_0, i_8_484_1486_0,
    i_8_484_1494_0, i_8_484_1506_0, i_8_484_1522_0, i_8_484_1531_0,
    i_8_484_1571_0, i_8_484_1649_0, i_8_484_1651_0, i_8_484_1665_0,
    i_8_484_1670_0, i_8_484_1681_0, i_8_484_1683_0, i_8_484_1693_0,
    i_8_484_1702_0, i_8_484_1729_0, i_8_484_1745_0, i_8_484_1747_0,
    i_8_484_1773_0, i_8_484_1774_0, i_8_484_1791_0, i_8_484_1794_0,
    i_8_484_1809_0, i_8_484_1813_0, i_8_484_1822_0, i_8_484_1846_0,
    i_8_484_1863_0, i_8_484_1870_0, i_8_484_1944_0, i_8_484_1945_0,
    i_8_484_1946_0, i_8_484_1947_0, i_8_484_1964_0, i_8_484_1965_0,
    i_8_484_1966_0, i_8_484_2007_0, i_8_484_2044_0, i_8_484_2045_0,
    i_8_484_2046_0, i_8_484_2061_0, i_8_484_2112_0, i_8_484_2116_0,
    i_8_484_2120_0, i_8_484_2125_0, i_8_484_2188_0, i_8_484_2230_0,
    i_8_484_2232_0, i_8_484_2260_0, i_8_484_2261_0, i_8_484_2263_0,
    o_8_484_0_0  );
  input  i_8_484_104_0, i_8_484_127_0, i_8_484_145_0, i_8_484_176_0,
    i_8_484_190_0, i_8_484_217_0, i_8_484_219_0, i_8_484_274_0,
    i_8_484_305_0, i_8_484_334_0, i_8_484_352_0, i_8_484_360_0,
    i_8_484_370_0, i_8_484_417_0, i_8_484_427_0, i_8_484_481_0,
    i_8_484_490_0, i_8_484_495_0, i_8_484_496_0, i_8_484_514_0,
    i_8_484_522_0, i_8_484_523_0, i_8_484_552_0, i_8_484_595_0,
    i_8_484_604_0, i_8_484_607_0, i_8_484_658_0, i_8_484_667_0,
    i_8_484_669_0, i_8_484_712_0, i_8_484_828_0, i_8_484_831_0,
    i_8_484_849_0, i_8_484_855_0, i_8_484_878_0, i_8_484_1027_0,
    i_8_484_1041_0, i_8_484_1071_0, i_8_484_1126_0, i_8_484_1129_0,
    i_8_484_1156_0, i_8_484_1174_0, i_8_484_1197_0, i_8_484_1225_0,
    i_8_484_1260_0, i_8_484_1282_0, i_8_484_1296_0, i_8_484_1297_0,
    i_8_484_1354_0, i_8_484_1387_0, i_8_484_1396_0, i_8_484_1486_0,
    i_8_484_1494_0, i_8_484_1506_0, i_8_484_1522_0, i_8_484_1531_0,
    i_8_484_1571_0, i_8_484_1649_0, i_8_484_1651_0, i_8_484_1665_0,
    i_8_484_1670_0, i_8_484_1681_0, i_8_484_1683_0, i_8_484_1693_0,
    i_8_484_1702_0, i_8_484_1729_0, i_8_484_1745_0, i_8_484_1747_0,
    i_8_484_1773_0, i_8_484_1774_0, i_8_484_1791_0, i_8_484_1794_0,
    i_8_484_1809_0, i_8_484_1813_0, i_8_484_1822_0, i_8_484_1846_0,
    i_8_484_1863_0, i_8_484_1870_0, i_8_484_1944_0, i_8_484_1945_0,
    i_8_484_1946_0, i_8_484_1947_0, i_8_484_1964_0, i_8_484_1965_0,
    i_8_484_1966_0, i_8_484_2007_0, i_8_484_2044_0, i_8_484_2045_0,
    i_8_484_2046_0, i_8_484_2061_0, i_8_484_2112_0, i_8_484_2116_0,
    i_8_484_2120_0, i_8_484_2125_0, i_8_484_2188_0, i_8_484_2230_0,
    i_8_484_2232_0, i_8_484_2260_0, i_8_484_2261_0, i_8_484_2263_0;
  output o_8_484_0_0;
  assign o_8_484_0_0 = 0;
endmodule



// Benchmark "kernel_8_485" written by ABC on Sun Jul 19 10:11:35 2020

module kernel_8_485 ( 
    i_8_485_11_0, i_8_485_52_0, i_8_485_84_0, i_8_485_93_0, i_8_485_153_0,
    i_8_485_172_0, i_8_485_174_0, i_8_485_241_0, i_8_485_245_0,
    i_8_485_300_0, i_8_485_306_0, i_8_485_345_0, i_8_485_346_0,
    i_8_485_354_0, i_8_485_363_0, i_8_485_381_0, i_8_485_384_0,
    i_8_485_385_0, i_8_485_450_0, i_8_485_457_0, i_8_485_507_0,
    i_8_485_523_0, i_8_485_526_0, i_8_485_528_0, i_8_485_609_0,
    i_8_485_612_0, i_8_485_615_0, i_8_485_634_0, i_8_485_642_0,
    i_8_485_660_0, i_8_485_675_0, i_8_485_694_0, i_8_485_702_0,
    i_8_485_705_0, i_8_485_709_0, i_8_485_764_0, i_8_485_768_0,
    i_8_485_795_0, i_8_485_804_0, i_8_485_822_0, i_8_485_880_0,
    i_8_485_921_0, i_8_485_924_0, i_8_485_930_0, i_8_485_967_0,
    i_8_485_993_0, i_8_485_1056_0, i_8_485_1170_0, i_8_485_1173_0,
    i_8_485_1174_0, i_8_485_1182_0, i_8_485_1189_0, i_8_485_1230_0,
    i_8_485_1233_0, i_8_485_1236_0, i_8_485_1239_0, i_8_485_1273_0,
    i_8_485_1288_0, i_8_485_1314_0, i_8_485_1332_0, i_8_485_1354_0,
    i_8_485_1371_0, i_8_485_1407_0, i_8_485_1440_0, i_8_485_1470_0,
    i_8_485_1489_0, i_8_485_1497_0, i_8_485_1560_0, i_8_485_1579_0,
    i_8_485_1605_0, i_8_485_1651_0, i_8_485_1654_0, i_8_485_1665_0,
    i_8_485_1686_0, i_8_485_1695_0, i_8_485_1758_0, i_8_485_1759_0,
    i_8_485_1777_0, i_8_485_1792_0, i_8_485_1807_0, i_8_485_1821_0,
    i_8_485_1824_0, i_8_485_1831_0, i_8_485_1858_0, i_8_485_1936_0,
    i_8_485_1938_0, i_8_485_2016_0, i_8_485_2019_0, i_8_485_2118_0,
    i_8_485_2146_0, i_8_485_2152_0, i_8_485_2158_0, i_8_485_2163_0,
    i_8_485_2172_0, i_8_485_2181_0, i_8_485_2182_0, i_8_485_2244_0,
    i_8_485_2245_0, i_8_485_2262_0, i_8_485_2283_0,
    o_8_485_0_0  );
  input  i_8_485_11_0, i_8_485_52_0, i_8_485_84_0, i_8_485_93_0,
    i_8_485_153_0, i_8_485_172_0, i_8_485_174_0, i_8_485_241_0,
    i_8_485_245_0, i_8_485_300_0, i_8_485_306_0, i_8_485_345_0,
    i_8_485_346_0, i_8_485_354_0, i_8_485_363_0, i_8_485_381_0,
    i_8_485_384_0, i_8_485_385_0, i_8_485_450_0, i_8_485_457_0,
    i_8_485_507_0, i_8_485_523_0, i_8_485_526_0, i_8_485_528_0,
    i_8_485_609_0, i_8_485_612_0, i_8_485_615_0, i_8_485_634_0,
    i_8_485_642_0, i_8_485_660_0, i_8_485_675_0, i_8_485_694_0,
    i_8_485_702_0, i_8_485_705_0, i_8_485_709_0, i_8_485_764_0,
    i_8_485_768_0, i_8_485_795_0, i_8_485_804_0, i_8_485_822_0,
    i_8_485_880_0, i_8_485_921_0, i_8_485_924_0, i_8_485_930_0,
    i_8_485_967_0, i_8_485_993_0, i_8_485_1056_0, i_8_485_1170_0,
    i_8_485_1173_0, i_8_485_1174_0, i_8_485_1182_0, i_8_485_1189_0,
    i_8_485_1230_0, i_8_485_1233_0, i_8_485_1236_0, i_8_485_1239_0,
    i_8_485_1273_0, i_8_485_1288_0, i_8_485_1314_0, i_8_485_1332_0,
    i_8_485_1354_0, i_8_485_1371_0, i_8_485_1407_0, i_8_485_1440_0,
    i_8_485_1470_0, i_8_485_1489_0, i_8_485_1497_0, i_8_485_1560_0,
    i_8_485_1579_0, i_8_485_1605_0, i_8_485_1651_0, i_8_485_1654_0,
    i_8_485_1665_0, i_8_485_1686_0, i_8_485_1695_0, i_8_485_1758_0,
    i_8_485_1759_0, i_8_485_1777_0, i_8_485_1792_0, i_8_485_1807_0,
    i_8_485_1821_0, i_8_485_1824_0, i_8_485_1831_0, i_8_485_1858_0,
    i_8_485_1936_0, i_8_485_1938_0, i_8_485_2016_0, i_8_485_2019_0,
    i_8_485_2118_0, i_8_485_2146_0, i_8_485_2152_0, i_8_485_2158_0,
    i_8_485_2163_0, i_8_485_2172_0, i_8_485_2181_0, i_8_485_2182_0,
    i_8_485_2244_0, i_8_485_2245_0, i_8_485_2262_0, i_8_485_2283_0;
  output o_8_485_0_0;
  assign o_8_485_0_0 = 0;
endmodule



// Benchmark "kernel_8_486" written by ABC on Sun Jul 19 10:11:36 2020

module kernel_8_486 ( 
    i_8_486_33_0, i_8_486_37_0, i_8_486_76_0, i_8_486_162_0, i_8_486_170_0,
    i_8_486_179_0, i_8_486_190_0, i_8_486_191_0, i_8_486_211_0,
    i_8_486_301_0, i_8_486_303_0, i_8_486_304_0, i_8_486_310_0,
    i_8_486_341_0, i_8_486_358_0, i_8_486_359_0, i_8_486_361_0,
    i_8_486_376_0, i_8_486_377_0, i_8_486_394_0, i_8_486_400_0,
    i_8_486_449_0, i_8_486_464_0, i_8_486_496_0, i_8_486_499_0,
    i_8_486_525_0, i_8_486_553_0, i_8_486_599_0, i_8_486_638_0,
    i_8_486_657_0, i_8_486_692_0, i_8_486_706_0, i_8_486_752_0,
    i_8_486_827_0, i_8_486_836_0, i_8_486_850_0, i_8_486_863_0,
    i_8_486_868_0, i_8_486_872_0, i_8_486_923_0, i_8_486_924_0,
    i_8_486_928_0, i_8_486_959_0, i_8_486_962_0, i_8_486_968_0,
    i_8_486_1003_0, i_8_486_1035_0, i_8_486_1079_0, i_8_486_1111_0,
    i_8_486_1126_0, i_8_486_1139_0, i_8_486_1227_0, i_8_486_1241_0,
    i_8_486_1258_0, i_8_486_1264_0, i_8_486_1266_0, i_8_486_1273_0,
    i_8_486_1274_0, i_8_486_1277_0, i_8_486_1312_0, i_8_486_1313_0,
    i_8_486_1346_0, i_8_486_1385_0, i_8_486_1400_0, i_8_486_1433_0,
    i_8_486_1437_0, i_8_486_1450_0, i_8_486_1467_0, i_8_486_1499_0,
    i_8_486_1552_0, i_8_486_1558_0, i_8_486_1598_0, i_8_486_1642_0,
    i_8_486_1654_0, i_8_486_1663_0, i_8_486_1678_0, i_8_486_1696_0,
    i_8_486_1702_0, i_8_486_1733_0, i_8_486_1750_0, i_8_486_1831_0,
    i_8_486_1870_0, i_8_486_1871_0, i_8_486_1877_0, i_8_486_1880_0,
    i_8_486_1885_0, i_8_486_1922_0, i_8_486_1996_0, i_8_486_2017_0,
    i_8_486_2048_0, i_8_486_2066_0, i_8_486_2069_0, i_8_486_2146_0,
    i_8_486_2147_0, i_8_486_2161_0, i_8_486_2186_0, i_8_486_2216_0,
    i_8_486_2237_0, i_8_486_2238_0, i_8_486_2285_0,
    o_8_486_0_0  );
  input  i_8_486_33_0, i_8_486_37_0, i_8_486_76_0, i_8_486_162_0,
    i_8_486_170_0, i_8_486_179_0, i_8_486_190_0, i_8_486_191_0,
    i_8_486_211_0, i_8_486_301_0, i_8_486_303_0, i_8_486_304_0,
    i_8_486_310_0, i_8_486_341_0, i_8_486_358_0, i_8_486_359_0,
    i_8_486_361_0, i_8_486_376_0, i_8_486_377_0, i_8_486_394_0,
    i_8_486_400_0, i_8_486_449_0, i_8_486_464_0, i_8_486_496_0,
    i_8_486_499_0, i_8_486_525_0, i_8_486_553_0, i_8_486_599_0,
    i_8_486_638_0, i_8_486_657_0, i_8_486_692_0, i_8_486_706_0,
    i_8_486_752_0, i_8_486_827_0, i_8_486_836_0, i_8_486_850_0,
    i_8_486_863_0, i_8_486_868_0, i_8_486_872_0, i_8_486_923_0,
    i_8_486_924_0, i_8_486_928_0, i_8_486_959_0, i_8_486_962_0,
    i_8_486_968_0, i_8_486_1003_0, i_8_486_1035_0, i_8_486_1079_0,
    i_8_486_1111_0, i_8_486_1126_0, i_8_486_1139_0, i_8_486_1227_0,
    i_8_486_1241_0, i_8_486_1258_0, i_8_486_1264_0, i_8_486_1266_0,
    i_8_486_1273_0, i_8_486_1274_0, i_8_486_1277_0, i_8_486_1312_0,
    i_8_486_1313_0, i_8_486_1346_0, i_8_486_1385_0, i_8_486_1400_0,
    i_8_486_1433_0, i_8_486_1437_0, i_8_486_1450_0, i_8_486_1467_0,
    i_8_486_1499_0, i_8_486_1552_0, i_8_486_1558_0, i_8_486_1598_0,
    i_8_486_1642_0, i_8_486_1654_0, i_8_486_1663_0, i_8_486_1678_0,
    i_8_486_1696_0, i_8_486_1702_0, i_8_486_1733_0, i_8_486_1750_0,
    i_8_486_1831_0, i_8_486_1870_0, i_8_486_1871_0, i_8_486_1877_0,
    i_8_486_1880_0, i_8_486_1885_0, i_8_486_1922_0, i_8_486_1996_0,
    i_8_486_2017_0, i_8_486_2048_0, i_8_486_2066_0, i_8_486_2069_0,
    i_8_486_2146_0, i_8_486_2147_0, i_8_486_2161_0, i_8_486_2186_0,
    i_8_486_2216_0, i_8_486_2237_0, i_8_486_2238_0, i_8_486_2285_0;
  output o_8_486_0_0;
  assign o_8_486_0_0 = 0;
endmodule



// Benchmark "kernel_8_487" written by ABC on Sun Jul 19 10:11:37 2020

module kernel_8_487 ( 
    i_8_487_24_0, i_8_487_39_0, i_8_487_49_0, i_8_487_52_0, i_8_487_85_0,
    i_8_487_97_0, i_8_487_170_0, i_8_487_175_0, i_8_487_181_0,
    i_8_487_189_0, i_8_487_193_0, i_8_487_238_0, i_8_487_263_0,
    i_8_487_277_0, i_8_487_300_0, i_8_487_302_0, i_8_487_313_0,
    i_8_487_340_0, i_8_487_345_0, i_8_487_378_0, i_8_487_403_0,
    i_8_487_494_0, i_8_487_556_0, i_8_487_603_0, i_8_487_613_0,
    i_8_487_634_0, i_8_487_637_0, i_8_487_676_0, i_8_487_687_0,
    i_8_487_698_0, i_8_487_700_0, i_8_487_706_0, i_8_487_707_0,
    i_8_487_748_0, i_8_487_769_0, i_8_487_798_0, i_8_487_840_0,
    i_8_487_849_0, i_8_487_855_0, i_8_487_879_0, i_8_487_883_0,
    i_8_487_924_0, i_8_487_925_0, i_8_487_931_0, i_8_487_934_0,
    i_8_487_970_0, i_8_487_990_0, i_8_487_1095_0, i_8_487_1146_0,
    i_8_487_1230_0, i_8_487_1236_0, i_8_487_1254_0, i_8_487_1273_0,
    i_8_487_1289_0, i_8_487_1339_0, i_8_487_1350_0, i_8_487_1355_0,
    i_8_487_1410_0, i_8_487_1455_0, i_8_487_1459_0, i_8_487_1489_0,
    i_8_487_1512_0, i_8_487_1536_0, i_8_487_1598_0, i_8_487_1606_0,
    i_8_487_1634_0, i_8_487_1749_0, i_8_487_1788_0, i_8_487_1824_0,
    i_8_487_1828_0, i_8_487_1831_0, i_8_487_1860_0, i_8_487_1884_0,
    i_8_487_1885_0, i_8_487_1908_0, i_8_487_1940_0, i_8_487_1947_0,
    i_8_487_1951_0, i_8_487_1986_0, i_8_487_2004_0, i_8_487_2019_0,
    i_8_487_2022_0, i_8_487_2091_0, i_8_487_2112_0, i_8_487_2149_0,
    i_8_487_2157_0, i_8_487_2172_0, i_8_487_2175_0, i_8_487_2182_0,
    i_8_487_2196_0, i_8_487_2202_0, i_8_487_2211_0, i_8_487_2227_0,
    i_8_487_2233_0, i_8_487_2235_0, i_8_487_2275_0, i_8_487_2283_0,
    i_8_487_2284_0, i_8_487_2292_0, i_8_487_2299_0,
    o_8_487_0_0  );
  input  i_8_487_24_0, i_8_487_39_0, i_8_487_49_0, i_8_487_52_0,
    i_8_487_85_0, i_8_487_97_0, i_8_487_170_0, i_8_487_175_0,
    i_8_487_181_0, i_8_487_189_0, i_8_487_193_0, i_8_487_238_0,
    i_8_487_263_0, i_8_487_277_0, i_8_487_300_0, i_8_487_302_0,
    i_8_487_313_0, i_8_487_340_0, i_8_487_345_0, i_8_487_378_0,
    i_8_487_403_0, i_8_487_494_0, i_8_487_556_0, i_8_487_603_0,
    i_8_487_613_0, i_8_487_634_0, i_8_487_637_0, i_8_487_676_0,
    i_8_487_687_0, i_8_487_698_0, i_8_487_700_0, i_8_487_706_0,
    i_8_487_707_0, i_8_487_748_0, i_8_487_769_0, i_8_487_798_0,
    i_8_487_840_0, i_8_487_849_0, i_8_487_855_0, i_8_487_879_0,
    i_8_487_883_0, i_8_487_924_0, i_8_487_925_0, i_8_487_931_0,
    i_8_487_934_0, i_8_487_970_0, i_8_487_990_0, i_8_487_1095_0,
    i_8_487_1146_0, i_8_487_1230_0, i_8_487_1236_0, i_8_487_1254_0,
    i_8_487_1273_0, i_8_487_1289_0, i_8_487_1339_0, i_8_487_1350_0,
    i_8_487_1355_0, i_8_487_1410_0, i_8_487_1455_0, i_8_487_1459_0,
    i_8_487_1489_0, i_8_487_1512_0, i_8_487_1536_0, i_8_487_1598_0,
    i_8_487_1606_0, i_8_487_1634_0, i_8_487_1749_0, i_8_487_1788_0,
    i_8_487_1824_0, i_8_487_1828_0, i_8_487_1831_0, i_8_487_1860_0,
    i_8_487_1884_0, i_8_487_1885_0, i_8_487_1908_0, i_8_487_1940_0,
    i_8_487_1947_0, i_8_487_1951_0, i_8_487_1986_0, i_8_487_2004_0,
    i_8_487_2019_0, i_8_487_2022_0, i_8_487_2091_0, i_8_487_2112_0,
    i_8_487_2149_0, i_8_487_2157_0, i_8_487_2172_0, i_8_487_2175_0,
    i_8_487_2182_0, i_8_487_2196_0, i_8_487_2202_0, i_8_487_2211_0,
    i_8_487_2227_0, i_8_487_2233_0, i_8_487_2235_0, i_8_487_2275_0,
    i_8_487_2283_0, i_8_487_2284_0, i_8_487_2292_0, i_8_487_2299_0;
  output o_8_487_0_0;
  assign o_8_487_0_0 = 0;
endmodule



// Benchmark "kernel_8_488" written by ABC on Sun Jul 19 10:11:39 2020

module kernel_8_488 ( 
    i_8_488_37_0, i_8_488_75_0, i_8_488_81_0, i_8_488_129_0, i_8_488_192_0,
    i_8_488_193_0, i_8_488_214_0, i_8_488_225_0, i_8_488_230_0,
    i_8_488_241_0, i_8_488_242_0, i_8_488_337_0, i_8_488_343_0,
    i_8_488_347_0, i_8_488_365_0, i_8_488_478_0, i_8_488_482_0,
    i_8_488_483_0, i_8_488_484_0, i_8_488_502_0, i_8_488_525_0,
    i_8_488_528_0, i_8_488_588_0, i_8_488_612_0, i_8_488_616_0,
    i_8_488_619_0, i_8_488_620_0, i_8_488_631_0, i_8_488_653_0,
    i_8_488_654_0, i_8_488_655_0, i_8_488_656_0, i_8_488_664_0,
    i_8_488_669_0, i_8_488_687_0, i_8_488_690_0, i_8_488_710_0,
    i_8_488_732_0, i_8_488_751_0, i_8_488_760_0, i_8_488_762_0,
    i_8_488_763_0, i_8_488_765_0, i_8_488_768_0, i_8_488_769_0,
    i_8_488_770_0, i_8_488_772_0, i_8_488_792_0, i_8_488_796_0,
    i_8_488_831_0, i_8_488_832_0, i_8_488_833_0, i_8_488_841_0,
    i_8_488_970_0, i_8_488_971_0, i_8_488_1031_0, i_8_488_1056_0,
    i_8_488_1156_0, i_8_488_1158_0, i_8_488_1159_0, i_8_488_1263_0,
    i_8_488_1264_0, i_8_488_1265_0, i_8_488_1272_0, i_8_488_1273_0,
    i_8_488_1274_0, i_8_488_1306_0, i_8_488_1329_0, i_8_488_1331_0,
    i_8_488_1350_0, i_8_488_1353_0, i_8_488_1358_0, i_8_488_1407_0,
    i_8_488_1767_0, i_8_488_1768_0, i_8_488_1770_0, i_8_488_1781_0,
    i_8_488_1834_0, i_8_488_1995_0, i_8_488_1996_0, i_8_488_2001_0,
    i_8_488_2078_0, i_8_488_2110_0, i_8_488_2118_0, i_8_488_2119_0,
    i_8_488_2136_0, i_8_488_2138_0, i_8_488_2150_0, i_8_488_2170_0,
    i_8_488_2171_0, i_8_488_2208_0, i_8_488_2215_0, i_8_488_2216_0,
    i_8_488_2224_0, i_8_488_2243_0, i_8_488_2245_0, i_8_488_2248_0,
    i_8_488_2249_0, i_8_488_2273_0, i_8_488_2289_0,
    o_8_488_0_0  );
  input  i_8_488_37_0, i_8_488_75_0, i_8_488_81_0, i_8_488_129_0,
    i_8_488_192_0, i_8_488_193_0, i_8_488_214_0, i_8_488_225_0,
    i_8_488_230_0, i_8_488_241_0, i_8_488_242_0, i_8_488_337_0,
    i_8_488_343_0, i_8_488_347_0, i_8_488_365_0, i_8_488_478_0,
    i_8_488_482_0, i_8_488_483_0, i_8_488_484_0, i_8_488_502_0,
    i_8_488_525_0, i_8_488_528_0, i_8_488_588_0, i_8_488_612_0,
    i_8_488_616_0, i_8_488_619_0, i_8_488_620_0, i_8_488_631_0,
    i_8_488_653_0, i_8_488_654_0, i_8_488_655_0, i_8_488_656_0,
    i_8_488_664_0, i_8_488_669_0, i_8_488_687_0, i_8_488_690_0,
    i_8_488_710_0, i_8_488_732_0, i_8_488_751_0, i_8_488_760_0,
    i_8_488_762_0, i_8_488_763_0, i_8_488_765_0, i_8_488_768_0,
    i_8_488_769_0, i_8_488_770_0, i_8_488_772_0, i_8_488_792_0,
    i_8_488_796_0, i_8_488_831_0, i_8_488_832_0, i_8_488_833_0,
    i_8_488_841_0, i_8_488_970_0, i_8_488_971_0, i_8_488_1031_0,
    i_8_488_1056_0, i_8_488_1156_0, i_8_488_1158_0, i_8_488_1159_0,
    i_8_488_1263_0, i_8_488_1264_0, i_8_488_1265_0, i_8_488_1272_0,
    i_8_488_1273_0, i_8_488_1274_0, i_8_488_1306_0, i_8_488_1329_0,
    i_8_488_1331_0, i_8_488_1350_0, i_8_488_1353_0, i_8_488_1358_0,
    i_8_488_1407_0, i_8_488_1767_0, i_8_488_1768_0, i_8_488_1770_0,
    i_8_488_1781_0, i_8_488_1834_0, i_8_488_1995_0, i_8_488_1996_0,
    i_8_488_2001_0, i_8_488_2078_0, i_8_488_2110_0, i_8_488_2118_0,
    i_8_488_2119_0, i_8_488_2136_0, i_8_488_2138_0, i_8_488_2150_0,
    i_8_488_2170_0, i_8_488_2171_0, i_8_488_2208_0, i_8_488_2215_0,
    i_8_488_2216_0, i_8_488_2224_0, i_8_488_2243_0, i_8_488_2245_0,
    i_8_488_2248_0, i_8_488_2249_0, i_8_488_2273_0, i_8_488_2289_0;
  output o_8_488_0_0;
  assign o_8_488_0_0 = ~((i_8_488_75_0 & ((~i_8_488_81_0 & ~i_8_488_343_0 & ~i_8_488_483_0 & i_8_488_1767_0) | (~i_8_488_347_0 & ~i_8_488_478_0 & ~i_8_488_502_0 & i_8_488_612_0 & ~i_8_488_690_0 & ~i_8_488_768_0 & ~i_8_488_1781_0 & ~i_8_488_2208_0))) | (~i_8_488_484_0 & ((~i_8_488_770_0 & ((i_8_488_193_0 & ((~i_8_488_343_0 & ~i_8_488_631_0 & ~i_8_488_768_0 & i_8_488_841_0 & ~i_8_488_1158_0 & ~i_8_488_2215_0) | (~i_8_488_37_0 & ~i_8_488_347_0 & ~i_8_488_664_0 & ~i_8_488_690_0 & ~i_8_488_732_0 & ~i_8_488_772_0 & ~i_8_488_1056_0 & ~i_8_488_2216_0 & ~i_8_488_2224_0))) | (~i_8_488_478_0 & ~i_8_488_483_0 & ~i_8_488_502_0 & ~i_8_488_792_0 & ~i_8_488_833_0 & ~i_8_488_1265_0 & ~i_8_488_1329_0 & ~i_8_488_1331_0 & i_8_488_1353_0 & ~i_8_488_1781_0 & ~i_8_488_2001_0 & ~i_8_488_2215_0 & ~i_8_488_2216_0 & ~i_8_488_2243_0))) | (~i_8_488_214_0 & ((~i_8_488_37_0 & ~i_8_488_365_0 & ~i_8_488_482_0 & ~i_8_488_483_0 & ~i_8_488_687_0 & ~i_8_488_763_0 & ~i_8_488_765_0 & ~i_8_488_841_0 & ~i_8_488_1056_0 & ~i_8_488_1273_0 & ~i_8_488_1274_0 & ~i_8_488_2078_0 & ~i_8_488_2215_0 & ~i_8_488_2243_0 & ~i_8_488_2273_0) | (~i_8_488_612_0 & i_8_488_653_0 & ~i_8_488_769_0 & i_8_488_1265_0 & ~i_8_488_1767_0 & ~i_8_488_2289_0))) | (~i_8_488_1834_0 & ((~i_8_488_37_0 & ~i_8_488_690_0 & ((~i_8_488_230_0 & ~i_8_488_337_0 & ~i_8_488_482_0 & ~i_8_488_612_0 & ~i_8_488_687_0 & ~i_8_488_765_0 & ~i_8_488_796_0 & ~i_8_488_1274_0 & ~i_8_488_1331_0 & i_8_488_1353_0 & ~i_8_488_1407_0 & ~i_8_488_2001_0 & ~i_8_488_2078_0 & ~i_8_488_2171_0) | (~i_8_488_762_0 & ~i_8_488_763_0 & ~i_8_488_1056_0 & i_8_488_1995_0 & i_8_488_1996_0 & ~i_8_488_2208_0))) | (~i_8_488_347_0 & ~i_8_488_478_0 & i_8_488_656_0 & ~i_8_488_2248_0))) | (~i_8_488_525_0 & ((~i_8_488_765_0 & ~i_8_488_796_0 & ~i_8_488_337_0 & ~i_8_488_762_0 & ~i_8_488_833_0 & ~i_8_488_1159_0 & i_8_488_1263_0 & ~i_8_488_1272_0 & ~i_8_488_2215_0) | (~i_8_488_347_0 & ~i_8_488_483_0 & i_8_488_631_0 & ~i_8_488_760_0 & ~i_8_488_769_0 & ~i_8_488_1056_0 & ~i_8_488_1996_0 & ~i_8_488_2216_0))) | (~i_8_488_765_0 & ~i_8_488_1156_0 & ~i_8_488_1306_0 & ~i_8_488_1329_0 & i_8_488_1768_0 & i_8_488_1996_0) | (i_8_488_482_0 & i_8_488_971_0 & ~i_8_488_1781_0 & ~i_8_488_2150_0 & ~i_8_488_2216_0 & ~i_8_488_2273_0))) | (~i_8_488_765_0 & ((~i_8_488_37_0 & ((~i_8_488_347_0 & ~i_8_488_588_0 & ~i_8_488_760_0 & ~i_8_488_971_0 & ~i_8_488_1263_0 & ~i_8_488_1353_0 & ~i_8_488_2138_0 & i_8_488_2224_0 & ~i_8_488_2245_0) | (~i_8_488_129_0 & ~i_8_488_528_0 & ~i_8_488_669_0 & ~i_8_488_1056_0 & i_8_488_1263_0 & ~i_8_488_1781_0 & ~i_8_488_2150_0 & ~i_8_488_2289_0))) | (~i_8_488_81_0 & ~i_8_488_2216_0 & ((~i_8_488_241_0 & ~i_8_488_483_0 & ~i_8_488_664_0 & ~i_8_488_768_0 & ~i_8_488_772_0 & ~i_8_488_1350_0 & i_8_488_1995_0) | (~i_8_488_192_0 & ~i_8_488_214_0 & ~i_8_488_482_0 & ~i_8_488_525_0 & ~i_8_488_690_0 & ~i_8_488_760_0 & ~i_8_488_796_0 & ~i_8_488_1056_0 & ~i_8_488_1274_0 & ~i_8_488_1329_0 & i_8_488_1768_0 & ~i_8_488_2119_0 & ~i_8_488_2249_0))) | (~i_8_488_478_0 & ~i_8_488_1273_0 & ((~i_8_488_241_0 & ~i_8_488_482_0 & ~i_8_488_612_0 & i_8_488_833_0 & ~i_8_488_1159_0 & ~i_8_488_1306_0 & ~i_8_488_1768_0 & ~i_8_488_1995_0) | (~i_8_488_483_0 & ~i_8_488_687_0 & ~i_8_488_772_0 & ~i_8_488_796_0 & ~i_8_488_1274_0 & i_8_488_2170_0 & ~i_8_488_2243_0))) | (~i_8_488_796_0 & ~i_8_488_2273_0 & ((~i_8_488_687_0 & ((~i_8_488_230_0 & ~i_8_488_482_0 & ~i_8_488_620_0 & ~i_8_488_762_0 & ~i_8_488_763_0 & ~i_8_488_1306_0 & i_8_488_1781_0 & ~i_8_488_2078_0) | (i_8_488_588_0 & i_8_488_732_0 & ~i_8_488_1770_0 & ~i_8_488_2150_0))) | (~i_8_488_225_0 & ~i_8_488_483_0 & ~i_8_488_653_0 & ~i_8_488_690_0 & ~i_8_488_762_0 & ~i_8_488_772_0 & ~i_8_488_1158_0 & ~i_8_488_1159_0 & ~i_8_488_1274_0 & ~i_8_488_1331_0 & i_8_488_1995_0 & ~i_8_488_2078_0 & ~i_8_488_2208_0))) | (~i_8_488_528_0 & i_8_488_656_0 & i_8_488_710_0 & ~i_8_488_1274_0 & ~i_8_488_1834_0) | (~i_8_488_129_0 & ~i_8_488_588_0 & ~i_8_488_772_0 & ~i_8_488_841_0 & ~i_8_488_1031_0 & i_8_488_1263_0 & ~i_8_488_1306_0 & ~i_8_488_1353_0 & ~i_8_488_2001_0 & ~i_8_488_2215_0))) | (~i_8_488_588_0 & ((~i_8_488_242_0 & ~i_8_488_528_0 & ~i_8_488_616_0 & i_8_488_669_0 & ~i_8_488_760_0 & ~i_8_488_1056_0 & ~i_8_488_1407_0) | (~i_8_488_690_0 & i_8_488_831_0 & ~i_8_488_1273_0 & ~i_8_488_1274_0 & i_8_488_1353_0 & ~i_8_488_2078_0))) | (~i_8_488_2224_0 & ((~i_8_488_242_0 & ~i_8_488_2216_0 & ((~i_8_488_483_0 & ~i_8_488_687_0 & ~i_8_488_772_0 & ~i_8_488_796_0 & i_8_488_1358_0) | (~i_8_488_760_0 & i_8_488_833_0 & i_8_488_2138_0))) | (~i_8_488_763_0 & ((i_8_488_365_0 & i_8_488_971_0 & ~i_8_488_1331_0 & ~i_8_488_1996_0) | (~i_8_488_337_0 & ~i_8_488_620_0 & ~i_8_488_690_0 & ~i_8_488_769_0 & i_8_488_970_0 & ~i_8_488_1329_0 & ~i_8_488_1767_0 & ~i_8_488_1768_0 & ~i_8_488_1834_0 & ~i_8_488_2215_0))) | (~i_8_488_241_0 & i_8_488_631_0 & ~i_8_488_687_0 & i_8_488_1768_0) | (~i_8_488_528_0 & i_8_488_751_0 & ~i_8_488_760_0 & ~i_8_488_792_0 & ~i_8_488_796_0 & i_8_488_841_0 & ~i_8_488_1158_0 & ~i_8_488_1781_0 & ~i_8_488_1996_0 & ~i_8_488_2118_0) | (~i_8_488_525_0 & ~i_8_488_612_0 & ~i_8_488_619_0 & i_8_488_1264_0 & ~i_8_488_1265_0 & ~i_8_488_1274_0 & ~i_8_488_1768_0 & ~i_8_488_2138_0 & ~i_8_488_2243_0))) | (i_8_488_365_0 & ((~i_8_488_482_0 & i_8_488_619_0 & ~i_8_488_732_0 & ~i_8_488_762_0 & ~i_8_488_1031_0 & ~i_8_488_1331_0) | (~i_8_488_81_0 & ~i_8_488_241_0 & ~i_8_488_763_0 & ~i_8_488_1272_0 & ~i_8_488_1273_0 & ~i_8_488_1274_0 & i_8_488_2170_0 & ~i_8_488_2215_0))) | (~i_8_488_81_0 & ((~i_8_488_528_0 & ~i_8_488_616_0 & ~i_8_488_347_0 & ~i_8_488_482_0 & ~i_8_488_763_0 & ~i_8_488_796_0 & i_8_488_832_0 & ~i_8_488_1329_0 & ~i_8_488_1353_0) | (~i_8_488_502_0 & ~i_8_488_612_0 & ~i_8_488_762_0 & ~i_8_488_768_0 & ~i_8_488_770_0 & ~i_8_488_831_0 & ~i_8_488_833_0 & ~i_8_488_841_0 & ~i_8_488_1158_0 & i_8_488_1264_0 & ~i_8_488_1273_0 & ~i_8_488_1306_0 & ~i_8_488_1331_0 & ~i_8_488_2001_0 & ~i_8_488_2078_0 & ~i_8_488_2119_0 & ~i_8_488_2249_0 & ~i_8_488_2273_0))) | (~i_8_488_483_0 & ((~i_8_488_241_0 & ((~i_8_488_129_0 & ~i_8_488_482_0 & ~i_8_488_525_0 & i_8_488_619_0 & ~i_8_488_760_0 & ~i_8_488_1274_0 & ~i_8_488_1781_0 & ~i_8_488_2110_0) | (~i_8_488_230_0 & ~i_8_488_347_0 & ~i_8_488_365_0 & ~i_8_488_664_0 & ~i_8_488_792_0 & ~i_8_488_970_0 & i_8_488_1264_0 & ~i_8_488_2138_0 & i_8_488_2170_0))) | (~i_8_488_772_0 & ~i_8_488_833_0 & ~i_8_488_1274_0 & ~i_8_488_1329_0 & ~i_8_488_2110_0 & i_8_488_2138_0 & i_8_488_2150_0))) | (~i_8_488_528_0 & ((i_8_488_655_0 & ~i_8_488_772_0 & ~i_8_488_1056_0 & ~i_8_488_2078_0 & ~i_8_488_2208_0 & ~i_8_488_1306_0 & ~i_8_488_2001_0) | (i_8_488_654_0 & ~i_8_488_762_0 & ~i_8_488_768_0 & i_8_488_841_0 & ~i_8_488_1995_0 & ~i_8_488_2215_0))) | (~i_8_488_616_0 & ((~i_8_488_478_0 & i_8_488_482_0 & i_8_488_1265_0 & i_8_488_1768_0) | (~i_8_488_762_0 & ~i_8_488_768_0 & ~i_8_488_75_0 & ~i_8_488_482_0 & ~i_8_488_792_0 & i_8_488_831_0 & ~i_8_488_970_0 & ~i_8_488_1350_0 & ~i_8_488_2110_0))) | (~i_8_488_482_0 & ((~i_8_488_687_0 & i_8_488_732_0 & i_8_488_832_0) | (~i_8_488_343_0 & ~i_8_488_690_0 & ~i_8_488_710_0 & ~i_8_488_763_0 & ~i_8_488_796_0 & i_8_488_2138_0))) | (~i_8_488_760_0 & ((~i_8_488_343_0 & ~i_8_488_664_0 & ~i_8_488_770_0 & ((i_8_488_751_0 & ~i_8_488_762_0 & ~i_8_488_792_0 & ~i_8_488_1306_0 & ~i_8_488_1770_0 & ~i_8_488_1996_0) | (~i_8_488_347_0 & ~i_8_488_631_0 & ~i_8_488_710_0 & ~i_8_488_2170_0 & i_8_488_2171_0))) | (~i_8_488_620_0 & ~i_8_488_796_0 & i_8_488_841_0 & ~i_8_488_1056_0 & ~i_8_488_1158_0 & ~i_8_488_1329_0 & i_8_488_2136_0 & ~i_8_488_2208_0))) | (~i_8_488_619_0 & i_8_488_620_0 & i_8_488_653_0 & ~i_8_488_772_0 & ~i_8_488_2138_0) | (~i_8_488_525_0 & ~i_8_488_620_0 & i_8_488_732_0 & ~i_8_488_769_0 & ~i_8_488_2001_0 & ~i_8_488_2216_0) | (i_8_488_2170_0 & i_8_488_2216_0 & i_8_488_2224_0 & i_8_488_2273_0 & ~i_8_488_2289_0));
endmodule



// Benchmark "kernel_8_489" written by ABC on Sun Jul 19 10:11:39 2020

module kernel_8_489 ( 
    i_8_489_52_0, i_8_489_82_0, i_8_489_86_0, i_8_489_97_0, i_8_489_104_0,
    i_8_489_138_0, i_8_489_139_0, i_8_489_140_0, i_8_489_165_0,
    i_8_489_232_0, i_8_489_258_0, i_8_489_262_0, i_8_489_299_0,
    i_8_489_301_0, i_8_489_302_0, i_8_489_346_0, i_8_489_354_0,
    i_8_489_365_0, i_8_489_486_0, i_8_489_509_0, i_8_489_528_0,
    i_8_489_579_0, i_8_489_584_0, i_8_489_590_0, i_8_489_604_0,
    i_8_489_659_0, i_8_489_675_0, i_8_489_677_0, i_8_489_698_0,
    i_8_489_704_0, i_8_489_707_0, i_8_489_716_0, i_8_489_729_0,
    i_8_489_782_0, i_8_489_799_0, i_8_489_827_0, i_8_489_851_0,
    i_8_489_930_0, i_8_489_967_0, i_8_489_971_0, i_8_489_1034_0,
    i_8_489_1108_0, i_8_489_1112_0, i_8_489_1135_0, i_8_489_1157_0,
    i_8_489_1220_0, i_8_489_1224_0, i_8_489_1236_0, i_8_489_1256_0,
    i_8_489_1272_0, i_8_489_1285_0, i_8_489_1298_0, i_8_489_1319_0,
    i_8_489_1404_0, i_8_489_1441_0, i_8_489_1443_0, i_8_489_1465_0,
    i_8_489_1537_0, i_8_489_1544_0, i_8_489_1558_0, i_8_489_1615_0,
    i_8_489_1628_0, i_8_489_1632_0, i_8_489_1644_0, i_8_489_1651_0,
    i_8_489_1652_0, i_8_489_1653_0, i_8_489_1667_0, i_8_489_1691_0,
    i_8_489_1705_0, i_8_489_1709_0, i_8_489_1783_0, i_8_489_1784_0,
    i_8_489_1787_0, i_8_489_1796_0, i_8_489_1804_0, i_8_489_1807_0,
    i_8_489_1838_0, i_8_489_1841_0, i_8_489_1859_0, i_8_489_1877_0,
    i_8_489_1884_0, i_8_489_1938_0, i_8_489_1948_0, i_8_489_1968_0,
    i_8_489_1995_0, i_8_489_2026_0, i_8_489_2059_0, i_8_489_2110_0,
    i_8_489_2111_0, i_8_489_2114_0, i_8_489_2119_0, i_8_489_2133_0,
    i_8_489_2155_0, i_8_489_2177_0, i_8_489_2183_0, i_8_489_2192_0,
    i_8_489_2231_0, i_8_489_2273_0, i_8_489_2286_0,
    o_8_489_0_0  );
  input  i_8_489_52_0, i_8_489_82_0, i_8_489_86_0, i_8_489_97_0,
    i_8_489_104_0, i_8_489_138_0, i_8_489_139_0, i_8_489_140_0,
    i_8_489_165_0, i_8_489_232_0, i_8_489_258_0, i_8_489_262_0,
    i_8_489_299_0, i_8_489_301_0, i_8_489_302_0, i_8_489_346_0,
    i_8_489_354_0, i_8_489_365_0, i_8_489_486_0, i_8_489_509_0,
    i_8_489_528_0, i_8_489_579_0, i_8_489_584_0, i_8_489_590_0,
    i_8_489_604_0, i_8_489_659_0, i_8_489_675_0, i_8_489_677_0,
    i_8_489_698_0, i_8_489_704_0, i_8_489_707_0, i_8_489_716_0,
    i_8_489_729_0, i_8_489_782_0, i_8_489_799_0, i_8_489_827_0,
    i_8_489_851_0, i_8_489_930_0, i_8_489_967_0, i_8_489_971_0,
    i_8_489_1034_0, i_8_489_1108_0, i_8_489_1112_0, i_8_489_1135_0,
    i_8_489_1157_0, i_8_489_1220_0, i_8_489_1224_0, i_8_489_1236_0,
    i_8_489_1256_0, i_8_489_1272_0, i_8_489_1285_0, i_8_489_1298_0,
    i_8_489_1319_0, i_8_489_1404_0, i_8_489_1441_0, i_8_489_1443_0,
    i_8_489_1465_0, i_8_489_1537_0, i_8_489_1544_0, i_8_489_1558_0,
    i_8_489_1615_0, i_8_489_1628_0, i_8_489_1632_0, i_8_489_1644_0,
    i_8_489_1651_0, i_8_489_1652_0, i_8_489_1653_0, i_8_489_1667_0,
    i_8_489_1691_0, i_8_489_1705_0, i_8_489_1709_0, i_8_489_1783_0,
    i_8_489_1784_0, i_8_489_1787_0, i_8_489_1796_0, i_8_489_1804_0,
    i_8_489_1807_0, i_8_489_1838_0, i_8_489_1841_0, i_8_489_1859_0,
    i_8_489_1877_0, i_8_489_1884_0, i_8_489_1938_0, i_8_489_1948_0,
    i_8_489_1968_0, i_8_489_1995_0, i_8_489_2026_0, i_8_489_2059_0,
    i_8_489_2110_0, i_8_489_2111_0, i_8_489_2114_0, i_8_489_2119_0,
    i_8_489_2133_0, i_8_489_2155_0, i_8_489_2177_0, i_8_489_2183_0,
    i_8_489_2192_0, i_8_489_2231_0, i_8_489_2273_0, i_8_489_2286_0;
  output o_8_489_0_0;
  assign o_8_489_0_0 = 0;
endmodule



// Benchmark "kernel_8_490" written by ABC on Sun Jul 19 10:11:40 2020

module kernel_8_490 ( 
    i_8_490_7_0, i_8_490_16_0, i_8_490_23_0, i_8_490_41_0, i_8_490_50_0,
    i_8_490_107_0, i_8_490_131_0, i_8_490_143_0, i_8_490_167_0,
    i_8_490_257_0, i_8_490_283_0, i_8_490_287_0, i_8_490_296_0,
    i_8_490_365_0, i_8_490_382_0, i_8_490_454_0, i_8_490_458_0,
    i_8_490_489_0, i_8_490_490_0, i_8_490_524_0, i_8_490_587_0,
    i_8_490_605_0, i_8_490_614_0, i_8_490_650_0, i_8_490_653_0,
    i_8_490_670_0, i_8_490_676_0, i_8_490_709_0, i_8_490_730_0,
    i_8_490_733_0, i_8_490_769_0, i_8_490_805_0, i_8_490_809_0,
    i_8_490_814_0, i_8_490_841_0, i_8_490_851_0, i_8_490_932_0,
    i_8_490_968_0, i_8_490_1067_0, i_8_490_1072_0, i_8_490_1109_0,
    i_8_490_1139_0, i_8_490_1229_0, i_8_490_1241_0, i_8_490_1274_0,
    i_8_490_1283_0, i_8_490_1292_0, i_8_490_1301_0, i_8_490_1322_0,
    i_8_490_1333_0, i_8_490_1385_0, i_8_490_1468_0, i_8_490_1489_0,
    i_8_490_1491_0, i_8_490_1553_0, i_8_490_1561_0, i_8_490_1574_0,
    i_8_490_1588_0, i_8_490_1603_0, i_8_490_1610_0, i_8_490_1625_0,
    i_8_490_1627_0, i_8_490_1628_0, i_8_490_1630_0, i_8_490_1633_0,
    i_8_490_1672_0, i_8_490_1679_0, i_8_490_1693_0, i_8_490_1700_0,
    i_8_490_1703_0, i_8_490_1747_0, i_8_490_1774_0, i_8_490_1781_0,
    i_8_490_1783_0, i_8_490_1822_0, i_8_490_1841_0, i_8_490_1847_0,
    i_8_490_1850_0, i_8_490_1885_0, i_8_490_1903_0, i_8_490_1963_0,
    i_8_490_1979_0, i_8_490_1988_0, i_8_490_1996_0, i_8_490_1997_0,
    i_8_490_2029_0, i_8_490_2039_0, i_8_490_2114_0, i_8_490_2119_0,
    i_8_490_2120_0, i_8_490_2134_0, i_8_490_2135_0, i_8_490_2147_0,
    i_8_490_2156_0, i_8_490_2170_0, i_8_490_2183_0, i_8_490_2187_0,
    i_8_490_2225_0, i_8_490_2243_0, i_8_490_2249_0,
    o_8_490_0_0  );
  input  i_8_490_7_0, i_8_490_16_0, i_8_490_23_0, i_8_490_41_0,
    i_8_490_50_0, i_8_490_107_0, i_8_490_131_0, i_8_490_143_0,
    i_8_490_167_0, i_8_490_257_0, i_8_490_283_0, i_8_490_287_0,
    i_8_490_296_0, i_8_490_365_0, i_8_490_382_0, i_8_490_454_0,
    i_8_490_458_0, i_8_490_489_0, i_8_490_490_0, i_8_490_524_0,
    i_8_490_587_0, i_8_490_605_0, i_8_490_614_0, i_8_490_650_0,
    i_8_490_653_0, i_8_490_670_0, i_8_490_676_0, i_8_490_709_0,
    i_8_490_730_0, i_8_490_733_0, i_8_490_769_0, i_8_490_805_0,
    i_8_490_809_0, i_8_490_814_0, i_8_490_841_0, i_8_490_851_0,
    i_8_490_932_0, i_8_490_968_0, i_8_490_1067_0, i_8_490_1072_0,
    i_8_490_1109_0, i_8_490_1139_0, i_8_490_1229_0, i_8_490_1241_0,
    i_8_490_1274_0, i_8_490_1283_0, i_8_490_1292_0, i_8_490_1301_0,
    i_8_490_1322_0, i_8_490_1333_0, i_8_490_1385_0, i_8_490_1468_0,
    i_8_490_1489_0, i_8_490_1491_0, i_8_490_1553_0, i_8_490_1561_0,
    i_8_490_1574_0, i_8_490_1588_0, i_8_490_1603_0, i_8_490_1610_0,
    i_8_490_1625_0, i_8_490_1627_0, i_8_490_1628_0, i_8_490_1630_0,
    i_8_490_1633_0, i_8_490_1672_0, i_8_490_1679_0, i_8_490_1693_0,
    i_8_490_1700_0, i_8_490_1703_0, i_8_490_1747_0, i_8_490_1774_0,
    i_8_490_1781_0, i_8_490_1783_0, i_8_490_1822_0, i_8_490_1841_0,
    i_8_490_1847_0, i_8_490_1850_0, i_8_490_1885_0, i_8_490_1903_0,
    i_8_490_1963_0, i_8_490_1979_0, i_8_490_1988_0, i_8_490_1996_0,
    i_8_490_1997_0, i_8_490_2029_0, i_8_490_2039_0, i_8_490_2114_0,
    i_8_490_2119_0, i_8_490_2120_0, i_8_490_2134_0, i_8_490_2135_0,
    i_8_490_2147_0, i_8_490_2156_0, i_8_490_2170_0, i_8_490_2183_0,
    i_8_490_2187_0, i_8_490_2225_0, i_8_490_2243_0, i_8_490_2249_0;
  output o_8_490_0_0;
  assign o_8_490_0_0 = 0;
endmodule



// Benchmark "kernel_8_491" written by ABC on Sun Jul 19 10:11:41 2020

module kernel_8_491 ( 
    i_8_491_4_0, i_8_491_34_0, i_8_491_85_0, i_8_491_86_0, i_8_491_88_0,
    i_8_491_187_0, i_8_491_246_0, i_8_491_263_0, i_8_491_284_0,
    i_8_491_325_0, i_8_491_329_0, i_8_491_361_0, i_8_491_364_0,
    i_8_491_366_0, i_8_491_371_0, i_8_491_454_0, i_8_491_488_0,
    i_8_491_523_0, i_8_491_588_0, i_8_491_589_0, i_8_491_599_0,
    i_8_491_625_0, i_8_491_634_0, i_8_491_637_0, i_8_491_660_0,
    i_8_491_679_0, i_8_491_695_0, i_8_491_697_0, i_8_491_724_0,
    i_8_491_734_0, i_8_491_772_0, i_8_491_778_0, i_8_491_840_0,
    i_8_491_869_0, i_8_491_881_0, i_8_491_964_0, i_8_491_1020_0,
    i_8_491_1030_0, i_8_491_1110_0, i_8_491_1118_0, i_8_491_1190_0,
    i_8_491_1192_0, i_8_491_1227_0, i_8_491_1228_0, i_8_491_1255_0,
    i_8_491_1265_0, i_8_491_1282_0, i_8_491_1283_0, i_8_491_1285_0,
    i_8_491_1299_0, i_8_491_1317_0, i_8_491_1354_0, i_8_491_1355_0,
    i_8_491_1360_0, i_8_491_1373_0, i_8_491_1435_0, i_8_491_1446_0,
    i_8_491_1471_0, i_8_491_1472_0, i_8_491_1561_0, i_8_491_1624_0,
    i_8_491_1625_0, i_8_491_1668_0, i_8_491_1671_0, i_8_491_1696_0,
    i_8_491_1700_0, i_8_491_1703_0, i_8_491_1723_0, i_8_491_1729_0,
    i_8_491_1743_0, i_8_491_1751_0, i_8_491_1754_0, i_8_491_1768_0,
    i_8_491_1772_0, i_8_491_1777_0, i_8_491_1820_0, i_8_491_1822_0,
    i_8_491_1855_0, i_8_491_1857_0, i_8_491_1858_0, i_8_491_1859_0,
    i_8_491_1870_0, i_8_491_1884_0, i_8_491_1904_0, i_8_491_1912_0,
    i_8_491_1992_0, i_8_491_1993_0, i_8_491_2120_0, i_8_491_2145_0,
    i_8_491_2148_0, i_8_491_2155_0, i_8_491_2191_0, i_8_491_2224_0,
    i_8_491_2244_0, i_8_491_2248_0, i_8_491_2263_0, i_8_491_2272_0,
    i_8_491_2281_0, i_8_491_2288_0, i_8_491_2290_0,
    o_8_491_0_0  );
  input  i_8_491_4_0, i_8_491_34_0, i_8_491_85_0, i_8_491_86_0,
    i_8_491_88_0, i_8_491_187_0, i_8_491_246_0, i_8_491_263_0,
    i_8_491_284_0, i_8_491_325_0, i_8_491_329_0, i_8_491_361_0,
    i_8_491_364_0, i_8_491_366_0, i_8_491_371_0, i_8_491_454_0,
    i_8_491_488_0, i_8_491_523_0, i_8_491_588_0, i_8_491_589_0,
    i_8_491_599_0, i_8_491_625_0, i_8_491_634_0, i_8_491_637_0,
    i_8_491_660_0, i_8_491_679_0, i_8_491_695_0, i_8_491_697_0,
    i_8_491_724_0, i_8_491_734_0, i_8_491_772_0, i_8_491_778_0,
    i_8_491_840_0, i_8_491_869_0, i_8_491_881_0, i_8_491_964_0,
    i_8_491_1020_0, i_8_491_1030_0, i_8_491_1110_0, i_8_491_1118_0,
    i_8_491_1190_0, i_8_491_1192_0, i_8_491_1227_0, i_8_491_1228_0,
    i_8_491_1255_0, i_8_491_1265_0, i_8_491_1282_0, i_8_491_1283_0,
    i_8_491_1285_0, i_8_491_1299_0, i_8_491_1317_0, i_8_491_1354_0,
    i_8_491_1355_0, i_8_491_1360_0, i_8_491_1373_0, i_8_491_1435_0,
    i_8_491_1446_0, i_8_491_1471_0, i_8_491_1472_0, i_8_491_1561_0,
    i_8_491_1624_0, i_8_491_1625_0, i_8_491_1668_0, i_8_491_1671_0,
    i_8_491_1696_0, i_8_491_1700_0, i_8_491_1703_0, i_8_491_1723_0,
    i_8_491_1729_0, i_8_491_1743_0, i_8_491_1751_0, i_8_491_1754_0,
    i_8_491_1768_0, i_8_491_1772_0, i_8_491_1777_0, i_8_491_1820_0,
    i_8_491_1822_0, i_8_491_1855_0, i_8_491_1857_0, i_8_491_1858_0,
    i_8_491_1859_0, i_8_491_1870_0, i_8_491_1884_0, i_8_491_1904_0,
    i_8_491_1912_0, i_8_491_1992_0, i_8_491_1993_0, i_8_491_2120_0,
    i_8_491_2145_0, i_8_491_2148_0, i_8_491_2155_0, i_8_491_2191_0,
    i_8_491_2224_0, i_8_491_2244_0, i_8_491_2248_0, i_8_491_2263_0,
    i_8_491_2272_0, i_8_491_2281_0, i_8_491_2288_0, i_8_491_2290_0;
  output o_8_491_0_0;
  assign o_8_491_0_0 = 0;
endmodule



// Benchmark "kernel_8_492" written by ABC on Sun Jul 19 10:11:42 2020

module kernel_8_492 ( 
    i_8_492_9_0, i_8_492_39_0, i_8_492_67_0, i_8_492_72_0, i_8_492_114_0,
    i_8_492_138_0, i_8_492_220_0, i_8_492_225_0, i_8_492_226_0,
    i_8_492_260_0, i_8_492_268_0, i_8_492_414_0, i_8_492_418_0,
    i_8_492_421_0, i_8_492_426_0, i_8_492_469_0, i_8_492_504_0,
    i_8_492_507_0, i_8_492_525_0, i_8_492_526_0, i_8_492_532_0,
    i_8_492_552_0, i_8_492_568_0, i_8_492_571_0, i_8_492_576_0,
    i_8_492_596_0, i_8_492_599_0, i_8_492_657_0, i_8_492_658_0,
    i_8_492_693_0, i_8_492_703_0, i_8_492_705_0, i_8_492_748_0,
    i_8_492_751_0, i_8_492_816_0, i_8_492_829_0, i_8_492_837_0,
    i_8_492_840_0, i_8_492_849_0, i_8_492_874_0, i_8_492_975_0,
    i_8_492_976_0, i_8_492_982_0, i_8_492_1050_0, i_8_492_1110_0,
    i_8_492_1161_0, i_8_492_1234_0, i_8_492_1237_0, i_8_492_1285_0,
    i_8_492_1286_0, i_8_492_1297_0, i_8_492_1300_0, i_8_492_1314_0,
    i_8_492_1315_0, i_8_492_1323_0, i_8_492_1350_0, i_8_492_1354_0,
    i_8_492_1362_0, i_8_492_1395_0, i_8_492_1432_0, i_8_492_1461_0,
    i_8_492_1462_0, i_8_492_1470_0, i_8_492_1476_0, i_8_492_1477_0,
    i_8_492_1481_0, i_8_492_1484_0, i_8_492_1489_0, i_8_492_1512_0,
    i_8_492_1524_0, i_8_492_1555_0, i_8_492_1621_0, i_8_492_1630_0,
    i_8_492_1669_0, i_8_492_1729_0, i_8_492_1734_0, i_8_492_1746_0,
    i_8_492_1747_0, i_8_492_1748_0, i_8_492_1764_0, i_8_492_1773_0,
    i_8_492_1777_0, i_8_492_1791_0, i_8_492_1794_0, i_8_492_1800_0,
    i_8_492_1819_0, i_8_492_1857_0, i_8_492_1893_0, i_8_492_1900_0,
    i_8_492_2053_0, i_8_492_2056_0, i_8_492_2083_0, i_8_492_2098_0,
    i_8_492_2125_0, i_8_492_2142_0, i_8_492_2152_0, i_8_492_2155_0,
    i_8_492_2242_0, i_8_492_2269_0, i_8_492_2270_0,
    o_8_492_0_0  );
  input  i_8_492_9_0, i_8_492_39_0, i_8_492_67_0, i_8_492_72_0,
    i_8_492_114_0, i_8_492_138_0, i_8_492_220_0, i_8_492_225_0,
    i_8_492_226_0, i_8_492_260_0, i_8_492_268_0, i_8_492_414_0,
    i_8_492_418_0, i_8_492_421_0, i_8_492_426_0, i_8_492_469_0,
    i_8_492_504_0, i_8_492_507_0, i_8_492_525_0, i_8_492_526_0,
    i_8_492_532_0, i_8_492_552_0, i_8_492_568_0, i_8_492_571_0,
    i_8_492_576_0, i_8_492_596_0, i_8_492_599_0, i_8_492_657_0,
    i_8_492_658_0, i_8_492_693_0, i_8_492_703_0, i_8_492_705_0,
    i_8_492_748_0, i_8_492_751_0, i_8_492_816_0, i_8_492_829_0,
    i_8_492_837_0, i_8_492_840_0, i_8_492_849_0, i_8_492_874_0,
    i_8_492_975_0, i_8_492_976_0, i_8_492_982_0, i_8_492_1050_0,
    i_8_492_1110_0, i_8_492_1161_0, i_8_492_1234_0, i_8_492_1237_0,
    i_8_492_1285_0, i_8_492_1286_0, i_8_492_1297_0, i_8_492_1300_0,
    i_8_492_1314_0, i_8_492_1315_0, i_8_492_1323_0, i_8_492_1350_0,
    i_8_492_1354_0, i_8_492_1362_0, i_8_492_1395_0, i_8_492_1432_0,
    i_8_492_1461_0, i_8_492_1462_0, i_8_492_1470_0, i_8_492_1476_0,
    i_8_492_1477_0, i_8_492_1481_0, i_8_492_1484_0, i_8_492_1489_0,
    i_8_492_1512_0, i_8_492_1524_0, i_8_492_1555_0, i_8_492_1621_0,
    i_8_492_1630_0, i_8_492_1669_0, i_8_492_1729_0, i_8_492_1734_0,
    i_8_492_1746_0, i_8_492_1747_0, i_8_492_1748_0, i_8_492_1764_0,
    i_8_492_1773_0, i_8_492_1777_0, i_8_492_1791_0, i_8_492_1794_0,
    i_8_492_1800_0, i_8_492_1819_0, i_8_492_1857_0, i_8_492_1893_0,
    i_8_492_1900_0, i_8_492_2053_0, i_8_492_2056_0, i_8_492_2083_0,
    i_8_492_2098_0, i_8_492_2125_0, i_8_492_2142_0, i_8_492_2152_0,
    i_8_492_2155_0, i_8_492_2242_0, i_8_492_2269_0, i_8_492_2270_0;
  output o_8_492_0_0;
  assign o_8_492_0_0 = 0;
endmodule



// Benchmark "kernel_8_493" written by ABC on Sun Jul 19 10:11:43 2020

module kernel_8_493 ( 
    i_8_493_30_0, i_8_493_33_0, i_8_493_80_0, i_8_493_86_0, i_8_493_88_0,
    i_8_493_142_0, i_8_493_166_0, i_8_493_190_0, i_8_493_258_0,
    i_8_493_265_0, i_8_493_266_0, i_8_493_268_0, i_8_493_269_0,
    i_8_493_296_0, i_8_493_301_0, i_8_493_302_0, i_8_493_304_0,
    i_8_493_337_0, i_8_493_385_0, i_8_493_454_0, i_8_493_455_0,
    i_8_493_470_0, i_8_493_474_0, i_8_493_485_0, i_8_493_520_0,
    i_8_493_525_0, i_8_493_528_0, i_8_493_554_0, i_8_493_556_0,
    i_8_493_571_0, i_8_493_592_0, i_8_493_593_0, i_8_493_607_0,
    i_8_493_609_0, i_8_493_627_0, i_8_493_634_0, i_8_493_638_0,
    i_8_493_664_0, i_8_493_674_0, i_8_493_680_0, i_8_493_693_0,
    i_8_493_719_0, i_8_493_727_0, i_8_493_841_0, i_8_493_880_0,
    i_8_493_1016_0, i_8_493_1030_0, i_8_493_1033_0, i_8_493_1115_0,
    i_8_493_1124_0, i_8_493_1131_0, i_8_493_1237_0, i_8_493_1241_0,
    i_8_493_1285_0, i_8_493_1286_0, i_8_493_1306_0, i_8_493_1349_0,
    i_8_493_1437_0, i_8_493_1453_0, i_8_493_1456_0, i_8_493_1457_0,
    i_8_493_1474_0, i_8_493_1535_0, i_8_493_1546_0, i_8_493_1556_0,
    i_8_493_1579_0, i_8_493_1601_0, i_8_493_1672_0, i_8_493_1677_0,
    i_8_493_1678_0, i_8_493_1706_0, i_8_493_1709_0, i_8_493_1742_0,
    i_8_493_1745_0, i_8_493_1808_0, i_8_493_1834_0, i_8_493_1844_0,
    i_8_493_1861_0, i_8_493_1906_0, i_8_493_1921_0, i_8_493_1922_0,
    i_8_493_1952_0, i_8_493_1969_0, i_8_493_1970_0, i_8_493_1996_0,
    i_8_493_2014_0, i_8_493_2023_0, i_8_493_2024_0, i_8_493_2111_0,
    i_8_493_2113_0, i_8_493_2122_0, i_8_493_2131_0, i_8_493_2132_0,
    i_8_493_2137_0, i_8_493_2156_0, i_8_493_2194_0, i_8_493_2195_0,
    i_8_493_2239_0, i_8_493_2276_0, i_8_493_2293_0,
    o_8_493_0_0  );
  input  i_8_493_30_0, i_8_493_33_0, i_8_493_80_0, i_8_493_86_0,
    i_8_493_88_0, i_8_493_142_0, i_8_493_166_0, i_8_493_190_0,
    i_8_493_258_0, i_8_493_265_0, i_8_493_266_0, i_8_493_268_0,
    i_8_493_269_0, i_8_493_296_0, i_8_493_301_0, i_8_493_302_0,
    i_8_493_304_0, i_8_493_337_0, i_8_493_385_0, i_8_493_454_0,
    i_8_493_455_0, i_8_493_470_0, i_8_493_474_0, i_8_493_485_0,
    i_8_493_520_0, i_8_493_525_0, i_8_493_528_0, i_8_493_554_0,
    i_8_493_556_0, i_8_493_571_0, i_8_493_592_0, i_8_493_593_0,
    i_8_493_607_0, i_8_493_609_0, i_8_493_627_0, i_8_493_634_0,
    i_8_493_638_0, i_8_493_664_0, i_8_493_674_0, i_8_493_680_0,
    i_8_493_693_0, i_8_493_719_0, i_8_493_727_0, i_8_493_841_0,
    i_8_493_880_0, i_8_493_1016_0, i_8_493_1030_0, i_8_493_1033_0,
    i_8_493_1115_0, i_8_493_1124_0, i_8_493_1131_0, i_8_493_1237_0,
    i_8_493_1241_0, i_8_493_1285_0, i_8_493_1286_0, i_8_493_1306_0,
    i_8_493_1349_0, i_8_493_1437_0, i_8_493_1453_0, i_8_493_1456_0,
    i_8_493_1457_0, i_8_493_1474_0, i_8_493_1535_0, i_8_493_1546_0,
    i_8_493_1556_0, i_8_493_1579_0, i_8_493_1601_0, i_8_493_1672_0,
    i_8_493_1677_0, i_8_493_1678_0, i_8_493_1706_0, i_8_493_1709_0,
    i_8_493_1742_0, i_8_493_1745_0, i_8_493_1808_0, i_8_493_1834_0,
    i_8_493_1844_0, i_8_493_1861_0, i_8_493_1906_0, i_8_493_1921_0,
    i_8_493_1922_0, i_8_493_1952_0, i_8_493_1969_0, i_8_493_1970_0,
    i_8_493_1996_0, i_8_493_2014_0, i_8_493_2023_0, i_8_493_2024_0,
    i_8_493_2111_0, i_8_493_2113_0, i_8_493_2122_0, i_8_493_2131_0,
    i_8_493_2132_0, i_8_493_2137_0, i_8_493_2156_0, i_8_493_2194_0,
    i_8_493_2195_0, i_8_493_2239_0, i_8_493_2276_0, i_8_493_2293_0;
  output o_8_493_0_0;
  assign o_8_493_0_0 = 0;
endmodule



// Benchmark "kernel_8_494" written by ABC on Sun Jul 19 10:11:44 2020

module kernel_8_494 ( 
    i_8_494_20_0, i_8_494_25_0, i_8_494_47_0, i_8_494_56_0, i_8_494_101_0,
    i_8_494_104_0, i_8_494_140_0, i_8_494_230_0, i_8_494_233_0,
    i_8_494_256_0, i_8_494_281_0, i_8_494_301_0, i_8_494_317_0,
    i_8_494_380_0, i_8_494_382_0, i_8_494_419_0, i_8_494_486_0,
    i_8_494_530_0, i_8_494_536_0, i_8_494_587_0, i_8_494_596_0,
    i_8_494_614_0, i_8_494_640_0, i_8_494_650_0, i_8_494_652_0,
    i_8_494_695_0, i_8_494_696_0, i_8_494_704_0, i_8_494_830_0,
    i_8_494_838_0, i_8_494_848_0, i_8_494_857_0, i_8_494_866_0,
    i_8_494_875_0, i_8_494_877_0, i_8_494_881_0, i_8_494_884_0,
    i_8_494_941_0, i_8_494_969_0, i_8_494_974_0, i_8_494_1103_0,
    i_8_494_1136_0, i_8_494_1139_0, i_8_494_1145_0, i_8_494_1202_0,
    i_8_494_1260_0, i_8_494_1297_0, i_8_494_1304_0, i_8_494_1317_0,
    i_8_494_1334_0, i_8_494_1342_0, i_8_494_1343_0, i_8_494_1351_0,
    i_8_494_1352_0, i_8_494_1355_0, i_8_494_1357_0, i_8_494_1397_0,
    i_8_494_1432_0, i_8_494_1433_0, i_8_494_1468_0, i_8_494_1487_0,
    i_8_494_1507_0, i_8_494_1525_0, i_8_494_1547_0, i_8_494_1561_0,
    i_8_494_1564_0, i_8_494_1604_0, i_8_494_1612_0, i_8_494_1688_0,
    i_8_494_1707_0, i_8_494_1715_0, i_8_494_1721_0, i_8_494_1746_0,
    i_8_494_1750_0, i_8_494_1753_0, i_8_494_1754_0, i_8_494_1756_0,
    i_8_494_1766_0, i_8_494_1768_0, i_8_494_1775_0, i_8_494_1785_0,
    i_8_494_1786_0, i_8_494_1792_0, i_8_494_1814_0, i_8_494_1823_0,
    i_8_494_1864_0, i_8_494_1883_0, i_8_494_1945_0, i_8_494_1964_0,
    i_8_494_1984_0, i_8_494_1991_0, i_8_494_1997_0, i_8_494_2054_0,
    i_8_494_2135_0, i_8_494_2153_0, i_8_494_2192_0, i_8_494_2225_0,
    i_8_494_2227_0, i_8_494_2234_0, i_8_494_2247_0,
    o_8_494_0_0  );
  input  i_8_494_20_0, i_8_494_25_0, i_8_494_47_0, i_8_494_56_0,
    i_8_494_101_0, i_8_494_104_0, i_8_494_140_0, i_8_494_230_0,
    i_8_494_233_0, i_8_494_256_0, i_8_494_281_0, i_8_494_301_0,
    i_8_494_317_0, i_8_494_380_0, i_8_494_382_0, i_8_494_419_0,
    i_8_494_486_0, i_8_494_530_0, i_8_494_536_0, i_8_494_587_0,
    i_8_494_596_0, i_8_494_614_0, i_8_494_640_0, i_8_494_650_0,
    i_8_494_652_0, i_8_494_695_0, i_8_494_696_0, i_8_494_704_0,
    i_8_494_830_0, i_8_494_838_0, i_8_494_848_0, i_8_494_857_0,
    i_8_494_866_0, i_8_494_875_0, i_8_494_877_0, i_8_494_881_0,
    i_8_494_884_0, i_8_494_941_0, i_8_494_969_0, i_8_494_974_0,
    i_8_494_1103_0, i_8_494_1136_0, i_8_494_1139_0, i_8_494_1145_0,
    i_8_494_1202_0, i_8_494_1260_0, i_8_494_1297_0, i_8_494_1304_0,
    i_8_494_1317_0, i_8_494_1334_0, i_8_494_1342_0, i_8_494_1343_0,
    i_8_494_1351_0, i_8_494_1352_0, i_8_494_1355_0, i_8_494_1357_0,
    i_8_494_1397_0, i_8_494_1432_0, i_8_494_1433_0, i_8_494_1468_0,
    i_8_494_1487_0, i_8_494_1507_0, i_8_494_1525_0, i_8_494_1547_0,
    i_8_494_1561_0, i_8_494_1564_0, i_8_494_1604_0, i_8_494_1612_0,
    i_8_494_1688_0, i_8_494_1707_0, i_8_494_1715_0, i_8_494_1721_0,
    i_8_494_1746_0, i_8_494_1750_0, i_8_494_1753_0, i_8_494_1754_0,
    i_8_494_1756_0, i_8_494_1766_0, i_8_494_1768_0, i_8_494_1775_0,
    i_8_494_1785_0, i_8_494_1786_0, i_8_494_1792_0, i_8_494_1814_0,
    i_8_494_1823_0, i_8_494_1864_0, i_8_494_1883_0, i_8_494_1945_0,
    i_8_494_1964_0, i_8_494_1984_0, i_8_494_1991_0, i_8_494_1997_0,
    i_8_494_2054_0, i_8_494_2135_0, i_8_494_2153_0, i_8_494_2192_0,
    i_8_494_2225_0, i_8_494_2227_0, i_8_494_2234_0, i_8_494_2247_0;
  output o_8_494_0_0;
  assign o_8_494_0_0 = 0;
endmodule



// Benchmark "kernel_8_495" written by ABC on Sun Jul 19 10:11:45 2020

module kernel_8_495 ( 
    i_8_495_34_0, i_8_495_58_0, i_8_495_72_0, i_8_495_77_0, i_8_495_79_0,
    i_8_495_80_0, i_8_495_120_0, i_8_495_143_0, i_8_495_151_0,
    i_8_495_230_0, i_8_495_400_0, i_8_495_422_0, i_8_495_426_0,
    i_8_495_429_0, i_8_495_431_0, i_8_495_457_0, i_8_495_522_0,
    i_8_495_538_0, i_8_495_539_0, i_8_495_556_0, i_8_495_561_0,
    i_8_495_611_0, i_8_495_613_0, i_8_495_630_0, i_8_495_634_0,
    i_8_495_638_0, i_8_495_646_0, i_8_495_655_0, i_8_495_660_0,
    i_8_495_661_0, i_8_495_673_0, i_8_495_703_0, i_8_495_704_0,
    i_8_495_707_0, i_8_495_719_0, i_8_495_749_0, i_8_495_752_0,
    i_8_495_755_0, i_8_495_836_0, i_8_495_873_0, i_8_495_921_0,
    i_8_495_967_0, i_8_495_970_0, i_8_495_976_0, i_8_495_994_0,
    i_8_495_1013_0, i_8_495_1015_0, i_8_495_1073_0, i_8_495_1075_0,
    i_8_495_1102_0, i_8_495_1133_0, i_8_495_1266_0, i_8_495_1300_0,
    i_8_495_1305_0, i_8_495_1337_0, i_8_495_1357_0, i_8_495_1399_0,
    i_8_495_1400_0, i_8_495_1436_0, i_8_495_1438_0, i_8_495_1439_0,
    i_8_495_1456_0, i_8_495_1480_0, i_8_495_1489_0, i_8_495_1490_0,
    i_8_495_1528_0, i_8_495_1542_0, i_8_495_1543_0, i_8_495_1544_0,
    i_8_495_1572_0, i_8_495_1651_0, i_8_495_1653_0, i_8_495_1677_0,
    i_8_495_1691_0, i_8_495_1700_0, i_8_495_1703_0, i_8_495_1707_0,
    i_8_495_1754_0, i_8_495_1770_0, i_8_495_1771_0, i_8_495_1774_0,
    i_8_495_1794_0, i_8_495_1795_0, i_8_495_1810_0, i_8_495_1823_0,
    i_8_495_1843_0, i_8_495_1891_0, i_8_495_1912_0, i_8_495_1951_0,
    i_8_495_1952_0, i_8_495_1957_0, i_8_495_1993_0, i_8_495_1996_0,
    i_8_495_2131_0, i_8_495_2148_0, i_8_495_2214_0, i_8_495_2215_0,
    i_8_495_2234_0, i_8_495_2287_0, i_8_495_2299_0,
    o_8_495_0_0  );
  input  i_8_495_34_0, i_8_495_58_0, i_8_495_72_0, i_8_495_77_0,
    i_8_495_79_0, i_8_495_80_0, i_8_495_120_0, i_8_495_143_0,
    i_8_495_151_0, i_8_495_230_0, i_8_495_400_0, i_8_495_422_0,
    i_8_495_426_0, i_8_495_429_0, i_8_495_431_0, i_8_495_457_0,
    i_8_495_522_0, i_8_495_538_0, i_8_495_539_0, i_8_495_556_0,
    i_8_495_561_0, i_8_495_611_0, i_8_495_613_0, i_8_495_630_0,
    i_8_495_634_0, i_8_495_638_0, i_8_495_646_0, i_8_495_655_0,
    i_8_495_660_0, i_8_495_661_0, i_8_495_673_0, i_8_495_703_0,
    i_8_495_704_0, i_8_495_707_0, i_8_495_719_0, i_8_495_749_0,
    i_8_495_752_0, i_8_495_755_0, i_8_495_836_0, i_8_495_873_0,
    i_8_495_921_0, i_8_495_967_0, i_8_495_970_0, i_8_495_976_0,
    i_8_495_994_0, i_8_495_1013_0, i_8_495_1015_0, i_8_495_1073_0,
    i_8_495_1075_0, i_8_495_1102_0, i_8_495_1133_0, i_8_495_1266_0,
    i_8_495_1300_0, i_8_495_1305_0, i_8_495_1337_0, i_8_495_1357_0,
    i_8_495_1399_0, i_8_495_1400_0, i_8_495_1436_0, i_8_495_1438_0,
    i_8_495_1439_0, i_8_495_1456_0, i_8_495_1480_0, i_8_495_1489_0,
    i_8_495_1490_0, i_8_495_1528_0, i_8_495_1542_0, i_8_495_1543_0,
    i_8_495_1544_0, i_8_495_1572_0, i_8_495_1651_0, i_8_495_1653_0,
    i_8_495_1677_0, i_8_495_1691_0, i_8_495_1700_0, i_8_495_1703_0,
    i_8_495_1707_0, i_8_495_1754_0, i_8_495_1770_0, i_8_495_1771_0,
    i_8_495_1774_0, i_8_495_1794_0, i_8_495_1795_0, i_8_495_1810_0,
    i_8_495_1823_0, i_8_495_1843_0, i_8_495_1891_0, i_8_495_1912_0,
    i_8_495_1951_0, i_8_495_1952_0, i_8_495_1957_0, i_8_495_1993_0,
    i_8_495_1996_0, i_8_495_2131_0, i_8_495_2148_0, i_8_495_2214_0,
    i_8_495_2215_0, i_8_495_2234_0, i_8_495_2287_0, i_8_495_2299_0;
  output o_8_495_0_0;
  assign o_8_495_0_0 = 0;
endmodule



// Benchmark "kernel_8_496" written by ABC on Sun Jul 19 10:11:46 2020

module kernel_8_496 ( 
    i_8_496_34_0, i_8_496_52_0, i_8_496_58_0, i_8_496_88_0, i_8_496_93_0,
    i_8_496_96_0, i_8_496_97_0, i_8_496_140_0, i_8_496_141_0,
    i_8_496_186_0, i_8_496_232_0, i_8_496_233_0, i_8_496_255_0,
    i_8_496_304_0, i_8_496_374_0, i_8_496_424_0, i_8_496_428_0,
    i_8_496_440_0, i_8_496_455_0, i_8_496_475_0, i_8_496_482_0,
    i_8_496_483_0, i_8_496_485_0, i_8_496_499_0, i_8_496_526_0,
    i_8_496_527_0, i_8_496_556_0, i_8_496_602_0, i_8_496_627_0,
    i_8_496_661_0, i_8_496_662_0, i_8_496_674_0, i_8_496_680_0,
    i_8_496_688_0, i_8_496_706_0, i_8_496_733_0, i_8_496_759_0,
    i_8_496_762_0, i_8_496_763_0, i_8_496_781_0, i_8_496_782_0,
    i_8_496_799_0, i_8_496_800_0, i_8_496_805_0, i_8_496_850_0,
    i_8_496_966_0, i_8_496_1050_0, i_8_496_1051_0, i_8_496_1071_0,
    i_8_496_1074_0, i_8_496_1075_0, i_8_496_1119_0, i_8_496_1120_0,
    i_8_496_1122_0, i_8_496_1136_0, i_8_496_1148_0, i_8_496_1191_0,
    i_8_496_1273_0, i_8_496_1299_0, i_8_496_1305_0, i_8_496_1324_0,
    i_8_496_1326_0, i_8_496_1390_0, i_8_496_1437_0, i_8_496_1450_0,
    i_8_496_1470_0, i_8_496_1506_0, i_8_496_1509_0, i_8_496_1533_0,
    i_8_496_1537_0, i_8_496_1545_0, i_8_496_1563_0, i_8_496_1570_0,
    i_8_496_1632_0, i_8_496_1652_0, i_8_496_1681_0, i_8_496_1682_0,
    i_8_496_1684_0, i_8_496_1751_0, i_8_496_1759_0, i_8_496_1763_0,
    i_8_496_1807_0, i_8_496_1811_0, i_8_496_1821_0, i_8_496_1876_0,
    i_8_496_1951_0, i_8_496_1982_0, i_8_496_1993_0, i_8_496_2003_0,
    i_8_496_2029_0, i_8_496_2055_0, i_8_496_2092_0, i_8_496_2093_0,
    i_8_496_2108_0, i_8_496_2146_0, i_8_496_2150_0, i_8_496_2210_0,
    i_8_496_2214_0, i_8_496_2215_0, i_8_496_2216_0,
    o_8_496_0_0  );
  input  i_8_496_34_0, i_8_496_52_0, i_8_496_58_0, i_8_496_88_0,
    i_8_496_93_0, i_8_496_96_0, i_8_496_97_0, i_8_496_140_0, i_8_496_141_0,
    i_8_496_186_0, i_8_496_232_0, i_8_496_233_0, i_8_496_255_0,
    i_8_496_304_0, i_8_496_374_0, i_8_496_424_0, i_8_496_428_0,
    i_8_496_440_0, i_8_496_455_0, i_8_496_475_0, i_8_496_482_0,
    i_8_496_483_0, i_8_496_485_0, i_8_496_499_0, i_8_496_526_0,
    i_8_496_527_0, i_8_496_556_0, i_8_496_602_0, i_8_496_627_0,
    i_8_496_661_0, i_8_496_662_0, i_8_496_674_0, i_8_496_680_0,
    i_8_496_688_0, i_8_496_706_0, i_8_496_733_0, i_8_496_759_0,
    i_8_496_762_0, i_8_496_763_0, i_8_496_781_0, i_8_496_782_0,
    i_8_496_799_0, i_8_496_800_0, i_8_496_805_0, i_8_496_850_0,
    i_8_496_966_0, i_8_496_1050_0, i_8_496_1051_0, i_8_496_1071_0,
    i_8_496_1074_0, i_8_496_1075_0, i_8_496_1119_0, i_8_496_1120_0,
    i_8_496_1122_0, i_8_496_1136_0, i_8_496_1148_0, i_8_496_1191_0,
    i_8_496_1273_0, i_8_496_1299_0, i_8_496_1305_0, i_8_496_1324_0,
    i_8_496_1326_0, i_8_496_1390_0, i_8_496_1437_0, i_8_496_1450_0,
    i_8_496_1470_0, i_8_496_1506_0, i_8_496_1509_0, i_8_496_1533_0,
    i_8_496_1537_0, i_8_496_1545_0, i_8_496_1563_0, i_8_496_1570_0,
    i_8_496_1632_0, i_8_496_1652_0, i_8_496_1681_0, i_8_496_1682_0,
    i_8_496_1684_0, i_8_496_1751_0, i_8_496_1759_0, i_8_496_1763_0,
    i_8_496_1807_0, i_8_496_1811_0, i_8_496_1821_0, i_8_496_1876_0,
    i_8_496_1951_0, i_8_496_1982_0, i_8_496_1993_0, i_8_496_2003_0,
    i_8_496_2029_0, i_8_496_2055_0, i_8_496_2092_0, i_8_496_2093_0,
    i_8_496_2108_0, i_8_496_2146_0, i_8_496_2150_0, i_8_496_2210_0,
    i_8_496_2214_0, i_8_496_2215_0, i_8_496_2216_0;
  output o_8_496_0_0;
  assign o_8_496_0_0 = 0;
endmodule



// Benchmark "kernel_8_497" written by ABC on Sun Jul 19 10:11:47 2020

module kernel_8_497 ( 
    i_8_497_3_0, i_8_497_31_0, i_8_497_82_0, i_8_497_103_0, i_8_497_165_0,
    i_8_497_208_0, i_8_497_246_0, i_8_497_248_0, i_8_497_282_0,
    i_8_497_298_0, i_8_497_328_0, i_8_497_436_0, i_8_497_450_0,
    i_8_497_486_0, i_8_497_489_0, i_8_497_550_0, i_8_497_588_0,
    i_8_497_589_0, i_8_497_597_0, i_8_497_622_0, i_8_497_633_0,
    i_8_497_634_0, i_8_497_642_0, i_8_497_643_0, i_8_497_651_0,
    i_8_497_669_0, i_8_497_670_0, i_8_497_672_0, i_8_497_678_0,
    i_8_497_703_0, i_8_497_721_0, i_8_497_732_0, i_8_497_733_0,
    i_8_497_754_0, i_8_497_778_0, i_8_497_785_0, i_8_497_817_0,
    i_8_497_826_0, i_8_497_831_0, i_8_497_874_0, i_8_497_886_0,
    i_8_497_931_0, i_8_497_958_0, i_8_497_963_0, i_8_497_970_0,
    i_8_497_973_0, i_8_497_976_0, i_8_497_985_0, i_8_497_991_0,
    i_8_497_1071_0, i_8_497_1072_0, i_8_497_1074_0, i_8_497_1130_0,
    i_8_497_1183_0, i_8_497_1236_0, i_8_497_1263_0, i_8_497_1270_0,
    i_8_497_1284_0, i_8_497_1285_0, i_8_497_1299_0, i_8_497_1357_0,
    i_8_497_1359_0, i_8_497_1362_0, i_8_497_1390_0, i_8_497_1439_0,
    i_8_497_1443_0, i_8_497_1470_0, i_8_497_1570_0, i_8_497_1575_0,
    i_8_497_1576_0, i_8_497_1588_0, i_8_497_1596_0, i_8_497_1632_0,
    i_8_497_1633_0, i_8_497_1677_0, i_8_497_1696_0, i_8_497_1699_0,
    i_8_497_1746_0, i_8_497_1747_0, i_8_497_1749_0, i_8_497_1768_0,
    i_8_497_1818_0, i_8_497_1822_0, i_8_497_1846_0, i_8_497_1848_0,
    i_8_497_1854_0, i_8_497_1855_0, i_8_497_1867_0, i_8_497_2010_0,
    i_8_497_2040_0, i_8_497_2080_0, i_8_497_2119_0, i_8_497_2134_0,
    i_8_497_2137_0, i_8_497_2147_0, i_8_497_2167_0, i_8_497_2169_0,
    i_8_497_2209_0, i_8_497_2214_0, i_8_497_2242_0,
    o_8_497_0_0  );
  input  i_8_497_3_0, i_8_497_31_0, i_8_497_82_0, i_8_497_103_0,
    i_8_497_165_0, i_8_497_208_0, i_8_497_246_0, i_8_497_248_0,
    i_8_497_282_0, i_8_497_298_0, i_8_497_328_0, i_8_497_436_0,
    i_8_497_450_0, i_8_497_486_0, i_8_497_489_0, i_8_497_550_0,
    i_8_497_588_0, i_8_497_589_0, i_8_497_597_0, i_8_497_622_0,
    i_8_497_633_0, i_8_497_634_0, i_8_497_642_0, i_8_497_643_0,
    i_8_497_651_0, i_8_497_669_0, i_8_497_670_0, i_8_497_672_0,
    i_8_497_678_0, i_8_497_703_0, i_8_497_721_0, i_8_497_732_0,
    i_8_497_733_0, i_8_497_754_0, i_8_497_778_0, i_8_497_785_0,
    i_8_497_817_0, i_8_497_826_0, i_8_497_831_0, i_8_497_874_0,
    i_8_497_886_0, i_8_497_931_0, i_8_497_958_0, i_8_497_963_0,
    i_8_497_970_0, i_8_497_973_0, i_8_497_976_0, i_8_497_985_0,
    i_8_497_991_0, i_8_497_1071_0, i_8_497_1072_0, i_8_497_1074_0,
    i_8_497_1130_0, i_8_497_1183_0, i_8_497_1236_0, i_8_497_1263_0,
    i_8_497_1270_0, i_8_497_1284_0, i_8_497_1285_0, i_8_497_1299_0,
    i_8_497_1357_0, i_8_497_1359_0, i_8_497_1362_0, i_8_497_1390_0,
    i_8_497_1439_0, i_8_497_1443_0, i_8_497_1470_0, i_8_497_1570_0,
    i_8_497_1575_0, i_8_497_1576_0, i_8_497_1588_0, i_8_497_1596_0,
    i_8_497_1632_0, i_8_497_1633_0, i_8_497_1677_0, i_8_497_1696_0,
    i_8_497_1699_0, i_8_497_1746_0, i_8_497_1747_0, i_8_497_1749_0,
    i_8_497_1768_0, i_8_497_1818_0, i_8_497_1822_0, i_8_497_1846_0,
    i_8_497_1848_0, i_8_497_1854_0, i_8_497_1855_0, i_8_497_1867_0,
    i_8_497_2010_0, i_8_497_2040_0, i_8_497_2080_0, i_8_497_2119_0,
    i_8_497_2134_0, i_8_497_2137_0, i_8_497_2147_0, i_8_497_2167_0,
    i_8_497_2169_0, i_8_497_2209_0, i_8_497_2214_0, i_8_497_2242_0;
  output o_8_497_0_0;
  assign o_8_497_0_0 = 0;
endmodule



// Benchmark "kernel_8_498" written by ABC on Sun Jul 19 10:11:48 2020

module kernel_8_498 ( 
    i_8_498_31_0, i_8_498_35_0, i_8_498_36_0, i_8_498_89_0, i_8_498_110_0,
    i_8_498_140_0, i_8_498_256_0, i_8_498_273_0, i_8_498_301_0,
    i_8_498_329_0, i_8_498_345_0, i_8_498_346_0, i_8_498_375_0,
    i_8_498_377_0, i_8_498_418_0, i_8_498_434_0, i_8_498_451_0,
    i_8_498_454_0, i_8_498_463_0, i_8_498_511_0, i_8_498_528_0,
    i_8_498_529_0, i_8_498_530_0, i_8_498_553_0, i_8_498_554_0,
    i_8_498_589_0, i_8_498_595_0, i_8_498_611_0, i_8_498_620_0,
    i_8_498_670_0, i_8_498_671_0, i_8_498_673_0, i_8_498_709_0,
    i_8_498_716_0, i_8_498_772_0, i_8_498_780_0, i_8_498_781_0,
    i_8_498_796_0, i_8_498_824_0, i_8_498_865_0, i_8_498_975_0,
    i_8_498_984_0, i_8_498_985_0, i_8_498_1014_0, i_8_498_1120_0,
    i_8_498_1131_0, i_8_498_1132_0, i_8_498_1158_0, i_8_498_1159_0,
    i_8_498_1218_0, i_8_498_1228_0, i_8_498_1249_0, i_8_498_1258_0,
    i_8_498_1268_0, i_8_498_1306_0, i_8_498_1307_0, i_8_498_1310_0,
    i_8_498_1387_0, i_8_498_1390_0, i_8_498_1397_0, i_8_498_1453_0,
    i_8_498_1470_0, i_8_498_1532_0, i_8_498_1533_0, i_8_498_1534_0,
    i_8_498_1540_0, i_8_498_1556_0, i_8_498_1597_0, i_8_498_1598_0,
    i_8_498_1607_0, i_8_498_1629_0, i_8_498_1669_0, i_8_498_1684_0,
    i_8_498_1762_0, i_8_498_1763_0, i_8_498_1808_0, i_8_498_1821_0,
    i_8_498_1840_0, i_8_498_1870_0, i_8_498_1874_0, i_8_498_1907_0,
    i_8_498_1948_0, i_8_498_1975_0, i_8_498_2019_0, i_8_498_2044_0,
    i_8_498_2065_0, i_8_498_2105_0, i_8_498_2126_0, i_8_498_2128_0,
    i_8_498_2140_0, i_8_498_2154_0, i_8_498_2172_0, i_8_498_2183_0,
    i_8_498_2188_0, i_8_498_2190_0, i_8_498_2191_0, i_8_498_2213_0,
    i_8_498_2215_0, i_8_498_2272_0, i_8_498_2289_0,
    o_8_498_0_0  );
  input  i_8_498_31_0, i_8_498_35_0, i_8_498_36_0, i_8_498_89_0,
    i_8_498_110_0, i_8_498_140_0, i_8_498_256_0, i_8_498_273_0,
    i_8_498_301_0, i_8_498_329_0, i_8_498_345_0, i_8_498_346_0,
    i_8_498_375_0, i_8_498_377_0, i_8_498_418_0, i_8_498_434_0,
    i_8_498_451_0, i_8_498_454_0, i_8_498_463_0, i_8_498_511_0,
    i_8_498_528_0, i_8_498_529_0, i_8_498_530_0, i_8_498_553_0,
    i_8_498_554_0, i_8_498_589_0, i_8_498_595_0, i_8_498_611_0,
    i_8_498_620_0, i_8_498_670_0, i_8_498_671_0, i_8_498_673_0,
    i_8_498_709_0, i_8_498_716_0, i_8_498_772_0, i_8_498_780_0,
    i_8_498_781_0, i_8_498_796_0, i_8_498_824_0, i_8_498_865_0,
    i_8_498_975_0, i_8_498_984_0, i_8_498_985_0, i_8_498_1014_0,
    i_8_498_1120_0, i_8_498_1131_0, i_8_498_1132_0, i_8_498_1158_0,
    i_8_498_1159_0, i_8_498_1218_0, i_8_498_1228_0, i_8_498_1249_0,
    i_8_498_1258_0, i_8_498_1268_0, i_8_498_1306_0, i_8_498_1307_0,
    i_8_498_1310_0, i_8_498_1387_0, i_8_498_1390_0, i_8_498_1397_0,
    i_8_498_1453_0, i_8_498_1470_0, i_8_498_1532_0, i_8_498_1533_0,
    i_8_498_1534_0, i_8_498_1540_0, i_8_498_1556_0, i_8_498_1597_0,
    i_8_498_1598_0, i_8_498_1607_0, i_8_498_1629_0, i_8_498_1669_0,
    i_8_498_1684_0, i_8_498_1762_0, i_8_498_1763_0, i_8_498_1808_0,
    i_8_498_1821_0, i_8_498_1840_0, i_8_498_1870_0, i_8_498_1874_0,
    i_8_498_1907_0, i_8_498_1948_0, i_8_498_1975_0, i_8_498_2019_0,
    i_8_498_2044_0, i_8_498_2065_0, i_8_498_2105_0, i_8_498_2126_0,
    i_8_498_2128_0, i_8_498_2140_0, i_8_498_2154_0, i_8_498_2172_0,
    i_8_498_2183_0, i_8_498_2188_0, i_8_498_2190_0, i_8_498_2191_0,
    i_8_498_2213_0, i_8_498_2215_0, i_8_498_2272_0, i_8_498_2289_0;
  output o_8_498_0_0;
  assign o_8_498_0_0 = 0;
endmodule



// Benchmark "kernel_8_499" written by ABC on Sun Jul 19 10:11:49 2020

module kernel_8_499 ( 
    i_8_499_52_0, i_8_499_75_0, i_8_499_86_0, i_8_499_116_0, i_8_499_131_0,
    i_8_499_190_0, i_8_499_191_0, i_8_499_193_0, i_8_499_258_0,
    i_8_499_274_0, i_8_499_307_0, i_8_499_318_0, i_8_499_320_0,
    i_8_499_360_0, i_8_499_362_0, i_8_499_365_0, i_8_499_453_0,
    i_8_499_499_0, i_8_499_522_0, i_8_499_523_0, i_8_499_525_0,
    i_8_499_526_0, i_8_499_527_0, i_8_499_528_0, i_8_499_588_0,
    i_8_499_590_0, i_8_499_631_0, i_8_499_639_0, i_8_499_657_0,
    i_8_499_659_0, i_8_499_660_0, i_8_499_675_0, i_8_499_676_0,
    i_8_499_677_0, i_8_499_678_0, i_8_499_712_0, i_8_499_716_0,
    i_8_499_719_0, i_8_499_760_0, i_8_499_761_0, i_8_499_837_0,
    i_8_499_838_0, i_8_499_840_0, i_8_499_881_0, i_8_499_968_0,
    i_8_499_970_0, i_8_499_974_0, i_8_499_990_0, i_8_499_994_0,
    i_8_499_997_0, i_8_499_1054_0, i_8_499_1128_0, i_8_499_1188_0,
    i_8_499_1224_0, i_8_499_1228_0, i_8_499_1229_0, i_8_499_1264_0,
    i_8_499_1267_0, i_8_499_1281_0, i_8_499_1282_0, i_8_499_1285_0,
    i_8_499_1319_0, i_8_499_1337_0, i_8_499_1404_0, i_8_499_1405_0,
    i_8_499_1436_0, i_8_499_1453_0, i_8_499_1532_0, i_8_499_1533_0,
    i_8_499_1534_0, i_8_499_1535_0, i_8_499_1593_0, i_8_499_1598_0,
    i_8_499_1633_0, i_8_499_1638_0, i_8_499_1650_0, i_8_499_1656_0,
    i_8_499_1658_0, i_8_499_1660_0, i_8_499_1661_0, i_8_499_1679_0,
    i_8_499_1783_0, i_8_499_1784_0, i_8_499_1821_0, i_8_499_1822_0,
    i_8_499_1872_0, i_8_499_1903_0, i_8_499_1975_0, i_8_499_2010_0,
    i_8_499_2012_0, i_8_499_2052_0, i_8_499_2090_0, i_8_499_2092_0,
    i_8_499_2093_0, i_8_499_2133_0, i_8_499_2174_0, i_8_499_2216_0,
    i_8_499_2244_0, i_8_499_2246_0, i_8_499_2247_0,
    o_8_499_0_0  );
  input  i_8_499_52_0, i_8_499_75_0, i_8_499_86_0, i_8_499_116_0,
    i_8_499_131_0, i_8_499_190_0, i_8_499_191_0, i_8_499_193_0,
    i_8_499_258_0, i_8_499_274_0, i_8_499_307_0, i_8_499_318_0,
    i_8_499_320_0, i_8_499_360_0, i_8_499_362_0, i_8_499_365_0,
    i_8_499_453_0, i_8_499_499_0, i_8_499_522_0, i_8_499_523_0,
    i_8_499_525_0, i_8_499_526_0, i_8_499_527_0, i_8_499_528_0,
    i_8_499_588_0, i_8_499_590_0, i_8_499_631_0, i_8_499_639_0,
    i_8_499_657_0, i_8_499_659_0, i_8_499_660_0, i_8_499_675_0,
    i_8_499_676_0, i_8_499_677_0, i_8_499_678_0, i_8_499_712_0,
    i_8_499_716_0, i_8_499_719_0, i_8_499_760_0, i_8_499_761_0,
    i_8_499_837_0, i_8_499_838_0, i_8_499_840_0, i_8_499_881_0,
    i_8_499_968_0, i_8_499_970_0, i_8_499_974_0, i_8_499_990_0,
    i_8_499_994_0, i_8_499_997_0, i_8_499_1054_0, i_8_499_1128_0,
    i_8_499_1188_0, i_8_499_1224_0, i_8_499_1228_0, i_8_499_1229_0,
    i_8_499_1264_0, i_8_499_1267_0, i_8_499_1281_0, i_8_499_1282_0,
    i_8_499_1285_0, i_8_499_1319_0, i_8_499_1337_0, i_8_499_1404_0,
    i_8_499_1405_0, i_8_499_1436_0, i_8_499_1453_0, i_8_499_1532_0,
    i_8_499_1533_0, i_8_499_1534_0, i_8_499_1535_0, i_8_499_1593_0,
    i_8_499_1598_0, i_8_499_1633_0, i_8_499_1638_0, i_8_499_1650_0,
    i_8_499_1656_0, i_8_499_1658_0, i_8_499_1660_0, i_8_499_1661_0,
    i_8_499_1679_0, i_8_499_1783_0, i_8_499_1784_0, i_8_499_1821_0,
    i_8_499_1822_0, i_8_499_1872_0, i_8_499_1903_0, i_8_499_1975_0,
    i_8_499_2010_0, i_8_499_2012_0, i_8_499_2052_0, i_8_499_2090_0,
    i_8_499_2092_0, i_8_499_2093_0, i_8_499_2133_0, i_8_499_2174_0,
    i_8_499_2216_0, i_8_499_2244_0, i_8_499_2246_0, i_8_499_2247_0;
  output o_8_499_0_0;
  assign o_8_499_0_0 = ~((~i_8_499_881_0 & ((~i_8_499_1337_0 & ((~i_8_499_52_0 & ((i_8_499_307_0 & ~i_8_499_678_0 & ~i_8_499_968_0 & ~i_8_499_1821_0 & ~i_8_499_2052_0) | (i_8_499_86_0 & ~i_8_499_362_0 & ~i_8_499_676_0 & ~i_8_499_838_0 & ~i_8_499_1267_0 & ~i_8_499_2244_0))) | (~i_8_499_116_0 & ~i_8_499_453_0 & ~i_8_499_499_0 & ~i_8_499_660_0 & ~i_8_499_677_0 & ~i_8_499_968_0 & ~i_8_499_1128_0 & ~i_8_499_1228_0 & i_8_499_1822_0 & ~i_8_499_2133_0 & ~i_8_499_2244_0 & ~i_8_499_2247_0))) | (~i_8_499_362_0 & ((~i_8_499_191_0 & ~i_8_499_590_0 & ~i_8_499_660_0 & ~i_8_499_1267_0 & ~i_8_499_1319_0 & i_8_499_2216_0) | (~i_8_499_318_0 & ~i_8_499_677_0 & i_8_499_1054_0 & i_8_499_1404_0 & ~i_8_499_2133_0 & ~i_8_499_2247_0))) | (~i_8_499_116_0 & ~i_8_499_190_0 & ~i_8_499_526_0 & ~i_8_499_678_0 & ~i_8_499_760_0 & ~i_8_499_968_0 & ~i_8_499_1228_0 & ~i_8_499_1285_0 & i_8_499_1436_0 & i_8_499_1679_0 & ~i_8_499_2052_0) | (i_8_499_86_0 & ~i_8_499_631_0 & ~i_8_499_837_0 & ~i_8_499_974_0 & ~i_8_499_1229_0 & i_8_499_1282_0 & ~i_8_499_2246_0))) | (~i_8_499_453_0 & ((~i_8_499_52_0 & ((~i_8_499_499_0 & ~i_8_499_523_0 & ~i_8_499_631_0 & ~i_8_499_675_0 & ~i_8_499_678_0 & ~i_8_499_968_0 & ~i_8_499_1598_0 & i_8_499_2092_0) | (i_8_499_528_0 & ~i_8_499_588_0 & i_8_499_1264_0 & ~i_8_499_2244_0))) | (~i_8_499_116_0 & ~i_8_499_258_0 & ((i_8_499_193_0 & i_8_499_528_0 & ~i_8_499_970_0 & ~i_8_499_1281_0) | (~i_8_499_365_0 & ~i_8_499_639_0 & ~i_8_499_675_0 & ~i_8_499_1229_0 & ~i_8_499_1267_0 & i_8_499_1404_0))) | (~i_8_499_131_0 & ((~i_8_499_193_0 & ~i_8_499_660_0 & ~i_8_499_838_0 & i_8_499_994_0 & ~i_8_499_1264_0 & ~i_8_499_1282_0 & ~i_8_499_1679_0) | (~i_8_499_307_0 & ~i_8_499_320_0 & ~i_8_499_588_0 & ~i_8_499_590_0 & ~i_8_499_676_0 & ~i_8_499_997_0 & ~i_8_499_1229_0 & i_8_499_1319_0 & ~i_8_499_1337_0 & ~i_8_499_1532_0 & ~i_8_499_1534_0 & ~i_8_499_1821_0 & ~i_8_499_2092_0 & ~i_8_499_2244_0 & ~i_8_499_2246_0))) | (i_8_499_193_0 & ~i_8_499_1264_0 & ~i_8_499_1282_0 & ((~i_8_499_588_0 & ~i_8_499_631_0 & ~i_8_499_660_0 & ~i_8_499_1228_0 & i_8_499_1822_0) | (~i_8_499_75_0 & ~i_8_499_678_0 & ~i_8_499_837_0 & ~i_8_499_840_0 & ~i_8_499_970_0 & ~i_8_499_997_0 & ~i_8_499_1822_0 & ~i_8_499_2133_0))) | (i_8_499_525_0 & ((~i_8_499_320_0 & ~i_8_499_590_0 & ~i_8_499_678_0 & ~i_8_499_1285_0 & i_8_499_1533_0) | (i_8_499_526_0 & ~i_8_499_840_0 & ~i_8_499_968_0 & ~i_8_499_1224_0 & ~i_8_499_2247_0))) | (~i_8_499_660_0 & ~i_8_499_838_0 & ~i_8_499_526_0 & i_8_499_528_0 & ~i_8_499_968_0 & ~i_8_499_1285_0 & ~i_8_499_1650_0 & ~i_8_499_1822_0) | (~i_8_499_676_0 & ~i_8_499_1337_0 & i_8_499_2092_0 & i_8_499_2093_0))) | (~i_8_499_75_0 & i_8_499_1535_0 & ((~i_8_499_590_0 & ~i_8_499_677_0 & ~i_8_499_1281_0 & ~i_8_499_1436_0) | (~i_8_499_320_0 & ~i_8_499_659_0 & ~i_8_499_675_0 & ~i_8_499_676_0 & ~i_8_499_970_0 & ~i_8_499_2133_0))) | (~i_8_499_2247_0 & ((~i_8_499_1285_0 & ((~i_8_499_52_0 & ((~i_8_499_258_0 & ~i_8_499_320_0 & ~i_8_499_365_0 & i_8_499_525_0 & ~i_8_499_590_0 & ~i_8_499_657_0 & ~i_8_499_760_0 & ~i_8_499_1633_0 & ~i_8_499_1784_0) | (i_8_499_190_0 & ~i_8_499_526_0 & ~i_8_499_588_0 & ~i_8_499_639_0 & ~i_8_499_660_0 & ~i_8_499_675_0 & ~i_8_499_1224_0 & ~i_8_499_1282_0 & ~i_8_499_1453_0 & ~i_8_499_1821_0 & ~i_8_499_2244_0 & ~i_8_499_2246_0))) | (~i_8_499_190_0 & ~i_8_499_840_0 & ~i_8_499_1282_0 & ~i_8_499_1650_0 & ((~i_8_499_258_0 & ~i_8_499_362_0 & ~i_8_499_659_0 & ~i_8_499_968_0 & ~i_8_499_1264_0 & ~i_8_499_1436_0 & ~i_8_499_1453_0 & ~i_8_499_1821_0 & ~i_8_499_2092_0 & ~i_8_499_2133_0) | (i_8_499_193_0 & ~i_8_499_526_0 & ~i_8_499_1281_0 & ~i_8_499_1822_0 & ~i_8_499_2246_0))))) | (~i_8_499_1228_0 & ((~i_8_499_677_0 & ~i_8_499_1319_0 & ((~i_8_499_522_0 & ~i_8_499_639_0 & ~i_8_499_712_0 & ~i_8_499_970_0 & ~i_8_499_1337_0 & i_8_499_1534_0 & ~i_8_499_1535_0 & ~i_8_499_2092_0) | (~i_8_499_116_0 & ~i_8_499_590_0 & ~i_8_499_974_0 & i_8_499_997_0 & ~i_8_499_1188_0 & ~i_8_499_1229_0 & ~i_8_499_1264_0 & ~i_8_499_1404_0 & ~i_8_499_1633_0 & ~i_8_499_1821_0 & ~i_8_499_2244_0))) | (~i_8_499_974_0 & ((~i_8_499_660_0 & ~i_8_499_1224_0 & ~i_8_499_1229_0 & i_8_499_1638_0) | (~i_8_499_318_0 & ~i_8_499_360_0 & ~i_8_499_588_0 & ~i_8_499_970_0 & i_8_499_1054_0 & ~i_8_499_1128_0 & ~i_8_499_1656_0 & ~i_8_499_2093_0 & ~i_8_499_2244_0))))) | (i_8_499_760_0 & i_8_499_761_0) | (~i_8_499_52_0 & i_8_499_274_0 & ~i_8_499_675_0 & ~i_8_499_840_0 & i_8_499_1281_0 & ~i_8_499_1319_0 & ~i_8_499_1337_0 & ~i_8_499_1679_0 & ~i_8_499_2010_0) | (i_8_499_131_0 & ~i_8_499_193_0 & ~i_8_499_365_0 & ~i_8_499_526_0 & ~i_8_499_712_0 & ~i_8_499_970_0 & ~i_8_499_1822_0 & ~i_8_499_2216_0 & ~i_8_499_2246_0))) | (~i_8_499_193_0 & ((~i_8_499_52_0 & i_8_499_522_0 & ~i_8_499_590_0 & ~i_8_499_639_0 & ~i_8_499_676_0 & ~i_8_499_837_0 & ~i_8_499_968_0 & ~i_8_499_970_0 & ~i_8_499_1224_0 & ~i_8_499_1229_0 & ~i_8_499_1453_0) | (~i_8_499_631_0 & ~i_8_499_675_0 & ~i_8_499_116_0 & ~i_8_499_258_0 & ~i_8_499_678_0 & ~i_8_499_1264_0 & i_8_499_1650_0 & i_8_499_1822_0 & ~i_8_499_2133_0))) | (~i_8_499_258_0 & ((~i_8_499_52_0 & i_8_499_525_0 & ~i_8_499_631_0 & ~i_8_499_1337_0 & i_8_499_1453_0) | (~i_8_499_318_0 & ~i_8_499_659_0 & ~i_8_499_970_0 & ~i_8_499_974_0 & i_8_499_1188_0 & ~i_8_499_1436_0 & ~i_8_499_1656_0 & ~i_8_499_2092_0 & ~i_8_499_2244_0))) | (i_8_499_522_0 & ((~i_8_499_588_0 & ~i_8_499_676_0 & ~i_8_499_677_0 & ~i_8_499_678_0 & i_8_499_1224_0) | (~i_8_499_52_0 & ~i_8_499_1224_0 & i_8_499_1534_0 & ~i_8_499_2244_0))) | (~i_8_499_525_0 & ((~i_8_499_116_0 & i_8_499_527_0 & ~i_8_499_659_0 & ~i_8_499_677_0 & ~i_8_499_837_0 & ~i_8_499_997_0 & ~i_8_499_1436_0) | (i_8_499_526_0 & ~i_8_499_676_0 & ~i_8_499_712_0 & ~i_8_499_838_0 & ~i_8_499_840_0 & ~i_8_499_968_0 & ~i_8_499_1285_0 & ~i_8_499_2244_0 & ~i_8_499_2246_0))) | (i_8_499_526_0 & ((~i_8_499_365_0 & i_8_499_523_0 & ~i_8_499_590_0 & ~i_8_499_840_0 & ~i_8_499_1224_0) | (i_8_499_525_0 & ~i_8_499_675_0 & ~i_8_499_968_0 & ~i_8_499_970_0 & ~i_8_499_1281_0 & ~i_8_499_1282_0 & ~i_8_499_1453_0))) | (~i_8_499_52_0 & ((~i_8_499_320_0 & ((~i_8_499_116_0 & i_8_499_527_0 & ~i_8_499_676_0 & ~i_8_499_974_0 & ~i_8_499_1264_0 & ~i_8_499_1267_0 & ~i_8_499_1282_0 & ~i_8_499_1650_0) | (~i_8_499_631_0 & ~i_8_499_677_0 & ~i_8_499_719_0 & ~i_8_499_1679_0 & i_8_499_2012_0 & ~i_8_499_2244_0))) | (~i_8_499_86_0 & i_8_499_527_0 & ~i_8_499_677_0 & ~i_8_499_760_0 & ~i_8_499_1319_0 & ~i_8_499_1337_0 & ~i_8_499_2174_0 & ~i_8_499_2244_0))) | (~i_8_499_678_0 & ((~i_8_499_677_0 & ((~i_8_499_116_0 & ((~i_8_499_639_0 & ~i_8_499_716_0 & ~i_8_499_970_0 & ~i_8_499_1282_0 & ~i_8_499_1650_0 & i_8_499_2090_0) | (~i_8_499_365_0 & ~i_8_499_675_0 & ~i_8_499_838_0 & ~i_8_499_1405_0 & ~i_8_499_1436_0 & ~i_8_499_1633_0 & i_8_499_1679_0 & ~i_8_499_1903_0 & ~i_8_499_2246_0))) | (~i_8_499_320_0 & i_8_499_719_0 & ~i_8_499_840_0 & i_8_499_1453_0 & ~i_8_499_2174_0))) | (~i_8_499_365_0 & ~i_8_499_1282_0 & i_8_499_1532_0))) | (~i_8_499_660_0 & ((~i_8_499_318_0 & ~i_8_499_1224_0 & i_8_499_1281_0 & ~i_8_499_1285_0 & i_8_499_1656_0) | (~i_8_499_365_0 & ~i_8_499_837_0 & ~i_8_499_838_0 & ~i_8_499_970_0 & ~i_8_499_1282_0 & i_8_499_1285_0 & i_8_499_1821_0))) | (~i_8_499_1282_0 & ((~i_8_499_1267_0 & i_8_499_1650_0 & i_8_499_1660_0) | (~i_8_499_659_0 & ~i_8_499_837_0 & ~i_8_499_1285_0 & ~i_8_499_1337_0 & i_8_499_2093_0))) | (~i_8_499_659_0 & ((i_8_499_719_0 & ~i_8_499_1228_0 & ~i_8_499_1281_0 & ~i_8_499_1285_0 & ~i_8_499_1319_0) | (i_8_499_1534_0 & ~i_8_499_1679_0 & ~i_8_499_1784_0 & ~i_8_499_1822_0 & ~i_8_499_2133_0 & ~i_8_499_2216_0))) | (~i_8_499_1285_0 & ((i_8_499_528_0 & ~i_8_499_657_0 & ~i_8_499_712_0 & ~i_8_499_968_0 & i_8_499_997_0 & ~i_8_499_1650_0) | (~i_8_499_499_0 & ~i_8_499_590_0 & ~i_8_499_1224_0 & ~i_8_499_1229_0 & ~i_8_499_1319_0 & i_8_499_1453_0 & ~i_8_499_1821_0 & ~i_8_499_1822_0 & ~i_8_499_2012_0 & ~i_8_499_2174_0 & ~i_8_499_2246_0))) | (i_8_499_2092_0 & i_8_499_2093_0 & i_8_499_2174_0 & ~i_8_499_2246_0) | (i_8_499_1660_0 & ~i_8_499_1822_0 & ~i_8_499_2133_0 & ~i_8_499_2174_0 & ~i_8_499_2244_0));
endmodule



// Benchmark "kernel_8_500" written by ABC on Sun Jul 19 10:11:50 2020

module kernel_8_500 ( 
    i_8_500_17_0, i_8_500_24_0, i_8_500_52_0, i_8_500_112_0, i_8_500_190_0,
    i_8_500_202_0, i_8_500_205_0, i_8_500_229_0, i_8_500_356_0,
    i_8_500_374_0, i_8_500_382_0, i_8_500_472_0, i_8_500_473_0,
    i_8_500_482_0, i_8_500_483_0, i_8_500_484_0, i_8_500_485_0,
    i_8_500_490_0, i_8_500_499_0, i_8_500_530_0, i_8_500_535_0,
    i_8_500_544_0, i_8_500_553_0, i_8_500_593_0, i_8_500_598_0,
    i_8_500_599_0, i_8_500_607_0, i_8_500_652_0, i_8_500_707_0,
    i_8_500_755_0, i_8_500_786_0, i_8_500_795_0, i_8_500_830_0,
    i_8_500_848_0, i_8_500_904_0, i_8_500_944_0, i_8_500_959_0,
    i_8_500_1001_0, i_8_500_1002_0, i_8_500_1012_0, i_8_500_1030_0,
    i_8_500_1135_0, i_8_500_1183_0, i_8_500_1184_0, i_8_500_1228_0,
    i_8_500_1294_0, i_8_500_1306_0, i_8_500_1340_0, i_8_500_1343_0,
    i_8_500_1346_0, i_8_500_1390_0, i_8_500_1433_0, i_8_500_1480_0,
    i_8_500_1525_0, i_8_500_1526_0, i_8_500_1562_0, i_8_500_1565_0,
    i_8_500_1600_0, i_8_500_1610_0, i_8_500_1639_0, i_8_500_1666_0,
    i_8_500_1671_0, i_8_500_1678_0, i_8_500_1687_0, i_8_500_1693_0,
    i_8_500_1694_0, i_8_500_1697_0, i_8_500_1705_0, i_8_500_1708_0,
    i_8_500_1724_0, i_8_500_1727_0, i_8_500_1751_0, i_8_500_1777_0,
    i_8_500_1806_0, i_8_500_1822_0, i_8_500_1826_0, i_8_500_1829_0,
    i_8_500_1858_0, i_8_500_1897_0, i_8_500_1921_0, i_8_500_1975_0,
    i_8_500_2003_0, i_8_500_2035_0, i_8_500_2038_0, i_8_500_2056_0,
    i_8_500_2093_0, i_8_500_2107_0, i_8_500_2125_0, i_8_500_2126_0,
    i_8_500_2134_0, i_8_500_2147_0, i_8_500_2183_0, i_8_500_2215_0,
    i_8_500_2236_0, i_8_500_2238_0, i_8_500_2242_0, i_8_500_2261_0,
    i_8_500_2272_0, i_8_500_2285_0, i_8_500_2294_0,
    o_8_500_0_0  );
  input  i_8_500_17_0, i_8_500_24_0, i_8_500_52_0, i_8_500_112_0,
    i_8_500_190_0, i_8_500_202_0, i_8_500_205_0, i_8_500_229_0,
    i_8_500_356_0, i_8_500_374_0, i_8_500_382_0, i_8_500_472_0,
    i_8_500_473_0, i_8_500_482_0, i_8_500_483_0, i_8_500_484_0,
    i_8_500_485_0, i_8_500_490_0, i_8_500_499_0, i_8_500_530_0,
    i_8_500_535_0, i_8_500_544_0, i_8_500_553_0, i_8_500_593_0,
    i_8_500_598_0, i_8_500_599_0, i_8_500_607_0, i_8_500_652_0,
    i_8_500_707_0, i_8_500_755_0, i_8_500_786_0, i_8_500_795_0,
    i_8_500_830_0, i_8_500_848_0, i_8_500_904_0, i_8_500_944_0,
    i_8_500_959_0, i_8_500_1001_0, i_8_500_1002_0, i_8_500_1012_0,
    i_8_500_1030_0, i_8_500_1135_0, i_8_500_1183_0, i_8_500_1184_0,
    i_8_500_1228_0, i_8_500_1294_0, i_8_500_1306_0, i_8_500_1340_0,
    i_8_500_1343_0, i_8_500_1346_0, i_8_500_1390_0, i_8_500_1433_0,
    i_8_500_1480_0, i_8_500_1525_0, i_8_500_1526_0, i_8_500_1562_0,
    i_8_500_1565_0, i_8_500_1600_0, i_8_500_1610_0, i_8_500_1639_0,
    i_8_500_1666_0, i_8_500_1671_0, i_8_500_1678_0, i_8_500_1687_0,
    i_8_500_1693_0, i_8_500_1694_0, i_8_500_1697_0, i_8_500_1705_0,
    i_8_500_1708_0, i_8_500_1724_0, i_8_500_1727_0, i_8_500_1751_0,
    i_8_500_1777_0, i_8_500_1806_0, i_8_500_1822_0, i_8_500_1826_0,
    i_8_500_1829_0, i_8_500_1858_0, i_8_500_1897_0, i_8_500_1921_0,
    i_8_500_1975_0, i_8_500_2003_0, i_8_500_2035_0, i_8_500_2038_0,
    i_8_500_2056_0, i_8_500_2093_0, i_8_500_2107_0, i_8_500_2125_0,
    i_8_500_2126_0, i_8_500_2134_0, i_8_500_2147_0, i_8_500_2183_0,
    i_8_500_2215_0, i_8_500_2236_0, i_8_500_2238_0, i_8_500_2242_0,
    i_8_500_2261_0, i_8_500_2272_0, i_8_500_2285_0, i_8_500_2294_0;
  output o_8_500_0_0;
  assign o_8_500_0_0 = 0;
endmodule



// Benchmark "kernel_8_501" written by ABC on Sun Jul 19 10:11:51 2020

module kernel_8_501 ( 
    i_8_501_30_0, i_8_501_31_0, i_8_501_40_0, i_8_501_41_0, i_8_501_43_0,
    i_8_501_47_0, i_8_501_54_0, i_8_501_55_0, i_8_501_58_0, i_8_501_67_0,
    i_8_501_73_0, i_8_501_100_0, i_8_501_159_0, i_8_501_162_0,
    i_8_501_191_0, i_8_501_217_0, i_8_501_297_0, i_8_501_324_0,
    i_8_501_361_0, i_8_501_363_0, i_8_501_364_0, i_8_501_382_0,
    i_8_501_423_0, i_8_501_424_0, i_8_501_501_0, i_8_501_550_0,
    i_8_501_577_0, i_8_501_586_0, i_8_501_589_0, i_8_501_634_0,
    i_8_501_658_0, i_8_501_675_0, i_8_501_703_0, i_8_501_705_0,
    i_8_501_706_0, i_8_501_751_0, i_8_501_832_0, i_8_501_837_0,
    i_8_501_840_0, i_8_501_843_0, i_8_501_846_0, i_8_501_847_0,
    i_8_501_855_0, i_8_501_856_0, i_8_501_874_0, i_8_501_882_0,
    i_8_501_894_0, i_8_501_895_0, i_8_501_1039_0, i_8_501_1112_0,
    i_8_501_1126_0, i_8_501_1129_0, i_8_501_1135_0, i_8_501_1143_0,
    i_8_501_1263_0, i_8_501_1264_0, i_8_501_1267_0, i_8_501_1279_0,
    i_8_501_1371_0, i_8_501_1407_0, i_8_501_1424_0, i_8_501_1438_0,
    i_8_501_1467_0, i_8_501_1468_0, i_8_501_1524_0, i_8_501_1629_0,
    i_8_501_1630_0, i_8_501_1651_0, i_8_501_1675_0, i_8_501_1677_0,
    i_8_501_1678_0, i_8_501_1705_0, i_8_501_1713_0, i_8_501_1756_0,
    i_8_501_1759_0, i_8_501_1767_0, i_8_501_1777_0, i_8_501_1786_0,
    i_8_501_1807_0, i_8_501_1862_0, i_8_501_1869_0, i_8_501_1899_0,
    i_8_501_1900_0, i_8_501_1970_0, i_8_501_1993_0, i_8_501_2052_0,
    i_8_501_2098_0, i_8_501_2106_0, i_8_501_2142_0, i_8_501_2146_0,
    i_8_501_2148_0, i_8_501_2149_0, i_8_501_2226_0, i_8_501_2232_0,
    i_8_501_2233_0, i_8_501_2235_0, i_8_501_2247_0, i_8_501_2248_0,
    i_8_501_2259_0, i_8_501_2262_0,
    o_8_501_0_0  );
  input  i_8_501_30_0, i_8_501_31_0, i_8_501_40_0, i_8_501_41_0,
    i_8_501_43_0, i_8_501_47_0, i_8_501_54_0, i_8_501_55_0, i_8_501_58_0,
    i_8_501_67_0, i_8_501_73_0, i_8_501_100_0, i_8_501_159_0,
    i_8_501_162_0, i_8_501_191_0, i_8_501_217_0, i_8_501_297_0,
    i_8_501_324_0, i_8_501_361_0, i_8_501_363_0, i_8_501_364_0,
    i_8_501_382_0, i_8_501_423_0, i_8_501_424_0, i_8_501_501_0,
    i_8_501_550_0, i_8_501_577_0, i_8_501_586_0, i_8_501_589_0,
    i_8_501_634_0, i_8_501_658_0, i_8_501_675_0, i_8_501_703_0,
    i_8_501_705_0, i_8_501_706_0, i_8_501_751_0, i_8_501_832_0,
    i_8_501_837_0, i_8_501_840_0, i_8_501_843_0, i_8_501_846_0,
    i_8_501_847_0, i_8_501_855_0, i_8_501_856_0, i_8_501_874_0,
    i_8_501_882_0, i_8_501_894_0, i_8_501_895_0, i_8_501_1039_0,
    i_8_501_1112_0, i_8_501_1126_0, i_8_501_1129_0, i_8_501_1135_0,
    i_8_501_1143_0, i_8_501_1263_0, i_8_501_1264_0, i_8_501_1267_0,
    i_8_501_1279_0, i_8_501_1371_0, i_8_501_1407_0, i_8_501_1424_0,
    i_8_501_1438_0, i_8_501_1467_0, i_8_501_1468_0, i_8_501_1524_0,
    i_8_501_1629_0, i_8_501_1630_0, i_8_501_1651_0, i_8_501_1675_0,
    i_8_501_1677_0, i_8_501_1678_0, i_8_501_1705_0, i_8_501_1713_0,
    i_8_501_1756_0, i_8_501_1759_0, i_8_501_1767_0, i_8_501_1777_0,
    i_8_501_1786_0, i_8_501_1807_0, i_8_501_1862_0, i_8_501_1869_0,
    i_8_501_1899_0, i_8_501_1900_0, i_8_501_1970_0, i_8_501_1993_0,
    i_8_501_2052_0, i_8_501_2098_0, i_8_501_2106_0, i_8_501_2142_0,
    i_8_501_2146_0, i_8_501_2148_0, i_8_501_2149_0, i_8_501_2226_0,
    i_8_501_2232_0, i_8_501_2233_0, i_8_501_2235_0, i_8_501_2247_0,
    i_8_501_2248_0, i_8_501_2259_0, i_8_501_2262_0;
  output o_8_501_0_0;
  assign o_8_501_0_0 = 0;
endmodule



// Benchmark "kernel_8_502" written by ABC on Sun Jul 19 10:11:52 2020

module kernel_8_502 ( 
    i_8_502_15_0, i_8_502_17_0, i_8_502_44_0, i_8_502_60_0, i_8_502_67_0,
    i_8_502_71_0, i_8_502_142_0, i_8_502_188_0, i_8_502_204_0,
    i_8_502_229_0, i_8_502_322_0, i_8_502_323_0, i_8_502_367_0,
    i_8_502_368_0, i_8_502_385_0, i_8_502_403_0, i_8_502_404_0,
    i_8_502_489_0, i_8_502_511_0, i_8_502_538_0, i_8_502_556_0,
    i_8_502_557_0, i_8_502_584_0, i_8_502_610_0, i_8_502_617_0,
    i_8_502_661_0, i_8_502_664_0, i_8_502_682_0, i_8_502_703_0,
    i_8_502_710_0, i_8_502_763_0, i_8_502_827_0, i_8_502_899_0,
    i_8_502_997_0, i_8_502_1006_0, i_8_502_1075_0, i_8_502_1105_0,
    i_8_502_1106_0, i_8_502_1113_0, i_8_502_1169_0, i_8_502_1180_0,
    i_8_502_1181_0, i_8_502_1186_0, i_8_502_1205_0, i_8_502_1261_0,
    i_8_502_1289_0, i_8_502_1340_0, i_8_502_1439_0, i_8_502_1444_0,
    i_8_502_1465_0, i_8_502_1471_0, i_8_502_1474_0, i_8_502_1483_0,
    i_8_502_1484_0, i_8_502_1501_0, i_8_502_1516_0, i_8_502_1520_0,
    i_8_502_1528_0, i_8_502_1529_0, i_8_502_1553_0, i_8_502_1561_0,
    i_8_502_1626_0, i_8_502_1632_0, i_8_502_1636_0, i_8_502_1646_0,
    i_8_502_1651_0, i_8_502_1663_0, i_8_502_1690_0, i_8_502_1699_0,
    i_8_502_1733_0, i_8_502_1753_0, i_8_502_1771_0, i_8_502_1787_0,
    i_8_502_1798_0, i_8_502_1800_0, i_8_502_1816_0, i_8_502_1898_0,
    i_8_502_1916_0, i_8_502_1942_0, i_8_502_1952_0, i_8_502_1958_0,
    i_8_502_1960_0, i_8_502_1966_0, i_8_502_1967_0, i_8_502_1969_0,
    i_8_502_1970_0, i_8_502_1988_0, i_8_502_2020_0, i_8_502_2060_0,
    i_8_502_2077_0, i_8_502_2104_0, i_8_502_2148_0, i_8_502_2172_0,
    i_8_502_2186_0, i_8_502_2194_0, i_8_502_2215_0, i_8_502_2218_0,
    i_8_502_2230_0, i_8_502_2239_0, i_8_502_2266_0,
    o_8_502_0_0  );
  input  i_8_502_15_0, i_8_502_17_0, i_8_502_44_0, i_8_502_60_0,
    i_8_502_67_0, i_8_502_71_0, i_8_502_142_0, i_8_502_188_0,
    i_8_502_204_0, i_8_502_229_0, i_8_502_322_0, i_8_502_323_0,
    i_8_502_367_0, i_8_502_368_0, i_8_502_385_0, i_8_502_403_0,
    i_8_502_404_0, i_8_502_489_0, i_8_502_511_0, i_8_502_538_0,
    i_8_502_556_0, i_8_502_557_0, i_8_502_584_0, i_8_502_610_0,
    i_8_502_617_0, i_8_502_661_0, i_8_502_664_0, i_8_502_682_0,
    i_8_502_703_0, i_8_502_710_0, i_8_502_763_0, i_8_502_827_0,
    i_8_502_899_0, i_8_502_997_0, i_8_502_1006_0, i_8_502_1075_0,
    i_8_502_1105_0, i_8_502_1106_0, i_8_502_1113_0, i_8_502_1169_0,
    i_8_502_1180_0, i_8_502_1181_0, i_8_502_1186_0, i_8_502_1205_0,
    i_8_502_1261_0, i_8_502_1289_0, i_8_502_1340_0, i_8_502_1439_0,
    i_8_502_1444_0, i_8_502_1465_0, i_8_502_1471_0, i_8_502_1474_0,
    i_8_502_1483_0, i_8_502_1484_0, i_8_502_1501_0, i_8_502_1516_0,
    i_8_502_1520_0, i_8_502_1528_0, i_8_502_1529_0, i_8_502_1553_0,
    i_8_502_1561_0, i_8_502_1626_0, i_8_502_1632_0, i_8_502_1636_0,
    i_8_502_1646_0, i_8_502_1651_0, i_8_502_1663_0, i_8_502_1690_0,
    i_8_502_1699_0, i_8_502_1733_0, i_8_502_1753_0, i_8_502_1771_0,
    i_8_502_1787_0, i_8_502_1798_0, i_8_502_1800_0, i_8_502_1816_0,
    i_8_502_1898_0, i_8_502_1916_0, i_8_502_1942_0, i_8_502_1952_0,
    i_8_502_1958_0, i_8_502_1960_0, i_8_502_1966_0, i_8_502_1967_0,
    i_8_502_1969_0, i_8_502_1970_0, i_8_502_1988_0, i_8_502_2020_0,
    i_8_502_2060_0, i_8_502_2077_0, i_8_502_2104_0, i_8_502_2148_0,
    i_8_502_2172_0, i_8_502_2186_0, i_8_502_2194_0, i_8_502_2215_0,
    i_8_502_2218_0, i_8_502_2230_0, i_8_502_2239_0, i_8_502_2266_0;
  output o_8_502_0_0;
  assign o_8_502_0_0 = ~((~i_8_502_584_0 & ((~i_8_502_44_0 & ((~i_8_502_682_0 & ~i_8_502_1444_0 & ~i_8_502_1465_0 & ~i_8_502_1484_0 & ~i_8_502_1916_0) | (~i_8_502_538_0 & ~i_8_502_899_0 & ~i_8_502_1340_0 & ~i_8_502_2104_0))) | (~i_8_502_2266_0 & ((~i_8_502_323_0 & i_8_502_617_0 & ~i_8_502_703_0 & ~i_8_502_1075_0 & ~i_8_502_1105_0 & ~i_8_502_1181_0 & ~i_8_502_1690_0 & ~i_8_502_1798_0 & ~i_8_502_2077_0 & ~i_8_502_2148_0) | (~i_8_502_322_0 & ~i_8_502_1113_0 & ~i_8_502_1186_0 & ~i_8_502_1205_0 & ~i_8_502_1465_0 & ~i_8_502_1501_0 & ~i_8_502_1528_0 & ~i_8_502_1561_0 & ~i_8_502_2239_0))))) | (~i_8_502_2194_0 & ((~i_8_502_71_0 & ((~i_8_502_827_0 & ~i_8_502_1186_0 & ~i_8_502_1484_0 & ~i_8_502_1632_0) | (~i_8_502_538_0 & ~i_8_502_1205_0 & ~i_8_502_1916_0 & ~i_8_502_1942_0 & ~i_8_502_1958_0))) | (~i_8_502_403_0 & ~i_8_502_1444_0 & ((~i_8_502_1205_0 & ~i_8_502_2020_0 & i_8_502_2172_0) | (~i_8_502_15_0 & ~i_8_502_1181_0 & ~i_8_502_1465_0 & ~i_8_502_1516_0 & ~i_8_502_1529_0 & ~i_8_502_1690_0 & ~i_8_502_1942_0 & ~i_8_502_2266_0))) | (~i_8_502_1960_0 & ((~i_8_502_404_0 & ~i_8_502_617_0 & ~i_8_502_1520_0 & i_8_502_1753_0 & ~i_8_502_1787_0 & ~i_8_502_1958_0) | (~i_8_502_229_0 & ~i_8_502_827_0 & ~i_8_502_899_0 & ~i_8_502_1465_0 & ~i_8_502_1553_0 & ~i_8_502_1898_0 & ~i_8_502_1916_0 & ~i_8_502_1967_0))))) | (i_8_502_1006_0 & ((~i_8_502_710_0 & ~i_8_502_1169_0 & ~i_8_502_1186_0 & ~i_8_502_1663_0 & i_8_502_1733_0) | (~i_8_502_367_0 & i_8_502_617_0 & ~i_8_502_682_0 & ~i_8_502_1181_0 & ~i_8_502_1561_0 & i_8_502_1753_0 & ~i_8_502_1960_0))) | (~i_8_502_1636_0 & ((~i_8_502_511_0 & ~i_8_502_664_0 & ~i_8_502_1105_0 & ~i_8_502_1113_0 & ~i_8_502_1516_0 & ~i_8_502_1520_0 & ~i_8_502_1690_0) | (i_8_502_368_0 & i_8_502_385_0 & ~i_8_502_1106_0 & ~i_8_502_1169_0 & ~i_8_502_1529_0 & ~i_8_502_1958_0))) | (~i_8_502_1529_0 & ((~i_8_502_142_0 & i_8_502_367_0 & i_8_502_1636_0 & ~i_8_502_1690_0) | (i_8_502_763_0 & ~i_8_502_1733_0))) | (~i_8_502_556_0 & ~i_8_502_557_0 & ~i_8_502_661_0 & ~i_8_502_827_0 & ~i_8_502_1483_0) | (~i_8_502_71_0 & ~i_8_502_899_0 & ~i_8_502_1465_0 & ~i_8_502_1753_0 & ~i_8_502_1787_0 & ~i_8_502_2020_0));
endmodule



// Benchmark "kernel_8_503" written by ABC on Sun Jul 19 10:11:53 2020

module kernel_8_503 ( 
    i_8_503_54_0, i_8_503_74_0, i_8_503_86_0, i_8_503_136_0, i_8_503_138_0,
    i_8_503_158_0, i_8_503_162_0, i_8_503_176_0, i_8_503_212_0,
    i_8_503_236_0, i_8_503_242_0, i_8_503_253_0, i_8_503_274_0,
    i_8_503_304_0, i_8_503_311_0, i_8_503_334_0, i_8_503_361_0,
    i_8_503_392_0, i_8_503_401_0, i_8_503_455_0, i_8_503_472_0,
    i_8_503_475_0, i_8_503_478_0, i_8_503_479_0, i_8_503_491_0,
    i_8_503_496_0, i_8_503_505_0, i_8_503_524_0, i_8_503_607_0,
    i_8_503_608_0, i_8_503_659_0, i_8_503_660_0, i_8_503_682_0,
    i_8_503_684_0, i_8_503_689_0, i_8_503_716_0, i_8_503_761_0,
    i_8_503_776_0, i_8_503_797_0, i_8_503_860_0, i_8_503_886_0,
    i_8_503_922_0, i_8_503_932_0, i_8_503_949_0, i_8_503_1058_0,
    i_8_503_1099_0, i_8_503_1112_0, i_8_503_1154_0, i_8_503_1175_0,
    i_8_503_1189_0, i_8_503_1190_0, i_8_503_1224_0, i_8_503_1233_0,
    i_8_503_1240_0, i_8_503_1256_0, i_8_503_1282_0, i_8_503_1283_0,
    i_8_503_1288_0, i_8_503_1308_0, i_8_503_1325_0, i_8_503_1326_0,
    i_8_503_1337_0, i_8_503_1409_0, i_8_503_1418_0, i_8_503_1439_0,
    i_8_503_1456_0, i_8_503_1468_0, i_8_503_1472_0, i_8_503_1480_0,
    i_8_503_1487_0, i_8_503_1605_0, i_8_503_1607_0, i_8_503_1631_0,
    i_8_503_1639_0, i_8_503_1650_0, i_8_503_1677_0, i_8_503_1696_0,
    i_8_503_1700_0, i_8_503_1713_0, i_8_503_1721_0, i_8_503_1760_0,
    i_8_503_1785_0, i_8_503_1820_0, i_8_503_1835_0, i_8_503_1936_0,
    i_8_503_1981_0, i_8_503_2003_0, i_8_503_2035_0, i_8_503_2039_0,
    i_8_503_2053_0, i_8_503_2075_0, i_8_503_2156_0, i_8_503_2159_0,
    i_8_503_2201_0, i_8_503_2210_0, i_8_503_2223_0, i_8_503_2231_0,
    i_8_503_2246_0, i_8_503_2261_0, i_8_503_2263_0,
    o_8_503_0_0  );
  input  i_8_503_54_0, i_8_503_74_0, i_8_503_86_0, i_8_503_136_0,
    i_8_503_138_0, i_8_503_158_0, i_8_503_162_0, i_8_503_176_0,
    i_8_503_212_0, i_8_503_236_0, i_8_503_242_0, i_8_503_253_0,
    i_8_503_274_0, i_8_503_304_0, i_8_503_311_0, i_8_503_334_0,
    i_8_503_361_0, i_8_503_392_0, i_8_503_401_0, i_8_503_455_0,
    i_8_503_472_0, i_8_503_475_0, i_8_503_478_0, i_8_503_479_0,
    i_8_503_491_0, i_8_503_496_0, i_8_503_505_0, i_8_503_524_0,
    i_8_503_607_0, i_8_503_608_0, i_8_503_659_0, i_8_503_660_0,
    i_8_503_682_0, i_8_503_684_0, i_8_503_689_0, i_8_503_716_0,
    i_8_503_761_0, i_8_503_776_0, i_8_503_797_0, i_8_503_860_0,
    i_8_503_886_0, i_8_503_922_0, i_8_503_932_0, i_8_503_949_0,
    i_8_503_1058_0, i_8_503_1099_0, i_8_503_1112_0, i_8_503_1154_0,
    i_8_503_1175_0, i_8_503_1189_0, i_8_503_1190_0, i_8_503_1224_0,
    i_8_503_1233_0, i_8_503_1240_0, i_8_503_1256_0, i_8_503_1282_0,
    i_8_503_1283_0, i_8_503_1288_0, i_8_503_1308_0, i_8_503_1325_0,
    i_8_503_1326_0, i_8_503_1337_0, i_8_503_1409_0, i_8_503_1418_0,
    i_8_503_1439_0, i_8_503_1456_0, i_8_503_1468_0, i_8_503_1472_0,
    i_8_503_1480_0, i_8_503_1487_0, i_8_503_1605_0, i_8_503_1607_0,
    i_8_503_1631_0, i_8_503_1639_0, i_8_503_1650_0, i_8_503_1677_0,
    i_8_503_1696_0, i_8_503_1700_0, i_8_503_1713_0, i_8_503_1721_0,
    i_8_503_1760_0, i_8_503_1785_0, i_8_503_1820_0, i_8_503_1835_0,
    i_8_503_1936_0, i_8_503_1981_0, i_8_503_2003_0, i_8_503_2035_0,
    i_8_503_2039_0, i_8_503_2053_0, i_8_503_2075_0, i_8_503_2156_0,
    i_8_503_2159_0, i_8_503_2201_0, i_8_503_2210_0, i_8_503_2223_0,
    i_8_503_2231_0, i_8_503_2246_0, i_8_503_2261_0, i_8_503_2263_0;
  output o_8_503_0_0;
  assign o_8_503_0_0 = 0;
endmodule



// Benchmark "kernel_8_504" written by ABC on Sun Jul 19 10:11:54 2020

module kernel_8_504 ( 
    i_8_504_51_0, i_8_504_73_0, i_8_504_111_0, i_8_504_114_0,
    i_8_504_228_0, i_8_504_229_0, i_8_504_286_0, i_8_504_297_0,
    i_8_504_303_0, i_8_504_384_0, i_8_504_399_0, i_8_504_403_0,
    i_8_504_420_0, i_8_504_550_0, i_8_504_585_0, i_8_504_593_0,
    i_8_504_600_0, i_8_504_601_0, i_8_504_610_0, i_8_504_657_0,
    i_8_504_664_0, i_8_504_667_0, i_8_504_668_0, i_8_504_683_0,
    i_8_504_699_0, i_8_504_700_0, i_8_504_701_0, i_8_504_702_0,
    i_8_504_711_0, i_8_504_780_0, i_8_504_781_0, i_8_504_790_0,
    i_8_504_816_0, i_8_504_822_0, i_8_504_823_0, i_8_504_825_0,
    i_8_504_835_0, i_8_504_843_0, i_8_504_844_0, i_8_504_845_0,
    i_8_504_856_0, i_8_504_861_0, i_8_504_870_0, i_8_504_880_0,
    i_8_504_889_0, i_8_504_892_0, i_8_504_928_0, i_8_504_931_0,
    i_8_504_939_0, i_8_504_940_0, i_8_504_1027_0, i_8_504_1041_0,
    i_8_504_1043_0, i_8_504_1107_0, i_8_504_1141_0, i_8_504_1146_0,
    i_8_504_1149_0, i_8_504_1166_0, i_8_504_1218_0, i_8_504_1242_0,
    i_8_504_1248_0, i_8_504_1284_0, i_8_504_1285_0, i_8_504_1305_0,
    i_8_504_1326_0, i_8_504_1335_0, i_8_504_1336_0, i_8_504_1353_0,
    i_8_504_1354_0, i_8_504_1356_0, i_8_504_1401_0, i_8_504_1425_0,
    i_8_504_1438_0, i_8_504_1473_0, i_8_504_1482_0, i_8_504_1510_0,
    i_8_504_1515_0, i_8_504_1546_0, i_8_504_1556_0, i_8_504_1606_0,
    i_8_504_1630_0, i_8_504_1633_0, i_8_504_1654_0, i_8_504_1714_0,
    i_8_504_1761_0, i_8_504_1776_0, i_8_504_1801_0, i_8_504_1839_0,
    i_8_504_1971_0, i_8_504_1981_0, i_8_504_1988_0, i_8_504_1997_0,
    i_8_504_2058_0, i_8_504_2074_0, i_8_504_2187_0, i_8_504_2214_0,
    i_8_504_2227_0, i_8_504_2248_0, i_8_504_2277_0, i_8_504_2299_0,
    o_8_504_0_0  );
  input  i_8_504_51_0, i_8_504_73_0, i_8_504_111_0, i_8_504_114_0,
    i_8_504_228_0, i_8_504_229_0, i_8_504_286_0, i_8_504_297_0,
    i_8_504_303_0, i_8_504_384_0, i_8_504_399_0, i_8_504_403_0,
    i_8_504_420_0, i_8_504_550_0, i_8_504_585_0, i_8_504_593_0,
    i_8_504_600_0, i_8_504_601_0, i_8_504_610_0, i_8_504_657_0,
    i_8_504_664_0, i_8_504_667_0, i_8_504_668_0, i_8_504_683_0,
    i_8_504_699_0, i_8_504_700_0, i_8_504_701_0, i_8_504_702_0,
    i_8_504_711_0, i_8_504_780_0, i_8_504_781_0, i_8_504_790_0,
    i_8_504_816_0, i_8_504_822_0, i_8_504_823_0, i_8_504_825_0,
    i_8_504_835_0, i_8_504_843_0, i_8_504_844_0, i_8_504_845_0,
    i_8_504_856_0, i_8_504_861_0, i_8_504_870_0, i_8_504_880_0,
    i_8_504_889_0, i_8_504_892_0, i_8_504_928_0, i_8_504_931_0,
    i_8_504_939_0, i_8_504_940_0, i_8_504_1027_0, i_8_504_1041_0,
    i_8_504_1043_0, i_8_504_1107_0, i_8_504_1141_0, i_8_504_1146_0,
    i_8_504_1149_0, i_8_504_1166_0, i_8_504_1218_0, i_8_504_1242_0,
    i_8_504_1248_0, i_8_504_1284_0, i_8_504_1285_0, i_8_504_1305_0,
    i_8_504_1326_0, i_8_504_1335_0, i_8_504_1336_0, i_8_504_1353_0,
    i_8_504_1354_0, i_8_504_1356_0, i_8_504_1401_0, i_8_504_1425_0,
    i_8_504_1438_0, i_8_504_1473_0, i_8_504_1482_0, i_8_504_1510_0,
    i_8_504_1515_0, i_8_504_1546_0, i_8_504_1556_0, i_8_504_1606_0,
    i_8_504_1630_0, i_8_504_1633_0, i_8_504_1654_0, i_8_504_1714_0,
    i_8_504_1761_0, i_8_504_1776_0, i_8_504_1801_0, i_8_504_1839_0,
    i_8_504_1971_0, i_8_504_1981_0, i_8_504_1988_0, i_8_504_1997_0,
    i_8_504_2058_0, i_8_504_2074_0, i_8_504_2187_0, i_8_504_2214_0,
    i_8_504_2227_0, i_8_504_2248_0, i_8_504_2277_0, i_8_504_2299_0;
  output o_8_504_0_0;
  assign o_8_504_0_0 = 0;
endmodule



// Benchmark "kernel_8_505" written by ABC on Sun Jul 19 10:11:55 2020

module kernel_8_505 ( 
    i_8_505_49_0, i_8_505_67_0, i_8_505_95_0, i_8_505_112_0, i_8_505_135_0,
    i_8_505_139_0, i_8_505_162_0, i_8_505_163_0, i_8_505_180_0,
    i_8_505_189_0, i_8_505_217_0, i_8_505_220_0, i_8_505_234_0,
    i_8_505_235_0, i_8_505_261_0, i_8_505_298_0, i_8_505_333_0,
    i_8_505_344_0, i_8_505_362_0, i_8_505_368_0, i_8_505_414_0,
    i_8_505_415_0, i_8_505_436_0, i_8_505_437_0, i_8_505_483_0,
    i_8_505_489_0, i_8_505_588_0, i_8_505_608_0, i_8_505_612_0,
    i_8_505_621_0, i_8_505_624_0, i_8_505_631_0, i_8_505_684_0,
    i_8_505_697_0, i_8_505_704_0, i_8_505_748_0, i_8_505_777_0,
    i_8_505_779_0, i_8_505_802_0, i_8_505_822_0, i_8_505_823_0,
    i_8_505_832_0, i_8_505_841_0, i_8_505_873_0, i_8_505_883_0,
    i_8_505_921_0, i_8_505_930_0, i_8_505_937_0, i_8_505_967_0,
    i_8_505_971_0, i_8_505_991_0, i_8_505_1011_0, i_8_505_1012_0,
    i_8_505_1038_0, i_8_505_1053_0, i_8_505_1056_0, i_8_505_1071_0,
    i_8_505_1104_0, i_8_505_1114_0, i_8_505_1170_0, i_8_505_1235_0,
    i_8_505_1278_0, i_8_505_1279_0, i_8_505_1284_0, i_8_505_1287_0,
    i_8_505_1288_0, i_8_505_1395_0, i_8_505_1404_0, i_8_505_1407_0,
    i_8_505_1434_0, i_8_505_1476_0, i_8_505_1488_0, i_8_505_1535_0,
    i_8_505_1539_0, i_8_505_1588_0, i_8_505_1740_0, i_8_505_1748_0,
    i_8_505_1756_0, i_8_505_1800_0, i_8_505_1804_0, i_8_505_1827_0,
    i_8_505_1828_0, i_8_505_1830_0, i_8_505_1864_0, i_8_505_1986_0,
    i_8_505_1992_0, i_8_505_2007_0, i_8_505_2019_0, i_8_505_2035_0,
    i_8_505_2037_0, i_8_505_2043_0, i_8_505_2044_0, i_8_505_2053_0,
    i_8_505_2070_0, i_8_505_2095_0, i_8_505_2133_0, i_8_505_2187_0,
    i_8_505_2206_0, i_8_505_2215_0, i_8_505_2268_0,
    o_8_505_0_0  );
  input  i_8_505_49_0, i_8_505_67_0, i_8_505_95_0, i_8_505_112_0,
    i_8_505_135_0, i_8_505_139_0, i_8_505_162_0, i_8_505_163_0,
    i_8_505_180_0, i_8_505_189_0, i_8_505_217_0, i_8_505_220_0,
    i_8_505_234_0, i_8_505_235_0, i_8_505_261_0, i_8_505_298_0,
    i_8_505_333_0, i_8_505_344_0, i_8_505_362_0, i_8_505_368_0,
    i_8_505_414_0, i_8_505_415_0, i_8_505_436_0, i_8_505_437_0,
    i_8_505_483_0, i_8_505_489_0, i_8_505_588_0, i_8_505_608_0,
    i_8_505_612_0, i_8_505_621_0, i_8_505_624_0, i_8_505_631_0,
    i_8_505_684_0, i_8_505_697_0, i_8_505_704_0, i_8_505_748_0,
    i_8_505_777_0, i_8_505_779_0, i_8_505_802_0, i_8_505_822_0,
    i_8_505_823_0, i_8_505_832_0, i_8_505_841_0, i_8_505_873_0,
    i_8_505_883_0, i_8_505_921_0, i_8_505_930_0, i_8_505_937_0,
    i_8_505_967_0, i_8_505_971_0, i_8_505_991_0, i_8_505_1011_0,
    i_8_505_1012_0, i_8_505_1038_0, i_8_505_1053_0, i_8_505_1056_0,
    i_8_505_1071_0, i_8_505_1104_0, i_8_505_1114_0, i_8_505_1170_0,
    i_8_505_1235_0, i_8_505_1278_0, i_8_505_1279_0, i_8_505_1284_0,
    i_8_505_1287_0, i_8_505_1288_0, i_8_505_1395_0, i_8_505_1404_0,
    i_8_505_1407_0, i_8_505_1434_0, i_8_505_1476_0, i_8_505_1488_0,
    i_8_505_1535_0, i_8_505_1539_0, i_8_505_1588_0, i_8_505_1740_0,
    i_8_505_1748_0, i_8_505_1756_0, i_8_505_1800_0, i_8_505_1804_0,
    i_8_505_1827_0, i_8_505_1828_0, i_8_505_1830_0, i_8_505_1864_0,
    i_8_505_1986_0, i_8_505_1992_0, i_8_505_2007_0, i_8_505_2019_0,
    i_8_505_2035_0, i_8_505_2037_0, i_8_505_2043_0, i_8_505_2044_0,
    i_8_505_2053_0, i_8_505_2070_0, i_8_505_2095_0, i_8_505_2133_0,
    i_8_505_2187_0, i_8_505_2206_0, i_8_505_2215_0, i_8_505_2268_0;
  output o_8_505_0_0;
  assign o_8_505_0_0 = ~((~i_8_505_112_0 & ((i_8_505_414_0 & ~i_8_505_1278_0 & ~i_8_505_1407_0) | (~i_8_505_930_0 & ~i_8_505_1053_0 & ~i_8_505_1279_0 & ~i_8_505_1992_0 & ~i_8_505_2037_0))) | (~i_8_505_135_0 & ((i_8_505_112_0 & ~i_8_505_608_0 & ~i_8_505_1071_0 & i_8_505_1114_0 & ~i_8_505_1827_0) | (~i_8_505_163_0 & ~i_8_505_588_0 & ~i_8_505_1053_0 & ~i_8_505_1284_0 & ~i_8_505_1588_0 & ~i_8_505_1830_0 & ~i_8_505_2053_0))) | (~i_8_505_49_0 & ((~i_8_505_139_0 & ((~i_8_505_612_0 & ~i_8_505_991_0 & ~i_8_505_1288_0 & ~i_8_505_1404_0 & i_8_505_1804_0) | (~i_8_505_163_0 & ~i_8_505_298_0 & ~i_8_505_841_0 & ~i_8_505_873_0 & ~i_8_505_921_0 & ~i_8_505_937_0 & ~i_8_505_971_0 & ~i_8_505_1038_0 & ~i_8_505_1827_0 & ~i_8_505_2043_0))) | (~i_8_505_162_0 & ~i_8_505_235_0 & ~i_8_505_1071_0 & ~i_8_505_1170_0 & ~i_8_505_1284_0 & ~i_8_505_1287_0 & ~i_8_505_2035_0))) | (~i_8_505_930_0 & ((~i_8_505_162_0 & ((~i_8_505_163_0 & ~i_8_505_234_0 & ~i_8_505_1287_0 & ~i_8_505_2019_0 & ~i_8_505_2035_0 & ~i_8_505_2037_0) | (i_8_505_217_0 & ~i_8_505_991_0 & ~i_8_505_1170_0 & ~i_8_505_1288_0 & ~i_8_505_1830_0 & ~i_8_505_2133_0))) | (~i_8_505_802_0 & ((~i_8_505_631_0 & ~i_8_505_1053_0 & ~i_8_505_1287_0 & ~i_8_505_1756_0 & ~i_8_505_2037_0) | (~i_8_505_180_0 & ~i_8_505_841_0 & ~i_8_505_1104_0 & ~i_8_505_1170_0 & ~i_8_505_1279_0 & ~i_8_505_1828_0 & ~i_8_505_2019_0 & ~i_8_505_2043_0))) | (~i_8_505_235_0 & ~i_8_505_483_0 & ~i_8_505_612_0 & ~i_8_505_1278_0 & ~i_8_505_1279_0 & ~i_8_505_2019_0))) | (~i_8_505_684_0 & ((~i_8_505_235_0 & ~i_8_505_802_0 & ((i_8_505_414_0 & ~i_8_505_1830_0) | (~i_8_505_333_0 & ~i_8_505_1104_0 & ~i_8_505_1407_0 & ~i_8_505_1804_0 & ~i_8_505_2187_0))) | (i_8_505_217_0 & ~i_8_505_1056_0 & ~i_8_505_1114_0 & ~i_8_505_1588_0 & ~i_8_505_1827_0) | (i_8_505_612_0 & i_8_505_832_0 & ~i_8_505_1038_0 & ~i_8_505_1287_0 & ~i_8_505_2019_0))) | (i_8_505_823_0 & (~i_8_505_1056_0 | i_8_505_2206_0)) | (~i_8_505_1740_0 & ((i_8_505_135_0 & i_8_505_489_0 & i_8_505_1284_0 & ~i_8_505_1287_0 & ~i_8_505_1288_0 & ~i_8_505_1404_0 & ~i_8_505_1800_0 & ~i_8_505_1804_0) | (i_8_505_624_0 & ~i_8_505_631_0 & ~i_8_505_937_0 & ~i_8_505_1864_0 & ~i_8_505_2070_0))) | (~i_8_505_483_0 & i_8_505_621_0 & ~i_8_505_802_0 & i_8_505_1800_0) | (i_8_505_220_0 & ~i_8_505_624_0 & ~i_8_505_991_0 & ~i_8_505_1284_0 & ~i_8_505_1828_0) | (~i_8_505_234_0 & i_8_505_362_0 & ~i_8_505_1827_0 & ~i_8_505_2037_0 & ~i_8_505_2206_0) | (~i_8_505_921_0 & ~i_8_505_1038_0 & ~i_8_505_1056_0 & ~i_8_505_1170_0 & ~i_8_505_1434_0 & ~i_8_505_1588_0 & ~i_8_505_1756_0 & ~i_8_505_1830_0 & ~i_8_505_2268_0));
endmodule



// Benchmark "kernel_8_506" written by ABC on Sun Jul 19 10:11:56 2020

module kernel_8_506 ( 
    i_8_506_28_0, i_8_506_38_0, i_8_506_64_0, i_8_506_65_0, i_8_506_139_0,
    i_8_506_165_0, i_8_506_173_0, i_8_506_212_0, i_8_506_227_0,
    i_8_506_260_0, i_8_506_308_0, i_8_506_325_0, i_8_506_332_0,
    i_8_506_335_0, i_8_506_338_0, i_8_506_344_0, i_8_506_365_0,
    i_8_506_368_0, i_8_506_404_0, i_8_506_421_0, i_8_506_428_0,
    i_8_506_455_0, i_8_506_490_0, i_8_506_493_0, i_8_506_494_0,
    i_8_506_553_0, i_8_506_583_0, i_8_506_584_0, i_8_506_606_0,
    i_8_506_689_0, i_8_506_707_0, i_8_506_719_0, i_8_506_730_0,
    i_8_506_734_0, i_8_506_797_0, i_8_506_800_0, i_8_506_815_0,
    i_8_506_818_0, i_8_506_853_0, i_8_506_854_0, i_8_506_876_0,
    i_8_506_884_0, i_8_506_923_0, i_8_506_931_0, i_8_506_935_0,
    i_8_506_956_0, i_8_506_971_0, i_8_506_1052_0, i_8_506_1060_0,
    i_8_506_1079_0, i_8_506_1094_0, i_8_506_1107_0, i_8_506_1114_0,
    i_8_506_1115_0, i_8_506_1172_0, i_8_506_1175_0, i_8_506_1238_0,
    i_8_506_1264_0, i_8_506_1265_0, i_8_506_1282_0, i_8_506_1290_0,
    i_8_506_1292_0, i_8_506_1308_0, i_8_506_1322_0, i_8_506_1330_0,
    i_8_506_1409_0, i_8_506_1411_0, i_8_506_1488_0, i_8_506_1520_0,
    i_8_506_1535_0, i_8_506_1586_0, i_8_506_1598_0, i_8_506_1655_0,
    i_8_506_1672_0, i_8_506_1703_0, i_8_506_1706_0, i_8_506_1709_0,
    i_8_506_1760_0, i_8_506_1821_0, i_8_506_1825_0, i_8_506_1922_0,
    i_8_506_1937_0, i_8_506_1951_0, i_8_506_1995_0, i_8_506_1996_0,
    i_8_506_2018_0, i_8_506_2021_0, i_8_506_2075_0, i_8_506_2111_0,
    i_8_506_2120_0, i_8_506_2170_0, i_8_506_2174_0, i_8_506_2180_0,
    i_8_506_2201_0, i_8_506_2209_0, i_8_506_2210_0, i_8_506_2227_0,
    i_8_506_2233_0, i_8_506_2239_0, i_8_506_2276_0,
    o_8_506_0_0  );
  input  i_8_506_28_0, i_8_506_38_0, i_8_506_64_0, i_8_506_65_0,
    i_8_506_139_0, i_8_506_165_0, i_8_506_173_0, i_8_506_212_0,
    i_8_506_227_0, i_8_506_260_0, i_8_506_308_0, i_8_506_325_0,
    i_8_506_332_0, i_8_506_335_0, i_8_506_338_0, i_8_506_344_0,
    i_8_506_365_0, i_8_506_368_0, i_8_506_404_0, i_8_506_421_0,
    i_8_506_428_0, i_8_506_455_0, i_8_506_490_0, i_8_506_493_0,
    i_8_506_494_0, i_8_506_553_0, i_8_506_583_0, i_8_506_584_0,
    i_8_506_606_0, i_8_506_689_0, i_8_506_707_0, i_8_506_719_0,
    i_8_506_730_0, i_8_506_734_0, i_8_506_797_0, i_8_506_800_0,
    i_8_506_815_0, i_8_506_818_0, i_8_506_853_0, i_8_506_854_0,
    i_8_506_876_0, i_8_506_884_0, i_8_506_923_0, i_8_506_931_0,
    i_8_506_935_0, i_8_506_956_0, i_8_506_971_0, i_8_506_1052_0,
    i_8_506_1060_0, i_8_506_1079_0, i_8_506_1094_0, i_8_506_1107_0,
    i_8_506_1114_0, i_8_506_1115_0, i_8_506_1172_0, i_8_506_1175_0,
    i_8_506_1238_0, i_8_506_1264_0, i_8_506_1265_0, i_8_506_1282_0,
    i_8_506_1290_0, i_8_506_1292_0, i_8_506_1308_0, i_8_506_1322_0,
    i_8_506_1330_0, i_8_506_1409_0, i_8_506_1411_0, i_8_506_1488_0,
    i_8_506_1520_0, i_8_506_1535_0, i_8_506_1586_0, i_8_506_1598_0,
    i_8_506_1655_0, i_8_506_1672_0, i_8_506_1703_0, i_8_506_1706_0,
    i_8_506_1709_0, i_8_506_1760_0, i_8_506_1821_0, i_8_506_1825_0,
    i_8_506_1922_0, i_8_506_1937_0, i_8_506_1951_0, i_8_506_1995_0,
    i_8_506_1996_0, i_8_506_2018_0, i_8_506_2021_0, i_8_506_2075_0,
    i_8_506_2111_0, i_8_506_2120_0, i_8_506_2170_0, i_8_506_2174_0,
    i_8_506_2180_0, i_8_506_2201_0, i_8_506_2209_0, i_8_506_2210_0,
    i_8_506_2227_0, i_8_506_2233_0, i_8_506_2239_0, i_8_506_2276_0;
  output o_8_506_0_0;
  assign o_8_506_0_0 = ~((~i_8_506_28_0 & ((~i_8_506_38_0 & ~i_8_506_344_0 & ~i_8_506_800_0 & ~i_8_506_1175_0 & ~i_8_506_1238_0 & ~i_8_506_1322_0 & ~i_8_506_1520_0 & ~i_8_506_1937_0) | (~i_8_506_212_0 & ~i_8_506_1094_0 & ~i_8_506_1172_0 & ~i_8_506_1292_0 & ~i_8_506_1488_0 & ~i_8_506_1709_0 & ~i_8_506_2018_0 & ~i_8_506_2210_0))) | (~i_8_506_65_0 & ((~i_8_506_173_0 & ~i_8_506_212_0 & ~i_8_506_335_0 & ~i_8_506_494_0 & ~i_8_506_1094_0 & ~i_8_506_1409_0) | (~i_8_506_404_0 & ~i_8_506_583_0 & i_8_506_1115_0 & ~i_8_506_2021_0 & i_8_506_2276_0))) | (~i_8_506_212_0 & ((~i_8_506_38_0 & ~i_8_506_260_0 & ~i_8_506_404_0 & i_8_506_428_0 & ~i_8_506_818_0 & ~i_8_506_1060_0 & ~i_8_506_1292_0 & ~i_8_506_2180_0 & ~i_8_506_2201_0) | (~i_8_506_2018_0 & ~i_8_506_2210_0 & ~i_8_506_689_0 & i_8_506_730_0))) | (~i_8_506_38_0 & ((~i_8_506_800_0 & i_8_506_1052_0 & ~i_8_506_1175_0 & ~i_8_506_2021_0) | (~i_8_506_173_0 & ~i_8_506_260_0 & ~i_8_506_428_0 & ~i_8_506_584_0 & ~i_8_506_923_0 & ~i_8_506_1703_0 & ~i_8_506_2209_0))) | (~i_8_506_797_0 & ((~i_8_506_455_0 & ((~i_8_506_584_0 & i_8_506_1996_0) | (~i_8_506_493_0 & ~i_8_506_956_0 & ~i_8_506_1322_0 & ~i_8_506_2180_0 & ~i_8_506_2233_0))) | (~i_8_506_1520_0 & ((~i_8_506_344_0 & ~i_8_506_815_0 & i_8_506_1238_0 & ~i_8_506_1292_0 & ~i_8_506_2174_0) | (~i_8_506_490_0 & ~i_8_506_935_0 & ~i_8_506_1172_0 & ~i_8_506_1322_0 & ~i_8_506_2180_0))) | (i_8_506_1292_0 & i_8_506_1996_0))) | (~i_8_506_689_0 & ((~i_8_506_730_0 & ~i_8_506_800_0 & ~i_8_506_971_0 & ~i_8_506_1238_0 & i_8_506_1282_0 & ~i_8_506_1409_0 & ~i_8_506_1937_0) | (~i_8_506_173_0 & ~i_8_506_428_0 & ~i_8_506_1703_0 & ~i_8_506_2018_0 & ~i_8_506_2111_0 & ~i_8_506_2201_0))) | (~i_8_506_2018_0 & ((~i_8_506_173_0 & ~i_8_506_2174_0 & ((~i_8_506_260_0 & ~i_8_506_730_0 & ~i_8_506_1175_0 & i_8_506_1922_0 & ~i_8_506_1996_0 & ~i_8_506_2201_0 & ~i_8_506_2210_0) | (~i_8_506_493_0 & ~i_8_506_923_0 & ~i_8_506_1172_0 & i_8_506_1282_0 & ~i_8_506_1411_0 & ~i_8_506_1535_0 & ~i_8_506_2276_0))) | (i_8_506_428_0 & ~i_8_506_935_0 & i_8_506_2120_0))) | (~i_8_506_956_0 & ((~i_8_506_338_0 & ~i_8_506_734_0 & ~i_8_506_1052_0 & ~i_8_506_1172_0 & ~i_8_506_1709_0 & ~i_8_506_2111_0) | (i_8_506_493_0 & ~i_8_506_1107_0 & ~i_8_506_1264_0 & ~i_8_506_1282_0 & ~i_8_506_1292_0 & ~i_8_506_1703_0 & ~i_8_506_2180_0))));
endmodule



// Benchmark "kernel_8_507" written by ABC on Sun Jul 19 10:11:57 2020

module kernel_8_507 ( 
    i_8_507_11_0, i_8_507_74_0, i_8_507_76_0, i_8_507_77_0, i_8_507_142_0,
    i_8_507_182_0, i_8_507_209_0, i_8_507_218_0, i_8_507_221_0,
    i_8_507_281_0, i_8_507_305_0, i_8_507_311_0, i_8_507_317_0,
    i_8_507_325_0, i_8_507_365_0, i_8_507_371_0, i_8_507_383_0,
    i_8_507_392_0, i_8_507_398_0, i_8_507_424_0, i_8_507_484_0,
    i_8_507_524_0, i_8_507_572_0, i_8_507_590_0, i_8_507_595_0,
    i_8_507_596_0, i_8_507_605_0, i_8_507_607_0, i_8_507_622_0,
    i_8_507_623_0, i_8_507_634_0, i_8_507_635_0, i_8_507_658_0,
    i_8_507_659_0, i_8_507_676_0, i_8_507_679_0, i_8_507_703_0,
    i_8_507_765_0, i_8_507_793_0, i_8_507_823_0, i_8_507_842_0,
    i_8_507_941_0, i_8_507_943_0, i_8_507_1102_0, i_8_507_1181_0,
    i_8_507_1198_0, i_8_507_1227_0, i_8_507_1235_0, i_8_507_1243_0,
    i_8_507_1244_0, i_8_507_1265_0, i_8_507_1267_0, i_8_507_1274_0,
    i_8_507_1282_0, i_8_507_1283_0, i_8_507_1337_0, i_8_507_1370_0,
    i_8_507_1396_0, i_8_507_1433_0, i_8_507_1451_0, i_8_507_1454_0,
    i_8_507_1478_0, i_8_507_1504_0, i_8_507_1507_0, i_8_507_1540_0,
    i_8_507_1544_0, i_8_507_1558_0, i_8_507_1565_0, i_8_507_1568_0,
    i_8_507_1570_0, i_8_507_1582_0, i_8_507_1631_0, i_8_507_1633_0,
    i_8_507_1649_0, i_8_507_1702_0, i_8_507_1733_0, i_8_507_1775_0,
    i_8_507_1777_0, i_8_507_1783_0, i_8_507_1786_0, i_8_507_1804_0,
    i_8_507_1817_0, i_8_507_1838_0, i_8_507_1841_0, i_8_507_1859_0,
    i_8_507_1886_0, i_8_507_1945_0, i_8_507_1946_0, i_8_507_1972_0,
    i_8_507_1973_0, i_8_507_2000_0, i_8_507_2044_0, i_8_507_2141_0,
    i_8_507_2155_0, i_8_507_2180_0, i_8_507_2206_0, i_8_507_2236_0,
    i_8_507_2245_0, i_8_507_2270_0, i_8_507_2285_0,
    o_8_507_0_0  );
  input  i_8_507_11_0, i_8_507_74_0, i_8_507_76_0, i_8_507_77_0,
    i_8_507_142_0, i_8_507_182_0, i_8_507_209_0, i_8_507_218_0,
    i_8_507_221_0, i_8_507_281_0, i_8_507_305_0, i_8_507_311_0,
    i_8_507_317_0, i_8_507_325_0, i_8_507_365_0, i_8_507_371_0,
    i_8_507_383_0, i_8_507_392_0, i_8_507_398_0, i_8_507_424_0,
    i_8_507_484_0, i_8_507_524_0, i_8_507_572_0, i_8_507_590_0,
    i_8_507_595_0, i_8_507_596_0, i_8_507_605_0, i_8_507_607_0,
    i_8_507_622_0, i_8_507_623_0, i_8_507_634_0, i_8_507_635_0,
    i_8_507_658_0, i_8_507_659_0, i_8_507_676_0, i_8_507_679_0,
    i_8_507_703_0, i_8_507_765_0, i_8_507_793_0, i_8_507_823_0,
    i_8_507_842_0, i_8_507_941_0, i_8_507_943_0, i_8_507_1102_0,
    i_8_507_1181_0, i_8_507_1198_0, i_8_507_1227_0, i_8_507_1235_0,
    i_8_507_1243_0, i_8_507_1244_0, i_8_507_1265_0, i_8_507_1267_0,
    i_8_507_1274_0, i_8_507_1282_0, i_8_507_1283_0, i_8_507_1337_0,
    i_8_507_1370_0, i_8_507_1396_0, i_8_507_1433_0, i_8_507_1451_0,
    i_8_507_1454_0, i_8_507_1478_0, i_8_507_1504_0, i_8_507_1507_0,
    i_8_507_1540_0, i_8_507_1544_0, i_8_507_1558_0, i_8_507_1565_0,
    i_8_507_1568_0, i_8_507_1570_0, i_8_507_1582_0, i_8_507_1631_0,
    i_8_507_1633_0, i_8_507_1649_0, i_8_507_1702_0, i_8_507_1733_0,
    i_8_507_1775_0, i_8_507_1777_0, i_8_507_1783_0, i_8_507_1786_0,
    i_8_507_1804_0, i_8_507_1817_0, i_8_507_1838_0, i_8_507_1841_0,
    i_8_507_1859_0, i_8_507_1886_0, i_8_507_1945_0, i_8_507_1946_0,
    i_8_507_1972_0, i_8_507_1973_0, i_8_507_2000_0, i_8_507_2044_0,
    i_8_507_2141_0, i_8_507_2155_0, i_8_507_2180_0, i_8_507_2206_0,
    i_8_507_2236_0, i_8_507_2245_0, i_8_507_2270_0, i_8_507_2285_0;
  output o_8_507_0_0;
  assign o_8_507_0_0 = 0;
endmodule



// Benchmark "kernel_8_508" written by ABC on Sun Jul 19 10:11:59 2020

module kernel_8_508 ( 
    i_8_508_116_0, i_8_508_157_0, i_8_508_160_0, i_8_508_262_0,
    i_8_508_270_0, i_8_508_351_0, i_8_508_365_0, i_8_508_368_0,
    i_8_508_429_0, i_8_508_477_0, i_8_508_479_0, i_8_508_480_0,
    i_8_508_482_0, i_8_508_483_0, i_8_508_484_0, i_8_508_485_0,
    i_8_508_492_0, i_8_508_493_0, i_8_508_498_0, i_8_508_522_0,
    i_8_508_523_0, i_8_508_524_0, i_8_508_525_0, i_8_508_527_0,
    i_8_508_624_0, i_8_508_655_0, i_8_508_662_0, i_8_508_696_0,
    i_8_508_702_0, i_8_508_704_0, i_8_508_705_0, i_8_508_707_0,
    i_8_508_748_0, i_8_508_750_0, i_8_508_759_0, i_8_508_760_0,
    i_8_508_761_0, i_8_508_762_0, i_8_508_763_0, i_8_508_764_0,
    i_8_508_837_0, i_8_508_838_0, i_8_508_839_0, i_8_508_840_0,
    i_8_508_842_0, i_8_508_844_0, i_8_508_845_0, i_8_508_879_0,
    i_8_508_954_0, i_8_508_955_0, i_8_508_956_0, i_8_508_990_0,
    i_8_508_991_0, i_8_508_993_0, i_8_508_1226_0, i_8_508_1227_0,
    i_8_508_1229_0, i_8_508_1232_0, i_8_508_1306_0, i_8_508_1353_0,
    i_8_508_1354_0, i_8_508_1355_0, i_8_508_1356_0, i_8_508_1434_0,
    i_8_508_1435_0, i_8_508_1439_0, i_8_508_1587_0, i_8_508_1678_0,
    i_8_508_1679_0, i_8_508_1682_0, i_8_508_1724_0, i_8_508_1726_0,
    i_8_508_1727_0, i_8_508_1738_0, i_8_508_1739_0, i_8_508_1754_0,
    i_8_508_1760_0, i_8_508_1762_0, i_8_508_1763_0, i_8_508_1774_0,
    i_8_508_1818_0, i_8_508_1819_0, i_8_508_1820_0, i_8_508_1821_0,
    i_8_508_1822_0, i_8_508_1823_0, i_8_508_1824_0, i_8_508_1825_0,
    i_8_508_1826_0, i_8_508_1925_0, i_8_508_1969_0, i_8_508_1994_0,
    i_8_508_1995_0, i_8_508_2051_0, i_8_508_2143_0, i_8_508_2145_0,
    i_8_508_2147_0, i_8_508_2149_0, i_8_508_2150_0, i_8_508_2215_0,
    o_8_508_0_0  );
  input  i_8_508_116_0, i_8_508_157_0, i_8_508_160_0, i_8_508_262_0,
    i_8_508_270_0, i_8_508_351_0, i_8_508_365_0, i_8_508_368_0,
    i_8_508_429_0, i_8_508_477_0, i_8_508_479_0, i_8_508_480_0,
    i_8_508_482_0, i_8_508_483_0, i_8_508_484_0, i_8_508_485_0,
    i_8_508_492_0, i_8_508_493_0, i_8_508_498_0, i_8_508_522_0,
    i_8_508_523_0, i_8_508_524_0, i_8_508_525_0, i_8_508_527_0,
    i_8_508_624_0, i_8_508_655_0, i_8_508_662_0, i_8_508_696_0,
    i_8_508_702_0, i_8_508_704_0, i_8_508_705_0, i_8_508_707_0,
    i_8_508_748_0, i_8_508_750_0, i_8_508_759_0, i_8_508_760_0,
    i_8_508_761_0, i_8_508_762_0, i_8_508_763_0, i_8_508_764_0,
    i_8_508_837_0, i_8_508_838_0, i_8_508_839_0, i_8_508_840_0,
    i_8_508_842_0, i_8_508_844_0, i_8_508_845_0, i_8_508_879_0,
    i_8_508_954_0, i_8_508_955_0, i_8_508_956_0, i_8_508_990_0,
    i_8_508_991_0, i_8_508_993_0, i_8_508_1226_0, i_8_508_1227_0,
    i_8_508_1229_0, i_8_508_1232_0, i_8_508_1306_0, i_8_508_1353_0,
    i_8_508_1354_0, i_8_508_1355_0, i_8_508_1356_0, i_8_508_1434_0,
    i_8_508_1435_0, i_8_508_1439_0, i_8_508_1587_0, i_8_508_1678_0,
    i_8_508_1679_0, i_8_508_1682_0, i_8_508_1724_0, i_8_508_1726_0,
    i_8_508_1727_0, i_8_508_1738_0, i_8_508_1739_0, i_8_508_1754_0,
    i_8_508_1760_0, i_8_508_1762_0, i_8_508_1763_0, i_8_508_1774_0,
    i_8_508_1818_0, i_8_508_1819_0, i_8_508_1820_0, i_8_508_1821_0,
    i_8_508_1822_0, i_8_508_1823_0, i_8_508_1824_0, i_8_508_1825_0,
    i_8_508_1826_0, i_8_508_1925_0, i_8_508_1969_0, i_8_508_1994_0,
    i_8_508_1995_0, i_8_508_2051_0, i_8_508_2143_0, i_8_508_2145_0,
    i_8_508_2147_0, i_8_508_2149_0, i_8_508_2150_0, i_8_508_2215_0;
  output o_8_508_0_0;
  assign o_8_508_0_0 = ~((~i_8_508_763_0 & ((~i_8_508_116_0 & ((~i_8_508_157_0 & ~i_8_508_479_0 & ~i_8_508_522_0 & ~i_8_508_759_0 & ~i_8_508_762_0 & i_8_508_838_0 & ~i_8_508_993_0 & ~i_8_508_1727_0) | (~i_8_508_480_0 & ~i_8_508_624_0 & ~i_8_508_1439_0 & i_8_508_1818_0))) | (~i_8_508_480_0 & ~i_8_508_1679_0 & ((~i_8_508_764_0 & i_8_508_1232_0 & ~i_8_508_1434_0 & ~i_8_508_1727_0) | (~i_8_508_1306_0 & ~i_8_508_1763_0 & i_8_508_1824_0 & ~i_8_508_1826_0))) | (~i_8_508_759_0 & ((~i_8_508_160_0 & ~i_8_508_524_0 & ~i_8_508_527_0 & ~i_8_508_761_0 & i_8_508_842_0 & i_8_508_845_0 & ~i_8_508_1678_0 & ~i_8_508_1760_0 & ~i_8_508_1763_0) | (~i_8_508_484_0 & ~i_8_508_498_0 & ~i_8_508_760_0 & i_8_508_1678_0 & i_8_508_2145_0))) | (i_8_508_365_0 & ~i_8_508_522_0 & ~i_8_508_624_0 & i_8_508_842_0 & ~i_8_508_956_0 & ~i_8_508_1738_0 & ~i_8_508_1760_0))) | (~i_8_508_485_0 & ((~i_8_508_479_0 & ~i_8_508_482_0 & ~i_8_508_483_0 & ~i_8_508_522_0 & ~i_8_508_762_0 & i_8_508_1354_0 & ~i_8_508_1682_0 & ~i_8_508_1763_0) | (i_8_508_368_0 & ~i_8_508_760_0 & ~i_8_508_993_0 & i_8_508_1826_0 & ~i_8_508_2051_0))) | (~i_8_508_527_0 & ((~i_8_508_493_0 & ((~i_8_508_270_0 & ~i_8_508_480_0 & ~i_8_508_522_0 & ~i_8_508_624_0 & ~i_8_508_762_0 & i_8_508_1434_0 & ~i_8_508_1679_0) | (~i_8_508_484_0 & ~i_8_508_760_0 & ~i_8_508_761_0 & ~i_8_508_842_0 & i_8_508_1682_0 & ~i_8_508_1760_0 & ~i_8_508_2051_0 & ~i_8_508_2145_0 & ~i_8_508_2215_0))) | (~i_8_508_524_0 & i_8_508_1229_0) | (~i_8_508_764_0 & ~i_8_508_839_0 & ~i_8_508_1356_0 & ~i_8_508_1435_0 & ~i_8_508_1726_0 & ~i_8_508_1754_0 & i_8_508_1925_0))) | (~i_8_508_477_0 & ((~i_8_508_1306_0 & ((~i_8_508_479_0 & ~i_8_508_525_0 & ((~i_8_508_484_0 & i_8_508_696_0 & ~i_8_508_991_0 & ~i_8_508_1355_0 & ~i_8_508_1587_0) | (~i_8_508_480_0 & ~i_8_508_483_0 & ~i_8_508_498_0 & ~i_8_508_624_0 & ~i_8_508_662_0 & ~i_8_508_764_0 & ~i_8_508_990_0 & ~i_8_508_1354_0 & ~i_8_508_1726_0 & ~i_8_508_1739_0 & ~i_8_508_1754_0 & ~i_8_508_1819_0 & ~i_8_508_2143_0))) | (~i_8_508_522_0 & ~i_8_508_759_0 & ~i_8_508_761_0 & ~i_8_508_993_0 & ~i_8_508_1682_0 & ~i_8_508_1739_0 & i_8_508_2150_0))) | (~i_8_508_1587_0 & ((~i_8_508_696_0 & ~i_8_508_761_0 & i_8_508_1435_0 & ~i_8_508_1439_0 & ~i_8_508_1739_0 & i_8_508_1820_0) | (~i_8_508_522_0 & i_8_508_1818_0 & ~i_8_508_1822_0 & i_8_508_2143_0))) | (~i_8_508_480_0 & ~i_8_508_483_0 & i_8_508_750_0) | (~i_8_508_523_0 & i_8_508_624_0 & ~i_8_508_662_0 & i_8_508_705_0 & ~i_8_508_1819_0 & ~i_8_508_2215_0))) | (~i_8_508_524_0 & ((~i_8_508_484_0 & ~i_8_508_525_0 & ~i_8_508_759_0 & ~i_8_508_1354_0 & i_8_508_1821_0) | (~i_8_508_483_0 & i_8_508_492_0 & ~i_8_508_993_0 & ~i_8_508_1754_0 & ~i_8_508_1824_0))) | (~i_8_508_523_0 & ((~i_8_508_157_0 & ((~i_8_508_482_0 & ~i_8_508_483_0 & ~i_8_508_705_0 & ~i_8_508_1738_0 & i_8_508_1819_0) | (~i_8_508_160_0 & i_8_508_1824_0 & ~i_8_508_1969_0))) | (~i_8_508_1678_0 & ~i_8_508_1760_0 & ((~i_8_508_480_0 & ~i_8_508_483_0 & ~i_8_508_761_0 & ~i_8_508_762_0 & ~i_8_508_764_0 & ~i_8_508_1435_0 & ~i_8_508_1682_0 & ~i_8_508_1739_0 & ~i_8_508_1762_0) | (~i_8_508_484_0 & i_8_508_844_0 & ~i_8_508_1439_0 & ~i_8_508_1821_0 & ~i_8_508_1969_0 & ~i_8_508_2215_0))) | (i_8_508_1227_0 & i_8_508_1821_0) | (i_8_508_522_0 & i_8_508_840_0 & ~i_8_508_2051_0))) | (~i_8_508_484_0 & ((~i_8_508_480_0 & ~i_8_508_1587_0 & ((~i_8_508_479_0 & ~i_8_508_990_0 & ~i_8_508_1434_0 & ~i_8_508_1435_0 & ~i_8_508_1754_0 & i_8_508_1774_0) | (~i_8_508_761_0 & i_8_508_1354_0 & i_8_508_2149_0))) | (i_8_508_704_0 & ~i_8_508_761_0 & ~i_8_508_879_0 & ~i_8_508_991_0))) | (~i_8_508_482_0 & ((~i_8_508_750_0 & ~i_8_508_762_0 & ~i_8_508_764_0 & ~i_8_508_1434_0 & ~i_8_508_1678_0 & ~i_8_508_1727_0 & i_8_508_1819_0) | (~i_8_508_157_0 & ~i_8_508_845_0 & i_8_508_1826_0 & i_8_508_2150_0))) | (~i_8_508_157_0 & ~i_8_508_761_0 & ~i_8_508_842_0 & ((i_8_508_705_0 & ~i_8_508_748_0 & ~i_8_508_764_0 & ~i_8_508_991_0 & ~i_8_508_993_0 & ~i_8_508_1354_0 & ~i_8_508_1738_0 & ~i_8_508_1774_0) | (~i_8_508_492_0 & ~i_8_508_762_0 & ~i_8_508_1724_0 & ~i_8_508_1823_0 & i_8_508_1825_0 & ~i_8_508_2215_0))) | (~i_8_508_525_0 & ~i_8_508_1353_0 & i_8_508_1356_0 & ~i_8_508_1439_0 & ~i_8_508_1726_0) | (~i_8_508_624_0 & ~i_8_508_662_0 & ~i_8_508_839_0 & i_8_508_842_0 & ~i_8_508_955_0 & i_8_508_1435_0 & i_8_508_2143_0) | (i_8_508_839_0 & i_8_508_1354_0 & i_8_508_2147_0) | (~i_8_508_990_0 & i_8_508_1824_0 & i_8_508_2149_0));
endmodule



// Benchmark "kernel_8_509" written by ABC on Sun Jul 19 10:12:00 2020

module kernel_8_509 ( 
    i_8_509_12_0, i_8_509_15_0, i_8_509_114_0, i_8_509_139_0,
    i_8_509_142_0, i_8_509_186_0, i_8_509_193_0, i_8_509_302_0,
    i_8_509_322_0, i_8_509_382_0, i_8_509_397_0, i_8_509_400_0,
    i_8_509_504_0, i_8_509_507_0, i_8_509_508_0, i_8_509_525_0,
    i_8_509_526_0, i_8_509_529_0, i_8_509_582_0, i_8_509_597_0,
    i_8_509_616_0, i_8_509_639_0, i_8_509_642_0, i_8_509_661_0,
    i_8_509_696_0, i_8_509_750_0, i_8_509_834_0, i_8_509_837_0,
    i_8_509_850_0, i_8_509_858_0, i_8_509_878_0, i_8_509_891_0,
    i_8_509_894_0, i_8_509_925_0, i_8_509_970_0, i_8_509_973_0,
    i_8_509_1037_0, i_8_509_1038_0, i_8_509_1104_0, i_8_509_1158_0,
    i_8_509_1260_0, i_8_509_1307_0, i_8_509_1317_0, i_8_509_1321_0,
    i_8_509_1362_0, i_8_509_1380_0, i_8_509_1399_0, i_8_509_1401_0,
    i_8_509_1425_0, i_8_509_1440_0, i_8_509_1442_0, i_8_509_1443_0,
    i_8_509_1461_0, i_8_509_1464_0, i_8_509_1468_0, i_8_509_1488_0,
    i_8_509_1503_0, i_8_509_1516_0, i_8_509_1533_0, i_8_509_1548_0,
    i_8_509_1549_0, i_8_509_1561_0, i_8_509_1570_0, i_8_509_1572_0,
    i_8_509_1573_0, i_8_509_1607_0, i_8_509_1678_0, i_8_509_1681_0,
    i_8_509_1686_0, i_8_509_1689_0, i_8_509_1693_0, i_8_509_1694_0,
    i_8_509_1696_0, i_8_509_1698_0, i_8_509_1699_0, i_8_509_1704_0,
    i_8_509_1722_0, i_8_509_1763_0, i_8_509_1765_0, i_8_509_1785_0,
    i_8_509_1794_0, i_8_509_1836_0, i_8_509_1839_0, i_8_509_1840_0,
    i_8_509_1848_0, i_8_509_1884_0, i_8_509_1911_0, i_8_509_1912_0,
    i_8_509_1935_0, i_8_509_1957_0, i_8_509_1962_0, i_8_509_1965_0,
    i_8_509_1971_0, i_8_509_1992_0, i_8_509_2055_0, i_8_509_2172_0,
    i_8_509_2226_0, i_8_509_2247_0, i_8_509_2248_0, i_8_509_2284_0,
    o_8_509_0_0  );
  input  i_8_509_12_0, i_8_509_15_0, i_8_509_114_0, i_8_509_139_0,
    i_8_509_142_0, i_8_509_186_0, i_8_509_193_0, i_8_509_302_0,
    i_8_509_322_0, i_8_509_382_0, i_8_509_397_0, i_8_509_400_0,
    i_8_509_504_0, i_8_509_507_0, i_8_509_508_0, i_8_509_525_0,
    i_8_509_526_0, i_8_509_529_0, i_8_509_582_0, i_8_509_597_0,
    i_8_509_616_0, i_8_509_639_0, i_8_509_642_0, i_8_509_661_0,
    i_8_509_696_0, i_8_509_750_0, i_8_509_834_0, i_8_509_837_0,
    i_8_509_850_0, i_8_509_858_0, i_8_509_878_0, i_8_509_891_0,
    i_8_509_894_0, i_8_509_925_0, i_8_509_970_0, i_8_509_973_0,
    i_8_509_1037_0, i_8_509_1038_0, i_8_509_1104_0, i_8_509_1158_0,
    i_8_509_1260_0, i_8_509_1307_0, i_8_509_1317_0, i_8_509_1321_0,
    i_8_509_1362_0, i_8_509_1380_0, i_8_509_1399_0, i_8_509_1401_0,
    i_8_509_1425_0, i_8_509_1440_0, i_8_509_1442_0, i_8_509_1443_0,
    i_8_509_1461_0, i_8_509_1464_0, i_8_509_1468_0, i_8_509_1488_0,
    i_8_509_1503_0, i_8_509_1516_0, i_8_509_1533_0, i_8_509_1548_0,
    i_8_509_1549_0, i_8_509_1561_0, i_8_509_1570_0, i_8_509_1572_0,
    i_8_509_1573_0, i_8_509_1607_0, i_8_509_1678_0, i_8_509_1681_0,
    i_8_509_1686_0, i_8_509_1689_0, i_8_509_1693_0, i_8_509_1694_0,
    i_8_509_1696_0, i_8_509_1698_0, i_8_509_1699_0, i_8_509_1704_0,
    i_8_509_1722_0, i_8_509_1763_0, i_8_509_1765_0, i_8_509_1785_0,
    i_8_509_1794_0, i_8_509_1836_0, i_8_509_1839_0, i_8_509_1840_0,
    i_8_509_1848_0, i_8_509_1884_0, i_8_509_1911_0, i_8_509_1912_0,
    i_8_509_1935_0, i_8_509_1957_0, i_8_509_1962_0, i_8_509_1965_0,
    i_8_509_1971_0, i_8_509_1992_0, i_8_509_2055_0, i_8_509_2172_0,
    i_8_509_2226_0, i_8_509_2247_0, i_8_509_2248_0, i_8_509_2284_0;
  output o_8_509_0_0;
  assign o_8_509_0_0 = ~((~i_8_509_1442_0 & ((~i_8_509_12_0 & ~i_8_509_1362_0 & ((~i_8_509_15_0 & ~i_8_509_397_0 & ~i_8_509_894_0 & ~i_8_509_1464_0 & ~i_8_509_1503_0 & ~i_8_509_1681_0 & ~i_8_509_1689_0 & ~i_8_509_1694_0 & ~i_8_509_1722_0 & ~i_8_509_1836_0 & ~i_8_509_1935_0 & ~i_8_509_1957_0) | (~i_8_509_114_0 & ~i_8_509_186_0 & ~i_8_509_322_0 & ~i_8_509_1561_0 & ~i_8_509_1573_0 & ~i_8_509_1693_0 & ~i_8_509_2055_0 & ~i_8_509_2247_0))) | (~i_8_509_114_0 & ~i_8_509_525_0 & ~i_8_509_639_0 & ~i_8_509_642_0 & i_8_509_696_0 & ~i_8_509_1686_0 & ~i_8_509_1722_0 & ~i_8_509_1839_0 & i_8_509_1962_0))) | (~i_8_509_582_0 & ((~i_8_509_12_0 & ~i_8_509_639_0 & ((i_8_509_525_0 & ~i_8_509_642_0 & ~i_8_509_925_0 & ~i_8_509_1443_0 & ~i_8_509_1957_0) | (~i_8_509_508_0 & ~i_8_509_891_0 & ~i_8_509_1037_0 & ~i_8_509_1317_0 & ~i_8_509_1401_0 & ~i_8_509_1689_0 & ~i_8_509_2172_0))) | (~i_8_509_139_0 & ~i_8_509_891_0 & ((~i_8_509_193_0 & ~i_8_509_302_0 & ~i_8_509_397_0 & ~i_8_509_750_0 & ~i_8_509_1037_0 & ~i_8_509_1443_0 & ~i_8_509_1678_0 & ~i_8_509_1696_0 & ~i_8_509_1699_0 & ~i_8_509_1884_0) | (i_8_509_193_0 & ~i_8_509_973_0 & ~i_8_509_1440_0 & ~i_8_509_1464_0 & ~i_8_509_1935_0 & i_8_509_2055_0))) | (~i_8_509_142_0 & ~i_8_509_834_0 & ~i_8_509_1399_0 & ~i_8_509_1440_0 & ~i_8_509_1516_0 & ~i_8_509_1549_0 & ~i_8_509_1572_0 & ~i_8_509_1704_0 & ~i_8_509_1794_0 & ~i_8_509_1840_0))) | (~i_8_509_12_0 & ((~i_8_509_322_0 & i_8_509_529_0 & ~i_8_509_973_0 & ~i_8_509_1836_0 & ~i_8_509_1912_0) | (~i_8_509_616_0 & ~i_8_509_639_0 & ~i_8_509_970_0 & ~i_8_509_1038_0 & ~i_8_509_1321_0 & i_8_509_1549_0 & ~i_8_509_1935_0))) | (~i_8_509_1693_0 & ((~i_8_509_322_0 & ((~i_8_509_973_0 & ~i_8_509_1037_0 & i_8_509_1681_0 & ~i_8_509_1765_0 & ~i_8_509_1884_0 & ~i_8_509_1935_0) | (~i_8_509_142_0 & ~i_8_509_639_0 & ~i_8_509_878_0 & ~i_8_509_1038_0 & ~i_8_509_1307_0 & ~i_8_509_1443_0 & ~i_8_509_1461_0 & ~i_8_509_1464_0 & ~i_8_509_1694_0 & ~i_8_509_1722_0 & ~i_8_509_1836_0 & ~i_8_509_1957_0))) | (~i_8_509_1461_0 & ~i_8_509_1839_0 & ((~i_8_509_894_0 & ~i_8_509_1380_0 & ~i_8_509_1443_0 & ~i_8_509_1488_0 & ~i_8_509_1572_0 & ~i_8_509_1794_0 & ~i_8_509_1840_0 & ~i_8_509_1912_0 & ~i_8_509_1935_0 & ~i_8_509_1957_0) | (~i_8_509_400_0 & i_8_509_526_0 & ~i_8_509_891_0 & ~i_8_509_1362_0 & ~i_8_509_1464_0 & ~i_8_509_1694_0 & ~i_8_509_2247_0))))) | (~i_8_509_1440_0 & ((~i_8_509_142_0 & ~i_8_509_1362_0 & ((~i_8_509_397_0 & ~i_8_509_400_0 & ~i_8_509_1686_0 & ~i_8_509_1722_0 & i_8_509_1965_0 & i_8_509_1992_0) | (~i_8_509_639_0 & ~i_8_509_661_0 & ~i_8_509_834_0 & ~i_8_509_1104_0 & ~i_8_509_1704_0 & ~i_8_509_1911_0 & ~i_8_509_1957_0 & ~i_8_509_2284_0))) | (~i_8_509_1992_0 & ((~i_8_509_1104_0 & ((~i_8_509_1037_0 & ~i_8_509_1158_0 & ~i_8_509_1260_0 & ~i_8_509_1516_0 & ~i_8_509_1699_0 & ~i_8_509_1839_0) | (~i_8_509_397_0 & ~i_8_509_894_0 & ~i_8_509_1321_0 & ~i_8_509_1464_0 & ~i_8_509_1573_0 & ~i_8_509_1694_0 & ~i_8_509_1794_0 & ~i_8_509_1935_0))) | (~i_8_509_400_0 & ~i_8_509_696_0 & ~i_8_509_1443_0 & ~i_8_509_1461_0 & ~i_8_509_1573_0 & ~i_8_509_1607_0 & ~i_8_509_1694_0 & ~i_8_509_1911_0 & ~i_8_509_1912_0 & ~i_8_509_2226_0))))) | (i_8_509_616_0 & ~i_8_509_1570_0 & ((~i_8_509_642_0 & ~i_8_509_837_0 & ~i_8_509_1681_0 & ~i_8_509_1698_0 & ~i_8_509_1699_0 & ~i_8_509_1840_0 & ~i_8_509_2226_0) | (~i_8_509_639_0 & ~i_8_509_1317_0 & ~i_8_509_1321_0 & ~i_8_509_1488_0 & ~i_8_509_1516_0 & ~i_8_509_1572_0 & ~i_8_509_1836_0 & ~i_8_509_1965_0 & ~i_8_509_2284_0))) | (~i_8_509_1516_0 & ~i_8_509_1698_0 & ((~i_8_509_508_0 & ~i_8_509_639_0 & ~i_8_509_894_0 & ~i_8_509_1038_0 & ~i_8_509_1573_0 & ~i_8_509_1681_0 & ~i_8_509_1785_0 & ~i_8_509_1839_0) | (~i_8_509_397_0 & ~i_8_509_837_0 & ~i_8_509_891_0 & ~i_8_509_970_0 & ~i_8_509_1686_0 & ~i_8_509_1689_0 & ~i_8_509_1794_0 & ~i_8_509_1957_0))) | (~i_8_509_400_0 & ~i_8_509_507_0 & ~i_8_509_526_0 & ~i_8_509_1461_0 & i_8_509_1678_0 & ~i_8_509_1686_0 & ~i_8_509_1696_0 & ~i_8_509_1911_0 & ~i_8_509_1962_0) | (i_8_509_526_0 & i_8_509_850_0 & i_8_509_1503_0 & ~i_8_509_2248_0));
endmodule



// Benchmark "kernel_8_510" written by ABC on Sun Jul 19 10:12:01 2020

module kernel_8_510 ( 
    i_8_510_22_0, i_8_510_23_0, i_8_510_40_0, i_8_510_77_0, i_8_510_107_0,
    i_8_510_184_0, i_8_510_259_0, i_8_510_346_0, i_8_510_359_0,
    i_8_510_368_0, i_8_510_454_0, i_8_510_499_0, i_8_510_541_0,
    i_8_510_552_0, i_8_510_607_0, i_8_510_634_0, i_8_510_644_0,
    i_8_510_656_0, i_8_510_664_0, i_8_510_671_0, i_8_510_680_0,
    i_8_510_682_0, i_8_510_683_0, i_8_510_707_0, i_8_510_725_0,
    i_8_510_727_0, i_8_510_728_0, i_8_510_755_0, i_8_510_778_0,
    i_8_510_818_0, i_8_510_824_0, i_8_510_835_0, i_8_510_841_0,
    i_8_510_844_0, i_8_510_860_0, i_8_510_869_0, i_8_510_876_0,
    i_8_510_877_0, i_8_510_938_0, i_8_510_980_0, i_8_510_1031_0,
    i_8_510_1034_0, i_8_510_1125_0, i_8_510_1127_0, i_8_510_1128_0,
    i_8_510_1131_0, i_8_510_1171_0, i_8_510_1178_0, i_8_510_1185_0,
    i_8_510_1214_0, i_8_510_1226_0, i_8_510_1267_0, i_8_510_1282_0,
    i_8_510_1286_0, i_8_510_1345_0, i_8_510_1358_0, i_8_510_1367_0,
    i_8_510_1394_0, i_8_510_1397_0, i_8_510_1400_0, i_8_510_1411_0,
    i_8_510_1519_0, i_8_510_1546_0, i_8_510_1551_0, i_8_510_1580_0,
    i_8_510_1592_0, i_8_510_1633_0, i_8_510_1641_0, i_8_510_1668_0,
    i_8_510_1671_0, i_8_510_1700_0, i_8_510_1709_0, i_8_510_1730_0,
    i_8_510_1752_0, i_8_510_1753_0, i_8_510_1769_0, i_8_510_1771_0,
    i_8_510_1775_0, i_8_510_1777_0, i_8_510_1779_0, i_8_510_1796_0,
    i_8_510_1801_0, i_8_510_1817_0, i_8_510_1822_0, i_8_510_1823_0,
    i_8_510_1824_0, i_8_510_1858_0, i_8_510_1859_0, i_8_510_2008_0,
    i_8_510_2109_0, i_8_510_2126_0, i_8_510_2142_0, i_8_510_2150_0,
    i_8_510_2152_0, i_8_510_2229_0, i_8_510_2246_0, i_8_510_2248_0,
    i_8_510_2257_0, i_8_510_2274_0, i_8_510_2293_0,
    o_8_510_0_0  );
  input  i_8_510_22_0, i_8_510_23_0, i_8_510_40_0, i_8_510_77_0,
    i_8_510_107_0, i_8_510_184_0, i_8_510_259_0, i_8_510_346_0,
    i_8_510_359_0, i_8_510_368_0, i_8_510_454_0, i_8_510_499_0,
    i_8_510_541_0, i_8_510_552_0, i_8_510_607_0, i_8_510_634_0,
    i_8_510_644_0, i_8_510_656_0, i_8_510_664_0, i_8_510_671_0,
    i_8_510_680_0, i_8_510_682_0, i_8_510_683_0, i_8_510_707_0,
    i_8_510_725_0, i_8_510_727_0, i_8_510_728_0, i_8_510_755_0,
    i_8_510_778_0, i_8_510_818_0, i_8_510_824_0, i_8_510_835_0,
    i_8_510_841_0, i_8_510_844_0, i_8_510_860_0, i_8_510_869_0,
    i_8_510_876_0, i_8_510_877_0, i_8_510_938_0, i_8_510_980_0,
    i_8_510_1031_0, i_8_510_1034_0, i_8_510_1125_0, i_8_510_1127_0,
    i_8_510_1128_0, i_8_510_1131_0, i_8_510_1171_0, i_8_510_1178_0,
    i_8_510_1185_0, i_8_510_1214_0, i_8_510_1226_0, i_8_510_1267_0,
    i_8_510_1282_0, i_8_510_1286_0, i_8_510_1345_0, i_8_510_1358_0,
    i_8_510_1367_0, i_8_510_1394_0, i_8_510_1397_0, i_8_510_1400_0,
    i_8_510_1411_0, i_8_510_1519_0, i_8_510_1546_0, i_8_510_1551_0,
    i_8_510_1580_0, i_8_510_1592_0, i_8_510_1633_0, i_8_510_1641_0,
    i_8_510_1668_0, i_8_510_1671_0, i_8_510_1700_0, i_8_510_1709_0,
    i_8_510_1730_0, i_8_510_1752_0, i_8_510_1753_0, i_8_510_1769_0,
    i_8_510_1771_0, i_8_510_1775_0, i_8_510_1777_0, i_8_510_1779_0,
    i_8_510_1796_0, i_8_510_1801_0, i_8_510_1817_0, i_8_510_1822_0,
    i_8_510_1823_0, i_8_510_1824_0, i_8_510_1858_0, i_8_510_1859_0,
    i_8_510_2008_0, i_8_510_2109_0, i_8_510_2126_0, i_8_510_2142_0,
    i_8_510_2150_0, i_8_510_2152_0, i_8_510_2229_0, i_8_510_2246_0,
    i_8_510_2248_0, i_8_510_2257_0, i_8_510_2274_0, i_8_510_2293_0;
  output o_8_510_0_0;
  assign o_8_510_0_0 = 0;
endmodule



// Benchmark "kernel_8_511" written by ABC on Sun Jul 19 10:12:02 2020

module kernel_8_511 ( 
    i_8_511_19_0, i_8_511_77_0, i_8_511_85_0, i_8_511_90_0, i_8_511_91_0,
    i_8_511_138_0, i_8_511_139_0, i_8_511_143_0, i_8_511_169_0,
    i_8_511_227_0, i_8_511_263_0, i_8_511_299_0, i_8_511_364_0,
    i_8_511_365_0, i_8_511_368_0, i_8_511_403_0, i_8_511_451_0,
    i_8_511_478_0, i_8_511_490_0, i_8_511_499_0, i_8_511_520_0,
    i_8_511_529_0, i_8_511_557_0, i_8_511_597_0, i_8_511_603_0,
    i_8_511_611_0, i_8_511_625_0, i_8_511_646_0, i_8_511_656_0,
    i_8_511_658_0, i_8_511_683_0, i_8_511_703_0, i_8_511_704_0,
    i_8_511_730_0, i_8_511_766_0, i_8_511_839_0, i_8_511_855_0,
    i_8_511_913_0, i_8_511_940_0, i_8_511_947_0, i_8_511_969_0,
    i_8_511_1114_0, i_8_511_1117_0, i_8_511_1186_0, i_8_511_1229_0,
    i_8_511_1261_0, i_8_511_1321_0, i_8_511_1325_0, i_8_511_1426_0,
    i_8_511_1434_0, i_8_511_1435_0, i_8_511_1468_0, i_8_511_1474_0,
    i_8_511_1475_0, i_8_511_1507_0, i_8_511_1534_0, i_8_511_1535_0,
    i_8_511_1544_0, i_8_511_1548_0, i_8_511_1574_0, i_8_511_1674_0,
    i_8_511_1680_0, i_8_511_1687_0, i_8_511_1700_0, i_8_511_1729_0,
    i_8_511_1750_0, i_8_511_1753_0, i_8_511_1754_0, i_8_511_1781_0,
    i_8_511_1784_0, i_8_511_1798_0, i_8_511_1802_0, i_8_511_1808_0,
    i_8_511_1824_0, i_8_511_1843_0, i_8_511_1844_0, i_8_511_1855_0,
    i_8_511_1857_0, i_8_511_1888_0, i_8_511_1889_0, i_8_511_1903_0,
    i_8_511_1968_0, i_8_511_1969_0, i_8_511_1993_0, i_8_511_1996_0,
    i_8_511_1997_0, i_8_511_2019_0, i_8_511_2087_0, i_8_511_2140_0,
    i_8_511_2145_0, i_8_511_2146_0, i_8_511_2152_0, i_8_511_2216_0,
    i_8_511_2226_0, i_8_511_2227_0, i_8_511_2233_0, i_8_511_2235_0,
    i_8_511_2246_0, i_8_511_2263_0, i_8_511_2287_0,
    o_8_511_0_0  );
  input  i_8_511_19_0, i_8_511_77_0, i_8_511_85_0, i_8_511_90_0,
    i_8_511_91_0, i_8_511_138_0, i_8_511_139_0, i_8_511_143_0,
    i_8_511_169_0, i_8_511_227_0, i_8_511_263_0, i_8_511_299_0,
    i_8_511_364_0, i_8_511_365_0, i_8_511_368_0, i_8_511_403_0,
    i_8_511_451_0, i_8_511_478_0, i_8_511_490_0, i_8_511_499_0,
    i_8_511_520_0, i_8_511_529_0, i_8_511_557_0, i_8_511_597_0,
    i_8_511_603_0, i_8_511_611_0, i_8_511_625_0, i_8_511_646_0,
    i_8_511_656_0, i_8_511_658_0, i_8_511_683_0, i_8_511_703_0,
    i_8_511_704_0, i_8_511_730_0, i_8_511_766_0, i_8_511_839_0,
    i_8_511_855_0, i_8_511_913_0, i_8_511_940_0, i_8_511_947_0,
    i_8_511_969_0, i_8_511_1114_0, i_8_511_1117_0, i_8_511_1186_0,
    i_8_511_1229_0, i_8_511_1261_0, i_8_511_1321_0, i_8_511_1325_0,
    i_8_511_1426_0, i_8_511_1434_0, i_8_511_1435_0, i_8_511_1468_0,
    i_8_511_1474_0, i_8_511_1475_0, i_8_511_1507_0, i_8_511_1534_0,
    i_8_511_1535_0, i_8_511_1544_0, i_8_511_1548_0, i_8_511_1574_0,
    i_8_511_1674_0, i_8_511_1680_0, i_8_511_1687_0, i_8_511_1700_0,
    i_8_511_1729_0, i_8_511_1750_0, i_8_511_1753_0, i_8_511_1754_0,
    i_8_511_1781_0, i_8_511_1784_0, i_8_511_1798_0, i_8_511_1802_0,
    i_8_511_1808_0, i_8_511_1824_0, i_8_511_1843_0, i_8_511_1844_0,
    i_8_511_1855_0, i_8_511_1857_0, i_8_511_1888_0, i_8_511_1889_0,
    i_8_511_1903_0, i_8_511_1968_0, i_8_511_1969_0, i_8_511_1993_0,
    i_8_511_1996_0, i_8_511_1997_0, i_8_511_2019_0, i_8_511_2087_0,
    i_8_511_2140_0, i_8_511_2145_0, i_8_511_2146_0, i_8_511_2152_0,
    i_8_511_2216_0, i_8_511_2226_0, i_8_511_2227_0, i_8_511_2233_0,
    i_8_511_2235_0, i_8_511_2246_0, i_8_511_2263_0, i_8_511_2287_0;
  output o_8_511_0_0;
  assign o_8_511_0_0 = 0;
endmodule



module kernel_8 (i_8_0, i_8_1, i_8_2, i_8_3, i_8_4, i_8_5, i_8_6, i_8_7, i_8_8, i_8_9, i_8_10, i_8_11, i_8_12, i_8_13, i_8_14, i_8_15, i_8_16, i_8_17, i_8_18, i_8_19, i_8_20, i_8_21, i_8_22, i_8_23, i_8_24, i_8_25, i_8_26, i_8_27, i_8_28, i_8_29, i_8_30, i_8_31, i_8_32, i_8_33, i_8_34, i_8_35, i_8_36, i_8_37, i_8_38, i_8_39, i_8_40, i_8_41, i_8_42, i_8_43, i_8_44, i_8_45, i_8_46, i_8_47, i_8_48, i_8_49, i_8_50, i_8_51, i_8_52, i_8_53, i_8_54, i_8_55, i_8_56, i_8_57, i_8_58, i_8_59, i_8_60, i_8_61, i_8_62, i_8_63, i_8_64, i_8_65, i_8_66, i_8_67, i_8_68, i_8_69, i_8_70, i_8_71, i_8_72, i_8_73, i_8_74, i_8_75, i_8_76, i_8_77, i_8_78, i_8_79, i_8_80, i_8_81, i_8_82, i_8_83, i_8_84, i_8_85, i_8_86, i_8_87, i_8_88, i_8_89, i_8_90, i_8_91, i_8_92, i_8_93, i_8_94, i_8_95, i_8_96, i_8_97, i_8_98, i_8_99, i_8_100, i_8_101, i_8_102, i_8_103, i_8_104, i_8_105, i_8_106, i_8_107, i_8_108, i_8_109, i_8_110, i_8_111, i_8_112, i_8_113, i_8_114, i_8_115, i_8_116, i_8_117, i_8_118, i_8_119, i_8_120, i_8_121, i_8_122, i_8_123, i_8_124, i_8_125, i_8_126, i_8_127, i_8_128, i_8_129, i_8_130, i_8_131, i_8_132, i_8_133, i_8_134, i_8_135, i_8_136, i_8_137, i_8_138, i_8_139, i_8_140, i_8_141, i_8_142, i_8_143, i_8_144, i_8_145, i_8_146, i_8_147, i_8_148, i_8_149, i_8_150, i_8_151, i_8_152, i_8_153, i_8_154, i_8_155, i_8_156, i_8_157, i_8_158, i_8_159, i_8_160, i_8_161, i_8_162, i_8_163, i_8_164, i_8_165, i_8_166, i_8_167, i_8_168, i_8_169, i_8_170, i_8_171, i_8_172, i_8_173, i_8_174, i_8_175, i_8_176, i_8_177, i_8_178, i_8_179, i_8_180, i_8_181, i_8_182, i_8_183, i_8_184, i_8_185, i_8_186, i_8_187, i_8_188, i_8_189, i_8_190, i_8_191, i_8_192, i_8_193, i_8_194, i_8_195, i_8_196, i_8_197, i_8_198, i_8_199, i_8_200, i_8_201, i_8_202, i_8_203, i_8_204, i_8_205, i_8_206, i_8_207, i_8_208, i_8_209, i_8_210, i_8_211, i_8_212, i_8_213, i_8_214, i_8_215, i_8_216, i_8_217, i_8_218, i_8_219, i_8_220, i_8_221, i_8_222, i_8_223, i_8_224, i_8_225, i_8_226, i_8_227, i_8_228, i_8_229, i_8_230, i_8_231, i_8_232, i_8_233, i_8_234, i_8_235, i_8_236, i_8_237, i_8_238, i_8_239, i_8_240, i_8_241, i_8_242, i_8_243, i_8_244, i_8_245, i_8_246, i_8_247, i_8_248, i_8_249, i_8_250, i_8_251, i_8_252, i_8_253, i_8_254, i_8_255, i_8_256, i_8_257, i_8_258, i_8_259, i_8_260, i_8_261, i_8_262, i_8_263, i_8_264, i_8_265, i_8_266, i_8_267, i_8_268, i_8_269, i_8_270, i_8_271, i_8_272, i_8_273, i_8_274, i_8_275, i_8_276, i_8_277, i_8_278, i_8_279, i_8_280, i_8_281, i_8_282, i_8_283, i_8_284, i_8_285, i_8_286, i_8_287, i_8_288, i_8_289, i_8_290, i_8_291, i_8_292, i_8_293, i_8_294, i_8_295, i_8_296, i_8_297, i_8_298, i_8_299, i_8_300, i_8_301, i_8_302, i_8_303, i_8_304, i_8_305, i_8_306, i_8_307, i_8_308, i_8_309, i_8_310, i_8_311, i_8_312, i_8_313, i_8_314, i_8_315, i_8_316, i_8_317, i_8_318, i_8_319, i_8_320, i_8_321, i_8_322, i_8_323, i_8_324, i_8_325, i_8_326, i_8_327, i_8_328, i_8_329, i_8_330, i_8_331, i_8_332, i_8_333, i_8_334, i_8_335, i_8_336, i_8_337, i_8_338, i_8_339, i_8_340, i_8_341, i_8_342, i_8_343, i_8_344, i_8_345, i_8_346, i_8_347, i_8_348, i_8_349, i_8_350, i_8_351, i_8_352, i_8_353, i_8_354, i_8_355, i_8_356, i_8_357, i_8_358, i_8_359, i_8_360, i_8_361, i_8_362, i_8_363, i_8_364, i_8_365, i_8_366, i_8_367, i_8_368, i_8_369, i_8_370, i_8_371, i_8_372, i_8_373, i_8_374, i_8_375, i_8_376, i_8_377, i_8_378, i_8_379, i_8_380, i_8_381, i_8_382, i_8_383, i_8_384, i_8_385, i_8_386, i_8_387, i_8_388, i_8_389, i_8_390, i_8_391, i_8_392, i_8_393, i_8_394, i_8_395, i_8_396, i_8_397, i_8_398, i_8_399, i_8_400, i_8_401, i_8_402, i_8_403, i_8_404, i_8_405, i_8_406, i_8_407, i_8_408, i_8_409, i_8_410, i_8_411, i_8_412, i_8_413, i_8_414, i_8_415, i_8_416, i_8_417, i_8_418, i_8_419, i_8_420, i_8_421, i_8_422, i_8_423, i_8_424, i_8_425, i_8_426, i_8_427, i_8_428, i_8_429, i_8_430, i_8_431, i_8_432, i_8_433, i_8_434, i_8_435, i_8_436, i_8_437, i_8_438, i_8_439, i_8_440, i_8_441, i_8_442, i_8_443, i_8_444, i_8_445, i_8_446, i_8_447, i_8_448, i_8_449, i_8_450, i_8_451, i_8_452, i_8_453, i_8_454, i_8_455, i_8_456, i_8_457, i_8_458, i_8_459, i_8_460, i_8_461, i_8_462, i_8_463, i_8_464, i_8_465, i_8_466, i_8_467, i_8_468, i_8_469, i_8_470, i_8_471, i_8_472, i_8_473, i_8_474, i_8_475, i_8_476, i_8_477, i_8_478, i_8_479, i_8_480, i_8_481, i_8_482, i_8_483, i_8_484, i_8_485, i_8_486, i_8_487, i_8_488, i_8_489, i_8_490, i_8_491, i_8_492, i_8_493, i_8_494, i_8_495, i_8_496, i_8_497, i_8_498, i_8_499, i_8_500, i_8_501, i_8_502, i_8_503, i_8_504, i_8_505, i_8_506, i_8_507, i_8_508, i_8_509, i_8_510, i_8_511, i_8_512, i_8_513, i_8_514, i_8_515, i_8_516, i_8_517, i_8_518, i_8_519, i_8_520, i_8_521, i_8_522, i_8_523, i_8_524, i_8_525, i_8_526, i_8_527, i_8_528, i_8_529, i_8_530, i_8_531, i_8_532, i_8_533, i_8_534, i_8_535, i_8_536, i_8_537, i_8_538, i_8_539, i_8_540, i_8_541, i_8_542, i_8_543, i_8_544, i_8_545, i_8_546, i_8_547, i_8_548, i_8_549, i_8_550, i_8_551, i_8_552, i_8_553, i_8_554, i_8_555, i_8_556, i_8_557, i_8_558, i_8_559, i_8_560, i_8_561, i_8_562, i_8_563, i_8_564, i_8_565, i_8_566, i_8_567, i_8_568, i_8_569, i_8_570, i_8_571, i_8_572, i_8_573, i_8_574, i_8_575, i_8_576, i_8_577, i_8_578, i_8_579, i_8_580, i_8_581, i_8_582, i_8_583, i_8_584, i_8_585, i_8_586, i_8_587, i_8_588, i_8_589, i_8_590, i_8_591, i_8_592, i_8_593, i_8_594, i_8_595, i_8_596, i_8_597, i_8_598, i_8_599, i_8_600, i_8_601, i_8_602, i_8_603, i_8_604, i_8_605, i_8_606, i_8_607, i_8_608, i_8_609, i_8_610, i_8_611, i_8_612, i_8_613, i_8_614, i_8_615, i_8_616, i_8_617, i_8_618, i_8_619, i_8_620, i_8_621, i_8_622, i_8_623, i_8_624, i_8_625, i_8_626, i_8_627, i_8_628, i_8_629, i_8_630, i_8_631, i_8_632, i_8_633, i_8_634, i_8_635, i_8_636, i_8_637, i_8_638, i_8_639, i_8_640, i_8_641, i_8_642, i_8_643, i_8_644, i_8_645, i_8_646, i_8_647, i_8_648, i_8_649, i_8_650, i_8_651, i_8_652, i_8_653, i_8_654, i_8_655, i_8_656, i_8_657, i_8_658, i_8_659, i_8_660, i_8_661, i_8_662, i_8_663, i_8_664, i_8_665, i_8_666, i_8_667, i_8_668, i_8_669, i_8_670, i_8_671, i_8_672, i_8_673, i_8_674, i_8_675, i_8_676, i_8_677, i_8_678, i_8_679, i_8_680, i_8_681, i_8_682, i_8_683, i_8_684, i_8_685, i_8_686, i_8_687, i_8_688, i_8_689, i_8_690, i_8_691, i_8_692, i_8_693, i_8_694, i_8_695, i_8_696, i_8_697, i_8_698, i_8_699, i_8_700, i_8_701, i_8_702, i_8_703, i_8_704, i_8_705, i_8_706, i_8_707, i_8_708, i_8_709, i_8_710, i_8_711, i_8_712, i_8_713, i_8_714, i_8_715, i_8_716, i_8_717, i_8_718, i_8_719, i_8_720, i_8_721, i_8_722, i_8_723, i_8_724, i_8_725, i_8_726, i_8_727, i_8_728, i_8_729, i_8_730, i_8_731, i_8_732, i_8_733, i_8_734, i_8_735, i_8_736, i_8_737, i_8_738, i_8_739, i_8_740, i_8_741, i_8_742, i_8_743, i_8_744, i_8_745, i_8_746, i_8_747, i_8_748, i_8_749, i_8_750, i_8_751, i_8_752, i_8_753, i_8_754, i_8_755, i_8_756, i_8_757, i_8_758, i_8_759, i_8_760, i_8_761, i_8_762, i_8_763, i_8_764, i_8_765, i_8_766, i_8_767, i_8_768, i_8_769, i_8_770, i_8_771, i_8_772, i_8_773, i_8_774, i_8_775, i_8_776, i_8_777, i_8_778, i_8_779, i_8_780, i_8_781, i_8_782, i_8_783, i_8_784, i_8_785, i_8_786, i_8_787, i_8_788, i_8_789, i_8_790, i_8_791, i_8_792, i_8_793, i_8_794, i_8_795, i_8_796, i_8_797, i_8_798, i_8_799, i_8_800, i_8_801, i_8_802, i_8_803, i_8_804, i_8_805, i_8_806, i_8_807, i_8_808, i_8_809, i_8_810, i_8_811, i_8_812, i_8_813, i_8_814, i_8_815, i_8_816, i_8_817, i_8_818, i_8_819, i_8_820, i_8_821, i_8_822, i_8_823, i_8_824, i_8_825, i_8_826, i_8_827, i_8_828, i_8_829, i_8_830, i_8_831, i_8_832, i_8_833, i_8_834, i_8_835, i_8_836, i_8_837, i_8_838, i_8_839, i_8_840, i_8_841, i_8_842, i_8_843, i_8_844, i_8_845, i_8_846, i_8_847, i_8_848, i_8_849, i_8_850, i_8_851, i_8_852, i_8_853, i_8_854, i_8_855, i_8_856, i_8_857, i_8_858, i_8_859, i_8_860, i_8_861, i_8_862, i_8_863, i_8_864, i_8_865, i_8_866, i_8_867, i_8_868, i_8_869, i_8_870, i_8_871, i_8_872, i_8_873, i_8_874, i_8_875, i_8_876, i_8_877, i_8_878, i_8_879, i_8_880, i_8_881, i_8_882, i_8_883, i_8_884, i_8_885, i_8_886, i_8_887, i_8_888, i_8_889, i_8_890, i_8_891, i_8_892, i_8_893, i_8_894, i_8_895, i_8_896, i_8_897, i_8_898, i_8_899, i_8_900, i_8_901, i_8_902, i_8_903, i_8_904, i_8_905, i_8_906, i_8_907, i_8_908, i_8_909, i_8_910, i_8_911, i_8_912, i_8_913, i_8_914, i_8_915, i_8_916, i_8_917, i_8_918, i_8_919, i_8_920, i_8_921, i_8_922, i_8_923, i_8_924, i_8_925, i_8_926, i_8_927, i_8_928, i_8_929, i_8_930, i_8_931, i_8_932, i_8_933, i_8_934, i_8_935, i_8_936, i_8_937, i_8_938, i_8_939, i_8_940, i_8_941, i_8_942, i_8_943, i_8_944, i_8_945, i_8_946, i_8_947, i_8_948, i_8_949, i_8_950, i_8_951, i_8_952, i_8_953, i_8_954, i_8_955, i_8_956, i_8_957, i_8_958, i_8_959, i_8_960, i_8_961, i_8_962, i_8_963, i_8_964, i_8_965, i_8_966, i_8_967, i_8_968, i_8_969, i_8_970, i_8_971, i_8_972, i_8_973, i_8_974, i_8_975, i_8_976, i_8_977, i_8_978, i_8_979, i_8_980, i_8_981, i_8_982, i_8_983, i_8_984, i_8_985, i_8_986, i_8_987, i_8_988, i_8_989, i_8_990, i_8_991, i_8_992, i_8_993, i_8_994, i_8_995, i_8_996, i_8_997, i_8_998, i_8_999, i_8_1000, i_8_1001, i_8_1002, i_8_1003, i_8_1004, i_8_1005, i_8_1006, i_8_1007, i_8_1008, i_8_1009, i_8_1010, i_8_1011, i_8_1012, i_8_1013, i_8_1014, i_8_1015, i_8_1016, i_8_1017, i_8_1018, i_8_1019, i_8_1020, i_8_1021, i_8_1022, i_8_1023, i_8_1024, i_8_1025, i_8_1026, i_8_1027, i_8_1028, i_8_1029, i_8_1030, i_8_1031, i_8_1032, i_8_1033, i_8_1034, i_8_1035, i_8_1036, i_8_1037, i_8_1038, i_8_1039, i_8_1040, i_8_1041, i_8_1042, i_8_1043, i_8_1044, i_8_1045, i_8_1046, i_8_1047, i_8_1048, i_8_1049, i_8_1050, i_8_1051, i_8_1052, i_8_1053, i_8_1054, i_8_1055, i_8_1056, i_8_1057, i_8_1058, i_8_1059, i_8_1060, i_8_1061, i_8_1062, i_8_1063, i_8_1064, i_8_1065, i_8_1066, i_8_1067, i_8_1068, i_8_1069, i_8_1070, i_8_1071, i_8_1072, i_8_1073, i_8_1074, i_8_1075, i_8_1076, i_8_1077, i_8_1078, i_8_1079, i_8_1080, i_8_1081, i_8_1082, i_8_1083, i_8_1084, i_8_1085, i_8_1086, i_8_1087, i_8_1088, i_8_1089, i_8_1090, i_8_1091, i_8_1092, i_8_1093, i_8_1094, i_8_1095, i_8_1096, i_8_1097, i_8_1098, i_8_1099, i_8_1100, i_8_1101, i_8_1102, i_8_1103, i_8_1104, i_8_1105, i_8_1106, i_8_1107, i_8_1108, i_8_1109, i_8_1110, i_8_1111, i_8_1112, i_8_1113, i_8_1114, i_8_1115, i_8_1116, i_8_1117, i_8_1118, i_8_1119, i_8_1120, i_8_1121, i_8_1122, i_8_1123, i_8_1124, i_8_1125, i_8_1126, i_8_1127, i_8_1128, i_8_1129, i_8_1130, i_8_1131, i_8_1132, i_8_1133, i_8_1134, i_8_1135, i_8_1136, i_8_1137, i_8_1138, i_8_1139, i_8_1140, i_8_1141, i_8_1142, i_8_1143, i_8_1144, i_8_1145, i_8_1146, i_8_1147, i_8_1148, i_8_1149, i_8_1150, i_8_1151, i_8_1152, i_8_1153, i_8_1154, i_8_1155, i_8_1156, i_8_1157, i_8_1158, i_8_1159, i_8_1160, i_8_1161, i_8_1162, i_8_1163, i_8_1164, i_8_1165, i_8_1166, i_8_1167, i_8_1168, i_8_1169, i_8_1170, i_8_1171, i_8_1172, i_8_1173, i_8_1174, i_8_1175, i_8_1176, i_8_1177, i_8_1178, i_8_1179, i_8_1180, i_8_1181, i_8_1182, i_8_1183, i_8_1184, i_8_1185, i_8_1186, i_8_1187, i_8_1188, i_8_1189, i_8_1190, i_8_1191, i_8_1192, i_8_1193, i_8_1194, i_8_1195, i_8_1196, i_8_1197, i_8_1198, i_8_1199, i_8_1200, i_8_1201, i_8_1202, i_8_1203, i_8_1204, i_8_1205, i_8_1206, i_8_1207, i_8_1208, i_8_1209, i_8_1210, i_8_1211, i_8_1212, i_8_1213, i_8_1214, i_8_1215, i_8_1216, i_8_1217, i_8_1218, i_8_1219, i_8_1220, i_8_1221, i_8_1222, i_8_1223, i_8_1224, i_8_1225, i_8_1226, i_8_1227, i_8_1228, i_8_1229, i_8_1230, i_8_1231, i_8_1232, i_8_1233, i_8_1234, i_8_1235, i_8_1236, i_8_1237, i_8_1238, i_8_1239, i_8_1240, i_8_1241, i_8_1242, i_8_1243, i_8_1244, i_8_1245, i_8_1246, i_8_1247, i_8_1248, i_8_1249, i_8_1250, i_8_1251, i_8_1252, i_8_1253, i_8_1254, i_8_1255, i_8_1256, i_8_1257, i_8_1258, i_8_1259, i_8_1260, i_8_1261, i_8_1262, i_8_1263, i_8_1264, i_8_1265, i_8_1266, i_8_1267, i_8_1268, i_8_1269, i_8_1270, i_8_1271, i_8_1272, i_8_1273, i_8_1274, i_8_1275, i_8_1276, i_8_1277, i_8_1278, i_8_1279, i_8_1280, i_8_1281, i_8_1282, i_8_1283, i_8_1284, i_8_1285, i_8_1286, i_8_1287, i_8_1288, i_8_1289, i_8_1290, i_8_1291, i_8_1292, i_8_1293, i_8_1294, i_8_1295, i_8_1296, i_8_1297, i_8_1298, i_8_1299, i_8_1300, i_8_1301, i_8_1302, i_8_1303, i_8_1304, i_8_1305, i_8_1306, i_8_1307, i_8_1308, i_8_1309, i_8_1310, i_8_1311, i_8_1312, i_8_1313, i_8_1314, i_8_1315, i_8_1316, i_8_1317, i_8_1318, i_8_1319, i_8_1320, i_8_1321, i_8_1322, i_8_1323, i_8_1324, i_8_1325, i_8_1326, i_8_1327, i_8_1328, i_8_1329, i_8_1330, i_8_1331, i_8_1332, i_8_1333, i_8_1334, i_8_1335, i_8_1336, i_8_1337, i_8_1338, i_8_1339, i_8_1340, i_8_1341, i_8_1342, i_8_1343, i_8_1344, i_8_1345, i_8_1346, i_8_1347, i_8_1348, i_8_1349, i_8_1350, i_8_1351, i_8_1352, i_8_1353, i_8_1354, i_8_1355, i_8_1356, i_8_1357, i_8_1358, i_8_1359, i_8_1360, i_8_1361, i_8_1362, i_8_1363, i_8_1364, i_8_1365, i_8_1366, i_8_1367, i_8_1368, i_8_1369, i_8_1370, i_8_1371, i_8_1372, i_8_1373, i_8_1374, i_8_1375, i_8_1376, i_8_1377, i_8_1378, i_8_1379, i_8_1380, i_8_1381, i_8_1382, i_8_1383, i_8_1384, i_8_1385, i_8_1386, i_8_1387, i_8_1388, i_8_1389, i_8_1390, i_8_1391, i_8_1392, i_8_1393, i_8_1394, i_8_1395, i_8_1396, i_8_1397, i_8_1398, i_8_1399, i_8_1400, i_8_1401, i_8_1402, i_8_1403, i_8_1404, i_8_1405, i_8_1406, i_8_1407, i_8_1408, i_8_1409, i_8_1410, i_8_1411, i_8_1412, i_8_1413, i_8_1414, i_8_1415, i_8_1416, i_8_1417, i_8_1418, i_8_1419, i_8_1420, i_8_1421, i_8_1422, i_8_1423, i_8_1424, i_8_1425, i_8_1426, i_8_1427, i_8_1428, i_8_1429, i_8_1430, i_8_1431, i_8_1432, i_8_1433, i_8_1434, i_8_1435, i_8_1436, i_8_1437, i_8_1438, i_8_1439, i_8_1440, i_8_1441, i_8_1442, i_8_1443, i_8_1444, i_8_1445, i_8_1446, i_8_1447, i_8_1448, i_8_1449, i_8_1450, i_8_1451, i_8_1452, i_8_1453, i_8_1454, i_8_1455, i_8_1456, i_8_1457, i_8_1458, i_8_1459, i_8_1460, i_8_1461, i_8_1462, i_8_1463, i_8_1464, i_8_1465, i_8_1466, i_8_1467, i_8_1468, i_8_1469, i_8_1470, i_8_1471, i_8_1472, i_8_1473, i_8_1474, i_8_1475, i_8_1476, i_8_1477, i_8_1478, i_8_1479, i_8_1480, i_8_1481, i_8_1482, i_8_1483, i_8_1484, i_8_1485, i_8_1486, i_8_1487, i_8_1488, i_8_1489, i_8_1490, i_8_1491, i_8_1492, i_8_1493, i_8_1494, i_8_1495, i_8_1496, i_8_1497, i_8_1498, i_8_1499, i_8_1500, i_8_1501, i_8_1502, i_8_1503, i_8_1504, i_8_1505, i_8_1506, i_8_1507, i_8_1508, i_8_1509, i_8_1510, i_8_1511, i_8_1512, i_8_1513, i_8_1514, i_8_1515, i_8_1516, i_8_1517, i_8_1518, i_8_1519, i_8_1520, i_8_1521, i_8_1522, i_8_1523, i_8_1524, i_8_1525, i_8_1526, i_8_1527, i_8_1528, i_8_1529, i_8_1530, i_8_1531, i_8_1532, i_8_1533, i_8_1534, i_8_1535, i_8_1536, i_8_1537, i_8_1538, i_8_1539, i_8_1540, i_8_1541, i_8_1542, i_8_1543, i_8_1544, i_8_1545, i_8_1546, i_8_1547, i_8_1548, i_8_1549, i_8_1550, i_8_1551, i_8_1552, i_8_1553, i_8_1554, i_8_1555, i_8_1556, i_8_1557, i_8_1558, i_8_1559, i_8_1560, i_8_1561, i_8_1562, i_8_1563, i_8_1564, i_8_1565, i_8_1566, i_8_1567, i_8_1568, i_8_1569, i_8_1570, i_8_1571, i_8_1572, i_8_1573, i_8_1574, i_8_1575, i_8_1576, i_8_1577, i_8_1578, i_8_1579, i_8_1580, i_8_1581, i_8_1582, i_8_1583, i_8_1584, i_8_1585, i_8_1586, i_8_1587, i_8_1588, i_8_1589, i_8_1590, i_8_1591, i_8_1592, i_8_1593, i_8_1594, i_8_1595, i_8_1596, i_8_1597, i_8_1598, i_8_1599, i_8_1600, i_8_1601, i_8_1602, i_8_1603, i_8_1604, i_8_1605, i_8_1606, i_8_1607, i_8_1608, i_8_1609, i_8_1610, i_8_1611, i_8_1612, i_8_1613, i_8_1614, i_8_1615, i_8_1616, i_8_1617, i_8_1618, i_8_1619, i_8_1620, i_8_1621, i_8_1622, i_8_1623, i_8_1624, i_8_1625, i_8_1626, i_8_1627, i_8_1628, i_8_1629, i_8_1630, i_8_1631, i_8_1632, i_8_1633, i_8_1634, i_8_1635, i_8_1636, i_8_1637, i_8_1638, i_8_1639, i_8_1640, i_8_1641, i_8_1642, i_8_1643, i_8_1644, i_8_1645, i_8_1646, i_8_1647, i_8_1648, i_8_1649, i_8_1650, i_8_1651, i_8_1652, i_8_1653, i_8_1654, i_8_1655, i_8_1656, i_8_1657, i_8_1658, i_8_1659, i_8_1660, i_8_1661, i_8_1662, i_8_1663, i_8_1664, i_8_1665, i_8_1666, i_8_1667, i_8_1668, i_8_1669, i_8_1670, i_8_1671, i_8_1672, i_8_1673, i_8_1674, i_8_1675, i_8_1676, i_8_1677, i_8_1678, i_8_1679, i_8_1680, i_8_1681, i_8_1682, i_8_1683, i_8_1684, i_8_1685, i_8_1686, i_8_1687, i_8_1688, i_8_1689, i_8_1690, i_8_1691, i_8_1692, i_8_1693, i_8_1694, i_8_1695, i_8_1696, i_8_1697, i_8_1698, i_8_1699, i_8_1700, i_8_1701, i_8_1702, i_8_1703, i_8_1704, i_8_1705, i_8_1706, i_8_1707, i_8_1708, i_8_1709, i_8_1710, i_8_1711, i_8_1712, i_8_1713, i_8_1714, i_8_1715, i_8_1716, i_8_1717, i_8_1718, i_8_1719, i_8_1720, i_8_1721, i_8_1722, i_8_1723, i_8_1724, i_8_1725, i_8_1726, i_8_1727, i_8_1728, i_8_1729, i_8_1730, i_8_1731, i_8_1732, i_8_1733, i_8_1734, i_8_1735, i_8_1736, i_8_1737, i_8_1738, i_8_1739, i_8_1740, i_8_1741, i_8_1742, i_8_1743, i_8_1744, i_8_1745, i_8_1746, i_8_1747, i_8_1748, i_8_1749, i_8_1750, i_8_1751, i_8_1752, i_8_1753, i_8_1754, i_8_1755, i_8_1756, i_8_1757, i_8_1758, i_8_1759, i_8_1760, i_8_1761, i_8_1762, i_8_1763, i_8_1764, i_8_1765, i_8_1766, i_8_1767, i_8_1768, i_8_1769, i_8_1770, i_8_1771, i_8_1772, i_8_1773, i_8_1774, i_8_1775, i_8_1776, i_8_1777, i_8_1778, i_8_1779, i_8_1780, i_8_1781, i_8_1782, i_8_1783, i_8_1784, i_8_1785, i_8_1786, i_8_1787, i_8_1788, i_8_1789, i_8_1790, i_8_1791, i_8_1792, i_8_1793, i_8_1794, i_8_1795, i_8_1796, i_8_1797, i_8_1798, i_8_1799, i_8_1800, i_8_1801, i_8_1802, i_8_1803, i_8_1804, i_8_1805, i_8_1806, i_8_1807, i_8_1808, i_8_1809, i_8_1810, i_8_1811, i_8_1812, i_8_1813, i_8_1814, i_8_1815, i_8_1816, i_8_1817, i_8_1818, i_8_1819, i_8_1820, i_8_1821, i_8_1822, i_8_1823, i_8_1824, i_8_1825, i_8_1826, i_8_1827, i_8_1828, i_8_1829, i_8_1830, i_8_1831, i_8_1832, i_8_1833, i_8_1834, i_8_1835, i_8_1836, i_8_1837, i_8_1838, i_8_1839, i_8_1840, i_8_1841, i_8_1842, i_8_1843, i_8_1844, i_8_1845, i_8_1846, i_8_1847, i_8_1848, i_8_1849, i_8_1850, i_8_1851, i_8_1852, i_8_1853, i_8_1854, i_8_1855, i_8_1856, i_8_1857, i_8_1858, i_8_1859, i_8_1860, i_8_1861, i_8_1862, i_8_1863, i_8_1864, i_8_1865, i_8_1866, i_8_1867, i_8_1868, i_8_1869, i_8_1870, i_8_1871, i_8_1872, i_8_1873, i_8_1874, i_8_1875, i_8_1876, i_8_1877, i_8_1878, i_8_1879, i_8_1880, i_8_1881, i_8_1882, i_8_1883, i_8_1884, i_8_1885, i_8_1886, i_8_1887, i_8_1888, i_8_1889, i_8_1890, i_8_1891, i_8_1892, i_8_1893, i_8_1894, i_8_1895, i_8_1896, i_8_1897, i_8_1898, i_8_1899, i_8_1900, i_8_1901, i_8_1902, i_8_1903, i_8_1904, i_8_1905, i_8_1906, i_8_1907, i_8_1908, i_8_1909, i_8_1910, i_8_1911, i_8_1912, i_8_1913, i_8_1914, i_8_1915, i_8_1916, i_8_1917, i_8_1918, i_8_1919, i_8_1920, i_8_1921, i_8_1922, i_8_1923, i_8_1924, i_8_1925, i_8_1926, i_8_1927, i_8_1928, i_8_1929, i_8_1930, i_8_1931, i_8_1932, i_8_1933, i_8_1934, i_8_1935, i_8_1936, i_8_1937, i_8_1938, i_8_1939, i_8_1940, i_8_1941, i_8_1942, i_8_1943, i_8_1944, i_8_1945, i_8_1946, i_8_1947, i_8_1948, i_8_1949, i_8_1950, i_8_1951, i_8_1952, i_8_1953, i_8_1954, i_8_1955, i_8_1956, i_8_1957, i_8_1958, i_8_1959, i_8_1960, i_8_1961, i_8_1962, i_8_1963, i_8_1964, i_8_1965, i_8_1966, i_8_1967, i_8_1968, i_8_1969, i_8_1970, i_8_1971, i_8_1972, i_8_1973, i_8_1974, i_8_1975, i_8_1976, i_8_1977, i_8_1978, i_8_1979, i_8_1980, i_8_1981, i_8_1982, i_8_1983, i_8_1984, i_8_1985, i_8_1986, i_8_1987, i_8_1988, i_8_1989, i_8_1990, i_8_1991, i_8_1992, i_8_1993, i_8_1994, i_8_1995, i_8_1996, i_8_1997, i_8_1998, i_8_1999, i_8_2000, i_8_2001, i_8_2002, i_8_2003, i_8_2004, i_8_2005, i_8_2006, i_8_2007, i_8_2008, i_8_2009, i_8_2010, i_8_2011, i_8_2012, i_8_2013, i_8_2014, i_8_2015, i_8_2016, i_8_2017, i_8_2018, i_8_2019, i_8_2020, i_8_2021, i_8_2022, i_8_2023, i_8_2024, i_8_2025, i_8_2026, i_8_2027, i_8_2028, i_8_2029, i_8_2030, i_8_2031, i_8_2032, i_8_2033, i_8_2034, i_8_2035, i_8_2036, i_8_2037, i_8_2038, i_8_2039, i_8_2040, i_8_2041, i_8_2042, i_8_2043, i_8_2044, i_8_2045, i_8_2046, i_8_2047, i_8_2048, i_8_2049, i_8_2050, i_8_2051, i_8_2052, i_8_2053, i_8_2054, i_8_2055, i_8_2056, i_8_2057, i_8_2058, i_8_2059, i_8_2060, i_8_2061, i_8_2062, i_8_2063, i_8_2064, i_8_2065, i_8_2066, i_8_2067, i_8_2068, i_8_2069, i_8_2070, i_8_2071, i_8_2072, i_8_2073, i_8_2074, i_8_2075, i_8_2076, i_8_2077, i_8_2078, i_8_2079, i_8_2080, i_8_2081, i_8_2082, i_8_2083, i_8_2084, i_8_2085, i_8_2086, i_8_2087, i_8_2088, i_8_2089, i_8_2090, i_8_2091, i_8_2092, i_8_2093, i_8_2094, i_8_2095, i_8_2096, i_8_2097, i_8_2098, i_8_2099, i_8_2100, i_8_2101, i_8_2102, i_8_2103, i_8_2104, i_8_2105, i_8_2106, i_8_2107, i_8_2108, i_8_2109, i_8_2110, i_8_2111, i_8_2112, i_8_2113, i_8_2114, i_8_2115, i_8_2116, i_8_2117, i_8_2118, i_8_2119, i_8_2120, i_8_2121, i_8_2122, i_8_2123, i_8_2124, i_8_2125, i_8_2126, i_8_2127, i_8_2128, i_8_2129, i_8_2130, i_8_2131, i_8_2132, i_8_2133, i_8_2134, i_8_2135, i_8_2136, i_8_2137, i_8_2138, i_8_2139, i_8_2140, i_8_2141, i_8_2142, i_8_2143, i_8_2144, i_8_2145, i_8_2146, i_8_2147, i_8_2148, i_8_2149, i_8_2150, i_8_2151, i_8_2152, i_8_2153, i_8_2154, i_8_2155, i_8_2156, i_8_2157, i_8_2158, i_8_2159, i_8_2160, i_8_2161, i_8_2162, i_8_2163, i_8_2164, i_8_2165, i_8_2166, i_8_2167, i_8_2168, i_8_2169, i_8_2170, i_8_2171, i_8_2172, i_8_2173, i_8_2174, i_8_2175, i_8_2176, i_8_2177, i_8_2178, i_8_2179, i_8_2180, i_8_2181, i_8_2182, i_8_2183, i_8_2184, i_8_2185, i_8_2186, i_8_2187, i_8_2188, i_8_2189, i_8_2190, i_8_2191, i_8_2192, i_8_2193, i_8_2194, i_8_2195, i_8_2196, i_8_2197, i_8_2198, i_8_2199, i_8_2200, i_8_2201, i_8_2202, i_8_2203, i_8_2204, i_8_2205, i_8_2206, i_8_2207, i_8_2208, i_8_2209, i_8_2210, i_8_2211, i_8_2212, i_8_2213, i_8_2214, i_8_2215, i_8_2216, i_8_2217, i_8_2218, i_8_2219, i_8_2220, i_8_2221, i_8_2222, i_8_2223, i_8_2224, i_8_2225, i_8_2226, i_8_2227, i_8_2228, i_8_2229, i_8_2230, i_8_2231, i_8_2232, i_8_2233, i_8_2234, i_8_2235, i_8_2236, i_8_2237, i_8_2238, i_8_2239, i_8_2240, i_8_2241, i_8_2242, i_8_2243, i_8_2244, i_8_2245, i_8_2246, i_8_2247, i_8_2248, i_8_2249, i_8_2250, i_8_2251, i_8_2252, i_8_2253, i_8_2254, i_8_2255, i_8_2256, i_8_2257, i_8_2258, i_8_2259, i_8_2260, i_8_2261, i_8_2262, i_8_2263, i_8_2264, i_8_2265, i_8_2266, i_8_2267, i_8_2268, i_8_2269, i_8_2270, i_8_2271, i_8_2272, i_8_2273, i_8_2274, i_8_2275, i_8_2276, i_8_2277, i_8_2278, i_8_2279, i_8_2280, i_8_2281, i_8_2282, i_8_2283, i_8_2284, i_8_2285, i_8_2286, i_8_2287, i_8_2288, i_8_2289, i_8_2290, i_8_2291, i_8_2292, i_8_2293, i_8_2294, i_8_2295, i_8_2296, i_8_2297, i_8_2298, i_8_2299, i_8_2300, i_8_2301, i_8_2302, i_8_2303, o_8_0, o_8_1, o_8_2, o_8_3, o_8_4, o_8_5, o_8_6, o_8_7, o_8_8, o_8_9, o_8_10, o_8_11, o_8_12, o_8_13, o_8_14, o_8_15, o_8_16, o_8_17, o_8_18, o_8_19, o_8_20, o_8_21, o_8_22, o_8_23, o_8_24, o_8_25, o_8_26, o_8_27, o_8_28, o_8_29, o_8_30, o_8_31, o_8_32, o_8_33, o_8_34, o_8_35, o_8_36, o_8_37, o_8_38, o_8_39, o_8_40, o_8_41, o_8_42, o_8_43, o_8_44, o_8_45, o_8_46, o_8_47, o_8_48, o_8_49, o_8_50, o_8_51, o_8_52, o_8_53, o_8_54, o_8_55, o_8_56, o_8_57, o_8_58, o_8_59, o_8_60, o_8_61, o_8_62, o_8_63, o_8_64, o_8_65, o_8_66, o_8_67, o_8_68, o_8_69, o_8_70, o_8_71, o_8_72, o_8_73, o_8_74, o_8_75, o_8_76, o_8_77, o_8_78, o_8_79, o_8_80, o_8_81, o_8_82, o_8_83, o_8_84, o_8_85, o_8_86, o_8_87, o_8_88, o_8_89, o_8_90, o_8_91, o_8_92, o_8_93, o_8_94, o_8_95, o_8_96, o_8_97, o_8_98, o_8_99, o_8_100, o_8_101, o_8_102, o_8_103, o_8_104, o_8_105, o_8_106, o_8_107, o_8_108, o_8_109, o_8_110, o_8_111, o_8_112, o_8_113, o_8_114, o_8_115, o_8_116, o_8_117, o_8_118, o_8_119, o_8_120, o_8_121, o_8_122, o_8_123, o_8_124, o_8_125, o_8_126, o_8_127, o_8_128, o_8_129, o_8_130, o_8_131, o_8_132, o_8_133, o_8_134, o_8_135, o_8_136, o_8_137, o_8_138, o_8_139, o_8_140, o_8_141, o_8_142, o_8_143, o_8_144, o_8_145, o_8_146, o_8_147, o_8_148, o_8_149, o_8_150, o_8_151, o_8_152, o_8_153, o_8_154, o_8_155, o_8_156, o_8_157, o_8_158, o_8_159, o_8_160, o_8_161, o_8_162, o_8_163, o_8_164, o_8_165, o_8_166, o_8_167, o_8_168, o_8_169, o_8_170, o_8_171, o_8_172, o_8_173, o_8_174, o_8_175, o_8_176, o_8_177, o_8_178, o_8_179, o_8_180, o_8_181, o_8_182, o_8_183, o_8_184, o_8_185, o_8_186, o_8_187, o_8_188, o_8_189, o_8_190, o_8_191, o_8_192, o_8_193, o_8_194, o_8_195, o_8_196, o_8_197, o_8_198, o_8_199, o_8_200, o_8_201, o_8_202, o_8_203, o_8_204, o_8_205, o_8_206, o_8_207, o_8_208, o_8_209, o_8_210, o_8_211, o_8_212, o_8_213, o_8_214, o_8_215, o_8_216, o_8_217, o_8_218, o_8_219, o_8_220, o_8_221, o_8_222, o_8_223, o_8_224, o_8_225, o_8_226, o_8_227, o_8_228, o_8_229, o_8_230, o_8_231, o_8_232, o_8_233, o_8_234, o_8_235, o_8_236, o_8_237, o_8_238, o_8_239, o_8_240, o_8_241, o_8_242, o_8_243, o_8_244, o_8_245, o_8_246, o_8_247, o_8_248, o_8_249, o_8_250, o_8_251, o_8_252, o_8_253, o_8_254, o_8_255, o_8_256, o_8_257, o_8_258, o_8_259, o_8_260, o_8_261, o_8_262, o_8_263, o_8_264, o_8_265, o_8_266, o_8_267, o_8_268, o_8_269, o_8_270, o_8_271, o_8_272, o_8_273, o_8_274, o_8_275, o_8_276, o_8_277, o_8_278, o_8_279, o_8_280, o_8_281, o_8_282, o_8_283, o_8_284, o_8_285, o_8_286, o_8_287, o_8_288, o_8_289, o_8_290, o_8_291, o_8_292, o_8_293, o_8_294, o_8_295, o_8_296, o_8_297, o_8_298, o_8_299, o_8_300, o_8_301, o_8_302, o_8_303, o_8_304, o_8_305, o_8_306, o_8_307, o_8_308, o_8_309, o_8_310, o_8_311, o_8_312, o_8_313, o_8_314, o_8_315, o_8_316, o_8_317, o_8_318, o_8_319, o_8_320, o_8_321, o_8_322, o_8_323, o_8_324, o_8_325, o_8_326, o_8_327, o_8_328, o_8_329, o_8_330, o_8_331, o_8_332, o_8_333, o_8_334, o_8_335, o_8_336, o_8_337, o_8_338, o_8_339, o_8_340, o_8_341, o_8_342, o_8_343, o_8_344, o_8_345, o_8_346, o_8_347, o_8_348, o_8_349, o_8_350, o_8_351, o_8_352, o_8_353, o_8_354, o_8_355, o_8_356, o_8_357, o_8_358, o_8_359, o_8_360, o_8_361, o_8_362, o_8_363, o_8_364, o_8_365, o_8_366, o_8_367, o_8_368, o_8_369, o_8_370, o_8_371, o_8_372, o_8_373, o_8_374, o_8_375, o_8_376, o_8_377, o_8_378, o_8_379, o_8_380, o_8_381, o_8_382, o_8_383, o_8_384, o_8_385, o_8_386, o_8_387, o_8_388, o_8_389, o_8_390, o_8_391, o_8_392, o_8_393, o_8_394, o_8_395, o_8_396, o_8_397, o_8_398, o_8_399, o_8_400, o_8_401, o_8_402, o_8_403, o_8_404, o_8_405, o_8_406, o_8_407, o_8_408, o_8_409, o_8_410, o_8_411, o_8_412, o_8_413, o_8_414, o_8_415, o_8_416, o_8_417, o_8_418, o_8_419, o_8_420, o_8_421, o_8_422, o_8_423, o_8_424, o_8_425, o_8_426, o_8_427, o_8_428, o_8_429, o_8_430, o_8_431, o_8_432, o_8_433, o_8_434, o_8_435, o_8_436, o_8_437, o_8_438, o_8_439, o_8_440, o_8_441, o_8_442, o_8_443, o_8_444, o_8_445, o_8_446, o_8_447, o_8_448, o_8_449, o_8_450, o_8_451, o_8_452, o_8_453, o_8_454, o_8_455, o_8_456, o_8_457, o_8_458, o_8_459, o_8_460, o_8_461, o_8_462, o_8_463, o_8_464, o_8_465, o_8_466, o_8_467, o_8_468, o_8_469, o_8_470, o_8_471, o_8_472, o_8_473, o_8_474, o_8_475, o_8_476, o_8_477, o_8_478, o_8_479, o_8_480, o_8_481, o_8_482, o_8_483, o_8_484, o_8_485, o_8_486, o_8_487, o_8_488, o_8_489, o_8_490, o_8_491, o_8_492, o_8_493, o_8_494, o_8_495, o_8_496, o_8_497, o_8_498, o_8_499, o_8_500, o_8_501, o_8_502, o_8_503, o_8_504, o_8_505, o_8_506, o_8_507, o_8_508, o_8_509, o_8_510, o_8_511);
input i_8_0, i_8_1, i_8_2, i_8_3, i_8_4, i_8_5, i_8_6, i_8_7, i_8_8, i_8_9, i_8_10, i_8_11, i_8_12, i_8_13, i_8_14, i_8_15, i_8_16, i_8_17, i_8_18, i_8_19, i_8_20, i_8_21, i_8_22, i_8_23, i_8_24, i_8_25, i_8_26, i_8_27, i_8_28, i_8_29, i_8_30, i_8_31, i_8_32, i_8_33, i_8_34, i_8_35, i_8_36, i_8_37, i_8_38, i_8_39, i_8_40, i_8_41, i_8_42, i_8_43, i_8_44, i_8_45, i_8_46, i_8_47, i_8_48, i_8_49, i_8_50, i_8_51, i_8_52, i_8_53, i_8_54, i_8_55, i_8_56, i_8_57, i_8_58, i_8_59, i_8_60, i_8_61, i_8_62, i_8_63, i_8_64, i_8_65, i_8_66, i_8_67, i_8_68, i_8_69, i_8_70, i_8_71, i_8_72, i_8_73, i_8_74, i_8_75, i_8_76, i_8_77, i_8_78, i_8_79, i_8_80, i_8_81, i_8_82, i_8_83, i_8_84, i_8_85, i_8_86, i_8_87, i_8_88, i_8_89, i_8_90, i_8_91, i_8_92, i_8_93, i_8_94, i_8_95, i_8_96, i_8_97, i_8_98, i_8_99, i_8_100, i_8_101, i_8_102, i_8_103, i_8_104, i_8_105, i_8_106, i_8_107, i_8_108, i_8_109, i_8_110, i_8_111, i_8_112, i_8_113, i_8_114, i_8_115, i_8_116, i_8_117, i_8_118, i_8_119, i_8_120, i_8_121, i_8_122, i_8_123, i_8_124, i_8_125, i_8_126, i_8_127, i_8_128, i_8_129, i_8_130, i_8_131, i_8_132, i_8_133, i_8_134, i_8_135, i_8_136, i_8_137, i_8_138, i_8_139, i_8_140, i_8_141, i_8_142, i_8_143, i_8_144, i_8_145, i_8_146, i_8_147, i_8_148, i_8_149, i_8_150, i_8_151, i_8_152, i_8_153, i_8_154, i_8_155, i_8_156, i_8_157, i_8_158, i_8_159, i_8_160, i_8_161, i_8_162, i_8_163, i_8_164, i_8_165, i_8_166, i_8_167, i_8_168, i_8_169, i_8_170, i_8_171, i_8_172, i_8_173, i_8_174, i_8_175, i_8_176, i_8_177, i_8_178, i_8_179, i_8_180, i_8_181, i_8_182, i_8_183, i_8_184, i_8_185, i_8_186, i_8_187, i_8_188, i_8_189, i_8_190, i_8_191, i_8_192, i_8_193, i_8_194, i_8_195, i_8_196, i_8_197, i_8_198, i_8_199, i_8_200, i_8_201, i_8_202, i_8_203, i_8_204, i_8_205, i_8_206, i_8_207, i_8_208, i_8_209, i_8_210, i_8_211, i_8_212, i_8_213, i_8_214, i_8_215, i_8_216, i_8_217, i_8_218, i_8_219, i_8_220, i_8_221, i_8_222, i_8_223, i_8_224, i_8_225, i_8_226, i_8_227, i_8_228, i_8_229, i_8_230, i_8_231, i_8_232, i_8_233, i_8_234, i_8_235, i_8_236, i_8_237, i_8_238, i_8_239, i_8_240, i_8_241, i_8_242, i_8_243, i_8_244, i_8_245, i_8_246, i_8_247, i_8_248, i_8_249, i_8_250, i_8_251, i_8_252, i_8_253, i_8_254, i_8_255, i_8_256, i_8_257, i_8_258, i_8_259, i_8_260, i_8_261, i_8_262, i_8_263, i_8_264, i_8_265, i_8_266, i_8_267, i_8_268, i_8_269, i_8_270, i_8_271, i_8_272, i_8_273, i_8_274, i_8_275, i_8_276, i_8_277, i_8_278, i_8_279, i_8_280, i_8_281, i_8_282, i_8_283, i_8_284, i_8_285, i_8_286, i_8_287, i_8_288, i_8_289, i_8_290, i_8_291, i_8_292, i_8_293, i_8_294, i_8_295, i_8_296, i_8_297, i_8_298, i_8_299, i_8_300, i_8_301, i_8_302, i_8_303, i_8_304, i_8_305, i_8_306, i_8_307, i_8_308, i_8_309, i_8_310, i_8_311, i_8_312, i_8_313, i_8_314, i_8_315, i_8_316, i_8_317, i_8_318, i_8_319, i_8_320, i_8_321, i_8_322, i_8_323, i_8_324, i_8_325, i_8_326, i_8_327, i_8_328, i_8_329, i_8_330, i_8_331, i_8_332, i_8_333, i_8_334, i_8_335, i_8_336, i_8_337, i_8_338, i_8_339, i_8_340, i_8_341, i_8_342, i_8_343, i_8_344, i_8_345, i_8_346, i_8_347, i_8_348, i_8_349, i_8_350, i_8_351, i_8_352, i_8_353, i_8_354, i_8_355, i_8_356, i_8_357, i_8_358, i_8_359, i_8_360, i_8_361, i_8_362, i_8_363, i_8_364, i_8_365, i_8_366, i_8_367, i_8_368, i_8_369, i_8_370, i_8_371, i_8_372, i_8_373, i_8_374, i_8_375, i_8_376, i_8_377, i_8_378, i_8_379, i_8_380, i_8_381, i_8_382, i_8_383, i_8_384, i_8_385, i_8_386, i_8_387, i_8_388, i_8_389, i_8_390, i_8_391, i_8_392, i_8_393, i_8_394, i_8_395, i_8_396, i_8_397, i_8_398, i_8_399, i_8_400, i_8_401, i_8_402, i_8_403, i_8_404, i_8_405, i_8_406, i_8_407, i_8_408, i_8_409, i_8_410, i_8_411, i_8_412, i_8_413, i_8_414, i_8_415, i_8_416, i_8_417, i_8_418, i_8_419, i_8_420, i_8_421, i_8_422, i_8_423, i_8_424, i_8_425, i_8_426, i_8_427, i_8_428, i_8_429, i_8_430, i_8_431, i_8_432, i_8_433, i_8_434, i_8_435, i_8_436, i_8_437, i_8_438, i_8_439, i_8_440, i_8_441, i_8_442, i_8_443, i_8_444, i_8_445, i_8_446, i_8_447, i_8_448, i_8_449, i_8_450, i_8_451, i_8_452, i_8_453, i_8_454, i_8_455, i_8_456, i_8_457, i_8_458, i_8_459, i_8_460, i_8_461, i_8_462, i_8_463, i_8_464, i_8_465, i_8_466, i_8_467, i_8_468, i_8_469, i_8_470, i_8_471, i_8_472, i_8_473, i_8_474, i_8_475, i_8_476, i_8_477, i_8_478, i_8_479, i_8_480, i_8_481, i_8_482, i_8_483, i_8_484, i_8_485, i_8_486, i_8_487, i_8_488, i_8_489, i_8_490, i_8_491, i_8_492, i_8_493, i_8_494, i_8_495, i_8_496, i_8_497, i_8_498, i_8_499, i_8_500, i_8_501, i_8_502, i_8_503, i_8_504, i_8_505, i_8_506, i_8_507, i_8_508, i_8_509, i_8_510, i_8_511, i_8_512, i_8_513, i_8_514, i_8_515, i_8_516, i_8_517, i_8_518, i_8_519, i_8_520, i_8_521, i_8_522, i_8_523, i_8_524, i_8_525, i_8_526, i_8_527, i_8_528, i_8_529, i_8_530, i_8_531, i_8_532, i_8_533, i_8_534, i_8_535, i_8_536, i_8_537, i_8_538, i_8_539, i_8_540, i_8_541, i_8_542, i_8_543, i_8_544, i_8_545, i_8_546, i_8_547, i_8_548, i_8_549, i_8_550, i_8_551, i_8_552, i_8_553, i_8_554, i_8_555, i_8_556, i_8_557, i_8_558, i_8_559, i_8_560, i_8_561, i_8_562, i_8_563, i_8_564, i_8_565, i_8_566, i_8_567, i_8_568, i_8_569, i_8_570, i_8_571, i_8_572, i_8_573, i_8_574, i_8_575, i_8_576, i_8_577, i_8_578, i_8_579, i_8_580, i_8_581, i_8_582, i_8_583, i_8_584, i_8_585, i_8_586, i_8_587, i_8_588, i_8_589, i_8_590, i_8_591, i_8_592, i_8_593, i_8_594, i_8_595, i_8_596, i_8_597, i_8_598, i_8_599, i_8_600, i_8_601, i_8_602, i_8_603, i_8_604, i_8_605, i_8_606, i_8_607, i_8_608, i_8_609, i_8_610, i_8_611, i_8_612, i_8_613, i_8_614, i_8_615, i_8_616, i_8_617, i_8_618, i_8_619, i_8_620, i_8_621, i_8_622, i_8_623, i_8_624, i_8_625, i_8_626, i_8_627, i_8_628, i_8_629, i_8_630, i_8_631, i_8_632, i_8_633, i_8_634, i_8_635, i_8_636, i_8_637, i_8_638, i_8_639, i_8_640, i_8_641, i_8_642, i_8_643, i_8_644, i_8_645, i_8_646, i_8_647, i_8_648, i_8_649, i_8_650, i_8_651, i_8_652, i_8_653, i_8_654, i_8_655, i_8_656, i_8_657, i_8_658, i_8_659, i_8_660, i_8_661, i_8_662, i_8_663, i_8_664, i_8_665, i_8_666, i_8_667, i_8_668, i_8_669, i_8_670, i_8_671, i_8_672, i_8_673, i_8_674, i_8_675, i_8_676, i_8_677, i_8_678, i_8_679, i_8_680, i_8_681, i_8_682, i_8_683, i_8_684, i_8_685, i_8_686, i_8_687, i_8_688, i_8_689, i_8_690, i_8_691, i_8_692, i_8_693, i_8_694, i_8_695, i_8_696, i_8_697, i_8_698, i_8_699, i_8_700, i_8_701, i_8_702, i_8_703, i_8_704, i_8_705, i_8_706, i_8_707, i_8_708, i_8_709, i_8_710, i_8_711, i_8_712, i_8_713, i_8_714, i_8_715, i_8_716, i_8_717, i_8_718, i_8_719, i_8_720, i_8_721, i_8_722, i_8_723, i_8_724, i_8_725, i_8_726, i_8_727, i_8_728, i_8_729, i_8_730, i_8_731, i_8_732, i_8_733, i_8_734, i_8_735, i_8_736, i_8_737, i_8_738, i_8_739, i_8_740, i_8_741, i_8_742, i_8_743, i_8_744, i_8_745, i_8_746, i_8_747, i_8_748, i_8_749, i_8_750, i_8_751, i_8_752, i_8_753, i_8_754, i_8_755, i_8_756, i_8_757, i_8_758, i_8_759, i_8_760, i_8_761, i_8_762, i_8_763, i_8_764, i_8_765, i_8_766, i_8_767, i_8_768, i_8_769, i_8_770, i_8_771, i_8_772, i_8_773, i_8_774, i_8_775, i_8_776, i_8_777, i_8_778, i_8_779, i_8_780, i_8_781, i_8_782, i_8_783, i_8_784, i_8_785, i_8_786, i_8_787, i_8_788, i_8_789, i_8_790, i_8_791, i_8_792, i_8_793, i_8_794, i_8_795, i_8_796, i_8_797, i_8_798, i_8_799, i_8_800, i_8_801, i_8_802, i_8_803, i_8_804, i_8_805, i_8_806, i_8_807, i_8_808, i_8_809, i_8_810, i_8_811, i_8_812, i_8_813, i_8_814, i_8_815, i_8_816, i_8_817, i_8_818, i_8_819, i_8_820, i_8_821, i_8_822, i_8_823, i_8_824, i_8_825, i_8_826, i_8_827, i_8_828, i_8_829, i_8_830, i_8_831, i_8_832, i_8_833, i_8_834, i_8_835, i_8_836, i_8_837, i_8_838, i_8_839, i_8_840, i_8_841, i_8_842, i_8_843, i_8_844, i_8_845, i_8_846, i_8_847, i_8_848, i_8_849, i_8_850, i_8_851, i_8_852, i_8_853, i_8_854, i_8_855, i_8_856, i_8_857, i_8_858, i_8_859, i_8_860, i_8_861, i_8_862, i_8_863, i_8_864, i_8_865, i_8_866, i_8_867, i_8_868, i_8_869, i_8_870, i_8_871, i_8_872, i_8_873, i_8_874, i_8_875, i_8_876, i_8_877, i_8_878, i_8_879, i_8_880, i_8_881, i_8_882, i_8_883, i_8_884, i_8_885, i_8_886, i_8_887, i_8_888, i_8_889, i_8_890, i_8_891, i_8_892, i_8_893, i_8_894, i_8_895, i_8_896, i_8_897, i_8_898, i_8_899, i_8_900, i_8_901, i_8_902, i_8_903, i_8_904, i_8_905, i_8_906, i_8_907, i_8_908, i_8_909, i_8_910, i_8_911, i_8_912, i_8_913, i_8_914, i_8_915, i_8_916, i_8_917, i_8_918, i_8_919, i_8_920, i_8_921, i_8_922, i_8_923, i_8_924, i_8_925, i_8_926, i_8_927, i_8_928, i_8_929, i_8_930, i_8_931, i_8_932, i_8_933, i_8_934, i_8_935, i_8_936, i_8_937, i_8_938, i_8_939, i_8_940, i_8_941, i_8_942, i_8_943, i_8_944, i_8_945, i_8_946, i_8_947, i_8_948, i_8_949, i_8_950, i_8_951, i_8_952, i_8_953, i_8_954, i_8_955, i_8_956, i_8_957, i_8_958, i_8_959, i_8_960, i_8_961, i_8_962, i_8_963, i_8_964, i_8_965, i_8_966, i_8_967, i_8_968, i_8_969, i_8_970, i_8_971, i_8_972, i_8_973, i_8_974, i_8_975, i_8_976, i_8_977, i_8_978, i_8_979, i_8_980, i_8_981, i_8_982, i_8_983, i_8_984, i_8_985, i_8_986, i_8_987, i_8_988, i_8_989, i_8_990, i_8_991, i_8_992, i_8_993, i_8_994, i_8_995, i_8_996, i_8_997, i_8_998, i_8_999, i_8_1000, i_8_1001, i_8_1002, i_8_1003, i_8_1004, i_8_1005, i_8_1006, i_8_1007, i_8_1008, i_8_1009, i_8_1010, i_8_1011, i_8_1012, i_8_1013, i_8_1014, i_8_1015, i_8_1016, i_8_1017, i_8_1018, i_8_1019, i_8_1020, i_8_1021, i_8_1022, i_8_1023, i_8_1024, i_8_1025, i_8_1026, i_8_1027, i_8_1028, i_8_1029, i_8_1030, i_8_1031, i_8_1032, i_8_1033, i_8_1034, i_8_1035, i_8_1036, i_8_1037, i_8_1038, i_8_1039, i_8_1040, i_8_1041, i_8_1042, i_8_1043, i_8_1044, i_8_1045, i_8_1046, i_8_1047, i_8_1048, i_8_1049, i_8_1050, i_8_1051, i_8_1052, i_8_1053, i_8_1054, i_8_1055, i_8_1056, i_8_1057, i_8_1058, i_8_1059, i_8_1060, i_8_1061, i_8_1062, i_8_1063, i_8_1064, i_8_1065, i_8_1066, i_8_1067, i_8_1068, i_8_1069, i_8_1070, i_8_1071, i_8_1072, i_8_1073, i_8_1074, i_8_1075, i_8_1076, i_8_1077, i_8_1078, i_8_1079, i_8_1080, i_8_1081, i_8_1082, i_8_1083, i_8_1084, i_8_1085, i_8_1086, i_8_1087, i_8_1088, i_8_1089, i_8_1090, i_8_1091, i_8_1092, i_8_1093, i_8_1094, i_8_1095, i_8_1096, i_8_1097, i_8_1098, i_8_1099, i_8_1100, i_8_1101, i_8_1102, i_8_1103, i_8_1104, i_8_1105, i_8_1106, i_8_1107, i_8_1108, i_8_1109, i_8_1110, i_8_1111, i_8_1112, i_8_1113, i_8_1114, i_8_1115, i_8_1116, i_8_1117, i_8_1118, i_8_1119, i_8_1120, i_8_1121, i_8_1122, i_8_1123, i_8_1124, i_8_1125, i_8_1126, i_8_1127, i_8_1128, i_8_1129, i_8_1130, i_8_1131, i_8_1132, i_8_1133, i_8_1134, i_8_1135, i_8_1136, i_8_1137, i_8_1138, i_8_1139, i_8_1140, i_8_1141, i_8_1142, i_8_1143, i_8_1144, i_8_1145, i_8_1146, i_8_1147, i_8_1148, i_8_1149, i_8_1150, i_8_1151, i_8_1152, i_8_1153, i_8_1154, i_8_1155, i_8_1156, i_8_1157, i_8_1158, i_8_1159, i_8_1160, i_8_1161, i_8_1162, i_8_1163, i_8_1164, i_8_1165, i_8_1166, i_8_1167, i_8_1168, i_8_1169, i_8_1170, i_8_1171, i_8_1172, i_8_1173, i_8_1174, i_8_1175, i_8_1176, i_8_1177, i_8_1178, i_8_1179, i_8_1180, i_8_1181, i_8_1182, i_8_1183, i_8_1184, i_8_1185, i_8_1186, i_8_1187, i_8_1188, i_8_1189, i_8_1190, i_8_1191, i_8_1192, i_8_1193, i_8_1194, i_8_1195, i_8_1196, i_8_1197, i_8_1198, i_8_1199, i_8_1200, i_8_1201, i_8_1202, i_8_1203, i_8_1204, i_8_1205, i_8_1206, i_8_1207, i_8_1208, i_8_1209, i_8_1210, i_8_1211, i_8_1212, i_8_1213, i_8_1214, i_8_1215, i_8_1216, i_8_1217, i_8_1218, i_8_1219, i_8_1220, i_8_1221, i_8_1222, i_8_1223, i_8_1224, i_8_1225, i_8_1226, i_8_1227, i_8_1228, i_8_1229, i_8_1230, i_8_1231, i_8_1232, i_8_1233, i_8_1234, i_8_1235, i_8_1236, i_8_1237, i_8_1238, i_8_1239, i_8_1240, i_8_1241, i_8_1242, i_8_1243, i_8_1244, i_8_1245, i_8_1246, i_8_1247, i_8_1248, i_8_1249, i_8_1250, i_8_1251, i_8_1252, i_8_1253, i_8_1254, i_8_1255, i_8_1256, i_8_1257, i_8_1258, i_8_1259, i_8_1260, i_8_1261, i_8_1262, i_8_1263, i_8_1264, i_8_1265, i_8_1266, i_8_1267, i_8_1268, i_8_1269, i_8_1270, i_8_1271, i_8_1272, i_8_1273, i_8_1274, i_8_1275, i_8_1276, i_8_1277, i_8_1278, i_8_1279, i_8_1280, i_8_1281, i_8_1282, i_8_1283, i_8_1284, i_8_1285, i_8_1286, i_8_1287, i_8_1288, i_8_1289, i_8_1290, i_8_1291, i_8_1292, i_8_1293, i_8_1294, i_8_1295, i_8_1296, i_8_1297, i_8_1298, i_8_1299, i_8_1300, i_8_1301, i_8_1302, i_8_1303, i_8_1304, i_8_1305, i_8_1306, i_8_1307, i_8_1308, i_8_1309, i_8_1310, i_8_1311, i_8_1312, i_8_1313, i_8_1314, i_8_1315, i_8_1316, i_8_1317, i_8_1318, i_8_1319, i_8_1320, i_8_1321, i_8_1322, i_8_1323, i_8_1324, i_8_1325, i_8_1326, i_8_1327, i_8_1328, i_8_1329, i_8_1330, i_8_1331, i_8_1332, i_8_1333, i_8_1334, i_8_1335, i_8_1336, i_8_1337, i_8_1338, i_8_1339, i_8_1340, i_8_1341, i_8_1342, i_8_1343, i_8_1344, i_8_1345, i_8_1346, i_8_1347, i_8_1348, i_8_1349, i_8_1350, i_8_1351, i_8_1352, i_8_1353, i_8_1354, i_8_1355, i_8_1356, i_8_1357, i_8_1358, i_8_1359, i_8_1360, i_8_1361, i_8_1362, i_8_1363, i_8_1364, i_8_1365, i_8_1366, i_8_1367, i_8_1368, i_8_1369, i_8_1370, i_8_1371, i_8_1372, i_8_1373, i_8_1374, i_8_1375, i_8_1376, i_8_1377, i_8_1378, i_8_1379, i_8_1380, i_8_1381, i_8_1382, i_8_1383, i_8_1384, i_8_1385, i_8_1386, i_8_1387, i_8_1388, i_8_1389, i_8_1390, i_8_1391, i_8_1392, i_8_1393, i_8_1394, i_8_1395, i_8_1396, i_8_1397, i_8_1398, i_8_1399, i_8_1400, i_8_1401, i_8_1402, i_8_1403, i_8_1404, i_8_1405, i_8_1406, i_8_1407, i_8_1408, i_8_1409, i_8_1410, i_8_1411, i_8_1412, i_8_1413, i_8_1414, i_8_1415, i_8_1416, i_8_1417, i_8_1418, i_8_1419, i_8_1420, i_8_1421, i_8_1422, i_8_1423, i_8_1424, i_8_1425, i_8_1426, i_8_1427, i_8_1428, i_8_1429, i_8_1430, i_8_1431, i_8_1432, i_8_1433, i_8_1434, i_8_1435, i_8_1436, i_8_1437, i_8_1438, i_8_1439, i_8_1440, i_8_1441, i_8_1442, i_8_1443, i_8_1444, i_8_1445, i_8_1446, i_8_1447, i_8_1448, i_8_1449, i_8_1450, i_8_1451, i_8_1452, i_8_1453, i_8_1454, i_8_1455, i_8_1456, i_8_1457, i_8_1458, i_8_1459, i_8_1460, i_8_1461, i_8_1462, i_8_1463, i_8_1464, i_8_1465, i_8_1466, i_8_1467, i_8_1468, i_8_1469, i_8_1470, i_8_1471, i_8_1472, i_8_1473, i_8_1474, i_8_1475, i_8_1476, i_8_1477, i_8_1478, i_8_1479, i_8_1480, i_8_1481, i_8_1482, i_8_1483, i_8_1484, i_8_1485, i_8_1486, i_8_1487, i_8_1488, i_8_1489, i_8_1490, i_8_1491, i_8_1492, i_8_1493, i_8_1494, i_8_1495, i_8_1496, i_8_1497, i_8_1498, i_8_1499, i_8_1500, i_8_1501, i_8_1502, i_8_1503, i_8_1504, i_8_1505, i_8_1506, i_8_1507, i_8_1508, i_8_1509, i_8_1510, i_8_1511, i_8_1512, i_8_1513, i_8_1514, i_8_1515, i_8_1516, i_8_1517, i_8_1518, i_8_1519, i_8_1520, i_8_1521, i_8_1522, i_8_1523, i_8_1524, i_8_1525, i_8_1526, i_8_1527, i_8_1528, i_8_1529, i_8_1530, i_8_1531, i_8_1532, i_8_1533, i_8_1534, i_8_1535, i_8_1536, i_8_1537, i_8_1538, i_8_1539, i_8_1540, i_8_1541, i_8_1542, i_8_1543, i_8_1544, i_8_1545, i_8_1546, i_8_1547, i_8_1548, i_8_1549, i_8_1550, i_8_1551, i_8_1552, i_8_1553, i_8_1554, i_8_1555, i_8_1556, i_8_1557, i_8_1558, i_8_1559, i_8_1560, i_8_1561, i_8_1562, i_8_1563, i_8_1564, i_8_1565, i_8_1566, i_8_1567, i_8_1568, i_8_1569, i_8_1570, i_8_1571, i_8_1572, i_8_1573, i_8_1574, i_8_1575, i_8_1576, i_8_1577, i_8_1578, i_8_1579, i_8_1580, i_8_1581, i_8_1582, i_8_1583, i_8_1584, i_8_1585, i_8_1586, i_8_1587, i_8_1588, i_8_1589, i_8_1590, i_8_1591, i_8_1592, i_8_1593, i_8_1594, i_8_1595, i_8_1596, i_8_1597, i_8_1598, i_8_1599, i_8_1600, i_8_1601, i_8_1602, i_8_1603, i_8_1604, i_8_1605, i_8_1606, i_8_1607, i_8_1608, i_8_1609, i_8_1610, i_8_1611, i_8_1612, i_8_1613, i_8_1614, i_8_1615, i_8_1616, i_8_1617, i_8_1618, i_8_1619, i_8_1620, i_8_1621, i_8_1622, i_8_1623, i_8_1624, i_8_1625, i_8_1626, i_8_1627, i_8_1628, i_8_1629, i_8_1630, i_8_1631, i_8_1632, i_8_1633, i_8_1634, i_8_1635, i_8_1636, i_8_1637, i_8_1638, i_8_1639, i_8_1640, i_8_1641, i_8_1642, i_8_1643, i_8_1644, i_8_1645, i_8_1646, i_8_1647, i_8_1648, i_8_1649, i_8_1650, i_8_1651, i_8_1652, i_8_1653, i_8_1654, i_8_1655, i_8_1656, i_8_1657, i_8_1658, i_8_1659, i_8_1660, i_8_1661, i_8_1662, i_8_1663, i_8_1664, i_8_1665, i_8_1666, i_8_1667, i_8_1668, i_8_1669, i_8_1670, i_8_1671, i_8_1672, i_8_1673, i_8_1674, i_8_1675, i_8_1676, i_8_1677, i_8_1678, i_8_1679, i_8_1680, i_8_1681, i_8_1682, i_8_1683, i_8_1684, i_8_1685, i_8_1686, i_8_1687, i_8_1688, i_8_1689, i_8_1690, i_8_1691, i_8_1692, i_8_1693, i_8_1694, i_8_1695, i_8_1696, i_8_1697, i_8_1698, i_8_1699, i_8_1700, i_8_1701, i_8_1702, i_8_1703, i_8_1704, i_8_1705, i_8_1706, i_8_1707, i_8_1708, i_8_1709, i_8_1710, i_8_1711, i_8_1712, i_8_1713, i_8_1714, i_8_1715, i_8_1716, i_8_1717, i_8_1718, i_8_1719, i_8_1720, i_8_1721, i_8_1722, i_8_1723, i_8_1724, i_8_1725, i_8_1726, i_8_1727, i_8_1728, i_8_1729, i_8_1730, i_8_1731, i_8_1732, i_8_1733, i_8_1734, i_8_1735, i_8_1736, i_8_1737, i_8_1738, i_8_1739, i_8_1740, i_8_1741, i_8_1742, i_8_1743, i_8_1744, i_8_1745, i_8_1746, i_8_1747, i_8_1748, i_8_1749, i_8_1750, i_8_1751, i_8_1752, i_8_1753, i_8_1754, i_8_1755, i_8_1756, i_8_1757, i_8_1758, i_8_1759, i_8_1760, i_8_1761, i_8_1762, i_8_1763, i_8_1764, i_8_1765, i_8_1766, i_8_1767, i_8_1768, i_8_1769, i_8_1770, i_8_1771, i_8_1772, i_8_1773, i_8_1774, i_8_1775, i_8_1776, i_8_1777, i_8_1778, i_8_1779, i_8_1780, i_8_1781, i_8_1782, i_8_1783, i_8_1784, i_8_1785, i_8_1786, i_8_1787, i_8_1788, i_8_1789, i_8_1790, i_8_1791, i_8_1792, i_8_1793, i_8_1794, i_8_1795, i_8_1796, i_8_1797, i_8_1798, i_8_1799, i_8_1800, i_8_1801, i_8_1802, i_8_1803, i_8_1804, i_8_1805, i_8_1806, i_8_1807, i_8_1808, i_8_1809, i_8_1810, i_8_1811, i_8_1812, i_8_1813, i_8_1814, i_8_1815, i_8_1816, i_8_1817, i_8_1818, i_8_1819, i_8_1820, i_8_1821, i_8_1822, i_8_1823, i_8_1824, i_8_1825, i_8_1826, i_8_1827, i_8_1828, i_8_1829, i_8_1830, i_8_1831, i_8_1832, i_8_1833, i_8_1834, i_8_1835, i_8_1836, i_8_1837, i_8_1838, i_8_1839, i_8_1840, i_8_1841, i_8_1842, i_8_1843, i_8_1844, i_8_1845, i_8_1846, i_8_1847, i_8_1848, i_8_1849, i_8_1850, i_8_1851, i_8_1852, i_8_1853, i_8_1854, i_8_1855, i_8_1856, i_8_1857, i_8_1858, i_8_1859, i_8_1860, i_8_1861, i_8_1862, i_8_1863, i_8_1864, i_8_1865, i_8_1866, i_8_1867, i_8_1868, i_8_1869, i_8_1870, i_8_1871, i_8_1872, i_8_1873, i_8_1874, i_8_1875, i_8_1876, i_8_1877, i_8_1878, i_8_1879, i_8_1880, i_8_1881, i_8_1882, i_8_1883, i_8_1884, i_8_1885, i_8_1886, i_8_1887, i_8_1888, i_8_1889, i_8_1890, i_8_1891, i_8_1892, i_8_1893, i_8_1894, i_8_1895, i_8_1896, i_8_1897, i_8_1898, i_8_1899, i_8_1900, i_8_1901, i_8_1902, i_8_1903, i_8_1904, i_8_1905, i_8_1906, i_8_1907, i_8_1908, i_8_1909, i_8_1910, i_8_1911, i_8_1912, i_8_1913, i_8_1914, i_8_1915, i_8_1916, i_8_1917, i_8_1918, i_8_1919, i_8_1920, i_8_1921, i_8_1922, i_8_1923, i_8_1924, i_8_1925, i_8_1926, i_8_1927, i_8_1928, i_8_1929, i_8_1930, i_8_1931, i_8_1932, i_8_1933, i_8_1934, i_8_1935, i_8_1936, i_8_1937, i_8_1938, i_8_1939, i_8_1940, i_8_1941, i_8_1942, i_8_1943, i_8_1944, i_8_1945, i_8_1946, i_8_1947, i_8_1948, i_8_1949, i_8_1950, i_8_1951, i_8_1952, i_8_1953, i_8_1954, i_8_1955, i_8_1956, i_8_1957, i_8_1958, i_8_1959, i_8_1960, i_8_1961, i_8_1962, i_8_1963, i_8_1964, i_8_1965, i_8_1966, i_8_1967, i_8_1968, i_8_1969, i_8_1970, i_8_1971, i_8_1972, i_8_1973, i_8_1974, i_8_1975, i_8_1976, i_8_1977, i_8_1978, i_8_1979, i_8_1980, i_8_1981, i_8_1982, i_8_1983, i_8_1984, i_8_1985, i_8_1986, i_8_1987, i_8_1988, i_8_1989, i_8_1990, i_8_1991, i_8_1992, i_8_1993, i_8_1994, i_8_1995, i_8_1996, i_8_1997, i_8_1998, i_8_1999, i_8_2000, i_8_2001, i_8_2002, i_8_2003, i_8_2004, i_8_2005, i_8_2006, i_8_2007, i_8_2008, i_8_2009, i_8_2010, i_8_2011, i_8_2012, i_8_2013, i_8_2014, i_8_2015, i_8_2016, i_8_2017, i_8_2018, i_8_2019, i_8_2020, i_8_2021, i_8_2022, i_8_2023, i_8_2024, i_8_2025, i_8_2026, i_8_2027, i_8_2028, i_8_2029, i_8_2030, i_8_2031, i_8_2032, i_8_2033, i_8_2034, i_8_2035, i_8_2036, i_8_2037, i_8_2038, i_8_2039, i_8_2040, i_8_2041, i_8_2042, i_8_2043, i_8_2044, i_8_2045, i_8_2046, i_8_2047, i_8_2048, i_8_2049, i_8_2050, i_8_2051, i_8_2052, i_8_2053, i_8_2054, i_8_2055, i_8_2056, i_8_2057, i_8_2058, i_8_2059, i_8_2060, i_8_2061, i_8_2062, i_8_2063, i_8_2064, i_8_2065, i_8_2066, i_8_2067, i_8_2068, i_8_2069, i_8_2070, i_8_2071, i_8_2072, i_8_2073, i_8_2074, i_8_2075, i_8_2076, i_8_2077, i_8_2078, i_8_2079, i_8_2080, i_8_2081, i_8_2082, i_8_2083, i_8_2084, i_8_2085, i_8_2086, i_8_2087, i_8_2088, i_8_2089, i_8_2090, i_8_2091, i_8_2092, i_8_2093, i_8_2094, i_8_2095, i_8_2096, i_8_2097, i_8_2098, i_8_2099, i_8_2100, i_8_2101, i_8_2102, i_8_2103, i_8_2104, i_8_2105, i_8_2106, i_8_2107, i_8_2108, i_8_2109, i_8_2110, i_8_2111, i_8_2112, i_8_2113, i_8_2114, i_8_2115, i_8_2116, i_8_2117, i_8_2118, i_8_2119, i_8_2120, i_8_2121, i_8_2122, i_8_2123, i_8_2124, i_8_2125, i_8_2126, i_8_2127, i_8_2128, i_8_2129, i_8_2130, i_8_2131, i_8_2132, i_8_2133, i_8_2134, i_8_2135, i_8_2136, i_8_2137, i_8_2138, i_8_2139, i_8_2140, i_8_2141, i_8_2142, i_8_2143, i_8_2144, i_8_2145, i_8_2146, i_8_2147, i_8_2148, i_8_2149, i_8_2150, i_8_2151, i_8_2152, i_8_2153, i_8_2154, i_8_2155, i_8_2156, i_8_2157, i_8_2158, i_8_2159, i_8_2160, i_8_2161, i_8_2162, i_8_2163, i_8_2164, i_8_2165, i_8_2166, i_8_2167, i_8_2168, i_8_2169, i_8_2170, i_8_2171, i_8_2172, i_8_2173, i_8_2174, i_8_2175, i_8_2176, i_8_2177, i_8_2178, i_8_2179, i_8_2180, i_8_2181, i_8_2182, i_8_2183, i_8_2184, i_8_2185, i_8_2186, i_8_2187, i_8_2188, i_8_2189, i_8_2190, i_8_2191, i_8_2192, i_8_2193, i_8_2194, i_8_2195, i_8_2196, i_8_2197, i_8_2198, i_8_2199, i_8_2200, i_8_2201, i_8_2202, i_8_2203, i_8_2204, i_8_2205, i_8_2206, i_8_2207, i_8_2208, i_8_2209, i_8_2210, i_8_2211, i_8_2212, i_8_2213, i_8_2214, i_8_2215, i_8_2216, i_8_2217, i_8_2218, i_8_2219, i_8_2220, i_8_2221, i_8_2222, i_8_2223, i_8_2224, i_8_2225, i_8_2226, i_8_2227, i_8_2228, i_8_2229, i_8_2230, i_8_2231, i_8_2232, i_8_2233, i_8_2234, i_8_2235, i_8_2236, i_8_2237, i_8_2238, i_8_2239, i_8_2240, i_8_2241, i_8_2242, i_8_2243, i_8_2244, i_8_2245, i_8_2246, i_8_2247, i_8_2248, i_8_2249, i_8_2250, i_8_2251, i_8_2252, i_8_2253, i_8_2254, i_8_2255, i_8_2256, i_8_2257, i_8_2258, i_8_2259, i_8_2260, i_8_2261, i_8_2262, i_8_2263, i_8_2264, i_8_2265, i_8_2266, i_8_2267, i_8_2268, i_8_2269, i_8_2270, i_8_2271, i_8_2272, i_8_2273, i_8_2274, i_8_2275, i_8_2276, i_8_2277, i_8_2278, i_8_2279, i_8_2280, i_8_2281, i_8_2282, i_8_2283, i_8_2284, i_8_2285, i_8_2286, i_8_2287, i_8_2288, i_8_2289, i_8_2290, i_8_2291, i_8_2292, i_8_2293, i_8_2294, i_8_2295, i_8_2296, i_8_2297, i_8_2298, i_8_2299, i_8_2300, i_8_2301, i_8_2302, i_8_2303;
output o_8_0, o_8_1, o_8_2, o_8_3, o_8_4, o_8_5, o_8_6, o_8_7, o_8_8, o_8_9, o_8_10, o_8_11, o_8_12, o_8_13, o_8_14, o_8_15, o_8_16, o_8_17, o_8_18, o_8_19, o_8_20, o_8_21, o_8_22, o_8_23, o_8_24, o_8_25, o_8_26, o_8_27, o_8_28, o_8_29, o_8_30, o_8_31, o_8_32, o_8_33, o_8_34, o_8_35, o_8_36, o_8_37, o_8_38, o_8_39, o_8_40, o_8_41, o_8_42, o_8_43, o_8_44, o_8_45, o_8_46, o_8_47, o_8_48, o_8_49, o_8_50, o_8_51, o_8_52, o_8_53, o_8_54, o_8_55, o_8_56, o_8_57, o_8_58, o_8_59, o_8_60, o_8_61, o_8_62, o_8_63, o_8_64, o_8_65, o_8_66, o_8_67, o_8_68, o_8_69, o_8_70, o_8_71, o_8_72, o_8_73, o_8_74, o_8_75, o_8_76, o_8_77, o_8_78, o_8_79, o_8_80, o_8_81, o_8_82, o_8_83, o_8_84, o_8_85, o_8_86, o_8_87, o_8_88, o_8_89, o_8_90, o_8_91, o_8_92, o_8_93, o_8_94, o_8_95, o_8_96, o_8_97, o_8_98, o_8_99, o_8_100, o_8_101, o_8_102, o_8_103, o_8_104, o_8_105, o_8_106, o_8_107, o_8_108, o_8_109, o_8_110, o_8_111, o_8_112, o_8_113, o_8_114, o_8_115, o_8_116, o_8_117, o_8_118, o_8_119, o_8_120, o_8_121, o_8_122, o_8_123, o_8_124, o_8_125, o_8_126, o_8_127, o_8_128, o_8_129, o_8_130, o_8_131, o_8_132, o_8_133, o_8_134, o_8_135, o_8_136, o_8_137, o_8_138, o_8_139, o_8_140, o_8_141, o_8_142, o_8_143, o_8_144, o_8_145, o_8_146, o_8_147, o_8_148, o_8_149, o_8_150, o_8_151, o_8_152, o_8_153, o_8_154, o_8_155, o_8_156, o_8_157, o_8_158, o_8_159, o_8_160, o_8_161, o_8_162, o_8_163, o_8_164, o_8_165, o_8_166, o_8_167, o_8_168, o_8_169, o_8_170, o_8_171, o_8_172, o_8_173, o_8_174, o_8_175, o_8_176, o_8_177, o_8_178, o_8_179, o_8_180, o_8_181, o_8_182, o_8_183, o_8_184, o_8_185, o_8_186, o_8_187, o_8_188, o_8_189, o_8_190, o_8_191, o_8_192, o_8_193, o_8_194, o_8_195, o_8_196, o_8_197, o_8_198, o_8_199, o_8_200, o_8_201, o_8_202, o_8_203, o_8_204, o_8_205, o_8_206, o_8_207, o_8_208, o_8_209, o_8_210, o_8_211, o_8_212, o_8_213, o_8_214, o_8_215, o_8_216, o_8_217, o_8_218, o_8_219, o_8_220, o_8_221, o_8_222, o_8_223, o_8_224, o_8_225, o_8_226, o_8_227, o_8_228, o_8_229, o_8_230, o_8_231, o_8_232, o_8_233, o_8_234, o_8_235, o_8_236, o_8_237, o_8_238, o_8_239, o_8_240, o_8_241, o_8_242, o_8_243, o_8_244, o_8_245, o_8_246, o_8_247, o_8_248, o_8_249, o_8_250, o_8_251, o_8_252, o_8_253, o_8_254, o_8_255, o_8_256, o_8_257, o_8_258, o_8_259, o_8_260, o_8_261, o_8_262, o_8_263, o_8_264, o_8_265, o_8_266, o_8_267, o_8_268, o_8_269, o_8_270, o_8_271, o_8_272, o_8_273, o_8_274, o_8_275, o_8_276, o_8_277, o_8_278, o_8_279, o_8_280, o_8_281, o_8_282, o_8_283, o_8_284, o_8_285, o_8_286, o_8_287, o_8_288, o_8_289, o_8_290, o_8_291, o_8_292, o_8_293, o_8_294, o_8_295, o_8_296, o_8_297, o_8_298, o_8_299, o_8_300, o_8_301, o_8_302, o_8_303, o_8_304, o_8_305, o_8_306, o_8_307, o_8_308, o_8_309, o_8_310, o_8_311, o_8_312, o_8_313, o_8_314, o_8_315, o_8_316, o_8_317, o_8_318, o_8_319, o_8_320, o_8_321, o_8_322, o_8_323, o_8_324, o_8_325, o_8_326, o_8_327, o_8_328, o_8_329, o_8_330, o_8_331, o_8_332, o_8_333, o_8_334, o_8_335, o_8_336, o_8_337, o_8_338, o_8_339, o_8_340, o_8_341, o_8_342, o_8_343, o_8_344, o_8_345, o_8_346, o_8_347, o_8_348, o_8_349, o_8_350, o_8_351, o_8_352, o_8_353, o_8_354, o_8_355, o_8_356, o_8_357, o_8_358, o_8_359, o_8_360, o_8_361, o_8_362, o_8_363, o_8_364, o_8_365, o_8_366, o_8_367, o_8_368, o_8_369, o_8_370, o_8_371, o_8_372, o_8_373, o_8_374, o_8_375, o_8_376, o_8_377, o_8_378, o_8_379, o_8_380, o_8_381, o_8_382, o_8_383, o_8_384, o_8_385, o_8_386, o_8_387, o_8_388, o_8_389, o_8_390, o_8_391, o_8_392, o_8_393, o_8_394, o_8_395, o_8_396, o_8_397, o_8_398, o_8_399, o_8_400, o_8_401, o_8_402, o_8_403, o_8_404, o_8_405, o_8_406, o_8_407, o_8_408, o_8_409, o_8_410, o_8_411, o_8_412, o_8_413, o_8_414, o_8_415, o_8_416, o_8_417, o_8_418, o_8_419, o_8_420, o_8_421, o_8_422, o_8_423, o_8_424, o_8_425, o_8_426, o_8_427, o_8_428, o_8_429, o_8_430, o_8_431, o_8_432, o_8_433, o_8_434, o_8_435, o_8_436, o_8_437, o_8_438, o_8_439, o_8_440, o_8_441, o_8_442, o_8_443, o_8_444, o_8_445, o_8_446, o_8_447, o_8_448, o_8_449, o_8_450, o_8_451, o_8_452, o_8_453, o_8_454, o_8_455, o_8_456, o_8_457, o_8_458, o_8_459, o_8_460, o_8_461, o_8_462, o_8_463, o_8_464, o_8_465, o_8_466, o_8_467, o_8_468, o_8_469, o_8_470, o_8_471, o_8_472, o_8_473, o_8_474, o_8_475, o_8_476, o_8_477, o_8_478, o_8_479, o_8_480, o_8_481, o_8_482, o_8_483, o_8_484, o_8_485, o_8_486, o_8_487, o_8_488, o_8_489, o_8_490, o_8_491, o_8_492, o_8_493, o_8_494, o_8_495, o_8_496, o_8_497, o_8_498, o_8_499, o_8_500, o_8_501, o_8_502, o_8_503, o_8_504, o_8_505, o_8_506, o_8_507, o_8_508, o_8_509, o_8_510, o_8_511;
	kernel_8_0 k_8_0(i_8_85, i_8_86, i_8_136, i_8_154, i_8_155, i_8_157, i_8_181, i_8_216, i_8_218, i_8_220, i_8_221, i_8_239, i_8_265, i_8_330, i_8_349, i_8_350, i_8_365, i_8_377, i_8_482, i_8_499, i_8_500, i_8_526, i_8_528, i_8_552, i_8_614, i_8_676, i_8_708, i_8_716, i_8_719, i_8_758, i_8_789, i_8_813, i_8_824, i_8_893, i_8_918, i_8_919, i_8_940, i_8_941, i_8_946, i_8_985, i_8_1026, i_8_1029, i_8_1030, i_8_1113, i_8_1114, i_8_1128, i_8_1134, i_8_1154, i_8_1157, i_8_1264, i_8_1305, i_8_1306, i_8_1307, i_8_1342, i_8_1343, i_8_1345, i_8_1346, i_8_1405, i_8_1410, i_8_1434, i_8_1437, i_8_1468, i_8_1474, i_8_1491, i_8_1508, i_8_1541, i_8_1547, i_8_1549, i_8_1550, i_8_1562, i_8_1633, i_8_1647, i_8_1649, i_8_1676, i_8_1678, i_8_1683, i_8_1702, i_8_1747, i_8_1749, i_8_1751, i_8_1786, i_8_1790, i_8_1805, i_8_1821, i_8_1825, i_8_1865, i_8_1868, i_8_1889, i_8_1949, i_8_1988, i_8_2043, i_8_2048, i_8_2216, i_8_2227, i_8_2243, i_8_2271, i_8_2273, i_8_2275, i_8_2290, i_8_2291, o_8_0);
	kernel_8_1 k_8_1(i_8_32, i_8_34, i_8_42, i_8_53, i_8_67, i_8_80, i_8_226, i_8_233, i_8_280, i_8_329, i_8_364, i_8_386, i_8_389, i_8_400, i_8_415, i_8_416, i_8_493, i_8_506, i_8_529, i_8_579, i_8_592, i_8_607, i_8_635, i_8_637, i_8_662, i_8_669, i_8_673, i_8_679, i_8_680, i_8_700, i_8_738, i_8_825, i_8_826, i_8_837, i_8_841, i_8_843, i_8_844, i_8_856, i_8_861, i_8_868, i_8_968, i_8_1012, i_8_1056, i_8_1071, i_8_1102, i_8_1105, i_8_1144, i_8_1189, i_8_1199, i_8_1240, i_8_1243, i_8_1263, i_8_1283, i_8_1300, i_8_1301, i_8_1316, i_8_1320, i_8_1363, i_8_1400, i_8_1439, i_8_1440, i_8_1445, i_8_1460, i_8_1464, i_8_1479, i_8_1480, i_8_1483, i_8_1505, i_8_1524, i_8_1542, i_8_1545, i_8_1571, i_8_1573, i_8_1633, i_8_1659, i_8_1687, i_8_1696, i_8_1767, i_8_1781, i_8_1782, i_8_1785, i_8_1793, i_8_1804, i_8_1858, i_8_1885, i_8_1929, i_8_1960, i_8_1984, i_8_1993, i_8_1996, i_8_2038, i_8_2047, i_8_2058, i_8_2110, i_8_2137, i_8_2143, i_8_2146, i_8_2155, i_8_2156, i_8_2248, o_8_1);
	kernel_8_2 k_8_2(i_8_2, i_8_11, i_8_40, i_8_55, i_8_73, i_8_101, i_8_135, i_8_181, i_8_192, i_8_195, i_8_225, i_8_228, i_8_306, i_8_315, i_8_321, i_8_361, i_8_368, i_8_388, i_8_493, i_8_504, i_8_508, i_8_509, i_8_534, i_8_550, i_8_568, i_8_577, i_8_622, i_8_640, i_8_675, i_8_697, i_8_704, i_8_747, i_8_865, i_8_866, i_8_873, i_8_874, i_8_949, i_8_950, i_8_977, i_8_978, i_8_1009, i_8_1066, i_8_1074, i_8_1099, i_8_1127, i_8_1203, i_8_1228, i_8_1243, i_8_1263, i_8_1266, i_8_1268, i_8_1282, i_8_1301, i_8_1328, i_8_1360, i_8_1403, i_8_1433, i_8_1477, i_8_1479, i_8_1488, i_8_1513, i_8_1515, i_8_1545, i_8_1567, i_8_1577, i_8_1580, i_8_1595, i_8_1598, i_8_1632, i_8_1634, i_8_1651, i_8_1674, i_8_1701, i_8_1702, i_8_1747, i_8_1753, i_8_1756, i_8_1757, i_8_1773, i_8_1787, i_8_1790, i_8_1809, i_8_1810, i_8_1824, i_8_1837, i_8_1946, i_8_1949, i_8_1953, i_8_1954, i_8_1995, i_8_2038, i_8_2070, i_8_2097, i_8_2098, i_8_2142, i_8_2172, i_8_2227, i_8_2281, i_8_2288, i_8_2292, o_8_2);
	kernel_8_3 k_8_3(i_8_72, i_8_103, i_8_126, i_8_147, i_8_202, i_8_208, i_8_262, i_8_273, i_8_275, i_8_318, i_8_378, i_8_383, i_8_397, i_8_420, i_8_441, i_8_476, i_8_492, i_8_507, i_8_514, i_8_577, i_8_580, i_8_630, i_8_665, i_8_668, i_8_679, i_8_702, i_8_800, i_8_838, i_8_841, i_8_847, i_8_910, i_8_926, i_8_948, i_8_955, i_8_966, i_8_1083, i_8_1111, i_8_1128, i_8_1153, i_8_1198, i_8_1224, i_8_1225, i_8_1269, i_8_1270, i_8_1281, i_8_1297, i_8_1335, i_8_1350, i_8_1385, i_8_1386, i_8_1387, i_8_1388, i_8_1405, i_8_1410, i_8_1461, i_8_1470, i_8_1478, i_8_1485, i_8_1494, i_8_1495, i_8_1521, i_8_1536, i_8_1537, i_8_1549, i_8_1650, i_8_1652, i_8_1675, i_8_1678, i_8_1686, i_8_1693, i_8_1701, i_8_1746, i_8_1747, i_8_1791, i_8_1803, i_8_1820, i_8_1821, i_8_1826, i_8_1841, i_8_1864, i_8_1926, i_8_1962, i_8_1992, i_8_2011, i_8_2044, i_8_2046, i_8_2136, i_8_2143, i_8_2149, i_8_2169, i_8_2170, i_8_2178, i_8_2226, i_8_2232, i_8_2234, i_8_2253, i_8_2256, i_8_2280, i_8_2295, i_8_2296, o_8_3);
	kernel_8_4 k_8_4(i_8_28, i_8_47, i_8_49, i_8_108, i_8_109, i_8_111, i_8_180, i_8_181, i_8_182, i_8_185, i_8_191, i_8_220, i_8_221, i_8_237, i_8_238, i_8_256, i_8_263, i_8_300, i_8_343, i_8_345, i_8_362, i_8_364, i_8_378, i_8_379, i_8_387, i_8_388, i_8_477, i_8_478, i_8_550, i_8_596, i_8_599, i_8_615, i_8_631, i_8_665, i_8_685, i_8_704, i_8_707, i_8_758, i_8_759, i_8_884, i_8_919, i_8_937, i_8_938, i_8_991, i_8_1089, i_8_1110, i_8_1117, i_8_1179, i_8_1180, i_8_1181, i_8_1189, i_8_1283, i_8_1288, i_8_1314, i_8_1334, i_8_1407, i_8_1409, i_8_1434, i_8_1435, i_8_1455, i_8_1467, i_8_1468, i_8_1476, i_8_1487, i_8_1506, i_8_1507, i_8_1542, i_8_1549, i_8_1554, i_8_1561, i_8_1631, i_8_1648, i_8_1651, i_8_1674, i_8_1675, i_8_1720, i_8_1724, i_8_1729, i_8_1739, i_8_1760, i_8_1778, i_8_1818, i_8_1819, i_8_1821, i_8_1827, i_8_1831, i_8_1857, i_8_1858, i_8_1864, i_8_1901, i_8_1948, i_8_1993, i_8_1996, i_8_2044, i_8_2143, i_8_2219, i_8_2245, i_8_2246, i_8_2281, i_8_2297, o_8_4);
	kernel_8_5 k_8_5(i_8_3, i_8_66, i_8_67, i_8_79, i_8_84, i_8_85, i_8_190, i_8_193, i_8_210, i_8_223, i_8_238, i_8_361, i_8_364, i_8_414, i_8_481, i_8_498, i_8_516, i_8_517, i_8_525, i_8_582, i_8_603, i_8_612, i_8_615, i_8_624, i_8_625, i_8_636, i_8_672, i_8_705, i_8_708, i_8_760, i_8_789, i_8_795, i_8_814, i_8_835, i_8_843, i_8_844, i_8_858, i_8_937, i_8_959, i_8_999, i_8_1002, i_8_1057, i_8_1059, i_8_1074, i_8_1114, i_8_1141, i_8_1168, i_8_1182, i_8_1183, i_8_1192, i_8_1219, i_8_1227, i_8_1236, i_8_1237, i_8_1239, i_8_1249, i_8_1275, i_8_1286, i_8_1300, i_8_1345, i_8_1348, i_8_1382, i_8_1407, i_8_1410, i_8_1497, i_8_1530, i_8_1533, i_8_1633, i_8_1650, i_8_1668, i_8_1689, i_8_1704, i_8_1741, i_8_1764, i_8_1818, i_8_1821, i_8_1839, i_8_1848, i_8_1857, i_8_1884, i_8_1885, i_8_1888, i_8_1896, i_8_2011, i_8_2037, i_8_2044, i_8_2047, i_8_2065, i_8_2104, i_8_2118, i_8_2119, i_8_2122, i_8_2146, i_8_2169, i_8_2174, i_8_2211, i_8_2214, i_8_2257, i_8_2290, i_8_2299, o_8_5);
	kernel_8_6 k_8_6(i_8_12, i_8_37, i_8_40, i_8_50, i_8_57, i_8_64, i_8_68, i_8_256, i_8_262, i_8_305, i_8_319, i_8_381, i_8_382, i_8_391, i_8_435, i_8_453, i_8_454, i_8_460, i_8_486, i_8_490, i_8_504, i_8_622, i_8_662, i_8_665, i_8_684, i_8_693, i_8_695, i_8_698, i_8_708, i_8_748, i_8_844, i_8_874, i_8_875, i_8_877, i_8_895, i_8_990, i_8_993, i_8_1034, i_8_1051, i_8_1054, i_8_1071, i_8_1114, i_8_1136, i_8_1198, i_8_1201, i_8_1225, i_8_1236, i_8_1237, i_8_1264, i_8_1265, i_8_1276, i_8_1282, i_8_1296, i_8_1328, i_8_1335, i_8_1354, i_8_1381, i_8_1383, i_8_1399, i_8_1404, i_8_1438, i_8_1461, i_8_1462, i_8_1486, i_8_1515, i_8_1530, i_8_1550, i_8_1623, i_8_1631, i_8_1632, i_8_1702, i_8_1746, i_8_1748, i_8_1754, i_8_1776, i_8_1791, i_8_1795, i_8_1812, i_8_1822, i_8_1836, i_8_1882, i_8_1903, i_8_1909, i_8_1911, i_8_1913, i_8_1936, i_8_1980, i_8_1992, i_8_1994, i_8_2038, i_8_2043, i_8_2044, i_8_2048, i_8_2055, i_8_2070, i_8_2106, i_8_2110, i_8_2142, i_8_2144, i_8_2296, o_8_6);
	kernel_8_7 k_8_7(i_8_12, i_8_13, i_8_46, i_8_52, i_8_78, i_8_139, i_8_159, i_8_211, i_8_237, i_8_262, i_8_264, i_8_265, i_8_285, i_8_322, i_8_328, i_8_336, i_8_337, i_8_381, i_8_384, i_8_400, i_8_417, i_8_420, i_8_421, i_8_471, i_8_510, i_8_556, i_8_573, i_8_574, i_8_580, i_8_660, i_8_687, i_8_688, i_8_697, i_8_753, i_8_807, i_8_822, i_8_894, i_8_895, i_8_898, i_8_919, i_8_966, i_8_975, i_8_976, i_8_1011, i_8_1012, i_8_1039, i_8_1041, i_8_1110, i_8_1113, i_8_1114, i_8_1239, i_8_1249, i_8_1260, i_8_1263, i_8_1267, i_8_1272, i_8_1273, i_8_1275, i_8_1282, i_8_1302, i_8_1303, i_8_1314, i_8_1315, i_8_1335, i_8_1338, i_8_1425, i_8_1426, i_8_1434, i_8_1437, i_8_1467, i_8_1510, i_8_1524, i_8_1525, i_8_1527, i_8_1528, i_8_1551, i_8_1554, i_8_1560, i_8_1572, i_8_1632, i_8_1668, i_8_1669, i_8_1722, i_8_1723, i_8_1726, i_8_1749, i_8_1768, i_8_1783, i_8_1797, i_8_1900, i_8_1939, i_8_1959, i_8_1969, i_8_1993, i_8_2154, i_8_2176, i_8_2229, i_8_2246, i_8_2249, i_8_2294, o_8_7);
	kernel_8_8 k_8_8(i_8_31, i_8_40, i_8_54, i_8_57, i_8_88, i_8_111, i_8_112, i_8_153, i_8_165, i_8_226, i_8_241, i_8_333, i_8_335, i_8_348, i_8_372, i_8_375, i_8_376, i_8_450, i_8_454, i_8_469, i_8_523, i_8_525, i_8_529, i_8_530, i_8_540, i_8_543, i_8_551, i_8_556, i_8_570, i_8_571, i_8_613, i_8_616, i_8_687, i_8_688, i_8_705, i_8_706, i_8_775, i_8_777, i_8_786, i_8_800, i_8_810, i_8_814, i_8_844, i_8_850, i_8_858, i_8_916, i_8_1056, i_8_1113, i_8_1114, i_8_1115, i_8_1124, i_8_1160, i_8_1182, i_8_1240, i_8_1267, i_8_1291, i_8_1292, i_8_1299, i_8_1308, i_8_1317, i_8_1323, i_8_1407, i_8_1490, i_8_1588, i_8_1596, i_8_1630, i_8_1651, i_8_1653, i_8_1654, i_8_1671, i_8_1696, i_8_1719, i_8_1722, i_8_1737, i_8_1741, i_8_1745, i_8_1749, i_8_1790, i_8_1840, i_8_1847, i_8_1856, i_8_1857, i_8_1884, i_8_1888, i_8_1946, i_8_1993, i_8_1997, i_8_2020, i_8_2022, i_8_2023, i_8_2037, i_8_2043, i_8_2044, i_8_2047, i_8_2050, i_8_2092, i_8_2123, i_8_2172, i_8_2233, i_8_2299, o_8_8);
	kernel_8_9 k_8_9(i_8_46, i_8_58, i_8_59, i_8_85, i_8_87, i_8_88, i_8_106, i_8_140, i_8_142, i_8_143, i_8_187, i_8_188, i_8_252, i_8_256, i_8_259, i_8_303, i_8_304, i_8_311, i_8_331, i_8_346, i_8_378, i_8_401, i_8_422, i_8_445, i_8_478, i_8_479, i_8_480, i_8_482, i_8_484, i_8_490, i_8_501, i_8_528, i_8_530, i_8_548, i_8_579, i_8_609, i_8_678, i_8_705, i_8_714, i_8_715, i_8_781, i_8_850, i_8_922, i_8_937, i_8_952, i_8_955, i_8_994, i_8_995, i_8_1030, i_8_1031, i_8_1075, i_8_1079, i_8_1112, i_8_1127, i_8_1243, i_8_1265, i_8_1270, i_8_1271, i_8_1274, i_8_1283, i_8_1306, i_8_1307, i_8_1390, i_8_1479, i_8_1492, i_8_1503, i_8_1521, i_8_1543, i_8_1544, i_8_1550, i_8_1574, i_8_1579, i_8_1653, i_8_1669, i_8_1684, i_8_1707, i_8_1716, i_8_1746, i_8_1750, i_8_1774, i_8_1779, i_8_1780, i_8_1804, i_8_1821, i_8_1894, i_8_1917, i_8_1920, i_8_2129, i_8_2130, i_8_2131, i_8_2143, i_8_2148, i_8_2214, i_8_2215, i_8_2218, i_8_2229, i_8_2235, i_8_2242, i_8_2281, i_8_2282, o_8_9);
	kernel_8_10 k_8_10(i_8_3, i_8_22, i_8_40, i_8_94, i_8_193, i_8_201, i_8_246, i_8_256, i_8_277, i_8_283, i_8_352, i_8_355, i_8_356, i_8_358, i_8_367, i_8_426, i_8_457, i_8_516, i_8_517, i_8_527, i_8_528, i_8_556, i_8_594, i_8_612, i_8_613, i_8_616, i_8_622, i_8_632, i_8_633, i_8_666, i_8_698, i_8_704, i_8_705, i_8_782, i_8_814, i_8_832, i_8_838, i_8_877, i_8_912, i_8_958, i_8_995, i_8_1128, i_8_1174, i_8_1192, i_8_1201, i_8_1228, i_8_1263, i_8_1284, i_8_1299, i_8_1305, i_8_1306, i_8_1307, i_8_1315, i_8_1354, i_8_1390, i_8_1467, i_8_1473, i_8_1497, i_8_1524, i_8_1525, i_8_1534, i_8_1570, i_8_1624, i_8_1635, i_8_1648, i_8_1678, i_8_1686, i_8_1696, i_8_1714, i_8_1746, i_8_1747, i_8_1752, i_8_1776, i_8_1791, i_8_1795, i_8_1801, i_8_1806, i_8_1818, i_8_1822, i_8_1848, i_8_1849, i_8_1876, i_8_1906, i_8_1918, i_8_1976, i_8_2014, i_8_2046, i_8_2047, i_8_2064, i_8_2065, i_8_2066, i_8_2091, i_8_2092, i_8_2119, i_8_2122, i_8_2155, i_8_2215, i_8_2216, i_8_2256, i_8_2291, o_8_10);
	kernel_8_11 k_8_11(i_8_64, i_8_79, i_8_111, i_8_141, i_8_197, i_8_231, i_8_262, i_8_265, i_8_311, i_8_326, i_8_329, i_8_364, i_8_367, i_8_379, i_8_392, i_8_401, i_8_419, i_8_424, i_8_439, i_8_475, i_8_486, i_8_499, i_8_509, i_8_525, i_8_528, i_8_529, i_8_557, i_8_571, i_8_616, i_8_625, i_8_631, i_8_635, i_8_656, i_8_659, i_8_661, i_8_673, i_8_700, i_8_703, i_8_718, i_8_724, i_8_725, i_8_734, i_8_754, i_8_771, i_8_824, i_8_835, i_8_837, i_8_838, i_8_840, i_8_841, i_8_968, i_8_1012, i_8_1110, i_8_1191, i_8_1229, i_8_1231, i_8_1246, i_8_1267, i_8_1301, i_8_1354, i_8_1355, i_8_1399, i_8_1411, i_8_1462, i_8_1471, i_8_1547, i_8_1571, i_8_1625, i_8_1647, i_8_1653, i_8_1655, i_8_1679, i_8_1696, i_8_1699, i_8_1747, i_8_1748, i_8_1750, i_8_1754, i_8_1769, i_8_1773, i_8_1795, i_8_1798, i_8_1819, i_8_1840, i_8_1849, i_8_1858, i_8_1912, i_8_1913, i_8_1952, i_8_1981, i_8_2011, i_8_2012, i_8_2048, i_8_2074, i_8_2095, i_8_2119, i_8_2136, i_8_2191, i_8_2257, i_8_2298, o_8_11);
	kernel_8_12 k_8_12(i_8_13, i_8_92, i_8_94, i_8_121, i_8_138, i_8_139, i_8_183, i_8_192, i_8_193, i_8_209, i_8_221, i_8_278, i_8_284, i_8_318, i_8_325, i_8_326, i_8_350, i_8_363, i_8_390, i_8_471, i_8_472, i_8_473, i_8_478, i_8_480, i_8_481, i_8_505, i_8_523, i_8_554, i_8_569, i_8_632, i_8_656, i_8_694, i_8_696, i_8_697, i_8_712, i_8_731, i_8_749, i_8_750, i_8_863, i_8_877, i_8_883, i_8_893, i_8_959, i_8_962, i_8_964, i_8_967, i_8_991, i_8_995, i_8_1027, i_8_1094, i_8_1120, i_8_1144, i_8_1201, i_8_1202, i_8_1234, i_8_1286, i_8_1309, i_8_1315, i_8_1316, i_8_1328, i_8_1342, i_8_1372, i_8_1382, i_8_1413, i_8_1432, i_8_1434, i_8_1442, i_8_1621, i_8_1625, i_8_1651, i_8_1665, i_8_1666, i_8_1696, i_8_1699, i_8_1705, i_8_1712, i_8_1749, i_8_1751, i_8_1805, i_8_1818, i_8_1857, i_8_1874, i_8_1981, i_8_1982, i_8_2008, i_8_2009, i_8_2025, i_8_2053, i_8_2083, i_8_2084, i_8_2090, i_8_2122, i_8_2123, i_8_2143, i_8_2170, i_8_2189, i_8_2227, i_8_2284, i_8_2285, i_8_2299, o_8_12);
	kernel_8_13 k_8_13(i_8_4, i_8_28, i_8_33, i_8_47, i_8_58, i_8_59, i_8_71, i_8_166, i_8_170, i_8_190, i_8_227, i_8_256, i_8_257, i_8_281, i_8_293, i_8_320, i_8_326, i_8_328, i_8_364, i_8_379, i_8_380, i_8_421, i_8_424, i_8_444, i_8_453, i_8_593, i_8_603, i_8_660, i_8_693, i_8_703, i_8_704, i_8_705, i_8_706, i_8_708, i_8_778, i_8_784, i_8_787, i_8_826, i_8_832, i_8_833, i_8_838, i_8_842, i_8_844, i_8_873, i_8_877, i_8_886, i_8_890, i_8_928, i_8_932, i_8_977, i_8_1083, i_8_1108, i_8_1115, i_8_1174, i_8_1180, i_8_1183, i_8_1234, i_8_1236, i_8_1271, i_8_1282, i_8_1286, i_8_1327, i_8_1352, i_8_1360, i_8_1435, i_8_1442, i_8_1472, i_8_1474, i_8_1498, i_8_1533, i_8_1597, i_8_1603, i_8_1607, i_8_1634, i_8_1673, i_8_1706, i_8_1746, i_8_1748, i_8_1764, i_8_1769, i_8_1789, i_8_1807, i_8_1813, i_8_1824, i_8_1881, i_8_1907, i_8_1965, i_8_1967, i_8_1984, i_8_1987, i_8_1989, i_8_2038, i_8_2052, i_8_2056, i_8_2060, i_8_2143, i_8_2150, i_8_2224, i_8_2263, i_8_2264, o_8_13);
	kernel_8_14 k_8_14(i_8_25, i_8_41, i_8_170, i_8_174, i_8_178, i_8_228, i_8_230, i_8_231, i_8_233, i_8_248, i_8_273, i_8_277, i_8_278, i_8_355, i_8_356, i_8_359, i_8_363, i_8_364, i_8_385, i_8_391, i_8_476, i_8_484, i_8_499, i_8_516, i_8_518, i_8_592, i_8_597, i_8_607, i_8_608, i_8_611, i_8_626, i_8_634, i_8_772, i_8_799, i_8_825, i_8_830, i_8_841, i_8_879, i_8_889, i_8_925, i_8_935, i_8_955, i_8_958, i_8_959, i_8_994, i_8_996, i_8_1039, i_8_1075, i_8_1076, i_8_1087, i_8_1178, i_8_1192, i_8_1228, i_8_1232, i_8_1241, i_8_1258, i_8_1273, i_8_1274, i_8_1277, i_8_1285, i_8_1385, i_8_1387, i_8_1391, i_8_1408, i_8_1412, i_8_1497, i_8_1525, i_8_1528, i_8_1546, i_8_1552, i_8_1645, i_8_1647, i_8_1650, i_8_1659, i_8_1680, i_8_1681, i_8_1726, i_8_1767, i_8_1768, i_8_1771, i_8_1800, i_8_1807, i_8_1849, i_8_1866, i_8_1870, i_8_1906, i_8_1919, i_8_1940, i_8_1967, i_8_1996, i_8_2040, i_8_2041, i_8_2066, i_8_2075, i_8_2146, i_8_2150, i_8_2159, i_8_2212, i_8_2219, i_8_2249, o_8_14);
	kernel_8_15 k_8_15(i_8_5, i_8_19, i_8_76, i_8_83, i_8_112, i_8_140, i_8_148, i_8_150, i_8_169, i_8_173, i_8_192, i_8_193, i_8_226, i_8_239, i_8_245, i_8_274, i_8_275, i_8_325, i_8_335, i_8_341, i_8_353, i_8_361, i_8_364, i_8_365, i_8_442, i_8_515, i_8_581, i_8_587, i_8_596, i_8_652, i_8_667, i_8_668, i_8_680, i_8_703, i_8_704, i_8_707, i_8_730, i_8_733, i_8_751, i_8_756, i_8_830, i_8_910, i_8_911, i_8_968, i_8_1111, i_8_1129, i_8_1171, i_8_1297, i_8_1355, i_8_1483, i_8_1495, i_8_1521, i_8_1522, i_8_1531, i_8_1549, i_8_1594, i_8_1634, i_8_1651, i_8_1652, i_8_1682, i_8_1694, i_8_1705, i_8_1748, i_8_1765, i_8_1766, i_8_1774, i_8_1777, i_8_1805, i_8_1818, i_8_1819, i_8_1821, i_8_1822, i_8_1826, i_8_1857, i_8_1864, i_8_1874, i_8_1881, i_8_1892, i_8_1946, i_8_1967, i_8_1991, i_8_1994, i_8_1995, i_8_1996, i_8_2008, i_8_2009, i_8_2011, i_8_2062, i_8_2063, i_8_2074, i_8_2146, i_8_2147, i_8_2215, i_8_2227, i_8_2255, i_8_2256, i_8_2258, i_8_2269, i_8_2294, i_8_2300, o_8_15);
	kernel_8_16 k_8_16(i_8_4, i_8_8, i_8_19, i_8_41, i_8_76, i_8_138, i_8_176, i_8_184, i_8_248, i_8_275, i_8_277, i_8_356, i_8_364, i_8_365, i_8_382, i_8_422, i_8_463, i_8_464, i_8_493, i_8_497, i_8_500, i_8_517, i_8_518, i_8_527, i_8_555, i_8_571, i_8_593, i_8_596, i_8_598, i_8_608, i_8_658, i_8_661, i_8_705, i_8_732, i_8_733, i_8_734, i_8_754, i_8_832, i_8_833, i_8_840, i_8_894, i_8_914, i_8_959, i_8_965, i_8_990, i_8_994, i_8_1073, i_8_1084, i_8_1175, i_8_1264, i_8_1298, i_8_1308, i_8_1331, i_8_1354, i_8_1358, i_8_1391, i_8_1466, i_8_1481, i_8_1484, i_8_1498, i_8_1499, i_8_1517, i_8_1534, i_8_1535, i_8_1597, i_8_1598, i_8_1654, i_8_1655, i_8_1660, i_8_1666, i_8_1678, i_8_1679, i_8_1695, i_8_1698, i_8_1777, i_8_1795, i_8_1812, i_8_1824, i_8_1826, i_8_1843, i_8_1849, i_8_1867, i_8_1876, i_8_1885, i_8_1894, i_8_1918, i_8_1951, i_8_1967, i_8_1995, i_8_2011, i_8_2039, i_8_2048, i_8_2172, i_8_2215, i_8_2227, i_8_2230, i_8_2234, i_8_2245, i_8_2284, i_8_2294, o_8_16);
	kernel_8_17 k_8_17(i_8_27, i_8_28, i_8_34, i_8_51, i_8_82, i_8_85, i_8_93, i_8_156, i_8_199, i_8_233, i_8_243, i_8_252, i_8_255, i_8_288, i_8_297, i_8_324, i_8_342, i_8_345, i_8_371, i_8_378, i_8_435, i_8_436, i_8_450, i_8_471, i_8_530, i_8_551, i_8_562, i_8_565, i_8_585, i_8_586, i_8_615, i_8_621, i_8_624, i_8_633, i_8_637, i_8_657, i_8_665, i_8_666, i_8_669, i_8_694, i_8_700, i_8_715, i_8_810, i_8_972, i_8_973, i_8_975, i_8_990, i_8_1011, i_8_1188, i_8_1215, i_8_1216, i_8_1219, i_8_1224, i_8_1233, i_8_1247, i_8_1263, i_8_1278, i_8_1279, i_8_1284, i_8_1326, i_8_1345, i_8_1375, i_8_1434, i_8_1443, i_8_1503, i_8_1539, i_8_1584, i_8_1585, i_8_1587, i_8_1593, i_8_1594, i_8_1633, i_8_1665, i_8_1680, i_8_1701, i_8_1710, i_8_1751, i_8_1758, i_8_1799, i_8_1831, i_8_1845, i_8_1848, i_8_1854, i_8_1890, i_8_1899, i_8_1963, i_8_2043, i_8_2046, i_8_2092, i_8_2106, i_8_2110, i_8_2124, i_8_2126, i_8_2178, i_8_2179, i_8_2187, i_8_2259, i_8_2260, i_8_2269, i_8_2277, o_8_17);
	kernel_8_18 k_8_18(i_8_12, i_8_13, i_8_14, i_8_31, i_8_41, i_8_67, i_8_88, i_8_114, i_8_122, i_8_136, i_8_150, i_8_175, i_8_178, i_8_193, i_8_202, i_8_211, i_8_274, i_8_276, i_8_277, i_8_292, i_8_354, i_8_362, i_8_401, i_8_410, i_8_421, i_8_427, i_8_507, i_8_534, i_8_535, i_8_544, i_8_553, i_8_571, i_8_574, i_8_616, i_8_633, i_8_634, i_8_653, i_8_660, i_8_662, i_8_676, i_8_680, i_8_697, i_8_700, i_8_703, i_8_707, i_8_729, i_8_732, i_8_804, i_8_826, i_8_864, i_8_866, i_8_867, i_8_868, i_8_973, i_8_976, i_8_1031, i_8_1084, i_8_1102, i_8_1108, i_8_1153, i_8_1155, i_8_1174, i_8_1243, i_8_1245, i_8_1278, i_8_1299, i_8_1301, i_8_1314, i_8_1315, i_8_1336, i_8_1372, i_8_1387, i_8_1398, i_8_1405, i_8_1423, i_8_1440, i_8_1477, i_8_1525, i_8_1549, i_8_1576, i_8_1606, i_8_1642, i_8_1665, i_8_1683, i_8_1689, i_8_1791, i_8_1805, i_8_1822, i_8_1826, i_8_1884, i_8_1938, i_8_1995, i_8_2119, i_8_2147, i_8_2148, i_8_2173, i_8_2181, i_8_2188, i_8_2244, i_8_2272, o_8_18);
	kernel_8_19 k_8_19(i_8_52, i_8_57, i_8_58, i_8_59, i_8_87, i_8_88, i_8_142, i_8_143, i_8_166, i_8_168, i_8_169, i_8_229, i_8_230, i_8_233, i_8_257, i_8_258, i_8_260, i_8_328, i_8_329, i_8_369, i_8_370, i_8_377, i_8_379, i_8_421, i_8_437, i_8_483, i_8_485, i_8_502, i_8_508, i_8_522, i_8_529, i_8_530, i_8_552, i_8_553, i_8_556, i_8_557, i_8_596, i_8_633, i_8_634, i_8_635, i_8_689, i_8_691, i_8_692, i_8_735, i_8_736, i_8_752, i_8_762, i_8_768, i_8_815, i_8_850, i_8_868, i_8_993, i_8_994, i_8_1050, i_8_1051, i_8_1052, i_8_1057, i_8_1073, i_8_1110, i_8_1112, i_8_1119, i_8_1120, i_8_1188, i_8_1189, i_8_1292, i_8_1305, i_8_1306, i_8_1307, i_8_1315, i_8_1317, i_8_1327, i_8_1407, i_8_1437, i_8_1438, i_8_1506, i_8_1516, i_8_1560, i_8_1574, i_8_1631, i_8_1632, i_8_1633, i_8_1680, i_8_1684, i_8_1723, i_8_1749, i_8_1750, i_8_1754, i_8_1823, i_8_1861, i_8_1919, i_8_1958, i_8_1959, i_8_1960, i_8_1992, i_8_2003, i_8_2005, i_8_2032, i_8_2057, i_8_2093, i_8_2096, o_8_19);
	kernel_8_20 k_8_20(i_8_16, i_8_37, i_8_79, i_8_80, i_8_147, i_8_158, i_8_197, i_8_226, i_8_229, i_8_230, i_8_233, i_8_310, i_8_364, i_8_404, i_8_418, i_8_430, i_8_456, i_8_471, i_8_579, i_8_583, i_8_598, i_8_611, i_8_638, i_8_645, i_8_652, i_8_656, i_8_662, i_8_670, i_8_700, i_8_702, i_8_780, i_8_825, i_8_843, i_8_861, i_8_862, i_8_881, i_8_899, i_8_967, i_8_1015, i_8_1043, i_8_1089, i_8_1112, i_8_1129, i_8_1131, i_8_1187, i_8_1228, i_8_1263, i_8_1285, i_8_1299, i_8_1303, i_8_1310, i_8_1339, i_8_1340, i_8_1353, i_8_1384, i_8_1403, i_8_1426, i_8_1439, i_8_1474, i_8_1488, i_8_1489, i_8_1520, i_8_1545, i_8_1551, i_8_1552, i_8_1624, i_8_1628, i_8_1642, i_8_1653, i_8_1681, i_8_1706, i_8_1752, i_8_1771, i_8_1789, i_8_1806, i_8_1807, i_8_1812, i_8_1831, i_8_1843, i_8_1844, i_8_1854, i_8_1870, i_8_1875, i_8_1921, i_8_1943, i_8_1974, i_8_1978, i_8_1987, i_8_1993, i_8_2041, i_8_2091, i_8_2092, i_8_2110, i_8_2141, i_8_2215, i_8_2229, i_8_2238, i_8_2253, i_8_2265, i_8_2301, o_8_20);
	kernel_8_21 k_8_21(i_8_28, i_8_29, i_8_60, i_8_138, i_8_139, i_8_158, i_8_159, i_8_166, i_8_193, i_8_229, i_8_230, i_8_232, i_8_363, i_8_364, i_8_365, i_8_366, i_8_368, i_8_381, i_8_484, i_8_510, i_8_528, i_8_657, i_8_661, i_8_687, i_8_688, i_8_690, i_8_691, i_8_692, i_8_695, i_8_707, i_8_709, i_8_762, i_8_763, i_8_764, i_8_822, i_8_827, i_8_844, i_8_845, i_8_868, i_8_994, i_8_1013, i_8_1026, i_8_1030, i_8_1033, i_8_1034, i_8_1051, i_8_1056, i_8_1059, i_8_1090, i_8_1115, i_8_1159, i_8_1160, i_8_1184, i_8_1255, i_8_1265, i_8_1296, i_8_1305, i_8_1306, i_8_1308, i_8_1310, i_8_1325, i_8_1344, i_8_1404, i_8_1556, i_8_1572, i_8_1634, i_8_1672, i_8_1674, i_8_1723, i_8_1741, i_8_1742, i_8_1743, i_8_1744, i_8_1745, i_8_1801, i_8_1805, i_8_1806, i_8_1808, i_8_1821, i_8_1822, i_8_1824, i_8_1825, i_8_1832, i_8_1834, i_8_1854, i_8_1918, i_8_2076, i_8_2119, i_8_2215, i_8_2216, i_8_2217, i_8_2224, i_8_2226, i_8_2233, i_8_2234, i_8_2271, i_8_2274, i_8_2275, i_8_2289, i_8_2290, o_8_21);
	kernel_8_22 k_8_22(i_8_9, i_8_49, i_8_118, i_8_126, i_8_300, i_8_360, i_8_361, i_8_382, i_8_390, i_8_391, i_8_399, i_8_400, i_8_417, i_8_426, i_8_453, i_8_504, i_8_505, i_8_558, i_8_559, i_8_561, i_8_568, i_8_639, i_8_640, i_8_660, i_8_661, i_8_676, i_8_679, i_8_696, i_8_697, i_8_702, i_8_766, i_8_783, i_8_784, i_8_847, i_8_891, i_8_892, i_8_969, i_8_999, i_8_1036, i_8_1045, i_8_1054, i_8_1102, i_8_1111, i_8_1130, i_8_1152, i_8_1179, i_8_1198, i_8_1234, i_8_1236, i_8_1263, i_8_1281, i_8_1295, i_8_1299, i_8_1339, i_8_1359, i_8_1360, i_8_1362, i_8_1363, i_8_1381, i_8_1399, i_8_1422, i_8_1423, i_8_1432, i_8_1440, i_8_1448, i_8_1450, i_8_1484, i_8_1486, i_8_1512, i_8_1513, i_8_1515, i_8_1521, i_8_1524, i_8_1551, i_8_1569, i_8_1639, i_8_1651, i_8_1656, i_8_1677, i_8_1678, i_8_1686, i_8_1746, i_8_1750, i_8_1767, i_8_1822, i_8_1839, i_8_1840, i_8_1845, i_8_1881, i_8_1974, i_8_1981, i_8_1992, i_8_2145, i_8_2147, i_8_2152, i_8_2190, i_8_2191, i_8_2224, i_8_2244, i_8_2245, o_8_22);
	kernel_8_23 k_8_23(i_8_22, i_8_37, i_8_40, i_8_52, i_8_75, i_8_82, i_8_85, i_8_94, i_8_123, i_8_126, i_8_165, i_8_175, i_8_214, i_8_255, i_8_288, i_8_346, i_8_355, i_8_364, i_8_373, i_8_382, i_8_383, i_8_400, i_8_427, i_8_453, i_8_484, i_8_500, i_8_551, i_8_555, i_8_586, i_8_587, i_8_589, i_8_595, i_8_598, i_8_606, i_8_607, i_8_662, i_8_679, i_8_696, i_8_702, i_8_709, i_8_786, i_8_799, i_8_868, i_8_880, i_8_955, i_8_975, i_8_1020, i_8_1069, i_8_1071, i_8_1072, i_8_1090, i_8_1119, i_8_1123, i_8_1221, i_8_1227, i_8_1267, i_8_1272, i_8_1291, i_8_1298, i_8_1305, i_8_1308, i_8_1324, i_8_1327, i_8_1365, i_8_1470, i_8_1542, i_8_1606, i_8_1614, i_8_1626, i_8_1686, i_8_1749, i_8_1794, i_8_1821, i_8_1822, i_8_1824, i_8_1825, i_8_1830, i_8_1849, i_8_1855, i_8_1935, i_8_1938, i_8_1944, i_8_1993, i_8_1996, i_8_2002, i_8_2075, i_8_2103, i_8_2137, i_8_2142, i_8_2182, i_8_2212, i_8_2226, i_8_2227, i_8_2232, i_8_2235, i_8_2236, i_8_2245, i_8_2263, i_8_2280, i_8_2281, o_8_23);
	kernel_8_24 k_8_24(i_8_34, i_8_69, i_8_78, i_8_79, i_8_115, i_8_133, i_8_169, i_8_250, i_8_312, i_8_337, i_8_380, i_8_384, i_8_475, i_8_500, i_8_501, i_8_511, i_8_519, i_8_525, i_8_528, i_8_539, i_8_553, i_8_555, i_8_574, i_8_583, i_8_600, i_8_628, i_8_637, i_8_664, i_8_673, i_8_733, i_8_750, i_8_834, i_8_843, i_8_916, i_8_1033, i_8_1087, i_8_1111, i_8_1177, i_8_1183, i_8_1245, i_8_1258, i_8_1273, i_8_1285, i_8_1291, i_8_1302, i_8_1303, i_8_1304, i_8_1365, i_8_1401, i_8_1407, i_8_1416, i_8_1438, i_8_1470, i_8_1489, i_8_1492, i_8_1501, i_8_1528, i_8_1536, i_8_1537, i_8_1544, i_8_1552, i_8_1608, i_8_1614, i_8_1653, i_8_1663, i_8_1672, i_8_1696, i_8_1702, i_8_1752, i_8_1762, i_8_1781, i_8_1794, i_8_1798, i_8_1816, i_8_1821, i_8_1851, i_8_1879, i_8_1884, i_8_1887, i_8_1898, i_8_1915, i_8_1951, i_8_1968, i_8_1970, i_8_2013, i_8_2041, i_8_2050, i_8_2064, i_8_2122, i_8_2153, i_8_2176, i_8_2186, i_8_2216, i_8_2218, i_8_2219, i_8_2228, i_8_2229, i_8_2247, i_8_2248, i_8_2257, o_8_24);
	kernel_8_25 k_8_25(i_8_20, i_8_27, i_8_44, i_8_48, i_8_54, i_8_87, i_8_108, i_8_115, i_8_220, i_8_304, i_8_325, i_8_345, i_8_355, i_8_365, i_8_489, i_8_491, i_8_553, i_8_571, i_8_606, i_8_607, i_8_613, i_8_617, i_8_643, i_8_651, i_8_655, i_8_675, i_8_694, i_8_698, i_8_701, i_8_782, i_8_791, i_8_802, i_8_876, i_8_882, i_8_993, i_8_1038, i_8_1040, i_8_1054, i_8_1071, i_8_1074, i_8_1093, i_8_1094, i_8_1098, i_8_1102, i_8_1125, i_8_1131, i_8_1137, i_8_1142, i_8_1146, i_8_1147, i_8_1164, i_8_1224, i_8_1237, i_8_1254, i_8_1313, i_8_1318, i_8_1322, i_8_1330, i_8_1351, i_8_1362, i_8_1422, i_8_1482, i_8_1526, i_8_1549, i_8_1600, i_8_1607, i_8_1621, i_8_1654, i_8_1677, i_8_1704, i_8_1737, i_8_1738, i_8_1739, i_8_1741, i_8_1770, i_8_1790, i_8_1804, i_8_1806, i_8_1808, i_8_1809, i_8_1821, i_8_1822, i_8_1949, i_8_1958, i_8_1966, i_8_1983, i_8_1995, i_8_2055, i_8_2058, i_8_2076, i_8_2097, i_8_2101, i_8_2104, i_8_2124, i_8_2154, i_8_2163, i_8_2173, i_8_2190, i_8_2191, i_8_2233, o_8_25);
	kernel_8_26 k_8_26(i_8_19, i_8_32, i_8_33, i_8_138, i_8_153, i_8_157, i_8_184, i_8_193, i_8_373, i_8_379, i_8_387, i_8_388, i_8_436, i_8_441, i_8_442, i_8_479, i_8_495, i_8_496, i_8_507, i_8_508, i_8_525, i_8_526, i_8_536, i_8_551, i_8_554, i_8_586, i_8_604, i_8_613, i_8_660, i_8_662, i_8_666, i_8_678, i_8_760, i_8_761, i_8_769, i_8_819, i_8_822, i_8_823, i_8_824, i_8_864, i_8_865, i_8_918, i_8_922, i_8_981, i_8_982, i_8_983, i_8_1008, i_8_1030, i_8_1108, i_8_1112, i_8_1129, i_8_1130, i_8_1153, i_8_1233, i_8_1236, i_8_1242, i_8_1243, i_8_1245, i_8_1246, i_8_1252, i_8_1263, i_8_1264, i_8_1278, i_8_1279, i_8_1323, i_8_1341, i_8_1400, i_8_1435, i_8_1503, i_8_1506, i_8_1513, i_8_1530, i_8_1531, i_8_1550, i_8_1561, i_8_1576, i_8_1594, i_8_1611, i_8_1614, i_8_1647, i_8_1667, i_8_1755, i_8_1756, i_8_1777, i_8_1785, i_8_1800, i_8_1837, i_8_1848, i_8_1890, i_8_1943, i_8_1999, i_8_2037, i_8_2043, i_8_2106, i_8_2107, i_8_2178, i_8_2223, i_8_2236, i_8_2237, i_8_2245, o_8_26);
	kernel_8_27 k_8_27(i_8_4, i_8_5, i_8_25, i_8_35, i_8_44, i_8_77, i_8_87, i_8_148, i_8_211, i_8_230, i_8_244, i_8_247, i_8_248, i_8_274, i_8_275, i_8_323, i_8_363, i_8_368, i_8_385, i_8_421, i_8_422, i_8_431, i_8_527, i_8_528, i_8_530, i_8_565, i_8_571, i_8_572, i_8_575, i_8_582, i_8_583, i_8_586, i_8_644, i_8_652, i_8_655, i_8_670, i_8_671, i_8_681, i_8_682, i_8_696, i_8_703, i_8_706, i_8_733, i_8_734, i_8_760, i_8_781, i_8_844, i_8_850, i_8_859, i_8_889, i_8_943, i_8_956, i_8_991, i_8_992, i_8_1105, i_8_1111, i_8_1129, i_8_1132, i_8_1172, i_8_1321, i_8_1329, i_8_1330, i_8_1354, i_8_1355, i_8_1358, i_8_1382, i_8_1399, i_8_1400, i_8_1465, i_8_1468, i_8_1480, i_8_1481, i_8_1518, i_8_1531, i_8_1535, i_8_1541, i_8_1598, i_8_1699, i_8_1703, i_8_1705, i_8_1753, i_8_1754, i_8_1772, i_8_1795, i_8_1796, i_8_1804, i_8_1807, i_8_1813, i_8_1843, i_8_1928, i_8_1960, i_8_2042, i_8_2065, i_8_2066, i_8_2194, i_8_2216, i_8_2244, i_8_2254, i_8_2255, i_8_2256, o_8_27);
	kernel_8_28 k_8_28(i_8_1, i_8_19, i_8_20, i_8_85, i_8_118, i_8_136, i_8_143, i_8_144, i_8_190, i_8_202, i_8_352, i_8_381, i_8_382, i_8_391, i_8_414, i_8_442, i_8_469, i_8_514, i_8_522, i_8_523, i_8_524, i_8_525, i_8_567, i_8_577, i_8_595, i_8_596, i_8_607, i_8_610, i_8_631, i_8_634, i_8_637, i_8_658, i_8_667, i_8_702, i_8_703, i_8_712, i_8_748, i_8_751, i_8_829, i_8_838, i_8_844, i_8_859, i_8_881, i_8_910, i_8_929, i_8_955, i_8_964, i_8_967, i_8_968, i_8_997, i_8_1179, i_8_1198, i_8_1234, i_8_1252, i_8_1282, i_8_1354, i_8_1387, i_8_1396, i_8_1467, i_8_1468, i_8_1486, i_8_1495, i_8_1507, i_8_1531, i_8_1533, i_8_1536, i_8_1594, i_8_1629, i_8_1639, i_8_1647, i_8_1657, i_8_1702, i_8_1703, i_8_1747, i_8_1757, i_8_1774, i_8_1775, i_8_1791, i_8_1792, i_8_1801, i_8_1802, i_8_1818, i_8_1819, i_8_1822, i_8_1846, i_8_1864, i_8_1873, i_8_1900, i_8_1910, i_8_1963, i_8_2008, i_8_2044, i_8_2062, i_8_2089, i_8_2116, i_8_2133, i_8_2134, i_8_2173, i_8_2227, i_8_2284, o_8_28);
	kernel_8_29 k_8_29(i_8_58, i_8_77, i_8_80, i_8_104, i_8_107, i_8_116, i_8_140, i_8_182, i_8_185, i_8_188, i_8_197, i_8_247, i_8_366, i_8_367, i_8_389, i_8_391, i_8_394, i_8_400, i_8_401, i_8_428, i_8_431, i_8_451, i_8_453, i_8_490, i_8_575, i_8_584, i_8_594, i_8_604, i_8_608, i_8_610, i_8_638, i_8_814, i_8_853, i_8_856, i_8_860, i_8_879, i_8_962, i_8_1012, i_8_1013, i_8_1015, i_8_1016, i_8_1029, i_8_1040, i_8_1105, i_8_1106, i_8_1129, i_8_1130, i_8_1142, i_8_1157, i_8_1160, i_8_1228, i_8_1322, i_8_1328, i_8_1331, i_8_1350, i_8_1407, i_8_1465, i_8_1493, i_8_1507, i_8_1510, i_8_1519, i_8_1538, i_8_1550, i_8_1553, i_8_1658, i_8_1688, i_8_1690, i_8_1697, i_8_1784, i_8_1817, i_8_1822, i_8_1838, i_8_1840, i_8_1844, i_8_1850, i_8_1860, i_8_1882, i_8_1885, i_8_1894, i_8_1895, i_8_1946, i_8_1966, i_8_2017, i_8_2038, i_8_2041, i_8_2072, i_8_2116, i_8_2119, i_8_2120, i_8_2126, i_8_2150, i_8_2154, i_8_2172, i_8_2177, i_8_2231, i_8_2263, i_8_2264, i_8_2266, i_8_2273, i_8_2276, o_8_29);
	kernel_8_30 k_8_30(i_8_32, i_8_49, i_8_50, i_8_87, i_8_95, i_8_116, i_8_143, i_8_167, i_8_176, i_8_220, i_8_227, i_8_304, i_8_347, i_8_361, i_8_378, i_8_383, i_8_385, i_8_416, i_8_425, i_8_490, i_8_525, i_8_527, i_8_550, i_8_553, i_8_581, i_8_614, i_8_653, i_8_656, i_8_671, i_8_677, i_8_687, i_8_689, i_8_695, i_8_749, i_8_794, i_8_796, i_8_797, i_8_806, i_8_830, i_8_838, i_8_932, i_8_956, i_8_991, i_8_994, i_8_1058, i_8_1101, i_8_1126, i_8_1127, i_8_1130, i_8_1175, i_8_1235, i_8_1256, i_8_1271, i_8_1277, i_8_1283, i_8_1285, i_8_1323, i_8_1340, i_8_1358, i_8_1382, i_8_1442, i_8_1453, i_8_1454, i_8_1471, i_8_1481, i_8_1489, i_8_1490, i_8_1536, i_8_1544, i_8_1552, i_8_1625, i_8_1639, i_8_1677, i_8_1697, i_8_1721, i_8_1741, i_8_1774, i_8_1775, i_8_1801, i_8_1823, i_8_1856, i_8_1868, i_8_1886, i_8_1889, i_8_1892, i_8_1943, i_8_1966, i_8_1991, i_8_2039, i_8_2050, i_8_2143, i_8_2146, i_8_2171, i_8_2192, i_8_2210, i_8_2215, i_8_2237, i_8_2261, i_8_2282, i_8_2291, o_8_30);
	kernel_8_31 k_8_31(i_8_10, i_8_37, i_8_73, i_8_114, i_8_169, i_8_172, i_8_363, i_8_364, i_8_373, i_8_442, i_8_454, i_8_471, i_8_486, i_8_487, i_8_493, i_8_507, i_8_522, i_8_526, i_8_535, i_8_555, i_8_580, i_8_616, i_8_656, i_8_664, i_8_669, i_8_684, i_8_694, i_8_696, i_8_697, i_8_704, i_8_766, i_8_837, i_8_840, i_8_841, i_8_847, i_8_913, i_8_948, i_8_949, i_8_955, i_8_956, i_8_1102, i_8_1103, i_8_1108, i_8_1110, i_8_1127, i_8_1129, i_8_1130, i_8_1224, i_8_1225, i_8_1227, i_8_1228, i_8_1281, i_8_1286, i_8_1305, i_8_1352, i_8_1357, i_8_1369, i_8_1390, i_8_1399, i_8_1456, i_8_1480, i_8_1489, i_8_1497, i_8_1516, i_8_1533, i_8_1549, i_8_1558, i_8_1673, i_8_1685, i_8_1704, i_8_1784, i_8_1794, i_8_1803, i_8_1805, i_8_1822, i_8_1824, i_8_1864, i_8_1885, i_8_1912, i_8_1917, i_8_1939, i_8_1957, i_8_1990, i_8_1993, i_8_2006, i_8_2021, i_8_2048, i_8_2133, i_8_2134, i_8_2143, i_8_2146, i_8_2147, i_8_2148, i_8_2165, i_8_2215, i_8_2232, i_8_2236, i_8_2242, i_8_2296, i_8_2299, o_8_31);
	kernel_8_32 k_8_32(i_8_22, i_8_39, i_8_196, i_8_232, i_8_300, i_8_303, i_8_304, i_8_330, i_8_360, i_8_364, i_8_365, i_8_367, i_8_368, i_8_420, i_8_421, i_8_448, i_8_457, i_8_510, i_8_511, i_8_520, i_8_525, i_8_528, i_8_605, i_8_606, i_8_658, i_8_660, i_8_700, i_8_751, i_8_762, i_8_781, i_8_782, i_8_795, i_8_823, i_8_835, i_8_842, i_8_843, i_8_852, i_8_996, i_8_997, i_8_1028, i_8_1050, i_8_1158, i_8_1159, i_8_1192, i_8_1249, i_8_1274, i_8_1282, i_8_1305, i_8_1308, i_8_1330, i_8_1382, i_8_1389, i_8_1391, i_8_1393, i_8_1432, i_8_1437, i_8_1438, i_8_1439, i_8_1545, i_8_1546, i_8_1554, i_8_1596, i_8_1635, i_8_1643, i_8_1679, i_8_1699, i_8_1700, i_8_1708, i_8_1764, i_8_1784, i_8_1818, i_8_1820, i_8_1840, i_8_1858, i_8_1875, i_8_1876, i_8_1879, i_8_1880, i_8_1887, i_8_2013, i_8_2014, i_8_2075, i_8_2077, i_8_2091, i_8_2092, i_8_2093, i_8_2095, i_8_2096, i_8_2122, i_8_2147, i_8_2154, i_8_2214, i_8_2215, i_8_2216, i_8_2218, i_8_2235, i_8_2236, i_8_2239, i_8_2244, i_8_2293, o_8_32);
	kernel_8_33 k_8_33(i_8_30, i_8_33, i_8_34, i_8_48, i_8_49, i_8_53, i_8_76, i_8_164, i_8_174, i_8_193, i_8_227, i_8_258, i_8_305, i_8_345, i_8_348, i_8_366, i_8_385, i_8_453, i_8_479, i_8_510, i_8_552, i_8_585, i_8_634, i_8_651, i_8_652, i_8_653, i_8_718, i_8_719, i_8_770, i_8_773, i_8_778, i_8_796, i_8_797, i_8_805, i_8_862, i_8_885, i_8_890, i_8_921, i_8_923, i_8_930, i_8_935, i_8_992, i_8_1091, i_8_1102, i_8_1159, i_8_1170, i_8_1258, i_8_1259, i_8_1263, i_8_1265, i_8_1274, i_8_1301, i_8_1302, i_8_1305, i_8_1330, i_8_1331, i_8_1355, i_8_1399, i_8_1408, i_8_1470, i_8_1471, i_8_1473, i_8_1489, i_8_1490, i_8_1549, i_8_1562, i_8_1587, i_8_1678, i_8_1700, i_8_1733, i_8_1753, i_8_1773, i_8_1774, i_8_1776, i_8_1778, i_8_1788, i_8_1805, i_8_1864, i_8_1939, i_8_1993, i_8_2017, i_8_2031, i_8_2048, i_8_2111, i_8_2172, i_8_2174, i_8_2175, i_8_2176, i_8_2177, i_8_2194, i_8_2200, i_8_2206, i_8_2244, i_8_2245, i_8_2246, i_8_2249, i_8_2264, i_8_2276, i_8_2291, i_8_2292, o_8_33);
	kernel_8_34 k_8_34(i_8_40, i_8_51, i_8_57, i_8_79, i_8_143, i_8_174, i_8_220, i_8_225, i_8_252, i_8_265, i_8_364, i_8_365, i_8_367, i_8_369, i_8_453, i_8_492, i_8_499, i_8_589, i_8_590, i_8_591, i_8_595, i_8_597, i_8_598, i_8_634, i_8_635, i_8_651, i_8_659, i_8_660, i_8_675, i_8_679, i_8_680, i_8_693, i_8_705, i_8_706, i_8_729, i_8_779, i_8_819, i_8_820, i_8_855, i_8_866, i_8_882, i_8_885, i_8_937, i_8_968, i_8_969, i_8_971, i_8_1035, i_8_1039, i_8_1137, i_8_1147, i_8_1164, i_8_1165, i_8_1182, i_8_1220, i_8_1227, i_8_1260, i_8_1262, i_8_1297, i_8_1318, i_8_1369, i_8_1389, i_8_1479, i_8_1507, i_8_1524, i_8_1545, i_8_1546, i_8_1547, i_8_1564, i_8_1607, i_8_1610, i_8_1614, i_8_1675, i_8_1677, i_8_1703, i_8_1714, i_8_1762, i_8_1807, i_8_1850, i_8_1885, i_8_1927, i_8_1981, i_8_1984, i_8_2004, i_8_2052, i_8_2056, i_8_2091, i_8_2100, i_8_2101, i_8_2133, i_8_2135, i_8_2155, i_8_2163, i_8_2173, i_8_2176, i_8_2214, i_8_2224, i_8_2227, i_8_2241, i_8_2244, i_8_2262, o_8_34);
	kernel_8_35 k_8_35(i_8_25, i_8_28, i_8_31, i_8_83, i_8_203, i_8_299, i_8_352, i_8_371, i_8_418, i_8_440, i_8_443, i_8_469, i_8_478, i_8_481, i_8_482, i_8_484, i_8_496, i_8_587, i_8_667, i_8_671, i_8_793, i_8_815, i_8_918, i_8_919, i_8_1003, i_8_1008, i_8_1013, i_8_1027, i_8_1108, i_8_1109, i_8_1125, i_8_1126, i_8_1127, i_8_1135, i_8_1139, i_8_1157, i_8_1217, i_8_1234, i_8_1256, i_8_1325, i_8_1346, i_8_1348, i_8_1435, i_8_1437, i_8_1468, i_8_1506, i_8_1521, i_8_1548, i_8_1556, i_8_1582, i_8_1603, i_8_1612, i_8_1640, i_8_1668, i_8_1669, i_8_1674, i_8_1675, i_8_1703, i_8_1704, i_8_1705, i_8_1714, i_8_1715, i_8_1717, i_8_1720, i_8_1746, i_8_1748, i_8_1749, i_8_1750, i_8_1751, i_8_1752, i_8_1776, i_8_1785, i_8_1791, i_8_1801, i_8_1808, i_8_1809, i_8_1812, i_8_1813, i_8_1838, i_8_1849, i_8_1859, i_8_1882, i_8_1918, i_8_1947, i_8_1951, i_8_1964, i_8_1986, i_8_1996, i_8_2000, i_8_2044, i_8_2107, i_8_2111, i_8_2125, i_8_2128, i_8_2143, i_8_2180, i_8_2188, i_8_2189, i_8_2245, i_8_2289, o_8_35);
	kernel_8_36 k_8_36(i_8_31, i_8_33, i_8_35, i_8_43, i_8_49, i_8_54, i_8_57, i_8_73, i_8_93, i_8_94, i_8_101, i_8_183, i_8_228, i_8_230, i_8_238, i_8_300, i_8_334, i_8_345, i_8_360, i_8_368, i_8_380, i_8_417, i_8_472, i_8_489, i_8_503, i_8_508, i_8_527, i_8_528, i_8_571, i_8_599, i_8_617, i_8_634, i_8_670, i_8_686, i_8_689, i_8_710, i_8_733, i_8_760, i_8_764, i_8_775, i_8_780, i_8_781, i_8_805, i_8_809, i_8_826, i_8_841, i_8_859, i_8_877, i_8_883, i_8_904, i_8_939, i_8_940, i_8_941, i_8_990, i_8_1075, i_8_1144, i_8_1160, i_8_1169, i_8_1228, i_8_1229, i_8_1236, i_8_1294, i_8_1300, i_8_1312, i_8_1331, i_8_1399, i_8_1467, i_8_1492, i_8_1506, i_8_1539, i_8_1585, i_8_1625, i_8_1632, i_8_1655, i_8_1678, i_8_1681, i_8_1682, i_8_1696, i_8_1697, i_8_1723, i_8_1741, i_8_1750, i_8_1753, i_8_1784, i_8_1813, i_8_1835, i_8_1903, i_8_1986, i_8_2058, i_8_2059, i_8_2098, i_8_2119, i_8_2137, i_8_2171, i_8_2173, i_8_2176, i_8_2191, i_8_2276, i_8_2296, i_8_2299, o_8_36);
	kernel_8_37 k_8_37(i_8_42, i_8_70, i_8_78, i_8_87, i_8_94, i_8_102, i_8_283, i_8_286, i_8_303, i_8_310, i_8_322, i_8_365, i_8_394, i_8_400, i_8_403, i_8_420, i_8_421, i_8_444, i_8_511, i_8_529, i_8_552, i_8_571, i_8_573, i_8_633, i_8_637, i_8_642, i_8_643, i_8_652, i_8_662, i_8_706, i_8_760, i_8_814, i_8_825, i_8_861, i_8_871, i_8_895, i_8_970, i_8_992, i_8_1071, i_8_1086, i_8_1104, i_8_1131, i_8_1156, i_8_1236, i_8_1262, i_8_1291, i_8_1318, i_8_1330, i_8_1338, i_8_1345, i_8_1365, i_8_1366, i_8_1393, i_8_1402, i_8_1407, i_8_1411, i_8_1425, i_8_1438, i_8_1464, i_8_1465, i_8_1471, i_8_1473, i_8_1479, i_8_1482, i_8_1483, i_8_1486, i_8_1515, i_8_1516, i_8_1518, i_8_1524, i_8_1527, i_8_1528, i_8_1536, i_8_1554, i_8_1635, i_8_1660, i_8_1669, i_8_1671, i_8_1676, i_8_1681, i_8_1690, i_8_1696, i_8_1704, i_8_1705, i_8_1707, i_8_1708, i_8_1779, i_8_1794, i_8_1823, i_8_1839, i_8_1840, i_8_1843, i_8_1914, i_8_1938, i_8_1977, i_8_2146, i_8_2149, i_8_2206, i_8_2223, i_8_2294, o_8_37);
	kernel_8_38 k_8_38(i_8_25, i_8_170, i_8_247, i_8_293, i_8_296, i_8_319, i_8_329, i_8_334, i_8_341, i_8_361, i_8_363, i_8_366, i_8_367, i_8_383, i_8_454, i_8_480, i_8_535, i_8_553, i_8_562, i_8_580, i_8_592, i_8_604, i_8_608, i_8_621, i_8_628, i_8_631, i_8_634, i_8_662, i_8_693, i_8_696, i_8_698, i_8_703, i_8_705, i_8_714, i_8_718, i_8_719, i_8_783, i_8_809, i_8_840, i_8_843, i_8_871, i_8_880, i_8_954, i_8_957, i_8_966, i_8_969, i_8_1015, i_8_1051, i_8_1075, i_8_1076, i_8_1115, i_8_1226, i_8_1228, i_8_1231, i_8_1240, i_8_1273, i_8_1285, i_8_1286, i_8_1321, i_8_1330, i_8_1372, i_8_1445, i_8_1456, i_8_1470, i_8_1518, i_8_1542, i_8_1552, i_8_1553, i_8_1560, i_8_1561, i_8_1563, i_8_1571, i_8_1591, i_8_1624, i_8_1632, i_8_1668, i_8_1680, i_8_1704, i_8_1708, i_8_1733, i_8_1808, i_8_1809, i_8_1825, i_8_1835, i_8_1854, i_8_1862, i_8_1870, i_8_1885, i_8_1912, i_8_1966, i_8_1992, i_8_1996, i_8_2132, i_8_2134, i_8_2147, i_8_2217, i_8_2244, i_8_2245, i_8_2248, i_8_2281, o_8_38);
	kernel_8_39 k_8_39(i_8_63, i_8_64, i_8_117, i_8_138, i_8_147, i_8_192, i_8_237, i_8_262, i_8_273, i_8_319, i_8_352, i_8_360, i_8_364, i_8_365, i_8_369, i_8_417, i_8_450, i_8_451, i_8_457, i_8_460, i_8_489, i_8_531, i_8_549, i_8_585, i_8_603, i_8_606, i_8_607, i_8_651, i_8_661, i_8_675, i_8_694, i_8_700, i_8_703, i_8_704, i_8_729, i_8_751, i_8_810, i_8_814, i_8_828, i_8_829, i_8_849, i_8_876, i_8_981, i_8_1063, i_8_1080, i_8_1101, i_8_1102, i_8_1114, i_8_1138, i_8_1162, i_8_1200, i_8_1260, i_8_1278, i_8_1296, i_8_1306, i_8_1324, i_8_1355, i_8_1377, i_8_1378, i_8_1386, i_8_1395, i_8_1396, i_8_1408, i_8_1452, i_8_1468, i_8_1486, i_8_1488, i_8_1503, i_8_1540, i_8_1548, i_8_1562, i_8_1624, i_8_1647, i_8_1650, i_8_1668, i_8_1674, i_8_1681, i_8_1702, i_8_1758, i_8_1764, i_8_1792, i_8_1801, i_8_1821, i_8_1824, i_8_1828, i_8_1857, i_8_1873, i_8_1885, i_8_1908, i_8_1944, i_8_1962, i_8_1972, i_8_1995, i_8_2007, i_8_2008, i_8_2089, i_8_2134, i_8_2148, i_8_2241, i_8_2295, o_8_39);
	kernel_8_40 k_8_40(i_8_8, i_8_39, i_8_66, i_8_89, i_8_168, i_8_169, i_8_175, i_8_183, i_8_187, i_8_191, i_8_324, i_8_425, i_8_450, i_8_456, i_8_489, i_8_524, i_8_528, i_8_529, i_8_530, i_8_552, i_8_553, i_8_589, i_8_601, i_8_615, i_8_636, i_8_685, i_8_690, i_8_691, i_8_699, i_8_700, i_8_705, i_8_707, i_8_737, i_8_763, i_8_798, i_8_837, i_8_838, i_8_843, i_8_881, i_8_892, i_8_957, i_8_966, i_8_995, i_8_1029, i_8_1030, i_8_1044, i_8_1076, i_8_1078, i_8_1096, i_8_1114, i_8_1205, i_8_1213, i_8_1230, i_8_1239, i_8_1273, i_8_1276, i_8_1284, i_8_1285, i_8_1340, i_8_1353, i_8_1362, i_8_1426, i_8_1446, i_8_1447, i_8_1452, i_8_1471, i_8_1490, i_8_1570, i_8_1605, i_8_1681, i_8_1689, i_8_1723, i_8_1751, i_8_1762, i_8_1773, i_8_1776, i_8_1777, i_8_1815, i_8_1852, i_8_1862, i_8_1903, i_8_1904, i_8_1941, i_8_1996, i_8_2005, i_8_2074, i_8_2113, i_8_2140, i_8_2145, i_8_2150, i_8_2174, i_8_2175, i_8_2185, i_8_2212, i_8_2226, i_8_2233, i_8_2234, i_8_2265, i_8_2267, i_8_2289, o_8_40);
	kernel_8_41 k_8_41(i_8_13, i_8_23, i_8_35, i_8_85, i_8_118, i_8_121, i_8_122, i_8_139, i_8_148, i_8_189, i_8_328, i_8_348, i_8_362, i_8_450, i_8_483, i_8_484, i_8_499, i_8_538, i_8_552, i_8_556, i_8_589, i_8_607, i_8_636, i_8_662, i_8_679, i_8_682, i_8_686, i_8_694, i_8_697, i_8_699, i_8_733, i_8_755, i_8_781, i_8_785, i_8_797, i_8_823, i_8_839, i_8_843, i_8_958, i_8_968, i_8_973, i_8_977, i_8_1027, i_8_1030, i_8_1036, i_8_1057, i_8_1087, i_8_1111, i_8_1113, i_8_1127, i_8_1133, i_8_1157, i_8_1183, i_8_1230, i_8_1251, i_8_1255, i_8_1300, i_8_1337, i_8_1355, i_8_1552, i_8_1564, i_8_1588, i_8_1610, i_8_1612, i_8_1622, i_8_1624, i_8_1627, i_8_1628, i_8_1639, i_8_1669, i_8_1684, i_8_1694, i_8_1748, i_8_1750, i_8_1759, i_8_1768, i_8_1769, i_8_1777, i_8_1778, i_8_1791, i_8_1802, i_8_1805, i_8_1816, i_8_1858, i_8_1926, i_8_1939, i_8_1996, i_8_2011, i_8_2134, i_8_2138, i_8_2149, i_8_2150, i_8_2173, i_8_2229, i_8_2230, i_8_2232, i_8_2245, i_8_2246, i_8_2247, i_8_2263, o_8_41);
	kernel_8_42 k_8_42(i_8_0, i_8_66, i_8_72, i_8_106, i_8_135, i_8_144, i_8_199, i_8_220, i_8_240, i_8_244, i_8_309, i_8_397, i_8_399, i_8_400, i_8_418, i_8_427, i_8_498, i_8_507, i_8_513, i_8_553, i_8_554, i_8_570, i_8_588, i_8_601, i_8_603, i_8_614, i_8_617, i_8_651, i_8_655, i_8_706, i_8_714, i_8_730, i_8_747, i_8_831, i_8_837, i_8_840, i_8_891, i_8_958, i_8_973, i_8_1108, i_8_1152, i_8_1170, i_8_1197, i_8_1200, i_8_1224, i_8_1236, i_8_1266, i_8_1294, i_8_1350, i_8_1353, i_8_1359, i_8_1363, i_8_1390, i_8_1399, i_8_1422, i_8_1431, i_8_1440, i_8_1461, i_8_1462, i_8_1467, i_8_1476, i_8_1494, i_8_1556, i_8_1632, i_8_1635, i_8_1692, i_8_1693, i_8_1722, i_8_1748, i_8_1749, i_8_1750, i_8_1751, i_8_1764, i_8_1782, i_8_1792, i_8_1805, i_8_1815, i_8_1822, i_8_1836, i_8_1840, i_8_1866, i_8_1881, i_8_1885, i_8_1917, i_8_1926, i_8_1947, i_8_1950, i_8_1974, i_8_1980, i_8_2007, i_8_2043, i_8_2044, i_8_2062, i_8_2116, i_8_2142, i_8_2143, i_8_2145, i_8_2146, i_8_2149, i_8_2248, o_8_42);
	kernel_8_43 k_8_43(i_8_3, i_8_30, i_8_31, i_8_34, i_8_42, i_8_94, i_8_99, i_8_100, i_8_117, i_8_120, i_8_126, i_8_220, i_8_274, i_8_279, i_8_288, i_8_309, i_8_315, i_8_345, i_8_348, i_8_356, i_8_378, i_8_381, i_8_384, i_8_402, i_8_427, i_8_432, i_8_433, i_8_435, i_8_442, i_8_517, i_8_527, i_8_530, i_8_547, i_8_660, i_8_665, i_8_723, i_8_774, i_8_814, i_8_819, i_8_841, i_8_861, i_8_894, i_8_913, i_8_967, i_8_972, i_8_981, i_8_999, i_8_1102, i_8_1200, i_8_1206, i_8_1251, i_8_1263, i_8_1266, i_8_1284, i_8_1372, i_8_1410, i_8_1434, i_8_1445, i_8_1453, i_8_1456, i_8_1491, i_8_1510, i_8_1539, i_8_1555, i_8_1565, i_8_1566, i_8_1584, i_8_1609, i_8_1611, i_8_1623, i_8_1627, i_8_1684, i_8_1755, i_8_1759, i_8_1776, i_8_1866, i_8_1873, i_8_1899, i_8_1902, i_8_1905, i_8_1936, i_8_1942, i_8_1975, i_8_1976, i_8_2001, i_8_2025, i_8_2062, i_8_2065, i_8_2080, i_8_2083, i_8_2115, i_8_2142, i_8_2143, i_8_2149, i_8_2169, i_8_2173, i_8_2187, i_8_2205, i_8_2209, i_8_2257, o_8_43);
	kernel_8_44 k_8_44(i_8_11, i_8_23, i_8_28, i_8_95, i_8_97, i_8_157, i_8_158, i_8_202, i_8_203, i_8_209, i_8_223, i_8_244, i_8_245, i_8_248, i_8_266, i_8_326, i_8_348, i_8_355, i_8_364, i_8_380, i_8_437, i_8_452, i_8_483, i_8_484, i_8_498, i_8_508, i_8_526, i_8_536, i_8_551, i_8_554, i_8_556, i_8_557, i_8_587, i_8_626, i_8_628, i_8_657, i_8_779, i_8_793, i_8_827, i_8_841, i_8_851, i_8_877, i_8_878, i_8_896, i_8_992, i_8_996, i_8_1012, i_8_1061, i_8_1066, i_8_1067, i_8_1084, i_8_1112, i_8_1115, i_8_1133, i_8_1148, i_8_1175, i_8_1246, i_8_1247, i_8_1261, i_8_1328, i_8_1346, i_8_1350, i_8_1417, i_8_1418, i_8_1451, i_8_1523, i_8_1525, i_8_1526, i_8_1550, i_8_1579, i_8_1613, i_8_1654, i_8_1667, i_8_1679, i_8_1681, i_8_1682, i_8_1729, i_8_1730, i_8_1733, i_8_1739, i_8_1747, i_8_1750, i_8_1753, i_8_1777, i_8_1778, i_8_1802, i_8_1808, i_8_1856, i_8_1867, i_8_1903, i_8_1904, i_8_1959, i_8_1990, i_8_1996, i_8_2011, i_8_2012, i_8_2077, i_8_2078, i_8_2153, i_8_2288, o_8_44);
	kernel_8_45 k_8_45(i_8_41, i_8_44, i_8_77, i_8_112, i_8_114, i_8_115, i_8_116, i_8_141, i_8_182, i_8_317, i_8_319, i_8_320, i_8_322, i_8_381, i_8_382, i_8_392, i_8_398, i_8_489, i_8_537, i_8_547, i_8_553, i_8_556, i_8_568, i_8_571, i_8_580, i_8_589, i_8_598, i_8_612, i_8_634, i_8_640, i_8_652, i_8_655, i_8_657, i_8_670, i_8_680, i_8_716, i_8_732, i_8_859, i_8_860, i_8_895, i_8_966, i_8_970, i_8_975, i_8_1102, i_8_1111, i_8_1187, i_8_1192, i_8_1193, i_8_1201, i_8_1225, i_8_1228, i_8_1243, i_8_1296, i_8_1316, i_8_1326, i_8_1327, i_8_1363, i_8_1384, i_8_1407, i_8_1423, i_8_1427, i_8_1435, i_8_1462, i_8_1463, i_8_1467, i_8_1469, i_8_1477, i_8_1481, i_8_1516, i_8_1546, i_8_1573, i_8_1625, i_8_1630, i_8_1633, i_8_1694, i_8_1697, i_8_1750, i_8_1765, i_8_1768, i_8_1771, i_8_1776, i_8_1783, i_8_1840, i_8_1885, i_8_1894, i_8_1906, i_8_1912, i_8_1918, i_8_1949, i_8_1957, i_8_1972, i_8_1975, i_8_1979, i_8_1984, i_8_2041, i_8_2069, i_8_2095, i_8_2135, i_8_2192, i_8_2226, o_8_45);
	kernel_8_46 k_8_46(i_8_77, i_8_107, i_8_250, i_8_259, i_8_284, i_8_296, i_8_322, i_8_323, i_8_368, i_8_431, i_8_457, i_8_490, i_8_494, i_8_530, i_8_587, i_8_593, i_8_599, i_8_628, i_8_643, i_8_653, i_8_661, i_8_673, i_8_681, i_8_691, i_8_697, i_8_698, i_8_707, i_8_719, i_8_728, i_8_736, i_8_763, i_8_775, i_8_809, i_8_815, i_8_817, i_8_838, i_8_842, i_8_845, i_8_881, i_8_970, i_8_971, i_8_1031, i_8_1033, i_8_1078, i_8_1205, i_8_1227, i_8_1228, i_8_1232, i_8_1238, i_8_1239, i_8_1240, i_8_1265, i_8_1268, i_8_1321, i_8_1350, i_8_1358, i_8_1363, i_8_1391, i_8_1407, i_8_1408, i_8_1432, i_8_1436, i_8_1475, i_8_1492, i_8_1519, i_8_1520, i_8_1527, i_8_1528, i_8_1570, i_8_1574, i_8_1591, i_8_1592, i_8_1625, i_8_1642, i_8_1706, i_8_1744, i_8_1754, i_8_1768, i_8_1771, i_8_1813, i_8_1822, i_8_1823, i_8_1826, i_8_1858, i_8_1859, i_8_1880, i_8_1885, i_8_1889, i_8_1982, i_8_1994, i_8_2029, i_8_2032, i_8_2077, i_8_2132, i_8_2149, i_8_2156, i_8_2195, i_8_2224, i_8_2285, i_8_2290, o_8_46);
	kernel_8_47 k_8_47(i_8_7, i_8_24, i_8_70, i_8_79, i_8_88, i_8_129, i_8_151, i_8_195, i_8_212, i_8_214, i_8_247, i_8_250, i_8_277, i_8_313, i_8_358, i_8_376, i_8_396, i_8_450, i_8_467, i_8_503, i_8_528, i_8_529, i_8_570, i_8_597, i_8_602, i_8_609, i_8_615, i_8_636, i_8_654, i_8_655, i_8_672, i_8_681, i_8_695, i_8_700, i_8_708, i_8_709, i_8_735, i_8_751, i_8_754, i_8_762, i_8_772, i_8_835, i_8_862, i_8_1060, i_8_1061, i_8_1069, i_8_1137, i_8_1155, i_8_1177, i_8_1227, i_8_1257, i_8_1266, i_8_1267, i_8_1300, i_8_1303, i_8_1357, i_8_1384, i_8_1393, i_8_1410, i_8_1455, i_8_1496, i_8_1498, i_8_1501, i_8_1534, i_8_1551, i_8_1552, i_8_1599, i_8_1645, i_8_1648, i_8_1653, i_8_1654, i_8_1662, i_8_1690, i_8_1735, i_8_1750, i_8_1813, i_8_1851, i_8_1852, i_8_1870, i_8_1914, i_8_1915, i_8_1920, i_8_1921, i_8_1968, i_8_1969, i_8_1996, i_8_2013, i_8_2014, i_8_2068, i_8_2095, i_8_2112, i_8_2122, i_8_2172, i_8_2175, i_8_2184, i_8_2185, i_8_2217, i_8_2218, i_8_2272, i_8_2292, o_8_47);
	kernel_8_48 k_8_48(i_8_22, i_8_82, i_8_104, i_8_263, i_8_292, i_8_302, i_8_303, i_8_346, i_8_347, i_8_377, i_8_418, i_8_463, i_8_464, i_8_476, i_8_482, i_8_500, i_8_503, i_8_547, i_8_554, i_8_556, i_8_557, i_8_589, i_8_593, i_8_597, i_8_599, i_8_625, i_8_674, i_8_716, i_8_796, i_8_827, i_8_892, i_8_895, i_8_1030, i_8_1114, i_8_1115, i_8_1121, i_8_1129, i_8_1130, i_8_1258, i_8_1271, i_8_1274, i_8_1283, i_8_1286, i_8_1307, i_8_1314, i_8_1323, i_8_1347, i_8_1350, i_8_1432, i_8_1453, i_8_1454, i_8_1470, i_8_1471, i_8_1472, i_8_1535, i_8_1587, i_8_1597, i_8_1604, i_8_1681, i_8_1706, i_8_1711, i_8_1714, i_8_1749, i_8_1763, i_8_1787, i_8_1790, i_8_1802, i_8_1807, i_8_1841, i_8_1854, i_8_1855, i_8_1867, i_8_1871, i_8_1895, i_8_1918, i_8_1919, i_8_1927, i_8_1948, i_8_1970, i_8_2033, i_8_2050, i_8_2051, i_8_2110, i_8_2111, i_8_2129, i_8_2134, i_8_2140, i_8_2183, i_8_2191, i_8_2192, i_8_2214, i_8_2215, i_8_2216, i_8_2230, i_8_2234, i_8_2247, i_8_2261, i_8_2273, i_8_2276, i_8_2290, o_8_48);
	kernel_8_49 k_8_49(i_8_22, i_8_39, i_8_53, i_8_126, i_8_147, i_8_318, i_8_319, i_8_320, i_8_321, i_8_322, i_8_323, i_8_336, i_8_342, i_8_396, i_8_397, i_8_424, i_8_425, i_8_427, i_8_439, i_8_547, i_8_552, i_8_561, i_8_571, i_8_580, i_8_588, i_8_589, i_8_596, i_8_603, i_8_604, i_8_610, i_8_611, i_8_658, i_8_676, i_8_695, i_8_750, i_8_766, i_8_777, i_8_841, i_8_865, i_8_875, i_8_894, i_8_969, i_8_976, i_8_1022, i_8_1100, i_8_1102, i_8_1103, i_8_1110, i_8_1180, i_8_1236, i_8_1237, i_8_1243, i_8_1264, i_8_1286, i_8_1327, i_8_1357, i_8_1362, i_8_1363, i_8_1380, i_8_1381, i_8_1399, i_8_1431, i_8_1432, i_8_1461, i_8_1463, i_8_1477, i_8_1514, i_8_1526, i_8_1536, i_8_1573, i_8_1605, i_8_1606, i_8_1626, i_8_1632, i_8_1681, i_8_1707, i_8_1735, i_8_1749, i_8_1750, i_8_1760, i_8_1766, i_8_1767, i_8_1781, i_8_1866, i_8_1884, i_8_1929, i_8_1930, i_8_1937, i_8_1957, i_8_1974, i_8_1975, i_8_1996, i_8_2091, i_8_2119, i_8_2143, i_8_2191, i_8_2244, i_8_2245, i_8_2246, i_8_2271, o_8_49);
	kernel_8_50 k_8_50(i_8_14, i_8_18, i_8_85, i_8_93, i_8_117, i_8_151, i_8_192, i_8_193, i_8_258, i_8_259, i_8_273, i_8_325, i_8_360, i_8_363, i_8_364, i_8_423, i_8_426, i_8_427, i_8_447, i_8_468, i_8_526, i_8_529, i_8_554, i_8_567, i_8_568, i_8_615, i_8_622, i_8_630, i_8_652, i_8_684, i_8_694, i_8_699, i_8_707, i_8_832, i_8_837, i_8_865, i_8_873, i_8_874, i_8_876, i_8_882, i_8_981, i_8_1023, i_8_1030, i_8_1036, i_8_1051, i_8_1089, i_8_1092, i_8_1102, i_8_1137, i_8_1138, i_8_1147, i_8_1237, i_8_1267, i_8_1314, i_8_1332, i_8_1349, i_8_1407, i_8_1455, i_8_1486, i_8_1597, i_8_1602, i_8_1605, i_8_1620, i_8_1638, i_8_1650, i_8_1696, i_8_1702, i_8_1765, i_8_1768, i_8_1774, i_8_1804, i_8_1807, i_8_1810, i_8_1818, i_8_1821, i_8_1857, i_8_1881, i_8_1882, i_8_1884, i_8_1893, i_8_1929, i_8_1938, i_8_2007, i_8_2044, i_8_2055, i_8_2066, i_8_2070, i_8_2079, i_8_2092, i_8_2097, i_8_2114, i_8_2124, i_8_2144, i_8_2146, i_8_2147, i_8_2152, i_8_2170, i_8_2241, i_8_2246, i_8_2294, o_8_50);
	kernel_8_51 k_8_51(i_8_26, i_8_69, i_8_88, i_8_176, i_8_193, i_8_197, i_8_204, i_8_205, i_8_206, i_8_214, i_8_215, i_8_278, i_8_345, i_8_358, i_8_359, i_8_364, i_8_367, i_8_377, i_8_379, i_8_383, i_8_384, i_8_398, i_8_449, i_8_458, i_8_475, i_8_500, i_8_503, i_8_520, i_8_521, i_8_530, i_8_575, i_8_592, i_8_593, i_8_619, i_8_634, i_8_673, i_8_674, i_8_692, i_8_719, i_8_772, i_8_773, i_8_818, i_8_826, i_8_833, i_8_881, i_8_890, i_8_959, i_8_995, i_8_1035, i_8_1043, i_8_1079, i_8_1087, i_8_1196, i_8_1232, i_8_1261, i_8_1264, i_8_1285, i_8_1294, i_8_1300, i_8_1304, i_8_1312, i_8_1353, i_8_1410, i_8_1439, i_8_1473, i_8_1501, i_8_1504, i_8_1544, i_8_1565, i_8_1646, i_8_1672, i_8_1673, i_8_1691, i_8_1699, i_8_1700, i_8_1717, i_8_1718, i_8_1722, i_8_1735, i_8_1771, i_8_1772, i_8_1789, i_8_1807, i_8_1816, i_8_1844, i_8_1853, i_8_1880, i_8_1886, i_8_1887, i_8_1948, i_8_2014, i_8_2015, i_8_2074, i_8_2152, i_8_2186, i_8_2194, i_8_2195, i_8_2218, i_8_2249, i_8_2267, o_8_51);
	kernel_8_52 k_8_52(i_8_3, i_8_17, i_8_20, i_8_21, i_8_29, i_8_31, i_8_37, i_8_53, i_8_87, i_8_88, i_8_104, i_8_263, i_8_290, i_8_307, i_8_316, i_8_335, i_8_348, i_8_363, i_8_379, i_8_380, i_8_402, i_8_417, i_8_483, i_8_489, i_8_528, i_8_529, i_8_586, i_8_587, i_8_605, i_8_621, i_8_634, i_8_649, i_8_660, i_8_675, i_8_693, i_8_703, i_8_721, i_8_730, i_8_791, i_8_824, i_8_841, i_8_843, i_8_874, i_8_888, i_8_918, i_8_923, i_8_950, i_8_968, i_8_974, i_8_1078, i_8_1120, i_8_1180, i_8_1222, i_8_1264, i_8_1276, i_8_1284, i_8_1290, i_8_1324, i_8_1334, i_8_1440, i_8_1469, i_8_1474, i_8_1504, i_8_1585, i_8_1680, i_8_1682, i_8_1698, i_8_1743, i_8_1745, i_8_1748, i_8_1752, i_8_1760, i_8_1764, i_8_1768, i_8_1773, i_8_1796, i_8_1817, i_8_1820, i_8_1854, i_8_1861, i_8_1901, i_8_1904, i_8_1981, i_8_1993, i_8_1999, i_8_2026, i_8_2071, i_8_2105, i_8_2117, i_8_2130, i_8_2139, i_8_2140, i_8_2141, i_8_2143, i_8_2187, i_8_2188, i_8_2234, i_8_2243, i_8_2287, i_8_2301, o_8_52);
	kernel_8_53 k_8_53(i_8_32, i_8_37, i_8_41, i_8_43, i_8_51, i_8_57, i_8_64, i_8_67, i_8_120, i_8_160, i_8_172, i_8_205, i_8_228, i_8_229, i_8_230, i_8_325, i_8_326, i_8_329, i_8_334, i_8_352, i_8_392, i_8_400, i_8_401, i_8_417, i_8_462, i_8_502, i_8_552, i_8_555, i_8_556, i_8_557, i_8_697, i_8_698, i_8_699, i_8_700, i_8_701, i_8_748, i_8_838, i_8_839, i_8_850, i_8_883, i_8_885, i_8_886, i_8_889, i_8_995, i_8_1012, i_8_1128, i_8_1129, i_8_1131, i_8_1133, i_8_1156, i_8_1158, i_8_1202, i_8_1203, i_8_1205, i_8_1236, i_8_1322, i_8_1328, i_8_1331, i_8_1381, i_8_1427, i_8_1489, i_8_1551, i_8_1552, i_8_1555, i_8_1682, i_8_1705, i_8_1709, i_8_1726, i_8_1732, i_8_1749, i_8_1751, i_8_1753, i_8_1797, i_8_1806, i_8_1807, i_8_1841, i_8_1912, i_8_1913, i_8_1914, i_8_1915, i_8_1916, i_8_1936, i_8_1939, i_8_1982, i_8_1983, i_8_1985, i_8_1992, i_8_1999, i_8_2017, i_8_2055, i_8_2057, i_8_2058, i_8_2059, i_8_2144, i_8_2146, i_8_2147, i_8_2154, i_8_2159, i_8_2177, i_8_2272, o_8_53);
	kernel_8_54 k_8_54(i_8_31, i_8_32, i_8_52, i_8_55, i_8_79, i_8_97, i_8_104, i_8_208, i_8_212, i_8_258, i_8_262, i_8_283, i_8_292, i_8_301, i_8_363, i_8_382, i_8_384, i_8_427, i_8_454, i_8_456, i_8_492, i_8_624, i_8_625, i_8_628, i_8_636, i_8_669, i_8_670, i_8_679, i_8_682, i_8_696, i_8_698, i_8_701, i_8_719, i_8_727, i_8_733, i_8_738, i_8_781, i_8_784, i_8_786, i_8_792, i_8_800, i_8_827, i_8_840, i_8_853, i_8_880, i_8_915, i_8_958, i_8_1029, i_8_1059, i_8_1108, i_8_1114, i_8_1138, i_8_1229, i_8_1249, i_8_1282, i_8_1285, i_8_1335, i_8_1354, i_8_1355, i_8_1381, i_8_1438, i_8_1444, i_8_1454, i_8_1542, i_8_1543, i_8_1565, i_8_1588, i_8_1591, i_8_1606, i_8_1683, i_8_1684, i_8_1700, i_8_1706, i_8_1732, i_8_1736, i_8_1762, i_8_1771, i_8_1794, i_8_1805, i_8_1808, i_8_1822, i_8_1823, i_8_1825, i_8_1858, i_8_1860, i_8_1867, i_8_1885, i_8_1912, i_8_1966, i_8_1983, i_8_1997, i_8_2147, i_8_2190, i_8_2193, i_8_2200, i_8_2215, i_8_2229, i_8_2247, i_8_2263, i_8_2284, o_8_54);
	kernel_8_55 k_8_55(i_8_6, i_8_23, i_8_30, i_8_41, i_8_65, i_8_68, i_8_85, i_8_86, i_8_137, i_8_142, i_8_145, i_8_175, i_8_176, i_8_199, i_8_205, i_8_247, i_8_282, i_8_335, i_8_355, i_8_356, i_8_364, i_8_368, i_8_437, i_8_440, i_8_444, i_8_445, i_8_497, i_8_517, i_8_527, i_8_550, i_8_588, i_8_597, i_8_615, i_8_661, i_8_682, i_8_699, i_8_707, i_8_710, i_8_713, i_8_715, i_8_727, i_8_728, i_8_770, i_8_914, i_8_958, i_8_971, i_8_992, i_8_1084, i_8_1127, i_8_1134, i_8_1229, i_8_1236, i_8_1267, i_8_1282, i_8_1305, i_8_1351, i_8_1363, i_8_1391, i_8_1407, i_8_1425, i_8_1437, i_8_1438, i_8_1447, i_8_1484, i_8_1487, i_8_1490, i_8_1525, i_8_1549, i_8_1598, i_8_1629, i_8_1642, i_8_1646, i_8_1654, i_8_1687, i_8_1700, i_8_1706, i_8_1745, i_8_1779, i_8_1781, i_8_1794, i_8_1813, i_8_1819, i_8_1820, i_8_1823, i_8_1837, i_8_1850, i_8_1873, i_8_1884, i_8_1916, i_8_1980, i_8_2004, i_8_2044, i_8_2046, i_8_2066, i_8_2090, i_8_2098, i_8_2147, i_8_2183, i_8_2238, i_8_2289, o_8_55);
	kernel_8_56 k_8_56(i_8_20, i_8_65, i_8_76, i_8_77, i_8_94, i_8_112, i_8_245, i_8_353, i_8_388, i_8_389, i_8_443, i_8_461, i_8_481, i_8_486, i_8_497, i_8_515, i_8_524, i_8_529, i_8_549, i_8_550, i_8_595, i_8_605, i_8_631, i_8_632, i_8_633, i_8_658, i_8_716, i_8_812, i_8_830, i_8_841, i_8_843, i_8_873, i_8_875, i_8_877, i_8_883, i_8_926, i_8_965, i_8_967, i_8_1040, i_8_1073, i_8_1127, i_8_1143, i_8_1144, i_8_1153, i_8_1171, i_8_1198, i_8_1199, i_8_1269, i_8_1283, i_8_1298, i_8_1315, i_8_1351, i_8_1382, i_8_1396, i_8_1397, i_8_1424, i_8_1431, i_8_1433, i_8_1451, i_8_1468, i_8_1495, i_8_1513, i_8_1514, i_8_1523, i_8_1532, i_8_1621, i_8_1649, i_8_1657, i_8_1658, i_8_1681, i_8_1702, i_8_1703, i_8_1730, i_8_1747, i_8_1773, i_8_1791, i_8_1792, i_8_1793, i_8_1823, i_8_1824, i_8_1864, i_8_1882, i_8_1909, i_8_1910, i_8_1936, i_8_1981, i_8_2044, i_8_2052, i_8_2053, i_8_2099, i_8_2117, i_8_2134, i_8_2143, i_8_2169, i_8_2171, i_8_2224, i_8_2234, i_8_2243, i_8_2254, i_8_2283, o_8_56);
	kernel_8_57 k_8_57(i_8_156, i_8_258, i_8_348, i_8_372, i_8_380, i_8_441, i_8_458, i_8_462, i_8_463, i_8_468, i_8_474, i_8_475, i_8_480, i_8_503, i_8_552, i_8_585, i_8_607, i_8_639, i_8_642, i_8_669, i_8_719, i_8_720, i_8_778, i_8_793, i_8_811, i_8_831, i_8_837, i_8_838, i_8_841, i_8_870, i_8_950, i_8_973, i_8_1011, i_8_1014, i_8_1066, i_8_1071, i_8_1072, i_8_1074, i_8_1075, i_8_1083, i_8_1084, i_8_1129, i_8_1134, i_8_1218, i_8_1225, i_8_1236, i_8_1237, i_8_1249, i_8_1252, i_8_1254, i_8_1255, i_8_1261, i_8_1263, i_8_1272, i_8_1283, i_8_1285, i_8_1288, i_8_1305, i_8_1306, i_8_1307, i_8_1378, i_8_1419, i_8_1452, i_8_1467, i_8_1519, i_8_1535, i_8_1542, i_8_1584, i_8_1587, i_8_1593, i_8_1596, i_8_1605, i_8_1606, i_8_1611, i_8_1624, i_8_1641, i_8_1659, i_8_1680, i_8_1704, i_8_1705, i_8_1718, i_8_1720, i_8_1747, i_8_1764, i_8_1767, i_8_1783, i_8_1803, i_8_1804, i_8_1805, i_8_1815, i_8_1828, i_8_1864, i_8_1981, i_8_2037, i_8_2124, i_8_2143, i_8_2146, i_8_2154, i_8_2272, i_8_2274, o_8_57);
	kernel_8_58 k_8_58(i_8_54, i_8_86, i_8_89, i_8_97, i_8_111, i_8_254, i_8_257, i_8_259, i_8_266, i_8_279, i_8_328, i_8_334, i_8_344, i_8_390, i_8_449, i_8_454, i_8_455, i_8_489, i_8_500, i_8_511, i_8_525, i_8_527, i_8_530, i_8_628, i_8_662, i_8_666, i_8_670, i_8_674, i_8_683, i_8_716, i_8_725, i_8_742, i_8_759, i_8_789, i_8_791, i_8_796, i_8_815, i_8_834, i_8_842, i_8_856, i_8_874, i_8_881, i_8_952, i_8_953, i_8_1030, i_8_1114, i_8_1120, i_8_1132, i_8_1138, i_8_1159, i_8_1160, i_8_1200, i_8_1236, i_8_1237, i_8_1238, i_8_1262, i_8_1283, i_8_1294, i_8_1321, i_8_1347, i_8_1406, i_8_1473, i_8_1527, i_8_1528, i_8_1536, i_8_1548, i_8_1588, i_8_1589, i_8_1634, i_8_1676, i_8_1700, i_8_1707, i_8_1717, i_8_1727, i_8_1729, i_8_1732, i_8_1751, i_8_1796, i_8_1807, i_8_1808, i_8_1814, i_8_1858, i_8_1859, i_8_1903, i_8_1904, i_8_1918, i_8_1921, i_8_1930, i_8_1976, i_8_1984, i_8_2011, i_8_2012, i_8_2028, i_8_2029, i_8_2032, i_8_2151, i_8_2174, i_8_2215, i_8_2216, i_8_2292, o_8_58);
	kernel_8_59 k_8_59(i_8_20, i_8_29, i_8_30, i_8_47, i_8_50, i_8_56, i_8_74, i_8_77, i_8_112, i_8_113, i_8_137, i_8_165, i_8_229, i_8_253, i_8_254, i_8_256, i_8_262, i_8_376, i_8_420, i_8_442, i_8_451, i_8_452, i_8_454, i_8_455, i_8_590, i_8_596, i_8_644, i_8_665, i_8_677, i_8_694, i_8_695, i_8_707, i_8_776, i_8_784, i_8_796, i_8_823, i_8_875, i_8_878, i_8_965, i_8_991, i_8_994, i_8_1038, i_8_1111, i_8_1120, i_8_1139, i_8_1163, i_8_1202, i_8_1226, i_8_1253, i_8_1255, i_8_1260, i_8_1289, i_8_1318, i_8_1334, i_8_1342, i_8_1379, i_8_1400, i_8_1487, i_8_1538, i_8_1546, i_8_1552, i_8_1559, i_8_1631, i_8_1637, i_8_1666, i_8_1675, i_8_1679, i_8_1681, i_8_1682, i_8_1687, i_8_1697, i_8_1701, i_8_1755, i_8_1757, i_8_1770, i_8_1772, i_8_1784, i_8_1789, i_8_1840, i_8_1882, i_8_1885, i_8_1904, i_8_1910, i_8_1918, i_8_1960, i_8_1984, i_8_1990, i_8_1994, i_8_1995, i_8_2033, i_8_2075, i_8_2099, i_8_2108, i_8_2136, i_8_2146, i_8_2156, i_8_2224, i_8_2233, i_8_2241, i_8_2260, o_8_59);
	kernel_8_60 k_8_60(i_8_25, i_8_41, i_8_44, i_8_88, i_8_116, i_8_248, i_8_283, i_8_363, i_8_365, i_8_389, i_8_400, i_8_419, i_8_422, i_8_430, i_8_472, i_8_473, i_8_493, i_8_508, i_8_517, i_8_527, i_8_574, i_8_575, i_8_580, i_8_581, i_8_592, i_8_593, i_8_604, i_8_608, i_8_661, i_8_679, i_8_680, i_8_693, i_8_697, i_8_751, i_8_752, i_8_781, i_8_824, i_8_833, i_8_839, i_8_841, i_8_848, i_8_881, i_8_882, i_8_886, i_8_895, i_8_955, i_8_1036, i_8_1040, i_8_1103, i_8_1111, i_8_1129, i_8_1184, i_8_1238, i_8_1241, i_8_1318, i_8_1325, i_8_1330, i_8_1337, i_8_1353, i_8_1358, i_8_1363, i_8_1364, i_8_1427, i_8_1436, i_8_1444, i_8_1480, i_8_1481, i_8_1490, i_8_1532, i_8_1552, i_8_1633, i_8_1651, i_8_1664, i_8_1682, i_8_1694, i_8_1697, i_8_1706, i_8_1733, i_8_1751, i_8_1772, i_8_1774, i_8_1775, i_8_1781, i_8_1784, i_8_1787, i_8_1790, i_8_1810, i_8_1855, i_8_1858, i_8_1859, i_8_1867, i_8_1877, i_8_1913, i_8_1975, i_8_1978, i_8_1997, i_8_2137, i_8_2150, i_8_2177, i_8_2249, o_8_60);
	kernel_8_61 k_8_61(i_8_11, i_8_19, i_8_21, i_8_22, i_8_102, i_8_219, i_8_224, i_8_265, i_8_306, i_8_391, i_8_398, i_8_404, i_8_429, i_8_437, i_8_464, i_8_487, i_8_488, i_8_530, i_8_538, i_8_565, i_8_583, i_8_590, i_8_601, i_8_610, i_8_646, i_8_657, i_8_661, i_8_664, i_8_696, i_8_709, i_8_749, i_8_754, i_8_781, i_8_783, i_8_797, i_8_799, i_8_842, i_8_858, i_8_869, i_8_894, i_8_994, i_8_1035, i_8_1065, i_8_1067, i_8_1137, i_8_1138, i_8_1139, i_8_1189, i_8_1190, i_8_1202, i_8_1249, i_8_1266, i_8_1292, i_8_1294, i_8_1298, i_8_1317, i_8_1363, i_8_1373, i_8_1425, i_8_1443, i_8_1444, i_8_1446, i_8_1508, i_8_1550, i_8_1605, i_8_1606, i_8_1607, i_8_1746, i_8_1747, i_8_1748, i_8_1752, i_8_1759, i_8_1771, i_8_1773, i_8_1778, i_8_1816, i_8_1823, i_8_1825, i_8_1831, i_8_1835, i_8_1841, i_8_1888, i_8_1907, i_8_1951, i_8_1963, i_8_1966, i_8_1972, i_8_1993, i_8_1995, i_8_2032, i_8_2043, i_8_2052, i_8_2053, i_8_2110, i_8_2166, i_8_2169, i_8_2225, i_8_2237, i_8_2244, i_8_2293, o_8_61);
	kernel_8_62 k_8_62(i_8_35, i_8_61, i_8_96, i_8_97, i_8_258, i_8_325, i_8_328, i_8_331, i_8_367, i_8_372, i_8_381, i_8_382, i_8_458, i_8_465, i_8_467, i_8_487, i_8_504, i_8_525, i_8_552, i_8_586, i_8_590, i_8_610, i_8_630, i_8_632, i_8_633, i_8_637, i_8_661, i_8_664, i_8_693, i_8_694, i_8_698, i_8_762, i_8_763, i_8_768, i_8_790, i_8_855, i_8_876, i_8_877, i_8_879, i_8_995, i_8_998, i_8_1137, i_8_1195, i_8_1236, i_8_1237, i_8_1239, i_8_1240, i_8_1261, i_8_1264, i_8_1285, i_8_1296, i_8_1297, i_8_1299, i_8_1333, i_8_1369, i_8_1396, i_8_1399, i_8_1410, i_8_1489, i_8_1535, i_8_1536, i_8_1538, i_8_1591, i_8_1599, i_8_1600, i_8_1602, i_8_1605, i_8_1629, i_8_1630, i_8_1704, i_8_1722, i_8_1744, i_8_1746, i_8_1791, i_8_1792, i_8_1795, i_8_1842, i_8_1843, i_8_1854, i_8_1855, i_8_1900, i_8_1903, i_8_1915, i_8_1947, i_8_1951, i_8_1969, i_8_2004, i_8_2047, i_8_2146, i_8_2154, i_8_2155, i_8_2156, i_8_2194, i_8_2218, i_8_2233, i_8_2246, i_8_2263, i_8_2264, i_8_2298, i_8_2299, o_8_62);
	kernel_8_63 k_8_63(i_8_26, i_8_77, i_8_89, i_8_160, i_8_161, i_8_224, i_8_259, i_8_286, i_8_296, i_8_312, i_8_337, i_8_349, i_8_367, i_8_404, i_8_422, i_8_457, i_8_485, i_8_525, i_8_526, i_8_556, i_8_606, i_8_628, i_8_636, i_8_682, i_8_694, i_8_696, i_8_718, i_8_763, i_8_818, i_8_843, i_8_844, i_8_872, i_8_898, i_8_926, i_8_951, i_8_952, i_8_953, i_8_958, i_8_980, i_8_1016, i_8_1033, i_8_1086, i_8_1106, i_8_1114, i_8_1151, i_8_1222, i_8_1223, i_8_1273, i_8_1274, i_8_1282, i_8_1286, i_8_1314, i_8_1324, i_8_1328, i_8_1393, i_8_1404, i_8_1411, i_8_1437, i_8_1447, i_8_1457, i_8_1471, i_8_1484, i_8_1524, i_8_1528, i_8_1534, i_8_1537, i_8_1546, i_8_1547, i_8_1574, i_8_1582, i_8_1591, i_8_1628, i_8_1636, i_8_1655, i_8_1658, i_8_1672, i_8_1690, i_8_1750, i_8_1753, i_8_1807, i_8_1815, i_8_1823, i_8_1825, i_8_1834, i_8_1840, i_8_1861, i_8_1870, i_8_1880, i_8_1888, i_8_1903, i_8_1905, i_8_1906, i_8_1907, i_8_1975, i_8_1986, i_8_2005, i_8_2049, i_8_2051, i_8_2060, i_8_2274, o_8_63);
	kernel_8_64 k_8_64(i_8_12, i_8_13, i_8_62, i_8_75, i_8_89, i_8_129, i_8_130, i_8_193, i_8_223, i_8_363, i_8_365, i_8_366, i_8_390, i_8_426, i_8_499, i_8_522, i_8_526, i_8_528, i_8_530, i_8_591, i_8_593, i_8_604, i_8_609, i_8_610, i_8_627, i_8_637, i_8_654, i_8_660, i_8_661, i_8_665, i_8_678, i_8_681, i_8_705, i_8_708, i_8_718, i_8_815, i_8_834, i_8_835, i_8_894, i_8_1032, i_8_1033, i_8_1078, i_8_1266, i_8_1272, i_8_1274, i_8_1302, i_8_1308, i_8_1338, i_8_1339, i_8_1340, i_8_1398, i_8_1403, i_8_1434, i_8_1439, i_8_1449, i_8_1461, i_8_1464, i_8_1507, i_8_1547, i_8_1599, i_8_1601, i_8_1625, i_8_1627, i_8_1636, i_8_1637, i_8_1641, i_8_1643, i_8_1662, i_8_1731, i_8_1734, i_8_1749, i_8_1779, i_8_1780, i_8_1787, i_8_1788, i_8_1789, i_8_1790, i_8_1804, i_8_1851, i_8_1853, i_8_1857, i_8_1860, i_8_1861, i_8_1866, i_8_1867, i_8_1869, i_8_1879, i_8_1905, i_8_1906, i_8_1907, i_8_1951, i_8_1952, i_8_2032, i_8_2040, i_8_2092, i_8_2093, i_8_2158, i_8_2215, i_8_2242, i_8_2249, o_8_64);
	kernel_8_65 k_8_65(i_8_43, i_8_53, i_8_76, i_8_127, i_8_145, i_8_196, i_8_210, i_8_284, i_8_301, i_8_319, i_8_325, i_8_328, i_8_347, i_8_361, i_8_384, i_8_390, i_8_453, i_8_454, i_8_508, i_8_526, i_8_562, i_8_583, i_8_599, i_8_608, i_8_611, i_8_643, i_8_656, i_8_658, i_8_664, i_8_695, i_8_697, i_8_709, i_8_710, i_8_775, i_8_792, i_8_839, i_8_840, i_8_895, i_8_926, i_8_967, i_8_968, i_8_1015, i_8_1074, i_8_1103, i_8_1106, i_8_1107, i_8_1115, i_8_1126, i_8_1183, i_8_1204, i_8_1231, i_8_1240, i_8_1263, i_8_1264, i_8_1267, i_8_1268, i_8_1286, i_8_1299, i_8_1339, i_8_1365, i_8_1410, i_8_1436, i_8_1444, i_8_1474, i_8_1490, i_8_1525, i_8_1546, i_8_1572, i_8_1603, i_8_1607, i_8_1609, i_8_1669, i_8_1690, i_8_1749, i_8_1751, i_8_1780, i_8_1786, i_8_1787, i_8_1806, i_8_1825, i_8_1886, i_8_1915, i_8_1930, i_8_1948, i_8_1949, i_8_1950, i_8_1992, i_8_1994, i_8_1995, i_8_2112, i_8_2142, i_8_2144, i_8_2147, i_8_2148, i_8_2150, i_8_2212, i_8_2260, i_8_2272, i_8_2290, i_8_2294, o_8_65);
	kernel_8_66 k_8_66(i_8_27, i_8_30, i_8_78, i_8_79, i_8_114, i_8_165, i_8_166, i_8_192, i_8_193, i_8_211, i_8_224, i_8_234, i_8_237, i_8_238, i_8_240, i_8_241, i_8_301, i_8_302, i_8_337, i_8_338, i_8_346, i_8_384, i_8_462, i_8_476, i_8_489, i_8_510, i_8_525, i_8_591, i_8_592, i_8_593, i_8_600, i_8_602, i_8_604, i_8_616, i_8_617, i_8_658, i_8_701, i_8_710, i_8_717, i_8_720, i_8_747, i_8_774, i_8_787, i_8_804, i_8_825, i_8_850, i_8_864, i_8_996, i_8_1047, i_8_1056, i_8_1120, i_8_1128, i_8_1260, i_8_1279, i_8_1284, i_8_1292, i_8_1306, i_8_1410, i_8_1412, i_8_1437, i_8_1438, i_8_1527, i_8_1528, i_8_1572, i_8_1611, i_8_1624, i_8_1625, i_8_1632, i_8_1633, i_8_1634, i_8_1635, i_8_1637, i_8_1653, i_8_1654, i_8_1655, i_8_1672, i_8_1699, i_8_1754, i_8_1782, i_8_1824, i_8_1832, i_8_1854, i_8_1857, i_8_1947, i_8_1983, i_8_1984, i_8_1992, i_8_1993, i_8_1994, i_8_1997, i_8_2031, i_8_2040, i_8_2076, i_8_2077, i_8_2088, i_8_2154, i_8_2212, i_8_2214, i_8_2259, i_8_2262, o_8_66);
	kernel_8_67 k_8_67(i_8_3, i_8_26, i_8_31, i_8_64, i_8_75, i_8_84, i_8_111, i_8_114, i_8_138, i_8_229, i_8_300, i_8_301, i_8_304, i_8_318, i_8_352, i_8_399, i_8_416, i_8_420, i_8_437, i_8_469, i_8_470, i_8_553, i_8_567, i_8_570, i_8_579, i_8_591, i_8_598, i_8_607, i_8_624, i_8_633, i_8_667, i_8_676, i_8_699, i_8_705, i_8_729, i_8_811, i_8_832, i_8_838, i_8_839, i_8_840, i_8_955, i_8_956, i_8_959, i_8_1101, i_8_1107, i_8_1152, i_8_1225, i_8_1228, i_8_1234, i_8_1296, i_8_1298, i_8_1318, i_8_1326, i_8_1335, i_8_1344, i_8_1353, i_8_1397, i_8_1399, i_8_1431, i_8_1432, i_8_1434, i_8_1440, i_8_1483, i_8_1487, i_8_1492, i_8_1495, i_8_1521, i_8_1624, i_8_1635, i_8_1642, i_8_1647, i_8_1686, i_8_1696, i_8_1705, i_8_1768, i_8_1779, i_8_1786, i_8_1804, i_8_1806, i_8_1807, i_8_1813, i_8_1827, i_8_1836, i_8_1848, i_8_1911, i_8_1915, i_8_1917, i_8_2038, i_8_2045, i_8_2056, i_8_2065, i_8_2073, i_8_2074, i_8_2090, i_8_2119, i_8_2120, i_8_2190, i_8_2244, i_8_2272, i_8_2297, o_8_67);
	kernel_8_68 k_8_68(i_8_29, i_8_49, i_8_52, i_8_95, i_8_131, i_8_173, i_8_328, i_8_337, i_8_364, i_8_371, i_8_373, i_8_434, i_8_445, i_8_454, i_8_475, i_8_510, i_8_527, i_8_528, i_8_596, i_8_630, i_8_667, i_8_717, i_8_753, i_8_760, i_8_777, i_8_780, i_8_826, i_8_827, i_8_840, i_8_841, i_8_842, i_8_843, i_8_844, i_8_886, i_8_901, i_8_943, i_8_977, i_8_1031, i_8_1046, i_8_1103, i_8_1248, i_8_1249, i_8_1259, i_8_1300, i_8_1401, i_8_1427, i_8_1434, i_8_1435, i_8_1438, i_8_1439, i_8_1450, i_8_1451, i_8_1471, i_8_1533, i_8_1534, i_8_1535, i_8_1543, i_8_1544, i_8_1547, i_8_1573, i_8_1606, i_8_1626, i_8_1627, i_8_1628, i_8_1634, i_8_1637, i_8_1648, i_8_1678, i_8_1679, i_8_1681, i_8_1682, i_8_1701, i_8_1705, i_8_1723, i_8_1748, i_8_1753, i_8_1758, i_8_1759, i_8_1760, i_8_1761, i_8_1762, i_8_1763, i_8_1767, i_8_1774, i_8_1777, i_8_1857, i_8_1877, i_8_1929, i_8_1940, i_8_1966, i_8_1980, i_8_1993, i_8_2003, i_8_2109, i_8_2110, i_8_2119, i_8_2150, i_8_2214, i_8_2215, i_8_2216, o_8_68);
	kernel_8_69 k_8_69(i_8_3, i_8_6, i_8_7, i_8_98, i_8_115, i_8_203, i_8_205, i_8_206, i_8_226, i_8_227, i_8_228, i_8_229, i_8_230, i_8_231, i_8_232, i_8_233, i_8_248, i_8_325, i_8_356, i_8_357, i_8_383, i_8_497, i_8_499, i_8_501, i_8_502, i_8_571, i_8_572, i_8_574, i_8_605, i_8_606, i_8_609, i_8_610, i_8_611, i_8_671, i_8_672, i_8_714, i_8_716, i_8_717, i_8_812, i_8_822, i_8_838, i_8_883, i_8_884, i_8_888, i_8_889, i_8_890, i_8_930, i_8_932, i_8_934, i_8_958, i_8_966, i_8_990, i_8_1047, i_8_1049, i_8_1175, i_8_1236, i_8_1256, i_8_1258, i_8_1272, i_8_1279, i_8_1300, i_8_1336, i_8_1446, i_8_1491, i_8_1642, i_8_1648, i_8_1720, i_8_1721, i_8_1724, i_8_1747, i_8_1768, i_8_1769, i_8_1789, i_8_1805, i_8_1807, i_8_1818, i_8_1849, i_8_1850, i_8_1858, i_8_1865, i_8_1866, i_8_1868, i_8_1871, i_8_1980, i_8_1982, i_8_1983, i_8_1995, i_8_2074, i_8_2104, i_8_2142, i_8_2143, i_8_2145, i_8_2153, i_8_2176, i_8_2245, i_8_2246, i_8_2275, i_8_2289, i_8_2290, i_8_2291, o_8_69);
	kernel_8_70 k_8_70(i_8_21, i_8_28, i_8_31, i_8_46, i_8_101, i_8_119, i_8_136, i_8_230, i_8_232, i_8_298, i_8_302, i_8_316, i_8_326, i_8_374, i_8_388, i_8_423, i_8_468, i_8_489, i_8_490, i_8_521, i_8_551, i_8_556, i_8_608, i_8_616, i_8_622, i_8_623, i_8_634, i_8_637, i_8_649, i_8_677, i_8_684, i_8_692, i_8_702, i_8_704, i_8_830, i_8_839, i_8_958, i_8_974, i_8_982, i_8_983, i_8_992, i_8_1000, i_8_1001, i_8_1037, i_8_1046, i_8_1089, i_8_1216, i_8_1262, i_8_1271, i_8_1309, i_8_1345, i_8_1370, i_8_1388, i_8_1423, i_8_1424, i_8_1433, i_8_1460, i_8_1462, i_8_1463, i_8_1478, i_8_1493, i_8_1495, i_8_1514, i_8_1522, i_8_1536, i_8_1550, i_8_1586, i_8_1600, i_8_1671, i_8_1674, i_8_1678, i_8_1711, i_8_1714, i_8_1721, i_8_1724, i_8_1746, i_8_1747, i_8_1784, i_8_1805, i_8_1808, i_8_1821, i_8_1823, i_8_1854, i_8_1891, i_8_1901, i_8_2008, i_8_2038, i_8_2039, i_8_2054, i_8_2065, i_8_2075, i_8_2098, i_8_2120, i_8_2143, i_8_2149, i_8_2215, i_8_2225, i_8_2230, i_8_2243, i_8_2260, o_8_70);
	kernel_8_71 k_8_71(i_8_22, i_8_29, i_8_80, i_8_112, i_8_139, i_8_148, i_8_221, i_8_224, i_8_256, i_8_296, i_8_304, i_8_305, i_8_329, i_8_377, i_8_414, i_8_457, i_8_485, i_8_486, i_8_549, i_8_550, i_8_551, i_8_554, i_8_578, i_8_585, i_8_586, i_8_587, i_8_590, i_8_596, i_8_605, i_8_612, i_8_638, i_8_662, i_8_675, i_8_676, i_8_677, i_8_699, i_8_716, i_8_719, i_8_784, i_8_790, i_8_821, i_8_822, i_8_838, i_8_839, i_8_851, i_8_864, i_8_865, i_8_946, i_8_983, i_8_1045, i_8_1046, i_8_1100, i_8_1130, i_8_1201, i_8_1233, i_8_1243, i_8_1267, i_8_1305, i_8_1308, i_8_1316, i_8_1355, i_8_1404, i_8_1405, i_8_1438, i_8_1453, i_8_1458, i_8_1477, i_8_1478, i_8_1486, i_8_1510, i_8_1550, i_8_1557, i_8_1558, i_8_1559, i_8_1603, i_8_1620, i_8_1647, i_8_1650, i_8_1669, i_8_1671, i_8_1694, i_8_1712, i_8_1730, i_8_1746, i_8_1757, i_8_1780, i_8_1792, i_8_1881, i_8_1882, i_8_1883, i_8_1944, i_8_1946, i_8_1965, i_8_1989, i_8_1990, i_8_2093, i_8_2135, i_8_2144, i_8_2268, i_8_2296, o_8_71);
	kernel_8_72 k_8_72(i_8_19, i_8_49, i_8_52, i_8_53, i_8_66, i_8_74, i_8_87, i_8_103, i_8_107, i_8_223, i_8_243, i_8_284, i_8_288, i_8_289, i_8_325, i_8_367, i_8_418, i_8_427, i_8_436, i_8_491, i_8_523, i_8_525, i_8_526, i_8_528, i_8_530, i_8_598, i_8_604, i_8_608, i_8_630, i_8_631, i_8_643, i_8_657, i_8_683, i_8_690, i_8_693, i_8_694, i_8_696, i_8_698, i_8_702, i_8_703, i_8_706, i_8_709, i_8_710, i_8_720, i_8_721, i_8_723, i_8_724, i_8_725, i_8_734, i_8_763, i_8_778, i_8_801, i_8_805, i_8_806, i_8_829, i_8_838, i_8_877, i_8_967, i_8_969, i_8_970, i_8_976, i_8_1026, i_8_1112, i_8_1183, i_8_1261, i_8_1262, i_8_1264, i_8_1282, i_8_1299, i_8_1317, i_8_1327, i_8_1352, i_8_1362, i_8_1400, i_8_1407, i_8_1408, i_8_1435, i_8_1445, i_8_1486, i_8_1544, i_8_1588, i_8_1622, i_8_1750, i_8_1776, i_8_1777, i_8_1855, i_8_1882, i_8_1885, i_8_1904, i_8_1964, i_8_1984, i_8_2025, i_8_2028, i_8_2038, i_8_2115, i_8_2116, i_8_2151, i_8_2191, i_8_2228, i_8_2241, o_8_72);
	kernel_8_73 k_8_73(i_8_32, i_8_33, i_8_48, i_8_52, i_8_58, i_8_61, i_8_85, i_8_120, i_8_141, i_8_170, i_8_183, i_8_222, i_8_223, i_8_259, i_8_295, i_8_301, i_8_312, i_8_328, i_8_373, i_8_391, i_8_440, i_8_480, i_8_481, i_8_483, i_8_500, i_8_502, i_8_507, i_8_527, i_8_530, i_8_556, i_8_594, i_8_607, i_8_687, i_8_690, i_8_759, i_8_786, i_8_787, i_8_789, i_8_800, i_8_844, i_8_849, i_8_862, i_8_868, i_8_876, i_8_947, i_8_994, i_8_1050, i_8_1060, i_8_1075, i_8_1120, i_8_1218, i_8_1219, i_8_1221, i_8_1222, i_8_1282, i_8_1305, i_8_1306, i_8_1307, i_8_1308, i_8_1314, i_8_1330, i_8_1345, i_8_1387, i_8_1390, i_8_1410, i_8_1471, i_8_1506, i_8_1509, i_8_1545, i_8_1547, i_8_1551, i_8_1555, i_8_1560, i_8_1570, i_8_1654, i_8_1677, i_8_1683, i_8_1707, i_8_1722, i_8_1726, i_8_1738, i_8_1740, i_8_1749, i_8_1750, i_8_1752, i_8_1753, i_8_1761, i_8_1788, i_8_1791, i_8_1804, i_8_1879, i_8_1906, i_8_2028, i_8_2046, i_8_2092, i_8_2145, i_8_2172, i_8_2215, i_8_2216, i_8_2285, o_8_73);
	kernel_8_74 k_8_74(i_8_82, i_8_136, i_8_139, i_8_157, i_8_208, i_8_255, i_8_289, i_8_297, i_8_339, i_8_343, i_8_387, i_8_388, i_8_392, i_8_445, i_8_450, i_8_451, i_8_460, i_8_507, i_8_508, i_8_529, i_8_540, i_8_549, i_8_595, i_8_598, i_8_603, i_8_604, i_8_610, i_8_621, i_8_669, i_8_679, i_8_711, i_8_712, i_8_716, i_8_735, i_8_748, i_8_760, i_8_765, i_8_766, i_8_770, i_8_793, i_8_814, i_8_828, i_8_844, i_8_877, i_8_907, i_8_939, i_8_946, i_8_994, i_8_1011, i_8_1012, i_8_1026, i_8_1071, i_8_1074, i_8_1081, i_8_1099, i_8_1108, i_8_1137, i_8_1251, i_8_1267, i_8_1323, i_8_1324, i_8_1344, i_8_1367, i_8_1441, i_8_1480, i_8_1503, i_8_1524, i_8_1548, i_8_1549, i_8_1552, i_8_1594, i_8_1597, i_8_1602, i_8_1605, i_8_1606, i_8_1611, i_8_1642, i_8_1648, i_8_1675, i_8_1681, i_8_1695, i_8_1701, i_8_1720, i_8_1730, i_8_1749, i_8_1776, i_8_1778, i_8_1779, i_8_1812, i_8_1819, i_8_1821, i_8_1890, i_8_1891, i_8_1947, i_8_1963, i_8_1994, i_8_2070, i_8_2140, i_8_2150, i_8_2214, o_8_74);
	kernel_8_75 k_8_75(i_8_33, i_8_35, i_8_40, i_8_42, i_8_78, i_8_105, i_8_142, i_8_150, i_8_172, i_8_184, i_8_190, i_8_193, i_8_223, i_8_313, i_8_321, i_8_330, i_8_364, i_8_417, i_8_420, i_8_453, i_8_507, i_8_510, i_8_524, i_8_528, i_8_537, i_8_555, i_8_571, i_8_601, i_8_607, i_8_664, i_8_665, i_8_687, i_8_696, i_8_701, i_8_753, i_8_799, i_8_837, i_8_840, i_8_844, i_8_845, i_8_877, i_8_897, i_8_945, i_8_946, i_8_951, i_8_952, i_8_978, i_8_993, i_8_1014, i_8_1015, i_8_1120, i_8_1129, i_8_1158, i_8_1239, i_8_1257, i_8_1330, i_8_1339, i_8_1425, i_8_1464, i_8_1469, i_8_1482, i_8_1515, i_8_1527, i_8_1528, i_8_1536, i_8_1549, i_8_1555, i_8_1560, i_8_1572, i_8_1617, i_8_1647, i_8_1653, i_8_1662, i_8_1686, i_8_1689, i_8_1752, i_8_1807, i_8_1822, i_8_1861, i_8_1884, i_8_1887, i_8_1894, i_8_1914, i_8_1933, i_8_1951, i_8_1983, i_8_1995, i_8_1996, i_8_2050, i_8_2095, i_8_2104, i_8_2116, i_8_2128, i_8_2139, i_8_2152, i_8_2153, i_8_2183, i_8_2190, i_8_2226, i_8_2248, o_8_75);
	kernel_8_76 k_8_76(i_8_1, i_8_77, i_8_115, i_8_318, i_8_319, i_8_362, i_8_368, i_8_398, i_8_464, i_8_505, i_8_526, i_8_571, i_8_575, i_8_578, i_8_580, i_8_581, i_8_587, i_8_589, i_8_595, i_8_607, i_8_610, i_8_634, i_8_636, i_8_637, i_8_692, i_8_707, i_8_784, i_8_840, i_8_844, i_8_883, i_8_892, i_8_967, i_8_995, i_8_1036, i_8_1037, i_8_1072, i_8_1103, i_8_1111, i_8_1127, i_8_1262, i_8_1264, i_8_1271, i_8_1298, i_8_1300, i_8_1315, i_8_1328, i_8_1334, i_8_1336, i_8_1337, i_8_1363, i_8_1400, i_8_1440, i_8_1441, i_8_1462, i_8_1471, i_8_1515, i_8_1524, i_8_1526, i_8_1544, i_8_1553, i_8_1558, i_8_1595, i_8_1603, i_8_1655, i_8_1684, i_8_1697, i_8_1700, i_8_1703, i_8_1706, i_8_1747, i_8_1748, i_8_1795, i_8_1819, i_8_1825, i_8_1867, i_8_1869, i_8_1871, i_8_1885, i_8_1888, i_8_1912, i_8_1913, i_8_1927, i_8_1950, i_8_2045, i_8_2122, i_8_2150, i_8_2154, i_8_2155, i_8_2157, i_8_2176, i_8_2190, i_8_2191, i_8_2218, i_8_2223, i_8_2224, i_8_2225, i_8_2243, i_8_2245, i_8_2286, i_8_2297, o_8_76);
	kernel_8_77 k_8_77(i_8_12, i_8_27, i_8_28, i_8_33, i_8_34, i_8_40, i_8_58, i_8_102, i_8_165, i_8_166, i_8_183, i_8_186, i_8_231, i_8_298, i_8_304, i_8_310, i_8_336, i_8_337, i_8_365, i_8_368, i_8_379, i_8_380, i_8_418, i_8_424, i_8_426, i_8_444, i_8_454, i_8_467, i_8_480, i_8_483, i_8_507, i_8_508, i_8_529, i_8_543, i_8_544, i_8_556, i_8_580, i_8_588, i_8_615, i_8_675, i_8_678, i_8_679, i_8_687, i_8_694, i_8_702, i_8_705, i_8_729, i_8_763, i_8_781, i_8_817, i_8_849, i_8_885, i_8_886, i_8_921, i_8_959, i_8_967, i_8_1054, i_8_1059, i_8_1103, i_8_1108, i_8_1192, i_8_1267, i_8_1284, i_8_1285, i_8_1290, i_8_1299, i_8_1326, i_8_1333, i_8_1354, i_8_1389, i_8_1395, i_8_1432, i_8_1468, i_8_1641, i_8_1649, i_8_1653, i_8_1690, i_8_1731, i_8_1740, i_8_1741, i_8_1769, i_8_1824, i_8_1825, i_8_1828, i_8_1831, i_8_1837, i_8_1884, i_8_1948, i_8_1983, i_8_1984, i_8_2002, i_8_2040, i_8_2047, i_8_2134, i_8_2146, i_8_2172, i_8_2214, i_8_2215, i_8_2248, i_8_2299, o_8_77);
	kernel_8_78 k_8_78(i_8_1, i_8_4, i_8_74, i_8_81, i_8_82, i_8_243, i_8_244, i_8_249, i_8_270, i_8_370, i_8_371, i_8_391, i_8_421, i_8_423, i_8_504, i_8_505, i_8_514, i_8_550, i_8_553, i_8_568, i_8_575, i_8_622, i_8_636, i_8_638, i_8_649, i_8_658, i_8_664, i_8_704, i_8_729, i_8_730, i_8_799, i_8_843, i_8_844, i_8_856, i_8_895, i_8_896, i_8_954, i_8_970, i_8_1005, i_8_1035, i_8_1071, i_8_1080, i_8_1098, i_8_1108, i_8_1156, i_8_1239, i_8_1260, i_8_1282, i_8_1297, i_8_1298, i_8_1318, i_8_1353, i_8_1359, i_8_1363, i_8_1396, i_8_1407, i_8_1426, i_8_1435, i_8_1469, i_8_1474, i_8_1481, i_8_1489, i_8_1494, i_8_1495, i_8_1516, i_8_1530, i_8_1531, i_8_1543, i_8_1552, i_8_1553, i_8_1555, i_8_1639, i_8_1651, i_8_1657, i_8_1672, i_8_1707, i_8_1746, i_8_1749, i_8_1750, i_8_1774, i_8_1780, i_8_1792, i_8_1819, i_8_1823, i_8_1846, i_8_1873, i_8_1877, i_8_1881, i_8_1888, i_8_1945, i_8_1948, i_8_2035, i_8_2044, i_8_2062, i_8_2074, i_8_2092, i_8_2122, i_8_2172, i_8_2173, i_8_2296, o_8_78);
	kernel_8_79 k_8_79(i_8_67, i_8_79, i_8_88, i_8_106, i_8_138, i_8_143, i_8_150, i_8_178, i_8_265, i_8_301, i_8_381, i_8_391, i_8_421, i_8_422, i_8_427, i_8_538, i_8_553, i_8_573, i_8_598, i_8_599, i_8_655, i_8_706, i_8_707, i_8_735, i_8_744, i_8_763, i_8_816, i_8_817, i_8_834, i_8_835, i_8_838, i_8_841, i_8_842, i_8_853, i_8_876, i_8_891, i_8_892, i_8_916, i_8_951, i_8_1087, i_8_1126, i_8_1127, i_8_1131, i_8_1135, i_8_1141, i_8_1178, i_8_1201, i_8_1267, i_8_1305, i_8_1306, i_8_1308, i_8_1338, i_8_1403, i_8_1410, i_8_1475, i_8_1481, i_8_1489, i_8_1492, i_8_1543, i_8_1544, i_8_1552, i_8_1601, i_8_1609, i_8_1645, i_8_1649, i_8_1651, i_8_1655, i_8_1690, i_8_1704, i_8_1709, i_8_1723, i_8_1750, i_8_1780, i_8_1814, i_8_1816, i_8_1824, i_8_1843, i_8_1855, i_8_1869, i_8_1885, i_8_1889, i_8_1912, i_8_1921, i_8_1957, i_8_1969, i_8_1976, i_8_1996, i_8_2023, i_8_2096, i_8_2119, i_8_2122, i_8_2141, i_8_2146, i_8_2150, i_8_2217, i_8_2218, i_8_2226, i_8_2227, i_8_2245, i_8_2299, o_8_79);
	kernel_8_80 k_8_80(i_8_38, i_8_41, i_8_50, i_8_57, i_8_60, i_8_62, i_8_95, i_8_166, i_8_239, i_8_260, i_8_300, i_8_319, i_8_335, i_8_338, i_8_365, i_8_382, i_8_421, i_8_425, i_8_427, i_8_437, i_8_490, i_8_493, i_8_496, i_8_497, i_8_552, i_8_554, i_8_555, i_8_556, i_8_584, i_8_604, i_8_613, i_8_653, i_8_658, i_8_676, i_8_700, i_8_751, i_8_755, i_8_761, i_8_799, i_8_800, i_8_803, i_8_932, i_8_968, i_8_1066, i_8_1073, i_8_1091, i_8_1156, i_8_1189, i_8_1264, i_8_1274, i_8_1282, i_8_1283, i_8_1285, i_8_1289, i_8_1292, i_8_1328, i_8_1355, i_8_1356, i_8_1382, i_8_1393, i_8_1409, i_8_1466, i_8_1472, i_8_1481, i_8_1552, i_8_1555, i_8_1562, i_8_1622, i_8_1625, i_8_1634, i_8_1651, i_8_1652, i_8_1655, i_8_1660, i_8_1669, i_8_1688, i_8_1706, i_8_1777, i_8_1781, i_8_1819, i_8_1828, i_8_1832, i_8_1867, i_8_1904, i_8_1939, i_8_1940, i_8_1943, i_8_1993, i_8_2005, i_8_2026, i_8_2107, i_8_2146, i_8_2153, i_8_2155, i_8_2156, i_8_2165, i_8_2179, i_8_2210, i_8_2225, i_8_2227, o_8_80);
	kernel_8_81 k_8_81(i_8_45, i_8_108, i_8_111, i_8_120, i_8_156, i_8_160, i_8_229, i_8_230, i_8_291, i_8_330, i_8_345, i_8_381, i_8_391, i_8_433, i_8_434, i_8_437, i_8_483, i_8_485, i_8_486, i_8_489, i_8_493, i_8_502, i_8_588, i_8_593, i_8_606, i_8_621, i_8_624, i_8_627, i_8_669, i_8_670, i_8_687, i_8_694, i_8_703, i_8_705, i_8_706, i_8_707, i_8_714, i_8_716, i_8_718, i_8_723, i_8_724, i_8_774, i_8_780, i_8_781, i_8_807, i_8_822, i_8_823, i_8_825, i_8_826, i_8_827, i_8_848, i_8_873, i_8_875, i_8_973, i_8_991, i_8_1015, i_8_1027, i_8_1029, i_8_1030, i_8_1059, i_8_1233, i_8_1254, i_8_1270, i_8_1288, i_8_1300, i_8_1318, i_8_1346, i_8_1356, i_8_1398, i_8_1399, i_8_1426, i_8_1437, i_8_1443, i_8_1587, i_8_1625, i_8_1645, i_8_1649, i_8_1652, i_8_1773, i_8_1803, i_8_1823, i_8_1824, i_8_1825, i_8_1854, i_8_1858, i_8_1864, i_8_1882, i_8_1884, i_8_1885, i_8_1951, i_8_1968, i_8_2026, i_8_2029, i_8_2073, i_8_2091, i_8_2122, i_8_2172, i_8_2242, i_8_2273, i_8_2290, o_8_81);
	kernel_8_82 k_8_82(i_8_18, i_8_31, i_8_89, i_8_93, i_8_200, i_8_211, i_8_230, i_8_301, i_8_343, i_8_374, i_8_378, i_8_379, i_8_440, i_8_453, i_8_454, i_8_462, i_8_476, i_8_551, i_8_557, i_8_568, i_8_572, i_8_588, i_8_596, i_8_601, i_8_611, i_8_615, i_8_616, i_8_621, i_8_633, i_8_660, i_8_672, i_8_693, i_8_732, i_8_772, i_8_779, i_8_795, i_8_796, i_8_811, i_8_846, i_8_847, i_8_850, i_8_855, i_8_856, i_8_946, i_8_980, i_8_1012, i_8_1027, i_8_1065, i_8_1088, i_8_1125, i_8_1128, i_8_1137, i_8_1183, i_8_1191, i_8_1255, i_8_1256, i_8_1281, i_8_1307, i_8_1309, i_8_1391, i_8_1437, i_8_1439, i_8_1450, i_8_1488, i_8_1489, i_8_1525, i_8_1528, i_8_1538, i_8_1541, i_8_1587, i_8_1588, i_8_1614, i_8_1624, i_8_1630, i_8_1632, i_8_1669, i_8_1702, i_8_1724, i_8_1728, i_8_1741, i_8_1742, i_8_1795, i_8_1808, i_8_1818, i_8_1839, i_8_1845, i_8_1858, i_8_1870, i_8_1884, i_8_1903, i_8_1906, i_8_1966, i_8_1995, i_8_2048, i_8_2151, i_8_2188, i_8_2216, i_8_2217, i_8_2291, i_8_2299, o_8_82);
	kernel_8_83 k_8_83(i_8_25, i_8_26, i_8_41, i_8_44, i_8_86, i_8_107, i_8_176, i_8_191, i_8_214, i_8_215, i_8_314, i_8_331, i_8_347, i_8_377, i_8_430, i_8_440, i_8_457, i_8_469, i_8_470, i_8_493, i_8_499, i_8_500, i_8_502, i_8_611, i_8_629, i_8_637, i_8_661, i_8_664, i_8_665, i_8_733, i_8_764, i_8_772, i_8_773, i_8_799, i_8_985, i_8_995, i_8_1012, i_8_1015, i_8_1024, i_8_1033, i_8_1060, i_8_1097, i_8_1132, i_8_1160, i_8_1175, i_8_1187, i_8_1258, i_8_1268, i_8_1310, i_8_1313, i_8_1348, i_8_1350, i_8_1358, i_8_1411, i_8_1412, i_8_1592, i_8_1596, i_8_1609, i_8_1636, i_8_1649, i_8_1655, i_8_1675, i_8_1691, i_8_1736, i_8_1753, i_8_1754, i_8_1858, i_8_1870, i_8_1871, i_8_1889, i_8_1897, i_8_1907, i_8_1917, i_8_1919, i_8_1922, i_8_1990, i_8_1995, i_8_2002, i_8_2005, i_8_2006, i_8_2023, i_8_2122, i_8_2123, i_8_2132, i_8_2158, i_8_2159, i_8_2164, i_8_2174, i_8_2176, i_8_2186, i_8_2195, i_8_2203, i_8_2215, i_8_2216, i_8_2218, i_8_2263, i_8_2276, i_8_2281, i_8_2284, i_8_2294, o_8_83);
	kernel_8_84 k_8_84(i_8_30, i_8_87, i_8_103, i_8_224, i_8_255, i_8_259, i_8_296, i_8_301, i_8_305, i_8_327, i_8_328, i_8_336, i_8_364, i_8_386, i_8_420, i_8_422, i_8_440, i_8_447, i_8_448, i_8_454, i_8_476, i_8_483, i_8_485, i_8_495, i_8_555, i_8_557, i_8_592, i_8_593, i_8_603, i_8_616, i_8_619, i_8_628, i_8_649, i_8_663, i_8_664, i_8_682, i_8_763, i_8_764, i_8_817, i_8_850, i_8_853, i_8_880, i_8_881, i_8_951, i_8_952, i_8_986, i_8_1032, i_8_1059, i_8_1071, i_8_1075, i_8_1114, i_8_1124, i_8_1307, i_8_1308, i_8_1311, i_8_1329, i_8_1330, i_8_1341, i_8_1349, i_8_1431, i_8_1432, i_8_1533, i_8_1537, i_8_1591, i_8_1600, i_8_1633, i_8_1637, i_8_1654, i_8_1671, i_8_1680, i_8_1723, i_8_1734, i_8_1743, i_8_1744, i_8_1749, i_8_1751, i_8_1786, i_8_1787, i_8_1790, i_8_1807, i_8_1837, i_8_1839, i_8_1844, i_8_1864, i_8_1867, i_8_1894, i_8_1951, i_8_1962, i_8_1965, i_8_1978, i_8_2013, i_8_2112, i_8_2131, i_8_2132, i_8_2146, i_8_2152, i_8_2194, i_8_2231, i_8_2239, i_8_2240, o_8_84);
	kernel_8_85 k_8_85(i_8_14, i_8_24, i_8_26, i_8_76, i_8_78, i_8_86, i_8_121, i_8_140, i_8_187, i_8_189, i_8_196, i_8_229, i_8_238, i_8_295, i_8_303, i_8_327, i_8_348, i_8_383, i_8_385, i_8_386, i_8_401, i_8_420, i_8_447, i_8_465, i_8_525, i_8_528, i_8_574, i_8_609, i_8_610, i_8_611, i_8_638, i_8_661, i_8_798, i_8_872, i_8_877, i_8_956, i_8_970, i_8_1006, i_8_1034, i_8_1102, i_8_1120, i_8_1123, i_8_1132, i_8_1159, i_8_1188, i_8_1192, i_8_1194, i_8_1197, i_8_1221, i_8_1237, i_8_1266, i_8_1285, i_8_1328, i_8_1330, i_8_1398, i_8_1422, i_8_1455, i_8_1456, i_8_1468, i_8_1469, i_8_1475, i_8_1493, i_8_1504, i_8_1509, i_8_1510, i_8_1542, i_8_1545, i_8_1546, i_8_1590, i_8_1600, i_8_1617, i_8_1618, i_8_1639, i_8_1640, i_8_1711, i_8_1750, i_8_1751, i_8_1816, i_8_1842, i_8_1843, i_8_1876, i_8_1877, i_8_1888, i_8_1894, i_8_1896, i_8_1905, i_8_1949, i_8_1988, i_8_1995, i_8_2041, i_8_2057, i_8_2112, i_8_2130, i_8_2135, i_8_2149, i_8_2156, i_8_2185, i_8_2193, i_8_2267, i_8_2274, o_8_85);
	kernel_8_86 k_8_86(i_8_7, i_8_40, i_8_64, i_8_76, i_8_79, i_8_139, i_8_150, i_8_151, i_8_190, i_8_214, i_8_230, i_8_304, i_8_322, i_8_364, i_8_376, i_8_394, i_8_395, i_8_400, i_8_401, i_8_420, i_8_421, i_8_422, i_8_446, i_8_479, i_8_482, i_8_483, i_8_485, i_8_490, i_8_526, i_8_530, i_8_570, i_8_574, i_8_592, i_8_593, i_8_594, i_8_596, i_8_602, i_8_611, i_8_639, i_8_642, i_8_705, i_8_715, i_8_728, i_8_751, i_8_762, i_8_814, i_8_827, i_8_843, i_8_844, i_8_845, i_8_859, i_8_886, i_8_895, i_8_899, i_8_925, i_8_1012, i_8_1027, i_8_1076, i_8_1101, i_8_1120, i_8_1229, i_8_1240, i_8_1271, i_8_1305, i_8_1308, i_8_1326, i_8_1328, i_8_1331, i_8_1335, i_8_1357, i_8_1416, i_8_1436, i_8_1437, i_8_1455, i_8_1465, i_8_1472, i_8_1480, i_8_1483, i_8_1547, i_8_1551, i_8_1573, i_8_1634, i_8_1636, i_8_1645, i_8_1654, i_8_1687, i_8_1707, i_8_1708, i_8_1723, i_8_1751, i_8_1754, i_8_1772, i_8_1808, i_8_1858, i_8_1912, i_8_1966, i_8_1996, i_8_2051, i_8_2152, i_8_2214, o_8_86);
	kernel_8_87 k_8_87(i_8_19, i_8_22, i_8_23, i_8_41, i_8_73, i_8_74, i_8_84, i_8_103, i_8_167, i_8_198, i_8_199, i_8_271, i_8_272, i_8_352, i_8_371, i_8_382, i_8_388, i_8_452, i_8_526, i_8_532, i_8_549, i_8_553, i_8_594, i_8_630, i_8_631, i_8_653, i_8_657, i_8_685, i_8_694, i_8_695, i_8_747, i_8_819, i_8_829, i_8_838, i_8_860, i_8_875, i_8_910, i_8_914, i_8_919, i_8_1029, i_8_1110, i_8_1111, i_8_1156, i_8_1198, i_8_1225, i_8_1233, i_8_1234, i_8_1268, i_8_1296, i_8_1297, i_8_1315, i_8_1318, i_8_1332, i_8_1354, i_8_1387, i_8_1390, i_8_1435, i_8_1458, i_8_1471, i_8_1477, i_8_1486, i_8_1530, i_8_1534, i_8_1540, i_8_1547, i_8_1548, i_8_1594, i_8_1595, i_8_1630, i_8_1631, i_8_1633, i_8_1639, i_8_1649, i_8_1657, i_8_1773, i_8_1782, i_8_1784, i_8_1791, i_8_1793, i_8_1818, i_8_1865, i_8_1873, i_8_1886, i_8_1909, i_8_1918, i_8_1944, i_8_1947, i_8_1964, i_8_1972, i_8_1980, i_8_2007, i_8_2063, i_8_2093, i_8_2107, i_8_2147, i_8_2157, i_8_2223, i_8_2233, i_8_2243, i_8_2287, o_8_87);
	kernel_8_88 k_8_88(i_8_93, i_8_94, i_8_107, i_8_143, i_8_197, i_8_223, i_8_266, i_8_283, i_8_284, i_8_288, i_8_296, i_8_299, i_8_305, i_8_319, i_8_322, i_8_328, i_8_368, i_8_382, i_8_404, i_8_431, i_8_437, i_8_489, i_8_492, i_8_553, i_8_557, i_8_593, i_8_599, i_8_628, i_8_637, i_8_643, i_8_656, i_8_661, i_8_664, i_8_724, i_8_727, i_8_781, i_8_782, i_8_790, i_8_791, i_8_824, i_8_827, i_8_840, i_8_843, i_8_845, i_8_930, i_8_931, i_8_953, i_8_976, i_8_991, i_8_1056, i_8_1075, i_8_1155, i_8_1157, i_8_1214, i_8_1240, i_8_1273, i_8_1283, i_8_1324, i_8_1345, i_8_1354, i_8_1366, i_8_1375, i_8_1390, i_8_1391, i_8_1454, i_8_1483, i_8_1490, i_8_1592, i_8_1647, i_8_1681, i_8_1751, i_8_1771, i_8_1789, i_8_1803, i_8_1806, i_8_1810, i_8_1837, i_8_1853, i_8_1859, i_8_1893, i_8_1903, i_8_1907, i_8_1949, i_8_1950, i_8_1994, i_8_1995, i_8_2046, i_8_2120, i_8_2129, i_8_2132, i_8_2150, i_8_2174, i_8_2177, i_8_2194, i_8_2195, i_8_2227, i_8_2248, i_8_2249, i_8_2282, i_8_2287, o_8_88);
	kernel_8_89 k_8_89(i_8_23, i_8_34, i_8_35, i_8_96, i_8_106, i_8_141, i_8_142, i_8_160, i_8_161, i_8_187, i_8_201, i_8_204, i_8_206, i_8_220, i_8_257, i_8_289, i_8_302, i_8_305, i_8_328, i_8_345, i_8_346, i_8_367, i_8_373, i_8_440, i_8_458, i_8_463, i_8_610, i_8_615, i_8_617, i_8_628, i_8_697, i_8_782, i_8_984, i_8_985, i_8_991, i_8_992, i_8_993, i_8_994, i_8_1014, i_8_1087, i_8_1112, i_8_1114, i_8_1135, i_8_1136, i_8_1138, i_8_1189, i_8_1192, i_8_1270, i_8_1271, i_8_1273, i_8_1306, i_8_1344, i_8_1397, i_8_1417, i_8_1434, i_8_1436, i_8_1438, i_8_1511, i_8_1537, i_8_1541, i_8_1542, i_8_1544, i_8_1564, i_8_1578, i_8_1612, i_8_1616, i_8_1629, i_8_1631, i_8_1714, i_8_1715, i_8_1723, i_8_1726, i_8_1727, i_8_1736, i_8_1801, i_8_1804, i_8_1807, i_8_1810, i_8_1812, i_8_1831, i_8_1838, i_8_1840, i_8_1841, i_8_1858, i_8_1922, i_8_2002, i_8_2015, i_8_2049, i_8_2050, i_8_2051, i_8_2134, i_8_2150, i_8_2182, i_8_2215, i_8_2230, i_8_2260, i_8_2261, i_8_2264, i_8_2272, i_8_2282, o_8_89);
	kernel_8_90 k_8_90(i_8_11, i_8_40, i_8_48, i_8_57, i_8_88, i_8_115, i_8_120, i_8_127, i_8_138, i_8_146, i_8_165, i_8_191, i_8_203, i_8_226, i_8_228, i_8_236, i_8_283, i_8_285, i_8_295, i_8_321, i_8_328, i_8_331, i_8_336, i_8_363, i_8_373, i_8_383, i_8_386, i_8_398, i_8_403, i_8_420, i_8_453, i_8_526, i_8_555, i_8_571, i_8_609, i_8_627, i_8_654, i_8_662, i_8_665, i_8_696, i_8_700, i_8_739, i_8_771, i_8_779, i_8_788, i_8_794, i_8_857, i_8_917, i_8_966, i_8_1059, i_8_1068, i_8_1118, i_8_1138, i_8_1235, i_8_1238, i_8_1253, i_8_1300, i_8_1319, i_8_1324, i_8_1353, i_8_1357, i_8_1408, i_8_1451, i_8_1455, i_8_1473, i_8_1534, i_8_1545, i_8_1547, i_8_1605, i_8_1606, i_8_1617, i_8_1623, i_8_1635, i_8_1649, i_8_1669, i_8_1708, i_8_1731, i_8_1732, i_8_1739, i_8_1770, i_8_1784, i_8_1830, i_8_1867, i_8_1886, i_8_1969, i_8_1983, i_8_2118, i_8_2127, i_8_2145, i_8_2149, i_8_2208, i_8_2211, i_8_2212, i_8_2218, i_8_2229, i_8_2238, i_8_2244, i_8_2245, i_8_2247, i_8_2248, o_8_90);
	kernel_8_91 k_8_91(i_8_22, i_8_25, i_8_28, i_8_63, i_8_67, i_8_80, i_8_144, i_8_172, i_8_303, i_8_318, i_8_351, i_8_352, i_8_360, i_8_364, i_8_379, i_8_401, i_8_421, i_8_441, i_8_513, i_8_514, i_8_522, i_8_557, i_8_571, i_8_631, i_8_644, i_8_657, i_8_666, i_8_667, i_8_676, i_8_697, i_8_702, i_8_703, i_8_766, i_8_824, i_8_846, i_8_880, i_8_949, i_8_955, i_8_956, i_8_1047, i_8_1057, i_8_1107, i_8_1115, i_8_1170, i_8_1180, i_8_1201, i_8_1228, i_8_1231, i_8_1269, i_8_1270, i_8_1296, i_8_1351, i_8_1353, i_8_1355, i_8_1386, i_8_1396, i_8_1404, i_8_1408, i_8_1434, i_8_1462, i_8_1463, i_8_1467, i_8_1494, i_8_1497, i_8_1535, i_8_1562, i_8_1631, i_8_1632, i_8_1634, i_8_1656, i_8_1701, i_8_1702, i_8_1746, i_8_1767, i_8_1768, i_8_1769, i_8_1780, i_8_1791, i_8_1794, i_8_1809, i_8_1822, i_8_1831, i_8_1845, i_8_1849, i_8_1863, i_8_1867, i_8_1872, i_8_1901, i_8_1944, i_8_1993, i_8_2034, i_8_2043, i_8_2065, i_8_2089, i_8_2135, i_8_2142, i_8_2147, i_8_2223, i_8_2226, i_8_2274, o_8_91);
	kernel_8_92 k_8_92(i_8_77, i_8_80, i_8_119, i_8_163, i_8_220, i_8_314, i_8_363, i_8_364, i_8_366, i_8_367, i_8_370, i_8_381, i_8_484, i_8_487, i_8_489, i_8_490, i_8_492, i_8_493, i_8_494, i_8_507, i_8_509, i_8_523, i_8_524, i_8_527, i_8_554, i_8_556, i_8_597, i_8_604, i_8_637, i_8_638, i_8_691, i_8_693, i_8_694, i_8_695, i_8_698, i_8_699, i_8_760, i_8_827, i_8_838, i_8_841, i_8_843, i_8_851, i_8_880, i_8_964, i_8_1027, i_8_1072, i_8_1110, i_8_1113, i_8_1255, i_8_1263, i_8_1265, i_8_1296, i_8_1301, i_8_1339, i_8_1355, i_8_1369, i_8_1370, i_8_1372, i_8_1373, i_8_1398, i_8_1399, i_8_1400, i_8_1437, i_8_1438, i_8_1439, i_8_1455, i_8_1468, i_8_1535, i_8_1620, i_8_1621, i_8_1623, i_8_1624, i_8_1625, i_8_1628, i_8_1629, i_8_1632, i_8_1634, i_8_1672, i_8_1693, i_8_1733, i_8_1746, i_8_1747, i_8_1748, i_8_1749, i_8_1752, i_8_1753, i_8_1763, i_8_1825, i_8_1826, i_8_1854, i_8_1861, i_8_1888, i_8_1900, i_8_1904, i_8_1945, i_8_1996, i_8_2171, i_8_2241, i_8_2246, i_8_2276, o_8_92);
	kernel_8_93 k_8_93(i_8_22, i_8_23, i_8_31, i_8_70, i_8_140, i_8_188, i_8_202, i_8_223, i_8_224, i_8_275, i_8_292, i_8_293, i_8_301, i_8_345, i_8_346, i_8_364, i_8_374, i_8_377, i_8_379, i_8_390, i_8_451, i_8_484, i_8_507, i_8_555, i_8_556, i_8_577, i_8_589, i_8_599, i_8_634, i_8_636, i_8_672, i_8_711, i_8_715, i_8_716, i_8_772, i_8_786, i_8_826, i_8_839, i_8_840, i_8_872, i_8_881, i_8_985, i_8_994, i_8_1029, i_8_1119, i_8_1120, i_8_1121, i_8_1124, i_8_1186, i_8_1192, i_8_1219, i_8_1220, i_8_1236, i_8_1256, i_8_1271, i_8_1274, i_8_1283, i_8_1299, i_8_1305, i_8_1306, i_8_1314, i_8_1328, i_8_1329, i_8_1331, i_8_1410, i_8_1467, i_8_1470, i_8_1478, i_8_1497, i_8_1506, i_8_1507, i_8_1508, i_8_1542, i_8_1573, i_8_1615, i_8_1653, i_8_1654, i_8_1669, i_8_1742, i_8_1752, i_8_1763, i_8_1788, i_8_1789, i_8_1790, i_8_1832, i_8_1857, i_8_1858, i_8_1859, i_8_1885, i_8_1985, i_8_2047, i_8_2137, i_8_2153, i_8_2214, i_8_2215, i_8_2216, i_8_2226, i_8_2249, i_8_2261, i_8_2273, o_8_93);
	kernel_8_94 k_8_94(i_8_13, i_8_43, i_8_115, i_8_139, i_8_143, i_8_152, i_8_153, i_8_201, i_8_226, i_8_233, i_8_356, i_8_382, i_8_392, i_8_455, i_8_458, i_8_522, i_8_526, i_8_572, i_8_591, i_8_592, i_8_595, i_8_596, i_8_635, i_8_652, i_8_656, i_8_659, i_8_661, i_8_671, i_8_688, i_8_706, i_8_733, i_8_759, i_8_760, i_8_838, i_8_860, i_8_923, i_8_959, i_8_1013, i_8_1032, i_8_1115, i_8_1156, i_8_1174, i_8_1188, i_8_1229, i_8_1232, i_8_1267, i_8_1268, i_8_1271, i_8_1297, i_8_1300, i_8_1305, i_8_1306, i_8_1307, i_8_1309, i_8_1331, i_8_1385, i_8_1390, i_8_1400, i_8_1438, i_8_1469, i_8_1470, i_8_1471, i_8_1478, i_8_1498, i_8_1531, i_8_1534, i_8_1535, i_8_1544, i_8_1645, i_8_1651, i_8_1679, i_8_1697, i_8_1706, i_8_1778, i_8_1798, i_8_1806, i_8_1807, i_8_1822, i_8_1823, i_8_1826, i_8_1868, i_8_1874, i_8_1883, i_8_1884, i_8_1886, i_8_1916, i_8_1960, i_8_1975, i_8_1992, i_8_2030, i_8_2041, i_8_2066, i_8_2120, i_8_2155, i_8_2173, i_8_2216, i_8_2230, i_8_2243, i_8_2248, i_8_2296, o_8_94);
	kernel_8_95 k_8_95(i_8_3, i_8_7, i_8_22, i_8_124, i_8_170, i_8_200, i_8_250, i_8_287, i_8_292, i_8_293, i_8_328, i_8_329, i_8_330, i_8_366, i_8_383, i_8_385, i_8_440, i_8_456, i_8_493, i_8_529, i_8_554, i_8_584, i_8_626, i_8_635, i_8_642, i_8_673, i_8_674, i_8_680, i_8_695, i_8_700, i_8_701, i_8_703, i_8_704, i_8_763, i_8_809, i_8_827, i_8_833, i_8_836, i_8_844, i_8_852, i_8_854, i_8_958, i_8_968, i_8_971, i_8_986, i_8_989, i_8_1154, i_8_1194, i_8_1227, i_8_1258, i_8_1259, i_8_1267, i_8_1270, i_8_1286, i_8_1299, i_8_1323, i_8_1350, i_8_1358, i_8_1436, i_8_1442, i_8_1468, i_8_1489, i_8_1493, i_8_1520, i_8_1538, i_8_1547, i_8_1574, i_8_1585, i_8_1588, i_8_1591, i_8_1650, i_8_1652, i_8_1675, i_8_1705, i_8_1724, i_8_1750, i_8_1769, i_8_1777, i_8_1781, i_8_1817, i_8_1820, i_8_1824, i_8_1834, i_8_1843, i_8_1860, i_8_1885, i_8_1892, i_8_1896, i_8_2032, i_8_2041, i_8_2042, i_8_2089, i_8_2146, i_8_2149, i_8_2155, i_8_2187, i_8_2191, i_8_2192, i_8_2244, i_8_2275, o_8_95);
	kernel_8_96 k_8_96(i_8_23, i_8_35, i_8_53, i_8_57, i_8_62, i_8_74, i_8_98, i_8_141, i_8_158, i_8_187, i_8_223, i_8_260, i_8_304, i_8_305, i_8_311, i_8_348, i_8_349, i_8_421, i_8_422, i_8_524, i_8_527, i_8_530, i_8_590, i_8_602, i_8_610, i_8_625, i_8_631, i_8_632, i_8_634, i_8_635, i_8_659, i_8_662, i_8_663, i_8_690, i_8_691, i_8_715, i_8_770, i_8_789, i_8_814, i_8_817, i_8_839, i_8_853, i_8_854, i_8_876, i_8_880, i_8_964, i_8_994, i_8_1016, i_8_1018, i_8_1032, i_8_1034, i_8_1052, i_8_1076, i_8_1129, i_8_1193, i_8_1264, i_8_1277, i_8_1299, i_8_1305, i_8_1327, i_8_1328, i_8_1331, i_8_1344, i_8_1346, i_8_1397, i_8_1411, i_8_1434, i_8_1438, i_8_1506, i_8_1507, i_8_1545, i_8_1546, i_8_1565, i_8_1574, i_8_1603, i_8_1624, i_8_1648, i_8_1654, i_8_1720, i_8_1723, i_8_1736, i_8_1742, i_8_1806, i_8_1808, i_8_1844, i_8_1888, i_8_1905, i_8_1906, i_8_1919, i_8_2017, i_8_2032, i_8_2072, i_8_2093, i_8_2134, i_8_2157, i_8_2165, i_8_2216, i_8_2239, i_8_2291, i_8_2292, o_8_96);
	kernel_8_97 k_8_97(i_8_60, i_8_61, i_8_69, i_8_70, i_8_115, i_8_132, i_8_171, i_8_186, i_8_189, i_8_190, i_8_213, i_8_214, i_8_295, i_8_296, i_8_303, i_8_304, i_8_339, i_8_378, i_8_382, i_8_420, i_8_456, i_8_469, i_8_492, i_8_582, i_8_591, i_8_606, i_8_619, i_8_633, i_8_637, i_8_658, i_8_665, i_8_753, i_8_898, i_8_924, i_8_1015, i_8_1073, i_8_1102, i_8_1105, i_8_1131, i_8_1141, i_8_1156, i_8_1176, i_8_1263, i_8_1267, i_8_1284, i_8_1286, i_8_1288, i_8_1304, i_8_1308, i_8_1332, i_8_1353, i_8_1356, i_8_1383, i_8_1402, i_8_1410, i_8_1482, i_8_1484, i_8_1528, i_8_1555, i_8_1591, i_8_1645, i_8_1671, i_8_1672, i_8_1673, i_8_1677, i_8_1681, i_8_1689, i_8_1707, i_8_1713, i_8_1714, i_8_1731, i_8_1732, i_8_1734, i_8_1746, i_8_1754, i_8_1762, i_8_1773, i_8_1779, i_8_1821, i_8_1843, i_8_1857, i_8_1860, i_8_1887, i_8_1888, i_8_1895, i_8_1942, i_8_1966, i_8_1986, i_8_1996, i_8_1997, i_8_2004, i_8_2014, i_8_2076, i_8_2149, i_8_2151, i_8_2173, i_8_2242, i_8_2250, i_8_2275, i_8_2292, o_8_97);
	kernel_8_98 k_8_98(i_8_12, i_8_52, i_8_70, i_8_115, i_8_139, i_8_141, i_8_228, i_8_230, i_8_231, i_8_314, i_8_319, i_8_334, i_8_342, i_8_345, i_8_363, i_8_366, i_8_384, i_8_400, i_8_420, i_8_430, i_8_504, i_8_525, i_8_538, i_8_553, i_8_557, i_8_570, i_8_571, i_8_581, i_8_583, i_8_588, i_8_600, i_8_601, i_8_603, i_8_628, i_8_634, i_8_651, i_8_657, i_8_696, i_8_700, i_8_704, i_8_732, i_8_777, i_8_781, i_8_819, i_8_831, i_8_840, i_8_842, i_8_843, i_8_875, i_8_877, i_8_879, i_8_895, i_8_947, i_8_993, i_8_1003, i_8_1105, i_8_1109, i_8_1115, i_8_1124, i_8_1156, i_8_1267, i_8_1282, i_8_1284, i_8_1315, i_8_1317, i_8_1320, i_8_1347, i_8_1354, i_8_1358, i_8_1366, i_8_1423, i_8_1426, i_8_1453, i_8_1462, i_8_1490, i_8_1509, i_8_1519, i_8_1524, i_8_1551, i_8_1633, i_8_1635, i_8_1680, i_8_1686, i_8_1690, i_8_1695, i_8_1699, i_8_1700, i_8_1703, i_8_1723, i_8_1770, i_8_1780, i_8_1884, i_8_1911, i_8_1956, i_8_1995, i_8_2132, i_8_2137, i_8_2151, i_8_2240, i_8_2275, o_8_98);
	kernel_8_99 k_8_99(i_8_13, i_8_34, i_8_35, i_8_57, i_8_67, i_8_97, i_8_127, i_8_129, i_8_255, i_8_299, i_8_310, i_8_344, i_8_364, i_8_365, i_8_422, i_8_423, i_8_480, i_8_483, i_8_517, i_8_523, i_8_528, i_8_530, i_8_545, i_8_571, i_8_580, i_8_607, i_8_608, i_8_631, i_8_649, i_8_679, i_8_680, i_8_705, i_8_707, i_8_799, i_8_826, i_8_839, i_8_857, i_8_866, i_8_964, i_8_993, i_8_994, i_8_1013, i_8_1050, i_8_1065, i_8_1110, i_8_1111, i_8_1153, i_8_1202, i_8_1237, i_8_1246, i_8_1267, i_8_1270, i_8_1305, i_8_1306, i_8_1307, i_8_1318, i_8_1324, i_8_1399, i_8_1423, i_8_1424, i_8_1437, i_8_1471, i_8_1472, i_8_1486, i_8_1525, i_8_1573, i_8_1574, i_8_1624, i_8_1630, i_8_1632, i_8_1673, i_8_1687, i_8_1705, i_8_1707, i_8_1743, i_8_1768, i_8_1784, i_8_1793, i_8_1795, i_8_1819, i_8_1820, i_8_1935, i_8_1937, i_8_1975, i_8_1995, i_8_2089, i_8_2090, i_8_2101, i_8_2104, i_8_2129, i_8_2145, i_8_2149, i_8_2156, i_8_2214, i_8_2216, i_8_2224, i_8_2225, i_8_2233, i_8_2245, i_8_2248, o_8_99);
	kernel_8_100 k_8_100(i_8_48, i_8_50, i_8_111, i_8_165, i_8_187, i_8_226, i_8_231, i_8_256, i_8_367, i_8_373, i_8_391, i_8_415, i_8_433, i_8_444, i_8_481, i_8_490, i_8_493, i_8_504, i_8_507, i_8_549, i_8_552, i_8_553, i_8_554, i_8_599, i_8_602, i_8_630, i_8_659, i_8_692, i_8_715, i_8_778, i_8_781, i_8_782, i_8_786, i_8_804, i_8_816, i_8_841, i_8_850, i_8_931, i_8_1047, i_8_1050, i_8_1051, i_8_1104, i_8_1110, i_8_1111, i_8_1120, i_8_1140, i_8_1162, i_8_1185, i_8_1236, i_8_1265, i_8_1270, i_8_1281, i_8_1282, i_8_1283, i_8_1285, i_8_1286, i_8_1306, i_8_1307, i_8_1327, i_8_1331, i_8_1390, i_8_1396, i_8_1404, i_8_1405, i_8_1407, i_8_1438, i_8_1506, i_8_1509, i_8_1536, i_8_1561, i_8_1590, i_8_1641, i_8_1649, i_8_1650, i_8_1719, i_8_1722, i_8_1724, i_8_1741, i_8_1846, i_8_1856, i_8_1857, i_8_1858, i_8_1866, i_8_1873, i_8_1884, i_8_1903, i_8_1904, i_8_1956, i_8_1958, i_8_2010, i_8_2016, i_8_2127, i_8_2140, i_8_2173, i_8_2214, i_8_2215, i_8_2216, i_8_2236, i_8_2261, i_8_2299, o_8_100);
	kernel_8_101 k_8_101(i_8_1, i_8_5, i_8_53, i_8_65, i_8_75, i_8_167, i_8_185, i_8_200, i_8_217, i_8_221, i_8_226, i_8_227, i_8_262, i_8_266, i_8_343, i_8_360, i_8_363, i_8_364, i_8_398, i_8_424, i_8_425, i_8_452, i_8_454, i_8_490, i_8_493, i_8_505, i_8_525, i_8_581, i_8_584, i_8_587, i_8_608, i_8_611, i_8_624, i_8_640, i_8_696, i_8_724, i_8_730, i_8_731, i_8_803, i_8_806, i_8_809, i_8_873, i_8_883, i_8_935, i_8_956, i_8_963, i_8_968, i_8_980, i_8_992, i_8_995, i_8_1073, i_8_1075, i_8_1076, i_8_1114, i_8_1127, i_8_1171, i_8_1229, i_8_1234, i_8_1238, i_8_1259, i_8_1274, i_8_1289, i_8_1298, i_8_1325, i_8_1355, i_8_1382, i_8_1385, i_8_1391, i_8_1441, i_8_1487, i_8_1492, i_8_1628, i_8_1636, i_8_1691, i_8_1703, i_8_1752, i_8_1759, i_8_1778, i_8_1792, i_8_1793, i_8_1823, i_8_1847, i_8_1850, i_8_1882, i_8_1909, i_8_1910, i_8_1980, i_8_1981, i_8_1982, i_8_1994, i_8_2018, i_8_2078, i_8_2099, i_8_2139, i_8_2140, i_8_2144, i_8_2147, i_8_2172, i_8_2213, i_8_2297, o_8_101);
	kernel_8_102 k_8_102(i_8_28, i_8_32, i_8_35, i_8_89, i_8_157, i_8_169, i_8_224, i_8_283, i_8_292, i_8_355, i_8_437, i_8_455, i_8_480, i_8_529, i_8_544, i_8_552, i_8_557, i_8_609, i_8_617, i_8_658, i_8_659, i_8_663, i_8_665, i_8_703, i_8_718, i_8_769, i_8_772, i_8_850, i_8_881, i_8_890, i_8_896, i_8_951, i_8_955, i_8_973, i_8_977, i_8_1013, i_8_1032, i_8_1048, i_8_1050, i_8_1066, i_8_1075, i_8_1084, i_8_1135, i_8_1137, i_8_1154, i_8_1157, i_8_1223, i_8_1246, i_8_1247, i_8_1249, i_8_1256, i_8_1258, i_8_1259, i_8_1265, i_8_1282, i_8_1283, i_8_1285, i_8_1297, i_8_1346, i_8_1350, i_8_1367, i_8_1436, i_8_1449, i_8_1453, i_8_1467, i_8_1468, i_8_1471, i_8_1482, i_8_1501, i_8_1502, i_8_1532, i_8_1549, i_8_1577, i_8_1580, i_8_1613, i_8_1679, i_8_1718, i_8_1731, i_8_1760, i_8_1771, i_8_1772, i_8_1776, i_8_1787, i_8_1855, i_8_1856, i_8_1928, i_8_1931, i_8_1948, i_8_1951, i_8_1960, i_8_2000, i_8_2030, i_8_2084, i_8_2143, i_8_2171, i_8_2179, i_8_2214, i_8_2263, i_8_2264, i_8_2290, o_8_102);
	kernel_8_103 k_8_103(i_8_23, i_8_26, i_8_33, i_8_34, i_8_35, i_8_61, i_8_73, i_8_87, i_8_114, i_8_168, i_8_189, i_8_190, i_8_223, i_8_240, i_8_241, i_8_340, i_8_375, i_8_437, i_8_469, i_8_470, i_8_483, i_8_484, i_8_525, i_8_527, i_8_574, i_8_575, i_8_602, i_8_619, i_8_636, i_8_637, i_8_679, i_8_690, i_8_691, i_8_763, i_8_781, i_8_826, i_8_861, i_8_889, i_8_934, i_8_943, i_8_944, i_8_970, i_8_994, i_8_995, i_8_1059, i_8_1060, i_8_1074, i_8_1111, i_8_1114, i_8_1185, i_8_1191, i_8_1260, i_8_1284, i_8_1285, i_8_1295, i_8_1303, i_8_1304, i_8_1305, i_8_1306, i_8_1339, i_8_1439, i_8_1492, i_8_1536, i_8_1564, i_8_1575, i_8_1576, i_8_1591, i_8_1647, i_8_1650, i_8_1653, i_8_1681, i_8_1699, i_8_1700, i_8_1723, i_8_1742, i_8_1743, i_8_1744, i_8_1745, i_8_1753, i_8_1762, i_8_1763, i_8_1780, i_8_1781, i_8_1834, i_8_1844, i_8_1885, i_8_1887, i_8_1889, i_8_2050, i_8_2059, i_8_2060, i_8_2074, i_8_2076, i_8_2123, i_8_2176, i_8_2218, i_8_2219, i_8_2220, i_8_2247, i_8_2302, o_8_103);
	kernel_8_104 k_8_104(i_8_12, i_8_63, i_8_72, i_8_73, i_8_84, i_8_181, i_8_298, i_8_301, i_8_318, i_8_319, i_8_334, i_8_343, i_8_361, i_8_387, i_8_418, i_8_469, i_8_492, i_8_504, i_8_505, i_8_523, i_8_540, i_8_558, i_8_577, i_8_579, i_8_588, i_8_603, i_8_630, i_8_640, i_8_651, i_8_652, i_8_657, i_8_660, i_8_678, i_8_687, i_8_707, i_8_757, i_8_819, i_8_823, i_8_839, i_8_842, i_8_856, i_8_882, i_8_886, i_8_941, i_8_954, i_8_969, i_8_1012, i_8_1026, i_8_1056, i_8_1071, i_8_1135, i_8_1153, i_8_1170, i_8_1197, i_8_1215, i_8_1225, i_8_1238, i_8_1261, i_8_1294, i_8_1381, i_8_1395, i_8_1398, i_8_1423, i_8_1479, i_8_1487, i_8_1506, i_8_1507, i_8_1512, i_8_1557, i_8_1570, i_8_1630, i_8_1654, i_8_1668, i_8_1671, i_8_1681, i_8_1728, i_8_1747, i_8_1794, i_8_1824, i_8_1825, i_8_1866, i_8_1918, i_8_1948, i_8_1962, i_8_1963, i_8_1989, i_8_1992, i_8_1997, i_8_2103, i_8_2106, i_8_2107, i_8_2115, i_8_2145, i_8_2149, i_8_2151, i_8_2152, i_8_2162, i_8_2190, i_8_2232, i_8_2245, o_8_104);
	kernel_8_105 k_8_105(i_8_32, i_8_33, i_8_141, i_8_142, i_8_146, i_8_189, i_8_196, i_8_318, i_8_358, i_8_393, i_8_399, i_8_421, i_8_462, i_8_502, i_8_516, i_8_524, i_8_594, i_8_597, i_8_604, i_8_624, i_8_679, i_8_702, i_8_782, i_8_789, i_8_811, i_8_834, i_8_867, i_8_941, i_8_970, i_8_993, i_8_1012, i_8_1014, i_8_1075, i_8_1108, i_8_1110, i_8_1128, i_8_1137, i_8_1167, i_8_1172, i_8_1230, i_8_1246, i_8_1272, i_8_1278, i_8_1300, i_8_1301, i_8_1306, i_8_1318, i_8_1326, i_8_1331, i_8_1337, i_8_1338, i_8_1355, i_8_1356, i_8_1411, i_8_1426, i_8_1437, i_8_1467, i_8_1480, i_8_1534, i_8_1546, i_8_1552, i_8_1596, i_8_1597, i_8_1642, i_8_1644, i_8_1645, i_8_1650, i_8_1672, i_8_1707, i_8_1721, i_8_1749, i_8_1785, i_8_1795, i_8_1800, i_8_1843, i_8_1852, i_8_1854, i_8_1858, i_8_1875, i_8_1885, i_8_1947, i_8_1974, i_8_1975, i_8_1986, i_8_2047, i_8_2064, i_8_2091, i_8_2094, i_8_2104, i_8_2119, i_8_2123, i_8_2143, i_8_2148, i_8_2150, i_8_2155, i_8_2169, i_8_2214, i_8_2216, i_8_2226, i_8_2244, o_8_105);
	kernel_8_106 k_8_106(i_8_34, i_8_71, i_8_80, i_8_88, i_8_107, i_8_115, i_8_194, i_8_228, i_8_241, i_8_242, i_8_278, i_8_304, i_8_379, i_8_381, i_8_385, i_8_424, i_8_484, i_8_489, i_8_490, i_8_492, i_8_523, i_8_529, i_8_610, i_8_634, i_8_637, i_8_658, i_8_682, i_8_694, i_8_706, i_8_715, i_8_717, i_8_723, i_8_735, i_8_738, i_8_798, i_8_799, i_8_817, i_8_853, i_8_880, i_8_994, i_8_1047, i_8_1048, i_8_1057, i_8_1066, i_8_1084, i_8_1105, i_8_1114, i_8_1116, i_8_1117, i_8_1147, i_8_1171, i_8_1225, i_8_1228, i_8_1235, i_8_1236, i_8_1278, i_8_1285, i_8_1288, i_8_1333, i_8_1354, i_8_1357, i_8_1438, i_8_1545, i_8_1552, i_8_1564, i_8_1605, i_8_1609, i_8_1615, i_8_1627, i_8_1646, i_8_1648, i_8_1663, i_8_1696, i_8_1753, i_8_1763, i_8_1771, i_8_1774, i_8_1785, i_8_1786, i_8_1821, i_8_1825, i_8_1843, i_8_1849, i_8_1855, i_8_1860, i_8_1887, i_8_1903, i_8_1914, i_8_1915, i_8_1986, i_8_1987, i_8_1988, i_8_1996, i_8_2041, i_8_2121, i_8_2122, i_8_2149, i_8_2157, i_8_2242, i_8_2292, o_8_106);
	kernel_8_107 k_8_107(i_8_31, i_8_50, i_8_86, i_8_167, i_8_230, i_8_233, i_8_234, i_8_326, i_8_335, i_8_338, i_8_365, i_8_368, i_8_380, i_8_386, i_8_400, i_8_419, i_8_424, i_8_425, i_8_428, i_8_440, i_8_449, i_8_451, i_8_452, i_8_494, i_8_499, i_8_500, i_8_581, i_8_613, i_8_614, i_8_617, i_8_655, i_8_694, i_8_698, i_8_706, i_8_707, i_8_733, i_8_767, i_8_770, i_8_796, i_8_797, i_8_839, i_8_842, i_8_845, i_8_878, i_8_932, i_8_956, i_8_968, i_8_1019, i_8_1022, i_8_1058, i_8_1097, i_8_1106, i_8_1157, i_8_1229, i_8_1235, i_8_1238, i_8_1253, i_8_1256, i_8_1264, i_8_1283, i_8_1292, i_8_1310, i_8_1404, i_8_1547, i_8_1588, i_8_1607, i_8_1628, i_8_1652, i_8_1673, i_8_1681, i_8_1706, i_8_1733, i_8_1763, i_8_1777, i_8_1819, i_8_1823, i_8_1825, i_8_1826, i_8_1858, i_8_1889, i_8_1940, i_8_1996, i_8_2003, i_8_2072, i_8_2108, i_8_2111, i_8_2134, i_8_2147, i_8_2149, i_8_2153, i_8_2156, i_8_2173, i_8_2180, i_8_2192, i_8_2200, i_8_2201, i_8_2225, i_8_2244, i_8_2273, i_8_2294, o_8_107);
	kernel_8_108 k_8_108(i_8_138, i_8_163, i_8_175, i_8_211, i_8_241, i_8_262, i_8_306, i_8_309, i_8_349, i_8_363, i_8_390, i_8_444, i_8_462, i_8_492, i_8_493, i_8_499, i_8_501, i_8_504, i_8_505, i_8_524, i_8_525, i_8_528, i_8_586, i_8_643, i_8_697, i_8_701, i_8_707, i_8_709, i_8_714, i_8_750, i_8_751, i_8_780, i_8_813, i_8_842, i_8_880, i_8_895, i_8_964, i_8_996, i_8_1013, i_8_1035, i_8_1040, i_8_1047, i_8_1071, i_8_1074, i_8_1084, i_8_1110, i_8_1113, i_8_1132, i_8_1157, i_8_1267, i_8_1303, i_8_1317, i_8_1326, i_8_1383, i_8_1401, i_8_1409, i_8_1422, i_8_1423, i_8_1443, i_8_1462, i_8_1465, i_8_1506, i_8_1507, i_8_1519, i_8_1533, i_8_1547, i_8_1548, i_8_1552, i_8_1553, i_8_1603, i_8_1623, i_8_1638, i_8_1672, i_8_1674, i_8_1683, i_8_1693, i_8_1701, i_8_1773, i_8_1775, i_8_1783, i_8_1832, i_8_1839, i_8_1840, i_8_1881, i_8_1882, i_8_1883, i_8_1885, i_8_1886, i_8_1888, i_8_1894, i_8_1900, i_8_1957, i_8_1984, i_8_2075, i_8_2088, i_8_2109, i_8_2148, i_8_2156, i_8_2173, i_8_2197, o_8_108);
	kernel_8_109 k_8_109(i_8_51, i_8_77, i_8_194, i_8_220, i_8_221, i_8_223, i_8_224, i_8_225, i_8_234, i_8_235, i_8_236, i_8_237, i_8_239, i_8_273, i_8_303, i_8_325, i_8_326, i_8_329, i_8_334, i_8_336, i_8_337, i_8_338, i_8_365, i_8_391, i_8_414, i_8_415, i_8_418, i_8_419, i_8_596, i_8_613, i_8_614, i_8_648, i_8_649, i_8_650, i_8_651, i_8_652, i_8_715, i_8_748, i_8_749, i_8_764, i_8_838, i_8_848, i_8_970, i_8_1032, i_8_1048, i_8_1050, i_8_1278, i_8_1287, i_8_1290, i_8_1291, i_8_1292, i_8_1303, i_8_1353, i_8_1355, i_8_1439, i_8_1545, i_8_1546, i_8_1547, i_8_1630, i_8_1631, i_8_1635, i_8_1675, i_8_1746, i_8_1759, i_8_1764, i_8_1767, i_8_1769, i_8_1773, i_8_1774, i_8_1775, i_8_1778, i_8_1808, i_8_1818, i_8_1819, i_8_1820, i_8_1827, i_8_1828, i_8_1829, i_8_1830, i_8_1831, i_8_1859, i_8_1883, i_8_1924, i_8_1949, i_8_1990, i_8_1992, i_8_1993, i_8_1994, i_8_2016, i_8_2017, i_8_2019, i_8_2028, i_8_2088, i_8_2133, i_8_2134, i_8_2152, i_8_2208, i_8_2209, i_8_2223, i_8_2290, o_8_109);
	kernel_8_110 k_8_110(i_8_0, i_8_19, i_8_20, i_8_36, i_8_46, i_8_47, i_8_100, i_8_111, i_8_136, i_8_189, i_8_347, i_8_379, i_8_398, i_8_425, i_8_487, i_8_496, i_8_527, i_8_595, i_8_607, i_8_633, i_8_634, i_8_709, i_8_766, i_8_767, i_8_838, i_8_874, i_8_879, i_8_884, i_8_919, i_8_922, i_8_966, i_8_968, i_8_991, i_8_992, i_8_1026, i_8_1036, i_8_1073, i_8_1135, i_8_1154, i_8_1180, i_8_1225, i_8_1226, i_8_1252, i_8_1253, i_8_1263, i_8_1265, i_8_1270, i_8_1279, i_8_1280, i_8_1399, i_8_1453, i_8_1468, i_8_1478, i_8_1486, i_8_1487, i_8_1493, i_8_1534, i_8_1558, i_8_1559, i_8_1603, i_8_1604, i_8_1634, i_8_1648, i_8_1649, i_8_1681, i_8_1710, i_8_1719, i_8_1746, i_8_1747, i_8_1748, i_8_1764, i_8_1768, i_8_1771, i_8_1779, i_8_1792, i_8_1803, i_8_1832, i_8_1882, i_8_1884, i_8_1886, i_8_1944, i_8_1946, i_8_1981, i_8_1991, i_8_1994, i_8_2008, i_8_2017, i_8_2054, i_8_2090, i_8_2106, i_8_2107, i_8_2108, i_8_2147, i_8_2153, i_8_2224, i_8_2242, i_8_2245, i_8_2270, i_8_2287, i_8_2288, o_8_110);
	kernel_8_111 k_8_111(i_8_10, i_8_37, i_8_49, i_8_76, i_8_107, i_8_189, i_8_223, i_8_253, i_8_301, i_8_361, i_8_363, i_8_365, i_8_389, i_8_398, i_8_426, i_8_440, i_8_490, i_8_526, i_8_532, i_8_577, i_8_580, i_8_589, i_8_590, i_8_604, i_8_607, i_8_631, i_8_632, i_8_633, i_8_634, i_8_665, i_8_671, i_8_676, i_8_680, i_8_738, i_8_740, i_8_805, i_8_824, i_8_832, i_8_837, i_8_838, i_8_839, i_8_955, i_8_965, i_8_1037, i_8_1051, i_8_1099, i_8_1103, i_8_1127, i_8_1136, i_8_1152, i_8_1181, i_8_1237, i_8_1238, i_8_1261, i_8_1262, i_8_1315, i_8_1325, i_8_1328, i_8_1382, i_8_1398, i_8_1407, i_8_1414, i_8_1433, i_8_1434, i_8_1442, i_8_1463, i_8_1470, i_8_1472, i_8_1478, i_8_1506, i_8_1513, i_8_1550, i_8_1624, i_8_1629, i_8_1641, i_8_1702, i_8_1724, i_8_1768, i_8_1784, i_8_1804, i_8_1818, i_8_1820, i_8_1822, i_8_1837, i_8_1839, i_8_1903, i_8_1994, i_8_2008, i_8_2009, i_8_2011, i_8_2038, i_8_2071, i_8_2089, i_8_2098, i_8_2225, i_8_2227, i_8_2244, i_8_2245, i_8_2263, i_8_2296, o_8_111);
	kernel_8_112 k_8_112(i_8_14, i_8_45, i_8_46, i_8_66, i_8_82, i_8_136, i_8_163, i_8_172, i_8_193, i_8_207, i_8_238, i_8_253, i_8_255, i_8_307, i_8_342, i_8_345, i_8_375, i_8_423, i_8_424, i_8_470, i_8_481, i_8_495, i_8_526, i_8_527, i_8_544, i_8_549, i_8_568, i_8_586, i_8_603, i_8_613, i_8_630, i_8_664, i_8_676, i_8_765, i_8_828, i_8_883, i_8_918, i_8_927, i_8_973, i_8_997, i_8_998, i_8_1009, i_8_1017, i_8_1044, i_8_1045, i_8_1053, i_8_1221, i_8_1228, i_8_1233, i_8_1269, i_8_1271, i_8_1288, i_8_1296, i_8_1297, i_8_1306, i_8_1314, i_8_1323, i_8_1413, i_8_1434, i_8_1435, i_8_1512, i_8_1524, i_8_1536, i_8_1541, i_8_1558, i_8_1566, i_8_1611, i_8_1630, i_8_1642, i_8_1648, i_8_1650, i_8_1680, i_8_1681, i_8_1682, i_8_1683, i_8_1695, i_8_1707, i_8_1729, i_8_1763, i_8_1764, i_8_1803, i_8_1822, i_8_1855, i_8_1884, i_8_1885, i_8_1886, i_8_1902, i_8_1998, i_8_2106, i_8_2119, i_8_2142, i_8_2145, i_8_2152, i_8_2154, i_8_2187, i_8_2196, i_8_2205, i_8_2259, i_8_2260, i_8_2269, o_8_112);
	kernel_8_113 k_8_113(i_8_38, i_8_40, i_8_43, i_8_81, i_8_84, i_8_115, i_8_148, i_8_151, i_8_163, i_8_190, i_8_194, i_8_245, i_8_346, i_8_347, i_8_352, i_8_417, i_8_464, i_8_469, i_8_470, i_8_483, i_8_489, i_8_490, i_8_522, i_8_526, i_8_538, i_8_552, i_8_555, i_8_595, i_8_598, i_8_634, i_8_648, i_8_695, i_8_697, i_8_700, i_8_702, i_8_706, i_8_733, i_8_734, i_8_770, i_8_790, i_8_793, i_8_813, i_8_833, i_8_881, i_8_893, i_8_896, i_8_926, i_8_998, i_8_1154, i_8_1161, i_8_1171, i_8_1223, i_8_1233, i_8_1238, i_8_1262, i_8_1288, i_8_1289, i_8_1292, i_8_1299, i_8_1306, i_8_1309, i_8_1311, i_8_1312, i_8_1352, i_8_1381, i_8_1384, i_8_1423, i_8_1442, i_8_1491, i_8_1498, i_8_1543, i_8_1549, i_8_1562, i_8_1637, i_8_1648, i_8_1653, i_8_1687, i_8_1688, i_8_1690, i_8_1701, i_8_1708, i_8_1748, i_8_1750, i_8_1753, i_8_1803, i_8_1806, i_8_1832, i_8_1840, i_8_1926, i_8_1960, i_8_1996, i_8_2038, i_8_2107, i_8_2203, i_8_2214, i_8_2217, i_8_2227, i_8_2273, i_8_2286, i_8_2290, o_8_113);
	kernel_8_114 k_8_114(i_8_16, i_8_17, i_8_43, i_8_67, i_8_68, i_8_115, i_8_143, i_8_187, i_8_223, i_8_301, i_8_322, i_8_363, i_8_366, i_8_367, i_8_368, i_8_382, i_8_403, i_8_416, i_8_430, i_8_475, i_8_476, i_8_511, i_8_529, i_8_539, i_8_592, i_8_603, i_8_606, i_8_608, i_8_609, i_8_610, i_8_611, i_8_634, i_8_637, i_8_643, i_8_655, i_8_660, i_8_664, i_8_682, i_8_840, i_8_842, i_8_843, i_8_844, i_8_845, i_8_881, i_8_895, i_8_970, i_8_977, i_8_1039, i_8_1106, i_8_1137, i_8_1184, i_8_1201, i_8_1264, i_8_1267, i_8_1282, i_8_1283, i_8_1285, i_8_1286, i_8_1301, i_8_1303, i_8_1318, i_8_1331, i_8_1340, i_8_1351, i_8_1366, i_8_1403, i_8_1426, i_8_1438, i_8_1465, i_8_1484, i_8_1493, i_8_1528, i_8_1529, i_8_1552, i_8_1555, i_8_1574, i_8_1649, i_8_1689, i_8_1690, i_8_1692, i_8_1697, i_8_1726, i_8_1771, i_8_1789, i_8_1794, i_8_1808, i_8_1840, i_8_1874, i_8_1885, i_8_1979, i_8_1981, i_8_2092, i_8_2096, i_8_2105, i_8_2173, i_8_2174, i_8_2227, i_8_2247, i_8_2248, i_8_2300, o_8_114);
	kernel_8_115 k_8_115(i_8_49, i_8_57, i_8_75, i_8_77, i_8_87, i_8_122, i_8_165, i_8_166, i_8_170, i_8_204, i_8_223, i_8_229, i_8_241, i_8_345, i_8_347, i_8_377, i_8_426, i_8_454, i_8_455, i_8_458, i_8_476, i_8_508, i_8_608, i_8_615, i_8_617, i_8_618, i_8_619, i_8_633, i_8_634, i_8_638, i_8_657, i_8_658, i_8_660, i_8_662, i_8_664, i_8_695, i_8_795, i_8_806, i_8_839, i_8_851, i_8_877, i_8_878, i_8_880, i_8_896, i_8_958, i_8_1012, i_8_1029, i_8_1030, i_8_1034, i_8_1037, i_8_1045, i_8_1071, i_8_1072, i_8_1076, i_8_1130, i_8_1166, i_8_1226, i_8_1228, i_8_1229, i_8_1240, i_8_1263, i_8_1264, i_8_1284, i_8_1293, i_8_1296, i_8_1298, i_8_1300, i_8_1301, i_8_1329, i_8_1453, i_8_1454, i_8_1455, i_8_1457, i_8_1506, i_8_1509, i_8_1510, i_8_1542, i_8_1543, i_8_1544, i_8_1550, i_8_1552, i_8_1607, i_8_1630, i_8_1806, i_8_1862, i_8_1893, i_8_1894, i_8_1895, i_8_1898, i_8_1951, i_8_2041, i_8_2096, i_8_2126, i_8_2128, i_8_2129, i_8_2143, i_8_2217, i_8_2218, i_8_2227, i_8_2273, o_8_115);
	kernel_8_116 k_8_116(i_8_160, i_8_186, i_8_257, i_8_293, i_8_331, i_8_373, i_8_381, i_8_394, i_8_430, i_8_462, i_8_463, i_8_464, i_8_528, i_8_529, i_8_553, i_8_556, i_8_592, i_8_593, i_8_599, i_8_607, i_8_608, i_8_615, i_8_636, i_8_653, i_8_661, i_8_665, i_8_710, i_8_760, i_8_780, i_8_782, i_8_795, i_8_817, i_8_827, i_8_833, i_8_838, i_8_955, i_8_998, i_8_1074, i_8_1078, i_8_1114, i_8_1160, i_8_1191, i_8_1231, i_8_1258, i_8_1285, i_8_1300, i_8_1318, i_8_1331, i_8_1382, i_8_1437, i_8_1438, i_8_1439, i_8_1452, i_8_1453, i_8_1480, i_8_1483, i_8_1506, i_8_1534, i_8_1535, i_8_1542, i_8_1547, i_8_1553, i_8_1562, i_8_1588, i_8_1592, i_8_1605, i_8_1615, i_8_1634, i_8_1715, i_8_1722, i_8_1762, i_8_1789, i_8_1799, i_8_1813, i_8_1822, i_8_1830, i_8_1839, i_8_1841, i_8_1867, i_8_1888, i_8_1893, i_8_1897, i_8_1898, i_8_1900, i_8_1922, i_8_1948, i_8_1965, i_8_1966, i_8_1995, i_8_1996, i_8_2001, i_8_2014, i_8_2109, i_8_2128, i_8_2163, i_8_2203, i_8_2216, i_8_2260, i_8_2264, i_8_2274, o_8_116);
	kernel_8_117 k_8_117(i_8_22, i_8_23, i_8_109, i_8_136, i_8_138, i_8_139, i_8_140, i_8_142, i_8_143, i_8_269, i_8_324, i_8_325, i_8_326, i_8_366, i_8_385, i_8_420, i_8_421, i_8_422, i_8_446, i_8_459, i_8_461, i_8_469, i_8_472, i_8_474, i_8_475, i_8_492, i_8_496, i_8_575, i_8_592, i_8_629, i_8_657, i_8_658, i_8_709, i_8_792, i_8_795, i_8_804, i_8_817, i_8_838, i_8_877, i_8_878, i_8_880, i_8_993, i_8_1078, i_8_1111, i_8_1114, i_8_1159, i_8_1185, i_8_1230, i_8_1279, i_8_1365, i_8_1393, i_8_1410, i_8_1426, i_8_1437, i_8_1471, i_8_1480, i_8_1482, i_8_1524, i_8_1607, i_8_1608, i_8_1609, i_8_1610, i_8_1652, i_8_1655, i_8_1677, i_8_1719, i_8_1724, i_8_1725, i_8_1732, i_8_1736, i_8_1747, i_8_1753, i_8_1787, i_8_1802, i_8_1805, i_8_1806, i_8_1856, i_8_1860, i_8_1886, i_8_1901, i_8_1903, i_8_1904, i_8_1945, i_8_1946, i_8_1948, i_8_1949, i_8_1951, i_8_1964, i_8_1967, i_8_1970, i_8_1992, i_8_2031, i_8_2109, i_8_2112, i_8_2137, i_8_2152, i_8_2153, i_8_2156, i_8_2158, i_8_2226, o_8_117);
	kernel_8_118 k_8_118(i_8_31, i_8_84, i_8_96, i_8_161, i_8_192, i_8_224, i_8_293, i_8_300, i_8_301, i_8_368, i_8_373, i_8_378, i_8_379, i_8_381, i_8_383, i_8_384, i_8_386, i_8_394, i_8_421, i_8_422, i_8_446, i_8_456, i_8_462, i_8_483, i_8_493, i_8_494, i_8_500, i_8_556, i_8_588, i_8_593, i_8_660, i_8_661, i_8_673, i_8_715, i_8_718, i_8_781, i_8_783, i_8_795, i_8_796, i_8_826, i_8_827, i_8_842, i_8_878, i_8_1012, i_8_1029, i_8_1077, i_8_1115, i_8_1120, i_8_1156, i_8_1191, i_8_1228, i_8_1229, i_8_1255, i_8_1274, i_8_1300, i_8_1331, i_8_1345, i_8_1346, i_8_1438, i_8_1457, i_8_1471, i_8_1534, i_8_1535, i_8_1548, i_8_1587, i_8_1597, i_8_1598, i_8_1606, i_8_1648, i_8_1649, i_8_1705, i_8_1751, i_8_1763, i_8_1804, i_8_1807, i_8_1808, i_8_1812, i_8_1822, i_8_1841, i_8_1844, i_8_1894, i_8_1903, i_8_1952, i_8_1966, i_8_2110, i_8_2113, i_8_2127, i_8_2132, i_8_2136, i_8_2139, i_8_2158, i_8_2172, i_8_2182, i_8_2190, i_8_2191, i_8_2195, i_8_2216, i_8_2227, i_8_2273, i_8_2276, o_8_118);
	kernel_8_119 k_8_119(i_8_50, i_8_139, i_8_224, i_8_225, i_8_230, i_8_323, i_8_363, i_8_365, i_8_385, i_8_394, i_8_402, i_8_403, i_8_489, i_8_550, i_8_554, i_8_569, i_8_604, i_8_606, i_8_626, i_8_632, i_8_638, i_8_644, i_8_664, i_8_665, i_8_675, i_8_679, i_8_697, i_8_700, i_8_781, i_8_785, i_8_823, i_8_833, i_8_839, i_8_858, i_8_873, i_8_876, i_8_893, i_8_898, i_8_959, i_8_968, i_8_992, i_8_1034, i_8_1040, i_8_1073, i_8_1094, i_8_1134, i_8_1137, i_8_1150, i_8_1202, i_8_1232, i_8_1264, i_8_1328, i_8_1340, i_8_1349, i_8_1366, i_8_1367, i_8_1372, i_8_1404, i_8_1436, i_8_1451, i_8_1465, i_8_1481, i_8_1490, i_8_1557, i_8_1558, i_8_1573, i_8_1629, i_8_1633, i_8_1634, i_8_1700, i_8_1704, i_8_1705, i_8_1709, i_8_1727, i_8_1733, i_8_1771, i_8_1772, i_8_1824, i_8_1825, i_8_1826, i_8_1884, i_8_1886, i_8_1888, i_8_1939, i_8_1940, i_8_1944, i_8_1960, i_8_1981, i_8_1997, i_8_2142, i_8_2155, i_8_2157, i_8_2225, i_8_2226, i_8_2231, i_8_2241, i_8_2248, i_8_2262, i_8_2282, i_8_2289, o_8_119);
	kernel_8_120 k_8_120(i_8_18, i_8_19, i_8_29, i_8_32, i_8_83, i_8_95, i_8_98, i_8_109, i_8_112, i_8_116, i_8_142, i_8_143, i_8_163, i_8_164, i_8_166, i_8_218, i_8_221, i_8_239, i_8_241, i_8_299, i_8_331, i_8_344, i_8_360, i_8_381, i_8_479, i_8_481, i_8_484, i_8_504, i_8_526, i_8_591, i_8_598, i_8_602, i_8_605, i_8_614, i_8_632, i_8_686, i_8_701, i_8_702, i_8_704, i_8_707, i_8_713, i_8_737, i_8_812, i_8_878, i_8_921, i_8_938, i_8_997, i_8_998, i_8_1012, i_8_1045, i_8_1048, i_8_1058, i_8_1091, i_8_1107, i_8_1117, i_8_1181, i_8_1235, i_8_1262, i_8_1265, i_8_1280, i_8_1282, i_8_1306, i_8_1355, i_8_1412, i_8_1434, i_8_1462, i_8_1534, i_8_1574, i_8_1586, i_8_1594, i_8_1679, i_8_1694, i_8_1696, i_8_1697, i_8_1724, i_8_1729, i_8_1739, i_8_1751, i_8_1754, i_8_1757, i_8_1804, i_8_1805, i_8_1814, i_8_1829, i_8_1856, i_8_1858, i_8_1867, i_8_1993, i_8_2036, i_8_2038, i_8_2039, i_8_2045, i_8_2047, i_8_2078, i_8_2096, i_8_2105, i_8_2117, i_8_2146, i_8_2187, i_8_2246, o_8_120);
	kernel_8_121 k_8_121(i_8_106, i_8_164, i_8_166, i_8_173, i_8_179, i_8_212, i_8_253, i_8_284, i_8_293, i_8_356, i_8_365, i_8_368, i_8_378, i_8_419, i_8_430, i_8_440, i_8_453, i_8_457, i_8_473, i_8_478, i_8_479, i_8_508, i_8_535, i_8_539, i_8_545, i_8_593, i_8_599, i_8_617, i_8_659, i_8_698, i_8_742, i_8_760, i_8_764, i_8_809, i_8_827, i_8_833, i_8_839, i_8_850, i_8_868, i_8_881, i_8_910, i_8_922, i_8_940, i_8_977, i_8_1045, i_8_1067, i_8_1075, i_8_1171, i_8_1208, i_8_1259, i_8_1264, i_8_1282, i_8_1344, i_8_1401, i_8_1417, i_8_1444, i_8_1454, i_8_1462, i_8_1508, i_8_1553, i_8_1574, i_8_1597, i_8_1640, i_8_1648, i_8_1666, i_8_1680, i_8_1702, i_8_1707, i_8_1731, i_8_1760, i_8_1779, i_8_1823, i_8_1826, i_8_1895, i_8_1903, i_8_1907, i_8_1920, i_8_1931, i_8_1993, i_8_1995, i_8_1996, i_8_2012, i_8_2117, i_8_2134, i_8_2137, i_8_2145, i_8_2146, i_8_2153, i_8_2156, i_8_2182, i_8_2185, i_8_2207, i_8_2210, i_8_2213, i_8_2215, i_8_2227, i_8_2245, i_8_2284, i_8_2288, i_8_2293, o_8_121);
	kernel_8_122 k_8_122(i_8_57, i_8_61, i_8_88, i_8_96, i_8_104, i_8_160, i_8_168, i_8_169, i_8_170, i_8_191, i_8_220, i_8_232, i_8_255, i_8_258, i_8_292, i_8_303, i_8_304, i_8_313, i_8_321, i_8_328, i_8_364, i_8_385, i_8_393, i_8_417, i_8_420, i_8_421, i_8_439, i_8_440, i_8_447, i_8_493, i_8_498, i_8_522, i_8_523, i_8_555, i_8_570, i_8_597, i_8_601, i_8_602, i_8_617, i_8_624, i_8_687, i_8_690, i_8_727, i_8_786, i_8_789, i_8_849, i_8_850, i_8_856, i_8_858, i_8_990, i_8_993, i_8_996, i_8_1050, i_8_1071, i_8_1075, i_8_1116, i_8_1122, i_8_1135, i_8_1188, i_8_1191, i_8_1222, i_8_1299, i_8_1305, i_8_1306, i_8_1307, i_8_1314, i_8_1318, i_8_1329, i_8_1346, i_8_1348, i_8_1470, i_8_1506, i_8_1509, i_8_1533, i_8_1536, i_8_1545, i_8_1561, i_8_1564, i_8_1570, i_8_1571, i_8_1574, i_8_1650, i_8_1651, i_8_1653, i_8_1681, i_8_1719, i_8_1727, i_8_1747, i_8_1750, i_8_1753, i_8_1795, i_8_1816, i_8_1956, i_8_1995, i_8_2031, i_8_2065, i_8_2122, i_8_2215, i_8_2226, i_8_2275, o_8_122);
	kernel_8_123 k_8_123(i_8_23, i_8_41, i_8_72, i_8_73, i_8_88, i_8_107, i_8_118, i_8_119, i_8_167, i_8_226, i_8_258, i_8_269, i_8_308, i_8_348, i_8_349, i_8_350, i_8_381, i_8_382, i_8_440, i_8_489, i_8_490, i_8_506, i_8_585, i_8_608, i_8_628, i_8_630, i_8_631, i_8_686, i_8_709, i_8_710, i_8_727, i_8_728, i_8_748, i_8_814, i_8_826, i_8_828, i_8_830, i_8_838, i_8_873, i_8_881, i_8_956, i_8_977, i_8_980, i_8_981, i_8_982, i_8_991, i_8_1027, i_8_1028, i_8_1029, i_8_1030, i_8_1031, i_8_1040, i_8_1058, i_8_1078, i_8_1161, i_8_1162, i_8_1226, i_8_1262, i_8_1279, i_8_1281, i_8_1296, i_8_1297, i_8_1300, i_8_1315, i_8_1319, i_8_1325, i_8_1327, i_8_1330, i_8_1334, i_8_1355, i_8_1437, i_8_1449, i_8_1467, i_8_1470, i_8_1471, i_8_1474, i_8_1705, i_8_1729, i_8_1746, i_8_1764, i_8_1765, i_8_1780, i_8_1787, i_8_1813, i_8_1832, i_8_1862, i_8_1888, i_8_1889, i_8_1949, i_8_1952, i_8_1965, i_8_2052, i_8_2059, i_8_2079, i_8_2114, i_8_2126, i_8_2140, i_8_2158, i_8_2241, i_8_2243, o_8_123);
	kernel_8_124 k_8_124(i_8_37, i_8_64, i_8_72, i_8_76, i_8_82, i_8_140, i_8_144, i_8_149, i_8_191, i_8_199, i_8_244, i_8_270, i_8_273, i_8_297, i_8_348, i_8_360, i_8_369, i_8_372, i_8_397, i_8_415, i_8_418, i_8_454, i_8_489, i_8_525, i_8_549, i_8_634, i_8_637, i_8_648, i_8_662, i_8_665, i_8_676, i_8_697, i_8_698, i_8_703, i_8_705, i_8_730, i_8_829, i_8_840, i_8_841, i_8_846, i_8_847, i_8_855, i_8_873, i_8_884, i_8_966, i_8_1027, i_8_1041, i_8_1042, i_8_1111, i_8_1112, i_8_1170, i_8_1224, i_8_1225, i_8_1235, i_8_1351, i_8_1387, i_8_1399, i_8_1458, i_8_1459, i_8_1479, i_8_1496, i_8_1522, i_8_1543, i_8_1550, i_8_1633, i_8_1638, i_8_1647, i_8_1648, i_8_1658, i_8_1682, i_8_1687, i_8_1705, i_8_1749, i_8_1765, i_8_1800, i_8_1810, i_8_1818, i_8_1819, i_8_1830, i_8_1845, i_8_1846, i_8_1864, i_8_1884, i_8_1885, i_8_1945, i_8_1996, i_8_2035, i_8_2038, i_8_2043, i_8_2044, i_8_2053, i_8_2125, i_8_2128, i_8_2141, i_8_2169, i_8_2173, i_8_2182, i_8_2253, i_8_2254, i_8_2255, o_8_124);
	kernel_8_125 k_8_125(i_8_13, i_8_52, i_8_103, i_8_112, i_8_130, i_8_142, i_8_165, i_8_199, i_8_221, i_8_237, i_8_254, i_8_334, i_8_361, i_8_391, i_8_424, i_8_453, i_8_455, i_8_459, i_8_475, i_8_492, i_8_507, i_8_523, i_8_544, i_8_598, i_8_607, i_8_624, i_8_654, i_8_659, i_8_660, i_8_662, i_8_685, i_8_695, i_8_696, i_8_699, i_8_704, i_8_755, i_8_760, i_8_765, i_8_786, i_8_797, i_8_806, i_8_840, i_8_841, i_8_895, i_8_926, i_8_931, i_8_940, i_8_966, i_8_1065, i_8_1108, i_8_1155, i_8_1197, i_8_1219, i_8_1237, i_8_1245, i_8_1258, i_8_1285, i_8_1290, i_8_1305, i_8_1321, i_8_1338, i_8_1398, i_8_1419, i_8_1426, i_8_1431, i_8_1433, i_8_1488, i_8_1527, i_8_1528, i_8_1650, i_8_1654, i_8_1682, i_8_1686, i_8_1689, i_8_1705, i_8_1801, i_8_1803, i_8_1804, i_8_1822, i_8_1825, i_8_1830, i_8_1831, i_8_1854, i_8_1855, i_8_1857, i_8_1858, i_8_1885, i_8_1980, i_8_1996, i_8_2092, i_8_2163, i_8_2203, i_8_2210, i_8_2224, i_8_2227, i_8_2260, i_8_2274, i_8_2281, i_8_2283, i_8_2290, o_8_125);
	kernel_8_126 k_8_126(i_8_14, i_8_47, i_8_53, i_8_121, i_8_224, i_8_233, i_8_247, i_8_268, i_8_295, i_8_305, i_8_346, i_8_367, i_8_395, i_8_437, i_8_455, i_8_502, i_8_536, i_8_568, i_8_608, i_8_650, i_8_673, i_8_685, i_8_716, i_8_732, i_8_752, i_8_874, i_8_877, i_8_884, i_8_950, i_8_992, i_8_1012, i_8_1039, i_8_1057, i_8_1114, i_8_1143, i_8_1162, i_8_1222, i_8_1237, i_8_1262, i_8_1286, i_8_1298, i_8_1306, i_8_1308, i_8_1311, i_8_1330, i_8_1331, i_8_1423, i_8_1455, i_8_1456, i_8_1474, i_8_1483, i_8_1486, i_8_1487, i_8_1537, i_8_1543, i_8_1546, i_8_1590, i_8_1600, i_8_1612, i_8_1637, i_8_1651, i_8_1672, i_8_1723, i_8_1730, i_8_1738, i_8_1744, i_8_1754, i_8_1761, i_8_1769, i_8_1772, i_8_1780, i_8_1781, i_8_1798, i_8_1803, i_8_1822, i_8_1843, i_8_1858, i_8_1903, i_8_1927, i_8_1978, i_8_1979, i_8_2003, i_8_2021, i_8_2024, i_8_2045, i_8_2053, i_8_2069, i_8_2083, i_8_2094, i_8_2102, i_8_2126, i_8_2130, i_8_2131, i_8_2149, i_8_2150, i_8_2171, i_8_2172, i_8_2174, i_8_2273, i_8_2299, o_8_126);
	kernel_8_127 k_8_127(i_8_94, i_8_111, i_8_124, i_8_190, i_8_191, i_8_223, i_8_231, i_8_248, i_8_301, i_8_328, i_8_346, i_8_365, i_8_368, i_8_376, i_8_420, i_8_439, i_8_445, i_8_455, i_8_471, i_8_492, i_8_499, i_8_522, i_8_523, i_8_530, i_8_591, i_8_597, i_8_634, i_8_637, i_8_645, i_8_660, i_8_673, i_8_681, i_8_696, i_8_697, i_8_770, i_8_841, i_8_871, i_8_877, i_8_879, i_8_880, i_8_888, i_8_924, i_8_958, i_8_961, i_8_969, i_8_976, i_8_993, i_8_1100, i_8_1105, i_8_1114, i_8_1137, i_8_1149, i_8_1189, i_8_1191, i_8_1192, i_8_1236, i_8_1239, i_8_1255, i_8_1266, i_8_1267, i_8_1281, i_8_1285, i_8_1356, i_8_1390, i_8_1444, i_8_1527, i_8_1535, i_8_1538, i_8_1545, i_8_1551, i_8_1596, i_8_1633, i_8_1634, i_8_1649, i_8_1741, i_8_1767, i_8_1770, i_8_1771, i_8_1779, i_8_1780, i_8_1814, i_8_1821, i_8_1840, i_8_1841, i_8_1859, i_8_1860, i_8_1861, i_8_1904, i_8_1991, i_8_2112, i_8_2137, i_8_2139, i_8_2141, i_8_2143, i_8_2146, i_8_2172, i_8_2215, i_8_2235, i_8_2247, i_8_2248, o_8_127);
	kernel_8_128 k_8_128(i_8_64, i_8_66, i_8_68, i_8_74, i_8_94, i_8_166, i_8_176, i_8_186, i_8_194, i_8_196, i_8_204, i_8_227, i_8_284, i_8_292, i_8_303, i_8_312, i_8_313, i_8_337, i_8_400, i_8_421, i_8_428, i_8_440, i_8_499, i_8_524, i_8_526, i_8_544, i_8_582, i_8_595, i_8_611, i_8_618, i_8_622, i_8_634, i_8_650, i_8_659, i_8_662, i_8_676, i_8_705, i_8_709, i_8_768, i_8_778, i_8_792, i_8_800, i_8_844, i_8_880, i_8_881, i_8_1023, i_8_1102, i_8_1104, i_8_1105, i_8_1123, i_8_1157, i_8_1162, i_8_1163, i_8_1219, i_8_1267, i_8_1317, i_8_1326, i_8_1383, i_8_1384, i_8_1427, i_8_1434, i_8_1437, i_8_1506, i_8_1551, i_8_1554, i_8_1555, i_8_1558, i_8_1559, i_8_1587, i_8_1609, i_8_1611, i_8_1681, i_8_1690, i_8_1743, i_8_1788, i_8_1822, i_8_1823, i_8_1880, i_8_1894, i_8_1913, i_8_1939, i_8_1940, i_8_1941, i_8_1942, i_8_1970, i_8_1974, i_8_1990, i_8_1999, i_8_2005, i_8_2092, i_8_2141, i_8_2156, i_8_2164, i_8_2166, i_8_2167, i_8_2183, i_8_2210, i_8_2216, i_8_2225, i_8_2279, o_8_128);
	kernel_8_129 k_8_129(i_8_22, i_8_48, i_8_64, i_8_72, i_8_73, i_8_74, i_8_76, i_8_90, i_8_94, i_8_136, i_8_171, i_8_194, i_8_197, i_8_297, i_8_325, i_8_505, i_8_550, i_8_585, i_8_586, i_8_588, i_8_595, i_8_621, i_8_622, i_8_624, i_8_630, i_8_631, i_8_632, i_8_652, i_8_653, i_8_684, i_8_702, i_8_703, i_8_707, i_8_820, i_8_829, i_8_969, i_8_990, i_8_991, i_8_1003, i_8_1012, i_8_1028, i_8_1029, i_8_1030, i_8_1031, i_8_1053, i_8_1054, i_8_1108, i_8_1198, i_8_1225, i_8_1263, i_8_1264, i_8_1265, i_8_1296, i_8_1297, i_8_1299, i_8_1351, i_8_1381, i_8_1395, i_8_1396, i_8_1398, i_8_1399, i_8_1400, i_8_1431, i_8_1449, i_8_1453, i_8_1454, i_8_1532, i_8_1621, i_8_1622, i_8_1701, i_8_1746, i_8_1767, i_8_1773, i_8_1776, i_8_1791, i_8_1802, i_8_1809, i_8_1818, i_8_1819, i_8_1821, i_8_1854, i_8_1855, i_8_1857, i_8_1899, i_8_1900, i_8_1903, i_8_1908, i_8_1911, i_8_1947, i_8_1948, i_8_1949, i_8_1963, i_8_1989, i_8_1992, i_8_1993, i_8_2134, i_8_2143, i_8_2246, i_8_2289, i_8_2294, o_8_129);
	kernel_8_130 k_8_130(i_8_22, i_8_25, i_8_37, i_8_54, i_8_184, i_8_208, i_8_243, i_8_247, i_8_301, i_8_310, i_8_323, i_8_346, i_8_365, i_8_368, i_8_375, i_8_376, i_8_438, i_8_451, i_8_487, i_8_490, i_8_493, i_8_499, i_8_525, i_8_529, i_8_556, i_8_557, i_8_600, i_8_637, i_8_645, i_8_661, i_8_667, i_8_673, i_8_711, i_8_719, i_8_760, i_8_773, i_8_788, i_8_820, i_8_841, i_8_869, i_8_881, i_8_919, i_8_931, i_8_941, i_8_977, i_8_1015, i_8_1153, i_8_1171, i_8_1187, i_8_1204, i_8_1222, i_8_1228, i_8_1238, i_8_1240, i_8_1255, i_8_1261, i_8_1309, i_8_1315, i_8_1349, i_8_1388, i_8_1407, i_8_1408, i_8_1409, i_8_1419, i_8_1438, i_8_1472, i_8_1501, i_8_1528, i_8_1543, i_8_1544, i_8_1553, i_8_1600, i_8_1606, i_8_1705, i_8_1732, i_8_1736, i_8_1787, i_8_1819, i_8_1824, i_8_1849, i_8_1871, i_8_1876, i_8_1927, i_8_1992, i_8_1993, i_8_1996, i_8_1999, i_8_2041, i_8_2124, i_8_2154, i_8_2155, i_8_2215, i_8_2217, i_8_2218, i_8_2273, i_8_2278, i_8_2284, i_8_2286, i_8_2287, i_8_2292, o_8_130);
	kernel_8_131 k_8_131(i_8_73, i_8_87, i_8_101, i_8_181, i_8_182, i_8_190, i_8_191, i_8_232, i_8_243, i_8_244, i_8_303, i_8_304, i_8_339, i_8_383, i_8_391, i_8_396, i_8_397, i_8_454, i_8_473, i_8_490, i_8_594, i_8_595, i_8_596, i_8_628, i_8_629, i_8_632, i_8_665, i_8_716, i_8_719, i_8_748, i_8_752, i_8_757, i_8_850, i_8_855, i_8_856, i_8_858, i_8_969, i_8_994, i_8_1033, i_8_1036, i_8_1047, i_8_1057, i_8_1073, i_8_1078, i_8_1099, i_8_1100, i_8_1262, i_8_1283, i_8_1291, i_8_1306, i_8_1307, i_8_1330, i_8_1354, i_8_1372, i_8_1405, i_8_1439, i_8_1459, i_8_1470, i_8_1505, i_8_1507, i_8_1521, i_8_1529, i_8_1538, i_8_1607, i_8_1647, i_8_1649, i_8_1670, i_8_1675, i_8_1683, i_8_1736, i_8_1805, i_8_1807, i_8_1809, i_8_1811, i_8_1837, i_8_1862, i_8_1882, i_8_1883, i_8_1937, i_8_1964, i_8_1982, i_8_1993, i_8_1994, i_8_2007, i_8_2057, i_8_2072, i_8_2106, i_8_2139, i_8_2140, i_8_2147, i_8_2153, i_8_2155, i_8_2156, i_8_2161, i_8_2180, i_8_2215, i_8_2241, i_8_2246, i_8_2267, i_8_2275, o_8_131);
	kernel_8_132 k_8_132(i_8_9, i_8_12, i_8_18, i_8_42, i_8_69, i_8_78, i_8_103, i_8_138, i_8_151, i_8_166, i_8_174, i_8_196, i_8_229, i_8_283, i_8_300, i_8_301, i_8_318, i_8_337, i_8_338, i_8_365, i_8_367, i_8_397, i_8_496, i_8_529, i_8_537, i_8_544, i_8_573, i_8_672, i_8_703, i_8_704, i_8_707, i_8_733, i_8_773, i_8_806, i_8_864, i_8_865, i_8_866, i_8_937, i_8_979, i_8_993, i_8_1003, i_8_1057, i_8_1074, i_8_1104, i_8_1105, i_8_1151, i_8_1224, i_8_1225, i_8_1228, i_8_1239, i_8_1258, i_8_1260, i_8_1261, i_8_1262, i_8_1291, i_8_1292, i_8_1323, i_8_1333, i_8_1335, i_8_1356, i_8_1384, i_8_1410, i_8_1412, i_8_1429, i_8_1449, i_8_1464, i_8_1468, i_8_1471, i_8_1491, i_8_1515, i_8_1527, i_8_1531, i_8_1562, i_8_1645, i_8_1653, i_8_1654, i_8_1686, i_8_1723, i_8_1746, i_8_1751, i_8_1807, i_8_1823, i_8_1858, i_8_1894, i_8_1907, i_8_1912, i_8_1956, i_8_1962, i_8_1963, i_8_1984, i_8_1995, i_8_2106, i_8_2145, i_8_2151, i_8_2152, i_8_2174, i_8_2200, i_8_2202, i_8_2245, i_8_2259, o_8_132);
	kernel_8_133 k_8_133(i_8_13, i_8_52, i_8_115, i_8_139, i_8_151, i_8_259, i_8_283, i_8_301, i_8_304, i_8_305, i_8_307, i_8_367, i_8_382, i_8_392, i_8_401, i_8_420, i_8_421, i_8_455, i_8_493, i_8_508, i_8_509, i_8_553, i_8_571, i_8_580, i_8_583, i_8_589, i_8_607, i_8_610, i_8_631, i_8_638, i_8_643, i_8_644, i_8_661, i_8_678, i_8_866, i_8_895, i_8_967, i_8_992, i_8_1012, i_8_1102, i_8_1103, i_8_1108, i_8_1111, i_8_1130, i_8_1157, i_8_1183, i_8_1201, i_8_1229, i_8_1246, i_8_1266, i_8_1267, i_8_1299, i_8_1301, i_8_1327, i_8_1328, i_8_1336, i_8_1355, i_8_1357, i_8_1435, i_8_1436, i_8_1441, i_8_1462, i_8_1463, i_8_1471, i_8_1477, i_8_1525, i_8_1526, i_8_1538, i_8_1541, i_8_1542, i_8_1552, i_8_1574, i_8_1632, i_8_1633, i_8_1642, i_8_1655, i_8_1678, i_8_1705, i_8_1749, i_8_1750, i_8_1753, i_8_1767, i_8_1776, i_8_1825, i_8_1841, i_8_1882, i_8_1894, i_8_1939, i_8_1940, i_8_1957, i_8_1958, i_8_1967, i_8_1975, i_8_1992, i_8_1995, i_8_1996, i_8_2136, i_8_2138, i_8_2210, i_8_2231, o_8_133);
	kernel_8_134 k_8_134(i_8_20, i_8_31, i_8_35, i_8_50, i_8_55, i_8_103, i_8_104, i_8_115, i_8_142, i_8_167, i_8_181, i_8_221, i_8_232, i_8_233, i_8_253, i_8_255, i_8_289, i_8_292, i_8_293, i_8_297, i_8_306, i_8_343, i_8_344, i_8_378, i_8_386, i_8_414, i_8_442, i_8_451, i_8_476, i_8_479, i_8_481, i_8_482, i_8_484, i_8_497, i_8_526, i_8_588, i_8_589, i_8_595, i_8_596, i_8_612, i_8_689, i_8_706, i_8_713, i_8_760, i_8_761, i_8_766, i_8_767, i_8_784, i_8_787, i_8_797, i_8_811, i_8_812, i_8_838, i_8_847, i_8_850, i_8_859, i_8_929, i_8_992, i_8_1058, i_8_1118, i_8_1183, i_8_1189, i_8_1216, i_8_1219, i_8_1238, i_8_1264, i_8_1265, i_8_1269, i_8_1271, i_8_1282, i_8_1291, i_8_1300, i_8_1306, i_8_1315, i_8_1318, i_8_1404, i_8_1470, i_8_1540, i_8_1550, i_8_1557, i_8_1558, i_8_1560, i_8_1562, i_8_1621, i_8_1633, i_8_1730, i_8_1739, i_8_1762, i_8_1786, i_8_1787, i_8_1831, i_8_1873, i_8_1904, i_8_1949, i_8_2029, i_8_2037, i_8_2089, i_8_2090, i_8_2093, i_8_2287, o_8_134);
	kernel_8_135 k_8_135(i_8_32, i_8_46, i_8_53, i_8_56, i_8_67, i_8_101, i_8_166, i_8_257, i_8_281, i_8_311, i_8_363, i_8_371, i_8_416, i_8_571, i_8_603, i_8_606, i_8_655, i_8_656, i_8_705, i_8_768, i_8_838, i_8_839, i_8_860, i_8_866, i_8_967, i_8_994, i_8_1056, i_8_1110, i_8_1111, i_8_1198, i_8_1217, i_8_1220, i_8_1229, i_8_1234, i_8_1265, i_8_1266, i_8_1267, i_8_1292, i_8_1318, i_8_1323, i_8_1326, i_8_1340, i_8_1351, i_8_1360, i_8_1367, i_8_1400, i_8_1427, i_8_1489, i_8_1504, i_8_1514, i_8_1522, i_8_1526, i_8_1548, i_8_1555, i_8_1557, i_8_1622, i_8_1630, i_8_1651, i_8_1665, i_8_1675, i_8_1684, i_8_1693, i_8_1703, i_8_1712, i_8_1757, i_8_1770, i_8_1777, i_8_1814, i_8_1818, i_8_1819, i_8_1820, i_8_1822, i_8_1825, i_8_1827, i_8_1856, i_8_1885, i_8_1891, i_8_1910, i_8_1966, i_8_1973, i_8_1975, i_8_1996, i_8_1997, i_8_2014, i_8_2097, i_8_2099, i_8_2128, i_8_2142, i_8_2146, i_8_2147, i_8_2148, i_8_2153, i_8_2197, i_8_2225, i_8_2244, i_8_2246, i_8_2258, i_8_2262, i_8_2272, i_8_2281, o_8_135);
	kernel_8_136 k_8_136(i_8_140, i_8_147, i_8_148, i_8_149, i_8_150, i_8_151, i_8_165, i_8_166, i_8_189, i_8_192, i_8_194, i_8_195, i_8_211, i_8_214, i_8_226, i_8_227, i_8_271, i_8_303, i_8_368, i_8_386, i_8_427, i_8_453, i_8_454, i_8_472, i_8_483, i_8_484, i_8_493, i_8_508, i_8_530, i_8_582, i_8_602, i_8_618, i_8_642, i_8_657, i_8_658, i_8_661, i_8_678, i_8_701, i_8_703, i_8_705, i_8_732, i_8_750, i_8_751, i_8_752, i_8_832, i_8_833, i_8_861, i_8_1003, i_8_1157, i_8_1160, i_8_1164, i_8_1256, i_8_1285, i_8_1327, i_8_1335, i_8_1336, i_8_1355, i_8_1356, i_8_1357, i_8_1399, i_8_1434, i_8_1436, i_8_1438, i_8_1439, i_8_1479, i_8_1481, i_8_1488, i_8_1593, i_8_1596, i_8_1599, i_8_1623, i_8_1644, i_8_1660, i_8_1662, i_8_1663, i_8_1749, i_8_1754, i_8_1773, i_8_1776, i_8_1787, i_8_1824, i_8_1837, i_8_1875, i_8_1886, i_8_1919, i_8_2003, i_8_2011, i_8_2012, i_8_2089, i_8_2091, i_8_2095, i_8_2119, i_8_2154, i_8_2170, i_8_2174, i_8_2177, i_8_2253, i_8_2256, i_8_2257, i_8_2258, o_8_136);
	kernel_8_137 k_8_137(i_8_33, i_8_85, i_8_114, i_8_141, i_8_159, i_8_165, i_8_186, i_8_204, i_8_220, i_8_222, i_8_223, i_8_230, i_8_231, i_8_240, i_8_298, i_8_420, i_8_476, i_8_501, i_8_546, i_8_549, i_8_550, i_8_609, i_8_625, i_8_636, i_8_700, i_8_762, i_8_777, i_8_780, i_8_824, i_8_825, i_8_834, i_8_868, i_8_870, i_8_877, i_8_878, i_8_879, i_8_888, i_8_895, i_8_949, i_8_991, i_8_993, i_8_994, i_8_995, i_8_1015, i_8_1027, i_8_1030, i_8_1073, i_8_1076, i_8_1086, i_8_1108, i_8_1112, i_8_1228, i_8_1266, i_8_1267, i_8_1281, i_8_1282, i_8_1284, i_8_1308, i_8_1329, i_8_1393, i_8_1402, i_8_1454, i_8_1470, i_8_1525, i_8_1527, i_8_1537, i_8_1544, i_8_1552, i_8_1553, i_8_1559, i_8_1653, i_8_1677, i_8_1678, i_8_1698, i_8_1705, i_8_1707, i_8_1721, i_8_1723, i_8_1725, i_8_1726, i_8_1729, i_8_1747, i_8_1779, i_8_1806, i_8_1808, i_8_1821, i_8_1834, i_8_1838, i_8_1867, i_8_1903, i_8_1948, i_8_2011, i_8_2046, i_8_2121, i_8_2139, i_8_2147, i_8_2149, i_8_2175, i_8_2214, i_8_2301, o_8_137);
	kernel_8_138 k_8_138(i_8_34, i_8_107, i_8_114, i_8_115, i_8_143, i_8_205, i_8_259, i_8_296, i_8_380, i_8_452, i_8_470, i_8_492, i_8_528, i_8_590, i_8_605, i_8_660, i_8_662, i_8_663, i_8_673, i_8_681, i_8_682, i_8_683, i_8_692, i_8_736, i_8_870, i_8_876, i_8_898, i_8_899, i_8_994, i_8_1026, i_8_1028, i_8_1075, i_8_1136, i_8_1157, i_8_1160, i_8_1224, i_8_1257, i_8_1258, i_8_1264, i_8_1273, i_8_1274, i_8_1276, i_8_1281, i_8_1340, i_8_1342, i_8_1343, i_8_1351, i_8_1355, i_8_1356, i_8_1403, i_8_1437, i_8_1438, i_8_1439, i_8_1444, i_8_1451, i_8_1489, i_8_1492, i_8_1503, i_8_1527, i_8_1529, i_8_1543, i_8_1562, i_8_1592, i_8_1599, i_8_1601, i_8_1603, i_8_1623, i_8_1625, i_8_1627, i_8_1628, i_8_1634, i_8_1636, i_8_1637, i_8_1645, i_8_1651, i_8_1675, i_8_1714, i_8_1716, i_8_1717, i_8_1748, i_8_1750, i_8_1751, i_8_1754, i_8_1818, i_8_1852, i_8_1857, i_8_1946, i_8_1964, i_8_1966, i_8_2128, i_8_2137, i_8_2138, i_8_2140, i_8_2141, i_8_2143, i_8_2144, i_8_2156, i_8_2214, i_8_2242, i_8_2288, o_8_138);
	kernel_8_139 k_8_139(i_8_39, i_8_42, i_8_44, i_8_49, i_8_66, i_8_69, i_8_70, i_8_93, i_8_105, i_8_175, i_8_202, i_8_333, i_8_355, i_8_367, i_8_372, i_8_384, i_8_426, i_8_444, i_8_454, i_8_481, i_8_484, i_8_540, i_8_601, i_8_634, i_8_652, i_8_662, i_8_687, i_8_703, i_8_769, i_8_784, i_8_801, i_8_822, i_8_866, i_8_883, i_8_930, i_8_931, i_8_939, i_8_949, i_8_966, i_8_981, i_8_1071, i_8_1081, i_8_1096, i_8_1110, i_8_1135, i_8_1170, i_8_1213, i_8_1228, i_8_1233, i_8_1263, i_8_1267, i_8_1284, i_8_1290, i_8_1294, i_8_1410, i_8_1425, i_8_1470, i_8_1488, i_8_1497, i_8_1524, i_8_1596, i_8_1611, i_8_1648, i_8_1650, i_8_1659, i_8_1678, i_8_1689, i_8_1696, i_8_1704, i_8_1705, i_8_1747, i_8_1764, i_8_1777, i_8_1806, i_8_1807, i_8_1821, i_8_1869, i_8_1875, i_8_1882, i_8_1918, i_8_1919, i_8_1949, i_8_1972, i_8_1992, i_8_1995, i_8_2008, i_8_2010, i_8_2056, i_8_2089, i_8_2146, i_8_2148, i_8_2172, i_8_2179, i_8_2181, i_8_2182, i_8_2226, i_8_2241, i_8_2280, i_8_2281, i_8_2299, o_8_139);
	kernel_8_140 k_8_140(i_8_31, i_8_77, i_8_89, i_8_161, i_8_170, i_8_224, i_8_229, i_8_233, i_8_259, i_8_305, i_8_347, i_8_359, i_8_366, i_8_458, i_8_481, i_8_493, i_8_525, i_8_526, i_8_530, i_8_557, i_8_593, i_8_601, i_8_604, i_8_663, i_8_665, i_8_692, i_8_698, i_8_699, i_8_719, i_8_763, i_8_826, i_8_827, i_8_845, i_8_869, i_8_880, i_8_896, i_8_974, i_8_994, i_8_1016, i_8_1031, i_8_1075, i_8_1097, i_8_1106, i_8_1115, i_8_1124, i_8_1133, i_8_1160, i_8_1184, i_8_1196, i_8_1232, i_8_1270, i_8_1277, i_8_1282, i_8_1285, i_8_1301, i_8_1349, i_8_1388, i_8_1441, i_8_1454, i_8_1457, i_8_1471, i_8_1472, i_8_1475, i_8_1484, i_8_1537, i_8_1546, i_8_1550, i_8_1553, i_8_1592, i_8_1633, i_8_1634, i_8_1636, i_8_1642, i_8_1647, i_8_1655, i_8_1678, i_8_1681, i_8_1682, i_8_1718, i_8_1733, i_8_1768, i_8_1807, i_8_1824, i_8_1826, i_8_1834, i_8_1840, i_8_1844, i_8_1870, i_8_1898, i_8_2008, i_8_2046, i_8_2111, i_8_2129, i_8_2132, i_8_2186, i_8_2194, i_8_2204, i_8_2249, i_8_2291, i_8_2294, o_8_140);
	kernel_8_141 k_8_141(i_8_18, i_8_34, i_8_35, i_8_81, i_8_84, i_8_93, i_8_94, i_8_143, i_8_221, i_8_244, i_8_288, i_8_298, i_8_301, i_8_344, i_8_346, i_8_369, i_8_374, i_8_383, i_8_415, i_8_434, i_8_459, i_8_460, i_8_471, i_8_481, i_8_482, i_8_485, i_8_522, i_8_526, i_8_550, i_8_613, i_8_615, i_8_622, i_8_715, i_8_756, i_8_780, i_8_793, i_8_812, i_8_844, i_8_874, i_8_895, i_8_946, i_8_977, i_8_988, i_8_1028, i_8_1029, i_8_1113, i_8_1153, i_8_1156, i_8_1216, i_8_1233, i_8_1235, i_8_1251, i_8_1269, i_8_1270, i_8_1283, i_8_1300, i_8_1315, i_8_1337, i_8_1434, i_8_1444, i_8_1468, i_8_1549, i_8_1584, i_8_1586, i_8_1596, i_8_1597, i_8_1602, i_8_1612, i_8_1615, i_8_1630, i_8_1657, i_8_1666, i_8_1678, i_8_1679, i_8_1707, i_8_1743, i_8_1753, i_8_1754, i_8_1762, i_8_1780, i_8_1783, i_8_1794, i_8_1805, i_8_1840, i_8_1858, i_8_1859, i_8_1918, i_8_1946, i_8_1950, i_8_1963, i_8_2050, i_8_2073, i_8_2125, i_8_2126, i_8_2139, i_8_2140, i_8_2179, i_8_2183, i_8_2227, i_8_2290, o_8_141);
	kernel_8_142 k_8_142(i_8_12, i_8_22, i_8_28, i_8_52, i_8_67, i_8_75, i_8_79, i_8_136, i_8_222, i_8_225, i_8_321, i_8_333, i_8_360, i_8_364, i_8_366, i_8_367, i_8_381, i_8_391, i_8_397, i_8_398, i_8_400, i_8_418, i_8_426, i_8_427, i_8_430, i_8_454, i_8_507, i_8_516, i_8_526, i_8_571, i_8_604, i_8_634, i_8_639, i_8_661, i_8_747, i_8_750, i_8_784, i_8_849, i_8_850, i_8_860, i_8_937, i_8_969, i_8_970, i_8_971, i_8_973, i_8_1102, i_8_1107, i_8_1109, i_8_1144, i_8_1153, i_8_1162, i_8_1196, i_8_1201, i_8_1224, i_8_1297, i_8_1300, i_8_1327, i_8_1336, i_8_1362, i_8_1365, i_8_1399, i_8_1422, i_8_1432, i_8_1436, i_8_1441, i_8_1461, i_8_1471, i_8_1477, i_8_1480, i_8_1491, i_8_1513, i_8_1558, i_8_1615, i_8_1633, i_8_1679, i_8_1683, i_8_1692, i_8_1701, i_8_1705, i_8_1714, i_8_1750, i_8_1764, i_8_1768, i_8_1774, i_8_1809, i_8_1839, i_8_1849, i_8_1912, i_8_1917, i_8_1926, i_8_1935, i_8_1972, i_8_2070, i_8_2073, i_8_2134, i_8_2145, i_8_2155, i_8_2169, i_8_2242, i_8_2244, o_8_142);
	kernel_8_143 k_8_143(i_8_41, i_8_44, i_8_48, i_8_54, i_8_57, i_8_66, i_8_103, i_8_108, i_8_150, i_8_189, i_8_203, i_8_225, i_8_226, i_8_252, i_8_253, i_8_297, i_8_378, i_8_390, i_8_433, i_8_534, i_8_553, i_8_594, i_8_604, i_8_610, i_8_612, i_8_639, i_8_648, i_8_652, i_8_658, i_8_675, i_8_696, i_8_699, i_8_700, i_8_763, i_8_780, i_8_846, i_8_849, i_8_855, i_8_857, i_8_858, i_8_880, i_8_967, i_8_982, i_8_988, i_8_1032, i_8_1059, i_8_1083, i_8_1134, i_8_1137, i_8_1152, i_8_1157, i_8_1196, i_8_1263, i_8_1278, i_8_1281, i_8_1300, i_8_1314, i_8_1326, i_8_1354, i_8_1357, i_8_1383, i_8_1461, i_8_1473, i_8_1512, i_8_1530, i_8_1542, i_8_1557, i_8_1558, i_8_1602, i_8_1605, i_8_1623, i_8_1656, i_8_1674, i_8_1683, i_8_1695, i_8_1710, i_8_1713, i_8_1755, i_8_1759, i_8_1773, i_8_1791, i_8_1803, i_8_1809, i_8_1818, i_8_1885, i_8_1980, i_8_1990, i_8_1992, i_8_1993, i_8_1996, i_8_2052, i_8_2076, i_8_2109, i_8_2156, i_8_2161, i_8_2232, i_8_2233, i_8_2235, i_8_2244, i_8_2253, o_8_143);
	kernel_8_144 k_8_144(i_8_11, i_8_35, i_8_49, i_8_59, i_8_77, i_8_111, i_8_226, i_8_229, i_8_230, i_8_231, i_8_282, i_8_293, i_8_310, i_8_325, i_8_337, i_8_342, i_8_343, i_8_345, i_8_364, i_8_370, i_8_373, i_8_423, i_8_443, i_8_450, i_8_454, i_8_479, i_8_481, i_8_482, i_8_499, i_8_505, i_8_522, i_8_526, i_8_544, i_8_549, i_8_554, i_8_613, i_8_662, i_8_687, i_8_688, i_8_697, i_8_704, i_8_715, i_8_769, i_8_783, i_8_786, i_8_795, i_8_815, i_8_832, i_8_840, i_8_875, i_8_931, i_8_932, i_8_954, i_8_955, i_8_973, i_8_985, i_8_1047, i_8_1057, i_8_1090, i_8_1099, i_8_1121, i_8_1123, i_8_1220, i_8_1243, i_8_1251, i_8_1266, i_8_1273, i_8_1274, i_8_1282, i_8_1305, i_8_1306, i_8_1328, i_8_1331, i_8_1346, i_8_1387, i_8_1401, i_8_1407, i_8_1537, i_8_1564, i_8_1571, i_8_1588, i_8_1612, i_8_1621, i_8_1629, i_8_1633, i_8_1651, i_8_1675, i_8_1721, i_8_1741, i_8_1804, i_8_1884, i_8_2003, i_8_2109, i_8_2145, i_8_2148, i_8_2191, i_8_2209, i_8_2215, i_8_2223, i_8_2289, o_8_144);
	kernel_8_145 k_8_145(i_8_24, i_8_52, i_8_67, i_8_165, i_8_210, i_8_231, i_8_232, i_8_301, i_8_310, i_8_325, i_8_336, i_8_342, i_8_349, i_8_354, i_8_363, i_8_366, i_8_367, i_8_426, i_8_430, i_8_475, i_8_492, i_8_498, i_8_529, i_8_552, i_8_580, i_8_588, i_8_598, i_8_604, i_8_606, i_8_607, i_8_609, i_8_610, i_8_612, i_8_615, i_8_651, i_8_660, i_8_681, i_8_702, i_8_735, i_8_768, i_8_780, i_8_795, i_8_876, i_8_921, i_8_927, i_8_958, i_8_1020, i_8_1053, i_8_1068, i_8_1074, i_8_1101, i_8_1156, i_8_1170, i_8_1173, i_8_1228, i_8_1236, i_8_1251, i_8_1254, i_8_1291, i_8_1292, i_8_1311, i_8_1317, i_8_1354, i_8_1454, i_8_1470, i_8_1489, i_8_1524, i_8_1560, i_8_1623, i_8_1641, i_8_1649, i_8_1650, i_8_1678, i_8_1704, i_8_1707, i_8_1800, i_8_1819, i_8_1821, i_8_1824, i_8_1825, i_8_1861, i_8_1884, i_8_1941, i_8_1966, i_8_2001, i_8_2004, i_8_2016, i_8_2019, i_8_2020, i_8_2037, i_8_2073, i_8_2113, i_8_2146, i_8_2181, i_8_2199, i_8_2208, i_8_2209, i_8_2226, i_8_2235, i_8_2244, o_8_145);
	kernel_8_146 k_8_146(i_8_4, i_8_13, i_8_22, i_8_53, i_8_67, i_8_97, i_8_184, i_8_239, i_8_246, i_8_263, i_8_298, i_8_327, i_8_364, i_8_365, i_8_368, i_8_437, i_8_455, i_8_464, i_8_473, i_8_507, i_8_517, i_8_518, i_8_534, i_8_535, i_8_553, i_8_571, i_8_589, i_8_592, i_8_595, i_8_615, i_8_624, i_8_632, i_8_634, i_8_652, i_8_660, i_8_661, i_8_663, i_8_665, i_8_682, i_8_706, i_8_751, i_8_841, i_8_869, i_8_938, i_8_941, i_8_958, i_8_965, i_8_977, i_8_1039, i_8_1042, i_8_1079, i_8_1102, i_8_1111, i_8_1122, i_8_1169, i_8_1210, i_8_1222, i_8_1223, i_8_1249, i_8_1267, i_8_1303, i_8_1318, i_8_1354, i_8_1381, i_8_1384, i_8_1397, i_8_1438, i_8_1456, i_8_1458, i_8_1469, i_8_1489, i_8_1513, i_8_1528, i_8_1532, i_8_1564, i_8_1641, i_8_1659, i_8_1687, i_8_1697, i_8_1729, i_8_1767, i_8_1774, i_8_1813, i_8_1824, i_8_1825, i_8_1826, i_8_1884, i_8_1885, i_8_1957, i_8_1992, i_8_1995, i_8_1996, i_8_2115, i_8_2119, i_8_2146, i_8_2226, i_8_2236, i_8_2242, i_8_2248, i_8_2299, o_8_146);
	kernel_8_147 k_8_147(i_8_28, i_8_97, i_8_98, i_8_136, i_8_224, i_8_356, i_8_370, i_8_376, i_8_424, i_8_426, i_8_427, i_8_463, i_8_475, i_8_476, i_8_488, i_8_491, i_8_493, i_8_502, i_8_563, i_8_570, i_8_592, i_8_625, i_8_632, i_8_666, i_8_679, i_8_683, i_8_696, i_8_697, i_8_705, i_8_725, i_8_757, i_8_773, i_8_778, i_8_781, i_8_783, i_8_786, i_8_787, i_8_790, i_8_812, i_8_826, i_8_829, i_8_838, i_8_841, i_8_842, i_8_847, i_8_848, i_8_869, i_8_874, i_8_917, i_8_932, i_8_1000, i_8_1057, i_8_1072, i_8_1135, i_8_1189, i_8_1234, i_8_1271, i_8_1328, i_8_1363, i_8_1369, i_8_1454, i_8_1457, i_8_1470, i_8_1524, i_8_1589, i_8_1607, i_8_1648, i_8_1655, i_8_1684, i_8_1696, i_8_1700, i_8_1729, i_8_1732, i_8_1749, i_8_1805, i_8_1846, i_8_1855, i_8_1856, i_8_1857, i_8_1858, i_8_1859, i_8_1861, i_8_1867, i_8_1888, i_8_1895, i_8_1898, i_8_1904, i_8_1981, i_8_2029, i_8_2072, i_8_2090, i_8_2174, i_8_2182, i_8_2183, i_8_2185, i_8_2191, i_8_2280, i_8_2290, i_8_2292, i_8_2294, o_8_147);
	kernel_8_148 k_8_148(i_8_9, i_8_70, i_8_118, i_8_123, i_8_127, i_8_164, i_8_180, i_8_218, i_8_228, i_8_236, i_8_271, i_8_313, i_8_352, i_8_378, i_8_388, i_8_425, i_8_433, i_8_438, i_8_531, i_8_551, i_8_553, i_8_567, i_8_603, i_8_621, i_8_649, i_8_698, i_8_804, i_8_831, i_8_832, i_8_837, i_8_848, i_8_878, i_8_885, i_8_921, i_8_930, i_8_981, i_8_982, i_8_984, i_8_985, i_8_990, i_8_994, i_8_999, i_8_1011, i_8_1012, i_8_1074, i_8_1089, i_8_1090, i_8_1128, i_8_1165, i_8_1183, i_8_1280, i_8_1291, i_8_1308, i_8_1317, i_8_1320, i_8_1387, i_8_1393, i_8_1401, i_8_1407, i_8_1424, i_8_1620, i_8_1621, i_8_1623, i_8_1641, i_8_1651, i_8_1654, i_8_1683, i_8_1686, i_8_1687, i_8_1728, i_8_1731, i_8_1734, i_8_1782, i_8_1794, i_8_1803, i_8_1829, i_8_1858, i_8_1864, i_8_1882, i_8_1884, i_8_1893, i_8_1896, i_8_1906, i_8_2055, i_8_2070, i_8_2073, i_8_2074, i_8_2083, i_8_2086, i_8_2092, i_8_2097, i_8_2148, i_8_2155, i_8_2215, i_8_2229, i_8_2232, i_8_2236, i_8_2247, i_8_2248, i_8_2258, o_8_148);
	kernel_8_149 k_8_149(i_8_34, i_8_44, i_8_87, i_8_106, i_8_159, i_8_160, i_8_161, i_8_168, i_8_204, i_8_205, i_8_214, i_8_222, i_8_258, i_8_340, i_8_345, i_8_417, i_8_463, i_8_464, i_8_474, i_8_478, i_8_480, i_8_483, i_8_524, i_8_526, i_8_557, i_8_594, i_8_601, i_8_619, i_8_629, i_8_661, i_8_664, i_8_718, i_8_726, i_8_748, i_8_749, i_8_764, i_8_773, i_8_834, i_8_907, i_8_925, i_8_952, i_8_984, i_8_985, i_8_988, i_8_997, i_8_1069, i_8_1072, i_8_1086, i_8_1087, i_8_1114, i_8_1137, i_8_1148, i_8_1174, i_8_1193, i_8_1199, i_8_1219, i_8_1254, i_8_1302, i_8_1320, i_8_1338, i_8_1420, i_8_1423, i_8_1426, i_8_1434, i_8_1484, i_8_1528, i_8_1537, i_8_1544, i_8_1549, i_8_1582, i_8_1610, i_8_1614, i_8_1615, i_8_1617, i_8_1633, i_8_1666, i_8_1680, i_8_1734, i_8_1735, i_8_1751, i_8_1752, i_8_1761, i_8_1799, i_8_1836, i_8_1869, i_8_1932, i_8_2001, i_8_2002, i_8_2004, i_8_2013, i_8_2014, i_8_2049, i_8_2073, i_8_2094, i_8_2113, i_8_2156, i_8_2175, i_8_2182, i_8_2266, i_8_2293, o_8_149);
	kernel_8_150 k_8_150(i_8_147, i_8_190, i_8_194, i_8_228, i_8_229, i_8_283, i_8_310, i_8_318, i_8_346, i_8_361, i_8_379, i_8_418, i_8_450, i_8_452, i_8_490, i_8_571, i_8_598, i_8_628, i_8_652, i_8_658, i_8_693, i_8_694, i_8_695, i_8_700, i_8_705, i_8_748, i_8_751, i_8_778, i_8_838, i_8_839, i_8_841, i_8_874, i_8_876, i_8_877, i_8_878, i_8_966, i_8_967, i_8_990, i_8_991, i_8_1000, i_8_1002, i_8_1034, i_8_1036, i_8_1037, i_8_1039, i_8_1046, i_8_1075, i_8_1147, i_8_1164, i_8_1226, i_8_1234, i_8_1268, i_8_1270, i_8_1283, i_8_1354, i_8_1355, i_8_1399, i_8_1407, i_8_1411, i_8_1452, i_8_1507, i_8_1524, i_8_1539, i_8_1540, i_8_1542, i_8_1605, i_8_1621, i_8_1622, i_8_1625, i_8_1629, i_8_1641, i_8_1642, i_8_1703, i_8_1729, i_8_1732, i_8_1767, i_8_1777, i_8_1807, i_8_1821, i_8_1822, i_8_1894, i_8_1903, i_8_1904, i_8_1936, i_8_1984, i_8_1992, i_8_1996, i_8_2009, i_8_2011, i_8_2014, i_8_2055, i_8_2056, i_8_2082, i_8_2083, i_8_2147, i_8_2151, i_8_2155, i_8_2170, i_8_2225, i_8_2272, o_8_150);
	kernel_8_151 k_8_151(i_8_11, i_8_33, i_8_51, i_8_67, i_8_74, i_8_96, i_8_120, i_8_137, i_8_142, i_8_159, i_8_191, i_8_254, i_8_262, i_8_310, i_8_312, i_8_346, i_8_348, i_8_372, i_8_441, i_8_448, i_8_456, i_8_484, i_8_492, i_8_524, i_8_598, i_8_600, i_8_601, i_8_690, i_8_691, i_8_718, i_8_734, i_8_735, i_8_736, i_8_799, i_8_800, i_8_826, i_8_838, i_8_923, i_8_946, i_8_1014, i_8_1015, i_8_1026, i_8_1060, i_8_1077, i_8_1113, i_8_1119, i_8_1120, i_8_1188, i_8_1231, i_8_1258, i_8_1273, i_8_1300, i_8_1305, i_8_1306, i_8_1324, i_8_1348, i_8_1387, i_8_1418, i_8_1425, i_8_1506, i_8_1507, i_8_1525, i_8_1578, i_8_1581, i_8_1582, i_8_1587, i_8_1588, i_8_1623, i_8_1632, i_8_1647, i_8_1648, i_8_1677, i_8_1686, i_8_1699, i_8_1720, i_8_1721, i_8_1740, i_8_1742, i_8_1749, i_8_1786, i_8_1789, i_8_1791, i_8_1876, i_8_1905, i_8_1906, i_8_1907, i_8_2004, i_8_2031, i_8_2049, i_8_2050, i_8_2092, i_8_2143, i_8_2155, i_8_2156, i_8_2157, i_8_2158, i_8_2182, i_8_2214, i_8_2219, i_8_2262, o_8_151);
	kernel_8_152 k_8_152(i_8_4, i_8_57, i_8_86, i_8_95, i_8_97, i_8_157, i_8_181, i_8_184, i_8_185, i_8_224, i_8_227, i_8_233, i_8_374, i_8_388, i_8_417, i_8_436, i_8_437, i_8_454, i_8_459, i_8_462, i_8_475, i_8_485, i_8_499, i_8_505, i_8_550, i_8_595, i_8_599, i_8_610, i_8_621, i_8_625, i_8_670, i_8_671, i_8_696, i_8_713, i_8_716, i_8_758, i_8_766, i_8_775, i_8_793, i_8_820, i_8_824, i_8_866, i_8_923, i_8_1009, i_8_1031, i_8_1081, i_8_1118, i_8_1180, i_8_1188, i_8_1204, i_8_1235, i_8_1255, i_8_1261, i_8_1269, i_8_1270, i_8_1280, i_8_1282, i_8_1283, i_8_1298, i_8_1308, i_8_1342, i_8_1346, i_8_1436, i_8_1450, i_8_1467, i_8_1469, i_8_1492, i_8_1503, i_8_1504, i_8_1539, i_8_1571, i_8_1597, i_8_1622, i_8_1679, i_8_1681, i_8_1746, i_8_1751, i_8_1752, i_8_1753, i_8_1781, i_8_1787, i_8_1789, i_8_1800, i_8_1805, i_8_1817, i_8_1855, i_8_1918, i_8_1948, i_8_1963, i_8_1966, i_8_2108, i_8_2109, i_8_2110, i_8_2139, i_8_2147, i_8_2244, i_8_2270, i_8_2272, i_8_2286, i_8_2290, o_8_152);
	kernel_8_153 k_8_153(i_8_51, i_8_53, i_8_124, i_8_125, i_8_168, i_8_169, i_8_170, i_8_172, i_8_177, i_8_330, i_8_341, i_8_348, i_8_368, i_8_378, i_8_379, i_8_384, i_8_393, i_8_418, i_8_420, i_8_422, i_8_469, i_8_499, i_8_598, i_8_659, i_8_704, i_8_753, i_8_778, i_8_879, i_8_898, i_8_985, i_8_987, i_8_988, i_8_994, i_8_1015, i_8_1040, i_8_1051, i_8_1111, i_8_1131, i_8_1132, i_8_1139, i_8_1140, i_8_1141, i_8_1168, i_8_1228, i_8_1236, i_8_1237, i_8_1261, i_8_1263, i_8_1275, i_8_1276, i_8_1277, i_8_1281, i_8_1284, i_8_1285, i_8_1286, i_8_1331, i_8_1381, i_8_1434, i_8_1446, i_8_1470, i_8_1471, i_8_1474, i_8_1475, i_8_1479, i_8_1482, i_8_1484, i_8_1511, i_8_1520, i_8_1527, i_8_1529, i_8_1536, i_8_1554, i_8_1588, i_8_1590, i_8_1635, i_8_1645, i_8_1654, i_8_1664, i_8_1671, i_8_1672, i_8_1734, i_8_1735, i_8_1762, i_8_1770, i_8_1783, i_8_1808, i_8_1862, i_8_1870, i_8_1969, i_8_1992, i_8_1993, i_8_2013, i_8_2015, i_8_2038, i_8_2048, i_8_2095, i_8_2122, i_8_2146, i_8_2147, i_8_2276, o_8_153);
	kernel_8_154 k_8_154(i_8_28, i_8_47, i_8_64, i_8_72, i_8_77, i_8_111, i_8_181, i_8_226, i_8_308, i_8_319, i_8_320, i_8_388, i_8_398, i_8_506, i_8_536, i_8_551, i_8_559, i_8_571, i_8_572, i_8_578, i_8_579, i_8_586, i_8_587, i_8_596, i_8_603, i_8_611, i_8_630, i_8_631, i_8_634, i_8_640, i_8_649, i_8_652, i_8_659, i_8_680, i_8_707, i_8_748, i_8_793, i_8_794, i_8_837, i_8_844, i_8_845, i_8_855, i_8_859, i_8_874, i_8_882, i_8_969, i_8_973, i_8_991, i_8_1073, i_8_1108, i_8_1128, i_8_1143, i_8_1170, i_8_1180, i_8_1199, i_8_1226, i_8_1243, i_8_1261, i_8_1264, i_8_1328, i_8_1405, i_8_1410, i_8_1459, i_8_1462, i_8_1469, i_8_1472, i_8_1478, i_8_1523, i_8_1536, i_8_1544, i_8_1625, i_8_1648, i_8_1650, i_8_1651, i_8_1682, i_8_1684, i_8_1694, i_8_1703, i_8_1748, i_8_1765, i_8_1777, i_8_1781, i_8_1782, i_8_1819, i_8_1820, i_8_1822, i_8_1823, i_8_1855, i_8_1881, i_8_1909, i_8_1936, i_8_1954, i_8_1994, i_8_2146, i_8_2147, i_8_2170, i_8_2191, i_8_2207, i_8_2225, i_8_2241, o_8_154);
	kernel_8_155 k_8_155(i_8_6, i_8_32, i_8_43, i_8_49, i_8_50, i_8_64, i_8_67, i_8_75, i_8_142, i_8_151, i_8_169, i_8_215, i_8_260, i_8_337, i_8_338, i_8_347, i_8_355, i_8_363, i_8_385, i_8_386, i_8_416, i_8_427, i_8_453, i_8_500, i_8_523, i_8_527, i_8_538, i_8_593, i_8_608, i_8_613, i_8_614, i_8_633, i_8_634, i_8_664, i_8_703, i_8_704, i_8_705, i_8_706, i_8_763, i_8_770, i_8_955, i_8_958, i_8_964, i_8_994, i_8_995, i_8_1078, i_8_1110, i_8_1125, i_8_1139, i_8_1154, i_8_1174, i_8_1175, i_8_1227, i_8_1228, i_8_1262, i_8_1299, i_8_1410, i_8_1417, i_8_1438, i_8_1453, i_8_1456, i_8_1475, i_8_1525, i_8_1531, i_8_1556, i_8_1600, i_8_1624, i_8_1648, i_8_1679, i_8_1682, i_8_1733, i_8_1785, i_8_1818, i_8_1819, i_8_1821, i_8_1824, i_8_1866, i_8_1877, i_8_1957, i_8_1967, i_8_1975, i_8_1995, i_8_2005, i_8_2013, i_8_2048, i_8_2057, i_8_2065, i_8_2094, i_8_2095, i_8_2143, i_8_2147, i_8_2148, i_8_2150, i_8_2157, i_8_2159, i_8_2171, i_8_2183, i_8_2226, i_8_2231, i_8_2266, o_8_155);
	kernel_8_156 k_8_156(i_8_35, i_8_37, i_8_77, i_8_87, i_8_111, i_8_140, i_8_229, i_8_235, i_8_259, i_8_304, i_8_355, i_8_382, i_8_418, i_8_419, i_8_442, i_8_445, i_8_446, i_8_464, i_8_490, i_8_504, i_8_505, i_8_506, i_8_507, i_8_508, i_8_509, i_8_528, i_8_610, i_8_621, i_8_625, i_8_665, i_8_698, i_8_748, i_8_780, i_8_781, i_8_845, i_8_876, i_8_880, i_8_885, i_8_967, i_8_1028, i_8_1030, i_8_1031, i_8_1136, i_8_1158, i_8_1192, i_8_1200, i_8_1201, i_8_1202, i_8_1225, i_8_1269, i_8_1281, i_8_1315, i_8_1325, i_8_1328, i_8_1350, i_8_1355, i_8_1387, i_8_1398, i_8_1399, i_8_1400, i_8_1437, i_8_1450, i_8_1453, i_8_1454, i_8_1537, i_8_1604, i_8_1623, i_8_1630, i_8_1631, i_8_1634, i_8_1650, i_8_1677, i_8_1678, i_8_1679, i_8_1701, i_8_1746, i_8_1751, i_8_1771, i_8_1792, i_8_1793, i_8_1794, i_8_1795, i_8_1855, i_8_1856, i_8_1858, i_8_1876, i_8_1877, i_8_1912, i_8_1980, i_8_1981, i_8_1984, i_8_1985, i_8_1993, i_8_2056, i_8_2057, i_8_2129, i_8_2143, i_8_2144, i_8_2156, i_8_2272, o_8_156);
	kernel_8_157 k_8_157(i_8_25, i_8_33, i_8_72, i_8_96, i_8_97, i_8_214, i_8_215, i_8_220, i_8_241, i_8_286, i_8_295, i_8_301, i_8_348, i_8_361, i_8_367, i_8_376, i_8_385, i_8_421, i_8_445, i_8_457, i_8_467, i_8_484, i_8_485, i_8_525, i_8_555, i_8_592, i_8_593, i_8_610, i_8_611, i_8_616, i_8_630, i_8_715, i_8_718, i_8_719, i_8_760, i_8_763, i_8_764, i_8_772, i_8_799, i_8_838, i_8_889, i_8_925, i_8_952, i_8_991, i_8_1012, i_8_1015, i_8_1016, i_8_1029, i_8_1030, i_8_1114, i_8_1124, i_8_1160, i_8_1237, i_8_1258, i_8_1263, i_8_1264, i_8_1273, i_8_1300, i_8_1305, i_8_1306, i_8_1331, i_8_1344, i_8_1363, i_8_1387, i_8_1438, i_8_1455, i_8_1456, i_8_1544, i_8_1600, i_8_1601, i_8_1632, i_8_1644, i_8_1680, i_8_1735, i_8_1748, i_8_1749, i_8_1754, i_8_1818, i_8_1867, i_8_1869, i_8_1894, i_8_1897, i_8_1903, i_8_1921, i_8_1922, i_8_1967, i_8_1969, i_8_2020, i_8_2056, i_8_2092, i_8_2114, i_8_2131, i_8_2157, i_8_2218, i_8_2266, i_8_2274, i_8_2275, i_8_2292, i_8_2293, i_8_2294, o_8_157);
	kernel_8_158 k_8_158(i_8_6, i_8_76, i_8_78, i_8_79, i_8_114, i_8_157, i_8_159, i_8_204, i_8_205, i_8_240, i_8_241, i_8_249, i_8_256, i_8_259, i_8_301, i_8_312, i_8_313, i_8_327, i_8_348, i_8_366, i_8_429, i_8_453, i_8_499, i_8_507, i_8_553, i_8_570, i_8_574, i_8_597, i_8_600, i_8_606, i_8_660, i_8_665, i_8_687, i_8_690, i_8_771, i_8_777, i_8_778, i_8_783, i_8_849, i_8_885, i_8_943, i_8_993, i_8_1028, i_8_1037, i_8_1048, i_8_1056, i_8_1059, i_8_1077, i_8_1104, i_8_1138, i_8_1146, i_8_1182, i_8_1227, i_8_1228, i_8_1294, i_8_1306, i_8_1371, i_8_1410, i_8_1436, i_8_1455, i_8_1510, i_8_1624, i_8_1626, i_8_1629, i_8_1644, i_8_1653, i_8_1654, i_8_1689, i_8_1705, i_8_1748, i_8_1750, i_8_1753, i_8_1754, i_8_1808, i_8_1823, i_8_1837, i_8_1860, i_8_1861, i_8_1863, i_8_1884, i_8_1887, i_8_1983, i_8_1984, i_8_1986, i_8_2046, i_8_2055, i_8_2058, i_8_2073, i_8_2074, i_8_2076, i_8_2085, i_8_2086, i_8_2141, i_8_2146, i_8_2150, i_8_2157, i_8_2217, i_8_2244, i_8_2274, i_8_2275, o_8_158);
	kernel_8_159 k_8_159(i_8_26, i_8_50, i_8_76, i_8_88, i_8_93, i_8_106, i_8_250, i_8_266, i_8_282, i_8_286, i_8_291, i_8_321, i_8_383, i_8_384, i_8_436, i_8_437, i_8_453, i_8_454, i_8_456, i_8_491, i_8_555, i_8_624, i_8_633, i_8_636, i_8_642, i_8_643, i_8_672, i_8_687, i_8_696, i_8_703, i_8_718, i_8_727, i_8_728, i_8_730, i_8_735, i_8_736, i_8_782, i_8_814, i_8_834, i_8_843, i_8_848, i_8_852, i_8_933, i_8_1074, i_8_1088, i_8_1138, i_8_1185, i_8_1213, i_8_1221, i_8_1222, i_8_1227, i_8_1228, i_8_1236, i_8_1237, i_8_1239, i_8_1266, i_8_1281, i_8_1290, i_8_1309, i_8_1349, i_8_1384, i_8_1390, i_8_1446, i_8_1455, i_8_1545, i_8_1561, i_8_1580, i_8_1617, i_8_1624, i_8_1653, i_8_1654, i_8_1704, i_8_1706, i_8_1723, i_8_1770, i_8_1808, i_8_1825, i_8_1843, i_8_1849, i_8_1860, i_8_1903, i_8_1989, i_8_1992, i_8_1995, i_8_2010, i_8_2019, i_8_2031, i_8_2040, i_8_2084, i_8_2131, i_8_2138, i_8_2147, i_8_2158, i_8_2173, i_8_2194, i_8_2226, i_8_2247, i_8_2263, i_8_2284, i_8_2289, o_8_159);
	kernel_8_160 k_8_160(i_8_31, i_8_34, i_8_35, i_8_46, i_8_52, i_8_53, i_8_59, i_8_80, i_8_94, i_8_95, i_8_98, i_8_115, i_8_184, i_8_232, i_8_233, i_8_304, i_8_314, i_8_329, i_8_349, i_8_381, i_8_425, i_8_454, i_8_455, i_8_503, i_8_552, i_8_556, i_8_557, i_8_614, i_8_696, i_8_698, i_8_706, i_8_956, i_8_967, i_8_968, i_8_992, i_8_994, i_8_1048, i_8_1049, i_8_1052, i_8_1075, i_8_1094, i_8_1110, i_8_1115, i_8_1135, i_8_1179, i_8_1183, i_8_1263, i_8_1271, i_8_1274, i_8_1282, i_8_1291, i_8_1306, i_8_1307, i_8_1325, i_8_1339, i_8_1348, i_8_1352, i_8_1355, i_8_1372, i_8_1388, i_8_1435, i_8_1436, i_8_1437, i_8_1438, i_8_1439, i_8_1506, i_8_1507, i_8_1535, i_8_1625, i_8_1627, i_8_1628, i_8_1636, i_8_1676, i_8_1677, i_8_1678, i_8_1679, i_8_1682, i_8_1750, i_8_1764, i_8_1784, i_8_1807, i_8_1822, i_8_1873, i_8_1876, i_8_1906, i_8_1907, i_8_1963, i_8_1966, i_8_1981, i_8_1982, i_8_2006, i_8_2032, i_8_2050, i_8_2093, i_8_2096, i_8_2109, i_8_2152, i_8_2216, i_8_2281, i_8_2282, o_8_160);
	kernel_8_161 k_8_161(i_8_20, i_8_23, i_8_43, i_8_88, i_8_121, i_8_131, i_8_194, i_8_230, i_8_232, i_8_247, i_8_278, i_8_310, i_8_311, i_8_314, i_8_325, i_8_363, i_8_367, i_8_393, i_8_419, i_8_430, i_8_473, i_8_492, i_8_634, i_8_693, i_8_706, i_8_709, i_8_751, i_8_790, i_8_799, i_8_825, i_8_831, i_8_838, i_8_842, i_8_844, i_8_850, i_8_878, i_8_879, i_8_880, i_8_886, i_8_887, i_8_953, i_8_964, i_8_968, i_8_970, i_8_986, i_8_994, i_8_1016, i_8_1039, i_8_1040, i_8_1048, i_8_1063, i_8_1075, i_8_1076, i_8_1102, i_8_1113, i_8_1127, i_8_1165, i_8_1239, i_8_1240, i_8_1246, i_8_1318, i_8_1336, i_8_1372, i_8_1399, i_8_1407, i_8_1470, i_8_1498, i_8_1528, i_8_1607, i_8_1609, i_8_1641, i_8_1645, i_8_1653, i_8_1690, i_8_1691, i_8_1704, i_8_1708, i_8_1733, i_8_1746, i_8_1751, i_8_1767, i_8_1769, i_8_1870, i_8_1884, i_8_1896, i_8_1906, i_8_1984, i_8_2039, i_8_2042, i_8_2066, i_8_2072, i_8_2075, i_8_2086, i_8_2089, i_8_2119, i_8_2153, i_8_2174, i_8_2227, i_8_2232, i_8_2275, o_8_161);
	kernel_8_162 k_8_162(i_8_23, i_8_25, i_8_138, i_8_139, i_8_140, i_8_141, i_8_143, i_8_194, i_8_228, i_8_282, i_8_286, i_8_287, i_8_318, i_8_320, i_8_398, i_8_404, i_8_440, i_8_504, i_8_580, i_8_583, i_8_641, i_8_642, i_8_694, i_8_727, i_8_823, i_8_858, i_8_859, i_8_873, i_8_877, i_8_882, i_8_885, i_8_972, i_8_973, i_8_974, i_8_976, i_8_977, i_8_979, i_8_980, i_8_1030, i_8_1040, i_8_1187, i_8_1198, i_8_1238, i_8_1362, i_8_1367, i_8_1410, i_8_1426, i_8_1427, i_8_1440, i_8_1443, i_8_1444, i_8_1447, i_8_1462, i_8_1470, i_8_1471, i_8_1525, i_8_1526, i_8_1529, i_8_1534, i_8_1600, i_8_1604, i_8_1606, i_8_1641, i_8_1669, i_8_1679, i_8_1697, i_8_1718, i_8_1726, i_8_1777, i_8_1808, i_8_1905, i_8_1944, i_8_1965, i_8_1966, i_8_1967, i_8_1969, i_8_1970, i_8_1975, i_8_1983, i_8_2011, i_8_2031, i_8_2052, i_8_2055, i_8_2056, i_8_2057, i_8_2109, i_8_2110, i_8_2112, i_8_2137, i_8_2154, i_8_2155, i_8_2159, i_8_2172, i_8_2173, i_8_2176, i_8_2232, i_8_2233, i_8_2234, i_8_2246, i_8_2249, o_8_162);
	kernel_8_163 k_8_163(i_8_103, i_8_140, i_8_220, i_8_226, i_8_230, i_8_247, i_8_256, i_8_262, i_8_299, i_8_304, i_8_314, i_8_316, i_8_326, i_8_363, i_8_367, i_8_381, i_8_418, i_8_428, i_8_454, i_8_455, i_8_553, i_8_581, i_8_582, i_8_584, i_8_599, i_8_635, i_8_793, i_8_823, i_8_839, i_8_840, i_8_844, i_8_845, i_8_859, i_8_874, i_8_881, i_8_882, i_8_891, i_8_994, i_8_1145, i_8_1147, i_8_1226, i_8_1229, i_8_1268, i_8_1282, i_8_1286, i_8_1319, i_8_1399, i_8_1403, i_8_1432, i_8_1435, i_8_1436, i_8_1438, i_8_1463, i_8_1470, i_8_1510, i_8_1562, i_8_1574, i_8_1668, i_8_1688, i_8_1690, i_8_1704, i_8_1774, i_8_1779, i_8_1786, i_8_1787, i_8_1805, i_8_1810, i_8_1819, i_8_1894, i_8_1963, i_8_1971, i_8_1975, i_8_1981, i_8_1983, i_8_1984, i_8_1994, i_8_2053, i_8_2056, i_8_2107, i_8_2108, i_8_2110, i_8_2134, i_8_2145, i_8_2146, i_8_2147, i_8_2148, i_8_2149, i_8_2155, i_8_2156, i_8_2158, i_8_2159, i_8_2169, i_8_2170, i_8_2223, i_8_2228, i_8_2229, i_8_2230, i_8_2234, i_8_2248, i_8_2263, o_8_163);
	kernel_8_164 k_8_164(i_8_21, i_8_33, i_8_34, i_8_35, i_8_85, i_8_93, i_8_96, i_8_156, i_8_165, i_8_202, i_8_220, i_8_222, i_8_223, i_8_255, i_8_262, i_8_277, i_8_291, i_8_300, i_8_301, i_8_345, i_8_393, i_8_420, i_8_474, i_8_475, i_8_493, i_8_500, i_8_501, i_8_503, i_8_547, i_8_552, i_8_555, i_8_588, i_8_589, i_8_624, i_8_657, i_8_670, i_8_715, i_8_716, i_8_723, i_8_759, i_8_768, i_8_781, i_8_823, i_8_877, i_8_1011, i_8_1029, i_8_1114, i_8_1115, i_8_1119, i_8_1128, i_8_1156, i_8_1159, i_8_1191, i_8_1254, i_8_1257, i_8_1258, i_8_1282, i_8_1344, i_8_1345, i_8_1347, i_8_1452, i_8_1453, i_8_1542, i_8_1551, i_8_1555, i_8_1587, i_8_1596, i_8_1597, i_8_1600, i_8_1611, i_8_1626, i_8_1651, i_8_1668, i_8_1680, i_8_1682, i_8_1708, i_8_1743, i_8_1760, i_8_1761, i_8_1762, i_8_1782, i_8_1804, i_8_1806, i_8_1839, i_8_1849, i_8_1867, i_8_1893, i_8_1894, i_8_1952, i_8_1992, i_8_1995, i_8_2031, i_8_2049, i_8_2110, i_8_2128, i_8_2190, i_8_2214, i_8_2215, i_8_2287, i_8_2289, o_8_164);
	kernel_8_165 k_8_165(i_8_20, i_8_38, i_8_44, i_8_106, i_8_184, i_8_214, i_8_226, i_8_257, i_8_263, i_8_270, i_8_288, i_8_289, i_8_297, i_8_344, i_8_353, i_8_370, i_8_380, i_8_388, i_8_416, i_8_443, i_8_452, i_8_462, i_8_475, i_8_535, i_8_625, i_8_627, i_8_638, i_8_661, i_8_663, i_8_665, i_8_695, i_8_696, i_8_713, i_8_724, i_8_756, i_8_759, i_8_792, i_8_793, i_8_817, i_8_869, i_8_875, i_8_876, i_8_927, i_8_971, i_8_982, i_8_988, i_8_992, i_8_999, i_8_1051, i_8_1110, i_8_1127, i_8_1156, i_8_1161, i_8_1217, i_8_1224, i_8_1236, i_8_1246, i_8_1252, i_8_1271, i_8_1281, i_8_1300, i_8_1341, i_8_1363, i_8_1367, i_8_1424, i_8_1427, i_8_1453, i_8_1469, i_8_1504, i_8_1560, i_8_1603, i_8_1604, i_8_1613, i_8_1631, i_8_1674, i_8_1687, i_8_1699, i_8_1714, i_8_1733, i_8_1750, i_8_1758, i_8_1762, i_8_1780, i_8_1791, i_8_1807, i_8_1838, i_8_1854, i_8_1920, i_8_1996, i_8_2018, i_8_2054, i_8_2056, i_8_2124, i_8_2129, i_8_2170, i_8_2171, i_8_2188, i_8_2223, i_8_2261, i_8_2270, o_8_165);
	kernel_8_166 k_8_166(i_8_13, i_8_28, i_8_44, i_8_79, i_8_80, i_8_106, i_8_115, i_8_140, i_8_185, i_8_227, i_8_320, i_8_322, i_8_323, i_8_349, i_8_391, i_8_401, i_8_421, i_8_431, i_8_455, i_8_486, i_8_500, i_8_536, i_8_556, i_8_557, i_8_572, i_8_607, i_8_623, i_8_635, i_8_653, i_8_655, i_8_656, i_8_670, i_8_674, i_8_702, i_8_703, i_8_826, i_8_827, i_8_838, i_8_839, i_8_877, i_8_881, i_8_896, i_8_956, i_8_970, i_8_971, i_8_991, i_8_1055, i_8_1111, i_8_1154, i_8_1202, i_8_1300, i_8_1301, i_8_1331, i_8_1336, i_8_1337, i_8_1366, i_8_1367, i_8_1400, i_8_1402, i_8_1435, i_8_1465, i_8_1474, i_8_1489, i_8_1493, i_8_1510, i_8_1517, i_8_1525, i_8_1526, i_8_1529, i_8_1548, i_8_1550, i_8_1553, i_8_1574, i_8_1622, i_8_1625, i_8_1630, i_8_1634, i_8_1651, i_8_1672, i_8_1753, i_8_1771, i_8_1774, i_8_1784, i_8_1795, i_8_1824, i_8_1825, i_8_1849, i_8_1886, i_8_1888, i_8_1937, i_8_1960, i_8_1968, i_8_1975, i_8_1995, i_8_2057, i_8_2072, i_8_2125, i_8_2146, i_8_2242, i_8_2285, o_8_166);
	kernel_8_167 k_8_167(i_8_76, i_8_115, i_8_137, i_8_184, i_8_279, i_8_299, i_8_320, i_8_322, i_8_392, i_8_423, i_8_427, i_8_429, i_8_483, i_8_487, i_8_489, i_8_496, i_8_553, i_8_574, i_8_580, i_8_581, i_8_588, i_8_606, i_8_607, i_8_630, i_8_633, i_8_640, i_8_641, i_8_651, i_8_655, i_8_661, i_8_676, i_8_703, i_8_706, i_8_742, i_8_744, i_8_755, i_8_841, i_8_842, i_8_895, i_8_971, i_8_973, i_8_974, i_8_1010, i_8_1020, i_8_1036, i_8_1039, i_8_1107, i_8_1109, i_8_1200, i_8_1201, i_8_1246, i_8_1247, i_8_1264, i_8_1267, i_8_1297, i_8_1315, i_8_1351, i_8_1363, i_8_1365, i_8_1382, i_8_1383, i_8_1416, i_8_1434, i_8_1435, i_8_1436, i_8_1438, i_8_1461, i_8_1462, i_8_1465, i_8_1469, i_8_1477, i_8_1487, i_8_1512, i_8_1547, i_8_1607, i_8_1630, i_8_1638, i_8_1707, i_8_1720, i_8_1802, i_8_1809, i_8_1825, i_8_1837, i_8_1838, i_8_1840, i_8_1912, i_8_1957, i_8_1981, i_8_1992, i_8_1994, i_8_1997, i_8_2119, i_8_2146, i_8_2147, i_8_2169, i_8_2170, i_8_2227, i_8_2247, i_8_2248, i_8_2289, o_8_167);
	kernel_8_168 k_8_168(i_8_19, i_8_20, i_8_58, i_8_78, i_8_79, i_8_94, i_8_114, i_8_289, i_8_298, i_8_325, i_8_353, i_8_360, i_8_370, i_8_383, i_8_417, i_8_459, i_8_460, i_8_461, i_8_482, i_8_490, i_8_526, i_8_549, i_8_553, i_8_615, i_8_621, i_8_622, i_8_623, i_8_627, i_8_628, i_8_629, i_8_661, i_8_667, i_8_696, i_8_703, i_8_712, i_8_779, i_8_792, i_8_830, i_8_832, i_8_841, i_8_885, i_8_938, i_8_971, i_8_977, i_8_990, i_8_992, i_8_997, i_8_1010, i_8_1110, i_8_1118, i_8_1127, i_8_1128, i_8_1225, i_8_1234, i_8_1278, i_8_1280, i_8_1316, i_8_1324, i_8_1341, i_8_1408, i_8_1411, i_8_1449, i_8_1450, i_8_1451, i_8_1504, i_8_1532, i_8_1533, i_8_1548, i_8_1549, i_8_1553, i_8_1594, i_8_1650, i_8_1749, i_8_1750, i_8_1758, i_8_1759, i_8_1775, i_8_1801, i_8_1838, i_8_1864, i_8_1865, i_8_1891, i_8_1909, i_8_1919, i_8_1963, i_8_1967, i_8_1985, i_8_1990, i_8_2106, i_8_2107, i_8_2126, i_8_2141, i_8_2142, i_8_2188, i_8_2224, i_8_2269, i_8_2270, i_8_2273, i_8_2286, i_8_2288, o_8_168);
	kernel_8_169 k_8_169(i_8_10, i_8_80, i_8_226, i_8_230, i_8_233, i_8_260, i_8_298, i_8_301, i_8_314, i_8_316, i_8_367, i_8_419, i_8_469, i_8_526, i_8_530, i_8_604, i_8_605, i_8_607, i_8_616, i_8_629, i_8_649, i_8_657, i_8_665, i_8_691, i_8_692, i_8_696, i_8_697, i_8_700, i_8_701, i_8_705, i_8_709, i_8_836, i_8_843, i_8_844, i_8_855, i_8_863, i_8_881, i_8_890, i_8_976, i_8_988, i_8_989, i_8_994, i_8_1006, i_8_1043, i_8_1052, i_8_1060, i_8_1097, i_8_1105, i_8_1150, i_8_1168, i_8_1219, i_8_1297, i_8_1325, i_8_1351, i_8_1411, i_8_1434, i_8_1462, i_8_1492, i_8_1504, i_8_1544, i_8_1551, i_8_1555, i_8_1565, i_8_1567, i_8_1609, i_8_1627, i_8_1628, i_8_1652, i_8_1663, i_8_1669, i_8_1674, i_8_1693, i_8_1709, i_8_1766, i_8_1780, i_8_1792, i_8_1798, i_8_1826, i_8_1837, i_8_1855, i_8_1858, i_8_1867, i_8_1880, i_8_1885, i_8_1888, i_8_1894, i_8_1897, i_8_1954, i_8_1990, i_8_2015, i_8_2071, i_8_2077, i_8_2078, i_8_2093, i_8_2095, i_8_2105, i_8_2136, i_8_2170, i_8_2259, i_8_2275, o_8_169);
	kernel_8_170 k_8_170(i_8_3, i_8_6, i_8_9, i_8_54, i_8_115, i_8_210, i_8_219, i_8_249, i_8_258, i_8_295, i_8_298, i_8_350, i_8_358, i_8_363, i_8_365, i_8_421, i_8_448, i_8_454, i_8_466, i_8_490, i_8_516, i_8_523, i_8_574, i_8_598, i_8_601, i_8_606, i_8_607, i_8_610, i_8_661, i_8_672, i_8_699, i_8_717, i_8_718, i_8_726, i_8_736, i_8_789, i_8_813, i_8_816, i_8_817, i_8_835, i_8_836, i_8_842, i_8_852, i_8_853, i_8_889, i_8_1015, i_8_1029, i_8_1031, i_8_1044, i_8_1074, i_8_1078, i_8_1087, i_8_1156, i_8_1204, i_8_1285, i_8_1308, i_8_1317, i_8_1392, i_8_1393, i_8_1394, i_8_1437, i_8_1446, i_8_1500, i_8_1636, i_8_1662, i_8_1695, i_8_1699, i_8_1763, i_8_1798, i_8_1808, i_8_1824, i_8_1848, i_8_1851, i_8_1858, i_8_1866, i_8_1870, i_8_1879, i_8_1881, i_8_1897, i_8_1920, i_8_2031, i_8_2059, i_8_2067, i_8_2068, i_8_2073, i_8_2074, i_8_2076, i_8_2077, i_8_2092, i_8_2112, i_8_2118, i_8_2121, i_8_2122, i_8_2154, i_8_2215, i_8_2235, i_8_2246, i_8_2283, i_8_2284, i_8_2293, o_8_170);
	kernel_8_171 k_8_171(i_8_53, i_8_58, i_8_62, i_8_83, i_8_115, i_8_136, i_8_142, i_8_143, i_8_147, i_8_195, i_8_225, i_8_227, i_8_238, i_8_262, i_8_364, i_8_418, i_8_491, i_8_493, i_8_555, i_8_556, i_8_557, i_8_575, i_8_781, i_8_782, i_8_786, i_8_964, i_8_976, i_8_993, i_8_994, i_8_996, i_8_1008, i_8_1051, i_8_1110, i_8_1111, i_8_1120, i_8_1121, i_8_1124, i_8_1191, i_8_1263, i_8_1281, i_8_1282, i_8_1284, i_8_1285, i_8_1305, i_8_1306, i_8_1307, i_8_1315, i_8_1330, i_8_1331, i_8_1344, i_8_1408, i_8_1409, i_8_1411, i_8_1435, i_8_1436, i_8_1437, i_8_1470, i_8_1474, i_8_1506, i_8_1507, i_8_1509, i_8_1545, i_8_1565, i_8_1573, i_8_1574, i_8_1590, i_8_1629, i_8_1653, i_8_1655, i_8_1682, i_8_1687, i_8_1700, i_8_1723, i_8_1740, i_8_1747, i_8_1804, i_8_1807, i_8_1875, i_8_1876, i_8_1888, i_8_1903, i_8_1925, i_8_1990, i_8_1991, i_8_1992, i_8_2005, i_8_2093, i_8_2102, i_8_2133, i_8_2147, i_8_2152, i_8_2155, i_8_2214, i_8_2215, i_8_2216, i_8_2242, i_8_2245, i_8_2246, i_8_2249, i_8_2260, o_8_171);
	kernel_8_172 k_8_172(i_8_53, i_8_59, i_8_62, i_8_63, i_8_98, i_8_139, i_8_143, i_8_188, i_8_259, i_8_260, i_8_287, i_8_304, i_8_346, i_8_360, i_8_366, i_8_376, i_8_385, i_8_422, i_8_438, i_8_448, i_8_457, i_8_460, i_8_461, i_8_485, i_8_502, i_8_508, i_8_511, i_8_512, i_8_529, i_8_587, i_8_599, i_8_749, i_8_763, i_8_764, i_8_790, i_8_824, i_8_851, i_8_854, i_8_880, i_8_958, i_8_994, i_8_995, i_8_997, i_8_1016, i_8_1051, i_8_1052, i_8_1075, i_8_1078, i_8_1079, i_8_1094, i_8_1103, i_8_1105, i_8_1114, i_8_1124, i_8_1130, i_8_1192, i_8_1193, i_8_1267, i_8_1306, i_8_1307, i_8_1310, i_8_1315, i_8_1350, i_8_1391, i_8_1394, i_8_1407, i_8_1508, i_8_1546, i_8_1553, i_8_1573, i_8_1574, i_8_1633, i_8_1653, i_8_1681, i_8_1690, i_8_1724, i_8_1726, i_8_1727, i_8_1753, i_8_1763, i_8_1837, i_8_1859, i_8_1862, i_8_1870, i_8_1879, i_8_1880, i_8_1888, i_8_1907, i_8_2002, i_8_2006, i_8_2033, i_8_2139, i_8_2154, i_8_2155, i_8_2170, i_8_2187, i_8_2197, i_8_2215, i_8_2237, i_8_2247, o_8_172);
	kernel_8_173 k_8_173(i_8_25, i_8_40, i_8_42, i_8_250, i_8_257, i_8_277, i_8_303, i_8_367, i_8_374, i_8_426, i_8_445, i_8_471, i_8_493, i_8_499, i_8_552, i_8_553, i_8_555, i_8_592, i_8_593, i_8_597, i_8_604, i_8_610, i_8_635, i_8_653, i_8_673, i_8_674, i_8_677, i_8_718, i_8_719, i_8_729, i_8_841, i_8_852, i_8_853, i_8_868, i_8_877, i_8_880, i_8_881, i_8_958, i_8_959, i_8_994, i_8_1035, i_8_1075, i_8_1078, i_8_1105, i_8_1113, i_8_1114, i_8_1186, i_8_1201, i_8_1203, i_8_1227, i_8_1230, i_8_1246, i_8_1263, i_8_1320, i_8_1345, i_8_1410, i_8_1411, i_8_1423, i_8_1440, i_8_1482, i_8_1483, i_8_1485, i_8_1488, i_8_1498, i_8_1529, i_8_1534, i_8_1536, i_8_1600, i_8_1601, i_8_1605, i_8_1644, i_8_1705, i_8_1715, i_8_1749, i_8_1813, i_8_1826, i_8_1853, i_8_1869, i_8_1870, i_8_1875, i_8_1878, i_8_1888, i_8_1918, i_8_1921, i_8_1951, i_8_1965, i_8_1974, i_8_1975, i_8_1983, i_8_1987, i_8_1997, i_8_2007, i_8_2049, i_8_2065, i_8_2068, i_8_2229, i_8_2231, i_8_2239, i_8_2242, i_8_2257, o_8_173);
	kernel_8_174 k_8_174(i_8_9, i_8_10, i_8_73, i_8_91, i_8_102, i_8_112, i_8_143, i_8_165, i_8_181, i_8_205, i_8_208, i_8_230, i_8_238, i_8_248, i_8_265, i_8_274, i_8_284, i_8_292, i_8_324, i_8_343, i_8_366, i_8_371, i_8_491, i_8_537, i_8_568, i_8_609, i_8_625, i_8_626, i_8_631, i_8_640, i_8_662, i_8_688, i_8_705, i_8_724, i_8_780, i_8_811, i_8_838, i_8_878, i_8_929, i_8_940, i_8_970, i_8_982, i_8_1009, i_8_1019, i_8_1053, i_8_1073, i_8_1100, i_8_1102, i_8_1104, i_8_1113, i_8_1152, i_8_1171, i_8_1172, i_8_1173, i_8_1192, i_8_1245, i_8_1258, i_8_1281, i_8_1297, i_8_1306, i_8_1312, i_8_1336, i_8_1368, i_8_1404, i_8_1475, i_8_1539, i_8_1554, i_8_1589, i_8_1668, i_8_1672, i_8_1675, i_8_1687, i_8_1690, i_8_1733, i_8_1758, i_8_1759, i_8_1789, i_8_1804, i_8_1831, i_8_1842, i_8_1846, i_8_1868, i_8_1873, i_8_1881, i_8_1889, i_8_1907, i_8_1937, i_8_1992, i_8_2070, i_8_2100, i_8_2129, i_8_2150, i_8_2151, i_8_2161, i_8_2205, i_8_2223, i_8_2241, i_8_2261, i_8_2287, i_8_2296, o_8_174);
	kernel_8_175 k_8_175(i_8_42, i_8_176, i_8_189, i_8_190, i_8_242, i_8_246, i_8_311, i_8_366, i_8_369, i_8_394, i_8_462, i_8_466, i_8_525, i_8_535, i_8_555, i_8_595, i_8_596, i_8_613, i_8_660, i_8_661, i_8_696, i_8_702, i_8_706, i_8_729, i_8_730, i_8_747, i_8_748, i_8_814, i_8_825, i_8_837, i_8_838, i_8_859, i_8_915, i_8_940, i_8_1126, i_8_1174, i_8_1182, i_8_1183, i_8_1198, i_8_1239, i_8_1241, i_8_1273, i_8_1282, i_8_1284, i_8_1299, i_8_1306, i_8_1318, i_8_1338, i_8_1434, i_8_1435, i_8_1442, i_8_1471, i_8_1479, i_8_1498, i_8_1509, i_8_1524, i_8_1525, i_8_1533, i_8_1540, i_8_1546, i_8_1606, i_8_1633, i_8_1641, i_8_1642, i_8_1647, i_8_1648, i_8_1687, i_8_1818, i_8_1821, i_8_1854, i_8_1858, i_8_1909, i_8_1915, i_8_1917, i_8_1930, i_8_1948, i_8_1962, i_8_1969, i_8_1992, i_8_2038, i_8_2047, i_8_2058, i_8_2065, i_8_2066, i_8_2089, i_8_2091, i_8_2119, i_8_2122, i_8_2136, i_8_2170, i_8_2172, i_8_2173, i_8_2200, i_8_2218, i_8_2221, i_8_2233, i_8_2248, i_8_2253, i_8_2274, i_8_2286, o_8_175);
	kernel_8_176 k_8_176(i_8_7, i_8_35, i_8_78, i_8_84, i_8_87, i_8_88, i_8_135, i_8_191, i_8_230, i_8_231, i_8_233, i_8_242, i_8_249, i_8_259, i_8_260, i_8_264, i_8_267, i_8_285, i_8_340, i_8_381, i_8_395, i_8_462, i_8_464, i_8_466, i_8_489, i_8_490, i_8_553, i_8_556, i_8_592, i_8_599, i_8_673, i_8_674, i_8_690, i_8_691, i_8_698, i_8_717, i_8_719, i_8_736, i_8_737, i_8_825, i_8_838, i_8_895, i_8_927, i_8_971, i_8_991, i_8_993, i_8_994, i_8_995, i_8_997, i_8_998, i_8_1047, i_8_1056, i_8_1060, i_8_1131, i_8_1132, i_8_1133, i_8_1137, i_8_1139, i_8_1186, i_8_1203, i_8_1204, i_8_1205, i_8_1236, i_8_1266, i_8_1293, i_8_1306, i_8_1315, i_8_1365, i_8_1385, i_8_1446, i_8_1457, i_8_1475, i_8_1547, i_8_1606, i_8_1623, i_8_1797, i_8_1798, i_8_1844, i_8_1911, i_8_1916, i_8_1918, i_8_1922, i_8_1981, i_8_1983, i_8_1985, i_8_2005, i_8_2053, i_8_2055, i_8_2059, i_8_2060, i_8_2069, i_8_2100, i_8_2145, i_8_2156, i_8_2175, i_8_2193, i_8_2195, i_8_2226, i_8_2263, i_8_2291, o_8_176);
	kernel_8_177 k_8_177(i_8_54, i_8_77, i_8_242, i_8_256, i_8_329, i_8_337, i_8_344, i_8_347, i_8_377, i_8_480, i_8_483, i_8_523, i_8_525, i_8_527, i_8_553, i_8_608, i_8_634, i_8_672, i_8_679, i_8_688, i_8_689, i_8_760, i_8_762, i_8_763, i_8_764, i_8_787, i_8_796, i_8_930, i_8_944, i_8_986, i_8_1030, i_8_1048, i_8_1049, i_8_1050, i_8_1051, i_8_1093, i_8_1112, i_8_1124, i_8_1227, i_8_1229, i_8_1236, i_8_1237, i_8_1268, i_8_1274, i_8_1281, i_8_1286, i_8_1295, i_8_1305, i_8_1307, i_8_1309, i_8_1317, i_8_1323, i_8_1328, i_8_1412, i_8_1435, i_8_1439, i_8_1537, i_8_1546, i_8_1547, i_8_1624, i_8_1643, i_8_1651, i_8_1679, i_8_1682, i_8_1696, i_8_1700, i_8_1720, i_8_1723, i_8_1724, i_8_1733, i_8_1742, i_8_1744, i_8_1745, i_8_1749, i_8_1750, i_8_1762, i_8_1763, i_8_1822, i_8_1832, i_8_1876, i_8_1877, i_8_1889, i_8_1903, i_8_1981, i_8_1984, i_8_1985, i_8_2041, i_8_2048, i_8_2057, i_8_2075, i_8_2084, i_8_2093, i_8_2148, i_8_2158, i_8_2164, i_8_2174, i_8_2216, i_8_2219, i_8_2230, i_8_2263, o_8_177);
	kernel_8_178 k_8_178(i_8_14, i_8_31, i_8_32, i_8_51, i_8_52, i_8_55, i_8_59, i_8_77, i_8_201, i_8_229, i_8_255, i_8_256, i_8_378, i_8_385, i_8_387, i_8_388, i_8_390, i_8_391, i_8_392, i_8_415, i_8_417, i_8_426, i_8_450, i_8_493, i_8_508, i_8_509, i_8_534, i_8_536, i_8_608, i_8_630, i_8_634, i_8_658, i_8_676, i_8_748, i_8_750, i_8_752, i_8_880, i_8_1010, i_8_1030, i_8_1127, i_8_1128, i_8_1129, i_8_1130, i_8_1200, i_8_1228, i_8_1234, i_8_1261, i_8_1282, i_8_1289, i_8_1328, i_8_1355, i_8_1358, i_8_1385, i_8_1405, i_8_1476, i_8_1477, i_8_1478, i_8_1479, i_8_1480, i_8_1486, i_8_1490, i_8_1506, i_8_1510, i_8_1540, i_8_1548, i_8_1550, i_8_1559, i_8_1603, i_8_1605, i_8_1607, i_8_1627, i_8_1677, i_8_1713, i_8_1810, i_8_1813, i_8_1822, i_8_1836, i_8_1841, i_8_1873, i_8_1882, i_8_1890, i_8_1891, i_8_1892, i_8_1893, i_8_1894, i_8_1895, i_8_1939, i_8_1984, i_8_1996, i_8_2053, i_8_2057, i_8_2089, i_8_2146, i_8_2147, i_8_2150, i_8_2151, i_8_2155, i_8_2261, i_8_2263, i_8_2276, o_8_178);
	kernel_8_179 k_8_179(i_8_30, i_8_31, i_8_40, i_8_51, i_8_75, i_8_78, i_8_81, i_8_102, i_8_120, i_8_165, i_8_166, i_8_363, i_8_364, i_8_373, i_8_426, i_8_450, i_8_492, i_8_582, i_8_588, i_8_607, i_8_612, i_8_633, i_8_654, i_8_660, i_8_665, i_8_676, i_8_696, i_8_699, i_8_700, i_8_714, i_8_723, i_8_754, i_8_804, i_8_807, i_8_822, i_8_825, i_8_832, i_8_841, i_8_865, i_8_877, i_8_930, i_8_941, i_8_964, i_8_966, i_8_993, i_8_994, i_8_1050, i_8_1056, i_8_1065, i_8_1071, i_8_1093, i_8_1108, i_8_1111, i_8_1138, i_8_1182, i_8_1201, i_8_1217, i_8_1273, i_8_1281, i_8_1326, i_8_1337, i_8_1351, i_8_1359, i_8_1372, i_8_1386, i_8_1432, i_8_1515, i_8_1542, i_8_1545, i_8_1563, i_8_1565, i_8_1587, i_8_1621, i_8_1632, i_8_1668, i_8_1677, i_8_1698, i_8_1699, i_8_1704, i_8_1716, i_8_1747, i_8_1752, i_8_1804, i_8_1819, i_8_1821, i_8_1845, i_8_1946, i_8_1981, i_8_1992, i_8_1995, i_8_1997, i_8_2045, i_8_2115, i_8_2118, i_8_2146, i_8_2149, i_8_2190, i_8_2226, i_8_2235, i_8_2259, o_8_179);
	kernel_8_180 k_8_180(i_8_39, i_8_76, i_8_85, i_8_138, i_8_139, i_8_169, i_8_183, i_8_190, i_8_222, i_8_226, i_8_300, i_8_318, i_8_333, i_8_360, i_8_363, i_8_382, i_8_384, i_8_389, i_8_400, i_8_507, i_8_508, i_8_510, i_8_525, i_8_571, i_8_591, i_8_606, i_8_631, i_8_659, i_8_672, i_8_678, i_8_679, i_8_695, i_8_697, i_8_841, i_8_844, i_8_876, i_8_895, i_8_955, i_8_1039, i_8_1056, i_8_1102, i_8_1105, i_8_1156, i_8_1166, i_8_1246, i_8_1276, i_8_1282, i_8_1304, i_8_1306, i_8_1317, i_8_1318, i_8_1321, i_8_1327, i_8_1330, i_8_1339, i_8_1383, i_8_1423, i_8_1426, i_8_1438, i_8_1461, i_8_1464, i_8_1506, i_8_1509, i_8_1511, i_8_1516, i_8_1519, i_8_1606, i_8_1630, i_8_1632, i_8_1633, i_8_1636, i_8_1642, i_8_1651, i_8_1681, i_8_1686, i_8_1687, i_8_1722, i_8_1723, i_8_1749, i_8_1770, i_8_1781, i_8_1794, i_8_1837, i_8_1849, i_8_1858, i_8_1890, i_8_1938, i_8_1939, i_8_1956, i_8_1957, i_8_1965, i_8_1996, i_8_2054, i_8_2059, i_8_2155, i_8_2174, i_8_2233, i_8_2244, i_8_2262, i_8_2272, o_8_180);
	kernel_8_181 k_8_181(i_8_38, i_8_65, i_8_86, i_8_143, i_8_163, i_8_184, i_8_190, i_8_230, i_8_300, i_8_305, i_8_334, i_8_347, i_8_362, i_8_364, i_8_382, i_8_416, i_8_429, i_8_442, i_8_451, i_8_454, i_8_493, i_8_524, i_8_536, i_8_572, i_8_611, i_8_653, i_8_658, i_8_662, i_8_665, i_8_680, i_8_693, i_8_696, i_8_698, i_8_699, i_8_704, i_8_706, i_8_710, i_8_716, i_8_751, i_8_773, i_8_799, i_8_823, i_8_850, i_8_866, i_8_881, i_8_964, i_8_965, i_8_967, i_8_977, i_8_1103, i_8_1180, i_8_1181, i_8_1192, i_8_1198, i_8_1226, i_8_1247, i_8_1266, i_8_1267, i_8_1283, i_8_1289, i_8_1295, i_8_1318, i_8_1328, i_8_1344, i_8_1364, i_8_1372, i_8_1400, i_8_1403, i_8_1404, i_8_1408, i_8_1410, i_8_1438, i_8_1450, i_8_1453, i_8_1562, i_8_1564, i_8_1655, i_8_1681, i_8_1690, i_8_1706, i_8_1777, i_8_1780, i_8_1784, i_8_1792, i_8_1825, i_8_1886, i_8_1903, i_8_1907, i_8_1975, i_8_1981, i_8_1993, i_8_1996, i_8_2056, i_8_2075, i_8_2146, i_8_2156, i_8_2165, i_8_2197, i_8_2229, i_8_2257, o_8_181);
	kernel_8_182 k_8_182(i_8_0, i_8_1, i_8_3, i_8_73, i_8_81, i_8_82, i_8_111, i_8_112, i_8_153, i_8_198, i_8_227, i_8_243, i_8_279, i_8_283, i_8_318, i_8_342, i_8_345, i_8_363, i_8_364, i_8_434, i_8_436, i_8_450, i_8_486, i_8_568, i_8_604, i_8_626, i_8_630, i_8_666, i_8_673, i_8_705, i_8_710, i_8_729, i_8_811, i_8_829, i_8_832, i_8_833, i_8_865, i_8_892, i_8_992, i_8_1028, i_8_1030, i_8_1033, i_8_1035, i_8_1081, i_8_1091, i_8_1172, i_8_1182, i_8_1198, i_8_1228, i_8_1233, i_8_1270, i_8_1293, i_8_1296, i_8_1299, i_8_1314, i_8_1351, i_8_1386, i_8_1404, i_8_1434, i_8_1506, i_8_1561, i_8_1587, i_8_1633, i_8_1641, i_8_1677, i_8_1720, i_8_1746, i_8_1749, i_8_1777, i_8_1780, i_8_1791, i_8_1801, i_8_1804, i_8_1813, i_8_1845, i_8_1846, i_8_1881, i_8_1890, i_8_1893, i_8_1912, i_8_1923, i_8_1935, i_8_1966, i_8_1971, i_8_1980, i_8_1992, i_8_2025, i_8_2034, i_8_2035, i_8_2055, i_8_2074, i_8_2115, i_8_2116, i_8_2128, i_8_2133, i_8_2134, i_8_2142, i_8_2145, i_8_2157, i_8_2274, o_8_182);
	kernel_8_183 k_8_183(i_8_1, i_8_95, i_8_103, i_8_104, i_8_106, i_8_143, i_8_214, i_8_219, i_8_220, i_8_243, i_8_244, i_8_265, i_8_310, i_8_346, i_8_377, i_8_395, i_8_419, i_8_422, i_8_427, i_8_438, i_8_440, i_8_446, i_8_460, i_8_474, i_8_484, i_8_505, i_8_522, i_8_584, i_8_599, i_8_627, i_8_689, i_8_691, i_8_706, i_8_707, i_8_718, i_8_780, i_8_872, i_8_926, i_8_931, i_8_932, i_8_978, i_8_1021, i_8_1030, i_8_1070, i_8_1074, i_8_1107, i_8_1108, i_8_1137, i_8_1159, i_8_1233, i_8_1265, i_8_1267, i_8_1364, i_8_1376, i_8_1382, i_8_1414, i_8_1434, i_8_1453, i_8_1531, i_8_1532, i_8_1533, i_8_1539, i_8_1548, i_8_1555, i_8_1592, i_8_1633, i_8_1642, i_8_1648, i_8_1677, i_8_1703, i_8_1706, i_8_1723, i_8_1758, i_8_1761, i_8_1819, i_8_1857, i_8_1889, i_8_1918, i_8_1963, i_8_2003, i_8_2010, i_8_2011, i_8_2028, i_8_2049, i_8_2057, i_8_2093, i_8_2114, i_8_2153, i_8_2154, i_8_2156, i_8_2165, i_8_2182, i_8_2183, i_8_2190, i_8_2214, i_8_2240, i_8_2270, i_8_2273, i_8_2294, i_8_2300, o_8_183);
	kernel_8_184 k_8_184(i_8_33, i_8_102, i_8_105, i_8_107, i_8_154, i_8_158, i_8_247, i_8_302, i_8_348, i_8_349, i_8_363, i_8_364, i_8_428, i_8_621, i_8_622, i_8_623, i_8_624, i_8_632, i_8_660, i_8_662, i_8_687, i_8_688, i_8_692, i_8_699, i_8_723, i_8_780, i_8_781, i_8_782, i_8_822, i_8_824, i_8_825, i_8_840, i_8_867, i_8_869, i_8_870, i_8_871, i_8_872, i_8_886, i_8_967, i_8_1008, i_8_1011, i_8_1026, i_8_1054, i_8_1056, i_8_1058, i_8_1060, i_8_1108, i_8_1192, i_8_1272, i_8_1274, i_8_1305, i_8_1306, i_8_1307, i_8_1341, i_8_1342, i_8_1407, i_8_1408, i_8_1409, i_8_1411, i_8_1431, i_8_1434, i_8_1437, i_8_1439, i_8_1449, i_8_1474, i_8_1625, i_8_1641, i_8_1642, i_8_1644, i_8_1648, i_8_1650, i_8_1652, i_8_1654, i_8_1676, i_8_1679, i_8_1681, i_8_1713, i_8_1716, i_8_1717, i_8_1720, i_8_1722, i_8_1723, i_8_1741, i_8_1750, i_8_1751, i_8_1758, i_8_1812, i_8_1828, i_8_1881, i_8_1882, i_8_1884, i_8_2088, i_8_2133, i_8_2136, i_8_2138, i_8_2143, i_8_2242, i_8_2249, i_8_2272, i_8_2288, o_8_184);
	kernel_8_185 k_8_185(i_8_19, i_8_43, i_8_44, i_8_99, i_8_136, i_8_138, i_8_187, i_8_225, i_8_262, i_8_334, i_8_336, i_8_365, i_8_369, i_8_370, i_8_379, i_8_423, i_8_427, i_8_439, i_8_492, i_8_497, i_8_505, i_8_554, i_8_568, i_8_588, i_8_594, i_8_597, i_8_604, i_8_630, i_8_639, i_8_652, i_8_661, i_8_675, i_8_678, i_8_695, i_8_705, i_8_833, i_8_837, i_8_846, i_8_850, i_8_855, i_8_882, i_8_883, i_8_937, i_8_966, i_8_1062, i_8_1071, i_8_1107, i_8_1110, i_8_1117, i_8_1135, i_8_1153, i_8_1191, i_8_1215, i_8_1226, i_8_1243, i_8_1269, i_8_1297, i_8_1351, i_8_1354, i_8_1355, i_8_1431, i_8_1434, i_8_1474, i_8_1486, i_8_1503, i_8_1602, i_8_1611, i_8_1629, i_8_1671, i_8_1681, i_8_1682, i_8_1696, i_8_1710, i_8_1711, i_8_1746, i_8_1755, i_8_1756, i_8_1767, i_8_1809, i_8_1812, i_8_1824, i_8_1836, i_8_1840, i_8_1867, i_8_1881, i_8_1882, i_8_1891, i_8_1945, i_8_1962, i_8_1963, i_8_1980, i_8_2038, i_8_2106, i_8_2107, i_8_2125, i_8_2149, i_8_2152, i_8_2156, i_8_2169, i_8_2242, o_8_185);
	kernel_8_186 k_8_186(i_8_22, i_8_34, i_8_98, i_8_107, i_8_114, i_8_130, i_8_131, i_8_165, i_8_166, i_8_256, i_8_320, i_8_322, i_8_345, i_8_375, i_8_390, i_8_397, i_8_398, i_8_439, i_8_450, i_8_451, i_8_457, i_8_492, i_8_508, i_8_530, i_8_580, i_8_606, i_8_608, i_8_626, i_8_639, i_8_643, i_8_660, i_8_665, i_8_675, i_8_707, i_8_748, i_8_750, i_8_778, i_8_811, i_8_838, i_8_853, i_8_883, i_8_888, i_8_921, i_8_955, i_8_1099, i_8_1102, i_8_1108, i_8_1134, i_8_1135, i_8_1231, i_8_1233, i_8_1236, i_8_1263, i_8_1273, i_8_1286, i_8_1300, i_8_1352, i_8_1360, i_8_1362, i_8_1384, i_8_1423, i_8_1441, i_8_1442, i_8_1461, i_8_1462, i_8_1471, i_8_1512, i_8_1559, i_8_1569, i_8_1570, i_8_1603, i_8_1615, i_8_1616, i_8_1618, i_8_1642, i_8_1643, i_8_1644, i_8_1719, i_8_1781, i_8_1783, i_8_1787, i_8_1822, i_8_1836, i_8_1849, i_8_1852, i_8_1935, i_8_1954, i_8_1958, i_8_1981, i_8_1993, i_8_2055, i_8_2077, i_8_2088, i_8_2120, i_8_2151, i_8_2163, i_8_2169, i_8_2170, i_8_2212, i_8_2296, o_8_186);
	kernel_8_187 k_8_187(i_8_23, i_8_52, i_8_81, i_8_93, i_8_111, i_8_114, i_8_115, i_8_117, i_8_118, i_8_162, i_8_165, i_8_166, i_8_173, i_8_279, i_8_318, i_8_346, i_8_349, i_8_382, i_8_392, i_8_433, i_8_486, i_8_493, i_8_556, i_8_562, i_8_621, i_8_628, i_8_630, i_8_666, i_8_696, i_8_697, i_8_712, i_8_715, i_8_716, i_8_718, i_8_720, i_8_762, i_8_819, i_8_826, i_8_845, i_8_846, i_8_928, i_8_956, i_8_985, i_8_996, i_8_1026, i_8_1057, i_8_1059, i_8_1060, i_8_1061, i_8_1065, i_8_1080, i_8_1114, i_8_1158, i_8_1164, i_8_1183, i_8_1226, i_8_1229, i_8_1258, i_8_1315, i_8_1353, i_8_1359, i_8_1467, i_8_1471, i_8_1565, i_8_1587, i_8_1608, i_8_1621, i_8_1642, i_8_1696, i_8_1699, i_8_1703, i_8_1704, i_8_1705, i_8_1728, i_8_1734, i_8_1752, i_8_1773, i_8_1800, i_8_1857, i_8_1860, i_8_1867, i_8_1885, i_8_1962, i_8_1967, i_8_1983, i_8_1984, i_8_1986, i_8_2017, i_8_2061, i_8_2115, i_8_2125, i_8_2142, i_8_2143, i_8_2145, i_8_2187, i_8_2192, i_8_2224, i_8_2225, i_8_2282, i_8_2292, o_8_187);
	kernel_8_188 k_8_188(i_8_33, i_8_53, i_8_55, i_8_57, i_8_63, i_8_86, i_8_97, i_8_98, i_8_141, i_8_223, i_8_256, i_8_260, i_8_313, i_8_314, i_8_328, i_8_346, i_8_362, i_8_363, i_8_373, i_8_379, i_8_439, i_8_481, i_8_507, i_8_525, i_8_528, i_8_529, i_8_530, i_8_553, i_8_556, i_8_557, i_8_598, i_8_602, i_8_633, i_8_657, i_8_658, i_8_691, i_8_692, i_8_703, i_8_705, i_8_789, i_8_800, i_8_853, i_8_854, i_8_855, i_8_880, i_8_946, i_8_1050, i_8_1072, i_8_1113, i_8_1120, i_8_1123, i_8_1124, i_8_1191, i_8_1223, i_8_1232, i_8_1263, i_8_1264, i_8_1274, i_8_1299, i_8_1305, i_8_1307, i_8_1309, i_8_1317, i_8_1318, i_8_1327, i_8_1331, i_8_1407, i_8_1450, i_8_1467, i_8_1470, i_8_1540, i_8_1545, i_8_1564, i_8_1573, i_8_1574, i_8_1576, i_8_1637, i_8_1675, i_8_1677, i_8_1678, i_8_1680, i_8_1741, i_8_1749, i_8_1790, i_8_1795, i_8_1808, i_8_1879, i_8_1884, i_8_1907, i_8_1995, i_8_1997, i_8_2031, i_8_2032, i_8_2095, i_8_2096, i_8_2104, i_8_2105, i_8_2222, i_8_2260, i_8_2275, o_8_188);
	kernel_8_189 k_8_189(i_8_61, i_8_80, i_8_87, i_8_88, i_8_160, i_8_165, i_8_174, i_8_177, i_8_196, i_8_256, i_8_268, i_8_309, i_8_312, i_8_313, i_8_331, i_8_356, i_8_376, i_8_395, i_8_418, i_8_517, i_8_520, i_8_522, i_8_529, i_8_530, i_8_535, i_8_550, i_8_652, i_8_696, i_8_701, i_8_704, i_8_709, i_8_718, i_8_751, i_8_832, i_8_835, i_8_841, i_8_853, i_8_862, i_8_873, i_8_916, i_8_933, i_8_940, i_8_1014, i_8_1043, i_8_1067, i_8_1111, i_8_1131, i_8_1158, i_8_1177, i_8_1204, i_8_1264, i_8_1273, i_8_1299, i_8_1300, i_8_1309, i_8_1317, i_8_1321, i_8_1348, i_8_1353, i_8_1366, i_8_1375, i_8_1381, i_8_1434, i_8_1446, i_8_1454, i_8_1498, i_8_1537, i_8_1553, i_8_1560, i_8_1618, i_8_1619, i_8_1668, i_8_1690, i_8_1707, i_8_1709, i_8_1768, i_8_1771, i_8_1818, i_8_1822, i_8_1824, i_8_1826, i_8_1840, i_8_1864, i_8_1870, i_8_1871, i_8_1995, i_8_2058, i_8_2112, i_8_2137, i_8_2139, i_8_2141, i_8_2147, i_8_2148, i_8_2151, i_8_2174, i_8_2185, i_8_2229, i_8_2240, i_8_2258, i_8_2274, o_8_189);
	kernel_8_190 k_8_190(i_8_71, i_8_142, i_8_143, i_8_154, i_8_173, i_8_202, i_8_203, i_8_205, i_8_208, i_8_268, i_8_275, i_8_278, i_8_341, i_8_345, i_8_346, i_8_348, i_8_377, i_8_380, i_8_495, i_8_496, i_8_497, i_8_522, i_8_523, i_8_524, i_8_553, i_8_555, i_8_607, i_8_609, i_8_620, i_8_652, i_8_696, i_8_700, i_8_837, i_8_838, i_8_839, i_8_841, i_8_868, i_8_879, i_8_881, i_8_980, i_8_1033, i_8_1049, i_8_1057, i_8_1088, i_8_1110, i_8_1128, i_8_1204, i_8_1281, i_8_1284, i_8_1285, i_8_1286, i_8_1302, i_8_1303, i_8_1322, i_8_1343, i_8_1396, i_8_1402, i_8_1430, i_8_1436, i_8_1528, i_8_1620, i_8_1708, i_8_1714, i_8_1727, i_8_1747, i_8_1762, i_8_1766, i_8_1778, i_8_1795, i_8_1798, i_8_1799, i_8_1800, i_8_1802, i_8_1803, i_8_1804, i_8_1805, i_8_1808, i_8_1826, i_8_1858, i_8_1861, i_8_1864, i_8_1865, i_8_1914, i_8_1915, i_8_1964, i_8_1970, i_8_1980, i_8_1983, i_8_2046, i_8_2047, i_8_2049, i_8_2065, i_8_2073, i_8_2125, i_8_2128, i_8_2237, i_8_2244, i_8_2286, i_8_2287, i_8_2289, o_8_190);
	kernel_8_191 k_8_191(i_8_22, i_8_25, i_8_52, i_8_54, i_8_60, i_8_138, i_8_160, i_8_193, i_8_262, i_8_336, i_8_341, i_8_354, i_8_376, i_8_385, i_8_403, i_8_457, i_8_499, i_8_529, i_8_555, i_8_573, i_8_604, i_8_607, i_8_609, i_8_653, i_8_675, i_8_678, i_8_688, i_8_798, i_8_799, i_8_837, i_8_838, i_8_843, i_8_849, i_8_881, i_8_922, i_8_924, i_8_933, i_8_968, i_8_970, i_8_991, i_8_993, i_8_995, i_8_1024, i_8_1043, i_8_1072, i_8_1075, i_8_1101, i_8_1112, i_8_1140, i_8_1155, i_8_1173, i_8_1194, i_8_1229, i_8_1263, i_8_1267, i_8_1284, i_8_1300, i_8_1301, i_8_1328, i_8_1331, i_8_1372, i_8_1384, i_8_1430, i_8_1442, i_8_1470, i_8_1473, i_8_1488, i_8_1527, i_8_1569, i_8_1570, i_8_1579, i_8_1609, i_8_1610, i_8_1624, i_8_1625, i_8_1629, i_8_1632, i_8_1644, i_8_1649, i_8_1700, i_8_1766, i_8_1788, i_8_1797, i_8_1818, i_8_1824, i_8_1828, i_8_1839, i_8_1893, i_8_1894, i_8_1942, i_8_1996, i_8_2019, i_8_2028, i_8_2112, i_8_2113, i_8_2152, i_8_2167, i_8_2231, i_8_2235, i_8_2241, o_8_191);
	kernel_8_192 k_8_192(i_8_33, i_8_88, i_8_114, i_8_266, i_8_293, i_8_374, i_8_377, i_8_383, i_8_386, i_8_440, i_8_463, i_8_476, i_8_482, i_8_485, i_8_500, i_8_524, i_8_530, i_8_571, i_8_574, i_8_616, i_8_617, i_8_624, i_8_634, i_8_674, i_8_760, i_8_762, i_8_781, i_8_787, i_8_826, i_8_841, i_8_878, i_8_886, i_8_895, i_8_936, i_8_939, i_8_945, i_8_946, i_8_995, i_8_1011, i_8_1013, i_8_1030, i_8_1114, i_8_1124, i_8_1140, i_8_1159, i_8_1192, i_8_1222, i_8_1237, i_8_1259, i_8_1264, i_8_1282, i_8_1283, i_8_1284, i_8_1285, i_8_1305, i_8_1306, i_8_1328, i_8_1331, i_8_1346, i_8_1438, i_8_1439, i_8_1441, i_8_1453, i_8_1470, i_8_1509, i_8_1534, i_8_1535, i_8_1544, i_8_1565, i_8_1632, i_8_1655, i_8_1681, i_8_1706, i_8_1732, i_8_1733, i_8_1742, i_8_1787, i_8_1841, i_8_1857, i_8_1859, i_8_1866, i_8_1867, i_8_1884, i_8_1885, i_8_1918, i_8_1919, i_8_1949, i_8_1952, i_8_1966, i_8_1967, i_8_2056, i_8_2111, i_8_2127, i_8_2128, i_8_2143, i_8_2156, i_8_2191, i_8_2192, i_8_2214, i_8_2276, o_8_192);
	kernel_8_193 k_8_193(i_8_33, i_8_39, i_8_45, i_8_55, i_8_104, i_8_114, i_8_119, i_8_190, i_8_226, i_8_327, i_8_364, i_8_367, i_8_423, i_8_426, i_8_450, i_8_481, i_8_525, i_8_526, i_8_530, i_8_549, i_8_570, i_8_588, i_8_612, i_8_659, i_8_661, i_8_665, i_8_684, i_8_695, i_8_697, i_8_700, i_8_706, i_8_747, i_8_769, i_8_777, i_8_792, i_8_832, i_8_877, i_8_882, i_8_981, i_8_990, i_8_996, i_8_1032, i_8_1044, i_8_1128, i_8_1135, i_8_1138, i_8_1143, i_8_1144, i_8_1148, i_8_1152, i_8_1188, i_8_1270, i_8_1278, i_8_1330, i_8_1360, i_8_1362, i_8_1368, i_8_1393, i_8_1404, i_8_1408, i_8_1413, i_8_1442, i_8_1480, i_8_1506, i_8_1530, i_8_1543, i_8_1620, i_8_1630, i_8_1632, i_8_1639, i_8_1648, i_8_1650, i_8_1668, i_8_1674, i_8_1701, i_8_1714, i_8_1719, i_8_1728, i_8_1764, i_8_1777, i_8_1821, i_8_1881, i_8_1900, i_8_1903, i_8_1935, i_8_1967, i_8_1971, i_8_1983, i_8_1984, i_8_2070, i_8_2108, i_8_2133, i_8_2146, i_8_2149, i_8_2150, i_8_2152, i_8_2227, i_8_2242, i_8_2244, i_8_2269, o_8_193);
	kernel_8_194 k_8_194(i_8_21, i_8_42, i_8_52, i_8_55, i_8_58, i_8_89, i_8_120, i_8_129, i_8_183, i_8_184, i_8_211, i_8_218, i_8_241, i_8_262, i_8_319, i_8_365, i_8_369, i_8_427, i_8_456, i_8_478, i_8_535, i_8_543, i_8_549, i_8_551, i_8_593, i_8_611, i_8_612, i_8_613, i_8_634, i_8_643, i_8_656, i_8_662, i_8_665, i_8_730, i_8_787, i_8_802, i_8_804, i_8_832, i_8_851, i_8_865, i_8_876, i_8_891, i_8_895, i_8_931, i_8_945, i_8_994, i_8_1101, i_8_1104, i_8_1115, i_8_1129, i_8_1240, i_8_1251, i_8_1256, i_8_1267, i_8_1268, i_8_1271, i_8_1291, i_8_1296, i_8_1329, i_8_1366, i_8_1378, i_8_1407, i_8_1435, i_8_1461, i_8_1465, i_8_1482, i_8_1544, i_8_1608, i_8_1620, i_8_1627, i_8_1651, i_8_1740, i_8_1747, i_8_1750, i_8_1760, i_8_1784, i_8_1787, i_8_1788, i_8_1789, i_8_1810, i_8_1840, i_8_1867, i_8_1899, i_8_1963, i_8_1966, i_8_1983, i_8_1984, i_8_1992, i_8_2068, i_8_2091, i_8_2104, i_8_2127, i_8_2158, i_8_2191, i_8_2216, i_8_2236, i_8_2240, i_8_2241, i_8_2246, i_8_2248, o_8_194);
	kernel_8_195 k_8_195(i_8_21, i_8_79, i_8_129, i_8_138, i_8_192, i_8_195, i_8_228, i_8_256, i_8_345, i_8_347, i_8_349, i_8_354, i_8_362, i_8_368, i_8_382, i_8_428, i_8_477, i_8_525, i_8_529, i_8_552, i_8_555, i_8_567, i_8_570, i_8_651, i_8_654, i_8_662, i_8_675, i_8_688, i_8_696, i_8_703, i_8_705, i_8_729, i_8_732, i_8_750, i_8_751, i_8_774, i_8_775, i_8_789, i_8_801, i_8_832, i_8_859, i_8_885, i_8_886, i_8_969, i_8_984, i_8_1002, i_8_1038, i_8_1051, i_8_1101, i_8_1119, i_8_1130, i_8_1137, i_8_1146, i_8_1164, i_8_1191, i_8_1356, i_8_1371, i_8_1395, i_8_1405, i_8_1435, i_8_1507, i_8_1524, i_8_1546, i_8_1547, i_8_1597, i_8_1606, i_8_1610, i_8_1626, i_8_1632, i_8_1650, i_8_1659, i_8_1677, i_8_1683, i_8_1722, i_8_1728, i_8_1731, i_8_1767, i_8_1768, i_8_1779, i_8_1780, i_8_1825, i_8_1858, i_8_1888, i_8_1938, i_8_1947, i_8_1978, i_8_1992, i_8_2056, i_8_2073, i_8_2091, i_8_2092, i_8_2097, i_8_2100, i_8_2142, i_8_2146, i_8_2172, i_8_2215, i_8_2258, i_8_2284, i_8_2298, o_8_195);
	kernel_8_196 k_8_196(i_8_0, i_8_3, i_8_67, i_8_73, i_8_75, i_8_84, i_8_111, i_8_114, i_8_126, i_8_184, i_8_192, i_8_194, i_8_246, i_8_274, i_8_301, i_8_305, i_8_345, i_8_354, i_8_364, i_8_388, i_8_397, i_8_418, i_8_453, i_8_462, i_8_463, i_8_495, i_8_572, i_8_578, i_8_588, i_8_592, i_8_604, i_8_615, i_8_641, i_8_642, i_8_648, i_8_652, i_8_659, i_8_669, i_8_676, i_8_699, i_8_733, i_8_748, i_8_756, i_8_833, i_8_841, i_8_866, i_8_886, i_8_913, i_8_1107, i_8_1201, i_8_1219, i_8_1225, i_8_1226, i_8_1234, i_8_1240, i_8_1279, i_8_1315, i_8_1335, i_8_1336, i_8_1353, i_8_1355, i_8_1363, i_8_1366, i_8_1375, i_8_1389, i_8_1390, i_8_1436, i_8_1492, i_8_1494, i_8_1508, i_8_1509, i_8_1533, i_8_1606, i_8_1633, i_8_1638, i_8_1641, i_8_1682, i_8_1697, i_8_1703, i_8_1747, i_8_1765, i_8_1787, i_8_1819, i_8_1820, i_8_1843, i_8_1848, i_8_1863, i_8_1866, i_8_1881, i_8_1884, i_8_1918, i_8_1927, i_8_2064, i_8_2133, i_8_2224, i_8_2232, i_8_2242, i_8_2245, i_8_2246, i_8_2281, o_8_196);
	kernel_8_197 k_8_197(i_8_66, i_8_75, i_8_88, i_8_114, i_8_148, i_8_165, i_8_174, i_8_193, i_8_202, i_8_228, i_8_300, i_8_312, i_8_336, i_8_349, i_8_354, i_8_366, i_8_418, i_8_426, i_8_429, i_8_453, i_8_489, i_8_508, i_8_522, i_8_535, i_8_574, i_8_582, i_8_606, i_8_608, i_8_615, i_8_657, i_8_665, i_8_700, i_8_701, i_8_705, i_8_730, i_8_759, i_8_772, i_8_835, i_8_840, i_8_841, i_8_858, i_8_865, i_8_870, i_8_912, i_8_921, i_8_969, i_8_1029, i_8_1034, i_8_1038, i_8_1068, i_8_1114, i_8_1123, i_8_1132, i_8_1134, i_8_1227, i_8_1232, i_8_1281, i_8_1305, i_8_1323, i_8_1372, i_8_1398, i_8_1470, i_8_1548, i_8_1571, i_8_1587, i_8_1623, i_8_1633, i_8_1686, i_8_1696, i_8_1699, i_8_1767, i_8_1773, i_8_1790, i_8_1794, i_8_1806, i_8_1822, i_8_1824, i_8_1840, i_8_1869, i_8_1929, i_8_1938, i_8_2004, i_8_2008, i_8_2010, i_8_2019, i_8_2073, i_8_2103, i_8_2109, i_8_2134, i_8_2144, i_8_2145, i_8_2147, i_8_2154, i_8_2158, i_8_2225, i_8_2226, i_8_2227, i_8_2229, i_8_2271, i_8_2281, o_8_197);
	kernel_8_198 k_8_198(i_8_58, i_8_73, i_8_76, i_8_77, i_8_115, i_8_116, i_8_137, i_8_140, i_8_181, i_8_184, i_8_221, i_8_231, i_8_256, i_8_301, i_8_320, i_8_389, i_8_419, i_8_431, i_8_482, i_8_496, i_8_509, i_8_524, i_8_526, i_8_527, i_8_572, i_8_590, i_8_608, i_8_611, i_8_655, i_8_658, i_8_694, i_8_696, i_8_737, i_8_760, i_8_761, i_8_776, i_8_824, i_8_837, i_8_838, i_8_850, i_8_928, i_8_1010, i_8_1100, i_8_1103, i_8_1129, i_8_1130, i_8_1229, i_8_1247, i_8_1268, i_8_1279, i_8_1295, i_8_1316, i_8_1319, i_8_1327, i_8_1334, i_8_1397, i_8_1423, i_8_1424, i_8_1442, i_8_1462, i_8_1463, i_8_1472, i_8_1478, i_8_1481, i_8_1493, i_8_1511, i_8_1514, i_8_1525, i_8_1526, i_8_1549, i_8_1550, i_8_1551, i_8_1559, i_8_1640, i_8_1643, i_8_1675, i_8_1676, i_8_1679, i_8_1684, i_8_1697, i_8_1700, i_8_1706, i_8_1721, i_8_1747, i_8_1780, i_8_1781, i_8_1787, i_8_1793, i_8_1810, i_8_1838, i_8_1840, i_8_1841, i_8_1885, i_8_1937, i_8_1949, i_8_1954, i_8_1968, i_8_2075, i_8_2135, i_8_2297, o_8_198);
	kernel_8_199 k_8_199(i_8_1, i_8_49, i_8_76, i_8_86, i_8_118, i_8_119, i_8_164, i_8_167, i_8_226, i_8_244, i_8_300, i_8_326, i_8_350, i_8_425, i_8_452, i_8_464, i_8_487, i_8_490, i_8_496, i_8_497, i_8_500, i_8_530, i_8_556, i_8_589, i_8_605, i_8_653, i_8_695, i_8_698, i_8_707, i_8_823, i_8_824, i_8_838, i_8_839, i_8_841, i_8_875, i_8_884, i_8_929, i_8_968, i_8_992, i_8_1001, i_8_1036, i_8_1037, i_8_1046, i_8_1052, i_8_1072, i_8_1075, i_8_1076, i_8_1163, i_8_1166, i_8_1226, i_8_1233, i_8_1270, i_8_1274, i_8_1280, i_8_1281, i_8_1282, i_8_1298, i_8_1318, i_8_1321, i_8_1327, i_8_1408, i_8_1432, i_8_1435, i_8_1436, i_8_1467, i_8_1468, i_8_1478, i_8_1496, i_8_1534, i_8_1543, i_8_1544, i_8_1657, i_8_1703, i_8_1733, i_8_1749, i_8_1751, i_8_1754, i_8_1760, i_8_1766, i_8_1769, i_8_1777, i_8_1811, i_8_1822, i_8_1850, i_8_1868, i_8_1974, i_8_1976, i_8_1982, i_8_1993, i_8_1994, i_8_2057, i_8_2102, i_8_2125, i_8_2135, i_8_2143, i_8_2153, i_8_2223, i_8_2225, i_8_2269, i_8_2273, o_8_199);
	kernel_8_200 k_8_200(i_8_25, i_8_50, i_8_53, i_8_111, i_8_114, i_8_115, i_8_116, i_8_123, i_8_124, i_8_175, i_8_179, i_8_219, i_8_220, i_8_221, i_8_224, i_8_257, i_8_383, i_8_453, i_8_455, i_8_457, i_8_458, i_8_523, i_8_571, i_8_572, i_8_575, i_8_601, i_8_602, i_8_607, i_8_657, i_8_658, i_8_689, i_8_702, i_8_703, i_8_704, i_8_768, i_8_775, i_8_776, i_8_798, i_8_883, i_8_887, i_8_888, i_8_932, i_8_959, i_8_961, i_8_966, i_8_1072, i_8_1167, i_8_1178, i_8_1179, i_8_1180, i_8_1227, i_8_1228, i_8_1229, i_8_1262, i_8_1263, i_8_1278, i_8_1296, i_8_1470, i_8_1474, i_8_1487, i_8_1490, i_8_1560, i_8_1563, i_8_1564, i_8_1584, i_8_1585, i_8_1587, i_8_1588, i_8_1623, i_8_1632, i_8_1683, i_8_1695, i_8_1696, i_8_1699, i_8_1700, i_8_1738, i_8_1746, i_8_1758, i_8_1770, i_8_1772, i_8_1787, i_8_1789, i_8_1818, i_8_1820, i_8_1821, i_8_1854, i_8_1857, i_8_1969, i_8_2009, i_8_2073, i_8_2129, i_8_2222, i_8_2224, i_8_2226, i_8_2237, i_8_2247, i_8_2248, i_8_2249, i_8_2261, i_8_2293, o_8_200);
	kernel_8_201 k_8_201(i_8_21, i_8_25, i_8_33, i_8_34, i_8_85, i_8_183, i_8_190, i_8_294, i_8_300, i_8_373, i_8_386, i_8_420, i_8_481, i_8_483, i_8_508, i_8_510, i_8_529, i_8_530, i_8_589, i_8_592, i_8_594, i_8_595, i_8_598, i_8_601, i_8_607, i_8_634, i_8_636, i_8_691, i_8_714, i_8_715, i_8_717, i_8_759, i_8_777, i_8_778, i_8_789, i_8_790, i_8_800, i_8_810, i_8_838, i_8_852, i_8_853, i_8_912, i_8_933, i_8_997, i_8_1005, i_8_1059, i_8_1093, i_8_1114, i_8_1123, i_8_1129, i_8_1159, i_8_1222, i_8_1277, i_8_1282, i_8_1285, i_8_1286, i_8_1307, i_8_1320, i_8_1321, i_8_1330, i_8_1366, i_8_1431, i_8_1451, i_8_1470, i_8_1471, i_8_1473, i_8_1474, i_8_1537, i_8_1543, i_8_1545, i_8_1548, i_8_1563, i_8_1570, i_8_1590, i_8_1668, i_8_1671, i_8_1681, i_8_1682, i_8_1723, i_8_1743, i_8_1749, i_8_1750, i_8_1753, i_8_1875, i_8_1876, i_8_1878, i_8_1920, i_8_1959, i_8_1960, i_8_1965, i_8_1969, i_8_1971, i_8_1995, i_8_2011, i_8_2137, i_8_2235, i_8_2253, i_8_2277, i_8_2284, i_8_2292, o_8_201);
	kernel_8_202 k_8_202(i_8_1, i_8_19, i_8_73, i_8_76, i_8_82, i_8_188, i_8_202, i_8_244, i_8_268, i_8_274, i_8_275, i_8_325, i_8_335, i_8_343, i_8_352, i_8_353, i_8_373, i_8_426, i_8_459, i_8_478, i_8_500, i_8_513, i_8_514, i_8_515, i_8_523, i_8_613, i_8_631, i_8_662, i_8_663, i_8_729, i_8_731, i_8_751, i_8_756, i_8_811, i_8_812, i_8_819, i_8_864, i_8_910, i_8_950, i_8_973, i_8_1029, i_8_1057, i_8_1072, i_8_1108, i_8_1170, i_8_1187, i_8_1188, i_8_1225, i_8_1226, i_8_1238, i_8_1261, i_8_1330, i_8_1355, i_8_1408, i_8_1429, i_8_1454, i_8_1468, i_8_1471, i_8_1494, i_8_1495, i_8_1496, i_8_1507, i_8_1509, i_8_1542, i_8_1561, i_8_1624, i_8_1641, i_8_1649, i_8_1656, i_8_1694, i_8_1702, i_8_1751, i_8_1800, i_8_1804, i_8_1810, i_8_1855, i_8_1864, i_8_1865, i_8_1873, i_8_1874, i_8_1963, i_8_1968, i_8_1973, i_8_1992, i_8_1994, i_8_2008, i_8_2045, i_8_2056, i_8_2062, i_8_2063, i_8_2071, i_8_2116, i_8_2117, i_8_2118, i_8_2130, i_8_2143, i_8_2170, i_8_2228, i_8_2234, i_8_2253, o_8_202);
	kernel_8_203 k_8_203(i_8_25, i_8_27, i_8_46, i_8_54, i_8_57, i_8_70, i_8_104, i_8_171, i_8_172, i_8_197, i_8_337, i_8_372, i_8_415, i_8_423, i_8_427, i_8_450, i_8_453, i_8_549, i_8_571, i_8_586, i_8_594, i_8_598, i_8_599, i_8_604, i_8_632, i_8_633, i_8_640, i_8_658, i_8_662, i_8_679, i_8_695, i_8_704, i_8_778, i_8_781, i_8_835, i_8_837, i_8_865, i_8_880, i_8_993, i_8_1035, i_8_1063, i_8_1137, i_8_1154, i_8_1178, i_8_1264, i_8_1281, i_8_1297, i_8_1298, i_8_1299, i_8_1367, i_8_1406, i_8_1470, i_8_1471, i_8_1557, i_8_1558, i_8_1559, i_8_1571, i_8_1602, i_8_1603, i_8_1611, i_8_1612, i_8_1629, i_8_1635, i_8_1646, i_8_1655, i_8_1686, i_8_1690, i_8_1710, i_8_1711, i_8_1713, i_8_1750, i_8_1753, i_8_1754, i_8_1755, i_8_1758, i_8_1759, i_8_1774, i_8_1780, i_8_1809, i_8_1819, i_8_1824, i_8_1889, i_8_1971, i_8_1980, i_8_1989, i_8_1993, i_8_1994, i_8_1996, i_8_2052, i_8_2053, i_8_2069, i_8_2106, i_8_2116, i_8_2147, i_8_2149, i_8_2223, i_8_2233, i_8_2235, i_8_2244, i_8_2259, o_8_203);
	kernel_8_204 k_8_204(i_8_32, i_8_73, i_8_82, i_8_88, i_8_90, i_8_104, i_8_182, i_8_216, i_8_217, i_8_220, i_8_244, i_8_300, i_8_319, i_8_349, i_8_364, i_8_369, i_8_380, i_8_385, i_8_388, i_8_460, i_8_471, i_8_496, i_8_515, i_8_528, i_8_552, i_8_555, i_8_623, i_8_657, i_8_659, i_8_664, i_8_665, i_8_693, i_8_711, i_8_737, i_8_778, i_8_779, i_8_783, i_8_793, i_8_830, i_8_844, i_8_874, i_8_967, i_8_970, i_8_998, i_8_1042, i_8_1071, i_8_1079, i_8_1104, i_8_1105, i_8_1110, i_8_1111, i_8_1151, i_8_1224, i_8_1225, i_8_1246, i_8_1260, i_8_1279, i_8_1281, i_8_1283, i_8_1306, i_8_1359, i_8_1397, i_8_1477, i_8_1486, i_8_1487, i_8_1522, i_8_1537, i_8_1538, i_8_1541, i_8_1549, i_8_1567, i_8_1594, i_8_1602, i_8_1649, i_8_1670, i_8_1680, i_8_1719, i_8_1720, i_8_1746, i_8_1752, i_8_1800, i_8_1803, i_8_1815, i_8_1816, i_8_1891, i_8_1910, i_8_1948, i_8_1962, i_8_1963, i_8_1969, i_8_1972, i_8_1989, i_8_2047, i_8_2071, i_8_2106, i_8_2107, i_8_2113, i_8_2133, i_8_2140, i_8_2141, o_8_204);
	kernel_8_205 k_8_205(i_8_34, i_8_85, i_8_158, i_8_181, i_8_184, i_8_203, i_8_217, i_8_220, i_8_233, i_8_237, i_8_238, i_8_255, i_8_304, i_8_371, i_8_374, i_8_380, i_8_382, i_8_385, i_8_423, i_8_437, i_8_453, i_8_477, i_8_478, i_8_481, i_8_482, i_8_484, i_8_485, i_8_498, i_8_499, i_8_505, i_8_523, i_8_526, i_8_532, i_8_564, i_8_634, i_8_661, i_8_684, i_8_703, i_8_757, i_8_759, i_8_760, i_8_761, i_8_767, i_8_780, i_8_811, i_8_823, i_8_830, i_8_869, i_8_892, i_8_904, i_8_1013, i_8_1030, i_8_1111, i_8_1112, i_8_1135, i_8_1174, i_8_1282, i_8_1294, i_8_1309, i_8_1328, i_8_1363, i_8_1366, i_8_1398, i_8_1506, i_8_1522, i_8_1537, i_8_1552, i_8_1565, i_8_1577, i_8_1605, i_8_1676, i_8_1678, i_8_1711, i_8_1723, i_8_1729, i_8_1730, i_8_1749, i_8_1752, i_8_1760, i_8_1805, i_8_1807, i_8_1818, i_8_1855, i_8_1903, i_8_1920, i_8_1947, i_8_1980, i_8_2020, i_8_2037, i_8_2038, i_8_2070, i_8_2093, i_8_2109, i_8_2150, i_8_2170, i_8_2218, i_8_2224, i_8_2237, i_8_2271, i_8_2286, o_8_205);
	kernel_8_206 k_8_206(i_8_22, i_8_41, i_8_52, i_8_53, i_8_76, i_8_103, i_8_130, i_8_138, i_8_168, i_8_169, i_8_319, i_8_354, i_8_365, i_8_373, i_8_382, i_8_386, i_8_394, i_8_429, i_8_430, i_8_454, i_8_492, i_8_493, i_8_495, i_8_507, i_8_538, i_8_544, i_8_556, i_8_565, i_8_610, i_8_637, i_8_679, i_8_694, i_8_724, i_8_747, i_8_766, i_8_823, i_8_835, i_8_847, i_8_962, i_8_970, i_8_1052, i_8_1065, i_8_1114, i_8_1115, i_8_1254, i_8_1257, i_8_1264, i_8_1265, i_8_1283, i_8_1315, i_8_1318, i_8_1354, i_8_1362, i_8_1363, i_8_1381, i_8_1384, i_8_1410, i_8_1413, i_8_1440, i_8_1455, i_8_1465, i_8_1467, i_8_1539, i_8_1542, i_8_1545, i_8_1553, i_8_1583, i_8_1669, i_8_1672, i_8_1687, i_8_1699, i_8_1731, i_8_1750, i_8_1801, i_8_1819, i_8_1823, i_8_1826, i_8_1850, i_8_1855, i_8_1859, i_8_1883, i_8_1972, i_8_1980, i_8_1986, i_8_2023, i_8_2073, i_8_2083, i_8_2126, i_8_2138, i_8_2146, i_8_2147, i_8_2191, i_8_2193, i_8_2224, i_8_2227, i_8_2243, i_8_2262, i_8_2278, i_8_2289, i_8_2292, o_8_206);
	kernel_8_207 k_8_207(i_8_18, i_8_37, i_8_39, i_8_49, i_8_63, i_8_81, i_8_102, i_8_147, i_8_175, i_8_189, i_8_198, i_8_220, i_8_252, i_8_261, i_8_270, i_8_297, i_8_302, i_8_306, i_8_363, i_8_426, i_8_489, i_8_531, i_8_534, i_8_539, i_8_552, i_8_568, i_8_634, i_8_639, i_8_648, i_8_651, i_8_666, i_8_674, i_8_679, i_8_697, i_8_712, i_8_748, i_8_823, i_8_841, i_8_844, i_8_862, i_8_865, i_8_891, i_8_963, i_8_966, i_8_1080, i_8_1098, i_8_1128, i_8_1133, i_8_1170, i_8_1171, i_8_1179, i_8_1224, i_8_1227, i_8_1233, i_8_1236, i_8_1237, i_8_1263, i_8_1281, i_8_1297, i_8_1326, i_8_1377, i_8_1381, i_8_1386, i_8_1395, i_8_1431, i_8_1458, i_8_1506, i_8_1534, i_8_1560, i_8_1630, i_8_1639, i_8_1647, i_8_1650, i_8_1651, i_8_1674, i_8_1696, i_8_1754, i_8_1764, i_8_1767, i_8_1803, i_8_1804, i_8_1818, i_8_1864, i_8_1866, i_8_1910, i_8_1918, i_8_1927, i_8_1947, i_8_1966, i_8_1988, i_8_2034, i_8_2043, i_8_2062, i_8_2142, i_8_2146, i_8_2169, i_8_2177, i_8_2232, i_8_2268, i_8_2289, o_8_207);
	kernel_8_208 k_8_208(i_8_7, i_8_26, i_8_88, i_8_179, i_8_219, i_8_232, i_8_240, i_8_250, i_8_266, i_8_287, i_8_292, i_8_332, i_8_348, i_8_349, i_8_386, i_8_463, i_8_466, i_8_467, i_8_502, i_8_520, i_8_526, i_8_527, i_8_556, i_8_594, i_8_610, i_8_627, i_8_656, i_8_662, i_8_672, i_8_673, i_8_698, i_8_717, i_8_718, i_8_754, i_8_782, i_8_798, i_8_799, i_8_808, i_8_843, i_8_879, i_8_926, i_8_992, i_8_994, i_8_995, i_8_997, i_8_998, i_8_1060, i_8_1077, i_8_1093, i_8_1139, i_8_1194, i_8_1205, i_8_1222, i_8_1258, i_8_1285, i_8_1286, i_8_1308, i_8_1316, i_8_1342, i_8_1357, i_8_1457, i_8_1474, i_8_1509, i_8_1538, i_8_1545, i_8_1546, i_8_1553, i_8_1555, i_8_1599, i_8_1601, i_8_1610, i_8_1647, i_8_1727, i_8_1751, i_8_1770, i_8_1832, i_8_1852, i_8_1853, i_8_1870, i_8_1897, i_8_1898, i_8_1921, i_8_1922, i_8_1925, i_8_1969, i_8_2014, i_8_2032, i_8_2074, i_8_2078, i_8_2113, i_8_2122, i_8_2131, i_8_2132, i_8_2150, i_8_2183, i_8_2219, i_8_2238, i_8_2249, i_8_2275, i_8_2293, o_8_208);
	kernel_8_209 k_8_209(i_8_33, i_8_52, i_8_155, i_8_221, i_8_256, i_8_289, i_8_297, i_8_298, i_8_342, i_8_343, i_8_369, i_8_370, i_8_371, i_8_378, i_8_379, i_8_388, i_8_389, i_8_415, i_8_441, i_8_453, i_8_459, i_8_460, i_8_461, i_8_472, i_8_544, i_8_549, i_8_604, i_8_609, i_8_610, i_8_613, i_8_625, i_8_711, i_8_712, i_8_715, i_8_756, i_8_782, i_8_783, i_8_792, i_8_793, i_8_846, i_8_867, i_8_998, i_8_1008, i_8_1013, i_8_1027, i_8_1117, i_8_1118, i_8_1125, i_8_1128, i_8_1130, i_8_1156, i_8_1233, i_8_1246, i_8_1249, i_8_1324, i_8_1333, i_8_1343, i_8_1419, i_8_1420, i_8_1421, i_8_1467, i_8_1488, i_8_1531, i_8_1532, i_8_1537, i_8_1539, i_8_1540, i_8_1565, i_8_1579, i_8_1594, i_8_1595, i_8_1609, i_8_1611, i_8_1649, i_8_1676, i_8_1731, i_8_1738, i_8_1750, i_8_1783, i_8_1793, i_8_1801, i_8_1802, i_8_1864, i_8_1866, i_8_1869, i_8_1885, i_8_1926, i_8_1947, i_8_1992, i_8_2124, i_8_2125, i_8_2136, i_8_2141, i_8_2179, i_8_2180, i_8_2187, i_8_2188, i_8_2273, i_8_2287, i_8_2298, o_8_209);
	kernel_8_210 k_8_210(i_8_32, i_8_47, i_8_49, i_8_65, i_8_91, i_8_92, i_8_103, i_8_236, i_8_320, i_8_326, i_8_362, i_8_380, i_8_383, i_8_388, i_8_417, i_8_424, i_8_452, i_8_490, i_8_493, i_8_512, i_8_578, i_8_604, i_8_635, i_8_640, i_8_658, i_8_668, i_8_676, i_8_677, i_8_686, i_8_701, i_8_703, i_8_705, i_8_731, i_8_767, i_8_778, i_8_841, i_8_844, i_8_929, i_8_955, i_8_967, i_8_968, i_8_1057, i_8_1112, i_8_1226, i_8_1261, i_8_1280, i_8_1316, i_8_1334, i_8_1352, i_8_1404, i_8_1442, i_8_1456, i_8_1468, i_8_1469, i_8_1473, i_8_1514, i_8_1530, i_8_1559, i_8_1604, i_8_1607, i_8_1612, i_8_1621, i_8_1622, i_8_1631, i_8_1648, i_8_1669, i_8_1678, i_8_1680, i_8_1684, i_8_1685, i_8_1693, i_8_1724, i_8_1730, i_8_1757, i_8_1768, i_8_1778, i_8_1783, i_8_1784, i_8_1818, i_8_1825, i_8_1864, i_8_1882, i_8_1946, i_8_1981, i_8_2000, i_8_2071, i_8_2075, i_8_2107, i_8_2133, i_8_2134, i_8_2147, i_8_2154, i_8_2156, i_8_2197, i_8_2198, i_8_2206, i_8_2224, i_8_2233, i_8_2260, i_8_2273, o_8_210);
	kernel_8_211 k_8_211(i_8_13, i_8_21, i_8_28, i_8_41, i_8_55, i_8_58, i_8_72, i_8_169, i_8_172, i_8_199, i_8_221, i_8_226, i_8_253, i_8_304, i_8_415, i_8_416, i_8_419, i_8_451, i_8_489, i_8_505, i_8_506, i_8_533, i_8_549, i_8_572, i_8_595, i_8_598, i_8_602, i_8_610, i_8_624, i_8_626, i_8_630, i_8_662, i_8_675, i_8_689, i_8_693, i_8_712, i_8_730, i_8_775, i_8_841, i_8_850, i_8_866, i_8_877, i_8_980, i_8_1073, i_8_1107, i_8_1135, i_8_1143, i_8_1199, i_8_1234, i_8_1260, i_8_1270, i_8_1278, i_8_1279, i_8_1282, i_8_1286, i_8_1298, i_8_1316, i_8_1387, i_8_1407, i_8_1408, i_8_1424, i_8_1438, i_8_1452, i_8_1470, i_8_1478, i_8_1481, i_8_1558, i_8_1607, i_8_1631, i_8_1632, i_8_1659, i_8_1684, i_8_1710, i_8_1747, i_8_1748, i_8_1766, i_8_1820, i_8_1821, i_8_1823, i_8_1854, i_8_1873, i_8_1882, i_8_1883, i_8_1885, i_8_1962, i_8_1966, i_8_1980, i_8_2017, i_8_2044, i_8_2088, i_8_2125, i_8_2135, i_8_2140, i_8_2151, i_8_2169, i_8_2232, i_8_2234, i_8_2261, i_8_2273, i_8_2296, o_8_211);
	kernel_8_212 k_8_212(i_8_13, i_8_16, i_8_31, i_8_57, i_8_66, i_8_75, i_8_94, i_8_98, i_8_124, i_8_188, i_8_229, i_8_232, i_8_304, i_8_339, i_8_360, i_8_367, i_8_384, i_8_385, i_8_399, i_8_400, i_8_420, i_8_466, i_8_525, i_8_574, i_8_591, i_8_592, i_8_608, i_8_655, i_8_678, i_8_681, i_8_750, i_8_817, i_8_843, i_8_844, i_8_852, i_8_853, i_8_861, i_8_879, i_8_883, i_8_961, i_8_967, i_8_1012, i_8_1128, i_8_1140, i_8_1141, i_8_1149, i_8_1150, i_8_1158, i_8_1186, i_8_1228, i_8_1231, i_8_1236, i_8_1263, i_8_1302, i_8_1317, i_8_1320, i_8_1321, i_8_1330, i_8_1331, i_8_1482, i_8_1553, i_8_1561, i_8_1606, i_8_1608, i_8_1636, i_8_1677, i_8_1680, i_8_1716, i_8_1722, i_8_1752, i_8_1763, i_8_1789, i_8_1795, i_8_1813, i_8_1816, i_8_1818, i_8_1860, i_8_1922, i_8_1951, i_8_1960, i_8_1995, i_8_2004, i_8_2058, i_8_2076, i_8_2094, i_8_2109, i_8_2136, i_8_2137, i_8_2142, i_8_2145, i_8_2147, i_8_2158, i_8_2176, i_8_2190, i_8_2238, i_8_2239, i_8_2244, i_8_2246, i_8_2248, i_8_2266, o_8_212);
	kernel_8_213 k_8_213(i_8_9, i_8_18, i_8_37, i_8_73, i_8_102, i_8_135, i_8_183, i_8_225, i_8_226, i_8_252, i_8_255, i_8_259, i_8_279, i_8_321, i_8_364, i_8_365, i_8_370, i_8_399, i_8_495, i_8_499, i_8_534, i_8_540, i_8_567, i_8_570, i_8_594, i_8_604, i_8_639, i_8_659, i_8_660, i_8_675, i_8_678, i_8_777, i_8_783, i_8_810, i_8_841, i_8_864, i_8_868, i_8_891, i_8_937, i_8_954, i_8_966, i_8_969, i_8_975, i_8_1036, i_8_1107, i_8_1110, i_8_1111, i_8_1125, i_8_1138, i_8_1179, i_8_1197, i_8_1225, i_8_1236, i_8_1242, i_8_1246, i_8_1261, i_8_1263, i_8_1264, i_8_1314, i_8_1335, i_8_1338, i_8_1342, i_8_1344, i_8_1377, i_8_1422, i_8_1424, i_8_1434, i_8_1435, i_8_1467, i_8_1468, i_8_1476, i_8_1480, i_8_1512, i_8_1516, i_8_1524, i_8_1539, i_8_1542, i_8_1555, i_8_1557, i_8_1629, i_8_1651, i_8_1705, i_8_1753, i_8_1755, i_8_1758, i_8_1759, i_8_1767, i_8_1773, i_8_1776, i_8_1789, i_8_1790, i_8_1950, i_8_1989, i_8_1996, i_8_2133, i_8_2145, i_8_2196, i_8_2232, i_8_2233, i_8_2271, o_8_213);
	kernel_8_214 k_8_214(i_8_18, i_8_21, i_8_57, i_8_120, i_8_141, i_8_142, i_8_169, i_8_192, i_8_237, i_8_266, i_8_269, i_8_285, i_8_348, i_8_385, i_8_426, i_8_430, i_8_492, i_8_527, i_8_530, i_8_555, i_8_580, i_8_611, i_8_637, i_8_642, i_8_665, i_8_696, i_8_706, i_8_709, i_8_734, i_8_772, i_8_832, i_8_839, i_8_843, i_8_867, i_8_957, i_8_958, i_8_966, i_8_1041, i_8_1042, i_8_1072, i_8_1130, i_8_1146, i_8_1149, i_8_1160, i_8_1167, i_8_1182, i_8_1227, i_8_1237, i_8_1284, i_8_1285, i_8_1299, i_8_1318, i_8_1358, i_8_1362, i_8_1443, i_8_1447, i_8_1479, i_8_1480, i_8_1483, i_8_1488, i_8_1489, i_8_1490, i_8_1560, i_8_1565, i_8_1605, i_8_1608, i_8_1679, i_8_1686, i_8_1719, i_8_1725, i_8_1770, i_8_1785, i_8_1812, i_8_1824, i_8_1825, i_8_1947, i_8_1956, i_8_1959, i_8_1983, i_8_2056, i_8_2070, i_8_2074, i_8_2112, i_8_2113, i_8_2139, i_8_2140, i_8_2147, i_8_2154, i_8_2158, i_8_2193, i_8_2203, i_8_2227, i_8_2229, i_8_2232, i_8_2235, i_8_2239, i_8_2262, i_8_2263, i_8_2289, i_8_2292, o_8_214);
	kernel_8_215 k_8_215(i_8_53, i_8_58, i_8_101, i_8_107, i_8_210, i_8_227, i_8_232, i_8_256, i_8_323, i_8_361, i_8_362, i_8_364, i_8_365, i_8_373, i_8_400, i_8_426, i_8_442, i_8_454, i_8_553, i_8_571, i_8_660, i_8_676, i_8_679, i_8_699, i_8_700, i_8_703, i_8_710, i_8_759, i_8_838, i_8_841, i_8_859, i_8_877, i_8_887, i_8_968, i_8_970, i_8_1017, i_8_1067, i_8_1147, i_8_1189, i_8_1228, i_8_1229, i_8_1231, i_8_1281, i_8_1297, i_8_1300, i_8_1301, i_8_1308, i_8_1318, i_8_1339, i_8_1343, i_8_1344, i_8_1345, i_8_1363, i_8_1397, i_8_1400, i_8_1441, i_8_1467, i_8_1486, i_8_1489, i_8_1526, i_8_1559, i_8_1562, i_8_1574, i_8_1606, i_8_1607, i_8_1633, i_8_1672, i_8_1677, i_8_1678, i_8_1718, i_8_1720, i_8_1731, i_8_1738, i_8_1747, i_8_1748, i_8_1760, i_8_1763, i_8_1820, i_8_1834, i_8_1972, i_8_1982, i_8_1989, i_8_1996, i_8_2055, i_8_2056, i_8_2057, i_8_2107, i_8_2110, i_8_2111, i_8_2126, i_8_2147, i_8_2156, i_8_2172, i_8_2225, i_8_2226, i_8_2227, i_8_2230, i_8_2242, i_8_2248, i_8_2286, o_8_215);
	kernel_8_216 k_8_216(i_8_2, i_8_6, i_8_7, i_8_34, i_8_106, i_8_108, i_8_169, i_8_260, i_8_285, i_8_286, i_8_294, i_8_295, i_8_323, i_8_328, i_8_337, i_8_347, i_8_431, i_8_439, i_8_440, i_8_547, i_8_583, i_8_602, i_8_609, i_8_628, i_8_654, i_8_705, i_8_715, i_8_719, i_8_726, i_8_781, i_8_789, i_8_808, i_8_814, i_8_817, i_8_819, i_8_826, i_8_850, i_8_851, i_8_853, i_8_879, i_8_899, i_8_925, i_8_933, i_8_969, i_8_970, i_8_975, i_8_1074, i_8_1115, i_8_1133, i_8_1149, i_8_1185, i_8_1186, i_8_1192, i_8_1201, i_8_1267, i_8_1273, i_8_1281, i_8_1282, i_8_1284, i_8_1295, i_8_1300, i_8_1302, i_8_1339, i_8_1354, i_8_1385, i_8_1390, i_8_1411, i_8_1440, i_8_1444, i_8_1473, i_8_1489, i_8_1591, i_8_1614, i_8_1617, i_8_1628, i_8_1648, i_8_1653, i_8_1655, i_8_1663, i_8_1678, i_8_1754, i_8_1792, i_8_1849, i_8_1891, i_8_1898, i_8_2028, i_8_2031, i_8_2070, i_8_2137, i_8_2139, i_8_2140, i_8_2141, i_8_2147, i_8_2148, i_8_2150, i_8_2151, i_8_2154, i_8_2205, i_8_2220, i_8_2247, o_8_216);
	kernel_8_217 k_8_217(i_8_15, i_8_20, i_8_21, i_8_41, i_8_65, i_8_115, i_8_226, i_8_299, i_8_316, i_8_319, i_8_363, i_8_415, i_8_418, i_8_447, i_8_460, i_8_483, i_8_495, i_8_497, i_8_532, i_8_550, i_8_553, i_8_568, i_8_577, i_8_596, i_8_608, i_8_635, i_8_650, i_8_705, i_8_729, i_8_760, i_8_818, i_8_859, i_8_879, i_8_880, i_8_918, i_8_968, i_8_976, i_8_1126, i_8_1132, i_8_1153, i_8_1171, i_8_1188, i_8_1198, i_8_1202, i_8_1226, i_8_1231, i_8_1234, i_8_1235, i_8_1261, i_8_1276, i_8_1324, i_8_1325, i_8_1328, i_8_1342, i_8_1353, i_8_1360, i_8_1378, i_8_1388, i_8_1396, i_8_1397, i_8_1432, i_8_1436, i_8_1459, i_8_1463, i_8_1468, i_8_1491, i_8_1511, i_8_1541, i_8_1556, i_8_1630, i_8_1643, i_8_1648, i_8_1679, i_8_1694, i_8_1714, i_8_1759, i_8_1778, i_8_1792, i_8_1819, i_8_1826, i_8_1838, i_8_1861, i_8_1873, i_8_1883, i_8_1946, i_8_1947, i_8_1972, i_8_1990, i_8_2061, i_8_2062, i_8_2065, i_8_2144, i_8_2145, i_8_2169, i_8_2170, i_8_2224, i_8_2242, i_8_2268, i_8_2269, i_8_2273, o_8_217);
	kernel_8_218 k_8_218(i_8_11, i_8_13, i_8_19, i_8_23, i_8_28, i_8_68, i_8_86, i_8_100, i_8_114, i_8_115, i_8_116, i_8_117, i_8_142, i_8_194, i_8_210, i_8_274, i_8_279, i_8_348, i_8_378, i_8_379, i_8_391, i_8_428, i_8_507, i_8_508, i_8_544, i_8_589, i_8_622, i_8_642, i_8_650, i_8_693, i_8_694, i_8_708, i_8_732, i_8_733, i_8_764, i_8_781, i_8_851, i_8_872, i_8_874, i_8_880, i_8_896, i_8_921, i_8_937, i_8_955, i_8_990, i_8_1027, i_8_1107, i_8_1114, i_8_1130, i_8_1134, i_8_1137, i_8_1139, i_8_1146, i_8_1224, i_8_1225, i_8_1260, i_8_1261, i_8_1264, i_8_1300, i_8_1315, i_8_1396, i_8_1400, i_8_1410, i_8_1422, i_8_1432, i_8_1492, i_8_1549, i_8_1611, i_8_1612, i_8_1633, i_8_1648, i_8_1668, i_8_1671, i_8_1681, i_8_1710, i_8_1718, i_8_1723, i_8_1751, i_8_1756, i_8_1775, i_8_1778, i_8_1803, i_8_1824, i_8_1840, i_8_1859, i_8_1868, i_8_1869, i_8_1884, i_8_1945, i_8_1946, i_8_1957, i_8_1989, i_8_2001, i_8_2053, i_8_2099, i_8_2138, i_8_2152, i_8_2197, i_8_2215, i_8_2263, o_8_218);
	kernel_8_219 k_8_219(i_8_22, i_8_24, i_8_34, i_8_39, i_8_67, i_8_158, i_8_180, i_8_223, i_8_229, i_8_262, i_8_300, i_8_370, i_8_379, i_8_381, i_8_426, i_8_440, i_8_534, i_8_535, i_8_592, i_8_602, i_8_610, i_8_613, i_8_628, i_8_655, i_8_660, i_8_695, i_8_703, i_8_704, i_8_706, i_8_727, i_8_753, i_8_771, i_8_816, i_8_838, i_8_840, i_8_843, i_8_849, i_8_850, i_8_853, i_8_869, i_8_876, i_8_877, i_8_940, i_8_979, i_8_980, i_8_984, i_8_993, i_8_1074, i_8_1126, i_8_1137, i_8_1157, i_8_1224, i_8_1225, i_8_1226, i_8_1227, i_8_1234, i_8_1263, i_8_1338, i_8_1346, i_8_1362, i_8_1379, i_8_1427, i_8_1467, i_8_1470, i_8_1506, i_8_1547, i_8_1549, i_8_1560, i_8_1574, i_8_1606, i_8_1615, i_8_1617, i_8_1650, i_8_1677, i_8_1686, i_8_1706, i_8_1729, i_8_1755, i_8_1759, i_8_1760, i_8_1787, i_8_1813, i_8_1824, i_8_1885, i_8_1974, i_8_1976, i_8_1983, i_8_1989, i_8_2002, i_8_2136, i_8_2143, i_8_2144, i_8_2146, i_8_2149, i_8_2158, i_8_2190, i_8_2191, i_8_2215, i_8_2226, i_8_2236, o_8_219);
	kernel_8_220 k_8_220(i_8_5, i_8_20, i_8_89, i_8_194, i_8_197, i_8_220, i_8_224, i_8_227, i_8_302, i_8_328, i_8_346, i_8_356, i_8_376, i_8_383, i_8_385, i_8_386, i_8_445, i_8_455, i_8_464, i_8_476, i_8_499, i_8_500, i_8_508, i_8_525, i_8_526, i_8_529, i_8_553, i_8_589, i_8_593, i_8_607, i_8_625, i_8_662, i_8_665, i_8_671, i_8_715, i_8_716, i_8_725, i_8_780, i_8_781, i_8_782, i_8_787, i_8_789, i_8_795, i_8_796, i_8_814, i_8_825, i_8_877, i_8_904, i_8_1012, i_8_1015, i_8_1030, i_8_1031, i_8_1086, i_8_1087, i_8_1132, i_8_1190, i_8_1193, i_8_1237, i_8_1256, i_8_1345, i_8_1436, i_8_1456, i_8_1457, i_8_1471, i_8_1540, i_8_1542, i_8_1544, i_8_1552, i_8_1579, i_8_1588, i_8_1598, i_8_1601, i_8_1607, i_8_1633, i_8_1636, i_8_1679, i_8_1714, i_8_1717, i_8_1732, i_8_1742, i_8_1754, i_8_1763, i_8_1894, i_8_1895, i_8_1918, i_8_1919, i_8_1933, i_8_1951, i_8_1967, i_8_1981, i_8_2005, i_8_2029, i_8_2047, i_8_2109, i_8_2112, i_8_2129, i_8_2171, i_8_2196, i_8_2289, i_8_2290, o_8_220);
	kernel_8_221 k_8_221(i_8_26, i_8_31, i_8_41, i_8_57, i_8_68, i_8_95, i_8_98, i_8_107, i_8_166, i_8_167, i_8_176, i_8_179, i_8_215, i_8_227, i_8_229, i_8_260, i_8_266, i_8_314, i_8_338, i_8_359, i_8_363, i_8_374, i_8_386, i_8_427, i_8_428, i_8_431, i_8_449, i_8_455, i_8_487, i_8_494, i_8_522, i_8_539, i_8_589, i_8_593, i_8_653, i_8_656, i_8_661, i_8_665, i_8_693, i_8_694, i_8_699, i_8_702, i_8_706, i_8_710, i_8_771, i_8_809, i_8_838, i_8_842, i_8_869, i_8_881, i_8_948, i_8_959, i_8_965, i_8_966, i_8_1022, i_8_1024, i_8_1129, i_8_1166, i_8_1175, i_8_1231, i_8_1241, i_8_1268, i_8_1321, i_8_1337, i_8_1373, i_8_1376, i_8_1402, i_8_1419, i_8_1435, i_8_1453, i_8_1456, i_8_1472, i_8_1526, i_8_1546, i_8_1562, i_8_1646, i_8_1655, i_8_1672, i_8_1673, i_8_1691, i_8_1706, i_8_1790, i_8_1821, i_8_1822, i_8_1823, i_8_1825, i_8_1832, i_8_1868, i_8_1870, i_8_1930, i_8_1965, i_8_2077, i_8_2078, i_8_2113, i_8_2145, i_8_2227, i_8_2249, i_8_2267, i_8_2276, i_8_2285, o_8_221);
	kernel_8_222 k_8_222(i_8_33, i_8_35, i_8_98, i_8_157, i_8_160, i_8_161, i_8_221, i_8_224, i_8_301, i_8_354, i_8_369, i_8_373, i_8_374, i_8_433, i_8_434, i_8_440, i_8_462, i_8_463, i_8_475, i_8_476, i_8_478, i_8_498, i_8_508, i_8_526, i_8_530, i_8_548, i_8_595, i_8_660, i_8_707, i_8_715, i_8_716, i_8_735, i_8_777, i_8_781, i_8_793, i_8_796, i_8_823, i_8_880, i_8_985, i_8_996, i_8_1009, i_8_1011, i_8_1012, i_8_1027, i_8_1085, i_8_1120, i_8_1121, i_8_1249, i_8_1256, i_8_1273, i_8_1285, i_8_1300, i_8_1344, i_8_1453, i_8_1456, i_8_1469, i_8_1471, i_8_1536, i_8_1540, i_8_1543, i_8_1544, i_8_1552, i_8_1553, i_8_1558, i_8_1574, i_8_1579, i_8_1587, i_8_1589, i_8_1597, i_8_1598, i_8_1629, i_8_1669, i_8_1714, i_8_1752, i_8_1780, i_8_1781, i_8_1783, i_8_1785, i_8_1807, i_8_1821, i_8_1840, i_8_1857, i_8_1858, i_8_1894, i_8_1895, i_8_1930, i_8_1950, i_8_1951, i_8_1974, i_8_1975, i_8_2102, i_8_2111, i_8_2128, i_8_2183, i_8_2191, i_8_2216, i_8_2224, i_8_2275, i_8_2289, i_8_2295, o_8_222);
	kernel_8_223 k_8_223(i_8_11, i_8_52, i_8_53, i_8_70, i_8_79, i_8_95, i_8_111, i_8_112, i_8_188, i_8_221, i_8_250, i_8_256, i_8_297, i_8_301, i_8_305, i_8_346, i_8_348, i_8_349, i_8_360, i_8_362, i_8_363, i_8_364, i_8_365, i_8_366, i_8_368, i_8_479, i_8_555, i_8_557, i_8_615, i_8_625, i_8_635, i_8_658, i_8_688, i_8_762, i_8_770, i_8_816, i_8_817, i_8_837, i_8_838, i_8_843, i_8_844, i_8_859, i_8_860, i_8_862, i_8_863, i_8_877, i_8_879, i_8_880, i_8_881, i_8_938, i_8_942, i_8_943, i_8_944, i_8_978, i_8_1030, i_8_1045, i_8_1086, i_8_1087, i_8_1113, i_8_1138, i_8_1148, i_8_1203, i_8_1301, i_8_1302, i_8_1306, i_8_1307, i_8_1410, i_8_1455, i_8_1456, i_8_1511, i_8_1533, i_8_1535, i_8_1543, i_8_1546, i_8_1649, i_8_1651, i_8_1764, i_8_1807, i_8_1888, i_8_1915, i_8_1918, i_8_1997, i_8_2013, i_8_2046, i_8_2048, i_8_2051, i_8_2111, i_8_2112, i_8_2113, i_8_2119, i_8_2121, i_8_2123, i_8_2132, i_8_2140, i_8_2213, i_8_2215, i_8_2216, i_8_2298, i_8_2299, i_8_2300, o_8_223);
	kernel_8_224 k_8_224(i_8_38, i_8_58, i_8_71, i_8_76, i_8_83, i_8_181, i_8_185, i_8_244, i_8_305, i_8_317, i_8_320, i_8_322, i_8_323, i_8_365, i_8_424, i_8_425, i_8_426, i_8_525, i_8_532, i_8_534, i_8_542, i_8_556, i_8_603, i_8_610, i_8_614, i_8_634, i_8_635, i_8_638, i_8_657, i_8_676, i_8_679, i_8_697, i_8_703, i_8_706, i_8_707, i_8_752, i_8_753, i_8_790, i_8_806, i_8_844, i_8_866, i_8_889, i_8_890, i_8_951, i_8_956, i_8_974, i_8_984, i_8_987, i_8_1003, i_8_1056, i_8_1060, i_8_1115, i_8_1138, i_8_1152, i_8_1166, i_8_1167, i_8_1190, i_8_1201, i_8_1225, i_8_1238, i_8_1247, i_8_1273, i_8_1282, i_8_1399, i_8_1415, i_8_1433, i_8_1439, i_8_1456, i_8_1463, i_8_1491, i_8_1507, i_8_1527, i_8_1546, i_8_1561, i_8_1606, i_8_1617, i_8_1678, i_8_1714, i_8_1722, i_8_1744, i_8_1784, i_8_1787, i_8_1791, i_8_1822, i_8_1826, i_8_1949, i_8_1957, i_8_1966, i_8_1967, i_8_1982, i_8_1985, i_8_1996, i_8_2047, i_8_2144, i_8_2153, i_8_2156, i_8_2188, i_8_2200, i_8_2226, i_8_2302, o_8_224);
	kernel_8_225 k_8_225(i_8_12, i_8_58, i_8_111, i_8_137, i_8_142, i_8_190, i_8_193, i_8_198, i_8_238, i_8_254, i_8_289, i_8_311, i_8_346, i_8_373, i_8_379, i_8_390, i_8_414, i_8_417, i_8_439, i_8_450, i_8_487, i_8_493, i_8_555, i_8_596, i_8_610, i_8_642, i_8_645, i_8_649, i_8_660, i_8_679, i_8_695, i_8_699, i_8_705, i_8_766, i_8_783, i_8_786, i_8_840, i_8_844, i_8_845, i_8_876, i_8_929, i_8_967, i_8_970, i_8_995, i_8_1064, i_8_1182, i_8_1185, i_8_1224, i_8_1226, i_8_1240, i_8_1255, i_8_1285, i_8_1288, i_8_1289, i_8_1300, i_8_1310, i_8_1314, i_8_1351, i_8_1354, i_8_1362, i_8_1381, i_8_1387, i_8_1461, i_8_1472, i_8_1481, i_8_1515, i_8_1540, i_8_1542, i_8_1545, i_8_1546, i_8_1632, i_8_1666, i_8_1671, i_8_1684, i_8_1693, i_8_1694, i_8_1699, i_8_1706, i_8_1747, i_8_1749, i_8_1758, i_8_1807, i_8_1826, i_8_1831, i_8_1855, i_8_1867, i_8_1887, i_8_1992, i_8_1993, i_8_2014, i_8_2071, i_8_2133, i_8_2142, i_8_2146, i_8_2151, i_8_2158, i_8_2226, i_8_2244, i_8_2278, i_8_2290, o_8_225);
	kernel_8_226 k_8_226(i_8_53, i_8_80, i_8_114, i_8_115, i_8_120, i_8_123, i_8_228, i_8_371, i_8_381, i_8_382, i_8_428, i_8_451, i_8_454, i_8_481, i_8_511, i_8_570, i_8_571, i_8_575, i_8_590, i_8_599, i_8_605, i_8_636, i_8_658, i_8_660, i_8_663, i_8_747, i_8_835, i_8_873, i_8_886, i_8_887, i_8_990, i_8_1028, i_8_1031, i_8_1044, i_8_1048, i_8_1061, i_8_1072, i_8_1073, i_8_1074, i_8_1111, i_8_1164, i_8_1187, i_8_1227, i_8_1228, i_8_1229, i_8_1230, i_8_1231, i_8_1309, i_8_1331, i_8_1338, i_8_1356, i_8_1370, i_8_1403, i_8_1411, i_8_1434, i_8_1467, i_8_1470, i_8_1472, i_8_1474, i_8_1489, i_8_1556, i_8_1621, i_8_1632, i_8_1633, i_8_1635, i_8_1637, i_8_1654, i_8_1655, i_8_1659, i_8_1702, i_8_1704, i_8_1705, i_8_1736, i_8_1746, i_8_1747, i_8_1749, i_8_1751, i_8_1752, i_8_1764, i_8_1803, i_8_1820, i_8_1823, i_8_1857, i_8_1862, i_8_1945, i_8_1950, i_8_1983, i_8_1984, i_8_1985, i_8_2058, i_8_2073, i_8_2078, i_8_2125, i_8_2144, i_8_2172, i_8_2173, i_8_2218, i_8_2227, i_8_2248, i_8_2276, o_8_226);
	kernel_8_227 k_8_227(i_8_65, i_8_107, i_8_115, i_8_140, i_8_172, i_8_173, i_8_269, i_8_284, i_8_293, i_8_323, i_8_353, i_8_360, i_8_368, i_8_382, i_8_398, i_8_452, i_8_489, i_8_490, i_8_492, i_8_530, i_8_590, i_8_614, i_8_634, i_8_706, i_8_707, i_8_764, i_8_797, i_8_833, i_8_845, i_8_858, i_8_859, i_8_868, i_8_922, i_8_969, i_8_1057, i_8_1058, i_8_1073, i_8_1100, i_8_1127, i_8_1129, i_8_1225, i_8_1226, i_8_1229, i_8_1262, i_8_1264, i_8_1298, i_8_1317, i_8_1325, i_8_1328, i_8_1366, i_8_1405, i_8_1406, i_8_1411, i_8_1435, i_8_1436, i_8_1456, i_8_1462, i_8_1463, i_8_1473, i_8_1522, i_8_1547, i_8_1549, i_8_1556, i_8_1622, i_8_1623, i_8_1633, i_8_1640, i_8_1730, i_8_1748, i_8_1757, i_8_1777, i_8_1784, i_8_1796, i_8_1823, i_8_1825, i_8_1832, i_8_1849, i_8_1867, i_8_1904, i_8_1957, i_8_1958, i_8_1975, i_8_1994, i_8_1996, i_8_1997, i_8_2003, i_8_2017, i_8_2020, i_8_2099, i_8_2117, i_8_2144, i_8_2150, i_8_2201, i_8_2225, i_8_2226, i_8_2244, i_8_2246, i_8_2249, i_8_2260, i_8_2287, o_8_227);
	kernel_8_228 k_8_228(i_8_21, i_8_25, i_8_44, i_8_79, i_8_84, i_8_247, i_8_248, i_8_265, i_8_320, i_8_323, i_8_338, i_8_367, i_8_368, i_8_395, i_8_422, i_8_430, i_8_469, i_8_511, i_8_516, i_8_517, i_8_527, i_8_552, i_8_571, i_8_574, i_8_575, i_8_584, i_8_591, i_8_593, i_8_597, i_8_599, i_8_611, i_8_634, i_8_647, i_8_683, i_8_704, i_8_710, i_8_733, i_8_763, i_8_788, i_8_824, i_8_832, i_8_842, i_8_858, i_8_861, i_8_941, i_8_971, i_8_1016, i_8_1106, i_8_1114, i_8_1129, i_8_1189, i_8_1205, i_8_1240, i_8_1267, i_8_1300, i_8_1304, i_8_1305, i_8_1366, i_8_1367, i_8_1403, i_8_1408, i_8_1410, i_8_1465, i_8_1466, i_8_1516, i_8_1517, i_8_1528, i_8_1533, i_8_1540, i_8_1588, i_8_1591, i_8_1653, i_8_1654, i_8_1691, i_8_1700, i_8_1750, i_8_1843, i_8_1844, i_8_1857, i_8_1868, i_8_1873, i_8_1876, i_8_1878, i_8_1886, i_8_1898, i_8_1916, i_8_1917, i_8_2011, i_8_2040, i_8_2048, i_8_2065, i_8_2128, i_8_2163, i_8_2173, i_8_2214, i_8_2231, i_8_2244, i_8_2245, i_8_2290, i_8_2298, o_8_228);
	kernel_8_229 k_8_229(i_8_40, i_8_59, i_8_64, i_8_83, i_8_104, i_8_140, i_8_163, i_8_220, i_8_221, i_8_229, i_8_247, i_8_281, i_8_283, i_8_326, i_8_363, i_8_364, i_8_381, i_8_434, i_8_451, i_8_481, i_8_487, i_8_504, i_8_505, i_8_522, i_8_524, i_8_526, i_8_527, i_8_528, i_8_589, i_8_594, i_8_598, i_8_609, i_8_610, i_8_623, i_8_659, i_8_662, i_8_685, i_8_689, i_8_694, i_8_696, i_8_706, i_8_716, i_8_725, i_8_760, i_8_823, i_8_838, i_8_845, i_8_996, i_8_1072, i_8_1100, i_8_1103, i_8_1180, i_8_1225, i_8_1234, i_8_1300, i_8_1309, i_8_1310, i_8_1352, i_8_1434, i_8_1438, i_8_1439, i_8_1589, i_8_1616, i_8_1625, i_8_1643, i_8_1674, i_8_1682, i_8_1720, i_8_1751, i_8_1752, i_8_1753, i_8_1771, i_8_1778, i_8_1810, i_8_1840, i_8_1856, i_8_1885, i_8_1901, i_8_1936, i_8_1949, i_8_1950, i_8_1968, i_8_1969, i_8_1990, i_8_2029, i_8_2041, i_8_2068, i_8_2089, i_8_2092, i_8_2129, i_8_2152, i_8_2153, i_8_2171, i_8_2173, i_8_2236, i_8_2237, i_8_2241, i_8_2246, i_8_2260, i_8_2261, o_8_229);
	kernel_8_230 k_8_230(i_8_43, i_8_96, i_8_114, i_8_140, i_8_143, i_8_156, i_8_158, i_8_185, i_8_188, i_8_217, i_8_218, i_8_224, i_8_227, i_8_253, i_8_301, i_8_329, i_8_414, i_8_461, i_8_482, i_8_485, i_8_489, i_8_496, i_8_505, i_8_522, i_8_523, i_8_524, i_8_525, i_8_528, i_8_530, i_8_592, i_8_609, i_8_614, i_8_624, i_8_630, i_8_632, i_8_661, i_8_696, i_8_697, i_8_700, i_8_701, i_8_711, i_8_713, i_8_714, i_8_715, i_8_716, i_8_719, i_8_768, i_8_812, i_8_837, i_8_839, i_8_840, i_8_1012, i_8_1121, i_8_1180, i_8_1181, i_8_1263, i_8_1284, i_8_1286, i_8_1297, i_8_1346, i_8_1382, i_8_1407, i_8_1411, i_8_1412, i_8_1504, i_8_1506, i_8_1624, i_8_1649, i_8_1651, i_8_1652, i_8_1655, i_8_1678, i_8_1747, i_8_1748, i_8_1749, i_8_1754, i_8_1825, i_8_1855, i_8_1881, i_8_1882, i_8_1901, i_8_1903, i_8_1981, i_8_1985, i_8_1992, i_8_1997, i_8_1999, i_8_2031, i_8_2037, i_8_2053, i_8_2056, i_8_2057, i_8_2089, i_8_2090, i_8_2143, i_8_2144, i_8_2150, i_8_2174, i_8_2218, i_8_2246, o_8_230);
	kernel_8_231 k_8_231(i_8_27, i_8_28, i_8_49, i_8_70, i_8_94, i_8_147, i_8_166, i_8_184, i_8_196, i_8_233, i_8_241, i_8_311, i_8_322, i_8_337, i_8_346, i_8_381, i_8_431, i_8_447, i_8_454, i_8_492, i_8_493, i_8_570, i_8_583, i_8_609, i_8_610, i_8_634, i_8_659, i_8_699, i_8_701, i_8_732, i_8_735, i_8_753, i_8_777, i_8_798, i_8_799, i_8_834, i_8_835, i_8_843, i_8_925, i_8_931, i_8_959, i_8_967, i_8_973, i_8_990, i_8_991, i_8_1020, i_8_1033, i_8_1059, i_8_1060, i_8_1102, i_8_1156, i_8_1236, i_8_1237, i_8_1263, i_8_1273, i_8_1296, i_8_1300, i_8_1373, i_8_1381, i_8_1407, i_8_1474, i_8_1488, i_8_1489, i_8_1491, i_8_1501, i_8_1564, i_8_1605, i_8_1606, i_8_1627, i_8_1628, i_8_1650, i_8_1661, i_8_1681, i_8_1705, i_8_1722, i_8_1758, i_8_1770, i_8_1826, i_8_1857, i_8_1884, i_8_1906, i_8_1969, i_8_2002, i_8_2004, i_8_2016, i_8_2046, i_8_2047, i_8_2102, i_8_2112, i_8_2145, i_8_2149, i_8_2163, i_8_2167, i_8_2173, i_8_2174, i_8_2208, i_8_2275, i_8_2281, i_8_2289, i_8_2298, o_8_231);
	kernel_8_232 k_8_232(i_8_22, i_8_23, i_8_31, i_8_34, i_8_35, i_8_85, i_8_106, i_8_107, i_8_232, i_8_247, i_8_295, i_8_345, i_8_346, i_8_348, i_8_386, i_8_394, i_8_426, i_8_443, i_8_458, i_8_480, i_8_482, i_8_524, i_8_526, i_8_527, i_8_529, i_8_554, i_8_555, i_8_602, i_8_609, i_8_611, i_8_628, i_8_631, i_8_633, i_8_634, i_8_707, i_8_732, i_8_761, i_8_763, i_8_771, i_8_783, i_8_799, i_8_800, i_8_811, i_8_814, i_8_815, i_8_838, i_8_931, i_8_934, i_8_965, i_8_986, i_8_991, i_8_1120, i_8_1189, i_8_1194, i_8_1219, i_8_1220, i_8_1223, i_8_1266, i_8_1267, i_8_1284, i_8_1311, i_8_1388, i_8_1391, i_8_1441, i_8_1525, i_8_1526, i_8_1535, i_8_1544, i_8_1545, i_8_1550, i_8_1554, i_8_1561, i_8_1633, i_8_1651, i_8_1676, i_8_1699, i_8_1722, i_8_1726, i_8_1733, i_8_1738, i_8_1740, i_8_1741, i_8_1748, i_8_1749, i_8_1753, i_8_1807, i_8_1819, i_8_1858, i_8_1867, i_8_1876, i_8_1897, i_8_1906, i_8_1956, i_8_1957, i_8_2150, i_8_2154, i_8_2215, i_8_2216, i_8_2218, i_8_2292, o_8_232);
	kernel_8_233 k_8_233(i_8_31, i_8_41, i_8_88, i_8_89, i_8_187, i_8_212, i_8_223, i_8_256, i_8_266, i_8_269, i_8_283, i_8_293, i_8_302, i_8_337, i_8_349, i_8_353, i_8_374, i_8_453, i_8_494, i_8_538, i_8_539, i_8_547, i_8_556, i_8_565, i_8_593, i_8_602, i_8_607, i_8_658, i_8_661, i_8_716, i_8_744, i_8_763, i_8_766, i_8_767, i_8_773, i_8_797, i_8_826, i_8_827, i_8_849, i_8_853, i_8_877, i_8_878, i_8_935, i_8_980, i_8_985, i_8_988, i_8_1012, i_8_1018, i_8_1030, i_8_1033, i_8_1041, i_8_1051, i_8_1069, i_8_1075, i_8_1091, i_8_1128, i_8_1129, i_8_1133, i_8_1139, i_8_1157, i_8_1226, i_8_1231, i_8_1237, i_8_1238, i_8_1249, i_8_1256, i_8_1262, i_8_1281, i_8_1318, i_8_1358, i_8_1363, i_8_1385, i_8_1453, i_8_1457, i_8_1543, i_8_1581, i_8_1627, i_8_1640, i_8_1652, i_8_1666, i_8_1700, i_8_1705, i_8_1708, i_8_1806, i_8_1855, i_8_1858, i_8_1868, i_8_1966, i_8_1995, i_8_1996, i_8_1997, i_8_2142, i_8_2158, i_8_2233, i_8_2268, i_8_2272, i_8_2273, i_8_2278, i_8_2282, i_8_2290, o_8_233);
	kernel_8_234 k_8_234(i_8_3, i_8_4, i_8_23, i_8_31, i_8_76, i_8_85, i_8_86, i_8_89, i_8_116, i_8_244, i_8_247, i_8_265, i_8_292, i_8_301, i_8_322, i_8_361, i_8_366, i_8_387, i_8_440, i_8_463, i_8_481, i_8_516, i_8_517, i_8_527, i_8_538, i_8_571, i_8_588, i_8_594, i_8_598, i_8_599, i_8_611, i_8_634, i_8_642, i_8_651, i_8_658, i_8_669, i_8_678, i_8_727, i_8_778, i_8_804, i_8_823, i_8_859, i_8_877, i_8_913, i_8_958, i_8_1012, i_8_1070, i_8_1210, i_8_1228, i_8_1239, i_8_1270, i_8_1390, i_8_1438, i_8_1439, i_8_1471, i_8_1489, i_8_1517, i_8_1533, i_8_1534, i_8_1571, i_8_1587, i_8_1588, i_8_1651, i_8_1659, i_8_1679, i_8_1702, i_8_1703, i_8_1706, i_8_1759, i_8_1763, i_8_1794, i_8_1795, i_8_1798, i_8_1820, i_8_1821, i_8_1822, i_8_1823, i_8_1840, i_8_1849, i_8_1876, i_8_1885, i_8_1903, i_8_1918, i_8_1948, i_8_1966, i_8_1967, i_8_1995, i_8_2028, i_8_2037, i_8_2053, i_8_2065, i_8_2119, i_8_2120, i_8_2154, i_8_2225, i_8_2226, i_8_2229, i_8_2256, i_8_2257, i_8_2281, o_8_234);
	kernel_8_235 k_8_235(i_8_16, i_8_53, i_8_111, i_8_148, i_8_194, i_8_227, i_8_230, i_8_259, i_8_260, i_8_283, i_8_383, i_8_401, i_8_417, i_8_427, i_8_493, i_8_508, i_8_556, i_8_574, i_8_575, i_8_579, i_8_591, i_8_592, i_8_598, i_8_599, i_8_665, i_8_706, i_8_751, i_8_786, i_8_798, i_8_826, i_8_838, i_8_841, i_8_977, i_8_984, i_8_1101, i_8_1102, i_8_1105, i_8_1108, i_8_1240, i_8_1270, i_8_1273, i_8_1274, i_8_1302, i_8_1330, i_8_1384, i_8_1385, i_8_1392, i_8_1396, i_8_1409, i_8_1433, i_8_1437, i_8_1439, i_8_1464, i_8_1483, i_8_1513, i_8_1519, i_8_1528, i_8_1552, i_8_1573, i_8_1574, i_8_1605, i_8_1606, i_8_1631, i_8_1632, i_8_1642, i_8_1671, i_8_1696, i_8_1699, i_8_1704, i_8_1707, i_8_1716, i_8_1732, i_8_1750, i_8_1768, i_8_1770, i_8_1791, i_8_1807, i_8_1813, i_8_1820, i_8_1888, i_8_1944, i_8_1945, i_8_1950, i_8_1954, i_8_1957, i_8_1960, i_8_1966, i_8_1975, i_8_1996, i_8_2056, i_8_2059, i_8_2093, i_8_2096, i_8_2134, i_8_2135, i_8_2157, i_8_2164, i_8_2214, i_8_2219, i_8_2257, o_8_235);
	kernel_8_236 k_8_236(i_8_36, i_8_37, i_8_64, i_8_112, i_8_166, i_8_167, i_8_193, i_8_194, i_8_221, i_8_226, i_8_300, i_8_362, i_8_373, i_8_385, i_8_397, i_8_420, i_8_421, i_8_484, i_8_489, i_8_493, i_8_522, i_8_525, i_8_526, i_8_529, i_8_606, i_8_607, i_8_608, i_8_613, i_8_662, i_8_698, i_8_700, i_8_701, i_8_707, i_8_710, i_8_801, i_8_802, i_8_803, i_8_806, i_8_809, i_8_843, i_8_844, i_8_854, i_8_932, i_8_935, i_8_972, i_8_993, i_8_995, i_8_1040, i_8_1047, i_8_1078, i_8_1113, i_8_1114, i_8_1115, i_8_1134, i_8_1233, i_8_1234, i_8_1259, i_8_1269, i_8_1271, i_8_1283, i_8_1286, i_8_1404, i_8_1489, i_8_1490, i_8_1507, i_8_1529, i_8_1585, i_8_1621, i_8_1624, i_8_1634, i_8_1650, i_8_1668, i_8_1678, i_8_1682, i_8_1710, i_8_1711, i_8_1748, i_8_1766, i_8_1775, i_8_1776, i_8_1777, i_8_1824, i_8_1854, i_8_1855, i_8_1862, i_8_1868, i_8_1881, i_8_1984, i_8_2021, i_8_2034, i_8_2035, i_8_2037, i_8_2039, i_8_2041, i_8_2092, i_8_2099, i_8_2147, i_8_2174, i_8_2237, i_8_2268, o_8_236);
	kernel_8_237 k_8_237(i_8_23, i_8_31, i_8_136, i_8_189, i_8_262, i_8_265, i_8_266, i_8_340, i_8_373, i_8_381, i_8_394, i_8_421, i_8_426, i_8_430, i_8_453, i_8_454, i_8_455, i_8_492, i_8_528, i_8_547, i_8_554, i_8_604, i_8_616, i_8_633, i_8_634, i_8_654, i_8_658, i_8_660, i_8_661, i_8_663, i_8_706, i_8_717, i_8_719, i_8_778, i_8_840, i_8_841, i_8_880, i_8_881, i_8_903, i_8_967, i_8_970, i_8_994, i_8_1024, i_8_1074, i_8_1081, i_8_1111, i_8_1121, i_8_1122, i_8_1129, i_8_1131, i_8_1198, i_8_1237, i_8_1249, i_8_1289, i_8_1292, i_8_1294, i_8_1321, i_8_1326, i_8_1357, i_8_1431, i_8_1434, i_8_1450, i_8_1471, i_8_1484, i_8_1489, i_8_1504, i_8_1519, i_8_1538, i_8_1542, i_8_1605, i_8_1625, i_8_1630, i_8_1632, i_8_1705, i_8_1743, i_8_1745, i_8_1749, i_8_1752, i_8_1753, i_8_1790, i_8_1804, i_8_1805, i_8_1813, i_8_1822, i_8_1823, i_8_1843, i_8_1849, i_8_1894, i_8_1922, i_8_1927, i_8_1947, i_8_1965, i_8_1992, i_8_2044, i_8_2093, i_8_2101, i_8_2146, i_8_2271, i_8_2289, i_8_2302, o_8_237);
	kernel_8_238 k_8_238(i_8_111, i_8_117, i_8_120, i_8_165, i_8_166, i_8_169, i_8_187, i_8_265, i_8_283, i_8_289, i_8_290, i_8_291, i_8_297, i_8_319, i_8_321, i_8_366, i_8_367, i_8_368, i_8_433, i_8_436, i_8_499, i_8_546, i_8_555, i_8_588, i_8_606, i_8_635, i_8_642, i_8_672, i_8_673, i_8_674, i_8_678, i_8_695, i_8_708, i_8_724, i_8_726, i_8_727, i_8_781, i_8_783, i_8_804, i_8_805, i_8_810, i_8_811, i_8_813, i_8_814, i_8_829, i_8_849, i_8_877, i_8_964, i_8_967, i_8_973, i_8_1011, i_8_1029, i_8_1030, i_8_1032, i_8_1119, i_8_1200, i_8_1239, i_8_1264, i_8_1299, i_8_1324, i_8_1345, i_8_1351, i_8_1441, i_8_1452, i_8_1491, i_8_1507, i_8_1533, i_8_1542, i_8_1546, i_8_1578, i_8_1587, i_8_1588, i_8_1623, i_8_1731, i_8_1749, i_8_1767, i_8_1770, i_8_1779, i_8_1782, i_8_1821, i_8_1824, i_8_1825, i_8_1846, i_8_1848, i_8_1851, i_8_1876, i_8_1903, i_8_1938, i_8_1993, i_8_1996, i_8_2029, i_8_2031, i_8_2037, i_8_2038, i_8_2074, i_8_2116, i_8_2128, i_8_2150, i_8_2190, i_8_2272, o_8_238);
	kernel_8_239 k_8_239(i_8_23, i_8_31, i_8_32, i_8_34, i_8_165, i_8_201, i_8_225, i_8_263, i_8_265, i_8_279, i_8_318, i_8_335, i_8_365, i_8_368, i_8_417, i_8_443, i_8_447, i_8_451, i_8_452, i_8_483, i_8_525, i_8_530, i_8_533, i_8_615, i_8_616, i_8_631, i_8_688, i_8_689, i_8_704, i_8_717, i_8_772, i_8_831, i_8_842, i_8_874, i_8_875, i_8_938, i_8_970, i_8_1054, i_8_1057, i_8_1075, i_8_1077, i_8_1078, i_8_1099, i_8_1225, i_8_1228, i_8_1246, i_8_1247, i_8_1261, i_8_1282, i_8_1305, i_8_1309, i_8_1385, i_8_1407, i_8_1410, i_8_1423, i_8_1435, i_8_1436, i_8_1437, i_8_1469, i_8_1472, i_8_1536, i_8_1562, i_8_1567, i_8_1591, i_8_1598, i_8_1607, i_8_1622, i_8_1626, i_8_1654, i_8_1675, i_8_1684, i_8_1702, i_8_1722, i_8_1723, i_8_1752, i_8_1810, i_8_1825, i_8_1837, i_8_1838, i_8_1841, i_8_1868, i_8_1870, i_8_1901, i_8_1930, i_8_1967, i_8_2045, i_8_2117, i_8_2126, i_8_2129, i_8_2143, i_8_2144, i_8_2209, i_8_2212, i_8_2214, i_8_2242, i_8_2246, i_8_2257, i_8_2264, i_8_2292, i_8_2303, o_8_239);
	kernel_8_240 k_8_240(i_8_11, i_8_84, i_8_87, i_8_96, i_8_97, i_8_102, i_8_107, i_8_222, i_8_223, i_8_240, i_8_255, i_8_282, i_8_300, i_8_301, i_8_375, i_8_444, i_8_453, i_8_454, i_8_475, i_8_483, i_8_485, i_8_555, i_8_588, i_8_596, i_8_601, i_8_613, i_8_621, i_8_714, i_8_717, i_8_720, i_8_759, i_8_771, i_8_780, i_8_795, i_8_811, i_8_813, i_8_825, i_8_840, i_8_889, i_8_972, i_8_1014, i_8_1026, i_8_1029, i_8_1049, i_8_1111, i_8_1113, i_8_1135, i_8_1137, i_8_1233, i_8_1255, i_8_1257, i_8_1281, i_8_1313, i_8_1438, i_8_1443, i_8_1482, i_8_1533, i_8_1534, i_8_1541, i_8_1542, i_8_1548, i_8_1555, i_8_1587, i_8_1588, i_8_1590, i_8_1668, i_8_1677, i_8_1725, i_8_1753, i_8_1761, i_8_1762, i_8_1780, i_8_1785, i_8_1788, i_8_1812, i_8_1813, i_8_1840, i_8_1867, i_8_1893, i_8_1914, i_8_1918, i_8_1923, i_8_1968, i_8_1969, i_8_1974, i_8_1995, i_8_2001, i_8_2031, i_8_2046, i_8_2050, i_8_2054, i_8_2130, i_8_2136, i_8_2181, i_8_2214, i_8_2215, i_8_2263, i_8_2271, i_8_2272, i_8_2284, o_8_240);
	kernel_8_241 k_8_241(i_8_36, i_8_63, i_8_189, i_8_190, i_8_191, i_8_192, i_8_193, i_8_194, i_8_223, i_8_237, i_8_238, i_8_258, i_8_300, i_8_325, i_8_327, i_8_328, i_8_360, i_8_393, i_8_529, i_8_615, i_8_618, i_8_624, i_8_628, i_8_665, i_8_689, i_8_696, i_8_716, i_8_781, i_8_837, i_8_842, i_8_844, i_8_849, i_8_853, i_8_861, i_8_862, i_8_874, i_8_875, i_8_877, i_8_878, i_8_937, i_8_939, i_8_970, i_8_996, i_8_1014, i_8_1015, i_8_1029, i_8_1030, i_8_1038, i_8_1050, i_8_1158, i_8_1231, i_8_1240, i_8_1263, i_8_1267, i_8_1269, i_8_1284, i_8_1285, i_8_1290, i_8_1291, i_8_1294, i_8_1315, i_8_1407, i_8_1408, i_8_1437, i_8_1444, i_8_1473, i_8_1492, i_8_1510, i_8_1530, i_8_1545, i_8_1546, i_8_1638, i_8_1647, i_8_1648, i_8_1651, i_8_1680, i_8_1700, i_8_1750, i_8_1768, i_8_1769, i_8_1779, i_8_1815, i_8_1822, i_8_1827, i_8_1830, i_8_1844, i_8_1881, i_8_1883, i_8_2037, i_8_2040, i_8_2070, i_8_2091, i_8_2156, i_8_2157, i_8_2158, i_8_2173, i_8_2218, i_8_2238, i_8_2239, i_8_2262, o_8_241);
	kernel_8_242 k_8_242(i_8_67, i_8_75, i_8_76, i_8_120, i_8_125, i_8_138, i_8_169, i_8_192, i_8_195, i_8_196, i_8_198, i_8_225, i_8_228, i_8_229, i_8_261, i_8_301, i_8_312, i_8_324, i_8_354, i_8_355, i_8_402, i_8_417, i_8_433, i_8_522, i_8_556, i_8_571, i_8_586, i_8_588, i_8_634, i_8_657, i_8_660, i_8_671, i_8_672, i_8_697, i_8_709, i_8_732, i_8_747, i_8_753, i_8_782, i_8_831, i_8_835, i_8_837, i_8_838, i_8_840, i_8_858, i_8_925, i_8_943, i_8_969, i_8_970, i_8_971, i_8_973, i_8_983, i_8_985, i_8_990, i_8_993, i_8_1003, i_8_1038, i_8_1129, i_8_1138, i_8_1144, i_8_1266, i_8_1282, i_8_1293, i_8_1299, i_8_1300, i_8_1368, i_8_1390, i_8_1445, i_8_1452, i_8_1457, i_8_1470, i_8_1480, i_8_1486, i_8_1524, i_8_1549, i_8_1551, i_8_1573, i_8_1605, i_8_1633, i_8_1641, i_8_1651, i_8_1663, i_8_1849, i_8_1857, i_8_1922, i_8_1938, i_8_1946, i_8_1965, i_8_1968, i_8_1983, i_8_1995, i_8_2025, i_8_2053, i_8_2073, i_8_2082, i_8_2146, i_8_2191, i_8_2232, i_8_2233, i_8_2276, o_8_242);
	kernel_8_243 k_8_243(i_8_39, i_8_42, i_8_49, i_8_58, i_8_82, i_8_115, i_8_117, i_8_148, i_8_151, i_8_166, i_8_221, i_8_241, i_8_273, i_8_275, i_8_343, i_8_356, i_8_370, i_8_432, i_8_444, i_8_453, i_8_461, i_8_476, i_8_477, i_8_517, i_8_523, i_8_524, i_8_545, i_8_621, i_8_667, i_8_668, i_8_712, i_8_760, i_8_769, i_8_776, i_8_790, i_8_805, i_8_813, i_8_861, i_8_868, i_8_923, i_8_944, i_8_993, i_8_1160, i_8_1184, i_8_1201, i_8_1254, i_8_1281, i_8_1282, i_8_1300, i_8_1301, i_8_1356, i_8_1382, i_8_1387, i_8_1435, i_8_1497, i_8_1498, i_8_1535, i_8_1542, i_8_1543, i_8_1585, i_8_1587, i_8_1588, i_8_1595, i_8_1604, i_8_1622, i_8_1650, i_8_1676, i_8_1681, i_8_1688, i_8_1720, i_8_1753, i_8_1759, i_8_1762, i_8_1808, i_8_1814, i_8_1848, i_8_1855, i_8_1872, i_8_1886, i_8_1945, i_8_1946, i_8_1982, i_8_1993, i_8_2001, i_8_2028, i_8_2041, i_8_2072, i_8_2073, i_8_2093, i_8_2107, i_8_2108, i_8_2122, i_8_2123, i_8_2126, i_8_2174, i_8_2245, i_8_2246, i_8_2271, i_8_2299, i_8_2300, o_8_243);
	kernel_8_244 k_8_244(i_8_0, i_8_78, i_8_84, i_8_94, i_8_103, i_8_120, i_8_126, i_8_135, i_8_156, i_8_184, i_8_190, i_8_217, i_8_255, i_8_297, i_8_328, i_8_364, i_8_381, i_8_451, i_8_454, i_8_480, i_8_493, i_8_525, i_8_544, i_8_549, i_8_553, i_8_561, i_8_580, i_8_589, i_8_595, i_8_610, i_8_622, i_8_628, i_8_631, i_8_640, i_8_661, i_8_679, i_8_682, i_8_715, i_8_718, i_8_733, i_8_786, i_8_792, i_8_832, i_8_841, i_8_842, i_8_847, i_8_850, i_8_911, i_8_964, i_8_967, i_8_976, i_8_1071, i_8_1072, i_8_1108, i_8_1111, i_8_1210, i_8_1255, i_8_1257, i_8_1264, i_8_1266, i_8_1270, i_8_1279, i_8_1297, i_8_1321, i_8_1326, i_8_1416, i_8_1435, i_8_1437, i_8_1438, i_8_1450, i_8_1453, i_8_1465, i_8_1551, i_8_1563, i_8_1564, i_8_1593, i_8_1625, i_8_1680, i_8_1722, i_8_1759, i_8_1762, i_8_1764, i_8_1802, i_8_1805, i_8_1809, i_8_1995, i_8_2026, i_8_2053, i_8_2116, i_8_2119, i_8_2125, i_8_2128, i_8_2223, i_8_2233, i_8_2242, i_8_2275, i_8_2280, i_8_2283, i_8_2286, i_8_2290, o_8_244);
	kernel_8_245 k_8_245(i_8_32, i_8_76, i_8_167, i_8_173, i_8_209, i_8_256, i_8_262, i_8_326, i_8_344, i_8_362, i_8_364, i_8_365, i_8_425, i_8_434, i_8_454, i_8_482, i_8_491, i_8_553, i_8_590, i_8_626, i_8_634, i_8_641, i_8_703, i_8_706, i_8_707, i_8_738, i_8_767, i_8_795, i_8_837, i_8_839, i_8_842, i_8_845, i_8_919, i_8_920, i_8_929, i_8_956, i_8_1055, i_8_1061, i_8_1067, i_8_1100, i_8_1114, i_8_1171, i_8_1172, i_8_1235, i_8_1264, i_8_1278, i_8_1282, i_8_1283, i_8_1316, i_8_1372, i_8_1379, i_8_1382, i_8_1413, i_8_1433, i_8_1478, i_8_1544, i_8_1559, i_8_1562, i_8_1565, i_8_1571, i_8_1613, i_8_1625, i_8_1633, i_8_1643, i_8_1685, i_8_1688, i_8_1694, i_8_1702, i_8_1703, i_8_1706, i_8_1711, i_8_1721, i_8_1765, i_8_1774, i_8_1775, i_8_1820, i_8_1821, i_8_1822, i_8_1832, i_8_1859, i_8_1863, i_8_1867, i_8_1882, i_8_1883, i_8_1982, i_8_2009, i_8_2017, i_8_2018, i_8_2108, i_8_2111, i_8_2144, i_8_2146, i_8_2147, i_8_2170, i_8_2192, i_8_2197, i_8_2198, i_8_2206, i_8_2242, i_8_2243, o_8_245);
	kernel_8_246 k_8_246(i_8_114, i_8_186, i_8_241, i_8_294, i_8_295, i_8_296, i_8_303, i_8_304, i_8_321, i_8_337, i_8_348, i_8_350, i_8_364, i_8_453, i_8_458, i_8_488, i_8_553, i_8_554, i_8_590, i_8_597, i_8_599, i_8_613, i_8_614, i_8_615, i_8_617, i_8_619, i_8_645, i_8_672, i_8_689, i_8_705, i_8_710, i_8_717, i_8_778, i_8_799, i_8_851, i_8_872, i_8_875, i_8_878, i_8_969, i_8_970, i_8_990, i_8_991, i_8_1031, i_8_1072, i_8_1074, i_8_1108, i_8_1112, i_8_1113, i_8_1119, i_8_1120, i_8_1121, i_8_1122, i_8_1123, i_8_1124, i_8_1229, i_8_1282, i_8_1306, i_8_1329, i_8_1330, i_8_1331, i_8_1407, i_8_1408, i_8_1411, i_8_1437, i_8_1489, i_8_1490, i_8_1509, i_8_1511, i_8_1545, i_8_1619, i_8_1650, i_8_1654, i_8_1672, i_8_1675, i_8_1677, i_8_1679, i_8_1790, i_8_1803, i_8_1806, i_8_1815, i_8_1823, i_8_1826, i_8_1866, i_8_1876, i_8_1884, i_8_1885, i_8_1983, i_8_1986, i_8_1988, i_8_2028, i_8_2056, i_8_2075, i_8_2090, i_8_2131, i_8_2193, i_8_2194, i_8_2219, i_8_2228, i_8_2249, i_8_2272, o_8_246);
	kernel_8_247 k_8_247(i_8_52, i_8_76, i_8_80, i_8_104, i_8_107, i_8_166, i_8_169, i_8_219, i_8_225, i_8_228, i_8_257, i_8_323, i_8_368, i_8_382, i_8_427, i_8_436, i_8_440, i_8_450, i_8_489, i_8_490, i_8_491, i_8_492, i_8_548, i_8_556, i_8_581, i_8_587, i_8_626, i_8_635, i_8_658, i_8_661, i_8_679, i_8_693, i_8_694, i_8_695, i_8_698, i_8_699, i_8_716, i_8_723, i_8_724, i_8_725, i_8_805, i_8_809, i_8_812, i_8_833, i_8_840, i_8_851, i_8_955, i_8_970, i_8_977, i_8_1031, i_8_1076, i_8_1111, i_8_1115, i_8_1184, i_8_1192, i_8_1210, i_8_1211, i_8_1226, i_8_1234, i_8_1255, i_8_1273, i_8_1280, i_8_1300, i_8_1301, i_8_1328, i_8_1360, i_8_1373, i_8_1391, i_8_1456, i_8_1471, i_8_1472, i_8_1577, i_8_1748, i_8_1773, i_8_1786, i_8_1789, i_8_1790, i_8_1818, i_8_1849, i_8_1850, i_8_1858, i_8_1867, i_8_1901, i_8_1904, i_8_1907, i_8_1979, i_8_1982, i_8_1996, i_8_2003, i_8_2029, i_8_2032, i_8_2038, i_8_2133, i_8_2134, i_8_2191, i_8_2200, i_8_2214, i_8_2223, i_8_2224, i_8_2273, o_8_247);
	kernel_8_248 k_8_248(i_8_31, i_8_39, i_8_42, i_8_51, i_8_55, i_8_96, i_8_97, i_8_169, i_8_256, i_8_258, i_8_300, i_8_307, i_8_319, i_8_331, i_8_334, i_8_360, i_8_363, i_8_417, i_8_418, i_8_421, i_8_440, i_8_481, i_8_483, i_8_484, i_8_529, i_8_587, i_8_588, i_8_601, i_8_628, i_8_653, i_8_661, i_8_669, i_8_680, i_8_691, i_8_707, i_8_747, i_8_748, i_8_786, i_8_789, i_8_823, i_8_839, i_8_842, i_8_844, i_8_845, i_8_868, i_8_894, i_8_993, i_8_994, i_8_996, i_8_1039, i_8_1050, i_8_1074, i_8_1075, i_8_1110, i_8_1112, i_8_1202, i_8_1227, i_8_1270, i_8_1274, i_8_1278, i_8_1282, i_8_1300, i_8_1307, i_8_1308, i_8_1359, i_8_1456, i_8_1462, i_8_1474, i_8_1507, i_8_1511, i_8_1516, i_8_1525, i_8_1540, i_8_1558, i_8_1561, i_8_1572, i_8_1633, i_8_1720, i_8_1726, i_8_1740, i_8_1749, i_8_1753, i_8_1775, i_8_1783, i_8_1796, i_8_1810, i_8_1828, i_8_1876, i_8_1906, i_8_1969, i_8_1991, i_8_2031, i_8_2136, i_8_2154, i_8_2191, i_8_2214, i_8_2218, i_8_2236, i_8_2243, i_8_2293, o_8_248);
	kernel_8_249 k_8_249(i_8_35, i_8_48, i_8_49, i_8_50, i_8_51, i_8_52, i_8_53, i_8_58, i_8_97, i_8_163, i_8_164, i_8_167, i_8_185, i_8_188, i_8_217, i_8_292, i_8_349, i_8_450, i_8_552, i_8_554, i_8_555, i_8_556, i_8_557, i_8_578, i_8_581, i_8_603, i_8_606, i_8_637, i_8_648, i_8_652, i_8_684, i_8_703, i_8_704, i_8_747, i_8_780, i_8_860, i_8_927, i_8_930, i_8_931, i_8_932, i_8_956, i_8_964, i_8_968, i_8_1050, i_8_1109, i_8_1110, i_8_1111, i_8_1112, i_8_1113, i_8_1114, i_8_1115, i_8_1125, i_8_1129, i_8_1256, i_8_1269, i_8_1270, i_8_1271, i_8_1335, i_8_1343, i_8_1388, i_8_1409, i_8_1437, i_8_1457, i_8_1533, i_8_1563, i_8_1564, i_8_1570, i_8_1651, i_8_1676, i_8_1678, i_8_1679, i_8_1682, i_8_1763, i_8_1773, i_8_1774, i_8_1775, i_8_1778, i_8_1819, i_8_1820, i_8_1917, i_8_1918, i_8_1947, i_8_1963, i_8_1964, i_8_1985, i_8_2004, i_8_2016, i_8_2046, i_8_2047, i_8_2049, i_8_2116, i_8_2153, i_8_2169, i_8_2171, i_8_2172, i_8_2173, i_8_2174, i_8_2247, i_8_2261, i_8_2291, o_8_249);
	kernel_8_250 k_8_250(i_8_3, i_8_12, i_8_18, i_8_21, i_8_22, i_8_52, i_8_66, i_8_75, i_8_114, i_8_147, i_8_192, i_8_202, i_8_226, i_8_273, i_8_274, i_8_276, i_8_321, i_8_354, i_8_375, i_8_400, i_8_516, i_8_526, i_8_574, i_8_579, i_8_590, i_8_598, i_8_616, i_8_619, i_8_633, i_8_643, i_8_649, i_8_651, i_8_693, i_8_696, i_8_701, i_8_703, i_8_732, i_8_780, i_8_831, i_8_841, i_8_858, i_8_861, i_8_977, i_8_1200, i_8_1228, i_8_1236, i_8_1237, i_8_1270, i_8_1296, i_8_1302, i_8_1317, i_8_1318, i_8_1323, i_8_1350, i_8_1353, i_8_1356, i_8_1389, i_8_1398, i_8_1408, i_8_1410, i_8_1423, i_8_1436, i_8_1488, i_8_1497, i_8_1505, i_8_1516, i_8_1534, i_8_1551, i_8_1569, i_8_1573, i_8_1639, i_8_1647, i_8_1659, i_8_1677, i_8_1701, i_8_1746, i_8_1753, i_8_1782, i_8_1813, i_8_1824, i_8_1839, i_8_1843, i_8_1866, i_8_1881, i_8_1884, i_8_1911, i_8_1917, i_8_1939, i_8_1944, i_8_1992, i_8_1993, i_8_2008, i_8_2010, i_8_2013, i_8_2046, i_8_2062, i_8_2064, i_8_2184, i_8_2215, i_8_2248, o_8_250);
	kernel_8_251 k_8_251(i_8_28, i_8_67, i_8_72, i_8_140, i_8_143, i_8_201, i_8_258, i_8_259, i_8_275, i_8_385, i_8_392, i_8_401, i_8_429, i_8_457, i_8_492, i_8_498, i_8_499, i_8_522, i_8_550, i_8_556, i_8_630, i_8_632, i_8_655, i_8_659, i_8_662, i_8_672, i_8_673, i_8_695, i_8_820, i_8_843, i_8_854, i_8_859, i_8_880, i_8_881, i_8_916, i_8_959, i_8_995, i_8_1075, i_8_1084, i_8_1087, i_8_1106, i_8_1108, i_8_1109, i_8_1113, i_8_1174, i_8_1201, i_8_1230, i_8_1238, i_8_1267, i_8_1273, i_8_1322, i_8_1330, i_8_1331, i_8_1333, i_8_1411, i_8_1426, i_8_1433, i_8_1471, i_8_1480, i_8_1484, i_8_1498, i_8_1528, i_8_1547, i_8_1561, i_8_1573, i_8_1598, i_8_1641, i_8_1653, i_8_1659, i_8_1705, i_8_1732, i_8_1748, i_8_1750, i_8_1753, i_8_1754, i_8_1762, i_8_1774, i_8_1816, i_8_1849, i_8_1852, i_8_1865, i_8_1867, i_8_1876, i_8_1882, i_8_1889, i_8_1895, i_8_1912, i_8_1921, i_8_1952, i_8_1966, i_8_1975, i_8_2048, i_8_2066, i_8_2092, i_8_2093, i_8_2119, i_8_2150, i_8_2229, i_8_2230, i_8_2299, o_8_251);
	kernel_8_252 k_8_252(i_8_3, i_8_8, i_8_22, i_8_50, i_8_78, i_8_80, i_8_114, i_8_125, i_8_177, i_8_185, i_8_192, i_8_204, i_8_223, i_8_224, i_8_232, i_8_292, i_8_420, i_8_456, i_8_457, i_8_462, i_8_480, i_8_483, i_8_517, i_8_535, i_8_555, i_8_557, i_8_591, i_8_592, i_8_593, i_8_608, i_8_690, i_8_715, i_8_727, i_8_756, i_8_815, i_8_850, i_8_853, i_8_951, i_8_995, i_8_1052, i_8_1142, i_8_1174, i_8_1179, i_8_1180, i_8_1228, i_8_1230, i_8_1237, i_8_1261, i_8_1283, i_8_1308, i_8_1311, i_8_1312, i_8_1314, i_8_1316, i_8_1325, i_8_1329, i_8_1330, i_8_1346, i_8_1364, i_8_1401, i_8_1448, i_8_1462, i_8_1492, i_8_1497, i_8_1504, i_8_1507, i_8_1508, i_8_1555, i_8_1629, i_8_1634, i_8_1647, i_8_1648, i_8_1654, i_8_1670, i_8_1678, i_8_1679, i_8_1682, i_8_1720, i_8_1751, i_8_1753, i_8_1754, i_8_1805, i_8_1812, i_8_1824, i_8_1947, i_8_1948, i_8_1949, i_8_1951, i_8_2005, i_8_2055, i_8_2077, i_8_2158, i_8_2185, i_8_2217, i_8_2235, i_8_2236, i_8_2253, i_8_2275, i_8_2278, i_8_2293, o_8_252);
	kernel_8_253 k_8_253(i_8_23, i_8_33, i_8_75, i_8_76, i_8_77, i_8_85, i_8_114, i_8_139, i_8_193, i_8_231, i_8_322, i_8_364, i_8_424, i_8_428, i_8_429, i_8_507, i_8_509, i_8_510, i_8_526, i_8_527, i_8_589, i_8_604, i_8_606, i_8_655, i_8_660, i_8_678, i_8_703, i_8_808, i_8_823, i_8_832, i_8_838, i_8_878, i_8_896, i_8_969, i_8_992, i_8_1012, i_8_1101, i_8_1155, i_8_1183, i_8_1189, i_8_1191, i_8_1229, i_8_1264, i_8_1266, i_8_1267, i_8_1282, i_8_1299, i_8_1318, i_8_1335, i_8_1336, i_8_1337, i_8_1366, i_8_1393, i_8_1399, i_8_1434, i_8_1437, i_8_1463, i_8_1508, i_8_1517, i_8_1519, i_8_1534, i_8_1543, i_8_1550, i_8_1625, i_8_1642, i_8_1686, i_8_1687, i_8_1689, i_8_1722, i_8_1723, i_8_1768, i_8_1770, i_8_1773, i_8_1774, i_8_1781, i_8_1782, i_8_1786, i_8_1804, i_8_1819, i_8_1822, i_8_1837, i_8_1848, i_8_1857, i_8_1858, i_8_1861, i_8_1866, i_8_1903, i_8_1938, i_8_1939, i_8_1995, i_8_1996, i_8_2029, i_8_2048, i_8_2118, i_8_2134, i_8_2149, i_8_2226, i_8_2245, i_8_2246, i_8_2247, o_8_253);
	kernel_8_254 k_8_254(i_8_22, i_8_88, i_8_141, i_8_203, i_8_206, i_8_229, i_8_240, i_8_257, i_8_265, i_8_310, i_8_328, i_8_337, i_8_345, i_8_355, i_8_373, i_8_382, i_8_426, i_8_427, i_8_430, i_8_455, i_8_457, i_8_490, i_8_505, i_8_524, i_8_554, i_8_556, i_8_565, i_8_569, i_8_604, i_8_626, i_8_627, i_8_676, i_8_710, i_8_752, i_8_761, i_8_770, i_8_778, i_8_836, i_8_938, i_8_951, i_8_1039, i_8_1088, i_8_1108, i_8_1112, i_8_1114, i_8_1115, i_8_1147, i_8_1264, i_8_1306, i_8_1329, i_8_1366, i_8_1369, i_8_1404, i_8_1407, i_8_1414, i_8_1433, i_8_1462, i_8_1480, i_8_1481, i_8_1490, i_8_1493, i_8_1543, i_8_1546, i_8_1552, i_8_1553, i_8_1562, i_8_1582, i_8_1651, i_8_1654, i_8_1677, i_8_1681, i_8_1706, i_8_1717, i_8_1723, i_8_1732, i_8_1733, i_8_1774, i_8_1778, i_8_1805, i_8_1814, i_8_1820, i_8_1821, i_8_1823, i_8_1826, i_8_1883, i_8_1888, i_8_1894, i_8_1903, i_8_1915, i_8_1957, i_8_1964, i_8_1984, i_8_1993, i_8_2105, i_8_2127, i_8_2150, i_8_2224, i_8_2266, i_8_2268, i_8_2290, o_8_254);
	kernel_8_255 k_8_255(i_8_54, i_8_63, i_8_84, i_8_145, i_8_191, i_8_255, i_8_285, i_8_303, i_8_318, i_8_383, i_8_385, i_8_386, i_8_420, i_8_423, i_8_438, i_8_445, i_8_450, i_8_453, i_8_499, i_8_507, i_8_508, i_8_523, i_8_529, i_8_537, i_8_564, i_8_628, i_8_633, i_8_637, i_8_648, i_8_664, i_8_696, i_8_709, i_8_760, i_8_763, i_8_768, i_8_777, i_8_782, i_8_865, i_8_894, i_8_895, i_8_933, i_8_969, i_8_975, i_8_996, i_8_1095, i_8_1098, i_8_1108, i_8_1110, i_8_1111, i_8_1113, i_8_1119, i_8_1237, i_8_1264, i_8_1269, i_8_1314, i_8_1317, i_8_1324, i_8_1365, i_8_1401, i_8_1450, i_8_1506, i_8_1512, i_8_1515, i_8_1533, i_8_1561, i_8_1629, i_8_1635, i_8_1636, i_8_1670, i_8_1677, i_8_1678, i_8_1680, i_8_1681, i_8_1683, i_8_1686, i_8_1701, i_8_1704, i_8_1746, i_8_1753, i_8_1773, i_8_1780, i_8_1790, i_8_1791, i_8_1804, i_8_1818, i_8_1819, i_8_1822, i_8_1825, i_8_1845, i_8_1858, i_8_1867, i_8_1881, i_8_1885, i_8_1917, i_8_2044, i_8_2125, i_8_2142, i_8_2145, i_8_2232, i_8_2233, o_8_255);
	kernel_8_256 k_8_256(i_8_22, i_8_37, i_8_40, i_8_49, i_8_94, i_8_124, i_8_157, i_8_165, i_8_166, i_8_213, i_8_256, i_8_287, i_8_292, i_8_328, i_8_337, i_8_361, i_8_363, i_8_427, i_8_453, i_8_492, i_8_571, i_8_583, i_8_599, i_8_627, i_8_682, i_8_703, i_8_706, i_8_744, i_8_759, i_8_772, i_8_773, i_8_787, i_8_805, i_8_823, i_8_842, i_8_876, i_8_880, i_8_955, i_8_967, i_8_979, i_8_1002, i_8_1040, i_8_1057, i_8_1066, i_8_1110, i_8_1111, i_8_1185, i_8_1227, i_8_1228, i_8_1229, i_8_1231, i_8_1249, i_8_1255, i_8_1257, i_8_1267, i_8_1279, i_8_1305, i_8_1327, i_8_1351, i_8_1357, i_8_1372, i_8_1375, i_8_1380, i_8_1381, i_8_1438, i_8_1447, i_8_1453, i_8_1455, i_8_1456, i_8_1467, i_8_1471, i_8_1578, i_8_1606, i_8_1614, i_8_1639, i_8_1651, i_8_1671, i_8_1696, i_8_1699, i_8_1701, i_8_1733, i_8_1749, i_8_1768, i_8_1821, i_8_1857, i_8_1939, i_8_1981, i_8_1992, i_8_2040, i_8_2055, i_8_2074, i_8_2164, i_8_2185, i_8_2200, i_8_2227, i_8_2238, i_8_2239, i_8_2259, i_8_2263, i_8_2284, o_8_256);
	kernel_8_257 k_8_257(i_8_37, i_8_82, i_8_165, i_8_210, i_8_262, i_8_265, i_8_279, i_8_307, i_8_336, i_8_358, i_8_384, i_8_393, i_8_394, i_8_421, i_8_456, i_8_489, i_8_492, i_8_498, i_8_527, i_8_549, i_8_591, i_8_622, i_8_625, i_8_636, i_8_637, i_8_642, i_8_658, i_8_660, i_8_663, i_8_673, i_8_688, i_8_696, i_8_699, i_8_701, i_8_729, i_8_747, i_8_751, i_8_837, i_8_843, i_8_874, i_8_882, i_8_921, i_8_930, i_8_973, i_8_983, i_8_1009, i_8_1050, i_8_1056, i_8_1071, i_8_1075, i_8_1084, i_8_1129, i_8_1182, i_8_1228, i_8_1234, i_8_1263, i_8_1278, i_8_1291, i_8_1296, i_8_1306, i_8_1357, i_8_1362, i_8_1383, i_8_1390, i_8_1399, i_8_1410, i_8_1411, i_8_1435, i_8_1440, i_8_1441, i_8_1479, i_8_1507, i_8_1548, i_8_1551, i_8_1565, i_8_1608, i_8_1681, i_8_1683, i_8_1687, i_8_1720, i_8_1729, i_8_1731, i_8_1746, i_8_1747, i_8_1752, i_8_1768, i_8_1824, i_8_1855, i_8_1884, i_8_1887, i_8_1980, i_8_1989, i_8_2019, i_8_2052, i_8_2070, i_8_2118, i_8_2142, i_8_2148, i_8_2226, i_8_2286, o_8_257);
	kernel_8_258 k_8_258(i_8_1, i_8_22, i_8_57, i_8_85, i_8_96, i_8_103, i_8_104, i_8_105, i_8_165, i_8_168, i_8_202, i_8_210, i_8_211, i_8_214, i_8_219, i_8_220, i_8_223, i_8_256, i_8_292, i_8_333, i_8_345, i_8_361, i_8_415, i_8_445, i_8_448, i_8_475, i_8_501, i_8_589, i_8_596, i_8_606, i_8_627, i_8_658, i_8_669, i_8_670, i_8_716, i_8_768, i_8_786, i_8_888, i_8_949, i_8_977, i_8_984, i_8_985, i_8_991, i_8_992, i_8_1084, i_8_1110, i_8_1113, i_8_1155, i_8_1216, i_8_1222, i_8_1232, i_8_1248, i_8_1267, i_8_1272, i_8_1344, i_8_1347, i_8_1402, i_8_1419, i_8_1420, i_8_1423, i_8_1428, i_8_1437, i_8_1467, i_8_1477, i_8_1489, i_8_1518, i_8_1524, i_8_1544, i_8_1555, i_8_1588, i_8_1615, i_8_1618, i_8_1636, i_8_1677, i_8_1678, i_8_1680, i_8_1704, i_8_1720, i_8_1749, i_8_1780, i_8_1783, i_8_1785, i_8_1786, i_8_1825, i_8_1855, i_8_1861, i_8_1902, i_8_1963, i_8_2009, i_8_2026, i_8_2126, i_8_2128, i_8_2139, i_8_2140, i_8_2143, i_8_2150, i_8_2152, i_8_2236, i_8_2293, i_8_2294, o_8_258);
	kernel_8_259 k_8_259(i_8_41, i_8_83, i_8_104, i_8_115, i_8_166, i_8_247, i_8_266, i_8_283, i_8_302, i_8_304, i_8_326, i_8_362, i_8_364, i_8_383, i_8_419, i_8_427, i_8_437, i_8_440, i_8_451, i_8_457, i_8_490, i_8_500, i_8_505, i_8_527, i_8_545, i_8_548, i_8_572, i_8_594, i_8_598, i_8_599, i_8_635, i_8_643, i_8_658, i_8_662, i_8_695, i_8_698, i_8_699, i_8_700, i_8_716, i_8_781, i_8_782, i_8_787, i_8_789, i_8_808, i_8_812, i_8_815, i_8_824, i_8_841, i_8_853, i_8_877, i_8_974, i_8_992, i_8_1061, i_8_1067, i_8_1211, i_8_1224, i_8_1228, i_8_1236, i_8_1253, i_8_1273, i_8_1296, i_8_1358, i_8_1365, i_8_1399, i_8_1426, i_8_1444, i_8_1471, i_8_1552, i_8_1589, i_8_1637, i_8_1697, i_8_1700, i_8_1705, i_8_1747, i_8_1768, i_8_1781, i_8_1783, i_8_1787, i_8_1805, i_8_1807, i_8_1851, i_8_1854, i_8_1855, i_8_1858, i_8_1859, i_8_1886, i_8_1949, i_8_1984, i_8_1993, i_8_1995, i_8_2029, i_8_2032, i_8_2090, i_8_2117, i_8_2134, i_8_2137, i_8_2155, i_8_2162, i_8_2191, i_8_2244, o_8_259);
	kernel_8_260 k_8_260(i_8_6, i_8_14, i_8_44, i_8_106, i_8_140, i_8_196, i_8_197, i_8_214, i_8_222, i_8_228, i_8_241, i_8_311, i_8_322, i_8_323, i_8_328, i_8_364, i_8_367, i_8_368, i_8_436, i_8_439, i_8_574, i_8_606, i_8_628, i_8_633, i_8_646, i_8_665, i_8_672, i_8_674, i_8_682, i_8_701, i_8_707, i_8_709, i_8_710, i_8_735, i_8_804, i_8_823, i_8_834, i_8_886, i_8_957, i_8_979, i_8_985, i_8_1060, i_8_1074, i_8_1105, i_8_1132, i_8_1158, i_8_1185, i_8_1236, i_8_1239, i_8_1266, i_8_1284, i_8_1310, i_8_1352, i_8_1353, i_8_1354, i_8_1357, i_8_1365, i_8_1374, i_8_1375, i_8_1384, i_8_1405, i_8_1426, i_8_1429, i_8_1480, i_8_1590, i_8_1623, i_8_1624, i_8_1636, i_8_1649, i_8_1671, i_8_1672, i_8_1731, i_8_1749, i_8_1752, i_8_1770, i_8_1797, i_8_1824, i_8_1825, i_8_1903, i_8_1905, i_8_1914, i_8_1942, i_8_2031, i_8_2056, i_8_2082, i_8_2128, i_8_2136, i_8_2148, i_8_2193, i_8_2194, i_8_2217, i_8_2230, i_8_2263, i_8_2269, i_8_2272, i_8_2273, i_8_2274, i_8_2275, i_8_2276, i_8_2290, o_8_260);
	kernel_8_261 k_8_261(i_8_14, i_8_50, i_8_55, i_8_58, i_8_141, i_8_143, i_8_157, i_8_159, i_8_187, i_8_259, i_8_310, i_8_373, i_8_378, i_8_429, i_8_437, i_8_442, i_8_445, i_8_474, i_8_481, i_8_526, i_8_582, i_8_596, i_8_601, i_8_607, i_8_627, i_8_691, i_8_693, i_8_710, i_8_714, i_8_717, i_8_760, i_8_778, i_8_818, i_8_884, i_8_913, i_8_941, i_8_956, i_8_1012, i_8_1048, i_8_1050, i_8_1056, i_8_1071, i_8_1088, i_8_1090, i_8_1116, i_8_1123, i_8_1133, i_8_1189, i_8_1241, i_8_1264, i_8_1267, i_8_1273, i_8_1276, i_8_1287, i_8_1295, i_8_1324, i_8_1326, i_8_1327, i_8_1335, i_8_1390, i_8_1435, i_8_1467, i_8_1472, i_8_1507, i_8_1545, i_8_1588, i_8_1599, i_8_1605, i_8_1629, i_8_1632, i_8_1653, i_8_1668, i_8_1719, i_8_1723, i_8_1746, i_8_1772, i_8_1784, i_8_1790, i_8_1797, i_8_1830, i_8_1831, i_8_1839, i_8_1877, i_8_1900, i_8_1917, i_8_1918, i_8_1919, i_8_1930, i_8_1939, i_8_1989, i_8_2028, i_8_2101, i_8_2112, i_8_2133, i_8_2185, i_8_2211, i_8_2241, i_8_2245, i_8_2270, i_8_2293, o_8_261);
	kernel_8_262 k_8_262(i_8_31, i_8_49, i_8_54, i_8_56, i_8_81, i_8_85, i_8_86, i_8_103, i_8_219, i_8_229, i_8_237, i_8_297, i_8_300, i_8_301, i_8_346, i_8_361, i_8_362, i_8_366, i_8_442, i_8_486, i_8_522, i_8_523, i_8_524, i_8_580, i_8_585, i_8_586, i_8_590, i_8_603, i_8_622, i_8_630, i_8_657, i_8_662, i_8_667, i_8_675, i_8_676, i_8_677, i_8_833, i_8_839, i_8_850, i_8_876, i_8_877, i_8_1048, i_8_1071, i_8_1072, i_8_1108, i_8_1189, i_8_1190, i_8_1225, i_8_1263, i_8_1264, i_8_1270, i_8_1271, i_8_1282, i_8_1283, i_8_1286, i_8_1296, i_8_1333, i_8_1334, i_8_1337, i_8_1353, i_8_1408, i_8_1409, i_8_1534, i_8_1550, i_8_1561, i_8_1620, i_8_1629, i_8_1631, i_8_1638, i_8_1648, i_8_1680, i_8_1728, i_8_1732, i_8_1768, i_8_1773, i_8_1774, i_8_1782, i_8_1784, i_8_1811, i_8_1818, i_8_1819, i_8_1830, i_8_1848, i_8_1855, i_8_1856, i_8_1888, i_8_1903, i_8_1904, i_8_1962, i_8_1982, i_8_1985, i_8_2037, i_8_2038, i_8_2133, i_8_2134, i_8_2147, i_8_2155, i_8_2245, i_8_2270, i_8_2293, o_8_262);
	kernel_8_263 k_8_263(i_8_20, i_8_36, i_8_135, i_8_253, i_8_280, i_8_297, i_8_364, i_8_396, i_8_432, i_8_480, i_8_530, i_8_544, i_8_585, i_8_595, i_8_615, i_8_621, i_8_630, i_8_636, i_8_657, i_8_666, i_8_667, i_8_675, i_8_682, i_8_703, i_8_720, i_8_721, i_8_724, i_8_765, i_8_801, i_8_804, i_8_822, i_8_847, i_8_866, i_8_868, i_8_879, i_8_892, i_8_955, i_8_965, i_8_967, i_8_985, i_8_991, i_8_1050, i_8_1071, i_8_1111, i_8_1188, i_8_1189, i_8_1233, i_8_1251, i_8_1261, i_8_1292, i_8_1300, i_8_1351, i_8_1353, i_8_1359, i_8_1365, i_8_1366, i_8_1367, i_8_1374, i_8_1382, i_8_1450, i_8_1467, i_8_1531, i_8_1536, i_8_1537, i_8_1549, i_8_1559, i_8_1565, i_8_1575, i_8_1584, i_8_1586, i_8_1588, i_8_1622, i_8_1624, i_8_1629, i_8_1639, i_8_1674, i_8_1680, i_8_1681, i_8_1697, i_8_1747, i_8_1750, i_8_1756, i_8_1762, i_8_1815, i_8_1837, i_8_1908, i_8_1944, i_8_1947, i_8_1982, i_8_2004, i_8_2107, i_8_2116, i_8_2125, i_8_2139, i_8_2147, i_8_2187, i_8_2188, i_8_2191, i_8_2255, i_8_2259, o_8_263);
	kernel_8_264 k_8_264(i_8_6, i_8_41, i_8_60, i_8_115, i_8_118, i_8_179, i_8_202, i_8_256, i_8_258, i_8_292, i_8_363, i_8_364, i_8_381, i_8_392, i_8_401, i_8_419, i_8_422, i_8_462, i_8_475, i_8_509, i_8_525, i_8_529, i_8_572, i_8_581, i_8_589, i_8_592, i_8_606, i_8_607, i_8_618, i_8_633, i_8_708, i_8_714, i_8_769, i_8_795, i_8_796, i_8_818, i_8_824, i_8_835, i_8_858, i_8_895, i_8_896, i_8_897, i_8_992, i_8_1040, i_8_1131, i_8_1132, i_8_1192, i_8_1202, i_8_1267, i_8_1278, i_8_1282, i_8_1286, i_8_1319, i_8_1328, i_8_1334, i_8_1382, i_8_1407, i_8_1427, i_8_1443, i_8_1448, i_8_1455, i_8_1481, i_8_1489, i_8_1490, i_8_1508, i_8_1550, i_8_1553, i_8_1578, i_8_1589, i_8_1597, i_8_1614, i_8_1632, i_8_1697, i_8_1705, i_8_1706, i_8_1751, i_8_1760, i_8_1762, i_8_1807, i_8_1808, i_8_1837, i_8_1841, i_8_1885, i_8_1888, i_8_1963, i_8_1994, i_8_2002, i_8_2011, i_8_2090, i_8_2111, i_8_2113, i_8_2127, i_8_2176, i_8_2177, i_8_2184, i_8_2188, i_8_2211, i_8_2262, i_8_2273, i_8_2291, o_8_264);
	kernel_8_265 k_8_265(i_8_1, i_8_2, i_8_19, i_8_31, i_8_60, i_8_115, i_8_116, i_8_198, i_8_266, i_8_269, i_8_284, i_8_293, i_8_346, i_8_349, i_8_366, i_8_378, i_8_380, i_8_385, i_8_427, i_8_437, i_8_445, i_8_446, i_8_463, i_8_464, i_8_488, i_8_492, i_8_556, i_8_572, i_8_586, i_8_590, i_8_599, i_8_614, i_8_649, i_8_658, i_8_660, i_8_665, i_8_673, i_8_674, i_8_716, i_8_718, i_8_725, i_8_735, i_8_782, i_8_796, i_8_827, i_8_841, i_8_956, i_8_976, i_8_997, i_8_998, i_8_1004, i_8_1007, i_8_1039, i_8_1058, i_8_1074, i_8_1114, i_8_1130, i_8_1211, i_8_1237, i_8_1259, i_8_1274, i_8_1281, i_8_1302, i_8_1355, i_8_1437, i_8_1525, i_8_1542, i_8_1543, i_8_1544, i_8_1546, i_8_1547, i_8_1589, i_8_1592, i_8_1598, i_8_1618, i_8_1634, i_8_1655, i_8_1669, i_8_1677, i_8_1699, i_8_1714, i_8_1723, i_8_1724, i_8_1730, i_8_1753, i_8_1780, i_8_1919, i_8_1922, i_8_1967, i_8_1970, i_8_2114, i_8_2120, i_8_2129, i_8_2149, i_8_2192, i_8_2195, i_8_2242, i_8_2263, i_8_2275, i_8_2294, o_8_265);
	kernel_8_266 k_8_266(i_8_39, i_8_40, i_8_49, i_8_82, i_8_90, i_8_120, i_8_192, i_8_300, i_8_318, i_8_321, i_8_322, i_8_391, i_8_399, i_8_415, i_8_418, i_8_428, i_8_453, i_8_507, i_8_532, i_8_552, i_8_571, i_8_572, i_8_574, i_8_595, i_8_606, i_8_639, i_8_651, i_8_657, i_8_660, i_8_678, i_8_706, i_8_829, i_8_831, i_8_840, i_8_925, i_8_964, i_8_967, i_8_969, i_8_972, i_8_975, i_8_984, i_8_993, i_8_1011, i_8_1039, i_8_1101, i_8_1104, i_8_1105, i_8_1111, i_8_1228, i_8_1239, i_8_1245, i_8_1257, i_8_1266, i_8_1397, i_8_1407, i_8_1435, i_8_1440, i_8_1452, i_8_1456, i_8_1461, i_8_1462, i_8_1464, i_8_1470, i_8_1474, i_8_1476, i_8_1479, i_8_1480, i_8_1488, i_8_1549, i_8_1551, i_8_1552, i_8_1624, i_8_1659, i_8_1704, i_8_1705, i_8_1719, i_8_1724, i_8_1731, i_8_1749, i_8_1767, i_8_1775, i_8_1779, i_8_1794, i_8_1795, i_8_1801, i_8_1820, i_8_1836, i_8_1839, i_8_1858, i_8_1859, i_8_1885, i_8_1911, i_8_1948, i_8_1956, i_8_2075, i_8_2173, i_8_2190, i_8_2226, i_8_2258, i_8_2278, o_8_266);
	kernel_8_267 k_8_267(i_8_50, i_8_52, i_8_58, i_8_59, i_8_71, i_8_89, i_8_97, i_8_118, i_8_142, i_8_157, i_8_160, i_8_204, i_8_205, i_8_210, i_8_212, i_8_214, i_8_223, i_8_241, i_8_244, i_8_258, i_8_346, i_8_373, i_8_419, i_8_440, i_8_476, i_8_498, i_8_499, i_8_500, i_8_502, i_8_522, i_8_588, i_8_589, i_8_605, i_8_662, i_8_715, i_8_730, i_8_765, i_8_781, i_8_784, i_8_877, i_8_904, i_8_907, i_8_925, i_8_975, i_8_986, i_8_1027, i_8_1074, i_8_1110, i_8_1186, i_8_1249, i_8_1250, i_8_1255, i_8_1281, i_8_1284, i_8_1341, i_8_1342, i_8_1420, i_8_1426, i_8_1435, i_8_1443, i_8_1470, i_8_1472, i_8_1492, i_8_1528, i_8_1541, i_8_1555, i_8_1588, i_8_1589, i_8_1596, i_8_1597, i_8_1598, i_8_1634, i_8_1647, i_8_1678, i_8_1699, i_8_1706, i_8_1711, i_8_1737, i_8_1753, i_8_1782, i_8_1796, i_8_1818, i_8_1819, i_8_1834, i_8_1844, i_8_1855, i_8_1867, i_8_1870, i_8_1903, i_8_1975, i_8_2046, i_8_2109, i_8_2110, i_8_2111, i_8_2143, i_8_2183, i_8_2190, i_8_2224, i_8_2244, i_8_2272, o_8_267);
	kernel_8_268 k_8_268(i_8_9, i_8_72, i_8_108, i_8_111, i_8_135, i_8_162, i_8_183, i_8_228, i_8_234, i_8_262, i_8_361, i_8_363, i_8_396, i_8_477, i_8_479, i_8_480, i_8_481, i_8_498, i_8_522, i_8_543, i_8_549, i_8_567, i_8_568, i_8_570, i_8_571, i_8_603, i_8_633, i_8_636, i_8_652, i_8_675, i_8_676, i_8_677, i_8_684, i_8_748, i_8_759, i_8_793, i_8_855, i_8_936, i_8_966, i_8_999, i_8_1010, i_8_1036, i_8_1183, i_8_1188, i_8_1228, i_8_1236, i_8_1263, i_8_1272, i_8_1296, i_8_1315, i_8_1323, i_8_1332, i_8_1434, i_8_1459, i_8_1476, i_8_1485, i_8_1486, i_8_1512, i_8_1521, i_8_1522, i_8_1553, i_8_1585, i_8_1596, i_8_1647, i_8_1650, i_8_1683, i_8_1696, i_8_1704, i_8_1719, i_8_1728, i_8_1737, i_8_1752, i_8_1755, i_8_1773, i_8_1774, i_8_1776, i_8_1804, i_8_1818, i_8_1827, i_8_1836, i_8_1837, i_8_1838, i_8_1839, i_8_1840, i_8_1846, i_8_1854, i_8_1881, i_8_1993, i_8_2070, i_8_2118, i_8_2133, i_8_2145, i_8_2146, i_8_2188, i_8_2214, i_8_2223, i_8_2241, i_8_2242, i_8_2262, i_8_2295, o_8_268);
	kernel_8_269 k_8_269(i_8_1, i_8_24, i_8_28, i_8_62, i_8_64, i_8_155, i_8_163, i_8_166, i_8_189, i_8_193, i_8_217, i_8_218, i_8_220, i_8_234, i_8_240, i_8_256, i_8_293, i_8_296, i_8_304, i_8_334, i_8_338, i_8_360, i_8_361, i_8_385, i_8_386, i_8_425, i_8_490, i_8_593, i_8_602, i_8_619, i_8_620, i_8_631, i_8_658, i_8_693, i_8_704, i_8_707, i_8_709, i_8_731, i_8_757, i_8_777, i_8_789, i_8_812, i_8_843, i_8_848, i_8_854, i_8_881, i_8_1123, i_8_1127, i_8_1154, i_8_1157, i_8_1179, i_8_1180, i_8_1181, i_8_1261, i_8_1271, i_8_1274, i_8_1277, i_8_1293, i_8_1302, i_8_1330, i_8_1341, i_8_1388, i_8_1391, i_8_1408, i_8_1410, i_8_1473, i_8_1474, i_8_1538, i_8_1545, i_8_1546, i_8_1548, i_8_1549, i_8_1586, i_8_1601, i_8_1604, i_8_1629, i_8_1654, i_8_1678, i_8_1720, i_8_1735, i_8_1776, i_8_1800, i_8_1818, i_8_1819, i_8_1846, i_8_1860, i_8_1887, i_8_2005, i_8_2051, i_8_2077, i_8_2116, i_8_2117, i_8_2150, i_8_2154, i_8_2155, i_8_2230, i_8_2269, i_8_2291, i_8_2295, i_8_2297, o_8_269);
	kernel_8_270 k_8_270(i_8_35, i_8_169, i_8_339, i_8_447, i_8_453, i_8_456, i_8_483, i_8_492, i_8_502, i_8_510, i_8_527, i_8_574, i_8_627, i_8_655, i_8_696, i_8_699, i_8_705, i_8_708, i_8_762, i_8_780, i_8_808, i_8_834, i_8_840, i_8_843, i_8_886, i_8_941, i_8_943, i_8_946, i_8_947, i_8_958, i_8_967, i_8_969, i_8_987, i_8_993, i_8_996, i_8_1032, i_8_1050, i_8_1060, i_8_1069, i_8_1093, i_8_1129, i_8_1168, i_8_1185, i_8_1186, i_8_1187, i_8_1232, i_8_1258, i_8_1285, i_8_1286, i_8_1306, i_8_1307, i_8_1310, i_8_1312, i_8_1336, i_8_1402, i_8_1410, i_8_1411, i_8_1438, i_8_1474, i_8_1490, i_8_1492, i_8_1510, i_8_1537, i_8_1538, i_8_1545, i_8_1554, i_8_1591, i_8_1624, i_8_1654, i_8_1655, i_8_1671, i_8_1725, i_8_1732, i_8_1734, i_8_1741, i_8_1744, i_8_1745, i_8_1762, i_8_1770, i_8_1788, i_8_1888, i_8_1896, i_8_1906, i_8_1984, i_8_2041, i_8_2058, i_8_2059, i_8_2073, i_8_2076, i_8_2092, i_8_2094, i_8_2095, i_8_2122, i_8_2132, i_8_2146, i_8_2218, i_8_2230, i_8_2236, i_8_2247, i_8_2302, o_8_270);
	kernel_8_271 k_8_271(i_8_50, i_8_112, i_8_114, i_8_218, i_8_253, i_8_255, i_8_301, i_8_316, i_8_343, i_8_361, i_8_418, i_8_426, i_8_427, i_8_453, i_8_454, i_8_455, i_8_505, i_8_532, i_8_586, i_8_595, i_8_639, i_8_648, i_8_650, i_8_651, i_8_657, i_8_661, i_8_675, i_8_676, i_8_677, i_8_706, i_8_713, i_8_820, i_8_849, i_8_850, i_8_875, i_8_886, i_8_892, i_8_991, i_8_992, i_8_1035, i_8_1054, i_8_1055, i_8_1102, i_8_1127, i_8_1217, i_8_1226, i_8_1234, i_8_1264, i_8_1270, i_8_1325, i_8_1327, i_8_1336, i_8_1424, i_8_1439, i_8_1452, i_8_1459, i_8_1462, i_8_1486, i_8_1487, i_8_1522, i_8_1524, i_8_1549, i_8_1603, i_8_1611, i_8_1612, i_8_1615, i_8_1629, i_8_1676, i_8_1680, i_8_1682, i_8_1693, i_8_1705, i_8_1747, i_8_1749, i_8_1769, i_8_1791, i_8_1810, i_8_1811, i_8_1825, i_8_1837, i_8_1881, i_8_1945, i_8_1946, i_8_1954, i_8_1957, i_8_1963, i_8_1966, i_8_1972, i_8_1981, i_8_1984, i_8_1990, i_8_2029, i_8_2054, i_8_2126, i_8_2223, i_8_2244, i_8_2245, i_8_2246, i_8_2260, i_8_2263, o_8_271);
	kernel_8_272 k_8_272(i_8_25, i_8_70, i_8_94, i_8_96, i_8_185, i_8_215, i_8_229, i_8_301, i_8_328, i_8_329, i_8_345, i_8_373, i_8_374, i_8_379, i_8_383, i_8_423, i_8_462, i_8_592, i_8_593, i_8_606, i_8_608, i_8_612, i_8_621, i_8_622, i_8_623, i_8_625, i_8_626, i_8_638, i_8_702, i_8_703, i_8_704, i_8_705, i_8_713, i_8_720, i_8_723, i_8_778, i_8_779, i_8_854, i_8_934, i_8_973, i_8_984, i_8_985, i_8_986, i_8_987, i_8_988, i_8_989, i_8_996, i_8_997, i_8_1027, i_8_1123, i_8_1191, i_8_1272, i_8_1273, i_8_1297, i_8_1305, i_8_1307, i_8_1330, i_8_1402, i_8_1410, i_8_1470, i_8_1471, i_8_1473, i_8_1483, i_8_1526, i_8_1529, i_8_1621, i_8_1623, i_8_1625, i_8_1626, i_8_1651, i_8_1661, i_8_1731, i_8_1733, i_8_1734, i_8_1735, i_8_1736, i_8_1752, i_8_1776, i_8_1789, i_8_1790, i_8_1818, i_8_1841, i_8_1857, i_8_1860, i_8_1862, i_8_1902, i_8_1950, i_8_1965, i_8_1967, i_8_1980, i_8_2015, i_8_2025, i_8_2026, i_8_2058, i_8_2070, i_8_2076, i_8_2154, i_8_2156, i_8_2169, i_8_2237, o_8_272);
	kernel_8_273 k_8_273(i_8_4, i_8_23, i_8_64, i_8_75, i_8_85, i_8_131, i_8_176, i_8_193, i_8_233, i_8_235, i_8_247, i_8_248, i_8_301, i_8_302, i_8_310, i_8_362, i_8_374, i_8_426, i_8_428, i_8_489, i_8_493, i_8_497, i_8_536, i_8_581, i_8_596, i_8_651, i_8_655, i_8_671, i_8_703, i_8_706, i_8_803, i_8_832, i_8_860, i_8_911, i_8_914, i_8_956, i_8_967, i_8_991, i_8_1030, i_8_1048, i_8_1085, i_8_1095, i_8_1112, i_8_1132, i_8_1135, i_8_1164, i_8_1190, i_8_1228, i_8_1271, i_8_1308, i_8_1324, i_8_1355, i_8_1397, i_8_1400, i_8_1405, i_8_1407, i_8_1408, i_8_1428, i_8_1468, i_8_1492, i_8_1493, i_8_1498, i_8_1532, i_8_1534, i_8_1535, i_8_1549, i_8_1632, i_8_1636, i_8_1642, i_8_1688, i_8_1781, i_8_1795, i_8_1804, i_8_1805, i_8_1807, i_8_1819, i_8_1821, i_8_1855, i_8_1868, i_8_1885, i_8_1905, i_8_1913, i_8_1919, i_8_1949, i_8_1992, i_8_1994, i_8_1996, i_8_2011, i_8_2047, i_8_2048, i_8_2063, i_8_2066, i_8_2119, i_8_2144, i_8_2145, i_8_2147, i_8_2149, i_8_2216, i_8_2234, i_8_2275, o_8_273);
	kernel_8_274 k_8_274(i_8_27, i_8_28, i_8_217, i_8_254, i_8_257, i_8_299, i_8_305, i_8_316, i_8_323, i_8_368, i_8_381, i_8_428, i_8_454, i_8_470, i_8_488, i_8_572, i_8_587, i_8_595, i_8_610, i_8_631, i_8_632, i_8_649, i_8_678, i_8_695, i_8_697, i_8_778, i_8_779, i_8_796, i_8_833, i_8_839, i_8_844, i_8_847, i_8_848, i_8_856, i_8_860, i_8_868, i_8_874, i_8_875, i_8_877, i_8_878, i_8_883, i_8_965, i_8_969, i_8_1136, i_8_1216, i_8_1226, i_8_1228, i_8_1255, i_8_1262, i_8_1281, i_8_1285, i_8_1298, i_8_1355, i_8_1410, i_8_1442, i_8_1449, i_8_1514, i_8_1516, i_8_1526, i_8_1543, i_8_1544, i_8_1547, i_8_1559, i_8_1561, i_8_1607, i_8_1615, i_8_1621, i_8_1630, i_8_1631, i_8_1634, i_8_1675, i_8_1703, i_8_1704, i_8_1714, i_8_1720, i_8_1756, i_8_1757, i_8_1759, i_8_1776, i_8_1810, i_8_1882, i_8_1972, i_8_1982, i_8_1990, i_8_1994, i_8_2054, i_8_2099, i_8_2102, i_8_2134, i_8_2136, i_8_2140, i_8_2156, i_8_2170, i_8_2225, i_8_2242, i_8_2243, i_8_2263, i_8_2264, i_8_2270, i_8_2291, o_8_274);
	kernel_8_275 k_8_275(i_8_20, i_8_38, i_8_47, i_8_50, i_8_55, i_8_56, i_8_65, i_8_92, i_8_115, i_8_173, i_8_189, i_8_236, i_8_299, i_8_304, i_8_308, i_8_335, i_8_352, i_8_362, i_8_379, i_8_380, i_8_387, i_8_418, i_8_425, i_8_452, i_8_524, i_8_530, i_8_578, i_8_586, i_8_587, i_8_658, i_8_666, i_8_704, i_8_779, i_8_793, i_8_801, i_8_803, i_8_829, i_8_848, i_8_880, i_8_883, i_8_884, i_8_919, i_8_927, i_8_928, i_8_992, i_8_994, i_8_1033, i_8_1054, i_8_1079, i_8_1091, i_8_1129, i_8_1145, i_8_1163, i_8_1226, i_8_1271, i_8_1283, i_8_1289, i_8_1297, i_8_1328, i_8_1333, i_8_1405, i_8_1406, i_8_1459, i_8_1505, i_8_1559, i_8_1603, i_8_1604, i_8_1747, i_8_1817, i_8_1823, i_8_1862, i_8_1864, i_8_1865, i_8_1883, i_8_1884, i_8_1886, i_8_1907, i_8_1918, i_8_1937, i_8_1992, i_8_1993, i_8_2008, i_8_2026, i_8_2030, i_8_2045, i_8_2052, i_8_2054, i_8_2096, i_8_2107, i_8_2132, i_8_2144, i_8_2152, i_8_2153, i_8_2180, i_8_2196, i_8_2197, i_8_2206, i_8_2210, i_8_2227, i_8_2287, o_8_275);
	kernel_8_276 k_8_276(i_8_14, i_8_26, i_8_27, i_8_54, i_8_57, i_8_87, i_8_168, i_8_169, i_8_189, i_8_228, i_8_259, i_8_300, i_8_338, i_8_344, i_8_346, i_8_360, i_8_383, i_8_403, i_8_427, i_8_428, i_8_455, i_8_555, i_8_574, i_8_635, i_8_659, i_8_694, i_8_700, i_8_705, i_8_706, i_8_708, i_8_762, i_8_791, i_8_798, i_8_799, i_8_874, i_8_920, i_8_929, i_8_997, i_8_998, i_8_1077, i_8_1103, i_8_1105, i_8_1192, i_8_1195, i_8_1239, i_8_1260, i_8_1265, i_8_1276, i_8_1283, i_8_1288, i_8_1289, i_8_1299, i_8_1308, i_8_1309, i_8_1318, i_8_1321, i_8_1348, i_8_1382, i_8_1385, i_8_1393, i_8_1410, i_8_1436, i_8_1451, i_8_1470, i_8_1549, i_8_1590, i_8_1591, i_8_1592, i_8_1623, i_8_1625, i_8_1639, i_8_1642, i_8_1649, i_8_1690, i_8_1743, i_8_1762, i_8_1823, i_8_1826, i_8_1885, i_8_1888, i_8_1940, i_8_1986, i_8_1993, i_8_2040, i_8_2055, i_8_2056, i_8_2059, i_8_2077, i_8_2132, i_8_2147, i_8_2177, i_8_2200, i_8_2210, i_8_2213, i_8_2217, i_8_2219, i_8_2239, i_8_2240, i_8_2301, i_8_2302, o_8_276);
	kernel_8_277 k_8_277(i_8_13, i_8_74, i_8_79, i_8_103, i_8_114, i_8_115, i_8_116, i_8_137, i_8_184, i_8_190, i_8_196, i_8_233, i_8_284, i_8_301, i_8_319, i_8_320, i_8_326, i_8_343, i_8_366, i_8_427, i_8_434, i_8_450, i_8_493, i_8_525, i_8_526, i_8_544, i_8_640, i_8_660, i_8_665, i_8_703, i_8_748, i_8_782, i_8_799, i_8_800, i_8_854, i_8_880, i_8_946, i_8_965, i_8_971, i_8_977, i_8_992, i_8_1051, i_8_1061, i_8_1110, i_8_1114, i_8_1228, i_8_1236, i_8_1246, i_8_1263, i_8_1294, i_8_1295, i_8_1316, i_8_1325, i_8_1328, i_8_1354, i_8_1363, i_8_1364, i_8_1417, i_8_1424, i_8_1432, i_8_1441, i_8_1462, i_8_1463, i_8_1468, i_8_1517, i_8_1522, i_8_1538, i_8_1552, i_8_1561, i_8_1614, i_8_1624, i_8_1651, i_8_1678, i_8_1694, i_8_1702, i_8_1730, i_8_1746, i_8_1747, i_8_1819, i_8_1855, i_8_1859, i_8_1913, i_8_1930, i_8_1939, i_8_1964, i_8_1982, i_8_1995, i_8_2008, i_8_2047, i_8_2074, i_8_2143, i_8_2149, i_8_2153, i_8_2156, i_8_2161, i_8_2170, i_8_2225, i_8_2245, i_8_2247, i_8_2249, o_8_277);
	kernel_8_278 k_8_278(i_8_19, i_8_25, i_8_35, i_8_48, i_8_93, i_8_139, i_8_141, i_8_142, i_8_246, i_8_310, i_8_349, i_8_453, i_8_455, i_8_481, i_8_485, i_8_491, i_8_522, i_8_525, i_8_526, i_8_527, i_8_529, i_8_530, i_8_535, i_8_544, i_8_546, i_8_563, i_8_593, i_8_625, i_8_638, i_8_655, i_8_661, i_8_691, i_8_693, i_8_697, i_8_739, i_8_762, i_8_763, i_8_764, i_8_771, i_8_825, i_8_874, i_8_882, i_8_943, i_8_949, i_8_968, i_8_994, i_8_996, i_8_1056, i_8_1059, i_8_1063, i_8_1066, i_8_1067, i_8_1129, i_8_1135, i_8_1138, i_8_1180, i_8_1192, i_8_1219, i_8_1237, i_8_1260, i_8_1268, i_8_1305, i_8_1306, i_8_1307, i_8_1308, i_8_1315, i_8_1322, i_8_1323, i_8_1421, i_8_1431, i_8_1510, i_8_1547, i_8_1564, i_8_1574, i_8_1606, i_8_1651, i_8_1670, i_8_1682, i_8_1696, i_8_1723, i_8_1732, i_8_1751, i_8_1752, i_8_1762, i_8_1795, i_8_1807, i_8_1842, i_8_1848, i_8_1885, i_8_1918, i_8_1947, i_8_1980, i_8_1994, i_8_2014, i_8_2150, i_8_2177, i_8_2183, i_8_2214, i_8_2223, i_8_2263, o_8_278);
	kernel_8_279 k_8_279(i_8_22, i_8_95, i_8_135, i_8_140, i_8_208, i_8_325, i_8_337, i_8_426, i_8_450, i_8_459, i_8_484, i_8_496, i_8_497, i_8_500, i_8_525, i_8_528, i_8_539, i_8_544, i_8_545, i_8_551, i_8_557, i_8_649, i_8_658, i_8_668, i_8_669, i_8_675, i_8_708, i_8_720, i_8_760, i_8_762, i_8_779, i_8_820, i_8_842, i_8_846, i_8_867, i_8_875, i_8_956, i_8_989, i_8_1010, i_8_1028, i_8_1107, i_8_1108, i_8_1109, i_8_1112, i_8_1151, i_8_1180, i_8_1231, i_8_1260, i_8_1263, i_8_1270, i_8_1279, i_8_1304, i_8_1315, i_8_1316, i_8_1324, i_8_1338, i_8_1343, i_8_1432, i_8_1435, i_8_1526, i_8_1534, i_8_1536, i_8_1537, i_8_1549, i_8_1565, i_8_1579, i_8_1585, i_8_1618, i_8_1619, i_8_1630, i_8_1662, i_8_1665, i_8_1679, i_8_1682, i_8_1705, i_8_1732, i_8_1735, i_8_1747, i_8_1754, i_8_1787, i_8_1790, i_8_1805, i_8_1821, i_8_1867, i_8_1887, i_8_1888, i_8_1898, i_8_1920, i_8_2013, i_8_2047, i_8_2073, i_8_2086, i_8_2087, i_8_2105, i_8_2141, i_8_2146, i_8_2216, i_8_2266, i_8_2288, i_8_2302, o_8_279);
	kernel_8_280 k_8_280(i_8_23, i_8_77, i_8_85, i_8_119, i_8_137, i_8_163, i_8_244, i_8_247, i_8_266, i_8_274, i_8_311, i_8_353, i_8_388, i_8_389, i_8_418, i_8_460, i_8_523, i_8_524, i_8_536, i_8_550, i_8_581, i_8_605, i_8_632, i_8_635, i_8_640, i_8_641, i_8_653, i_8_670, i_8_685, i_8_694, i_8_728, i_8_733, i_8_802, i_8_831, i_8_838, i_8_841, i_8_859, i_8_883, i_8_977, i_8_991, i_8_992, i_8_1054, i_8_1172, i_8_1199, i_8_1225, i_8_1243, i_8_1246, i_8_1247, i_8_1263, i_8_1279, i_8_1319, i_8_1354, i_8_1355, i_8_1388, i_8_1405, i_8_1408, i_8_1468, i_8_1486, i_8_1487, i_8_1496, i_8_1506, i_8_1507, i_8_1531, i_8_1542, i_8_1544, i_8_1595, i_8_1634, i_8_1648, i_8_1702, i_8_1748, i_8_1780, i_8_1801, i_8_1805, i_8_1818, i_8_1822, i_8_1847, i_8_1885, i_8_1913, i_8_1939, i_8_1940, i_8_1966, i_8_1980, i_8_1981, i_8_1993, i_8_2009, i_8_2038, i_8_2045, i_8_2052, i_8_2062, i_8_2065, i_8_2089, i_8_2122, i_8_2123, i_8_2149, i_8_2152, i_8_2227, i_8_2228, i_8_2241, i_8_2254, i_8_2256, o_8_280);
	kernel_8_281 k_8_281(i_8_24, i_8_25, i_8_52, i_8_62, i_8_76, i_8_169, i_8_204, i_8_223, i_8_328, i_8_333, i_8_348, i_8_376, i_8_384, i_8_400, i_8_429, i_8_455, i_8_490, i_8_494, i_8_503, i_8_522, i_8_526, i_8_574, i_8_583, i_8_588, i_8_592, i_8_608, i_8_613, i_8_616, i_8_642, i_8_661, i_8_750, i_8_754, i_8_759, i_8_771, i_8_773, i_8_789, i_8_845, i_8_854, i_8_895, i_8_941, i_8_944, i_8_966, i_8_998, i_8_1050, i_8_1086, i_8_1110, i_8_1111, i_8_1113, i_8_1114, i_8_1120, i_8_1123, i_8_1162, i_8_1265, i_8_1305, i_8_1308, i_8_1321, i_8_1331, i_8_1339, i_8_1348, i_8_1383, i_8_1399, i_8_1425, i_8_1426, i_8_1429, i_8_1471, i_8_1474, i_8_1509, i_8_1510, i_8_1527, i_8_1564, i_8_1565, i_8_1570, i_8_1588, i_8_1635, i_8_1636, i_8_1650, i_8_1651, i_8_1654, i_8_1689, i_8_1704, i_8_1752, i_8_1821, i_8_1822, i_8_1858, i_8_1860, i_8_1870, i_8_1876, i_8_1897, i_8_1906, i_8_1907, i_8_1978, i_8_1993, i_8_2041, i_8_2074, i_8_2091, i_8_2093, i_8_2215, i_8_2217, i_8_2227, i_8_2235, o_8_281);
	kernel_8_282 k_8_282(i_8_17, i_8_175, i_8_186, i_8_193, i_8_219, i_8_220, i_8_258, i_8_326, i_8_328, i_8_366, i_8_399, i_8_401, i_8_499, i_8_510, i_8_511, i_8_516, i_8_526, i_8_543, i_8_544, i_8_556, i_8_587, i_8_592, i_8_598, i_8_600, i_8_633, i_8_656, i_8_697, i_8_704, i_8_739, i_8_742, i_8_781, i_8_785, i_8_792, i_8_812, i_8_818, i_8_823, i_8_841, i_8_879, i_8_1014, i_8_1016, i_8_1051, i_8_1110, i_8_1123, i_8_1137, i_8_1155, i_8_1156, i_8_1158, i_8_1193, i_8_1236, i_8_1258, i_8_1274, i_8_1275, i_8_1279, i_8_1297, i_8_1302, i_8_1307, i_8_1314, i_8_1322, i_8_1330, i_8_1335, i_8_1338, i_8_1403, i_8_1462, i_8_1468, i_8_1472, i_8_1498, i_8_1560, i_8_1565, i_8_1608, i_8_1609, i_8_1636, i_8_1652, i_8_1653, i_8_1703, i_8_1706, i_8_1712, i_8_1749, i_8_1762, i_8_1774, i_8_1778, i_8_1833, i_8_1852, i_8_1886, i_8_1888, i_8_1950, i_8_1972, i_8_2055, i_8_2058, i_8_2113, i_8_2119, i_8_2157, i_8_2167, i_8_2170, i_8_2203, i_8_2211, i_8_2219, i_8_2230, i_8_2239, i_8_2244, i_8_2283, o_8_282);
	kernel_8_283 k_8_283(i_8_20, i_8_27, i_8_56, i_8_58, i_8_59, i_8_112, i_8_113, i_8_137, i_8_142, i_8_143, i_8_184, i_8_221, i_8_226, i_8_254, i_8_257, i_8_299, i_8_301, i_8_304, i_8_320, i_8_329, i_8_425, i_8_451, i_8_452, i_8_454, i_8_478, i_8_479, i_8_524, i_8_554, i_8_586, i_8_605, i_8_632, i_8_634, i_8_640, i_8_649, i_8_662, i_8_680, i_8_706, i_8_713, i_8_779, i_8_830, i_8_838, i_8_848, i_8_883, i_8_929, i_8_965, i_8_968, i_8_1049, i_8_1064, i_8_1099, i_8_1135, i_8_1136, i_8_1138, i_8_1160, i_8_1220, i_8_1228, i_8_1264, i_8_1279, i_8_1315, i_8_1366, i_8_1404, i_8_1451, i_8_1467, i_8_1471, i_8_1475, i_8_1514, i_8_1544, i_8_1631, i_8_1633, i_8_1676, i_8_1678, i_8_1687, i_8_1703, i_8_1719, i_8_1759, i_8_1769, i_8_1774, i_8_1804, i_8_1820, i_8_1856, i_8_1858, i_8_1885, i_8_1964, i_8_1976, i_8_1981, i_8_1982, i_8_1990, i_8_1991, i_8_1993, i_8_1997, i_8_2047, i_8_2072, i_8_2074, i_8_2099, i_8_2142, i_8_2144, i_8_2147, i_8_2228, i_8_2245, i_8_2279, i_8_2290, o_8_283);
	kernel_8_284 k_8_284(i_8_33, i_8_52, i_8_55, i_8_84, i_8_85, i_8_87, i_8_94, i_8_151, i_8_201, i_8_202, i_8_210, i_8_219, i_8_249, i_8_255, i_8_297, i_8_326, i_8_345, i_8_374, i_8_383, i_8_440, i_8_443, i_8_454, i_8_455, i_8_461, i_8_463, i_8_472, i_8_501, i_8_540, i_8_550, i_8_552, i_8_589, i_8_590, i_8_625, i_8_626, i_8_672, i_8_714, i_8_726, i_8_778, i_8_813, i_8_822, i_8_831, i_8_878, i_8_903, i_8_948, i_8_949, i_8_985, i_8_991, i_8_994, i_8_1029, i_8_1039, i_8_1053, i_8_1071, i_8_1083, i_8_1085, i_8_1112, i_8_1121, i_8_1138, i_8_1219, i_8_1240, i_8_1256, i_8_1259, i_8_1270, i_8_1274, i_8_1282, i_8_1283, i_8_1328, i_8_1395, i_8_1454, i_8_1472, i_8_1479, i_8_1480, i_8_1508, i_8_1509, i_8_1533, i_8_1541, i_8_1549, i_8_1555, i_8_1597, i_8_1607, i_8_1614, i_8_1615, i_8_1627, i_8_1738, i_8_1754, i_8_1759, i_8_1838, i_8_1841, i_8_1858, i_8_1864, i_8_1929, i_8_1975, i_8_2010, i_8_2047, i_8_2048, i_8_2049, i_8_2091, i_8_2109, i_8_2191, i_8_2223, i_8_2247, o_8_284);
	kernel_8_285 k_8_285(i_8_17, i_8_48, i_8_49, i_8_51, i_8_85, i_8_93, i_8_96, i_8_114, i_8_139, i_8_142, i_8_143, i_8_177, i_8_183, i_8_186, i_8_193, i_8_196, i_8_231, i_8_257, i_8_344, i_8_345, i_8_348, i_8_354, i_8_357, i_8_361, i_8_433, i_8_444, i_8_456, i_8_494, i_8_573, i_8_582, i_8_601, i_8_654, i_8_660, i_8_703, i_8_748, i_8_768, i_8_774, i_8_825, i_8_843, i_8_924, i_8_933, i_8_958, i_8_966, i_8_967, i_8_969, i_8_1059, i_8_1071, i_8_1113, i_8_1119, i_8_1121, i_8_1126, i_8_1155, i_8_1166, i_8_1182, i_8_1183, i_8_1191, i_8_1232, i_8_1305, i_8_1307, i_8_1320, i_8_1329, i_8_1362, i_8_1366, i_8_1372, i_8_1407, i_8_1411, i_8_1470, i_8_1492, i_8_1560, i_8_1563, i_8_1564, i_8_1574, i_8_1641, i_8_1644, i_8_1648, i_8_1652, i_8_1655, i_8_1681, i_8_1689, i_8_1776, i_8_1833, i_8_1842, i_8_1877, i_8_1965, i_8_1996, i_8_2004, i_8_2073, i_8_2112, i_8_2143, i_8_2149, i_8_2157, i_8_2211, i_8_2214, i_8_2215, i_8_2216, i_8_2218, i_8_2229, i_8_2230, i_8_2232, i_8_2244, o_8_285);
	kernel_8_286 k_8_286(i_8_20, i_8_33, i_8_49, i_8_63, i_8_80, i_8_82, i_8_84, i_8_139, i_8_141, i_8_157, i_8_265, i_8_282, i_8_284, i_8_285, i_8_292, i_8_319, i_8_321, i_8_324, i_8_380, i_8_403, i_8_404, i_8_436, i_8_465, i_8_534, i_8_552, i_8_581, i_8_582, i_8_601, i_8_608, i_8_610, i_8_625, i_8_633, i_8_678, i_8_708, i_8_716, i_8_723, i_8_726, i_8_736, i_8_737, i_8_795, i_8_813, i_8_870, i_8_922, i_8_931, i_8_951, i_8_980, i_8_985, i_8_991, i_8_1012, i_8_1030, i_8_1032, i_8_1110, i_8_1112, i_8_1182, i_8_1185, i_8_1236, i_8_1239, i_8_1240, i_8_1260, i_8_1261, i_8_1285, i_8_1331, i_8_1383, i_8_1401, i_8_1436, i_8_1443, i_8_1570, i_8_1614, i_8_1623, i_8_1635, i_8_1649, i_8_1675, i_8_1680, i_8_1722, i_8_1734, i_8_1736, i_8_1749, i_8_1822, i_8_1848, i_8_1858, i_8_1863, i_8_1902, i_8_1903, i_8_1911, i_8_1915, i_8_1948, i_8_1957, i_8_1960, i_8_2014, i_8_2015, i_8_2029, i_8_2031, i_8_2058, i_8_2136, i_8_2152, i_8_2153, i_8_2163, i_8_2241, i_8_2262, i_8_2266, o_8_286);
	kernel_8_287 k_8_287(i_8_41, i_8_77, i_8_80, i_8_194, i_8_202, i_8_203, i_8_247, i_8_278, i_8_301, i_8_356, i_8_358, i_8_364, i_8_367, i_8_391, i_8_392, i_8_424, i_8_460, i_8_499, i_8_527, i_8_529, i_8_536, i_8_593, i_8_607, i_8_608, i_8_610, i_8_612, i_8_614, i_8_635, i_8_638, i_8_642, i_8_648, i_8_656, i_8_664, i_8_679, i_8_703, i_8_704, i_8_706, i_8_710, i_8_812, i_8_832, i_8_833, i_8_835, i_8_840, i_8_842, i_8_857, i_8_869, i_8_873, i_8_875, i_8_956, i_8_967, i_8_970, i_8_1053, i_8_1133, i_8_1154, i_8_1174, i_8_1192, i_8_1228, i_8_1267, i_8_1285, i_8_1286, i_8_1315, i_8_1352, i_8_1382, i_8_1400, i_8_1404, i_8_1436, i_8_1438, i_8_1496, i_8_1508, i_8_1532, i_8_1551, i_8_1574, i_8_1607, i_8_1660, i_8_1670, i_8_1702, i_8_1703, i_8_1750, i_8_1751, i_8_1775, i_8_1803, i_8_1823, i_8_1825, i_8_1913, i_8_1951, i_8_1967, i_8_1996, i_8_2012, i_8_2052, i_8_2065, i_8_2107, i_8_2120, i_8_2129, i_8_2144, i_8_2145, i_8_2224, i_8_2247, i_8_2297, i_8_2299, i_8_2300, o_8_287);
	kernel_8_288 k_8_288(i_8_19, i_8_30, i_8_31, i_8_32, i_8_53, i_8_85, i_8_103, i_8_109, i_8_111, i_8_153, i_8_163, i_8_228, i_8_236, i_8_238, i_8_326, i_8_373, i_8_378, i_8_439, i_8_471, i_8_480, i_8_549, i_8_568, i_8_569, i_8_610, i_8_613, i_8_615, i_8_684, i_8_692, i_8_698, i_8_703, i_8_705, i_8_759, i_8_847, i_8_858, i_8_882, i_8_937, i_8_939, i_8_956, i_8_985, i_8_1008, i_8_1038, i_8_1039, i_8_1041, i_8_1042, i_8_1069, i_8_1118, i_8_1120, i_8_1183, i_8_1188, i_8_1260, i_8_1288, i_8_1291, i_8_1296, i_8_1306, i_8_1411, i_8_1432, i_8_1433, i_8_1435, i_8_1449, i_8_1454, i_8_1472, i_8_1532, i_8_1574, i_8_1622, i_8_1676, i_8_1696, i_8_1719, i_8_1720, i_8_1740, i_8_1746, i_8_1770, i_8_1808, i_8_1821, i_8_1828, i_8_1830, i_8_1854, i_8_1855, i_8_1881, i_8_1882, i_8_1884, i_8_1892, i_8_1901, i_8_1903, i_8_1962, i_8_1982, i_8_2044, i_8_2047, i_8_2074, i_8_2144, i_8_2147, i_8_2149, i_8_2170, i_8_2172, i_8_2190, i_8_2215, i_8_2229, i_8_2242, i_8_2272, i_8_2296, i_8_2297, o_8_288);
	kernel_8_289 k_8_289(i_8_24, i_8_26, i_8_33, i_8_57, i_8_61, i_8_88, i_8_105, i_8_142, i_8_168, i_8_177, i_8_196, i_8_228, i_8_258, i_8_303, i_8_333, i_8_336, i_8_369, i_8_393, i_8_394, i_8_420, i_8_426, i_8_465, i_8_492, i_8_539, i_8_591, i_8_595, i_8_597, i_8_600, i_8_610, i_8_642, i_8_661, i_8_690, i_8_703, i_8_708, i_8_733, i_8_754, i_8_780, i_8_840, i_8_852, i_8_867, i_8_876, i_8_888, i_8_924, i_8_958, i_8_982, i_8_993, i_8_1041, i_8_1105, i_8_1132, i_8_1176, i_8_1203, i_8_1227, i_8_1230, i_8_1231, i_8_1262, i_8_1263, i_8_1264, i_8_1281, i_8_1284, i_8_1311, i_8_1326, i_8_1362, i_8_1366, i_8_1389, i_8_1398, i_8_1407, i_8_1437, i_8_1440, i_8_1473, i_8_1501, i_8_1626, i_8_1674, i_8_1707, i_8_1749, i_8_1753, i_8_1770, i_8_1779, i_8_1786, i_8_1789, i_8_1812, i_8_1869, i_8_1875, i_8_1914, i_8_1965, i_8_1981, i_8_1983, i_8_1995, i_8_2067, i_8_2103, i_8_2136, i_8_2145, i_8_2148, i_8_2149, i_8_2151, i_8_2152, i_8_2154, i_8_2230, i_8_2235, i_8_2262, i_8_2293, o_8_289);
	kernel_8_290 k_8_290(i_8_9, i_8_135, i_8_138, i_8_139, i_8_151, i_8_173, i_8_181, i_8_233, i_8_302, i_8_392, i_8_394, i_8_398, i_8_401, i_8_423, i_8_424, i_8_463, i_8_476, i_8_506, i_8_528, i_8_532, i_8_538, i_8_554, i_8_568, i_8_576, i_8_657, i_8_670, i_8_702, i_8_748, i_8_815, i_8_829, i_8_833, i_8_839, i_8_842, i_8_890, i_8_936, i_8_964, i_8_968, i_8_970, i_8_1052, i_8_1197, i_8_1198, i_8_1199, i_8_1202, i_8_1228, i_8_1235, i_8_1253, i_8_1291, i_8_1296, i_8_1300, i_8_1314, i_8_1315, i_8_1382, i_8_1398, i_8_1400, i_8_1403, i_8_1404, i_8_1407, i_8_1436, i_8_1459, i_8_1460, i_8_1467, i_8_1486, i_8_1494, i_8_1512, i_8_1524, i_8_1525, i_8_1538, i_8_1539, i_8_1650, i_8_1684, i_8_1707, i_8_1708, i_8_1719, i_8_1720, i_8_1727, i_8_1745, i_8_1756, i_8_1786, i_8_1809, i_8_1825, i_8_1826, i_8_1840, i_8_1861, i_8_1882, i_8_1935, i_8_1952, i_8_1974, i_8_2012, i_8_2072, i_8_2096, i_8_2120, i_8_2126, i_8_2152, i_8_2170, i_8_2171, i_8_2177, i_8_2233, i_8_2253, i_8_2295, i_8_2297, o_8_290);
	kernel_8_291 k_8_291(i_8_9, i_8_31, i_8_87, i_8_88, i_8_92, i_8_111, i_8_112, i_8_135, i_8_147, i_8_189, i_8_268, i_8_280, i_8_281, i_8_295, i_8_304, i_8_339, i_8_345, i_8_347, i_8_353, i_8_370, i_8_389, i_8_396, i_8_397, i_8_415, i_8_416, i_8_418, i_8_424, i_8_448, i_8_453, i_8_489, i_8_508, i_8_522, i_8_550, i_8_568, i_8_569, i_8_657, i_8_658, i_8_701, i_8_747, i_8_766, i_8_842, i_8_844, i_8_847, i_8_892, i_8_937, i_8_938, i_8_966, i_8_1009, i_8_1010, i_8_1033, i_8_1065, i_8_1098, i_8_1109, i_8_1142, i_8_1152, i_8_1198, i_8_1281, i_8_1294, i_8_1305, i_8_1352, i_8_1393, i_8_1404, i_8_1422, i_8_1423, i_8_1487, i_8_1521, i_8_1522, i_8_1523, i_8_1530, i_8_1543, i_8_1548, i_8_1549, i_8_1604, i_8_1634, i_8_1649, i_8_1669, i_8_1670, i_8_1683, i_8_1721, i_8_1757, i_8_1765, i_8_1773, i_8_1803, i_8_1855, i_8_1889, i_8_1935, i_8_1936, i_8_1954, i_8_1955, i_8_2017, i_8_2026, i_8_2039, i_8_2161, i_8_2173, i_8_2206, i_8_2226, i_8_2243, i_8_2256, i_8_2271, i_8_2297, o_8_291);
	kernel_8_292 k_8_292(i_8_3, i_8_35, i_8_42, i_8_43, i_8_44, i_8_66, i_8_79, i_8_129, i_8_138, i_8_141, i_8_150, i_8_190, i_8_202, i_8_355, i_8_384, i_8_421, i_8_498, i_8_499, i_8_500, i_8_507, i_8_553, i_8_554, i_8_594, i_8_607, i_8_624, i_8_642, i_8_643, i_8_656, i_8_789, i_8_811, i_8_828, i_8_831, i_8_840, i_8_876, i_8_877, i_8_880, i_8_958, i_8_1005, i_8_1039, i_8_1053, i_8_1083, i_8_1132, i_8_1155, i_8_1156, i_8_1200, i_8_1230, i_8_1272, i_8_1317, i_8_1318, i_8_1321, i_8_1326, i_8_1350, i_8_1372, i_8_1384, i_8_1385, i_8_1389, i_8_1390, i_8_1393, i_8_1399, i_8_1402, i_8_1449, i_8_1473, i_8_1483, i_8_1485, i_8_1486, i_8_1498, i_8_1503, i_8_1524, i_8_1533, i_8_1599, i_8_1615, i_8_1652, i_8_1654, i_8_1696, i_8_1753, i_8_1828, i_8_1876, i_8_1887, i_8_1897, i_8_1915, i_8_1950, i_8_1981, i_8_1996, i_8_2010, i_8_2011, i_8_2023, i_8_2035, i_8_2043, i_8_2053, i_8_2068, i_8_2082, i_8_2089, i_8_2093, i_8_2122, i_8_2150, i_8_2173, i_8_2185, i_8_2237, i_8_2249, i_8_2284, o_8_292);
	kernel_8_293 k_8_293(i_8_50, i_8_60, i_8_61, i_8_62, i_8_96, i_8_125, i_8_141, i_8_143, i_8_185, i_8_189, i_8_229, i_8_259, i_8_260, i_8_303, i_8_308, i_8_349, i_8_365, i_8_366, i_8_382, i_8_420, i_8_427, i_8_448, i_8_449, i_8_456, i_8_457, i_8_511, i_8_555, i_8_556, i_8_591, i_8_592, i_8_602, i_8_617, i_8_622, i_8_633, i_8_636, i_8_768, i_8_789, i_8_790, i_8_795, i_8_818, i_8_826, i_8_827, i_8_845, i_8_857, i_8_881, i_8_969, i_8_970, i_8_995, i_8_1051, i_8_1076, i_8_1124, i_8_1228, i_8_1237, i_8_1268, i_8_1282, i_8_1283, i_8_1284, i_8_1285, i_8_1286, i_8_1295, i_8_1314, i_8_1319, i_8_1331, i_8_1407, i_8_1408, i_8_1439, i_8_1473, i_8_1474, i_8_1484, i_8_1541, i_8_1547, i_8_1574, i_8_1601, i_8_1605, i_8_1626, i_8_1635, i_8_1648, i_8_1649, i_8_1653, i_8_1669, i_8_1679, i_8_1724, i_8_1736, i_8_1747, i_8_1773, i_8_1857, i_8_1948, i_8_2031, i_8_2033, i_8_2046, i_8_2095, i_8_2096, i_8_2151, i_8_2152, i_8_2217, i_8_2218, i_8_2219, i_8_2226, i_8_2243, i_8_2286, o_8_293);
	kernel_8_294 k_8_294(i_8_13, i_8_63, i_8_66, i_8_75, i_8_129, i_8_183, i_8_204, i_8_237, i_8_309, i_8_336, i_8_345, i_8_354, i_8_450, i_8_453, i_8_475, i_8_489, i_8_490, i_8_504, i_8_552, i_8_555, i_8_591, i_8_597, i_8_608, i_8_637, i_8_658, i_8_662, i_8_664, i_8_682, i_8_690, i_8_697, i_8_728, i_8_765, i_8_768, i_8_769, i_8_771, i_8_795, i_8_804, i_8_825, i_8_921, i_8_930, i_8_933, i_8_970, i_8_1029, i_8_1056, i_8_1060, i_8_1072, i_8_1074, i_8_1089, i_8_1168, i_8_1173, i_8_1176, i_8_1254, i_8_1264, i_8_1266, i_8_1267, i_8_1275, i_8_1297, i_8_1305, i_8_1440, i_8_1470, i_8_1536, i_8_1554, i_8_1560, i_8_1563, i_8_1596, i_8_1605, i_8_1621, i_8_1641, i_8_1645, i_8_1668, i_8_1680, i_8_1704, i_8_1737, i_8_1747, i_8_1759, i_8_1767, i_8_1770, i_8_1778, i_8_1821, i_8_1830, i_8_1831, i_8_1857, i_8_1861, i_8_1875, i_8_1879, i_8_1885, i_8_1929, i_8_1965, i_8_2017, i_8_2019, i_8_2059, i_8_2119, i_8_2148, i_8_2169, i_8_2182, i_8_2184, i_8_2194, i_8_2211, i_8_2215, i_8_2291, o_8_294);
	kernel_8_295 k_8_295(i_8_1, i_8_22, i_8_73, i_8_75, i_8_115, i_8_137, i_8_148, i_8_226, i_8_229, i_8_302, i_8_319, i_8_364, i_8_380, i_8_388, i_8_400, i_8_425, i_8_454, i_8_490, i_8_497, i_8_508, i_8_528, i_8_552, i_8_599, i_8_602, i_8_605, i_8_607, i_8_635, i_8_641, i_8_659, i_8_660, i_8_676, i_8_680, i_8_695, i_8_696, i_8_706, i_8_710, i_8_757, i_8_814, i_8_815, i_8_860, i_8_968, i_8_1013, i_8_1103, i_8_1108, i_8_1111, i_8_1202, i_8_1228, i_8_1264, i_8_1273, i_8_1307, i_8_1311, i_8_1328, i_8_1358, i_8_1387, i_8_1388, i_8_1414, i_8_1424, i_8_1432, i_8_1462, i_8_1463, i_8_1466, i_8_1474, i_8_1478, i_8_1511, i_8_1517, i_8_1526, i_8_1557, i_8_1633, i_8_1648, i_8_1667, i_8_1678, i_8_1691, i_8_1697, i_8_1750, i_8_1766, i_8_1769, i_8_1772, i_8_1775, i_8_1787, i_8_1789, i_8_1792, i_8_1807, i_8_1811, i_8_1841, i_8_1846, i_8_1910, i_8_1927, i_8_1940, i_8_1958, i_8_1964, i_8_1972, i_8_1976, i_8_1981, i_8_1982, i_8_1997, i_8_2002, i_8_2020, i_8_2055, i_8_2119, i_8_2149, o_8_295);
	kernel_8_296 k_8_296(i_8_0, i_8_1, i_8_104, i_8_155, i_8_163, i_8_216, i_8_232, i_8_233, i_8_262, i_8_289, i_8_325, i_8_326, i_8_366, i_8_432, i_8_433, i_8_480, i_8_481, i_8_486, i_8_489, i_8_550, i_8_556, i_8_603, i_8_621, i_8_630, i_8_694, i_8_695, i_8_696, i_8_697, i_8_701, i_8_709, i_8_721, i_8_783, i_8_802, i_8_811, i_8_812, i_8_820, i_8_825, i_8_827, i_8_840, i_8_865, i_8_874, i_8_967, i_8_970, i_8_973, i_8_996, i_8_1071, i_8_1154, i_8_1180, i_8_1207, i_8_1208, i_8_1224, i_8_1233, i_8_1234, i_8_1260, i_8_1270, i_8_1352, i_8_1360, i_8_1367, i_8_1387, i_8_1399, i_8_1435, i_8_1452, i_8_1537, i_8_1542, i_8_1548, i_8_1571, i_8_1584, i_8_1585, i_8_1622, i_8_1624, i_8_1650, i_8_1651, i_8_1720, i_8_1747, i_8_1770, i_8_1774, i_8_1818, i_8_1864, i_8_1874, i_8_1989, i_8_2025, i_8_2026, i_8_2034, i_8_2035, i_8_2038, i_8_2088, i_8_2116, i_8_2144, i_8_2147, i_8_2152, i_8_2153, i_8_2155, i_8_2188, i_8_2269, i_8_2272, i_8_2279, i_8_2281, i_8_2286, i_8_2289, i_8_2297, o_8_296);
	kernel_8_297 k_8_297(i_8_29, i_8_82, i_8_100, i_8_154, i_8_162, i_8_171, i_8_175, i_8_190, i_8_218, i_8_257, i_8_259, i_8_266, i_8_281, i_8_339, i_8_379, i_8_380, i_8_427, i_8_436, i_8_437, i_8_459, i_8_478, i_8_572, i_8_587, i_8_598, i_8_621, i_8_626, i_8_684, i_8_696, i_8_703, i_8_707, i_8_716, i_8_757, i_8_761, i_8_775, i_8_778, i_8_802, i_8_821, i_8_876, i_8_991, i_8_992, i_8_1108, i_8_1111, i_8_1135, i_8_1136, i_8_1153, i_8_1157, i_8_1170, i_8_1180, i_8_1261, i_8_1279, i_8_1283, i_8_1306, i_8_1325, i_8_1352, i_8_1370, i_8_1381, i_8_1405, i_8_1407, i_8_1418, i_8_1433, i_8_1460, i_8_1472, i_8_1481, i_8_1487, i_8_1551, i_8_1568, i_8_1603, i_8_1611, i_8_1625, i_8_1642, i_8_1669, i_8_1675, i_8_1697, i_8_1737, i_8_1753, i_8_1759, i_8_1773, i_8_1774, i_8_1801, i_8_1805, i_8_1811, i_8_1823, i_8_1928, i_8_1946, i_8_1981, i_8_1992, i_8_1994, i_8_2054, i_8_2107, i_8_2112, i_8_2150, i_8_2151, i_8_2152, i_8_2189, i_8_2225, i_8_2241, i_8_2259, i_8_2287, i_8_2288, i_8_2299, o_8_297);
	kernel_8_298 k_8_298(i_8_0, i_8_1, i_8_40, i_8_79, i_8_83, i_8_104, i_8_112, i_8_143, i_8_166, i_8_167, i_8_190, i_8_208, i_8_259, i_8_265, i_8_280, i_8_281, i_8_289, i_8_290, i_8_299, i_8_308, i_8_310, i_8_317, i_8_319, i_8_418, i_8_424, i_8_437, i_8_451, i_8_488, i_8_585, i_8_589, i_8_641, i_8_651, i_8_670, i_8_693, i_8_701, i_8_703, i_8_704, i_8_710, i_8_730, i_8_767, i_8_778, i_8_779, i_8_824, i_8_847, i_8_929, i_8_967, i_8_976, i_8_991, i_8_992, i_8_1028, i_8_1180, i_8_1234, i_8_1235, i_8_1256, i_8_1262, i_8_1283, i_8_1300, i_8_1316, i_8_1330, i_8_1352, i_8_1360, i_8_1384, i_8_1405, i_8_1438, i_8_1441, i_8_1442, i_8_1459, i_8_1486, i_8_1507, i_8_1541, i_8_1558, i_8_1585, i_8_1586, i_8_1639, i_8_1651, i_8_1682, i_8_1765, i_8_1766, i_8_1811, i_8_1823, i_8_1824, i_8_1838, i_8_1846, i_8_1982, i_8_1993, i_8_1994, i_8_1999, i_8_2026, i_8_2053, i_8_2074, i_8_2125, i_8_2126, i_8_2147, i_8_2158, i_8_2188, i_8_2189, i_8_2196, i_8_2224, i_8_2233, i_8_2242, o_8_298);
	kernel_8_299 k_8_299(i_8_31, i_8_89, i_8_96, i_8_98, i_8_196, i_8_237, i_8_240, i_8_241, i_8_295, i_8_296, i_8_312, i_8_324, i_8_349, i_8_372, i_8_424, i_8_480, i_8_528, i_8_529, i_8_556, i_8_605, i_8_733, i_8_735, i_8_736, i_8_763, i_8_778, i_8_779, i_8_781, i_8_789, i_8_797, i_8_815, i_8_837, i_8_862, i_8_940, i_8_941, i_8_943, i_8_947, i_8_996, i_8_1005, i_8_1012, i_8_1015, i_8_1060, i_8_1114, i_8_1115, i_8_1127, i_8_1130, i_8_1195, i_8_1219, i_8_1223, i_8_1292, i_8_1294, i_8_1306, i_8_1307, i_8_1310, i_8_1311, i_8_1314, i_8_1336, i_8_1410, i_8_1438, i_8_1472, i_8_1537, i_8_1538, i_8_1544, i_8_1597, i_8_1609, i_8_1632, i_8_1645, i_8_1649, i_8_1667, i_8_1668, i_8_1677, i_8_1707, i_8_1722, i_8_1723, i_8_1724, i_8_1743, i_8_1763, i_8_1814, i_8_1815, i_8_1816, i_8_1825, i_8_1831, i_8_1894, i_8_1907, i_8_1919, i_8_1970, i_8_2003, i_8_2041, i_8_2047, i_8_2109, i_8_2121, i_8_2174, i_8_2177, i_8_2202, i_8_2203, i_8_2212, i_8_2215, i_8_2256, i_8_2257, i_8_2274, i_8_2298, o_8_299);
	kernel_8_300 k_8_300(i_8_22, i_8_23, i_8_53, i_8_115, i_8_121, i_8_142, i_8_143, i_8_188, i_8_212, i_8_229, i_8_304, i_8_382, i_8_383, i_8_384, i_8_385, i_8_386, i_8_419, i_8_421, i_8_422, i_8_464, i_8_484, i_8_485, i_8_556, i_8_572, i_8_575, i_8_591, i_8_598, i_8_599, i_8_637, i_8_673, i_8_695, i_8_832, i_8_841, i_8_854, i_8_880, i_8_896, i_8_966, i_8_968, i_8_995, i_8_1015, i_8_1039, i_8_1040, i_8_1132, i_8_1225, i_8_1228, i_8_1232, i_8_1233, i_8_1255, i_8_1258, i_8_1259, i_8_1273, i_8_1277, i_8_1283, i_8_1284, i_8_1427, i_8_1438, i_8_1472, i_8_1474, i_8_1475, i_8_1481, i_8_1484, i_8_1490, i_8_1525, i_8_1526, i_8_1528, i_8_1529, i_8_1553, i_8_1556, i_8_1621, i_8_1643, i_8_1649, i_8_1655, i_8_1688, i_8_1696, i_8_1697, i_8_1723, i_8_1726, i_8_1727, i_8_1752, i_8_1771, i_8_1776, i_8_1795, i_8_1904, i_8_1944, i_8_1966, i_8_1973, i_8_2014, i_8_2038, i_8_2050, i_8_2093, i_8_2137, i_8_2150, i_8_2153, i_8_2155, i_8_2156, i_8_2158, i_8_2203, i_8_2233, i_8_2272, i_8_2275, o_8_300);
	kernel_8_301 k_8_301(i_8_40, i_8_41, i_8_43, i_8_44, i_8_97, i_8_118, i_8_170, i_8_178, i_8_239, i_8_242, i_8_256, i_8_259, i_8_260, i_8_269, i_8_301, i_8_304, i_8_305, i_8_347, i_8_363, i_8_377, i_8_380, i_8_401, i_8_430, i_8_453, i_8_454, i_8_456, i_8_494, i_8_528, i_8_584, i_8_634, i_8_638, i_8_647, i_8_662, i_8_679, i_8_680, i_8_692, i_8_698, i_8_709, i_8_796, i_8_842, i_8_855, i_8_886, i_8_955, i_8_1060, i_8_1080, i_8_1125, i_8_1192, i_8_1228, i_8_1237, i_8_1261, i_8_1274, i_8_1282, i_8_1285, i_8_1295, i_8_1308, i_8_1310, i_8_1336, i_8_1352, i_8_1354, i_8_1373, i_8_1411, i_8_1416, i_8_1419, i_8_1456, i_8_1457, i_8_1610, i_8_1615, i_8_1642, i_8_1645, i_8_1673, i_8_1690, i_8_1691, i_8_1703, i_8_1787, i_8_1855, i_8_1857, i_8_1859, i_8_1886, i_8_1922, i_8_1940, i_8_1970, i_8_1982, i_8_1989, i_8_1993, i_8_2003, i_8_2005, i_8_2006, i_8_2056, i_8_2113, i_8_2114, i_8_2154, i_8_2156, i_8_2159, i_8_2201, i_8_2213, i_8_2223, i_8_2257, i_8_2261, i_8_2284, i_8_2285, o_8_301);
	kernel_8_302 k_8_302(i_8_28, i_8_40, i_8_227, i_8_259, i_8_275, i_8_318, i_8_335, i_8_348, i_8_390, i_8_398, i_8_401, i_8_418, i_8_422, i_8_427, i_8_451, i_8_506, i_8_508, i_8_509, i_8_552, i_8_553, i_8_554, i_8_572, i_8_603, i_8_604, i_8_631, i_8_638, i_8_651, i_8_705, i_8_707, i_8_710, i_8_749, i_8_884, i_8_895, i_8_896, i_8_1011, i_8_1040, i_8_1052, i_8_1058, i_8_1103, i_8_1106, i_8_1107, i_8_1112, i_8_1138, i_8_1139, i_8_1154, i_8_1180, i_8_1202, i_8_1235, i_8_1238, i_8_1244, i_8_1279, i_8_1305, i_8_1319, i_8_1362, i_8_1364, i_8_1422, i_8_1427, i_8_1429, i_8_1436, i_8_1458, i_8_1461, i_8_1462, i_8_1463, i_8_1471, i_8_1479, i_8_1480, i_8_1487, i_8_1508, i_8_1511, i_8_1512, i_8_1515, i_8_1524, i_8_1551, i_8_1569, i_8_1678, i_8_1702, i_8_1705, i_8_1706, i_8_1774, i_8_1776, i_8_1784, i_8_1795, i_8_1836, i_8_1839, i_8_1841, i_8_1892, i_8_1919, i_8_1955, i_8_1974, i_8_1997, i_8_2057, i_8_2075, i_8_2151, i_8_2155, i_8_2223, i_8_2224, i_8_2225, i_8_2245, i_8_2248, i_8_2249, o_8_302);
	kernel_8_303 k_8_303(i_8_20, i_8_107, i_8_240, i_8_255, i_8_324, i_8_325, i_8_328, i_8_345, i_8_348, i_8_380, i_8_382, i_8_391, i_8_440, i_8_460, i_8_469, i_8_474, i_8_478, i_8_483, i_8_507, i_8_523, i_8_524, i_8_527, i_8_549, i_8_551, i_8_552, i_8_599, i_8_604, i_8_637, i_8_712, i_8_715, i_8_732, i_8_757, i_8_763, i_8_778, i_8_800, i_8_943, i_8_945, i_8_946, i_8_947, i_8_990, i_8_997, i_8_1050, i_8_1072, i_8_1075, i_8_1110, i_8_1114, i_8_1117, i_8_1130, i_8_1169, i_8_1176, i_8_1190, i_8_1238, i_8_1257, i_8_1273, i_8_1284, i_8_1315, i_8_1323, i_8_1324, i_8_1326, i_8_1347, i_8_1387, i_8_1417, i_8_1438, i_8_1441, i_8_1452, i_8_1506, i_8_1530, i_8_1534, i_8_1562, i_8_1649, i_8_1671, i_8_1681, i_8_1716, i_8_1722, i_8_1723, i_8_1726, i_8_1732, i_8_1746, i_8_1833, i_8_1841, i_8_1854, i_8_1864, i_8_1887, i_8_1894, i_8_1949, i_8_1965, i_8_1992, i_8_2002, i_8_2028, i_8_2031, i_8_2032, i_8_2051, i_8_2064, i_8_2092, i_8_2115, i_8_2175, i_8_2215, i_8_2216, i_8_2219, i_8_2283, o_8_303);
	kernel_8_304 k_8_304(i_8_19, i_8_39, i_8_87, i_8_111, i_8_112, i_8_113, i_8_219, i_8_245, i_8_266, i_8_269, i_8_286, i_8_287, i_8_295, i_8_296, i_8_304, i_8_305, i_8_381, i_8_383, i_8_427, i_8_428, i_8_429, i_8_430, i_8_431, i_8_504, i_8_524, i_8_567, i_8_568, i_8_569, i_8_577, i_8_578, i_8_606, i_8_607, i_8_635, i_8_705, i_8_708, i_8_709, i_8_710, i_8_713, i_8_715, i_8_726, i_8_816, i_8_817, i_8_838, i_8_846, i_8_847, i_8_878, i_8_1078, i_8_1179, i_8_1180, i_8_1181, i_8_1189, i_8_1266, i_8_1315, i_8_1329, i_8_1359, i_8_1365, i_8_1394, i_8_1399, i_8_1467, i_8_1468, i_8_1469, i_8_1470, i_8_1472, i_8_1522, i_8_1534, i_8_1565, i_8_1621, i_8_1683, i_8_1684, i_8_1693, i_8_1694, i_8_1730, i_8_1747, i_8_1749, i_8_1765, i_8_1777, i_8_1780, i_8_1784, i_8_1785, i_8_1786, i_8_1787, i_8_1825, i_8_1826, i_8_1854, i_8_1873, i_8_1874, i_8_1889, i_8_1920, i_8_1946, i_8_2060, i_8_2070, i_8_2071, i_8_2088, i_8_2138, i_8_2139, i_8_2226, i_8_2227, i_8_2233, i_8_2243, i_8_2274, o_8_304);
	kernel_8_305 k_8_305(i_8_21, i_8_30, i_8_31, i_8_35, i_8_53, i_8_57, i_8_114, i_8_116, i_8_142, i_8_143, i_8_171, i_8_188, i_8_192, i_8_225, i_8_238, i_8_246, i_8_395, i_8_415, i_8_422, i_8_446, i_8_585, i_8_598, i_8_599, i_8_611, i_8_698, i_8_701, i_8_716, i_8_759, i_8_780, i_8_781, i_8_815, i_8_818, i_8_823, i_8_841, i_8_845, i_8_849, i_8_853, i_8_888, i_8_959, i_8_964, i_8_1016, i_8_1030, i_8_1034, i_8_1050, i_8_1051, i_8_1060, i_8_1114, i_8_1121, i_8_1160, i_8_1182, i_8_1183, i_8_1281, i_8_1282, i_8_1283, i_8_1284, i_8_1291, i_8_1300, i_8_1305, i_8_1306, i_8_1307, i_8_1330, i_8_1344, i_8_1347, i_8_1390, i_8_1391, i_8_1410, i_8_1437, i_8_1438, i_8_1453, i_8_1470, i_8_1471, i_8_1552, i_8_1574, i_8_1652, i_8_1677, i_8_1683, i_8_1699, i_8_1754, i_8_1875, i_8_1876, i_8_1877, i_8_1984, i_8_1988, i_8_1991, i_8_1992, i_8_1995, i_8_2033, i_8_2071, i_8_2076, i_8_2093, i_8_2114, i_8_2132, i_8_2151, i_8_2214, i_8_2215, i_8_2216, i_8_2237, i_8_2245, i_8_2261, i_8_2290, o_8_305);
	kernel_8_306 k_8_306(i_8_9, i_8_10, i_8_47, i_8_112, i_8_118, i_8_136, i_8_137, i_8_139, i_8_140, i_8_221, i_8_230, i_8_265, i_8_316, i_8_383, i_8_391, i_8_398, i_8_414, i_8_415, i_8_417, i_8_425, i_8_427, i_8_478, i_8_481, i_8_510, i_8_522, i_8_524, i_8_526, i_8_528, i_8_553, i_8_554, i_8_568, i_8_577, i_8_585, i_8_632, i_8_640, i_8_651, i_8_704, i_8_730, i_8_784, i_8_792, i_8_793, i_8_823, i_8_837, i_8_847, i_8_859, i_8_874, i_8_887, i_8_892, i_8_964, i_8_991, i_8_1036, i_8_1072, i_8_1111, i_8_1199, i_8_1237, i_8_1315, i_8_1324, i_8_1352, i_8_1354, i_8_1360, i_8_1372, i_8_1388, i_8_1396, i_8_1438, i_8_1458, i_8_1459, i_8_1470, i_8_1477, i_8_1513, i_8_1521, i_8_1540, i_8_1566, i_8_1567, i_8_1571, i_8_1603, i_8_1630, i_8_1684, i_8_1693, i_8_1720, i_8_1751, i_8_1776, i_8_1777, i_8_1778, i_8_1781, i_8_1786, i_8_1837, i_8_1864, i_8_1885, i_8_1900, i_8_1935, i_8_1936, i_8_1954, i_8_1972, i_8_1993, i_8_2026, i_8_2092, i_8_2138, i_8_2147, i_8_2170, i_8_2241, o_8_306);
	kernel_8_307 k_8_307(i_8_85, i_8_88, i_8_91, i_8_181, i_8_189, i_8_190, i_8_220, i_8_292, i_8_305, i_8_370, i_8_372, i_8_417, i_8_418, i_8_476, i_8_481, i_8_483, i_8_546, i_8_556, i_8_595, i_8_634, i_8_648, i_8_672, i_8_703, i_8_705, i_8_728, i_8_759, i_8_764, i_8_797, i_8_811, i_8_855, i_8_872, i_8_898, i_8_899, i_8_966, i_8_991, i_8_1000, i_8_1030, i_8_1060, i_8_1061, i_8_1111, i_8_1121, i_8_1179, i_8_1191, i_8_1285, i_8_1291, i_8_1296, i_8_1297, i_8_1305, i_8_1316, i_8_1319, i_8_1323, i_8_1327, i_8_1455, i_8_1456, i_8_1469, i_8_1490, i_8_1509, i_8_1528, i_8_1529, i_8_1531, i_8_1544, i_8_1553, i_8_1561, i_8_1588, i_8_1603, i_8_1618, i_8_1669, i_8_1678, i_8_1718, i_8_1737, i_8_1738, i_8_1752, i_8_1753, i_8_1754, i_8_1761, i_8_1803, i_8_1805, i_8_1808, i_8_1839, i_8_1857, i_8_1867, i_8_1874, i_8_1904, i_8_1906, i_8_1911, i_8_1933, i_8_1981, i_8_2006, i_8_2032, i_8_2046, i_8_2047, i_8_2116, i_8_2142, i_8_2152, i_8_2153, i_8_2216, i_8_2218, i_8_2254, i_8_2290, i_8_2296, o_8_307);
	kernel_8_308 k_8_308(i_8_22, i_8_23, i_8_28, i_8_50, i_8_140, i_8_202, i_8_260, i_8_262, i_8_263, i_8_281, i_8_289, i_8_291, i_8_301, i_8_302, i_8_322, i_8_345, i_8_346, i_8_362, i_8_375, i_8_381, i_8_382, i_8_391, i_8_460, i_8_505, i_8_517, i_8_523, i_8_525, i_8_526, i_8_529, i_8_553, i_8_670, i_8_702, i_8_763, i_8_769, i_8_775, i_8_804, i_8_805, i_8_832, i_8_892, i_8_905, i_8_968, i_8_971, i_8_1067, i_8_1074, i_8_1138, i_8_1173, i_8_1182, i_8_1233, i_8_1254, i_8_1255, i_8_1260, i_8_1273, i_8_1279, i_8_1281, i_8_1282, i_8_1286, i_8_1300, i_8_1327, i_8_1384, i_8_1424, i_8_1435, i_8_1452, i_8_1467, i_8_1490, i_8_1498, i_8_1528, i_8_1533, i_8_1542, i_8_1555, i_8_1587, i_8_1597, i_8_1606, i_8_1630, i_8_1631, i_8_1632, i_8_1654, i_8_1660, i_8_1690, i_8_1696, i_8_1719, i_8_1720, i_8_1723, i_8_1724, i_8_1740, i_8_1762, i_8_1792, i_8_1808, i_8_1820, i_8_1837, i_8_1876, i_8_1990, i_8_2047, i_8_2089, i_8_2118, i_8_2126, i_8_2143, i_8_2154, i_8_2188, i_8_2234, i_8_2290, o_8_308);
	kernel_8_309 k_8_309(i_8_46, i_8_52, i_8_87, i_8_142, i_8_171, i_8_172, i_8_210, i_8_259, i_8_294, i_8_334, i_8_364, i_8_376, i_8_381, i_8_383, i_8_390, i_8_436, i_8_487, i_8_489, i_8_492, i_8_532, i_8_534, i_8_550, i_8_551, i_8_576, i_8_581, i_8_585, i_8_609, i_8_630, i_8_676, i_8_684, i_8_699, i_8_736, i_8_765, i_8_766, i_8_769, i_8_792, i_8_795, i_8_839, i_8_841, i_8_879, i_8_880, i_8_919, i_8_927, i_8_930, i_8_965, i_8_966, i_8_991, i_8_1036, i_8_1053, i_8_1171, i_8_1233, i_8_1234, i_8_1255, i_8_1263, i_8_1266, i_8_1288, i_8_1308, i_8_1315, i_8_1316, i_8_1393, i_8_1455, i_8_1471, i_8_1544, i_8_1558, i_8_1642, i_8_1650, i_8_1668, i_8_1669, i_8_1683, i_8_1702, i_8_1729, i_8_1749, i_8_1777, i_8_1821, i_8_1828, i_8_1854, i_8_1857, i_8_1858, i_8_1861, i_8_1885, i_8_1938, i_8_1947, i_8_1950, i_8_1981, i_8_1989, i_8_2001, i_8_2016, i_8_2017, i_8_2056, i_8_2106, i_8_2139, i_8_2152, i_8_2155, i_8_2182, i_8_2196, i_8_2199, i_8_2205, i_8_2259, i_8_2272, i_8_2277, o_8_309);
	kernel_8_310 k_8_310(i_8_22, i_8_54, i_8_64, i_8_219, i_8_220, i_8_283, i_8_319, i_8_321, i_8_397, i_8_424, i_8_441, i_8_496, i_8_504, i_8_524, i_8_526, i_8_571, i_8_580, i_8_589, i_8_596, i_8_613, i_8_622, i_8_642, i_8_659, i_8_660, i_8_675, i_8_676, i_8_699, i_8_700, i_8_707, i_8_730, i_8_750, i_8_751, i_8_766, i_8_812, i_8_814, i_8_822, i_8_837, i_8_838, i_8_874, i_8_877, i_8_883, i_8_914, i_8_919, i_8_938, i_8_959, i_8_1036, i_8_1071, i_8_1072, i_8_1108, i_8_1129, i_8_1153, i_8_1198, i_8_1201, i_8_1237, i_8_1243, i_8_1260, i_8_1265, i_8_1266, i_8_1318, i_8_1327, i_8_1335, i_8_1338, i_8_1355, i_8_1381, i_8_1441, i_8_1462, i_8_1480, i_8_1524, i_8_1539, i_8_1544, i_8_1630, i_8_1646, i_8_1647, i_8_1651, i_8_1667, i_8_1676, i_8_1687, i_8_1701, i_8_1702, i_8_1707, i_8_1747, i_8_1749, i_8_1765, i_8_1796, i_8_1800, i_8_1855, i_8_1864, i_8_1868, i_8_1957, i_8_1989, i_8_1993, i_8_1996, i_8_2044, i_8_2106, i_8_2148, i_8_2154, i_8_2226, i_8_2245, i_8_2290, i_8_2298, o_8_310);
	kernel_8_311 k_8_311(i_8_4, i_8_76, i_8_77, i_8_104, i_8_121, i_8_130, i_8_263, i_8_356, i_8_360, i_8_427, i_8_445, i_8_455, i_8_496, i_8_497, i_8_517, i_8_526, i_8_551, i_8_554, i_8_572, i_8_597, i_8_609, i_8_611, i_8_612, i_8_647, i_8_656, i_8_661, i_8_680, i_8_707, i_8_749, i_8_751, i_8_828, i_8_832, i_8_836, i_8_837, i_8_840, i_8_845, i_8_850, i_8_913, i_8_958, i_8_963, i_8_1003, i_8_1108, i_8_1109, i_8_1111, i_8_1129, i_8_1130, i_8_1154, i_8_1156, i_8_1177, i_8_1229, i_8_1234, i_8_1270, i_8_1299, i_8_1318, i_8_1322, i_8_1325, i_8_1390, i_8_1391, i_8_1399, i_8_1455, i_8_1460, i_8_1470, i_8_1493, i_8_1498, i_8_1598, i_8_1634, i_8_1643, i_8_1652, i_8_1706, i_8_1747, i_8_1757, i_8_1784, i_8_1807, i_8_1818, i_8_1844, i_8_1846, i_8_1849, i_8_1930, i_8_1972, i_8_1992, i_8_1993, i_8_2040, i_8_2041, i_8_2044, i_8_2065, i_8_2123, i_8_2134, i_8_2141, i_8_2145, i_8_2147, i_8_2149, i_8_2150, i_8_2159, i_8_2174, i_8_2176, i_8_2183, i_8_2228, i_8_2231, i_8_2248, i_8_2273, o_8_311);
	kernel_8_312 k_8_312(i_8_23, i_8_26, i_8_34, i_8_120, i_8_139, i_8_148, i_8_202, i_8_239, i_8_275, i_8_278, i_8_308, i_8_310, i_8_365, i_8_384, i_8_425, i_8_453, i_8_490, i_8_491, i_8_522, i_8_523, i_8_552, i_8_553, i_8_569, i_8_608, i_8_612, i_8_667, i_8_734, i_8_748, i_8_760, i_8_767, i_8_771, i_8_787, i_8_800, i_8_814, i_8_828, i_8_838, i_8_844, i_8_874, i_8_964, i_8_970, i_8_985, i_8_993, i_8_996, i_8_1021, i_8_1050, i_8_1067, i_8_1084, i_8_1102, i_8_1131, i_8_1135, i_8_1234, i_8_1238, i_8_1264, i_8_1267, i_8_1284, i_8_1305, i_8_1357, i_8_1381, i_8_1400, i_8_1408, i_8_1432, i_8_1437, i_8_1452, i_8_1508, i_8_1531, i_8_1544, i_8_1607, i_8_1643, i_8_1666, i_8_1667, i_8_1669, i_8_1671, i_8_1678, i_8_1747, i_8_1754, i_8_1757, i_8_1810, i_8_1822, i_8_1843, i_8_1883, i_8_1887, i_8_1927, i_8_1966, i_8_2000, i_8_2008, i_8_2009, i_8_2023, i_8_2070, i_8_2084, i_8_2143, i_8_2151, i_8_2153, i_8_2164, i_8_2165, i_8_2170, i_8_2176, i_8_2224, i_8_2245, i_8_2264, i_8_2273, o_8_312);
	kernel_8_313 k_8_313(i_8_18, i_8_41, i_8_59, i_8_88, i_8_115, i_8_143, i_8_188, i_8_234, i_8_266, i_8_283, i_8_284, i_8_361, i_8_362, i_8_379, i_8_383, i_8_481, i_8_493, i_8_524, i_8_525, i_8_554, i_8_569, i_8_610, i_8_635, i_8_679, i_8_682, i_8_693, i_8_698, i_8_704, i_8_709, i_8_724, i_8_735, i_8_754, i_8_762, i_8_771, i_8_773, i_8_787, i_8_789, i_8_799, i_8_841, i_8_958, i_8_964, i_8_970, i_8_1075, i_8_1106, i_8_1109, i_8_1256, i_8_1268, i_8_1301, i_8_1305, i_8_1351, i_8_1363, i_8_1399, i_8_1436, i_8_1455, i_8_1467, i_8_1471, i_8_1481, i_8_1489, i_8_1490, i_8_1529, i_8_1534, i_8_1606, i_8_1644, i_8_1649, i_8_1652, i_8_1670, i_8_1689, i_8_1703, i_8_1723, i_8_1725, i_8_1751, i_8_1752, i_8_1759, i_8_1765, i_8_1795, i_8_1804, i_8_1826, i_8_1838, i_8_1848, i_8_1849, i_8_1866, i_8_1867, i_8_1882, i_8_1886, i_8_1912, i_8_1919, i_8_1982, i_8_2001, i_8_2028, i_8_2075, i_8_2092, i_8_2142, i_8_2194, i_8_2224, i_8_2229, i_8_2230, i_8_2232, i_8_2242, i_8_2248, i_8_2264, o_8_313);
	kernel_8_314 k_8_314(i_8_33, i_8_85, i_8_100, i_8_135, i_8_183, i_8_207, i_8_208, i_8_209, i_8_217, i_8_220, i_8_223, i_8_304, i_8_326, i_8_362, i_8_450, i_8_452, i_8_493, i_8_498, i_8_514, i_8_523, i_8_540, i_8_605, i_8_612, i_8_621, i_8_631, i_8_632, i_8_634, i_8_715, i_8_721, i_8_725, i_8_734, i_8_759, i_8_766, i_8_767, i_8_769, i_8_779, i_8_796, i_8_833, i_8_864, i_8_880, i_8_883, i_8_901, i_8_903, i_8_918, i_8_947, i_8_983, i_8_991, i_8_1031, i_8_1066, i_8_1072, i_8_1073, i_8_1172, i_8_1174, i_8_1246, i_8_1247, i_8_1256, i_8_1288, i_8_1324, i_8_1417, i_8_1538, i_8_1555, i_8_1556, i_8_1561, i_8_1565, i_8_1576, i_8_1606, i_8_1613, i_8_1665, i_8_1670, i_8_1675, i_8_1681, i_8_1684, i_8_1703, i_8_1710, i_8_1711, i_8_1712, i_8_1716, i_8_1721, i_8_1730, i_8_1746, i_8_1752, i_8_1783, i_8_1811, i_8_1819, i_8_1822, i_8_1823, i_8_1855, i_8_1963, i_8_1972, i_8_1999, i_8_2000, i_8_2107, i_8_2139, i_8_2144, i_8_2147, i_8_2215, i_8_2243, i_8_2255, i_8_2289, i_8_2293, o_8_314);
	kernel_8_315 k_8_315(i_8_10, i_8_38, i_8_49, i_8_82, i_8_93, i_8_111, i_8_181, i_8_216, i_8_217, i_8_315, i_8_316, i_8_317, i_8_324, i_8_325, i_8_360, i_8_397, i_8_416, i_8_505, i_8_522, i_8_523, i_8_550, i_8_576, i_8_577, i_8_595, i_8_603, i_8_604, i_8_640, i_8_653, i_8_659, i_8_667, i_8_706, i_8_730, i_8_731, i_8_748, i_8_799, i_8_841, i_8_874, i_8_1010, i_8_1036, i_8_1108, i_8_1135, i_8_1136, i_8_1153, i_8_1156, i_8_1233, i_8_1234, i_8_1243, i_8_1244, i_8_1260, i_8_1269, i_8_1278, i_8_1296, i_8_1297, i_8_1324, i_8_1333, i_8_1360, i_8_1363, i_8_1388, i_8_1407, i_8_1423, i_8_1431, i_8_1450, i_8_1455, i_8_1459, i_8_1462, i_8_1468, i_8_1470, i_8_1471, i_8_1476, i_8_1489, i_8_1512, i_8_1513, i_8_1522, i_8_1523, i_8_1544, i_8_1594, i_8_1604, i_8_1675, i_8_1684, i_8_1693, i_8_1710, i_8_1774, i_8_1822, i_8_1837, i_8_1881, i_8_1888, i_8_1936, i_8_1971, i_8_1972, i_8_1990, i_8_1992, i_8_2043, i_8_2104, i_8_2133, i_8_2169, i_8_2187, i_8_2259, i_8_2260, i_8_2287, i_8_2291, o_8_315);
	kernel_8_316 k_8_316(i_8_30, i_8_31, i_8_37, i_8_82, i_8_84, i_8_114, i_8_115, i_8_128, i_8_136, i_8_143, i_8_150, i_8_194, i_8_247, i_8_382, i_8_383, i_8_386, i_8_389, i_8_391, i_8_398, i_8_419, i_8_433, i_8_491, i_8_496, i_8_497, i_8_517, i_8_556, i_8_605, i_8_607, i_8_614, i_8_631, i_8_634, i_8_638, i_8_661, i_8_747, i_8_786, i_8_842, i_8_850, i_8_858, i_8_931, i_8_940, i_8_959, i_8_964, i_8_1072, i_8_1082, i_8_1125, i_8_1135, i_8_1228, i_8_1237, i_8_1262, i_8_1264, i_8_1274, i_8_1304, i_8_1309, i_8_1355, i_8_1388, i_8_1400, i_8_1434, i_8_1435, i_8_1462, i_8_1509, i_8_1522, i_8_1525, i_8_1531, i_8_1642, i_8_1647, i_8_1667, i_8_1675, i_8_1697, i_8_1702, i_8_1717, i_8_1747, i_8_1760, i_8_1766, i_8_1792, i_8_1805, i_8_1808, i_8_1823, i_8_1826, i_8_1865, i_8_1866, i_8_1918, i_8_1948, i_8_1972, i_8_1997, i_8_2060, i_8_2110, i_8_2134, i_8_2138, i_8_2141, i_8_2144, i_8_2154, i_8_2155, i_8_2170, i_8_2209, i_8_2215, i_8_2218, i_8_2255, i_8_2281, i_8_2286, i_8_2298, o_8_316);
	kernel_8_317 k_8_317(i_8_22, i_8_165, i_8_208, i_8_262, i_8_264, i_8_265, i_8_279, i_8_282, i_8_285, i_8_292, i_8_295, i_8_310, i_8_319, i_8_321, i_8_397, i_8_436, i_8_439, i_8_450, i_8_525, i_8_526, i_8_639, i_8_706, i_8_727, i_8_747, i_8_807, i_8_808, i_8_883, i_8_966, i_8_969, i_8_1035, i_8_1182, i_8_1191, i_8_1198, i_8_1227, i_8_1236, i_8_1264, i_8_1267, i_8_1290, i_8_1305, i_8_1310, i_8_1351, i_8_1354, i_8_1357, i_8_1359, i_8_1362, i_8_1365, i_8_1398, i_8_1440, i_8_1446, i_8_1456, i_8_1468, i_8_1470, i_8_1474, i_8_1489, i_8_1491, i_8_1524, i_8_1533, i_8_1536, i_8_1547, i_8_1560, i_8_1570, i_8_1627, i_8_1641, i_8_1645, i_8_1649, i_8_1674, i_8_1677, i_8_1678, i_8_1695, i_8_1696, i_8_1704, i_8_1713, i_8_1767, i_8_1780, i_8_1789, i_8_1791, i_8_1820, i_8_1822, i_8_1826, i_8_1836, i_8_1861, i_8_1876, i_8_1956, i_8_1987, i_8_1995, i_8_2028, i_8_2056, i_8_2112, i_8_2133, i_8_2136, i_8_2149, i_8_2154, i_8_2164, i_8_2172, i_8_2190, i_8_2193, i_8_2194, i_8_2228, i_8_2248, i_8_2260, o_8_317);
	kernel_8_318 k_8_318(i_8_27, i_8_33, i_8_34, i_8_54, i_8_84, i_8_96, i_8_106, i_8_156, i_8_157, i_8_201, i_8_202, i_8_219, i_8_246, i_8_265, i_8_274, i_8_292, i_8_324, i_8_325, i_8_360, i_8_383, i_8_440, i_8_445, i_8_475, i_8_484, i_8_498, i_8_508, i_8_523, i_8_546, i_8_552, i_8_556, i_8_591, i_8_606, i_8_625, i_8_627, i_8_657, i_8_658, i_8_660, i_8_661, i_8_676, i_8_714, i_8_723, i_8_757, i_8_759, i_8_760, i_8_768, i_8_795, i_8_822, i_8_823, i_8_837, i_8_840, i_8_895, i_8_949, i_8_1050, i_8_1087, i_8_1107, i_8_1113, i_8_1114, i_8_1130, i_8_1134, i_8_1135, i_8_1155, i_8_1267, i_8_1305, i_8_1320, i_8_1346, i_8_1387, i_8_1408, i_8_1420, i_8_1470, i_8_1480, i_8_1524, i_8_1525, i_8_1551, i_8_1579, i_8_1589, i_8_1606, i_8_1629, i_8_1705, i_8_1716, i_8_1746, i_8_1781, i_8_1805, i_8_1809, i_8_1839, i_8_1858, i_8_1859, i_8_1902, i_8_1966, i_8_2001, i_8_2011, i_8_2028, i_8_2031, i_8_2043, i_8_2049, i_8_2127, i_8_2146, i_8_2187, i_8_2188, i_8_2263, i_8_2286, o_8_318);
	kernel_8_319 k_8_319(i_8_34, i_8_80, i_8_85, i_8_125, i_8_139, i_8_142, i_8_151, i_8_194, i_8_197, i_8_230, i_8_365, i_8_373, i_8_427, i_8_430, i_8_454, i_8_490, i_8_491, i_8_538, i_8_556, i_8_584, i_8_605, i_8_616, i_8_628, i_8_629, i_8_662, i_8_665, i_8_677, i_8_694, i_8_696, i_8_697, i_8_698, i_8_725, i_8_731, i_8_736, i_8_755, i_8_782, i_8_784, i_8_808, i_8_838, i_8_842, i_8_843, i_8_844, i_8_845, i_8_869, i_8_952, i_8_989, i_8_995, i_8_1139, i_8_1142, i_8_1151, i_8_1241, i_8_1260, i_8_1283, i_8_1301, i_8_1331, i_8_1355, i_8_1376, i_8_1388, i_8_1411, i_8_1412, i_8_1450, i_8_1472, i_8_1483, i_8_1484, i_8_1529, i_8_1615, i_8_1664, i_8_1691, i_8_1701, i_8_1709, i_8_1732, i_8_1751, i_8_1771, i_8_1823, i_8_1825, i_8_1846, i_8_1858, i_8_1859, i_8_1886, i_8_1904, i_8_1961, i_8_1966, i_8_1990, i_8_1997, i_8_2012, i_8_2015, i_8_2060, i_8_2075, i_8_2087, i_8_2096, i_8_2129, i_8_2148, i_8_2153, i_8_2174, i_8_2176, i_8_2177, i_8_2236, i_8_2263, i_8_2275, i_8_2289, o_8_319);
	kernel_8_320 k_8_320(i_8_31, i_8_50, i_8_57, i_8_60, i_8_75, i_8_101, i_8_131, i_8_168, i_8_190, i_8_301, i_8_311, i_8_322, i_8_356, i_8_361, i_8_371, i_8_384, i_8_427, i_8_455, i_8_461, i_8_538, i_8_539, i_8_548, i_8_553, i_8_581, i_8_582, i_8_608, i_8_613, i_8_638, i_8_644, i_8_653, i_8_655, i_8_664, i_8_683, i_8_695, i_8_701, i_8_745, i_8_752, i_8_755, i_8_779, i_8_781, i_8_820, i_8_827, i_8_884, i_8_886, i_8_944, i_8_955, i_8_1006, i_8_1039, i_8_1127, i_8_1226, i_8_1246, i_8_1247, i_8_1267, i_8_1268, i_8_1282, i_8_1283, i_8_1301, i_8_1302, i_8_1303, i_8_1339, i_8_1350, i_8_1353, i_8_1432, i_8_1455, i_8_1603, i_8_1607, i_8_1608, i_8_1633, i_8_1668, i_8_1699, i_8_1709, i_8_1718, i_8_1737, i_8_1759, i_8_1768, i_8_1777, i_8_1780, i_8_1789, i_8_1807, i_8_1810, i_8_1903, i_8_1904, i_8_1912, i_8_1939, i_8_1973, i_8_1981, i_8_1984, i_8_1992, i_8_2039, i_8_2048, i_8_2107, i_8_2145, i_8_2155, i_8_2156, i_8_2173, i_8_2195, i_8_2249, i_8_2270, i_8_2290, i_8_2294, o_8_320);
	kernel_8_321 k_8_321(i_8_49, i_8_51, i_8_52, i_8_70, i_8_132, i_8_159, i_8_168, i_8_177, i_8_191, i_8_213, i_8_214, i_8_215, i_8_273, i_8_285, i_8_292, i_8_294, i_8_300, i_8_303, i_8_304, i_8_328, i_8_339, i_8_340, i_8_357, i_8_382, i_8_429, i_8_431, i_8_456, i_8_501, i_8_528, i_8_552, i_8_592, i_8_606, i_8_607, i_8_610, i_8_615, i_8_638, i_8_646, i_8_660, i_8_707, i_8_753, i_8_754, i_8_768, i_8_771, i_8_772, i_8_881, i_8_924, i_8_925, i_8_933, i_8_991, i_8_1093, i_8_1158, i_8_1159, i_8_1176, i_8_1195, i_8_1230, i_8_1267, i_8_1299, i_8_1313, i_8_1338, i_8_1347, i_8_1385, i_8_1410, i_8_1422, i_8_1489, i_8_1493, i_8_1528, i_8_1534, i_8_1553, i_8_1649, i_8_1671, i_8_1687, i_8_1731, i_8_1735, i_8_1770, i_8_1771, i_8_1818, i_8_1823, i_8_1824, i_8_1826, i_8_1831, i_8_1863, i_8_1885, i_8_1995, i_8_2004, i_8_2005, i_8_2022, i_8_2038, i_8_2074, i_8_2130, i_8_2153, i_8_2155, i_8_2157, i_8_2182, i_8_2184, i_8_2202, i_8_2211, i_8_2212, i_8_2229, i_8_2263, i_8_2292, o_8_321);
	kernel_8_322 k_8_322(i_8_1, i_8_31, i_8_34, i_8_54, i_8_55, i_8_58, i_8_93, i_8_94, i_8_138, i_8_169, i_8_220, i_8_241, i_8_255, i_8_256, i_8_265, i_8_292, i_8_360, i_8_362, i_8_363, i_8_381, i_8_382, i_8_442, i_8_458, i_8_489, i_8_499, i_8_523, i_8_547, i_8_594, i_8_625, i_8_633, i_8_657, i_8_706, i_8_732, i_8_736, i_8_751, i_8_786, i_8_805, i_8_811, i_8_838, i_8_840, i_8_871, i_8_873, i_8_958, i_8_976, i_8_995, i_8_1071, i_8_1074, i_8_1182, i_8_1225, i_8_1240, i_8_1347, i_8_1360, i_8_1387, i_8_1403, i_8_1453, i_8_1471, i_8_1506, i_8_1524, i_8_1579, i_8_1615, i_8_1621, i_8_1630, i_8_1678, i_8_1681, i_8_1734, i_8_1743, i_8_1749, i_8_1750, i_8_1759, i_8_1760, i_8_1765, i_8_1768, i_8_1774, i_8_1777, i_8_1790, i_8_1821, i_8_1848, i_8_1849, i_8_1856, i_8_1857, i_8_1858, i_8_1902, i_8_1903, i_8_1946, i_8_1984, i_8_1995, i_8_2028, i_8_2029, i_8_2031, i_8_2092, i_8_2098, i_8_2119, i_8_2128, i_8_2129, i_8_2133, i_8_2134, i_8_2232, i_8_2245, i_8_2248, i_8_2259, o_8_322);
	kernel_8_323 k_8_323(i_8_85, i_8_88, i_8_121, i_8_193, i_8_222, i_8_223, i_8_266, i_8_272, i_8_288, i_8_345, i_8_348, i_8_374, i_8_391, i_8_419, i_8_424, i_8_426, i_8_427, i_8_444, i_8_451, i_8_457, i_8_491, i_8_526, i_8_589, i_8_590, i_8_595, i_8_599, i_8_625, i_8_649, i_8_652, i_8_666, i_8_679, i_8_685, i_8_709, i_8_715, i_8_761, i_8_798, i_8_815, i_8_820, i_8_838, i_8_847, i_8_909, i_8_996, i_8_1040, i_8_1047, i_8_1048, i_8_1084, i_8_1139, i_8_1141, i_8_1219, i_8_1228, i_8_1264, i_8_1269, i_8_1280, i_8_1309, i_8_1360, i_8_1373, i_8_1398, i_8_1407, i_8_1426, i_8_1440, i_8_1473, i_8_1498, i_8_1535, i_8_1544, i_8_1555, i_8_1638, i_8_1651, i_8_1680, i_8_1681, i_8_1731, i_8_1741, i_8_1761, i_8_1804, i_8_1810, i_8_1857, i_8_1883, i_8_1885, i_8_1930, i_8_1948, i_8_1959, i_8_1980, i_8_1993, i_8_2025, i_8_2059, i_8_2066, i_8_2106, i_8_2111, i_8_2134, i_8_2150, i_8_2152, i_8_2172, i_8_2221, i_8_2227, i_8_2235, i_8_2245, i_8_2258, i_8_2263, i_8_2273, i_8_2275, i_8_2281, o_8_323);
	kernel_8_324 k_8_324(i_8_6, i_8_11, i_8_14, i_8_43, i_8_61, i_8_78, i_8_79, i_8_80, i_8_85, i_8_87, i_8_105, i_8_106, i_8_124, i_8_141, i_8_142, i_8_258, i_8_268, i_8_285, i_8_294, i_8_295, i_8_309, i_8_336, i_8_339, i_8_345, i_8_364, i_8_370, i_8_525, i_8_529, i_8_555, i_8_564, i_8_595, i_8_598, i_8_601, i_8_608, i_8_609, i_8_624, i_8_634, i_8_642, i_8_645, i_8_654, i_8_660, i_8_664, i_8_688, i_8_708, i_8_718, i_8_726, i_8_753, i_8_768, i_8_783, i_8_789, i_8_825, i_8_834, i_8_835, i_8_840, i_8_853, i_8_870, i_8_939, i_8_950, i_8_958, i_8_1012, i_8_1116, i_8_1164, i_8_1185, i_8_1213, i_8_1299, i_8_1309, i_8_1317, i_8_1330, i_8_1357, i_8_1375, i_8_1380, i_8_1409, i_8_1437, i_8_1438, i_8_1446, i_8_1473, i_8_1542, i_8_1546, i_8_1565, i_8_1588, i_8_1590, i_8_1600, i_8_1734, i_8_1779, i_8_1857, i_8_1861, i_8_1905, i_8_1906, i_8_2034, i_8_2037, i_8_2049, i_8_2073, i_8_2085, i_8_2090, i_8_2121, i_8_2172, i_8_2191, i_8_2193, i_8_2235, i_8_2268, o_8_324);
	kernel_8_325 k_8_325(i_8_41, i_8_65, i_8_82, i_8_91, i_8_92, i_8_128, i_8_131, i_8_136, i_8_137, i_8_140, i_8_142, i_8_163, i_8_181, i_8_189, i_8_212, i_8_236, i_8_282, i_8_307, i_8_308, i_8_316, i_8_335, i_8_344, i_8_380, i_8_446, i_8_451, i_8_452, i_8_486, i_8_491, i_8_527, i_8_542, i_8_553, i_8_554, i_8_595, i_8_604, i_8_614, i_8_622, i_8_652, i_8_661, i_8_686, i_8_696, i_8_700, i_8_703, i_8_730, i_8_731, i_8_792, i_8_837, i_8_838, i_8_841, i_8_852, i_8_878, i_8_929, i_8_932, i_8_956, i_8_965, i_8_973, i_8_1018, i_8_1035, i_8_1061, i_8_1115, i_8_1271, i_8_1283, i_8_1297, i_8_1315, i_8_1325, i_8_1328, i_8_1367, i_8_1373, i_8_1449, i_8_1621, i_8_1622, i_8_1639, i_8_1682, i_8_1686, i_8_1707, i_8_1715, i_8_1729, i_8_1733, i_8_1744, i_8_1760, i_8_1764, i_8_1828, i_8_1838, i_8_1882, i_8_1900, i_8_1937, i_8_1949, i_8_2017, i_8_2020, i_8_2108, i_8_2110, i_8_2144, i_8_2146, i_8_2153, i_8_2180, i_8_2198, i_8_2206, i_8_2212, i_8_2246, i_8_2264, i_8_2270, o_8_325);
	kernel_8_326 k_8_326(i_8_21, i_8_22, i_8_32, i_8_73, i_8_103, i_8_148, i_8_150, i_8_190, i_8_202, i_8_247, i_8_275, i_8_355, i_8_365, i_8_373, i_8_382, i_8_383, i_8_386, i_8_426, i_8_445, i_8_469, i_8_490, i_8_499, i_8_517, i_8_652, i_8_704, i_8_733, i_8_751, i_8_752, i_8_777, i_8_814, i_8_832, i_8_837, i_8_846, i_8_913, i_8_941, i_8_967, i_8_1069, i_8_1072, i_8_1112, i_8_1174, i_8_1202, i_8_1224, i_8_1233, i_8_1264, i_8_1284, i_8_1350, i_8_1394, i_8_1399, i_8_1404, i_8_1452, i_8_1479, i_8_1497, i_8_1531, i_8_1552, i_8_1597, i_8_1625, i_8_1648, i_8_1649, i_8_1657, i_8_1660, i_8_1676, i_8_1677, i_8_1705, i_8_1746, i_8_1792, i_8_1805, i_8_1806, i_8_1808, i_8_1812, i_8_1821, i_8_1840, i_8_1848, i_8_1849, i_8_1850, i_8_1864, i_8_1866, i_8_1890, i_8_1917, i_8_1928, i_8_1951, i_8_1952, i_8_1966, i_8_1972, i_8_1989, i_8_1997, i_8_2011, i_8_2038, i_8_2088, i_8_2089, i_8_2145, i_8_2146, i_8_2148, i_8_2149, i_8_2150, i_8_2155, i_8_2224, i_8_2233, i_8_2257, i_8_2273, i_8_2299, o_8_326);
	kernel_8_327 k_8_327(i_8_34, i_8_54, i_8_55, i_8_86, i_8_87, i_8_96, i_8_103, i_8_142, i_8_167, i_8_201, i_8_202, i_8_223, i_8_255, i_8_369, i_8_415, i_8_421, i_8_441, i_8_456, i_8_471, i_8_479, i_8_500, i_8_526, i_8_528, i_8_530, i_8_552, i_8_553, i_8_601, i_8_625, i_8_660, i_8_714, i_8_772, i_8_795, i_8_815, i_8_827, i_8_868, i_8_888, i_8_895, i_8_1012, i_8_1028, i_8_1051, i_8_1059, i_8_1061, i_8_1084, i_8_1112, i_8_1156, i_8_1188, i_8_1198, i_8_1215, i_8_1249, i_8_1259, i_8_1266, i_8_1274, i_8_1277, i_8_1281, i_8_1325, i_8_1390, i_8_1417, i_8_1435, i_8_1438, i_8_1449, i_8_1471, i_8_1480, i_8_1536, i_8_1549, i_8_1551, i_8_1552, i_8_1579, i_8_1627, i_8_1629, i_8_1633, i_8_1668, i_8_1675, i_8_1681, i_8_1682, i_8_1707, i_8_1726, i_8_1731, i_8_1732, i_8_1744, i_8_1749, i_8_1753, i_8_1758, i_8_1813, i_8_1855, i_8_1858, i_8_1872, i_8_1873, i_8_1889, i_8_1894, i_8_1902, i_8_2002, i_8_2074, i_8_2136, i_8_2154, i_8_2191, i_8_2212, i_8_2228, i_8_2259, i_8_2271, i_8_2272, o_8_327);
	kernel_8_328 k_8_328(i_8_22, i_8_64, i_8_67, i_8_94, i_8_114, i_8_193, i_8_194, i_8_226, i_8_275, i_8_283, i_8_297, i_8_361, i_8_382, i_8_391, i_8_416, i_8_426, i_8_484, i_8_492, i_8_493, i_8_505, i_8_518, i_8_535, i_8_546, i_8_567, i_8_631, i_8_635, i_8_652, i_8_660, i_8_691, i_8_693, i_8_709, i_8_739, i_8_750, i_8_751, i_8_814, i_8_815, i_8_837, i_8_851, i_8_865, i_8_904, i_8_964, i_8_970, i_8_1012, i_8_1033, i_8_1072, i_8_1102, i_8_1134, i_8_1135, i_8_1171, i_8_1192, i_8_1202, i_8_1229, i_8_1249, i_8_1278, i_8_1282, i_8_1283, i_8_1286, i_8_1306, i_8_1391, i_8_1397, i_8_1439, i_8_1450, i_8_1477, i_8_1478, i_8_1489, i_8_1526, i_8_1546, i_8_1552, i_8_1582, i_8_1606, i_8_1640, i_8_1660, i_8_1673, i_8_1704, i_8_1769, i_8_1784, i_8_1819, i_8_1840, i_8_1849, i_8_1885, i_8_1902, i_8_1957, i_8_1981, i_8_1997, i_8_2011, i_8_2014, i_8_2145, i_8_2149, i_8_2171, i_8_2174, i_8_2214, i_8_2216, i_8_2242, i_8_2245, i_8_2255, i_8_2258, i_8_2262, i_8_2289, i_8_2300, i_8_2303, o_8_328);
	kernel_8_329 k_8_329(i_8_22, i_8_23, i_8_28, i_8_29, i_8_56, i_8_67, i_8_74, i_8_79, i_8_162, i_8_172, i_8_181, i_8_191, i_8_193, i_8_198, i_8_218, i_8_226, i_8_227, i_8_229, i_8_231, i_8_299, i_8_302, i_8_370, i_8_379, i_8_383, i_8_414, i_8_415, i_8_424, i_8_434, i_8_463, i_8_488, i_8_492, i_8_493, i_8_592, i_8_604, i_8_605, i_8_658, i_8_679, i_8_823, i_8_837, i_8_838, i_8_839, i_8_842, i_8_859, i_8_869, i_8_873, i_8_883, i_8_955, i_8_965, i_8_971, i_8_1041, i_8_1104, i_8_1129, i_8_1175, i_8_1189, i_8_1237, i_8_1279, i_8_1297, i_8_1307, i_8_1328, i_8_1341, i_8_1360, i_8_1382, i_8_1441, i_8_1471, i_8_1472, i_8_1564, i_8_1573, i_8_1585, i_8_1603, i_8_1604, i_8_1622, i_8_1634, i_8_1652, i_8_1688, i_8_1756, i_8_1774, i_8_1775, i_8_1805, i_8_1809, i_8_1843, i_8_1873, i_8_1874, i_8_1882, i_8_1909, i_8_1982, i_8_1989, i_8_1991, i_8_1995, i_8_2052, i_8_2054, i_8_2065, i_8_2140, i_8_2145, i_8_2170, i_8_2171, i_8_2214, i_8_2215, i_8_2216, i_8_2233, i_8_2243, o_8_329);
	kernel_8_330 k_8_330(i_8_58, i_8_104, i_8_106, i_8_107, i_8_110, i_8_163, i_8_256, i_8_257, i_8_346, i_8_368, i_8_377, i_8_378, i_8_384, i_8_385, i_8_396, i_8_398, i_8_451, i_8_453, i_8_493, i_8_580, i_8_601, i_8_642, i_8_648, i_8_702, i_8_732, i_8_748, i_8_751, i_8_752, i_8_847, i_8_868, i_8_965, i_8_1058, i_8_1134, i_8_1135, i_8_1137, i_8_1138, i_8_1153, i_8_1192, i_8_1228, i_8_1233, i_8_1234, i_8_1273, i_8_1274, i_8_1314, i_8_1319, i_8_1324, i_8_1326, i_8_1328, i_8_1353, i_8_1408, i_8_1440, i_8_1486, i_8_1490, i_8_1506, i_8_1507, i_8_1533, i_8_1534, i_8_1551, i_8_1613, i_8_1614, i_8_1615, i_8_1616, i_8_1630, i_8_1652, i_8_1686, i_8_1688, i_8_1691, i_8_1710, i_8_1711, i_8_1712, i_8_1713, i_8_1714, i_8_1715, i_8_1810, i_8_1811, i_8_1812, i_8_1813, i_8_1831, i_8_1836, i_8_1837, i_8_1838, i_8_1839, i_8_1840, i_8_1841, i_8_1862, i_8_1885, i_8_1894, i_8_1895, i_8_1939, i_8_1986, i_8_2093, i_8_2099, i_8_2133, i_8_2134, i_8_2171, i_8_2260, i_8_2262, i_8_2263, i_8_2264, i_8_2298, o_8_330);
	kernel_8_331 k_8_331(i_8_48, i_8_63, i_8_64, i_8_121, i_8_152, i_8_171, i_8_219, i_8_226, i_8_294, i_8_295, i_8_304, i_8_324, i_8_340, i_8_354, i_8_374, i_8_382, i_8_384, i_8_385, i_8_430, i_8_489, i_8_492, i_8_552, i_8_554, i_8_583, i_8_591, i_8_592, i_8_600, i_8_642, i_8_655, i_8_661, i_8_662, i_8_687, i_8_710, i_8_733, i_8_750, i_8_795, i_8_798, i_8_879, i_8_881, i_8_926, i_8_935, i_8_990, i_8_1032, i_8_1110, i_8_1152, i_8_1170, i_8_1188, i_8_1224, i_8_1257, i_8_1258, i_8_1259, i_8_1266, i_8_1267, i_8_1272, i_8_1276, i_8_1284, i_8_1285, i_8_1286, i_8_1330, i_8_1371, i_8_1375, i_8_1389, i_8_1443, i_8_1455, i_8_1552, i_8_1554, i_8_1607, i_8_1633, i_8_1635, i_8_1647, i_8_1653, i_8_1678, i_8_1686, i_8_1723, i_8_1730, i_8_1736, i_8_1747, i_8_1751, i_8_1777, i_8_1778, i_8_1869, i_8_1950, i_8_2013, i_8_2048, i_8_2056, i_8_2078, i_8_2095, i_8_2097, i_8_2112, i_8_2114, i_8_2131, i_8_2142, i_8_2157, i_8_2176, i_8_2185, i_8_2194, i_8_2222, i_8_2223, i_8_2249, i_8_2266, o_8_331);
	kernel_8_332 k_8_332(i_8_12, i_8_30, i_8_72, i_8_82, i_8_83, i_8_119, i_8_135, i_8_139, i_8_153, i_8_156, i_8_201, i_8_202, i_8_207, i_8_216, i_8_219, i_8_220, i_8_267, i_8_282, i_8_324, i_8_333, i_8_343, i_8_373, i_8_384, i_8_432, i_8_495, i_8_498, i_8_533, i_8_550, i_8_552, i_8_585, i_8_595, i_8_609, i_8_612, i_8_621, i_8_636, i_8_637, i_8_669, i_8_720, i_8_774, i_8_775, i_8_777, i_8_804, i_8_821, i_8_823, i_8_847, i_8_867, i_8_875, i_8_876, i_8_891, i_8_932, i_8_963, i_8_965, i_8_972, i_8_981, i_8_991, i_8_994, i_8_1008, i_8_1009, i_8_1011, i_8_1083, i_8_1129, i_8_1145, i_8_1155, i_8_1171, i_8_1245, i_8_1255, i_8_1270, i_8_1275, i_8_1288, i_8_1296, i_8_1312, i_8_1341, i_8_1342, i_8_1428, i_8_1432, i_8_1443, i_8_1516, i_8_1521, i_8_1524, i_8_1548, i_8_1549, i_8_1611, i_8_1669, i_8_1675, i_8_1705, i_8_1775, i_8_1800, i_8_1801, i_8_1839, i_8_1919, i_8_1945, i_8_1999, i_8_2038, i_8_2107, i_8_2117, i_8_2146, i_8_2269, i_8_2281, i_8_2286, i_8_2291, o_8_332);
	kernel_8_333 k_8_333(i_8_34, i_8_35, i_8_50, i_8_53, i_8_60, i_8_65, i_8_95, i_8_125, i_8_143, i_8_169, i_8_233, i_8_242, i_8_278, i_8_347, i_8_350, i_8_360, i_8_365, i_8_401, i_8_431, i_8_454, i_8_455, i_8_553, i_8_557, i_8_581, i_8_590, i_8_607, i_8_613, i_8_614, i_8_638, i_8_656, i_8_661, i_8_662, i_8_679, i_8_680, i_8_697, i_8_700, i_8_701, i_8_707, i_8_711, i_8_731, i_8_759, i_8_779, i_8_782, i_8_793, i_8_799, i_8_844, i_8_969, i_8_1030, i_8_1103, i_8_1129, i_8_1146, i_8_1154, i_8_1157, i_8_1172, i_8_1175, i_8_1264, i_8_1265, i_8_1274, i_8_1292, i_8_1305, i_8_1373, i_8_1411, i_8_1412, i_8_1472, i_8_1493, i_8_1508, i_8_1525, i_8_1562, i_8_1607, i_8_1609, i_8_1628, i_8_1648, i_8_1649, i_8_1655, i_8_1664, i_8_1679, i_8_1698, i_8_1778, i_8_1803, i_8_1819, i_8_1823, i_8_1832, i_8_1854, i_8_1859, i_8_1886, i_8_1906, i_8_1967, i_8_1984, i_8_1985, i_8_1996, i_8_2018, i_8_2096, i_8_2146, i_8_2156, i_8_2183, i_8_2210, i_8_2219, i_8_2227, i_8_2244, i_8_2276, o_8_333);
	kernel_8_334 k_8_334(i_8_53, i_8_86, i_8_87, i_8_97, i_8_139, i_8_230, i_8_255, i_8_258, i_8_260, i_8_327, i_8_328, i_8_329, i_8_362, i_8_363, i_8_457, i_8_462, i_8_463, i_8_464, i_8_466, i_8_474, i_8_476, i_8_500, i_8_523, i_8_526, i_8_528, i_8_530, i_8_555, i_8_617, i_8_660, i_8_661, i_8_663, i_8_672, i_8_674, i_8_682, i_8_732, i_8_762, i_8_763, i_8_840, i_8_841, i_8_842, i_8_845, i_8_958, i_8_977, i_8_996, i_8_997, i_8_1052, i_8_1086, i_8_1113, i_8_1114, i_8_1133, i_8_1139, i_8_1156, i_8_1326, i_8_1327, i_8_1410, i_8_1527, i_8_1528, i_8_1535, i_8_1596, i_8_1598, i_8_1599, i_8_1600, i_8_1645, i_8_1654, i_8_1669, i_8_1762, i_8_1768, i_8_1771, i_8_1788, i_8_1802, i_8_1806, i_8_1807, i_8_1808, i_8_1867, i_8_1868, i_8_1870, i_8_1902, i_8_1903, i_8_1904, i_8_1918, i_8_1919, i_8_1921, i_8_1922, i_8_1949, i_8_1950, i_8_1952, i_8_1965, i_8_1969, i_8_1980, i_8_1983, i_8_2064, i_8_2118, i_8_2120, i_8_2121, i_8_2214, i_8_2216, i_8_2218, i_8_2219, i_8_2245, i_8_2267, o_8_334);
	kernel_8_335 k_8_335(i_8_34, i_8_53, i_8_80, i_8_115, i_8_143, i_8_189, i_8_190, i_8_191, i_8_193, i_8_252, i_8_292, i_8_301, i_8_302, i_8_305, i_8_345, i_8_346, i_8_362, i_8_378, i_8_379, i_8_380, i_8_381, i_8_383, i_8_463, i_8_468, i_8_469, i_8_492, i_8_522, i_8_550, i_8_591, i_8_606, i_8_607, i_8_608, i_8_610, i_8_611, i_8_627, i_8_663, i_8_664, i_8_689, i_8_712, i_8_726, i_8_735, i_8_764, i_8_834, i_8_989, i_8_997, i_8_998, i_8_1086, i_8_1111, i_8_1112, i_8_1125, i_8_1235, i_8_1261, i_8_1273, i_8_1274, i_8_1286, i_8_1306, i_8_1410, i_8_1435, i_8_1436, i_8_1470, i_8_1471, i_8_1528, i_8_1529, i_8_1533, i_8_1537, i_8_1605, i_8_1617, i_8_1624, i_8_1660, i_8_1680, i_8_1681, i_8_1751, i_8_1758, i_8_1803, i_8_1804, i_8_1824, i_8_1863, i_8_1865, i_8_1887, i_8_1984, i_8_1991, i_8_1992, i_8_1996, i_8_2034, i_8_2073, i_8_2109, i_8_2139, i_8_2140, i_8_2141, i_8_2149, i_8_2151, i_8_2153, i_8_2154, i_8_2155, i_8_2156, i_8_2157, i_8_2214, i_8_2215, i_8_2216, i_8_2275, o_8_335);
	kernel_8_336 k_8_336(i_8_11, i_8_19, i_8_27, i_8_34, i_8_73, i_8_74, i_8_83, i_8_101, i_8_141, i_8_298, i_8_325, i_8_326, i_8_364, i_8_367, i_8_450, i_8_486, i_8_562, i_8_577, i_8_579, i_8_589, i_8_611, i_8_639, i_8_640, i_8_657, i_8_663, i_8_676, i_8_684, i_8_694, i_8_707, i_8_708, i_8_712, i_8_713, i_8_721, i_8_729, i_8_733, i_8_791, i_8_822, i_8_837, i_8_844, i_8_855, i_8_967, i_8_996, i_8_1026, i_8_1129, i_8_1134, i_8_1179, i_8_1183, i_8_1206, i_8_1243, i_8_1252, i_8_1261, i_8_1285, i_8_1286, i_8_1296, i_8_1395, i_8_1398, i_8_1473, i_8_1480, i_8_1507, i_8_1513, i_8_1516, i_8_1530, i_8_1534, i_8_1555, i_8_1563, i_8_1595, i_8_1605, i_8_1625, i_8_1668, i_8_1675, i_8_1680, i_8_1707, i_8_1710, i_8_1711, i_8_1745, i_8_1754, i_8_1756, i_8_1757, i_8_1789, i_8_1802, i_8_1810, i_8_1819, i_8_1826, i_8_1854, i_8_1883, i_8_1900, i_8_1989, i_8_1990, i_8_2011, i_8_2017, i_8_2025, i_8_2088, i_8_2137, i_8_2147, i_8_2152, i_8_2206, i_8_2245, i_8_2246, i_8_2265, i_8_2292, o_8_336);
	kernel_8_337 k_8_337(i_8_5, i_8_20, i_8_49, i_8_64, i_8_83, i_8_89, i_8_101, i_8_257, i_8_263, i_8_275, i_8_290, i_8_301, i_8_303, i_8_366, i_8_367, i_8_368, i_8_380, i_8_382, i_8_401, i_8_434, i_8_440, i_8_452, i_8_455, i_8_476, i_8_486, i_8_491, i_8_506, i_8_518, i_8_528, i_8_547, i_8_586, i_8_590, i_8_626, i_8_632, i_8_634, i_8_658, i_8_670, i_8_671, i_8_694, i_8_703, i_8_706, i_8_716, i_8_803, i_8_824, i_8_830, i_8_839, i_8_844, i_8_845, i_8_877, i_8_1012, i_8_1028, i_8_1130, i_8_1225, i_8_1256, i_8_1286, i_8_1350, i_8_1355, i_8_1388, i_8_1420, i_8_1442, i_8_1445, i_8_1456, i_8_1471, i_8_1531, i_8_1532, i_8_1536, i_8_1537, i_8_1544, i_8_1576, i_8_1585, i_8_1615, i_8_1621, i_8_1622, i_8_1747, i_8_1751, i_8_1753, i_8_1768, i_8_1782, i_8_1802, i_8_1819, i_8_1838, i_8_1846, i_8_1847, i_8_1850, i_8_1892, i_8_1895, i_8_1963, i_8_1964, i_8_1990, i_8_1993, i_8_2000, i_8_2012, i_8_2047, i_8_2063, i_8_2111, i_8_2117, i_8_2141, i_8_2170, i_8_2227, i_8_2237, o_8_337);
	kernel_8_338 k_8_338(i_8_19, i_8_37, i_8_47, i_8_67, i_8_72, i_8_73, i_8_83, i_8_119, i_8_163, i_8_208, i_8_209, i_8_253, i_8_307, i_8_362, i_8_398, i_8_424, i_8_487, i_8_489, i_8_497, i_8_500, i_8_524, i_8_526, i_8_612, i_8_625, i_8_662, i_8_685, i_8_688, i_8_694, i_8_695, i_8_729, i_8_752, i_8_760, i_8_767, i_8_777, i_8_796, i_8_829, i_8_830, i_8_833, i_8_837, i_8_839, i_8_865, i_8_878, i_8_956, i_8_965, i_8_970, i_8_971, i_8_974, i_8_998, i_8_1018, i_8_1057, i_8_1073, i_8_1102, i_8_1171, i_8_1172, i_8_1234, i_8_1235, i_8_1267, i_8_1288, i_8_1289, i_8_1294, i_8_1307, i_8_1378, i_8_1400, i_8_1405, i_8_1453, i_8_1468, i_8_1471, i_8_1555, i_8_1559, i_8_1620, i_8_1639, i_8_1647, i_8_1682, i_8_1712, i_8_1733, i_8_1754, i_8_1760, i_8_1762, i_8_1775, i_8_1792, i_8_1883, i_8_1885, i_8_1928, i_8_1989, i_8_1997, i_8_2053, i_8_2054, i_8_2055, i_8_2107, i_8_2146, i_8_2147, i_8_2148, i_8_2149, i_8_2155, i_8_2162, i_8_2180, i_8_2210, i_8_2224, i_8_2225, i_8_2288, o_8_338);
	kernel_8_339 k_8_339(i_8_138, i_8_146, i_8_148, i_8_189, i_8_227, i_8_229, i_8_273, i_8_302, i_8_359, i_8_366, i_8_392, i_8_432, i_8_455, i_8_464, i_8_470, i_8_475, i_8_490, i_8_503, i_8_512, i_8_529, i_8_551, i_8_583, i_8_592, i_8_595, i_8_610, i_8_614, i_8_637, i_8_656, i_8_679, i_8_718, i_8_751, i_8_812, i_8_819, i_8_827, i_8_860, i_8_863, i_8_866, i_8_874, i_8_914, i_8_917, i_8_985, i_8_1046, i_8_1055, i_8_1058, i_8_1174, i_8_1181, i_8_1188, i_8_1205, i_8_1243, i_8_1298, i_8_1305, i_8_1306, i_8_1311, i_8_1329, i_8_1334, i_8_1343, i_8_1354, i_8_1391, i_8_1410, i_8_1420, i_8_1470, i_8_1471, i_8_1487, i_8_1498, i_8_1502, i_8_1541, i_8_1554, i_8_1559, i_8_1637, i_8_1642, i_8_1647, i_8_1667, i_8_1675, i_8_1676, i_8_1703, i_8_1750, i_8_1751, i_8_1766, i_8_1780, i_8_1784, i_8_1838, i_8_1844, i_8_1919, i_8_1930, i_8_1973, i_8_1989, i_8_1993, i_8_1997, i_8_2000, i_8_2042, i_8_2056, i_8_2065, i_8_2066, i_8_2147, i_8_2191, i_8_2234, i_8_2242, i_8_2248, i_8_2249, i_8_2268, o_8_339);
	kernel_8_340 k_8_340(i_8_10, i_8_18, i_8_28, i_8_49, i_8_73, i_8_135, i_8_156, i_8_183, i_8_229, i_8_252, i_8_265, i_8_288, i_8_370, i_8_387, i_8_421, i_8_435, i_8_472, i_8_473, i_8_493, i_8_507, i_8_543, i_8_546, i_8_550, i_8_595, i_8_608, i_8_611, i_8_625, i_8_633, i_8_660, i_8_661, i_8_663, i_8_684, i_8_687, i_8_690, i_8_711, i_8_756, i_8_765, i_8_769, i_8_781, i_8_783, i_8_786, i_8_806, i_8_819, i_8_820, i_8_822, i_8_847, i_8_865, i_8_873, i_8_891, i_8_892, i_8_946, i_8_975, i_8_984, i_8_1009, i_8_1065, i_8_1107, i_8_1126, i_8_1127, i_8_1144, i_8_1159, i_8_1215, i_8_1245, i_8_1260, i_8_1286, i_8_1305, i_8_1341, i_8_1416, i_8_1417, i_8_1440, i_8_1471, i_8_1549, i_8_1557, i_8_1565, i_8_1629, i_8_1633, i_8_1671, i_8_1674, i_8_1677, i_8_1682, i_8_1702, i_8_1710, i_8_1719, i_8_1737, i_8_1750, i_8_1758, i_8_1783, i_8_1788, i_8_1803, i_8_1808, i_8_1854, i_8_1857, i_8_1861, i_8_1893, i_8_1995, i_8_2025, i_8_2089, i_8_2110, i_8_2181, i_8_2298, i_8_2299, o_8_340);
	kernel_8_341 k_8_341(i_8_27, i_8_45, i_8_49, i_8_82, i_8_111, i_8_162, i_8_190, i_8_216, i_8_217, i_8_220, i_8_223, i_8_229, i_8_237, i_8_253, i_8_257, i_8_325, i_8_361, i_8_363, i_8_364, i_8_388, i_8_414, i_8_425, i_8_436, i_8_451, i_8_452, i_8_461, i_8_493, i_8_570, i_8_571, i_8_607, i_8_608, i_8_631, i_8_661, i_8_687, i_8_694, i_8_732, i_8_735, i_8_756, i_8_758, i_8_767, i_8_803, i_8_811, i_8_840, i_8_841, i_8_842, i_8_856, i_8_876, i_8_919, i_8_936, i_8_937, i_8_938, i_8_991, i_8_995, i_8_996, i_8_1008, i_8_1155, i_8_1179, i_8_1180, i_8_1181, i_8_1182, i_8_1189, i_8_1224, i_8_1234, i_8_1282, i_8_1305, i_8_1333, i_8_1335, i_8_1407, i_8_1467, i_8_1486, i_8_1492, i_8_1493, i_8_1549, i_8_1621, i_8_1631, i_8_1635, i_8_1649, i_8_1674, i_8_1692, i_8_1694, i_8_1730, i_8_1740, i_8_1748, i_8_1758, i_8_1759, i_8_1783, i_8_1797, i_8_1819, i_8_1821, i_8_1822, i_8_1993, i_8_2029, i_8_2054, i_8_2073, i_8_2187, i_8_2245, i_8_2271, i_8_2295, i_8_2296, i_8_2297, o_8_341);
	kernel_8_342 k_8_342(i_8_25, i_8_34, i_8_81, i_8_87, i_8_89, i_8_93, i_8_106, i_8_160, i_8_183, i_8_262, i_8_291, i_8_307, i_8_328, i_8_378, i_8_403, i_8_433, i_8_462, i_8_503, i_8_523, i_8_554, i_8_572, i_8_595, i_8_621, i_8_624, i_8_633, i_8_634, i_8_637, i_8_669, i_8_670, i_8_690, i_8_707, i_8_712, i_8_756, i_8_762, i_8_767, i_8_777, i_8_778, i_8_783, i_8_803, i_8_823, i_8_873, i_8_971, i_8_973, i_8_987, i_8_1026, i_8_1029, i_8_1111, i_8_1119, i_8_1171, i_8_1172, i_8_1219, i_8_1236, i_8_1254, i_8_1282, i_8_1285, i_8_1305, i_8_1314, i_8_1317, i_8_1402, i_8_1424, i_8_1441, i_8_1474, i_8_1476, i_8_1482, i_8_1545, i_8_1547, i_8_1563, i_8_1579, i_8_1585, i_8_1587, i_8_1600, i_8_1651, i_8_1663, i_8_1668, i_8_1671, i_8_1680, i_8_1681, i_8_1695, i_8_1698, i_8_1708, i_8_1746, i_8_1751, i_8_1792, i_8_1804, i_8_1822, i_8_1841, i_8_1902, i_8_1912, i_8_1947, i_8_2107, i_8_2109, i_8_2128, i_8_2136, i_8_2146, i_8_2190, i_8_2226, i_8_2244, i_8_2291, i_8_2292, i_8_2295, o_8_342);
	kernel_8_343 k_8_343(i_8_36, i_8_135, i_8_172, i_8_193, i_8_226, i_8_261, i_8_309, i_8_321, i_8_345, i_8_364, i_8_396, i_8_414, i_8_417, i_8_418, i_8_422, i_8_453, i_8_472, i_8_480, i_8_504, i_8_507, i_8_508, i_8_522, i_8_523, i_8_525, i_8_534, i_8_552, i_8_567, i_8_571, i_8_573, i_8_579, i_8_582, i_8_604, i_8_625, i_8_696, i_8_702, i_8_751, i_8_756, i_8_759, i_8_823, i_8_891, i_8_963, i_8_1009, i_8_1098, i_8_1103, i_8_1128, i_8_1134, i_8_1179, i_8_1197, i_8_1234, i_8_1263, i_8_1266, i_8_1314, i_8_1362, i_8_1422, i_8_1440, i_8_1461, i_8_1464, i_8_1465, i_8_1485, i_8_1512, i_8_1513, i_8_1521, i_8_1522, i_8_1540, i_8_1544, i_8_1569, i_8_1597, i_8_1606, i_8_1629, i_8_1665, i_8_1692, i_8_1693, i_8_1696, i_8_1723, i_8_1765, i_8_1784, i_8_1794, i_8_1803, i_8_1804, i_8_1830, i_8_1836, i_8_1840, i_8_1887, i_8_1899, i_8_1911, i_8_1927, i_8_1935, i_8_1938, i_8_1956, i_8_1974, i_8_1992, i_8_1993, i_8_2070, i_8_2079, i_8_2107, i_8_2141, i_8_2151, i_8_2163, i_8_2208, i_8_2232, o_8_343);
	kernel_8_344 k_8_344(i_8_34, i_8_76, i_8_103, i_8_115, i_8_119, i_8_121, i_8_166, i_8_167, i_8_220, i_8_229, i_8_245, i_8_281, i_8_301, i_8_320, i_8_323, i_8_324, i_8_326, i_8_338, i_8_371, i_8_437, i_8_504, i_8_523, i_8_525, i_8_527, i_8_529, i_8_543, i_8_562, i_8_563, i_8_566, i_8_583, i_8_604, i_8_605, i_8_626, i_8_679, i_8_722, i_8_729, i_8_760, i_8_761, i_8_785, i_8_795, i_8_796, i_8_806, i_8_832, i_8_840, i_8_932, i_8_1049, i_8_1072, i_8_1073, i_8_1109, i_8_1111, i_8_1127, i_8_1154, i_8_1180, i_8_1277, i_8_1282, i_8_1298, i_8_1334, i_8_1346, i_8_1360, i_8_1361, i_8_1364, i_8_1381, i_8_1450, i_8_1454, i_8_1469, i_8_1477, i_8_1478, i_8_1481, i_8_1543, i_8_1544, i_8_1552, i_8_1553, i_8_1684, i_8_1701, i_8_1711, i_8_1733, i_8_1747, i_8_1767, i_8_1768, i_8_1787, i_8_1822, i_8_1846, i_8_1856, i_8_1859, i_8_1864, i_8_1919, i_8_1943, i_8_1975, i_8_1996, i_8_2056, i_8_2074, i_8_2075, i_8_2133, i_8_2141, i_8_2156, i_8_2171, i_8_2192, i_8_2223, i_8_2282, i_8_2296, o_8_344);
	kernel_8_345 k_8_345(i_8_84, i_8_85, i_8_96, i_8_106, i_8_138, i_8_245, i_8_291, i_8_294, i_8_304, i_8_327, i_8_372, i_8_375, i_8_381, i_8_384, i_8_385, i_8_419, i_8_436, i_8_462, i_8_475, i_8_480, i_8_481, i_8_483, i_8_523, i_8_526, i_8_598, i_8_599, i_8_601, i_8_672, i_8_699, i_8_759, i_8_780, i_8_781, i_8_795, i_8_813, i_8_826, i_8_843, i_8_879, i_8_940, i_8_969, i_8_985, i_8_1014, i_8_1032, i_8_1086, i_8_1115, i_8_1119, i_8_1132, i_8_1159, i_8_1218, i_8_1225, i_8_1248, i_8_1257, i_8_1284, i_8_1315, i_8_1327, i_8_1344, i_8_1389, i_8_1506, i_8_1524, i_8_1537, i_8_1542, i_8_1543, i_8_1545, i_8_1551, i_8_1590, i_8_1597, i_8_1606, i_8_1627, i_8_1632, i_8_1633, i_8_1680, i_8_1690, i_8_1698, i_8_1719, i_8_1722, i_8_1741, i_8_1752, i_8_1761, i_8_1803, i_8_1812, i_8_1813, i_8_1840, i_8_1841, i_8_1857, i_8_1866, i_8_1872, i_8_1875, i_8_1921, i_8_1950, i_8_2092, i_8_2110, i_8_2112, i_8_2113, i_8_2127, i_8_2131, i_8_2184, i_8_2185, i_8_2190, i_8_2214, i_8_2215, i_8_2289, o_8_345);
	kernel_8_346 k_8_346(i_8_9, i_8_27, i_8_37, i_8_81, i_8_102, i_8_104, i_8_111, i_8_136, i_8_147, i_8_180, i_8_189, i_8_219, i_8_243, i_8_262, i_8_315, i_8_337, i_8_366, i_8_378, i_8_381, i_8_398, i_8_467, i_8_505, i_8_510, i_8_531, i_8_567, i_8_570, i_8_588, i_8_596, i_8_603, i_8_604, i_8_639, i_8_649, i_8_662, i_8_707, i_8_731, i_8_822, i_8_841, i_8_877, i_8_879, i_8_880, i_8_884, i_8_891, i_8_966, i_8_998, i_8_1008, i_8_1049, i_8_1098, i_8_1108, i_8_1109, i_8_1127, i_8_1140, i_8_1154, i_8_1171, i_8_1231, i_8_1233, i_8_1234, i_8_1276, i_8_1323, i_8_1324, i_8_1351, i_8_1354, i_8_1359, i_8_1404, i_8_1436, i_8_1457, i_8_1458, i_8_1476, i_8_1480, i_8_1491, i_8_1503, i_8_1522, i_8_1567, i_8_1602, i_8_1630, i_8_1683, i_8_1686, i_8_1696, i_8_1758, i_8_1764, i_8_1800, i_8_1810, i_8_1836, i_8_1837, i_8_1882, i_8_1890, i_8_1908, i_8_1936, i_8_1990, i_8_1992, i_8_2037, i_8_2066, i_8_2070, i_8_2071, i_8_2124, i_8_2145, i_8_2234, i_8_2244, i_8_2247, i_8_2269, i_8_2271, o_8_346);
	kernel_8_347 k_8_347(i_8_79, i_8_84, i_8_85, i_8_88, i_8_168, i_8_193, i_8_224, i_8_295, i_8_303, i_8_323, i_8_364, i_8_499, i_8_500, i_8_525, i_8_526, i_8_527, i_8_528, i_8_529, i_8_530, i_8_591, i_8_592, i_8_593, i_8_606, i_8_629, i_8_634, i_8_660, i_8_665, i_8_670, i_8_678, i_8_679, i_8_682, i_8_683, i_8_707, i_8_708, i_8_763, i_8_807, i_8_813, i_8_842, i_8_964, i_8_1057, i_8_1058, i_8_1076, i_8_1192, i_8_1193, i_8_1266, i_8_1268, i_8_1272, i_8_1274, i_8_1299, i_8_1309, i_8_1339, i_8_1340, i_8_1353, i_8_1354, i_8_1390, i_8_1433, i_8_1437, i_8_1455, i_8_1485, i_8_1534, i_8_1536, i_8_1627, i_8_1632, i_8_1633, i_8_1634, i_8_1642, i_8_1732, i_8_1750, i_8_1752, i_8_1770, i_8_1771, i_8_1778, i_8_1783, i_8_1784, i_8_1785, i_8_1787, i_8_1789, i_8_1790, i_8_1822, i_8_1858, i_8_1859, i_8_1860, i_8_1861, i_8_1862, i_8_1866, i_8_1869, i_8_1905, i_8_1906, i_8_1975, i_8_1978, i_8_1996, i_8_2041, i_8_2136, i_8_2137, i_8_2214, i_8_2215, i_8_2226, i_8_2248, i_8_2249, i_8_2284, o_8_347);
	kernel_8_348 k_8_348(i_8_32, i_8_58, i_8_84, i_8_85, i_8_92, i_8_94, i_8_101, i_8_103, i_8_140, i_8_155, i_8_185, i_8_299, i_8_372, i_8_373, i_8_380, i_8_419, i_8_437, i_8_441, i_8_460, i_8_461, i_8_482, i_8_522, i_8_529, i_8_572, i_8_587, i_8_613, i_8_622, i_8_623, i_8_667, i_8_668, i_8_697, i_8_713, i_8_715, i_8_716, i_8_722, i_8_731, i_8_756, i_8_757, i_8_767, i_8_779, i_8_793, i_8_821, i_8_842, i_8_866, i_8_1010, i_8_1028, i_8_1043, i_8_1135, i_8_1153, i_8_1154, i_8_1157, i_8_1253, i_8_1279, i_8_1280, i_8_1305, i_8_1306, i_8_1313, i_8_1323, i_8_1342, i_8_1343, i_8_1435, i_8_1436, i_8_1452, i_8_1504, i_8_1505, i_8_1542, i_8_1550, i_8_1562, i_8_1603, i_8_1613, i_8_1630, i_8_1676, i_8_1697, i_8_1711, i_8_1748, i_8_1749, i_8_1759, i_8_1802, i_8_1818, i_8_1856, i_8_1886, i_8_1892, i_8_1964, i_8_1973, i_8_1985, i_8_1994, i_8_2036, i_8_2075, i_8_2108, i_8_2134, i_8_2141, i_8_2143, i_8_2144, i_8_2145, i_8_2153, i_8_2171, i_8_2188, i_8_2246, i_8_2272, i_8_2288, o_8_348);
	kernel_8_349 k_8_349(i_8_6, i_8_24, i_8_25, i_8_78, i_8_115, i_8_177, i_8_249, i_8_250, i_8_265, i_8_349, i_8_355, i_8_357, i_8_373, i_8_384, i_8_385, i_8_395, i_8_445, i_8_465, i_8_475, i_8_481, i_8_493, i_8_501, i_8_520, i_8_522, i_8_556, i_8_580, i_8_673, i_8_710, i_8_762, i_8_770, i_8_771, i_8_807, i_8_842, i_8_850, i_8_856, i_8_861, i_8_889, i_8_944, i_8_967, i_8_968, i_8_1057, i_8_1059, i_8_1060, i_8_1087, i_8_1194, i_8_1227, i_8_1230, i_8_1239, i_8_1266, i_8_1272, i_8_1275, i_8_1276, i_8_1285, i_8_1299, i_8_1307, i_8_1317, i_8_1393, i_8_1399, i_8_1402, i_8_1404, i_8_1419, i_8_1432, i_8_1472, i_8_1473, i_8_1536, i_8_1538, i_8_1553, i_8_1632, i_8_1636, i_8_1654, i_8_1663, i_8_1699, i_8_1704, i_8_1716, i_8_1749, i_8_1808, i_8_1860, i_8_1862, i_8_1868, i_8_1879, i_8_1885, i_8_1888, i_8_1921, i_8_1929, i_8_1960, i_8_1969, i_8_1975, i_8_1995, i_8_2047, i_8_2058, i_8_2059, i_8_2068, i_8_2073, i_8_2076, i_8_2145, i_8_2158, i_8_2176, i_8_2219, i_8_2299, i_8_2302, o_8_349);
	kernel_8_350 k_8_350(i_8_10, i_8_13, i_8_38, i_8_40, i_8_41, i_8_47, i_8_50, i_8_73, i_8_91, i_8_136, i_8_143, i_8_182, i_8_193, i_8_239, i_8_254, i_8_334, i_8_344, i_8_362, i_8_364, i_8_397, i_8_398, i_8_423, i_8_425, i_8_427, i_8_428, i_8_451, i_8_452, i_8_490, i_8_491, i_8_532, i_8_533, i_8_578, i_8_595, i_8_608, i_8_612, i_8_613, i_8_640, i_8_641, i_8_675, i_8_676, i_8_677, i_8_694, i_8_695, i_8_699, i_8_700, i_8_748, i_8_775, i_8_782, i_8_796, i_8_839, i_8_844, i_8_856, i_8_857, i_8_858, i_8_878, i_8_973, i_8_1034, i_8_1036, i_8_1057, i_8_1154, i_8_1156, i_8_1226, i_8_1235, i_8_1236, i_8_1243, i_8_1292, i_8_1314, i_8_1315, i_8_1325, i_8_1411, i_8_1468, i_8_1489, i_8_1490, i_8_1564, i_8_1624, i_8_1632, i_8_1669, i_8_1694, i_8_1764, i_8_1765, i_8_1767, i_8_1783, i_8_1786, i_8_1818, i_8_1819, i_8_1830, i_8_1837, i_8_1885, i_8_1940, i_8_1969, i_8_2110, i_8_2111, i_8_2133, i_8_2147, i_8_2148, i_8_2152, i_8_2165, i_8_2225, i_8_2236, i_8_2263, o_8_350);
	kernel_8_351 k_8_351(i_8_22, i_8_29, i_8_34, i_8_56, i_8_57, i_8_73, i_8_95, i_8_136, i_8_184, i_8_231, i_8_253, i_8_254, i_8_259, i_8_305, i_8_365, i_8_378, i_8_398, i_8_424, i_8_454, i_8_469, i_8_505, i_8_506, i_8_554, i_8_581, i_8_586, i_8_609, i_8_622, i_8_637, i_8_639, i_8_678, i_8_680, i_8_704, i_8_706, i_8_709, i_8_710, i_8_730, i_8_751, i_8_778, i_8_785, i_8_839, i_8_856, i_8_866, i_8_875, i_8_965, i_8_1063, i_8_1064, i_8_1099, i_8_1102, i_8_1103, i_8_1130, i_8_1145, i_8_1265, i_8_1283, i_8_1297, i_8_1298, i_8_1299, i_8_1355, i_8_1360, i_8_1366, i_8_1385, i_8_1393, i_8_1397, i_8_1402, i_8_1431, i_8_1434, i_8_1462, i_8_1463, i_8_1471, i_8_1548, i_8_1559, i_8_1632, i_8_1633, i_8_1688, i_8_1705, i_8_1786, i_8_1789, i_8_1795, i_8_1812, i_8_1821, i_8_1886, i_8_1888, i_8_1889, i_8_1891, i_8_1940, i_8_1963, i_8_1989, i_8_2056, i_8_2101, i_8_2107, i_8_2131, i_8_2132, i_8_2153, i_8_2170, i_8_2225, i_8_2234, i_8_2244, i_8_2246, i_8_2261, i_8_2263, i_8_2264, o_8_351);
	kernel_8_352 k_8_352(i_8_18, i_8_21, i_8_33, i_8_34, i_8_52, i_8_105, i_8_114, i_8_173, i_8_203, i_8_223, i_8_300, i_8_307, i_8_319, i_8_356, i_8_372, i_8_374, i_8_381, i_8_391, i_8_392, i_8_497, i_8_518, i_8_594, i_8_597, i_8_600, i_8_604, i_8_608, i_8_610, i_8_640, i_8_657, i_8_661, i_8_668, i_8_675, i_8_678, i_8_681, i_8_748, i_8_776, i_8_850, i_8_860, i_8_867, i_8_870, i_8_871, i_8_878, i_8_896, i_8_974, i_8_986, i_8_1037, i_8_1085, i_8_1101, i_8_1102, i_8_1125, i_8_1126, i_8_1136, i_8_1140, i_8_1218, i_8_1228, i_8_1317, i_8_1362, i_8_1382, i_8_1443, i_8_1459, i_8_1462, i_8_1470, i_8_1499, i_8_1514, i_8_1517, i_8_1533, i_8_1557, i_8_1596, i_8_1605, i_8_1680, i_8_1688, i_8_1701, i_8_1702, i_8_1713, i_8_1733, i_8_1747, i_8_1748, i_8_1761, i_8_1762, i_8_1776, i_8_1782, i_8_1783, i_8_1810, i_8_1812, i_8_1817, i_8_1821, i_8_1890, i_8_1891, i_8_1903, i_8_1910, i_8_1947, i_8_1981, i_8_2056, i_8_2107, i_8_2129, i_8_2154, i_8_2201, i_8_2235, i_8_2241, i_8_2262, o_8_352);
	kernel_8_353 k_8_353(i_8_17, i_8_40, i_8_45, i_8_65, i_8_68, i_8_142, i_8_184, i_8_187, i_8_205, i_8_222, i_8_228, i_8_237, i_8_243, i_8_252, i_8_281, i_8_298, i_8_322, i_8_335, i_8_360, i_8_382, i_8_417, i_8_426, i_8_451, i_8_471, i_8_505, i_8_514, i_8_549, i_8_556, i_8_583, i_8_584, i_8_637, i_8_655, i_8_681, i_8_738, i_8_749, i_8_763, i_8_770, i_8_778, i_8_796, i_8_797, i_8_840, i_8_842, i_8_917, i_8_940, i_8_941, i_8_1053, i_8_1112, i_8_1137, i_8_1147, i_8_1155, i_8_1227, i_8_1234, i_8_1245, i_8_1246, i_8_1256, i_8_1280, i_8_1285, i_8_1286, i_8_1288, i_8_1296, i_8_1331, i_8_1332, i_8_1335, i_8_1336, i_8_1365, i_8_1367, i_8_1384, i_8_1400, i_8_1440, i_8_1464, i_8_1467, i_8_1528, i_8_1556, i_8_1606, i_8_1678, i_8_1689, i_8_1696, i_8_1702, i_8_1706, i_8_1714, i_8_1722, i_8_1745, i_8_1753, i_8_1754, i_8_1784, i_8_1787, i_8_1822, i_8_1883, i_8_1902, i_8_1963, i_8_1975, i_8_1996, i_8_2001, i_8_2073, i_8_2097, i_8_2106, i_8_2170, i_8_2224, i_8_2259, i_8_2280, o_8_353);
	kernel_8_354 k_8_354(i_8_16, i_8_34, i_8_185, i_8_257, i_8_281, i_8_283, i_8_338, i_8_383, i_8_391, i_8_392, i_8_400, i_8_418, i_8_450, i_8_451, i_8_509, i_8_554, i_8_557, i_8_563, i_8_569, i_8_583, i_8_633, i_8_644, i_8_652, i_8_653, i_8_663, i_8_700, i_8_703, i_8_704, i_8_751, i_8_769, i_8_782, i_8_785, i_8_823, i_8_827, i_8_842, i_8_866, i_8_874, i_8_895, i_8_958, i_8_969, i_8_1012, i_8_1013, i_8_1036, i_8_1109, i_8_1129, i_8_1132, i_8_1201, i_8_1285, i_8_1300, i_8_1303, i_8_1328, i_8_1357, i_8_1382, i_8_1411, i_8_1435, i_8_1436, i_8_1452, i_8_1468, i_8_1477, i_8_1478, i_8_1489, i_8_1511, i_8_1525, i_8_1526, i_8_1547, i_8_1553, i_8_1571, i_8_1603, i_8_1679, i_8_1696, i_8_1705, i_8_1706, i_8_1723, i_8_1750, i_8_1784, i_8_1794, i_8_1796, i_8_1807, i_8_1821, i_8_1822, i_8_1824, i_8_1840, i_8_1841, i_8_1868, i_8_1886, i_8_1894, i_8_1895, i_8_1912, i_8_1939, i_8_1976, i_8_1982, i_8_2074, i_8_2075, i_8_2154, i_8_2159, i_8_2182, i_8_2224, i_8_2227, i_8_2248, i_8_2276, o_8_354);
	kernel_8_355 k_8_355(i_8_50, i_8_59, i_8_76, i_8_85, i_8_104, i_8_107, i_8_118, i_8_218, i_8_304, i_8_322, i_8_362, i_8_367, i_8_368, i_8_374, i_8_385, i_8_414, i_8_453, i_8_488, i_8_524, i_8_530, i_8_547, i_8_556, i_8_557, i_8_608, i_8_611, i_8_616, i_8_633, i_8_634, i_8_652, i_8_655, i_8_656, i_8_657, i_8_661, i_8_662, i_8_665, i_8_697, i_8_700, i_8_707, i_8_760, i_8_769, i_8_772, i_8_827, i_8_844, i_8_869, i_8_877, i_8_886, i_8_943, i_8_956, i_8_958, i_8_959, i_8_965, i_8_970, i_8_977, i_8_991, i_8_1039, i_8_1115, i_8_1138, i_8_1256, i_8_1267, i_8_1268, i_8_1319, i_8_1348, i_8_1439, i_8_1453, i_8_1474, i_8_1489, i_8_1516, i_8_1525, i_8_1544, i_8_1546, i_8_1555, i_8_1562, i_8_1673, i_8_1732, i_8_1765, i_8_1787, i_8_1795, i_8_1813, i_8_1822, i_8_1859, i_8_1877, i_8_1887, i_8_1909, i_8_1915, i_8_1993, i_8_1996, i_8_2056, i_8_2090, i_8_2092, i_8_2093, i_8_2102, i_8_2125, i_8_2129, i_8_2135, i_8_2149, i_8_2156, i_8_2173, i_8_2227, i_8_2233, i_8_2245, o_8_355);
	kernel_8_356 k_8_356(i_8_39, i_8_88, i_8_136, i_8_159, i_8_183, i_8_187, i_8_265, i_8_285, i_8_295, i_8_300, i_8_322, i_8_331, i_8_363, i_8_364, i_8_368, i_8_393, i_8_399, i_8_420, i_8_426, i_8_459, i_8_510, i_8_565, i_8_591, i_8_592, i_8_594, i_8_598, i_8_608, i_8_612, i_8_660, i_8_673, i_8_681, i_8_683, i_8_703, i_8_707, i_8_736, i_8_750, i_8_809, i_8_826, i_8_832, i_8_835, i_8_838, i_8_841, i_8_843, i_8_850, i_8_927, i_8_1024, i_8_1050, i_8_1052, i_8_1055, i_8_1060, i_8_1132, i_8_1165, i_8_1200, i_8_1229, i_8_1231, i_8_1236, i_8_1240, i_8_1326, i_8_1375, i_8_1376, i_8_1381, i_8_1384, i_8_1402, i_8_1426, i_8_1456, i_8_1510, i_8_1524, i_8_1549, i_8_1552, i_8_1600, i_8_1635, i_8_1680, i_8_1686, i_8_1687, i_8_1704, i_8_1705, i_8_1796, i_8_1798, i_8_1819, i_8_1842, i_8_1884, i_8_1938, i_8_1939, i_8_1978, i_8_2048, i_8_2113, i_8_2121, i_8_2122, i_8_2131, i_8_2132, i_8_2140, i_8_2145, i_8_2147, i_8_2153, i_8_2172, i_8_2173, i_8_2224, i_8_2247, i_8_2256, i_8_2293, o_8_356);
	kernel_8_357 k_8_357(i_8_30, i_8_112, i_8_119, i_8_194, i_8_220, i_8_223, i_8_289, i_8_298, i_8_317, i_8_343, i_8_344, i_8_380, i_8_382, i_8_431, i_8_442, i_8_451, i_8_453, i_8_463, i_8_496, i_8_498, i_8_529, i_8_549, i_8_605, i_8_610, i_8_611, i_8_622, i_8_668, i_8_686, i_8_697, i_8_704, i_8_707, i_8_711, i_8_752, i_8_765, i_8_792, i_8_794, i_8_820, i_8_823, i_8_837, i_8_840, i_8_875, i_8_991, i_8_1004, i_8_1045, i_8_1046, i_8_1077, i_8_1103, i_8_1107, i_8_1111, i_8_1117, i_8_1139, i_8_1253, i_8_1271, i_8_1297, i_8_1324, i_8_1335, i_8_1355, i_8_1449, i_8_1451, i_8_1468, i_8_1478, i_8_1507, i_8_1536, i_8_1537, i_8_1541, i_8_1544, i_8_1549, i_8_1550, i_8_1594, i_8_1602, i_8_1620, i_8_1643, i_8_1649, i_8_1674, i_8_1749, i_8_1751, i_8_1801, i_8_1821, i_8_1856, i_8_1859, i_8_1863, i_8_1891, i_8_1901, i_8_1927, i_8_1962, i_8_2072, i_8_2089, i_8_2090, i_8_2107, i_8_2124, i_8_2125, i_8_2126, i_8_2132, i_8_2146, i_8_2242, i_8_2254, i_8_2268, i_8_2269, i_8_2270, i_8_2287, o_8_357);
	kernel_8_358 k_8_358(i_8_104, i_8_153, i_8_154, i_8_155, i_8_158, i_8_160, i_8_205, i_8_206, i_8_221, i_8_435, i_8_471, i_8_480, i_8_489, i_8_499, i_8_500, i_8_572, i_8_592, i_8_606, i_8_610, i_8_624, i_8_684, i_8_688, i_8_699, i_8_714, i_8_716, i_8_717, i_8_729, i_8_778, i_8_779, i_8_780, i_8_782, i_8_787, i_8_837, i_8_838, i_8_867, i_8_869, i_8_871, i_8_879, i_8_881, i_8_998, i_8_1008, i_8_1012, i_8_1026, i_8_1027, i_8_1031, i_8_1044, i_8_1112, i_8_1135, i_8_1154, i_8_1155, i_8_1229, i_8_1297, i_8_1300, i_8_1305, i_8_1306, i_8_1314, i_8_1341, i_8_1342, i_8_1343, i_8_1345, i_8_1346, i_8_1349, i_8_1355, i_8_1407, i_8_1434, i_8_1435, i_8_1436, i_8_1455, i_8_1542, i_8_1545, i_8_1548, i_8_1550, i_8_1551, i_8_1624, i_8_1647, i_8_1651, i_8_1652, i_8_1677, i_8_1682, i_8_1741, i_8_1748, i_8_1779, i_8_1803, i_8_1866, i_8_1884, i_8_1925, i_8_1945, i_8_1962, i_8_1983, i_8_1992, i_8_1994, i_8_1996, i_8_2049, i_8_2051, i_8_2147, i_8_2245, i_8_2271, i_8_2286, i_8_2290, i_8_2291, o_8_358);
	kernel_8_359 k_8_359(i_8_10, i_8_20, i_8_35, i_8_65, i_8_73, i_8_74, i_8_77, i_8_106, i_8_113, i_8_124, i_8_266, i_8_302, i_8_322, i_8_323, i_8_361, i_8_362, i_8_364, i_8_365, i_8_368, i_8_392, i_8_398, i_8_428, i_8_445, i_8_487, i_8_505, i_8_506, i_8_509, i_8_578, i_8_590, i_8_604, i_8_605, i_8_607, i_8_608, i_8_641, i_8_661, i_8_671, i_8_677, i_8_680, i_8_727, i_8_758, i_8_781, i_8_817, i_8_824, i_8_826, i_8_955, i_8_974, i_8_1037, i_8_1040, i_8_1109, i_8_1114, i_8_1127, i_8_1181, i_8_1183, i_8_1199, i_8_1225, i_8_1229, i_8_1244, i_8_1264, i_8_1265, i_8_1280, i_8_1295, i_8_1307, i_8_1315, i_8_1316, i_8_1325, i_8_1361, i_8_1397, i_8_1424, i_8_1436, i_8_1438, i_8_1460, i_8_1463, i_8_1465, i_8_1492, i_8_1510, i_8_1514, i_8_1522, i_8_1525, i_8_1549, i_8_1550, i_8_1553, i_8_1630, i_8_1631, i_8_1634, i_8_1679, i_8_1702, i_8_1747, i_8_1748, i_8_1792, i_8_1805, i_8_1819, i_8_1822, i_8_1838, i_8_1883, i_8_1976, i_8_1982, i_8_1993, i_8_2135, i_8_2245, i_8_2246, o_8_359);
	kernel_8_360 k_8_360(i_8_26, i_8_63, i_8_76, i_8_192, i_8_279, i_8_318, i_8_324, i_8_327, i_8_350, i_8_367, i_8_373, i_8_383, i_8_391, i_8_450, i_8_504, i_8_526, i_8_531, i_8_556, i_8_557, i_8_562, i_8_585, i_8_589, i_8_602, i_8_603, i_8_604, i_8_607, i_8_630, i_8_631, i_8_639, i_8_675, i_8_676, i_8_700, i_8_702, i_8_703, i_8_706, i_8_793, i_8_838, i_8_937, i_8_968, i_8_1008, i_8_1036, i_8_1047, i_8_1106, i_8_1179, i_8_1197, i_8_1200, i_8_1225, i_8_1246, i_8_1261, i_8_1264, i_8_1296, i_8_1298, i_8_1299, i_8_1315, i_8_1327, i_8_1341, i_8_1354, i_8_1359, i_8_1362, i_8_1422, i_8_1423, i_8_1433, i_8_1434, i_8_1440, i_8_1461, i_8_1476, i_8_1512, i_8_1513, i_8_1515, i_8_1522, i_8_1539, i_8_1543, i_8_1564, i_8_1632, i_8_1651, i_8_1682, i_8_1701, i_8_1747, i_8_1748, i_8_1773, i_8_1786, i_8_1791, i_8_1810, i_8_1829, i_8_1887, i_8_1953, i_8_1957, i_8_1989, i_8_2011, i_8_2072, i_8_2132, i_8_2140, i_8_2142, i_8_2144, i_8_2145, i_8_2146, i_8_2154, i_8_2223, i_8_2226, i_8_2227, o_8_360);
	kernel_8_361 k_8_361(i_8_0, i_8_63, i_8_84, i_8_139, i_8_283, i_8_381, i_8_383, i_8_423, i_8_482, i_8_499, i_8_516, i_8_520, i_8_525, i_8_526, i_8_527, i_8_528, i_8_549, i_8_579, i_8_609, i_8_700, i_8_704, i_8_705, i_8_751, i_8_777, i_8_778, i_8_850, i_8_937, i_8_968, i_8_970, i_8_1010, i_8_1047, i_8_1074, i_8_1117, i_8_1127, i_8_1128, i_8_1138, i_8_1180, i_8_1227, i_8_1263, i_8_1279, i_8_1283, i_8_1286, i_8_1294, i_8_1296, i_8_1297, i_8_1332, i_8_1359, i_8_1395, i_8_1434, i_8_1437, i_8_1438, i_8_1456, i_8_1457, i_8_1467, i_8_1469, i_8_1486, i_8_1489, i_8_1494, i_8_1531, i_8_1585, i_8_1600, i_8_1601, i_8_1602, i_8_1603, i_8_1620, i_8_1638, i_8_1664, i_8_1686, i_8_1728, i_8_1746, i_8_1748, i_8_1756, i_8_1758, i_8_1765, i_8_1768, i_8_1787, i_8_1789, i_8_1792, i_8_1804, i_8_1805, i_8_1807, i_8_1808, i_8_1873, i_8_1881, i_8_1948, i_8_1951, i_8_1963, i_8_1965, i_8_1966, i_8_1970, i_8_2047, i_8_2068, i_8_2101, i_8_2133, i_8_2136, i_8_2140, i_8_2149, i_8_2226, i_8_2273, i_8_2295, o_8_361);
	kernel_8_362 k_8_362(i_8_25, i_8_33, i_8_62, i_8_98, i_8_140, i_8_160, i_8_192, i_8_197, i_8_224, i_8_250, i_8_268, i_8_291, i_8_338, i_8_357, i_8_359, i_8_384, i_8_420, i_8_458, i_8_464, i_8_480, i_8_485, i_8_503, i_8_522, i_8_528, i_8_570, i_8_629, i_8_709, i_8_715, i_8_726, i_8_764, i_8_787, i_8_817, i_8_907, i_8_922, i_8_924, i_8_952, i_8_985, i_8_987, i_8_1075, i_8_1113, i_8_1124, i_8_1128, i_8_1132, i_8_1137, i_8_1138, i_8_1140, i_8_1194, i_8_1419, i_8_1420, i_8_1421, i_8_1429, i_8_1437, i_8_1455, i_8_1483, i_8_1527, i_8_1543, i_8_1545, i_8_1554, i_8_1601, i_8_1609, i_8_1617, i_8_1618, i_8_1635, i_8_1663, i_8_1671, i_8_1672, i_8_1717, i_8_1732, i_8_1733, i_8_1743, i_8_1744, i_8_1750, i_8_1762, i_8_1797, i_8_1808, i_8_1821, i_8_1839, i_8_1872, i_8_1875, i_8_1877, i_8_1880, i_8_1906, i_8_1921, i_8_1922, i_8_1929, i_8_1966, i_8_1967, i_8_1984, i_8_2031, i_8_2049, i_8_2055, i_8_2059, i_8_2096, i_8_2112, i_8_2120, i_8_2154, i_8_2218, i_8_2219, i_8_2229, i_8_2274, o_8_362);
	kernel_8_363 k_8_363(i_8_31, i_8_38, i_8_83, i_8_139, i_8_217, i_8_229, i_8_281, i_8_304, i_8_379, i_8_388, i_8_416, i_8_425, i_8_439, i_8_442, i_8_443, i_8_453, i_8_473, i_8_550, i_8_571, i_8_585, i_8_586, i_8_587, i_8_604, i_8_605, i_8_608, i_8_611, i_8_622, i_8_631, i_8_638, i_8_667, i_8_669, i_8_677, i_8_685, i_8_704, i_8_736, i_8_749, i_8_821, i_8_830, i_8_839, i_8_864, i_8_967, i_8_968, i_8_1009, i_8_1031, i_8_1100, i_8_1118, i_8_1130, i_8_1154, i_8_1180, i_8_1181, i_8_1225, i_8_1226, i_8_1234, i_8_1235, i_8_1270, i_8_1280, i_8_1316, i_8_1327, i_8_1334, i_8_1406, i_8_1439, i_8_1460, i_8_1534, i_8_1536, i_8_1549, i_8_1555, i_8_1595, i_8_1658, i_8_1670, i_8_1681, i_8_1709, i_8_1745, i_8_1757, i_8_1758, i_8_1759, i_8_1774, i_8_1837, i_8_1838, i_8_1841, i_8_1891, i_8_1892, i_8_1895, i_8_1936, i_8_1963, i_8_1964, i_8_2008, i_8_2026, i_8_2037, i_8_2072, i_8_2108, i_8_2110, i_8_2140, i_8_2142, i_8_2143, i_8_2145, i_8_2152, i_8_2171, i_8_2188, i_8_2189, i_8_2191, o_8_363);
	kernel_8_364 k_8_364(i_8_12, i_8_44, i_8_66, i_8_106, i_8_115, i_8_133, i_8_139, i_8_172, i_8_256, i_8_273, i_8_283, i_8_309, i_8_321, i_8_381, i_8_399, i_8_400, i_8_471, i_8_498, i_8_524, i_8_549, i_8_555, i_8_571, i_8_577, i_8_591, i_8_608, i_8_630, i_8_635, i_8_642, i_8_666, i_8_672, i_8_681, i_8_707, i_8_750, i_8_780, i_8_825, i_8_841, i_8_845, i_8_966, i_8_967, i_8_1035, i_8_1038, i_8_1039, i_8_1042, i_8_1072, i_8_1074, i_8_1225, i_8_1227, i_8_1236, i_8_1237, i_8_1246, i_8_1263, i_8_1270, i_8_1300, i_8_1314, i_8_1317, i_8_1318, i_8_1327, i_8_1330, i_8_1338, i_8_1362, i_8_1372, i_8_1390, i_8_1422, i_8_1437, i_8_1442, i_8_1464, i_8_1465, i_8_1506, i_8_1525, i_8_1527, i_8_1545, i_8_1564, i_8_1573, i_8_1623, i_8_1636, i_8_1641, i_8_1651, i_8_1678, i_8_1681, i_8_1698, i_8_1782, i_8_1787, i_8_1824, i_8_1893, i_8_1912, i_8_1938, i_8_1960, i_8_1969, i_8_1975, i_8_1977, i_8_1984, i_8_2071, i_8_2179, i_8_2208, i_8_2226, i_8_2231, i_8_2246, i_8_2247, i_8_2271, i_8_2298, o_8_364);
	kernel_8_365 k_8_365(i_8_18, i_8_19, i_8_47, i_8_51, i_8_54, i_8_55, i_8_58, i_8_138, i_8_216, i_8_228, i_8_229, i_8_252, i_8_272, i_8_292, i_8_350, i_8_363, i_8_399, i_8_427, i_8_433, i_8_436, i_8_457, i_8_552, i_8_597, i_8_615, i_8_621, i_8_631, i_8_657, i_8_664, i_8_665, i_8_689, i_8_697, i_8_699, i_8_709, i_8_716, i_8_729, i_8_730, i_8_759, i_8_783, i_8_792, i_8_847, i_8_880, i_8_990, i_8_998, i_8_1027, i_8_1045, i_8_1047, i_8_1077, i_8_1090, i_8_1109, i_8_1117, i_8_1129, i_8_1188, i_8_1233, i_8_1266, i_8_1270, i_8_1317, i_8_1369, i_8_1436, i_8_1441, i_8_1449, i_8_1452, i_8_1467, i_8_1468, i_8_1505, i_8_1534, i_8_1539, i_8_1546, i_8_1562, i_8_1591, i_8_1603, i_8_1611, i_8_1620, i_8_1629, i_8_1658, i_8_1666, i_8_1676, i_8_1678, i_8_1679, i_8_1681, i_8_1682, i_8_1740, i_8_1802, i_8_1855, i_8_1856, i_8_1873, i_8_1989, i_8_1991, i_8_2029, i_8_2035, i_8_2046, i_8_2053, i_8_2093, i_8_2125, i_8_2138, i_8_2139, i_8_2156, i_8_2232, i_8_2259, i_8_2261, i_8_2286, o_8_365);
	kernel_8_366 k_8_366(i_8_30, i_8_33, i_8_53, i_8_79, i_8_84, i_8_118, i_8_138, i_8_165, i_8_184, i_8_187, i_8_192, i_8_210, i_8_240, i_8_241, i_8_301, i_8_336, i_8_369, i_8_381, i_8_382, i_8_439, i_8_472, i_8_522, i_8_543, i_8_573, i_8_608, i_8_638, i_8_760, i_8_771, i_8_774, i_8_810, i_8_811, i_8_858, i_8_861, i_8_878, i_8_879, i_8_939, i_8_940, i_8_968, i_8_984, i_8_1059, i_8_1060, i_8_1133, i_8_1138, i_8_1182, i_8_1188, i_8_1191, i_8_1264, i_8_1266, i_8_1269, i_8_1282, i_8_1287, i_8_1288, i_8_1291, i_8_1293, i_8_1305, i_8_1326, i_8_1333, i_8_1386, i_8_1387, i_8_1403, i_8_1407, i_8_1411, i_8_1489, i_8_1531, i_8_1545, i_8_1553, i_8_1600, i_8_1614, i_8_1633, i_8_1678, i_8_1681, i_8_1713, i_8_1719, i_8_1720, i_8_1731, i_8_1734, i_8_1747, i_8_1758, i_8_1759, i_8_1771, i_8_1783, i_8_1790, i_8_1796, i_8_1804, i_8_1822, i_8_1839, i_8_1857, i_8_1885, i_8_1918, i_8_1981, i_8_1998, i_8_2022, i_8_2047, i_8_2056, i_8_2124, i_8_2149, i_8_2169, i_8_2223, i_8_2235, i_8_2298, o_8_366);
	kernel_8_367 k_8_367(i_8_51, i_8_97, i_8_120, i_8_138, i_8_163, i_8_193, i_8_202, i_8_233, i_8_246, i_8_252, i_8_256, i_8_264, i_8_282, i_8_291, i_8_292, i_8_293, i_8_321, i_8_328, i_8_330, i_8_345, i_8_346, i_8_364, i_8_394, i_8_437, i_8_439, i_8_450, i_8_455, i_8_456, i_8_480, i_8_598, i_8_601, i_8_612, i_8_616, i_8_672, i_8_701, i_8_702, i_8_706, i_8_709, i_8_715, i_8_723, i_8_786, i_8_797, i_8_822, i_8_826, i_8_874, i_8_966, i_8_969, i_8_972, i_8_995, i_8_1050, i_8_1061, i_8_1074, i_8_1080, i_8_1081, i_8_1119, i_8_1182, i_8_1234, i_8_1237, i_8_1273, i_8_1347, i_8_1354, i_8_1389, i_8_1390, i_8_1408, i_8_1411, i_8_1437, i_8_1439, i_8_1452, i_8_1464, i_8_1527, i_8_1545, i_8_1546, i_8_1570, i_8_1573, i_8_1632, i_8_1681, i_8_1719, i_8_1746, i_8_1758, i_8_1759, i_8_1867, i_8_1884, i_8_1885, i_8_1887, i_8_1902, i_8_1948, i_8_1992, i_8_1995, i_8_2028, i_8_2031, i_8_2056, i_8_2058, i_8_2077, i_8_2128, i_8_2140, i_8_2156, i_8_2190, i_8_2215, i_8_2216, i_8_2270, o_8_367);
	kernel_8_368 k_8_368(i_8_13, i_8_50, i_8_139, i_8_170, i_8_188, i_8_192, i_8_226, i_8_229, i_8_257, i_8_263, i_8_277, i_8_278, i_8_283, i_8_365, i_8_383, i_8_385, i_8_425, i_8_449, i_8_454, i_8_457, i_8_490, i_8_493, i_8_526, i_8_528, i_8_530, i_8_544, i_8_606, i_8_613, i_8_617, i_8_631, i_8_632, i_8_655, i_8_656, i_8_661, i_8_703, i_8_709, i_8_710, i_8_785, i_8_798, i_8_854, i_8_866, i_8_892, i_8_935, i_8_977, i_8_1019, i_8_1023, i_8_1060, i_8_1075, i_8_1103, i_8_1163, i_8_1174, i_8_1228, i_8_1280, i_8_1282, i_8_1307, i_8_1334, i_8_1379, i_8_1414, i_8_1424, i_8_1471, i_8_1538, i_8_1558, i_8_1610, i_8_1642, i_8_1655, i_8_1685, i_8_1705, i_8_1750, i_8_1811, i_8_1849, i_8_1910, i_8_1913, i_8_1946, i_8_1952, i_8_1964, i_8_1973, i_8_1978, i_8_1982, i_8_1997, i_8_2006, i_8_2009, i_8_2038, i_8_2039, i_8_2091, i_8_2095, i_8_2126, i_8_2144, i_8_2146, i_8_2164, i_8_2168, i_8_2171, i_8_2173, i_8_2183, i_8_2186, i_8_2228, i_8_2239, i_8_2249, i_8_2259, i_8_2268, i_8_2293, o_8_368);
	kernel_8_369 k_8_369(i_8_37, i_8_52, i_8_80, i_8_89, i_8_130, i_8_139, i_8_166, i_8_192, i_8_304, i_8_325, i_8_356, i_8_367, i_8_368, i_8_464, i_8_483, i_8_486, i_8_487, i_8_489, i_8_517, i_8_518, i_8_526, i_8_527, i_8_595, i_8_608, i_8_613, i_8_621, i_8_696, i_8_699, i_8_705, i_8_748, i_8_750, i_8_757, i_8_760, i_8_761, i_8_829, i_8_840, i_8_841, i_8_869, i_8_967, i_8_981, i_8_982, i_8_990, i_8_1074, i_8_1075, i_8_1076, i_8_1084, i_8_1128, i_8_1224, i_8_1234, i_8_1264, i_8_1265, i_8_1268, i_8_1273, i_8_1282, i_8_1305, i_8_1327, i_8_1331, i_8_1358, i_8_1408, i_8_1476, i_8_1481, i_8_1498, i_8_1499, i_8_1548, i_8_1557, i_8_1579, i_8_1613, i_8_1642, i_8_1648, i_8_1670, i_8_1710, i_8_1729, i_8_1746, i_8_1748, i_8_1753, i_8_1754, i_8_1779, i_8_1783, i_8_1787, i_8_1795, i_8_1800, i_8_1821, i_8_1858, i_8_1867, i_8_1877, i_8_1900, i_8_1999, i_8_2003, i_8_2008, i_8_2026, i_8_2047, i_8_2080, i_8_2154, i_8_2170, i_8_2174, i_8_2215, i_8_2216, i_8_2246, i_8_2253, i_8_2260, o_8_369);
	kernel_8_370 k_8_370(i_8_4, i_8_18, i_8_20, i_8_35, i_8_40, i_8_41, i_8_88, i_8_114, i_8_115, i_8_166, i_8_184, i_8_275, i_8_307, i_8_319, i_8_320, i_8_335, i_8_343, i_8_364, i_8_418, i_8_419, i_8_427, i_8_453, i_8_454, i_8_508, i_8_526, i_8_554, i_8_572, i_8_590, i_8_599, i_8_613, i_8_614, i_8_635, i_8_638, i_8_640, i_8_671, i_8_695, i_8_769, i_8_882, i_8_893, i_8_991, i_8_1033, i_8_1040, i_8_1061, i_8_1084, i_8_1112, i_8_1115, i_8_1129, i_8_1130, i_8_1174, i_8_1226, i_8_1229, i_8_1240, i_8_1270, i_8_1298, i_8_1300, i_8_1396, i_8_1397, i_8_1408, i_8_1481, i_8_1498, i_8_1526, i_8_1532, i_8_1544, i_8_1546, i_8_1552, i_8_1630, i_8_1640, i_8_1642, i_8_1648, i_8_1651, i_8_1661, i_8_1663, i_8_1693, i_8_1694, i_8_1705, i_8_1707, i_8_1750, i_8_1754, i_8_1779, i_8_1807, i_8_1858, i_8_1883, i_8_1885, i_8_1886, i_8_1949, i_8_1966, i_8_1968, i_8_2000, i_8_2054, i_8_2093, i_8_2094, i_8_2135, i_8_2139, i_8_2140, i_8_2170, i_8_2171, i_8_2192, i_8_2233, i_8_2257, i_8_2258, o_8_370);
	kernel_8_371 k_8_371(i_8_14, i_8_60, i_8_61, i_8_76, i_8_140, i_8_188, i_8_263, i_8_341, i_8_362, i_8_422, i_8_457, i_8_491, i_8_494, i_8_512, i_8_523, i_8_575, i_8_607, i_8_610, i_8_633, i_8_652, i_8_700, i_8_709, i_8_719, i_8_736, i_8_773, i_8_781, i_8_787, i_8_788, i_8_863, i_8_871, i_8_912, i_8_998, i_8_1075, i_8_1106, i_8_1111, i_8_1112, i_8_1114, i_8_1115, i_8_1157, i_8_1202, i_8_1204, i_8_1229, i_8_1231, i_8_1240, i_8_1247, i_8_1263, i_8_1300, i_8_1319, i_8_1322, i_8_1329, i_8_1331, i_8_1334, i_8_1397, i_8_1401, i_8_1402, i_8_1403, i_8_1435, i_8_1439, i_8_1445, i_8_1466, i_8_1490, i_8_1528, i_8_1552, i_8_1555, i_8_1597, i_8_1640, i_8_1645, i_8_1667, i_8_1679, i_8_1703, i_8_1717, i_8_1724, i_8_1748, i_8_1751, i_8_1762, i_8_1771, i_8_1778, i_8_1787, i_8_1808, i_8_1825, i_8_1835, i_8_1841, i_8_1848, i_8_1884, i_8_1888, i_8_1895, i_8_1948, i_8_1952, i_8_1966, i_8_1992, i_8_2012, i_8_2138, i_8_2140, i_8_2144, i_8_2147, i_8_2236, i_8_2237, i_8_2249, i_8_2264, i_8_2290, o_8_371);
	kernel_8_372 k_8_372(i_8_34, i_8_88, i_8_96, i_8_143, i_8_258, i_8_330, i_8_331, i_8_332, i_8_349, i_8_363, i_8_366, i_8_385, i_8_448, i_8_449, i_8_466, i_8_485, i_8_502, i_8_522, i_8_523, i_8_524, i_8_527, i_8_553, i_8_556, i_8_557, i_8_599, i_8_601, i_8_663, i_8_871, i_8_898, i_8_926, i_8_988, i_8_989, i_8_993, i_8_994, i_8_996, i_8_1015, i_8_1016, i_8_1032, i_8_1069, i_8_1074, i_8_1087, i_8_1088, i_8_1112, i_8_1120, i_8_1138, i_8_1140, i_8_1195, i_8_1258, i_8_1264, i_8_1265, i_8_1282, i_8_1286, i_8_1307, i_8_1309, i_8_1456, i_8_1528, i_8_1536, i_8_1543, i_8_1552, i_8_1555, i_8_1556, i_8_1574, i_8_1610, i_8_1617, i_8_1628, i_8_1635, i_8_1636, i_8_1637, i_8_1651, i_8_1652, i_8_1671, i_8_1672, i_8_1673, i_8_1679, i_8_1699, i_8_1700, i_8_1704, i_8_1717, i_8_1735, i_8_1736, i_8_1750, i_8_1809, i_8_1810, i_8_1858, i_8_1861, i_8_1905, i_8_1906, i_8_1933, i_8_1934, i_8_1992, i_8_1994, i_8_1995, i_8_2005, i_8_2006, i_8_2015, i_8_2114, i_8_2146, i_8_2215, i_8_2266, i_8_2267, o_8_372);
	kernel_8_373 k_8_373(i_8_0, i_8_1, i_8_31, i_8_81, i_8_82, i_8_83, i_8_84, i_8_102, i_8_111, i_8_184, i_8_203, i_8_244, i_8_259, i_8_280, i_8_306, i_8_307, i_8_342, i_8_343, i_8_346, i_8_349, i_8_350, i_8_360, i_8_388, i_8_423, i_8_424, i_8_450, i_8_460, i_8_599, i_8_603, i_8_630, i_8_632, i_8_634, i_8_661, i_8_702, i_8_706, i_8_710, i_8_711, i_8_712, i_8_756, i_8_757, i_8_758, i_8_779, i_8_780, i_8_811, i_8_838, i_8_858, i_8_993, i_8_996, i_8_1035, i_8_1078, i_8_1093, i_8_1098, i_8_1099, i_8_1100, i_8_1101, i_8_1103, i_8_1110, i_8_1115, i_8_1260, i_8_1266, i_8_1314, i_8_1328, i_8_1331, i_8_1388, i_8_1438, i_8_1507, i_8_1516, i_8_1532, i_8_1533, i_8_1642, i_8_1678, i_8_1679, i_8_1683, i_8_1684, i_8_1685, i_8_1759, i_8_1763, i_8_1779, i_8_1804, i_8_1805, i_8_1826, i_8_1935, i_8_1936, i_8_1937, i_8_1938, i_8_1939, i_8_1964, i_8_1969, i_8_2026, i_8_2115, i_8_2116, i_8_2117, i_8_2136, i_8_2137, i_8_2138, i_8_2229, i_8_2245, i_8_2248, i_8_2260, i_8_2270, o_8_373);
	kernel_8_374 k_8_374(i_8_6, i_8_7, i_8_37, i_8_41, i_8_64, i_8_111, i_8_130, i_8_172, i_8_178, i_8_263, i_8_297, i_8_301, i_8_307, i_8_316, i_8_319, i_8_355, i_8_356, i_8_361, i_8_363, i_8_414, i_8_424, i_8_447, i_8_527, i_8_532, i_8_568, i_8_612, i_8_624, i_8_639, i_8_661, i_8_664, i_8_667, i_8_675, i_8_682, i_8_684, i_8_704, i_8_796, i_8_837, i_8_838, i_8_853, i_8_870, i_8_874, i_8_975, i_8_1008, i_8_1053, i_8_1099, i_8_1126, i_8_1145, i_8_1174, i_8_1225, i_8_1233, i_8_1241, i_8_1285, i_8_1296, i_8_1297, i_8_1331, i_8_1337, i_8_1350, i_8_1380, i_8_1383, i_8_1446, i_8_1467, i_8_1488, i_8_1510, i_8_1522, i_8_1614, i_8_1631, i_8_1638, i_8_1645, i_8_1705, i_8_1707, i_8_1750, i_8_1764, i_8_1768, i_8_1773, i_8_1781, i_8_1809, i_8_1819, i_8_1855, i_8_1887, i_8_1891, i_8_1929, i_8_1935, i_8_1948, i_8_1953, i_8_2012, i_8_2016, i_8_2044, i_8_2053, i_8_2061, i_8_2071, i_8_2079, i_8_2080, i_8_2134, i_8_2140, i_8_2167, i_8_2185, i_8_2216, i_8_2230, i_8_2236, i_8_2284, o_8_374);
	kernel_8_375 k_8_375(i_8_21, i_8_45, i_8_73, i_8_129, i_8_130, i_8_147, i_8_150, i_8_192, i_8_193, i_8_222, i_8_329, i_8_355, i_8_378, i_8_385, i_8_462, i_8_472, i_8_493, i_8_516, i_8_517, i_8_519, i_8_525, i_8_549, i_8_606, i_8_613, i_8_624, i_8_631, i_8_652, i_8_658, i_8_659, i_8_661, i_8_694, i_8_703, i_8_705, i_8_715, i_8_733, i_8_831, i_8_832, i_8_876, i_8_879, i_8_925, i_8_963, i_8_1000, i_8_1003, i_8_1059, i_8_1086, i_8_1158, i_8_1164, i_8_1192, i_8_1224, i_8_1266, i_8_1281, i_8_1284, i_8_1302, i_8_1335, i_8_1336, i_8_1348, i_8_1354, i_8_1390, i_8_1435, i_8_1438, i_8_1455, i_8_1464, i_8_1489, i_8_1498, i_8_1539, i_8_1593, i_8_1596, i_8_1621, i_8_1641, i_8_1650, i_8_1659, i_8_1660, i_8_1662, i_8_1696, i_8_1704, i_8_1740, i_8_1743, i_8_1750, i_8_1875, i_8_1876, i_8_1881, i_8_1974, i_8_2010, i_8_2011, i_8_2046, i_8_2047, i_8_2057, i_8_2064, i_8_2092, i_8_2118, i_8_2146, i_8_2169, i_8_2172, i_8_2173, i_8_2185, i_8_2209, i_8_2253, i_8_2254, i_8_2256, i_8_2257, o_8_375);
	kernel_8_376 k_8_376(i_8_11, i_8_27, i_8_32, i_8_51, i_8_97, i_8_141, i_8_142, i_8_169, i_8_223, i_8_224, i_8_230, i_8_259, i_8_260, i_8_346, i_8_372, i_8_418, i_8_440, i_8_480, i_8_501, i_8_505, i_8_507, i_8_523, i_8_524, i_8_555, i_8_556, i_8_591, i_8_598, i_8_602, i_8_617, i_8_649, i_8_687, i_8_692, i_8_702, i_8_705, i_8_750, i_8_760, i_8_762, i_8_763, i_8_838, i_8_843, i_8_844, i_8_850, i_8_886, i_8_958, i_8_969, i_8_994, i_8_1032, i_8_1051, i_8_1074, i_8_1075, i_8_1077, i_8_1094, i_8_1096, i_8_1123, i_8_1124, i_8_1191, i_8_1222, i_8_1282, i_8_1285, i_8_1305, i_8_1306, i_8_1316, i_8_1318, i_8_1330, i_8_1331, i_8_1386, i_8_1387, i_8_1390, i_8_1410, i_8_1411, i_8_1470, i_8_1471, i_8_1507, i_8_1509, i_8_1533, i_8_1548, i_8_1560, i_8_1564, i_8_1573, i_8_1574, i_8_1635, i_8_1655, i_8_1680, i_8_1681, i_8_1682, i_8_1704, i_8_1722, i_8_1723, i_8_1821, i_8_1834, i_8_1858, i_8_1906, i_8_2032, i_8_2119, i_8_2122, i_8_2145, i_8_2211, i_8_2214, i_8_2215, i_8_2216, o_8_376);
	kernel_8_377 k_8_377(i_8_3, i_8_6, i_8_7, i_8_19, i_8_36, i_8_84, i_8_87, i_8_184, i_8_193, i_8_230, i_8_246, i_8_247, i_8_249, i_8_250, i_8_347, i_8_350, i_8_360, i_8_361, i_8_427, i_8_430, i_8_439, i_8_499, i_8_518, i_8_525, i_8_528, i_8_571, i_8_573, i_8_597, i_8_601, i_8_606, i_8_607, i_8_608, i_8_654, i_8_661, i_8_669, i_8_672, i_8_685, i_8_703, i_8_706, i_8_717, i_8_718, i_8_726, i_8_762, i_8_777, i_8_813, i_8_814, i_8_816, i_8_817, i_8_831, i_8_832, i_8_838, i_8_1071, i_8_1074, i_8_1084, i_8_1155, i_8_1159, i_8_1192, i_8_1285, i_8_1291, i_8_1295, i_8_1389, i_8_1392, i_8_1434, i_8_1497, i_8_1498, i_8_1542, i_8_1573, i_8_1658, i_8_1696, i_8_1749, i_8_1763, i_8_1819, i_8_1830, i_8_1833, i_8_1848, i_8_1851, i_8_1852, i_8_1866, i_8_1915, i_8_1938, i_8_1946, i_8_1947, i_8_1963, i_8_1974, i_8_1984, i_8_1985, i_8_2028, i_8_2031, i_8_2037, i_8_2047, i_8_2056, i_8_2064, i_8_2073, i_8_2076, i_8_2091, i_8_2095, i_8_2113, i_8_2118, i_8_2246, i_8_2281, o_8_377);
	kernel_8_378 k_8_378(i_8_33, i_8_96, i_8_97, i_8_114, i_8_211, i_8_258, i_8_259, i_8_294, i_8_297, i_8_298, i_8_330, i_8_367, i_8_421, i_8_442, i_8_444, i_8_445, i_8_457, i_8_476, i_8_483, i_8_484, i_8_525, i_8_555, i_8_568, i_8_602, i_8_607, i_8_609, i_8_660, i_8_661, i_8_662, i_8_705, i_8_706, i_8_780, i_8_781, i_8_834, i_8_840, i_8_867, i_8_877, i_8_886, i_8_990, i_8_993, i_8_1026, i_8_1060, i_8_1071, i_8_1072, i_8_1074, i_8_1084, i_8_1111, i_8_1113, i_8_1141, i_8_1239, i_8_1261, i_8_1274, i_8_1283, i_8_1284, i_8_1285, i_8_1327, i_8_1392, i_8_1393, i_8_1408, i_8_1435, i_8_1437, i_8_1438, i_8_1507, i_8_1538, i_8_1584, i_8_1587, i_8_1590, i_8_1591, i_8_1598, i_8_1632, i_8_1633, i_8_1679, i_8_1699, i_8_1741, i_8_1744, i_8_1759, i_8_1761, i_8_1762, i_8_1821, i_8_1824, i_8_1825, i_8_1862, i_8_1902, i_8_1918, i_8_1989, i_8_1996, i_8_2058, i_8_2076, i_8_2089, i_8_2111, i_8_2114, i_8_2125, i_8_2187, i_8_2214, i_8_2215, i_8_2248, i_8_2249, i_8_2262, i_8_2295, i_8_2303, o_8_378);
	kernel_8_379 k_8_379(i_8_3, i_8_4, i_8_39, i_8_67, i_8_147, i_8_192, i_8_201, i_8_228, i_8_244, i_8_246, i_8_247, i_8_307, i_8_378, i_8_379, i_8_390, i_8_418, i_8_427, i_8_469, i_8_472, i_8_481, i_8_495, i_8_507, i_8_516, i_8_555, i_8_571, i_8_594, i_8_598, i_8_634, i_8_659, i_8_707, i_8_748, i_8_753, i_8_759, i_8_762, i_8_813, i_8_840, i_8_858, i_8_867, i_8_913, i_8_954, i_8_955, i_8_963, i_8_967, i_8_1030, i_8_1036, i_8_1071, i_8_1173, i_8_1191, i_8_1200, i_8_1203, i_8_1236, i_8_1269, i_8_1270, i_8_1296, i_8_1336, i_8_1353, i_8_1354, i_8_1389, i_8_1390, i_8_1401, i_8_1407, i_8_1485, i_8_1489, i_8_1494, i_8_1495, i_8_1497, i_8_1534, i_8_1597, i_8_1641, i_8_1651, i_8_1659, i_8_1696, i_8_1748, i_8_1750, i_8_1777, i_8_1794, i_8_1836, i_8_1848, i_8_1849, i_8_1855, i_8_1863, i_8_1872, i_8_1873, i_8_1882, i_8_1888, i_8_1911, i_8_1948, i_8_1950, i_8_1965, i_8_1971, i_8_2010, i_8_2047, i_8_2065, i_8_2091, i_8_2119, i_8_2146, i_8_2149, i_8_2229, i_8_2233, i_8_2256, o_8_379);
	kernel_8_380 k_8_380(i_8_28, i_8_31, i_8_54, i_8_56, i_8_118, i_8_218, i_8_221, i_8_227, i_8_253, i_8_365, i_8_417, i_8_451, i_8_478, i_8_480, i_8_481, i_8_500, i_8_507, i_8_545, i_8_552, i_8_553, i_8_582, i_8_594, i_8_599, i_8_604, i_8_606, i_8_607, i_8_608, i_8_612, i_8_649, i_8_655, i_8_660, i_8_715, i_8_756, i_8_768, i_8_781, i_8_789, i_8_795, i_8_847, i_8_903, i_8_981, i_8_1008, i_8_1059, i_8_1060, i_8_1110, i_8_1111, i_8_1127, i_8_1130, i_8_1234, i_8_1260, i_8_1261, i_8_1292, i_8_1297, i_8_1307, i_8_1344, i_8_1345, i_8_1350, i_8_1379, i_8_1401, i_8_1416, i_8_1431, i_8_1443, i_8_1468, i_8_1541, i_8_1552, i_8_1555, i_8_1578, i_8_1588, i_8_1603, i_8_1680, i_8_1752, i_8_1753, i_8_1755, i_8_1756, i_8_1775, i_8_1783, i_8_1784, i_8_1788, i_8_1789, i_8_1801, i_8_1810, i_8_1822, i_8_1825, i_8_1837, i_8_1945, i_8_1946, i_8_1949, i_8_1973, i_8_1998, i_8_2050, i_8_2133, i_8_2142, i_8_2152, i_8_2153, i_8_2170, i_8_2214, i_8_2224, i_8_2227, i_8_2232, i_8_2287, i_8_2292, o_8_380);
	kernel_8_381 k_8_381(i_8_32, i_8_51, i_8_95, i_8_97, i_8_114, i_8_115, i_8_141, i_8_258, i_8_331, i_8_332, i_8_377, i_8_383, i_8_421, i_8_457, i_8_462, i_8_463, i_8_476, i_8_479, i_8_482, i_8_527, i_8_553, i_8_556, i_8_606, i_8_608, i_8_661, i_8_662, i_8_663, i_8_682, i_8_782, i_8_817, i_8_818, i_8_840, i_8_841, i_8_847, i_8_851, i_8_1074, i_8_1077, i_8_1239, i_8_1240, i_8_1259, i_8_1283, i_8_1292, i_8_1307, i_8_1437, i_8_1438, i_8_1439, i_8_1534, i_8_1535, i_8_1540, i_8_1551, i_8_1588, i_8_1589, i_8_1590, i_8_1591, i_8_1592, i_8_1600, i_8_1615, i_8_1616, i_8_1633, i_8_1634, i_8_1636, i_8_1637, i_8_1671, i_8_1679, i_8_1680, i_8_1742, i_8_1744, i_8_1751, i_8_1760, i_8_1761, i_8_1762, i_8_1763, i_8_1825, i_8_1826, i_8_1834, i_8_1839, i_8_1843, i_8_1879, i_8_1904, i_8_1922, i_8_1967, i_8_1985, i_8_1993, i_8_1994, i_8_1997, i_8_2056, i_8_2059, i_8_2090, i_8_2107, i_8_2130, i_8_2149, i_8_2172, i_8_2190, i_8_2214, i_8_2215, i_8_2216, i_8_2219, i_8_2264, i_8_2296, i_8_2303, o_8_381);
	kernel_8_382 k_8_382(i_8_28, i_8_57, i_8_87, i_8_143, i_8_214, i_8_264, i_8_268, i_8_269, i_8_328, i_8_349, i_8_360, i_8_376, i_8_378, i_8_379, i_8_381, i_8_384, i_8_417, i_8_463, i_8_481, i_8_490, i_8_500, i_8_529, i_8_589, i_8_590, i_8_592, i_8_599, i_8_608, i_8_611, i_8_615, i_8_616, i_8_628, i_8_633, i_8_637, i_8_638, i_8_661, i_8_664, i_8_670, i_8_682, i_8_715, i_8_716, i_8_760, i_8_769, i_8_778, i_8_823, i_8_843, i_8_870, i_8_871, i_8_898, i_8_899, i_8_984, i_8_985, i_8_1016, i_8_1079, i_8_1086, i_8_1110, i_8_1111, i_8_1114, i_8_1189, i_8_1236, i_8_1250, i_8_1281, i_8_1305, i_8_1307, i_8_1328, i_8_1345, i_8_1347, i_8_1449, i_8_1455, i_8_1456, i_8_1492, i_8_1534, i_8_1538, i_8_1579, i_8_1605, i_8_1606, i_8_1607, i_8_1608, i_8_1609, i_8_1644, i_8_1671, i_8_1706, i_8_1725, i_8_1726, i_8_1749, i_8_1763, i_8_1779, i_8_1823, i_8_1834, i_8_1870, i_8_1952, i_8_2012, i_8_2014, i_8_2050, i_8_2092, i_8_2129, i_8_2173, i_8_2199, i_8_2275, i_8_2293, i_8_2294, o_8_382);
	kernel_8_383 k_8_383(i_8_12, i_8_31, i_8_58, i_8_64, i_8_136, i_8_180, i_8_185, i_8_221, i_8_226, i_8_289, i_8_301, i_8_335, i_8_386, i_8_389, i_8_397, i_8_423, i_8_427, i_8_433, i_8_453, i_8_479, i_8_507, i_8_517, i_8_530, i_8_557, i_8_587, i_8_614, i_8_652, i_8_657, i_8_661, i_8_676, i_8_677, i_8_758, i_8_790, i_8_821, i_8_847, i_8_848, i_8_865, i_8_868, i_8_875, i_8_881, i_8_882, i_8_883, i_8_884, i_8_998, i_8_1049, i_8_1103, i_8_1106, i_8_1110, i_8_1115, i_8_1156, i_8_1199, i_8_1237, i_8_1255, i_8_1265, i_8_1286, i_8_1296, i_8_1298, i_8_1333, i_8_1340, i_8_1403, i_8_1408, i_8_1423, i_8_1435, i_8_1481, i_8_1507, i_8_1508, i_8_1539, i_8_1545, i_8_1558, i_8_1561, i_8_1581, i_8_1631, i_8_1642, i_8_1682, i_8_1683, i_8_1684, i_8_1737, i_8_1749, i_8_1750, i_8_1767, i_8_1771, i_8_1772, i_8_1778, i_8_1846, i_8_1881, i_8_1884, i_8_1885, i_8_1888, i_8_1947, i_8_1981, i_8_1992, i_8_2045, i_8_2098, i_8_2126, i_8_2170, i_8_2173, i_8_2268, i_8_2296, i_8_2297, i_8_2299, o_8_383);
	kernel_8_384 k_8_384(i_8_11, i_8_80, i_8_85, i_8_120, i_8_121, i_8_143, i_8_147, i_8_184, i_8_191, i_8_316, i_8_317, i_8_360, i_8_361, i_8_366, i_8_368, i_8_386, i_8_435, i_8_500, i_8_508, i_8_532, i_8_533, i_8_535, i_8_580, i_8_604, i_8_633, i_8_644, i_8_653, i_8_656, i_8_662, i_8_732, i_8_733, i_8_748, i_8_749, i_8_787, i_8_826, i_8_829, i_8_831, i_8_850, i_8_872, i_8_873, i_8_893, i_8_1037, i_8_1103, i_8_1138, i_8_1153, i_8_1202, i_8_1227, i_8_1240, i_8_1241, i_8_1244, i_8_1256, i_8_1319, i_8_1327, i_8_1336, i_8_1354, i_8_1364, i_8_1424, i_8_1456, i_8_1457, i_8_1462, i_8_1463, i_8_1471, i_8_1478, i_8_1493, i_8_1514, i_8_1522, i_8_1526, i_8_1540, i_8_1544, i_8_1570, i_8_1571, i_8_1591, i_8_1675, i_8_1696, i_8_1702, i_8_1703, i_8_1748, i_8_1766, i_8_1781, i_8_1783, i_8_1821, i_8_1844, i_8_1858, i_8_1882, i_8_1883, i_8_1892, i_8_1936, i_8_1954, i_8_1958, i_8_1975, i_8_1976, i_8_1985, i_8_1992, i_8_2044, i_8_2146, i_8_2155, i_8_2227, i_8_2231, i_8_2246, i_8_2257, o_8_384);
	kernel_8_385 k_8_385(i_8_20, i_8_35, i_8_85, i_8_94, i_8_224, i_8_264, i_8_269, i_8_323, i_8_356, i_8_370, i_8_445, i_8_453, i_8_460, i_8_506, i_8_538, i_8_554, i_8_556, i_8_565, i_8_620, i_8_647, i_8_658, i_8_662, i_8_698, i_8_708, i_8_718, i_8_721, i_8_733, i_8_734, i_8_779, i_8_793, i_8_843, i_8_923, i_8_935, i_8_950, i_8_953, i_8_977, i_8_988, i_8_989, i_8_994, i_8_997, i_8_998, i_8_1060, i_8_1105, i_8_1139, i_8_1183, i_8_1203, i_8_1234, i_8_1259, i_8_1260, i_8_1261, i_8_1268, i_8_1282, i_8_1283, i_8_1286, i_8_1319, i_8_1321, i_8_1325, i_8_1327, i_8_1328, i_8_1332, i_8_1366, i_8_1416, i_8_1418, i_8_1450, i_8_1452, i_8_1470, i_8_1481, i_8_1526, i_8_1532, i_8_1538, i_8_1553, i_8_1603, i_8_1604, i_8_1723, i_8_1754, i_8_1770, i_8_1771, i_8_1772, i_8_1788, i_8_1796, i_8_1813, i_8_1823, i_8_1931, i_8_1964, i_8_1983, i_8_1988, i_8_1989, i_8_2042, i_8_2067, i_8_2069, i_8_2077, i_8_2078, i_8_2113, i_8_2114, i_8_2136, i_8_2218, i_8_2226, i_8_2264, i_8_2294, i_8_2299, o_8_385);
	kernel_8_386 k_8_386(i_8_19, i_8_31, i_8_32, i_8_54, i_8_55, i_8_81, i_8_84, i_8_100, i_8_107, i_8_117, i_8_205, i_8_255, i_8_256, i_8_297, i_8_304, i_8_423, i_8_495, i_8_502, i_8_530, i_8_549, i_8_554, i_8_576, i_8_586, i_8_589, i_8_603, i_8_606, i_8_607, i_8_627, i_8_628, i_8_631, i_8_632, i_8_677, i_8_703, i_8_730, i_8_735, i_8_764, i_8_823, i_8_846, i_8_855, i_8_864, i_8_865, i_8_882, i_8_883, i_8_945, i_8_948, i_8_1033, i_8_1034, i_8_1062, i_8_1063, i_8_1111, i_8_1125, i_8_1134, i_8_1143, i_8_1144, i_8_1152, i_8_1171, i_8_1226, i_8_1233, i_8_1297, i_8_1299, i_8_1305, i_8_1332, i_8_1333, i_8_1403, i_8_1431, i_8_1432, i_8_1436, i_8_1467, i_8_1530, i_8_1543, i_8_1602, i_8_1615, i_8_1623, i_8_1631, i_8_1650, i_8_1652, i_8_1660, i_8_1693, i_8_1702, i_8_1710, i_8_1747, i_8_1755, i_8_1756, i_8_1762, i_8_1774, i_8_1776, i_8_1793, i_8_1809, i_8_1815, i_8_1872, i_8_1963, i_8_1980, i_8_2137, i_8_2143, i_8_2151, i_8_2196, i_8_2224, i_8_2234, i_8_2242, i_8_2245, o_8_386);
	kernel_8_387 k_8_387(i_8_14, i_8_30, i_8_98, i_8_102, i_8_103, i_8_107, i_8_114, i_8_216, i_8_223, i_8_297, i_8_300, i_8_345, i_8_361, i_8_362, i_8_365, i_8_367, i_8_391, i_8_418, i_8_444, i_8_453, i_8_525, i_8_530, i_8_535, i_8_546, i_8_552, i_8_589, i_8_591, i_8_607, i_8_609, i_8_630, i_8_637, i_8_659, i_8_665, i_8_694, i_8_697, i_8_723, i_8_738, i_8_780, i_8_781, i_8_786, i_8_822, i_8_842, i_8_874, i_8_894, i_8_958, i_8_970, i_8_987, i_8_1071, i_8_1107, i_8_1138, i_8_1145, i_8_1159, i_8_1204, i_8_1227, i_8_1228, i_8_1264, i_8_1279, i_8_1282, i_8_1285, i_8_1344, i_8_1426, i_8_1437, i_8_1438, i_8_1461, i_8_1525, i_8_1542, i_8_1552, i_8_1563, i_8_1564, i_8_1614, i_8_1635, i_8_1668, i_8_1681, i_8_1701, i_8_1719, i_8_1749, i_8_1761, i_8_1765, i_8_1773, i_8_1780, i_8_1782, i_8_1785, i_8_1786, i_8_1815, i_8_1843, i_8_2109, i_8_2110, i_8_2134, i_8_2139, i_8_2147, i_8_2157, i_8_2158, i_8_2184, i_8_2190, i_8_2215, i_8_2226, i_8_2232, i_8_2233, i_8_2265, i_8_2287, o_8_387);
	kernel_8_388 k_8_388(i_8_4, i_8_7, i_8_86, i_8_89, i_8_121, i_8_151, i_8_197, i_8_202, i_8_214, i_8_220, i_8_247, i_8_248, i_8_301, i_8_342, i_8_346, i_8_367, i_8_376, i_8_400, i_8_401, i_8_440, i_8_455, i_8_516, i_8_517, i_8_527, i_8_529, i_8_530, i_8_571, i_8_659, i_8_683, i_8_688, i_8_699, i_8_701, i_8_727, i_8_728, i_8_763, i_8_781, i_8_815, i_8_818, i_8_835, i_8_862, i_8_982, i_8_985, i_8_1003, i_8_1004, i_8_1045, i_8_1114, i_8_1153, i_8_1155, i_8_1157, i_8_1186, i_8_1281, i_8_1328, i_8_1330, i_8_1331, i_8_1342, i_8_1344, i_8_1358, i_8_1365, i_8_1434, i_8_1473, i_8_1474, i_8_1490, i_8_1535, i_8_1565, i_8_1610, i_8_1634, i_8_1642, i_8_1661, i_8_1662, i_8_1732, i_8_1733, i_8_1750, i_8_1753, i_8_1786, i_8_1787, i_8_1804, i_8_1806, i_8_1807, i_8_1840, i_8_1858, i_8_1861, i_8_1885, i_8_1975, i_8_1997, i_8_2011, i_8_2012, i_8_2032, i_8_2113, i_8_2120, i_8_2122, i_8_2123, i_8_2159, i_8_2174, i_8_2200, i_8_2215, i_8_2216, i_8_2225, i_8_2254, i_8_2289, i_8_2294, o_8_388);
	kernel_8_389 k_8_389(i_8_47, i_8_92, i_8_101, i_8_112, i_8_164, i_8_172, i_8_226, i_8_232, i_8_307, i_8_308, i_8_334, i_8_335, i_8_345, i_8_350, i_8_352, i_8_353, i_8_362, i_8_374, i_8_380, i_8_418, i_8_424, i_8_451, i_8_452, i_8_479, i_8_488, i_8_550, i_8_551, i_8_568, i_8_685, i_8_695, i_8_703, i_8_796, i_8_805, i_8_928, i_8_1018, i_8_1035, i_8_1054, i_8_1055, i_8_1057, i_8_1099, i_8_1100, i_8_1181, i_8_1229, i_8_1253, i_8_1274, i_8_1280, i_8_1289, i_8_1292, i_8_1297, i_8_1309, i_8_1315, i_8_1370, i_8_1378, i_8_1379, i_8_1381, i_8_1382, i_8_1408, i_8_1436, i_8_1443, i_8_1521, i_8_1549, i_8_1558, i_8_1559, i_8_1562, i_8_1603, i_8_1607, i_8_1624, i_8_1639, i_8_1640, i_8_1649, i_8_1650, i_8_1694, i_8_1702, i_8_1703, i_8_1752, i_8_1804, i_8_1820, i_8_1822, i_8_1829, i_8_1847, i_8_1855, i_8_1937, i_8_2002, i_8_2035, i_8_2036, i_8_2063, i_8_2072, i_8_2107, i_8_2143, i_8_2144, i_8_2152, i_8_2153, i_8_2197, i_8_2198, i_8_2207, i_8_2215, i_8_2225, i_8_2241, i_8_2245, i_8_2287, o_8_389);
	kernel_8_390 k_8_390(i_8_53, i_8_193, i_8_238, i_8_255, i_8_256, i_8_258, i_8_259, i_8_260, i_8_289, i_8_299, i_8_364, i_8_366, i_8_367, i_8_379, i_8_380, i_8_382, i_8_393, i_8_394, i_8_395, i_8_446, i_8_457, i_8_465, i_8_475, i_8_555, i_8_585, i_8_587, i_8_606, i_8_612, i_8_613, i_8_614, i_8_615, i_8_616, i_8_658, i_8_660, i_8_661, i_8_697, i_8_702, i_8_711, i_8_712, i_8_813, i_8_814, i_8_815, i_8_816, i_8_817, i_8_820, i_8_955, i_8_990, i_8_992, i_8_1026, i_8_1072, i_8_1074, i_8_1076, i_8_1077, i_8_1111, i_8_1112, i_8_1159, i_8_1230, i_8_1232, i_8_1260, i_8_1264, i_8_1268, i_8_1299, i_8_1455, i_8_1457, i_8_1491, i_8_1492, i_8_1539, i_8_1542, i_8_1543, i_8_1554, i_8_1601, i_8_1637, i_8_1650, i_8_1651, i_8_1652, i_8_1685, i_8_1700, i_8_1735, i_8_1779, i_8_1780, i_8_1896, i_8_1897, i_8_1898, i_8_1904, i_8_1915, i_8_2008, i_8_2031, i_8_2053, i_8_2077, i_8_2111, i_8_2127, i_8_2128, i_8_2130, i_8_2171, i_8_2187, i_8_2188, i_8_2189, i_8_2264, i_8_2267, i_8_2291, o_8_390);
	kernel_8_391 k_8_391(i_8_18, i_8_22, i_8_26, i_8_41, i_8_67, i_8_115, i_8_130, i_8_139, i_8_179, i_8_197, i_8_204, i_8_262, i_8_266, i_8_273, i_8_305, i_8_355, i_8_385, i_8_428, i_8_429, i_8_445, i_8_457, i_8_458, i_8_460, i_8_464, i_8_481, i_8_509, i_8_535, i_8_538, i_8_583, i_8_599, i_8_626, i_8_657, i_8_661, i_8_664, i_8_682, i_8_694, i_8_710, i_8_715, i_8_769, i_8_790, i_8_838, i_8_887, i_8_896, i_8_911, i_8_1041, i_8_1075, i_8_1076, i_8_1115, i_8_1133, i_8_1175, i_8_1192, i_8_1229, i_8_1232, i_8_1241, i_8_1296, i_8_1315, i_8_1318, i_8_1354, i_8_1386, i_8_1387, i_8_1395, i_8_1398, i_8_1399, i_8_1403, i_8_1407, i_8_1434, i_8_1436, i_8_1490, i_8_1494, i_8_1495, i_8_1498, i_8_1529, i_8_1634, i_8_1656, i_8_1702, i_8_1703, i_8_1706, i_8_1750, i_8_1768, i_8_1773, i_8_1795, i_8_1796, i_8_1819, i_8_1820, i_8_1826, i_8_1863, i_8_1919, i_8_1976, i_8_2007, i_8_2062, i_8_2138, i_8_2144, i_8_2147, i_8_2149, i_8_2216, i_8_2232, i_8_2237, i_8_2245, i_8_2246, i_8_2253, o_8_391);
	kernel_8_392 k_8_392(i_8_4, i_8_67, i_8_140, i_8_148, i_8_169, i_8_202, i_8_203, i_8_248, i_8_274, i_8_334, i_8_362, i_8_364, i_8_373, i_8_422, i_8_445, i_8_454, i_8_464, i_8_473, i_8_493, i_8_529, i_8_535, i_8_547, i_8_553, i_8_608, i_8_634, i_8_706, i_8_707, i_8_736, i_8_739, i_8_760, i_8_790, i_8_814, i_8_835, i_8_860, i_8_873, i_8_916, i_8_971, i_8_1067, i_8_1103, i_8_1114, i_8_1115, i_8_1129, i_8_1130, i_8_1201, i_8_1267, i_8_1301, i_8_1305, i_8_1306, i_8_1357, i_8_1399, i_8_1400, i_8_1407, i_8_1419, i_8_1435, i_8_1468, i_8_1489, i_8_1490, i_8_1492, i_8_1499, i_8_1546, i_8_1564, i_8_1573, i_8_1580, i_8_1595, i_8_1606, i_8_1633, i_8_1634, i_8_1705, i_8_1706, i_8_1729, i_8_1733, i_8_1774, i_8_1778, i_8_1782, i_8_1805, i_8_1810, i_8_1822, i_8_1823, i_8_1825, i_8_1826, i_8_1885, i_8_1886, i_8_1888, i_8_1904, i_8_1939, i_8_1981, i_8_1982, i_8_1985, i_8_2135, i_8_2145, i_8_2147, i_8_2150, i_8_2233, i_8_2249, i_8_2254, i_8_2258, i_8_2263, i_8_2266, i_8_2293, i_8_2299, o_8_392);
	kernel_8_393 k_8_393(i_8_4, i_8_9, i_8_24, i_8_40, i_8_43, i_8_53, i_8_70, i_8_85, i_8_94, i_8_104, i_8_141, i_8_157, i_8_159, i_8_160, i_8_192, i_8_241, i_8_265, i_8_293, i_8_346, i_8_355, i_8_371, i_8_391, i_8_394, i_8_417, i_8_418, i_8_420, i_8_421, i_8_427, i_8_428, i_8_433, i_8_481, i_8_483, i_8_493, i_8_535, i_8_553, i_8_557, i_8_605, i_8_608, i_8_627, i_8_628, i_8_633, i_8_662, i_8_672, i_8_704, i_8_709, i_8_769, i_8_825, i_8_849, i_8_850, i_8_922, i_8_938, i_8_943, i_8_951, i_8_968, i_8_976, i_8_991, i_8_1030, i_8_1113, i_8_1158, i_8_1201, i_8_1203, i_8_1258, i_8_1305, i_8_1307, i_8_1471, i_8_1489, i_8_1490, i_8_1534, i_8_1639, i_8_1654, i_8_1659, i_8_1671, i_8_1700, i_8_1702, i_8_1703, i_8_1704, i_8_1708, i_8_1729, i_8_1750, i_8_1781, i_8_1808, i_8_1819, i_8_1822, i_8_1824, i_8_1826, i_8_1974, i_8_1997, i_8_2001, i_8_2029, i_8_2047, i_8_2092, i_8_2146, i_8_2170, i_8_2182, i_8_2183, i_8_2214, i_8_2215, i_8_2247, i_8_2258, i_8_2281, o_8_393);
	kernel_8_394 k_8_394(i_8_15, i_8_23, i_8_43, i_8_66, i_8_79, i_8_98, i_8_118, i_8_169, i_8_191, i_8_257, i_8_265, i_8_266, i_8_268, i_8_282, i_8_283, i_8_287, i_8_296, i_8_299, i_8_338, i_8_340, i_8_382, i_8_430, i_8_454, i_8_456, i_8_491, i_8_492, i_8_493, i_8_502, i_8_529, i_8_530, i_8_583, i_8_588, i_8_592, i_8_615, i_8_628, i_8_672, i_8_673, i_8_690, i_8_693, i_8_711, i_8_716, i_8_718, i_8_719, i_8_750, i_8_769, i_8_770, i_8_772, i_8_789, i_8_795, i_8_822, i_8_842, i_8_843, i_8_845, i_8_880, i_8_894, i_8_954, i_8_1012, i_8_1021, i_8_1024, i_8_1033, i_8_1074, i_8_1078, i_8_1079, i_8_1087, i_8_1220, i_8_1242, i_8_1249, i_8_1254, i_8_1257, i_8_1258, i_8_1259, i_8_1267, i_8_1270, i_8_1295, i_8_1297, i_8_1310, i_8_1353, i_8_1417, i_8_1434, i_8_1457, i_8_1464, i_8_1617, i_8_1639, i_8_1650, i_8_1696, i_8_1704, i_8_1706, i_8_1728, i_8_1763, i_8_1927, i_8_1929, i_8_1936, i_8_2022, i_8_2023, i_8_2194, i_8_2195, i_8_2212, i_8_2262, i_8_2266, i_8_2281, o_8_394);
	kernel_8_395 k_8_395(i_8_5, i_8_69, i_8_78, i_8_79, i_8_88, i_8_114, i_8_159, i_8_204, i_8_205, i_8_206, i_8_249, i_8_251, i_8_277, i_8_278, i_8_286, i_8_305, i_8_332, i_8_348, i_8_349, i_8_350, i_8_355, i_8_358, i_8_363, i_8_393, i_8_404, i_8_422, i_8_445, i_8_446, i_8_519, i_8_528, i_8_555, i_8_592, i_8_601, i_8_602, i_8_615, i_8_618, i_8_619, i_8_696, i_8_706, i_8_726, i_8_762, i_8_818, i_8_836, i_8_840, i_8_845, i_8_849, i_8_868, i_8_880, i_8_918, i_8_951, i_8_961, i_8_1015, i_8_1060, i_8_1075, i_8_1086, i_8_1087, i_8_1088, i_8_1115, i_8_1178, i_8_1203, i_8_1258, i_8_1284, i_8_1286, i_8_1328, i_8_1410, i_8_1438, i_8_1456, i_8_1457, i_8_1502, i_8_1543, i_8_1591, i_8_1592, i_8_1617, i_8_1661, i_8_1749, i_8_1752, i_8_1753, i_8_1772, i_8_1797, i_8_1799, i_8_1808, i_8_1815, i_8_1816, i_8_1835, i_8_1853, i_8_1896, i_8_1897, i_8_1941, i_8_1969, i_8_1978, i_8_2004, i_8_2013, i_8_2014, i_8_2058, i_8_2059, i_8_2069, i_8_2152, i_8_2193, i_8_2194, i_8_2218, o_8_395);
	kernel_8_396 k_8_396(i_8_43, i_8_55, i_8_61, i_8_96, i_8_106, i_8_121, i_8_142, i_8_249, i_8_255, i_8_295, i_8_300, i_8_301, i_8_321, i_8_328, i_8_330, i_8_340, i_8_367, i_8_429, i_8_436, i_8_439, i_8_440, i_8_457, i_8_460, i_8_484, i_8_486, i_8_489, i_8_492, i_8_588, i_8_593, i_8_618, i_8_624, i_8_627, i_8_635, i_8_661, i_8_664, i_8_672, i_8_708, i_8_717, i_8_736, i_8_768, i_8_807, i_8_808, i_8_835, i_8_840, i_8_845, i_8_873, i_8_970, i_8_979, i_8_993, i_8_1104, i_8_1105, i_8_1115, i_8_1152, i_8_1183, i_8_1228, i_8_1239, i_8_1258, i_8_1270, i_8_1354, i_8_1357, i_8_1393, i_8_1401, i_8_1428, i_8_1440, i_8_1447, i_8_1545, i_8_1588, i_8_1591, i_8_1681, i_8_1701, i_8_1705, i_8_1752, i_8_1754, i_8_1767, i_8_1768, i_8_1770, i_8_1777, i_8_1788, i_8_1789, i_8_1824, i_8_1825, i_8_1854, i_8_1857, i_8_1858, i_8_1861, i_8_1907, i_8_1942, i_8_1990, i_8_1995, i_8_2028, i_8_2031, i_8_2058, i_8_2091, i_8_2100, i_8_2109, i_8_2131, i_8_2133, i_8_2193, i_8_2194, i_8_2278, o_8_396);
	kernel_8_397 k_8_397(i_8_22, i_8_79, i_8_142, i_8_196, i_8_229, i_8_232, i_8_266, i_8_309, i_8_312, i_8_348, i_8_366, i_8_385, i_8_401, i_8_489, i_8_571, i_8_572, i_8_582, i_8_589, i_8_606, i_8_625, i_8_654, i_8_655, i_8_679, i_8_696, i_8_697, i_8_698, i_8_699, i_8_700, i_8_701, i_8_705, i_8_708, i_8_733, i_8_751, i_8_835, i_8_840, i_8_843, i_8_864, i_8_880, i_8_886, i_8_966, i_8_968, i_8_1041, i_8_1049, i_8_1093, i_8_1132, i_8_1147, i_8_1148, i_8_1168, i_8_1227, i_8_1230, i_8_1231, i_8_1267, i_8_1305, i_8_1317, i_8_1318, i_8_1357, i_8_1358, i_8_1373, i_8_1375, i_8_1390, i_8_1405, i_8_1449, i_8_1491, i_8_1492, i_8_1525, i_8_1543, i_8_1552, i_8_1599, i_8_1600, i_8_1624, i_8_1641, i_8_1642, i_8_1654, i_8_1655, i_8_1663, i_8_1751, i_8_1779, i_8_1780, i_8_1824, i_8_1825, i_8_1857, i_8_1860, i_8_1874, i_8_1904, i_8_1929, i_8_1939, i_8_1982, i_8_1992, i_8_2075, i_8_2086, i_8_2092, i_8_2093, i_8_2149, i_8_2152, i_8_2167, i_8_2174, i_8_2233, i_8_2244, i_8_2257, i_8_2273, o_8_397);
	kernel_8_398 k_8_398(i_8_19, i_8_109, i_8_139, i_8_238, i_8_300, i_8_310, i_8_372, i_8_373, i_8_375, i_8_381, i_8_383, i_8_419, i_8_431, i_8_460, i_8_463, i_8_479, i_8_480, i_8_506, i_8_510, i_8_529, i_8_549, i_8_552, i_8_553, i_8_590, i_8_603, i_8_606, i_8_613, i_8_706, i_8_796, i_8_858, i_8_867, i_8_868, i_8_878, i_8_976, i_8_991, i_8_1030, i_8_1084, i_8_1127, i_8_1130, i_8_1158, i_8_1188, i_8_1189, i_8_1192, i_8_1255, i_8_1279, i_8_1283, i_8_1325, i_8_1326, i_8_1327, i_8_1480, i_8_1507, i_8_1524, i_8_1533, i_8_1534, i_8_1535, i_8_1596, i_8_1597, i_8_1605, i_8_1606, i_8_1616, i_8_1660, i_8_1676, i_8_1681, i_8_1701, i_8_1733, i_8_1746, i_8_1779, i_8_1781, i_8_1782, i_8_1789, i_8_1790, i_8_1805, i_8_1806, i_8_1815, i_8_1821, i_8_1836, i_8_1837, i_8_1840, i_8_1844, i_8_1864, i_8_1891, i_8_1894, i_8_1901, i_8_1917, i_8_1919, i_8_1921, i_8_1951, i_8_1965, i_8_2053, i_8_2117, i_8_2127, i_8_2128, i_8_2169, i_8_2176, i_8_2179, i_8_2232, i_8_2244, i_8_2294, i_8_2297, i_8_2303, o_8_398);
	kernel_8_399 k_8_399(i_8_27, i_8_33, i_8_34, i_8_35, i_8_61, i_8_62, i_8_79, i_8_80, i_8_140, i_8_187, i_8_191, i_8_239, i_8_256, i_8_269, i_8_296, i_8_347, i_8_349, i_8_350, i_8_401, i_8_482, i_8_507, i_8_524, i_8_554, i_8_615, i_8_633, i_8_637, i_8_638, i_8_700, i_8_701, i_8_705, i_8_706, i_8_714, i_8_754, i_8_850, i_8_861, i_8_862, i_8_880, i_8_887, i_8_888, i_8_889, i_8_890, i_8_944, i_8_991, i_8_992, i_8_995, i_8_1016, i_8_1028, i_8_1050, i_8_1057, i_8_1060, i_8_1106, i_8_1131, i_8_1132, i_8_1157, i_8_1186, i_8_1187, i_8_1267, i_8_1268, i_8_1286, i_8_1297, i_8_1303, i_8_1322, i_8_1400, i_8_1483, i_8_1504, i_8_1505, i_8_1543, i_8_1545, i_8_1553, i_8_1556, i_8_1591, i_8_1648, i_8_1650, i_8_1690, i_8_1697, i_8_1751, i_8_1760, i_8_1762, i_8_1763, i_8_1857, i_8_1859, i_8_1886, i_8_1888, i_8_1898, i_8_1904, i_8_1949, i_8_1970, i_8_1985, i_8_1991, i_8_2015, i_8_2137, i_8_2146, i_8_2150, i_8_2159, i_8_2219, i_8_2241, i_8_2243, i_8_2248, i_8_2249, i_8_2263, o_8_399);
	kernel_8_400 k_8_400(i_8_9, i_8_12, i_8_20, i_8_50, i_8_74, i_8_101, i_8_140, i_8_149, i_8_165, i_8_254, i_8_290, i_8_299, i_8_304, i_8_362, i_8_364, i_8_379, i_8_380, i_8_423, i_8_424, i_8_490, i_8_554, i_8_578, i_8_582, i_8_583, i_8_598, i_8_605, i_8_640, i_8_650, i_8_653, i_8_677, i_8_679, i_8_695, i_8_697, i_8_731, i_8_775, i_8_776, i_8_787, i_8_794, i_8_803, i_8_842, i_8_850, i_8_878, i_8_883, i_8_936, i_8_965, i_8_971, i_8_1037, i_8_1199, i_8_1231, i_8_1255, i_8_1271, i_8_1282, i_8_1299, i_8_1313, i_8_1316, i_8_1339, i_8_1345, i_8_1378, i_8_1397, i_8_1433, i_8_1457, i_8_1471, i_8_1538, i_8_1557, i_8_1571, i_8_1607, i_8_1622, i_8_1629, i_8_1703, i_8_1715, i_8_1750, i_8_1755, i_8_1756, i_8_1768, i_8_1777, i_8_1791, i_8_1818, i_8_1819, i_8_1823, i_8_1832, i_8_1888, i_8_1973, i_8_1981, i_8_1993, i_8_2052, i_8_2054, i_8_2072, i_8_2099, i_8_2106, i_8_2108, i_8_2135, i_8_2143, i_8_2155, i_8_2170, i_8_2188, i_8_2230, i_8_2243, i_8_2264, i_8_2295, i_8_2298, o_8_400);
	kernel_8_401 k_8_401(i_8_30, i_8_31, i_8_84, i_8_88, i_8_111, i_8_114, i_8_165, i_8_238, i_8_240, i_8_372, i_8_386, i_8_390, i_8_421, i_8_427, i_8_437, i_8_474, i_8_475, i_8_483, i_8_520, i_8_522, i_8_540, i_8_553, i_8_571, i_8_574, i_8_598, i_8_606, i_8_633, i_8_693, i_8_694, i_8_706, i_8_709, i_8_712, i_8_759, i_8_762, i_8_763, i_8_778, i_8_799, i_8_839, i_8_888, i_8_940, i_8_943, i_8_966, i_8_994, i_8_1056, i_8_1059, i_8_1090, i_8_1102, i_8_1182, i_8_1185, i_8_1281, i_8_1293, i_8_1300, i_8_1305, i_8_1309, i_8_1318, i_8_1345, i_8_1390, i_8_1438, i_8_1516, i_8_1533, i_8_1534, i_8_1563, i_8_1590, i_8_1603, i_8_1614, i_8_1624, i_8_1654, i_8_1686, i_8_1690, i_8_1731, i_8_1735, i_8_1747, i_8_1749, i_8_1751, i_8_1753, i_8_1762, i_8_1780, i_8_1789, i_8_1804, i_8_1824, i_8_1825, i_8_1831, i_8_1917, i_8_1929, i_8_1996, i_8_2019, i_8_2047, i_8_2058, i_8_2077, i_8_2118, i_8_2122, i_8_2124, i_8_2142, i_8_2150, i_8_2173, i_8_2224, i_8_2260, i_8_2290, i_8_2295, i_8_2299, o_8_401);
	kernel_8_402 k_8_402(i_8_55, i_8_78, i_8_95, i_8_97, i_8_105, i_8_106, i_8_107, i_8_141, i_8_220, i_8_223, i_8_228, i_8_229, i_8_256, i_8_276, i_8_379, i_8_492, i_8_573, i_8_580, i_8_583, i_8_597, i_8_636, i_8_658, i_8_661, i_8_663, i_8_664, i_8_672, i_8_700, i_8_704, i_8_733, i_8_763, i_8_781, i_8_822, i_8_858, i_8_861, i_8_871, i_8_894, i_8_925, i_8_969, i_8_975, i_8_976, i_8_1107, i_8_1108, i_8_1122, i_8_1228, i_8_1237, i_8_1272, i_8_1302, i_8_1322, i_8_1348, i_8_1393, i_8_1470, i_8_1473, i_8_1479, i_8_1483, i_8_1506, i_8_1509, i_8_1524, i_8_1561, i_8_1563, i_8_1606, i_8_1617, i_8_1618, i_8_1620, i_8_1677, i_8_1700, i_8_1702, i_8_1704, i_8_1750, i_8_1771, i_8_1785, i_8_1786, i_8_1810, i_8_1812, i_8_1833, i_8_1842, i_8_1866, i_8_1878, i_8_1885, i_8_1947, i_8_1949, i_8_1962, i_8_1965, i_8_1968, i_8_1974, i_8_1983, i_8_1986, i_8_1988, i_8_1992, i_8_2055, i_8_2112, i_8_2148, i_8_2154, i_8_2172, i_8_2175, i_8_2185, i_8_2188, i_8_2202, i_8_2229, i_8_2262, i_8_2278, o_8_402);
	kernel_8_403 k_8_403(i_8_25, i_8_39, i_8_51, i_8_66, i_8_67, i_8_143, i_8_195, i_8_219, i_8_228, i_8_230, i_8_267, i_8_269, i_8_286, i_8_287, i_8_313, i_8_402, i_8_403, i_8_423, i_8_467, i_8_492, i_8_522, i_8_526, i_8_527, i_8_551, i_8_582, i_8_583, i_8_588, i_8_619, i_8_652, i_8_654, i_8_665, i_8_703, i_8_726, i_8_807, i_8_823, i_8_840, i_8_843, i_8_844, i_8_876, i_8_883, i_8_886, i_8_897, i_8_898, i_8_922, i_8_924, i_8_930, i_8_931, i_8_933, i_8_964, i_8_978, i_8_979, i_8_980, i_8_1030, i_8_1074, i_8_1276, i_8_1307, i_8_1428, i_8_1429, i_8_1438, i_8_1446, i_8_1447, i_8_1455, i_8_1534, i_8_1535, i_8_1599, i_8_1624, i_8_1632, i_8_1671, i_8_1672, i_8_1725, i_8_1733, i_8_1744, i_8_1748, i_8_1773, i_8_1774, i_8_1803, i_8_1857, i_8_1903, i_8_1941, i_8_1950, i_8_1962, i_8_1968, i_8_1969, i_8_2004, i_8_2100, i_8_2104, i_8_2143, i_8_2158, i_8_2172, i_8_2174, i_8_2175, i_8_2176, i_8_2177, i_8_2209, i_8_2233, i_8_2245, i_8_2262, i_8_2263, i_8_2265, i_8_2271, o_8_403);
	kernel_8_404 k_8_404(i_8_25, i_8_31, i_8_35, i_8_86, i_8_160, i_8_188, i_8_205, i_8_295, i_8_296, i_8_332, i_8_377, i_8_457, i_8_463, i_8_483, i_8_484, i_8_502, i_8_508, i_8_528, i_8_529, i_8_539, i_8_553, i_8_556, i_8_626, i_8_629, i_8_636, i_8_664, i_8_692, i_8_716, i_8_718, i_8_719, i_8_727, i_8_735, i_8_760, i_8_762, i_8_769, i_8_772, i_8_870, i_8_871, i_8_880, i_8_897, i_8_926, i_8_951, i_8_978, i_8_988, i_8_989, i_8_993, i_8_994, i_8_995, i_8_1032, i_8_1033, i_8_1034, i_8_1093, i_8_1113, i_8_1114, i_8_1203, i_8_1230, i_8_1239, i_8_1293, i_8_1330, i_8_1347, i_8_1407, i_8_1452, i_8_1482, i_8_1484, i_8_1509, i_8_1528, i_8_1529, i_8_1601, i_8_1618, i_8_1680, i_8_1705, i_8_1708, i_8_1716, i_8_1717, i_8_1718, i_8_1730, i_8_1735, i_8_1743, i_8_1762, i_8_1778, i_8_1784, i_8_1798, i_8_1808, i_8_1822, i_8_1905, i_8_1920, i_8_1929, i_8_1933, i_8_1969, i_8_1985, i_8_2013, i_8_2015, i_8_2029, i_8_2113, i_8_2140, i_8_2145, i_8_2146, i_8_2191, i_8_2230, i_8_2272, o_8_404);
	kernel_8_405 k_8_405(i_8_1, i_8_2, i_8_82, i_8_83, i_8_95, i_8_101, i_8_104, i_8_154, i_8_221, i_8_244, i_8_281, i_8_289, i_8_290, i_8_292, i_8_293, i_8_326, i_8_342, i_8_343, i_8_363, i_8_382, i_8_401, i_8_419, i_8_434, i_8_437, i_8_440, i_8_454, i_8_478, i_8_479, i_8_545, i_8_585, i_8_607, i_8_608, i_8_613, i_8_622, i_8_623, i_8_625, i_8_631, i_8_659, i_8_666, i_8_667, i_8_682, i_8_703, i_8_704, i_8_713, i_8_721, i_8_722, i_8_776, i_8_784, i_8_796, i_8_823, i_8_830, i_8_832, i_8_833, i_8_838, i_8_843, i_8_868, i_8_968, i_8_974, i_8_977, i_8_1031, i_8_1040, i_8_1049, i_8_1112, i_8_1161, i_8_1180, i_8_1181, i_8_1208, i_8_1238, i_8_1265, i_8_1298, i_8_1355, i_8_1373, i_8_1388, i_8_1435, i_8_1547, i_8_1565, i_8_1576, i_8_1585, i_8_1586, i_8_1679, i_8_1750, i_8_1783, i_8_1801, i_8_1807, i_8_1855, i_8_1858, i_8_1876, i_8_1900, i_8_1904, i_8_1985, i_8_1991, i_8_1992, i_8_1994, i_8_2036, i_8_2093, i_8_2110, i_8_2143, i_8_2146, i_8_2182, i_8_2279, o_8_405);
	kernel_8_406 k_8_406(i_8_3, i_8_23, i_8_51, i_8_52, i_8_58, i_8_68, i_8_97, i_8_98, i_8_140, i_8_142, i_8_160, i_8_219, i_8_241, i_8_247, i_8_304, i_8_311, i_8_328, i_8_329, i_8_346, i_8_347, i_8_388, i_8_437, i_8_440, i_8_507, i_8_528, i_8_555, i_8_580, i_8_599, i_8_600, i_8_606, i_8_608, i_8_610, i_8_634, i_8_642, i_8_655, i_8_705, i_8_706, i_8_709, i_8_716, i_8_723, i_8_724, i_8_760, i_8_813, i_8_814, i_8_815, i_8_836, i_8_840, i_8_875, i_8_970, i_8_971, i_8_1034, i_8_1050, i_8_1051, i_8_1071, i_8_1114, i_8_1241, i_8_1281, i_8_1292, i_8_1305, i_8_1306, i_8_1316, i_8_1355, i_8_1389, i_8_1391, i_8_1407, i_8_1409, i_8_1410, i_8_1411, i_8_1471, i_8_1507, i_8_1531, i_8_1570, i_8_1573, i_8_1574, i_8_1642, i_8_1653, i_8_1664, i_8_1678, i_8_1679, i_8_1719, i_8_1731, i_8_1760, i_8_1784, i_8_1820, i_8_1887, i_8_1948, i_8_1963, i_8_1983, i_8_1997, i_8_2028, i_8_2031, i_8_2056, i_8_2057, i_8_2109, i_8_2151, i_8_2154, i_8_2156, i_8_2190, i_8_2216, i_8_2282, o_8_406);
	kernel_8_407 k_8_407(i_8_22, i_8_34, i_8_52, i_8_53, i_8_58, i_8_69, i_8_94, i_8_97, i_8_103, i_8_106, i_8_107, i_8_135, i_8_214, i_8_223, i_8_224, i_8_241, i_8_255, i_8_256, i_8_257, i_8_304, i_8_429, i_8_453, i_8_454, i_8_507, i_8_527, i_8_586, i_8_598, i_8_606, i_8_607, i_8_633, i_8_658, i_8_660, i_8_661, i_8_663, i_8_664, i_8_678, i_8_679, i_8_688, i_8_736, i_8_766, i_8_782, i_8_825, i_8_850, i_8_868, i_8_871, i_8_922, i_8_969, i_8_990, i_8_1051, i_8_1060, i_8_1066, i_8_1071, i_8_1137, i_8_1138, i_8_1268, i_8_1351, i_8_1431, i_8_1444, i_8_1453, i_8_1454, i_8_1490, i_8_1533, i_8_1535, i_8_1549, i_8_1561, i_8_1564, i_8_1596, i_8_1614, i_8_1618, i_8_1633, i_8_1713, i_8_1714, i_8_1742, i_8_1750, i_8_1813, i_8_1839, i_8_1840, i_8_1841, i_8_1860, i_8_1884, i_8_1887, i_8_1893, i_8_1894, i_8_1904, i_8_1969, i_8_1987, i_8_2002, i_8_2005, i_8_2077, i_8_2111, i_8_2127, i_8_2129, i_8_2131, i_8_2137, i_8_2200, i_8_2215, i_8_2227, i_8_2236, i_8_2260, i_8_2263, o_8_407);
	kernel_8_408 k_8_408(i_8_21, i_8_76, i_8_84, i_8_91, i_8_159, i_8_224, i_8_325, i_8_329, i_8_345, i_8_367, i_8_381, i_8_382, i_8_384, i_8_390, i_8_391, i_8_399, i_8_462, i_8_463, i_8_478, i_8_483, i_8_484, i_8_501, i_8_525, i_8_526, i_8_529, i_8_621, i_8_669, i_8_673, i_8_685, i_8_753, i_8_759, i_8_760, i_8_768, i_8_823, i_8_827, i_8_840, i_8_841, i_8_892, i_8_992, i_8_1031, i_8_1075, i_8_1159, i_8_1191, i_8_1204, i_8_1218, i_8_1249, i_8_1254, i_8_1255, i_8_1272, i_8_1273, i_8_1274, i_8_1281, i_8_1303, i_8_1326, i_8_1358, i_8_1401, i_8_1402, i_8_1470, i_8_1506, i_8_1539, i_8_1542, i_8_1554, i_8_1587, i_8_1597, i_8_1600, i_8_1605, i_8_1633, i_8_1647, i_8_1680, i_8_1720, i_8_1741, i_8_1761, i_8_1762, i_8_1803, i_8_1807, i_8_1821, i_8_1839, i_8_1866, i_8_1867, i_8_1875, i_8_1893, i_8_1899, i_8_1917, i_8_1918, i_8_1921, i_8_1947, i_8_1950, i_8_1965, i_8_1967, i_8_2030, i_8_2033, i_8_2049, i_8_2088, i_8_2110, i_8_2150, i_8_2181, i_8_2190, i_8_2191, i_8_2215, i_8_2229, o_8_408);
	kernel_8_409 k_8_409(i_8_9, i_8_12, i_8_33, i_8_61, i_8_63, i_8_72, i_8_75, i_8_135, i_8_180, i_8_181, i_8_208, i_8_279, i_8_318, i_8_397, i_8_399, i_8_417, i_8_426, i_8_427, i_8_450, i_8_453, i_8_495, i_8_504, i_8_525, i_8_528, i_8_535, i_8_570, i_8_573, i_8_579, i_8_585, i_8_589, i_8_658, i_8_660, i_8_661, i_8_662, i_8_702, i_8_748, i_8_751, i_8_777, i_8_783, i_8_797, i_8_822, i_8_829, i_8_838, i_8_841, i_8_858, i_8_865, i_8_867, i_8_877, i_8_973, i_8_1101, i_8_1107, i_8_1152, i_8_1153, i_8_1198, i_8_1293, i_8_1294, i_8_1314, i_8_1326, i_8_1332, i_8_1354, i_8_1355, i_8_1363, i_8_1395, i_8_1398, i_8_1422, i_8_1425, i_8_1440, i_8_1467, i_8_1480, i_8_1515, i_8_1521, i_8_1522, i_8_1539, i_8_1551, i_8_1611, i_8_1629, i_8_1689, i_8_1701, i_8_1705, i_8_1746, i_8_1764, i_8_1791, i_8_1794, i_8_1803, i_8_1818, i_8_1822, i_8_1836, i_8_1837, i_8_1891, i_8_1956, i_8_1974, i_8_1992, i_8_1996, i_8_2008, i_8_2052, i_8_2133, i_8_2147, i_8_2223, i_8_2243, i_8_2273, o_8_409);
	kernel_8_410 k_8_410(i_8_4, i_8_21, i_8_24, i_8_53, i_8_89, i_8_115, i_8_175, i_8_188, i_8_193, i_8_255, i_8_256, i_8_277, i_8_310, i_8_313, i_8_336, i_8_355, i_8_356, i_8_364, i_8_463, i_8_516, i_8_517, i_8_571, i_8_580, i_8_604, i_8_615, i_8_616, i_8_617, i_8_652, i_8_669, i_8_671, i_8_678, i_8_697, i_8_708, i_8_815, i_8_831, i_8_832, i_8_840, i_8_842, i_8_846, i_8_991, i_8_1057, i_8_1126, i_8_1131, i_8_1156, i_8_1159, i_8_1173, i_8_1183, i_8_1201, i_8_1237, i_8_1273, i_8_1284, i_8_1285, i_8_1305, i_8_1306, i_8_1336, i_8_1353, i_8_1393, i_8_1470, i_8_1490, i_8_1498, i_8_1499, i_8_1525, i_8_1526, i_8_1534, i_8_1597, i_8_1629, i_8_1653, i_8_1659, i_8_1660, i_8_1696, i_8_1697, i_8_1724, i_8_1746, i_8_1771, i_8_1780, i_8_1802, i_8_1806, i_8_1807, i_8_1808, i_8_1825, i_8_1857, i_8_1858, i_8_1866, i_8_1876, i_8_1906, i_8_1919, i_8_1949, i_8_1969, i_8_1974, i_8_2038, i_8_2047, i_8_2048, i_8_2050, i_8_2066, i_8_2092, i_8_2108, i_8_2137, i_8_2147, i_8_2154, i_8_2257, o_8_410);
	kernel_8_411 k_8_411(i_8_18, i_8_96, i_8_106, i_8_196, i_8_222, i_8_225, i_8_258, i_8_348, i_8_364, i_8_365, i_8_421, i_8_439, i_8_486, i_8_610, i_8_627, i_8_635, i_8_648, i_8_651, i_8_654, i_8_664, i_8_682, i_8_693, i_8_697, i_8_700, i_8_706, i_8_708, i_8_726, i_8_729, i_8_732, i_8_733, i_8_747, i_8_751, i_8_769, i_8_777, i_8_842, i_8_874, i_8_876, i_8_877, i_8_880, i_8_882, i_8_967, i_8_969, i_8_981, i_8_984, i_8_990, i_8_996, i_8_1030, i_8_1128, i_8_1173, i_8_1174, i_8_1224, i_8_1372, i_8_1410, i_8_1470, i_8_1483, i_8_1527, i_8_1530, i_8_1533, i_8_1540, i_8_1542, i_8_1546, i_8_1548, i_8_1555, i_8_1624, i_8_1642, i_8_1659, i_8_1663, i_8_1683, i_8_1686, i_8_1691, i_8_1696, i_8_1701, i_8_1705, i_8_1725, i_8_1734, i_8_1759, i_8_1767, i_8_1809, i_8_1812, i_8_1824, i_8_1855, i_8_1885, i_8_1962, i_8_1965, i_8_1986, i_8_1995, i_8_2007, i_8_2070, i_8_2083, i_8_2088, i_8_2091, i_8_2104, i_8_2146, i_8_2223, i_8_2236, i_8_2242, i_8_2247, i_8_2253, i_8_2254, i_8_2262, o_8_411);
	kernel_8_412 k_8_412(i_8_59, i_8_60, i_8_105, i_8_107, i_8_108, i_8_184, i_8_225, i_8_226, i_8_228, i_8_229, i_8_258, i_8_285, i_8_337, i_8_349, i_8_367, i_8_393, i_8_484, i_8_485, i_8_504, i_8_505, i_8_526, i_8_592, i_8_600, i_8_602, i_8_630, i_8_701, i_8_750, i_8_780, i_8_850, i_8_851, i_8_876, i_8_879, i_8_882, i_8_1013, i_8_1016, i_8_1032, i_8_1102, i_8_1138, i_8_1155, i_8_1203, i_8_1231, i_8_1237, i_8_1238, i_8_1240, i_8_1241, i_8_1261, i_8_1274, i_8_1311, i_8_1314, i_8_1315, i_8_1317, i_8_1322, i_8_1326, i_8_1331, i_8_1353, i_8_1354, i_8_1361, i_8_1479, i_8_1484, i_8_1490, i_8_1542, i_8_1548, i_8_1551, i_8_1552, i_8_1553, i_8_1556, i_8_1653, i_8_1689, i_8_1691, i_8_1697, i_8_1701, i_8_1708, i_8_1713, i_8_1715, i_8_1716, i_8_1717, i_8_1726, i_8_1813, i_8_1814, i_8_1816, i_8_1825, i_8_1859, i_8_1884, i_8_1885, i_8_1887, i_8_1888, i_8_1938, i_8_1939, i_8_1940, i_8_1941, i_8_1980, i_8_1995, i_8_2053, i_8_2115, i_8_2140, i_8_2169, i_8_2170, i_8_2287, i_8_2290, i_8_2301, o_8_412);
	kernel_8_413 k_8_413(i_8_17, i_8_20, i_8_41, i_8_89, i_8_113, i_8_167, i_8_197, i_8_201, i_8_233, i_8_242, i_8_248, i_8_347, i_8_352, i_8_361, i_8_362, i_8_365, i_8_374, i_8_386, i_8_427, i_8_441, i_8_454, i_8_488, i_8_524, i_8_527, i_8_581, i_8_595, i_8_609, i_8_652, i_8_657, i_8_659, i_8_676, i_8_677, i_8_693, i_8_698, i_8_703, i_8_709, i_8_729, i_8_734, i_8_761, i_8_764, i_8_778, i_8_833, i_8_835, i_8_838, i_8_839, i_8_848, i_8_850, i_8_862, i_8_869, i_8_878, i_8_881, i_8_887, i_8_941, i_8_959, i_8_1075, i_8_1076, i_8_1118, i_8_1136, i_8_1193, i_8_1237, i_8_1262, i_8_1283, i_8_1325, i_8_1342, i_8_1357, i_8_1411, i_8_1414, i_8_1474, i_8_1477, i_8_1478, i_8_1526, i_8_1534, i_8_1543, i_8_1552, i_8_1589, i_8_1603, i_8_1612, i_8_1625, i_8_1631, i_8_1697, i_8_1712, i_8_1736, i_8_1741, i_8_1742, i_8_1863, i_8_1886, i_8_1889, i_8_1895, i_8_1901, i_8_1964, i_8_1982, i_8_1985, i_8_2007, i_8_2011, i_8_2075, i_8_2077, i_8_2134, i_8_2147, i_8_2150, i_8_2156, o_8_413);
	kernel_8_414 k_8_414(i_8_3, i_8_4, i_8_27, i_8_44, i_8_51, i_8_57, i_8_75, i_8_117, i_8_165, i_8_168, i_8_192, i_8_193, i_8_221, i_8_255, i_8_265, i_8_282, i_8_292, i_8_300, i_8_337, i_8_339, i_8_346, i_8_363, i_8_364, i_8_366, i_8_368, i_8_381, i_8_382, i_8_417, i_8_436, i_8_439, i_8_455, i_8_479, i_8_480, i_8_523, i_8_525, i_8_526, i_8_528, i_8_595, i_8_615, i_8_624, i_8_633, i_8_642, i_8_661, i_8_665, i_8_672, i_8_678, i_8_694, i_8_705, i_8_715, i_8_723, i_8_759, i_8_804, i_8_837, i_8_840, i_8_841, i_8_844, i_8_876, i_8_966, i_8_969, i_8_971, i_8_1072, i_8_1074, i_8_1182, i_8_1199, i_8_1227, i_8_1231, i_8_1254, i_8_1263, i_8_1301, i_8_1305, i_8_1336, i_8_1357, i_8_1551, i_8_1570, i_8_1574, i_8_1587, i_8_1623, i_8_1624, i_8_1641, i_8_1644, i_8_1677, i_8_1717, i_8_1731, i_8_1749, i_8_1807, i_8_1830, i_8_1857, i_8_1866, i_8_1903, i_8_1992, i_8_1995, i_8_2028, i_8_2036, i_8_2056, i_8_2090, i_8_2133, i_8_2190, i_8_2194, i_8_2293, i_8_2301, o_8_414);
	kernel_8_415 k_8_415(i_8_13, i_8_38, i_8_40, i_8_75, i_8_113, i_8_135, i_8_193, i_8_226, i_8_262, i_8_264, i_8_308, i_8_320, i_8_361, i_8_362, i_8_422, i_8_490, i_8_509, i_8_514, i_8_520, i_8_535, i_8_543, i_8_544, i_8_580, i_8_604, i_8_612, i_8_613, i_8_634, i_8_653, i_8_656, i_8_748, i_8_751, i_8_756, i_8_766, i_8_800, i_8_802, i_8_815, i_8_837, i_8_881, i_8_896, i_8_937, i_8_967, i_8_968, i_8_974, i_8_1071, i_8_1085, i_8_1102, i_8_1117, i_8_1163, i_8_1228, i_8_1253, i_8_1260, i_8_1262, i_8_1270, i_8_1273, i_8_1295, i_8_1432, i_8_1463, i_8_1495, i_8_1496, i_8_1498, i_8_1514, i_8_1516, i_8_1519, i_8_1526, i_8_1531, i_8_1596, i_8_1638, i_8_1651, i_8_1676, i_8_1682, i_8_1688, i_8_1694, i_8_1702, i_8_1729, i_8_1747, i_8_1760, i_8_1769, i_8_1773, i_8_1784, i_8_1819, i_8_1822, i_8_1837, i_8_1873, i_8_1881, i_8_1884, i_8_1891, i_8_1912, i_8_1927, i_8_1939, i_8_1965, i_8_1971, i_8_1980, i_8_2017, i_8_2054, i_8_2072, i_8_2146, i_8_2152, i_8_2244, i_8_2246, i_8_2270, o_8_415);
	kernel_8_416 k_8_416(i_8_27, i_8_31, i_8_34, i_8_96, i_8_97, i_8_114, i_8_115, i_8_116, i_8_166, i_8_184, i_8_224, i_8_241, i_8_300, i_8_303, i_8_367, i_8_369, i_8_381, i_8_382, i_8_421, i_8_492, i_8_508, i_8_525, i_8_572, i_8_588, i_8_616, i_8_633, i_8_634, i_8_662, i_8_701, i_8_703, i_8_704, i_8_706, i_8_707, i_8_714, i_8_754, i_8_778, i_8_859, i_8_887, i_8_940, i_8_941, i_8_994, i_8_1030, i_8_1096, i_8_1113, i_8_1114, i_8_1120, i_8_1159, i_8_1182, i_8_1183, i_8_1186, i_8_1188, i_8_1197, i_8_1284, i_8_1292, i_8_1299, i_8_1307, i_8_1308, i_8_1330, i_8_1411, i_8_1412, i_8_1437, i_8_1535, i_8_1545, i_8_1551, i_8_1591, i_8_1635, i_8_1642, i_8_1654, i_8_1678, i_8_1684, i_8_1696, i_8_1731, i_8_1741, i_8_1742, i_8_1744, i_8_1751, i_8_1762, i_8_1785, i_8_1821, i_8_1825, i_8_1831, i_8_1858, i_8_1939, i_8_2047, i_8_2050, i_8_2075, i_8_2119, i_8_2122, i_8_2123, i_8_2153, i_8_2157, i_8_2172, i_8_2189, i_8_2214, i_8_2215, i_8_2217, i_8_2218, i_8_2245, i_8_2248, i_8_2303, o_8_416);
	kernel_8_417 k_8_417(i_8_12, i_8_52, i_8_114, i_8_193, i_8_220, i_8_226, i_8_279, i_8_318, i_8_319, i_8_321, i_8_365, i_8_397, i_8_399, i_8_400, i_8_402, i_8_427, i_8_428, i_8_440, i_8_471, i_8_490, i_8_492, i_8_525, i_8_582, i_8_583, i_8_584, i_8_612, i_8_639, i_8_642, i_8_645, i_8_646, i_8_660, i_8_748, i_8_759, i_8_762, i_8_799, i_8_808, i_8_843, i_8_844, i_8_852, i_8_855, i_8_877, i_8_933, i_8_934, i_8_966, i_8_967, i_8_1179, i_8_1228, i_8_1240, i_8_1257, i_8_1263, i_8_1281, i_8_1284, i_8_1285, i_8_1303, i_8_1307, i_8_1318, i_8_1330, i_8_1359, i_8_1366, i_8_1435, i_8_1438, i_8_1440, i_8_1443, i_8_1456, i_8_1461, i_8_1464, i_8_1470, i_8_1493, i_8_1559, i_8_1564, i_8_1662, i_8_1677, i_8_1713, i_8_1717, i_8_1756, i_8_1876, i_8_1893, i_8_1935, i_8_1939, i_8_1966, i_8_1997, i_8_2041, i_8_2057, i_8_2091, i_8_2134, i_8_2146, i_8_2147, i_8_2149, i_8_2154, i_8_2170, i_8_2171, i_8_2173, i_8_2174, i_8_2175, i_8_2177, i_8_2185, i_8_2193, i_8_2194, i_8_2216, i_8_2232, o_8_417);
	kernel_8_418 k_8_418(i_8_21, i_8_30, i_8_139, i_8_140, i_8_184, i_8_193, i_8_229, i_8_246, i_8_247, i_8_262, i_8_274, i_8_292, i_8_356, i_8_373, i_8_417, i_8_420, i_8_430, i_8_461, i_8_462, i_8_463, i_8_474, i_8_517, i_8_529, i_8_557, i_8_571, i_8_612, i_8_615, i_8_634, i_8_671, i_8_678, i_8_681, i_8_703, i_8_715, i_8_730, i_8_761, i_8_792, i_8_793, i_8_795, i_8_837, i_8_849, i_8_880, i_8_959, i_8_993, i_8_996, i_8_997, i_8_1081, i_8_1114, i_8_1157, i_8_1159, i_8_1192, i_8_1236, i_8_1237, i_8_1259, i_8_1270, i_8_1274, i_8_1281, i_8_1283, i_8_1284, i_8_1300, i_8_1307, i_8_1326, i_8_1387, i_8_1468, i_8_1483, i_8_1493, i_8_1539, i_8_1542, i_8_1546, i_8_1597, i_8_1598, i_8_1659, i_8_1731, i_8_1752, i_8_1776, i_8_1785, i_8_1803, i_8_1804, i_8_1812, i_8_1818, i_8_1820, i_8_1855, i_8_1867, i_8_1874, i_8_1876, i_8_1894, i_8_1912, i_8_1918, i_8_1919, i_8_1997, i_8_2007, i_8_2045, i_8_2065, i_8_2093, i_8_2109, i_8_2137, i_8_2158, i_8_2192, i_8_2254, i_8_2257, i_8_2291, o_8_418);
	kernel_8_419 k_8_419(i_8_44, i_8_93, i_8_95, i_8_131, i_8_174, i_8_175, i_8_185, i_8_223, i_8_241, i_8_264, i_8_276, i_8_282, i_8_302, i_8_309, i_8_310, i_8_312, i_8_314, i_8_338, i_8_391, i_8_430, i_8_527, i_8_591, i_8_592, i_8_593, i_8_607, i_8_617, i_8_626, i_8_655, i_8_661, i_8_663, i_8_664, i_8_692, i_8_822, i_8_826, i_8_827, i_8_838, i_8_955, i_8_959, i_8_969, i_8_970, i_8_996, i_8_1003, i_8_1047, i_8_1049, i_8_1060, i_8_1061, i_8_1092, i_8_1110, i_8_1159, i_8_1191, i_8_1192, i_8_1193, i_8_1236, i_8_1263, i_8_1264, i_8_1265, i_8_1278, i_8_1279, i_8_1280, i_8_1282, i_8_1300, i_8_1306, i_8_1308, i_8_1366, i_8_1410, i_8_1411, i_8_1412, i_8_1434, i_8_1435, i_8_1436, i_8_1471, i_8_1641, i_8_1643, i_8_1644, i_8_1645, i_8_1646, i_8_1653, i_8_1655, i_8_1662, i_8_1663, i_8_1664, i_8_1715, i_8_1819, i_8_1877, i_8_1899, i_8_1964, i_8_2073, i_8_2093, i_8_2135, i_8_2136, i_8_2141, i_8_2164, i_8_2175, i_8_2193, i_8_2215, i_8_2216, i_8_2219, i_8_2263, i_8_2264, i_8_2290, o_8_419);
	kernel_8_420 k_8_420(i_8_22, i_8_34, i_8_47, i_8_50, i_8_61, i_8_154, i_8_161, i_8_208, i_8_211, i_8_212, i_8_214, i_8_290, i_8_293, i_8_296, i_8_335, i_8_391, i_8_424, i_8_425, i_8_451, i_8_452, i_8_463, i_8_658, i_8_662, i_8_673, i_8_704, i_8_749, i_8_828, i_8_829, i_8_923, i_8_952, i_8_955, i_8_1027, i_8_1036, i_8_1135, i_8_1136, i_8_1138, i_8_1139, i_8_1225, i_8_1233, i_8_1272, i_8_1276, i_8_1286, i_8_1351, i_8_1354, i_8_1355, i_8_1357, i_8_1358, i_8_1361, i_8_1469, i_8_1486, i_8_1487, i_8_1506, i_8_1532, i_8_1533, i_8_1535, i_8_1544, i_8_1550, i_8_1558, i_8_1559, i_8_1603, i_8_1604, i_8_1702, i_8_1711, i_8_1714, i_8_1715, i_8_1719, i_8_1720, i_8_1821, i_8_1861, i_8_1881, i_8_1886, i_8_1895, i_8_1944, i_8_1985, i_8_1993, i_8_2002, i_8_2003, i_8_2005, i_8_2006, i_8_2045, i_8_2053, i_8_2117, i_8_2129, i_8_2142, i_8_2146, i_8_2153, i_8_2154, i_8_2179, i_8_2188, i_8_2191, i_8_2200, i_8_2210, i_8_2225, i_8_2227, i_8_2246, i_8_2260, i_8_2261, i_8_2263, i_8_2264, i_8_2273, o_8_420);
	kernel_8_421 k_8_421(i_8_34, i_8_76, i_8_91, i_8_95, i_8_154, i_8_234, i_8_252, i_8_305, i_8_334, i_8_337, i_8_352, i_8_353, i_8_365, i_8_371, i_8_443, i_8_469, i_8_492, i_8_496, i_8_497, i_8_499, i_8_526, i_8_527, i_8_557, i_8_586, i_8_589, i_8_602, i_8_609, i_8_613, i_8_614, i_8_631, i_8_634, i_8_659, i_8_691, i_8_703, i_8_706, i_8_760, i_8_775, i_8_799, i_8_812, i_8_833, i_8_836, i_8_841, i_8_842, i_8_844, i_8_866, i_8_896, i_8_902, i_8_932, i_8_946, i_8_947, i_8_958, i_8_967, i_8_982, i_8_1057, i_8_1058, i_8_1225, i_8_1229, i_8_1247, i_8_1292, i_8_1318, i_8_1322, i_8_1349, i_8_1435, i_8_1436, i_8_1468, i_8_1485, i_8_1525, i_8_1538, i_8_1543, i_8_1553, i_8_1654, i_8_1655, i_8_1682, i_8_1723, i_8_1729, i_8_1733, i_8_1753, i_8_1784, i_8_1786, i_8_1787, i_8_1822, i_8_1871, i_8_1886, i_8_1972, i_8_1984, i_8_1992, i_8_1993, i_8_2005, i_8_2044, i_8_2125, i_8_2143, i_8_2144, i_8_2146, i_8_2147, i_8_2155, i_8_2200, i_8_2224, i_8_2245, i_8_2289, i_8_2294, o_8_421);
	kernel_8_422 k_8_422(i_8_38, i_8_47, i_8_55, i_8_64, i_8_65, i_8_73, i_8_77, i_8_107, i_8_127, i_8_140, i_8_236, i_8_262, i_8_263, i_8_309, i_8_312, i_8_319, i_8_344, i_8_360, i_8_371, i_8_373, i_8_374, i_8_388, i_8_389, i_8_398, i_8_416, i_8_419, i_8_424, i_8_451, i_8_457, i_8_529, i_8_533, i_8_545, i_8_559, i_8_577, i_8_580, i_8_589, i_8_610, i_8_632, i_8_693, i_8_694, i_8_698, i_8_702, i_8_721, i_8_749, i_8_782, i_8_838, i_8_866, i_8_929, i_8_967, i_8_968, i_8_973, i_8_978, i_8_1081, i_8_1127, i_8_1153, i_8_1172, i_8_1198, i_8_1234, i_8_1235, i_8_1279, i_8_1298, i_8_1315, i_8_1336, i_8_1351, i_8_1366, i_8_1379, i_8_1398, i_8_1406, i_8_1414, i_8_1442, i_8_1462, i_8_1468, i_8_1469, i_8_1487, i_8_1514, i_8_1605, i_8_1669, i_8_1684, i_8_1685, i_8_1688, i_8_1712, i_8_1777, i_8_1793, i_8_1801, i_8_1819, i_8_1820, i_8_1821, i_8_1837, i_8_1883, i_8_1910, i_8_1936, i_8_1939, i_8_1990, i_8_2005, i_8_2032, i_8_2059, i_8_2072, i_8_2189, i_8_2265, i_8_2296, o_8_422);
	kernel_8_423 k_8_423(i_8_89, i_8_166, i_8_194, i_8_195, i_8_197, i_8_260, i_8_314, i_8_381, i_8_384, i_8_385, i_8_386, i_8_451, i_8_458, i_8_485, i_8_539, i_8_556, i_8_575, i_8_598, i_8_602, i_8_607, i_8_611, i_8_619, i_8_633, i_8_635, i_8_662, i_8_670, i_8_716, i_8_736, i_8_751, i_8_754, i_8_835, i_8_841, i_8_844, i_8_863, i_8_877, i_8_986, i_8_994, i_8_1039, i_8_1040, i_8_1042, i_8_1043, i_8_1051, i_8_1052, i_8_1074, i_8_1079, i_8_1106, i_8_1177, i_8_1227, i_8_1229, i_8_1231, i_8_1236, i_8_1262, i_8_1263, i_8_1264, i_8_1284, i_8_1294, i_8_1302, i_8_1402, i_8_1412, i_8_1475, i_8_1484, i_8_1493, i_8_1528, i_8_1529, i_8_1561, i_8_1562, i_8_1655, i_8_1663, i_8_1677, i_8_1679, i_8_1682, i_8_1689, i_8_1700, i_8_1724, i_8_1727, i_8_1751, i_8_1752, i_8_1771, i_8_1790, i_8_1807, i_8_1816, i_8_1825, i_8_1867, i_8_1871, i_8_1880, i_8_1888, i_8_1889, i_8_1967, i_8_1995, i_8_2014, i_8_2074, i_8_2075, i_8_2129, i_8_2132, i_8_2143, i_8_2195, i_8_2210, i_8_2239, i_8_2248, i_8_2249, o_8_423);
	kernel_8_424 k_8_424(i_8_36, i_8_41, i_8_67, i_8_72, i_8_73, i_8_74, i_8_76, i_8_104, i_8_136, i_8_173, i_8_220, i_8_244, i_8_304, i_8_352, i_8_353, i_8_356, i_8_361, i_8_365, i_8_389, i_8_426, i_8_427, i_8_470, i_8_490, i_8_505, i_8_514, i_8_515, i_8_526, i_8_527, i_8_569, i_8_582, i_8_587, i_8_596, i_8_603, i_8_611, i_8_623, i_8_676, i_8_679, i_8_748, i_8_757, i_8_793, i_8_826, i_8_829, i_8_847, i_8_866, i_8_911, i_8_1127, i_8_1161, i_8_1172, i_8_1199, i_8_1250, i_8_1316, i_8_1378, i_8_1397, i_8_1404, i_8_1468, i_8_1495, i_8_1531, i_8_1533, i_8_1534, i_8_1537, i_8_1538, i_8_1595, i_8_1639, i_8_1648, i_8_1657, i_8_1682, i_8_1694, i_8_1701, i_8_1706, i_8_1743, i_8_1754, i_8_1764, i_8_1802, i_8_1810, i_8_1838, i_8_1843, i_8_1846, i_8_1886, i_8_1909, i_8_1910, i_8_1948, i_8_1970, i_8_1972, i_8_1991, i_8_2063, i_8_2064, i_8_2093, i_8_2142, i_8_2144, i_8_2147, i_8_2150, i_8_2206, i_8_2242, i_8_2254, i_8_2255, i_8_2256, i_8_2273, i_8_2282, i_8_2293, i_8_2296, o_8_424);
	kernel_8_425 k_8_425(i_8_7, i_8_8, i_8_11, i_8_76, i_8_79, i_8_89, i_8_121, i_8_169, i_8_227, i_8_269, i_8_296, i_8_322, i_8_332, i_8_364, i_8_365, i_8_366, i_8_368, i_8_379, i_8_383, i_8_421, i_8_429, i_8_448, i_8_455, i_8_484, i_8_491, i_8_492, i_8_493, i_8_599, i_8_605, i_8_629, i_8_647, i_8_658, i_8_661, i_8_664, i_8_670, i_8_683, i_8_696, i_8_698, i_8_719, i_8_727, i_8_748, i_8_771, i_8_815, i_8_818, i_8_827, i_8_893, i_8_977, i_8_996, i_8_998, i_8_1025, i_8_1078, i_8_1126, i_8_1127, i_8_1186, i_8_1214, i_8_1241, i_8_1294, i_8_1301, i_8_1309, i_8_1318, i_8_1325, i_8_1358, i_8_1366, i_8_1388, i_8_1391, i_8_1394, i_8_1410, i_8_1411, i_8_1430, i_8_1591, i_8_1627, i_8_1628, i_8_1649, i_8_1655, i_8_1675, i_8_1679, i_8_1689, i_8_1699, i_8_1771, i_8_1779, i_8_1784, i_8_1807, i_8_1852, i_8_1862, i_8_1907, i_8_1954, i_8_1988, i_8_2032, i_8_2060, i_8_2089, i_8_2092, i_8_2122, i_8_2146, i_8_2149, i_8_2152, i_8_2153, i_8_2175, i_8_2180, i_8_2195, i_8_2219, o_8_425);
	kernel_8_426 k_8_426(i_8_21, i_8_48, i_8_78, i_8_106, i_8_114, i_8_115, i_8_143, i_8_157, i_8_190, i_8_265, i_8_288, i_8_366, i_8_381, i_8_400, i_8_452, i_8_454, i_8_469, i_8_508, i_8_527, i_8_550, i_8_554, i_8_557, i_8_579, i_8_581, i_8_583, i_8_584, i_8_601, i_8_633, i_8_634, i_8_642, i_8_643, i_8_653, i_8_660, i_8_662, i_8_679, i_8_680, i_8_683, i_8_702, i_8_710, i_8_720, i_8_751, i_8_754, i_8_819, i_8_826, i_8_827, i_8_851, i_8_868, i_8_895, i_8_940, i_8_961, i_8_971, i_8_993, i_8_1013, i_8_1039, i_8_1041, i_8_1115, i_8_1137, i_8_1146, i_8_1149, i_8_1198, i_8_1229, i_8_1236, i_8_1263, i_8_1267, i_8_1295, i_8_1300, i_8_1398, i_8_1431, i_8_1435, i_8_1436, i_8_1437, i_8_1463, i_8_1465, i_8_1470, i_8_1489, i_8_1491, i_8_1560, i_8_1679, i_8_1702, i_8_1750, i_8_1759, i_8_1767, i_8_1769, i_8_1774, i_8_1783, i_8_1795, i_8_1829, i_8_1837, i_8_1939, i_8_1947, i_8_1957, i_8_1983, i_8_2036, i_8_2055, i_8_2110, i_8_2134, i_8_2226, i_8_2235, i_8_2246, i_8_2263, o_8_426);
	kernel_8_427 k_8_427(i_8_8, i_8_29, i_8_34, i_8_44, i_8_94, i_8_115, i_8_130, i_8_190, i_8_194, i_8_203, i_8_206, i_8_230, i_8_247, i_8_259, i_8_262, i_8_275, i_8_278, i_8_292, i_8_311, i_8_325, i_8_429, i_8_430, i_8_445, i_8_453, i_8_454, i_8_462, i_8_475, i_8_528, i_8_552, i_8_588, i_8_607, i_8_608, i_8_661, i_8_664, i_8_673, i_8_681, i_8_704, i_8_761, i_8_792, i_8_844, i_8_959, i_8_968, i_8_972, i_8_1087, i_8_1102, i_8_1112, i_8_1131, i_8_1132, i_8_1134, i_8_1159, i_8_1175, i_8_1231, i_8_1274, i_8_1312, i_8_1346, i_8_1370, i_8_1383, i_8_1385, i_8_1392, i_8_1407, i_8_1426, i_8_1482, i_8_1498, i_8_1534, i_8_1537, i_8_1553, i_8_1597, i_8_1598, i_8_1601, i_8_1615, i_8_1642, i_8_1645, i_8_1687, i_8_1748, i_8_1769, i_8_1770, i_8_1777, i_8_1779, i_8_1836, i_8_1842, i_8_1849, i_8_1852, i_8_1873, i_8_1877, i_8_1886, i_8_1887, i_8_1894, i_8_1919, i_8_1969, i_8_1983, i_8_1985, i_8_2024, i_8_2069, i_8_2084, i_8_2174, i_8_2177, i_8_2183, i_8_2191, i_8_2258, i_8_2275, o_8_427);
	kernel_8_428 k_8_428(i_8_20, i_8_22, i_8_23, i_8_24, i_8_40, i_8_52, i_8_67, i_8_91, i_8_114, i_8_142, i_8_175, i_8_193, i_8_200, i_8_244, i_8_273, i_8_274, i_8_356, i_8_365, i_8_368, i_8_382, i_8_385, i_8_430, i_8_468, i_8_469, i_8_571, i_8_599, i_8_651, i_8_703, i_8_706, i_8_707, i_8_730, i_8_751, i_8_814, i_8_853, i_8_856, i_8_883, i_8_955, i_8_1053, i_8_1066, i_8_1102, i_8_1105, i_8_1111, i_8_1123, i_8_1182, i_8_1228, i_8_1303, i_8_1343, i_8_1351, i_8_1390, i_8_1391, i_8_1400, i_8_1414, i_8_1453, i_8_1470, i_8_1473, i_8_1510, i_8_1542, i_8_1606, i_8_1633, i_8_1638, i_8_1642, i_8_1650, i_8_1653, i_8_1687, i_8_1694, i_8_1705, i_8_1732, i_8_1764, i_8_1771, i_8_1807, i_8_1808, i_8_1821, i_8_1873, i_8_1881, i_8_1882, i_8_1906, i_8_1913, i_8_1918, i_8_1939, i_8_1942, i_8_1949, i_8_1990, i_8_1991, i_8_2011, i_8_2065, i_8_2088, i_8_2091, i_8_2112, i_8_2120, i_8_2149, i_8_2153, i_8_2182, i_8_2183, i_8_2206, i_8_2207, i_8_2223, i_8_2233, i_8_2244, i_8_2272, i_8_2302, o_8_428);
	kernel_8_429 k_8_429(i_8_30, i_8_33, i_8_34, i_8_36, i_8_39, i_8_63, i_8_75, i_8_87, i_8_126, i_8_172, i_8_175, i_8_180, i_8_210, i_8_220, i_8_227, i_8_237, i_8_256, i_8_301, i_8_306, i_8_309, i_8_328, i_8_336, i_8_351, i_8_378, i_8_451, i_8_472, i_8_489, i_8_490, i_8_525, i_8_550, i_8_579, i_8_589, i_8_606, i_8_607, i_8_610, i_8_624, i_8_634, i_8_660, i_8_664, i_8_694, i_8_705, i_8_760, i_8_768, i_8_843, i_8_883, i_8_886, i_8_921, i_8_924, i_8_954, i_8_967, i_8_970, i_8_985, i_8_990, i_8_1026, i_8_1032, i_8_1056, i_8_1089, i_8_1170, i_8_1188, i_8_1227, i_8_1228, i_8_1233, i_8_1254, i_8_1275, i_8_1301, i_8_1329, i_8_1345, i_8_1371, i_8_1380, i_8_1461, i_8_1541, i_8_1557, i_8_1560, i_8_1638, i_8_1650, i_8_1671, i_8_1677, i_8_1701, i_8_1704, i_8_1749, i_8_1751, i_8_1768, i_8_1774, i_8_1780, i_8_1803, i_8_1827, i_8_1863, i_8_1888, i_8_1905, i_8_1906, i_8_2108, i_8_2133, i_8_2154, i_8_2158, i_8_2163, i_8_2178, i_8_2181, i_8_2245, i_8_2272, i_8_2289, o_8_429);
	kernel_8_430 k_8_430(i_8_3, i_8_28, i_8_33, i_8_36, i_8_57, i_8_94, i_8_106, i_8_168, i_8_224, i_8_259, i_8_323, i_8_361, i_8_390, i_8_470, i_8_498, i_8_507, i_8_523, i_8_582, i_8_597, i_8_607, i_8_642, i_8_651, i_8_654, i_8_659, i_8_678, i_8_681, i_8_751, i_8_786, i_8_845, i_8_861, i_8_870, i_8_871, i_8_885, i_8_940, i_8_1013, i_8_1038, i_8_1039, i_8_1084, i_8_1111, i_8_1114, i_8_1128, i_8_1129, i_8_1159, i_8_1182, i_8_1194, i_8_1258, i_8_1266, i_8_1272, i_8_1317, i_8_1338, i_8_1395, i_8_1410, i_8_1425, i_8_1434, i_8_1437, i_8_1438, i_8_1448, i_8_1464, i_8_1471, i_8_1483, i_8_1489, i_8_1492, i_8_1515, i_8_1516, i_8_1548, i_8_1551, i_8_1605, i_8_1623, i_8_1633, i_8_1683, i_8_1716, i_8_1722, i_8_1752, i_8_1759, i_8_1768, i_8_1794, i_8_1803, i_8_1812, i_8_1822, i_8_1824, i_8_1839, i_8_1840, i_8_1855, i_8_1881, i_8_1888, i_8_1938, i_8_1947, i_8_1965, i_8_1984, i_8_1987, i_8_2133, i_8_2147, i_8_2148, i_8_2154, i_8_2157, i_8_2158, i_8_2229, i_8_2233, i_8_2246, i_8_2248, o_8_430);
	kernel_8_431 k_8_431(i_8_115, i_8_143, i_8_169, i_8_191, i_8_260, i_8_296, i_8_311, i_8_316, i_8_395, i_8_459, i_8_466, i_8_467, i_8_484, i_8_485, i_8_494, i_8_511, i_8_520, i_8_523, i_8_526, i_8_527, i_8_528, i_8_529, i_8_537, i_8_557, i_8_664, i_8_715, i_8_718, i_8_719, i_8_763, i_8_764, i_8_771, i_8_772, i_8_782, i_8_835, i_8_844, i_8_869, i_8_915, i_8_949, i_8_959, i_8_967, i_8_1040, i_8_1050, i_8_1114, i_8_1124, i_8_1223, i_8_1267, i_8_1277, i_8_1283, i_8_1308, i_8_1309, i_8_1319, i_8_1328, i_8_1330, i_8_1331, i_8_1346, i_8_1392, i_8_1402, i_8_1439, i_8_1447, i_8_1493, i_8_1501, i_8_1534, i_8_1537, i_8_1538, i_8_1555, i_8_1600, i_8_1601, i_8_1633, i_8_1651, i_8_1681, i_8_1682, i_8_1723, i_8_1732, i_8_1735, i_8_1768, i_8_1771, i_8_1796, i_8_1799, i_8_1825, i_8_1843, i_8_1871, i_8_1886, i_8_1916, i_8_1920, i_8_1921, i_8_1950, i_8_1979, i_8_1995, i_8_2014, i_8_2015, i_8_2032, i_8_2068, i_8_2095, i_8_2114, i_8_2122, i_8_2185, i_8_2218, i_8_2240, i_8_2247, i_8_2302, o_8_431);
	kernel_8_432 k_8_432(i_8_52, i_8_57, i_8_84, i_8_141, i_8_142, i_8_143, i_8_192, i_8_225, i_8_255, i_8_328, i_8_370, i_8_373, i_8_382, i_8_417, i_8_480, i_8_481, i_8_483, i_8_484, i_8_500, i_8_507, i_8_510, i_8_522, i_8_526, i_8_528, i_8_530, i_8_544, i_8_596, i_8_602, i_8_610, i_8_651, i_8_656, i_8_661, i_8_702, i_8_759, i_8_760, i_8_763, i_8_777, i_8_778, i_8_789, i_8_796, i_8_813, i_8_814, i_8_836, i_8_842, i_8_871, i_8_879, i_8_904, i_8_949, i_8_993, i_8_1011, i_8_1016, i_8_1050, i_8_1074, i_8_1135, i_8_1177, i_8_1272, i_8_1284, i_8_1305, i_8_1306, i_8_1344, i_8_1348, i_8_1349, i_8_1357, i_8_1419, i_8_1437, i_8_1506, i_8_1527, i_8_1544, i_8_1545, i_8_1547, i_8_1573, i_8_1630, i_8_1633, i_8_1644, i_8_1668, i_8_1677, i_8_1679, i_8_1682, i_8_1710, i_8_1714, i_8_1717, i_8_1718, i_8_1722, i_8_1726, i_8_1732, i_8_1753, i_8_1867, i_8_1868, i_8_1906, i_8_1950, i_8_1997, i_8_2028, i_8_2101, i_8_2104, i_8_2128, i_8_2130, i_8_2131, i_8_2214, i_8_2215, i_8_2216, o_8_432);
	kernel_8_433 k_8_433(i_8_30, i_8_49, i_8_81, i_8_106, i_8_138, i_8_141, i_8_142, i_8_183, i_8_255, i_8_256, i_8_328, i_8_352, i_8_355, i_8_374, i_8_418, i_8_442, i_8_445, i_8_450, i_8_453, i_8_481, i_8_494, i_8_497, i_8_547, i_8_616, i_8_663, i_8_691, i_8_702, i_8_703, i_8_706, i_8_736, i_8_765, i_8_786, i_8_811, i_8_814, i_8_815, i_8_819, i_8_828, i_8_848, i_8_867, i_8_868, i_8_869, i_8_895, i_8_922, i_8_949, i_8_950, i_8_953, i_8_969, i_8_972, i_8_973, i_8_976, i_8_982, i_8_984, i_8_994, i_8_1011, i_8_1027, i_8_1074, i_8_1134, i_8_1155, i_8_1267, i_8_1273, i_8_1305, i_8_1325, i_8_1336, i_8_1342, i_8_1442, i_8_1468, i_8_1525, i_8_1559, i_8_1564, i_8_1617, i_8_1713, i_8_1714, i_8_1717, i_8_1726, i_8_1731, i_8_1732, i_8_1750, i_8_1753, i_8_1754, i_8_1786, i_8_1789, i_8_1802, i_8_1812, i_8_1813, i_8_1864, i_8_1903, i_8_1904, i_8_1930, i_8_1952, i_8_2007, i_8_2010, i_8_2011, i_8_2068, i_8_2069, i_8_2093, i_8_2131, i_8_2136, i_8_2214, i_8_2215, i_8_2244, o_8_433);
	kernel_8_434 k_8_434(i_8_48, i_8_49, i_8_66, i_8_67, i_8_72, i_8_78, i_8_93, i_8_107, i_8_114, i_8_130, i_8_138, i_8_166, i_8_174, i_8_178, i_8_183, i_8_191, i_8_237, i_8_304, i_8_321, i_8_334, i_8_336, i_8_337, i_8_361, i_8_381, i_8_382, i_8_399, i_8_400, i_8_579, i_8_607, i_8_608, i_8_642, i_8_651, i_8_693, i_8_694, i_8_705, i_8_729, i_8_795, i_8_831, i_8_864, i_8_882, i_8_930, i_8_954, i_8_969, i_8_1020, i_8_1092, i_8_1093, i_8_1128, i_8_1255, i_8_1263, i_8_1287, i_8_1300, i_8_1306, i_8_1311, i_8_1314, i_8_1317, i_8_1354, i_8_1388, i_8_1400, i_8_1448, i_8_1469, i_8_1493, i_8_1524, i_8_1527, i_8_1545, i_8_1560, i_8_1686, i_8_1687, i_8_1704, i_8_1706, i_8_1749, i_8_1821, i_8_1825, i_8_1830, i_8_1840, i_8_1846, i_8_1848, i_8_1851, i_8_1855, i_8_1869, i_8_1893, i_8_1938, i_8_1993, i_8_1995, i_8_2038, i_8_2040, i_8_2041, i_8_2056, i_8_2077, i_8_2145, i_8_2154, i_8_2155, i_8_2157, i_8_2181, i_8_2199, i_8_2200, i_8_2202, i_8_2220, i_8_2246, i_8_2275, i_8_2299, o_8_434);
	kernel_8_435 k_8_435(i_8_18, i_8_31, i_8_32, i_8_154, i_8_208, i_8_220, i_8_289, i_8_326, i_8_370, i_8_371, i_8_373, i_8_374, i_8_426, i_8_445, i_8_473, i_8_478, i_8_485, i_8_496, i_8_522, i_8_524, i_8_578, i_8_586, i_8_604, i_8_610, i_8_611, i_8_625, i_8_631, i_8_657, i_8_667, i_8_668, i_8_671, i_8_711, i_8_712, i_8_713, i_8_757, i_8_776, i_8_783, i_8_787, i_8_792, i_8_793, i_8_821, i_8_855, i_8_892, i_8_938, i_8_947, i_8_1112, i_8_1127, i_8_1130, i_8_1216, i_8_1225, i_8_1246, i_8_1247, i_8_1252, i_8_1260, i_8_1264, i_8_1279, i_8_1280, i_8_1297, i_8_1317, i_8_1318, i_8_1323, i_8_1431, i_8_1434, i_8_1450, i_8_1451, i_8_1503, i_8_1504, i_8_1505, i_8_1522, i_8_1585, i_8_1586, i_8_1595, i_8_1631, i_8_1634, i_8_1666, i_8_1681, i_8_1696, i_8_1713, i_8_1739, i_8_1752, i_8_1753, i_8_1759, i_8_1776, i_8_1802, i_8_1824, i_8_1837, i_8_1854, i_8_1856, i_8_1890, i_8_1891, i_8_1948, i_8_1965, i_8_2047, i_8_2125, i_8_2126, i_8_2147, i_8_2189, i_8_2245, i_8_2270, i_8_2286, o_8_435);
	kernel_8_436 k_8_436(i_8_18, i_8_48, i_8_78, i_8_117, i_8_141, i_8_142, i_8_219, i_8_259, i_8_310, i_8_322, i_8_336, i_8_345, i_8_346, i_8_348, i_8_360, i_8_363, i_8_367, i_8_378, i_8_381, i_8_400, i_8_402, i_8_417, i_8_427, i_8_454, i_8_493, i_8_499, i_8_579, i_8_603, i_8_615, i_8_643, i_8_654, i_8_658, i_8_660, i_8_675, i_8_696, i_8_702, i_8_750, i_8_795, i_8_799, i_8_849, i_8_873, i_8_889, i_8_991, i_8_1020, i_8_1056, i_8_1059, i_8_1092, i_8_1104, i_8_1115, i_8_1146, i_8_1152, i_8_1158, i_8_1266, i_8_1283, i_8_1284, i_8_1291, i_8_1314, i_8_1323, i_8_1383, i_8_1426, i_8_1439, i_8_1440, i_8_1444, i_8_1473, i_8_1597, i_8_1602, i_8_1633, i_8_1644, i_8_1671, i_8_1688, i_8_1699, i_8_1702, i_8_1704, i_8_1723, i_8_1749, i_8_1753, i_8_1803, i_8_1818, i_8_1830, i_8_1836, i_8_1840, i_8_1857, i_8_1885, i_8_1887, i_8_1899, i_8_1944, i_8_1947, i_8_1980, i_8_1981, i_8_2004, i_8_2184, i_8_2223, i_8_2227, i_8_2229, i_8_2238, i_8_2247, i_8_2248, i_8_2271, i_8_2277, i_8_2287, o_8_436);
	kernel_8_437 k_8_437(i_8_9, i_8_58, i_8_86, i_8_136, i_8_138, i_8_139, i_8_165, i_8_223, i_8_363, i_8_370, i_8_374, i_8_375, i_8_385, i_8_417, i_8_468, i_8_480, i_8_499, i_8_507, i_8_527, i_8_529, i_8_547, i_8_554, i_8_597, i_8_624, i_8_625, i_8_715, i_8_716, i_8_760, i_8_761, i_8_762, i_8_769, i_8_868, i_8_873, i_8_906, i_8_912, i_8_935, i_8_938, i_8_945, i_8_966, i_8_1029, i_8_1046, i_8_1050, i_8_1052, i_8_1074, i_8_1104, i_8_1111, i_8_1114, i_8_1128, i_8_1129, i_8_1222, i_8_1317, i_8_1323, i_8_1330, i_8_1346, i_8_1348, i_8_1378, i_8_1380, i_8_1438, i_8_1456, i_8_1459, i_8_1490, i_8_1506, i_8_1539, i_8_1542, i_8_1556, i_8_1560, i_8_1637, i_8_1667, i_8_1669, i_8_1678, i_8_1682, i_8_1704, i_8_1707, i_8_1722, i_8_1726, i_8_1753, i_8_1762, i_8_1785, i_8_1799, i_8_1863, i_8_1918, i_8_1919, i_8_1934, i_8_1977, i_8_1996, i_8_2006, i_8_2028, i_8_2101, i_8_2112, i_8_2119, i_8_2129, i_8_2141, i_8_2190, i_8_2209, i_8_2211, i_8_2217, i_8_2276, i_8_2290, i_8_2293, i_8_2294, o_8_437);
	kernel_8_438 k_8_438(i_8_6, i_8_21, i_8_25, i_8_35, i_8_78, i_8_79, i_8_87, i_8_120, i_8_121, i_8_123, i_8_141, i_8_171, i_8_193, i_8_195, i_8_214, i_8_264, i_8_268, i_8_286, i_8_321, i_8_489, i_8_492, i_8_582, i_8_591, i_8_601, i_8_627, i_8_628, i_8_636, i_8_645, i_8_672, i_8_693, i_8_703, i_8_706, i_8_735, i_8_813, i_8_825, i_8_834, i_8_835, i_8_860, i_8_876, i_8_888, i_8_969, i_8_978, i_8_979, i_8_994, i_8_1032, i_8_1033, i_8_1131, i_8_1167, i_8_1185, i_8_1187, i_8_1191, i_8_1213, i_8_1230, i_8_1257, i_8_1264, i_8_1275, i_8_1276, i_8_1281, i_8_1329, i_8_1330, i_8_1349, i_8_1362, i_8_1365, i_8_1404, i_8_1407, i_8_1452, i_8_1455, i_8_1474, i_8_1489, i_8_1491, i_8_1554, i_8_1573, i_8_1578, i_8_1582, i_8_1590, i_8_1651, i_8_1668, i_8_1689, i_8_1749, i_8_1786, i_8_1822, i_8_1858, i_8_1860, i_8_1861, i_8_1907, i_8_1965, i_8_1995, i_8_2013, i_8_2058, i_8_2096, i_8_2140, i_8_2145, i_8_2151, i_8_2152, i_8_2155, i_8_2172, i_8_2193, i_8_2194, i_8_2202, i_8_2247, o_8_438);
	kernel_8_439 k_8_439(i_8_51, i_8_52, i_8_57, i_8_60, i_8_61, i_8_62, i_8_85, i_8_142, i_8_216, i_8_226, i_8_229, i_8_230, i_8_255, i_8_257, i_8_258, i_8_259, i_8_260, i_8_301, i_8_329, i_8_379, i_8_389, i_8_426, i_8_453, i_8_485, i_8_554, i_8_556, i_8_557, i_8_597, i_8_602, i_8_678, i_8_786, i_8_851, i_8_852, i_8_853, i_8_877, i_8_971, i_8_991, i_8_992, i_8_1013, i_8_1050, i_8_1052, i_8_1112, i_8_1120, i_8_1124, i_8_1129, i_8_1137, i_8_1159, i_8_1238, i_8_1261, i_8_1281, i_8_1286, i_8_1315, i_8_1316, i_8_1342, i_8_1407, i_8_1410, i_8_1411, i_8_1449, i_8_1489, i_8_1490, i_8_1535, i_8_1537, i_8_1545, i_8_1549, i_8_1551, i_8_1552, i_8_1553, i_8_1561, i_8_1564, i_8_1615, i_8_1625, i_8_1632, i_8_1633, i_8_1652, i_8_1653, i_8_1655, i_8_1696, i_8_1782, i_8_1789, i_8_1805, i_8_1813, i_8_1855, i_8_1858, i_8_1884, i_8_1885, i_8_1887, i_8_1888, i_8_1889, i_8_1944, i_8_1996, i_8_2028, i_8_2032, i_8_2048, i_8_2073, i_8_2139, i_8_2143, i_8_2147, i_8_2216, i_8_2236, i_8_2273, o_8_439);
	kernel_8_440 k_8_440(i_8_13, i_8_77, i_8_80, i_8_140, i_8_167, i_8_184, i_8_221, i_8_233, i_8_253, i_8_254, i_8_259, i_8_263, i_8_281, i_8_284, i_8_302, i_8_304, i_8_322, i_8_335, i_8_364, i_8_376, i_8_400, i_8_437, i_8_439, i_8_440, i_8_488, i_8_494, i_8_578, i_8_580, i_8_590, i_8_619, i_8_625, i_8_626, i_8_643, i_8_662, i_8_664, i_8_698, i_8_702, i_8_707, i_8_712, i_8_716, i_8_725, i_8_732, i_8_808, i_8_812, i_8_853, i_8_869, i_8_878, i_8_942, i_8_968, i_8_1027, i_8_1057, i_8_1067, i_8_1075, i_8_1143, i_8_1192, i_8_1211, i_8_1220, i_8_1241, i_8_1277, i_8_1282, i_8_1323, i_8_1370, i_8_1411, i_8_1436, i_8_1453, i_8_1480, i_8_1489, i_8_1552, i_8_1561, i_8_1618, i_8_1625, i_8_1697, i_8_1716, i_8_1723, i_8_1729, i_8_1769, i_8_1779, i_8_1780, i_8_1801, i_8_1808, i_8_1825, i_8_1849, i_8_1855, i_8_1904, i_8_1945, i_8_1970, i_8_1993, i_8_2039, i_8_2083, i_8_2111, i_8_2129, i_8_2191, i_8_2192, i_8_2228, i_8_2245, i_8_2247, i_8_2248, i_8_2261, i_8_2282, i_8_2301, o_8_440);
	kernel_8_441 k_8_441(i_8_19, i_8_22, i_8_23, i_8_107, i_8_125, i_8_144, i_8_176, i_8_221, i_8_223, i_8_224, i_8_266, i_8_281, i_8_296, i_8_329, i_8_349, i_8_418, i_8_428, i_8_437, i_8_439, i_8_440, i_8_490, i_8_491, i_8_492, i_8_493, i_8_499, i_8_527, i_8_530, i_8_611, i_8_632, i_8_671, i_8_698, i_8_700, i_8_702, i_8_703, i_8_704, i_8_705, i_8_706, i_8_707, i_8_710, i_8_728, i_8_736, i_8_809, i_8_827, i_8_836, i_8_841, i_8_842, i_8_844, i_8_845, i_8_964, i_8_971, i_8_1047, i_8_1073, i_8_1103, i_8_1157, i_8_1183, i_8_1184, i_8_1300, i_8_1310, i_8_1358, i_8_1363, i_8_1390, i_8_1405, i_8_1411, i_8_1434, i_8_1442, i_8_1471, i_8_1473, i_8_1546, i_8_1565, i_8_1589, i_8_1592, i_8_1607, i_8_1628, i_8_1633, i_8_1643, i_8_1650, i_8_1681, i_8_1694, i_8_1733, i_8_1751, i_8_1771, i_8_1778, i_8_1817, i_8_1850, i_8_1862, i_8_1867, i_8_1871, i_8_1991, i_8_2026, i_8_2028, i_8_2030, i_8_2032, i_8_2074, i_8_2111, i_8_2120, i_8_2140, i_8_2189, i_8_2191, i_8_2192, i_8_2243, o_8_441);
	kernel_8_442 k_8_442(i_8_7, i_8_29, i_8_49, i_8_58, i_8_89, i_8_96, i_8_97, i_8_113, i_8_169, i_8_174, i_8_184, i_8_232, i_8_239, i_8_254, i_8_259, i_8_268, i_8_292, i_8_297, i_8_329, i_8_335, i_8_371, i_8_374, i_8_418, i_8_432, i_8_443, i_8_468, i_8_479, i_8_481, i_8_500, i_8_508, i_8_510, i_8_524, i_8_525, i_8_528, i_8_529, i_8_556, i_8_572, i_8_595, i_8_600, i_8_636, i_8_659, i_8_665, i_8_690, i_8_705, i_8_735, i_8_770, i_8_789, i_8_849, i_8_857, i_8_875, i_8_1039, i_8_1075, i_8_1093, i_8_1189, i_8_1190, i_8_1200, i_8_1219, i_8_1277, i_8_1293, i_8_1297, i_8_1307, i_8_1348, i_8_1408, i_8_1410, i_8_1437, i_8_1471, i_8_1487, i_8_1531, i_8_1536, i_8_1545, i_8_1586, i_8_1624, i_8_1633, i_8_1634, i_8_1669, i_8_1696, i_8_1704, i_8_1724, i_8_1739, i_8_1742, i_8_1768, i_8_1779, i_8_1794, i_8_1795, i_8_1799, i_8_1874, i_8_1906, i_8_1918, i_8_1957, i_8_1958, i_8_1965, i_8_1969, i_8_1981, i_8_2019, i_8_2032, i_8_2116, i_8_2122, i_8_2149, i_8_2236, i_8_2246, o_8_442);
	kernel_8_443 k_8_443(i_8_11, i_8_48, i_8_103, i_8_112, i_8_125, i_8_134, i_8_280, i_8_301, i_8_335, i_8_349, i_8_367, i_8_377, i_8_385, i_8_390, i_8_399, i_8_428, i_8_430, i_8_454, i_8_458, i_8_569, i_8_576, i_8_588, i_8_589, i_8_604, i_8_628, i_8_653, i_8_655, i_8_658, i_8_736, i_8_819, i_8_893, i_8_934, i_8_985, i_8_988, i_8_995, i_8_1033, i_8_1036, i_8_1043, i_8_1078, i_8_1093, i_8_1108, i_8_1109, i_8_1180, i_8_1229, i_8_1232, i_8_1265, i_8_1284, i_8_1285, i_8_1286, i_8_1315, i_8_1319, i_8_1331, i_8_1356, i_8_1363, i_8_1399, i_8_1432, i_8_1459, i_8_1484, i_8_1486, i_8_1514, i_8_1527, i_8_1528, i_8_1548, i_8_1558, i_8_1624, i_8_1638, i_8_1652, i_8_1654, i_8_1658, i_8_1676, i_8_1687, i_8_1706, i_8_1748, i_8_1749, i_8_1765, i_8_1825, i_8_1834, i_8_1836, i_8_1837, i_8_1855, i_8_1860, i_8_1861, i_8_1888, i_8_1902, i_8_1909, i_8_1980, i_8_1992, i_8_2013, i_8_2087, i_8_2093, i_8_2101, i_8_2106, i_8_2132, i_8_2144, i_8_2146, i_8_2147, i_8_2150, i_8_2224, i_8_2245, i_8_2275, o_8_443);
	kernel_8_444 k_8_444(i_8_31, i_8_70, i_8_89, i_8_96, i_8_191, i_8_194, i_8_204, i_8_205, i_8_292, i_8_293, i_8_311, i_8_328, i_8_343, i_8_358, i_8_376, i_8_383, i_8_422, i_8_456, i_8_477, i_8_552, i_8_587, i_8_596, i_8_601, i_8_609, i_8_610, i_8_613, i_8_619, i_8_672, i_8_760, i_8_772, i_8_780, i_8_818, i_8_874, i_8_875, i_8_877, i_8_898, i_8_899, i_8_916, i_8_946, i_8_951, i_8_976, i_8_985, i_8_987, i_8_989, i_8_1030, i_8_1108, i_8_1110, i_8_1132, i_8_1141, i_8_1194, i_8_1223, i_8_1256, i_8_1257, i_8_1259, i_8_1262, i_8_1277, i_8_1281, i_8_1284, i_8_1430, i_8_1438, i_8_1455, i_8_1471, i_8_1483, i_8_1484, i_8_1527, i_8_1552, i_8_1553, i_8_1558, i_8_1582, i_8_1603, i_8_1606, i_8_1637, i_8_1672, i_8_1680, i_8_1699, i_8_1734, i_8_1735, i_8_1743, i_8_1745, i_8_1775, i_8_1779, i_8_1784, i_8_1788, i_8_1797, i_8_1815, i_8_1821, i_8_1822, i_8_1823, i_8_1839, i_8_1855, i_8_1867, i_8_1964, i_8_1982, i_8_2013, i_8_2014, i_8_2050, i_8_2108, i_8_2130, i_8_2193, i_8_2290, o_8_444);
	kernel_8_445 k_8_445(i_8_7, i_8_18, i_8_59, i_8_112, i_8_136, i_8_142, i_8_154, i_8_162, i_8_163, i_8_220, i_8_222, i_8_225, i_8_300, i_8_330, i_8_378, i_8_382, i_8_493, i_8_516, i_8_522, i_8_530, i_8_576, i_8_580, i_8_589, i_8_590, i_8_600, i_8_628, i_8_631, i_8_639, i_8_640, i_8_648, i_8_649, i_8_658, i_8_675, i_8_693, i_8_694, i_8_703, i_8_708, i_8_729, i_8_747, i_8_748, i_8_820, i_8_829, i_8_877, i_8_886, i_8_956, i_8_973, i_8_990, i_8_993, i_8_999, i_8_1034, i_8_1107, i_8_1108, i_8_1125, i_8_1152, i_8_1156, i_8_1161, i_8_1162, i_8_1261, i_8_1275, i_8_1327, i_8_1335, i_8_1352, i_8_1355, i_8_1407, i_8_1433, i_8_1485, i_8_1486, i_8_1530, i_8_1593, i_8_1596, i_8_1609, i_8_1656, i_8_1659, i_8_1680, i_8_1681, i_8_1753, i_8_1773, i_8_1784, i_8_1804, i_8_1818, i_8_1819, i_8_1852, i_8_1853, i_8_1971, i_8_1972, i_8_1992, i_8_2007, i_8_2008, i_8_2043, i_8_2088, i_8_2089, i_8_2093, i_8_2098, i_8_2123, i_8_2145, i_8_2170, i_8_2206, i_8_2226, i_8_2253, i_8_2254, o_8_445);
	kernel_8_446 k_8_446(i_8_10, i_8_114, i_8_115, i_8_120, i_8_121, i_8_125, i_8_171, i_8_193, i_8_196, i_8_223, i_8_232, i_8_292, i_8_349, i_8_365, i_8_422, i_8_426, i_8_472, i_8_475, i_8_507, i_8_556, i_8_572, i_8_602, i_8_625, i_8_679, i_8_696, i_8_698, i_8_724, i_8_732, i_8_784, i_8_787, i_8_814, i_8_832, i_8_843, i_8_862, i_8_877, i_8_885, i_8_930, i_8_967, i_8_976, i_8_984, i_8_994, i_8_995, i_8_1003, i_8_1030, i_8_1040, i_8_1047, i_8_1057, i_8_1126, i_8_1179, i_8_1281, i_8_1315, i_8_1355, i_8_1372, i_8_1436, i_8_1453, i_8_1456, i_8_1484, i_8_1551, i_8_1553, i_8_1623, i_8_1624, i_8_1642, i_8_1650, i_8_1651, i_8_1652, i_8_1653, i_8_1655, i_8_1663, i_8_1696, i_8_1697, i_8_1699, i_8_1747, i_8_1767, i_8_1771, i_8_1804, i_8_1808, i_8_1821, i_8_1823, i_8_1826, i_8_1839, i_8_1867, i_8_1893, i_8_1967, i_8_1992, i_8_2073, i_8_2096, i_8_2100, i_8_2101, i_8_2109, i_8_2119, i_8_2126, i_8_2128, i_8_2134, i_8_2172, i_8_2173, i_8_2176, i_8_2230, i_8_2244, i_8_2245, i_8_2258, o_8_446);
	kernel_8_447 k_8_447(i_8_138, i_8_232, i_8_233, i_8_360, i_8_361, i_8_365, i_8_366, i_8_368, i_8_372, i_8_378, i_8_382, i_8_422, i_8_426, i_8_427, i_8_428, i_8_474, i_8_477, i_8_478, i_8_479, i_8_480, i_8_482, i_8_492, i_8_493, i_8_592, i_8_612, i_8_670, i_8_671, i_8_673, i_8_674, i_8_684, i_8_687, i_8_689, i_8_691, i_8_695, i_8_696, i_8_697, i_8_703, i_8_704, i_8_757, i_8_758, i_8_763, i_8_837, i_8_838, i_8_839, i_8_878, i_8_955, i_8_1060, i_8_1079, i_8_1129, i_8_1132, i_8_1159, i_8_1185, i_8_1224, i_8_1226, i_8_1231, i_8_1273, i_8_1282, i_8_1303, i_8_1305, i_8_1306, i_8_1307, i_8_1332, i_8_1352, i_8_1456, i_8_1477, i_8_1552, i_8_1587, i_8_1719, i_8_1720, i_8_1722, i_8_1737, i_8_1740, i_8_1746, i_8_1807, i_8_1808, i_8_1818, i_8_1820, i_8_1821, i_8_1824, i_8_1832, i_8_1902, i_8_1951, i_8_1967, i_8_1981, i_8_1985, i_8_2143, i_8_2149, i_8_2150, i_8_2223, i_8_2226, i_8_2229, i_8_2272, i_8_2275, i_8_2276, i_8_2289, i_8_2290, i_8_2299, i_8_2300, i_8_2301, i_8_2303, o_8_447);
	kernel_8_448 k_8_448(i_8_19, i_8_31, i_8_37, i_8_46, i_8_50, i_8_60, i_8_114, i_8_172, i_8_175, i_8_238, i_8_271, i_8_307, i_8_311, i_8_334, i_8_343, i_8_365, i_8_379, i_8_397, i_8_417, i_8_418, i_8_424, i_8_439, i_8_443, i_8_526, i_8_527, i_8_550, i_8_571, i_8_572, i_8_592, i_8_611, i_8_630, i_8_661, i_8_664, i_8_680, i_8_688, i_8_695, i_8_700, i_8_705, i_8_707, i_8_736, i_8_760, i_8_796, i_8_797, i_8_805, i_8_839, i_8_841, i_8_842, i_8_861, i_8_863, i_8_886, i_8_941, i_8_955, i_8_956, i_8_963, i_8_964, i_8_1018, i_8_1059, i_8_1066, i_8_1071, i_8_1090, i_8_1101, i_8_1179, i_8_1183, i_8_1226, i_8_1282, i_8_1291, i_8_1305, i_8_1336, i_8_1407, i_8_1408, i_8_1435, i_8_1542, i_8_1545, i_8_1561, i_8_1562, i_8_1587, i_8_1588, i_8_1610, i_8_1618, i_8_1634, i_8_1679, i_8_1697, i_8_1731, i_8_1733, i_8_1765, i_8_1818, i_8_1859, i_8_1888, i_8_1992, i_8_1996, i_8_2017, i_8_2056, i_8_2075, i_8_2145, i_8_2149, i_8_2152, i_8_2155, i_8_2156, i_8_2197, i_8_2209, o_8_448);
	kernel_8_449 k_8_449(i_8_28, i_8_38, i_8_107, i_8_142, i_8_171, i_8_213, i_8_214, i_8_272, i_8_292, i_8_295, i_8_298, i_8_300, i_8_301, i_8_302, i_8_307, i_8_308, i_8_310, i_8_314, i_8_338, i_8_351, i_8_420, i_8_421, i_8_430, i_8_483, i_8_489, i_8_492, i_8_496, i_8_498, i_8_528, i_8_589, i_8_591, i_8_592, i_8_605, i_8_606, i_8_631, i_8_633, i_8_635, i_8_677, i_8_679, i_8_689, i_8_706, i_8_709, i_8_766, i_8_780, i_8_830, i_8_849, i_8_925, i_8_954, i_8_985, i_8_1033, i_8_1138, i_8_1156, i_8_1263, i_8_1264, i_8_1267, i_8_1274, i_8_1283, i_8_1286, i_8_1332, i_8_1333, i_8_1335, i_8_1551, i_8_1558, i_8_1561, i_8_1595, i_8_1650, i_8_1651, i_8_1657, i_8_1658, i_8_1659, i_8_1671, i_8_1719, i_8_1740, i_8_1763, i_8_1779, i_8_1789, i_8_1801, i_8_1803, i_8_1805, i_8_1826, i_8_1861, i_8_1863, i_8_1989, i_8_1994, i_8_2004, i_8_2007, i_8_2010, i_8_2013, i_8_2150, i_8_2155, i_8_2164, i_8_2165, i_8_2253, i_8_2255, i_8_2256, i_8_2268, i_8_2272, i_8_2273, i_8_2275, i_8_2286, o_8_449);
	kernel_8_450 k_8_450(i_8_35, i_8_43, i_8_88, i_8_114, i_8_115, i_8_124, i_8_130, i_8_148, i_8_193, i_8_194, i_8_338, i_8_363, i_8_371, i_8_377, i_8_421, i_8_455, i_8_494, i_8_509, i_8_534, i_8_553, i_8_556, i_8_616, i_8_637, i_8_653, i_8_656, i_8_694, i_8_697, i_8_833, i_8_959, i_8_992, i_8_1027, i_8_1037, i_8_1110, i_8_1111, i_8_1127, i_8_1130, i_8_1132, i_8_1202, i_8_1204, i_8_1224, i_8_1226, i_8_1306, i_8_1307, i_8_1310, i_8_1312, i_8_1399, i_8_1400, i_8_1444, i_8_1455, i_8_1462, i_8_1471, i_8_1472, i_8_1486, i_8_1490, i_8_1524, i_8_1547, i_8_1549, i_8_1550, i_8_1552, i_8_1562, i_8_1634, i_8_1641, i_8_1660, i_8_1669, i_8_1748, i_8_1750, i_8_1771, i_8_1795, i_8_1805, i_8_1810, i_8_1823, i_8_1824, i_8_1825, i_8_1881, i_8_1886, i_8_1895, i_8_1939, i_8_1951, i_8_1973, i_8_1976, i_8_2009, i_8_2011, i_8_2012, i_8_2045, i_8_2090, i_8_2098, i_8_2101, i_8_2122, i_8_2137, i_8_2143, i_8_2146, i_8_2150, i_8_2167, i_8_2170, i_8_2171, i_8_2194, i_8_2201, i_8_2236, i_8_2242, i_8_2245, o_8_450);
	kernel_8_451 k_8_451(i_8_18, i_8_27, i_8_40, i_8_46, i_8_90, i_8_166, i_8_171, i_8_173, i_8_191, i_8_207, i_8_227, i_8_288, i_8_343, i_8_361, i_8_378, i_8_396, i_8_397, i_8_415, i_8_423, i_8_490, i_8_498, i_8_522, i_8_523, i_8_594, i_8_608, i_8_612, i_8_615, i_8_648, i_8_684, i_8_690, i_8_694, i_8_703, i_8_766, i_8_795, i_8_810, i_8_827, i_8_829, i_8_838, i_8_858, i_8_883, i_8_927, i_8_954, i_8_963, i_8_965, i_8_993, i_8_1017, i_8_1053, i_8_1054, i_8_1107, i_8_1143, i_8_1171, i_8_1224, i_8_1225, i_8_1261, i_8_1269, i_8_1278, i_8_1279, i_8_1287, i_8_1288, i_8_1297, i_8_1377, i_8_1380, i_8_1435, i_8_1467, i_8_1489, i_8_1548, i_8_1603, i_8_1629, i_8_1638, i_8_1641, i_8_1693, i_8_1720, i_8_1722, i_8_1729, i_8_1737, i_8_1740, i_8_1741, i_8_1869, i_8_1884, i_8_1936, i_8_1993, i_8_1994, i_8_1998, i_8_2034, i_8_2052, i_8_2053, i_8_2055, i_8_2089, i_8_2101, i_8_2102, i_8_2106, i_8_2140, i_8_2169, i_8_2172, i_8_2178, i_8_2196, i_8_2223, i_8_2225, i_8_2226, i_8_2296, o_8_451);
	kernel_8_452 k_8_452(i_8_44, i_8_45, i_8_60, i_8_69, i_8_70, i_8_90, i_8_106, i_8_166, i_8_194, i_8_224, i_8_225, i_8_226, i_8_227, i_8_241, i_8_301, i_8_340, i_8_341, i_8_348, i_8_362, i_8_402, i_8_528, i_8_529, i_8_601, i_8_602, i_8_628, i_8_630, i_8_631, i_8_632, i_8_651, i_8_652, i_8_653, i_8_654, i_8_660, i_8_665, i_8_672, i_8_691, i_8_717, i_8_719, i_8_765, i_8_768, i_8_795, i_8_836, i_8_839, i_8_844, i_8_853, i_8_857, i_8_877, i_8_880, i_8_881, i_8_1033, i_8_1042, i_8_1105, i_8_1132, i_8_1155, i_8_1156, i_8_1295, i_8_1314, i_8_1321, i_8_1322, i_8_1329, i_8_1330, i_8_1331, i_8_1338, i_8_1339, i_8_1356, i_8_1383, i_8_1384, i_8_1389, i_8_1407, i_8_1410, i_8_1435, i_8_1625, i_8_1673, i_8_1705, i_8_1708, i_8_1776, i_8_1818, i_8_1819, i_8_1821, i_8_1830, i_8_1834, i_8_1835, i_8_1844, i_8_1862, i_8_1942, i_8_1987, i_8_1995, i_8_1996, i_8_2016, i_8_2022, i_8_2095, i_8_2096, i_8_2109, i_8_2112, i_8_2113, i_8_2151, i_8_2171, i_8_2178, i_8_2227, i_8_2244, o_8_452);
	kernel_8_453 k_8_453(i_8_21, i_8_24, i_8_30, i_8_39, i_8_43, i_8_115, i_8_120, i_8_121, i_8_124, i_8_129, i_8_140, i_8_150, i_8_160, i_8_175, i_8_273, i_8_276, i_8_309, i_8_310, i_8_324, i_8_345, i_8_348, i_8_351, i_8_354, i_8_365, i_8_378, i_8_387, i_8_426, i_8_529, i_8_553, i_8_555, i_8_624, i_8_625, i_8_643, i_8_652, i_8_654, i_8_672, i_8_673, i_8_697, i_8_741, i_8_762, i_8_768, i_8_829, i_8_833, i_8_841, i_8_848, i_8_854, i_8_877, i_8_881, i_8_915, i_8_943, i_8_944, i_8_951, i_8_954, i_8_969, i_8_987, i_8_1012, i_8_1203, i_8_1270, i_8_1271, i_8_1285, i_8_1324, i_8_1410, i_8_1432, i_8_1474, i_8_1479, i_8_1482, i_8_1492, i_8_1545, i_8_1546, i_8_1571, i_8_1580, i_8_1605, i_8_1606, i_8_1623, i_8_1641, i_8_1644, i_8_1660, i_8_1705, i_8_1749, i_8_1765, i_8_1806, i_8_1821, i_8_1848, i_8_1912, i_8_1951, i_8_1962, i_8_1969, i_8_1971, i_8_2011, i_8_2046, i_8_2064, i_8_2086, i_8_2094, i_8_2104, i_8_2215, i_8_2224, i_8_2245, i_8_2257, i_8_2272, i_8_2298, o_8_453);
	kernel_8_454 k_8_454(i_8_37, i_8_38, i_8_59, i_8_64, i_8_65, i_8_172, i_8_173, i_8_182, i_8_225, i_8_227, i_8_319, i_8_325, i_8_353, i_8_379, i_8_380, i_8_401, i_8_493, i_8_584, i_8_617, i_8_620, i_8_657, i_8_665, i_8_703, i_8_704, i_8_707, i_8_765, i_8_777, i_8_840, i_8_842, i_8_873, i_8_875, i_8_877, i_8_882, i_8_884, i_8_932, i_8_956, i_8_965, i_8_991, i_8_993, i_8_995, i_8_1026, i_8_1028, i_8_1031, i_8_1073, i_8_1103, i_8_1171, i_8_1172, i_8_1175, i_8_1199, i_8_1225, i_8_1234, i_8_1238, i_8_1315, i_8_1354, i_8_1381, i_8_1382, i_8_1397, i_8_1434, i_8_1439, i_8_1460, i_8_1468, i_8_1469, i_8_1489, i_8_1505, i_8_1543, i_8_1544, i_8_1552, i_8_1648, i_8_1654, i_8_1675, i_8_1676, i_8_1678, i_8_1679, i_8_1702, i_8_1703, i_8_1706, i_8_1746, i_8_1749, i_8_1777, i_8_1778, i_8_1792, i_8_1804, i_8_1819, i_8_1820, i_8_1823, i_8_1855, i_8_1910, i_8_1913, i_8_1918, i_8_1936, i_8_1943, i_8_2053, i_8_2099, i_8_2143, i_8_2144, i_8_2147, i_8_2168, i_8_2183, i_8_2210, i_8_2287, o_8_454);
	kernel_8_455 k_8_455(i_8_7, i_8_26, i_8_79, i_8_86, i_8_134, i_8_140, i_8_184, i_8_206, i_8_250, i_8_314, i_8_359, i_8_366, i_8_401, i_8_499, i_8_521, i_8_529, i_8_539, i_8_556, i_8_575, i_8_583, i_8_601, i_8_611, i_8_652, i_8_656, i_8_664, i_8_665, i_8_719, i_8_737, i_8_754, i_8_763, i_8_781, i_8_789, i_8_844, i_8_886, i_8_896, i_8_917, i_8_923, i_8_959, i_8_962, i_8_968, i_8_1015, i_8_1075, i_8_1078, i_8_1088, i_8_1195, i_8_1196, i_8_1201, i_8_1205, i_8_1230, i_8_1339, i_8_1384, i_8_1385, i_8_1393, i_8_1394, i_8_1403, i_8_1410, i_8_1466, i_8_1484, i_8_1492, i_8_1502, i_8_1517, i_8_1528, i_8_1573, i_8_1601, i_8_1636, i_8_1646, i_8_1652, i_8_1663, i_8_1664, i_8_1700, i_8_1717, i_8_1718, i_8_1727, i_8_1753, i_8_1781, i_8_1826, i_8_1844, i_8_1852, i_8_1879, i_8_1880, i_8_1885, i_8_1922, i_8_1929, i_8_1939, i_8_1979, i_8_2015, i_8_2060, i_8_2065, i_8_2094, i_8_2146, i_8_2149, i_8_2150, i_8_2174, i_8_2177, i_8_2185, i_8_2214, i_8_2217, i_8_2218, i_8_2231, i_8_2240, o_8_455);
	kernel_8_456 k_8_456(i_8_12, i_8_22, i_8_28, i_8_31, i_8_33, i_8_50, i_8_54, i_8_55, i_8_56, i_8_76, i_8_103, i_8_105, i_8_136, i_8_139, i_8_195, i_8_299, i_8_430, i_8_441, i_8_523, i_8_529, i_8_543, i_8_552, i_8_606, i_8_608, i_8_610, i_8_615, i_8_631, i_8_652, i_8_678, i_8_708, i_8_729, i_8_750, i_8_751, i_8_760, i_8_762, i_8_783, i_8_811, i_8_814, i_8_840, i_8_860, i_8_876, i_8_891, i_8_940, i_8_1050, i_8_1090, i_8_1104, i_8_1108, i_8_1111, i_8_1112, i_8_1139, i_8_1246, i_8_1254, i_8_1255, i_8_1294, i_8_1308, i_8_1309, i_8_1314, i_8_1324, i_8_1331, i_8_1334, i_8_1337, i_8_1362, i_8_1399, i_8_1422, i_8_1435, i_8_1441, i_8_1477, i_8_1480, i_8_1512, i_8_1513, i_8_1615, i_8_1632, i_8_1634, i_8_1635, i_8_1680, i_8_1682, i_8_1705, i_8_1714, i_8_1746, i_8_1756, i_8_1757, i_8_1784, i_8_1857, i_8_1885, i_8_1902, i_8_1904, i_8_1912, i_8_1926, i_8_1948, i_8_1975, i_8_1981, i_8_1993, i_8_2029, i_8_2053, i_8_2098, i_8_2149, i_8_2236, i_8_2273, i_8_2286, i_8_2295, o_8_456);
	kernel_8_457 k_8_457(i_8_19, i_8_46, i_8_67, i_8_70, i_8_88, i_8_136, i_8_232, i_8_252, i_8_255, i_8_343, i_8_350, i_8_378, i_8_379, i_8_429, i_8_430, i_8_450, i_8_454, i_8_484, i_8_496, i_8_507, i_8_556, i_8_585, i_8_586, i_8_610, i_8_634, i_8_655, i_8_699, i_8_702, i_8_703, i_8_708, i_8_709, i_8_718, i_8_733, i_8_814, i_8_841, i_8_879, i_8_880, i_8_889, i_8_978, i_8_979, i_8_996, i_8_1032, i_8_1078, i_8_1140, i_8_1141, i_8_1144, i_8_1149, i_8_1150, i_8_1168, i_8_1171, i_8_1227, i_8_1239, i_8_1240, i_8_1251, i_8_1264, i_8_1273, i_8_1275, i_8_1278, i_8_1356, i_8_1357, i_8_1359, i_8_1410, i_8_1412, i_8_1547, i_8_1602, i_8_1603, i_8_1604, i_8_1632, i_8_1637, i_8_1779, i_8_1803, i_8_1819, i_8_1824, i_8_1869, i_8_1986, i_8_1996, i_8_2058, i_8_2059, i_8_2107, i_8_2146, i_8_2148, i_8_2149, i_8_2150, i_8_2152, i_8_2157, i_8_2175, i_8_2176, i_8_2233, i_8_2238, i_8_2241, i_8_2242, i_8_2243, i_8_2244, i_8_2248, i_8_2260, i_8_2263, i_8_2272, i_8_2273, i_8_2301, i_8_2302, o_8_457);
	kernel_8_458 k_8_458(i_8_87, i_8_88, i_8_93, i_8_157, i_8_187, i_8_192, i_8_206, i_8_221, i_8_255, i_8_259, i_8_263, i_8_275, i_8_295, i_8_304, i_8_322, i_8_363, i_8_367, i_8_392, i_8_414, i_8_415, i_8_445, i_8_456, i_8_464, i_8_466, i_8_483, i_8_525, i_8_528, i_8_556, i_8_602, i_8_606, i_8_625, i_8_627, i_8_652, i_8_663, i_8_673, i_8_718, i_8_769, i_8_795, i_8_798, i_8_799, i_8_840, i_8_854, i_8_855, i_8_876, i_8_879, i_8_881, i_8_895, i_8_990, i_8_993, i_8_1033, i_8_1113, i_8_1114, i_8_1159, i_8_1216, i_8_1218, i_8_1263, i_8_1322, i_8_1325, i_8_1331, i_8_1349, i_8_1438, i_8_1443, i_8_1444, i_8_1447, i_8_1524, i_8_1528, i_8_1543, i_8_1555, i_8_1571, i_8_1587, i_8_1590, i_8_1600, i_8_1617, i_8_1648, i_8_1736, i_8_1744, i_8_1786, i_8_1807, i_8_1843, i_8_1844, i_8_1930, i_8_1951, i_8_1989, i_8_2025, i_8_2028, i_8_2050, i_8_2109, i_8_2110, i_8_2131, i_8_2184, i_8_2185, i_8_2186, i_8_2193, i_8_2214, i_8_2215, i_8_2217, i_8_2224, i_8_2235, i_8_2239, i_8_2293, o_8_458);
	kernel_8_459 k_8_459(i_8_86, i_8_148, i_8_157, i_8_201, i_8_203, i_8_207, i_8_221, i_8_231, i_8_232, i_8_298, i_8_300, i_8_340, i_8_342, i_8_350, i_8_370, i_8_388, i_8_454, i_8_473, i_8_479, i_8_484, i_8_485, i_8_498, i_8_525, i_8_543, i_8_552, i_8_574, i_8_625, i_8_659, i_8_663, i_8_666, i_8_667, i_8_678, i_8_704, i_8_708, i_8_762, i_8_768, i_8_778, i_8_779, i_8_829, i_8_867, i_8_949, i_8_984, i_8_991, i_8_1003, i_8_1013, i_8_1030, i_8_1031, i_8_1090, i_8_1104, i_8_1106, i_8_1108, i_8_1117, i_8_1129, i_8_1204, i_8_1217, i_8_1219, i_8_1220, i_8_1327, i_8_1345, i_8_1346, i_8_1358, i_8_1402, i_8_1417, i_8_1443, i_8_1514, i_8_1544, i_8_1563, i_8_1564, i_8_1578, i_8_1594, i_8_1597, i_8_1611, i_8_1613, i_8_1630, i_8_1669, i_8_1677, i_8_1707, i_8_1710, i_8_1713, i_8_1722, i_8_1735, i_8_1774, i_8_1798, i_8_1802, i_8_1826, i_8_1867, i_8_1872, i_8_1899, i_8_2047, i_8_2048, i_8_2049, i_8_2055, i_8_2070, i_8_2074, i_8_2088, i_8_2106, i_8_2227, i_8_2260, i_8_2286, i_8_2299, o_8_459);
	kernel_8_460 k_8_460(i_8_23, i_8_41, i_8_73, i_8_106, i_8_187, i_8_189, i_8_193, i_8_217, i_8_243, i_8_364, i_8_390, i_8_411, i_8_423, i_8_424, i_8_425, i_8_426, i_8_454, i_8_468, i_8_472, i_8_490, i_8_572, i_8_583, i_8_610, i_8_652, i_8_665, i_8_676, i_8_679, i_8_705, i_8_738, i_8_752, i_8_775, i_8_808, i_8_837, i_8_856, i_8_867, i_8_876, i_8_882, i_8_883, i_8_931, i_8_984, i_8_994, i_8_1039, i_8_1040, i_8_1048, i_8_1057, i_8_1123, i_8_1126, i_8_1138, i_8_1162, i_8_1174, i_8_1200, i_8_1223, i_8_1226, i_8_1239, i_8_1242, i_8_1245, i_8_1286, i_8_1294, i_8_1311, i_8_1348, i_8_1362, i_8_1363, i_8_1396, i_8_1431, i_8_1456, i_8_1539, i_8_1546, i_8_1547, i_8_1563, i_8_1564, i_8_1574, i_8_1601, i_8_1624, i_8_1639, i_8_1642, i_8_1655, i_8_1659, i_8_1679, i_8_1702, i_8_1713, i_8_1746, i_8_1783, i_8_1802, i_8_1861, i_8_1885, i_8_1920, i_8_1974, i_8_1981, i_8_1984, i_8_1992, i_8_2031, i_8_2083, i_8_2091, i_8_2137, i_8_2155, i_8_2164, i_8_2246, i_8_2247, i_8_2272, i_8_2275, o_8_460);
	kernel_8_461 k_8_461(i_8_30, i_8_143, i_8_214, i_8_215, i_8_219, i_8_259, i_8_268, i_8_347, i_8_350, i_8_377, i_8_378, i_8_383, i_8_385, i_8_430, i_8_456, i_8_468, i_8_469, i_8_556, i_8_557, i_8_606, i_8_615, i_8_618, i_8_627, i_8_646, i_8_663, i_8_772, i_8_780, i_8_796, i_8_871, i_8_881, i_8_898, i_8_899, i_8_921, i_8_952, i_8_953, i_8_975, i_8_978, i_8_979, i_8_1015, i_8_1027, i_8_1045, i_8_1051, i_8_1057, i_8_1140, i_8_1159, i_8_1185, i_8_1194, i_8_1204, i_8_1237, i_8_1239, i_8_1272, i_8_1282, i_8_1285, i_8_1286, i_8_1339, i_8_1429, i_8_1435, i_8_1438, i_8_1446, i_8_1447, i_8_1474, i_8_1506, i_8_1507, i_8_1527, i_8_1528, i_8_1529, i_8_1534, i_8_1538, i_8_1545, i_8_1555, i_8_1635, i_8_1645, i_8_1652, i_8_1671, i_8_1672, i_8_1735, i_8_1753, i_8_1779, i_8_1786, i_8_1798, i_8_1807, i_8_1840, i_8_1860, i_8_1867, i_8_1941, i_8_1942, i_8_1969, i_8_1987, i_8_2002, i_8_2004, i_8_2014, i_8_2113, i_8_2139, i_8_2151, i_8_2158, i_8_2219, i_8_2264, i_8_2267, i_8_2274, i_8_2293, o_8_461);
	kernel_8_462 k_8_462(i_8_21, i_8_30, i_8_86, i_8_87, i_8_142, i_8_169, i_8_185, i_8_187, i_8_193, i_8_213, i_8_233, i_8_255, i_8_256, i_8_260, i_8_292, i_8_295, i_8_346, i_8_376, i_8_417, i_8_418, i_8_445, i_8_453, i_8_456, i_8_464, i_8_481, i_8_485, i_8_503, i_8_510, i_8_522, i_8_525, i_8_526, i_8_530, i_8_556, i_8_592, i_8_601, i_8_704, i_8_705, i_8_717, i_8_761, i_8_763, i_8_764, i_8_789, i_8_798, i_8_894, i_8_952, i_8_993, i_8_996, i_8_998, i_8_1050, i_8_1074, i_8_1078, i_8_1121, i_8_1123, i_8_1124, i_8_1159, i_8_1191, i_8_1305, i_8_1306, i_8_1307, i_8_1308, i_8_1310, i_8_1328, i_8_1411, i_8_1419, i_8_1444, i_8_1447, i_8_1471, i_8_1510, i_8_1543, i_8_1544, i_8_1545, i_8_1578, i_8_1633, i_8_1642, i_8_1707, i_8_1723, i_8_1730, i_8_1733, i_8_1741, i_8_1752, i_8_1779, i_8_1790, i_8_1805, i_8_1812, i_8_1813, i_8_1889, i_8_1906, i_8_1960, i_8_1993, i_8_2049, i_8_2104, i_8_2144, i_8_2218, i_8_2222, i_8_2236, i_8_2247, i_8_2263, i_8_2275, i_8_2292, i_8_2294, o_8_462);
	kernel_8_463 k_8_463(i_8_3, i_8_48, i_8_53, i_8_106, i_8_120, i_8_156, i_8_197, i_8_258, i_8_265, i_8_282, i_8_285, i_8_376, i_8_397, i_8_409, i_8_412, i_8_439, i_8_454, i_8_456, i_8_488, i_8_490, i_8_534, i_8_546, i_8_588, i_8_591, i_8_621, i_8_624, i_8_625, i_8_628, i_8_654, i_8_658, i_8_661, i_8_663, i_8_664, i_8_673, i_8_675, i_8_682, i_8_693, i_8_703, i_8_732, i_8_735, i_8_742, i_8_780, i_8_835, i_8_841, i_8_879, i_8_943, i_8_971, i_8_985, i_8_991, i_8_1019, i_8_1025, i_8_1029, i_8_1066, i_8_1110, i_8_1213, i_8_1257, i_8_1281, i_8_1292, i_8_1362, i_8_1371, i_8_1380, i_8_1451, i_8_1488, i_8_1543, i_8_1544, i_8_1547, i_8_1561, i_8_1675, i_8_1689, i_8_1699, i_8_1704, i_8_1705, i_8_1753, i_8_1770, i_8_1776, i_8_1806, i_8_1807, i_8_1815, i_8_1821, i_8_1830, i_8_1848, i_8_1849, i_8_1857, i_8_1858, i_8_1866, i_8_1911, i_8_1951, i_8_1995, i_8_2010, i_8_2037, i_8_2041, i_8_2082, i_8_2112, i_8_2149, i_8_2193, i_8_2233, i_8_2235, i_8_2236, i_8_2242, i_8_2272, o_8_463);
	kernel_8_464 k_8_464(i_8_33, i_8_34, i_8_70, i_8_76, i_8_77, i_8_141, i_8_187, i_8_191, i_8_205, i_8_214, i_8_215, i_8_224, i_8_267, i_8_268, i_8_292, i_8_330, i_8_332, i_8_340, i_8_358, i_8_446, i_8_448, i_8_456, i_8_457, i_8_463, i_8_468, i_8_486, i_8_557, i_8_603, i_8_618, i_8_619, i_8_627, i_8_637, i_8_661, i_8_664, i_8_719, i_8_772, i_8_787, i_8_825, i_8_855, i_8_879, i_8_898, i_8_899, i_8_925, i_8_952, i_8_953, i_8_987, i_8_988, i_8_998, i_8_1014, i_8_1015, i_8_1016, i_8_1113, i_8_1114, i_8_1128, i_8_1131, i_8_1132, i_8_1141, i_8_1186, i_8_1195, i_8_1429, i_8_1430, i_8_1441, i_8_1455, i_8_1510, i_8_1516, i_8_1537, i_8_1556, i_8_1601, i_8_1618, i_8_1648, i_8_1672, i_8_1673, i_8_1699, i_8_1734, i_8_1741, i_8_1745, i_8_1780, i_8_1781, i_8_1817, i_8_1857, i_8_1907, i_8_1933, i_8_1934, i_8_1951, i_8_2005, i_8_2006, i_8_2013, i_8_2014, i_8_2015, i_8_2050, i_8_2051, i_8_2096, i_8_2130, i_8_2131, i_8_2132, i_8_2139, i_8_2152, i_8_2263, i_8_2274, i_8_2293, o_8_464);
	kernel_8_465 k_8_465(i_8_25, i_8_76, i_8_77, i_8_79, i_8_185, i_8_211, i_8_259, i_8_349, i_8_362, i_8_365, i_8_367, i_8_368, i_8_401, i_8_458, i_8_484, i_8_532, i_8_539, i_8_572, i_8_589, i_8_598, i_8_608, i_8_628, i_8_643, i_8_647, i_8_653, i_8_656, i_8_679, i_8_697, i_8_778, i_8_781, i_8_782, i_8_784, i_8_796, i_8_815, i_8_817, i_8_833, i_8_838, i_8_839, i_8_851, i_8_853, i_8_862, i_8_878, i_8_959, i_8_1067, i_8_1070, i_8_1075, i_8_1134, i_8_1222, i_8_1254, i_8_1264, i_8_1282, i_8_1283, i_8_1286, i_8_1304, i_8_1305, i_8_1327, i_8_1337, i_8_1379, i_8_1391, i_8_1423, i_8_1427, i_8_1436, i_8_1444, i_8_1463, i_8_1466, i_8_1484, i_8_1514, i_8_1549, i_8_1613, i_8_1619, i_8_1630, i_8_1633, i_8_1688, i_8_1706, i_8_1721, i_8_1750, i_8_1751, i_8_1799, i_8_1803, i_8_1807, i_8_1877, i_8_1883, i_8_1898, i_8_1927, i_8_1951, i_8_1988, i_8_1993, i_8_1994, i_8_2006, i_8_2024, i_8_2093, i_8_2140, i_8_2144, i_8_2147, i_8_2158, i_8_2159, i_8_2229, i_8_2261, i_8_2263, i_8_2267, o_8_465);
	kernel_8_466 k_8_466(i_8_39, i_8_52, i_8_66, i_8_69, i_8_139, i_8_169, i_8_174, i_8_183, i_8_192, i_8_210, i_8_232, i_8_264, i_8_270, i_8_291, i_8_295, i_8_327, i_8_345, i_8_348, i_8_366, i_8_384, i_8_445, i_8_462, i_8_466, i_8_528, i_8_552, i_8_554, i_8_598, i_8_633, i_8_662, i_8_664, i_8_674, i_8_687, i_8_699, i_8_704, i_8_768, i_8_770, i_8_777, i_8_843, i_8_858, i_8_877, i_8_880, i_8_990, i_8_993, i_8_1056, i_8_1107, i_8_1113, i_8_1119, i_8_1155, i_8_1156, i_8_1158, i_8_1159, i_8_1173, i_8_1185, i_8_1191, i_8_1230, i_8_1231, i_8_1233, i_8_1237, i_8_1272, i_8_1302, i_8_1317, i_8_1324, i_8_1380, i_8_1452, i_8_1470, i_8_1509, i_8_1540, i_8_1542, i_8_1596, i_8_1600, i_8_1633, i_8_1704, i_8_1731, i_8_1740, i_8_1753, i_8_1806, i_8_1816, i_8_1830, i_8_1843, i_8_1879, i_8_1906, i_8_1948, i_8_1966, i_8_1969, i_8_1975, i_8_1989, i_8_1995, i_8_2109, i_8_2112, i_8_2114, i_8_2145, i_8_2152, i_8_2155, i_8_2158, i_8_2181, i_8_2182, i_8_2190, i_8_2211, i_8_2226, i_8_2275, o_8_466);
	kernel_8_467 k_8_467(i_8_32, i_8_34, i_8_87, i_8_107, i_8_160, i_8_213, i_8_220, i_8_224, i_8_256, i_8_302, i_8_327, i_8_328, i_8_383, i_8_418, i_8_421, i_8_440, i_8_442, i_8_463, i_8_472, i_8_485, i_8_502, i_8_510, i_8_526, i_8_547, i_8_599, i_8_616, i_8_625, i_8_627, i_8_637, i_8_658, i_8_716, i_8_723, i_8_726, i_8_759, i_8_760, i_8_769, i_8_773, i_8_781, i_8_782, i_8_795, i_8_814, i_8_850, i_8_880, i_8_881, i_8_895, i_8_896, i_8_898, i_8_1012, i_8_1013, i_8_1029, i_8_1109, i_8_1115, i_8_1156, i_8_1159, i_8_1318, i_8_1345, i_8_1347, i_8_1348, i_8_1452, i_8_1453, i_8_1471, i_8_1472, i_8_1537, i_8_1544, i_8_1552, i_8_1579, i_8_1599, i_8_1603, i_8_1615, i_8_1633, i_8_1670, i_8_1681, i_8_1714, i_8_1715, i_8_1717, i_8_1726, i_8_1727, i_8_1748, i_8_1759, i_8_1762, i_8_1805, i_8_1860, i_8_1883, i_8_1895, i_8_1903, i_8_1931, i_8_1965, i_8_1995, i_8_2002, i_8_2012, i_8_2031, i_8_2049, i_8_2050, i_8_2110, i_8_2111, i_8_2136, i_8_2145, i_8_2146, i_8_2149, i_8_2215, o_8_467);
	kernel_8_468 k_8_468(i_8_13, i_8_35, i_8_41, i_8_87, i_8_142, i_8_187, i_8_189, i_8_190, i_8_214, i_8_224, i_8_228, i_8_300, i_8_347, i_8_368, i_8_377, i_8_381, i_8_383, i_8_429, i_8_431, i_8_444, i_8_454, i_8_457, i_8_488, i_8_505, i_8_510, i_8_511, i_8_557, i_8_605, i_8_629, i_8_661, i_8_682, i_8_688, i_8_696, i_8_699, i_8_700, i_8_707, i_8_710, i_8_719, i_8_743, i_8_764, i_8_815, i_8_845, i_8_868, i_8_869, i_8_877, i_8_951, i_8_971, i_8_977, i_8_980, i_8_1065, i_8_1106, i_8_1112, i_8_1132, i_8_1184, i_8_1193, i_8_1225, i_8_1232, i_8_1240, i_8_1249, i_8_1268, i_8_1344, i_8_1353, i_8_1417, i_8_1433, i_8_1519, i_8_1537, i_8_1544, i_8_1564, i_8_1581, i_8_1637, i_8_1650, i_8_1654, i_8_1673, i_8_1707, i_8_1717, i_8_1732, i_8_1792, i_8_1808, i_8_1815, i_8_1822, i_8_1861, i_8_1888, i_8_1922, i_8_1933, i_8_1947, i_8_2046, i_8_2056, i_8_2092, i_8_2111, i_8_2112, i_8_2131, i_8_2136, i_8_2137, i_8_2147, i_8_2214, i_8_2218, i_8_2219, i_8_2231, i_8_2244, i_8_2247, o_8_468);
	kernel_8_469 k_8_469(i_8_11, i_8_26, i_8_51, i_8_77, i_8_86, i_8_107, i_8_165, i_8_246, i_8_255, i_8_256, i_8_262, i_8_303, i_8_310, i_8_318, i_8_321, i_8_361, i_8_368, i_8_436, i_8_492, i_8_535, i_8_552, i_8_579, i_8_580, i_8_595, i_8_598, i_8_609, i_8_624, i_8_625, i_8_636, i_8_639, i_8_657, i_8_660, i_8_661, i_8_675, i_8_678, i_8_696, i_8_705, i_8_715, i_8_778, i_8_786, i_8_791, i_8_823, i_8_843, i_8_844, i_8_846, i_8_847, i_8_850, i_8_968, i_8_1040, i_8_1061, i_8_1074, i_8_1139, i_8_1146, i_8_1229, i_8_1233, i_8_1246, i_8_1255, i_8_1273, i_8_1284, i_8_1303, i_8_1317, i_8_1336, i_8_1359, i_8_1362, i_8_1387, i_8_1396, i_8_1455, i_8_1458, i_8_1470, i_8_1471, i_8_1489, i_8_1543, i_8_1545, i_8_1547, i_8_1570, i_8_1696, i_8_1697, i_8_1702, i_8_1733, i_8_1767, i_8_1804, i_8_1819, i_8_1839, i_8_1884, i_8_1885, i_8_1902, i_8_1911, i_8_1912, i_8_1997, i_8_2028, i_8_2095, i_8_2096, i_8_2129, i_8_2133, i_8_2140, i_8_2173, i_8_2191, i_8_2194, i_8_2284, i_8_2289, o_8_469);
	kernel_8_470 k_8_470(i_8_19, i_8_21, i_8_28, i_8_30, i_8_34, i_8_37, i_8_229, i_8_340, i_8_364, i_8_365, i_8_366, i_8_468, i_8_469, i_8_478, i_8_480, i_8_487, i_8_490, i_8_528, i_8_540, i_8_567, i_8_568, i_8_611, i_8_612, i_8_622, i_8_652, i_8_656, i_8_685, i_8_709, i_8_755, i_8_766, i_8_789, i_8_844, i_8_875, i_8_928, i_8_983, i_8_992, i_8_997, i_8_999, i_8_1029, i_8_1042, i_8_1099, i_8_1127, i_8_1225, i_8_1226, i_8_1261, i_8_1262, i_8_1271, i_8_1277, i_8_1280, i_8_1283, i_8_1288, i_8_1297, i_8_1324, i_8_1325, i_8_1378, i_8_1379, i_8_1407, i_8_1468, i_8_1486, i_8_1495, i_8_1536, i_8_1538, i_8_1541, i_8_1549, i_8_1675, i_8_1681, i_8_1682, i_8_1696, i_8_1741, i_8_1752, i_8_1765, i_8_1772, i_8_1817, i_8_1820, i_8_1825, i_8_1827, i_8_1867, i_8_1888, i_8_1889, i_8_1900, i_8_1946, i_8_1971, i_8_1975, i_8_2000, i_8_2015, i_8_2052, i_8_2053, i_8_2130, i_8_2132, i_8_2133, i_8_2139, i_8_2145, i_8_2152, i_8_2224, i_8_2230, i_8_2242, i_8_2243, i_8_2246, i_8_2270, i_8_2273, o_8_470);
	kernel_8_471 k_8_471(i_8_64, i_8_141, i_8_165, i_8_238, i_8_265, i_8_297, i_8_334, i_8_352, i_8_361, i_8_379, i_8_399, i_8_400, i_8_418, i_8_453, i_8_481, i_8_493, i_8_524, i_8_525, i_8_526, i_8_541, i_8_550, i_8_552, i_8_553, i_8_570, i_8_571, i_8_580, i_8_589, i_8_606, i_8_659, i_8_661, i_8_662, i_8_687, i_8_688, i_8_708, i_8_760, i_8_804, i_8_837, i_8_840, i_8_874, i_8_990, i_8_1057, i_8_1058, i_8_1111, i_8_1183, i_8_1200, i_8_1238, i_8_1266, i_8_1267, i_8_1271, i_8_1288, i_8_1291, i_8_1308, i_8_1399, i_8_1411, i_8_1416, i_8_1432, i_8_1437, i_8_1441, i_8_1462, i_8_1515, i_8_1544, i_8_1546, i_8_1547, i_8_1555, i_8_1561, i_8_1564, i_8_1602, i_8_1605, i_8_1611, i_8_1612, i_8_1641, i_8_1679, i_8_1692, i_8_1696, i_8_1714, i_8_1730, i_8_1732, i_8_1786, i_8_1790, i_8_1805, i_8_1809, i_8_1820, i_8_1830, i_8_1938, i_8_1948, i_8_1981, i_8_1992, i_8_1995, i_8_2071, i_8_2073, i_8_2092, i_8_2135, i_8_2142, i_8_2145, i_8_2216, i_8_2223, i_8_2234, i_8_2242, i_8_2244, i_8_2286, o_8_471);
	kernel_8_472 k_8_472(i_8_96, i_8_111, i_8_114, i_8_137, i_8_189, i_8_190, i_8_193, i_8_204, i_8_211, i_8_220, i_8_258, i_8_259, i_8_330, i_8_363, i_8_382, i_8_393, i_8_394, i_8_427, i_8_440, i_8_447, i_8_456, i_8_492, i_8_495, i_8_510, i_8_511, i_8_556, i_8_601, i_8_609, i_8_610, i_8_631, i_8_659, i_8_673, i_8_706, i_8_726, i_8_750, i_8_789, i_8_813, i_8_856, i_8_876, i_8_889, i_8_933, i_8_934, i_8_958, i_8_987, i_8_994, i_8_1029, i_8_1052, i_8_1074, i_8_1087, i_8_1113, i_8_1114, i_8_1124, i_8_1221, i_8_1273, i_8_1281, i_8_1282, i_8_1285, i_8_1301, i_8_1305, i_8_1308, i_8_1331, i_8_1390, i_8_1410, i_8_1435, i_8_1439, i_8_1473, i_8_1493, i_8_1536, i_8_1542, i_8_1573, i_8_1599, i_8_1617, i_8_1635, i_8_1651, i_8_1653, i_8_1669, i_8_1678, i_8_1679, i_8_1681, i_8_1698, i_8_1710, i_8_1725, i_8_1740, i_8_1763, i_8_1851, i_8_1857, i_8_1879, i_8_1905, i_8_1906, i_8_1986, i_8_1987, i_8_1996, i_8_2031, i_8_2037, i_8_2058, i_8_2059, i_8_2107, i_8_2155, i_8_2217, i_8_2283, o_8_472);
	kernel_8_473 k_8_473(i_8_86, i_8_88, i_8_143, i_8_160, i_8_169, i_8_170, i_8_212, i_8_221, i_8_266, i_8_269, i_8_296, i_8_311, i_8_329, i_8_440, i_8_454, i_8_455, i_8_464, i_8_481, i_8_485, i_8_493, i_8_494, i_8_502, i_8_553, i_8_554, i_8_593, i_8_606, i_8_625, i_8_626, i_8_637, i_8_661, i_8_714, i_8_716, i_8_727, i_8_769, i_8_781, i_8_782, i_8_787, i_8_833, i_8_836, i_8_844, i_8_854, i_8_872, i_8_881, i_8_896, i_8_949, i_8_977, i_8_995, i_8_1013, i_8_1067, i_8_1087, i_8_1112, i_8_1114, i_8_1159, i_8_1160, i_8_1228, i_8_1229, i_8_1250, i_8_1336, i_8_1346, i_8_1358, i_8_1401, i_8_1421, i_8_1439, i_8_1444, i_8_1451, i_8_1526, i_8_1546, i_8_1563, i_8_1579, i_8_1580, i_8_1598, i_8_1616, i_8_1625, i_8_1637, i_8_1670, i_8_1679, i_8_1700, i_8_1732, i_8_1750, i_8_1762, i_8_1805, i_8_1825, i_8_1840, i_8_1859, i_8_1862, i_8_1868, i_8_1965, i_8_2002, i_8_2003, i_8_2030, i_8_2032, i_8_2051, i_8_2132, i_8_2141, i_8_2148, i_8_2150, i_8_2151, i_8_2170, i_8_2223, i_8_2290, o_8_473);
	kernel_8_474 k_8_474(i_8_30, i_8_72, i_8_82, i_8_84, i_8_104, i_8_147, i_8_190, i_8_219, i_8_368, i_8_382, i_8_427, i_8_440, i_8_441, i_8_550, i_8_568, i_8_586, i_8_606, i_8_641, i_8_664, i_8_688, i_8_692, i_8_700, i_8_729, i_8_730, i_8_732, i_8_749, i_8_752, i_8_778, i_8_794, i_8_802, i_8_803, i_8_817, i_8_823, i_8_829, i_8_840, i_8_842, i_8_864, i_8_896, i_8_965, i_8_994, i_8_1003, i_8_1009, i_8_1128, i_8_1129, i_8_1156, i_8_1190, i_8_1198, i_8_1229, i_8_1233, i_8_1237, i_8_1261, i_8_1283, i_8_1285, i_8_1295, i_8_1296, i_8_1327, i_8_1351, i_8_1359, i_8_1360, i_8_1362, i_8_1397, i_8_1423, i_8_1432, i_8_1456, i_8_1469, i_8_1481, i_8_1503, i_8_1506, i_8_1513, i_8_1526, i_8_1534, i_8_1548, i_8_1550, i_8_1582, i_8_1672, i_8_1679, i_8_1705, i_8_1721, i_8_1745, i_8_1765, i_8_1804, i_8_1819, i_8_1838, i_8_1877, i_8_1894, i_8_1909, i_8_1910, i_8_1936, i_8_1962, i_8_1972, i_8_1973, i_8_1992, i_8_2072, i_8_2147, i_8_2149, i_8_2224, i_8_2225, i_8_2226, i_8_2273, i_8_2287, o_8_474);
	kernel_8_475 k_8_475(i_8_31, i_8_49, i_8_56, i_8_104, i_8_117, i_8_125, i_8_169, i_8_188, i_8_198, i_8_230, i_8_418, i_8_423, i_8_490, i_8_496, i_8_511, i_8_523, i_8_524, i_8_527, i_8_556, i_8_590, i_8_608, i_8_610, i_8_625, i_8_631, i_8_637, i_8_659, i_8_664, i_8_698, i_8_699, i_8_710, i_8_742, i_8_747, i_8_772, i_8_786, i_8_789, i_8_790, i_8_850, i_8_857, i_8_963, i_8_966, i_8_971, i_8_1043, i_8_1059, i_8_1067, i_8_1078, i_8_1139, i_8_1148, i_8_1160, i_8_1197, i_8_1214, i_8_1233, i_8_1250, i_8_1251, i_8_1279, i_8_1306, i_8_1328, i_8_1354, i_8_1358, i_8_1359, i_8_1426, i_8_1432, i_8_1485, i_8_1490, i_8_1525, i_8_1543, i_8_1544, i_8_1547, i_8_1552, i_8_1630, i_8_1636, i_8_1669, i_8_1674, i_8_1680, i_8_1681, i_8_1682, i_8_1753, i_8_1764, i_8_1778, i_8_1790, i_8_1795, i_8_1801, i_8_1818, i_8_1822, i_8_1837, i_8_1849, i_8_1851, i_8_1888, i_8_1960, i_8_2057, i_8_2105, i_8_2125, i_8_2149, i_8_2150, i_8_2161, i_8_2227, i_8_2229, i_8_2242, i_8_2246, i_8_2254, i_8_2278, o_8_475);
	kernel_8_476 k_8_476(i_8_16, i_8_24, i_8_25, i_8_26, i_8_43, i_8_52, i_8_77, i_8_88, i_8_176, i_8_177, i_8_178, i_8_204, i_8_276, i_8_277, i_8_286, i_8_303, i_8_314, i_8_328, i_8_329, i_8_339, i_8_348, i_8_354, i_8_357, i_8_358, i_8_359, i_8_363, i_8_368, i_8_370, i_8_384, i_8_385, i_8_458, i_8_484, i_8_492, i_8_499, i_8_519, i_8_574, i_8_575, i_8_601, i_8_611, i_8_618, i_8_628, i_8_629, i_8_699, i_8_701, i_8_708, i_8_709, i_8_856, i_8_863, i_8_958, i_8_961, i_8_1015, i_8_1033, i_8_1040, i_8_1042, i_8_1096, i_8_1112, i_8_1176, i_8_1177, i_8_1178, i_8_1195, i_8_1231, i_8_1232, i_8_1274, i_8_1293, i_8_1294, i_8_1295, i_8_1309, i_8_1363, i_8_1365, i_8_1366, i_8_1367, i_8_1457, i_8_1474, i_8_1475, i_8_1564, i_8_1565, i_8_1590, i_8_1603, i_8_1709, i_8_1725, i_8_1726, i_8_1727, i_8_1761, i_8_1770, i_8_1771, i_8_1776, i_8_1825, i_8_1861, i_8_1921, i_8_2052, i_8_2067, i_8_2113, i_8_2157, i_8_2158, i_8_2194, i_8_2213, i_8_2219, i_8_2229, i_8_2239, i_8_2245, o_8_476);
	kernel_8_477 k_8_477(i_8_10, i_8_18, i_8_31, i_8_64, i_8_65, i_8_68, i_8_112, i_8_117, i_8_118, i_8_195, i_8_221, i_8_224, i_8_227, i_8_307, i_8_317, i_8_320, i_8_346, i_8_362, i_8_364, i_8_373, i_8_418, i_8_419, i_8_505, i_8_506, i_8_551, i_8_590, i_8_605, i_8_632, i_8_635, i_8_640, i_8_641, i_8_649, i_8_707, i_8_735, i_8_749, i_8_811, i_8_829, i_8_838, i_8_839, i_8_841, i_8_846, i_8_847, i_8_974, i_8_991, i_8_1035, i_8_1048, i_8_1071, i_8_1081, i_8_1109, i_8_1134, i_8_1135, i_8_1161, i_8_1215, i_8_1229, i_8_1296, i_8_1325, i_8_1360, i_8_1382, i_8_1387, i_8_1423, i_8_1424, i_8_1436, i_8_1460, i_8_1462, i_8_1463, i_8_1471, i_8_1507, i_8_1514, i_8_1522, i_8_1539, i_8_1570, i_8_1571, i_8_1634, i_8_1694, i_8_1703, i_8_1775, i_8_1781, i_8_1838, i_8_1886, i_8_1887, i_8_1888, i_8_1955, i_8_1957, i_8_1970, i_8_1973, i_8_1976, i_8_1982, i_8_1991, i_8_2011, i_8_2052, i_8_2089, i_8_2090, i_8_2097, i_8_2098, i_8_2135, i_8_2188, i_8_2224, i_8_2252, i_8_2255, i_8_2269, o_8_477);
	kernel_8_478 k_8_478(i_8_18, i_8_21, i_8_22, i_8_27, i_8_30, i_8_31, i_8_32, i_8_54, i_8_57, i_8_99, i_8_100, i_8_141, i_8_201, i_8_202, i_8_216, i_8_255, i_8_262, i_8_298, i_8_300, i_8_318, i_8_319, i_8_379, i_8_417, i_8_418, i_8_426, i_8_543, i_8_544, i_8_555, i_8_572, i_8_580, i_8_604, i_8_630, i_8_640, i_8_652, i_8_702, i_8_707, i_8_747, i_8_792, i_8_858, i_8_859, i_8_882, i_8_900, i_8_936, i_8_937, i_8_963, i_8_966, i_8_1035, i_8_1065, i_8_1076, i_8_1161, i_8_1240, i_8_1315, i_8_1319, i_8_1332, i_8_1358, i_8_1359, i_8_1360, i_8_1362, i_8_1395, i_8_1398, i_8_1416, i_8_1462, i_8_1463, i_8_1467, i_8_1472, i_8_1521, i_8_1629, i_8_1630, i_8_1674, i_8_1675, i_8_1676, i_8_1677, i_8_1683, i_8_1710, i_8_1711, i_8_1713, i_8_1812, i_8_1836, i_8_1839, i_8_1926, i_8_1927, i_8_1944, i_8_1945, i_8_1947, i_8_1951, i_8_1962, i_8_1983, i_8_2008, i_8_2119, i_8_2133, i_8_2144, i_8_2154, i_8_2157, i_8_2169, i_8_2196, i_8_2224, i_8_2226, i_8_2232, i_8_2233, i_8_2259, o_8_478);
	kernel_8_479 k_8_479(i_8_35, i_8_74, i_8_89, i_8_107, i_8_142, i_8_189, i_8_190, i_8_222, i_8_259, i_8_331, i_8_379, i_8_386, i_8_392, i_8_445, i_8_457, i_8_481, i_8_502, i_8_522, i_8_555, i_8_556, i_8_597, i_8_634, i_8_645, i_8_664, i_8_696, i_8_699, i_8_706, i_8_762, i_8_817, i_8_818, i_8_826, i_8_897, i_8_906, i_8_925, i_8_943, i_8_951, i_8_979, i_8_980, i_8_987, i_8_988, i_8_997, i_8_1012, i_8_1014, i_8_1015, i_8_1029, i_8_1113, i_8_1122, i_8_1131, i_8_1140, i_8_1186, i_8_1303, i_8_1308, i_8_1327, i_8_1330, i_8_1338, i_8_1348, i_8_1350, i_8_1453, i_8_1455, i_8_1489, i_8_1510, i_8_1527, i_8_1599, i_8_1608, i_8_1617, i_8_1618, i_8_1632, i_8_1651, i_8_1673, i_8_1681, i_8_1686, i_8_1704, i_8_1708, i_8_1716, i_8_1717, i_8_1732, i_8_1750, i_8_1812, i_8_1861, i_8_1862, i_8_1869, i_8_1870, i_8_1876, i_8_1904, i_8_1918, i_8_1949, i_8_1950, i_8_1981, i_8_1993, i_8_2001, i_8_2005, i_8_2049, i_8_2090, i_8_2093, i_8_2107, i_8_2139, i_8_2140, i_8_2184, i_8_2193, i_8_2265, o_8_479);
	kernel_8_480 k_8_480(i_8_13, i_8_21, i_8_22, i_8_58, i_8_66, i_8_109, i_8_114, i_8_138, i_8_194, i_8_219, i_8_220, i_8_279, i_8_285, i_8_321, i_8_325, i_8_328, i_8_345, i_8_364, i_8_384, i_8_396, i_8_400, i_8_486, i_8_492, i_8_527, i_8_530, i_8_552, i_8_555, i_8_573, i_8_589, i_8_594, i_8_595, i_8_606, i_8_608, i_8_615, i_8_696, i_8_777, i_8_822, i_8_838, i_8_874, i_8_877, i_8_880, i_8_883, i_8_891, i_8_894, i_8_969, i_8_970, i_8_972, i_8_1029, i_8_1036, i_8_1092, i_8_1111, i_8_1137, i_8_1146, i_8_1152, i_8_1155, i_8_1197, i_8_1255, i_8_1263, i_8_1317, i_8_1324, i_8_1336, i_8_1396, i_8_1400, i_8_1422, i_8_1423, i_8_1425, i_8_1440, i_8_1443, i_8_1461, i_8_1462, i_8_1481, i_8_1518, i_8_1524, i_8_1525, i_8_1548, i_8_1549, i_8_1587, i_8_1605, i_8_1638, i_8_1639, i_8_1695, i_8_1722, i_8_1724, i_8_1746, i_8_1783, i_8_1813, i_8_1839, i_8_1935, i_8_1967, i_8_1974, i_8_1995, i_8_2011, i_8_2053, i_8_2060, i_8_2110, i_8_2111, i_8_2232, i_8_2233, i_8_2247, i_8_2298, o_8_480);
	kernel_8_481 k_8_481(i_8_31, i_8_70, i_8_187, i_8_188, i_8_259, i_8_301, i_8_305, i_8_367, i_8_368, i_8_430, i_8_454, i_8_493, i_8_505, i_8_512, i_8_556, i_8_565, i_8_584, i_8_593, i_8_596, i_8_599, i_8_607, i_8_610, i_8_627, i_8_630, i_8_631, i_8_634, i_8_643, i_8_654, i_8_682, i_8_707, i_8_778, i_8_781, i_8_782, i_8_796, i_8_842, i_8_844, i_8_865, i_8_890, i_8_965, i_8_976, i_8_977, i_8_1042, i_8_1069, i_8_1105, i_8_1167, i_8_1183, i_8_1201, i_8_1222, i_8_1228, i_8_1244, i_8_1246, i_8_1262, i_8_1264, i_8_1297, i_8_1300, i_8_1313, i_8_1318, i_8_1331, i_8_1427, i_8_1465, i_8_1468, i_8_1471, i_8_1474, i_8_1483, i_8_1516, i_8_1525, i_8_1543, i_8_1552, i_8_1675, i_8_1688, i_8_1694, i_8_1705, i_8_1750, i_8_1752, i_8_1771, i_8_1772, i_8_1783, i_8_1792, i_8_1795, i_8_1821, i_8_1837, i_8_1843, i_8_1888, i_8_1912, i_8_1937, i_8_1943, i_8_1959, i_8_1996, i_8_2047, i_8_2063, i_8_2077, i_8_2132, i_8_2139, i_8_2149, i_8_2155, i_8_2165, i_8_2223, i_8_2227, i_8_2233, i_8_2248, o_8_481);
	kernel_8_482 k_8_482(i_8_49, i_8_65, i_8_114, i_8_168, i_8_211, i_8_212, i_8_219, i_8_223, i_8_227, i_8_252, i_8_353, i_8_372, i_8_422, i_8_453, i_8_456, i_8_472, i_8_481, i_8_483, i_8_496, i_8_526, i_8_552, i_8_555, i_8_573, i_8_628, i_8_636, i_8_661, i_8_698, i_8_708, i_8_807, i_8_840, i_8_861, i_8_888, i_8_923, i_8_929, i_8_942, i_8_993, i_8_996, i_8_1102, i_8_1113, i_8_1114, i_8_1123, i_8_1171, i_8_1172, i_8_1185, i_8_1215, i_8_1224, i_8_1225, i_8_1260, i_8_1261, i_8_1263, i_8_1281, i_8_1282, i_8_1284, i_8_1287, i_8_1288, i_8_1293, i_8_1299, i_8_1308, i_8_1318, i_8_1324, i_8_1338, i_8_1386, i_8_1389, i_8_1395, i_8_1534, i_8_1542, i_8_1590, i_8_1591, i_8_1623, i_8_1626, i_8_1645, i_8_1653, i_8_1677, i_8_1680, i_8_1686, i_8_1689, i_8_1690, i_8_1698, i_8_1722, i_8_1735, i_8_1740, i_8_1741, i_8_1820, i_8_1822, i_8_1887, i_8_1914, i_8_1969, i_8_1996, i_8_2016, i_8_2018, i_8_2077, i_8_2121, i_8_2146, i_8_2155, i_8_2175, i_8_2244, i_8_2247, i_8_2259, i_8_2266, i_8_2287, o_8_482);
	kernel_8_483 k_8_483(i_8_19, i_8_77, i_8_116, i_8_143, i_8_151, i_8_189, i_8_247, i_8_302, i_8_310, i_8_319, i_8_322, i_8_323, i_8_346, i_8_361, i_8_427, i_8_481, i_8_489, i_8_492, i_8_498, i_8_508, i_8_523, i_8_536, i_8_553, i_8_556, i_8_572, i_8_575, i_8_580, i_8_584, i_8_607, i_8_636, i_8_637, i_8_643, i_8_644, i_8_650, i_8_682, i_8_703, i_8_705, i_8_751, i_8_841, i_8_928, i_8_941, i_8_973, i_8_1015, i_8_1083, i_8_1115, i_8_1237, i_8_1282, i_8_1315, i_8_1328, i_8_1339, i_8_1382, i_8_1403, i_8_1436, i_8_1445, i_8_1462, i_8_1463, i_8_1477, i_8_1507, i_8_1508, i_8_1510, i_8_1511, i_8_1520, i_8_1535, i_8_1552, i_8_1555, i_8_1628, i_8_1633, i_8_1648, i_8_1690, i_8_1691, i_8_1694, i_8_1700, i_8_1750, i_8_1751, i_8_1753, i_8_1754, i_8_1771, i_8_1772, i_8_1822, i_8_1840, i_8_1841, i_8_1864, i_8_1894, i_8_1912, i_8_1940, i_8_1952, i_8_1974, i_8_1983, i_8_1997, i_8_2075, i_8_2104, i_8_2137, i_8_2138, i_8_2140, i_8_2147, i_8_2153, i_8_2158, i_8_2216, i_8_2230, i_8_2289, o_8_483);
	kernel_8_484 k_8_484(i_8_104, i_8_127, i_8_145, i_8_176, i_8_190, i_8_217, i_8_219, i_8_274, i_8_305, i_8_334, i_8_352, i_8_360, i_8_370, i_8_417, i_8_427, i_8_481, i_8_490, i_8_495, i_8_496, i_8_514, i_8_522, i_8_523, i_8_552, i_8_595, i_8_604, i_8_607, i_8_658, i_8_667, i_8_669, i_8_712, i_8_828, i_8_831, i_8_849, i_8_855, i_8_878, i_8_1027, i_8_1041, i_8_1071, i_8_1126, i_8_1129, i_8_1156, i_8_1174, i_8_1197, i_8_1225, i_8_1260, i_8_1282, i_8_1296, i_8_1297, i_8_1354, i_8_1387, i_8_1396, i_8_1486, i_8_1494, i_8_1506, i_8_1522, i_8_1531, i_8_1571, i_8_1649, i_8_1651, i_8_1665, i_8_1670, i_8_1681, i_8_1683, i_8_1693, i_8_1702, i_8_1729, i_8_1745, i_8_1747, i_8_1773, i_8_1774, i_8_1791, i_8_1794, i_8_1809, i_8_1813, i_8_1822, i_8_1846, i_8_1863, i_8_1870, i_8_1944, i_8_1945, i_8_1946, i_8_1947, i_8_1964, i_8_1965, i_8_1966, i_8_2007, i_8_2044, i_8_2045, i_8_2046, i_8_2061, i_8_2112, i_8_2116, i_8_2120, i_8_2125, i_8_2188, i_8_2230, i_8_2232, i_8_2260, i_8_2261, i_8_2263, o_8_484);
	kernel_8_485 k_8_485(i_8_11, i_8_52, i_8_84, i_8_93, i_8_153, i_8_172, i_8_174, i_8_241, i_8_245, i_8_300, i_8_306, i_8_345, i_8_346, i_8_354, i_8_363, i_8_381, i_8_384, i_8_385, i_8_450, i_8_457, i_8_507, i_8_523, i_8_526, i_8_528, i_8_609, i_8_612, i_8_615, i_8_634, i_8_642, i_8_660, i_8_675, i_8_694, i_8_702, i_8_705, i_8_709, i_8_764, i_8_768, i_8_795, i_8_804, i_8_822, i_8_880, i_8_921, i_8_924, i_8_930, i_8_967, i_8_993, i_8_1056, i_8_1170, i_8_1173, i_8_1174, i_8_1182, i_8_1189, i_8_1230, i_8_1233, i_8_1236, i_8_1239, i_8_1273, i_8_1288, i_8_1314, i_8_1332, i_8_1354, i_8_1371, i_8_1407, i_8_1440, i_8_1470, i_8_1489, i_8_1497, i_8_1560, i_8_1579, i_8_1605, i_8_1651, i_8_1654, i_8_1665, i_8_1686, i_8_1695, i_8_1758, i_8_1759, i_8_1777, i_8_1792, i_8_1807, i_8_1821, i_8_1824, i_8_1831, i_8_1858, i_8_1936, i_8_1938, i_8_2016, i_8_2019, i_8_2118, i_8_2146, i_8_2152, i_8_2158, i_8_2163, i_8_2172, i_8_2181, i_8_2182, i_8_2244, i_8_2245, i_8_2262, i_8_2283, o_8_485);
	kernel_8_486 k_8_486(i_8_33, i_8_37, i_8_76, i_8_162, i_8_170, i_8_179, i_8_190, i_8_191, i_8_211, i_8_301, i_8_303, i_8_304, i_8_310, i_8_341, i_8_358, i_8_359, i_8_361, i_8_376, i_8_377, i_8_394, i_8_400, i_8_449, i_8_464, i_8_496, i_8_499, i_8_525, i_8_553, i_8_599, i_8_638, i_8_657, i_8_692, i_8_706, i_8_752, i_8_827, i_8_836, i_8_850, i_8_863, i_8_868, i_8_872, i_8_923, i_8_924, i_8_928, i_8_959, i_8_962, i_8_968, i_8_1003, i_8_1035, i_8_1079, i_8_1111, i_8_1126, i_8_1139, i_8_1227, i_8_1241, i_8_1258, i_8_1264, i_8_1266, i_8_1273, i_8_1274, i_8_1277, i_8_1312, i_8_1313, i_8_1346, i_8_1385, i_8_1400, i_8_1433, i_8_1437, i_8_1450, i_8_1467, i_8_1499, i_8_1552, i_8_1558, i_8_1598, i_8_1642, i_8_1654, i_8_1663, i_8_1678, i_8_1696, i_8_1702, i_8_1733, i_8_1750, i_8_1831, i_8_1870, i_8_1871, i_8_1877, i_8_1880, i_8_1885, i_8_1922, i_8_1996, i_8_2017, i_8_2048, i_8_2066, i_8_2069, i_8_2146, i_8_2147, i_8_2161, i_8_2186, i_8_2216, i_8_2237, i_8_2238, i_8_2285, o_8_486);
	kernel_8_487 k_8_487(i_8_24, i_8_39, i_8_49, i_8_52, i_8_85, i_8_97, i_8_170, i_8_175, i_8_181, i_8_189, i_8_193, i_8_238, i_8_263, i_8_277, i_8_300, i_8_302, i_8_313, i_8_340, i_8_345, i_8_378, i_8_403, i_8_494, i_8_556, i_8_603, i_8_613, i_8_634, i_8_637, i_8_676, i_8_687, i_8_698, i_8_700, i_8_706, i_8_707, i_8_748, i_8_769, i_8_798, i_8_840, i_8_849, i_8_855, i_8_879, i_8_883, i_8_924, i_8_925, i_8_931, i_8_934, i_8_970, i_8_990, i_8_1095, i_8_1146, i_8_1230, i_8_1236, i_8_1254, i_8_1273, i_8_1289, i_8_1339, i_8_1350, i_8_1355, i_8_1410, i_8_1455, i_8_1459, i_8_1489, i_8_1512, i_8_1536, i_8_1598, i_8_1606, i_8_1634, i_8_1749, i_8_1788, i_8_1824, i_8_1828, i_8_1831, i_8_1860, i_8_1884, i_8_1885, i_8_1908, i_8_1940, i_8_1947, i_8_1951, i_8_1986, i_8_2004, i_8_2019, i_8_2022, i_8_2091, i_8_2112, i_8_2149, i_8_2157, i_8_2172, i_8_2175, i_8_2182, i_8_2196, i_8_2202, i_8_2211, i_8_2227, i_8_2233, i_8_2235, i_8_2275, i_8_2283, i_8_2284, i_8_2292, i_8_2299, o_8_487);
	kernel_8_488 k_8_488(i_8_37, i_8_75, i_8_81, i_8_129, i_8_192, i_8_193, i_8_214, i_8_225, i_8_230, i_8_241, i_8_242, i_8_337, i_8_343, i_8_347, i_8_365, i_8_478, i_8_482, i_8_483, i_8_484, i_8_502, i_8_525, i_8_528, i_8_588, i_8_612, i_8_616, i_8_619, i_8_620, i_8_631, i_8_653, i_8_654, i_8_655, i_8_656, i_8_664, i_8_669, i_8_687, i_8_690, i_8_710, i_8_732, i_8_751, i_8_760, i_8_762, i_8_763, i_8_765, i_8_768, i_8_769, i_8_770, i_8_772, i_8_792, i_8_796, i_8_831, i_8_832, i_8_833, i_8_841, i_8_970, i_8_971, i_8_1031, i_8_1056, i_8_1156, i_8_1158, i_8_1159, i_8_1263, i_8_1264, i_8_1265, i_8_1272, i_8_1273, i_8_1274, i_8_1306, i_8_1329, i_8_1331, i_8_1350, i_8_1353, i_8_1358, i_8_1407, i_8_1767, i_8_1768, i_8_1770, i_8_1781, i_8_1834, i_8_1995, i_8_1996, i_8_2001, i_8_2078, i_8_2110, i_8_2118, i_8_2119, i_8_2136, i_8_2138, i_8_2150, i_8_2170, i_8_2171, i_8_2208, i_8_2215, i_8_2216, i_8_2224, i_8_2243, i_8_2245, i_8_2248, i_8_2249, i_8_2273, i_8_2289, o_8_488);
	kernel_8_489 k_8_489(i_8_52, i_8_82, i_8_86, i_8_97, i_8_104, i_8_138, i_8_139, i_8_140, i_8_165, i_8_232, i_8_258, i_8_262, i_8_299, i_8_301, i_8_302, i_8_346, i_8_354, i_8_365, i_8_486, i_8_509, i_8_528, i_8_579, i_8_584, i_8_590, i_8_604, i_8_659, i_8_675, i_8_677, i_8_698, i_8_704, i_8_707, i_8_716, i_8_729, i_8_782, i_8_799, i_8_827, i_8_851, i_8_930, i_8_967, i_8_971, i_8_1034, i_8_1108, i_8_1112, i_8_1135, i_8_1157, i_8_1220, i_8_1224, i_8_1236, i_8_1256, i_8_1272, i_8_1285, i_8_1298, i_8_1319, i_8_1404, i_8_1441, i_8_1443, i_8_1465, i_8_1537, i_8_1544, i_8_1558, i_8_1615, i_8_1628, i_8_1632, i_8_1644, i_8_1651, i_8_1652, i_8_1653, i_8_1667, i_8_1691, i_8_1705, i_8_1709, i_8_1783, i_8_1784, i_8_1787, i_8_1796, i_8_1804, i_8_1807, i_8_1838, i_8_1841, i_8_1859, i_8_1877, i_8_1884, i_8_1938, i_8_1948, i_8_1968, i_8_1995, i_8_2026, i_8_2059, i_8_2110, i_8_2111, i_8_2114, i_8_2119, i_8_2133, i_8_2155, i_8_2177, i_8_2183, i_8_2192, i_8_2231, i_8_2273, i_8_2286, o_8_489);
	kernel_8_490 k_8_490(i_8_7, i_8_16, i_8_23, i_8_41, i_8_50, i_8_107, i_8_131, i_8_143, i_8_167, i_8_257, i_8_283, i_8_287, i_8_296, i_8_365, i_8_382, i_8_454, i_8_458, i_8_489, i_8_490, i_8_524, i_8_587, i_8_605, i_8_614, i_8_650, i_8_653, i_8_670, i_8_676, i_8_709, i_8_730, i_8_733, i_8_769, i_8_805, i_8_809, i_8_814, i_8_841, i_8_851, i_8_932, i_8_968, i_8_1067, i_8_1072, i_8_1109, i_8_1139, i_8_1229, i_8_1241, i_8_1274, i_8_1283, i_8_1292, i_8_1301, i_8_1322, i_8_1333, i_8_1385, i_8_1468, i_8_1489, i_8_1491, i_8_1553, i_8_1561, i_8_1574, i_8_1588, i_8_1603, i_8_1610, i_8_1625, i_8_1627, i_8_1628, i_8_1630, i_8_1633, i_8_1672, i_8_1679, i_8_1693, i_8_1700, i_8_1703, i_8_1747, i_8_1774, i_8_1781, i_8_1783, i_8_1822, i_8_1841, i_8_1847, i_8_1850, i_8_1885, i_8_1903, i_8_1963, i_8_1979, i_8_1988, i_8_1996, i_8_1997, i_8_2029, i_8_2039, i_8_2114, i_8_2119, i_8_2120, i_8_2134, i_8_2135, i_8_2147, i_8_2156, i_8_2170, i_8_2183, i_8_2187, i_8_2225, i_8_2243, i_8_2249, o_8_490);
	kernel_8_491 k_8_491(i_8_4, i_8_34, i_8_85, i_8_86, i_8_88, i_8_187, i_8_246, i_8_263, i_8_284, i_8_325, i_8_329, i_8_361, i_8_364, i_8_366, i_8_371, i_8_454, i_8_488, i_8_523, i_8_588, i_8_589, i_8_599, i_8_625, i_8_634, i_8_637, i_8_660, i_8_679, i_8_695, i_8_697, i_8_724, i_8_734, i_8_772, i_8_778, i_8_840, i_8_869, i_8_881, i_8_964, i_8_1020, i_8_1030, i_8_1110, i_8_1118, i_8_1190, i_8_1192, i_8_1227, i_8_1228, i_8_1255, i_8_1265, i_8_1282, i_8_1283, i_8_1285, i_8_1299, i_8_1317, i_8_1354, i_8_1355, i_8_1360, i_8_1373, i_8_1435, i_8_1446, i_8_1471, i_8_1472, i_8_1561, i_8_1624, i_8_1625, i_8_1668, i_8_1671, i_8_1696, i_8_1700, i_8_1703, i_8_1723, i_8_1729, i_8_1743, i_8_1751, i_8_1754, i_8_1768, i_8_1772, i_8_1777, i_8_1820, i_8_1822, i_8_1855, i_8_1857, i_8_1858, i_8_1859, i_8_1870, i_8_1884, i_8_1904, i_8_1912, i_8_1992, i_8_1993, i_8_2120, i_8_2145, i_8_2148, i_8_2155, i_8_2191, i_8_2224, i_8_2244, i_8_2248, i_8_2263, i_8_2272, i_8_2281, i_8_2288, i_8_2290, o_8_491);
	kernel_8_492 k_8_492(i_8_9, i_8_39, i_8_67, i_8_72, i_8_114, i_8_138, i_8_220, i_8_225, i_8_226, i_8_260, i_8_268, i_8_414, i_8_418, i_8_421, i_8_426, i_8_469, i_8_504, i_8_507, i_8_525, i_8_526, i_8_532, i_8_552, i_8_568, i_8_571, i_8_576, i_8_596, i_8_599, i_8_657, i_8_658, i_8_693, i_8_703, i_8_705, i_8_748, i_8_751, i_8_816, i_8_829, i_8_837, i_8_840, i_8_849, i_8_874, i_8_975, i_8_976, i_8_982, i_8_1050, i_8_1110, i_8_1161, i_8_1234, i_8_1237, i_8_1285, i_8_1286, i_8_1297, i_8_1300, i_8_1314, i_8_1315, i_8_1323, i_8_1350, i_8_1354, i_8_1362, i_8_1395, i_8_1432, i_8_1461, i_8_1462, i_8_1470, i_8_1476, i_8_1477, i_8_1481, i_8_1484, i_8_1489, i_8_1512, i_8_1524, i_8_1555, i_8_1621, i_8_1630, i_8_1669, i_8_1729, i_8_1734, i_8_1746, i_8_1747, i_8_1748, i_8_1764, i_8_1773, i_8_1777, i_8_1791, i_8_1794, i_8_1800, i_8_1819, i_8_1857, i_8_1893, i_8_1900, i_8_2053, i_8_2056, i_8_2083, i_8_2098, i_8_2125, i_8_2142, i_8_2152, i_8_2155, i_8_2242, i_8_2269, i_8_2270, o_8_492);
	kernel_8_493 k_8_493(i_8_30, i_8_33, i_8_80, i_8_86, i_8_88, i_8_142, i_8_166, i_8_190, i_8_258, i_8_265, i_8_266, i_8_268, i_8_269, i_8_296, i_8_301, i_8_302, i_8_304, i_8_337, i_8_385, i_8_454, i_8_455, i_8_470, i_8_474, i_8_485, i_8_520, i_8_525, i_8_528, i_8_554, i_8_556, i_8_571, i_8_592, i_8_593, i_8_607, i_8_609, i_8_627, i_8_634, i_8_638, i_8_664, i_8_674, i_8_680, i_8_693, i_8_719, i_8_727, i_8_841, i_8_880, i_8_1016, i_8_1030, i_8_1033, i_8_1115, i_8_1124, i_8_1131, i_8_1237, i_8_1241, i_8_1285, i_8_1286, i_8_1306, i_8_1349, i_8_1437, i_8_1453, i_8_1456, i_8_1457, i_8_1474, i_8_1535, i_8_1546, i_8_1556, i_8_1579, i_8_1601, i_8_1672, i_8_1677, i_8_1678, i_8_1706, i_8_1709, i_8_1742, i_8_1745, i_8_1808, i_8_1834, i_8_1844, i_8_1861, i_8_1906, i_8_1921, i_8_1922, i_8_1952, i_8_1969, i_8_1970, i_8_1996, i_8_2014, i_8_2023, i_8_2024, i_8_2111, i_8_2113, i_8_2122, i_8_2131, i_8_2132, i_8_2137, i_8_2156, i_8_2194, i_8_2195, i_8_2239, i_8_2276, i_8_2293, o_8_493);
	kernel_8_494 k_8_494(i_8_20, i_8_25, i_8_47, i_8_56, i_8_101, i_8_104, i_8_140, i_8_230, i_8_233, i_8_256, i_8_281, i_8_301, i_8_317, i_8_380, i_8_382, i_8_419, i_8_486, i_8_530, i_8_536, i_8_587, i_8_596, i_8_614, i_8_640, i_8_650, i_8_652, i_8_695, i_8_696, i_8_704, i_8_830, i_8_838, i_8_848, i_8_857, i_8_866, i_8_875, i_8_877, i_8_881, i_8_884, i_8_941, i_8_969, i_8_974, i_8_1103, i_8_1136, i_8_1139, i_8_1145, i_8_1202, i_8_1260, i_8_1297, i_8_1304, i_8_1317, i_8_1334, i_8_1342, i_8_1343, i_8_1351, i_8_1352, i_8_1355, i_8_1357, i_8_1397, i_8_1432, i_8_1433, i_8_1468, i_8_1487, i_8_1507, i_8_1525, i_8_1547, i_8_1561, i_8_1564, i_8_1604, i_8_1612, i_8_1688, i_8_1707, i_8_1715, i_8_1721, i_8_1746, i_8_1750, i_8_1753, i_8_1754, i_8_1756, i_8_1766, i_8_1768, i_8_1775, i_8_1785, i_8_1786, i_8_1792, i_8_1814, i_8_1823, i_8_1864, i_8_1883, i_8_1945, i_8_1964, i_8_1984, i_8_1991, i_8_1997, i_8_2054, i_8_2135, i_8_2153, i_8_2192, i_8_2225, i_8_2227, i_8_2234, i_8_2247, o_8_494);
	kernel_8_495 k_8_495(i_8_34, i_8_58, i_8_72, i_8_77, i_8_79, i_8_80, i_8_120, i_8_143, i_8_151, i_8_230, i_8_400, i_8_422, i_8_426, i_8_429, i_8_431, i_8_457, i_8_522, i_8_538, i_8_539, i_8_556, i_8_561, i_8_611, i_8_613, i_8_630, i_8_634, i_8_638, i_8_646, i_8_655, i_8_660, i_8_661, i_8_673, i_8_703, i_8_704, i_8_707, i_8_719, i_8_749, i_8_752, i_8_755, i_8_836, i_8_873, i_8_921, i_8_967, i_8_970, i_8_976, i_8_994, i_8_1013, i_8_1015, i_8_1073, i_8_1075, i_8_1102, i_8_1133, i_8_1266, i_8_1300, i_8_1305, i_8_1337, i_8_1357, i_8_1399, i_8_1400, i_8_1436, i_8_1438, i_8_1439, i_8_1456, i_8_1480, i_8_1489, i_8_1490, i_8_1528, i_8_1542, i_8_1543, i_8_1544, i_8_1572, i_8_1651, i_8_1653, i_8_1677, i_8_1691, i_8_1700, i_8_1703, i_8_1707, i_8_1754, i_8_1770, i_8_1771, i_8_1774, i_8_1794, i_8_1795, i_8_1810, i_8_1823, i_8_1843, i_8_1891, i_8_1912, i_8_1951, i_8_1952, i_8_1957, i_8_1993, i_8_1996, i_8_2131, i_8_2148, i_8_2214, i_8_2215, i_8_2234, i_8_2287, i_8_2299, o_8_495);
	kernel_8_496 k_8_496(i_8_34, i_8_52, i_8_58, i_8_88, i_8_93, i_8_96, i_8_97, i_8_140, i_8_141, i_8_186, i_8_232, i_8_233, i_8_255, i_8_304, i_8_374, i_8_424, i_8_428, i_8_440, i_8_455, i_8_475, i_8_482, i_8_483, i_8_485, i_8_499, i_8_526, i_8_527, i_8_556, i_8_602, i_8_627, i_8_661, i_8_662, i_8_674, i_8_680, i_8_688, i_8_706, i_8_733, i_8_759, i_8_762, i_8_763, i_8_781, i_8_782, i_8_799, i_8_800, i_8_805, i_8_850, i_8_966, i_8_1050, i_8_1051, i_8_1071, i_8_1074, i_8_1075, i_8_1119, i_8_1120, i_8_1122, i_8_1136, i_8_1148, i_8_1191, i_8_1273, i_8_1299, i_8_1305, i_8_1324, i_8_1326, i_8_1390, i_8_1437, i_8_1450, i_8_1470, i_8_1506, i_8_1509, i_8_1533, i_8_1537, i_8_1545, i_8_1563, i_8_1570, i_8_1632, i_8_1652, i_8_1681, i_8_1682, i_8_1684, i_8_1751, i_8_1759, i_8_1763, i_8_1807, i_8_1811, i_8_1821, i_8_1876, i_8_1951, i_8_1982, i_8_1993, i_8_2003, i_8_2029, i_8_2055, i_8_2092, i_8_2093, i_8_2108, i_8_2146, i_8_2150, i_8_2210, i_8_2214, i_8_2215, i_8_2216, o_8_496);
	kernel_8_497 k_8_497(i_8_3, i_8_31, i_8_82, i_8_103, i_8_165, i_8_208, i_8_246, i_8_248, i_8_282, i_8_298, i_8_328, i_8_436, i_8_450, i_8_486, i_8_489, i_8_550, i_8_588, i_8_589, i_8_597, i_8_622, i_8_633, i_8_634, i_8_642, i_8_643, i_8_651, i_8_669, i_8_670, i_8_672, i_8_678, i_8_703, i_8_721, i_8_732, i_8_733, i_8_754, i_8_778, i_8_785, i_8_817, i_8_826, i_8_831, i_8_874, i_8_886, i_8_931, i_8_958, i_8_963, i_8_970, i_8_973, i_8_976, i_8_985, i_8_991, i_8_1071, i_8_1072, i_8_1074, i_8_1130, i_8_1183, i_8_1236, i_8_1263, i_8_1270, i_8_1284, i_8_1285, i_8_1299, i_8_1357, i_8_1359, i_8_1362, i_8_1390, i_8_1439, i_8_1443, i_8_1470, i_8_1570, i_8_1575, i_8_1576, i_8_1588, i_8_1596, i_8_1632, i_8_1633, i_8_1677, i_8_1696, i_8_1699, i_8_1746, i_8_1747, i_8_1749, i_8_1768, i_8_1818, i_8_1822, i_8_1846, i_8_1848, i_8_1854, i_8_1855, i_8_1867, i_8_2010, i_8_2040, i_8_2080, i_8_2119, i_8_2134, i_8_2137, i_8_2147, i_8_2167, i_8_2169, i_8_2209, i_8_2214, i_8_2242, o_8_497);
	kernel_8_498 k_8_498(i_8_31, i_8_35, i_8_36, i_8_89, i_8_110, i_8_140, i_8_256, i_8_273, i_8_301, i_8_329, i_8_345, i_8_346, i_8_375, i_8_377, i_8_418, i_8_434, i_8_451, i_8_454, i_8_463, i_8_511, i_8_528, i_8_529, i_8_530, i_8_553, i_8_554, i_8_589, i_8_595, i_8_611, i_8_620, i_8_670, i_8_671, i_8_673, i_8_709, i_8_716, i_8_772, i_8_780, i_8_781, i_8_796, i_8_824, i_8_865, i_8_975, i_8_984, i_8_985, i_8_1014, i_8_1120, i_8_1131, i_8_1132, i_8_1158, i_8_1159, i_8_1218, i_8_1228, i_8_1249, i_8_1258, i_8_1268, i_8_1306, i_8_1307, i_8_1310, i_8_1387, i_8_1390, i_8_1397, i_8_1453, i_8_1470, i_8_1532, i_8_1533, i_8_1534, i_8_1540, i_8_1556, i_8_1597, i_8_1598, i_8_1607, i_8_1629, i_8_1669, i_8_1684, i_8_1762, i_8_1763, i_8_1808, i_8_1821, i_8_1840, i_8_1870, i_8_1874, i_8_1907, i_8_1948, i_8_1975, i_8_2019, i_8_2044, i_8_2065, i_8_2105, i_8_2126, i_8_2128, i_8_2140, i_8_2154, i_8_2172, i_8_2183, i_8_2188, i_8_2190, i_8_2191, i_8_2213, i_8_2215, i_8_2272, i_8_2289, o_8_498);
	kernel_8_499 k_8_499(i_8_52, i_8_75, i_8_86, i_8_116, i_8_131, i_8_190, i_8_191, i_8_193, i_8_258, i_8_274, i_8_307, i_8_318, i_8_320, i_8_360, i_8_362, i_8_365, i_8_453, i_8_499, i_8_522, i_8_523, i_8_525, i_8_526, i_8_527, i_8_528, i_8_588, i_8_590, i_8_631, i_8_639, i_8_657, i_8_659, i_8_660, i_8_675, i_8_676, i_8_677, i_8_678, i_8_712, i_8_716, i_8_719, i_8_760, i_8_761, i_8_837, i_8_838, i_8_840, i_8_881, i_8_968, i_8_970, i_8_974, i_8_990, i_8_994, i_8_997, i_8_1054, i_8_1128, i_8_1188, i_8_1224, i_8_1228, i_8_1229, i_8_1264, i_8_1267, i_8_1281, i_8_1282, i_8_1285, i_8_1319, i_8_1337, i_8_1404, i_8_1405, i_8_1436, i_8_1453, i_8_1532, i_8_1533, i_8_1534, i_8_1535, i_8_1593, i_8_1598, i_8_1633, i_8_1638, i_8_1650, i_8_1656, i_8_1658, i_8_1660, i_8_1661, i_8_1679, i_8_1783, i_8_1784, i_8_1821, i_8_1822, i_8_1872, i_8_1903, i_8_1975, i_8_2010, i_8_2012, i_8_2052, i_8_2090, i_8_2092, i_8_2093, i_8_2133, i_8_2174, i_8_2216, i_8_2244, i_8_2246, i_8_2247, o_8_499);
	kernel_8_500 k_8_500(i_8_17, i_8_24, i_8_52, i_8_112, i_8_190, i_8_202, i_8_205, i_8_229, i_8_356, i_8_374, i_8_382, i_8_472, i_8_473, i_8_482, i_8_483, i_8_484, i_8_485, i_8_490, i_8_499, i_8_530, i_8_535, i_8_544, i_8_553, i_8_593, i_8_598, i_8_599, i_8_607, i_8_652, i_8_707, i_8_755, i_8_786, i_8_795, i_8_830, i_8_848, i_8_904, i_8_944, i_8_959, i_8_1001, i_8_1002, i_8_1012, i_8_1030, i_8_1135, i_8_1183, i_8_1184, i_8_1228, i_8_1294, i_8_1306, i_8_1340, i_8_1343, i_8_1346, i_8_1390, i_8_1433, i_8_1480, i_8_1525, i_8_1526, i_8_1562, i_8_1565, i_8_1600, i_8_1610, i_8_1639, i_8_1666, i_8_1671, i_8_1678, i_8_1687, i_8_1693, i_8_1694, i_8_1697, i_8_1705, i_8_1708, i_8_1724, i_8_1727, i_8_1751, i_8_1777, i_8_1806, i_8_1822, i_8_1826, i_8_1829, i_8_1858, i_8_1897, i_8_1921, i_8_1975, i_8_2003, i_8_2035, i_8_2038, i_8_2056, i_8_2093, i_8_2107, i_8_2125, i_8_2126, i_8_2134, i_8_2147, i_8_2183, i_8_2215, i_8_2236, i_8_2238, i_8_2242, i_8_2261, i_8_2272, i_8_2285, i_8_2294, o_8_500);
	kernel_8_501 k_8_501(i_8_30, i_8_31, i_8_40, i_8_41, i_8_43, i_8_47, i_8_54, i_8_55, i_8_58, i_8_67, i_8_73, i_8_100, i_8_159, i_8_162, i_8_191, i_8_217, i_8_297, i_8_324, i_8_361, i_8_363, i_8_364, i_8_382, i_8_423, i_8_424, i_8_501, i_8_550, i_8_577, i_8_586, i_8_589, i_8_634, i_8_658, i_8_675, i_8_703, i_8_705, i_8_706, i_8_751, i_8_832, i_8_837, i_8_840, i_8_843, i_8_846, i_8_847, i_8_855, i_8_856, i_8_874, i_8_882, i_8_894, i_8_895, i_8_1039, i_8_1112, i_8_1126, i_8_1129, i_8_1135, i_8_1143, i_8_1263, i_8_1264, i_8_1267, i_8_1279, i_8_1371, i_8_1407, i_8_1424, i_8_1438, i_8_1467, i_8_1468, i_8_1524, i_8_1629, i_8_1630, i_8_1651, i_8_1675, i_8_1677, i_8_1678, i_8_1705, i_8_1713, i_8_1756, i_8_1759, i_8_1767, i_8_1777, i_8_1786, i_8_1807, i_8_1862, i_8_1869, i_8_1899, i_8_1900, i_8_1970, i_8_1993, i_8_2052, i_8_2098, i_8_2106, i_8_2142, i_8_2146, i_8_2148, i_8_2149, i_8_2226, i_8_2232, i_8_2233, i_8_2235, i_8_2247, i_8_2248, i_8_2259, i_8_2262, o_8_501);
	kernel_8_502 k_8_502(i_8_15, i_8_17, i_8_44, i_8_60, i_8_67, i_8_71, i_8_142, i_8_188, i_8_204, i_8_229, i_8_322, i_8_323, i_8_367, i_8_368, i_8_385, i_8_403, i_8_404, i_8_489, i_8_511, i_8_538, i_8_556, i_8_557, i_8_584, i_8_610, i_8_617, i_8_661, i_8_664, i_8_682, i_8_703, i_8_710, i_8_763, i_8_827, i_8_899, i_8_997, i_8_1006, i_8_1075, i_8_1105, i_8_1106, i_8_1113, i_8_1169, i_8_1180, i_8_1181, i_8_1186, i_8_1205, i_8_1261, i_8_1289, i_8_1340, i_8_1439, i_8_1444, i_8_1465, i_8_1471, i_8_1474, i_8_1483, i_8_1484, i_8_1501, i_8_1516, i_8_1520, i_8_1528, i_8_1529, i_8_1553, i_8_1561, i_8_1626, i_8_1632, i_8_1636, i_8_1646, i_8_1651, i_8_1663, i_8_1690, i_8_1699, i_8_1733, i_8_1753, i_8_1771, i_8_1787, i_8_1798, i_8_1800, i_8_1816, i_8_1898, i_8_1916, i_8_1942, i_8_1952, i_8_1958, i_8_1960, i_8_1966, i_8_1967, i_8_1969, i_8_1970, i_8_1988, i_8_2020, i_8_2060, i_8_2077, i_8_2104, i_8_2148, i_8_2172, i_8_2186, i_8_2194, i_8_2215, i_8_2218, i_8_2230, i_8_2239, i_8_2266, o_8_502);
	kernel_8_503 k_8_503(i_8_54, i_8_74, i_8_86, i_8_136, i_8_138, i_8_158, i_8_162, i_8_176, i_8_212, i_8_236, i_8_242, i_8_253, i_8_274, i_8_304, i_8_311, i_8_334, i_8_361, i_8_392, i_8_401, i_8_455, i_8_472, i_8_475, i_8_478, i_8_479, i_8_491, i_8_496, i_8_505, i_8_524, i_8_607, i_8_608, i_8_659, i_8_660, i_8_682, i_8_684, i_8_689, i_8_716, i_8_761, i_8_776, i_8_797, i_8_860, i_8_886, i_8_922, i_8_932, i_8_949, i_8_1058, i_8_1099, i_8_1112, i_8_1154, i_8_1175, i_8_1189, i_8_1190, i_8_1224, i_8_1233, i_8_1240, i_8_1256, i_8_1282, i_8_1283, i_8_1288, i_8_1308, i_8_1325, i_8_1326, i_8_1337, i_8_1409, i_8_1418, i_8_1439, i_8_1456, i_8_1468, i_8_1472, i_8_1480, i_8_1487, i_8_1605, i_8_1607, i_8_1631, i_8_1639, i_8_1650, i_8_1677, i_8_1696, i_8_1700, i_8_1713, i_8_1721, i_8_1760, i_8_1785, i_8_1820, i_8_1835, i_8_1936, i_8_1981, i_8_2003, i_8_2035, i_8_2039, i_8_2053, i_8_2075, i_8_2156, i_8_2159, i_8_2201, i_8_2210, i_8_2223, i_8_2231, i_8_2246, i_8_2261, i_8_2263, o_8_503);
	kernel_8_504 k_8_504(i_8_51, i_8_73, i_8_111, i_8_114, i_8_228, i_8_229, i_8_286, i_8_297, i_8_303, i_8_384, i_8_399, i_8_403, i_8_420, i_8_550, i_8_585, i_8_593, i_8_600, i_8_601, i_8_610, i_8_657, i_8_664, i_8_667, i_8_668, i_8_683, i_8_699, i_8_700, i_8_701, i_8_702, i_8_711, i_8_780, i_8_781, i_8_790, i_8_816, i_8_822, i_8_823, i_8_825, i_8_835, i_8_843, i_8_844, i_8_845, i_8_856, i_8_861, i_8_870, i_8_880, i_8_889, i_8_892, i_8_928, i_8_931, i_8_939, i_8_940, i_8_1027, i_8_1041, i_8_1043, i_8_1107, i_8_1141, i_8_1146, i_8_1149, i_8_1166, i_8_1218, i_8_1242, i_8_1248, i_8_1284, i_8_1285, i_8_1305, i_8_1326, i_8_1335, i_8_1336, i_8_1353, i_8_1354, i_8_1356, i_8_1401, i_8_1425, i_8_1438, i_8_1473, i_8_1482, i_8_1510, i_8_1515, i_8_1546, i_8_1556, i_8_1606, i_8_1630, i_8_1633, i_8_1654, i_8_1714, i_8_1761, i_8_1776, i_8_1801, i_8_1839, i_8_1971, i_8_1981, i_8_1988, i_8_1997, i_8_2058, i_8_2074, i_8_2187, i_8_2214, i_8_2227, i_8_2248, i_8_2277, i_8_2299, o_8_504);
	kernel_8_505 k_8_505(i_8_49, i_8_67, i_8_95, i_8_112, i_8_135, i_8_139, i_8_162, i_8_163, i_8_180, i_8_189, i_8_217, i_8_220, i_8_234, i_8_235, i_8_261, i_8_298, i_8_333, i_8_344, i_8_362, i_8_368, i_8_414, i_8_415, i_8_436, i_8_437, i_8_483, i_8_489, i_8_588, i_8_608, i_8_612, i_8_621, i_8_624, i_8_631, i_8_684, i_8_697, i_8_704, i_8_748, i_8_777, i_8_779, i_8_802, i_8_822, i_8_823, i_8_832, i_8_841, i_8_873, i_8_883, i_8_921, i_8_930, i_8_937, i_8_967, i_8_971, i_8_991, i_8_1011, i_8_1012, i_8_1038, i_8_1053, i_8_1056, i_8_1071, i_8_1104, i_8_1114, i_8_1170, i_8_1235, i_8_1278, i_8_1279, i_8_1284, i_8_1287, i_8_1288, i_8_1395, i_8_1404, i_8_1407, i_8_1434, i_8_1476, i_8_1488, i_8_1535, i_8_1539, i_8_1588, i_8_1740, i_8_1748, i_8_1756, i_8_1800, i_8_1804, i_8_1827, i_8_1828, i_8_1830, i_8_1864, i_8_1986, i_8_1992, i_8_2007, i_8_2019, i_8_2035, i_8_2037, i_8_2043, i_8_2044, i_8_2053, i_8_2070, i_8_2095, i_8_2133, i_8_2187, i_8_2206, i_8_2215, i_8_2268, o_8_505);
	kernel_8_506 k_8_506(i_8_28, i_8_38, i_8_64, i_8_65, i_8_139, i_8_165, i_8_173, i_8_212, i_8_227, i_8_260, i_8_308, i_8_325, i_8_332, i_8_335, i_8_338, i_8_344, i_8_365, i_8_368, i_8_404, i_8_421, i_8_428, i_8_455, i_8_490, i_8_493, i_8_494, i_8_553, i_8_583, i_8_584, i_8_606, i_8_689, i_8_707, i_8_719, i_8_730, i_8_734, i_8_797, i_8_800, i_8_815, i_8_818, i_8_853, i_8_854, i_8_876, i_8_884, i_8_923, i_8_931, i_8_935, i_8_956, i_8_971, i_8_1052, i_8_1060, i_8_1079, i_8_1094, i_8_1107, i_8_1114, i_8_1115, i_8_1172, i_8_1175, i_8_1238, i_8_1264, i_8_1265, i_8_1282, i_8_1290, i_8_1292, i_8_1308, i_8_1322, i_8_1330, i_8_1409, i_8_1411, i_8_1488, i_8_1520, i_8_1535, i_8_1586, i_8_1598, i_8_1655, i_8_1672, i_8_1703, i_8_1706, i_8_1709, i_8_1760, i_8_1821, i_8_1825, i_8_1922, i_8_1937, i_8_1951, i_8_1995, i_8_1996, i_8_2018, i_8_2021, i_8_2075, i_8_2111, i_8_2120, i_8_2170, i_8_2174, i_8_2180, i_8_2201, i_8_2209, i_8_2210, i_8_2227, i_8_2233, i_8_2239, i_8_2276, o_8_506);
	kernel_8_507 k_8_507(i_8_11, i_8_74, i_8_76, i_8_77, i_8_142, i_8_182, i_8_209, i_8_218, i_8_221, i_8_281, i_8_305, i_8_311, i_8_317, i_8_325, i_8_365, i_8_371, i_8_383, i_8_392, i_8_398, i_8_424, i_8_484, i_8_524, i_8_572, i_8_590, i_8_595, i_8_596, i_8_605, i_8_607, i_8_622, i_8_623, i_8_634, i_8_635, i_8_658, i_8_659, i_8_676, i_8_679, i_8_703, i_8_765, i_8_793, i_8_823, i_8_842, i_8_941, i_8_943, i_8_1102, i_8_1181, i_8_1198, i_8_1227, i_8_1235, i_8_1243, i_8_1244, i_8_1265, i_8_1267, i_8_1274, i_8_1282, i_8_1283, i_8_1337, i_8_1370, i_8_1396, i_8_1433, i_8_1451, i_8_1454, i_8_1478, i_8_1504, i_8_1507, i_8_1540, i_8_1544, i_8_1558, i_8_1565, i_8_1568, i_8_1570, i_8_1582, i_8_1631, i_8_1633, i_8_1649, i_8_1702, i_8_1733, i_8_1775, i_8_1777, i_8_1783, i_8_1786, i_8_1804, i_8_1817, i_8_1838, i_8_1841, i_8_1859, i_8_1886, i_8_1945, i_8_1946, i_8_1972, i_8_1973, i_8_2000, i_8_2044, i_8_2141, i_8_2155, i_8_2180, i_8_2206, i_8_2236, i_8_2245, i_8_2270, i_8_2285, o_8_507);
	kernel_8_508 k_8_508(i_8_116, i_8_157, i_8_160, i_8_262, i_8_270, i_8_351, i_8_365, i_8_368, i_8_429, i_8_477, i_8_479, i_8_480, i_8_482, i_8_483, i_8_484, i_8_485, i_8_492, i_8_493, i_8_498, i_8_522, i_8_523, i_8_524, i_8_525, i_8_527, i_8_624, i_8_655, i_8_662, i_8_696, i_8_702, i_8_704, i_8_705, i_8_707, i_8_748, i_8_750, i_8_759, i_8_760, i_8_761, i_8_762, i_8_763, i_8_764, i_8_837, i_8_838, i_8_839, i_8_840, i_8_842, i_8_844, i_8_845, i_8_879, i_8_954, i_8_955, i_8_956, i_8_990, i_8_991, i_8_993, i_8_1226, i_8_1227, i_8_1229, i_8_1232, i_8_1306, i_8_1353, i_8_1354, i_8_1355, i_8_1356, i_8_1434, i_8_1435, i_8_1439, i_8_1587, i_8_1678, i_8_1679, i_8_1682, i_8_1724, i_8_1726, i_8_1727, i_8_1738, i_8_1739, i_8_1754, i_8_1760, i_8_1762, i_8_1763, i_8_1774, i_8_1818, i_8_1819, i_8_1820, i_8_1821, i_8_1822, i_8_1823, i_8_1824, i_8_1825, i_8_1826, i_8_1925, i_8_1969, i_8_1994, i_8_1995, i_8_2051, i_8_2143, i_8_2145, i_8_2147, i_8_2149, i_8_2150, i_8_2215, o_8_508);
	kernel_8_509 k_8_509(i_8_12, i_8_15, i_8_114, i_8_139, i_8_142, i_8_186, i_8_193, i_8_302, i_8_322, i_8_382, i_8_397, i_8_400, i_8_504, i_8_507, i_8_508, i_8_525, i_8_526, i_8_529, i_8_582, i_8_597, i_8_616, i_8_639, i_8_642, i_8_661, i_8_696, i_8_750, i_8_834, i_8_837, i_8_850, i_8_858, i_8_878, i_8_891, i_8_894, i_8_925, i_8_970, i_8_973, i_8_1037, i_8_1038, i_8_1104, i_8_1158, i_8_1260, i_8_1307, i_8_1317, i_8_1321, i_8_1362, i_8_1380, i_8_1399, i_8_1401, i_8_1425, i_8_1440, i_8_1442, i_8_1443, i_8_1461, i_8_1464, i_8_1468, i_8_1488, i_8_1503, i_8_1516, i_8_1533, i_8_1548, i_8_1549, i_8_1561, i_8_1570, i_8_1572, i_8_1573, i_8_1607, i_8_1678, i_8_1681, i_8_1686, i_8_1689, i_8_1693, i_8_1694, i_8_1696, i_8_1698, i_8_1699, i_8_1704, i_8_1722, i_8_1763, i_8_1765, i_8_1785, i_8_1794, i_8_1836, i_8_1839, i_8_1840, i_8_1848, i_8_1884, i_8_1911, i_8_1912, i_8_1935, i_8_1957, i_8_1962, i_8_1965, i_8_1971, i_8_1992, i_8_2055, i_8_2172, i_8_2226, i_8_2247, i_8_2248, i_8_2284, o_8_509);
	kernel_8_510 k_8_510(i_8_22, i_8_23, i_8_40, i_8_77, i_8_107, i_8_184, i_8_259, i_8_346, i_8_359, i_8_368, i_8_454, i_8_499, i_8_541, i_8_552, i_8_607, i_8_634, i_8_644, i_8_656, i_8_664, i_8_671, i_8_680, i_8_682, i_8_683, i_8_707, i_8_725, i_8_727, i_8_728, i_8_755, i_8_778, i_8_818, i_8_824, i_8_835, i_8_841, i_8_844, i_8_860, i_8_869, i_8_876, i_8_877, i_8_938, i_8_980, i_8_1031, i_8_1034, i_8_1125, i_8_1127, i_8_1128, i_8_1131, i_8_1171, i_8_1178, i_8_1185, i_8_1214, i_8_1226, i_8_1267, i_8_1282, i_8_1286, i_8_1345, i_8_1358, i_8_1367, i_8_1394, i_8_1397, i_8_1400, i_8_1411, i_8_1519, i_8_1546, i_8_1551, i_8_1580, i_8_1592, i_8_1633, i_8_1641, i_8_1668, i_8_1671, i_8_1700, i_8_1709, i_8_1730, i_8_1752, i_8_1753, i_8_1769, i_8_1771, i_8_1775, i_8_1777, i_8_1779, i_8_1796, i_8_1801, i_8_1817, i_8_1822, i_8_1823, i_8_1824, i_8_1858, i_8_1859, i_8_2008, i_8_2109, i_8_2126, i_8_2142, i_8_2150, i_8_2152, i_8_2229, i_8_2246, i_8_2248, i_8_2257, i_8_2274, i_8_2293, o_8_510);
	kernel_8_511 k_8_511(i_8_19, i_8_77, i_8_85, i_8_90, i_8_91, i_8_138, i_8_139, i_8_143, i_8_169, i_8_227, i_8_263, i_8_299, i_8_364, i_8_365, i_8_368, i_8_403, i_8_451, i_8_478, i_8_490, i_8_499, i_8_520, i_8_529, i_8_557, i_8_597, i_8_603, i_8_611, i_8_625, i_8_646, i_8_656, i_8_658, i_8_683, i_8_703, i_8_704, i_8_730, i_8_766, i_8_839, i_8_855, i_8_913, i_8_940, i_8_947, i_8_969, i_8_1114, i_8_1117, i_8_1186, i_8_1229, i_8_1261, i_8_1321, i_8_1325, i_8_1426, i_8_1434, i_8_1435, i_8_1468, i_8_1474, i_8_1475, i_8_1507, i_8_1534, i_8_1535, i_8_1544, i_8_1548, i_8_1574, i_8_1674, i_8_1680, i_8_1687, i_8_1700, i_8_1729, i_8_1750, i_8_1753, i_8_1754, i_8_1781, i_8_1784, i_8_1798, i_8_1802, i_8_1808, i_8_1824, i_8_1843, i_8_1844, i_8_1855, i_8_1857, i_8_1888, i_8_1889, i_8_1903, i_8_1968, i_8_1969, i_8_1993, i_8_1996, i_8_1997, i_8_2019, i_8_2087, i_8_2140, i_8_2145, i_8_2146, i_8_2152, i_8_2216, i_8_2226, i_8_2227, i_8_2233, i_8_2235, i_8_2246, i_8_2263, i_8_2287, o_8_511);
endmodule


module kernel_8_wrapper (input ap_clk, ap_rst, ap_ce, ap_start, ap_continue,
                        input [2303:0] in_reg,
                        output ap_idle, ap_done, ap_ready,
                        output out_reg_ap_vld,
                        output reg [511:0] out_reg);

  wire ce = ap_ce;
  reg i_8_0, i_8_1, i_8_2, i_8_3, i_8_4, i_8_5, i_8_6, i_8_7, i_8_8, i_8_9, i_8_10, i_8_11, i_8_12, i_8_13, i_8_14, i_8_15, i_8_16, i_8_17, i_8_18, i_8_19, i_8_20, i_8_21, i_8_22, i_8_23, i_8_24, i_8_25, i_8_26, i_8_27, i_8_28, i_8_29, i_8_30, i_8_31, i_8_32, i_8_33, i_8_34, i_8_35, i_8_36, i_8_37, i_8_38, i_8_39, i_8_40, i_8_41, i_8_42, i_8_43, i_8_44, i_8_45, i_8_46, i_8_47, i_8_48, i_8_49, i_8_50, i_8_51, i_8_52, i_8_53, i_8_54, i_8_55, i_8_56, i_8_57, i_8_58, i_8_59, i_8_60, i_8_61, i_8_62, i_8_63, i_8_64, i_8_65, i_8_66, i_8_67, i_8_68, i_8_69, i_8_70, i_8_71, i_8_72, i_8_73, i_8_74, i_8_75, i_8_76, i_8_77, i_8_78, i_8_79, i_8_80, i_8_81, i_8_82, i_8_83, i_8_84, i_8_85, i_8_86, i_8_87, i_8_88, i_8_89, i_8_90, i_8_91, i_8_92, i_8_93, i_8_94, i_8_95, i_8_96, i_8_97, i_8_98, i_8_99, i_8_100, i_8_101, i_8_102, i_8_103, i_8_104, i_8_105, i_8_106, i_8_107, i_8_108, i_8_109, i_8_110, i_8_111, i_8_112, i_8_113, i_8_114, i_8_115, i_8_116, i_8_117, i_8_118, i_8_119, i_8_120, i_8_121, i_8_122, i_8_123, i_8_124, i_8_125, i_8_126, i_8_127, i_8_128, i_8_129, i_8_130, i_8_131, i_8_132, i_8_133, i_8_134, i_8_135, i_8_136, i_8_137, i_8_138, i_8_139, i_8_140, i_8_141, i_8_142, i_8_143, i_8_144, i_8_145, i_8_146, i_8_147, i_8_148, i_8_149, i_8_150, i_8_151, i_8_152, i_8_153, i_8_154, i_8_155, i_8_156, i_8_157, i_8_158, i_8_159, i_8_160, i_8_161, i_8_162, i_8_163, i_8_164, i_8_165, i_8_166, i_8_167, i_8_168, i_8_169, i_8_170, i_8_171, i_8_172, i_8_173, i_8_174, i_8_175, i_8_176, i_8_177, i_8_178, i_8_179, i_8_180, i_8_181, i_8_182, i_8_183, i_8_184, i_8_185, i_8_186, i_8_187, i_8_188, i_8_189, i_8_190, i_8_191, i_8_192, i_8_193, i_8_194, i_8_195, i_8_196, i_8_197, i_8_198, i_8_199, i_8_200, i_8_201, i_8_202, i_8_203, i_8_204, i_8_205, i_8_206, i_8_207, i_8_208, i_8_209, i_8_210, i_8_211, i_8_212, i_8_213, i_8_214, i_8_215, i_8_216, i_8_217, i_8_218, i_8_219, i_8_220, i_8_221, i_8_222, i_8_223, i_8_224, i_8_225, i_8_226, i_8_227, i_8_228, i_8_229, i_8_230, i_8_231, i_8_232, i_8_233, i_8_234, i_8_235, i_8_236, i_8_237, i_8_238, i_8_239, i_8_240, i_8_241, i_8_242, i_8_243, i_8_244, i_8_245, i_8_246, i_8_247, i_8_248, i_8_249, i_8_250, i_8_251, i_8_252, i_8_253, i_8_254, i_8_255, i_8_256, i_8_257, i_8_258, i_8_259, i_8_260, i_8_261, i_8_262, i_8_263, i_8_264, i_8_265, i_8_266, i_8_267, i_8_268, i_8_269, i_8_270, i_8_271, i_8_272, i_8_273, i_8_274, i_8_275, i_8_276, i_8_277, i_8_278, i_8_279, i_8_280, i_8_281, i_8_282, i_8_283, i_8_284, i_8_285, i_8_286, i_8_287, i_8_288, i_8_289, i_8_290, i_8_291, i_8_292, i_8_293, i_8_294, i_8_295, i_8_296, i_8_297, i_8_298, i_8_299, i_8_300, i_8_301, i_8_302, i_8_303, i_8_304, i_8_305, i_8_306, i_8_307, i_8_308, i_8_309, i_8_310, i_8_311, i_8_312, i_8_313, i_8_314, i_8_315, i_8_316, i_8_317, i_8_318, i_8_319, i_8_320, i_8_321, i_8_322, i_8_323, i_8_324, i_8_325, i_8_326, i_8_327, i_8_328, i_8_329, i_8_330, i_8_331, i_8_332, i_8_333, i_8_334, i_8_335, i_8_336, i_8_337, i_8_338, i_8_339, i_8_340, i_8_341, i_8_342, i_8_343, i_8_344, i_8_345, i_8_346, i_8_347, i_8_348, i_8_349, i_8_350, i_8_351, i_8_352, i_8_353, i_8_354, i_8_355, i_8_356, i_8_357, i_8_358, i_8_359, i_8_360, i_8_361, i_8_362, i_8_363, i_8_364, i_8_365, i_8_366, i_8_367, i_8_368, i_8_369, i_8_370, i_8_371, i_8_372, i_8_373, i_8_374, i_8_375, i_8_376, i_8_377, i_8_378, i_8_379, i_8_380, i_8_381, i_8_382, i_8_383, i_8_384, i_8_385, i_8_386, i_8_387, i_8_388, i_8_389, i_8_390, i_8_391, i_8_392, i_8_393, i_8_394, i_8_395, i_8_396, i_8_397, i_8_398, i_8_399, i_8_400, i_8_401, i_8_402, i_8_403, i_8_404, i_8_405, i_8_406, i_8_407, i_8_408, i_8_409, i_8_410, i_8_411, i_8_412, i_8_413, i_8_414, i_8_415, i_8_416, i_8_417, i_8_418, i_8_419, i_8_420, i_8_421, i_8_422, i_8_423, i_8_424, i_8_425, i_8_426, i_8_427, i_8_428, i_8_429, i_8_430, i_8_431, i_8_432, i_8_433, i_8_434, i_8_435, i_8_436, i_8_437, i_8_438, i_8_439, i_8_440, i_8_441, i_8_442, i_8_443, i_8_444, i_8_445, i_8_446, i_8_447, i_8_448, i_8_449, i_8_450, i_8_451, i_8_452, i_8_453, i_8_454, i_8_455, i_8_456, i_8_457, i_8_458, i_8_459, i_8_460, i_8_461, i_8_462, i_8_463, i_8_464, i_8_465, i_8_466, i_8_467, i_8_468, i_8_469, i_8_470, i_8_471, i_8_472, i_8_473, i_8_474, i_8_475, i_8_476, i_8_477, i_8_478, i_8_479, i_8_480, i_8_481, i_8_482, i_8_483, i_8_484, i_8_485, i_8_486, i_8_487, i_8_488, i_8_489, i_8_490, i_8_491, i_8_492, i_8_493, i_8_494, i_8_495, i_8_496, i_8_497, i_8_498, i_8_499, i_8_500, i_8_501, i_8_502, i_8_503, i_8_504, i_8_505, i_8_506, i_8_507, i_8_508, i_8_509, i_8_510, i_8_511, i_8_512, i_8_513, i_8_514, i_8_515, i_8_516, i_8_517, i_8_518, i_8_519, i_8_520, i_8_521, i_8_522, i_8_523, i_8_524, i_8_525, i_8_526, i_8_527, i_8_528, i_8_529, i_8_530, i_8_531, i_8_532, i_8_533, i_8_534, i_8_535, i_8_536, i_8_537, i_8_538, i_8_539, i_8_540, i_8_541, i_8_542, i_8_543, i_8_544, i_8_545, i_8_546, i_8_547, i_8_548, i_8_549, i_8_550, i_8_551, i_8_552, i_8_553, i_8_554, i_8_555, i_8_556, i_8_557, i_8_558, i_8_559, i_8_560, i_8_561, i_8_562, i_8_563, i_8_564, i_8_565, i_8_566, i_8_567, i_8_568, i_8_569, i_8_570, i_8_571, i_8_572, i_8_573, i_8_574, i_8_575, i_8_576, i_8_577, i_8_578, i_8_579, i_8_580, i_8_581, i_8_582, i_8_583, i_8_584, i_8_585, i_8_586, i_8_587, i_8_588, i_8_589, i_8_590, i_8_591, i_8_592, i_8_593, i_8_594, i_8_595, i_8_596, i_8_597, i_8_598, i_8_599, i_8_600, i_8_601, i_8_602, i_8_603, i_8_604, i_8_605, i_8_606, i_8_607, i_8_608, i_8_609, i_8_610, i_8_611, i_8_612, i_8_613, i_8_614, i_8_615, i_8_616, i_8_617, i_8_618, i_8_619, i_8_620, i_8_621, i_8_622, i_8_623, i_8_624, i_8_625, i_8_626, i_8_627, i_8_628, i_8_629, i_8_630, i_8_631, i_8_632, i_8_633, i_8_634, i_8_635, i_8_636, i_8_637, i_8_638, i_8_639, i_8_640, i_8_641, i_8_642, i_8_643, i_8_644, i_8_645, i_8_646, i_8_647, i_8_648, i_8_649, i_8_650, i_8_651, i_8_652, i_8_653, i_8_654, i_8_655, i_8_656, i_8_657, i_8_658, i_8_659, i_8_660, i_8_661, i_8_662, i_8_663, i_8_664, i_8_665, i_8_666, i_8_667, i_8_668, i_8_669, i_8_670, i_8_671, i_8_672, i_8_673, i_8_674, i_8_675, i_8_676, i_8_677, i_8_678, i_8_679, i_8_680, i_8_681, i_8_682, i_8_683, i_8_684, i_8_685, i_8_686, i_8_687, i_8_688, i_8_689, i_8_690, i_8_691, i_8_692, i_8_693, i_8_694, i_8_695, i_8_696, i_8_697, i_8_698, i_8_699, i_8_700, i_8_701, i_8_702, i_8_703, i_8_704, i_8_705, i_8_706, i_8_707, i_8_708, i_8_709, i_8_710, i_8_711, i_8_712, i_8_713, i_8_714, i_8_715, i_8_716, i_8_717, i_8_718, i_8_719, i_8_720, i_8_721, i_8_722, i_8_723, i_8_724, i_8_725, i_8_726, i_8_727, i_8_728, i_8_729, i_8_730, i_8_731, i_8_732, i_8_733, i_8_734, i_8_735, i_8_736, i_8_737, i_8_738, i_8_739, i_8_740, i_8_741, i_8_742, i_8_743, i_8_744, i_8_745, i_8_746, i_8_747, i_8_748, i_8_749, i_8_750, i_8_751, i_8_752, i_8_753, i_8_754, i_8_755, i_8_756, i_8_757, i_8_758, i_8_759, i_8_760, i_8_761, i_8_762, i_8_763, i_8_764, i_8_765, i_8_766, i_8_767, i_8_768, i_8_769, i_8_770, i_8_771, i_8_772, i_8_773, i_8_774, i_8_775, i_8_776, i_8_777, i_8_778, i_8_779, i_8_780, i_8_781, i_8_782, i_8_783, i_8_784, i_8_785, i_8_786, i_8_787, i_8_788, i_8_789, i_8_790, i_8_791, i_8_792, i_8_793, i_8_794, i_8_795, i_8_796, i_8_797, i_8_798, i_8_799, i_8_800, i_8_801, i_8_802, i_8_803, i_8_804, i_8_805, i_8_806, i_8_807, i_8_808, i_8_809, i_8_810, i_8_811, i_8_812, i_8_813, i_8_814, i_8_815, i_8_816, i_8_817, i_8_818, i_8_819, i_8_820, i_8_821, i_8_822, i_8_823, i_8_824, i_8_825, i_8_826, i_8_827, i_8_828, i_8_829, i_8_830, i_8_831, i_8_832, i_8_833, i_8_834, i_8_835, i_8_836, i_8_837, i_8_838, i_8_839, i_8_840, i_8_841, i_8_842, i_8_843, i_8_844, i_8_845, i_8_846, i_8_847, i_8_848, i_8_849, i_8_850, i_8_851, i_8_852, i_8_853, i_8_854, i_8_855, i_8_856, i_8_857, i_8_858, i_8_859, i_8_860, i_8_861, i_8_862, i_8_863, i_8_864, i_8_865, i_8_866, i_8_867, i_8_868, i_8_869, i_8_870, i_8_871, i_8_872, i_8_873, i_8_874, i_8_875, i_8_876, i_8_877, i_8_878, i_8_879, i_8_880, i_8_881, i_8_882, i_8_883, i_8_884, i_8_885, i_8_886, i_8_887, i_8_888, i_8_889, i_8_890, i_8_891, i_8_892, i_8_893, i_8_894, i_8_895, i_8_896, i_8_897, i_8_898, i_8_899, i_8_900, i_8_901, i_8_902, i_8_903, i_8_904, i_8_905, i_8_906, i_8_907, i_8_908, i_8_909, i_8_910, i_8_911, i_8_912, i_8_913, i_8_914, i_8_915, i_8_916, i_8_917, i_8_918, i_8_919, i_8_920, i_8_921, i_8_922, i_8_923, i_8_924, i_8_925, i_8_926, i_8_927, i_8_928, i_8_929, i_8_930, i_8_931, i_8_932, i_8_933, i_8_934, i_8_935, i_8_936, i_8_937, i_8_938, i_8_939, i_8_940, i_8_941, i_8_942, i_8_943, i_8_944, i_8_945, i_8_946, i_8_947, i_8_948, i_8_949, i_8_950, i_8_951, i_8_952, i_8_953, i_8_954, i_8_955, i_8_956, i_8_957, i_8_958, i_8_959, i_8_960, i_8_961, i_8_962, i_8_963, i_8_964, i_8_965, i_8_966, i_8_967, i_8_968, i_8_969, i_8_970, i_8_971, i_8_972, i_8_973, i_8_974, i_8_975, i_8_976, i_8_977, i_8_978, i_8_979, i_8_980, i_8_981, i_8_982, i_8_983, i_8_984, i_8_985, i_8_986, i_8_987, i_8_988, i_8_989, i_8_990, i_8_991, i_8_992, i_8_993, i_8_994, i_8_995, i_8_996, i_8_997, i_8_998, i_8_999, i_8_1000, i_8_1001, i_8_1002, i_8_1003, i_8_1004, i_8_1005, i_8_1006, i_8_1007, i_8_1008, i_8_1009, i_8_1010, i_8_1011, i_8_1012, i_8_1013, i_8_1014, i_8_1015, i_8_1016, i_8_1017, i_8_1018, i_8_1019, i_8_1020, i_8_1021, i_8_1022, i_8_1023, i_8_1024, i_8_1025, i_8_1026, i_8_1027, i_8_1028, i_8_1029, i_8_1030, i_8_1031, i_8_1032, i_8_1033, i_8_1034, i_8_1035, i_8_1036, i_8_1037, i_8_1038, i_8_1039, i_8_1040, i_8_1041, i_8_1042, i_8_1043, i_8_1044, i_8_1045, i_8_1046, i_8_1047, i_8_1048, i_8_1049, i_8_1050, i_8_1051, i_8_1052, i_8_1053, i_8_1054, i_8_1055, i_8_1056, i_8_1057, i_8_1058, i_8_1059, i_8_1060, i_8_1061, i_8_1062, i_8_1063, i_8_1064, i_8_1065, i_8_1066, i_8_1067, i_8_1068, i_8_1069, i_8_1070, i_8_1071, i_8_1072, i_8_1073, i_8_1074, i_8_1075, i_8_1076, i_8_1077, i_8_1078, i_8_1079, i_8_1080, i_8_1081, i_8_1082, i_8_1083, i_8_1084, i_8_1085, i_8_1086, i_8_1087, i_8_1088, i_8_1089, i_8_1090, i_8_1091, i_8_1092, i_8_1093, i_8_1094, i_8_1095, i_8_1096, i_8_1097, i_8_1098, i_8_1099, i_8_1100, i_8_1101, i_8_1102, i_8_1103, i_8_1104, i_8_1105, i_8_1106, i_8_1107, i_8_1108, i_8_1109, i_8_1110, i_8_1111, i_8_1112, i_8_1113, i_8_1114, i_8_1115, i_8_1116, i_8_1117, i_8_1118, i_8_1119, i_8_1120, i_8_1121, i_8_1122, i_8_1123, i_8_1124, i_8_1125, i_8_1126, i_8_1127, i_8_1128, i_8_1129, i_8_1130, i_8_1131, i_8_1132, i_8_1133, i_8_1134, i_8_1135, i_8_1136, i_8_1137, i_8_1138, i_8_1139, i_8_1140, i_8_1141, i_8_1142, i_8_1143, i_8_1144, i_8_1145, i_8_1146, i_8_1147, i_8_1148, i_8_1149, i_8_1150, i_8_1151, i_8_1152, i_8_1153, i_8_1154, i_8_1155, i_8_1156, i_8_1157, i_8_1158, i_8_1159, i_8_1160, i_8_1161, i_8_1162, i_8_1163, i_8_1164, i_8_1165, i_8_1166, i_8_1167, i_8_1168, i_8_1169, i_8_1170, i_8_1171, i_8_1172, i_8_1173, i_8_1174, i_8_1175, i_8_1176, i_8_1177, i_8_1178, i_8_1179, i_8_1180, i_8_1181, i_8_1182, i_8_1183, i_8_1184, i_8_1185, i_8_1186, i_8_1187, i_8_1188, i_8_1189, i_8_1190, i_8_1191, i_8_1192, i_8_1193, i_8_1194, i_8_1195, i_8_1196, i_8_1197, i_8_1198, i_8_1199, i_8_1200, i_8_1201, i_8_1202, i_8_1203, i_8_1204, i_8_1205, i_8_1206, i_8_1207, i_8_1208, i_8_1209, i_8_1210, i_8_1211, i_8_1212, i_8_1213, i_8_1214, i_8_1215, i_8_1216, i_8_1217, i_8_1218, i_8_1219, i_8_1220, i_8_1221, i_8_1222, i_8_1223, i_8_1224, i_8_1225, i_8_1226, i_8_1227, i_8_1228, i_8_1229, i_8_1230, i_8_1231, i_8_1232, i_8_1233, i_8_1234, i_8_1235, i_8_1236, i_8_1237, i_8_1238, i_8_1239, i_8_1240, i_8_1241, i_8_1242, i_8_1243, i_8_1244, i_8_1245, i_8_1246, i_8_1247, i_8_1248, i_8_1249, i_8_1250, i_8_1251, i_8_1252, i_8_1253, i_8_1254, i_8_1255, i_8_1256, i_8_1257, i_8_1258, i_8_1259, i_8_1260, i_8_1261, i_8_1262, i_8_1263, i_8_1264, i_8_1265, i_8_1266, i_8_1267, i_8_1268, i_8_1269, i_8_1270, i_8_1271, i_8_1272, i_8_1273, i_8_1274, i_8_1275, i_8_1276, i_8_1277, i_8_1278, i_8_1279, i_8_1280, i_8_1281, i_8_1282, i_8_1283, i_8_1284, i_8_1285, i_8_1286, i_8_1287, i_8_1288, i_8_1289, i_8_1290, i_8_1291, i_8_1292, i_8_1293, i_8_1294, i_8_1295, i_8_1296, i_8_1297, i_8_1298, i_8_1299, i_8_1300, i_8_1301, i_8_1302, i_8_1303, i_8_1304, i_8_1305, i_8_1306, i_8_1307, i_8_1308, i_8_1309, i_8_1310, i_8_1311, i_8_1312, i_8_1313, i_8_1314, i_8_1315, i_8_1316, i_8_1317, i_8_1318, i_8_1319, i_8_1320, i_8_1321, i_8_1322, i_8_1323, i_8_1324, i_8_1325, i_8_1326, i_8_1327, i_8_1328, i_8_1329, i_8_1330, i_8_1331, i_8_1332, i_8_1333, i_8_1334, i_8_1335, i_8_1336, i_8_1337, i_8_1338, i_8_1339, i_8_1340, i_8_1341, i_8_1342, i_8_1343, i_8_1344, i_8_1345, i_8_1346, i_8_1347, i_8_1348, i_8_1349, i_8_1350, i_8_1351, i_8_1352, i_8_1353, i_8_1354, i_8_1355, i_8_1356, i_8_1357, i_8_1358, i_8_1359, i_8_1360, i_8_1361, i_8_1362, i_8_1363, i_8_1364, i_8_1365, i_8_1366, i_8_1367, i_8_1368, i_8_1369, i_8_1370, i_8_1371, i_8_1372, i_8_1373, i_8_1374, i_8_1375, i_8_1376, i_8_1377, i_8_1378, i_8_1379, i_8_1380, i_8_1381, i_8_1382, i_8_1383, i_8_1384, i_8_1385, i_8_1386, i_8_1387, i_8_1388, i_8_1389, i_8_1390, i_8_1391, i_8_1392, i_8_1393, i_8_1394, i_8_1395, i_8_1396, i_8_1397, i_8_1398, i_8_1399, i_8_1400, i_8_1401, i_8_1402, i_8_1403, i_8_1404, i_8_1405, i_8_1406, i_8_1407, i_8_1408, i_8_1409, i_8_1410, i_8_1411, i_8_1412, i_8_1413, i_8_1414, i_8_1415, i_8_1416, i_8_1417, i_8_1418, i_8_1419, i_8_1420, i_8_1421, i_8_1422, i_8_1423, i_8_1424, i_8_1425, i_8_1426, i_8_1427, i_8_1428, i_8_1429, i_8_1430, i_8_1431, i_8_1432, i_8_1433, i_8_1434, i_8_1435, i_8_1436, i_8_1437, i_8_1438, i_8_1439, i_8_1440, i_8_1441, i_8_1442, i_8_1443, i_8_1444, i_8_1445, i_8_1446, i_8_1447, i_8_1448, i_8_1449, i_8_1450, i_8_1451, i_8_1452, i_8_1453, i_8_1454, i_8_1455, i_8_1456, i_8_1457, i_8_1458, i_8_1459, i_8_1460, i_8_1461, i_8_1462, i_8_1463, i_8_1464, i_8_1465, i_8_1466, i_8_1467, i_8_1468, i_8_1469, i_8_1470, i_8_1471, i_8_1472, i_8_1473, i_8_1474, i_8_1475, i_8_1476, i_8_1477, i_8_1478, i_8_1479, i_8_1480, i_8_1481, i_8_1482, i_8_1483, i_8_1484, i_8_1485, i_8_1486, i_8_1487, i_8_1488, i_8_1489, i_8_1490, i_8_1491, i_8_1492, i_8_1493, i_8_1494, i_8_1495, i_8_1496, i_8_1497, i_8_1498, i_8_1499, i_8_1500, i_8_1501, i_8_1502, i_8_1503, i_8_1504, i_8_1505, i_8_1506, i_8_1507, i_8_1508, i_8_1509, i_8_1510, i_8_1511, i_8_1512, i_8_1513, i_8_1514, i_8_1515, i_8_1516, i_8_1517, i_8_1518, i_8_1519, i_8_1520, i_8_1521, i_8_1522, i_8_1523, i_8_1524, i_8_1525, i_8_1526, i_8_1527, i_8_1528, i_8_1529, i_8_1530, i_8_1531, i_8_1532, i_8_1533, i_8_1534, i_8_1535, i_8_1536, i_8_1537, i_8_1538, i_8_1539, i_8_1540, i_8_1541, i_8_1542, i_8_1543, i_8_1544, i_8_1545, i_8_1546, i_8_1547, i_8_1548, i_8_1549, i_8_1550, i_8_1551, i_8_1552, i_8_1553, i_8_1554, i_8_1555, i_8_1556, i_8_1557, i_8_1558, i_8_1559, i_8_1560, i_8_1561, i_8_1562, i_8_1563, i_8_1564, i_8_1565, i_8_1566, i_8_1567, i_8_1568, i_8_1569, i_8_1570, i_8_1571, i_8_1572, i_8_1573, i_8_1574, i_8_1575, i_8_1576, i_8_1577, i_8_1578, i_8_1579, i_8_1580, i_8_1581, i_8_1582, i_8_1583, i_8_1584, i_8_1585, i_8_1586, i_8_1587, i_8_1588, i_8_1589, i_8_1590, i_8_1591, i_8_1592, i_8_1593, i_8_1594, i_8_1595, i_8_1596, i_8_1597, i_8_1598, i_8_1599, i_8_1600, i_8_1601, i_8_1602, i_8_1603, i_8_1604, i_8_1605, i_8_1606, i_8_1607, i_8_1608, i_8_1609, i_8_1610, i_8_1611, i_8_1612, i_8_1613, i_8_1614, i_8_1615, i_8_1616, i_8_1617, i_8_1618, i_8_1619, i_8_1620, i_8_1621, i_8_1622, i_8_1623, i_8_1624, i_8_1625, i_8_1626, i_8_1627, i_8_1628, i_8_1629, i_8_1630, i_8_1631, i_8_1632, i_8_1633, i_8_1634, i_8_1635, i_8_1636, i_8_1637, i_8_1638, i_8_1639, i_8_1640, i_8_1641, i_8_1642, i_8_1643, i_8_1644, i_8_1645, i_8_1646, i_8_1647, i_8_1648, i_8_1649, i_8_1650, i_8_1651, i_8_1652, i_8_1653, i_8_1654, i_8_1655, i_8_1656, i_8_1657, i_8_1658, i_8_1659, i_8_1660, i_8_1661, i_8_1662, i_8_1663, i_8_1664, i_8_1665, i_8_1666, i_8_1667, i_8_1668, i_8_1669, i_8_1670, i_8_1671, i_8_1672, i_8_1673, i_8_1674, i_8_1675, i_8_1676, i_8_1677, i_8_1678, i_8_1679, i_8_1680, i_8_1681, i_8_1682, i_8_1683, i_8_1684, i_8_1685, i_8_1686, i_8_1687, i_8_1688, i_8_1689, i_8_1690, i_8_1691, i_8_1692, i_8_1693, i_8_1694, i_8_1695, i_8_1696, i_8_1697, i_8_1698, i_8_1699, i_8_1700, i_8_1701, i_8_1702, i_8_1703, i_8_1704, i_8_1705, i_8_1706, i_8_1707, i_8_1708, i_8_1709, i_8_1710, i_8_1711, i_8_1712, i_8_1713, i_8_1714, i_8_1715, i_8_1716, i_8_1717, i_8_1718, i_8_1719, i_8_1720, i_8_1721, i_8_1722, i_8_1723, i_8_1724, i_8_1725, i_8_1726, i_8_1727, i_8_1728, i_8_1729, i_8_1730, i_8_1731, i_8_1732, i_8_1733, i_8_1734, i_8_1735, i_8_1736, i_8_1737, i_8_1738, i_8_1739, i_8_1740, i_8_1741, i_8_1742, i_8_1743, i_8_1744, i_8_1745, i_8_1746, i_8_1747, i_8_1748, i_8_1749, i_8_1750, i_8_1751, i_8_1752, i_8_1753, i_8_1754, i_8_1755, i_8_1756, i_8_1757, i_8_1758, i_8_1759, i_8_1760, i_8_1761, i_8_1762, i_8_1763, i_8_1764, i_8_1765, i_8_1766, i_8_1767, i_8_1768, i_8_1769, i_8_1770, i_8_1771, i_8_1772, i_8_1773, i_8_1774, i_8_1775, i_8_1776, i_8_1777, i_8_1778, i_8_1779, i_8_1780, i_8_1781, i_8_1782, i_8_1783, i_8_1784, i_8_1785, i_8_1786, i_8_1787, i_8_1788, i_8_1789, i_8_1790, i_8_1791, i_8_1792, i_8_1793, i_8_1794, i_8_1795, i_8_1796, i_8_1797, i_8_1798, i_8_1799, i_8_1800, i_8_1801, i_8_1802, i_8_1803, i_8_1804, i_8_1805, i_8_1806, i_8_1807, i_8_1808, i_8_1809, i_8_1810, i_8_1811, i_8_1812, i_8_1813, i_8_1814, i_8_1815, i_8_1816, i_8_1817, i_8_1818, i_8_1819, i_8_1820, i_8_1821, i_8_1822, i_8_1823, i_8_1824, i_8_1825, i_8_1826, i_8_1827, i_8_1828, i_8_1829, i_8_1830, i_8_1831, i_8_1832, i_8_1833, i_8_1834, i_8_1835, i_8_1836, i_8_1837, i_8_1838, i_8_1839, i_8_1840, i_8_1841, i_8_1842, i_8_1843, i_8_1844, i_8_1845, i_8_1846, i_8_1847, i_8_1848, i_8_1849, i_8_1850, i_8_1851, i_8_1852, i_8_1853, i_8_1854, i_8_1855, i_8_1856, i_8_1857, i_8_1858, i_8_1859, i_8_1860, i_8_1861, i_8_1862, i_8_1863, i_8_1864, i_8_1865, i_8_1866, i_8_1867, i_8_1868, i_8_1869, i_8_1870, i_8_1871, i_8_1872, i_8_1873, i_8_1874, i_8_1875, i_8_1876, i_8_1877, i_8_1878, i_8_1879, i_8_1880, i_8_1881, i_8_1882, i_8_1883, i_8_1884, i_8_1885, i_8_1886, i_8_1887, i_8_1888, i_8_1889, i_8_1890, i_8_1891, i_8_1892, i_8_1893, i_8_1894, i_8_1895, i_8_1896, i_8_1897, i_8_1898, i_8_1899, i_8_1900, i_8_1901, i_8_1902, i_8_1903, i_8_1904, i_8_1905, i_8_1906, i_8_1907, i_8_1908, i_8_1909, i_8_1910, i_8_1911, i_8_1912, i_8_1913, i_8_1914, i_8_1915, i_8_1916, i_8_1917, i_8_1918, i_8_1919, i_8_1920, i_8_1921, i_8_1922, i_8_1923, i_8_1924, i_8_1925, i_8_1926, i_8_1927, i_8_1928, i_8_1929, i_8_1930, i_8_1931, i_8_1932, i_8_1933, i_8_1934, i_8_1935, i_8_1936, i_8_1937, i_8_1938, i_8_1939, i_8_1940, i_8_1941, i_8_1942, i_8_1943, i_8_1944, i_8_1945, i_8_1946, i_8_1947, i_8_1948, i_8_1949, i_8_1950, i_8_1951, i_8_1952, i_8_1953, i_8_1954, i_8_1955, i_8_1956, i_8_1957, i_8_1958, i_8_1959, i_8_1960, i_8_1961, i_8_1962, i_8_1963, i_8_1964, i_8_1965, i_8_1966, i_8_1967, i_8_1968, i_8_1969, i_8_1970, i_8_1971, i_8_1972, i_8_1973, i_8_1974, i_8_1975, i_8_1976, i_8_1977, i_8_1978, i_8_1979, i_8_1980, i_8_1981, i_8_1982, i_8_1983, i_8_1984, i_8_1985, i_8_1986, i_8_1987, i_8_1988, i_8_1989, i_8_1990, i_8_1991, i_8_1992, i_8_1993, i_8_1994, i_8_1995, i_8_1996, i_8_1997, i_8_1998, i_8_1999, i_8_2000, i_8_2001, i_8_2002, i_8_2003, i_8_2004, i_8_2005, i_8_2006, i_8_2007, i_8_2008, i_8_2009, i_8_2010, i_8_2011, i_8_2012, i_8_2013, i_8_2014, i_8_2015, i_8_2016, i_8_2017, i_8_2018, i_8_2019, i_8_2020, i_8_2021, i_8_2022, i_8_2023, i_8_2024, i_8_2025, i_8_2026, i_8_2027, i_8_2028, i_8_2029, i_8_2030, i_8_2031, i_8_2032, i_8_2033, i_8_2034, i_8_2035, i_8_2036, i_8_2037, i_8_2038, i_8_2039, i_8_2040, i_8_2041, i_8_2042, i_8_2043, i_8_2044, i_8_2045, i_8_2046, i_8_2047, i_8_2048, i_8_2049, i_8_2050, i_8_2051, i_8_2052, i_8_2053, i_8_2054, i_8_2055, i_8_2056, i_8_2057, i_8_2058, i_8_2059, i_8_2060, i_8_2061, i_8_2062, i_8_2063, i_8_2064, i_8_2065, i_8_2066, i_8_2067, i_8_2068, i_8_2069, i_8_2070, i_8_2071, i_8_2072, i_8_2073, i_8_2074, i_8_2075, i_8_2076, i_8_2077, i_8_2078, i_8_2079, i_8_2080, i_8_2081, i_8_2082, i_8_2083, i_8_2084, i_8_2085, i_8_2086, i_8_2087, i_8_2088, i_8_2089, i_8_2090, i_8_2091, i_8_2092, i_8_2093, i_8_2094, i_8_2095, i_8_2096, i_8_2097, i_8_2098, i_8_2099, i_8_2100, i_8_2101, i_8_2102, i_8_2103, i_8_2104, i_8_2105, i_8_2106, i_8_2107, i_8_2108, i_8_2109, i_8_2110, i_8_2111, i_8_2112, i_8_2113, i_8_2114, i_8_2115, i_8_2116, i_8_2117, i_8_2118, i_8_2119, i_8_2120, i_8_2121, i_8_2122, i_8_2123, i_8_2124, i_8_2125, i_8_2126, i_8_2127, i_8_2128, i_8_2129, i_8_2130, i_8_2131, i_8_2132, i_8_2133, i_8_2134, i_8_2135, i_8_2136, i_8_2137, i_8_2138, i_8_2139, i_8_2140, i_8_2141, i_8_2142, i_8_2143, i_8_2144, i_8_2145, i_8_2146, i_8_2147, i_8_2148, i_8_2149, i_8_2150, i_8_2151, i_8_2152, i_8_2153, i_8_2154, i_8_2155, i_8_2156, i_8_2157, i_8_2158, i_8_2159, i_8_2160, i_8_2161, i_8_2162, i_8_2163, i_8_2164, i_8_2165, i_8_2166, i_8_2167, i_8_2168, i_8_2169, i_8_2170, i_8_2171, i_8_2172, i_8_2173, i_8_2174, i_8_2175, i_8_2176, i_8_2177, i_8_2178, i_8_2179, i_8_2180, i_8_2181, i_8_2182, i_8_2183, i_8_2184, i_8_2185, i_8_2186, i_8_2187, i_8_2188, i_8_2189, i_8_2190, i_8_2191, i_8_2192, i_8_2193, i_8_2194, i_8_2195, i_8_2196, i_8_2197, i_8_2198, i_8_2199, i_8_2200, i_8_2201, i_8_2202, i_8_2203, i_8_2204, i_8_2205, i_8_2206, i_8_2207, i_8_2208, i_8_2209, i_8_2210, i_8_2211, i_8_2212, i_8_2213, i_8_2214, i_8_2215, i_8_2216, i_8_2217, i_8_2218, i_8_2219, i_8_2220, i_8_2221, i_8_2222, i_8_2223, i_8_2224, i_8_2225, i_8_2226, i_8_2227, i_8_2228, i_8_2229, i_8_2230, i_8_2231, i_8_2232, i_8_2233, i_8_2234, i_8_2235, i_8_2236, i_8_2237, i_8_2238, i_8_2239, i_8_2240, i_8_2241, i_8_2242, i_8_2243, i_8_2244, i_8_2245, i_8_2246, i_8_2247, i_8_2248, i_8_2249, i_8_2250, i_8_2251, i_8_2252, i_8_2253, i_8_2254, i_8_2255, i_8_2256, i_8_2257, i_8_2258, i_8_2259, i_8_2260, i_8_2261, i_8_2262, i_8_2263, i_8_2264, i_8_2265, i_8_2266, i_8_2267, i_8_2268, i_8_2269, i_8_2270, i_8_2271, i_8_2272, i_8_2273, i_8_2274, i_8_2275, i_8_2276, i_8_2277, i_8_2278, i_8_2279, i_8_2280, i_8_2281, i_8_2282, i_8_2283, i_8_2284, i_8_2285, i_8_2286, i_8_2287, i_8_2288, i_8_2289, i_8_2290, i_8_2291, i_8_2292, i_8_2293, i_8_2294, i_8_2295, i_8_2296, i_8_2297, i_8_2298, i_8_2299, i_8_2300, i_8_2301, i_8_2302, i_8_2303;
  reg dly1, dly2;
  wire o_8_0, o_8_1, o_8_2, o_8_3, o_8_4, o_8_5, o_8_6, o_8_7, o_8_8, o_8_9, o_8_10, o_8_11, o_8_12, o_8_13, o_8_14, o_8_15, o_8_16, o_8_17, o_8_18, o_8_19, o_8_20, o_8_21, o_8_22, o_8_23, o_8_24, o_8_25, o_8_26, o_8_27, o_8_28, o_8_29, o_8_30, o_8_31, o_8_32, o_8_33, o_8_34, o_8_35, o_8_36, o_8_37, o_8_38, o_8_39, o_8_40, o_8_41, o_8_42, o_8_43, o_8_44, o_8_45, o_8_46, o_8_47, o_8_48, o_8_49, o_8_50, o_8_51, o_8_52, o_8_53, o_8_54, o_8_55, o_8_56, o_8_57, o_8_58, o_8_59, o_8_60, o_8_61, o_8_62, o_8_63, o_8_64, o_8_65, o_8_66, o_8_67, o_8_68, o_8_69, o_8_70, o_8_71, o_8_72, o_8_73, o_8_74, o_8_75, o_8_76, o_8_77, o_8_78, o_8_79, o_8_80, o_8_81, o_8_82, o_8_83, o_8_84, o_8_85, o_8_86, o_8_87, o_8_88, o_8_89, o_8_90, o_8_91, o_8_92, o_8_93, o_8_94, o_8_95, o_8_96, o_8_97, o_8_98, o_8_99, o_8_100, o_8_101, o_8_102, o_8_103, o_8_104, o_8_105, o_8_106, o_8_107, o_8_108, o_8_109, o_8_110, o_8_111, o_8_112, o_8_113, o_8_114, o_8_115, o_8_116, o_8_117, o_8_118, o_8_119, o_8_120, o_8_121, o_8_122, o_8_123, o_8_124, o_8_125, o_8_126, o_8_127, o_8_128, o_8_129, o_8_130, o_8_131, o_8_132, o_8_133, o_8_134, o_8_135, o_8_136, o_8_137, o_8_138, o_8_139, o_8_140, o_8_141, o_8_142, o_8_143, o_8_144, o_8_145, o_8_146, o_8_147, o_8_148, o_8_149, o_8_150, o_8_151, o_8_152, o_8_153, o_8_154, o_8_155, o_8_156, o_8_157, o_8_158, o_8_159, o_8_160, o_8_161, o_8_162, o_8_163, o_8_164, o_8_165, o_8_166, o_8_167, o_8_168, o_8_169, o_8_170, o_8_171, o_8_172, o_8_173, o_8_174, o_8_175, o_8_176, o_8_177, o_8_178, o_8_179, o_8_180, o_8_181, o_8_182, o_8_183, o_8_184, o_8_185, o_8_186, o_8_187, o_8_188, o_8_189, o_8_190, o_8_191, o_8_192, o_8_193, o_8_194, o_8_195, o_8_196, o_8_197, o_8_198, o_8_199, o_8_200, o_8_201, o_8_202, o_8_203, o_8_204, o_8_205, o_8_206, o_8_207, o_8_208, o_8_209, o_8_210, o_8_211, o_8_212, o_8_213, o_8_214, o_8_215, o_8_216, o_8_217, o_8_218, o_8_219, o_8_220, o_8_221, o_8_222, o_8_223, o_8_224, o_8_225, o_8_226, o_8_227, o_8_228, o_8_229, o_8_230, o_8_231, o_8_232, o_8_233, o_8_234, o_8_235, o_8_236, o_8_237, o_8_238, o_8_239, o_8_240, o_8_241, o_8_242, o_8_243, o_8_244, o_8_245, o_8_246, o_8_247, o_8_248, o_8_249, o_8_250, o_8_251, o_8_252, o_8_253, o_8_254, o_8_255, o_8_256, o_8_257, o_8_258, o_8_259, o_8_260, o_8_261, o_8_262, o_8_263, o_8_264, o_8_265, o_8_266, o_8_267, o_8_268, o_8_269, o_8_270, o_8_271, o_8_272, o_8_273, o_8_274, o_8_275, o_8_276, o_8_277, o_8_278, o_8_279, o_8_280, o_8_281, o_8_282, o_8_283, o_8_284, o_8_285, o_8_286, o_8_287, o_8_288, o_8_289, o_8_290, o_8_291, o_8_292, o_8_293, o_8_294, o_8_295, o_8_296, o_8_297, o_8_298, o_8_299, o_8_300, o_8_301, o_8_302, o_8_303, o_8_304, o_8_305, o_8_306, o_8_307, o_8_308, o_8_309, o_8_310, o_8_311, o_8_312, o_8_313, o_8_314, o_8_315, o_8_316, o_8_317, o_8_318, o_8_319, o_8_320, o_8_321, o_8_322, o_8_323, o_8_324, o_8_325, o_8_326, o_8_327, o_8_328, o_8_329, o_8_330, o_8_331, o_8_332, o_8_333, o_8_334, o_8_335, o_8_336, o_8_337, o_8_338, o_8_339, o_8_340, o_8_341, o_8_342, o_8_343, o_8_344, o_8_345, o_8_346, o_8_347, o_8_348, o_8_349, o_8_350, o_8_351, o_8_352, o_8_353, o_8_354, o_8_355, o_8_356, o_8_357, o_8_358, o_8_359, o_8_360, o_8_361, o_8_362, o_8_363, o_8_364, o_8_365, o_8_366, o_8_367, o_8_368, o_8_369, o_8_370, o_8_371, o_8_372, o_8_373, o_8_374, o_8_375, o_8_376, o_8_377, o_8_378, o_8_379, o_8_380, o_8_381, o_8_382, o_8_383, o_8_384, o_8_385, o_8_386, o_8_387, o_8_388, o_8_389, o_8_390, o_8_391, o_8_392, o_8_393, o_8_394, o_8_395, o_8_396, o_8_397, o_8_398, o_8_399, o_8_400, o_8_401, o_8_402, o_8_403, o_8_404, o_8_405, o_8_406, o_8_407, o_8_408, o_8_409, o_8_410, o_8_411, o_8_412, o_8_413, o_8_414, o_8_415, o_8_416, o_8_417, o_8_418, o_8_419, o_8_420, o_8_421, o_8_422, o_8_423, o_8_424, o_8_425, o_8_426, o_8_427, o_8_428, o_8_429, o_8_430, o_8_431, o_8_432, o_8_433, o_8_434, o_8_435, o_8_436, o_8_437, o_8_438, o_8_439, o_8_440, o_8_441, o_8_442, o_8_443, o_8_444, o_8_445, o_8_446, o_8_447, o_8_448, o_8_449, o_8_450, o_8_451, o_8_452, o_8_453, o_8_454, o_8_455, o_8_456, o_8_457, o_8_458, o_8_459, o_8_460, o_8_461, o_8_462, o_8_463, o_8_464, o_8_465, o_8_466, o_8_467, o_8_468, o_8_469, o_8_470, o_8_471, o_8_472, o_8_473, o_8_474, o_8_475, o_8_476, o_8_477, o_8_478, o_8_479, o_8_480, o_8_481, o_8_482, o_8_483, o_8_484, o_8_485, o_8_486, o_8_487, o_8_488, o_8_489, o_8_490, o_8_491, o_8_492, o_8_493, o_8_494, o_8_495, o_8_496, o_8_497, o_8_498, o_8_499, o_8_500, o_8_501, o_8_502, o_8_503, o_8_504, o_8_505, o_8_506, o_8_507, o_8_508, o_8_509, o_8_510, o_8_511;

  kernel_8 kernel_nulla( i_8_0, i_8_1, i_8_2, i_8_3, i_8_4, i_8_5, i_8_6, i_8_7, i_8_8, i_8_9, i_8_10, i_8_11, i_8_12, i_8_13, i_8_14, i_8_15, i_8_16, i_8_17, i_8_18, i_8_19, i_8_20, i_8_21, i_8_22, i_8_23, i_8_24, i_8_25, i_8_26, i_8_27, i_8_28, i_8_29, i_8_30, i_8_31, i_8_32, i_8_33, i_8_34, i_8_35, i_8_36, i_8_37, i_8_38, i_8_39, i_8_40, i_8_41, i_8_42, i_8_43, i_8_44, i_8_45, i_8_46, i_8_47, i_8_48, i_8_49, i_8_50, i_8_51, i_8_52, i_8_53, i_8_54, i_8_55, i_8_56, i_8_57, i_8_58, i_8_59, i_8_60, i_8_61, i_8_62, i_8_63, i_8_64, i_8_65, i_8_66, i_8_67, i_8_68, i_8_69, i_8_70, i_8_71, i_8_72, i_8_73, i_8_74, i_8_75, i_8_76, i_8_77, i_8_78, i_8_79, i_8_80, i_8_81, i_8_82, i_8_83, i_8_84, i_8_85, i_8_86, i_8_87, i_8_88, i_8_89, i_8_90, i_8_91, i_8_92, i_8_93, i_8_94, i_8_95, i_8_96, i_8_97, i_8_98, i_8_99, i_8_100, i_8_101, i_8_102, i_8_103, i_8_104, i_8_105, i_8_106, i_8_107, i_8_108, i_8_109, i_8_110, i_8_111, i_8_112, i_8_113, i_8_114, i_8_115, i_8_116, i_8_117, i_8_118, i_8_119, i_8_120, i_8_121, i_8_122, i_8_123, i_8_124, i_8_125, i_8_126, i_8_127, i_8_128, i_8_129, i_8_130, i_8_131, i_8_132, i_8_133, i_8_134, i_8_135, i_8_136, i_8_137, i_8_138, i_8_139, i_8_140, i_8_141, i_8_142, i_8_143, i_8_144, i_8_145, i_8_146, i_8_147, i_8_148, i_8_149, i_8_150, i_8_151, i_8_152, i_8_153, i_8_154, i_8_155, i_8_156, i_8_157, i_8_158, i_8_159, i_8_160, i_8_161, i_8_162, i_8_163, i_8_164, i_8_165, i_8_166, i_8_167, i_8_168, i_8_169, i_8_170, i_8_171, i_8_172, i_8_173, i_8_174, i_8_175, i_8_176, i_8_177, i_8_178, i_8_179, i_8_180, i_8_181, i_8_182, i_8_183, i_8_184, i_8_185, i_8_186, i_8_187, i_8_188, i_8_189, i_8_190, i_8_191, i_8_192, i_8_193, i_8_194, i_8_195, i_8_196, i_8_197, i_8_198, i_8_199, i_8_200, i_8_201, i_8_202, i_8_203, i_8_204, i_8_205, i_8_206, i_8_207, i_8_208, i_8_209, i_8_210, i_8_211, i_8_212, i_8_213, i_8_214, i_8_215, i_8_216, i_8_217, i_8_218, i_8_219, i_8_220, i_8_221, i_8_222, i_8_223, i_8_224, i_8_225, i_8_226, i_8_227, i_8_228, i_8_229, i_8_230, i_8_231, i_8_232, i_8_233, i_8_234, i_8_235, i_8_236, i_8_237, i_8_238, i_8_239, i_8_240, i_8_241, i_8_242, i_8_243, i_8_244, i_8_245, i_8_246, i_8_247, i_8_248, i_8_249, i_8_250, i_8_251, i_8_252, i_8_253, i_8_254, i_8_255, i_8_256, i_8_257, i_8_258, i_8_259, i_8_260, i_8_261, i_8_262, i_8_263, i_8_264, i_8_265, i_8_266, i_8_267, i_8_268, i_8_269, i_8_270, i_8_271, i_8_272, i_8_273, i_8_274, i_8_275, i_8_276, i_8_277, i_8_278, i_8_279, i_8_280, i_8_281, i_8_282, i_8_283, i_8_284, i_8_285, i_8_286, i_8_287, i_8_288, i_8_289, i_8_290, i_8_291, i_8_292, i_8_293, i_8_294, i_8_295, i_8_296, i_8_297, i_8_298, i_8_299, i_8_300, i_8_301, i_8_302, i_8_303, i_8_304, i_8_305, i_8_306, i_8_307, i_8_308, i_8_309, i_8_310, i_8_311, i_8_312, i_8_313, i_8_314, i_8_315, i_8_316, i_8_317, i_8_318, i_8_319, i_8_320, i_8_321, i_8_322, i_8_323, i_8_324, i_8_325, i_8_326, i_8_327, i_8_328, i_8_329, i_8_330, i_8_331, i_8_332, i_8_333, i_8_334, i_8_335, i_8_336, i_8_337, i_8_338, i_8_339, i_8_340, i_8_341, i_8_342, i_8_343, i_8_344, i_8_345, i_8_346, i_8_347, i_8_348, i_8_349, i_8_350, i_8_351, i_8_352, i_8_353, i_8_354, i_8_355, i_8_356, i_8_357, i_8_358, i_8_359, i_8_360, i_8_361, i_8_362, i_8_363, i_8_364, i_8_365, i_8_366, i_8_367, i_8_368, i_8_369, i_8_370, i_8_371, i_8_372, i_8_373, i_8_374, i_8_375, i_8_376, i_8_377, i_8_378, i_8_379, i_8_380, i_8_381, i_8_382, i_8_383, i_8_384, i_8_385, i_8_386, i_8_387, i_8_388, i_8_389, i_8_390, i_8_391, i_8_392, i_8_393, i_8_394, i_8_395, i_8_396, i_8_397, i_8_398, i_8_399, i_8_400, i_8_401, i_8_402, i_8_403, i_8_404, i_8_405, i_8_406, i_8_407, i_8_408, i_8_409, i_8_410, i_8_411, i_8_412, i_8_413, i_8_414, i_8_415, i_8_416, i_8_417, i_8_418, i_8_419, i_8_420, i_8_421, i_8_422, i_8_423, i_8_424, i_8_425, i_8_426, i_8_427, i_8_428, i_8_429, i_8_430, i_8_431, i_8_432, i_8_433, i_8_434, i_8_435, i_8_436, i_8_437, i_8_438, i_8_439, i_8_440, i_8_441, i_8_442, i_8_443, i_8_444, i_8_445, i_8_446, i_8_447, i_8_448, i_8_449, i_8_450, i_8_451, i_8_452, i_8_453, i_8_454, i_8_455, i_8_456, i_8_457, i_8_458, i_8_459, i_8_460, i_8_461, i_8_462, i_8_463, i_8_464, i_8_465, i_8_466, i_8_467, i_8_468, i_8_469, i_8_470, i_8_471, i_8_472, i_8_473, i_8_474, i_8_475, i_8_476, i_8_477, i_8_478, i_8_479, i_8_480, i_8_481, i_8_482, i_8_483, i_8_484, i_8_485, i_8_486, i_8_487, i_8_488, i_8_489, i_8_490, i_8_491, i_8_492, i_8_493, i_8_494, i_8_495, i_8_496, i_8_497, i_8_498, i_8_499, i_8_500, i_8_501, i_8_502, i_8_503, i_8_504, i_8_505, i_8_506, i_8_507, i_8_508, i_8_509, i_8_510, i_8_511, i_8_512, i_8_513, i_8_514, i_8_515, i_8_516, i_8_517, i_8_518, i_8_519, i_8_520, i_8_521, i_8_522, i_8_523, i_8_524, i_8_525, i_8_526, i_8_527, i_8_528, i_8_529, i_8_530, i_8_531, i_8_532, i_8_533, i_8_534, i_8_535, i_8_536, i_8_537, i_8_538, i_8_539, i_8_540, i_8_541, i_8_542, i_8_543, i_8_544, i_8_545, i_8_546, i_8_547, i_8_548, i_8_549, i_8_550, i_8_551, i_8_552, i_8_553, i_8_554, i_8_555, i_8_556, i_8_557, i_8_558, i_8_559, i_8_560, i_8_561, i_8_562, i_8_563, i_8_564, i_8_565, i_8_566, i_8_567, i_8_568, i_8_569, i_8_570, i_8_571, i_8_572, i_8_573, i_8_574, i_8_575, i_8_576, i_8_577, i_8_578, i_8_579, i_8_580, i_8_581, i_8_582, i_8_583, i_8_584, i_8_585, i_8_586, i_8_587, i_8_588, i_8_589, i_8_590, i_8_591, i_8_592, i_8_593, i_8_594, i_8_595, i_8_596, i_8_597, i_8_598, i_8_599, i_8_600, i_8_601, i_8_602, i_8_603, i_8_604, i_8_605, i_8_606, i_8_607, i_8_608, i_8_609, i_8_610, i_8_611, i_8_612, i_8_613, i_8_614, i_8_615, i_8_616, i_8_617, i_8_618, i_8_619, i_8_620, i_8_621, i_8_622, i_8_623, i_8_624, i_8_625, i_8_626, i_8_627, i_8_628, i_8_629, i_8_630, i_8_631, i_8_632, i_8_633, i_8_634, i_8_635, i_8_636, i_8_637, i_8_638, i_8_639, i_8_640, i_8_641, i_8_642, i_8_643, i_8_644, i_8_645, i_8_646, i_8_647, i_8_648, i_8_649, i_8_650, i_8_651, i_8_652, i_8_653, i_8_654, i_8_655, i_8_656, i_8_657, i_8_658, i_8_659, i_8_660, i_8_661, i_8_662, i_8_663, i_8_664, i_8_665, i_8_666, i_8_667, i_8_668, i_8_669, i_8_670, i_8_671, i_8_672, i_8_673, i_8_674, i_8_675, i_8_676, i_8_677, i_8_678, i_8_679, i_8_680, i_8_681, i_8_682, i_8_683, i_8_684, i_8_685, i_8_686, i_8_687, i_8_688, i_8_689, i_8_690, i_8_691, i_8_692, i_8_693, i_8_694, i_8_695, i_8_696, i_8_697, i_8_698, i_8_699, i_8_700, i_8_701, i_8_702, i_8_703, i_8_704, i_8_705, i_8_706, i_8_707, i_8_708, i_8_709, i_8_710, i_8_711, i_8_712, i_8_713, i_8_714, i_8_715, i_8_716, i_8_717, i_8_718, i_8_719, i_8_720, i_8_721, i_8_722, i_8_723, i_8_724, i_8_725, i_8_726, i_8_727, i_8_728, i_8_729, i_8_730, i_8_731, i_8_732, i_8_733, i_8_734, i_8_735, i_8_736, i_8_737, i_8_738, i_8_739, i_8_740, i_8_741, i_8_742, i_8_743, i_8_744, i_8_745, i_8_746, i_8_747, i_8_748, i_8_749, i_8_750, i_8_751, i_8_752, i_8_753, i_8_754, i_8_755, i_8_756, i_8_757, i_8_758, i_8_759, i_8_760, i_8_761, i_8_762, i_8_763, i_8_764, i_8_765, i_8_766, i_8_767, i_8_768, i_8_769, i_8_770, i_8_771, i_8_772, i_8_773, i_8_774, i_8_775, i_8_776, i_8_777, i_8_778, i_8_779, i_8_780, i_8_781, i_8_782, i_8_783, i_8_784, i_8_785, i_8_786, i_8_787, i_8_788, i_8_789, i_8_790, i_8_791, i_8_792, i_8_793, i_8_794, i_8_795, i_8_796, i_8_797, i_8_798, i_8_799, i_8_800, i_8_801, i_8_802, i_8_803, i_8_804, i_8_805, i_8_806, i_8_807, i_8_808, i_8_809, i_8_810, i_8_811, i_8_812, i_8_813, i_8_814, i_8_815, i_8_816, i_8_817, i_8_818, i_8_819, i_8_820, i_8_821, i_8_822, i_8_823, i_8_824, i_8_825, i_8_826, i_8_827, i_8_828, i_8_829, i_8_830, i_8_831, i_8_832, i_8_833, i_8_834, i_8_835, i_8_836, i_8_837, i_8_838, i_8_839, i_8_840, i_8_841, i_8_842, i_8_843, i_8_844, i_8_845, i_8_846, i_8_847, i_8_848, i_8_849, i_8_850, i_8_851, i_8_852, i_8_853, i_8_854, i_8_855, i_8_856, i_8_857, i_8_858, i_8_859, i_8_860, i_8_861, i_8_862, i_8_863, i_8_864, i_8_865, i_8_866, i_8_867, i_8_868, i_8_869, i_8_870, i_8_871, i_8_872, i_8_873, i_8_874, i_8_875, i_8_876, i_8_877, i_8_878, i_8_879, i_8_880, i_8_881, i_8_882, i_8_883, i_8_884, i_8_885, i_8_886, i_8_887, i_8_888, i_8_889, i_8_890, i_8_891, i_8_892, i_8_893, i_8_894, i_8_895, i_8_896, i_8_897, i_8_898, i_8_899, i_8_900, i_8_901, i_8_902, i_8_903, i_8_904, i_8_905, i_8_906, i_8_907, i_8_908, i_8_909, i_8_910, i_8_911, i_8_912, i_8_913, i_8_914, i_8_915, i_8_916, i_8_917, i_8_918, i_8_919, i_8_920, i_8_921, i_8_922, i_8_923, i_8_924, i_8_925, i_8_926, i_8_927, i_8_928, i_8_929, i_8_930, i_8_931, i_8_932, i_8_933, i_8_934, i_8_935, i_8_936, i_8_937, i_8_938, i_8_939, i_8_940, i_8_941, i_8_942, i_8_943, i_8_944, i_8_945, i_8_946, i_8_947, i_8_948, i_8_949, i_8_950, i_8_951, i_8_952, i_8_953, i_8_954, i_8_955, i_8_956, i_8_957, i_8_958, i_8_959, i_8_960, i_8_961, i_8_962, i_8_963, i_8_964, i_8_965, i_8_966, i_8_967, i_8_968, i_8_969, i_8_970, i_8_971, i_8_972, i_8_973, i_8_974, i_8_975, i_8_976, i_8_977, i_8_978, i_8_979, i_8_980, i_8_981, i_8_982, i_8_983, i_8_984, i_8_985, i_8_986, i_8_987, i_8_988, i_8_989, i_8_990, i_8_991, i_8_992, i_8_993, i_8_994, i_8_995, i_8_996, i_8_997, i_8_998, i_8_999, i_8_1000, i_8_1001, i_8_1002, i_8_1003, i_8_1004, i_8_1005, i_8_1006, i_8_1007, i_8_1008, i_8_1009, i_8_1010, i_8_1011, i_8_1012, i_8_1013, i_8_1014, i_8_1015, i_8_1016, i_8_1017, i_8_1018, i_8_1019, i_8_1020, i_8_1021, i_8_1022, i_8_1023, i_8_1024, i_8_1025, i_8_1026, i_8_1027, i_8_1028, i_8_1029, i_8_1030, i_8_1031, i_8_1032, i_8_1033, i_8_1034, i_8_1035, i_8_1036, i_8_1037, i_8_1038, i_8_1039, i_8_1040, i_8_1041, i_8_1042, i_8_1043, i_8_1044, i_8_1045, i_8_1046, i_8_1047, i_8_1048, i_8_1049, i_8_1050, i_8_1051, i_8_1052, i_8_1053, i_8_1054, i_8_1055, i_8_1056, i_8_1057, i_8_1058, i_8_1059, i_8_1060, i_8_1061, i_8_1062, i_8_1063, i_8_1064, i_8_1065, i_8_1066, i_8_1067, i_8_1068, i_8_1069, i_8_1070, i_8_1071, i_8_1072, i_8_1073, i_8_1074, i_8_1075, i_8_1076, i_8_1077, i_8_1078, i_8_1079, i_8_1080, i_8_1081, i_8_1082, i_8_1083, i_8_1084, i_8_1085, i_8_1086, i_8_1087, i_8_1088, i_8_1089, i_8_1090, i_8_1091, i_8_1092, i_8_1093, i_8_1094, i_8_1095, i_8_1096, i_8_1097, i_8_1098, i_8_1099, i_8_1100, i_8_1101, i_8_1102, i_8_1103, i_8_1104, i_8_1105, i_8_1106, i_8_1107, i_8_1108, i_8_1109, i_8_1110, i_8_1111, i_8_1112, i_8_1113, i_8_1114, i_8_1115, i_8_1116, i_8_1117, i_8_1118, i_8_1119, i_8_1120, i_8_1121, i_8_1122, i_8_1123, i_8_1124, i_8_1125, i_8_1126, i_8_1127, i_8_1128, i_8_1129, i_8_1130, i_8_1131, i_8_1132, i_8_1133, i_8_1134, i_8_1135, i_8_1136, i_8_1137, i_8_1138, i_8_1139, i_8_1140, i_8_1141, i_8_1142, i_8_1143, i_8_1144, i_8_1145, i_8_1146, i_8_1147, i_8_1148, i_8_1149, i_8_1150, i_8_1151, i_8_1152, i_8_1153, i_8_1154, i_8_1155, i_8_1156, i_8_1157, i_8_1158, i_8_1159, i_8_1160, i_8_1161, i_8_1162, i_8_1163, i_8_1164, i_8_1165, i_8_1166, i_8_1167, i_8_1168, i_8_1169, i_8_1170, i_8_1171, i_8_1172, i_8_1173, i_8_1174, i_8_1175, i_8_1176, i_8_1177, i_8_1178, i_8_1179, i_8_1180, i_8_1181, i_8_1182, i_8_1183, i_8_1184, i_8_1185, i_8_1186, i_8_1187, i_8_1188, i_8_1189, i_8_1190, i_8_1191, i_8_1192, i_8_1193, i_8_1194, i_8_1195, i_8_1196, i_8_1197, i_8_1198, i_8_1199, i_8_1200, i_8_1201, i_8_1202, i_8_1203, i_8_1204, i_8_1205, i_8_1206, i_8_1207, i_8_1208, i_8_1209, i_8_1210, i_8_1211, i_8_1212, i_8_1213, i_8_1214, i_8_1215, i_8_1216, i_8_1217, i_8_1218, i_8_1219, i_8_1220, i_8_1221, i_8_1222, i_8_1223, i_8_1224, i_8_1225, i_8_1226, i_8_1227, i_8_1228, i_8_1229, i_8_1230, i_8_1231, i_8_1232, i_8_1233, i_8_1234, i_8_1235, i_8_1236, i_8_1237, i_8_1238, i_8_1239, i_8_1240, i_8_1241, i_8_1242, i_8_1243, i_8_1244, i_8_1245, i_8_1246, i_8_1247, i_8_1248, i_8_1249, i_8_1250, i_8_1251, i_8_1252, i_8_1253, i_8_1254, i_8_1255, i_8_1256, i_8_1257, i_8_1258, i_8_1259, i_8_1260, i_8_1261, i_8_1262, i_8_1263, i_8_1264, i_8_1265, i_8_1266, i_8_1267, i_8_1268, i_8_1269, i_8_1270, i_8_1271, i_8_1272, i_8_1273, i_8_1274, i_8_1275, i_8_1276, i_8_1277, i_8_1278, i_8_1279, i_8_1280, i_8_1281, i_8_1282, i_8_1283, i_8_1284, i_8_1285, i_8_1286, i_8_1287, i_8_1288, i_8_1289, i_8_1290, i_8_1291, i_8_1292, i_8_1293, i_8_1294, i_8_1295, i_8_1296, i_8_1297, i_8_1298, i_8_1299, i_8_1300, i_8_1301, i_8_1302, i_8_1303, i_8_1304, i_8_1305, i_8_1306, i_8_1307, i_8_1308, i_8_1309, i_8_1310, i_8_1311, i_8_1312, i_8_1313, i_8_1314, i_8_1315, i_8_1316, i_8_1317, i_8_1318, i_8_1319, i_8_1320, i_8_1321, i_8_1322, i_8_1323, i_8_1324, i_8_1325, i_8_1326, i_8_1327, i_8_1328, i_8_1329, i_8_1330, i_8_1331, i_8_1332, i_8_1333, i_8_1334, i_8_1335, i_8_1336, i_8_1337, i_8_1338, i_8_1339, i_8_1340, i_8_1341, i_8_1342, i_8_1343, i_8_1344, i_8_1345, i_8_1346, i_8_1347, i_8_1348, i_8_1349, i_8_1350, i_8_1351, i_8_1352, i_8_1353, i_8_1354, i_8_1355, i_8_1356, i_8_1357, i_8_1358, i_8_1359, i_8_1360, i_8_1361, i_8_1362, i_8_1363, i_8_1364, i_8_1365, i_8_1366, i_8_1367, i_8_1368, i_8_1369, i_8_1370, i_8_1371, i_8_1372, i_8_1373, i_8_1374, i_8_1375, i_8_1376, i_8_1377, i_8_1378, i_8_1379, i_8_1380, i_8_1381, i_8_1382, i_8_1383, i_8_1384, i_8_1385, i_8_1386, i_8_1387, i_8_1388, i_8_1389, i_8_1390, i_8_1391, i_8_1392, i_8_1393, i_8_1394, i_8_1395, i_8_1396, i_8_1397, i_8_1398, i_8_1399, i_8_1400, i_8_1401, i_8_1402, i_8_1403, i_8_1404, i_8_1405, i_8_1406, i_8_1407, i_8_1408, i_8_1409, i_8_1410, i_8_1411, i_8_1412, i_8_1413, i_8_1414, i_8_1415, i_8_1416, i_8_1417, i_8_1418, i_8_1419, i_8_1420, i_8_1421, i_8_1422, i_8_1423, i_8_1424, i_8_1425, i_8_1426, i_8_1427, i_8_1428, i_8_1429, i_8_1430, i_8_1431, i_8_1432, i_8_1433, i_8_1434, i_8_1435, i_8_1436, i_8_1437, i_8_1438, i_8_1439, i_8_1440, i_8_1441, i_8_1442, i_8_1443, i_8_1444, i_8_1445, i_8_1446, i_8_1447, i_8_1448, i_8_1449, i_8_1450, i_8_1451, i_8_1452, i_8_1453, i_8_1454, i_8_1455, i_8_1456, i_8_1457, i_8_1458, i_8_1459, i_8_1460, i_8_1461, i_8_1462, i_8_1463, i_8_1464, i_8_1465, i_8_1466, i_8_1467, i_8_1468, i_8_1469, i_8_1470, i_8_1471, i_8_1472, i_8_1473, i_8_1474, i_8_1475, i_8_1476, i_8_1477, i_8_1478, i_8_1479, i_8_1480, i_8_1481, i_8_1482, i_8_1483, i_8_1484, i_8_1485, i_8_1486, i_8_1487, i_8_1488, i_8_1489, i_8_1490, i_8_1491, i_8_1492, i_8_1493, i_8_1494, i_8_1495, i_8_1496, i_8_1497, i_8_1498, i_8_1499, i_8_1500, i_8_1501, i_8_1502, i_8_1503, i_8_1504, i_8_1505, i_8_1506, i_8_1507, i_8_1508, i_8_1509, i_8_1510, i_8_1511, i_8_1512, i_8_1513, i_8_1514, i_8_1515, i_8_1516, i_8_1517, i_8_1518, i_8_1519, i_8_1520, i_8_1521, i_8_1522, i_8_1523, i_8_1524, i_8_1525, i_8_1526, i_8_1527, i_8_1528, i_8_1529, i_8_1530, i_8_1531, i_8_1532, i_8_1533, i_8_1534, i_8_1535, i_8_1536, i_8_1537, i_8_1538, i_8_1539, i_8_1540, i_8_1541, i_8_1542, i_8_1543, i_8_1544, i_8_1545, i_8_1546, i_8_1547, i_8_1548, i_8_1549, i_8_1550, i_8_1551, i_8_1552, i_8_1553, i_8_1554, i_8_1555, i_8_1556, i_8_1557, i_8_1558, i_8_1559, i_8_1560, i_8_1561, i_8_1562, i_8_1563, i_8_1564, i_8_1565, i_8_1566, i_8_1567, i_8_1568, i_8_1569, i_8_1570, i_8_1571, i_8_1572, i_8_1573, i_8_1574, i_8_1575, i_8_1576, i_8_1577, i_8_1578, i_8_1579, i_8_1580, i_8_1581, i_8_1582, i_8_1583, i_8_1584, i_8_1585, i_8_1586, i_8_1587, i_8_1588, i_8_1589, i_8_1590, i_8_1591, i_8_1592, i_8_1593, i_8_1594, i_8_1595, i_8_1596, i_8_1597, i_8_1598, i_8_1599, i_8_1600, i_8_1601, i_8_1602, i_8_1603, i_8_1604, i_8_1605, i_8_1606, i_8_1607, i_8_1608, i_8_1609, i_8_1610, i_8_1611, i_8_1612, i_8_1613, i_8_1614, i_8_1615, i_8_1616, i_8_1617, i_8_1618, i_8_1619, i_8_1620, i_8_1621, i_8_1622, i_8_1623, i_8_1624, i_8_1625, i_8_1626, i_8_1627, i_8_1628, i_8_1629, i_8_1630, i_8_1631, i_8_1632, i_8_1633, i_8_1634, i_8_1635, i_8_1636, i_8_1637, i_8_1638, i_8_1639, i_8_1640, i_8_1641, i_8_1642, i_8_1643, i_8_1644, i_8_1645, i_8_1646, i_8_1647, i_8_1648, i_8_1649, i_8_1650, i_8_1651, i_8_1652, i_8_1653, i_8_1654, i_8_1655, i_8_1656, i_8_1657, i_8_1658, i_8_1659, i_8_1660, i_8_1661, i_8_1662, i_8_1663, i_8_1664, i_8_1665, i_8_1666, i_8_1667, i_8_1668, i_8_1669, i_8_1670, i_8_1671, i_8_1672, i_8_1673, i_8_1674, i_8_1675, i_8_1676, i_8_1677, i_8_1678, i_8_1679, i_8_1680, i_8_1681, i_8_1682, i_8_1683, i_8_1684, i_8_1685, i_8_1686, i_8_1687, i_8_1688, i_8_1689, i_8_1690, i_8_1691, i_8_1692, i_8_1693, i_8_1694, i_8_1695, i_8_1696, i_8_1697, i_8_1698, i_8_1699, i_8_1700, i_8_1701, i_8_1702, i_8_1703, i_8_1704, i_8_1705, i_8_1706, i_8_1707, i_8_1708, i_8_1709, i_8_1710, i_8_1711, i_8_1712, i_8_1713, i_8_1714, i_8_1715, i_8_1716, i_8_1717, i_8_1718, i_8_1719, i_8_1720, i_8_1721, i_8_1722, i_8_1723, i_8_1724, i_8_1725, i_8_1726, i_8_1727, i_8_1728, i_8_1729, i_8_1730, i_8_1731, i_8_1732, i_8_1733, i_8_1734, i_8_1735, i_8_1736, i_8_1737, i_8_1738, i_8_1739, i_8_1740, i_8_1741, i_8_1742, i_8_1743, i_8_1744, i_8_1745, i_8_1746, i_8_1747, i_8_1748, i_8_1749, i_8_1750, i_8_1751, i_8_1752, i_8_1753, i_8_1754, i_8_1755, i_8_1756, i_8_1757, i_8_1758, i_8_1759, i_8_1760, i_8_1761, i_8_1762, i_8_1763, i_8_1764, i_8_1765, i_8_1766, i_8_1767, i_8_1768, i_8_1769, i_8_1770, i_8_1771, i_8_1772, i_8_1773, i_8_1774, i_8_1775, i_8_1776, i_8_1777, i_8_1778, i_8_1779, i_8_1780, i_8_1781, i_8_1782, i_8_1783, i_8_1784, i_8_1785, i_8_1786, i_8_1787, i_8_1788, i_8_1789, i_8_1790, i_8_1791, i_8_1792, i_8_1793, i_8_1794, i_8_1795, i_8_1796, i_8_1797, i_8_1798, i_8_1799, i_8_1800, i_8_1801, i_8_1802, i_8_1803, i_8_1804, i_8_1805, i_8_1806, i_8_1807, i_8_1808, i_8_1809, i_8_1810, i_8_1811, i_8_1812, i_8_1813, i_8_1814, i_8_1815, i_8_1816, i_8_1817, i_8_1818, i_8_1819, i_8_1820, i_8_1821, i_8_1822, i_8_1823, i_8_1824, i_8_1825, i_8_1826, i_8_1827, i_8_1828, i_8_1829, i_8_1830, i_8_1831, i_8_1832, i_8_1833, i_8_1834, i_8_1835, i_8_1836, i_8_1837, i_8_1838, i_8_1839, i_8_1840, i_8_1841, i_8_1842, i_8_1843, i_8_1844, i_8_1845, i_8_1846, i_8_1847, i_8_1848, i_8_1849, i_8_1850, i_8_1851, i_8_1852, i_8_1853, i_8_1854, i_8_1855, i_8_1856, i_8_1857, i_8_1858, i_8_1859, i_8_1860, i_8_1861, i_8_1862, i_8_1863, i_8_1864, i_8_1865, i_8_1866, i_8_1867, i_8_1868, i_8_1869, i_8_1870, i_8_1871, i_8_1872, i_8_1873, i_8_1874, i_8_1875, i_8_1876, i_8_1877, i_8_1878, i_8_1879, i_8_1880, i_8_1881, i_8_1882, i_8_1883, i_8_1884, i_8_1885, i_8_1886, i_8_1887, i_8_1888, i_8_1889, i_8_1890, i_8_1891, i_8_1892, i_8_1893, i_8_1894, i_8_1895, i_8_1896, i_8_1897, i_8_1898, i_8_1899, i_8_1900, i_8_1901, i_8_1902, i_8_1903, i_8_1904, i_8_1905, i_8_1906, i_8_1907, i_8_1908, i_8_1909, i_8_1910, i_8_1911, i_8_1912, i_8_1913, i_8_1914, i_8_1915, i_8_1916, i_8_1917, i_8_1918, i_8_1919, i_8_1920, i_8_1921, i_8_1922, i_8_1923, i_8_1924, i_8_1925, i_8_1926, i_8_1927, i_8_1928, i_8_1929, i_8_1930, i_8_1931, i_8_1932, i_8_1933, i_8_1934, i_8_1935, i_8_1936, i_8_1937, i_8_1938, i_8_1939, i_8_1940, i_8_1941, i_8_1942, i_8_1943, i_8_1944, i_8_1945, i_8_1946, i_8_1947, i_8_1948, i_8_1949, i_8_1950, i_8_1951, i_8_1952, i_8_1953, i_8_1954, i_8_1955, i_8_1956, i_8_1957, i_8_1958, i_8_1959, i_8_1960, i_8_1961, i_8_1962, i_8_1963, i_8_1964, i_8_1965, i_8_1966, i_8_1967, i_8_1968, i_8_1969, i_8_1970, i_8_1971, i_8_1972, i_8_1973, i_8_1974, i_8_1975, i_8_1976, i_8_1977, i_8_1978, i_8_1979, i_8_1980, i_8_1981, i_8_1982, i_8_1983, i_8_1984, i_8_1985, i_8_1986, i_8_1987, i_8_1988, i_8_1989, i_8_1990, i_8_1991, i_8_1992, i_8_1993, i_8_1994, i_8_1995, i_8_1996, i_8_1997, i_8_1998, i_8_1999, i_8_2000, i_8_2001, i_8_2002, i_8_2003, i_8_2004, i_8_2005, i_8_2006, i_8_2007, i_8_2008, i_8_2009, i_8_2010, i_8_2011, i_8_2012, i_8_2013, i_8_2014, i_8_2015, i_8_2016, i_8_2017, i_8_2018, i_8_2019, i_8_2020, i_8_2021, i_8_2022, i_8_2023, i_8_2024, i_8_2025, i_8_2026, i_8_2027, i_8_2028, i_8_2029, i_8_2030, i_8_2031, i_8_2032, i_8_2033, i_8_2034, i_8_2035, i_8_2036, i_8_2037, i_8_2038, i_8_2039, i_8_2040, i_8_2041, i_8_2042, i_8_2043, i_8_2044, i_8_2045, i_8_2046, i_8_2047, i_8_2048, i_8_2049, i_8_2050, i_8_2051, i_8_2052, i_8_2053, i_8_2054, i_8_2055, i_8_2056, i_8_2057, i_8_2058, i_8_2059, i_8_2060, i_8_2061, i_8_2062, i_8_2063, i_8_2064, i_8_2065, i_8_2066, i_8_2067, i_8_2068, i_8_2069, i_8_2070, i_8_2071, i_8_2072, i_8_2073, i_8_2074, i_8_2075, i_8_2076, i_8_2077, i_8_2078, i_8_2079, i_8_2080, i_8_2081, i_8_2082, i_8_2083, i_8_2084, i_8_2085, i_8_2086, i_8_2087, i_8_2088, i_8_2089, i_8_2090, i_8_2091, i_8_2092, i_8_2093, i_8_2094, i_8_2095, i_8_2096, i_8_2097, i_8_2098, i_8_2099, i_8_2100, i_8_2101, i_8_2102, i_8_2103, i_8_2104, i_8_2105, i_8_2106, i_8_2107, i_8_2108, i_8_2109, i_8_2110, i_8_2111, i_8_2112, i_8_2113, i_8_2114, i_8_2115, i_8_2116, i_8_2117, i_8_2118, i_8_2119, i_8_2120, i_8_2121, i_8_2122, i_8_2123, i_8_2124, i_8_2125, i_8_2126, i_8_2127, i_8_2128, i_8_2129, i_8_2130, i_8_2131, i_8_2132, i_8_2133, i_8_2134, i_8_2135, i_8_2136, i_8_2137, i_8_2138, i_8_2139, i_8_2140, i_8_2141, i_8_2142, i_8_2143, i_8_2144, i_8_2145, i_8_2146, i_8_2147, i_8_2148, i_8_2149, i_8_2150, i_8_2151, i_8_2152, i_8_2153, i_8_2154, i_8_2155, i_8_2156, i_8_2157, i_8_2158, i_8_2159, i_8_2160, i_8_2161, i_8_2162, i_8_2163, i_8_2164, i_8_2165, i_8_2166, i_8_2167, i_8_2168, i_8_2169, i_8_2170, i_8_2171, i_8_2172, i_8_2173, i_8_2174, i_8_2175, i_8_2176, i_8_2177, i_8_2178, i_8_2179, i_8_2180, i_8_2181, i_8_2182, i_8_2183, i_8_2184, i_8_2185, i_8_2186, i_8_2187, i_8_2188, i_8_2189, i_8_2190, i_8_2191, i_8_2192, i_8_2193, i_8_2194, i_8_2195, i_8_2196, i_8_2197, i_8_2198, i_8_2199, i_8_2200, i_8_2201, i_8_2202, i_8_2203, i_8_2204, i_8_2205, i_8_2206, i_8_2207, i_8_2208, i_8_2209, i_8_2210, i_8_2211, i_8_2212, i_8_2213, i_8_2214, i_8_2215, i_8_2216, i_8_2217, i_8_2218, i_8_2219, i_8_2220, i_8_2221, i_8_2222, i_8_2223, i_8_2224, i_8_2225, i_8_2226, i_8_2227, i_8_2228, i_8_2229, i_8_2230, i_8_2231, i_8_2232, i_8_2233, i_8_2234, i_8_2235, i_8_2236, i_8_2237, i_8_2238, i_8_2239, i_8_2240, i_8_2241, i_8_2242, i_8_2243, i_8_2244, i_8_2245, i_8_2246, i_8_2247, i_8_2248, i_8_2249, i_8_2250, i_8_2251, i_8_2252, i_8_2253, i_8_2254, i_8_2255, i_8_2256, i_8_2257, i_8_2258, i_8_2259, i_8_2260, i_8_2261, i_8_2262, i_8_2263, i_8_2264, i_8_2265, i_8_2266, i_8_2267, i_8_2268, i_8_2269, i_8_2270, i_8_2271, i_8_2272, i_8_2273, i_8_2274, i_8_2275, i_8_2276, i_8_2277, i_8_2278, i_8_2279, i_8_2280, i_8_2281, i_8_2282, i_8_2283, i_8_2284, i_8_2285, i_8_2286, i_8_2287, i_8_2288, i_8_2289, i_8_2290, i_8_2291, i_8_2292, i_8_2293, i_8_2294, i_8_2295, i_8_2296, i_8_2297, i_8_2298, i_8_2299, i_8_2300, i_8_2301, i_8_2302, i_8_2303, o_8_0, o_8_1, o_8_2, o_8_3, o_8_4, o_8_5, o_8_6, o_8_7, o_8_8, o_8_9, o_8_10, o_8_11, o_8_12, o_8_13, o_8_14, o_8_15, o_8_16, o_8_17, o_8_18, o_8_19, o_8_20, o_8_21, o_8_22, o_8_23, o_8_24, o_8_25, o_8_26, o_8_27, o_8_28, o_8_29, o_8_30, o_8_31, o_8_32, o_8_33, o_8_34, o_8_35, o_8_36, o_8_37, o_8_38, o_8_39, o_8_40, o_8_41, o_8_42, o_8_43, o_8_44, o_8_45, o_8_46, o_8_47, o_8_48, o_8_49, o_8_50, o_8_51, o_8_52, o_8_53, o_8_54, o_8_55, o_8_56, o_8_57, o_8_58, o_8_59, o_8_60, o_8_61, o_8_62, o_8_63, o_8_64, o_8_65, o_8_66, o_8_67, o_8_68, o_8_69, o_8_70, o_8_71, o_8_72, o_8_73, o_8_74, o_8_75, o_8_76, o_8_77, o_8_78, o_8_79, o_8_80, o_8_81, o_8_82, o_8_83, o_8_84, o_8_85, o_8_86, o_8_87, o_8_88, o_8_89, o_8_90, o_8_91, o_8_92, o_8_93, o_8_94, o_8_95, o_8_96, o_8_97, o_8_98, o_8_99, o_8_100, o_8_101, o_8_102, o_8_103, o_8_104, o_8_105, o_8_106, o_8_107, o_8_108, o_8_109, o_8_110, o_8_111, o_8_112, o_8_113, o_8_114, o_8_115, o_8_116, o_8_117, o_8_118, o_8_119, o_8_120, o_8_121, o_8_122, o_8_123, o_8_124, o_8_125, o_8_126, o_8_127, o_8_128, o_8_129, o_8_130, o_8_131, o_8_132, o_8_133, o_8_134, o_8_135, o_8_136, o_8_137, o_8_138, o_8_139, o_8_140, o_8_141, o_8_142, o_8_143, o_8_144, o_8_145, o_8_146, o_8_147, o_8_148, o_8_149, o_8_150, o_8_151, o_8_152, o_8_153, o_8_154, o_8_155, o_8_156, o_8_157, o_8_158, o_8_159, o_8_160, o_8_161, o_8_162, o_8_163, o_8_164, o_8_165, o_8_166, o_8_167, o_8_168, o_8_169, o_8_170, o_8_171, o_8_172, o_8_173, o_8_174, o_8_175, o_8_176, o_8_177, o_8_178, o_8_179, o_8_180, o_8_181, o_8_182, o_8_183, o_8_184, o_8_185, o_8_186, o_8_187, o_8_188, o_8_189, o_8_190, o_8_191, o_8_192, o_8_193, o_8_194, o_8_195, o_8_196, o_8_197, o_8_198, o_8_199, o_8_200, o_8_201, o_8_202, o_8_203, o_8_204, o_8_205, o_8_206, o_8_207, o_8_208, o_8_209, o_8_210, o_8_211, o_8_212, o_8_213, o_8_214, o_8_215, o_8_216, o_8_217, o_8_218, o_8_219, o_8_220, o_8_221, o_8_222, o_8_223, o_8_224, o_8_225, o_8_226, o_8_227, o_8_228, o_8_229, o_8_230, o_8_231, o_8_232, o_8_233, o_8_234, o_8_235, o_8_236, o_8_237, o_8_238, o_8_239, o_8_240, o_8_241, o_8_242, o_8_243, o_8_244, o_8_245, o_8_246, o_8_247, o_8_248, o_8_249, o_8_250, o_8_251, o_8_252, o_8_253, o_8_254, o_8_255, o_8_256, o_8_257, o_8_258, o_8_259, o_8_260, o_8_261, o_8_262, o_8_263, o_8_264, o_8_265, o_8_266, o_8_267, o_8_268, o_8_269, o_8_270, o_8_271, o_8_272, o_8_273, o_8_274, o_8_275, o_8_276, o_8_277, o_8_278, o_8_279, o_8_280, o_8_281, o_8_282, o_8_283, o_8_284, o_8_285, o_8_286, o_8_287, o_8_288, o_8_289, o_8_290, o_8_291, o_8_292, o_8_293, o_8_294, o_8_295, o_8_296, o_8_297, o_8_298, o_8_299, o_8_300, o_8_301, o_8_302, o_8_303, o_8_304, o_8_305, o_8_306, o_8_307, o_8_308, o_8_309, o_8_310, o_8_311, o_8_312, o_8_313, o_8_314, o_8_315, o_8_316, o_8_317, o_8_318, o_8_319, o_8_320, o_8_321, o_8_322, o_8_323, o_8_324, o_8_325, o_8_326, o_8_327, o_8_328, o_8_329, o_8_330, o_8_331, o_8_332, o_8_333, o_8_334, o_8_335, o_8_336, o_8_337, o_8_338, o_8_339, o_8_340, o_8_341, o_8_342, o_8_343, o_8_344, o_8_345, o_8_346, o_8_347, o_8_348, o_8_349, o_8_350, o_8_351, o_8_352, o_8_353, o_8_354, o_8_355, o_8_356, o_8_357, o_8_358, o_8_359, o_8_360, o_8_361, o_8_362, o_8_363, o_8_364, o_8_365, o_8_366, o_8_367, o_8_368, o_8_369, o_8_370, o_8_371, o_8_372, o_8_373, o_8_374, o_8_375, o_8_376, o_8_377, o_8_378, o_8_379, o_8_380, o_8_381, o_8_382, o_8_383, o_8_384, o_8_385, o_8_386, o_8_387, o_8_388, o_8_389, o_8_390, o_8_391, o_8_392, o_8_393, o_8_394, o_8_395, o_8_396, o_8_397, o_8_398, o_8_399, o_8_400, o_8_401, o_8_402, o_8_403, o_8_404, o_8_405, o_8_406, o_8_407, o_8_408, o_8_409, o_8_410, o_8_411, o_8_412, o_8_413, o_8_414, o_8_415, o_8_416, o_8_417, o_8_418, o_8_419, o_8_420, o_8_421, o_8_422, o_8_423, o_8_424, o_8_425, o_8_426, o_8_427, o_8_428, o_8_429, o_8_430, o_8_431, o_8_432, o_8_433, o_8_434, o_8_435, o_8_436, o_8_437, o_8_438, o_8_439, o_8_440, o_8_441, o_8_442, o_8_443, o_8_444, o_8_445, o_8_446, o_8_447, o_8_448, o_8_449, o_8_450, o_8_451, o_8_452, o_8_453, o_8_454, o_8_455, o_8_456, o_8_457, o_8_458, o_8_459, o_8_460, o_8_461, o_8_462, o_8_463, o_8_464, o_8_465, o_8_466, o_8_467, o_8_468, o_8_469, o_8_470, o_8_471, o_8_472, o_8_473, o_8_474, o_8_475, o_8_476, o_8_477, o_8_478, o_8_479, o_8_480, o_8_481, o_8_482, o_8_483, o_8_484, o_8_485, o_8_486, o_8_487, o_8_488, o_8_489, o_8_490, o_8_491, o_8_492, o_8_493, o_8_494, o_8_495, o_8_496, o_8_497, o_8_498, o_8_499, o_8_500, o_8_501, o_8_502, o_8_503, o_8_504, o_8_505, o_8_506, o_8_507, o_8_508, o_8_509, o_8_510, o_8_511);

  always @ (posedge ap_clk)
    if (ap_rst)
      begin
        out_reg <= 0;
        i_8_0 <= 0;
        i_8_1 <= 0;
        i_8_2 <= 0;
        i_8_3 <= 0;
        i_8_4 <= 0;
        i_8_5 <= 0;
        i_8_6 <= 0;
        i_8_7 <= 0;
        i_8_8 <= 0;
        i_8_9 <= 0;
        i_8_10 <= 0;
        i_8_11 <= 0;
        i_8_12 <= 0;
        i_8_13 <= 0;
        i_8_14 <= 0;
        i_8_15 <= 0;
        i_8_16 <= 0;
        i_8_17 <= 0;
        i_8_18 <= 0;
        i_8_19 <= 0;
        i_8_20 <= 0;
        i_8_21 <= 0;
        i_8_22 <= 0;
        i_8_23 <= 0;
        i_8_24 <= 0;
        i_8_25 <= 0;
        i_8_26 <= 0;
        i_8_27 <= 0;
        i_8_28 <= 0;
        i_8_29 <= 0;
        i_8_30 <= 0;
        i_8_31 <= 0;
        i_8_32 <= 0;
        i_8_33 <= 0;
        i_8_34 <= 0;
        i_8_35 <= 0;
        i_8_36 <= 0;
        i_8_37 <= 0;
        i_8_38 <= 0;
        i_8_39 <= 0;
        i_8_40 <= 0;
        i_8_41 <= 0;
        i_8_42 <= 0;
        i_8_43 <= 0;
        i_8_44 <= 0;
        i_8_45 <= 0;
        i_8_46 <= 0;
        i_8_47 <= 0;
        i_8_48 <= 0;
        i_8_49 <= 0;
        i_8_50 <= 0;
        i_8_51 <= 0;
        i_8_52 <= 0;
        i_8_53 <= 0;
        i_8_54 <= 0;
        i_8_55 <= 0;
        i_8_56 <= 0;
        i_8_57 <= 0;
        i_8_58 <= 0;
        i_8_59 <= 0;
        i_8_60 <= 0;
        i_8_61 <= 0;
        i_8_62 <= 0;
        i_8_63 <= 0;
        i_8_64 <= 0;
        i_8_65 <= 0;
        i_8_66 <= 0;
        i_8_67 <= 0;
        i_8_68 <= 0;
        i_8_69 <= 0;
        i_8_70 <= 0;
        i_8_71 <= 0;
        i_8_72 <= 0;
        i_8_73 <= 0;
        i_8_74 <= 0;
        i_8_75 <= 0;
        i_8_76 <= 0;
        i_8_77 <= 0;
        i_8_78 <= 0;
        i_8_79 <= 0;
        i_8_80 <= 0;
        i_8_81 <= 0;
        i_8_82 <= 0;
        i_8_83 <= 0;
        i_8_84 <= 0;
        i_8_85 <= 0;
        i_8_86 <= 0;
        i_8_87 <= 0;
        i_8_88 <= 0;
        i_8_89 <= 0;
        i_8_90 <= 0;
        i_8_91 <= 0;
        i_8_92 <= 0;
        i_8_93 <= 0;
        i_8_94 <= 0;
        i_8_95 <= 0;
        i_8_96 <= 0;
        i_8_97 <= 0;
        i_8_98 <= 0;
        i_8_99 <= 0;
        i_8_100 <= 0;
        i_8_101 <= 0;
        i_8_102 <= 0;
        i_8_103 <= 0;
        i_8_104 <= 0;
        i_8_105 <= 0;
        i_8_106 <= 0;
        i_8_107 <= 0;
        i_8_108 <= 0;
        i_8_109 <= 0;
        i_8_110 <= 0;
        i_8_111 <= 0;
        i_8_112 <= 0;
        i_8_113 <= 0;
        i_8_114 <= 0;
        i_8_115 <= 0;
        i_8_116 <= 0;
        i_8_117 <= 0;
        i_8_118 <= 0;
        i_8_119 <= 0;
        i_8_120 <= 0;
        i_8_121 <= 0;
        i_8_122 <= 0;
        i_8_123 <= 0;
        i_8_124 <= 0;
        i_8_125 <= 0;
        i_8_126 <= 0;
        i_8_127 <= 0;
        i_8_128 <= 0;
        i_8_129 <= 0;
        i_8_130 <= 0;
        i_8_131 <= 0;
        i_8_132 <= 0;
        i_8_133 <= 0;
        i_8_134 <= 0;
        i_8_135 <= 0;
        i_8_136 <= 0;
        i_8_137 <= 0;
        i_8_138 <= 0;
        i_8_139 <= 0;
        i_8_140 <= 0;
        i_8_141 <= 0;
        i_8_142 <= 0;
        i_8_143 <= 0;
        i_8_144 <= 0;
        i_8_145 <= 0;
        i_8_146 <= 0;
        i_8_147 <= 0;
        i_8_148 <= 0;
        i_8_149 <= 0;
        i_8_150 <= 0;
        i_8_151 <= 0;
        i_8_152 <= 0;
        i_8_153 <= 0;
        i_8_154 <= 0;
        i_8_155 <= 0;
        i_8_156 <= 0;
        i_8_157 <= 0;
        i_8_158 <= 0;
        i_8_159 <= 0;
        i_8_160 <= 0;
        i_8_161 <= 0;
        i_8_162 <= 0;
        i_8_163 <= 0;
        i_8_164 <= 0;
        i_8_165 <= 0;
        i_8_166 <= 0;
        i_8_167 <= 0;
        i_8_168 <= 0;
        i_8_169 <= 0;
        i_8_170 <= 0;
        i_8_171 <= 0;
        i_8_172 <= 0;
        i_8_173 <= 0;
        i_8_174 <= 0;
        i_8_175 <= 0;
        i_8_176 <= 0;
        i_8_177 <= 0;
        i_8_178 <= 0;
        i_8_179 <= 0;
        i_8_180 <= 0;
        i_8_181 <= 0;
        i_8_182 <= 0;
        i_8_183 <= 0;
        i_8_184 <= 0;
        i_8_185 <= 0;
        i_8_186 <= 0;
        i_8_187 <= 0;
        i_8_188 <= 0;
        i_8_189 <= 0;
        i_8_190 <= 0;
        i_8_191 <= 0;
        i_8_192 <= 0;
        i_8_193 <= 0;
        i_8_194 <= 0;
        i_8_195 <= 0;
        i_8_196 <= 0;
        i_8_197 <= 0;
        i_8_198 <= 0;
        i_8_199 <= 0;
        i_8_200 <= 0;
        i_8_201 <= 0;
        i_8_202 <= 0;
        i_8_203 <= 0;
        i_8_204 <= 0;
        i_8_205 <= 0;
        i_8_206 <= 0;
        i_8_207 <= 0;
        i_8_208 <= 0;
        i_8_209 <= 0;
        i_8_210 <= 0;
        i_8_211 <= 0;
        i_8_212 <= 0;
        i_8_213 <= 0;
        i_8_214 <= 0;
        i_8_215 <= 0;
        i_8_216 <= 0;
        i_8_217 <= 0;
        i_8_218 <= 0;
        i_8_219 <= 0;
        i_8_220 <= 0;
        i_8_221 <= 0;
        i_8_222 <= 0;
        i_8_223 <= 0;
        i_8_224 <= 0;
        i_8_225 <= 0;
        i_8_226 <= 0;
        i_8_227 <= 0;
        i_8_228 <= 0;
        i_8_229 <= 0;
        i_8_230 <= 0;
        i_8_231 <= 0;
        i_8_232 <= 0;
        i_8_233 <= 0;
        i_8_234 <= 0;
        i_8_235 <= 0;
        i_8_236 <= 0;
        i_8_237 <= 0;
        i_8_238 <= 0;
        i_8_239 <= 0;
        i_8_240 <= 0;
        i_8_241 <= 0;
        i_8_242 <= 0;
        i_8_243 <= 0;
        i_8_244 <= 0;
        i_8_245 <= 0;
        i_8_246 <= 0;
        i_8_247 <= 0;
        i_8_248 <= 0;
        i_8_249 <= 0;
        i_8_250 <= 0;
        i_8_251 <= 0;
        i_8_252 <= 0;
        i_8_253 <= 0;
        i_8_254 <= 0;
        i_8_255 <= 0;
        i_8_256 <= 0;
        i_8_257 <= 0;
        i_8_258 <= 0;
        i_8_259 <= 0;
        i_8_260 <= 0;
        i_8_261 <= 0;
        i_8_262 <= 0;
        i_8_263 <= 0;
        i_8_264 <= 0;
        i_8_265 <= 0;
        i_8_266 <= 0;
        i_8_267 <= 0;
        i_8_268 <= 0;
        i_8_269 <= 0;
        i_8_270 <= 0;
        i_8_271 <= 0;
        i_8_272 <= 0;
        i_8_273 <= 0;
        i_8_274 <= 0;
        i_8_275 <= 0;
        i_8_276 <= 0;
        i_8_277 <= 0;
        i_8_278 <= 0;
        i_8_279 <= 0;
        i_8_280 <= 0;
        i_8_281 <= 0;
        i_8_282 <= 0;
        i_8_283 <= 0;
        i_8_284 <= 0;
        i_8_285 <= 0;
        i_8_286 <= 0;
        i_8_287 <= 0;
        i_8_288 <= 0;
        i_8_289 <= 0;
        i_8_290 <= 0;
        i_8_291 <= 0;
        i_8_292 <= 0;
        i_8_293 <= 0;
        i_8_294 <= 0;
        i_8_295 <= 0;
        i_8_296 <= 0;
        i_8_297 <= 0;
        i_8_298 <= 0;
        i_8_299 <= 0;
        i_8_300 <= 0;
        i_8_301 <= 0;
        i_8_302 <= 0;
        i_8_303 <= 0;
        i_8_304 <= 0;
        i_8_305 <= 0;
        i_8_306 <= 0;
        i_8_307 <= 0;
        i_8_308 <= 0;
        i_8_309 <= 0;
        i_8_310 <= 0;
        i_8_311 <= 0;
        i_8_312 <= 0;
        i_8_313 <= 0;
        i_8_314 <= 0;
        i_8_315 <= 0;
        i_8_316 <= 0;
        i_8_317 <= 0;
        i_8_318 <= 0;
        i_8_319 <= 0;
        i_8_320 <= 0;
        i_8_321 <= 0;
        i_8_322 <= 0;
        i_8_323 <= 0;
        i_8_324 <= 0;
        i_8_325 <= 0;
        i_8_326 <= 0;
        i_8_327 <= 0;
        i_8_328 <= 0;
        i_8_329 <= 0;
        i_8_330 <= 0;
        i_8_331 <= 0;
        i_8_332 <= 0;
        i_8_333 <= 0;
        i_8_334 <= 0;
        i_8_335 <= 0;
        i_8_336 <= 0;
        i_8_337 <= 0;
        i_8_338 <= 0;
        i_8_339 <= 0;
        i_8_340 <= 0;
        i_8_341 <= 0;
        i_8_342 <= 0;
        i_8_343 <= 0;
        i_8_344 <= 0;
        i_8_345 <= 0;
        i_8_346 <= 0;
        i_8_347 <= 0;
        i_8_348 <= 0;
        i_8_349 <= 0;
        i_8_350 <= 0;
        i_8_351 <= 0;
        i_8_352 <= 0;
        i_8_353 <= 0;
        i_8_354 <= 0;
        i_8_355 <= 0;
        i_8_356 <= 0;
        i_8_357 <= 0;
        i_8_358 <= 0;
        i_8_359 <= 0;
        i_8_360 <= 0;
        i_8_361 <= 0;
        i_8_362 <= 0;
        i_8_363 <= 0;
        i_8_364 <= 0;
        i_8_365 <= 0;
        i_8_366 <= 0;
        i_8_367 <= 0;
        i_8_368 <= 0;
        i_8_369 <= 0;
        i_8_370 <= 0;
        i_8_371 <= 0;
        i_8_372 <= 0;
        i_8_373 <= 0;
        i_8_374 <= 0;
        i_8_375 <= 0;
        i_8_376 <= 0;
        i_8_377 <= 0;
        i_8_378 <= 0;
        i_8_379 <= 0;
        i_8_380 <= 0;
        i_8_381 <= 0;
        i_8_382 <= 0;
        i_8_383 <= 0;
        i_8_384 <= 0;
        i_8_385 <= 0;
        i_8_386 <= 0;
        i_8_387 <= 0;
        i_8_388 <= 0;
        i_8_389 <= 0;
        i_8_390 <= 0;
        i_8_391 <= 0;
        i_8_392 <= 0;
        i_8_393 <= 0;
        i_8_394 <= 0;
        i_8_395 <= 0;
        i_8_396 <= 0;
        i_8_397 <= 0;
        i_8_398 <= 0;
        i_8_399 <= 0;
        i_8_400 <= 0;
        i_8_401 <= 0;
        i_8_402 <= 0;
        i_8_403 <= 0;
        i_8_404 <= 0;
        i_8_405 <= 0;
        i_8_406 <= 0;
        i_8_407 <= 0;
        i_8_408 <= 0;
        i_8_409 <= 0;
        i_8_410 <= 0;
        i_8_411 <= 0;
        i_8_412 <= 0;
        i_8_413 <= 0;
        i_8_414 <= 0;
        i_8_415 <= 0;
        i_8_416 <= 0;
        i_8_417 <= 0;
        i_8_418 <= 0;
        i_8_419 <= 0;
        i_8_420 <= 0;
        i_8_421 <= 0;
        i_8_422 <= 0;
        i_8_423 <= 0;
        i_8_424 <= 0;
        i_8_425 <= 0;
        i_8_426 <= 0;
        i_8_427 <= 0;
        i_8_428 <= 0;
        i_8_429 <= 0;
        i_8_430 <= 0;
        i_8_431 <= 0;
        i_8_432 <= 0;
        i_8_433 <= 0;
        i_8_434 <= 0;
        i_8_435 <= 0;
        i_8_436 <= 0;
        i_8_437 <= 0;
        i_8_438 <= 0;
        i_8_439 <= 0;
        i_8_440 <= 0;
        i_8_441 <= 0;
        i_8_442 <= 0;
        i_8_443 <= 0;
        i_8_444 <= 0;
        i_8_445 <= 0;
        i_8_446 <= 0;
        i_8_447 <= 0;
        i_8_448 <= 0;
        i_8_449 <= 0;
        i_8_450 <= 0;
        i_8_451 <= 0;
        i_8_452 <= 0;
        i_8_453 <= 0;
        i_8_454 <= 0;
        i_8_455 <= 0;
        i_8_456 <= 0;
        i_8_457 <= 0;
        i_8_458 <= 0;
        i_8_459 <= 0;
        i_8_460 <= 0;
        i_8_461 <= 0;
        i_8_462 <= 0;
        i_8_463 <= 0;
        i_8_464 <= 0;
        i_8_465 <= 0;
        i_8_466 <= 0;
        i_8_467 <= 0;
        i_8_468 <= 0;
        i_8_469 <= 0;
        i_8_470 <= 0;
        i_8_471 <= 0;
        i_8_472 <= 0;
        i_8_473 <= 0;
        i_8_474 <= 0;
        i_8_475 <= 0;
        i_8_476 <= 0;
        i_8_477 <= 0;
        i_8_478 <= 0;
        i_8_479 <= 0;
        i_8_480 <= 0;
        i_8_481 <= 0;
        i_8_482 <= 0;
        i_8_483 <= 0;
        i_8_484 <= 0;
        i_8_485 <= 0;
        i_8_486 <= 0;
        i_8_487 <= 0;
        i_8_488 <= 0;
        i_8_489 <= 0;
        i_8_490 <= 0;
        i_8_491 <= 0;
        i_8_492 <= 0;
        i_8_493 <= 0;
        i_8_494 <= 0;
        i_8_495 <= 0;
        i_8_496 <= 0;
        i_8_497 <= 0;
        i_8_498 <= 0;
        i_8_499 <= 0;
        i_8_500 <= 0;
        i_8_501 <= 0;
        i_8_502 <= 0;
        i_8_503 <= 0;
        i_8_504 <= 0;
        i_8_505 <= 0;
        i_8_506 <= 0;
        i_8_507 <= 0;
        i_8_508 <= 0;
        i_8_509 <= 0;
        i_8_510 <= 0;
        i_8_511 <= 0;
        i_8_512 <= 0;
        i_8_513 <= 0;
        i_8_514 <= 0;
        i_8_515 <= 0;
        i_8_516 <= 0;
        i_8_517 <= 0;
        i_8_518 <= 0;
        i_8_519 <= 0;
        i_8_520 <= 0;
        i_8_521 <= 0;
        i_8_522 <= 0;
        i_8_523 <= 0;
        i_8_524 <= 0;
        i_8_525 <= 0;
        i_8_526 <= 0;
        i_8_527 <= 0;
        i_8_528 <= 0;
        i_8_529 <= 0;
        i_8_530 <= 0;
        i_8_531 <= 0;
        i_8_532 <= 0;
        i_8_533 <= 0;
        i_8_534 <= 0;
        i_8_535 <= 0;
        i_8_536 <= 0;
        i_8_537 <= 0;
        i_8_538 <= 0;
        i_8_539 <= 0;
        i_8_540 <= 0;
        i_8_541 <= 0;
        i_8_542 <= 0;
        i_8_543 <= 0;
        i_8_544 <= 0;
        i_8_545 <= 0;
        i_8_546 <= 0;
        i_8_547 <= 0;
        i_8_548 <= 0;
        i_8_549 <= 0;
        i_8_550 <= 0;
        i_8_551 <= 0;
        i_8_552 <= 0;
        i_8_553 <= 0;
        i_8_554 <= 0;
        i_8_555 <= 0;
        i_8_556 <= 0;
        i_8_557 <= 0;
        i_8_558 <= 0;
        i_8_559 <= 0;
        i_8_560 <= 0;
        i_8_561 <= 0;
        i_8_562 <= 0;
        i_8_563 <= 0;
        i_8_564 <= 0;
        i_8_565 <= 0;
        i_8_566 <= 0;
        i_8_567 <= 0;
        i_8_568 <= 0;
        i_8_569 <= 0;
        i_8_570 <= 0;
        i_8_571 <= 0;
        i_8_572 <= 0;
        i_8_573 <= 0;
        i_8_574 <= 0;
        i_8_575 <= 0;
        i_8_576 <= 0;
        i_8_577 <= 0;
        i_8_578 <= 0;
        i_8_579 <= 0;
        i_8_580 <= 0;
        i_8_581 <= 0;
        i_8_582 <= 0;
        i_8_583 <= 0;
        i_8_584 <= 0;
        i_8_585 <= 0;
        i_8_586 <= 0;
        i_8_587 <= 0;
        i_8_588 <= 0;
        i_8_589 <= 0;
        i_8_590 <= 0;
        i_8_591 <= 0;
        i_8_592 <= 0;
        i_8_593 <= 0;
        i_8_594 <= 0;
        i_8_595 <= 0;
        i_8_596 <= 0;
        i_8_597 <= 0;
        i_8_598 <= 0;
        i_8_599 <= 0;
        i_8_600 <= 0;
        i_8_601 <= 0;
        i_8_602 <= 0;
        i_8_603 <= 0;
        i_8_604 <= 0;
        i_8_605 <= 0;
        i_8_606 <= 0;
        i_8_607 <= 0;
        i_8_608 <= 0;
        i_8_609 <= 0;
        i_8_610 <= 0;
        i_8_611 <= 0;
        i_8_612 <= 0;
        i_8_613 <= 0;
        i_8_614 <= 0;
        i_8_615 <= 0;
        i_8_616 <= 0;
        i_8_617 <= 0;
        i_8_618 <= 0;
        i_8_619 <= 0;
        i_8_620 <= 0;
        i_8_621 <= 0;
        i_8_622 <= 0;
        i_8_623 <= 0;
        i_8_624 <= 0;
        i_8_625 <= 0;
        i_8_626 <= 0;
        i_8_627 <= 0;
        i_8_628 <= 0;
        i_8_629 <= 0;
        i_8_630 <= 0;
        i_8_631 <= 0;
        i_8_632 <= 0;
        i_8_633 <= 0;
        i_8_634 <= 0;
        i_8_635 <= 0;
        i_8_636 <= 0;
        i_8_637 <= 0;
        i_8_638 <= 0;
        i_8_639 <= 0;
        i_8_640 <= 0;
        i_8_641 <= 0;
        i_8_642 <= 0;
        i_8_643 <= 0;
        i_8_644 <= 0;
        i_8_645 <= 0;
        i_8_646 <= 0;
        i_8_647 <= 0;
        i_8_648 <= 0;
        i_8_649 <= 0;
        i_8_650 <= 0;
        i_8_651 <= 0;
        i_8_652 <= 0;
        i_8_653 <= 0;
        i_8_654 <= 0;
        i_8_655 <= 0;
        i_8_656 <= 0;
        i_8_657 <= 0;
        i_8_658 <= 0;
        i_8_659 <= 0;
        i_8_660 <= 0;
        i_8_661 <= 0;
        i_8_662 <= 0;
        i_8_663 <= 0;
        i_8_664 <= 0;
        i_8_665 <= 0;
        i_8_666 <= 0;
        i_8_667 <= 0;
        i_8_668 <= 0;
        i_8_669 <= 0;
        i_8_670 <= 0;
        i_8_671 <= 0;
        i_8_672 <= 0;
        i_8_673 <= 0;
        i_8_674 <= 0;
        i_8_675 <= 0;
        i_8_676 <= 0;
        i_8_677 <= 0;
        i_8_678 <= 0;
        i_8_679 <= 0;
        i_8_680 <= 0;
        i_8_681 <= 0;
        i_8_682 <= 0;
        i_8_683 <= 0;
        i_8_684 <= 0;
        i_8_685 <= 0;
        i_8_686 <= 0;
        i_8_687 <= 0;
        i_8_688 <= 0;
        i_8_689 <= 0;
        i_8_690 <= 0;
        i_8_691 <= 0;
        i_8_692 <= 0;
        i_8_693 <= 0;
        i_8_694 <= 0;
        i_8_695 <= 0;
        i_8_696 <= 0;
        i_8_697 <= 0;
        i_8_698 <= 0;
        i_8_699 <= 0;
        i_8_700 <= 0;
        i_8_701 <= 0;
        i_8_702 <= 0;
        i_8_703 <= 0;
        i_8_704 <= 0;
        i_8_705 <= 0;
        i_8_706 <= 0;
        i_8_707 <= 0;
        i_8_708 <= 0;
        i_8_709 <= 0;
        i_8_710 <= 0;
        i_8_711 <= 0;
        i_8_712 <= 0;
        i_8_713 <= 0;
        i_8_714 <= 0;
        i_8_715 <= 0;
        i_8_716 <= 0;
        i_8_717 <= 0;
        i_8_718 <= 0;
        i_8_719 <= 0;
        i_8_720 <= 0;
        i_8_721 <= 0;
        i_8_722 <= 0;
        i_8_723 <= 0;
        i_8_724 <= 0;
        i_8_725 <= 0;
        i_8_726 <= 0;
        i_8_727 <= 0;
        i_8_728 <= 0;
        i_8_729 <= 0;
        i_8_730 <= 0;
        i_8_731 <= 0;
        i_8_732 <= 0;
        i_8_733 <= 0;
        i_8_734 <= 0;
        i_8_735 <= 0;
        i_8_736 <= 0;
        i_8_737 <= 0;
        i_8_738 <= 0;
        i_8_739 <= 0;
        i_8_740 <= 0;
        i_8_741 <= 0;
        i_8_742 <= 0;
        i_8_743 <= 0;
        i_8_744 <= 0;
        i_8_745 <= 0;
        i_8_746 <= 0;
        i_8_747 <= 0;
        i_8_748 <= 0;
        i_8_749 <= 0;
        i_8_750 <= 0;
        i_8_751 <= 0;
        i_8_752 <= 0;
        i_8_753 <= 0;
        i_8_754 <= 0;
        i_8_755 <= 0;
        i_8_756 <= 0;
        i_8_757 <= 0;
        i_8_758 <= 0;
        i_8_759 <= 0;
        i_8_760 <= 0;
        i_8_761 <= 0;
        i_8_762 <= 0;
        i_8_763 <= 0;
        i_8_764 <= 0;
        i_8_765 <= 0;
        i_8_766 <= 0;
        i_8_767 <= 0;
        i_8_768 <= 0;
        i_8_769 <= 0;
        i_8_770 <= 0;
        i_8_771 <= 0;
        i_8_772 <= 0;
        i_8_773 <= 0;
        i_8_774 <= 0;
        i_8_775 <= 0;
        i_8_776 <= 0;
        i_8_777 <= 0;
        i_8_778 <= 0;
        i_8_779 <= 0;
        i_8_780 <= 0;
        i_8_781 <= 0;
        i_8_782 <= 0;
        i_8_783 <= 0;
        i_8_784 <= 0;
        i_8_785 <= 0;
        i_8_786 <= 0;
        i_8_787 <= 0;
        i_8_788 <= 0;
        i_8_789 <= 0;
        i_8_790 <= 0;
        i_8_791 <= 0;
        i_8_792 <= 0;
        i_8_793 <= 0;
        i_8_794 <= 0;
        i_8_795 <= 0;
        i_8_796 <= 0;
        i_8_797 <= 0;
        i_8_798 <= 0;
        i_8_799 <= 0;
        i_8_800 <= 0;
        i_8_801 <= 0;
        i_8_802 <= 0;
        i_8_803 <= 0;
        i_8_804 <= 0;
        i_8_805 <= 0;
        i_8_806 <= 0;
        i_8_807 <= 0;
        i_8_808 <= 0;
        i_8_809 <= 0;
        i_8_810 <= 0;
        i_8_811 <= 0;
        i_8_812 <= 0;
        i_8_813 <= 0;
        i_8_814 <= 0;
        i_8_815 <= 0;
        i_8_816 <= 0;
        i_8_817 <= 0;
        i_8_818 <= 0;
        i_8_819 <= 0;
        i_8_820 <= 0;
        i_8_821 <= 0;
        i_8_822 <= 0;
        i_8_823 <= 0;
        i_8_824 <= 0;
        i_8_825 <= 0;
        i_8_826 <= 0;
        i_8_827 <= 0;
        i_8_828 <= 0;
        i_8_829 <= 0;
        i_8_830 <= 0;
        i_8_831 <= 0;
        i_8_832 <= 0;
        i_8_833 <= 0;
        i_8_834 <= 0;
        i_8_835 <= 0;
        i_8_836 <= 0;
        i_8_837 <= 0;
        i_8_838 <= 0;
        i_8_839 <= 0;
        i_8_840 <= 0;
        i_8_841 <= 0;
        i_8_842 <= 0;
        i_8_843 <= 0;
        i_8_844 <= 0;
        i_8_845 <= 0;
        i_8_846 <= 0;
        i_8_847 <= 0;
        i_8_848 <= 0;
        i_8_849 <= 0;
        i_8_850 <= 0;
        i_8_851 <= 0;
        i_8_852 <= 0;
        i_8_853 <= 0;
        i_8_854 <= 0;
        i_8_855 <= 0;
        i_8_856 <= 0;
        i_8_857 <= 0;
        i_8_858 <= 0;
        i_8_859 <= 0;
        i_8_860 <= 0;
        i_8_861 <= 0;
        i_8_862 <= 0;
        i_8_863 <= 0;
        i_8_864 <= 0;
        i_8_865 <= 0;
        i_8_866 <= 0;
        i_8_867 <= 0;
        i_8_868 <= 0;
        i_8_869 <= 0;
        i_8_870 <= 0;
        i_8_871 <= 0;
        i_8_872 <= 0;
        i_8_873 <= 0;
        i_8_874 <= 0;
        i_8_875 <= 0;
        i_8_876 <= 0;
        i_8_877 <= 0;
        i_8_878 <= 0;
        i_8_879 <= 0;
        i_8_880 <= 0;
        i_8_881 <= 0;
        i_8_882 <= 0;
        i_8_883 <= 0;
        i_8_884 <= 0;
        i_8_885 <= 0;
        i_8_886 <= 0;
        i_8_887 <= 0;
        i_8_888 <= 0;
        i_8_889 <= 0;
        i_8_890 <= 0;
        i_8_891 <= 0;
        i_8_892 <= 0;
        i_8_893 <= 0;
        i_8_894 <= 0;
        i_8_895 <= 0;
        i_8_896 <= 0;
        i_8_897 <= 0;
        i_8_898 <= 0;
        i_8_899 <= 0;
        i_8_900 <= 0;
        i_8_901 <= 0;
        i_8_902 <= 0;
        i_8_903 <= 0;
        i_8_904 <= 0;
        i_8_905 <= 0;
        i_8_906 <= 0;
        i_8_907 <= 0;
        i_8_908 <= 0;
        i_8_909 <= 0;
        i_8_910 <= 0;
        i_8_911 <= 0;
        i_8_912 <= 0;
        i_8_913 <= 0;
        i_8_914 <= 0;
        i_8_915 <= 0;
        i_8_916 <= 0;
        i_8_917 <= 0;
        i_8_918 <= 0;
        i_8_919 <= 0;
        i_8_920 <= 0;
        i_8_921 <= 0;
        i_8_922 <= 0;
        i_8_923 <= 0;
        i_8_924 <= 0;
        i_8_925 <= 0;
        i_8_926 <= 0;
        i_8_927 <= 0;
        i_8_928 <= 0;
        i_8_929 <= 0;
        i_8_930 <= 0;
        i_8_931 <= 0;
        i_8_932 <= 0;
        i_8_933 <= 0;
        i_8_934 <= 0;
        i_8_935 <= 0;
        i_8_936 <= 0;
        i_8_937 <= 0;
        i_8_938 <= 0;
        i_8_939 <= 0;
        i_8_940 <= 0;
        i_8_941 <= 0;
        i_8_942 <= 0;
        i_8_943 <= 0;
        i_8_944 <= 0;
        i_8_945 <= 0;
        i_8_946 <= 0;
        i_8_947 <= 0;
        i_8_948 <= 0;
        i_8_949 <= 0;
        i_8_950 <= 0;
        i_8_951 <= 0;
        i_8_952 <= 0;
        i_8_953 <= 0;
        i_8_954 <= 0;
        i_8_955 <= 0;
        i_8_956 <= 0;
        i_8_957 <= 0;
        i_8_958 <= 0;
        i_8_959 <= 0;
        i_8_960 <= 0;
        i_8_961 <= 0;
        i_8_962 <= 0;
        i_8_963 <= 0;
        i_8_964 <= 0;
        i_8_965 <= 0;
        i_8_966 <= 0;
        i_8_967 <= 0;
        i_8_968 <= 0;
        i_8_969 <= 0;
        i_8_970 <= 0;
        i_8_971 <= 0;
        i_8_972 <= 0;
        i_8_973 <= 0;
        i_8_974 <= 0;
        i_8_975 <= 0;
        i_8_976 <= 0;
        i_8_977 <= 0;
        i_8_978 <= 0;
        i_8_979 <= 0;
        i_8_980 <= 0;
        i_8_981 <= 0;
        i_8_982 <= 0;
        i_8_983 <= 0;
        i_8_984 <= 0;
        i_8_985 <= 0;
        i_8_986 <= 0;
        i_8_987 <= 0;
        i_8_988 <= 0;
        i_8_989 <= 0;
        i_8_990 <= 0;
        i_8_991 <= 0;
        i_8_992 <= 0;
        i_8_993 <= 0;
        i_8_994 <= 0;
        i_8_995 <= 0;
        i_8_996 <= 0;
        i_8_997 <= 0;
        i_8_998 <= 0;
        i_8_999 <= 0;
        i_8_1000 <= 0;
        i_8_1001 <= 0;
        i_8_1002 <= 0;
        i_8_1003 <= 0;
        i_8_1004 <= 0;
        i_8_1005 <= 0;
        i_8_1006 <= 0;
        i_8_1007 <= 0;
        i_8_1008 <= 0;
        i_8_1009 <= 0;
        i_8_1010 <= 0;
        i_8_1011 <= 0;
        i_8_1012 <= 0;
        i_8_1013 <= 0;
        i_8_1014 <= 0;
        i_8_1015 <= 0;
        i_8_1016 <= 0;
        i_8_1017 <= 0;
        i_8_1018 <= 0;
        i_8_1019 <= 0;
        i_8_1020 <= 0;
        i_8_1021 <= 0;
        i_8_1022 <= 0;
        i_8_1023 <= 0;
        i_8_1024 <= 0;
        i_8_1025 <= 0;
        i_8_1026 <= 0;
        i_8_1027 <= 0;
        i_8_1028 <= 0;
        i_8_1029 <= 0;
        i_8_1030 <= 0;
        i_8_1031 <= 0;
        i_8_1032 <= 0;
        i_8_1033 <= 0;
        i_8_1034 <= 0;
        i_8_1035 <= 0;
        i_8_1036 <= 0;
        i_8_1037 <= 0;
        i_8_1038 <= 0;
        i_8_1039 <= 0;
        i_8_1040 <= 0;
        i_8_1041 <= 0;
        i_8_1042 <= 0;
        i_8_1043 <= 0;
        i_8_1044 <= 0;
        i_8_1045 <= 0;
        i_8_1046 <= 0;
        i_8_1047 <= 0;
        i_8_1048 <= 0;
        i_8_1049 <= 0;
        i_8_1050 <= 0;
        i_8_1051 <= 0;
        i_8_1052 <= 0;
        i_8_1053 <= 0;
        i_8_1054 <= 0;
        i_8_1055 <= 0;
        i_8_1056 <= 0;
        i_8_1057 <= 0;
        i_8_1058 <= 0;
        i_8_1059 <= 0;
        i_8_1060 <= 0;
        i_8_1061 <= 0;
        i_8_1062 <= 0;
        i_8_1063 <= 0;
        i_8_1064 <= 0;
        i_8_1065 <= 0;
        i_8_1066 <= 0;
        i_8_1067 <= 0;
        i_8_1068 <= 0;
        i_8_1069 <= 0;
        i_8_1070 <= 0;
        i_8_1071 <= 0;
        i_8_1072 <= 0;
        i_8_1073 <= 0;
        i_8_1074 <= 0;
        i_8_1075 <= 0;
        i_8_1076 <= 0;
        i_8_1077 <= 0;
        i_8_1078 <= 0;
        i_8_1079 <= 0;
        i_8_1080 <= 0;
        i_8_1081 <= 0;
        i_8_1082 <= 0;
        i_8_1083 <= 0;
        i_8_1084 <= 0;
        i_8_1085 <= 0;
        i_8_1086 <= 0;
        i_8_1087 <= 0;
        i_8_1088 <= 0;
        i_8_1089 <= 0;
        i_8_1090 <= 0;
        i_8_1091 <= 0;
        i_8_1092 <= 0;
        i_8_1093 <= 0;
        i_8_1094 <= 0;
        i_8_1095 <= 0;
        i_8_1096 <= 0;
        i_8_1097 <= 0;
        i_8_1098 <= 0;
        i_8_1099 <= 0;
        i_8_1100 <= 0;
        i_8_1101 <= 0;
        i_8_1102 <= 0;
        i_8_1103 <= 0;
        i_8_1104 <= 0;
        i_8_1105 <= 0;
        i_8_1106 <= 0;
        i_8_1107 <= 0;
        i_8_1108 <= 0;
        i_8_1109 <= 0;
        i_8_1110 <= 0;
        i_8_1111 <= 0;
        i_8_1112 <= 0;
        i_8_1113 <= 0;
        i_8_1114 <= 0;
        i_8_1115 <= 0;
        i_8_1116 <= 0;
        i_8_1117 <= 0;
        i_8_1118 <= 0;
        i_8_1119 <= 0;
        i_8_1120 <= 0;
        i_8_1121 <= 0;
        i_8_1122 <= 0;
        i_8_1123 <= 0;
        i_8_1124 <= 0;
        i_8_1125 <= 0;
        i_8_1126 <= 0;
        i_8_1127 <= 0;
        i_8_1128 <= 0;
        i_8_1129 <= 0;
        i_8_1130 <= 0;
        i_8_1131 <= 0;
        i_8_1132 <= 0;
        i_8_1133 <= 0;
        i_8_1134 <= 0;
        i_8_1135 <= 0;
        i_8_1136 <= 0;
        i_8_1137 <= 0;
        i_8_1138 <= 0;
        i_8_1139 <= 0;
        i_8_1140 <= 0;
        i_8_1141 <= 0;
        i_8_1142 <= 0;
        i_8_1143 <= 0;
        i_8_1144 <= 0;
        i_8_1145 <= 0;
        i_8_1146 <= 0;
        i_8_1147 <= 0;
        i_8_1148 <= 0;
        i_8_1149 <= 0;
        i_8_1150 <= 0;
        i_8_1151 <= 0;
        i_8_1152 <= 0;
        i_8_1153 <= 0;
        i_8_1154 <= 0;
        i_8_1155 <= 0;
        i_8_1156 <= 0;
        i_8_1157 <= 0;
        i_8_1158 <= 0;
        i_8_1159 <= 0;
        i_8_1160 <= 0;
        i_8_1161 <= 0;
        i_8_1162 <= 0;
        i_8_1163 <= 0;
        i_8_1164 <= 0;
        i_8_1165 <= 0;
        i_8_1166 <= 0;
        i_8_1167 <= 0;
        i_8_1168 <= 0;
        i_8_1169 <= 0;
        i_8_1170 <= 0;
        i_8_1171 <= 0;
        i_8_1172 <= 0;
        i_8_1173 <= 0;
        i_8_1174 <= 0;
        i_8_1175 <= 0;
        i_8_1176 <= 0;
        i_8_1177 <= 0;
        i_8_1178 <= 0;
        i_8_1179 <= 0;
        i_8_1180 <= 0;
        i_8_1181 <= 0;
        i_8_1182 <= 0;
        i_8_1183 <= 0;
        i_8_1184 <= 0;
        i_8_1185 <= 0;
        i_8_1186 <= 0;
        i_8_1187 <= 0;
        i_8_1188 <= 0;
        i_8_1189 <= 0;
        i_8_1190 <= 0;
        i_8_1191 <= 0;
        i_8_1192 <= 0;
        i_8_1193 <= 0;
        i_8_1194 <= 0;
        i_8_1195 <= 0;
        i_8_1196 <= 0;
        i_8_1197 <= 0;
        i_8_1198 <= 0;
        i_8_1199 <= 0;
        i_8_1200 <= 0;
        i_8_1201 <= 0;
        i_8_1202 <= 0;
        i_8_1203 <= 0;
        i_8_1204 <= 0;
        i_8_1205 <= 0;
        i_8_1206 <= 0;
        i_8_1207 <= 0;
        i_8_1208 <= 0;
        i_8_1209 <= 0;
        i_8_1210 <= 0;
        i_8_1211 <= 0;
        i_8_1212 <= 0;
        i_8_1213 <= 0;
        i_8_1214 <= 0;
        i_8_1215 <= 0;
        i_8_1216 <= 0;
        i_8_1217 <= 0;
        i_8_1218 <= 0;
        i_8_1219 <= 0;
        i_8_1220 <= 0;
        i_8_1221 <= 0;
        i_8_1222 <= 0;
        i_8_1223 <= 0;
        i_8_1224 <= 0;
        i_8_1225 <= 0;
        i_8_1226 <= 0;
        i_8_1227 <= 0;
        i_8_1228 <= 0;
        i_8_1229 <= 0;
        i_8_1230 <= 0;
        i_8_1231 <= 0;
        i_8_1232 <= 0;
        i_8_1233 <= 0;
        i_8_1234 <= 0;
        i_8_1235 <= 0;
        i_8_1236 <= 0;
        i_8_1237 <= 0;
        i_8_1238 <= 0;
        i_8_1239 <= 0;
        i_8_1240 <= 0;
        i_8_1241 <= 0;
        i_8_1242 <= 0;
        i_8_1243 <= 0;
        i_8_1244 <= 0;
        i_8_1245 <= 0;
        i_8_1246 <= 0;
        i_8_1247 <= 0;
        i_8_1248 <= 0;
        i_8_1249 <= 0;
        i_8_1250 <= 0;
        i_8_1251 <= 0;
        i_8_1252 <= 0;
        i_8_1253 <= 0;
        i_8_1254 <= 0;
        i_8_1255 <= 0;
        i_8_1256 <= 0;
        i_8_1257 <= 0;
        i_8_1258 <= 0;
        i_8_1259 <= 0;
        i_8_1260 <= 0;
        i_8_1261 <= 0;
        i_8_1262 <= 0;
        i_8_1263 <= 0;
        i_8_1264 <= 0;
        i_8_1265 <= 0;
        i_8_1266 <= 0;
        i_8_1267 <= 0;
        i_8_1268 <= 0;
        i_8_1269 <= 0;
        i_8_1270 <= 0;
        i_8_1271 <= 0;
        i_8_1272 <= 0;
        i_8_1273 <= 0;
        i_8_1274 <= 0;
        i_8_1275 <= 0;
        i_8_1276 <= 0;
        i_8_1277 <= 0;
        i_8_1278 <= 0;
        i_8_1279 <= 0;
        i_8_1280 <= 0;
        i_8_1281 <= 0;
        i_8_1282 <= 0;
        i_8_1283 <= 0;
        i_8_1284 <= 0;
        i_8_1285 <= 0;
        i_8_1286 <= 0;
        i_8_1287 <= 0;
        i_8_1288 <= 0;
        i_8_1289 <= 0;
        i_8_1290 <= 0;
        i_8_1291 <= 0;
        i_8_1292 <= 0;
        i_8_1293 <= 0;
        i_8_1294 <= 0;
        i_8_1295 <= 0;
        i_8_1296 <= 0;
        i_8_1297 <= 0;
        i_8_1298 <= 0;
        i_8_1299 <= 0;
        i_8_1300 <= 0;
        i_8_1301 <= 0;
        i_8_1302 <= 0;
        i_8_1303 <= 0;
        i_8_1304 <= 0;
        i_8_1305 <= 0;
        i_8_1306 <= 0;
        i_8_1307 <= 0;
        i_8_1308 <= 0;
        i_8_1309 <= 0;
        i_8_1310 <= 0;
        i_8_1311 <= 0;
        i_8_1312 <= 0;
        i_8_1313 <= 0;
        i_8_1314 <= 0;
        i_8_1315 <= 0;
        i_8_1316 <= 0;
        i_8_1317 <= 0;
        i_8_1318 <= 0;
        i_8_1319 <= 0;
        i_8_1320 <= 0;
        i_8_1321 <= 0;
        i_8_1322 <= 0;
        i_8_1323 <= 0;
        i_8_1324 <= 0;
        i_8_1325 <= 0;
        i_8_1326 <= 0;
        i_8_1327 <= 0;
        i_8_1328 <= 0;
        i_8_1329 <= 0;
        i_8_1330 <= 0;
        i_8_1331 <= 0;
        i_8_1332 <= 0;
        i_8_1333 <= 0;
        i_8_1334 <= 0;
        i_8_1335 <= 0;
        i_8_1336 <= 0;
        i_8_1337 <= 0;
        i_8_1338 <= 0;
        i_8_1339 <= 0;
        i_8_1340 <= 0;
        i_8_1341 <= 0;
        i_8_1342 <= 0;
        i_8_1343 <= 0;
        i_8_1344 <= 0;
        i_8_1345 <= 0;
        i_8_1346 <= 0;
        i_8_1347 <= 0;
        i_8_1348 <= 0;
        i_8_1349 <= 0;
        i_8_1350 <= 0;
        i_8_1351 <= 0;
        i_8_1352 <= 0;
        i_8_1353 <= 0;
        i_8_1354 <= 0;
        i_8_1355 <= 0;
        i_8_1356 <= 0;
        i_8_1357 <= 0;
        i_8_1358 <= 0;
        i_8_1359 <= 0;
        i_8_1360 <= 0;
        i_8_1361 <= 0;
        i_8_1362 <= 0;
        i_8_1363 <= 0;
        i_8_1364 <= 0;
        i_8_1365 <= 0;
        i_8_1366 <= 0;
        i_8_1367 <= 0;
        i_8_1368 <= 0;
        i_8_1369 <= 0;
        i_8_1370 <= 0;
        i_8_1371 <= 0;
        i_8_1372 <= 0;
        i_8_1373 <= 0;
        i_8_1374 <= 0;
        i_8_1375 <= 0;
        i_8_1376 <= 0;
        i_8_1377 <= 0;
        i_8_1378 <= 0;
        i_8_1379 <= 0;
        i_8_1380 <= 0;
        i_8_1381 <= 0;
        i_8_1382 <= 0;
        i_8_1383 <= 0;
        i_8_1384 <= 0;
        i_8_1385 <= 0;
        i_8_1386 <= 0;
        i_8_1387 <= 0;
        i_8_1388 <= 0;
        i_8_1389 <= 0;
        i_8_1390 <= 0;
        i_8_1391 <= 0;
        i_8_1392 <= 0;
        i_8_1393 <= 0;
        i_8_1394 <= 0;
        i_8_1395 <= 0;
        i_8_1396 <= 0;
        i_8_1397 <= 0;
        i_8_1398 <= 0;
        i_8_1399 <= 0;
        i_8_1400 <= 0;
        i_8_1401 <= 0;
        i_8_1402 <= 0;
        i_8_1403 <= 0;
        i_8_1404 <= 0;
        i_8_1405 <= 0;
        i_8_1406 <= 0;
        i_8_1407 <= 0;
        i_8_1408 <= 0;
        i_8_1409 <= 0;
        i_8_1410 <= 0;
        i_8_1411 <= 0;
        i_8_1412 <= 0;
        i_8_1413 <= 0;
        i_8_1414 <= 0;
        i_8_1415 <= 0;
        i_8_1416 <= 0;
        i_8_1417 <= 0;
        i_8_1418 <= 0;
        i_8_1419 <= 0;
        i_8_1420 <= 0;
        i_8_1421 <= 0;
        i_8_1422 <= 0;
        i_8_1423 <= 0;
        i_8_1424 <= 0;
        i_8_1425 <= 0;
        i_8_1426 <= 0;
        i_8_1427 <= 0;
        i_8_1428 <= 0;
        i_8_1429 <= 0;
        i_8_1430 <= 0;
        i_8_1431 <= 0;
        i_8_1432 <= 0;
        i_8_1433 <= 0;
        i_8_1434 <= 0;
        i_8_1435 <= 0;
        i_8_1436 <= 0;
        i_8_1437 <= 0;
        i_8_1438 <= 0;
        i_8_1439 <= 0;
        i_8_1440 <= 0;
        i_8_1441 <= 0;
        i_8_1442 <= 0;
        i_8_1443 <= 0;
        i_8_1444 <= 0;
        i_8_1445 <= 0;
        i_8_1446 <= 0;
        i_8_1447 <= 0;
        i_8_1448 <= 0;
        i_8_1449 <= 0;
        i_8_1450 <= 0;
        i_8_1451 <= 0;
        i_8_1452 <= 0;
        i_8_1453 <= 0;
        i_8_1454 <= 0;
        i_8_1455 <= 0;
        i_8_1456 <= 0;
        i_8_1457 <= 0;
        i_8_1458 <= 0;
        i_8_1459 <= 0;
        i_8_1460 <= 0;
        i_8_1461 <= 0;
        i_8_1462 <= 0;
        i_8_1463 <= 0;
        i_8_1464 <= 0;
        i_8_1465 <= 0;
        i_8_1466 <= 0;
        i_8_1467 <= 0;
        i_8_1468 <= 0;
        i_8_1469 <= 0;
        i_8_1470 <= 0;
        i_8_1471 <= 0;
        i_8_1472 <= 0;
        i_8_1473 <= 0;
        i_8_1474 <= 0;
        i_8_1475 <= 0;
        i_8_1476 <= 0;
        i_8_1477 <= 0;
        i_8_1478 <= 0;
        i_8_1479 <= 0;
        i_8_1480 <= 0;
        i_8_1481 <= 0;
        i_8_1482 <= 0;
        i_8_1483 <= 0;
        i_8_1484 <= 0;
        i_8_1485 <= 0;
        i_8_1486 <= 0;
        i_8_1487 <= 0;
        i_8_1488 <= 0;
        i_8_1489 <= 0;
        i_8_1490 <= 0;
        i_8_1491 <= 0;
        i_8_1492 <= 0;
        i_8_1493 <= 0;
        i_8_1494 <= 0;
        i_8_1495 <= 0;
        i_8_1496 <= 0;
        i_8_1497 <= 0;
        i_8_1498 <= 0;
        i_8_1499 <= 0;
        i_8_1500 <= 0;
        i_8_1501 <= 0;
        i_8_1502 <= 0;
        i_8_1503 <= 0;
        i_8_1504 <= 0;
        i_8_1505 <= 0;
        i_8_1506 <= 0;
        i_8_1507 <= 0;
        i_8_1508 <= 0;
        i_8_1509 <= 0;
        i_8_1510 <= 0;
        i_8_1511 <= 0;
        i_8_1512 <= 0;
        i_8_1513 <= 0;
        i_8_1514 <= 0;
        i_8_1515 <= 0;
        i_8_1516 <= 0;
        i_8_1517 <= 0;
        i_8_1518 <= 0;
        i_8_1519 <= 0;
        i_8_1520 <= 0;
        i_8_1521 <= 0;
        i_8_1522 <= 0;
        i_8_1523 <= 0;
        i_8_1524 <= 0;
        i_8_1525 <= 0;
        i_8_1526 <= 0;
        i_8_1527 <= 0;
        i_8_1528 <= 0;
        i_8_1529 <= 0;
        i_8_1530 <= 0;
        i_8_1531 <= 0;
        i_8_1532 <= 0;
        i_8_1533 <= 0;
        i_8_1534 <= 0;
        i_8_1535 <= 0;
        i_8_1536 <= 0;
        i_8_1537 <= 0;
        i_8_1538 <= 0;
        i_8_1539 <= 0;
        i_8_1540 <= 0;
        i_8_1541 <= 0;
        i_8_1542 <= 0;
        i_8_1543 <= 0;
        i_8_1544 <= 0;
        i_8_1545 <= 0;
        i_8_1546 <= 0;
        i_8_1547 <= 0;
        i_8_1548 <= 0;
        i_8_1549 <= 0;
        i_8_1550 <= 0;
        i_8_1551 <= 0;
        i_8_1552 <= 0;
        i_8_1553 <= 0;
        i_8_1554 <= 0;
        i_8_1555 <= 0;
        i_8_1556 <= 0;
        i_8_1557 <= 0;
        i_8_1558 <= 0;
        i_8_1559 <= 0;
        i_8_1560 <= 0;
        i_8_1561 <= 0;
        i_8_1562 <= 0;
        i_8_1563 <= 0;
        i_8_1564 <= 0;
        i_8_1565 <= 0;
        i_8_1566 <= 0;
        i_8_1567 <= 0;
        i_8_1568 <= 0;
        i_8_1569 <= 0;
        i_8_1570 <= 0;
        i_8_1571 <= 0;
        i_8_1572 <= 0;
        i_8_1573 <= 0;
        i_8_1574 <= 0;
        i_8_1575 <= 0;
        i_8_1576 <= 0;
        i_8_1577 <= 0;
        i_8_1578 <= 0;
        i_8_1579 <= 0;
        i_8_1580 <= 0;
        i_8_1581 <= 0;
        i_8_1582 <= 0;
        i_8_1583 <= 0;
        i_8_1584 <= 0;
        i_8_1585 <= 0;
        i_8_1586 <= 0;
        i_8_1587 <= 0;
        i_8_1588 <= 0;
        i_8_1589 <= 0;
        i_8_1590 <= 0;
        i_8_1591 <= 0;
        i_8_1592 <= 0;
        i_8_1593 <= 0;
        i_8_1594 <= 0;
        i_8_1595 <= 0;
        i_8_1596 <= 0;
        i_8_1597 <= 0;
        i_8_1598 <= 0;
        i_8_1599 <= 0;
        i_8_1600 <= 0;
        i_8_1601 <= 0;
        i_8_1602 <= 0;
        i_8_1603 <= 0;
        i_8_1604 <= 0;
        i_8_1605 <= 0;
        i_8_1606 <= 0;
        i_8_1607 <= 0;
        i_8_1608 <= 0;
        i_8_1609 <= 0;
        i_8_1610 <= 0;
        i_8_1611 <= 0;
        i_8_1612 <= 0;
        i_8_1613 <= 0;
        i_8_1614 <= 0;
        i_8_1615 <= 0;
        i_8_1616 <= 0;
        i_8_1617 <= 0;
        i_8_1618 <= 0;
        i_8_1619 <= 0;
        i_8_1620 <= 0;
        i_8_1621 <= 0;
        i_8_1622 <= 0;
        i_8_1623 <= 0;
        i_8_1624 <= 0;
        i_8_1625 <= 0;
        i_8_1626 <= 0;
        i_8_1627 <= 0;
        i_8_1628 <= 0;
        i_8_1629 <= 0;
        i_8_1630 <= 0;
        i_8_1631 <= 0;
        i_8_1632 <= 0;
        i_8_1633 <= 0;
        i_8_1634 <= 0;
        i_8_1635 <= 0;
        i_8_1636 <= 0;
        i_8_1637 <= 0;
        i_8_1638 <= 0;
        i_8_1639 <= 0;
        i_8_1640 <= 0;
        i_8_1641 <= 0;
        i_8_1642 <= 0;
        i_8_1643 <= 0;
        i_8_1644 <= 0;
        i_8_1645 <= 0;
        i_8_1646 <= 0;
        i_8_1647 <= 0;
        i_8_1648 <= 0;
        i_8_1649 <= 0;
        i_8_1650 <= 0;
        i_8_1651 <= 0;
        i_8_1652 <= 0;
        i_8_1653 <= 0;
        i_8_1654 <= 0;
        i_8_1655 <= 0;
        i_8_1656 <= 0;
        i_8_1657 <= 0;
        i_8_1658 <= 0;
        i_8_1659 <= 0;
        i_8_1660 <= 0;
        i_8_1661 <= 0;
        i_8_1662 <= 0;
        i_8_1663 <= 0;
        i_8_1664 <= 0;
        i_8_1665 <= 0;
        i_8_1666 <= 0;
        i_8_1667 <= 0;
        i_8_1668 <= 0;
        i_8_1669 <= 0;
        i_8_1670 <= 0;
        i_8_1671 <= 0;
        i_8_1672 <= 0;
        i_8_1673 <= 0;
        i_8_1674 <= 0;
        i_8_1675 <= 0;
        i_8_1676 <= 0;
        i_8_1677 <= 0;
        i_8_1678 <= 0;
        i_8_1679 <= 0;
        i_8_1680 <= 0;
        i_8_1681 <= 0;
        i_8_1682 <= 0;
        i_8_1683 <= 0;
        i_8_1684 <= 0;
        i_8_1685 <= 0;
        i_8_1686 <= 0;
        i_8_1687 <= 0;
        i_8_1688 <= 0;
        i_8_1689 <= 0;
        i_8_1690 <= 0;
        i_8_1691 <= 0;
        i_8_1692 <= 0;
        i_8_1693 <= 0;
        i_8_1694 <= 0;
        i_8_1695 <= 0;
        i_8_1696 <= 0;
        i_8_1697 <= 0;
        i_8_1698 <= 0;
        i_8_1699 <= 0;
        i_8_1700 <= 0;
        i_8_1701 <= 0;
        i_8_1702 <= 0;
        i_8_1703 <= 0;
        i_8_1704 <= 0;
        i_8_1705 <= 0;
        i_8_1706 <= 0;
        i_8_1707 <= 0;
        i_8_1708 <= 0;
        i_8_1709 <= 0;
        i_8_1710 <= 0;
        i_8_1711 <= 0;
        i_8_1712 <= 0;
        i_8_1713 <= 0;
        i_8_1714 <= 0;
        i_8_1715 <= 0;
        i_8_1716 <= 0;
        i_8_1717 <= 0;
        i_8_1718 <= 0;
        i_8_1719 <= 0;
        i_8_1720 <= 0;
        i_8_1721 <= 0;
        i_8_1722 <= 0;
        i_8_1723 <= 0;
        i_8_1724 <= 0;
        i_8_1725 <= 0;
        i_8_1726 <= 0;
        i_8_1727 <= 0;
        i_8_1728 <= 0;
        i_8_1729 <= 0;
        i_8_1730 <= 0;
        i_8_1731 <= 0;
        i_8_1732 <= 0;
        i_8_1733 <= 0;
        i_8_1734 <= 0;
        i_8_1735 <= 0;
        i_8_1736 <= 0;
        i_8_1737 <= 0;
        i_8_1738 <= 0;
        i_8_1739 <= 0;
        i_8_1740 <= 0;
        i_8_1741 <= 0;
        i_8_1742 <= 0;
        i_8_1743 <= 0;
        i_8_1744 <= 0;
        i_8_1745 <= 0;
        i_8_1746 <= 0;
        i_8_1747 <= 0;
        i_8_1748 <= 0;
        i_8_1749 <= 0;
        i_8_1750 <= 0;
        i_8_1751 <= 0;
        i_8_1752 <= 0;
        i_8_1753 <= 0;
        i_8_1754 <= 0;
        i_8_1755 <= 0;
        i_8_1756 <= 0;
        i_8_1757 <= 0;
        i_8_1758 <= 0;
        i_8_1759 <= 0;
        i_8_1760 <= 0;
        i_8_1761 <= 0;
        i_8_1762 <= 0;
        i_8_1763 <= 0;
        i_8_1764 <= 0;
        i_8_1765 <= 0;
        i_8_1766 <= 0;
        i_8_1767 <= 0;
        i_8_1768 <= 0;
        i_8_1769 <= 0;
        i_8_1770 <= 0;
        i_8_1771 <= 0;
        i_8_1772 <= 0;
        i_8_1773 <= 0;
        i_8_1774 <= 0;
        i_8_1775 <= 0;
        i_8_1776 <= 0;
        i_8_1777 <= 0;
        i_8_1778 <= 0;
        i_8_1779 <= 0;
        i_8_1780 <= 0;
        i_8_1781 <= 0;
        i_8_1782 <= 0;
        i_8_1783 <= 0;
        i_8_1784 <= 0;
        i_8_1785 <= 0;
        i_8_1786 <= 0;
        i_8_1787 <= 0;
        i_8_1788 <= 0;
        i_8_1789 <= 0;
        i_8_1790 <= 0;
        i_8_1791 <= 0;
        i_8_1792 <= 0;
        i_8_1793 <= 0;
        i_8_1794 <= 0;
        i_8_1795 <= 0;
        i_8_1796 <= 0;
        i_8_1797 <= 0;
        i_8_1798 <= 0;
        i_8_1799 <= 0;
        i_8_1800 <= 0;
        i_8_1801 <= 0;
        i_8_1802 <= 0;
        i_8_1803 <= 0;
        i_8_1804 <= 0;
        i_8_1805 <= 0;
        i_8_1806 <= 0;
        i_8_1807 <= 0;
        i_8_1808 <= 0;
        i_8_1809 <= 0;
        i_8_1810 <= 0;
        i_8_1811 <= 0;
        i_8_1812 <= 0;
        i_8_1813 <= 0;
        i_8_1814 <= 0;
        i_8_1815 <= 0;
        i_8_1816 <= 0;
        i_8_1817 <= 0;
        i_8_1818 <= 0;
        i_8_1819 <= 0;
        i_8_1820 <= 0;
        i_8_1821 <= 0;
        i_8_1822 <= 0;
        i_8_1823 <= 0;
        i_8_1824 <= 0;
        i_8_1825 <= 0;
        i_8_1826 <= 0;
        i_8_1827 <= 0;
        i_8_1828 <= 0;
        i_8_1829 <= 0;
        i_8_1830 <= 0;
        i_8_1831 <= 0;
        i_8_1832 <= 0;
        i_8_1833 <= 0;
        i_8_1834 <= 0;
        i_8_1835 <= 0;
        i_8_1836 <= 0;
        i_8_1837 <= 0;
        i_8_1838 <= 0;
        i_8_1839 <= 0;
        i_8_1840 <= 0;
        i_8_1841 <= 0;
        i_8_1842 <= 0;
        i_8_1843 <= 0;
        i_8_1844 <= 0;
        i_8_1845 <= 0;
        i_8_1846 <= 0;
        i_8_1847 <= 0;
        i_8_1848 <= 0;
        i_8_1849 <= 0;
        i_8_1850 <= 0;
        i_8_1851 <= 0;
        i_8_1852 <= 0;
        i_8_1853 <= 0;
        i_8_1854 <= 0;
        i_8_1855 <= 0;
        i_8_1856 <= 0;
        i_8_1857 <= 0;
        i_8_1858 <= 0;
        i_8_1859 <= 0;
        i_8_1860 <= 0;
        i_8_1861 <= 0;
        i_8_1862 <= 0;
        i_8_1863 <= 0;
        i_8_1864 <= 0;
        i_8_1865 <= 0;
        i_8_1866 <= 0;
        i_8_1867 <= 0;
        i_8_1868 <= 0;
        i_8_1869 <= 0;
        i_8_1870 <= 0;
        i_8_1871 <= 0;
        i_8_1872 <= 0;
        i_8_1873 <= 0;
        i_8_1874 <= 0;
        i_8_1875 <= 0;
        i_8_1876 <= 0;
        i_8_1877 <= 0;
        i_8_1878 <= 0;
        i_8_1879 <= 0;
        i_8_1880 <= 0;
        i_8_1881 <= 0;
        i_8_1882 <= 0;
        i_8_1883 <= 0;
        i_8_1884 <= 0;
        i_8_1885 <= 0;
        i_8_1886 <= 0;
        i_8_1887 <= 0;
        i_8_1888 <= 0;
        i_8_1889 <= 0;
        i_8_1890 <= 0;
        i_8_1891 <= 0;
        i_8_1892 <= 0;
        i_8_1893 <= 0;
        i_8_1894 <= 0;
        i_8_1895 <= 0;
        i_8_1896 <= 0;
        i_8_1897 <= 0;
        i_8_1898 <= 0;
        i_8_1899 <= 0;
        i_8_1900 <= 0;
        i_8_1901 <= 0;
        i_8_1902 <= 0;
        i_8_1903 <= 0;
        i_8_1904 <= 0;
        i_8_1905 <= 0;
        i_8_1906 <= 0;
        i_8_1907 <= 0;
        i_8_1908 <= 0;
        i_8_1909 <= 0;
        i_8_1910 <= 0;
        i_8_1911 <= 0;
        i_8_1912 <= 0;
        i_8_1913 <= 0;
        i_8_1914 <= 0;
        i_8_1915 <= 0;
        i_8_1916 <= 0;
        i_8_1917 <= 0;
        i_8_1918 <= 0;
        i_8_1919 <= 0;
        i_8_1920 <= 0;
        i_8_1921 <= 0;
        i_8_1922 <= 0;
        i_8_1923 <= 0;
        i_8_1924 <= 0;
        i_8_1925 <= 0;
        i_8_1926 <= 0;
        i_8_1927 <= 0;
        i_8_1928 <= 0;
        i_8_1929 <= 0;
        i_8_1930 <= 0;
        i_8_1931 <= 0;
        i_8_1932 <= 0;
        i_8_1933 <= 0;
        i_8_1934 <= 0;
        i_8_1935 <= 0;
        i_8_1936 <= 0;
        i_8_1937 <= 0;
        i_8_1938 <= 0;
        i_8_1939 <= 0;
        i_8_1940 <= 0;
        i_8_1941 <= 0;
        i_8_1942 <= 0;
        i_8_1943 <= 0;
        i_8_1944 <= 0;
        i_8_1945 <= 0;
        i_8_1946 <= 0;
        i_8_1947 <= 0;
        i_8_1948 <= 0;
        i_8_1949 <= 0;
        i_8_1950 <= 0;
        i_8_1951 <= 0;
        i_8_1952 <= 0;
        i_8_1953 <= 0;
        i_8_1954 <= 0;
        i_8_1955 <= 0;
        i_8_1956 <= 0;
        i_8_1957 <= 0;
        i_8_1958 <= 0;
        i_8_1959 <= 0;
        i_8_1960 <= 0;
        i_8_1961 <= 0;
        i_8_1962 <= 0;
        i_8_1963 <= 0;
        i_8_1964 <= 0;
        i_8_1965 <= 0;
        i_8_1966 <= 0;
        i_8_1967 <= 0;
        i_8_1968 <= 0;
        i_8_1969 <= 0;
        i_8_1970 <= 0;
        i_8_1971 <= 0;
        i_8_1972 <= 0;
        i_8_1973 <= 0;
        i_8_1974 <= 0;
        i_8_1975 <= 0;
        i_8_1976 <= 0;
        i_8_1977 <= 0;
        i_8_1978 <= 0;
        i_8_1979 <= 0;
        i_8_1980 <= 0;
        i_8_1981 <= 0;
        i_8_1982 <= 0;
        i_8_1983 <= 0;
        i_8_1984 <= 0;
        i_8_1985 <= 0;
        i_8_1986 <= 0;
        i_8_1987 <= 0;
        i_8_1988 <= 0;
        i_8_1989 <= 0;
        i_8_1990 <= 0;
        i_8_1991 <= 0;
        i_8_1992 <= 0;
        i_8_1993 <= 0;
        i_8_1994 <= 0;
        i_8_1995 <= 0;
        i_8_1996 <= 0;
        i_8_1997 <= 0;
        i_8_1998 <= 0;
        i_8_1999 <= 0;
        i_8_2000 <= 0;
        i_8_2001 <= 0;
        i_8_2002 <= 0;
        i_8_2003 <= 0;
        i_8_2004 <= 0;
        i_8_2005 <= 0;
        i_8_2006 <= 0;
        i_8_2007 <= 0;
        i_8_2008 <= 0;
        i_8_2009 <= 0;
        i_8_2010 <= 0;
        i_8_2011 <= 0;
        i_8_2012 <= 0;
        i_8_2013 <= 0;
        i_8_2014 <= 0;
        i_8_2015 <= 0;
        i_8_2016 <= 0;
        i_8_2017 <= 0;
        i_8_2018 <= 0;
        i_8_2019 <= 0;
        i_8_2020 <= 0;
        i_8_2021 <= 0;
        i_8_2022 <= 0;
        i_8_2023 <= 0;
        i_8_2024 <= 0;
        i_8_2025 <= 0;
        i_8_2026 <= 0;
        i_8_2027 <= 0;
        i_8_2028 <= 0;
        i_8_2029 <= 0;
        i_8_2030 <= 0;
        i_8_2031 <= 0;
        i_8_2032 <= 0;
        i_8_2033 <= 0;
        i_8_2034 <= 0;
        i_8_2035 <= 0;
        i_8_2036 <= 0;
        i_8_2037 <= 0;
        i_8_2038 <= 0;
        i_8_2039 <= 0;
        i_8_2040 <= 0;
        i_8_2041 <= 0;
        i_8_2042 <= 0;
        i_8_2043 <= 0;
        i_8_2044 <= 0;
        i_8_2045 <= 0;
        i_8_2046 <= 0;
        i_8_2047 <= 0;
        i_8_2048 <= 0;
        i_8_2049 <= 0;
        i_8_2050 <= 0;
        i_8_2051 <= 0;
        i_8_2052 <= 0;
        i_8_2053 <= 0;
        i_8_2054 <= 0;
        i_8_2055 <= 0;
        i_8_2056 <= 0;
        i_8_2057 <= 0;
        i_8_2058 <= 0;
        i_8_2059 <= 0;
        i_8_2060 <= 0;
        i_8_2061 <= 0;
        i_8_2062 <= 0;
        i_8_2063 <= 0;
        i_8_2064 <= 0;
        i_8_2065 <= 0;
        i_8_2066 <= 0;
        i_8_2067 <= 0;
        i_8_2068 <= 0;
        i_8_2069 <= 0;
        i_8_2070 <= 0;
        i_8_2071 <= 0;
        i_8_2072 <= 0;
        i_8_2073 <= 0;
        i_8_2074 <= 0;
        i_8_2075 <= 0;
        i_8_2076 <= 0;
        i_8_2077 <= 0;
        i_8_2078 <= 0;
        i_8_2079 <= 0;
        i_8_2080 <= 0;
        i_8_2081 <= 0;
        i_8_2082 <= 0;
        i_8_2083 <= 0;
        i_8_2084 <= 0;
        i_8_2085 <= 0;
        i_8_2086 <= 0;
        i_8_2087 <= 0;
        i_8_2088 <= 0;
        i_8_2089 <= 0;
        i_8_2090 <= 0;
        i_8_2091 <= 0;
        i_8_2092 <= 0;
        i_8_2093 <= 0;
        i_8_2094 <= 0;
        i_8_2095 <= 0;
        i_8_2096 <= 0;
        i_8_2097 <= 0;
        i_8_2098 <= 0;
        i_8_2099 <= 0;
        i_8_2100 <= 0;
        i_8_2101 <= 0;
        i_8_2102 <= 0;
        i_8_2103 <= 0;
        i_8_2104 <= 0;
        i_8_2105 <= 0;
        i_8_2106 <= 0;
        i_8_2107 <= 0;
        i_8_2108 <= 0;
        i_8_2109 <= 0;
        i_8_2110 <= 0;
        i_8_2111 <= 0;
        i_8_2112 <= 0;
        i_8_2113 <= 0;
        i_8_2114 <= 0;
        i_8_2115 <= 0;
        i_8_2116 <= 0;
        i_8_2117 <= 0;
        i_8_2118 <= 0;
        i_8_2119 <= 0;
        i_8_2120 <= 0;
        i_8_2121 <= 0;
        i_8_2122 <= 0;
        i_8_2123 <= 0;
        i_8_2124 <= 0;
        i_8_2125 <= 0;
        i_8_2126 <= 0;
        i_8_2127 <= 0;
        i_8_2128 <= 0;
        i_8_2129 <= 0;
        i_8_2130 <= 0;
        i_8_2131 <= 0;
        i_8_2132 <= 0;
        i_8_2133 <= 0;
        i_8_2134 <= 0;
        i_8_2135 <= 0;
        i_8_2136 <= 0;
        i_8_2137 <= 0;
        i_8_2138 <= 0;
        i_8_2139 <= 0;
        i_8_2140 <= 0;
        i_8_2141 <= 0;
        i_8_2142 <= 0;
        i_8_2143 <= 0;
        i_8_2144 <= 0;
        i_8_2145 <= 0;
        i_8_2146 <= 0;
        i_8_2147 <= 0;
        i_8_2148 <= 0;
        i_8_2149 <= 0;
        i_8_2150 <= 0;
        i_8_2151 <= 0;
        i_8_2152 <= 0;
        i_8_2153 <= 0;
        i_8_2154 <= 0;
        i_8_2155 <= 0;
        i_8_2156 <= 0;
        i_8_2157 <= 0;
        i_8_2158 <= 0;
        i_8_2159 <= 0;
        i_8_2160 <= 0;
        i_8_2161 <= 0;
        i_8_2162 <= 0;
        i_8_2163 <= 0;
        i_8_2164 <= 0;
        i_8_2165 <= 0;
        i_8_2166 <= 0;
        i_8_2167 <= 0;
        i_8_2168 <= 0;
        i_8_2169 <= 0;
        i_8_2170 <= 0;
        i_8_2171 <= 0;
        i_8_2172 <= 0;
        i_8_2173 <= 0;
        i_8_2174 <= 0;
        i_8_2175 <= 0;
        i_8_2176 <= 0;
        i_8_2177 <= 0;
        i_8_2178 <= 0;
        i_8_2179 <= 0;
        i_8_2180 <= 0;
        i_8_2181 <= 0;
        i_8_2182 <= 0;
        i_8_2183 <= 0;
        i_8_2184 <= 0;
        i_8_2185 <= 0;
        i_8_2186 <= 0;
        i_8_2187 <= 0;
        i_8_2188 <= 0;
        i_8_2189 <= 0;
        i_8_2190 <= 0;
        i_8_2191 <= 0;
        i_8_2192 <= 0;
        i_8_2193 <= 0;
        i_8_2194 <= 0;
        i_8_2195 <= 0;
        i_8_2196 <= 0;
        i_8_2197 <= 0;
        i_8_2198 <= 0;
        i_8_2199 <= 0;
        i_8_2200 <= 0;
        i_8_2201 <= 0;
        i_8_2202 <= 0;
        i_8_2203 <= 0;
        i_8_2204 <= 0;
        i_8_2205 <= 0;
        i_8_2206 <= 0;
        i_8_2207 <= 0;
        i_8_2208 <= 0;
        i_8_2209 <= 0;
        i_8_2210 <= 0;
        i_8_2211 <= 0;
        i_8_2212 <= 0;
        i_8_2213 <= 0;
        i_8_2214 <= 0;
        i_8_2215 <= 0;
        i_8_2216 <= 0;
        i_8_2217 <= 0;
        i_8_2218 <= 0;
        i_8_2219 <= 0;
        i_8_2220 <= 0;
        i_8_2221 <= 0;
        i_8_2222 <= 0;
        i_8_2223 <= 0;
        i_8_2224 <= 0;
        i_8_2225 <= 0;
        i_8_2226 <= 0;
        i_8_2227 <= 0;
        i_8_2228 <= 0;
        i_8_2229 <= 0;
        i_8_2230 <= 0;
        i_8_2231 <= 0;
        i_8_2232 <= 0;
        i_8_2233 <= 0;
        i_8_2234 <= 0;
        i_8_2235 <= 0;
        i_8_2236 <= 0;
        i_8_2237 <= 0;
        i_8_2238 <= 0;
        i_8_2239 <= 0;
        i_8_2240 <= 0;
        i_8_2241 <= 0;
        i_8_2242 <= 0;
        i_8_2243 <= 0;
        i_8_2244 <= 0;
        i_8_2245 <= 0;
        i_8_2246 <= 0;
        i_8_2247 <= 0;
        i_8_2248 <= 0;
        i_8_2249 <= 0;
        i_8_2250 <= 0;
        i_8_2251 <= 0;
        i_8_2252 <= 0;
        i_8_2253 <= 0;
        i_8_2254 <= 0;
        i_8_2255 <= 0;
        i_8_2256 <= 0;
        i_8_2257 <= 0;
        i_8_2258 <= 0;
        i_8_2259 <= 0;
        i_8_2260 <= 0;
        i_8_2261 <= 0;
        i_8_2262 <= 0;
        i_8_2263 <= 0;
        i_8_2264 <= 0;
        i_8_2265 <= 0;
        i_8_2266 <= 0;
        i_8_2267 <= 0;
        i_8_2268 <= 0;
        i_8_2269 <= 0;
        i_8_2270 <= 0;
        i_8_2271 <= 0;
        i_8_2272 <= 0;
        i_8_2273 <= 0;
        i_8_2274 <= 0;
        i_8_2275 <= 0;
        i_8_2276 <= 0;
        i_8_2277 <= 0;
        i_8_2278 <= 0;
        i_8_2279 <= 0;
        i_8_2280 <= 0;
        i_8_2281 <= 0;
        i_8_2282 <= 0;
        i_8_2283 <= 0;
        i_8_2284 <= 0;
        i_8_2285 <= 0;
        i_8_2286 <= 0;
        i_8_2287 <= 0;
        i_8_2288 <= 0;
        i_8_2289 <= 0;
        i_8_2290 <= 0;
        i_8_2291 <= 0;
        i_8_2292 <= 0;
        i_8_2293 <= 0;
        i_8_2294 <= 0;
        i_8_2295 <= 0;
        i_8_2296 <= 0;
        i_8_2297 <= 0;
        i_8_2298 <= 0;
        i_8_2299 <= 0;
        i_8_2300 <= 0;
        i_8_2301 <= 0;
        i_8_2302 <= 0;
        i_8_2303 <= 0;
        dly1 <= 0;
        dly2 <= 0;
      end
    else if (ce)
      begin
        out_reg <= { o_8_511, o_8_510, o_8_509, o_8_508, o_8_507, o_8_506, o_8_505, o_8_504, o_8_503, o_8_502, o_8_501, o_8_500, o_8_499, o_8_498, o_8_497, o_8_496, o_8_495, o_8_494, o_8_493, o_8_492, o_8_491, o_8_490, o_8_489, o_8_488, o_8_487, o_8_486, o_8_485, o_8_484, o_8_483, o_8_482, o_8_481, o_8_480, o_8_479, o_8_478, o_8_477, o_8_476, o_8_475, o_8_474, o_8_473, o_8_472, o_8_471, o_8_470, o_8_469, o_8_468, o_8_467, o_8_466, o_8_465, o_8_464, o_8_463, o_8_462, o_8_461, o_8_460, o_8_459, o_8_458, o_8_457, o_8_456, o_8_455, o_8_454, o_8_453, o_8_452, o_8_451, o_8_450, o_8_449, o_8_448, o_8_447, o_8_446, o_8_445, o_8_444, o_8_443, o_8_442, o_8_441, o_8_440, o_8_439, o_8_438, o_8_437, o_8_436, o_8_435, o_8_434, o_8_433, o_8_432, o_8_431, o_8_430, o_8_429, o_8_428, o_8_427, o_8_426, o_8_425, o_8_424, o_8_423, o_8_422, o_8_421, o_8_420, o_8_419, o_8_418, o_8_417, o_8_416, o_8_415, o_8_414, o_8_413, o_8_412, o_8_411, o_8_410, o_8_409, o_8_408, o_8_407, o_8_406, o_8_405, o_8_404, o_8_403, o_8_402, o_8_401, o_8_400, o_8_399, o_8_398, o_8_397, o_8_396, o_8_395, o_8_394, o_8_393, o_8_392, o_8_391, o_8_390, o_8_389, o_8_388, o_8_387, o_8_386, o_8_385, o_8_384, o_8_383, o_8_382, o_8_381, o_8_380, o_8_379, o_8_378, o_8_377, o_8_376, o_8_375, o_8_374, o_8_373, o_8_372, o_8_371, o_8_370, o_8_369, o_8_368, o_8_367, o_8_366, o_8_365, o_8_364, o_8_363, o_8_362, o_8_361, o_8_360, o_8_359, o_8_358, o_8_357, o_8_356, o_8_355, o_8_354, o_8_353, o_8_352, o_8_351, o_8_350, o_8_349, o_8_348, o_8_347, o_8_346, o_8_345, o_8_344, o_8_343, o_8_342, o_8_341, o_8_340, o_8_339, o_8_338, o_8_337, o_8_336, o_8_335, o_8_334, o_8_333, o_8_332, o_8_331, o_8_330, o_8_329, o_8_328, o_8_327, o_8_326, o_8_325, o_8_324, o_8_323, o_8_322, o_8_321, o_8_320, o_8_319, o_8_318, o_8_317, o_8_316, o_8_315, o_8_314, o_8_313, o_8_312, o_8_311, o_8_310, o_8_309, o_8_308, o_8_307, o_8_306, o_8_305, o_8_304, o_8_303, o_8_302, o_8_301, o_8_300, o_8_299, o_8_298, o_8_297, o_8_296, o_8_295, o_8_294, o_8_293, o_8_292, o_8_291, o_8_290, o_8_289, o_8_288, o_8_287, o_8_286, o_8_285, o_8_284, o_8_283, o_8_282, o_8_281, o_8_280, o_8_279, o_8_278, o_8_277, o_8_276, o_8_275, o_8_274, o_8_273, o_8_272, o_8_271, o_8_270, o_8_269, o_8_268, o_8_267, o_8_266, o_8_265, o_8_264, o_8_263, o_8_262, o_8_261, o_8_260, o_8_259, o_8_258, o_8_257, o_8_256, o_8_255, o_8_254, o_8_253, o_8_252, o_8_251, o_8_250, o_8_249, o_8_248, o_8_247, o_8_246, o_8_245, o_8_244, o_8_243, o_8_242, o_8_241, o_8_240, o_8_239, o_8_238, o_8_237, o_8_236, o_8_235, o_8_234, o_8_233, o_8_232, o_8_231, o_8_230, o_8_229, o_8_228, o_8_227, o_8_226, o_8_225, o_8_224, o_8_223, o_8_222, o_8_221, o_8_220, o_8_219, o_8_218, o_8_217, o_8_216, o_8_215, o_8_214, o_8_213, o_8_212, o_8_211, o_8_210, o_8_209, o_8_208, o_8_207, o_8_206, o_8_205, o_8_204, o_8_203, o_8_202, o_8_201, o_8_200, o_8_199, o_8_198, o_8_197, o_8_196, o_8_195, o_8_194, o_8_193, o_8_192, o_8_191, o_8_190, o_8_189, o_8_188, o_8_187, o_8_186, o_8_185, o_8_184, o_8_183, o_8_182, o_8_181, o_8_180, o_8_179, o_8_178, o_8_177, o_8_176, o_8_175, o_8_174, o_8_173, o_8_172, o_8_171, o_8_170, o_8_169, o_8_168, o_8_167, o_8_166, o_8_165, o_8_164, o_8_163, o_8_162, o_8_161, o_8_160, o_8_159, o_8_158, o_8_157, o_8_156, o_8_155, o_8_154, o_8_153, o_8_152, o_8_151, o_8_150, o_8_149, o_8_148, o_8_147, o_8_146, o_8_145, o_8_144, o_8_143, o_8_142, o_8_141, o_8_140, o_8_139, o_8_138, o_8_137, o_8_136, o_8_135, o_8_134, o_8_133, o_8_132, o_8_131, o_8_130, o_8_129, o_8_128, o_8_127, o_8_126, o_8_125, o_8_124, o_8_123, o_8_122, o_8_121, o_8_120, o_8_119, o_8_118, o_8_117, o_8_116, o_8_115, o_8_114, o_8_113, o_8_112, o_8_111, o_8_110, o_8_109, o_8_108, o_8_107, o_8_106, o_8_105, o_8_104, o_8_103, o_8_102, o_8_101, o_8_100, o_8_99, o_8_98, o_8_97, o_8_96, o_8_95, o_8_94, o_8_93, o_8_92, o_8_91, o_8_90, o_8_89, o_8_88, o_8_87, o_8_86, o_8_85, o_8_84, o_8_83, o_8_82, o_8_81, o_8_80, o_8_79, o_8_78, o_8_77, o_8_76, o_8_75, o_8_74, o_8_73, o_8_72, o_8_71, o_8_70, o_8_69, o_8_68, o_8_67, o_8_66, o_8_65, o_8_64, o_8_63, o_8_62, o_8_61, o_8_60, o_8_59, o_8_58, o_8_57, o_8_56, o_8_55, o_8_54, o_8_53, o_8_52, o_8_51, o_8_50, o_8_49, o_8_48, o_8_47, o_8_46, o_8_45, o_8_44, o_8_43, o_8_42, o_8_41, o_8_40, o_8_39, o_8_38, o_8_37, o_8_36, o_8_35, o_8_34, o_8_33, o_8_32, o_8_31, o_8_30, o_8_29, o_8_28, o_8_27, o_8_26, o_8_25, o_8_24, o_8_23, o_8_22, o_8_21, o_8_20, o_8_19, o_8_18, o_8_17, o_8_16, o_8_15, o_8_14, o_8_13, o_8_12, o_8_11, o_8_10, o_8_9, o_8_8, o_8_7, o_8_6, o_8_5, o_8_4, o_8_3, o_8_2, o_8_1, o_8_0};
        i_8_0 <= in_reg[0];
        i_8_1 <= in_reg[256];
        i_8_2 <= in_reg[512];
        i_8_3 <= in_reg[768];
        i_8_4 <= in_reg[1024];
        i_8_5 <= in_reg[1280];
        i_8_6 <= in_reg[1536];
        i_8_7 <= in_reg[1792];
        i_8_8 <= in_reg[2048];
        i_8_9 <= in_reg[1];
        i_8_10 <= in_reg[257];
        i_8_11 <= in_reg[513];
        i_8_12 <= in_reg[769];
        i_8_13 <= in_reg[1025];
        i_8_14 <= in_reg[1281];
        i_8_15 <= in_reg[1537];
        i_8_16 <= in_reg[1793];
        i_8_17 <= in_reg[2049];
        i_8_18 <= in_reg[2];
        i_8_19 <= in_reg[258];
        i_8_20 <= in_reg[514];
        i_8_21 <= in_reg[770];
        i_8_22 <= in_reg[1026];
        i_8_23 <= in_reg[1282];
        i_8_24 <= in_reg[1538];
        i_8_25 <= in_reg[1794];
        i_8_26 <= in_reg[2050];
        i_8_27 <= in_reg[3];
        i_8_28 <= in_reg[259];
        i_8_29 <= in_reg[515];
        i_8_30 <= in_reg[771];
        i_8_31 <= in_reg[1027];
        i_8_32 <= in_reg[1283];
        i_8_33 <= in_reg[1539];
        i_8_34 <= in_reg[1795];
        i_8_35 <= in_reg[2051];
        i_8_36 <= in_reg[4];
        i_8_37 <= in_reg[260];
        i_8_38 <= in_reg[516];
        i_8_39 <= in_reg[772];
        i_8_40 <= in_reg[1028];
        i_8_41 <= in_reg[1284];
        i_8_42 <= in_reg[1540];
        i_8_43 <= in_reg[1796];
        i_8_44 <= in_reg[2052];
        i_8_45 <= in_reg[5];
        i_8_46 <= in_reg[261];
        i_8_47 <= in_reg[517];
        i_8_48 <= in_reg[773];
        i_8_49 <= in_reg[1029];
        i_8_50 <= in_reg[1285];
        i_8_51 <= in_reg[1541];
        i_8_52 <= in_reg[1797];
        i_8_53 <= in_reg[2053];
        i_8_54 <= in_reg[6];
        i_8_55 <= in_reg[262];
        i_8_56 <= in_reg[518];
        i_8_57 <= in_reg[774];
        i_8_58 <= in_reg[1030];
        i_8_59 <= in_reg[1286];
        i_8_60 <= in_reg[1542];
        i_8_61 <= in_reg[1798];
        i_8_62 <= in_reg[2054];
        i_8_63 <= in_reg[7];
        i_8_64 <= in_reg[263];
        i_8_65 <= in_reg[519];
        i_8_66 <= in_reg[775];
        i_8_67 <= in_reg[1031];
        i_8_68 <= in_reg[1287];
        i_8_69 <= in_reg[1543];
        i_8_70 <= in_reg[1799];
        i_8_71 <= in_reg[2055];
        i_8_72 <= in_reg[8];
        i_8_73 <= in_reg[264];
        i_8_74 <= in_reg[520];
        i_8_75 <= in_reg[776];
        i_8_76 <= in_reg[1032];
        i_8_77 <= in_reg[1288];
        i_8_78 <= in_reg[1544];
        i_8_79 <= in_reg[1800];
        i_8_80 <= in_reg[2056];
        i_8_81 <= in_reg[9];
        i_8_82 <= in_reg[265];
        i_8_83 <= in_reg[521];
        i_8_84 <= in_reg[777];
        i_8_85 <= in_reg[1033];
        i_8_86 <= in_reg[1289];
        i_8_87 <= in_reg[1545];
        i_8_88 <= in_reg[1801];
        i_8_89 <= in_reg[2057];
        i_8_90 <= in_reg[10];
        i_8_91 <= in_reg[266];
        i_8_92 <= in_reg[522];
        i_8_93 <= in_reg[778];
        i_8_94 <= in_reg[1034];
        i_8_95 <= in_reg[1290];
        i_8_96 <= in_reg[1546];
        i_8_97 <= in_reg[1802];
        i_8_98 <= in_reg[2058];
        i_8_99 <= in_reg[11];
        i_8_100 <= in_reg[267];
        i_8_101 <= in_reg[523];
        i_8_102 <= in_reg[779];
        i_8_103 <= in_reg[1035];
        i_8_104 <= in_reg[1291];
        i_8_105 <= in_reg[1547];
        i_8_106 <= in_reg[1803];
        i_8_107 <= in_reg[2059];
        i_8_108 <= in_reg[12];
        i_8_109 <= in_reg[268];
        i_8_110 <= in_reg[524];
        i_8_111 <= in_reg[780];
        i_8_112 <= in_reg[1036];
        i_8_113 <= in_reg[1292];
        i_8_114 <= in_reg[1548];
        i_8_115 <= in_reg[1804];
        i_8_116 <= in_reg[2060];
        i_8_117 <= in_reg[13];
        i_8_118 <= in_reg[269];
        i_8_119 <= in_reg[525];
        i_8_120 <= in_reg[781];
        i_8_121 <= in_reg[1037];
        i_8_122 <= in_reg[1293];
        i_8_123 <= in_reg[1549];
        i_8_124 <= in_reg[1805];
        i_8_125 <= in_reg[2061];
        i_8_126 <= in_reg[14];
        i_8_127 <= in_reg[270];
        i_8_128 <= in_reg[526];
        i_8_129 <= in_reg[782];
        i_8_130 <= in_reg[1038];
        i_8_131 <= in_reg[1294];
        i_8_132 <= in_reg[1550];
        i_8_133 <= in_reg[1806];
        i_8_134 <= in_reg[2062];
        i_8_135 <= in_reg[15];
        i_8_136 <= in_reg[271];
        i_8_137 <= in_reg[527];
        i_8_138 <= in_reg[783];
        i_8_139 <= in_reg[1039];
        i_8_140 <= in_reg[1295];
        i_8_141 <= in_reg[1551];
        i_8_142 <= in_reg[1807];
        i_8_143 <= in_reg[2063];
        i_8_144 <= in_reg[16];
        i_8_145 <= in_reg[272];
        i_8_146 <= in_reg[528];
        i_8_147 <= in_reg[784];
        i_8_148 <= in_reg[1040];
        i_8_149 <= in_reg[1296];
        i_8_150 <= in_reg[1552];
        i_8_151 <= in_reg[1808];
        i_8_152 <= in_reg[2064];
        i_8_153 <= in_reg[17];
        i_8_154 <= in_reg[273];
        i_8_155 <= in_reg[529];
        i_8_156 <= in_reg[785];
        i_8_157 <= in_reg[1041];
        i_8_158 <= in_reg[1297];
        i_8_159 <= in_reg[1553];
        i_8_160 <= in_reg[1809];
        i_8_161 <= in_reg[2065];
        i_8_162 <= in_reg[18];
        i_8_163 <= in_reg[274];
        i_8_164 <= in_reg[530];
        i_8_165 <= in_reg[786];
        i_8_166 <= in_reg[1042];
        i_8_167 <= in_reg[1298];
        i_8_168 <= in_reg[1554];
        i_8_169 <= in_reg[1810];
        i_8_170 <= in_reg[2066];
        i_8_171 <= in_reg[19];
        i_8_172 <= in_reg[275];
        i_8_173 <= in_reg[531];
        i_8_174 <= in_reg[787];
        i_8_175 <= in_reg[1043];
        i_8_176 <= in_reg[1299];
        i_8_177 <= in_reg[1555];
        i_8_178 <= in_reg[1811];
        i_8_179 <= in_reg[2067];
        i_8_180 <= in_reg[20];
        i_8_181 <= in_reg[276];
        i_8_182 <= in_reg[532];
        i_8_183 <= in_reg[788];
        i_8_184 <= in_reg[1044];
        i_8_185 <= in_reg[1300];
        i_8_186 <= in_reg[1556];
        i_8_187 <= in_reg[1812];
        i_8_188 <= in_reg[2068];
        i_8_189 <= in_reg[21];
        i_8_190 <= in_reg[277];
        i_8_191 <= in_reg[533];
        i_8_192 <= in_reg[789];
        i_8_193 <= in_reg[1045];
        i_8_194 <= in_reg[1301];
        i_8_195 <= in_reg[1557];
        i_8_196 <= in_reg[1813];
        i_8_197 <= in_reg[2069];
        i_8_198 <= in_reg[22];
        i_8_199 <= in_reg[278];
        i_8_200 <= in_reg[534];
        i_8_201 <= in_reg[790];
        i_8_202 <= in_reg[1046];
        i_8_203 <= in_reg[1302];
        i_8_204 <= in_reg[1558];
        i_8_205 <= in_reg[1814];
        i_8_206 <= in_reg[2070];
        i_8_207 <= in_reg[23];
        i_8_208 <= in_reg[279];
        i_8_209 <= in_reg[535];
        i_8_210 <= in_reg[791];
        i_8_211 <= in_reg[1047];
        i_8_212 <= in_reg[1303];
        i_8_213 <= in_reg[1559];
        i_8_214 <= in_reg[1815];
        i_8_215 <= in_reg[2071];
        i_8_216 <= in_reg[24];
        i_8_217 <= in_reg[280];
        i_8_218 <= in_reg[536];
        i_8_219 <= in_reg[792];
        i_8_220 <= in_reg[1048];
        i_8_221 <= in_reg[1304];
        i_8_222 <= in_reg[1560];
        i_8_223 <= in_reg[1816];
        i_8_224 <= in_reg[2072];
        i_8_225 <= in_reg[25];
        i_8_226 <= in_reg[281];
        i_8_227 <= in_reg[537];
        i_8_228 <= in_reg[793];
        i_8_229 <= in_reg[1049];
        i_8_230 <= in_reg[1305];
        i_8_231 <= in_reg[1561];
        i_8_232 <= in_reg[1817];
        i_8_233 <= in_reg[2073];
        i_8_234 <= in_reg[26];
        i_8_235 <= in_reg[282];
        i_8_236 <= in_reg[538];
        i_8_237 <= in_reg[794];
        i_8_238 <= in_reg[1050];
        i_8_239 <= in_reg[1306];
        i_8_240 <= in_reg[1562];
        i_8_241 <= in_reg[1818];
        i_8_242 <= in_reg[2074];
        i_8_243 <= in_reg[27];
        i_8_244 <= in_reg[283];
        i_8_245 <= in_reg[539];
        i_8_246 <= in_reg[795];
        i_8_247 <= in_reg[1051];
        i_8_248 <= in_reg[1307];
        i_8_249 <= in_reg[1563];
        i_8_250 <= in_reg[1819];
        i_8_251 <= in_reg[2075];
        i_8_252 <= in_reg[28];
        i_8_253 <= in_reg[284];
        i_8_254 <= in_reg[540];
        i_8_255 <= in_reg[796];
        i_8_256 <= in_reg[1052];
        i_8_257 <= in_reg[1308];
        i_8_258 <= in_reg[1564];
        i_8_259 <= in_reg[1820];
        i_8_260 <= in_reg[2076];
        i_8_261 <= in_reg[29];
        i_8_262 <= in_reg[285];
        i_8_263 <= in_reg[541];
        i_8_264 <= in_reg[797];
        i_8_265 <= in_reg[1053];
        i_8_266 <= in_reg[1309];
        i_8_267 <= in_reg[1565];
        i_8_268 <= in_reg[1821];
        i_8_269 <= in_reg[2077];
        i_8_270 <= in_reg[30];
        i_8_271 <= in_reg[286];
        i_8_272 <= in_reg[542];
        i_8_273 <= in_reg[798];
        i_8_274 <= in_reg[1054];
        i_8_275 <= in_reg[1310];
        i_8_276 <= in_reg[1566];
        i_8_277 <= in_reg[1822];
        i_8_278 <= in_reg[2078];
        i_8_279 <= in_reg[31];
        i_8_280 <= in_reg[287];
        i_8_281 <= in_reg[543];
        i_8_282 <= in_reg[799];
        i_8_283 <= in_reg[1055];
        i_8_284 <= in_reg[1311];
        i_8_285 <= in_reg[1567];
        i_8_286 <= in_reg[1823];
        i_8_287 <= in_reg[2079];
        i_8_288 <= in_reg[32];
        i_8_289 <= in_reg[288];
        i_8_290 <= in_reg[544];
        i_8_291 <= in_reg[800];
        i_8_292 <= in_reg[1056];
        i_8_293 <= in_reg[1312];
        i_8_294 <= in_reg[1568];
        i_8_295 <= in_reg[1824];
        i_8_296 <= in_reg[2080];
        i_8_297 <= in_reg[33];
        i_8_298 <= in_reg[289];
        i_8_299 <= in_reg[545];
        i_8_300 <= in_reg[801];
        i_8_301 <= in_reg[1057];
        i_8_302 <= in_reg[1313];
        i_8_303 <= in_reg[1569];
        i_8_304 <= in_reg[1825];
        i_8_305 <= in_reg[2081];
        i_8_306 <= in_reg[34];
        i_8_307 <= in_reg[290];
        i_8_308 <= in_reg[546];
        i_8_309 <= in_reg[802];
        i_8_310 <= in_reg[1058];
        i_8_311 <= in_reg[1314];
        i_8_312 <= in_reg[1570];
        i_8_313 <= in_reg[1826];
        i_8_314 <= in_reg[2082];
        i_8_315 <= in_reg[35];
        i_8_316 <= in_reg[291];
        i_8_317 <= in_reg[547];
        i_8_318 <= in_reg[803];
        i_8_319 <= in_reg[1059];
        i_8_320 <= in_reg[1315];
        i_8_321 <= in_reg[1571];
        i_8_322 <= in_reg[1827];
        i_8_323 <= in_reg[2083];
        i_8_324 <= in_reg[36];
        i_8_325 <= in_reg[292];
        i_8_326 <= in_reg[548];
        i_8_327 <= in_reg[804];
        i_8_328 <= in_reg[1060];
        i_8_329 <= in_reg[1316];
        i_8_330 <= in_reg[1572];
        i_8_331 <= in_reg[1828];
        i_8_332 <= in_reg[2084];
        i_8_333 <= in_reg[37];
        i_8_334 <= in_reg[293];
        i_8_335 <= in_reg[549];
        i_8_336 <= in_reg[805];
        i_8_337 <= in_reg[1061];
        i_8_338 <= in_reg[1317];
        i_8_339 <= in_reg[1573];
        i_8_340 <= in_reg[1829];
        i_8_341 <= in_reg[2085];
        i_8_342 <= in_reg[38];
        i_8_343 <= in_reg[294];
        i_8_344 <= in_reg[550];
        i_8_345 <= in_reg[806];
        i_8_346 <= in_reg[1062];
        i_8_347 <= in_reg[1318];
        i_8_348 <= in_reg[1574];
        i_8_349 <= in_reg[1830];
        i_8_350 <= in_reg[2086];
        i_8_351 <= in_reg[39];
        i_8_352 <= in_reg[295];
        i_8_353 <= in_reg[551];
        i_8_354 <= in_reg[807];
        i_8_355 <= in_reg[1063];
        i_8_356 <= in_reg[1319];
        i_8_357 <= in_reg[1575];
        i_8_358 <= in_reg[1831];
        i_8_359 <= in_reg[2087];
        i_8_360 <= in_reg[40];
        i_8_361 <= in_reg[296];
        i_8_362 <= in_reg[552];
        i_8_363 <= in_reg[808];
        i_8_364 <= in_reg[1064];
        i_8_365 <= in_reg[1320];
        i_8_366 <= in_reg[1576];
        i_8_367 <= in_reg[1832];
        i_8_368 <= in_reg[2088];
        i_8_369 <= in_reg[41];
        i_8_370 <= in_reg[297];
        i_8_371 <= in_reg[553];
        i_8_372 <= in_reg[809];
        i_8_373 <= in_reg[1065];
        i_8_374 <= in_reg[1321];
        i_8_375 <= in_reg[1577];
        i_8_376 <= in_reg[1833];
        i_8_377 <= in_reg[2089];
        i_8_378 <= in_reg[42];
        i_8_379 <= in_reg[298];
        i_8_380 <= in_reg[554];
        i_8_381 <= in_reg[810];
        i_8_382 <= in_reg[1066];
        i_8_383 <= in_reg[1322];
        i_8_384 <= in_reg[1578];
        i_8_385 <= in_reg[1834];
        i_8_386 <= in_reg[2090];
        i_8_387 <= in_reg[43];
        i_8_388 <= in_reg[299];
        i_8_389 <= in_reg[555];
        i_8_390 <= in_reg[811];
        i_8_391 <= in_reg[1067];
        i_8_392 <= in_reg[1323];
        i_8_393 <= in_reg[1579];
        i_8_394 <= in_reg[1835];
        i_8_395 <= in_reg[2091];
        i_8_396 <= in_reg[44];
        i_8_397 <= in_reg[300];
        i_8_398 <= in_reg[556];
        i_8_399 <= in_reg[812];
        i_8_400 <= in_reg[1068];
        i_8_401 <= in_reg[1324];
        i_8_402 <= in_reg[1580];
        i_8_403 <= in_reg[1836];
        i_8_404 <= in_reg[2092];
        i_8_405 <= in_reg[45];
        i_8_406 <= in_reg[301];
        i_8_407 <= in_reg[557];
        i_8_408 <= in_reg[813];
        i_8_409 <= in_reg[1069];
        i_8_410 <= in_reg[1325];
        i_8_411 <= in_reg[1581];
        i_8_412 <= in_reg[1837];
        i_8_413 <= in_reg[2093];
        i_8_414 <= in_reg[46];
        i_8_415 <= in_reg[302];
        i_8_416 <= in_reg[558];
        i_8_417 <= in_reg[814];
        i_8_418 <= in_reg[1070];
        i_8_419 <= in_reg[1326];
        i_8_420 <= in_reg[1582];
        i_8_421 <= in_reg[1838];
        i_8_422 <= in_reg[2094];
        i_8_423 <= in_reg[47];
        i_8_424 <= in_reg[303];
        i_8_425 <= in_reg[559];
        i_8_426 <= in_reg[815];
        i_8_427 <= in_reg[1071];
        i_8_428 <= in_reg[1327];
        i_8_429 <= in_reg[1583];
        i_8_430 <= in_reg[1839];
        i_8_431 <= in_reg[2095];
        i_8_432 <= in_reg[48];
        i_8_433 <= in_reg[304];
        i_8_434 <= in_reg[560];
        i_8_435 <= in_reg[816];
        i_8_436 <= in_reg[1072];
        i_8_437 <= in_reg[1328];
        i_8_438 <= in_reg[1584];
        i_8_439 <= in_reg[1840];
        i_8_440 <= in_reg[2096];
        i_8_441 <= in_reg[49];
        i_8_442 <= in_reg[305];
        i_8_443 <= in_reg[561];
        i_8_444 <= in_reg[817];
        i_8_445 <= in_reg[1073];
        i_8_446 <= in_reg[1329];
        i_8_447 <= in_reg[1585];
        i_8_448 <= in_reg[1841];
        i_8_449 <= in_reg[2097];
        i_8_450 <= in_reg[50];
        i_8_451 <= in_reg[306];
        i_8_452 <= in_reg[562];
        i_8_453 <= in_reg[818];
        i_8_454 <= in_reg[1074];
        i_8_455 <= in_reg[1330];
        i_8_456 <= in_reg[1586];
        i_8_457 <= in_reg[1842];
        i_8_458 <= in_reg[2098];
        i_8_459 <= in_reg[51];
        i_8_460 <= in_reg[307];
        i_8_461 <= in_reg[563];
        i_8_462 <= in_reg[819];
        i_8_463 <= in_reg[1075];
        i_8_464 <= in_reg[1331];
        i_8_465 <= in_reg[1587];
        i_8_466 <= in_reg[1843];
        i_8_467 <= in_reg[2099];
        i_8_468 <= in_reg[52];
        i_8_469 <= in_reg[308];
        i_8_470 <= in_reg[564];
        i_8_471 <= in_reg[820];
        i_8_472 <= in_reg[1076];
        i_8_473 <= in_reg[1332];
        i_8_474 <= in_reg[1588];
        i_8_475 <= in_reg[1844];
        i_8_476 <= in_reg[2100];
        i_8_477 <= in_reg[53];
        i_8_478 <= in_reg[309];
        i_8_479 <= in_reg[565];
        i_8_480 <= in_reg[821];
        i_8_481 <= in_reg[1077];
        i_8_482 <= in_reg[1333];
        i_8_483 <= in_reg[1589];
        i_8_484 <= in_reg[1845];
        i_8_485 <= in_reg[2101];
        i_8_486 <= in_reg[54];
        i_8_487 <= in_reg[310];
        i_8_488 <= in_reg[566];
        i_8_489 <= in_reg[822];
        i_8_490 <= in_reg[1078];
        i_8_491 <= in_reg[1334];
        i_8_492 <= in_reg[1590];
        i_8_493 <= in_reg[1846];
        i_8_494 <= in_reg[2102];
        i_8_495 <= in_reg[55];
        i_8_496 <= in_reg[311];
        i_8_497 <= in_reg[567];
        i_8_498 <= in_reg[823];
        i_8_499 <= in_reg[1079];
        i_8_500 <= in_reg[1335];
        i_8_501 <= in_reg[1591];
        i_8_502 <= in_reg[1847];
        i_8_503 <= in_reg[2103];
        i_8_504 <= in_reg[56];
        i_8_505 <= in_reg[312];
        i_8_506 <= in_reg[568];
        i_8_507 <= in_reg[824];
        i_8_508 <= in_reg[1080];
        i_8_509 <= in_reg[1336];
        i_8_510 <= in_reg[1592];
        i_8_511 <= in_reg[1848];
        i_8_512 <= in_reg[2104];
        i_8_513 <= in_reg[57];
        i_8_514 <= in_reg[313];
        i_8_515 <= in_reg[569];
        i_8_516 <= in_reg[825];
        i_8_517 <= in_reg[1081];
        i_8_518 <= in_reg[1337];
        i_8_519 <= in_reg[1593];
        i_8_520 <= in_reg[1849];
        i_8_521 <= in_reg[2105];
        i_8_522 <= in_reg[58];
        i_8_523 <= in_reg[314];
        i_8_524 <= in_reg[570];
        i_8_525 <= in_reg[826];
        i_8_526 <= in_reg[1082];
        i_8_527 <= in_reg[1338];
        i_8_528 <= in_reg[1594];
        i_8_529 <= in_reg[1850];
        i_8_530 <= in_reg[2106];
        i_8_531 <= in_reg[59];
        i_8_532 <= in_reg[315];
        i_8_533 <= in_reg[571];
        i_8_534 <= in_reg[827];
        i_8_535 <= in_reg[1083];
        i_8_536 <= in_reg[1339];
        i_8_537 <= in_reg[1595];
        i_8_538 <= in_reg[1851];
        i_8_539 <= in_reg[2107];
        i_8_540 <= in_reg[60];
        i_8_541 <= in_reg[316];
        i_8_542 <= in_reg[572];
        i_8_543 <= in_reg[828];
        i_8_544 <= in_reg[1084];
        i_8_545 <= in_reg[1340];
        i_8_546 <= in_reg[1596];
        i_8_547 <= in_reg[1852];
        i_8_548 <= in_reg[2108];
        i_8_549 <= in_reg[61];
        i_8_550 <= in_reg[317];
        i_8_551 <= in_reg[573];
        i_8_552 <= in_reg[829];
        i_8_553 <= in_reg[1085];
        i_8_554 <= in_reg[1341];
        i_8_555 <= in_reg[1597];
        i_8_556 <= in_reg[1853];
        i_8_557 <= in_reg[2109];
        i_8_558 <= in_reg[62];
        i_8_559 <= in_reg[318];
        i_8_560 <= in_reg[574];
        i_8_561 <= in_reg[830];
        i_8_562 <= in_reg[1086];
        i_8_563 <= in_reg[1342];
        i_8_564 <= in_reg[1598];
        i_8_565 <= in_reg[1854];
        i_8_566 <= in_reg[2110];
        i_8_567 <= in_reg[63];
        i_8_568 <= in_reg[319];
        i_8_569 <= in_reg[575];
        i_8_570 <= in_reg[831];
        i_8_571 <= in_reg[1087];
        i_8_572 <= in_reg[1343];
        i_8_573 <= in_reg[1599];
        i_8_574 <= in_reg[1855];
        i_8_575 <= in_reg[2111];
        i_8_576 <= in_reg[64];
        i_8_577 <= in_reg[320];
        i_8_578 <= in_reg[576];
        i_8_579 <= in_reg[832];
        i_8_580 <= in_reg[1088];
        i_8_581 <= in_reg[1344];
        i_8_582 <= in_reg[1600];
        i_8_583 <= in_reg[1856];
        i_8_584 <= in_reg[2112];
        i_8_585 <= in_reg[65];
        i_8_586 <= in_reg[321];
        i_8_587 <= in_reg[577];
        i_8_588 <= in_reg[833];
        i_8_589 <= in_reg[1089];
        i_8_590 <= in_reg[1345];
        i_8_591 <= in_reg[1601];
        i_8_592 <= in_reg[1857];
        i_8_593 <= in_reg[2113];
        i_8_594 <= in_reg[66];
        i_8_595 <= in_reg[322];
        i_8_596 <= in_reg[578];
        i_8_597 <= in_reg[834];
        i_8_598 <= in_reg[1090];
        i_8_599 <= in_reg[1346];
        i_8_600 <= in_reg[1602];
        i_8_601 <= in_reg[1858];
        i_8_602 <= in_reg[2114];
        i_8_603 <= in_reg[67];
        i_8_604 <= in_reg[323];
        i_8_605 <= in_reg[579];
        i_8_606 <= in_reg[835];
        i_8_607 <= in_reg[1091];
        i_8_608 <= in_reg[1347];
        i_8_609 <= in_reg[1603];
        i_8_610 <= in_reg[1859];
        i_8_611 <= in_reg[2115];
        i_8_612 <= in_reg[68];
        i_8_613 <= in_reg[324];
        i_8_614 <= in_reg[580];
        i_8_615 <= in_reg[836];
        i_8_616 <= in_reg[1092];
        i_8_617 <= in_reg[1348];
        i_8_618 <= in_reg[1604];
        i_8_619 <= in_reg[1860];
        i_8_620 <= in_reg[2116];
        i_8_621 <= in_reg[69];
        i_8_622 <= in_reg[325];
        i_8_623 <= in_reg[581];
        i_8_624 <= in_reg[837];
        i_8_625 <= in_reg[1093];
        i_8_626 <= in_reg[1349];
        i_8_627 <= in_reg[1605];
        i_8_628 <= in_reg[1861];
        i_8_629 <= in_reg[2117];
        i_8_630 <= in_reg[70];
        i_8_631 <= in_reg[326];
        i_8_632 <= in_reg[582];
        i_8_633 <= in_reg[838];
        i_8_634 <= in_reg[1094];
        i_8_635 <= in_reg[1350];
        i_8_636 <= in_reg[1606];
        i_8_637 <= in_reg[1862];
        i_8_638 <= in_reg[2118];
        i_8_639 <= in_reg[71];
        i_8_640 <= in_reg[327];
        i_8_641 <= in_reg[583];
        i_8_642 <= in_reg[839];
        i_8_643 <= in_reg[1095];
        i_8_644 <= in_reg[1351];
        i_8_645 <= in_reg[1607];
        i_8_646 <= in_reg[1863];
        i_8_647 <= in_reg[2119];
        i_8_648 <= in_reg[72];
        i_8_649 <= in_reg[328];
        i_8_650 <= in_reg[584];
        i_8_651 <= in_reg[840];
        i_8_652 <= in_reg[1096];
        i_8_653 <= in_reg[1352];
        i_8_654 <= in_reg[1608];
        i_8_655 <= in_reg[1864];
        i_8_656 <= in_reg[2120];
        i_8_657 <= in_reg[73];
        i_8_658 <= in_reg[329];
        i_8_659 <= in_reg[585];
        i_8_660 <= in_reg[841];
        i_8_661 <= in_reg[1097];
        i_8_662 <= in_reg[1353];
        i_8_663 <= in_reg[1609];
        i_8_664 <= in_reg[1865];
        i_8_665 <= in_reg[2121];
        i_8_666 <= in_reg[74];
        i_8_667 <= in_reg[330];
        i_8_668 <= in_reg[586];
        i_8_669 <= in_reg[842];
        i_8_670 <= in_reg[1098];
        i_8_671 <= in_reg[1354];
        i_8_672 <= in_reg[1610];
        i_8_673 <= in_reg[1866];
        i_8_674 <= in_reg[2122];
        i_8_675 <= in_reg[75];
        i_8_676 <= in_reg[331];
        i_8_677 <= in_reg[587];
        i_8_678 <= in_reg[843];
        i_8_679 <= in_reg[1099];
        i_8_680 <= in_reg[1355];
        i_8_681 <= in_reg[1611];
        i_8_682 <= in_reg[1867];
        i_8_683 <= in_reg[2123];
        i_8_684 <= in_reg[76];
        i_8_685 <= in_reg[332];
        i_8_686 <= in_reg[588];
        i_8_687 <= in_reg[844];
        i_8_688 <= in_reg[1100];
        i_8_689 <= in_reg[1356];
        i_8_690 <= in_reg[1612];
        i_8_691 <= in_reg[1868];
        i_8_692 <= in_reg[2124];
        i_8_693 <= in_reg[77];
        i_8_694 <= in_reg[333];
        i_8_695 <= in_reg[589];
        i_8_696 <= in_reg[845];
        i_8_697 <= in_reg[1101];
        i_8_698 <= in_reg[1357];
        i_8_699 <= in_reg[1613];
        i_8_700 <= in_reg[1869];
        i_8_701 <= in_reg[2125];
        i_8_702 <= in_reg[78];
        i_8_703 <= in_reg[334];
        i_8_704 <= in_reg[590];
        i_8_705 <= in_reg[846];
        i_8_706 <= in_reg[1102];
        i_8_707 <= in_reg[1358];
        i_8_708 <= in_reg[1614];
        i_8_709 <= in_reg[1870];
        i_8_710 <= in_reg[2126];
        i_8_711 <= in_reg[79];
        i_8_712 <= in_reg[335];
        i_8_713 <= in_reg[591];
        i_8_714 <= in_reg[847];
        i_8_715 <= in_reg[1103];
        i_8_716 <= in_reg[1359];
        i_8_717 <= in_reg[1615];
        i_8_718 <= in_reg[1871];
        i_8_719 <= in_reg[2127];
        i_8_720 <= in_reg[80];
        i_8_721 <= in_reg[336];
        i_8_722 <= in_reg[592];
        i_8_723 <= in_reg[848];
        i_8_724 <= in_reg[1104];
        i_8_725 <= in_reg[1360];
        i_8_726 <= in_reg[1616];
        i_8_727 <= in_reg[1872];
        i_8_728 <= in_reg[2128];
        i_8_729 <= in_reg[81];
        i_8_730 <= in_reg[337];
        i_8_731 <= in_reg[593];
        i_8_732 <= in_reg[849];
        i_8_733 <= in_reg[1105];
        i_8_734 <= in_reg[1361];
        i_8_735 <= in_reg[1617];
        i_8_736 <= in_reg[1873];
        i_8_737 <= in_reg[2129];
        i_8_738 <= in_reg[82];
        i_8_739 <= in_reg[338];
        i_8_740 <= in_reg[594];
        i_8_741 <= in_reg[850];
        i_8_742 <= in_reg[1106];
        i_8_743 <= in_reg[1362];
        i_8_744 <= in_reg[1618];
        i_8_745 <= in_reg[1874];
        i_8_746 <= in_reg[2130];
        i_8_747 <= in_reg[83];
        i_8_748 <= in_reg[339];
        i_8_749 <= in_reg[595];
        i_8_750 <= in_reg[851];
        i_8_751 <= in_reg[1107];
        i_8_752 <= in_reg[1363];
        i_8_753 <= in_reg[1619];
        i_8_754 <= in_reg[1875];
        i_8_755 <= in_reg[2131];
        i_8_756 <= in_reg[84];
        i_8_757 <= in_reg[340];
        i_8_758 <= in_reg[596];
        i_8_759 <= in_reg[852];
        i_8_760 <= in_reg[1108];
        i_8_761 <= in_reg[1364];
        i_8_762 <= in_reg[1620];
        i_8_763 <= in_reg[1876];
        i_8_764 <= in_reg[2132];
        i_8_765 <= in_reg[85];
        i_8_766 <= in_reg[341];
        i_8_767 <= in_reg[597];
        i_8_768 <= in_reg[853];
        i_8_769 <= in_reg[1109];
        i_8_770 <= in_reg[1365];
        i_8_771 <= in_reg[1621];
        i_8_772 <= in_reg[1877];
        i_8_773 <= in_reg[2133];
        i_8_774 <= in_reg[86];
        i_8_775 <= in_reg[342];
        i_8_776 <= in_reg[598];
        i_8_777 <= in_reg[854];
        i_8_778 <= in_reg[1110];
        i_8_779 <= in_reg[1366];
        i_8_780 <= in_reg[1622];
        i_8_781 <= in_reg[1878];
        i_8_782 <= in_reg[2134];
        i_8_783 <= in_reg[87];
        i_8_784 <= in_reg[343];
        i_8_785 <= in_reg[599];
        i_8_786 <= in_reg[855];
        i_8_787 <= in_reg[1111];
        i_8_788 <= in_reg[1367];
        i_8_789 <= in_reg[1623];
        i_8_790 <= in_reg[1879];
        i_8_791 <= in_reg[2135];
        i_8_792 <= in_reg[88];
        i_8_793 <= in_reg[344];
        i_8_794 <= in_reg[600];
        i_8_795 <= in_reg[856];
        i_8_796 <= in_reg[1112];
        i_8_797 <= in_reg[1368];
        i_8_798 <= in_reg[1624];
        i_8_799 <= in_reg[1880];
        i_8_800 <= in_reg[2136];
        i_8_801 <= in_reg[89];
        i_8_802 <= in_reg[345];
        i_8_803 <= in_reg[601];
        i_8_804 <= in_reg[857];
        i_8_805 <= in_reg[1113];
        i_8_806 <= in_reg[1369];
        i_8_807 <= in_reg[1625];
        i_8_808 <= in_reg[1881];
        i_8_809 <= in_reg[2137];
        i_8_810 <= in_reg[90];
        i_8_811 <= in_reg[346];
        i_8_812 <= in_reg[602];
        i_8_813 <= in_reg[858];
        i_8_814 <= in_reg[1114];
        i_8_815 <= in_reg[1370];
        i_8_816 <= in_reg[1626];
        i_8_817 <= in_reg[1882];
        i_8_818 <= in_reg[2138];
        i_8_819 <= in_reg[91];
        i_8_820 <= in_reg[347];
        i_8_821 <= in_reg[603];
        i_8_822 <= in_reg[859];
        i_8_823 <= in_reg[1115];
        i_8_824 <= in_reg[1371];
        i_8_825 <= in_reg[1627];
        i_8_826 <= in_reg[1883];
        i_8_827 <= in_reg[2139];
        i_8_828 <= in_reg[92];
        i_8_829 <= in_reg[348];
        i_8_830 <= in_reg[604];
        i_8_831 <= in_reg[860];
        i_8_832 <= in_reg[1116];
        i_8_833 <= in_reg[1372];
        i_8_834 <= in_reg[1628];
        i_8_835 <= in_reg[1884];
        i_8_836 <= in_reg[2140];
        i_8_837 <= in_reg[93];
        i_8_838 <= in_reg[349];
        i_8_839 <= in_reg[605];
        i_8_840 <= in_reg[861];
        i_8_841 <= in_reg[1117];
        i_8_842 <= in_reg[1373];
        i_8_843 <= in_reg[1629];
        i_8_844 <= in_reg[1885];
        i_8_845 <= in_reg[2141];
        i_8_846 <= in_reg[94];
        i_8_847 <= in_reg[350];
        i_8_848 <= in_reg[606];
        i_8_849 <= in_reg[862];
        i_8_850 <= in_reg[1118];
        i_8_851 <= in_reg[1374];
        i_8_852 <= in_reg[1630];
        i_8_853 <= in_reg[1886];
        i_8_854 <= in_reg[2142];
        i_8_855 <= in_reg[95];
        i_8_856 <= in_reg[351];
        i_8_857 <= in_reg[607];
        i_8_858 <= in_reg[863];
        i_8_859 <= in_reg[1119];
        i_8_860 <= in_reg[1375];
        i_8_861 <= in_reg[1631];
        i_8_862 <= in_reg[1887];
        i_8_863 <= in_reg[2143];
        i_8_864 <= in_reg[96];
        i_8_865 <= in_reg[352];
        i_8_866 <= in_reg[608];
        i_8_867 <= in_reg[864];
        i_8_868 <= in_reg[1120];
        i_8_869 <= in_reg[1376];
        i_8_870 <= in_reg[1632];
        i_8_871 <= in_reg[1888];
        i_8_872 <= in_reg[2144];
        i_8_873 <= in_reg[97];
        i_8_874 <= in_reg[353];
        i_8_875 <= in_reg[609];
        i_8_876 <= in_reg[865];
        i_8_877 <= in_reg[1121];
        i_8_878 <= in_reg[1377];
        i_8_879 <= in_reg[1633];
        i_8_880 <= in_reg[1889];
        i_8_881 <= in_reg[2145];
        i_8_882 <= in_reg[98];
        i_8_883 <= in_reg[354];
        i_8_884 <= in_reg[610];
        i_8_885 <= in_reg[866];
        i_8_886 <= in_reg[1122];
        i_8_887 <= in_reg[1378];
        i_8_888 <= in_reg[1634];
        i_8_889 <= in_reg[1890];
        i_8_890 <= in_reg[2146];
        i_8_891 <= in_reg[99];
        i_8_892 <= in_reg[355];
        i_8_893 <= in_reg[611];
        i_8_894 <= in_reg[867];
        i_8_895 <= in_reg[1123];
        i_8_896 <= in_reg[1379];
        i_8_897 <= in_reg[1635];
        i_8_898 <= in_reg[1891];
        i_8_899 <= in_reg[2147];
        i_8_900 <= in_reg[100];
        i_8_901 <= in_reg[356];
        i_8_902 <= in_reg[612];
        i_8_903 <= in_reg[868];
        i_8_904 <= in_reg[1124];
        i_8_905 <= in_reg[1380];
        i_8_906 <= in_reg[1636];
        i_8_907 <= in_reg[1892];
        i_8_908 <= in_reg[2148];
        i_8_909 <= in_reg[101];
        i_8_910 <= in_reg[357];
        i_8_911 <= in_reg[613];
        i_8_912 <= in_reg[869];
        i_8_913 <= in_reg[1125];
        i_8_914 <= in_reg[1381];
        i_8_915 <= in_reg[1637];
        i_8_916 <= in_reg[1893];
        i_8_917 <= in_reg[2149];
        i_8_918 <= in_reg[102];
        i_8_919 <= in_reg[358];
        i_8_920 <= in_reg[614];
        i_8_921 <= in_reg[870];
        i_8_922 <= in_reg[1126];
        i_8_923 <= in_reg[1382];
        i_8_924 <= in_reg[1638];
        i_8_925 <= in_reg[1894];
        i_8_926 <= in_reg[2150];
        i_8_927 <= in_reg[103];
        i_8_928 <= in_reg[359];
        i_8_929 <= in_reg[615];
        i_8_930 <= in_reg[871];
        i_8_931 <= in_reg[1127];
        i_8_932 <= in_reg[1383];
        i_8_933 <= in_reg[1639];
        i_8_934 <= in_reg[1895];
        i_8_935 <= in_reg[2151];
        i_8_936 <= in_reg[104];
        i_8_937 <= in_reg[360];
        i_8_938 <= in_reg[616];
        i_8_939 <= in_reg[872];
        i_8_940 <= in_reg[1128];
        i_8_941 <= in_reg[1384];
        i_8_942 <= in_reg[1640];
        i_8_943 <= in_reg[1896];
        i_8_944 <= in_reg[2152];
        i_8_945 <= in_reg[105];
        i_8_946 <= in_reg[361];
        i_8_947 <= in_reg[617];
        i_8_948 <= in_reg[873];
        i_8_949 <= in_reg[1129];
        i_8_950 <= in_reg[1385];
        i_8_951 <= in_reg[1641];
        i_8_952 <= in_reg[1897];
        i_8_953 <= in_reg[2153];
        i_8_954 <= in_reg[106];
        i_8_955 <= in_reg[362];
        i_8_956 <= in_reg[618];
        i_8_957 <= in_reg[874];
        i_8_958 <= in_reg[1130];
        i_8_959 <= in_reg[1386];
        i_8_960 <= in_reg[1642];
        i_8_961 <= in_reg[1898];
        i_8_962 <= in_reg[2154];
        i_8_963 <= in_reg[107];
        i_8_964 <= in_reg[363];
        i_8_965 <= in_reg[619];
        i_8_966 <= in_reg[875];
        i_8_967 <= in_reg[1131];
        i_8_968 <= in_reg[1387];
        i_8_969 <= in_reg[1643];
        i_8_970 <= in_reg[1899];
        i_8_971 <= in_reg[2155];
        i_8_972 <= in_reg[108];
        i_8_973 <= in_reg[364];
        i_8_974 <= in_reg[620];
        i_8_975 <= in_reg[876];
        i_8_976 <= in_reg[1132];
        i_8_977 <= in_reg[1388];
        i_8_978 <= in_reg[1644];
        i_8_979 <= in_reg[1900];
        i_8_980 <= in_reg[2156];
        i_8_981 <= in_reg[109];
        i_8_982 <= in_reg[365];
        i_8_983 <= in_reg[621];
        i_8_984 <= in_reg[877];
        i_8_985 <= in_reg[1133];
        i_8_986 <= in_reg[1389];
        i_8_987 <= in_reg[1645];
        i_8_988 <= in_reg[1901];
        i_8_989 <= in_reg[2157];
        i_8_990 <= in_reg[110];
        i_8_991 <= in_reg[366];
        i_8_992 <= in_reg[622];
        i_8_993 <= in_reg[878];
        i_8_994 <= in_reg[1134];
        i_8_995 <= in_reg[1390];
        i_8_996 <= in_reg[1646];
        i_8_997 <= in_reg[1902];
        i_8_998 <= in_reg[2158];
        i_8_999 <= in_reg[111];
        i_8_1000 <= in_reg[367];
        i_8_1001 <= in_reg[623];
        i_8_1002 <= in_reg[879];
        i_8_1003 <= in_reg[1135];
        i_8_1004 <= in_reg[1391];
        i_8_1005 <= in_reg[1647];
        i_8_1006 <= in_reg[1903];
        i_8_1007 <= in_reg[2159];
        i_8_1008 <= in_reg[112];
        i_8_1009 <= in_reg[368];
        i_8_1010 <= in_reg[624];
        i_8_1011 <= in_reg[880];
        i_8_1012 <= in_reg[1136];
        i_8_1013 <= in_reg[1392];
        i_8_1014 <= in_reg[1648];
        i_8_1015 <= in_reg[1904];
        i_8_1016 <= in_reg[2160];
        i_8_1017 <= in_reg[113];
        i_8_1018 <= in_reg[369];
        i_8_1019 <= in_reg[625];
        i_8_1020 <= in_reg[881];
        i_8_1021 <= in_reg[1137];
        i_8_1022 <= in_reg[1393];
        i_8_1023 <= in_reg[1649];
        i_8_1024 <= in_reg[1905];
        i_8_1025 <= in_reg[2161];
        i_8_1026 <= in_reg[114];
        i_8_1027 <= in_reg[370];
        i_8_1028 <= in_reg[626];
        i_8_1029 <= in_reg[882];
        i_8_1030 <= in_reg[1138];
        i_8_1031 <= in_reg[1394];
        i_8_1032 <= in_reg[1650];
        i_8_1033 <= in_reg[1906];
        i_8_1034 <= in_reg[2162];
        i_8_1035 <= in_reg[115];
        i_8_1036 <= in_reg[371];
        i_8_1037 <= in_reg[627];
        i_8_1038 <= in_reg[883];
        i_8_1039 <= in_reg[1139];
        i_8_1040 <= in_reg[1395];
        i_8_1041 <= in_reg[1651];
        i_8_1042 <= in_reg[1907];
        i_8_1043 <= in_reg[2163];
        i_8_1044 <= in_reg[116];
        i_8_1045 <= in_reg[372];
        i_8_1046 <= in_reg[628];
        i_8_1047 <= in_reg[884];
        i_8_1048 <= in_reg[1140];
        i_8_1049 <= in_reg[1396];
        i_8_1050 <= in_reg[1652];
        i_8_1051 <= in_reg[1908];
        i_8_1052 <= in_reg[2164];
        i_8_1053 <= in_reg[117];
        i_8_1054 <= in_reg[373];
        i_8_1055 <= in_reg[629];
        i_8_1056 <= in_reg[885];
        i_8_1057 <= in_reg[1141];
        i_8_1058 <= in_reg[1397];
        i_8_1059 <= in_reg[1653];
        i_8_1060 <= in_reg[1909];
        i_8_1061 <= in_reg[2165];
        i_8_1062 <= in_reg[118];
        i_8_1063 <= in_reg[374];
        i_8_1064 <= in_reg[630];
        i_8_1065 <= in_reg[886];
        i_8_1066 <= in_reg[1142];
        i_8_1067 <= in_reg[1398];
        i_8_1068 <= in_reg[1654];
        i_8_1069 <= in_reg[1910];
        i_8_1070 <= in_reg[2166];
        i_8_1071 <= in_reg[119];
        i_8_1072 <= in_reg[375];
        i_8_1073 <= in_reg[631];
        i_8_1074 <= in_reg[887];
        i_8_1075 <= in_reg[1143];
        i_8_1076 <= in_reg[1399];
        i_8_1077 <= in_reg[1655];
        i_8_1078 <= in_reg[1911];
        i_8_1079 <= in_reg[2167];
        i_8_1080 <= in_reg[120];
        i_8_1081 <= in_reg[376];
        i_8_1082 <= in_reg[632];
        i_8_1083 <= in_reg[888];
        i_8_1084 <= in_reg[1144];
        i_8_1085 <= in_reg[1400];
        i_8_1086 <= in_reg[1656];
        i_8_1087 <= in_reg[1912];
        i_8_1088 <= in_reg[2168];
        i_8_1089 <= in_reg[121];
        i_8_1090 <= in_reg[377];
        i_8_1091 <= in_reg[633];
        i_8_1092 <= in_reg[889];
        i_8_1093 <= in_reg[1145];
        i_8_1094 <= in_reg[1401];
        i_8_1095 <= in_reg[1657];
        i_8_1096 <= in_reg[1913];
        i_8_1097 <= in_reg[2169];
        i_8_1098 <= in_reg[122];
        i_8_1099 <= in_reg[378];
        i_8_1100 <= in_reg[634];
        i_8_1101 <= in_reg[890];
        i_8_1102 <= in_reg[1146];
        i_8_1103 <= in_reg[1402];
        i_8_1104 <= in_reg[1658];
        i_8_1105 <= in_reg[1914];
        i_8_1106 <= in_reg[2170];
        i_8_1107 <= in_reg[123];
        i_8_1108 <= in_reg[379];
        i_8_1109 <= in_reg[635];
        i_8_1110 <= in_reg[891];
        i_8_1111 <= in_reg[1147];
        i_8_1112 <= in_reg[1403];
        i_8_1113 <= in_reg[1659];
        i_8_1114 <= in_reg[1915];
        i_8_1115 <= in_reg[2171];
        i_8_1116 <= in_reg[124];
        i_8_1117 <= in_reg[380];
        i_8_1118 <= in_reg[636];
        i_8_1119 <= in_reg[892];
        i_8_1120 <= in_reg[1148];
        i_8_1121 <= in_reg[1404];
        i_8_1122 <= in_reg[1660];
        i_8_1123 <= in_reg[1916];
        i_8_1124 <= in_reg[2172];
        i_8_1125 <= in_reg[125];
        i_8_1126 <= in_reg[381];
        i_8_1127 <= in_reg[637];
        i_8_1128 <= in_reg[893];
        i_8_1129 <= in_reg[1149];
        i_8_1130 <= in_reg[1405];
        i_8_1131 <= in_reg[1661];
        i_8_1132 <= in_reg[1917];
        i_8_1133 <= in_reg[2173];
        i_8_1134 <= in_reg[126];
        i_8_1135 <= in_reg[382];
        i_8_1136 <= in_reg[638];
        i_8_1137 <= in_reg[894];
        i_8_1138 <= in_reg[1150];
        i_8_1139 <= in_reg[1406];
        i_8_1140 <= in_reg[1662];
        i_8_1141 <= in_reg[1918];
        i_8_1142 <= in_reg[2174];
        i_8_1143 <= in_reg[127];
        i_8_1144 <= in_reg[383];
        i_8_1145 <= in_reg[639];
        i_8_1146 <= in_reg[895];
        i_8_1147 <= in_reg[1151];
        i_8_1148 <= in_reg[1407];
        i_8_1149 <= in_reg[1663];
        i_8_1150 <= in_reg[1919];
        i_8_1151 <= in_reg[2175];
        i_8_1152 <= in_reg[128];
        i_8_1153 <= in_reg[384];
        i_8_1154 <= in_reg[640];
        i_8_1155 <= in_reg[896];
        i_8_1156 <= in_reg[1152];
        i_8_1157 <= in_reg[1408];
        i_8_1158 <= in_reg[1664];
        i_8_1159 <= in_reg[1920];
        i_8_1160 <= in_reg[2176];
        i_8_1161 <= in_reg[129];
        i_8_1162 <= in_reg[385];
        i_8_1163 <= in_reg[641];
        i_8_1164 <= in_reg[897];
        i_8_1165 <= in_reg[1153];
        i_8_1166 <= in_reg[1409];
        i_8_1167 <= in_reg[1665];
        i_8_1168 <= in_reg[1921];
        i_8_1169 <= in_reg[2177];
        i_8_1170 <= in_reg[130];
        i_8_1171 <= in_reg[386];
        i_8_1172 <= in_reg[642];
        i_8_1173 <= in_reg[898];
        i_8_1174 <= in_reg[1154];
        i_8_1175 <= in_reg[1410];
        i_8_1176 <= in_reg[1666];
        i_8_1177 <= in_reg[1922];
        i_8_1178 <= in_reg[2178];
        i_8_1179 <= in_reg[131];
        i_8_1180 <= in_reg[387];
        i_8_1181 <= in_reg[643];
        i_8_1182 <= in_reg[899];
        i_8_1183 <= in_reg[1155];
        i_8_1184 <= in_reg[1411];
        i_8_1185 <= in_reg[1667];
        i_8_1186 <= in_reg[1923];
        i_8_1187 <= in_reg[2179];
        i_8_1188 <= in_reg[132];
        i_8_1189 <= in_reg[388];
        i_8_1190 <= in_reg[644];
        i_8_1191 <= in_reg[900];
        i_8_1192 <= in_reg[1156];
        i_8_1193 <= in_reg[1412];
        i_8_1194 <= in_reg[1668];
        i_8_1195 <= in_reg[1924];
        i_8_1196 <= in_reg[2180];
        i_8_1197 <= in_reg[133];
        i_8_1198 <= in_reg[389];
        i_8_1199 <= in_reg[645];
        i_8_1200 <= in_reg[901];
        i_8_1201 <= in_reg[1157];
        i_8_1202 <= in_reg[1413];
        i_8_1203 <= in_reg[1669];
        i_8_1204 <= in_reg[1925];
        i_8_1205 <= in_reg[2181];
        i_8_1206 <= in_reg[134];
        i_8_1207 <= in_reg[390];
        i_8_1208 <= in_reg[646];
        i_8_1209 <= in_reg[902];
        i_8_1210 <= in_reg[1158];
        i_8_1211 <= in_reg[1414];
        i_8_1212 <= in_reg[1670];
        i_8_1213 <= in_reg[1926];
        i_8_1214 <= in_reg[2182];
        i_8_1215 <= in_reg[135];
        i_8_1216 <= in_reg[391];
        i_8_1217 <= in_reg[647];
        i_8_1218 <= in_reg[903];
        i_8_1219 <= in_reg[1159];
        i_8_1220 <= in_reg[1415];
        i_8_1221 <= in_reg[1671];
        i_8_1222 <= in_reg[1927];
        i_8_1223 <= in_reg[2183];
        i_8_1224 <= in_reg[136];
        i_8_1225 <= in_reg[392];
        i_8_1226 <= in_reg[648];
        i_8_1227 <= in_reg[904];
        i_8_1228 <= in_reg[1160];
        i_8_1229 <= in_reg[1416];
        i_8_1230 <= in_reg[1672];
        i_8_1231 <= in_reg[1928];
        i_8_1232 <= in_reg[2184];
        i_8_1233 <= in_reg[137];
        i_8_1234 <= in_reg[393];
        i_8_1235 <= in_reg[649];
        i_8_1236 <= in_reg[905];
        i_8_1237 <= in_reg[1161];
        i_8_1238 <= in_reg[1417];
        i_8_1239 <= in_reg[1673];
        i_8_1240 <= in_reg[1929];
        i_8_1241 <= in_reg[2185];
        i_8_1242 <= in_reg[138];
        i_8_1243 <= in_reg[394];
        i_8_1244 <= in_reg[650];
        i_8_1245 <= in_reg[906];
        i_8_1246 <= in_reg[1162];
        i_8_1247 <= in_reg[1418];
        i_8_1248 <= in_reg[1674];
        i_8_1249 <= in_reg[1930];
        i_8_1250 <= in_reg[2186];
        i_8_1251 <= in_reg[139];
        i_8_1252 <= in_reg[395];
        i_8_1253 <= in_reg[651];
        i_8_1254 <= in_reg[907];
        i_8_1255 <= in_reg[1163];
        i_8_1256 <= in_reg[1419];
        i_8_1257 <= in_reg[1675];
        i_8_1258 <= in_reg[1931];
        i_8_1259 <= in_reg[2187];
        i_8_1260 <= in_reg[140];
        i_8_1261 <= in_reg[396];
        i_8_1262 <= in_reg[652];
        i_8_1263 <= in_reg[908];
        i_8_1264 <= in_reg[1164];
        i_8_1265 <= in_reg[1420];
        i_8_1266 <= in_reg[1676];
        i_8_1267 <= in_reg[1932];
        i_8_1268 <= in_reg[2188];
        i_8_1269 <= in_reg[141];
        i_8_1270 <= in_reg[397];
        i_8_1271 <= in_reg[653];
        i_8_1272 <= in_reg[909];
        i_8_1273 <= in_reg[1165];
        i_8_1274 <= in_reg[1421];
        i_8_1275 <= in_reg[1677];
        i_8_1276 <= in_reg[1933];
        i_8_1277 <= in_reg[2189];
        i_8_1278 <= in_reg[142];
        i_8_1279 <= in_reg[398];
        i_8_1280 <= in_reg[654];
        i_8_1281 <= in_reg[910];
        i_8_1282 <= in_reg[1166];
        i_8_1283 <= in_reg[1422];
        i_8_1284 <= in_reg[1678];
        i_8_1285 <= in_reg[1934];
        i_8_1286 <= in_reg[2190];
        i_8_1287 <= in_reg[143];
        i_8_1288 <= in_reg[399];
        i_8_1289 <= in_reg[655];
        i_8_1290 <= in_reg[911];
        i_8_1291 <= in_reg[1167];
        i_8_1292 <= in_reg[1423];
        i_8_1293 <= in_reg[1679];
        i_8_1294 <= in_reg[1935];
        i_8_1295 <= in_reg[2191];
        i_8_1296 <= in_reg[144];
        i_8_1297 <= in_reg[400];
        i_8_1298 <= in_reg[656];
        i_8_1299 <= in_reg[912];
        i_8_1300 <= in_reg[1168];
        i_8_1301 <= in_reg[1424];
        i_8_1302 <= in_reg[1680];
        i_8_1303 <= in_reg[1936];
        i_8_1304 <= in_reg[2192];
        i_8_1305 <= in_reg[145];
        i_8_1306 <= in_reg[401];
        i_8_1307 <= in_reg[657];
        i_8_1308 <= in_reg[913];
        i_8_1309 <= in_reg[1169];
        i_8_1310 <= in_reg[1425];
        i_8_1311 <= in_reg[1681];
        i_8_1312 <= in_reg[1937];
        i_8_1313 <= in_reg[2193];
        i_8_1314 <= in_reg[146];
        i_8_1315 <= in_reg[402];
        i_8_1316 <= in_reg[658];
        i_8_1317 <= in_reg[914];
        i_8_1318 <= in_reg[1170];
        i_8_1319 <= in_reg[1426];
        i_8_1320 <= in_reg[1682];
        i_8_1321 <= in_reg[1938];
        i_8_1322 <= in_reg[2194];
        i_8_1323 <= in_reg[147];
        i_8_1324 <= in_reg[403];
        i_8_1325 <= in_reg[659];
        i_8_1326 <= in_reg[915];
        i_8_1327 <= in_reg[1171];
        i_8_1328 <= in_reg[1427];
        i_8_1329 <= in_reg[1683];
        i_8_1330 <= in_reg[1939];
        i_8_1331 <= in_reg[2195];
        i_8_1332 <= in_reg[148];
        i_8_1333 <= in_reg[404];
        i_8_1334 <= in_reg[660];
        i_8_1335 <= in_reg[916];
        i_8_1336 <= in_reg[1172];
        i_8_1337 <= in_reg[1428];
        i_8_1338 <= in_reg[1684];
        i_8_1339 <= in_reg[1940];
        i_8_1340 <= in_reg[2196];
        i_8_1341 <= in_reg[149];
        i_8_1342 <= in_reg[405];
        i_8_1343 <= in_reg[661];
        i_8_1344 <= in_reg[917];
        i_8_1345 <= in_reg[1173];
        i_8_1346 <= in_reg[1429];
        i_8_1347 <= in_reg[1685];
        i_8_1348 <= in_reg[1941];
        i_8_1349 <= in_reg[2197];
        i_8_1350 <= in_reg[150];
        i_8_1351 <= in_reg[406];
        i_8_1352 <= in_reg[662];
        i_8_1353 <= in_reg[918];
        i_8_1354 <= in_reg[1174];
        i_8_1355 <= in_reg[1430];
        i_8_1356 <= in_reg[1686];
        i_8_1357 <= in_reg[1942];
        i_8_1358 <= in_reg[2198];
        i_8_1359 <= in_reg[151];
        i_8_1360 <= in_reg[407];
        i_8_1361 <= in_reg[663];
        i_8_1362 <= in_reg[919];
        i_8_1363 <= in_reg[1175];
        i_8_1364 <= in_reg[1431];
        i_8_1365 <= in_reg[1687];
        i_8_1366 <= in_reg[1943];
        i_8_1367 <= in_reg[2199];
        i_8_1368 <= in_reg[152];
        i_8_1369 <= in_reg[408];
        i_8_1370 <= in_reg[664];
        i_8_1371 <= in_reg[920];
        i_8_1372 <= in_reg[1176];
        i_8_1373 <= in_reg[1432];
        i_8_1374 <= in_reg[1688];
        i_8_1375 <= in_reg[1944];
        i_8_1376 <= in_reg[2200];
        i_8_1377 <= in_reg[153];
        i_8_1378 <= in_reg[409];
        i_8_1379 <= in_reg[665];
        i_8_1380 <= in_reg[921];
        i_8_1381 <= in_reg[1177];
        i_8_1382 <= in_reg[1433];
        i_8_1383 <= in_reg[1689];
        i_8_1384 <= in_reg[1945];
        i_8_1385 <= in_reg[2201];
        i_8_1386 <= in_reg[154];
        i_8_1387 <= in_reg[410];
        i_8_1388 <= in_reg[666];
        i_8_1389 <= in_reg[922];
        i_8_1390 <= in_reg[1178];
        i_8_1391 <= in_reg[1434];
        i_8_1392 <= in_reg[1690];
        i_8_1393 <= in_reg[1946];
        i_8_1394 <= in_reg[2202];
        i_8_1395 <= in_reg[155];
        i_8_1396 <= in_reg[411];
        i_8_1397 <= in_reg[667];
        i_8_1398 <= in_reg[923];
        i_8_1399 <= in_reg[1179];
        i_8_1400 <= in_reg[1435];
        i_8_1401 <= in_reg[1691];
        i_8_1402 <= in_reg[1947];
        i_8_1403 <= in_reg[2203];
        i_8_1404 <= in_reg[156];
        i_8_1405 <= in_reg[412];
        i_8_1406 <= in_reg[668];
        i_8_1407 <= in_reg[924];
        i_8_1408 <= in_reg[1180];
        i_8_1409 <= in_reg[1436];
        i_8_1410 <= in_reg[1692];
        i_8_1411 <= in_reg[1948];
        i_8_1412 <= in_reg[2204];
        i_8_1413 <= in_reg[157];
        i_8_1414 <= in_reg[413];
        i_8_1415 <= in_reg[669];
        i_8_1416 <= in_reg[925];
        i_8_1417 <= in_reg[1181];
        i_8_1418 <= in_reg[1437];
        i_8_1419 <= in_reg[1693];
        i_8_1420 <= in_reg[1949];
        i_8_1421 <= in_reg[2205];
        i_8_1422 <= in_reg[158];
        i_8_1423 <= in_reg[414];
        i_8_1424 <= in_reg[670];
        i_8_1425 <= in_reg[926];
        i_8_1426 <= in_reg[1182];
        i_8_1427 <= in_reg[1438];
        i_8_1428 <= in_reg[1694];
        i_8_1429 <= in_reg[1950];
        i_8_1430 <= in_reg[2206];
        i_8_1431 <= in_reg[159];
        i_8_1432 <= in_reg[415];
        i_8_1433 <= in_reg[671];
        i_8_1434 <= in_reg[927];
        i_8_1435 <= in_reg[1183];
        i_8_1436 <= in_reg[1439];
        i_8_1437 <= in_reg[1695];
        i_8_1438 <= in_reg[1951];
        i_8_1439 <= in_reg[2207];
        i_8_1440 <= in_reg[160];
        i_8_1441 <= in_reg[416];
        i_8_1442 <= in_reg[672];
        i_8_1443 <= in_reg[928];
        i_8_1444 <= in_reg[1184];
        i_8_1445 <= in_reg[1440];
        i_8_1446 <= in_reg[1696];
        i_8_1447 <= in_reg[1952];
        i_8_1448 <= in_reg[2208];
        i_8_1449 <= in_reg[161];
        i_8_1450 <= in_reg[417];
        i_8_1451 <= in_reg[673];
        i_8_1452 <= in_reg[929];
        i_8_1453 <= in_reg[1185];
        i_8_1454 <= in_reg[1441];
        i_8_1455 <= in_reg[1697];
        i_8_1456 <= in_reg[1953];
        i_8_1457 <= in_reg[2209];
        i_8_1458 <= in_reg[162];
        i_8_1459 <= in_reg[418];
        i_8_1460 <= in_reg[674];
        i_8_1461 <= in_reg[930];
        i_8_1462 <= in_reg[1186];
        i_8_1463 <= in_reg[1442];
        i_8_1464 <= in_reg[1698];
        i_8_1465 <= in_reg[1954];
        i_8_1466 <= in_reg[2210];
        i_8_1467 <= in_reg[163];
        i_8_1468 <= in_reg[419];
        i_8_1469 <= in_reg[675];
        i_8_1470 <= in_reg[931];
        i_8_1471 <= in_reg[1187];
        i_8_1472 <= in_reg[1443];
        i_8_1473 <= in_reg[1699];
        i_8_1474 <= in_reg[1955];
        i_8_1475 <= in_reg[2211];
        i_8_1476 <= in_reg[164];
        i_8_1477 <= in_reg[420];
        i_8_1478 <= in_reg[676];
        i_8_1479 <= in_reg[932];
        i_8_1480 <= in_reg[1188];
        i_8_1481 <= in_reg[1444];
        i_8_1482 <= in_reg[1700];
        i_8_1483 <= in_reg[1956];
        i_8_1484 <= in_reg[2212];
        i_8_1485 <= in_reg[165];
        i_8_1486 <= in_reg[421];
        i_8_1487 <= in_reg[677];
        i_8_1488 <= in_reg[933];
        i_8_1489 <= in_reg[1189];
        i_8_1490 <= in_reg[1445];
        i_8_1491 <= in_reg[1701];
        i_8_1492 <= in_reg[1957];
        i_8_1493 <= in_reg[2213];
        i_8_1494 <= in_reg[166];
        i_8_1495 <= in_reg[422];
        i_8_1496 <= in_reg[678];
        i_8_1497 <= in_reg[934];
        i_8_1498 <= in_reg[1190];
        i_8_1499 <= in_reg[1446];
        i_8_1500 <= in_reg[1702];
        i_8_1501 <= in_reg[1958];
        i_8_1502 <= in_reg[2214];
        i_8_1503 <= in_reg[167];
        i_8_1504 <= in_reg[423];
        i_8_1505 <= in_reg[679];
        i_8_1506 <= in_reg[935];
        i_8_1507 <= in_reg[1191];
        i_8_1508 <= in_reg[1447];
        i_8_1509 <= in_reg[1703];
        i_8_1510 <= in_reg[1959];
        i_8_1511 <= in_reg[2215];
        i_8_1512 <= in_reg[168];
        i_8_1513 <= in_reg[424];
        i_8_1514 <= in_reg[680];
        i_8_1515 <= in_reg[936];
        i_8_1516 <= in_reg[1192];
        i_8_1517 <= in_reg[1448];
        i_8_1518 <= in_reg[1704];
        i_8_1519 <= in_reg[1960];
        i_8_1520 <= in_reg[2216];
        i_8_1521 <= in_reg[169];
        i_8_1522 <= in_reg[425];
        i_8_1523 <= in_reg[681];
        i_8_1524 <= in_reg[937];
        i_8_1525 <= in_reg[1193];
        i_8_1526 <= in_reg[1449];
        i_8_1527 <= in_reg[1705];
        i_8_1528 <= in_reg[1961];
        i_8_1529 <= in_reg[2217];
        i_8_1530 <= in_reg[170];
        i_8_1531 <= in_reg[426];
        i_8_1532 <= in_reg[682];
        i_8_1533 <= in_reg[938];
        i_8_1534 <= in_reg[1194];
        i_8_1535 <= in_reg[1450];
        i_8_1536 <= in_reg[1706];
        i_8_1537 <= in_reg[1962];
        i_8_1538 <= in_reg[2218];
        i_8_1539 <= in_reg[171];
        i_8_1540 <= in_reg[427];
        i_8_1541 <= in_reg[683];
        i_8_1542 <= in_reg[939];
        i_8_1543 <= in_reg[1195];
        i_8_1544 <= in_reg[1451];
        i_8_1545 <= in_reg[1707];
        i_8_1546 <= in_reg[1963];
        i_8_1547 <= in_reg[2219];
        i_8_1548 <= in_reg[172];
        i_8_1549 <= in_reg[428];
        i_8_1550 <= in_reg[684];
        i_8_1551 <= in_reg[940];
        i_8_1552 <= in_reg[1196];
        i_8_1553 <= in_reg[1452];
        i_8_1554 <= in_reg[1708];
        i_8_1555 <= in_reg[1964];
        i_8_1556 <= in_reg[2220];
        i_8_1557 <= in_reg[173];
        i_8_1558 <= in_reg[429];
        i_8_1559 <= in_reg[685];
        i_8_1560 <= in_reg[941];
        i_8_1561 <= in_reg[1197];
        i_8_1562 <= in_reg[1453];
        i_8_1563 <= in_reg[1709];
        i_8_1564 <= in_reg[1965];
        i_8_1565 <= in_reg[2221];
        i_8_1566 <= in_reg[174];
        i_8_1567 <= in_reg[430];
        i_8_1568 <= in_reg[686];
        i_8_1569 <= in_reg[942];
        i_8_1570 <= in_reg[1198];
        i_8_1571 <= in_reg[1454];
        i_8_1572 <= in_reg[1710];
        i_8_1573 <= in_reg[1966];
        i_8_1574 <= in_reg[2222];
        i_8_1575 <= in_reg[175];
        i_8_1576 <= in_reg[431];
        i_8_1577 <= in_reg[687];
        i_8_1578 <= in_reg[943];
        i_8_1579 <= in_reg[1199];
        i_8_1580 <= in_reg[1455];
        i_8_1581 <= in_reg[1711];
        i_8_1582 <= in_reg[1967];
        i_8_1583 <= in_reg[2223];
        i_8_1584 <= in_reg[176];
        i_8_1585 <= in_reg[432];
        i_8_1586 <= in_reg[688];
        i_8_1587 <= in_reg[944];
        i_8_1588 <= in_reg[1200];
        i_8_1589 <= in_reg[1456];
        i_8_1590 <= in_reg[1712];
        i_8_1591 <= in_reg[1968];
        i_8_1592 <= in_reg[2224];
        i_8_1593 <= in_reg[177];
        i_8_1594 <= in_reg[433];
        i_8_1595 <= in_reg[689];
        i_8_1596 <= in_reg[945];
        i_8_1597 <= in_reg[1201];
        i_8_1598 <= in_reg[1457];
        i_8_1599 <= in_reg[1713];
        i_8_1600 <= in_reg[1969];
        i_8_1601 <= in_reg[2225];
        i_8_1602 <= in_reg[178];
        i_8_1603 <= in_reg[434];
        i_8_1604 <= in_reg[690];
        i_8_1605 <= in_reg[946];
        i_8_1606 <= in_reg[1202];
        i_8_1607 <= in_reg[1458];
        i_8_1608 <= in_reg[1714];
        i_8_1609 <= in_reg[1970];
        i_8_1610 <= in_reg[2226];
        i_8_1611 <= in_reg[179];
        i_8_1612 <= in_reg[435];
        i_8_1613 <= in_reg[691];
        i_8_1614 <= in_reg[947];
        i_8_1615 <= in_reg[1203];
        i_8_1616 <= in_reg[1459];
        i_8_1617 <= in_reg[1715];
        i_8_1618 <= in_reg[1971];
        i_8_1619 <= in_reg[2227];
        i_8_1620 <= in_reg[180];
        i_8_1621 <= in_reg[436];
        i_8_1622 <= in_reg[692];
        i_8_1623 <= in_reg[948];
        i_8_1624 <= in_reg[1204];
        i_8_1625 <= in_reg[1460];
        i_8_1626 <= in_reg[1716];
        i_8_1627 <= in_reg[1972];
        i_8_1628 <= in_reg[2228];
        i_8_1629 <= in_reg[181];
        i_8_1630 <= in_reg[437];
        i_8_1631 <= in_reg[693];
        i_8_1632 <= in_reg[949];
        i_8_1633 <= in_reg[1205];
        i_8_1634 <= in_reg[1461];
        i_8_1635 <= in_reg[1717];
        i_8_1636 <= in_reg[1973];
        i_8_1637 <= in_reg[2229];
        i_8_1638 <= in_reg[182];
        i_8_1639 <= in_reg[438];
        i_8_1640 <= in_reg[694];
        i_8_1641 <= in_reg[950];
        i_8_1642 <= in_reg[1206];
        i_8_1643 <= in_reg[1462];
        i_8_1644 <= in_reg[1718];
        i_8_1645 <= in_reg[1974];
        i_8_1646 <= in_reg[2230];
        i_8_1647 <= in_reg[183];
        i_8_1648 <= in_reg[439];
        i_8_1649 <= in_reg[695];
        i_8_1650 <= in_reg[951];
        i_8_1651 <= in_reg[1207];
        i_8_1652 <= in_reg[1463];
        i_8_1653 <= in_reg[1719];
        i_8_1654 <= in_reg[1975];
        i_8_1655 <= in_reg[2231];
        i_8_1656 <= in_reg[184];
        i_8_1657 <= in_reg[440];
        i_8_1658 <= in_reg[696];
        i_8_1659 <= in_reg[952];
        i_8_1660 <= in_reg[1208];
        i_8_1661 <= in_reg[1464];
        i_8_1662 <= in_reg[1720];
        i_8_1663 <= in_reg[1976];
        i_8_1664 <= in_reg[2232];
        i_8_1665 <= in_reg[185];
        i_8_1666 <= in_reg[441];
        i_8_1667 <= in_reg[697];
        i_8_1668 <= in_reg[953];
        i_8_1669 <= in_reg[1209];
        i_8_1670 <= in_reg[1465];
        i_8_1671 <= in_reg[1721];
        i_8_1672 <= in_reg[1977];
        i_8_1673 <= in_reg[2233];
        i_8_1674 <= in_reg[186];
        i_8_1675 <= in_reg[442];
        i_8_1676 <= in_reg[698];
        i_8_1677 <= in_reg[954];
        i_8_1678 <= in_reg[1210];
        i_8_1679 <= in_reg[1466];
        i_8_1680 <= in_reg[1722];
        i_8_1681 <= in_reg[1978];
        i_8_1682 <= in_reg[2234];
        i_8_1683 <= in_reg[187];
        i_8_1684 <= in_reg[443];
        i_8_1685 <= in_reg[699];
        i_8_1686 <= in_reg[955];
        i_8_1687 <= in_reg[1211];
        i_8_1688 <= in_reg[1467];
        i_8_1689 <= in_reg[1723];
        i_8_1690 <= in_reg[1979];
        i_8_1691 <= in_reg[2235];
        i_8_1692 <= in_reg[188];
        i_8_1693 <= in_reg[444];
        i_8_1694 <= in_reg[700];
        i_8_1695 <= in_reg[956];
        i_8_1696 <= in_reg[1212];
        i_8_1697 <= in_reg[1468];
        i_8_1698 <= in_reg[1724];
        i_8_1699 <= in_reg[1980];
        i_8_1700 <= in_reg[2236];
        i_8_1701 <= in_reg[189];
        i_8_1702 <= in_reg[445];
        i_8_1703 <= in_reg[701];
        i_8_1704 <= in_reg[957];
        i_8_1705 <= in_reg[1213];
        i_8_1706 <= in_reg[1469];
        i_8_1707 <= in_reg[1725];
        i_8_1708 <= in_reg[1981];
        i_8_1709 <= in_reg[2237];
        i_8_1710 <= in_reg[190];
        i_8_1711 <= in_reg[446];
        i_8_1712 <= in_reg[702];
        i_8_1713 <= in_reg[958];
        i_8_1714 <= in_reg[1214];
        i_8_1715 <= in_reg[1470];
        i_8_1716 <= in_reg[1726];
        i_8_1717 <= in_reg[1982];
        i_8_1718 <= in_reg[2238];
        i_8_1719 <= in_reg[191];
        i_8_1720 <= in_reg[447];
        i_8_1721 <= in_reg[703];
        i_8_1722 <= in_reg[959];
        i_8_1723 <= in_reg[1215];
        i_8_1724 <= in_reg[1471];
        i_8_1725 <= in_reg[1727];
        i_8_1726 <= in_reg[1983];
        i_8_1727 <= in_reg[2239];
        i_8_1728 <= in_reg[192];
        i_8_1729 <= in_reg[448];
        i_8_1730 <= in_reg[704];
        i_8_1731 <= in_reg[960];
        i_8_1732 <= in_reg[1216];
        i_8_1733 <= in_reg[1472];
        i_8_1734 <= in_reg[1728];
        i_8_1735 <= in_reg[1984];
        i_8_1736 <= in_reg[2240];
        i_8_1737 <= in_reg[193];
        i_8_1738 <= in_reg[449];
        i_8_1739 <= in_reg[705];
        i_8_1740 <= in_reg[961];
        i_8_1741 <= in_reg[1217];
        i_8_1742 <= in_reg[1473];
        i_8_1743 <= in_reg[1729];
        i_8_1744 <= in_reg[1985];
        i_8_1745 <= in_reg[2241];
        i_8_1746 <= in_reg[194];
        i_8_1747 <= in_reg[450];
        i_8_1748 <= in_reg[706];
        i_8_1749 <= in_reg[962];
        i_8_1750 <= in_reg[1218];
        i_8_1751 <= in_reg[1474];
        i_8_1752 <= in_reg[1730];
        i_8_1753 <= in_reg[1986];
        i_8_1754 <= in_reg[2242];
        i_8_1755 <= in_reg[195];
        i_8_1756 <= in_reg[451];
        i_8_1757 <= in_reg[707];
        i_8_1758 <= in_reg[963];
        i_8_1759 <= in_reg[1219];
        i_8_1760 <= in_reg[1475];
        i_8_1761 <= in_reg[1731];
        i_8_1762 <= in_reg[1987];
        i_8_1763 <= in_reg[2243];
        i_8_1764 <= in_reg[196];
        i_8_1765 <= in_reg[452];
        i_8_1766 <= in_reg[708];
        i_8_1767 <= in_reg[964];
        i_8_1768 <= in_reg[1220];
        i_8_1769 <= in_reg[1476];
        i_8_1770 <= in_reg[1732];
        i_8_1771 <= in_reg[1988];
        i_8_1772 <= in_reg[2244];
        i_8_1773 <= in_reg[197];
        i_8_1774 <= in_reg[453];
        i_8_1775 <= in_reg[709];
        i_8_1776 <= in_reg[965];
        i_8_1777 <= in_reg[1221];
        i_8_1778 <= in_reg[1477];
        i_8_1779 <= in_reg[1733];
        i_8_1780 <= in_reg[1989];
        i_8_1781 <= in_reg[2245];
        i_8_1782 <= in_reg[198];
        i_8_1783 <= in_reg[454];
        i_8_1784 <= in_reg[710];
        i_8_1785 <= in_reg[966];
        i_8_1786 <= in_reg[1222];
        i_8_1787 <= in_reg[1478];
        i_8_1788 <= in_reg[1734];
        i_8_1789 <= in_reg[1990];
        i_8_1790 <= in_reg[2246];
        i_8_1791 <= in_reg[199];
        i_8_1792 <= in_reg[455];
        i_8_1793 <= in_reg[711];
        i_8_1794 <= in_reg[967];
        i_8_1795 <= in_reg[1223];
        i_8_1796 <= in_reg[1479];
        i_8_1797 <= in_reg[1735];
        i_8_1798 <= in_reg[1991];
        i_8_1799 <= in_reg[2247];
        i_8_1800 <= in_reg[200];
        i_8_1801 <= in_reg[456];
        i_8_1802 <= in_reg[712];
        i_8_1803 <= in_reg[968];
        i_8_1804 <= in_reg[1224];
        i_8_1805 <= in_reg[1480];
        i_8_1806 <= in_reg[1736];
        i_8_1807 <= in_reg[1992];
        i_8_1808 <= in_reg[2248];
        i_8_1809 <= in_reg[201];
        i_8_1810 <= in_reg[457];
        i_8_1811 <= in_reg[713];
        i_8_1812 <= in_reg[969];
        i_8_1813 <= in_reg[1225];
        i_8_1814 <= in_reg[1481];
        i_8_1815 <= in_reg[1737];
        i_8_1816 <= in_reg[1993];
        i_8_1817 <= in_reg[2249];
        i_8_1818 <= in_reg[202];
        i_8_1819 <= in_reg[458];
        i_8_1820 <= in_reg[714];
        i_8_1821 <= in_reg[970];
        i_8_1822 <= in_reg[1226];
        i_8_1823 <= in_reg[1482];
        i_8_1824 <= in_reg[1738];
        i_8_1825 <= in_reg[1994];
        i_8_1826 <= in_reg[2250];
        i_8_1827 <= in_reg[203];
        i_8_1828 <= in_reg[459];
        i_8_1829 <= in_reg[715];
        i_8_1830 <= in_reg[971];
        i_8_1831 <= in_reg[1227];
        i_8_1832 <= in_reg[1483];
        i_8_1833 <= in_reg[1739];
        i_8_1834 <= in_reg[1995];
        i_8_1835 <= in_reg[2251];
        i_8_1836 <= in_reg[204];
        i_8_1837 <= in_reg[460];
        i_8_1838 <= in_reg[716];
        i_8_1839 <= in_reg[972];
        i_8_1840 <= in_reg[1228];
        i_8_1841 <= in_reg[1484];
        i_8_1842 <= in_reg[1740];
        i_8_1843 <= in_reg[1996];
        i_8_1844 <= in_reg[2252];
        i_8_1845 <= in_reg[205];
        i_8_1846 <= in_reg[461];
        i_8_1847 <= in_reg[717];
        i_8_1848 <= in_reg[973];
        i_8_1849 <= in_reg[1229];
        i_8_1850 <= in_reg[1485];
        i_8_1851 <= in_reg[1741];
        i_8_1852 <= in_reg[1997];
        i_8_1853 <= in_reg[2253];
        i_8_1854 <= in_reg[206];
        i_8_1855 <= in_reg[462];
        i_8_1856 <= in_reg[718];
        i_8_1857 <= in_reg[974];
        i_8_1858 <= in_reg[1230];
        i_8_1859 <= in_reg[1486];
        i_8_1860 <= in_reg[1742];
        i_8_1861 <= in_reg[1998];
        i_8_1862 <= in_reg[2254];
        i_8_1863 <= in_reg[207];
        i_8_1864 <= in_reg[463];
        i_8_1865 <= in_reg[719];
        i_8_1866 <= in_reg[975];
        i_8_1867 <= in_reg[1231];
        i_8_1868 <= in_reg[1487];
        i_8_1869 <= in_reg[1743];
        i_8_1870 <= in_reg[1999];
        i_8_1871 <= in_reg[2255];
        i_8_1872 <= in_reg[208];
        i_8_1873 <= in_reg[464];
        i_8_1874 <= in_reg[720];
        i_8_1875 <= in_reg[976];
        i_8_1876 <= in_reg[1232];
        i_8_1877 <= in_reg[1488];
        i_8_1878 <= in_reg[1744];
        i_8_1879 <= in_reg[2000];
        i_8_1880 <= in_reg[2256];
        i_8_1881 <= in_reg[209];
        i_8_1882 <= in_reg[465];
        i_8_1883 <= in_reg[721];
        i_8_1884 <= in_reg[977];
        i_8_1885 <= in_reg[1233];
        i_8_1886 <= in_reg[1489];
        i_8_1887 <= in_reg[1745];
        i_8_1888 <= in_reg[2001];
        i_8_1889 <= in_reg[2257];
        i_8_1890 <= in_reg[210];
        i_8_1891 <= in_reg[466];
        i_8_1892 <= in_reg[722];
        i_8_1893 <= in_reg[978];
        i_8_1894 <= in_reg[1234];
        i_8_1895 <= in_reg[1490];
        i_8_1896 <= in_reg[1746];
        i_8_1897 <= in_reg[2002];
        i_8_1898 <= in_reg[2258];
        i_8_1899 <= in_reg[211];
        i_8_1900 <= in_reg[467];
        i_8_1901 <= in_reg[723];
        i_8_1902 <= in_reg[979];
        i_8_1903 <= in_reg[1235];
        i_8_1904 <= in_reg[1491];
        i_8_1905 <= in_reg[1747];
        i_8_1906 <= in_reg[2003];
        i_8_1907 <= in_reg[2259];
        i_8_1908 <= in_reg[212];
        i_8_1909 <= in_reg[468];
        i_8_1910 <= in_reg[724];
        i_8_1911 <= in_reg[980];
        i_8_1912 <= in_reg[1236];
        i_8_1913 <= in_reg[1492];
        i_8_1914 <= in_reg[1748];
        i_8_1915 <= in_reg[2004];
        i_8_1916 <= in_reg[2260];
        i_8_1917 <= in_reg[213];
        i_8_1918 <= in_reg[469];
        i_8_1919 <= in_reg[725];
        i_8_1920 <= in_reg[981];
        i_8_1921 <= in_reg[1237];
        i_8_1922 <= in_reg[1493];
        i_8_1923 <= in_reg[1749];
        i_8_1924 <= in_reg[2005];
        i_8_1925 <= in_reg[2261];
        i_8_1926 <= in_reg[214];
        i_8_1927 <= in_reg[470];
        i_8_1928 <= in_reg[726];
        i_8_1929 <= in_reg[982];
        i_8_1930 <= in_reg[1238];
        i_8_1931 <= in_reg[1494];
        i_8_1932 <= in_reg[1750];
        i_8_1933 <= in_reg[2006];
        i_8_1934 <= in_reg[2262];
        i_8_1935 <= in_reg[215];
        i_8_1936 <= in_reg[471];
        i_8_1937 <= in_reg[727];
        i_8_1938 <= in_reg[983];
        i_8_1939 <= in_reg[1239];
        i_8_1940 <= in_reg[1495];
        i_8_1941 <= in_reg[1751];
        i_8_1942 <= in_reg[2007];
        i_8_1943 <= in_reg[2263];
        i_8_1944 <= in_reg[216];
        i_8_1945 <= in_reg[472];
        i_8_1946 <= in_reg[728];
        i_8_1947 <= in_reg[984];
        i_8_1948 <= in_reg[1240];
        i_8_1949 <= in_reg[1496];
        i_8_1950 <= in_reg[1752];
        i_8_1951 <= in_reg[2008];
        i_8_1952 <= in_reg[2264];
        i_8_1953 <= in_reg[217];
        i_8_1954 <= in_reg[473];
        i_8_1955 <= in_reg[729];
        i_8_1956 <= in_reg[985];
        i_8_1957 <= in_reg[1241];
        i_8_1958 <= in_reg[1497];
        i_8_1959 <= in_reg[1753];
        i_8_1960 <= in_reg[2009];
        i_8_1961 <= in_reg[2265];
        i_8_1962 <= in_reg[218];
        i_8_1963 <= in_reg[474];
        i_8_1964 <= in_reg[730];
        i_8_1965 <= in_reg[986];
        i_8_1966 <= in_reg[1242];
        i_8_1967 <= in_reg[1498];
        i_8_1968 <= in_reg[1754];
        i_8_1969 <= in_reg[2010];
        i_8_1970 <= in_reg[2266];
        i_8_1971 <= in_reg[219];
        i_8_1972 <= in_reg[475];
        i_8_1973 <= in_reg[731];
        i_8_1974 <= in_reg[987];
        i_8_1975 <= in_reg[1243];
        i_8_1976 <= in_reg[1499];
        i_8_1977 <= in_reg[1755];
        i_8_1978 <= in_reg[2011];
        i_8_1979 <= in_reg[2267];
        i_8_1980 <= in_reg[220];
        i_8_1981 <= in_reg[476];
        i_8_1982 <= in_reg[732];
        i_8_1983 <= in_reg[988];
        i_8_1984 <= in_reg[1244];
        i_8_1985 <= in_reg[1500];
        i_8_1986 <= in_reg[1756];
        i_8_1987 <= in_reg[2012];
        i_8_1988 <= in_reg[2268];
        i_8_1989 <= in_reg[221];
        i_8_1990 <= in_reg[477];
        i_8_1991 <= in_reg[733];
        i_8_1992 <= in_reg[989];
        i_8_1993 <= in_reg[1245];
        i_8_1994 <= in_reg[1501];
        i_8_1995 <= in_reg[1757];
        i_8_1996 <= in_reg[2013];
        i_8_1997 <= in_reg[2269];
        i_8_1998 <= in_reg[222];
        i_8_1999 <= in_reg[478];
        i_8_2000 <= in_reg[734];
        i_8_2001 <= in_reg[990];
        i_8_2002 <= in_reg[1246];
        i_8_2003 <= in_reg[1502];
        i_8_2004 <= in_reg[1758];
        i_8_2005 <= in_reg[2014];
        i_8_2006 <= in_reg[2270];
        i_8_2007 <= in_reg[223];
        i_8_2008 <= in_reg[479];
        i_8_2009 <= in_reg[735];
        i_8_2010 <= in_reg[991];
        i_8_2011 <= in_reg[1247];
        i_8_2012 <= in_reg[1503];
        i_8_2013 <= in_reg[1759];
        i_8_2014 <= in_reg[2015];
        i_8_2015 <= in_reg[2271];
        i_8_2016 <= in_reg[224];
        i_8_2017 <= in_reg[480];
        i_8_2018 <= in_reg[736];
        i_8_2019 <= in_reg[992];
        i_8_2020 <= in_reg[1248];
        i_8_2021 <= in_reg[1504];
        i_8_2022 <= in_reg[1760];
        i_8_2023 <= in_reg[2016];
        i_8_2024 <= in_reg[2272];
        i_8_2025 <= in_reg[225];
        i_8_2026 <= in_reg[481];
        i_8_2027 <= in_reg[737];
        i_8_2028 <= in_reg[993];
        i_8_2029 <= in_reg[1249];
        i_8_2030 <= in_reg[1505];
        i_8_2031 <= in_reg[1761];
        i_8_2032 <= in_reg[2017];
        i_8_2033 <= in_reg[2273];
        i_8_2034 <= in_reg[226];
        i_8_2035 <= in_reg[482];
        i_8_2036 <= in_reg[738];
        i_8_2037 <= in_reg[994];
        i_8_2038 <= in_reg[1250];
        i_8_2039 <= in_reg[1506];
        i_8_2040 <= in_reg[1762];
        i_8_2041 <= in_reg[2018];
        i_8_2042 <= in_reg[2274];
        i_8_2043 <= in_reg[227];
        i_8_2044 <= in_reg[483];
        i_8_2045 <= in_reg[739];
        i_8_2046 <= in_reg[995];
        i_8_2047 <= in_reg[1251];
        i_8_2048 <= in_reg[1507];
        i_8_2049 <= in_reg[1763];
        i_8_2050 <= in_reg[2019];
        i_8_2051 <= in_reg[2275];
        i_8_2052 <= in_reg[228];
        i_8_2053 <= in_reg[484];
        i_8_2054 <= in_reg[740];
        i_8_2055 <= in_reg[996];
        i_8_2056 <= in_reg[1252];
        i_8_2057 <= in_reg[1508];
        i_8_2058 <= in_reg[1764];
        i_8_2059 <= in_reg[2020];
        i_8_2060 <= in_reg[2276];
        i_8_2061 <= in_reg[229];
        i_8_2062 <= in_reg[485];
        i_8_2063 <= in_reg[741];
        i_8_2064 <= in_reg[997];
        i_8_2065 <= in_reg[1253];
        i_8_2066 <= in_reg[1509];
        i_8_2067 <= in_reg[1765];
        i_8_2068 <= in_reg[2021];
        i_8_2069 <= in_reg[2277];
        i_8_2070 <= in_reg[230];
        i_8_2071 <= in_reg[486];
        i_8_2072 <= in_reg[742];
        i_8_2073 <= in_reg[998];
        i_8_2074 <= in_reg[1254];
        i_8_2075 <= in_reg[1510];
        i_8_2076 <= in_reg[1766];
        i_8_2077 <= in_reg[2022];
        i_8_2078 <= in_reg[2278];
        i_8_2079 <= in_reg[231];
        i_8_2080 <= in_reg[487];
        i_8_2081 <= in_reg[743];
        i_8_2082 <= in_reg[999];
        i_8_2083 <= in_reg[1255];
        i_8_2084 <= in_reg[1511];
        i_8_2085 <= in_reg[1767];
        i_8_2086 <= in_reg[2023];
        i_8_2087 <= in_reg[2279];
        i_8_2088 <= in_reg[232];
        i_8_2089 <= in_reg[488];
        i_8_2090 <= in_reg[744];
        i_8_2091 <= in_reg[1000];
        i_8_2092 <= in_reg[1256];
        i_8_2093 <= in_reg[1512];
        i_8_2094 <= in_reg[1768];
        i_8_2095 <= in_reg[2024];
        i_8_2096 <= in_reg[2280];
        i_8_2097 <= in_reg[233];
        i_8_2098 <= in_reg[489];
        i_8_2099 <= in_reg[745];
        i_8_2100 <= in_reg[1001];
        i_8_2101 <= in_reg[1257];
        i_8_2102 <= in_reg[1513];
        i_8_2103 <= in_reg[1769];
        i_8_2104 <= in_reg[2025];
        i_8_2105 <= in_reg[2281];
        i_8_2106 <= in_reg[234];
        i_8_2107 <= in_reg[490];
        i_8_2108 <= in_reg[746];
        i_8_2109 <= in_reg[1002];
        i_8_2110 <= in_reg[1258];
        i_8_2111 <= in_reg[1514];
        i_8_2112 <= in_reg[1770];
        i_8_2113 <= in_reg[2026];
        i_8_2114 <= in_reg[2282];
        i_8_2115 <= in_reg[235];
        i_8_2116 <= in_reg[491];
        i_8_2117 <= in_reg[747];
        i_8_2118 <= in_reg[1003];
        i_8_2119 <= in_reg[1259];
        i_8_2120 <= in_reg[1515];
        i_8_2121 <= in_reg[1771];
        i_8_2122 <= in_reg[2027];
        i_8_2123 <= in_reg[2283];
        i_8_2124 <= in_reg[236];
        i_8_2125 <= in_reg[492];
        i_8_2126 <= in_reg[748];
        i_8_2127 <= in_reg[1004];
        i_8_2128 <= in_reg[1260];
        i_8_2129 <= in_reg[1516];
        i_8_2130 <= in_reg[1772];
        i_8_2131 <= in_reg[2028];
        i_8_2132 <= in_reg[2284];
        i_8_2133 <= in_reg[237];
        i_8_2134 <= in_reg[493];
        i_8_2135 <= in_reg[749];
        i_8_2136 <= in_reg[1005];
        i_8_2137 <= in_reg[1261];
        i_8_2138 <= in_reg[1517];
        i_8_2139 <= in_reg[1773];
        i_8_2140 <= in_reg[2029];
        i_8_2141 <= in_reg[2285];
        i_8_2142 <= in_reg[238];
        i_8_2143 <= in_reg[494];
        i_8_2144 <= in_reg[750];
        i_8_2145 <= in_reg[1006];
        i_8_2146 <= in_reg[1262];
        i_8_2147 <= in_reg[1518];
        i_8_2148 <= in_reg[1774];
        i_8_2149 <= in_reg[2030];
        i_8_2150 <= in_reg[2286];
        i_8_2151 <= in_reg[239];
        i_8_2152 <= in_reg[495];
        i_8_2153 <= in_reg[751];
        i_8_2154 <= in_reg[1007];
        i_8_2155 <= in_reg[1263];
        i_8_2156 <= in_reg[1519];
        i_8_2157 <= in_reg[1775];
        i_8_2158 <= in_reg[2031];
        i_8_2159 <= in_reg[2287];
        i_8_2160 <= in_reg[240];
        i_8_2161 <= in_reg[496];
        i_8_2162 <= in_reg[752];
        i_8_2163 <= in_reg[1008];
        i_8_2164 <= in_reg[1264];
        i_8_2165 <= in_reg[1520];
        i_8_2166 <= in_reg[1776];
        i_8_2167 <= in_reg[2032];
        i_8_2168 <= in_reg[2288];
        i_8_2169 <= in_reg[241];
        i_8_2170 <= in_reg[497];
        i_8_2171 <= in_reg[753];
        i_8_2172 <= in_reg[1009];
        i_8_2173 <= in_reg[1265];
        i_8_2174 <= in_reg[1521];
        i_8_2175 <= in_reg[1777];
        i_8_2176 <= in_reg[2033];
        i_8_2177 <= in_reg[2289];
        i_8_2178 <= in_reg[242];
        i_8_2179 <= in_reg[498];
        i_8_2180 <= in_reg[754];
        i_8_2181 <= in_reg[1010];
        i_8_2182 <= in_reg[1266];
        i_8_2183 <= in_reg[1522];
        i_8_2184 <= in_reg[1778];
        i_8_2185 <= in_reg[2034];
        i_8_2186 <= in_reg[2290];
        i_8_2187 <= in_reg[243];
        i_8_2188 <= in_reg[499];
        i_8_2189 <= in_reg[755];
        i_8_2190 <= in_reg[1011];
        i_8_2191 <= in_reg[1267];
        i_8_2192 <= in_reg[1523];
        i_8_2193 <= in_reg[1779];
        i_8_2194 <= in_reg[2035];
        i_8_2195 <= in_reg[2291];
        i_8_2196 <= in_reg[244];
        i_8_2197 <= in_reg[500];
        i_8_2198 <= in_reg[756];
        i_8_2199 <= in_reg[1012];
        i_8_2200 <= in_reg[1268];
        i_8_2201 <= in_reg[1524];
        i_8_2202 <= in_reg[1780];
        i_8_2203 <= in_reg[2036];
        i_8_2204 <= in_reg[2292];
        i_8_2205 <= in_reg[245];
        i_8_2206 <= in_reg[501];
        i_8_2207 <= in_reg[757];
        i_8_2208 <= in_reg[1013];
        i_8_2209 <= in_reg[1269];
        i_8_2210 <= in_reg[1525];
        i_8_2211 <= in_reg[1781];
        i_8_2212 <= in_reg[2037];
        i_8_2213 <= in_reg[2293];
        i_8_2214 <= in_reg[246];
        i_8_2215 <= in_reg[502];
        i_8_2216 <= in_reg[758];
        i_8_2217 <= in_reg[1014];
        i_8_2218 <= in_reg[1270];
        i_8_2219 <= in_reg[1526];
        i_8_2220 <= in_reg[1782];
        i_8_2221 <= in_reg[2038];
        i_8_2222 <= in_reg[2294];
        i_8_2223 <= in_reg[247];
        i_8_2224 <= in_reg[503];
        i_8_2225 <= in_reg[759];
        i_8_2226 <= in_reg[1015];
        i_8_2227 <= in_reg[1271];
        i_8_2228 <= in_reg[1527];
        i_8_2229 <= in_reg[1783];
        i_8_2230 <= in_reg[2039];
        i_8_2231 <= in_reg[2295];
        i_8_2232 <= in_reg[248];
        i_8_2233 <= in_reg[504];
        i_8_2234 <= in_reg[760];
        i_8_2235 <= in_reg[1016];
        i_8_2236 <= in_reg[1272];
        i_8_2237 <= in_reg[1528];
        i_8_2238 <= in_reg[1784];
        i_8_2239 <= in_reg[2040];
        i_8_2240 <= in_reg[2296];
        i_8_2241 <= in_reg[249];
        i_8_2242 <= in_reg[505];
        i_8_2243 <= in_reg[761];
        i_8_2244 <= in_reg[1017];
        i_8_2245 <= in_reg[1273];
        i_8_2246 <= in_reg[1529];
        i_8_2247 <= in_reg[1785];
        i_8_2248 <= in_reg[2041];
        i_8_2249 <= in_reg[2297];
        i_8_2250 <= in_reg[250];
        i_8_2251 <= in_reg[506];
        i_8_2252 <= in_reg[762];
        i_8_2253 <= in_reg[1018];
        i_8_2254 <= in_reg[1274];
        i_8_2255 <= in_reg[1530];
        i_8_2256 <= in_reg[1786];
        i_8_2257 <= in_reg[2042];
        i_8_2258 <= in_reg[2298];
        i_8_2259 <= in_reg[251];
        i_8_2260 <= in_reg[507];
        i_8_2261 <= in_reg[763];
        i_8_2262 <= in_reg[1019];
        i_8_2263 <= in_reg[1275];
        i_8_2264 <= in_reg[1531];
        i_8_2265 <= in_reg[1787];
        i_8_2266 <= in_reg[2043];
        i_8_2267 <= in_reg[2299];
        i_8_2268 <= in_reg[252];
        i_8_2269 <= in_reg[508];
        i_8_2270 <= in_reg[764];
        i_8_2271 <= in_reg[1020];
        i_8_2272 <= in_reg[1276];
        i_8_2273 <= in_reg[1532];
        i_8_2274 <= in_reg[1788];
        i_8_2275 <= in_reg[2044];
        i_8_2276 <= in_reg[2300];
        i_8_2277 <= in_reg[253];
        i_8_2278 <= in_reg[509];
        i_8_2279 <= in_reg[765];
        i_8_2280 <= in_reg[1021];
        i_8_2281 <= in_reg[1277];
        i_8_2282 <= in_reg[1533];
        i_8_2283 <= in_reg[1789];
        i_8_2284 <= in_reg[2045];
        i_8_2285 <= in_reg[2301];
        i_8_2286 <= in_reg[254];
        i_8_2287 <= in_reg[510];
        i_8_2288 <= in_reg[766];
        i_8_2289 <= in_reg[1022];
        i_8_2290 <= in_reg[1278];
        i_8_2291 <= in_reg[1534];
        i_8_2292 <= in_reg[1790];
        i_8_2293 <= in_reg[2046];
        i_8_2294 <= in_reg[2302];
        i_8_2295 <= in_reg[255];
        i_8_2296 <= in_reg[511];
        i_8_2297 <= in_reg[767];
        i_8_2298 <= in_reg[1023];
        i_8_2299 <= in_reg[1279];
        i_8_2300 <= in_reg[1535];
        i_8_2301 <= in_reg[1791];
        i_8_2302 <= in_reg[2047];
        i_8_2303 <= in_reg[2303];
        dly1 <= ap_start;
        dly2 <= dly1;
      end

  assign out_reg_ap_vld = dly2;
  assign ap_ready = dly2;
  assign ap_done = dly2;
  assign ap_idle = ~ap_start;

endmodule
